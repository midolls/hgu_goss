magic
tech sky130A
magscale 1 2
timestamp 1699539897
<< nwell >>
rect -270 -1139 1830 -767
rect -166 -2078 1830 -1757
rect -178 -2419 1830 -2078
rect -178 -2420 1795 -2419
<< pwell >>
rect -159 -1379 1791 -1197
rect 1728 -1417 1762 -1379
rect -97 -1517 -63 -1479
rect 636 -1517 670 -1479
rect 1176 -1517 1210 -1479
rect 1728 -1517 1762 -1479
rect -127 -1673 147 -1517
rect 177 -1699 699 -1517
rect 717 -1699 1239 -1517
rect 1269 -1699 1791 -1517
rect -139 -2659 135 -2503
rect 137 -2659 411 -2503
rect 413 -2659 687 -2503
rect 689 -2659 963 -2503
rect 965 -2659 1239 -2503
rect 1241 -2659 1515 -2503
rect 1517 -2659 1791 -2503
rect -109 -2697 -75 -2659
rect 167 -2697 201 -2659
rect 443 -2697 477 -2659
rect 899 -2697 933 -2659
rect 995 -2697 1029 -2659
rect 1451 -2697 1485 -2659
rect 1547 -2697 1581 -2659
<< scnmos >>
rect -81 -1353 -51 -1223
rect 3 -1353 33 -1223
rect 87 -1353 117 -1223
rect 171 -1353 201 -1223
rect 255 -1353 285 -1223
rect 339 -1353 369 -1223
rect 423 -1353 453 -1223
rect 507 -1353 537 -1223
rect 591 -1353 621 -1223
rect 675 -1353 705 -1223
rect 759 -1353 789 -1223
rect 843 -1353 873 -1223
rect 927 -1353 957 -1223
rect 1011 -1353 1041 -1223
rect 1095 -1353 1125 -1223
rect 1179 -1353 1209 -1223
rect 1263 -1353 1293 -1223
rect 1347 -1353 1377 -1223
rect 1431 -1353 1461 -1223
rect 1515 -1353 1545 -1223
rect 1599 -1353 1629 -1223
rect 1683 -1353 1713 -1223
rect -49 -1647 -19 -1543
rect 39 -1647 69 -1543
rect 255 -1673 285 -1543
rect 339 -1673 369 -1543
rect 423 -1673 453 -1543
rect 507 -1673 537 -1543
rect 591 -1673 621 -1543
rect 795 -1673 825 -1543
rect 879 -1673 909 -1543
rect 963 -1673 993 -1543
rect 1047 -1673 1077 -1543
rect 1131 -1673 1161 -1543
rect 1347 -1673 1377 -1543
rect 1431 -1673 1461 -1543
rect 1515 -1673 1545 -1543
rect 1599 -1673 1629 -1543
rect 1683 -1673 1713 -1543
rect -61 -2633 -31 -2529
rect 27 -2633 57 -2529
rect 215 -2633 245 -2529
rect 303 -2633 333 -2529
rect 491 -2633 521 -2529
rect 579 -2633 609 -2529
rect 767 -2633 797 -2529
rect 855 -2633 885 -2529
rect 1043 -2633 1073 -2529
rect 1131 -2633 1161 -2529
rect 1319 -2633 1349 -2529
rect 1407 -2633 1437 -2529
rect 1595 -2633 1625 -2529
rect 1683 -2633 1713 -2529
<< scpmoshvt >>
rect -81 -1103 -51 -903
rect 3 -1103 33 -903
rect 87 -1103 117 -903
rect 171 -1103 201 -903
rect 255 -1103 285 -903
rect 339 -1103 369 -903
rect 423 -1103 453 -903
rect 507 -1103 537 -903
rect 591 -1103 621 -903
rect 675 -1103 705 -903
rect 759 -1103 789 -903
rect 843 -1103 873 -903
rect 927 -1103 957 -903
rect 1011 -1103 1041 -903
rect 1095 -1103 1125 -903
rect 1179 -1103 1209 -903
rect 1263 -1103 1293 -903
rect 1347 -1103 1377 -903
rect 1431 -1103 1461 -903
rect 1515 -1103 1545 -903
rect 1599 -1103 1629 -903
rect 1683 -1103 1713 -903
rect -49 -1993 -19 -1835
rect 39 -1993 69 -1835
rect 255 -1993 285 -1793
rect 339 -1993 369 -1793
rect 423 -1993 453 -1793
rect 507 -1993 537 -1793
rect 591 -1993 621 -1793
rect 795 -1993 825 -1793
rect 879 -1993 909 -1793
rect 963 -1993 993 -1793
rect 1047 -1993 1077 -1793
rect 1131 -1993 1161 -1793
rect 1347 -1993 1377 -1793
rect 1431 -1993 1461 -1793
rect 1515 -1993 1545 -1793
rect 1599 -1993 1629 -1793
rect 1683 -1993 1713 -1793
rect -61 -2341 -31 -2183
rect 27 -2341 57 -2183
rect 215 -2341 245 -2183
rect 303 -2341 333 -2183
rect 491 -2341 521 -2183
rect 579 -2341 609 -2183
rect 767 -2341 797 -2183
rect 855 -2341 885 -2183
rect 1043 -2341 1073 -2183
rect 1131 -2341 1161 -2183
rect 1319 -2341 1349 -2183
rect 1407 -2341 1437 -2183
rect 1595 -2341 1625 -2183
rect 1683 -2341 1713 -2183
<< ndiff >>
rect -133 -1303 -81 -1223
rect -133 -1337 -125 -1303
rect -91 -1337 -81 -1303
rect -133 -1353 -81 -1337
rect -51 -1235 3 -1223
rect -51 -1269 -41 -1235
rect -7 -1269 3 -1235
rect -51 -1303 3 -1269
rect -51 -1337 -41 -1303
rect -7 -1337 3 -1303
rect -51 -1353 3 -1337
rect 33 -1303 87 -1223
rect 33 -1337 43 -1303
rect 77 -1337 87 -1303
rect 33 -1353 87 -1337
rect 117 -1235 171 -1223
rect 117 -1269 127 -1235
rect 161 -1269 171 -1235
rect 117 -1303 171 -1269
rect 117 -1337 127 -1303
rect 161 -1337 171 -1303
rect 117 -1353 171 -1337
rect 201 -1303 255 -1223
rect 201 -1337 211 -1303
rect 245 -1337 255 -1303
rect 201 -1353 255 -1337
rect 285 -1235 339 -1223
rect 285 -1269 295 -1235
rect 329 -1269 339 -1235
rect 285 -1303 339 -1269
rect 285 -1337 295 -1303
rect 329 -1337 339 -1303
rect 285 -1353 339 -1337
rect 369 -1303 423 -1223
rect 369 -1337 379 -1303
rect 413 -1337 423 -1303
rect 369 -1353 423 -1337
rect 453 -1235 507 -1223
rect 453 -1269 463 -1235
rect 497 -1269 507 -1235
rect 453 -1303 507 -1269
rect 453 -1337 463 -1303
rect 497 -1337 507 -1303
rect 453 -1353 507 -1337
rect 537 -1303 591 -1223
rect 537 -1337 547 -1303
rect 581 -1337 591 -1303
rect 537 -1353 591 -1337
rect 621 -1235 675 -1223
rect 621 -1269 631 -1235
rect 665 -1269 675 -1235
rect 621 -1303 675 -1269
rect 621 -1337 631 -1303
rect 665 -1337 675 -1303
rect 621 -1353 675 -1337
rect 705 -1303 759 -1223
rect 705 -1337 715 -1303
rect 749 -1337 759 -1303
rect 705 -1353 759 -1337
rect 789 -1235 843 -1223
rect 789 -1269 799 -1235
rect 833 -1269 843 -1235
rect 789 -1303 843 -1269
rect 789 -1337 799 -1303
rect 833 -1337 843 -1303
rect 789 -1353 843 -1337
rect 873 -1303 927 -1223
rect 873 -1337 883 -1303
rect 917 -1337 927 -1303
rect 873 -1353 927 -1337
rect 957 -1235 1011 -1223
rect 957 -1269 967 -1235
rect 1001 -1269 1011 -1235
rect 957 -1303 1011 -1269
rect 957 -1337 967 -1303
rect 1001 -1337 1011 -1303
rect 957 -1353 1011 -1337
rect 1041 -1303 1095 -1223
rect 1041 -1337 1051 -1303
rect 1085 -1337 1095 -1303
rect 1041 -1353 1095 -1337
rect 1125 -1235 1179 -1223
rect 1125 -1269 1135 -1235
rect 1169 -1269 1179 -1235
rect 1125 -1303 1179 -1269
rect 1125 -1337 1135 -1303
rect 1169 -1337 1179 -1303
rect 1125 -1353 1179 -1337
rect 1209 -1303 1263 -1223
rect 1209 -1337 1219 -1303
rect 1253 -1337 1263 -1303
rect 1209 -1353 1263 -1337
rect 1293 -1235 1347 -1223
rect 1293 -1269 1303 -1235
rect 1337 -1269 1347 -1235
rect 1293 -1303 1347 -1269
rect 1293 -1337 1303 -1303
rect 1337 -1337 1347 -1303
rect 1293 -1353 1347 -1337
rect 1377 -1303 1431 -1223
rect 1377 -1337 1387 -1303
rect 1421 -1337 1431 -1303
rect 1377 -1353 1431 -1337
rect 1461 -1235 1515 -1223
rect 1461 -1269 1471 -1235
rect 1505 -1269 1515 -1235
rect 1461 -1303 1515 -1269
rect 1461 -1337 1471 -1303
rect 1505 -1337 1515 -1303
rect 1461 -1353 1515 -1337
rect 1545 -1303 1599 -1223
rect 1545 -1337 1555 -1303
rect 1589 -1337 1599 -1303
rect 1545 -1353 1599 -1337
rect 1629 -1235 1683 -1223
rect 1629 -1269 1639 -1235
rect 1673 -1269 1683 -1235
rect 1629 -1303 1683 -1269
rect 1629 -1337 1639 -1303
rect 1673 -1337 1683 -1303
rect 1629 -1353 1683 -1337
rect 1713 -1235 1765 -1223
rect 1713 -1269 1723 -1235
rect 1757 -1269 1765 -1235
rect 1713 -1303 1765 -1269
rect 1713 -1337 1723 -1303
rect 1757 -1337 1765 -1303
rect 1713 -1353 1765 -1337
rect -101 -1568 -49 -1543
rect -101 -1602 -93 -1568
rect -59 -1602 -49 -1568
rect -101 -1647 -49 -1602
rect -19 -1555 39 -1543
rect -19 -1589 -7 -1555
rect 27 -1589 39 -1555
rect -19 -1647 39 -1589
rect 69 -1585 121 -1543
rect 69 -1619 79 -1585
rect 113 -1619 121 -1585
rect 69 -1647 121 -1619
rect 203 -1555 255 -1543
rect 203 -1589 211 -1555
rect 245 -1589 255 -1555
rect 203 -1623 255 -1589
rect 203 -1657 211 -1623
rect 245 -1657 255 -1623
rect 203 -1673 255 -1657
rect 285 -1591 339 -1543
rect 285 -1625 295 -1591
rect 329 -1625 339 -1591
rect 285 -1673 339 -1625
rect 369 -1559 423 -1543
rect 369 -1593 379 -1559
rect 413 -1593 423 -1559
rect 369 -1673 423 -1593
rect 453 -1591 507 -1543
rect 453 -1625 463 -1591
rect 497 -1625 507 -1591
rect 453 -1673 507 -1625
rect 537 -1559 591 -1543
rect 537 -1593 547 -1559
rect 581 -1593 591 -1559
rect 537 -1673 591 -1593
rect 621 -1591 673 -1543
rect 621 -1625 631 -1591
rect 665 -1625 673 -1591
rect 621 -1673 673 -1625
rect 743 -1555 795 -1543
rect 743 -1589 751 -1555
rect 785 -1589 795 -1555
rect 743 -1623 795 -1589
rect 743 -1657 751 -1623
rect 785 -1657 795 -1623
rect 743 -1673 795 -1657
rect 825 -1591 879 -1543
rect 825 -1625 835 -1591
rect 869 -1625 879 -1591
rect 825 -1673 879 -1625
rect 909 -1559 963 -1543
rect 909 -1593 919 -1559
rect 953 -1593 963 -1559
rect 909 -1673 963 -1593
rect 993 -1591 1047 -1543
rect 993 -1625 1003 -1591
rect 1037 -1625 1047 -1591
rect 993 -1673 1047 -1625
rect 1077 -1559 1131 -1543
rect 1077 -1593 1087 -1559
rect 1121 -1593 1131 -1559
rect 1077 -1673 1131 -1593
rect 1161 -1591 1213 -1543
rect 1161 -1625 1171 -1591
rect 1205 -1625 1213 -1591
rect 1161 -1673 1213 -1625
rect 1295 -1555 1347 -1543
rect 1295 -1589 1303 -1555
rect 1337 -1589 1347 -1555
rect 1295 -1623 1347 -1589
rect 1295 -1657 1303 -1623
rect 1337 -1657 1347 -1623
rect 1295 -1673 1347 -1657
rect 1377 -1591 1431 -1543
rect 1377 -1625 1387 -1591
rect 1421 -1625 1431 -1591
rect 1377 -1673 1431 -1625
rect 1461 -1559 1515 -1543
rect 1461 -1593 1471 -1559
rect 1505 -1593 1515 -1559
rect 1461 -1673 1515 -1593
rect 1545 -1591 1599 -1543
rect 1545 -1625 1555 -1591
rect 1589 -1625 1599 -1591
rect 1545 -1673 1599 -1625
rect 1629 -1559 1683 -1543
rect 1629 -1593 1639 -1559
rect 1673 -1593 1683 -1559
rect 1629 -1673 1683 -1593
rect 1713 -1591 1765 -1543
rect 1713 -1625 1723 -1591
rect 1757 -1625 1765 -1591
rect 1713 -1673 1765 -1625
rect -113 -2574 -61 -2529
rect -113 -2608 -105 -2574
rect -71 -2608 -61 -2574
rect -113 -2633 -61 -2608
rect -31 -2587 27 -2529
rect -31 -2621 -19 -2587
rect 15 -2621 27 -2587
rect -31 -2633 27 -2621
rect 57 -2557 109 -2529
rect 57 -2591 67 -2557
rect 101 -2591 109 -2557
rect 57 -2633 109 -2591
rect 163 -2574 215 -2529
rect 163 -2608 171 -2574
rect 205 -2608 215 -2574
rect 163 -2633 215 -2608
rect 245 -2587 303 -2529
rect 245 -2621 257 -2587
rect 291 -2621 303 -2587
rect 245 -2633 303 -2621
rect 333 -2557 385 -2529
rect 333 -2591 343 -2557
rect 377 -2591 385 -2557
rect 333 -2633 385 -2591
rect 439 -2574 491 -2529
rect 439 -2608 447 -2574
rect 481 -2608 491 -2574
rect 439 -2633 491 -2608
rect 521 -2587 579 -2529
rect 521 -2621 533 -2587
rect 567 -2621 579 -2587
rect 521 -2633 579 -2621
rect 609 -2557 661 -2529
rect 609 -2591 619 -2557
rect 653 -2591 661 -2557
rect 609 -2633 661 -2591
rect 715 -2557 767 -2529
rect 715 -2591 723 -2557
rect 757 -2591 767 -2557
rect 715 -2633 767 -2591
rect 797 -2587 855 -2529
rect 797 -2621 809 -2587
rect 843 -2621 855 -2587
rect 797 -2633 855 -2621
rect 885 -2574 937 -2529
rect 885 -2608 895 -2574
rect 929 -2608 937 -2574
rect 885 -2633 937 -2608
rect 991 -2574 1043 -2529
rect 991 -2608 999 -2574
rect 1033 -2608 1043 -2574
rect 991 -2633 1043 -2608
rect 1073 -2587 1131 -2529
rect 1073 -2621 1085 -2587
rect 1119 -2621 1131 -2587
rect 1073 -2633 1131 -2621
rect 1161 -2557 1213 -2529
rect 1161 -2591 1171 -2557
rect 1205 -2591 1213 -2557
rect 1161 -2633 1213 -2591
rect 1267 -2557 1319 -2529
rect 1267 -2591 1275 -2557
rect 1309 -2591 1319 -2557
rect 1267 -2633 1319 -2591
rect 1349 -2587 1407 -2529
rect 1349 -2621 1361 -2587
rect 1395 -2621 1407 -2587
rect 1349 -2633 1407 -2621
rect 1437 -2574 1489 -2529
rect 1437 -2608 1447 -2574
rect 1481 -2608 1489 -2574
rect 1437 -2633 1489 -2608
rect 1543 -2574 1595 -2529
rect 1543 -2608 1551 -2574
rect 1585 -2608 1595 -2574
rect 1543 -2633 1595 -2608
rect 1625 -2587 1683 -2529
rect 1625 -2621 1637 -2587
rect 1671 -2621 1683 -2587
rect 1625 -2633 1683 -2621
rect 1713 -2557 1765 -2529
rect 1713 -2591 1723 -2557
rect 1757 -2591 1765 -2557
rect 1713 -2633 1765 -2591
<< pdiff >>
rect -133 -915 -81 -903
rect -133 -949 -125 -915
rect -91 -949 -81 -915
rect -133 -983 -81 -949
rect -133 -1017 -125 -983
rect -91 -1017 -81 -983
rect -133 -1103 -81 -1017
rect -51 -921 3 -903
rect -51 -955 -41 -921
rect -7 -955 3 -921
rect -51 -989 3 -955
rect -51 -1023 -41 -989
rect -7 -1023 3 -989
rect -51 -1057 3 -1023
rect -51 -1091 -41 -1057
rect -7 -1091 3 -1057
rect -51 -1103 3 -1091
rect 33 -915 87 -903
rect 33 -949 43 -915
rect 77 -949 87 -915
rect 33 -983 87 -949
rect 33 -1017 43 -983
rect 77 -1017 87 -983
rect 33 -1103 87 -1017
rect 117 -921 171 -903
rect 117 -955 127 -921
rect 161 -955 171 -921
rect 117 -989 171 -955
rect 117 -1023 127 -989
rect 161 -1023 171 -989
rect 117 -1057 171 -1023
rect 117 -1091 127 -1057
rect 161 -1091 171 -1057
rect 117 -1103 171 -1091
rect 201 -915 255 -903
rect 201 -949 211 -915
rect 245 -949 255 -915
rect 201 -983 255 -949
rect 201 -1017 211 -983
rect 245 -1017 255 -983
rect 201 -1103 255 -1017
rect 285 -921 339 -903
rect 285 -955 295 -921
rect 329 -955 339 -921
rect 285 -989 339 -955
rect 285 -1023 295 -989
rect 329 -1023 339 -989
rect 285 -1057 339 -1023
rect 285 -1091 295 -1057
rect 329 -1091 339 -1057
rect 285 -1103 339 -1091
rect 369 -915 423 -903
rect 369 -949 379 -915
rect 413 -949 423 -915
rect 369 -983 423 -949
rect 369 -1017 379 -983
rect 413 -1017 423 -983
rect 369 -1103 423 -1017
rect 453 -921 507 -903
rect 453 -955 463 -921
rect 497 -955 507 -921
rect 453 -989 507 -955
rect 453 -1023 463 -989
rect 497 -1023 507 -989
rect 453 -1057 507 -1023
rect 453 -1091 463 -1057
rect 497 -1091 507 -1057
rect 453 -1103 507 -1091
rect 537 -915 591 -903
rect 537 -949 547 -915
rect 581 -949 591 -915
rect 537 -983 591 -949
rect 537 -1017 547 -983
rect 581 -1017 591 -983
rect 537 -1103 591 -1017
rect 621 -921 675 -903
rect 621 -955 631 -921
rect 665 -955 675 -921
rect 621 -989 675 -955
rect 621 -1023 631 -989
rect 665 -1023 675 -989
rect 621 -1057 675 -1023
rect 621 -1091 631 -1057
rect 665 -1091 675 -1057
rect 621 -1103 675 -1091
rect 705 -915 759 -903
rect 705 -949 715 -915
rect 749 -949 759 -915
rect 705 -983 759 -949
rect 705 -1017 715 -983
rect 749 -1017 759 -983
rect 705 -1103 759 -1017
rect 789 -921 843 -903
rect 789 -955 799 -921
rect 833 -955 843 -921
rect 789 -989 843 -955
rect 789 -1023 799 -989
rect 833 -1023 843 -989
rect 789 -1057 843 -1023
rect 789 -1091 799 -1057
rect 833 -1091 843 -1057
rect 789 -1103 843 -1091
rect 873 -915 927 -903
rect 873 -949 883 -915
rect 917 -949 927 -915
rect 873 -983 927 -949
rect 873 -1017 883 -983
rect 917 -1017 927 -983
rect 873 -1103 927 -1017
rect 957 -921 1011 -903
rect 957 -955 967 -921
rect 1001 -955 1011 -921
rect 957 -989 1011 -955
rect 957 -1023 967 -989
rect 1001 -1023 1011 -989
rect 957 -1057 1011 -1023
rect 957 -1091 967 -1057
rect 1001 -1091 1011 -1057
rect 957 -1103 1011 -1091
rect 1041 -915 1095 -903
rect 1041 -949 1051 -915
rect 1085 -949 1095 -915
rect 1041 -983 1095 -949
rect 1041 -1017 1051 -983
rect 1085 -1017 1095 -983
rect 1041 -1103 1095 -1017
rect 1125 -921 1179 -903
rect 1125 -955 1135 -921
rect 1169 -955 1179 -921
rect 1125 -989 1179 -955
rect 1125 -1023 1135 -989
rect 1169 -1023 1179 -989
rect 1125 -1057 1179 -1023
rect 1125 -1091 1135 -1057
rect 1169 -1091 1179 -1057
rect 1125 -1103 1179 -1091
rect 1209 -915 1263 -903
rect 1209 -949 1219 -915
rect 1253 -949 1263 -915
rect 1209 -983 1263 -949
rect 1209 -1017 1219 -983
rect 1253 -1017 1263 -983
rect 1209 -1103 1263 -1017
rect 1293 -921 1347 -903
rect 1293 -955 1303 -921
rect 1337 -955 1347 -921
rect 1293 -989 1347 -955
rect 1293 -1023 1303 -989
rect 1337 -1023 1347 -989
rect 1293 -1057 1347 -1023
rect 1293 -1091 1303 -1057
rect 1337 -1091 1347 -1057
rect 1293 -1103 1347 -1091
rect 1377 -915 1431 -903
rect 1377 -949 1387 -915
rect 1421 -949 1431 -915
rect 1377 -983 1431 -949
rect 1377 -1017 1387 -983
rect 1421 -1017 1431 -983
rect 1377 -1103 1431 -1017
rect 1461 -921 1515 -903
rect 1461 -955 1471 -921
rect 1505 -955 1515 -921
rect 1461 -989 1515 -955
rect 1461 -1023 1471 -989
rect 1505 -1023 1515 -989
rect 1461 -1057 1515 -1023
rect 1461 -1091 1471 -1057
rect 1505 -1091 1515 -1057
rect 1461 -1103 1515 -1091
rect 1545 -915 1599 -903
rect 1545 -949 1555 -915
rect 1589 -949 1599 -915
rect 1545 -983 1599 -949
rect 1545 -1017 1555 -983
rect 1589 -1017 1599 -983
rect 1545 -1103 1599 -1017
rect 1629 -921 1683 -903
rect 1629 -955 1639 -921
rect 1673 -955 1683 -921
rect 1629 -989 1683 -955
rect 1629 -1023 1639 -989
rect 1673 -1023 1683 -989
rect 1629 -1057 1683 -1023
rect 1629 -1091 1639 -1057
rect 1673 -1091 1683 -1057
rect 1629 -1103 1683 -1091
rect 1713 -915 1765 -903
rect 1713 -949 1723 -915
rect 1757 -949 1765 -915
rect 1713 -983 1765 -949
rect 1713 -1017 1723 -983
rect 1757 -1017 1765 -983
rect 1713 -1051 1765 -1017
rect 1713 -1085 1723 -1051
rect 1757 -1085 1765 -1051
rect 1713 -1103 1765 -1085
rect 203 -1811 255 -1793
rect -101 -1871 -49 -1835
rect -101 -1905 -93 -1871
rect -59 -1905 -49 -1871
rect -101 -1939 -49 -1905
rect -101 -1973 -93 -1939
rect -59 -1973 -49 -1939
rect -101 -1993 -49 -1973
rect -19 -1871 39 -1835
rect -19 -1905 -7 -1871
rect 27 -1905 39 -1871
rect -19 -1939 39 -1905
rect -19 -1973 -7 -1939
rect 27 -1973 39 -1939
rect -19 -1993 39 -1973
rect 69 -1858 121 -1835
rect 69 -1892 79 -1858
rect 113 -1892 121 -1858
rect 69 -1939 121 -1892
rect 69 -1973 79 -1939
rect 113 -1973 121 -1939
rect 69 -1993 121 -1973
rect 203 -1845 211 -1811
rect 245 -1845 255 -1811
rect 203 -1879 255 -1845
rect 203 -1913 211 -1879
rect 245 -1913 255 -1879
rect 203 -1947 255 -1913
rect 203 -1981 211 -1947
rect 245 -1981 255 -1947
rect 203 -1993 255 -1981
rect 285 -1830 339 -1793
rect 285 -1864 295 -1830
rect 329 -1864 339 -1830
rect 285 -1925 339 -1864
rect 285 -1959 295 -1925
rect 329 -1959 339 -1925
rect 285 -1993 339 -1959
rect 369 -1879 423 -1793
rect 369 -1913 379 -1879
rect 413 -1913 423 -1879
rect 369 -1947 423 -1913
rect 369 -1981 379 -1947
rect 413 -1981 423 -1947
rect 369 -1993 423 -1981
rect 453 -1830 507 -1793
rect 453 -1864 463 -1830
rect 497 -1864 507 -1830
rect 453 -1925 507 -1864
rect 453 -1959 463 -1925
rect 497 -1959 507 -1925
rect 453 -1993 507 -1959
rect 537 -1879 591 -1793
rect 537 -1913 547 -1879
rect 581 -1913 591 -1879
rect 537 -1947 591 -1913
rect 537 -1981 547 -1947
rect 581 -1981 591 -1947
rect 537 -1993 591 -1981
rect 621 -1805 673 -1793
rect 621 -1839 631 -1805
rect 665 -1839 673 -1805
rect 621 -1873 673 -1839
rect 621 -1907 631 -1873
rect 665 -1907 673 -1873
rect 621 -1941 673 -1907
rect 621 -1975 631 -1941
rect 665 -1975 673 -1941
rect 621 -1993 673 -1975
rect 743 -1811 795 -1793
rect 743 -1845 751 -1811
rect 785 -1845 795 -1811
rect 743 -1879 795 -1845
rect 743 -1913 751 -1879
rect 785 -1913 795 -1879
rect 743 -1947 795 -1913
rect 743 -1981 751 -1947
rect 785 -1981 795 -1947
rect 743 -1993 795 -1981
rect 825 -1830 879 -1793
rect 825 -1864 835 -1830
rect 869 -1864 879 -1830
rect 825 -1925 879 -1864
rect 825 -1959 835 -1925
rect 869 -1959 879 -1925
rect 825 -1993 879 -1959
rect 909 -1879 963 -1793
rect 909 -1913 919 -1879
rect 953 -1913 963 -1879
rect 909 -1947 963 -1913
rect 909 -1981 919 -1947
rect 953 -1981 963 -1947
rect 909 -1993 963 -1981
rect 993 -1830 1047 -1793
rect 993 -1864 1003 -1830
rect 1037 -1864 1047 -1830
rect 993 -1925 1047 -1864
rect 993 -1959 1003 -1925
rect 1037 -1959 1047 -1925
rect 993 -1993 1047 -1959
rect 1077 -1879 1131 -1793
rect 1077 -1913 1087 -1879
rect 1121 -1913 1131 -1879
rect 1077 -1947 1131 -1913
rect 1077 -1981 1087 -1947
rect 1121 -1981 1131 -1947
rect 1077 -1993 1131 -1981
rect 1161 -1805 1213 -1793
rect 1161 -1839 1171 -1805
rect 1205 -1839 1213 -1805
rect 1161 -1873 1213 -1839
rect 1161 -1907 1171 -1873
rect 1205 -1907 1213 -1873
rect 1161 -1941 1213 -1907
rect 1161 -1975 1171 -1941
rect 1205 -1975 1213 -1941
rect 1161 -1993 1213 -1975
rect 1295 -1811 1347 -1793
rect 1295 -1845 1303 -1811
rect 1337 -1845 1347 -1811
rect 1295 -1879 1347 -1845
rect 1295 -1913 1303 -1879
rect 1337 -1913 1347 -1879
rect 1295 -1947 1347 -1913
rect 1295 -1981 1303 -1947
rect 1337 -1981 1347 -1947
rect 1295 -1993 1347 -1981
rect 1377 -1830 1431 -1793
rect 1377 -1864 1387 -1830
rect 1421 -1864 1431 -1830
rect 1377 -1925 1431 -1864
rect 1377 -1959 1387 -1925
rect 1421 -1959 1431 -1925
rect 1377 -1993 1431 -1959
rect 1461 -1879 1515 -1793
rect 1461 -1913 1471 -1879
rect 1505 -1913 1515 -1879
rect 1461 -1947 1515 -1913
rect 1461 -1981 1471 -1947
rect 1505 -1981 1515 -1947
rect 1461 -1993 1515 -1981
rect 1545 -1830 1599 -1793
rect 1545 -1864 1555 -1830
rect 1589 -1864 1599 -1830
rect 1545 -1925 1599 -1864
rect 1545 -1959 1555 -1925
rect 1589 -1959 1599 -1925
rect 1545 -1993 1599 -1959
rect 1629 -1879 1683 -1793
rect 1629 -1913 1639 -1879
rect 1673 -1913 1683 -1879
rect 1629 -1947 1683 -1913
rect 1629 -1981 1639 -1947
rect 1673 -1981 1683 -1947
rect 1629 -1993 1683 -1981
rect 1713 -1805 1765 -1793
rect 1713 -1839 1723 -1805
rect 1757 -1839 1765 -1805
rect 1713 -1873 1765 -1839
rect 1713 -1907 1723 -1873
rect 1757 -1907 1765 -1873
rect 1713 -1941 1765 -1907
rect 1713 -1975 1723 -1941
rect 1757 -1975 1765 -1941
rect 1713 -1993 1765 -1975
rect -113 -2203 -61 -2183
rect -113 -2237 -105 -2203
rect -71 -2237 -61 -2203
rect -113 -2271 -61 -2237
rect -113 -2305 -105 -2271
rect -71 -2305 -61 -2271
rect -113 -2341 -61 -2305
rect -31 -2203 27 -2183
rect -31 -2237 -19 -2203
rect 15 -2237 27 -2203
rect -31 -2271 27 -2237
rect -31 -2305 -19 -2271
rect 15 -2305 27 -2271
rect -31 -2341 27 -2305
rect 57 -2203 109 -2183
rect 57 -2237 67 -2203
rect 101 -2237 109 -2203
rect 57 -2284 109 -2237
rect 57 -2318 67 -2284
rect 101 -2318 109 -2284
rect 57 -2341 109 -2318
rect 163 -2203 215 -2183
rect 163 -2237 171 -2203
rect 205 -2237 215 -2203
rect 163 -2271 215 -2237
rect 163 -2305 171 -2271
rect 205 -2305 215 -2271
rect 163 -2341 215 -2305
rect 245 -2203 303 -2183
rect 245 -2237 257 -2203
rect 291 -2237 303 -2203
rect 245 -2271 303 -2237
rect 245 -2305 257 -2271
rect 291 -2305 303 -2271
rect 245 -2341 303 -2305
rect 333 -2203 385 -2183
rect 333 -2237 343 -2203
rect 377 -2237 385 -2203
rect 333 -2284 385 -2237
rect 333 -2318 343 -2284
rect 377 -2318 385 -2284
rect 333 -2341 385 -2318
rect 439 -2203 491 -2183
rect 439 -2237 447 -2203
rect 481 -2237 491 -2203
rect 439 -2271 491 -2237
rect 439 -2305 447 -2271
rect 481 -2305 491 -2271
rect 439 -2341 491 -2305
rect 521 -2203 579 -2183
rect 521 -2237 533 -2203
rect 567 -2237 579 -2203
rect 521 -2271 579 -2237
rect 521 -2305 533 -2271
rect 567 -2305 579 -2271
rect 521 -2341 579 -2305
rect 609 -2203 661 -2183
rect 609 -2237 619 -2203
rect 653 -2237 661 -2203
rect 609 -2284 661 -2237
rect 609 -2318 619 -2284
rect 653 -2318 661 -2284
rect 609 -2341 661 -2318
rect 715 -2203 767 -2183
rect 715 -2237 723 -2203
rect 757 -2237 767 -2203
rect 715 -2284 767 -2237
rect 715 -2318 723 -2284
rect 757 -2318 767 -2284
rect 715 -2341 767 -2318
rect 797 -2203 855 -2183
rect 797 -2237 809 -2203
rect 843 -2237 855 -2203
rect 797 -2271 855 -2237
rect 797 -2305 809 -2271
rect 843 -2305 855 -2271
rect 797 -2341 855 -2305
rect 885 -2203 937 -2183
rect 885 -2237 895 -2203
rect 929 -2237 937 -2203
rect 885 -2271 937 -2237
rect 885 -2305 895 -2271
rect 929 -2305 937 -2271
rect 885 -2341 937 -2305
rect 991 -2203 1043 -2183
rect 991 -2237 999 -2203
rect 1033 -2237 1043 -2203
rect 991 -2271 1043 -2237
rect 991 -2305 999 -2271
rect 1033 -2305 1043 -2271
rect 991 -2341 1043 -2305
rect 1073 -2203 1131 -2183
rect 1073 -2237 1085 -2203
rect 1119 -2237 1131 -2203
rect 1073 -2271 1131 -2237
rect 1073 -2305 1085 -2271
rect 1119 -2305 1131 -2271
rect 1073 -2341 1131 -2305
rect 1161 -2203 1213 -2183
rect 1161 -2237 1171 -2203
rect 1205 -2237 1213 -2203
rect 1161 -2284 1213 -2237
rect 1161 -2318 1171 -2284
rect 1205 -2318 1213 -2284
rect 1161 -2341 1213 -2318
rect 1267 -2203 1319 -2183
rect 1267 -2237 1275 -2203
rect 1309 -2237 1319 -2203
rect 1267 -2284 1319 -2237
rect 1267 -2318 1275 -2284
rect 1309 -2318 1319 -2284
rect 1267 -2341 1319 -2318
rect 1349 -2203 1407 -2183
rect 1349 -2237 1361 -2203
rect 1395 -2237 1407 -2203
rect 1349 -2271 1407 -2237
rect 1349 -2305 1361 -2271
rect 1395 -2305 1407 -2271
rect 1349 -2341 1407 -2305
rect 1437 -2203 1489 -2183
rect 1437 -2237 1447 -2203
rect 1481 -2237 1489 -2203
rect 1437 -2271 1489 -2237
rect 1437 -2305 1447 -2271
rect 1481 -2305 1489 -2271
rect 1437 -2341 1489 -2305
rect 1543 -2203 1595 -2183
rect 1543 -2237 1551 -2203
rect 1585 -2237 1595 -2203
rect 1543 -2271 1595 -2237
rect 1543 -2305 1551 -2271
rect 1585 -2305 1595 -2271
rect 1543 -2341 1595 -2305
rect 1625 -2203 1683 -2183
rect 1625 -2237 1637 -2203
rect 1671 -2237 1683 -2203
rect 1625 -2271 1683 -2237
rect 1625 -2305 1637 -2271
rect 1671 -2305 1683 -2271
rect 1625 -2341 1683 -2305
rect 1713 -2203 1765 -2183
rect 1713 -2237 1723 -2203
rect 1757 -2237 1765 -2203
rect 1713 -2284 1765 -2237
rect 1713 -2318 1723 -2284
rect 1757 -2318 1765 -2284
rect 1713 -2341 1765 -2318
<< ndiffc >>
rect -125 -1337 -91 -1303
rect -41 -1269 -7 -1235
rect -41 -1337 -7 -1303
rect 43 -1337 77 -1303
rect 127 -1269 161 -1235
rect 127 -1337 161 -1303
rect 211 -1337 245 -1303
rect 295 -1269 329 -1235
rect 295 -1337 329 -1303
rect 379 -1337 413 -1303
rect 463 -1269 497 -1235
rect 463 -1337 497 -1303
rect 547 -1337 581 -1303
rect 631 -1269 665 -1235
rect 631 -1337 665 -1303
rect 715 -1337 749 -1303
rect 799 -1269 833 -1235
rect 799 -1337 833 -1303
rect 883 -1337 917 -1303
rect 967 -1269 1001 -1235
rect 967 -1337 1001 -1303
rect 1051 -1337 1085 -1303
rect 1135 -1269 1169 -1235
rect 1135 -1337 1169 -1303
rect 1219 -1337 1253 -1303
rect 1303 -1269 1337 -1235
rect 1303 -1337 1337 -1303
rect 1387 -1337 1421 -1303
rect 1471 -1269 1505 -1235
rect 1471 -1337 1505 -1303
rect 1555 -1337 1589 -1303
rect 1639 -1269 1673 -1235
rect 1639 -1337 1673 -1303
rect 1723 -1269 1757 -1235
rect 1723 -1337 1757 -1303
rect -93 -1602 -59 -1568
rect -7 -1589 27 -1555
rect 79 -1619 113 -1585
rect 211 -1589 245 -1555
rect 211 -1657 245 -1623
rect 295 -1625 329 -1591
rect 379 -1593 413 -1559
rect 463 -1625 497 -1591
rect 547 -1593 581 -1559
rect 631 -1625 665 -1591
rect 751 -1589 785 -1555
rect 751 -1657 785 -1623
rect 835 -1625 869 -1591
rect 919 -1593 953 -1559
rect 1003 -1625 1037 -1591
rect 1087 -1593 1121 -1559
rect 1171 -1625 1205 -1591
rect 1303 -1589 1337 -1555
rect 1303 -1657 1337 -1623
rect 1387 -1625 1421 -1591
rect 1471 -1593 1505 -1559
rect 1555 -1625 1589 -1591
rect 1639 -1593 1673 -1559
rect 1723 -1625 1757 -1591
rect -105 -2608 -71 -2574
rect -19 -2621 15 -2587
rect 67 -2591 101 -2557
rect 171 -2608 205 -2574
rect 257 -2621 291 -2587
rect 343 -2591 377 -2557
rect 447 -2608 481 -2574
rect 533 -2621 567 -2587
rect 619 -2591 653 -2557
rect 723 -2591 757 -2557
rect 809 -2621 843 -2587
rect 895 -2608 929 -2574
rect 999 -2608 1033 -2574
rect 1085 -2621 1119 -2587
rect 1171 -2591 1205 -2557
rect 1275 -2591 1309 -2557
rect 1361 -2621 1395 -2587
rect 1447 -2608 1481 -2574
rect 1551 -2608 1585 -2574
rect 1637 -2621 1671 -2587
rect 1723 -2591 1757 -2557
<< pdiffc >>
rect -125 -949 -91 -915
rect -125 -1017 -91 -983
rect -41 -955 -7 -921
rect -41 -1023 -7 -989
rect -41 -1091 -7 -1057
rect 43 -949 77 -915
rect 43 -1017 77 -983
rect 127 -955 161 -921
rect 127 -1023 161 -989
rect 127 -1091 161 -1057
rect 211 -949 245 -915
rect 211 -1017 245 -983
rect 295 -955 329 -921
rect 295 -1023 329 -989
rect 295 -1091 329 -1057
rect 379 -949 413 -915
rect 379 -1017 413 -983
rect 463 -955 497 -921
rect 463 -1023 497 -989
rect 463 -1091 497 -1057
rect 547 -949 581 -915
rect 547 -1017 581 -983
rect 631 -955 665 -921
rect 631 -1023 665 -989
rect 631 -1091 665 -1057
rect 715 -949 749 -915
rect 715 -1017 749 -983
rect 799 -955 833 -921
rect 799 -1023 833 -989
rect 799 -1091 833 -1057
rect 883 -949 917 -915
rect 883 -1017 917 -983
rect 967 -955 1001 -921
rect 967 -1023 1001 -989
rect 967 -1091 1001 -1057
rect 1051 -949 1085 -915
rect 1051 -1017 1085 -983
rect 1135 -955 1169 -921
rect 1135 -1023 1169 -989
rect 1135 -1091 1169 -1057
rect 1219 -949 1253 -915
rect 1219 -1017 1253 -983
rect 1303 -955 1337 -921
rect 1303 -1023 1337 -989
rect 1303 -1091 1337 -1057
rect 1387 -949 1421 -915
rect 1387 -1017 1421 -983
rect 1471 -955 1505 -921
rect 1471 -1023 1505 -989
rect 1471 -1091 1505 -1057
rect 1555 -949 1589 -915
rect 1555 -1017 1589 -983
rect 1639 -955 1673 -921
rect 1639 -1023 1673 -989
rect 1639 -1091 1673 -1057
rect 1723 -949 1757 -915
rect 1723 -1017 1757 -983
rect 1723 -1085 1757 -1051
rect -93 -1905 -59 -1871
rect -93 -1973 -59 -1939
rect -7 -1905 27 -1871
rect -7 -1973 27 -1939
rect 79 -1892 113 -1858
rect 79 -1973 113 -1939
rect 211 -1845 245 -1811
rect 211 -1913 245 -1879
rect 211 -1981 245 -1947
rect 295 -1864 329 -1830
rect 295 -1959 329 -1925
rect 379 -1913 413 -1879
rect 379 -1981 413 -1947
rect 463 -1864 497 -1830
rect 463 -1959 497 -1925
rect 547 -1913 581 -1879
rect 547 -1981 581 -1947
rect 631 -1839 665 -1805
rect 631 -1907 665 -1873
rect 631 -1975 665 -1941
rect 751 -1845 785 -1811
rect 751 -1913 785 -1879
rect 751 -1981 785 -1947
rect 835 -1864 869 -1830
rect 835 -1959 869 -1925
rect 919 -1913 953 -1879
rect 919 -1981 953 -1947
rect 1003 -1864 1037 -1830
rect 1003 -1959 1037 -1925
rect 1087 -1913 1121 -1879
rect 1087 -1981 1121 -1947
rect 1171 -1839 1205 -1805
rect 1171 -1907 1205 -1873
rect 1171 -1975 1205 -1941
rect 1303 -1845 1337 -1811
rect 1303 -1913 1337 -1879
rect 1303 -1981 1337 -1947
rect 1387 -1864 1421 -1830
rect 1387 -1959 1421 -1925
rect 1471 -1913 1505 -1879
rect 1471 -1981 1505 -1947
rect 1555 -1864 1589 -1830
rect 1555 -1959 1589 -1925
rect 1639 -1913 1673 -1879
rect 1639 -1981 1673 -1947
rect 1723 -1839 1757 -1805
rect 1723 -1907 1757 -1873
rect 1723 -1975 1757 -1941
rect -105 -2237 -71 -2203
rect -105 -2305 -71 -2271
rect -19 -2237 15 -2203
rect -19 -2305 15 -2271
rect 67 -2237 101 -2203
rect 67 -2318 101 -2284
rect 171 -2237 205 -2203
rect 171 -2305 205 -2271
rect 257 -2237 291 -2203
rect 257 -2305 291 -2271
rect 343 -2237 377 -2203
rect 343 -2318 377 -2284
rect 447 -2237 481 -2203
rect 447 -2305 481 -2271
rect 533 -2237 567 -2203
rect 533 -2305 567 -2271
rect 619 -2237 653 -2203
rect 619 -2318 653 -2284
rect 723 -2237 757 -2203
rect 723 -2318 757 -2284
rect 809 -2237 843 -2203
rect 809 -2305 843 -2271
rect 895 -2237 929 -2203
rect 895 -2305 929 -2271
rect 999 -2237 1033 -2203
rect 999 -2305 1033 -2271
rect 1085 -2237 1119 -2203
rect 1085 -2305 1119 -2271
rect 1171 -2237 1205 -2203
rect 1171 -2318 1205 -2284
rect 1275 -2237 1309 -2203
rect 1275 -2318 1309 -2284
rect 1361 -2237 1395 -2203
rect 1361 -2305 1395 -2271
rect 1447 -2237 1481 -2203
rect 1447 -2305 1481 -2271
rect 1551 -2237 1585 -2203
rect 1551 -2305 1585 -2271
rect 1637 -2237 1671 -2203
rect 1637 -2305 1671 -2271
rect 1723 -2237 1757 -2203
rect 1723 -2318 1757 -2284
<< psubdiff >>
rect -118 -1463 -89 -1429
rect -55 -1430 85 -1429
rect -55 -1463 -5 -1430
rect -118 -1464 -5 -1463
rect 29 -1463 85 -1430
rect 119 -1463 177 -1429
rect 211 -1430 545 -1429
rect 211 -1463 267 -1430
rect 29 -1464 267 -1463
rect 301 -1464 361 -1430
rect 395 -1464 452 -1430
rect 486 -1463 545 -1430
rect 579 -1430 1453 -1429
rect 579 -1463 636 -1430
rect 486 -1464 636 -1463
rect 670 -1464 716 -1430
rect 750 -1464 809 -1430
rect 843 -1464 901 -1430
rect 935 -1464 994 -1430
rect 1028 -1464 1085 -1430
rect 1119 -1464 1177 -1430
rect 1211 -1464 1270 -1430
rect 1304 -1464 1361 -1430
rect 1395 -1463 1453 -1430
rect 1487 -1430 1790 -1429
rect 1487 -1463 1545 -1430
rect 1395 -1464 1545 -1463
rect 1579 -1464 1640 -1430
rect 1674 -1464 1728 -1430
rect 1762 -1464 1790 -1430
rect -133 -2698 -19 -2697
rect -133 -2732 -109 -2698
rect -75 -2731 -19 -2698
rect 15 -2731 73 -2697
rect 107 -2731 165 -2697
rect 199 -2731 257 -2697
rect 291 -2731 349 -2697
rect 383 -2731 441 -2697
rect 475 -2731 533 -2697
rect 567 -2731 625 -2697
rect 659 -2731 717 -2697
rect 751 -2731 809 -2697
rect 843 -2731 901 -2697
rect 935 -2731 993 -2697
rect 1027 -2731 1085 -2697
rect 1119 -2731 1177 -2697
rect 1211 -2698 1361 -2697
rect 1211 -2731 1269 -2698
rect -75 -2732 1269 -2731
rect 1303 -2731 1361 -2698
rect 1395 -2731 1453 -2697
rect 1487 -2731 1545 -2697
rect 1579 -2731 1637 -2697
rect 1671 -2731 1717 -2697
rect 1751 -2731 1775 -2697
rect 1303 -2732 1775 -2731
<< nsubdiff >>
rect -151 -805 1757 -804
rect -151 -839 -111 -805
rect -77 -839 -19 -805
rect 15 -839 73 -805
rect 107 -839 165 -805
rect 199 -839 257 -805
rect 291 -839 349 -805
rect 383 -839 441 -805
rect 475 -839 533 -805
rect 567 -839 625 -805
rect 659 -839 717 -805
rect 751 -839 809 -805
rect 843 -839 901 -805
rect 935 -839 993 -805
rect 1027 -839 1085 -805
rect 1119 -839 1177 -805
rect 1211 -839 1269 -805
rect 1303 -839 1361 -805
rect 1395 -839 1453 -805
rect 1487 -839 1545 -805
rect 1579 -839 1637 -805
rect 1671 -839 1757 -805
rect -125 -2105 -101 -2071
rect -67 -2072 269 -2071
rect -67 -2105 -5 -2072
rect -125 -2106 -5 -2105
rect 29 -2106 88 -2072
rect 122 -2106 177 -2072
rect 211 -2105 269 -2072
rect 303 -2072 453 -2071
rect 303 -2105 360 -2072
rect 211 -2106 360 -2105
rect 394 -2105 453 -2072
rect 487 -2105 545 -2071
rect 579 -2072 809 -2071
rect 579 -2105 639 -2072
rect 394 -2106 639 -2105
rect 673 -2106 718 -2072
rect 752 -2105 809 -2072
rect 843 -2072 1637 -2071
rect 843 -2105 901 -2072
rect 752 -2106 901 -2105
rect 935 -2106 993 -2072
rect 1027 -2106 1085 -2072
rect 1119 -2106 1176 -2072
rect 1210 -2106 1269 -2072
rect 1303 -2106 1362 -2072
rect 1396 -2106 1454 -2072
rect 1488 -2106 1545 -2072
rect 1579 -2105 1637 -2072
rect 1671 -2105 1724 -2071
rect 1758 -2105 1783 -2071
rect 1579 -2106 1783 -2105
<< psubdiffcont >>
rect -89 -1463 -55 -1429
rect -5 -1464 29 -1430
rect 85 -1463 119 -1429
rect 177 -1463 211 -1429
rect 267 -1464 301 -1430
rect 361 -1464 395 -1430
rect 452 -1464 486 -1430
rect 545 -1463 579 -1429
rect 636 -1464 670 -1430
rect 716 -1464 750 -1430
rect 809 -1464 843 -1430
rect 901 -1464 935 -1430
rect 994 -1464 1028 -1430
rect 1085 -1464 1119 -1430
rect 1177 -1464 1211 -1430
rect 1270 -1464 1304 -1430
rect 1361 -1464 1395 -1430
rect 1453 -1463 1487 -1429
rect 1545 -1464 1579 -1430
rect 1640 -1464 1674 -1430
rect 1728 -1464 1762 -1430
rect -109 -2732 -75 -2698
rect -19 -2731 15 -2697
rect 73 -2731 107 -2697
rect 165 -2731 199 -2697
rect 257 -2731 291 -2697
rect 349 -2731 383 -2697
rect 441 -2731 475 -2697
rect 533 -2731 567 -2697
rect 625 -2731 659 -2697
rect 717 -2731 751 -2697
rect 809 -2731 843 -2697
rect 901 -2731 935 -2697
rect 993 -2731 1027 -2697
rect 1085 -2731 1119 -2697
rect 1177 -2731 1211 -2697
rect 1269 -2732 1303 -2698
rect 1361 -2731 1395 -2697
rect 1453 -2731 1487 -2697
rect 1545 -2731 1579 -2697
rect 1637 -2731 1671 -2697
rect 1717 -2731 1751 -2697
<< nsubdiffcont >>
rect -111 -839 -77 -805
rect -19 -839 15 -805
rect 73 -839 107 -805
rect 165 -839 199 -805
rect 257 -839 291 -805
rect 349 -839 383 -805
rect 441 -839 475 -805
rect 533 -839 567 -805
rect 625 -839 659 -805
rect 717 -839 751 -805
rect 809 -839 843 -805
rect 901 -839 935 -805
rect 993 -839 1027 -805
rect 1085 -839 1119 -805
rect 1177 -839 1211 -805
rect 1269 -839 1303 -805
rect 1361 -839 1395 -805
rect 1453 -839 1487 -805
rect 1545 -839 1579 -805
rect 1637 -839 1671 -805
rect -101 -2105 -67 -2071
rect -5 -2106 29 -2072
rect 88 -2106 122 -2072
rect 177 -2106 211 -2072
rect 269 -2105 303 -2071
rect 360 -2106 394 -2072
rect 453 -2105 487 -2071
rect 545 -2105 579 -2071
rect 639 -2106 673 -2072
rect 718 -2106 752 -2072
rect 809 -2105 843 -2071
rect 901 -2106 935 -2072
rect 993 -2106 1027 -2072
rect 1085 -2106 1119 -2072
rect 1176 -2106 1210 -2072
rect 1269 -2106 1303 -2072
rect 1362 -2106 1396 -2072
rect 1454 -2106 1488 -2072
rect 1545 -2106 1579 -2072
rect 1637 -2105 1671 -2071
rect 1724 -2105 1758 -2071
<< poly >>
rect -81 -903 -51 -877
rect 3 -903 33 -877
rect 87 -903 117 -877
rect 171 -903 201 -877
rect 255 -903 285 -877
rect 339 -903 369 -877
rect 423 -903 453 -877
rect 507 -903 537 -877
rect 591 -903 621 -877
rect 675 -903 705 -877
rect 759 -903 789 -877
rect 843 -903 873 -877
rect 927 -903 957 -877
rect 1011 -903 1041 -877
rect 1095 -903 1125 -877
rect 1179 -903 1209 -877
rect 1263 -903 1293 -877
rect 1347 -903 1377 -877
rect 1431 -903 1461 -877
rect 1515 -903 1545 -877
rect 1599 -903 1629 -877
rect 1683 -903 1713 -877
rect -81 -1141 -51 -1103
rect 3 -1141 33 -1103
rect 87 -1141 117 -1103
rect 171 -1141 201 -1103
rect 255 -1141 285 -1103
rect 339 -1141 369 -1103
rect 423 -1141 453 -1103
rect 507 -1141 537 -1103
rect 591 -1141 621 -1103
rect 675 -1141 705 -1103
rect 759 -1141 789 -1103
rect 843 -1141 873 -1103
rect 927 -1141 957 -1103
rect 1011 -1141 1041 -1103
rect 1095 -1141 1125 -1103
rect 1179 -1141 1209 -1103
rect -85 -1151 1209 -1141
rect -85 -1185 -69 -1151
rect -35 -1185 -1 -1151
rect 33 -1185 67 -1151
rect 101 -1185 135 -1151
rect 169 -1185 203 -1151
rect 237 -1185 271 -1151
rect 305 -1185 339 -1151
rect 373 -1185 407 -1151
rect 441 -1185 475 -1151
rect 509 -1185 543 -1151
rect 577 -1185 611 -1151
rect 645 -1185 679 -1151
rect 713 -1185 747 -1151
rect 781 -1185 815 -1151
rect 849 -1185 883 -1151
rect 917 -1185 951 -1151
rect 985 -1185 1019 -1151
rect 1053 -1185 1087 -1151
rect 1121 -1185 1155 -1151
rect 1189 -1185 1209 -1151
rect -85 -1195 1209 -1185
rect -81 -1223 -51 -1195
rect 3 -1223 33 -1195
rect 87 -1223 117 -1195
rect 171 -1223 201 -1195
rect 255 -1223 285 -1195
rect 339 -1223 369 -1195
rect 423 -1223 453 -1195
rect 507 -1223 537 -1195
rect 591 -1223 621 -1195
rect 675 -1223 705 -1195
rect 759 -1223 789 -1195
rect 843 -1223 873 -1195
rect 927 -1223 957 -1195
rect 1011 -1223 1041 -1195
rect 1095 -1223 1125 -1195
rect 1179 -1223 1209 -1195
rect 1263 -1141 1293 -1103
rect 1347 -1141 1377 -1103
rect 1431 -1141 1461 -1103
rect 1515 -1141 1545 -1103
rect 1599 -1141 1629 -1103
rect 1683 -1141 1713 -1103
rect 1263 -1151 1713 -1141
rect 1263 -1185 1315 -1151
rect 1349 -1185 1383 -1151
rect 1417 -1185 1451 -1151
rect 1485 -1185 1519 -1151
rect 1553 -1185 1587 -1151
rect 1621 -1185 1655 -1151
rect 1689 -1185 1713 -1151
rect 1263 -1195 1713 -1185
rect 1263 -1223 1293 -1195
rect 1347 -1223 1377 -1195
rect 1431 -1223 1461 -1195
rect 1515 -1223 1545 -1195
rect 1599 -1223 1629 -1195
rect 1683 -1223 1713 -1195
rect -81 -1379 -51 -1353
rect 3 -1379 33 -1353
rect 87 -1379 117 -1353
rect 171 -1379 201 -1353
rect 255 -1379 285 -1353
rect 339 -1379 369 -1353
rect 423 -1379 453 -1353
rect 507 -1379 537 -1353
rect 591 -1379 621 -1353
rect 675 -1379 705 -1353
rect 759 -1379 789 -1353
rect 843 -1379 873 -1353
rect 927 -1379 957 -1353
rect 1011 -1379 1041 -1353
rect 1095 -1379 1125 -1353
rect 1179 -1379 1209 -1353
rect 1263 -1379 1293 -1353
rect 1347 -1379 1377 -1353
rect 1431 -1379 1461 -1353
rect 1515 -1379 1545 -1353
rect 1599 -1379 1629 -1353
rect 1683 -1379 1713 -1353
rect -49 -1543 -19 -1517
rect 39 -1543 69 -1517
rect 255 -1543 285 -1517
rect 339 -1543 369 -1517
rect 423 -1543 453 -1517
rect 507 -1543 537 -1517
rect 591 -1543 621 -1517
rect 795 -1543 825 -1517
rect 879 -1543 909 -1517
rect 963 -1543 993 -1517
rect 1047 -1543 1077 -1517
rect 1131 -1543 1161 -1517
rect 1347 -1543 1377 -1517
rect 1431 -1543 1461 -1517
rect 1515 -1543 1545 -1517
rect 1599 -1543 1629 -1517
rect 1683 -1543 1713 -1517
rect -49 -1662 -19 -1647
rect -55 -1686 -19 -1662
rect -55 -1695 -25 -1686
rect -101 -1711 -25 -1695
rect 39 -1708 69 -1647
rect 255 -1701 285 -1673
rect 339 -1701 369 -1673
rect 423 -1701 453 -1673
rect 507 -1701 537 -1673
rect 591 -1699 621 -1673
rect -101 -1745 -91 -1711
rect -57 -1745 -25 -1711
rect -101 -1761 -25 -1745
rect -55 -1796 -25 -1761
rect 17 -1724 71 -1708
rect 17 -1758 27 -1724
rect 61 -1758 71 -1724
rect 17 -1774 71 -1758
rect 255 -1711 538 -1701
rect 255 -1745 488 -1711
rect 522 -1745 538 -1711
rect 255 -1755 538 -1745
rect 591 -1711 672 -1699
rect 591 -1745 622 -1711
rect 656 -1745 672 -1711
rect -55 -1820 -19 -1796
rect -49 -1835 -19 -1820
rect 39 -1835 69 -1774
rect 255 -1793 285 -1755
rect 339 -1793 369 -1755
rect 423 -1793 453 -1755
rect 507 -1793 537 -1755
rect 591 -1757 672 -1745
rect 795 -1701 825 -1673
rect 879 -1701 909 -1673
rect 963 -1701 993 -1673
rect 1047 -1701 1077 -1673
rect 1131 -1699 1161 -1673
rect 795 -1711 1078 -1701
rect 795 -1745 1028 -1711
rect 1062 -1745 1078 -1711
rect 795 -1755 1078 -1745
rect 1131 -1711 1212 -1699
rect 1131 -1745 1162 -1711
rect 1196 -1745 1212 -1711
rect 591 -1793 621 -1757
rect 795 -1793 825 -1755
rect 879 -1793 909 -1755
rect 963 -1793 993 -1755
rect 1047 -1793 1077 -1755
rect 1131 -1757 1212 -1745
rect 1347 -1701 1377 -1673
rect 1431 -1701 1461 -1673
rect 1515 -1701 1545 -1673
rect 1599 -1701 1629 -1673
rect 1683 -1699 1713 -1673
rect 1347 -1711 1630 -1701
rect 1347 -1745 1580 -1711
rect 1614 -1745 1630 -1711
rect 1347 -1755 1630 -1745
rect 1683 -1711 1764 -1699
rect 1683 -1745 1714 -1711
rect 1748 -1745 1764 -1711
rect 1131 -1793 1161 -1757
rect 1347 -1793 1377 -1755
rect 1431 -1793 1461 -1755
rect 1515 -1793 1545 -1755
rect 1599 -1793 1629 -1755
rect 1683 -1757 1764 -1745
rect 1683 -1793 1713 -1757
rect -49 -2019 -19 -1993
rect 39 -2019 69 -1993
rect 255 -2019 285 -1993
rect 339 -2019 369 -1993
rect 423 -2019 453 -1993
rect 507 -2019 537 -1993
rect 591 -2019 621 -1993
rect 795 -2019 825 -1993
rect 879 -2019 909 -1993
rect 963 -2019 993 -1993
rect 1047 -2019 1077 -1993
rect 1131 -2019 1161 -1993
rect 1347 -2019 1377 -1993
rect 1431 -2019 1461 -1993
rect 1515 -2019 1545 -1993
rect 1599 -2019 1629 -1993
rect 1683 -2019 1713 -1993
rect -61 -2183 -31 -2157
rect 27 -2183 57 -2157
rect 215 -2183 245 -2157
rect 303 -2183 333 -2157
rect 491 -2183 521 -2157
rect 579 -2183 609 -2157
rect 767 -2183 797 -2157
rect 855 -2183 885 -2157
rect 1043 -2183 1073 -2157
rect 1131 -2183 1161 -2157
rect 1319 -2183 1349 -2157
rect 1407 -2183 1437 -2157
rect 1595 -2183 1625 -2157
rect 1683 -2183 1713 -2157
rect -61 -2356 -31 -2341
rect -67 -2380 -31 -2356
rect -67 -2415 -37 -2380
rect 27 -2402 57 -2341
rect 215 -2356 245 -2341
rect 209 -2380 245 -2356
rect -113 -2431 -37 -2415
rect -113 -2465 -103 -2431
rect -69 -2465 -37 -2431
rect -113 -2481 -37 -2465
rect 5 -2418 59 -2402
rect 209 -2415 239 -2380
rect 303 -2402 333 -2341
rect 491 -2356 521 -2341
rect 485 -2380 521 -2356
rect 5 -2452 15 -2418
rect 49 -2452 59 -2418
rect 5 -2468 59 -2452
rect 163 -2431 239 -2415
rect 163 -2465 173 -2431
rect 207 -2465 239 -2431
rect -67 -2490 -37 -2481
rect -67 -2514 -31 -2490
rect -61 -2529 -31 -2514
rect 27 -2529 57 -2468
rect 163 -2481 239 -2465
rect 281 -2418 335 -2402
rect 485 -2415 515 -2380
rect 579 -2402 609 -2341
rect 767 -2402 797 -2341
rect 855 -2356 885 -2341
rect 1043 -2356 1073 -2341
rect 855 -2380 891 -2356
rect 281 -2452 291 -2418
rect 325 -2452 335 -2418
rect 281 -2468 335 -2452
rect 439 -2431 515 -2415
rect 439 -2465 449 -2431
rect 483 -2465 515 -2431
rect 209 -2490 239 -2481
rect 209 -2514 245 -2490
rect 215 -2529 245 -2514
rect 303 -2529 333 -2468
rect 439 -2481 515 -2465
rect 557 -2418 611 -2402
rect 557 -2452 567 -2418
rect 601 -2452 611 -2418
rect 557 -2468 611 -2452
rect 765 -2418 819 -2402
rect 765 -2452 775 -2418
rect 809 -2452 819 -2418
rect 765 -2468 819 -2452
rect 861 -2415 891 -2380
rect 1037 -2380 1073 -2356
rect 1037 -2415 1067 -2380
rect 1131 -2402 1161 -2341
rect 1319 -2402 1349 -2341
rect 1407 -2356 1437 -2341
rect 1595 -2356 1625 -2341
rect 1407 -2380 1443 -2356
rect 861 -2431 937 -2415
rect 861 -2465 893 -2431
rect 927 -2465 937 -2431
rect 485 -2490 515 -2481
rect 485 -2514 521 -2490
rect 491 -2529 521 -2514
rect 579 -2529 609 -2468
rect 767 -2529 797 -2468
rect 861 -2481 937 -2465
rect 991 -2431 1067 -2415
rect 991 -2465 1001 -2431
rect 1035 -2465 1067 -2431
rect 991 -2481 1067 -2465
rect 1109 -2418 1163 -2402
rect 1109 -2452 1119 -2418
rect 1153 -2452 1163 -2418
rect 1109 -2468 1163 -2452
rect 1317 -2418 1371 -2402
rect 1317 -2452 1327 -2418
rect 1361 -2452 1371 -2418
rect 1317 -2468 1371 -2452
rect 1413 -2415 1443 -2380
rect 1589 -2380 1625 -2356
rect 1589 -2415 1619 -2380
rect 1683 -2402 1713 -2341
rect 1413 -2431 1489 -2415
rect 1413 -2465 1445 -2431
rect 1479 -2465 1489 -2431
rect 861 -2490 891 -2481
rect 855 -2514 891 -2490
rect 1037 -2490 1067 -2481
rect 1037 -2514 1073 -2490
rect 855 -2529 885 -2514
rect 1043 -2529 1073 -2514
rect 1131 -2529 1161 -2468
rect 1319 -2529 1349 -2468
rect 1413 -2481 1489 -2465
rect 1543 -2431 1619 -2415
rect 1543 -2465 1553 -2431
rect 1587 -2465 1619 -2431
rect 1543 -2481 1619 -2465
rect 1661 -2418 1715 -2402
rect 1661 -2452 1671 -2418
rect 1705 -2452 1715 -2418
rect 1661 -2468 1715 -2452
rect 1413 -2490 1443 -2481
rect 1407 -2514 1443 -2490
rect 1589 -2490 1619 -2481
rect 1589 -2514 1625 -2490
rect 1407 -2529 1437 -2514
rect 1595 -2529 1625 -2514
rect 1683 -2529 1713 -2468
rect -61 -2659 -31 -2633
rect 27 -2659 57 -2633
rect 215 -2659 245 -2633
rect 303 -2659 333 -2633
rect 491 -2659 521 -2633
rect 579 -2659 609 -2633
rect 767 -2659 797 -2633
rect 855 -2659 885 -2633
rect 1043 -2659 1073 -2633
rect 1131 -2659 1161 -2633
rect 1319 -2659 1349 -2633
rect 1407 -2659 1437 -2633
rect 1595 -2659 1625 -2633
rect 1683 -2659 1713 -2633
<< polycont >>
rect -69 -1185 -35 -1151
rect -1 -1185 33 -1151
rect 67 -1185 101 -1151
rect 135 -1185 169 -1151
rect 203 -1185 237 -1151
rect 271 -1185 305 -1151
rect 339 -1185 373 -1151
rect 407 -1185 441 -1151
rect 475 -1185 509 -1151
rect 543 -1185 577 -1151
rect 611 -1185 645 -1151
rect 679 -1185 713 -1151
rect 747 -1185 781 -1151
rect 815 -1185 849 -1151
rect 883 -1185 917 -1151
rect 951 -1185 985 -1151
rect 1019 -1185 1053 -1151
rect 1087 -1185 1121 -1151
rect 1155 -1185 1189 -1151
rect 1315 -1185 1349 -1151
rect 1383 -1185 1417 -1151
rect 1451 -1185 1485 -1151
rect 1519 -1185 1553 -1151
rect 1587 -1185 1621 -1151
rect 1655 -1185 1689 -1151
rect -91 -1745 -57 -1711
rect 27 -1758 61 -1724
rect 488 -1745 522 -1711
rect 622 -1745 656 -1711
rect 1028 -1745 1062 -1711
rect 1162 -1745 1196 -1711
rect 1580 -1745 1614 -1711
rect 1714 -1745 1748 -1711
rect -103 -2465 -69 -2431
rect 15 -2452 49 -2418
rect 173 -2465 207 -2431
rect 291 -2452 325 -2418
rect 449 -2465 483 -2431
rect 567 -2452 601 -2418
rect 775 -2452 809 -2418
rect 893 -2465 927 -2431
rect 1001 -2465 1035 -2431
rect 1119 -2452 1153 -2418
rect 1327 -2452 1361 -2418
rect 1445 -2465 1479 -2431
rect 1553 -2465 1587 -2431
rect 1671 -2452 1705 -2418
<< locali >>
rect -232 -805 1792 -804
rect -232 -839 -111 -805
rect -232 -873 -203 -839
rect -169 -873 -111 -839
rect -77 -873 -19 -805
rect 15 -873 73 -805
rect 107 -873 165 -805
rect 199 -873 257 -805
rect 291 -873 349 -805
rect 383 -873 441 -805
rect 475 -873 533 -805
rect 567 -873 625 -805
rect 659 -873 717 -805
rect 751 -873 809 -805
rect 843 -873 901 -805
rect 935 -873 993 -805
rect 1027 -873 1085 -805
rect 1119 -873 1177 -805
rect 1211 -873 1269 -805
rect 1303 -873 1361 -805
rect 1395 -873 1453 -805
rect 1487 -873 1545 -805
rect 1579 -873 1637 -805
rect 1671 -839 1792 -805
rect 1671 -873 1729 -839
rect 1763 -873 1792 -839
rect -125 -915 -91 -873
rect -215 -1077 -160 -928
rect -125 -983 -91 -949
rect -125 -1033 -91 -1017
rect -57 -921 9 -907
rect -57 -955 -41 -921
rect -7 -955 9 -921
rect -57 -989 9 -955
rect -57 -1023 -41 -989
rect -7 -1023 9 -989
rect -57 -1057 9 -1023
rect 43 -915 77 -873
rect 43 -983 77 -949
rect 43 -1033 77 -1017
rect 111 -921 177 -907
rect 111 -955 127 -921
rect 161 -955 177 -921
rect 111 -989 177 -955
rect 111 -1023 127 -989
rect 161 -1023 177 -989
rect -57 -1077 -41 -1057
rect -215 -1091 -41 -1077
rect -7 -1077 9 -1057
rect 111 -1057 177 -1023
rect 211 -915 245 -873
rect 211 -983 245 -949
rect 211 -1033 245 -1017
rect 279 -921 345 -907
rect 279 -955 295 -921
rect 329 -955 345 -921
rect 279 -989 345 -955
rect 279 -1023 295 -989
rect 329 -1023 345 -989
rect 111 -1077 127 -1057
rect -7 -1091 127 -1077
rect 161 -1077 177 -1057
rect 279 -1057 345 -1023
rect 379 -915 413 -873
rect 379 -983 413 -949
rect 379 -1033 413 -1017
rect 447 -921 513 -907
rect 447 -955 463 -921
rect 497 -955 513 -921
rect 447 -989 513 -955
rect 447 -1023 463 -989
rect 497 -1023 513 -989
rect 279 -1077 295 -1057
rect 161 -1091 295 -1077
rect 329 -1077 345 -1057
rect 447 -1057 513 -1023
rect 547 -915 581 -873
rect 547 -983 581 -949
rect 547 -1033 581 -1017
rect 615 -921 681 -907
rect 615 -955 631 -921
rect 665 -955 681 -921
rect 615 -989 681 -955
rect 615 -1023 631 -989
rect 665 -1023 681 -989
rect 447 -1077 463 -1057
rect 329 -1091 463 -1077
rect 497 -1077 513 -1057
rect 615 -1057 681 -1023
rect 715 -915 749 -873
rect 715 -983 749 -949
rect 715 -1033 749 -1017
rect 783 -921 849 -907
rect 783 -955 799 -921
rect 833 -955 849 -921
rect 783 -989 849 -955
rect 783 -1023 799 -989
rect 833 -1023 849 -989
rect 615 -1077 631 -1057
rect 497 -1091 631 -1077
rect 665 -1077 681 -1057
rect 783 -1057 849 -1023
rect 883 -915 917 -873
rect 883 -983 917 -949
rect 883 -1033 917 -1017
rect 951 -921 1017 -907
rect 951 -955 967 -921
rect 1001 -955 1017 -921
rect 951 -989 1017 -955
rect 951 -1023 967 -989
rect 1001 -1023 1017 -989
rect 783 -1077 799 -1057
rect 665 -1091 799 -1077
rect 833 -1077 849 -1057
rect 951 -1057 1017 -1023
rect 1051 -915 1085 -873
rect 1051 -983 1085 -949
rect 1051 -1033 1085 -1017
rect 1119 -921 1185 -907
rect 1119 -955 1135 -921
rect 1169 -955 1185 -921
rect 1119 -989 1185 -955
rect 1119 -1023 1135 -989
rect 1169 -1023 1185 -989
rect 951 -1077 967 -1057
rect 833 -1091 967 -1077
rect 1001 -1077 1017 -1057
rect 1119 -1057 1185 -1023
rect 1219 -915 1253 -873
rect 1219 -983 1253 -949
rect 1219 -1033 1253 -1017
rect 1287 -921 1353 -907
rect 1287 -955 1303 -921
rect 1337 -955 1353 -921
rect 1287 -989 1353 -955
rect 1287 -1023 1303 -989
rect 1337 -1023 1353 -989
rect 1119 -1077 1135 -1057
rect 1001 -1091 1135 -1077
rect 1169 -1091 1185 -1057
rect 1287 -1057 1353 -1023
rect 1387 -915 1421 -873
rect 1387 -983 1421 -949
rect 1387 -1033 1421 -1017
rect 1455 -921 1521 -907
rect 1455 -955 1471 -921
rect 1505 -955 1521 -921
rect 1455 -989 1521 -955
rect 1455 -1023 1471 -989
rect 1505 -1023 1521 -989
rect 1287 -1077 1303 -1057
rect -215 -1111 1185 -1091
rect 1219 -1091 1303 -1077
rect 1337 -1077 1353 -1057
rect 1455 -1057 1521 -1023
rect 1555 -915 1589 -873
rect 1555 -983 1589 -949
rect 1555 -1033 1589 -1017
rect 1623 -921 1689 -907
rect 1623 -955 1639 -921
rect 1673 -955 1689 -921
rect 1623 -989 1689 -955
rect 1623 -1023 1639 -989
rect 1673 -1023 1689 -989
rect 1455 -1077 1471 -1057
rect 1337 -1091 1471 -1077
rect 1505 -1077 1521 -1057
rect 1623 -1057 1689 -1023
rect 1623 -1077 1639 -1057
rect 1505 -1091 1639 -1077
rect 1673 -1091 1689 -1057
rect 1219 -1111 1689 -1091
rect 1723 -915 1757 -873
rect 1723 -983 1757 -949
rect 1723 -1051 1757 -1017
rect 1723 -1111 1757 -1085
rect -215 -1142 -139 -1111
rect -215 -1176 -200 -1142
rect -166 -1176 -139 -1142
rect 1219 -1145 1254 -1111
rect -215 -1219 -139 -1176
rect -90 -1151 1254 -1145
rect -90 -1185 -69 -1151
rect -35 -1185 -1 -1151
rect 33 -1185 67 -1151
rect 101 -1185 135 -1151
rect 169 -1185 203 -1151
rect 237 -1185 271 -1151
rect 305 -1185 339 -1151
rect 373 -1185 407 -1151
rect 441 -1185 475 -1151
rect 509 -1185 543 -1151
rect 577 -1185 611 -1151
rect 645 -1185 679 -1151
rect 713 -1185 747 -1151
rect 781 -1185 815 -1151
rect 849 -1185 883 -1151
rect 917 -1185 951 -1151
rect 985 -1185 1019 -1151
rect 1053 -1185 1087 -1151
rect 1121 -1185 1155 -1151
rect 1189 -1185 1254 -1151
rect 1295 -1149 1775 -1145
rect 1295 -1151 1419 -1149
rect 1453 -1151 1775 -1149
rect 1295 -1185 1315 -1151
rect 1349 -1185 1383 -1151
rect 1417 -1183 1419 -1151
rect 1417 -1185 1451 -1183
rect 1485 -1185 1519 -1151
rect 1553 -1185 1587 -1151
rect 1621 -1185 1655 -1151
rect 1689 -1185 1775 -1151
rect 1219 -1219 1254 -1185
rect -215 -1235 1185 -1219
rect -215 -1253 -41 -1235
rect -215 -1327 -160 -1253
rect -57 -1269 -41 -1253
rect -7 -1253 127 -1235
rect -7 -1269 9 -1253
rect -125 -1303 -91 -1287
rect -125 -1383 -91 -1337
rect -57 -1303 9 -1269
rect 111 -1269 127 -1253
rect 161 -1253 295 -1235
rect 161 -1269 177 -1253
rect -57 -1337 -41 -1303
rect -7 -1337 9 -1303
rect -57 -1348 9 -1337
rect 43 -1303 77 -1287
rect 43 -1383 77 -1337
rect 111 -1303 177 -1269
rect 279 -1269 295 -1253
rect 329 -1253 463 -1235
rect 329 -1269 345 -1253
rect 111 -1337 127 -1303
rect 161 -1337 177 -1303
rect 111 -1348 177 -1337
rect 211 -1303 245 -1287
rect 211 -1383 245 -1337
rect 279 -1303 345 -1269
rect 447 -1269 463 -1253
rect 497 -1253 631 -1235
rect 497 -1269 513 -1253
rect 279 -1337 295 -1303
rect 329 -1337 345 -1303
rect 279 -1348 345 -1337
rect 379 -1303 413 -1287
rect 379 -1383 413 -1337
rect 447 -1303 513 -1269
rect 615 -1269 631 -1253
rect 665 -1253 799 -1235
rect 665 -1269 681 -1253
rect 447 -1337 463 -1303
rect 497 -1337 513 -1303
rect 447 -1348 513 -1337
rect 547 -1303 581 -1287
rect 547 -1383 581 -1337
rect 615 -1303 681 -1269
rect 783 -1269 799 -1253
rect 833 -1253 967 -1235
rect 833 -1269 849 -1253
rect 615 -1337 631 -1303
rect 665 -1337 681 -1303
rect 615 -1348 681 -1337
rect 715 -1303 749 -1287
rect 715 -1383 749 -1337
rect 783 -1303 849 -1269
rect 951 -1269 967 -1253
rect 1001 -1253 1135 -1235
rect 1001 -1269 1017 -1253
rect 783 -1337 799 -1303
rect 833 -1337 849 -1303
rect 783 -1348 849 -1337
rect 883 -1303 917 -1287
rect 799 -1349 833 -1348
rect 883 -1383 917 -1337
rect 951 -1303 1017 -1269
rect 1119 -1269 1135 -1253
rect 1169 -1269 1185 -1235
rect 1219 -1235 1689 -1219
rect 1219 -1253 1303 -1235
rect 951 -1337 967 -1303
rect 1001 -1337 1017 -1303
rect 951 -1348 1017 -1337
rect 1051 -1303 1085 -1287
rect 967 -1349 1001 -1348
rect 1051 -1383 1085 -1337
rect 1119 -1303 1185 -1269
rect 1287 -1269 1303 -1253
rect 1337 -1253 1471 -1235
rect 1337 -1269 1353 -1253
rect 1119 -1337 1135 -1303
rect 1169 -1337 1185 -1303
rect 1119 -1348 1185 -1337
rect 1135 -1349 1185 -1348
rect 1219 -1303 1253 -1287
rect 1219 -1383 1253 -1337
rect 1287 -1303 1353 -1269
rect 1455 -1269 1471 -1253
rect 1505 -1253 1639 -1235
rect 1505 -1269 1521 -1253
rect 1287 -1337 1303 -1303
rect 1337 -1337 1353 -1303
rect 1287 -1348 1353 -1337
rect 1387 -1303 1421 -1287
rect 1387 -1383 1421 -1337
rect 1455 -1303 1521 -1269
rect 1623 -1269 1639 -1253
rect 1673 -1269 1689 -1235
rect 1455 -1337 1471 -1303
rect 1505 -1337 1521 -1303
rect 1455 -1348 1521 -1337
rect 1555 -1303 1589 -1287
rect 1555 -1383 1589 -1337
rect 1623 -1303 1689 -1269
rect 1623 -1337 1639 -1303
rect 1673 -1337 1689 -1303
rect 1623 -1348 1689 -1337
rect 1723 -1235 1757 -1219
rect 1723 -1303 1757 -1269
rect 1723 -1383 1757 -1337
rect -232 -1417 -203 -1383
rect -169 -1417 -111 -1383
rect -77 -1417 -19 -1383
rect 15 -1417 73 -1383
rect 107 -1417 165 -1383
rect 199 -1417 257 -1383
rect 291 -1417 349 -1383
rect 383 -1417 441 -1383
rect 475 -1417 533 -1383
rect 567 -1417 625 -1383
rect 659 -1417 717 -1383
rect 751 -1417 809 -1383
rect 843 -1417 901 -1383
rect 935 -1417 993 -1383
rect 1027 -1417 1085 -1383
rect 1119 -1417 1177 -1383
rect 1211 -1417 1269 -1383
rect 1303 -1417 1361 -1383
rect 1395 -1417 1453 -1383
rect 1487 -1417 1545 -1383
rect 1579 -1417 1637 -1383
rect 1671 -1417 1729 -1383
rect 1763 -1417 1792 -1383
rect -128 -1429 1792 -1417
rect -128 -1463 -89 -1429
rect -55 -1430 85 -1429
rect -55 -1463 -5 -1430
rect -128 -1464 -5 -1463
rect 29 -1463 85 -1430
rect 119 -1463 177 -1429
rect 211 -1430 545 -1429
rect 211 -1463 267 -1430
rect 29 -1464 267 -1463
rect 301 -1464 361 -1430
rect 395 -1464 452 -1430
rect 486 -1463 545 -1430
rect 579 -1430 1453 -1429
rect 579 -1463 636 -1430
rect 486 -1464 636 -1463
rect 670 -1464 716 -1430
rect 750 -1464 809 -1430
rect 843 -1464 901 -1430
rect 935 -1464 994 -1430
rect 1028 -1464 1085 -1430
rect 1119 -1464 1177 -1430
rect 1211 -1464 1270 -1430
rect 1304 -1464 1361 -1430
rect 1395 -1463 1453 -1430
rect 1487 -1430 1792 -1429
rect 1487 -1463 1545 -1430
rect 1395 -1464 1545 -1463
rect 1579 -1464 1640 -1430
rect 1674 -1464 1728 -1430
rect 1762 -1464 1792 -1430
rect -128 -1479 1792 -1464
rect -128 -1513 -99 -1479
rect -65 -1513 -7 -1479
rect 27 -1513 85 -1479
rect 119 -1513 177 -1479
rect 211 -1513 269 -1479
rect 303 -1513 361 -1479
rect 395 -1513 453 -1479
rect 487 -1513 545 -1479
rect 579 -1513 637 -1479
rect 671 -1513 717 -1479
rect 751 -1513 809 -1479
rect 843 -1513 901 -1479
rect 935 -1513 993 -1479
rect 1027 -1513 1085 -1479
rect 1119 -1513 1177 -1479
rect 1211 -1513 1269 -1479
rect 1303 -1513 1361 -1479
rect 1395 -1513 1453 -1479
rect 1487 -1513 1545 -1479
rect 1579 -1513 1637 -1479
rect 1671 -1513 1729 -1479
rect 1763 -1513 1792 -1479
rect -93 -1568 -59 -1547
rect -23 -1555 43 -1513
rect -23 -1589 -7 -1555
rect 27 -1589 43 -1555
rect 79 -1585 131 -1547
rect -93 -1623 -59 -1602
rect 113 -1619 131 -1585
rect -93 -1657 40 -1623
rect 79 -1648 131 -1619
rect -107 -1711 -39 -1693
rect -107 -1745 -97 -1711
rect -57 -1745 -39 -1711
rect -107 -1767 -39 -1745
rect 6 -1708 40 -1657
rect 6 -1724 61 -1708
rect 6 -1758 27 -1724
rect 6 -1774 61 -1758
rect 6 -1803 40 -1774
rect -95 -1837 40 -1803
rect 95 -1808 131 -1648
rect 195 -1555 261 -1513
rect 195 -1589 211 -1555
rect 245 -1589 261 -1555
rect 195 -1623 261 -1589
rect 195 -1657 211 -1623
rect 245 -1657 261 -1623
rect 195 -1673 261 -1657
rect 295 -1591 329 -1547
rect 363 -1559 429 -1513
rect 363 -1593 379 -1559
rect 413 -1593 429 -1559
rect 363 -1609 429 -1593
rect 463 -1591 497 -1547
rect 295 -1643 329 -1625
rect 547 -1559 595 -1513
rect 581 -1593 595 -1559
rect 547 -1609 595 -1593
rect 631 -1591 665 -1547
rect 463 -1643 497 -1625
rect 631 -1643 665 -1625
rect 295 -1677 497 -1643
rect 538 -1677 665 -1643
rect 735 -1555 801 -1513
rect 735 -1589 751 -1555
rect 785 -1589 801 -1555
rect 735 -1623 801 -1589
rect 735 -1657 751 -1623
rect 785 -1657 801 -1623
rect 735 -1673 801 -1657
rect 835 -1591 869 -1547
rect 903 -1559 969 -1513
rect 903 -1593 919 -1559
rect 953 -1593 969 -1559
rect 903 -1609 969 -1593
rect 1003 -1591 1037 -1547
rect 835 -1643 869 -1625
rect 1087 -1559 1135 -1513
rect 1121 -1593 1135 -1559
rect 1087 -1609 1135 -1593
rect 1171 -1591 1205 -1547
rect 1003 -1643 1037 -1625
rect 1171 -1643 1205 -1625
rect 835 -1677 1037 -1643
rect 1078 -1677 1205 -1643
rect 1287 -1555 1353 -1513
rect 1287 -1589 1303 -1555
rect 1337 -1589 1353 -1555
rect 1287 -1623 1353 -1589
rect 1287 -1657 1303 -1623
rect 1337 -1657 1353 -1623
rect 1287 -1673 1353 -1657
rect 1387 -1591 1421 -1547
rect 1455 -1559 1521 -1513
rect 1455 -1593 1471 -1559
rect 1505 -1593 1521 -1559
rect 1455 -1609 1521 -1593
rect 1555 -1591 1589 -1547
rect 1387 -1643 1421 -1625
rect 1639 -1559 1687 -1513
rect 1673 -1593 1687 -1559
rect 1639 -1609 1687 -1593
rect 1723 -1591 1757 -1547
rect 1555 -1643 1589 -1625
rect 1723 -1643 1757 -1625
rect 1387 -1677 1589 -1643
rect 1630 -1677 1757 -1643
rect 295 -1714 394 -1677
rect 538 -1711 572 -1677
rect 295 -1748 302 -1714
rect 336 -1748 394 -1714
rect 472 -1745 488 -1711
rect 522 -1745 572 -1711
rect 295 -1785 394 -1748
rect -95 -1871 -59 -1837
rect 77 -1858 131 -1808
rect -95 -1905 -93 -1871
rect -95 -1939 -59 -1905
rect -95 -1973 -93 -1939
rect -95 -1989 -59 -1973
rect -23 -1905 -7 -1871
rect 27 -1905 43 -1871
rect -23 -1939 43 -1905
rect -23 -1973 -7 -1939
rect 27 -1973 43 -1939
rect -23 -2023 43 -1973
rect 77 -1892 79 -1858
rect 113 -1892 131 -1858
rect 77 -1939 131 -1892
rect 77 -1973 79 -1939
rect 113 -1973 131 -1939
rect 77 -1989 131 -1973
rect 195 -1811 261 -1793
rect 195 -1845 211 -1811
rect 245 -1845 261 -1811
rect 195 -1879 261 -1845
rect 195 -1913 211 -1879
rect 245 -1913 261 -1879
rect 195 -1947 261 -1913
rect 195 -1981 211 -1947
rect 245 -1981 261 -1947
rect 195 -2023 261 -1981
rect 295 -1819 497 -1785
rect 295 -1830 329 -1819
rect 463 -1830 497 -1819
rect 538 -1793 572 -1745
rect 606 -1745 622 -1711
rect 656 -1718 682 -1711
rect 606 -1752 632 -1745
rect 666 -1752 682 -1718
rect 606 -1759 682 -1752
rect 835 -1720 934 -1677
rect 1078 -1711 1112 -1677
rect 835 -1754 872 -1720
rect 906 -1754 934 -1720
rect 1012 -1745 1028 -1711
rect 1062 -1745 1112 -1711
rect 835 -1785 934 -1754
rect 538 -1805 681 -1793
rect 538 -1827 631 -1805
rect 295 -1925 329 -1864
rect 295 -1989 329 -1959
rect 363 -1879 429 -1863
rect 363 -1913 379 -1879
rect 413 -1913 429 -1879
rect 363 -1947 429 -1913
rect 363 -1981 379 -1947
rect 413 -1981 429 -1947
rect 363 -2023 429 -1981
rect 615 -1839 631 -1827
rect 665 -1839 681 -1805
rect 463 -1925 497 -1864
rect 463 -1989 497 -1959
rect 533 -1879 581 -1863
rect 533 -1913 547 -1879
rect 533 -1947 581 -1913
rect 533 -1981 547 -1947
rect 533 -2023 581 -1981
rect 615 -1873 681 -1839
rect 615 -1907 631 -1873
rect 665 -1907 681 -1873
rect 615 -1941 681 -1907
rect 615 -1975 631 -1941
rect 665 -1975 681 -1941
rect 615 -1989 681 -1975
rect 735 -1811 801 -1793
rect 735 -1845 751 -1811
rect 785 -1845 801 -1811
rect 735 -1879 801 -1845
rect 735 -1913 751 -1879
rect 785 -1913 801 -1879
rect 735 -1947 801 -1913
rect 735 -1981 751 -1947
rect 785 -1981 801 -1947
rect 735 -2023 801 -1981
rect 835 -1819 1037 -1785
rect 835 -1830 869 -1819
rect 1003 -1830 1037 -1819
rect 1078 -1793 1112 -1745
rect 1146 -1723 1162 -1711
rect 1146 -1757 1160 -1723
rect 1196 -1745 1222 -1711
rect 1194 -1757 1222 -1745
rect 1146 -1759 1222 -1757
rect 1387 -1713 1486 -1677
rect 1630 -1711 1664 -1677
rect 1387 -1747 1425 -1713
rect 1459 -1747 1486 -1713
rect 1564 -1745 1580 -1711
rect 1614 -1745 1664 -1711
rect 1387 -1785 1486 -1747
rect 1078 -1805 1221 -1793
rect 1078 -1827 1171 -1805
rect 835 -1925 869 -1864
rect 835 -1989 869 -1959
rect 903 -1879 969 -1863
rect 903 -1913 919 -1879
rect 953 -1913 969 -1879
rect 903 -1947 969 -1913
rect 903 -1981 919 -1947
rect 953 -1981 969 -1947
rect 903 -2023 969 -1981
rect 1155 -1839 1171 -1827
rect 1205 -1839 1221 -1805
rect 1003 -1925 1037 -1864
rect 1003 -1989 1037 -1959
rect 1073 -1879 1121 -1863
rect 1073 -1913 1087 -1879
rect 1073 -1947 1121 -1913
rect 1073 -1981 1087 -1947
rect 1073 -2023 1121 -1981
rect 1155 -1873 1221 -1839
rect 1155 -1907 1171 -1873
rect 1205 -1907 1221 -1873
rect 1155 -1941 1221 -1907
rect 1155 -1975 1171 -1941
rect 1205 -1975 1221 -1941
rect 1155 -1989 1221 -1975
rect 1287 -1811 1353 -1793
rect 1287 -1845 1303 -1811
rect 1337 -1845 1353 -1811
rect 1287 -1879 1353 -1845
rect 1287 -1913 1303 -1879
rect 1337 -1913 1353 -1879
rect 1287 -1947 1353 -1913
rect 1287 -1981 1303 -1947
rect 1337 -1981 1353 -1947
rect 1287 -2023 1353 -1981
rect 1387 -1819 1589 -1785
rect 1387 -1830 1421 -1819
rect 1555 -1830 1589 -1819
rect 1630 -1793 1664 -1745
rect 1698 -1720 1714 -1711
rect 1698 -1754 1712 -1720
rect 1748 -1745 1774 -1711
rect 1746 -1754 1774 -1745
rect 1698 -1759 1774 -1754
rect 1630 -1805 1773 -1793
rect 1630 -1827 1723 -1805
rect 1387 -1925 1421 -1864
rect 1387 -1989 1421 -1959
rect 1455 -1879 1521 -1863
rect 1455 -1913 1471 -1879
rect 1505 -1913 1521 -1879
rect 1455 -1947 1521 -1913
rect 1455 -1981 1471 -1947
rect 1505 -1981 1521 -1947
rect 1455 -2023 1521 -1981
rect 1707 -1839 1723 -1827
rect 1757 -1839 1773 -1805
rect 1555 -1925 1589 -1864
rect 1555 -1989 1589 -1959
rect 1625 -1879 1673 -1863
rect 1625 -1913 1639 -1879
rect 1625 -1947 1673 -1913
rect 1625 -1981 1639 -1947
rect 1625 -2023 1673 -1981
rect 1707 -1873 1773 -1839
rect 1707 -1907 1723 -1873
rect 1757 -1907 1773 -1873
rect 1707 -1941 1773 -1907
rect 1707 -1975 1723 -1941
rect 1757 -1975 1773 -1941
rect 1707 -1989 1773 -1975
rect -128 -2057 -99 -2023
rect -65 -2057 -7 -2023
rect 27 -2057 85 -2023
rect 119 -2057 177 -2023
rect 211 -2057 269 -2023
rect 303 -2057 361 -2023
rect 395 -2057 453 -2023
rect 487 -2057 545 -2023
rect 579 -2057 637 -2023
rect 671 -2057 717 -2023
rect 751 -2057 809 -2023
rect 843 -2057 901 -2023
rect 935 -2057 993 -2023
rect 1027 -2057 1085 -2023
rect 1119 -2057 1177 -2023
rect 1211 -2057 1269 -2023
rect 1303 -2057 1361 -2023
rect 1395 -2057 1453 -2023
rect 1487 -2057 1545 -2023
rect 1579 -2057 1637 -2023
rect 1671 -2057 1729 -2023
rect 1763 -2057 1792 -2023
rect -128 -2071 1792 -2057
rect -128 -2105 -101 -2071
rect -67 -2072 269 -2071
rect -67 -2105 -5 -2072
rect -128 -2106 -5 -2105
rect 29 -2106 88 -2072
rect 122 -2106 177 -2072
rect 211 -2105 269 -2072
rect 303 -2072 453 -2071
rect 303 -2105 360 -2072
rect 211 -2106 360 -2105
rect 394 -2105 453 -2072
rect 487 -2105 545 -2071
rect 579 -2072 809 -2071
rect 579 -2105 639 -2072
rect 394 -2106 639 -2105
rect 673 -2106 718 -2072
rect 752 -2105 809 -2072
rect 843 -2072 1637 -2071
rect 843 -2105 901 -2072
rect 752 -2106 901 -2105
rect 935 -2106 993 -2072
rect 1027 -2106 1085 -2072
rect 1119 -2106 1176 -2072
rect 1210 -2106 1269 -2072
rect 1303 -2106 1362 -2072
rect 1396 -2106 1454 -2072
rect 1488 -2106 1545 -2072
rect 1579 -2105 1637 -2072
rect 1671 -2105 1724 -2071
rect 1758 -2105 1792 -2071
rect 1579 -2106 1792 -2105
rect -128 -2119 1792 -2106
rect -140 -2153 -111 -2119
rect -77 -2153 -19 -2119
rect 15 -2153 73 -2119
rect 107 -2153 165 -2119
rect 199 -2153 257 -2119
rect 291 -2153 349 -2119
rect 383 -2153 441 -2119
rect 475 -2153 533 -2119
rect 567 -2153 625 -2119
rect 659 -2153 717 -2119
rect 751 -2153 809 -2119
rect 843 -2153 901 -2119
rect 935 -2153 993 -2119
rect 1027 -2153 1085 -2119
rect 1119 -2153 1177 -2119
rect 1211 -2153 1269 -2119
rect 1303 -2153 1361 -2119
rect 1395 -2153 1453 -2119
rect 1487 -2153 1545 -2119
rect 1579 -2153 1637 -2119
rect 1671 -2153 1729 -2119
rect 1763 -2153 1792 -2119
rect -107 -2203 -71 -2187
rect -107 -2237 -105 -2203
rect -107 -2271 -71 -2237
rect -107 -2305 -105 -2271
rect -35 -2203 31 -2153
rect -35 -2237 -19 -2203
rect 15 -2237 31 -2203
rect -35 -2271 31 -2237
rect -35 -2305 -19 -2271
rect 15 -2305 31 -2271
rect 65 -2203 119 -2187
rect 65 -2237 67 -2203
rect 101 -2237 119 -2203
rect 65 -2276 119 -2237
rect 65 -2284 78 -2276
rect -107 -2339 -71 -2305
rect 65 -2318 67 -2284
rect 112 -2310 119 -2276
rect 101 -2318 119 -2310
rect -107 -2373 28 -2339
rect 65 -2368 119 -2318
rect -6 -2402 28 -2373
rect -119 -2431 -51 -2409
rect -119 -2433 -103 -2431
rect -119 -2467 -110 -2433
rect -69 -2465 -51 -2431
rect -76 -2467 -51 -2465
rect -119 -2483 -51 -2467
rect -6 -2418 49 -2402
rect -6 -2452 15 -2418
rect -6 -2468 49 -2452
rect -6 -2519 28 -2468
rect -105 -2553 28 -2519
rect 83 -2528 119 -2368
rect 169 -2203 205 -2187
rect 169 -2237 171 -2203
rect 169 -2271 205 -2237
rect 169 -2305 171 -2271
rect 241 -2203 307 -2153
rect 241 -2237 257 -2203
rect 291 -2237 307 -2203
rect 241 -2271 307 -2237
rect 241 -2305 257 -2271
rect 291 -2305 307 -2271
rect 341 -2203 395 -2187
rect 341 -2237 343 -2203
rect 377 -2237 395 -2203
rect 341 -2273 395 -2237
rect 341 -2284 353 -2273
rect 169 -2339 205 -2305
rect 341 -2318 343 -2284
rect 387 -2307 395 -2273
rect 377 -2318 395 -2307
rect 169 -2373 304 -2339
rect 341 -2368 395 -2318
rect 270 -2402 304 -2373
rect 157 -2431 225 -2409
rect 157 -2433 173 -2431
rect 157 -2467 166 -2433
rect 207 -2465 225 -2431
rect 200 -2467 225 -2465
rect 157 -2483 225 -2467
rect 270 -2418 325 -2402
rect 270 -2452 291 -2418
rect 270 -2468 325 -2452
rect 270 -2519 304 -2468
rect -105 -2574 -71 -2553
rect 67 -2557 119 -2528
rect -105 -2629 -71 -2608
rect -35 -2621 -19 -2587
rect 15 -2621 31 -2587
rect -35 -2663 31 -2621
rect 101 -2591 119 -2557
rect 67 -2629 119 -2591
rect 171 -2553 304 -2519
rect 359 -2528 395 -2368
rect 445 -2203 481 -2187
rect 445 -2237 447 -2203
rect 445 -2271 481 -2237
rect 445 -2305 447 -2271
rect 517 -2203 583 -2153
rect 517 -2237 533 -2203
rect 567 -2237 583 -2203
rect 517 -2271 583 -2237
rect 517 -2305 533 -2271
rect 567 -2305 583 -2271
rect 617 -2203 671 -2187
rect 617 -2237 619 -2203
rect 653 -2237 671 -2203
rect 617 -2273 671 -2237
rect 617 -2284 627 -2273
rect 445 -2339 481 -2305
rect 617 -2318 619 -2284
rect 661 -2307 671 -2273
rect 653 -2318 671 -2307
rect 445 -2373 580 -2339
rect 617 -2368 671 -2318
rect 546 -2402 580 -2373
rect 433 -2431 501 -2409
rect 433 -2433 449 -2431
rect 433 -2467 442 -2433
rect 483 -2465 501 -2431
rect 476 -2467 501 -2465
rect 433 -2483 501 -2467
rect 546 -2418 601 -2402
rect 546 -2452 567 -2418
rect 546 -2468 601 -2452
rect 546 -2519 580 -2468
rect 171 -2574 205 -2553
rect 343 -2557 395 -2528
rect 171 -2629 205 -2608
rect 241 -2621 257 -2587
rect 291 -2621 307 -2587
rect 241 -2663 307 -2621
rect 377 -2591 395 -2557
rect 343 -2629 395 -2591
rect 447 -2553 580 -2519
rect 635 -2528 671 -2368
rect 447 -2574 481 -2553
rect 619 -2557 671 -2528
rect 447 -2629 481 -2608
rect 517 -2621 533 -2587
rect 567 -2621 583 -2587
rect 517 -2663 583 -2621
rect 653 -2591 671 -2557
rect 619 -2629 671 -2591
rect 705 -2203 759 -2187
rect 705 -2237 723 -2203
rect 757 -2237 759 -2203
rect 705 -2284 759 -2237
rect 705 -2318 723 -2284
rect 757 -2318 759 -2284
rect 793 -2203 859 -2153
rect 793 -2237 809 -2203
rect 843 -2237 859 -2203
rect 793 -2271 859 -2237
rect 793 -2305 809 -2271
rect 843 -2305 859 -2271
rect 895 -2203 931 -2187
rect 929 -2237 931 -2203
rect 895 -2271 931 -2237
rect 929 -2305 931 -2271
rect 705 -2368 759 -2318
rect 895 -2339 931 -2305
rect 705 -2528 741 -2368
rect 796 -2373 931 -2339
rect 997 -2203 1033 -2187
rect 997 -2237 999 -2203
rect 997 -2271 1033 -2237
rect 997 -2305 999 -2271
rect 1069 -2203 1135 -2153
rect 1069 -2237 1085 -2203
rect 1119 -2237 1135 -2203
rect 1069 -2271 1135 -2237
rect 1069 -2305 1085 -2271
rect 1119 -2305 1135 -2271
rect 1169 -2203 1223 -2187
rect 1169 -2237 1171 -2203
rect 1205 -2237 1223 -2203
rect 1169 -2270 1223 -2237
rect 1169 -2284 1185 -2270
rect 997 -2339 1033 -2305
rect 1169 -2318 1171 -2284
rect 1219 -2304 1223 -2270
rect 1205 -2318 1223 -2304
rect 997 -2373 1132 -2339
rect 1169 -2368 1223 -2318
rect 796 -2402 830 -2373
rect 775 -2418 830 -2402
rect 1098 -2402 1132 -2373
rect 809 -2452 830 -2418
rect 775 -2468 830 -2452
rect 796 -2519 830 -2468
rect 875 -2431 943 -2409
rect 875 -2465 893 -2431
rect 933 -2465 943 -2431
rect 875 -2483 943 -2465
rect 985 -2431 1053 -2409
rect 985 -2465 994 -2431
rect 1035 -2465 1053 -2431
rect 985 -2483 1053 -2465
rect 1098 -2418 1153 -2402
rect 1098 -2452 1119 -2418
rect 1098 -2468 1153 -2452
rect 1098 -2519 1132 -2468
rect 705 -2557 757 -2528
rect 796 -2553 929 -2519
rect 705 -2591 723 -2557
rect 895 -2574 929 -2553
rect 705 -2629 757 -2591
rect 793 -2621 809 -2587
rect 843 -2621 859 -2587
rect 793 -2663 859 -2621
rect 895 -2629 929 -2608
rect 999 -2553 1132 -2519
rect 1187 -2528 1223 -2368
rect 999 -2574 1033 -2553
rect 1171 -2557 1223 -2528
rect 999 -2629 1033 -2608
rect 1069 -2621 1085 -2587
rect 1119 -2621 1135 -2587
rect 1069 -2663 1135 -2621
rect 1205 -2591 1223 -2557
rect 1171 -2629 1223 -2591
rect 1257 -2203 1311 -2187
rect 1257 -2237 1275 -2203
rect 1309 -2237 1311 -2203
rect 1257 -2284 1311 -2237
rect 1257 -2318 1275 -2284
rect 1309 -2318 1311 -2284
rect 1345 -2203 1411 -2153
rect 1345 -2237 1361 -2203
rect 1395 -2237 1411 -2203
rect 1345 -2271 1411 -2237
rect 1345 -2305 1361 -2271
rect 1395 -2305 1411 -2271
rect 1447 -2203 1483 -2187
rect 1481 -2237 1483 -2203
rect 1447 -2271 1483 -2237
rect 1481 -2305 1483 -2271
rect 1257 -2368 1311 -2318
rect 1447 -2339 1483 -2305
rect 1257 -2528 1293 -2368
rect 1348 -2373 1483 -2339
rect 1549 -2203 1585 -2187
rect 1549 -2237 1551 -2203
rect 1549 -2271 1585 -2237
rect 1549 -2305 1551 -2271
rect 1621 -2203 1687 -2153
rect 1621 -2237 1637 -2203
rect 1671 -2237 1687 -2203
rect 1621 -2271 1687 -2237
rect 1621 -2305 1637 -2271
rect 1671 -2305 1687 -2271
rect 1721 -2203 1775 -2187
rect 1721 -2237 1723 -2203
rect 1757 -2237 1775 -2203
rect 1721 -2272 1775 -2237
rect 1721 -2284 1733 -2272
rect 1549 -2339 1585 -2305
rect 1721 -2318 1723 -2284
rect 1767 -2306 1775 -2272
rect 1757 -2318 1775 -2306
rect 1549 -2373 1684 -2339
rect 1721 -2368 1775 -2318
rect 1348 -2402 1382 -2373
rect 1327 -2418 1382 -2402
rect 1650 -2402 1684 -2373
rect 1361 -2452 1382 -2418
rect 1327 -2468 1382 -2452
rect 1348 -2519 1382 -2468
rect 1427 -2431 1495 -2409
rect 1427 -2465 1445 -2431
rect 1485 -2465 1495 -2431
rect 1427 -2483 1495 -2465
rect 1537 -2431 1605 -2409
rect 1537 -2465 1547 -2431
rect 1587 -2465 1605 -2431
rect 1537 -2483 1605 -2465
rect 1650 -2418 1705 -2402
rect 1650 -2452 1671 -2418
rect 1650 -2468 1705 -2452
rect 1650 -2519 1684 -2468
rect 1257 -2557 1309 -2528
rect 1348 -2553 1481 -2519
rect 1257 -2591 1275 -2557
rect 1447 -2574 1481 -2553
rect 1257 -2629 1309 -2591
rect 1345 -2621 1361 -2587
rect 1395 -2621 1411 -2587
rect 1345 -2663 1411 -2621
rect 1447 -2629 1481 -2608
rect 1551 -2553 1684 -2519
rect 1739 -2528 1775 -2368
rect 1551 -2574 1585 -2553
rect 1723 -2557 1775 -2528
rect 1551 -2629 1585 -2608
rect 1621 -2621 1637 -2587
rect 1671 -2621 1687 -2587
rect 1621 -2663 1687 -2621
rect 1757 -2591 1775 -2557
rect 1723 -2629 1775 -2591
rect -140 -2697 -111 -2663
rect -77 -2697 -19 -2663
rect -140 -2698 -19 -2697
rect -140 -2732 -109 -2698
rect -75 -2731 -19 -2698
rect 15 -2731 73 -2663
rect 107 -2731 165 -2663
rect 199 -2731 257 -2663
rect 291 -2731 349 -2663
rect 383 -2731 441 -2663
rect 475 -2731 533 -2663
rect 567 -2731 625 -2663
rect 659 -2731 717 -2663
rect 751 -2731 809 -2663
rect 843 -2731 901 -2663
rect 935 -2731 993 -2663
rect 1027 -2731 1085 -2663
rect 1119 -2731 1177 -2663
rect 1211 -2697 1269 -2663
rect 1303 -2697 1361 -2663
rect 1211 -2698 1361 -2697
rect 1211 -2731 1269 -2698
rect -75 -2732 1269 -2731
rect 1303 -2731 1361 -2698
rect 1395 -2731 1453 -2663
rect 1487 -2731 1545 -2663
rect 1579 -2731 1637 -2663
rect 1671 -2697 1729 -2663
rect 1763 -2697 1792 -2663
rect 1671 -2731 1717 -2697
rect 1751 -2731 1792 -2697
rect 1303 -2732 1792 -2731
rect -140 -2733 1792 -2732
<< viali >>
rect -203 -873 -169 -839
rect -111 -873 -77 -839
rect -19 -873 15 -839
rect 73 -873 107 -839
rect 165 -873 199 -839
rect 257 -873 291 -839
rect 349 -873 383 -839
rect 441 -873 475 -839
rect 533 -873 567 -839
rect 625 -873 659 -839
rect 717 -873 751 -839
rect 809 -873 843 -839
rect 901 -873 935 -839
rect 993 -873 1027 -839
rect 1085 -873 1119 -839
rect 1177 -873 1211 -839
rect 1269 -873 1303 -839
rect 1361 -873 1395 -839
rect 1453 -873 1487 -839
rect 1545 -873 1579 -839
rect 1637 -873 1671 -839
rect 1729 -873 1763 -839
rect -200 -1176 -166 -1142
rect 1419 -1151 1453 -1149
rect 1419 -1183 1451 -1151
rect 1451 -1183 1453 -1151
rect -203 -1417 -169 -1383
rect -111 -1417 -77 -1383
rect -19 -1417 15 -1383
rect 73 -1417 107 -1383
rect 165 -1417 199 -1383
rect 257 -1417 291 -1383
rect 349 -1417 383 -1383
rect 441 -1417 475 -1383
rect 533 -1417 567 -1383
rect 625 -1417 659 -1383
rect 717 -1417 751 -1383
rect 809 -1417 843 -1383
rect 901 -1417 935 -1383
rect 993 -1417 1027 -1383
rect 1085 -1417 1119 -1383
rect 1177 -1417 1211 -1383
rect 1269 -1417 1303 -1383
rect 1361 -1417 1395 -1383
rect 1453 -1417 1487 -1383
rect 1545 -1417 1579 -1383
rect 1637 -1417 1671 -1383
rect 1729 -1417 1763 -1383
rect -99 -1513 -65 -1479
rect -7 -1513 27 -1479
rect 85 -1513 119 -1479
rect 177 -1513 211 -1479
rect 269 -1513 303 -1479
rect 361 -1513 395 -1479
rect 453 -1513 487 -1479
rect 545 -1513 579 -1479
rect 637 -1513 671 -1479
rect 717 -1513 751 -1479
rect 809 -1513 843 -1479
rect 901 -1513 935 -1479
rect 993 -1513 1027 -1479
rect 1085 -1513 1119 -1479
rect 1177 -1513 1211 -1479
rect 1269 -1513 1303 -1479
rect 1361 -1513 1395 -1479
rect 1453 -1513 1487 -1479
rect 1545 -1513 1579 -1479
rect 1637 -1513 1671 -1479
rect 1729 -1513 1763 -1479
rect -97 -1745 -91 -1711
rect -91 -1745 -63 -1711
rect 302 -1748 336 -1714
rect 632 -1745 656 -1718
rect 656 -1745 666 -1718
rect 632 -1752 666 -1745
rect 872 -1754 906 -1720
rect 1160 -1745 1162 -1723
rect 1162 -1745 1194 -1723
rect 1160 -1757 1194 -1745
rect 1425 -1747 1459 -1713
rect 1712 -1745 1714 -1720
rect 1714 -1745 1746 -1720
rect 1712 -1754 1746 -1745
rect -99 -2057 -65 -2023
rect -7 -2057 27 -2023
rect 85 -2057 119 -2023
rect 177 -2057 211 -2023
rect 269 -2057 303 -2023
rect 361 -2057 395 -2023
rect 453 -2057 487 -2023
rect 545 -2057 579 -2023
rect 637 -2057 671 -2023
rect 717 -2057 751 -2023
rect 809 -2057 843 -2023
rect 901 -2057 935 -2023
rect 993 -2057 1027 -2023
rect 1085 -2057 1119 -2023
rect 1177 -2057 1211 -2023
rect 1269 -2057 1303 -2023
rect 1361 -2057 1395 -2023
rect 1453 -2057 1487 -2023
rect 1545 -2057 1579 -2023
rect 1637 -2057 1671 -2023
rect 1729 -2057 1763 -2023
rect -111 -2153 -77 -2119
rect -19 -2153 15 -2119
rect 73 -2153 107 -2119
rect 165 -2153 199 -2119
rect 257 -2153 291 -2119
rect 349 -2153 383 -2119
rect 441 -2153 475 -2119
rect 533 -2153 567 -2119
rect 625 -2153 659 -2119
rect 717 -2153 751 -2119
rect 809 -2153 843 -2119
rect 901 -2153 935 -2119
rect 993 -2153 1027 -2119
rect 1085 -2153 1119 -2119
rect 1177 -2153 1211 -2119
rect 1269 -2153 1303 -2119
rect 1361 -2153 1395 -2119
rect 1453 -2153 1487 -2119
rect 1545 -2153 1579 -2119
rect 1637 -2153 1671 -2119
rect 1729 -2153 1763 -2119
rect 78 -2284 112 -2276
rect 78 -2310 101 -2284
rect 101 -2310 112 -2284
rect -110 -2465 -103 -2433
rect -103 -2465 -76 -2433
rect -110 -2467 -76 -2465
rect 353 -2284 387 -2273
rect 353 -2307 377 -2284
rect 377 -2307 387 -2284
rect 166 -2465 173 -2433
rect 173 -2465 200 -2433
rect 166 -2467 200 -2465
rect 627 -2284 661 -2273
rect 627 -2307 653 -2284
rect 653 -2307 661 -2284
rect 442 -2465 449 -2433
rect 449 -2465 476 -2433
rect 442 -2467 476 -2465
rect 1185 -2284 1219 -2270
rect 1185 -2304 1205 -2284
rect 1205 -2304 1219 -2284
rect 899 -2465 927 -2431
rect 927 -2465 933 -2431
rect 994 -2465 1001 -2431
rect 1001 -2465 1028 -2431
rect 1733 -2284 1767 -2272
rect 1733 -2306 1757 -2284
rect 1757 -2306 1767 -2284
rect 1451 -2465 1479 -2431
rect 1479 -2465 1485 -2431
rect 1547 -2465 1553 -2431
rect 1553 -2465 1581 -2431
rect -111 -2697 -77 -2663
rect -19 -2697 15 -2663
rect 73 -2697 107 -2663
rect 165 -2697 199 -2663
rect 257 -2697 291 -2663
rect 349 -2697 383 -2663
rect 441 -2697 475 -2663
rect 533 -2697 567 -2663
rect 625 -2697 659 -2663
rect 717 -2697 751 -2663
rect 809 -2697 843 -2663
rect 901 -2697 935 -2663
rect 993 -2697 1027 -2663
rect 1085 -2697 1119 -2663
rect 1177 -2697 1211 -2663
rect 1269 -2697 1303 -2663
rect 1361 -2697 1395 -2663
rect 1453 -2697 1487 -2663
rect 1545 -2697 1579 -2663
rect 1637 -2697 1671 -2663
rect 1729 -2697 1763 -2663
<< metal1 >>
rect -19 -808 15 -805
rect 73 -808 107 -805
rect 165 -808 199 -805
rect 257 -808 291 -805
rect 349 -808 383 -805
rect 441 -808 475 -805
rect 533 -808 567 -805
rect 625 -808 659 -805
rect 717 -808 751 -805
rect 809 -808 843 -805
rect 901 -808 935 -805
rect 993 -808 1027 -805
rect 1085 -808 1119 -805
rect 1177 -808 1211 -805
rect 1269 -808 1303 -805
rect 1361 -808 1395 -805
rect 1453 -808 1487 -805
rect 1545 -808 1579 -805
rect 1637 -808 1671 -805
rect -232 -825 1792 -808
rect -232 -828 1375 -825
rect -232 -829 1175 -828
rect -232 -839 974 -829
rect 1026 -839 1175 -829
rect 1227 -839 1375 -828
rect 1427 -826 1792 -825
rect 1427 -839 1599 -826
rect 1651 -839 1792 -826
rect -232 -873 -203 -839
rect -169 -873 -111 -839
rect -77 -873 -19 -839
rect 15 -873 73 -839
rect 107 -873 165 -839
rect 199 -873 257 -839
rect 291 -873 349 -839
rect 383 -873 441 -839
rect 475 -873 533 -839
rect 567 -873 625 -839
rect 659 -873 717 -839
rect 751 -873 809 -839
rect 843 -873 901 -839
rect 935 -873 974 -839
rect 1027 -873 1085 -839
rect 1119 -873 1175 -839
rect 1227 -873 1269 -839
rect 1303 -873 1361 -839
rect 1427 -873 1453 -839
rect 1487 -873 1545 -839
rect 1579 -873 1599 -839
rect 1671 -873 1729 -839
rect 1763 -873 1792 -839
rect -232 -881 974 -873
rect 1026 -880 1175 -873
rect 1227 -877 1375 -873
rect 1427 -877 1599 -873
rect 1227 -878 1599 -877
rect 1651 -878 1792 -873
rect 1227 -880 1792 -878
rect 1026 -881 1792 -880
rect -232 -904 1792 -881
rect -209 -1133 -157 -1127
rect -209 -1191 -157 -1185
rect 1410 -1140 1462 -1134
rect 1410 -1198 1462 -1192
rect -232 -1383 1792 -1352
rect -232 -1417 -203 -1383
rect -169 -1417 -111 -1383
rect -77 -1417 -19 -1383
rect 15 -1417 73 -1383
rect 107 -1417 165 -1383
rect 199 -1417 257 -1383
rect 291 -1417 349 -1383
rect 383 -1417 441 -1383
rect 475 -1417 533 -1383
rect 567 -1417 625 -1383
rect 659 -1417 717 -1383
rect 751 -1417 809 -1383
rect 843 -1417 901 -1383
rect 935 -1417 993 -1383
rect 1027 -1417 1085 -1383
rect 1119 -1417 1177 -1383
rect 1211 -1417 1269 -1383
rect 1303 -1417 1361 -1383
rect 1395 -1417 1453 -1383
rect 1487 -1417 1545 -1383
rect 1579 -1417 1637 -1383
rect 1671 -1417 1729 -1383
rect 1763 -1417 1792 -1383
rect -232 -1419 1792 -1417
rect -232 -1422 432 -1419
rect -232 -1448 -61 -1422
rect -128 -1474 -61 -1448
rect -9 -1471 432 -1422
rect 484 -1420 1792 -1419
rect 484 -1471 618 -1420
rect -9 -1472 618 -1471
rect 670 -1472 1792 -1420
rect -9 -1474 1792 -1472
rect -128 -1479 1792 -1474
rect -128 -1513 -99 -1479
rect -65 -1513 -7 -1479
rect 27 -1513 85 -1479
rect 119 -1513 177 -1479
rect 211 -1513 269 -1479
rect 303 -1513 361 -1479
rect 395 -1513 453 -1479
rect 487 -1513 545 -1479
rect 579 -1513 637 -1479
rect 671 -1513 717 -1479
rect 751 -1513 809 -1479
rect 843 -1513 901 -1479
rect 935 -1513 993 -1479
rect 1027 -1513 1085 -1479
rect 1119 -1513 1177 -1479
rect 1211 -1513 1269 -1479
rect 1303 -1513 1361 -1479
rect 1395 -1513 1453 -1479
rect 1487 -1513 1545 -1479
rect 1579 -1513 1637 -1479
rect 1671 -1513 1729 -1479
rect 1763 -1513 1792 -1479
rect -128 -1544 1792 -1513
rect -108 -1711 -51 -1544
rect -108 -1745 -97 -1711
rect -63 -1745 -51 -1711
rect -108 -1757 -51 -1745
rect 201 -1705 253 -1699
rect 295 -1709 349 -1706
rect 253 -1714 349 -1709
rect 253 -1748 302 -1714
rect 336 -1748 349 -1714
rect 253 -1752 349 -1748
rect 295 -1755 349 -1752
rect 623 -1709 675 -1703
rect 1416 -1704 1468 -1698
rect 201 -1763 253 -1757
rect 623 -1767 675 -1761
rect 863 -1711 915 -1705
rect 863 -1769 915 -1763
rect 1151 -1714 1203 -1708
rect 1416 -1762 1468 -1756
rect 1703 -1711 1755 -1705
rect 1151 -1772 1203 -1766
rect 1703 -1769 1755 -1763
rect -128 -2023 1792 -1992
rect -128 -2057 -99 -2023
rect -65 -2057 -7 -2023
rect 27 -2057 85 -2023
rect 119 -2057 177 -2023
rect 211 -2057 269 -2023
rect 303 -2057 361 -2023
rect 395 -2057 453 -2023
rect 487 -2057 545 -2023
rect 579 -2057 637 -2023
rect 671 -2057 717 -2023
rect 751 -2057 809 -2023
rect 843 -2057 901 -2023
rect 935 -2057 993 -2023
rect 1027 -2057 1085 -2023
rect 1119 -2057 1177 -2023
rect 1211 -2057 1269 -2023
rect 1303 -2057 1361 -2023
rect 1395 -2057 1453 -2023
rect 1487 -2057 1545 -2023
rect 1579 -2057 1637 -2023
rect 1671 -2057 1729 -2023
rect 1763 -2057 1792 -2023
rect -128 -2061 1792 -2057
rect -128 -2062 1064 -2061
rect -128 -2088 879 -2062
rect -140 -2114 879 -2088
rect 931 -2113 1064 -2062
rect 1116 -2113 1254 -2061
rect 1306 -2062 1792 -2061
rect 1306 -2113 1438 -2062
rect 931 -2114 1438 -2113
rect 1490 -2065 1792 -2062
rect 1490 -2114 1622 -2065
rect -140 -2117 1622 -2114
rect 1674 -2117 1792 -2065
rect -140 -2119 1792 -2117
rect -140 -2153 -111 -2119
rect -77 -2153 -19 -2119
rect 15 -2153 73 -2119
rect 107 -2153 165 -2119
rect 199 -2153 257 -2119
rect 291 -2153 349 -2119
rect 383 -2153 441 -2119
rect 475 -2153 533 -2119
rect 567 -2153 625 -2119
rect 659 -2153 717 -2119
rect 751 -2153 809 -2119
rect 843 -2153 901 -2119
rect 935 -2153 993 -2119
rect 1027 -2153 1085 -2119
rect 1119 -2153 1177 -2119
rect 1211 -2153 1269 -2119
rect 1303 -2153 1361 -2119
rect 1395 -2153 1453 -2119
rect 1487 -2153 1545 -2119
rect 1579 -2153 1637 -2119
rect 1671 -2153 1729 -2119
rect 1763 -2153 1792 -2119
rect -140 -2184 1792 -2153
rect 69 -2267 121 -2261
rect 69 -2325 121 -2319
rect 344 -2264 396 -2258
rect 344 -2322 396 -2316
rect 618 -2264 670 -2258
rect 618 -2322 670 -2316
rect 1176 -2261 1228 -2255
rect 1176 -2319 1228 -2313
rect 1724 -2263 1776 -2257
rect 1724 -2321 1776 -2315
rect -119 -2424 -67 -2418
rect -119 -2482 -67 -2476
rect 157 -2424 209 -2418
rect 157 -2482 209 -2476
rect 433 -2424 485 -2418
rect 433 -2482 485 -2476
rect 887 -2431 944 -2419
rect 887 -2465 899 -2431
rect 933 -2465 944 -2431
rect 887 -2632 944 -2465
rect 985 -2422 1037 -2416
rect 985 -2480 1037 -2474
rect 1439 -2431 1496 -2419
rect 1439 -2465 1451 -2431
rect 1485 -2465 1496 -2431
rect 1439 -2632 1496 -2465
rect 1538 -2422 1590 -2416
rect 1538 -2480 1590 -2474
rect -140 -2654 1792 -2632
rect -140 -2663 11 -2654
rect 63 -2658 1792 -2654
rect 63 -2663 270 -2658
rect 322 -2663 575 -2658
rect 627 -2663 1792 -2658
rect -140 -2697 -111 -2663
rect -77 -2697 -19 -2663
rect 63 -2697 73 -2663
rect 107 -2697 165 -2663
rect 199 -2697 257 -2663
rect 322 -2697 349 -2663
rect 383 -2697 441 -2663
rect 475 -2697 533 -2663
rect 567 -2697 575 -2663
rect 659 -2697 717 -2663
rect 751 -2697 809 -2663
rect 843 -2697 901 -2663
rect 935 -2697 993 -2663
rect 1027 -2697 1085 -2663
rect 1119 -2697 1177 -2663
rect 1211 -2697 1269 -2663
rect 1303 -2697 1361 -2663
rect 1395 -2697 1453 -2663
rect 1487 -2697 1545 -2663
rect 1579 -2697 1637 -2663
rect 1671 -2697 1729 -2663
rect 1763 -2697 1792 -2663
rect -140 -2706 11 -2697
rect 63 -2706 270 -2697
rect -140 -2710 270 -2706
rect 322 -2710 575 -2697
rect 627 -2710 1792 -2697
rect -140 -2728 1792 -2710
rect -19 -2731 15 -2728
rect 73 -2731 107 -2728
rect 165 -2731 199 -2728
rect 257 -2731 291 -2728
rect 349 -2731 383 -2728
rect 441 -2731 475 -2728
rect 533 -2731 567 -2728
rect 625 -2731 659 -2728
rect 717 -2731 751 -2728
rect 809 -2731 843 -2728
rect 901 -2731 935 -2728
rect 993 -2731 1027 -2728
rect 1085 -2731 1119 -2728
rect 1177 -2731 1211 -2728
rect 1269 -2732 1303 -2728
rect 1361 -2731 1395 -2728
rect 1453 -2731 1487 -2728
rect 1545 -2731 1579 -2728
rect 1637 -2731 1671 -2728
rect 1716 -2731 1750 -2728
<< via1 >>
rect 974 -839 1026 -829
rect 1175 -839 1227 -828
rect 1375 -839 1427 -825
rect 1599 -839 1651 -826
rect 974 -873 993 -839
rect 993 -873 1026 -839
rect 1175 -873 1177 -839
rect 1177 -873 1211 -839
rect 1211 -873 1227 -839
rect 1375 -873 1395 -839
rect 1395 -873 1427 -839
rect 1599 -873 1637 -839
rect 1637 -873 1651 -839
rect 974 -881 1026 -873
rect 1175 -880 1227 -873
rect 1375 -877 1427 -873
rect 1599 -878 1651 -873
rect -209 -1142 -157 -1133
rect -209 -1176 -200 -1142
rect -200 -1176 -166 -1142
rect -166 -1176 -157 -1142
rect -209 -1185 -157 -1176
rect 1410 -1149 1462 -1140
rect 1410 -1183 1419 -1149
rect 1419 -1183 1453 -1149
rect 1453 -1183 1462 -1149
rect 1410 -1192 1462 -1183
rect -61 -1474 -9 -1422
rect 432 -1471 484 -1419
rect 618 -1472 670 -1420
rect 201 -1757 253 -1705
rect 623 -1718 675 -1709
rect 623 -1752 632 -1718
rect 632 -1752 666 -1718
rect 666 -1752 675 -1718
rect 623 -1761 675 -1752
rect 863 -1720 915 -1711
rect 863 -1754 872 -1720
rect 872 -1754 906 -1720
rect 906 -1754 915 -1720
rect 863 -1763 915 -1754
rect 1151 -1723 1203 -1714
rect 1151 -1757 1160 -1723
rect 1160 -1757 1194 -1723
rect 1194 -1757 1203 -1723
rect 1151 -1766 1203 -1757
rect 1416 -1713 1468 -1704
rect 1416 -1747 1425 -1713
rect 1425 -1747 1459 -1713
rect 1459 -1747 1468 -1713
rect 1416 -1756 1468 -1747
rect 1703 -1720 1755 -1711
rect 1703 -1754 1712 -1720
rect 1712 -1754 1746 -1720
rect 1746 -1754 1755 -1720
rect 1703 -1763 1755 -1754
rect 879 -2114 931 -2062
rect 1064 -2113 1116 -2061
rect 1254 -2113 1306 -2061
rect 1438 -2114 1490 -2062
rect 1622 -2117 1674 -2065
rect 69 -2276 121 -2267
rect 69 -2310 78 -2276
rect 78 -2310 112 -2276
rect 112 -2310 121 -2276
rect 69 -2319 121 -2310
rect 344 -2273 396 -2264
rect 344 -2307 353 -2273
rect 353 -2307 387 -2273
rect 387 -2307 396 -2273
rect 344 -2316 396 -2307
rect 618 -2273 670 -2264
rect 618 -2307 627 -2273
rect 627 -2307 661 -2273
rect 661 -2307 670 -2273
rect 618 -2316 670 -2307
rect 1176 -2270 1228 -2261
rect 1176 -2304 1185 -2270
rect 1185 -2304 1219 -2270
rect 1219 -2304 1228 -2270
rect 1176 -2313 1228 -2304
rect 1724 -2272 1776 -2263
rect 1724 -2306 1733 -2272
rect 1733 -2306 1767 -2272
rect 1767 -2306 1776 -2272
rect 1724 -2315 1776 -2306
rect -119 -2433 -67 -2424
rect -119 -2467 -110 -2433
rect -110 -2467 -76 -2433
rect -76 -2467 -67 -2433
rect -119 -2476 -67 -2467
rect 157 -2433 209 -2424
rect 157 -2467 166 -2433
rect 166 -2467 200 -2433
rect 200 -2467 209 -2433
rect 157 -2476 209 -2467
rect 433 -2433 485 -2424
rect 433 -2467 442 -2433
rect 442 -2467 476 -2433
rect 476 -2467 485 -2433
rect 433 -2476 485 -2467
rect 985 -2431 1037 -2422
rect 985 -2465 994 -2431
rect 994 -2465 1028 -2431
rect 1028 -2465 1037 -2431
rect 985 -2474 1037 -2465
rect 1538 -2431 1590 -2422
rect 1538 -2465 1547 -2431
rect 1547 -2465 1581 -2431
rect 1581 -2465 1590 -2431
rect 1538 -2474 1590 -2465
rect 11 -2663 63 -2654
rect 270 -2663 322 -2658
rect 575 -2663 627 -2658
rect 11 -2697 15 -2663
rect 15 -2697 63 -2663
rect 270 -2697 291 -2663
rect 291 -2697 322 -2663
rect 575 -2697 625 -2663
rect 625 -2697 627 -2663
rect 11 -2706 63 -2697
rect 270 -2710 322 -2697
rect 575 -2710 627 -2697
<< metal2 >>
rect -204 -1127 -163 -714
rect -209 -1133 -157 -1127
rect -209 -1191 -157 -1185
rect -72 -1476 -63 -1420
rect -7 -1476 2 -1420
rect 74 -2261 115 -714
rect 206 -1699 247 -714
rect 201 -1705 253 -1699
rect 201 -1763 253 -1757
rect 350 -2258 391 -714
rect 421 -1473 430 -1417
rect 486 -1473 495 -1417
rect 607 -1474 616 -1418
rect 672 -1474 681 -1418
rect 623 -1709 675 -1703
rect 869 -1705 910 -714
rect 963 -883 972 -827
rect 1028 -883 1037 -827
rect 1164 -882 1173 -826
rect 1229 -882 1238 -826
rect 1364 -879 1373 -823
rect 1429 -879 1438 -823
rect 1588 -880 1597 -824
rect 1653 -880 1662 -824
rect 1410 -1140 1462 -1134
rect 1462 -1192 1466 -1170
rect 1410 -1198 1466 -1192
rect 1416 -1698 1466 -1198
rect 1416 -1704 1468 -1698
rect 621 -1761 623 -1730
rect 621 -1767 675 -1761
rect 863 -1711 915 -1705
rect 621 -2258 671 -1767
rect 863 -1769 915 -1763
rect 1151 -1714 1203 -1708
rect 1203 -1766 1215 -1735
rect 1416 -1762 1468 -1756
rect 1703 -1711 1755 -1705
rect 1151 -1772 1215 -1766
rect 1755 -1763 1765 -1736
rect 1703 -1769 1765 -1763
rect 868 -2116 877 -2060
rect 933 -2116 942 -2060
rect 1053 -2115 1062 -2059
rect 1118 -2115 1127 -2059
rect 69 -2267 121 -2261
rect 69 -2325 121 -2319
rect 344 -2264 396 -2258
rect 344 -2322 396 -2316
rect 618 -2264 671 -2258
rect 670 -2298 671 -2264
rect 1165 -2255 1215 -1772
rect 1243 -2115 1252 -2059
rect 1308 -2115 1317 -2059
rect 1427 -2116 1436 -2060
rect 1492 -2116 1501 -2060
rect 1611 -2119 1620 -2063
rect 1676 -2119 1685 -2063
rect 1165 -2261 1228 -2255
rect 1165 -2303 1176 -2261
rect 618 -2322 670 -2316
rect 1715 -2257 1765 -1769
rect 1715 -2263 1776 -2257
rect 1715 -2304 1724 -2263
rect 1176 -2319 1228 -2313
rect 1724 -2321 1776 -2315
rect -119 -2424 -67 -2418
rect -119 -2482 -67 -2476
rect 157 -2424 209 -2418
rect 157 -2482 209 -2476
rect 433 -2424 485 -2418
rect 433 -2482 485 -2476
rect 985 -2422 1037 -2416
rect 985 -2480 1037 -2474
rect 1538 -2422 1590 -2416
rect 1538 -2480 1590 -2474
rect -106 -2798 -78 -2482
rect 0 -2708 9 -2652
rect 65 -2708 74 -2652
rect 171 -2798 199 -2482
rect 259 -2712 268 -2656
rect 324 -2712 333 -2656
rect 446 -2793 474 -2482
rect 564 -2712 573 -2656
rect 629 -2712 638 -2656
rect 991 -2788 1019 -2480
rect 1550 -2793 1578 -2480
<< via2 >>
rect -63 -1422 -7 -1420
rect -63 -1474 -61 -1422
rect -61 -1474 -9 -1422
rect -9 -1474 -7 -1422
rect -63 -1476 -7 -1474
rect 430 -1419 486 -1417
rect 430 -1471 432 -1419
rect 432 -1471 484 -1419
rect 484 -1471 486 -1419
rect 430 -1473 486 -1471
rect 616 -1420 672 -1418
rect 616 -1472 618 -1420
rect 618 -1472 670 -1420
rect 670 -1472 672 -1420
rect 616 -1474 672 -1472
rect 972 -829 1028 -827
rect 972 -881 974 -829
rect 974 -881 1026 -829
rect 1026 -881 1028 -829
rect 972 -883 1028 -881
rect 1173 -828 1229 -826
rect 1173 -880 1175 -828
rect 1175 -880 1227 -828
rect 1227 -880 1229 -828
rect 1173 -882 1229 -880
rect 1373 -825 1429 -823
rect 1373 -877 1375 -825
rect 1375 -877 1427 -825
rect 1427 -877 1429 -825
rect 1373 -879 1429 -877
rect 1597 -826 1653 -824
rect 1597 -878 1599 -826
rect 1599 -878 1651 -826
rect 1651 -878 1653 -826
rect 1597 -880 1653 -878
rect 877 -2062 933 -2060
rect 877 -2114 879 -2062
rect 879 -2114 931 -2062
rect 931 -2114 933 -2062
rect 877 -2116 933 -2114
rect 1062 -2061 1118 -2059
rect 1062 -2113 1064 -2061
rect 1064 -2113 1116 -2061
rect 1116 -2113 1118 -2061
rect 1062 -2115 1118 -2113
rect 1252 -2061 1308 -2059
rect 1252 -2113 1254 -2061
rect 1254 -2113 1306 -2061
rect 1306 -2113 1308 -2061
rect 1252 -2115 1308 -2113
rect 1436 -2062 1492 -2060
rect 1436 -2114 1438 -2062
rect 1438 -2114 1490 -2062
rect 1490 -2114 1492 -2062
rect 1436 -2116 1492 -2114
rect 1620 -2065 1676 -2063
rect 1620 -2117 1622 -2065
rect 1622 -2117 1674 -2065
rect 1674 -2117 1676 -2065
rect 1620 -2119 1676 -2117
rect 9 -2654 65 -2652
rect 9 -2706 11 -2654
rect 11 -2706 63 -2654
rect 63 -2706 65 -2654
rect 9 -2708 65 -2706
rect 268 -2658 324 -2656
rect 268 -2710 270 -2658
rect 270 -2710 322 -2658
rect 322 -2710 324 -2658
rect 268 -2712 324 -2710
rect 573 -2658 629 -2656
rect 573 -2710 575 -2658
rect 575 -2710 627 -2658
rect 627 -2710 629 -2658
rect 573 -2712 629 -2710
<< metal3 >>
rect 942 -824 1066 -818
rect 942 -888 968 -824
rect 1032 -888 1066 -824
rect 942 -896 1066 -888
rect 1143 -823 1267 -817
rect 1143 -887 1169 -823
rect 1233 -887 1267 -823
rect 1143 -895 1267 -887
rect 1343 -820 1467 -814
rect 1343 -884 1369 -820
rect 1433 -884 1467 -820
rect 1343 -892 1467 -884
rect 1567 -821 1691 -815
rect 1567 -885 1593 -821
rect 1657 -885 1691 -821
rect 1567 -893 1691 -885
rect -93 -1417 31 -1411
rect -93 -1481 -67 -1417
rect -3 -1481 31 -1417
rect -93 -1489 31 -1481
rect 400 -1414 524 -1408
rect 400 -1478 426 -1414
rect 490 -1478 524 -1414
rect 400 -1486 524 -1478
rect 586 -1415 710 -1409
rect 586 -1479 612 -1415
rect 676 -1479 710 -1415
rect 586 -1487 710 -1479
rect 847 -2057 971 -2051
rect 847 -2121 873 -2057
rect 937 -2121 971 -2057
rect 847 -2129 971 -2121
rect 1032 -2056 1156 -2050
rect 1032 -2120 1058 -2056
rect 1122 -2120 1156 -2056
rect 1032 -2128 1156 -2120
rect 1222 -2056 1346 -2050
rect 1222 -2120 1248 -2056
rect 1312 -2120 1346 -2056
rect 1222 -2128 1346 -2120
rect 1406 -2057 1530 -2051
rect 1406 -2121 1432 -2057
rect 1496 -2121 1530 -2057
rect 1406 -2129 1530 -2121
rect 1590 -2060 1714 -2054
rect 1590 -2124 1616 -2060
rect 1680 -2124 1714 -2060
rect 1590 -2132 1714 -2124
rect -21 -2649 103 -2643
rect -21 -2713 5 -2649
rect 69 -2713 103 -2649
rect -21 -2721 103 -2713
rect 238 -2653 362 -2647
rect 238 -2717 264 -2653
rect 328 -2717 362 -2653
rect 238 -2725 362 -2717
rect 543 -2653 667 -2647
rect 543 -2717 569 -2653
rect 633 -2717 667 -2653
rect 543 -2725 667 -2717
<< via3 >>
rect 968 -827 1032 -824
rect 968 -883 972 -827
rect 972 -883 1028 -827
rect 1028 -883 1032 -827
rect 968 -888 1032 -883
rect 1169 -826 1233 -823
rect 1169 -882 1173 -826
rect 1173 -882 1229 -826
rect 1229 -882 1233 -826
rect 1169 -887 1233 -882
rect 1369 -823 1433 -820
rect 1369 -879 1373 -823
rect 1373 -879 1429 -823
rect 1429 -879 1433 -823
rect 1369 -884 1433 -879
rect 1593 -824 1657 -821
rect 1593 -880 1597 -824
rect 1597 -880 1653 -824
rect 1653 -880 1657 -824
rect 1593 -885 1657 -880
rect -67 -1420 -3 -1417
rect -67 -1476 -63 -1420
rect -63 -1476 -7 -1420
rect -7 -1476 -3 -1420
rect -67 -1481 -3 -1476
rect 426 -1417 490 -1414
rect 426 -1473 430 -1417
rect 430 -1473 486 -1417
rect 486 -1473 490 -1417
rect 426 -1478 490 -1473
rect 612 -1418 676 -1415
rect 612 -1474 616 -1418
rect 616 -1474 672 -1418
rect 672 -1474 676 -1418
rect 612 -1479 676 -1474
rect 873 -2060 937 -2057
rect 873 -2116 877 -2060
rect 877 -2116 933 -2060
rect 933 -2116 937 -2060
rect 873 -2121 937 -2116
rect 1058 -2059 1122 -2056
rect 1058 -2115 1062 -2059
rect 1062 -2115 1118 -2059
rect 1118 -2115 1122 -2059
rect 1058 -2120 1122 -2115
rect 1248 -2059 1312 -2056
rect 1248 -2115 1252 -2059
rect 1252 -2115 1308 -2059
rect 1308 -2115 1312 -2059
rect 1248 -2120 1312 -2115
rect 1432 -2060 1496 -2057
rect 1432 -2116 1436 -2060
rect 1436 -2116 1492 -2060
rect 1492 -2116 1496 -2060
rect 1432 -2121 1496 -2116
rect 1616 -2063 1680 -2060
rect 1616 -2119 1620 -2063
rect 1620 -2119 1676 -2063
rect 1676 -2119 1680 -2063
rect 1616 -2124 1680 -2119
rect 5 -2652 69 -2649
rect 5 -2708 9 -2652
rect 9 -2708 65 -2652
rect 65 -2708 69 -2652
rect 5 -2713 69 -2708
rect 264 -2656 328 -2653
rect 264 -2712 268 -2656
rect 268 -2712 324 -2656
rect 324 -2712 328 -2656
rect 264 -2717 328 -2712
rect 569 -2656 633 -2653
rect 569 -2712 573 -2656
rect 573 -2712 629 -2656
rect 629 -2712 633 -2656
rect 569 -2717 633 -2712
<< metal4 >>
rect -233 -1414 746 -804
rect -233 -1417 426 -1414
rect -233 -1481 -67 -1417
rect -3 -1478 426 -1417
rect 490 -1415 746 -1414
rect 490 -1478 612 -1415
rect -3 -1479 612 -1478
rect 676 -1479 746 -1415
rect -3 -1481 746 -1479
rect -233 -2649 746 -1481
rect -233 -2713 5 -2649
rect 69 -2653 746 -2649
rect 69 -2713 264 -2653
rect -233 -2717 264 -2713
rect 328 -2717 569 -2653
rect 633 -2717 746 -2653
rect -233 -2732 746 -2717
rect 826 -820 1795 -808
rect 826 -823 1369 -820
rect 826 -824 1169 -823
rect 826 -888 968 -824
rect 1032 -887 1169 -824
rect 1233 -884 1369 -823
rect 1433 -821 1795 -820
rect 1433 -884 1593 -821
rect 1233 -885 1593 -884
rect 1657 -885 1795 -821
rect 1233 -887 1795 -885
rect 1032 -888 1795 -887
rect 826 -2056 1795 -888
rect 826 -2057 1058 -2056
rect 826 -2121 873 -2057
rect 937 -2120 1058 -2057
rect 1122 -2120 1248 -2056
rect 1312 -2057 1795 -2056
rect 1312 -2120 1432 -2057
rect 937 -2121 1432 -2120
rect 1496 -2060 1795 -2057
rect 1496 -2121 1616 -2060
rect 826 -2124 1616 -2121
rect 1680 -2124 1795 -2060
rect 826 -2736 1795 -2124
<< labels >>
flabel metal4 1680 -2736 1795 -808 0 FreeSans 320 0 0 0 VDD
port 0 nsew
flabel metal4 -233 -2732 -67 -804 0 FreeSans 320 0 0 0 VSS
port 1 nsew
flabel metal2 1550 -2793 1578 -2474 0 FreeSans 320 0 0 0 sar_val<7>
port 2 nsew
flabel metal2 991 -2788 1019 -2474 0 FreeSans 320 0 0 0 sar_val<6>
port 3 nsew
flabel metal2 446 -2793 474 -2476 0 FreeSans 320 0 0 0 sar_val<5>
port 4 nsew
flabel metal2 171 -2798 199 -2476 0 FreeSans 320 0 0 0 sar_val<4>
port 5 nsew
flabel metal2 -106 -2798 -78 -2476 0 FreeSans 320 0 0 0 sar_val<3>
port 6 nsew
flabel metal2 -204 -1133 -163 -714 0 FreeSans 320 0 0 0 sw<6>
port 7 nsew
flabel metal2 74 -2267 115 -714 0 FreeSans 320 0 0 0 sw<2>
port 8 nsew
flabel metal2 350 -2264 391 -714 0 FreeSans 320 0 0 0 sw<3>
port 9 nsew
flabel metal2 206 -1705 247 -714 0 FreeSans 320 0 0 0 sw<4>
port 10 nsew
flabel metal2 869 -1711 910 -714 0 FreeSans 320 0 0 0 sw<5>
port 11 nsew
flabel metal1 -97 -1513 -63 -1479 0 FreeSans 200 0 0 0 x7.VGND
flabel metal1 -99 -2057 -65 -2023 0 FreeSans 200 0 0 0 x7.VPWR
flabel locali -99 -2057 -65 -2023 0 FreeSans 200 0 0 0 x7.VPWR
flabel locali -97 -1513 -63 -1479 0 FreeSans 200 0 0 0 x7.VGND
flabel locali 83 -1615 117 -1581 0 FreeSans 200 0 0 0 x7.X
flabel locali 83 -1887 117 -1853 0 FreeSans 200 0 0 0 x7.X
flabel locali 83 -1955 117 -1921 0 FreeSans 200 0 0 0 x7.X
flabel locali -99 -1751 -65 -1717 0 FreeSans 200 0 0 0 x7.A
flabel nwell -99 -2057 -65 -2023 0 FreeSans 200 0 0 0 x7.VPB
flabel pwell -97 -1513 -63 -1479 0 FreeSans 200 0 0 0 x7.VNB
rlabel comment -128 -1496 -128 -1496 2 x7.buf_1
rlabel metal1 -128 -1544 148 -1448 5 x7.VGND
rlabel metal1 -128 -2088 148 -1992 5 x7.VPWR
flabel metal1 167 -2697 201 -2663 0 FreeSans 200 0 0 0 x6.VGND
flabel metal1 165 -2153 199 -2119 0 FreeSans 200 0 0 0 x6.VPWR
flabel locali 165 -2153 199 -2119 0 FreeSans 200 0 0 0 x6.VPWR
flabel locali 167 -2697 201 -2663 0 FreeSans 200 0 0 0 x6.VGND
flabel locali 347 -2595 381 -2561 0 FreeSans 200 0 0 0 x6.X
flabel locali 347 -2323 381 -2289 0 FreeSans 200 0 0 0 x6.X
flabel locali 347 -2255 381 -2221 0 FreeSans 200 0 0 0 x6.X
flabel locali 165 -2459 199 -2425 0 FreeSans 200 0 0 0 x6.A
flabel nwell 165 -2153 199 -2119 0 FreeSans 200 0 0 0 x6.VPB
flabel pwell 167 -2697 201 -2663 0 FreeSans 200 0 0 0 x6.VNB
rlabel comment 136 -2680 136 -2680 4 x6.buf_1
rlabel metal1 136 -2728 412 -2632 1 x6.VGND
rlabel metal1 136 -2184 412 -2088 1 x6.VPWR
flabel metal1 -109 -2697 -75 -2663 0 FreeSans 200 0 0 0 x5.VGND
flabel metal1 -111 -2153 -77 -2119 0 FreeSans 200 0 0 0 x5.VPWR
flabel locali -111 -2153 -77 -2119 0 FreeSans 200 0 0 0 x5.VPWR
flabel locali -109 -2697 -75 -2663 0 FreeSans 200 0 0 0 x5.VGND
flabel locali 71 -2595 105 -2561 0 FreeSans 200 0 0 0 x5.X
flabel locali 71 -2323 105 -2289 0 FreeSans 200 0 0 0 x5.X
flabel locali 71 -2255 105 -2221 0 FreeSans 200 0 0 0 x5.X
flabel locali -111 -2459 -77 -2425 0 FreeSans 200 0 0 0 x5.A
flabel nwell -111 -2153 -77 -2119 0 FreeSans 200 0 0 0 x5.VPB
flabel pwell -109 -2697 -75 -2663 0 FreeSans 200 0 0 0 x5.VNB
rlabel comment -140 -2680 -140 -2680 4 x5.buf_1
rlabel metal1 -140 -2728 136 -2632 1 x5.VGND
rlabel metal1 -140 -2184 136 -2088 1 x5.VPWR
flabel metal1 636 -2057 670 -2023 0 FreeSans 200 0 0 0 x2.VPWR
flabel metal1 636 -1513 670 -1479 0 FreeSans 200 0 0 0 x2.VGND
flabel locali 360 -1751 394 -1717 0 FreeSans 200 0 0 0 x2.X
flabel locali 360 -1819 394 -1785 0 FreeSans 200 0 0 0 x2.X
flabel locali 360 -1683 394 -1649 0 FreeSans 200 0 0 0 x2.X
flabel locali 636 -2057 670 -2023 0 FreeSans 200 0 0 0 x2.VPWR
flabel locali 636 -1513 670 -1479 0 FreeSans 200 0 0 0 x2.VGND
flabel locali 636 -1751 670 -1717 0 FreeSans 200 0 0 0 x2.A
flabel nwell 636 -2057 670 -2023 0 FreeSans 200 0 0 0 x2.VPB
flabel pwell 636 -1513 670 -1479 0 FreeSans 200 0 0 0 x2.VNB
rlabel comment 700 -1496 700 -1496 8 x2.buf_4
rlabel metal1 148 -1544 700 -1448 5 x2.VGND
rlabel metal1 148 -2088 700 -1992 5 x2.VPWR
flabel metal1 899 -2697 933 -2663 0 FreeSans 200 0 0 0 x12.VGND
flabel metal1 901 -2153 935 -2119 0 FreeSans 200 0 0 0 x12.VPWR
flabel locali 901 -2153 935 -2119 0 FreeSans 200 0 0 0 x12.VPWR
flabel locali 899 -2697 933 -2663 0 FreeSans 200 0 0 0 x12.VGND
flabel locali 719 -2595 753 -2561 0 FreeSans 200 0 0 0 x12.X
flabel locali 719 -2323 753 -2289 0 FreeSans 200 0 0 0 x12.X
flabel locali 719 -2255 753 -2221 0 FreeSans 200 0 0 0 x12.X
flabel locali 901 -2459 935 -2425 0 FreeSans 200 0 0 0 x12.A
flabel nwell 901 -2153 935 -2119 0 FreeSans 200 0 0 0 x12.VPB
flabel pwell 899 -2697 933 -2663 0 FreeSans 200 0 0 0 x12.VNB
rlabel comment 964 -2680 964 -2680 6 x12.buf_1
rlabel metal1 688 -2728 964 -2632 1 x12.VGND
rlabel metal1 688 -2184 964 -2088 1 x12.VPWR
flabel metal1 443 -2697 477 -2663 0 FreeSans 200 0 0 0 x4.VGND
flabel metal1 441 -2153 475 -2119 0 FreeSans 200 0 0 0 x4.VPWR
flabel locali 441 -2153 475 -2119 0 FreeSans 200 0 0 0 x4.VPWR
flabel locali 443 -2697 477 -2663 0 FreeSans 200 0 0 0 x4.VGND
flabel locali 623 -2595 657 -2561 0 FreeSans 200 0 0 0 x4.X
flabel locali 623 -2323 657 -2289 0 FreeSans 200 0 0 0 x4.X
flabel locali 623 -2255 657 -2221 0 FreeSans 200 0 0 0 x4.X
flabel locali 441 -2459 475 -2425 0 FreeSans 200 0 0 0 x4.A
flabel nwell 441 -2153 475 -2119 0 FreeSans 200 0 0 0 x4.VPB
flabel pwell 443 -2697 477 -2663 0 FreeSans 200 0 0 0 x4.VNB
rlabel comment 412 -2680 412 -2680 4 x4.buf_1
rlabel metal1 412 -2728 688 -2632 1 x4.VGND
rlabel metal1 412 -2184 688 -2088 1 x4.VPWR
flabel metal1 995 -2697 1029 -2663 0 FreeSans 200 0 0 0 x3.VGND
flabel metal1 993 -2153 1027 -2119 0 FreeSans 200 0 0 0 x3.VPWR
flabel locali 993 -2153 1027 -2119 0 FreeSans 200 0 0 0 x3.VPWR
flabel locali 995 -2697 1029 -2663 0 FreeSans 200 0 0 0 x3.VGND
flabel locali 1175 -2595 1209 -2561 0 FreeSans 200 0 0 0 x3.X
flabel locali 1175 -2323 1209 -2289 0 FreeSans 200 0 0 0 x3.X
flabel locali 1175 -2255 1209 -2221 0 FreeSans 200 0 0 0 x3.X
flabel locali 993 -2459 1027 -2425 0 FreeSans 200 0 0 0 x3.A
flabel nwell 993 -2153 1027 -2119 0 FreeSans 200 0 0 0 x3.VPB
flabel pwell 995 -2697 1029 -2663 0 FreeSans 200 0 0 0 x3.VNB
rlabel comment 964 -2680 964 -2680 4 x3.buf_1
rlabel metal1 964 -2728 1240 -2632 1 x3.VGND
rlabel metal1 964 -2184 1240 -2088 1 x3.VPWR
flabel metal1 1176 -2057 1210 -2023 0 FreeSans 200 0 0 0 x1.VPWR
flabel metal1 1176 -1513 1210 -1479 0 FreeSans 200 0 0 0 x1.VGND
flabel locali 900 -1751 934 -1717 0 FreeSans 200 0 0 0 x1.X
flabel locali 900 -1819 934 -1785 0 FreeSans 200 0 0 0 x1.X
flabel locali 900 -1683 934 -1649 0 FreeSans 200 0 0 0 x1.X
flabel locali 1176 -2057 1210 -2023 0 FreeSans 200 0 0 0 x1.VPWR
flabel locali 1176 -1513 1210 -1479 0 FreeSans 200 0 0 0 x1.VGND
flabel locali 1176 -1751 1210 -1717 0 FreeSans 200 0 0 0 x1.A
flabel nwell 1176 -2057 1210 -2023 0 FreeSans 200 0 0 0 x1.VPB
flabel pwell 1176 -1513 1210 -1479 0 FreeSans 200 0 0 0 x1.VNB
rlabel comment 1240 -1496 1240 -1496 8 x1.buf_4
rlabel metal1 688 -1544 1240 -1448 5 x1.VGND
rlabel metal1 688 -2088 1240 -1992 5 x1.VPWR
flabel metal1 1728 -2057 1762 -2023 0 FreeSans 200 0 0 0 x10.VPWR
flabel metal1 1728 -1513 1762 -1479 0 FreeSans 200 0 0 0 x10.VGND
flabel locali 1452 -1751 1486 -1717 0 FreeSans 200 0 0 0 x10.X
flabel locali 1452 -1819 1486 -1785 0 FreeSans 200 0 0 0 x10.X
flabel locali 1452 -1683 1486 -1649 0 FreeSans 200 0 0 0 x10.X
flabel locali 1728 -2057 1762 -2023 0 FreeSans 200 0 0 0 x10.VPWR
flabel locali 1728 -1513 1762 -1479 0 FreeSans 200 0 0 0 x10.VGND
flabel locali 1728 -1751 1762 -1717 0 FreeSans 200 0 0 0 x10.A
flabel nwell 1728 -2057 1762 -2023 0 FreeSans 200 0 0 0 x10.VPB
flabel pwell 1728 -1513 1762 -1479 0 FreeSans 200 0 0 0 x10.VNB
rlabel comment 1792 -1496 1792 -1496 8 x10.buf_4
rlabel metal1 1240 -1544 1792 -1448 5 x10.VGND
rlabel metal1 1240 -2088 1792 -1992 5 x10.VPWR
flabel metal1 1547 -2697 1581 -2663 0 FreeSans 200 0 0 0 x9.VGND
flabel metal1 1545 -2153 1579 -2119 0 FreeSans 200 0 0 0 x9.VPWR
flabel locali 1545 -2153 1579 -2119 0 FreeSans 200 0 0 0 x9.VPWR
flabel locali 1547 -2697 1581 -2663 0 FreeSans 200 0 0 0 x9.VGND
flabel locali 1727 -2595 1761 -2561 0 FreeSans 200 0 0 0 x9.X
flabel locali 1727 -2323 1761 -2289 0 FreeSans 200 0 0 0 x9.X
flabel locali 1727 -2255 1761 -2221 0 FreeSans 200 0 0 0 x9.X
flabel locali 1545 -2459 1579 -2425 0 FreeSans 200 0 0 0 x9.A
flabel nwell 1545 -2153 1579 -2119 0 FreeSans 200 0 0 0 x9.VPB
flabel pwell 1547 -2697 1581 -2663 0 FreeSans 200 0 0 0 x9.VNB
rlabel comment 1516 -2680 1516 -2680 4 x9.buf_1
rlabel metal1 1516 -2728 1792 -2632 1 x9.VGND
rlabel metal1 1516 -2184 1792 -2088 1 x9.VPWR
flabel metal1 1451 -2697 1485 -2663 0 FreeSans 200 0 0 0 x8.VGND
flabel metal1 1453 -2153 1487 -2119 0 FreeSans 200 0 0 0 x8.VPWR
flabel locali 1453 -2153 1487 -2119 0 FreeSans 200 0 0 0 x8.VPWR
flabel locali 1451 -2697 1485 -2663 0 FreeSans 200 0 0 0 x8.VGND
flabel locali 1271 -2595 1305 -2561 0 FreeSans 200 0 0 0 x8.X
flabel locali 1271 -2323 1305 -2289 0 FreeSans 200 0 0 0 x8.X
flabel locali 1271 -2255 1305 -2221 0 FreeSans 200 0 0 0 x8.X
flabel locali 1453 -2459 1487 -2425 0 FreeSans 200 0 0 0 x8.A
flabel nwell 1453 -2153 1487 -2119 0 FreeSans 200 0 0 0 x8.VPB
flabel pwell 1451 -2697 1485 -2663 0 FreeSans 200 0 0 0 x8.VNB
rlabel comment 1516 -2680 1516 -2680 6 x8.buf_1
rlabel metal1 1240 -2728 1516 -2632 1 x8.VGND
rlabel metal1 1240 -2184 1516 -2088 1 x8.VPWR
flabel locali 1360 -1179 1394 -1145 0 FreeSans 200 0 0 0 x11.A
flabel locali 1452 -1179 1486 -1145 0 FreeSans 200 0 0 0 x11.A
flabel locali -203 -1179 -169 -1145 0 FreeSans 200 0 0 0 x11.X
flabel locali -203 -1111 -169 -1077 0 FreeSans 200 0 0 0 x11.X
flabel pwell 1728 -1417 1762 -1383 0 FreeSans 200 0 0 0 x11.VNB
flabel nwell 1728 -873 1762 -839 0 FreeSans 200 0 0 0 x11.VPB
flabel metal1 1728 -1417 1762 -1383 0 FreeSans 200 0 0 0 x11.VGND
flabel metal1 1728 -873 1762 -839 0 FreeSans 200 0 0 0 x11.VPWR
rlabel comment 1792 -1400 1792 -1400 6 x11.buf_16
rlabel metal1 -232 -1448 1792 -1352 1 x11.VGND
rlabel metal1 -232 -904 1792 -808 1 x11.VPWR
<< end >>
