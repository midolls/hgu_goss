magic
tech sky130A
magscale 1 2
timestamp 1697348449
<< error_s >>
rect 1699 1092 1734 1101
rect 1663 1067 1734 1092
rect 1060 1051 1095 1056
rect 1024 1022 1095 1051
rect 1024 583 1094 1022
rect 1024 547 1077 583
rect 1663 530 1733 1067
rect 2395 856 2429 910
rect 2817 892 2852 897
rect 2781 863 2852 892
rect 1663 494 1716 530
rect 2414 477 2429 856
rect 2448 822 2483 856
rect 2448 477 2482 822
rect 2594 754 2652 760
rect 2594 720 2606 754
rect 2594 714 2652 720
rect 2594 560 2652 566
rect 2594 526 2606 560
rect 2594 520 2652 526
rect 2448 443 2463 477
rect 2781 424 2851 863
rect 2963 795 3021 801
rect 2963 761 2975 795
rect 3133 786 3167 801
rect 3555 786 3590 791
rect 2963 755 3021 761
rect 3133 750 3203 786
rect 3519 757 3590 786
rect 3870 764 3905 782
rect 4293 764 4327 782
rect 3870 757 3941 764
rect 3150 716 3221 750
rect 2963 507 3021 513
rect 2963 473 2975 507
rect 2963 467 3021 473
rect 2781 388 2834 424
rect 3150 371 3220 716
rect 3332 648 3390 654
rect 3332 614 3344 648
rect 3332 608 3390 614
rect 3332 454 3390 460
rect 3332 420 3344 454
rect 3332 414 3390 420
rect 3150 335 3203 371
rect 3519 318 3589 757
rect 3871 728 3941 757
rect 3701 689 3759 695
rect 3888 694 3959 728
rect 3701 655 3713 689
rect 3701 649 3759 655
rect 3701 401 3759 407
rect 3701 367 3713 401
rect 3701 361 3759 367
rect 3519 282 3572 318
rect 3888 265 3958 694
rect 4070 626 4128 632
rect 4070 592 4082 626
rect 4070 586 4128 592
rect 4070 348 4128 354
rect 4070 314 4082 348
rect 4070 308 4128 314
rect 3888 229 3941 265
rect 4257 212 4327 764
rect 4439 743 4497 749
rect 4439 709 4451 743
rect 4439 703 4497 709
rect 5789 563 5853 575
rect 6211 563 6275 575
rect 6633 563 6697 575
rect 7055 563 7119 575
rect 7477 563 7541 575
rect 7899 563 7963 575
rect 8321 563 8385 575
rect 8743 563 8807 575
rect 9165 563 9229 575
rect 9587 563 9651 575
rect 10009 563 10073 575
rect 10431 563 10495 575
rect 10853 563 10917 575
rect 11275 563 11339 575
rect 11697 563 11761 575
rect 12119 563 12183 575
rect 12541 563 12605 575
rect 12963 563 13027 575
rect 13385 563 13449 575
rect 13807 563 13871 575
rect 14229 563 14293 575
rect 14651 563 14715 575
rect 15073 563 15137 575
rect 15495 563 15559 575
rect 15917 563 15981 575
rect 16339 563 16403 575
rect 16761 563 16825 575
rect 17183 563 17247 575
rect 17605 563 17669 575
rect 18027 563 18091 575
rect 18449 563 18513 575
rect 18871 563 18935 575
rect 19293 563 19357 575
rect 19715 563 19779 575
rect 20137 563 20201 575
rect 20559 563 20623 575
rect 20981 563 21045 575
rect 21403 563 21467 575
rect 21825 563 21889 575
rect 22247 563 22311 575
rect 22669 563 22733 575
rect 23091 563 23155 575
rect 23513 563 23577 575
rect 23935 563 23999 575
rect 24357 563 24421 575
rect 24779 563 24843 575
rect 25201 563 25265 575
rect 25623 563 25687 575
rect 26045 563 26109 575
rect 26467 563 26531 575
rect 26889 563 26953 575
rect 27311 563 27375 575
rect 27733 563 27797 575
rect 28155 563 28219 575
rect 28577 563 28641 575
rect 28999 563 29063 575
rect 29421 563 29485 575
rect 29843 563 29907 575
rect 30265 563 30329 575
rect 30687 563 30751 575
rect 31109 563 31173 575
rect 31531 563 31595 575
rect 31953 563 32017 575
rect 32375 563 32439 575
rect 32797 563 32861 575
rect 33219 563 33283 575
rect 33641 563 33705 575
rect 34063 563 34127 575
rect 34485 563 34549 575
rect 34907 563 34971 575
rect 35329 563 35393 575
rect 35751 563 35815 575
rect 36173 563 36237 575
rect 36595 563 36659 575
rect 37017 563 37081 575
rect 37439 563 37503 575
rect 37861 563 37925 575
rect 38283 563 38347 575
rect 38705 563 38769 575
rect 39127 563 39191 575
rect 39549 563 39613 575
rect 39971 563 40035 575
rect 40393 563 40457 575
rect 40815 563 40879 575
rect 41237 563 41301 575
rect 41659 563 41723 575
rect 42081 563 42145 575
rect 42503 563 42567 575
rect 42925 563 42989 575
rect 43347 563 43411 575
rect 43769 563 43833 575
rect 44191 563 44255 575
rect 44613 563 44677 575
rect 45035 563 45099 575
rect 45457 563 45521 575
rect 45879 563 45943 575
rect 46301 563 46365 575
rect 46723 563 46787 575
rect 47145 563 47209 575
rect 47567 563 47631 575
rect 47989 563 48053 575
rect 48411 563 48475 575
rect 48833 563 48897 575
rect 49255 563 49319 575
rect 49677 563 49741 575
rect 50099 563 50163 575
rect 50521 563 50585 575
rect 50943 563 51007 575
rect 51365 563 51429 575
rect 51787 563 51851 575
rect 52209 563 52273 575
rect 52631 563 52695 575
rect 53053 563 53117 575
rect 53475 563 53539 575
rect 53897 563 53961 575
rect 54319 563 54383 575
rect 54741 563 54805 575
rect 55163 563 55227 575
rect 55585 563 55649 575
rect 56007 563 56071 575
rect 56429 563 56493 575
rect 56851 563 56915 575
rect 57273 563 57337 575
rect 57695 563 57759 575
rect 58117 563 58181 575
rect 58539 563 58603 575
rect 58961 563 59025 575
rect 59383 563 59447 575
rect 59805 563 59869 575
rect 60227 563 60291 575
rect 60649 563 60713 575
rect 61071 563 61135 575
rect 61493 563 61557 575
rect 61915 563 61979 575
rect 62337 563 62401 575
rect 62759 563 62823 575
rect 63181 563 63245 575
rect 63603 563 63667 575
rect 64025 563 64089 575
rect 64447 563 64511 575
rect 64869 563 64933 575
rect 65291 563 65355 575
rect 65713 563 65777 575
rect 66135 563 66199 575
rect 66557 563 66621 575
rect 66979 563 67043 575
rect 67401 563 67465 575
rect 67823 563 67887 575
rect 68245 563 68309 575
rect 68667 563 68731 575
rect 69089 563 69153 575
rect 69511 563 69575 575
rect 69933 563 69997 575
rect 70355 563 70419 575
rect 70777 563 70841 575
rect 71199 563 71263 575
rect 71621 563 71685 575
rect 72043 563 72107 575
rect 72465 563 72529 575
rect 72887 563 72951 575
rect 73309 563 73373 575
rect 73731 563 73795 575
rect 74153 563 74217 575
rect 74575 563 74639 575
rect 74997 563 75061 575
rect 75419 563 75483 575
rect 75841 563 75905 575
rect 76263 563 76327 575
rect 76685 563 76749 575
rect 77107 563 77171 575
rect 77529 563 77593 575
rect 77951 563 78015 575
rect 78373 563 78437 575
rect 78795 563 78859 575
rect 79217 563 79281 575
rect 79639 563 79703 575
rect 80061 563 80125 575
rect 80483 563 80547 575
rect 80905 563 80969 575
rect 81327 563 81391 575
rect 81749 563 81813 575
rect 82171 563 82235 575
rect 82593 563 82657 575
rect 83015 563 83079 575
rect 83437 563 83501 575
rect 83859 563 83923 575
rect 84281 563 84345 575
rect 84703 563 84767 575
rect 85125 563 85189 575
rect 85547 563 85611 575
rect 85969 563 86033 575
rect 86391 563 86455 575
rect 86813 563 86877 575
rect 87235 563 87299 575
rect 87657 563 87721 575
rect 88079 563 88143 575
rect 88501 563 88565 575
rect 88923 563 88987 575
rect 89345 563 89409 575
rect 89767 563 89831 575
rect 90189 563 90253 575
rect 90611 563 90675 575
rect 91033 563 91097 575
rect 91455 563 91519 575
rect 91877 563 91941 575
rect 92299 563 92363 575
rect 92721 563 92785 575
rect 93143 563 93207 575
rect 93565 563 93629 575
rect 93987 563 94051 575
rect 94409 563 94473 575
rect 94831 563 94895 575
rect 95253 563 95317 575
rect 95675 563 95739 575
rect 96097 563 96161 575
rect 96519 563 96583 575
rect 96941 563 97005 575
rect 97363 563 97427 575
rect 97785 563 97849 575
rect 98207 563 98271 575
rect 98629 563 98693 575
rect 99051 563 99115 575
rect 99473 563 99537 575
rect 99895 563 99959 575
rect 100317 563 100381 575
rect 100739 563 100803 575
rect 101161 563 101225 575
rect 101583 563 101647 575
rect 102005 563 102069 575
rect 102427 563 102491 575
rect 102849 563 102913 575
rect 103271 563 103335 575
rect 103693 563 103757 575
rect 104115 563 104179 575
rect 104537 563 104601 575
rect 104959 563 105023 575
rect 105381 563 105445 575
rect 105803 563 105867 575
rect 106225 563 106289 575
rect 106647 563 106711 575
rect 107069 563 107133 575
rect 107491 563 107555 575
rect 107913 563 107977 575
rect 108335 563 108399 575
rect 108757 563 108821 575
rect 109179 563 109243 575
rect 109601 563 109665 575
rect 110023 563 110087 575
rect 110445 563 110509 575
rect 110867 563 110931 575
rect 111289 563 111353 575
rect 111711 563 111775 575
rect 112133 563 112197 575
rect 112555 563 112619 575
rect 5563 495 5709 563
rect 5853 523 5869 563
rect 4861 489 4919 495
rect 5283 489 5341 495
rect 5563 489 5763 495
rect 4861 455 4873 489
rect 5283 455 5295 489
rect 5563 455 5717 489
rect 4861 449 4919 455
rect 5283 449 5341 455
rect 5563 449 5763 455
rect 4439 295 4497 301
rect 4439 261 4451 295
rect 4439 255 4497 261
rect 4257 176 4310 212
rect 5563 163 5709 449
rect 5789 203 5869 523
rect 5853 164 5869 203
rect 5789 163 5869 164
rect 5985 495 6131 563
rect 6275 523 6291 563
rect 5985 489 6185 495
rect 5985 455 6139 489
rect 5985 449 6185 455
rect 5985 163 6131 449
rect 6211 203 6291 523
rect 6275 164 6291 203
rect 6211 163 6291 164
rect 6407 495 6553 563
rect 6697 523 6713 563
rect 6407 489 6607 495
rect 6407 455 6561 489
rect 6407 449 6607 455
rect 6407 163 6553 449
rect 6633 203 6713 523
rect 6697 164 6713 203
rect 6633 163 6713 164
rect 6829 495 6975 563
rect 7119 523 7135 563
rect 6829 489 7029 495
rect 6829 455 6983 489
rect 6829 449 7029 455
rect 6829 163 6975 449
rect 7055 203 7135 523
rect 7119 164 7135 203
rect 7055 163 7135 164
rect 7251 495 7397 563
rect 7541 523 7557 563
rect 7251 489 7451 495
rect 7251 455 7405 489
rect 7251 449 7451 455
rect 7251 163 7397 449
rect 7477 203 7557 523
rect 7541 164 7557 203
rect 7477 163 7557 164
rect 7673 495 7819 563
rect 7963 523 7979 563
rect 7673 489 7873 495
rect 7673 455 7827 489
rect 7673 449 7873 455
rect 7673 163 7819 449
rect 7899 203 7979 523
rect 7963 164 7979 203
rect 7899 163 7979 164
rect 8095 495 8241 563
rect 8385 523 8401 563
rect 8095 489 8295 495
rect 8095 455 8249 489
rect 8095 449 8295 455
rect 8095 163 8241 449
rect 8321 203 8401 523
rect 8385 164 8401 203
rect 8321 163 8401 164
rect 8517 495 8663 563
rect 8807 523 8823 563
rect 8517 489 8717 495
rect 8517 455 8671 489
rect 8517 449 8717 455
rect 8517 163 8663 449
rect 8743 203 8823 523
rect 8807 164 8823 203
rect 8743 163 8823 164
rect 8939 495 9085 563
rect 9229 523 9245 563
rect 8939 489 9139 495
rect 8939 455 9093 489
rect 8939 449 9139 455
rect 8939 163 9085 449
rect 9165 203 9245 523
rect 9229 164 9245 203
rect 9165 163 9245 164
rect 9361 495 9507 563
rect 9651 523 9667 563
rect 9361 489 9561 495
rect 9361 455 9515 489
rect 9361 449 9561 455
rect 9361 163 9507 449
rect 9587 203 9667 523
rect 9651 164 9667 203
rect 9587 163 9667 164
rect 9783 495 9929 563
rect 10073 523 10089 563
rect 9783 489 9983 495
rect 9783 455 9937 489
rect 9783 449 9983 455
rect 9783 163 9929 449
rect 10009 203 10089 523
rect 10073 164 10089 203
rect 10009 163 10089 164
rect 10205 495 10351 563
rect 10495 523 10511 563
rect 10205 489 10405 495
rect 10205 455 10359 489
rect 10205 449 10405 455
rect 10205 163 10351 449
rect 10431 203 10511 523
rect 10495 164 10511 203
rect 10431 163 10511 164
rect 10627 495 10773 563
rect 10917 523 10933 563
rect 10627 489 10827 495
rect 10627 455 10781 489
rect 10627 449 10827 455
rect 10627 163 10773 449
rect 10853 203 10933 523
rect 10917 164 10933 203
rect 10853 163 10933 164
rect 11049 495 11195 563
rect 11339 523 11355 563
rect 11049 489 11249 495
rect 11049 455 11203 489
rect 11049 449 11249 455
rect 11049 163 11195 449
rect 11275 203 11355 523
rect 11339 164 11355 203
rect 11275 163 11355 164
rect 11471 495 11617 563
rect 11761 523 11777 563
rect 11471 489 11671 495
rect 11471 455 11625 489
rect 11471 449 11671 455
rect 11471 163 11617 449
rect 11697 203 11777 523
rect 11761 164 11777 203
rect 11697 163 11777 164
rect 11893 495 12039 563
rect 12183 523 12199 563
rect 11893 489 12093 495
rect 11893 455 12047 489
rect 11893 449 12093 455
rect 11893 163 12039 449
rect 12119 203 12199 523
rect 12183 164 12199 203
rect 12119 163 12199 164
rect 12315 495 12461 563
rect 12605 523 12621 563
rect 12315 489 12515 495
rect 12315 455 12469 489
rect 12315 449 12515 455
rect 12315 163 12461 449
rect 12541 203 12621 523
rect 12605 164 12621 203
rect 12541 163 12621 164
rect 12737 495 12883 563
rect 13027 523 13043 563
rect 12737 489 12937 495
rect 12737 455 12891 489
rect 12737 449 12937 455
rect 12737 163 12883 449
rect 12963 203 13043 523
rect 13027 164 13043 203
rect 12963 163 13043 164
rect 13159 495 13305 563
rect 13449 523 13465 563
rect 13159 489 13359 495
rect 13159 455 13313 489
rect 13159 449 13359 455
rect 13159 163 13305 449
rect 13385 203 13465 523
rect 13449 164 13465 203
rect 13385 163 13465 164
rect 13581 495 13727 563
rect 13871 523 13887 563
rect 13581 489 13781 495
rect 13581 455 13735 489
rect 13581 449 13781 455
rect 13581 163 13727 449
rect 13807 203 13887 523
rect 13871 164 13887 203
rect 13807 163 13887 164
rect 14003 495 14149 563
rect 14293 523 14309 563
rect 14003 489 14203 495
rect 14003 455 14157 489
rect 14003 449 14203 455
rect 14003 163 14149 449
rect 14229 203 14309 523
rect 14293 164 14309 203
rect 14229 163 14309 164
rect 14425 495 14571 563
rect 14715 523 14731 563
rect 14425 489 14625 495
rect 14425 455 14579 489
rect 14425 449 14625 455
rect 14425 163 14571 449
rect 14651 203 14731 523
rect 14715 164 14731 203
rect 14651 163 14731 164
rect 14847 495 14993 563
rect 15137 523 15153 563
rect 14847 489 15047 495
rect 14847 455 15001 489
rect 14847 449 15047 455
rect 14847 163 14993 449
rect 15073 203 15153 523
rect 15137 164 15153 203
rect 15073 163 15153 164
rect 15269 495 15415 563
rect 15559 523 15575 563
rect 15269 489 15469 495
rect 15269 455 15423 489
rect 15269 449 15469 455
rect 15269 163 15415 449
rect 15495 203 15575 523
rect 15559 164 15575 203
rect 15495 163 15575 164
rect 15691 495 15837 563
rect 15981 523 15997 563
rect 15691 489 15891 495
rect 15691 455 15845 489
rect 15691 449 15891 455
rect 15691 163 15837 449
rect 15917 203 15997 523
rect 15981 164 15997 203
rect 15917 163 15997 164
rect 16113 495 16259 563
rect 16403 523 16419 563
rect 16113 489 16313 495
rect 16113 455 16267 489
rect 16113 449 16313 455
rect 16113 163 16259 449
rect 16339 203 16419 523
rect 16403 164 16419 203
rect 16339 163 16419 164
rect 16535 495 16681 563
rect 16825 523 16841 563
rect 16535 489 16735 495
rect 16535 455 16689 489
rect 16535 449 16735 455
rect 16535 163 16681 449
rect 16761 203 16841 523
rect 16825 164 16841 203
rect 16761 163 16841 164
rect 16957 495 17103 563
rect 17247 523 17263 563
rect 16957 489 17157 495
rect 16957 455 17111 489
rect 16957 449 17157 455
rect 16957 163 17103 449
rect 17183 203 17263 523
rect 17247 164 17263 203
rect 17183 163 17263 164
rect 17379 495 17525 563
rect 17669 523 17685 563
rect 17379 489 17579 495
rect 17379 455 17533 489
rect 17379 449 17579 455
rect 17379 163 17525 449
rect 17605 203 17685 523
rect 17669 164 17685 203
rect 17605 163 17685 164
rect 17801 495 17947 563
rect 18091 523 18107 563
rect 17801 489 18001 495
rect 17801 455 17955 489
rect 17801 449 18001 455
rect 17801 163 17947 449
rect 18027 203 18107 523
rect 18091 164 18107 203
rect 18027 163 18107 164
rect 18223 495 18369 563
rect 18513 523 18529 563
rect 18223 489 18423 495
rect 18223 455 18377 489
rect 18223 449 18423 455
rect 18223 163 18369 449
rect 18449 203 18529 523
rect 18513 164 18529 203
rect 18449 163 18529 164
rect 18645 495 18791 563
rect 18935 523 18951 563
rect 18645 489 18845 495
rect 18645 455 18799 489
rect 18645 449 18845 455
rect 18645 163 18791 449
rect 18871 203 18951 523
rect 18935 164 18951 203
rect 18871 163 18951 164
rect 19067 495 19213 563
rect 19357 523 19373 563
rect 19067 489 19267 495
rect 19067 455 19221 489
rect 19067 449 19267 455
rect 19067 163 19213 449
rect 19293 203 19373 523
rect 19357 164 19373 203
rect 19293 163 19373 164
rect 19489 495 19635 563
rect 19779 523 19795 563
rect 19489 489 19689 495
rect 19489 455 19643 489
rect 19489 449 19689 455
rect 19489 163 19635 449
rect 19715 203 19795 523
rect 19779 164 19795 203
rect 19715 163 19795 164
rect 19911 495 20057 563
rect 20201 523 20217 563
rect 19911 489 20111 495
rect 19911 455 20065 489
rect 19911 449 20111 455
rect 19911 163 20057 449
rect 20137 203 20217 523
rect 20201 164 20217 203
rect 20137 163 20217 164
rect 20333 495 20479 563
rect 20623 523 20639 563
rect 20333 489 20533 495
rect 20333 455 20487 489
rect 20333 449 20533 455
rect 20333 163 20479 449
rect 20559 203 20639 523
rect 20623 164 20639 203
rect 20559 163 20639 164
rect 20755 495 20901 563
rect 21045 523 21061 563
rect 20755 489 20955 495
rect 20755 455 20909 489
rect 20755 449 20955 455
rect 20755 163 20901 449
rect 20981 203 21061 523
rect 21045 164 21061 203
rect 20981 163 21061 164
rect 21177 495 21323 563
rect 21467 523 21483 563
rect 21177 489 21377 495
rect 21177 455 21331 489
rect 21177 449 21377 455
rect 21177 163 21323 449
rect 21403 203 21483 523
rect 21467 164 21483 203
rect 21403 163 21483 164
rect 21599 495 21745 563
rect 21889 523 21905 563
rect 21599 489 21799 495
rect 21599 455 21753 489
rect 21599 449 21799 455
rect 21599 163 21745 449
rect 21825 203 21905 523
rect 21889 164 21905 203
rect 21825 163 21905 164
rect 22021 495 22167 563
rect 22311 523 22327 563
rect 22021 489 22221 495
rect 22021 455 22175 489
rect 22021 449 22221 455
rect 22021 163 22167 449
rect 22247 203 22327 523
rect 22311 164 22327 203
rect 22247 163 22327 164
rect 22443 495 22589 563
rect 22733 523 22749 563
rect 22443 489 22643 495
rect 22443 455 22597 489
rect 22443 449 22643 455
rect 22443 163 22589 449
rect 22669 203 22749 523
rect 22733 164 22749 203
rect 22669 163 22749 164
rect 22865 495 23011 563
rect 23155 523 23171 563
rect 22865 489 23065 495
rect 22865 455 23019 489
rect 22865 449 23065 455
rect 22865 163 23011 449
rect 23091 203 23171 523
rect 23155 164 23171 203
rect 23091 163 23171 164
rect 23287 495 23433 563
rect 23577 523 23593 563
rect 23287 489 23487 495
rect 23287 455 23441 489
rect 23287 449 23487 455
rect 23287 163 23433 449
rect 23513 203 23593 523
rect 23577 164 23593 203
rect 23513 163 23593 164
rect 23709 495 23855 563
rect 23999 523 24015 563
rect 23709 489 23909 495
rect 23709 455 23863 489
rect 23709 449 23909 455
rect 23709 163 23855 449
rect 23935 203 24015 523
rect 23999 164 24015 203
rect 23935 163 24015 164
rect 24131 495 24277 563
rect 24421 523 24437 563
rect 24131 489 24331 495
rect 24131 455 24285 489
rect 24131 449 24331 455
rect 24131 163 24277 449
rect 24357 203 24437 523
rect 24421 164 24437 203
rect 24357 163 24437 164
rect 24553 495 24699 563
rect 24843 523 24859 563
rect 24553 489 24753 495
rect 24553 455 24707 489
rect 24553 449 24753 455
rect 24553 163 24699 449
rect 24779 203 24859 523
rect 24843 164 24859 203
rect 24779 163 24859 164
rect 24975 495 25121 563
rect 25265 523 25281 563
rect 24975 489 25175 495
rect 24975 455 25129 489
rect 24975 449 25175 455
rect 24975 163 25121 449
rect 25201 203 25281 523
rect 25265 164 25281 203
rect 25201 163 25281 164
rect 25397 495 25543 563
rect 25687 523 25703 563
rect 25397 489 25597 495
rect 25397 455 25551 489
rect 25397 449 25597 455
rect 25397 163 25543 449
rect 25623 203 25703 523
rect 25687 164 25703 203
rect 25623 163 25703 164
rect 25819 495 25965 563
rect 26109 523 26125 563
rect 25819 489 26019 495
rect 25819 455 25973 489
rect 25819 449 26019 455
rect 25819 163 25965 449
rect 26045 203 26125 523
rect 26109 164 26125 203
rect 26045 163 26125 164
rect 26241 495 26387 563
rect 26531 523 26547 563
rect 26241 489 26441 495
rect 26241 455 26395 489
rect 26241 449 26441 455
rect 26241 163 26387 449
rect 26467 203 26547 523
rect 26531 164 26547 203
rect 26467 163 26547 164
rect 26663 495 26809 563
rect 26953 523 26969 563
rect 26663 489 26863 495
rect 26663 455 26817 489
rect 26663 449 26863 455
rect 26663 163 26809 449
rect 26889 203 26969 523
rect 26953 164 26969 203
rect 26889 163 26969 164
rect 27085 495 27231 563
rect 27375 523 27391 563
rect 27085 489 27285 495
rect 27085 455 27239 489
rect 27085 449 27285 455
rect 27085 163 27231 449
rect 27311 203 27391 523
rect 27375 164 27391 203
rect 27311 163 27391 164
rect 27507 495 27653 563
rect 27797 523 27813 563
rect 27507 489 27707 495
rect 27507 455 27661 489
rect 27507 449 27707 455
rect 27507 163 27653 449
rect 27733 203 27813 523
rect 27797 164 27813 203
rect 27733 163 27813 164
rect 27929 495 28075 563
rect 28219 523 28235 563
rect 27929 489 28129 495
rect 27929 455 28083 489
rect 27929 449 28129 455
rect 27929 163 28075 449
rect 28155 203 28235 523
rect 28219 164 28235 203
rect 28155 163 28235 164
rect 28351 495 28497 563
rect 28641 523 28657 563
rect 28351 489 28551 495
rect 28351 455 28505 489
rect 28351 449 28551 455
rect 28351 163 28497 449
rect 28577 203 28657 523
rect 28641 164 28657 203
rect 28577 163 28657 164
rect 28773 495 28919 563
rect 29063 523 29079 563
rect 28773 489 28973 495
rect 28773 455 28927 489
rect 28773 449 28973 455
rect 28773 163 28919 449
rect 28999 203 29079 523
rect 29063 164 29079 203
rect 28999 163 29079 164
rect 29195 495 29341 563
rect 29485 523 29501 563
rect 29195 489 29395 495
rect 29195 455 29349 489
rect 29195 449 29395 455
rect 29195 163 29341 449
rect 29421 203 29501 523
rect 29485 164 29501 203
rect 29421 163 29501 164
rect 29617 495 29763 563
rect 29907 523 29923 563
rect 29617 489 29817 495
rect 29617 455 29771 489
rect 29617 449 29817 455
rect 29617 163 29763 449
rect 29843 203 29923 523
rect 29907 164 29923 203
rect 29843 163 29923 164
rect 30039 495 30185 563
rect 30329 523 30345 563
rect 30039 489 30239 495
rect 30039 455 30193 489
rect 30039 449 30239 455
rect 30039 163 30185 449
rect 30265 203 30345 523
rect 30329 164 30345 203
rect 30265 163 30345 164
rect 30461 495 30607 563
rect 30751 523 30767 563
rect 30461 489 30661 495
rect 30461 455 30615 489
rect 30461 449 30661 455
rect 30461 163 30607 449
rect 30687 203 30767 523
rect 30751 164 30767 203
rect 30687 163 30767 164
rect 30883 495 31029 563
rect 31173 523 31189 563
rect 30883 489 31083 495
rect 30883 455 31037 489
rect 30883 449 31083 455
rect 30883 163 31029 449
rect 31109 203 31189 523
rect 31173 164 31189 203
rect 31109 163 31189 164
rect 31305 495 31451 563
rect 31595 523 31611 563
rect 31305 489 31505 495
rect 31305 455 31459 489
rect 31305 449 31505 455
rect 31305 163 31451 449
rect 31531 203 31611 523
rect 31595 164 31611 203
rect 31531 163 31611 164
rect 31727 495 31873 563
rect 32017 523 32033 563
rect 31727 489 31927 495
rect 31727 455 31881 489
rect 31727 449 31927 455
rect 31727 163 31873 449
rect 31953 203 32033 523
rect 32017 164 32033 203
rect 31953 163 32033 164
rect 32149 495 32295 563
rect 32439 523 32455 563
rect 32149 489 32349 495
rect 32149 455 32303 489
rect 32149 449 32349 455
rect 32149 163 32295 449
rect 32375 203 32455 523
rect 32439 164 32455 203
rect 32375 163 32455 164
rect 32571 495 32717 563
rect 32861 523 32877 563
rect 32571 489 32771 495
rect 32571 455 32725 489
rect 32571 449 32771 455
rect 32571 163 32717 449
rect 32797 203 32877 523
rect 32861 164 32877 203
rect 32797 163 32877 164
rect 32993 495 33139 563
rect 33283 523 33299 563
rect 32993 489 33193 495
rect 32993 455 33147 489
rect 32993 449 33193 455
rect 32993 163 33139 449
rect 33219 203 33299 523
rect 33283 164 33299 203
rect 33219 163 33299 164
rect 33415 495 33561 563
rect 33705 523 33721 563
rect 33415 489 33615 495
rect 33415 455 33569 489
rect 33415 449 33615 455
rect 33415 163 33561 449
rect 33641 203 33721 523
rect 33705 164 33721 203
rect 33641 163 33721 164
rect 33837 495 33983 563
rect 34127 523 34143 563
rect 33837 489 34037 495
rect 33837 455 33991 489
rect 33837 449 34037 455
rect 33837 163 33983 449
rect 34063 203 34143 523
rect 34127 164 34143 203
rect 34063 163 34143 164
rect 34259 495 34405 563
rect 34549 523 34565 563
rect 34259 489 34459 495
rect 34259 455 34413 489
rect 34259 449 34459 455
rect 34259 163 34405 449
rect 34485 203 34565 523
rect 34549 164 34565 203
rect 34485 163 34565 164
rect 34681 495 34827 563
rect 34971 523 34987 563
rect 34681 489 34881 495
rect 34681 455 34835 489
rect 34681 449 34881 455
rect 34681 163 34827 449
rect 34907 203 34987 523
rect 34971 164 34987 203
rect 34907 163 34987 164
rect 35103 495 35249 563
rect 35393 523 35409 563
rect 35103 489 35303 495
rect 35103 455 35257 489
rect 35103 449 35303 455
rect 35103 163 35249 449
rect 35329 203 35409 523
rect 35393 164 35409 203
rect 35329 163 35409 164
rect 35525 495 35671 563
rect 35815 523 35831 563
rect 35525 489 35725 495
rect 35525 455 35679 489
rect 35525 449 35725 455
rect 35525 163 35671 449
rect 35751 203 35831 523
rect 35815 164 35831 203
rect 35751 163 35831 164
rect 35947 495 36093 563
rect 36237 523 36253 563
rect 35947 489 36147 495
rect 35947 455 36101 489
rect 35947 449 36147 455
rect 35947 163 36093 449
rect 36173 203 36253 523
rect 36237 164 36253 203
rect 36173 163 36253 164
rect 36369 495 36515 563
rect 36659 523 36675 563
rect 36369 489 36569 495
rect 36369 455 36523 489
rect 36369 449 36569 455
rect 36369 163 36515 449
rect 36595 203 36675 523
rect 36659 164 36675 203
rect 36595 163 36675 164
rect 36791 495 36937 563
rect 37081 523 37097 563
rect 36791 489 36991 495
rect 36791 455 36945 489
rect 36791 449 36991 455
rect 36791 163 36937 449
rect 37017 203 37097 523
rect 37081 164 37097 203
rect 37017 163 37097 164
rect 37213 495 37359 563
rect 37503 523 37519 563
rect 37213 489 37413 495
rect 37213 455 37367 489
rect 37213 449 37413 455
rect 37213 163 37359 449
rect 37439 203 37519 523
rect 37503 164 37519 203
rect 37439 163 37519 164
rect 37635 495 37781 563
rect 37925 523 37941 563
rect 37635 489 37835 495
rect 37635 455 37789 489
rect 37635 449 37835 455
rect 37635 163 37781 449
rect 37861 203 37941 523
rect 37925 164 37941 203
rect 37861 163 37941 164
rect 38057 495 38203 563
rect 38347 523 38363 563
rect 38057 489 38257 495
rect 38057 455 38211 489
rect 38057 449 38257 455
rect 38057 163 38203 449
rect 38283 203 38363 523
rect 38347 164 38363 203
rect 38283 163 38363 164
rect 38479 495 38625 563
rect 38769 523 38785 563
rect 38479 489 38679 495
rect 38479 455 38633 489
rect 38479 449 38679 455
rect 38479 163 38625 449
rect 38705 203 38785 523
rect 38769 164 38785 203
rect 38705 163 38785 164
rect 38901 495 39047 563
rect 39191 523 39207 563
rect 38901 489 39101 495
rect 38901 455 39055 489
rect 38901 449 39101 455
rect 38901 163 39047 449
rect 39127 203 39207 523
rect 39191 164 39207 203
rect 39127 163 39207 164
rect 39323 495 39469 563
rect 39613 523 39629 563
rect 39323 489 39523 495
rect 39323 455 39477 489
rect 39323 449 39523 455
rect 39323 163 39469 449
rect 39549 203 39629 523
rect 39613 164 39629 203
rect 39549 163 39629 164
rect 39745 495 39891 563
rect 40035 523 40051 563
rect 39745 489 39945 495
rect 39745 455 39899 489
rect 39745 449 39945 455
rect 39745 163 39891 449
rect 39971 203 40051 523
rect 40035 164 40051 203
rect 39971 163 40051 164
rect 40167 495 40313 563
rect 40457 523 40473 563
rect 40167 489 40367 495
rect 40167 455 40321 489
rect 40167 449 40367 455
rect 40167 163 40313 449
rect 40393 203 40473 523
rect 40457 164 40473 203
rect 40393 163 40473 164
rect 40589 495 40735 563
rect 40879 523 40895 563
rect 40589 489 40789 495
rect 40589 455 40743 489
rect 40589 449 40789 455
rect 40589 163 40735 449
rect 40815 203 40895 523
rect 40879 164 40895 203
rect 40815 163 40895 164
rect 41011 495 41157 563
rect 41301 523 41317 563
rect 41011 489 41211 495
rect 41011 455 41165 489
rect 41011 449 41211 455
rect 41011 163 41157 449
rect 41237 203 41317 523
rect 41301 164 41317 203
rect 41237 163 41317 164
rect 41433 495 41579 563
rect 41723 523 41739 563
rect 41433 489 41633 495
rect 41433 455 41587 489
rect 41433 449 41633 455
rect 41433 163 41579 449
rect 41659 203 41739 523
rect 41723 164 41739 203
rect 41659 163 41739 164
rect 41855 495 42001 563
rect 42145 523 42161 563
rect 41855 489 42055 495
rect 41855 455 42009 489
rect 41855 449 42055 455
rect 41855 163 42001 449
rect 42081 203 42161 523
rect 42145 164 42161 203
rect 42081 163 42161 164
rect 42277 495 42423 563
rect 42567 523 42583 563
rect 42277 489 42477 495
rect 42277 455 42431 489
rect 42277 449 42477 455
rect 42277 163 42423 449
rect 42503 203 42583 523
rect 42567 164 42583 203
rect 42503 163 42583 164
rect 42699 495 42845 563
rect 42989 523 43005 563
rect 42699 489 42899 495
rect 42699 455 42853 489
rect 42699 449 42899 455
rect 42699 163 42845 449
rect 42925 203 43005 523
rect 42989 164 43005 203
rect 42925 163 43005 164
rect 43121 495 43267 563
rect 43411 523 43427 563
rect 43121 489 43321 495
rect 43121 455 43275 489
rect 43121 449 43321 455
rect 43121 163 43267 449
rect 43347 203 43427 523
rect 43411 164 43427 203
rect 43347 163 43427 164
rect 43543 495 43689 563
rect 43833 523 43849 563
rect 43543 489 43743 495
rect 43543 455 43697 489
rect 43543 449 43743 455
rect 43543 163 43689 449
rect 43769 203 43849 523
rect 43833 164 43849 203
rect 43769 163 43849 164
rect 43965 495 44111 563
rect 44255 523 44271 563
rect 43965 489 44165 495
rect 43965 455 44119 489
rect 43965 449 44165 455
rect 43965 163 44111 449
rect 44191 203 44271 523
rect 44255 164 44271 203
rect 44191 163 44271 164
rect 44387 495 44533 563
rect 44677 523 44693 563
rect 44387 489 44587 495
rect 44387 455 44541 489
rect 44387 449 44587 455
rect 44387 163 44533 449
rect 44613 203 44693 523
rect 44677 164 44693 203
rect 44613 163 44693 164
rect 44809 495 44955 563
rect 45099 523 45115 563
rect 44809 489 45009 495
rect 44809 455 44963 489
rect 44809 449 45009 455
rect 44809 163 44955 449
rect 45035 203 45115 523
rect 45099 164 45115 203
rect 45035 163 45115 164
rect 45231 495 45377 563
rect 45521 523 45537 563
rect 45231 489 45431 495
rect 45231 455 45385 489
rect 45231 449 45431 455
rect 45231 163 45377 449
rect 45457 203 45537 523
rect 45521 164 45537 203
rect 45457 163 45537 164
rect 45653 495 45799 563
rect 45943 523 45959 563
rect 45653 489 45853 495
rect 45653 455 45807 489
rect 45653 449 45853 455
rect 45653 163 45799 449
rect 45879 203 45959 523
rect 45943 164 45959 203
rect 45879 163 45959 164
rect 46075 495 46221 563
rect 46365 523 46381 563
rect 46075 489 46275 495
rect 46075 455 46229 489
rect 46075 449 46275 455
rect 46075 163 46221 449
rect 46301 203 46381 523
rect 46365 164 46381 203
rect 46301 163 46381 164
rect 46497 495 46643 563
rect 46787 523 46803 563
rect 46497 489 46697 495
rect 46497 455 46651 489
rect 46497 449 46697 455
rect 46497 163 46643 449
rect 46723 203 46803 523
rect 46787 164 46803 203
rect 46723 163 46803 164
rect 46919 495 47065 563
rect 47209 523 47225 563
rect 46919 489 47119 495
rect 46919 455 47073 489
rect 46919 449 47119 455
rect 46919 163 47065 449
rect 47145 203 47225 523
rect 47209 164 47225 203
rect 47145 163 47225 164
rect 47341 495 47487 563
rect 47631 523 47647 563
rect 47341 489 47541 495
rect 47341 455 47495 489
rect 47341 449 47541 455
rect 47341 163 47487 449
rect 47567 203 47647 523
rect 47631 164 47647 203
rect 47567 163 47647 164
rect 47763 495 47909 563
rect 48053 523 48069 563
rect 47763 489 47963 495
rect 47763 455 47917 489
rect 47763 449 47963 455
rect 47763 163 47909 449
rect 47989 203 48069 523
rect 48053 164 48069 203
rect 47989 163 48069 164
rect 48185 495 48331 563
rect 48475 523 48491 563
rect 48185 489 48385 495
rect 48185 455 48339 489
rect 48185 449 48385 455
rect 48185 163 48331 449
rect 48411 203 48491 523
rect 48475 164 48491 203
rect 48411 163 48491 164
rect 48607 495 48753 563
rect 48897 523 48913 563
rect 48607 489 48807 495
rect 48607 455 48761 489
rect 48607 449 48807 455
rect 48607 163 48753 449
rect 48833 203 48913 523
rect 48897 164 48913 203
rect 48833 163 48913 164
rect 49029 495 49175 563
rect 49319 523 49335 563
rect 49029 489 49229 495
rect 49029 455 49183 489
rect 49029 449 49229 455
rect 49029 163 49175 449
rect 49255 203 49335 523
rect 49319 164 49335 203
rect 49255 163 49335 164
rect 49451 495 49597 563
rect 49741 523 49757 563
rect 49451 489 49651 495
rect 49451 455 49605 489
rect 49451 449 49651 455
rect 49451 163 49597 449
rect 49677 203 49757 523
rect 49741 164 49757 203
rect 49677 163 49757 164
rect 49873 495 50019 563
rect 50163 523 50179 563
rect 49873 489 50073 495
rect 49873 455 50027 489
rect 49873 449 50073 455
rect 49873 163 50019 449
rect 50099 203 50179 523
rect 50163 164 50179 203
rect 50099 163 50179 164
rect 50295 495 50441 563
rect 50585 523 50601 563
rect 50295 489 50495 495
rect 50295 455 50449 489
rect 50295 449 50495 455
rect 50295 163 50441 449
rect 50521 203 50601 523
rect 50585 164 50601 203
rect 50521 163 50601 164
rect 50717 495 50863 563
rect 51007 523 51023 563
rect 50717 489 50917 495
rect 50717 455 50871 489
rect 50717 449 50917 455
rect 50717 163 50863 449
rect 50943 203 51023 523
rect 51007 164 51023 203
rect 50943 163 51023 164
rect 51139 495 51285 563
rect 51429 523 51445 563
rect 51139 489 51339 495
rect 51139 455 51293 489
rect 51139 449 51339 455
rect 51139 163 51285 449
rect 51365 203 51445 523
rect 51429 164 51445 203
rect 51365 163 51445 164
rect 51561 495 51707 563
rect 51851 523 51867 563
rect 51561 489 51761 495
rect 51561 455 51715 489
rect 51561 449 51761 455
rect 51561 163 51707 449
rect 51787 203 51867 523
rect 51851 164 51867 203
rect 51787 163 51867 164
rect 51983 495 52129 563
rect 52273 523 52289 563
rect 51983 489 52183 495
rect 51983 455 52137 489
rect 51983 449 52183 455
rect 51983 163 52129 449
rect 52209 203 52289 523
rect 52273 164 52289 203
rect 52209 163 52289 164
rect 52405 495 52551 563
rect 52695 523 52711 563
rect 52405 489 52605 495
rect 52405 455 52559 489
rect 52405 449 52605 455
rect 52405 163 52551 449
rect 52631 203 52711 523
rect 52695 164 52711 203
rect 52631 163 52711 164
rect 52827 495 52973 563
rect 53117 523 53133 563
rect 52827 489 53027 495
rect 52827 455 52981 489
rect 52827 449 53027 455
rect 52827 163 52973 449
rect 53053 203 53133 523
rect 53117 164 53133 203
rect 53053 163 53133 164
rect 53249 495 53395 563
rect 53539 523 53555 563
rect 53249 489 53449 495
rect 53249 455 53403 489
rect 53249 449 53449 455
rect 53249 163 53395 449
rect 53475 203 53555 523
rect 53539 164 53555 203
rect 53475 163 53555 164
rect 53671 495 53817 563
rect 53961 523 53977 563
rect 53671 489 53871 495
rect 53671 455 53825 489
rect 53671 449 53871 455
rect 53671 163 53817 449
rect 53897 203 53977 523
rect 53961 164 53977 203
rect 53897 163 53977 164
rect 54093 495 54239 563
rect 54383 523 54399 563
rect 54093 489 54293 495
rect 54093 455 54247 489
rect 54093 449 54293 455
rect 54093 163 54239 449
rect 54319 203 54399 523
rect 54383 164 54399 203
rect 54319 163 54399 164
rect 54515 495 54661 563
rect 54805 523 54821 563
rect 54515 489 54715 495
rect 54515 455 54669 489
rect 54515 449 54715 455
rect 54515 163 54661 449
rect 54741 203 54821 523
rect 54805 164 54821 203
rect 54741 163 54821 164
rect 54937 495 55083 563
rect 55227 523 55243 563
rect 54937 489 55137 495
rect 54937 455 55091 489
rect 54937 449 55137 455
rect 54937 163 55083 449
rect 55163 203 55243 523
rect 55227 164 55243 203
rect 55163 163 55243 164
rect 55359 495 55505 563
rect 55649 523 55665 563
rect 55359 489 55559 495
rect 55359 455 55513 489
rect 55359 449 55559 455
rect 55359 163 55505 449
rect 55585 203 55665 523
rect 55649 164 55665 203
rect 55585 163 55665 164
rect 55781 495 55927 563
rect 56071 523 56087 563
rect 55781 489 55981 495
rect 55781 455 55935 489
rect 55781 449 55981 455
rect 55781 163 55927 449
rect 56007 203 56087 523
rect 56071 164 56087 203
rect 56007 163 56087 164
rect 56203 495 56349 563
rect 56493 523 56509 563
rect 56203 489 56403 495
rect 56203 455 56357 489
rect 56203 449 56403 455
rect 56203 163 56349 449
rect 56429 203 56509 523
rect 56493 164 56509 203
rect 56429 163 56509 164
rect 56625 495 56771 563
rect 56915 523 56931 563
rect 56625 489 56825 495
rect 56625 455 56779 489
rect 56625 449 56825 455
rect 56625 163 56771 449
rect 56851 203 56931 523
rect 56915 164 56931 203
rect 56851 163 56931 164
rect 57047 495 57193 563
rect 57337 523 57353 563
rect 57047 489 57247 495
rect 57047 455 57201 489
rect 57047 449 57247 455
rect 57047 163 57193 449
rect 57273 203 57353 523
rect 57337 164 57353 203
rect 57273 163 57353 164
rect 57469 495 57615 563
rect 57759 523 57775 563
rect 57469 489 57669 495
rect 57469 455 57623 489
rect 57469 449 57669 455
rect 57469 163 57615 449
rect 57695 203 57775 523
rect 57759 164 57775 203
rect 57695 163 57775 164
rect 57891 495 58037 563
rect 58181 523 58197 563
rect 57891 489 58091 495
rect 57891 455 58045 489
rect 57891 449 58091 455
rect 57891 163 58037 449
rect 58117 203 58197 523
rect 58181 164 58197 203
rect 58117 163 58197 164
rect 58313 495 58459 563
rect 58603 523 58619 563
rect 58313 489 58513 495
rect 58313 455 58467 489
rect 58313 449 58513 455
rect 58313 163 58459 449
rect 58539 203 58619 523
rect 58603 164 58619 203
rect 58539 163 58619 164
rect 58735 495 58881 563
rect 59025 523 59041 563
rect 58735 489 58935 495
rect 58735 455 58889 489
rect 58735 449 58935 455
rect 58735 163 58881 449
rect 58961 203 59041 523
rect 59025 164 59041 203
rect 58961 163 59041 164
rect 59157 495 59303 563
rect 59447 523 59463 563
rect 59157 489 59357 495
rect 59157 455 59311 489
rect 59157 449 59357 455
rect 59157 163 59303 449
rect 59383 203 59463 523
rect 59447 164 59463 203
rect 59383 163 59463 164
rect 59579 495 59725 563
rect 59869 523 59885 563
rect 59579 489 59779 495
rect 59579 455 59733 489
rect 59579 449 59779 455
rect 59579 163 59725 449
rect 59805 203 59885 523
rect 59869 164 59885 203
rect 59805 163 59885 164
rect 60001 495 60147 563
rect 60291 523 60307 563
rect 60001 489 60201 495
rect 60001 455 60155 489
rect 60001 449 60201 455
rect 60001 163 60147 449
rect 60227 203 60307 523
rect 60291 164 60307 203
rect 60227 163 60307 164
rect 60423 495 60569 563
rect 60713 523 60729 563
rect 60423 489 60623 495
rect 60423 455 60577 489
rect 60423 449 60623 455
rect 60423 163 60569 449
rect 60649 203 60729 523
rect 60713 164 60729 203
rect 60649 163 60729 164
rect 60845 495 60991 563
rect 61135 523 61151 563
rect 60845 489 61045 495
rect 60845 455 60999 489
rect 60845 449 61045 455
rect 60845 163 60991 449
rect 61071 203 61151 523
rect 61135 164 61151 203
rect 61071 163 61151 164
rect 61267 495 61413 563
rect 61557 523 61573 563
rect 61267 489 61467 495
rect 61267 455 61421 489
rect 61267 449 61467 455
rect 61267 163 61413 449
rect 61493 203 61573 523
rect 61557 164 61573 203
rect 61493 163 61573 164
rect 61689 495 61835 563
rect 61979 523 61995 563
rect 61689 489 61889 495
rect 61689 455 61843 489
rect 61689 449 61889 455
rect 61689 163 61835 449
rect 61915 203 61995 523
rect 61979 164 61995 203
rect 61915 163 61995 164
rect 62111 495 62257 563
rect 62401 523 62417 563
rect 62111 489 62311 495
rect 62111 455 62265 489
rect 62111 449 62311 455
rect 62111 163 62257 449
rect 62337 203 62417 523
rect 62401 164 62417 203
rect 62337 163 62417 164
rect 62533 495 62679 563
rect 62823 523 62839 563
rect 62533 489 62733 495
rect 62533 455 62687 489
rect 62533 449 62733 455
rect 62533 163 62679 449
rect 62759 203 62839 523
rect 62823 164 62839 203
rect 62759 163 62839 164
rect 62955 495 63101 563
rect 63245 523 63261 563
rect 62955 489 63155 495
rect 62955 455 63109 489
rect 62955 449 63155 455
rect 62955 163 63101 449
rect 63181 203 63261 523
rect 63245 164 63261 203
rect 63181 163 63261 164
rect 63377 495 63523 563
rect 63667 523 63683 563
rect 63377 489 63577 495
rect 63377 455 63531 489
rect 63377 449 63577 455
rect 63377 163 63523 449
rect 63603 203 63683 523
rect 63667 164 63683 203
rect 63603 163 63683 164
rect 63799 495 63945 563
rect 64089 523 64105 563
rect 63799 489 63999 495
rect 63799 455 63953 489
rect 63799 449 63999 455
rect 63799 163 63945 449
rect 64025 203 64105 523
rect 64089 164 64105 203
rect 64025 163 64105 164
rect 64221 495 64367 563
rect 64511 523 64527 563
rect 64221 489 64421 495
rect 64221 455 64375 489
rect 64221 449 64421 455
rect 64221 163 64367 449
rect 64447 203 64527 523
rect 64511 164 64527 203
rect 64447 163 64527 164
rect 64643 495 64789 563
rect 64933 523 64949 563
rect 64643 489 64843 495
rect 64643 455 64797 489
rect 64643 449 64843 455
rect 64643 163 64789 449
rect 64869 203 64949 523
rect 64933 164 64949 203
rect 64869 163 64949 164
rect 65065 495 65211 563
rect 65355 523 65371 563
rect 65065 489 65265 495
rect 65065 455 65219 489
rect 65065 449 65265 455
rect 65065 163 65211 449
rect 65291 203 65371 523
rect 65355 164 65371 203
rect 65291 163 65371 164
rect 65487 495 65633 563
rect 65777 523 65793 563
rect 65487 489 65687 495
rect 65487 455 65641 489
rect 65487 449 65687 455
rect 65487 163 65633 449
rect 65713 203 65793 523
rect 65777 164 65793 203
rect 65713 163 65793 164
rect 65909 495 66055 563
rect 66199 523 66215 563
rect 65909 489 66109 495
rect 65909 455 66063 489
rect 65909 449 66109 455
rect 65909 163 66055 449
rect 66135 203 66215 523
rect 66199 164 66215 203
rect 66135 163 66215 164
rect 66331 495 66477 563
rect 66621 523 66637 563
rect 66331 489 66531 495
rect 66331 455 66485 489
rect 66331 449 66531 455
rect 66331 163 66477 449
rect 66557 203 66637 523
rect 66621 164 66637 203
rect 66557 163 66637 164
rect 66753 495 66899 563
rect 67043 523 67059 563
rect 66753 489 66953 495
rect 66753 455 66907 489
rect 66753 449 66953 455
rect 66753 163 66899 449
rect 66979 203 67059 523
rect 67043 164 67059 203
rect 66979 163 67059 164
rect 67175 495 67321 563
rect 67465 523 67481 563
rect 67175 489 67375 495
rect 67175 455 67329 489
rect 67175 449 67375 455
rect 67175 163 67321 449
rect 67401 203 67481 523
rect 67465 164 67481 203
rect 67401 163 67481 164
rect 67597 495 67743 563
rect 67887 523 67903 563
rect 67597 489 67797 495
rect 67597 455 67751 489
rect 67597 449 67797 455
rect 67597 163 67743 449
rect 67823 203 67903 523
rect 67887 164 67903 203
rect 67823 163 67903 164
rect 68019 495 68165 563
rect 68309 523 68325 563
rect 68019 489 68219 495
rect 68019 455 68173 489
rect 68019 449 68219 455
rect 68019 163 68165 449
rect 68245 203 68325 523
rect 68309 164 68325 203
rect 68245 163 68325 164
rect 68441 495 68587 563
rect 68731 523 68747 563
rect 68441 489 68641 495
rect 68441 455 68595 489
rect 68441 449 68641 455
rect 68441 163 68587 449
rect 68667 203 68747 523
rect 68731 164 68747 203
rect 68667 163 68747 164
rect 68863 495 69009 563
rect 69153 523 69169 563
rect 68863 489 69063 495
rect 68863 455 69017 489
rect 68863 449 69063 455
rect 68863 163 69009 449
rect 69089 203 69169 523
rect 69153 164 69169 203
rect 69089 163 69169 164
rect 69285 495 69431 563
rect 69575 523 69591 563
rect 69285 489 69485 495
rect 69285 455 69439 489
rect 69285 449 69485 455
rect 69285 163 69431 449
rect 69511 203 69591 523
rect 69575 164 69591 203
rect 69511 163 69591 164
rect 69707 495 69853 563
rect 69997 523 70013 563
rect 69707 489 69907 495
rect 69707 455 69861 489
rect 69707 449 69907 455
rect 69707 163 69853 449
rect 69933 203 70013 523
rect 69997 164 70013 203
rect 69933 163 70013 164
rect 70129 495 70275 563
rect 70419 523 70435 563
rect 70129 489 70329 495
rect 70129 455 70283 489
rect 70129 449 70329 455
rect 70129 163 70275 449
rect 70355 203 70435 523
rect 70419 164 70435 203
rect 70355 163 70435 164
rect 70551 495 70697 563
rect 70841 523 70857 563
rect 70551 489 70751 495
rect 70551 455 70705 489
rect 70551 449 70751 455
rect 70551 163 70697 449
rect 70777 203 70857 523
rect 70841 164 70857 203
rect 70777 163 70857 164
rect 70973 495 71119 563
rect 71263 523 71279 563
rect 70973 489 71173 495
rect 70973 455 71127 489
rect 70973 449 71173 455
rect 70973 163 71119 449
rect 71199 203 71279 523
rect 71263 164 71279 203
rect 71199 163 71279 164
rect 71395 495 71541 563
rect 71685 523 71701 563
rect 71395 489 71595 495
rect 71395 455 71549 489
rect 71395 449 71595 455
rect 71395 163 71541 449
rect 71621 203 71701 523
rect 71685 164 71701 203
rect 71621 163 71701 164
rect 71817 495 71963 563
rect 72107 523 72123 563
rect 71817 489 72017 495
rect 71817 455 71971 489
rect 71817 449 72017 455
rect 71817 163 71963 449
rect 72043 203 72123 523
rect 72107 164 72123 203
rect 72043 163 72123 164
rect 72239 495 72385 563
rect 72529 523 72545 563
rect 72239 489 72439 495
rect 72239 455 72393 489
rect 72239 449 72439 455
rect 72239 163 72385 449
rect 72465 203 72545 523
rect 72529 164 72545 203
rect 72465 163 72545 164
rect 72661 495 72807 563
rect 72951 523 72967 563
rect 72661 489 72861 495
rect 72661 455 72815 489
rect 72661 449 72861 455
rect 72661 163 72807 449
rect 72887 203 72967 523
rect 72951 164 72967 203
rect 72887 163 72967 164
rect 73083 495 73229 563
rect 73373 523 73389 563
rect 73083 489 73283 495
rect 73083 455 73237 489
rect 73083 449 73283 455
rect 73083 163 73229 449
rect 73309 203 73389 523
rect 73373 164 73389 203
rect 73309 163 73389 164
rect 73505 495 73651 563
rect 73795 523 73811 563
rect 73505 489 73705 495
rect 73505 455 73659 489
rect 73505 449 73705 455
rect 73505 163 73651 449
rect 73731 203 73811 523
rect 73795 164 73811 203
rect 73731 163 73811 164
rect 73927 495 74073 563
rect 74217 523 74233 563
rect 73927 489 74127 495
rect 73927 455 74081 489
rect 73927 449 74127 455
rect 73927 163 74073 449
rect 74153 203 74233 523
rect 74217 164 74233 203
rect 74153 163 74233 164
rect 74349 495 74495 563
rect 74639 523 74655 563
rect 74349 489 74549 495
rect 74349 455 74503 489
rect 74349 449 74549 455
rect 74349 163 74495 449
rect 74575 203 74655 523
rect 74639 164 74655 203
rect 74575 163 74655 164
rect 74771 495 74917 563
rect 75061 523 75077 563
rect 74771 489 74971 495
rect 74771 455 74925 489
rect 74771 449 74971 455
rect 74771 163 74917 449
rect 74997 203 75077 523
rect 75061 164 75077 203
rect 74997 163 75077 164
rect 75193 495 75339 563
rect 75483 523 75499 563
rect 75193 489 75393 495
rect 75193 455 75347 489
rect 75193 449 75393 455
rect 75193 163 75339 449
rect 75419 203 75499 523
rect 75483 164 75499 203
rect 75419 163 75499 164
rect 75615 495 75761 563
rect 75905 523 75921 563
rect 75615 489 75815 495
rect 75615 455 75769 489
rect 75615 449 75815 455
rect 75615 163 75761 449
rect 75841 203 75921 523
rect 75905 164 75921 203
rect 75841 163 75921 164
rect 76037 495 76183 563
rect 76327 523 76343 563
rect 76037 489 76237 495
rect 76037 455 76191 489
rect 76037 449 76237 455
rect 76037 163 76183 449
rect 76263 203 76343 523
rect 76327 164 76343 203
rect 76263 163 76343 164
rect 76459 495 76605 563
rect 76749 523 76765 563
rect 76459 489 76659 495
rect 76459 455 76613 489
rect 76459 449 76659 455
rect 76459 163 76605 449
rect 76685 203 76765 523
rect 76749 164 76765 203
rect 76685 163 76765 164
rect 76881 495 77027 563
rect 77171 523 77187 563
rect 76881 489 77081 495
rect 76881 455 77035 489
rect 76881 449 77081 455
rect 76881 163 77027 449
rect 77107 203 77187 523
rect 77171 164 77187 203
rect 77107 163 77187 164
rect 77303 495 77449 563
rect 77593 523 77609 563
rect 77303 489 77503 495
rect 77303 455 77457 489
rect 77303 449 77503 455
rect 77303 163 77449 449
rect 77529 203 77609 523
rect 77593 164 77609 203
rect 77529 163 77609 164
rect 77725 495 77871 563
rect 78015 523 78031 563
rect 77725 489 77925 495
rect 77725 455 77879 489
rect 77725 449 77925 455
rect 77725 163 77871 449
rect 77951 203 78031 523
rect 78015 164 78031 203
rect 77951 163 78031 164
rect 78147 495 78293 563
rect 78437 523 78453 563
rect 78147 489 78347 495
rect 78147 455 78301 489
rect 78147 449 78347 455
rect 78147 163 78293 449
rect 78373 203 78453 523
rect 78437 164 78453 203
rect 78373 163 78453 164
rect 78569 495 78715 563
rect 78859 523 78875 563
rect 78569 489 78769 495
rect 78569 455 78723 489
rect 78569 449 78769 455
rect 78569 163 78715 449
rect 78795 203 78875 523
rect 78859 164 78875 203
rect 78795 163 78875 164
rect 78991 495 79137 563
rect 79281 523 79297 563
rect 78991 489 79191 495
rect 78991 455 79145 489
rect 78991 449 79191 455
rect 78991 163 79137 449
rect 79217 203 79297 523
rect 79281 164 79297 203
rect 79217 163 79297 164
rect 79413 495 79559 563
rect 79703 523 79719 563
rect 79413 489 79613 495
rect 79413 455 79567 489
rect 79413 449 79613 455
rect 79413 163 79559 449
rect 79639 203 79719 523
rect 79703 164 79719 203
rect 79639 163 79719 164
rect 79835 495 79981 563
rect 80125 523 80141 563
rect 79835 489 80035 495
rect 79835 455 79989 489
rect 79835 449 80035 455
rect 79835 163 79981 449
rect 80061 203 80141 523
rect 80125 164 80141 203
rect 80061 163 80141 164
rect 80257 495 80403 563
rect 80547 523 80563 563
rect 80257 489 80457 495
rect 80257 455 80411 489
rect 80257 449 80457 455
rect 80257 163 80403 449
rect 80483 203 80563 523
rect 80547 164 80563 203
rect 80483 163 80563 164
rect 80679 495 80825 563
rect 80969 523 80985 563
rect 80679 489 80879 495
rect 80679 455 80833 489
rect 80679 449 80879 455
rect 80679 163 80825 449
rect 80905 203 80985 523
rect 80969 164 80985 203
rect 80905 163 80985 164
rect 81101 495 81247 563
rect 81391 523 81407 563
rect 81101 489 81301 495
rect 81101 455 81255 489
rect 81101 449 81301 455
rect 81101 163 81247 449
rect 81327 203 81407 523
rect 81391 164 81407 203
rect 81327 163 81407 164
rect 81523 495 81669 563
rect 81813 523 81829 563
rect 81523 489 81723 495
rect 81523 455 81677 489
rect 81523 449 81723 455
rect 81523 163 81669 449
rect 81749 203 81829 523
rect 81813 164 81829 203
rect 81749 163 81829 164
rect 81945 495 82091 563
rect 82235 523 82251 563
rect 81945 489 82145 495
rect 81945 455 82099 489
rect 81945 449 82145 455
rect 81945 163 82091 449
rect 82171 203 82251 523
rect 82235 164 82251 203
rect 82171 163 82251 164
rect 82367 495 82513 563
rect 82657 523 82673 563
rect 82367 489 82567 495
rect 82367 455 82521 489
rect 82367 449 82567 455
rect 82367 163 82513 449
rect 82593 203 82673 523
rect 82657 164 82673 203
rect 82593 163 82673 164
rect 82789 495 82935 563
rect 83079 523 83095 563
rect 82789 489 82989 495
rect 82789 455 82943 489
rect 82789 449 82989 455
rect 82789 163 82935 449
rect 83015 203 83095 523
rect 83079 164 83095 203
rect 83015 163 83095 164
rect 83211 495 83357 563
rect 83501 523 83517 563
rect 83211 489 83411 495
rect 83211 455 83365 489
rect 83211 449 83411 455
rect 83211 163 83357 449
rect 83437 203 83517 523
rect 83501 164 83517 203
rect 83437 163 83517 164
rect 83633 495 83779 563
rect 83923 523 83939 563
rect 83633 489 83833 495
rect 83633 455 83787 489
rect 83633 449 83833 455
rect 83633 163 83779 449
rect 83859 203 83939 523
rect 83923 164 83939 203
rect 83859 163 83939 164
rect 84055 495 84201 563
rect 84345 523 84361 563
rect 84055 489 84255 495
rect 84055 455 84209 489
rect 84055 449 84255 455
rect 84055 163 84201 449
rect 84281 203 84361 523
rect 84345 164 84361 203
rect 84281 163 84361 164
rect 84477 495 84623 563
rect 84767 523 84783 563
rect 84477 489 84677 495
rect 84477 455 84631 489
rect 84477 449 84677 455
rect 84477 163 84623 449
rect 84703 203 84783 523
rect 84767 164 84783 203
rect 84703 163 84783 164
rect 84899 495 85045 563
rect 85189 523 85205 563
rect 84899 489 85099 495
rect 84899 455 85053 489
rect 84899 449 85099 455
rect 84899 163 85045 449
rect 85125 203 85205 523
rect 85189 164 85205 203
rect 85125 163 85205 164
rect 85321 495 85467 563
rect 85611 523 85627 563
rect 85321 489 85521 495
rect 85321 455 85475 489
rect 85321 449 85521 455
rect 85321 163 85467 449
rect 85547 203 85627 523
rect 85611 164 85627 203
rect 85547 163 85627 164
rect 85743 495 85889 563
rect 86033 523 86049 563
rect 85743 489 85943 495
rect 85743 455 85897 489
rect 85743 449 85943 455
rect 85743 163 85889 449
rect 85969 203 86049 523
rect 86033 164 86049 203
rect 85969 163 86049 164
rect 86165 495 86311 563
rect 86455 523 86471 563
rect 86165 489 86365 495
rect 86165 455 86319 489
rect 86165 449 86365 455
rect 86165 163 86311 449
rect 86391 203 86471 523
rect 86455 164 86471 203
rect 86391 163 86471 164
rect 86587 495 86733 563
rect 86877 523 86893 563
rect 86587 489 86787 495
rect 86587 455 86741 489
rect 86587 449 86787 455
rect 86587 163 86733 449
rect 86813 203 86893 523
rect 86877 164 86893 203
rect 86813 163 86893 164
rect 87009 495 87155 563
rect 87299 523 87315 563
rect 87009 489 87209 495
rect 87009 455 87163 489
rect 87009 449 87209 455
rect 87009 163 87155 449
rect 87235 203 87315 523
rect 87299 164 87315 203
rect 87235 163 87315 164
rect 87431 495 87577 563
rect 87721 523 87737 563
rect 87431 489 87631 495
rect 87431 455 87585 489
rect 87431 449 87631 455
rect 87431 163 87577 449
rect 87657 203 87737 523
rect 87721 164 87737 203
rect 87657 163 87737 164
rect 87853 495 87999 563
rect 88143 523 88159 563
rect 87853 489 88053 495
rect 87853 455 88007 489
rect 87853 449 88053 455
rect 87853 163 87999 449
rect 88079 203 88159 523
rect 88143 164 88159 203
rect 88079 163 88159 164
rect 88275 495 88421 563
rect 88565 523 88581 563
rect 88275 489 88475 495
rect 88275 455 88429 489
rect 88275 449 88475 455
rect 88275 163 88421 449
rect 88501 203 88581 523
rect 88565 164 88581 203
rect 88501 163 88581 164
rect 88697 495 88843 563
rect 88987 523 89003 563
rect 88697 489 88897 495
rect 88697 455 88851 489
rect 88697 449 88897 455
rect 88697 163 88843 449
rect 88923 203 89003 523
rect 88987 164 89003 203
rect 88923 163 89003 164
rect 89119 495 89265 563
rect 89409 523 89425 563
rect 89119 489 89319 495
rect 89119 455 89273 489
rect 89119 449 89319 455
rect 89119 163 89265 449
rect 89345 203 89425 523
rect 89409 164 89425 203
rect 89345 163 89425 164
rect 89541 495 89687 563
rect 89831 523 89847 563
rect 89541 489 89741 495
rect 89541 455 89695 489
rect 89541 449 89741 455
rect 89541 163 89687 449
rect 89767 203 89847 523
rect 89831 164 89847 203
rect 89767 163 89847 164
rect 89963 495 90109 563
rect 90253 523 90269 563
rect 89963 489 90163 495
rect 89963 455 90117 489
rect 89963 449 90163 455
rect 89963 163 90109 449
rect 90189 203 90269 523
rect 90253 164 90269 203
rect 90189 163 90269 164
rect 90385 495 90531 563
rect 90675 523 90691 563
rect 90385 489 90585 495
rect 90385 455 90539 489
rect 90385 449 90585 455
rect 90385 163 90531 449
rect 90611 203 90691 523
rect 90675 164 90691 203
rect 90611 163 90691 164
rect 90807 495 90953 563
rect 91097 523 91113 563
rect 90807 489 91007 495
rect 90807 455 90961 489
rect 90807 449 91007 455
rect 90807 163 90953 449
rect 91033 203 91113 523
rect 91097 164 91113 203
rect 91033 163 91113 164
rect 91229 495 91375 563
rect 91519 523 91535 563
rect 91229 489 91429 495
rect 91229 455 91383 489
rect 91229 449 91429 455
rect 91229 163 91375 449
rect 91455 203 91535 523
rect 91519 164 91535 203
rect 91455 163 91535 164
rect 91651 495 91797 563
rect 91941 523 91957 563
rect 91651 489 91851 495
rect 91651 455 91805 489
rect 91651 449 91851 455
rect 91651 163 91797 449
rect 91877 203 91957 523
rect 91941 164 91957 203
rect 91877 163 91957 164
rect 92073 495 92219 563
rect 92363 523 92379 563
rect 92073 489 92273 495
rect 92073 455 92227 489
rect 92073 449 92273 455
rect 92073 163 92219 449
rect 92299 203 92379 523
rect 92363 164 92379 203
rect 92299 163 92379 164
rect 92495 495 92641 563
rect 92785 523 92801 563
rect 92495 489 92695 495
rect 92495 455 92649 489
rect 92495 449 92695 455
rect 92495 163 92641 449
rect 92721 203 92801 523
rect 92785 164 92801 203
rect 92721 163 92801 164
rect 92917 495 93063 563
rect 93207 523 93223 563
rect 92917 489 93117 495
rect 92917 455 93071 489
rect 92917 449 93117 455
rect 92917 163 93063 449
rect 93143 203 93223 523
rect 93207 164 93223 203
rect 93143 163 93223 164
rect 93339 495 93485 563
rect 93629 523 93645 563
rect 93339 489 93539 495
rect 93339 455 93493 489
rect 93339 449 93539 455
rect 93339 163 93485 449
rect 93565 203 93645 523
rect 93629 164 93645 203
rect 93565 163 93645 164
rect 93761 495 93907 563
rect 94051 523 94067 563
rect 93761 489 93961 495
rect 93761 455 93915 489
rect 93761 449 93961 455
rect 93761 163 93907 449
rect 93987 203 94067 523
rect 94051 164 94067 203
rect 93987 163 94067 164
rect 94183 495 94329 563
rect 94473 523 94489 563
rect 94183 489 94383 495
rect 94183 455 94337 489
rect 94183 449 94383 455
rect 94183 163 94329 449
rect 94409 203 94489 523
rect 94473 164 94489 203
rect 94409 163 94489 164
rect 94605 495 94751 563
rect 94895 523 94911 563
rect 94605 489 94805 495
rect 94605 455 94759 489
rect 94605 449 94805 455
rect 94605 163 94751 449
rect 94831 203 94911 523
rect 94895 164 94911 203
rect 94831 163 94911 164
rect 95027 495 95173 563
rect 95317 523 95333 563
rect 95027 489 95227 495
rect 95027 455 95181 489
rect 95027 449 95227 455
rect 95027 163 95173 449
rect 95253 203 95333 523
rect 95317 164 95333 203
rect 95253 163 95333 164
rect 95449 495 95595 563
rect 95739 523 95755 563
rect 95449 489 95649 495
rect 95449 455 95603 489
rect 95449 449 95649 455
rect 95449 163 95595 449
rect 95675 203 95755 523
rect 95739 164 95755 203
rect 95675 163 95755 164
rect 95871 495 96017 563
rect 96161 523 96177 563
rect 95871 489 96071 495
rect 95871 455 96025 489
rect 95871 449 96071 455
rect 95871 163 96017 449
rect 96097 203 96177 523
rect 96161 164 96177 203
rect 96097 163 96177 164
rect 96293 495 96439 563
rect 96583 523 96599 563
rect 96293 489 96493 495
rect 96293 455 96447 489
rect 96293 449 96493 455
rect 96293 163 96439 449
rect 96519 203 96599 523
rect 96583 164 96599 203
rect 96519 163 96599 164
rect 96715 495 96861 563
rect 97005 523 97021 563
rect 96715 489 96915 495
rect 96715 455 96869 489
rect 96715 449 96915 455
rect 96715 163 96861 449
rect 96941 203 97021 523
rect 97005 164 97021 203
rect 96941 163 97021 164
rect 97137 495 97283 563
rect 97427 523 97443 563
rect 97137 489 97337 495
rect 97137 455 97291 489
rect 97137 449 97337 455
rect 97137 163 97283 449
rect 97363 203 97443 523
rect 97427 164 97443 203
rect 97363 163 97443 164
rect 97559 495 97705 563
rect 97849 523 97865 563
rect 97559 489 97759 495
rect 97559 455 97713 489
rect 97559 449 97759 455
rect 97559 163 97705 449
rect 97785 203 97865 523
rect 97849 164 97865 203
rect 97785 163 97865 164
rect 97981 495 98127 563
rect 98271 523 98287 563
rect 97981 489 98181 495
rect 97981 455 98135 489
rect 97981 449 98181 455
rect 97981 163 98127 449
rect 98207 203 98287 523
rect 98271 164 98287 203
rect 98207 163 98287 164
rect 98403 495 98549 563
rect 98693 523 98709 563
rect 98403 489 98603 495
rect 98403 455 98557 489
rect 98403 449 98603 455
rect 98403 163 98549 449
rect 98629 203 98709 523
rect 98693 164 98709 203
rect 98629 163 98709 164
rect 98825 495 98971 563
rect 99115 523 99131 563
rect 98825 489 99025 495
rect 98825 455 98979 489
rect 98825 449 99025 455
rect 98825 163 98971 449
rect 99051 203 99131 523
rect 99115 164 99131 203
rect 99051 163 99131 164
rect 99247 495 99393 563
rect 99537 523 99553 563
rect 99247 489 99447 495
rect 99247 455 99401 489
rect 99247 449 99447 455
rect 99247 163 99393 449
rect 99473 203 99553 523
rect 99537 164 99553 203
rect 99473 163 99553 164
rect 99669 495 99815 563
rect 99959 523 99975 563
rect 99669 489 99869 495
rect 99669 455 99823 489
rect 99669 449 99869 455
rect 99669 163 99815 449
rect 99895 203 99975 523
rect 99959 164 99975 203
rect 99895 163 99975 164
rect 100091 495 100237 563
rect 100381 523 100397 563
rect 100091 489 100291 495
rect 100091 455 100245 489
rect 100091 449 100291 455
rect 100091 163 100237 449
rect 100317 203 100397 523
rect 100381 164 100397 203
rect 100317 163 100397 164
rect 100513 495 100659 563
rect 100803 523 100819 563
rect 100513 489 100713 495
rect 100513 455 100667 489
rect 100513 449 100713 455
rect 100513 163 100659 449
rect 100739 203 100819 523
rect 100803 164 100819 203
rect 100739 163 100819 164
rect 100935 495 101081 563
rect 101225 523 101241 563
rect 100935 489 101135 495
rect 100935 455 101089 489
rect 100935 449 101135 455
rect 100935 163 101081 449
rect 101161 203 101241 523
rect 101225 164 101241 203
rect 101161 163 101241 164
rect 101357 495 101503 563
rect 101647 523 101663 563
rect 101357 489 101557 495
rect 101357 455 101511 489
rect 101357 449 101557 455
rect 101357 163 101503 449
rect 101583 203 101663 523
rect 101647 164 101663 203
rect 101583 163 101663 164
rect 101779 495 101925 563
rect 102069 523 102085 563
rect 101779 489 101979 495
rect 101779 455 101933 489
rect 101779 449 101979 455
rect 101779 163 101925 449
rect 102005 203 102085 523
rect 102069 164 102085 203
rect 102005 163 102085 164
rect 102201 495 102347 563
rect 102491 523 102507 563
rect 102201 489 102401 495
rect 102201 455 102355 489
rect 102201 449 102401 455
rect 102201 163 102347 449
rect 102427 203 102507 523
rect 102491 164 102507 203
rect 102427 163 102507 164
rect 102623 495 102769 563
rect 102913 523 102929 563
rect 102623 489 102823 495
rect 102623 455 102777 489
rect 102623 449 102823 455
rect 102623 163 102769 449
rect 102849 203 102929 523
rect 102913 164 102929 203
rect 102849 163 102929 164
rect 103045 495 103191 563
rect 103335 523 103351 563
rect 103045 489 103245 495
rect 103045 455 103199 489
rect 103045 449 103245 455
rect 103045 163 103191 449
rect 103271 203 103351 523
rect 103335 164 103351 203
rect 103271 163 103351 164
rect 103467 495 103613 563
rect 103757 523 103773 563
rect 103467 489 103667 495
rect 103467 455 103621 489
rect 103467 449 103667 455
rect 103467 163 103613 449
rect 103693 203 103773 523
rect 103757 164 103773 203
rect 103693 163 103773 164
rect 103889 495 104035 563
rect 104179 523 104195 563
rect 103889 489 104089 495
rect 103889 455 104043 489
rect 103889 449 104089 455
rect 103889 163 104035 449
rect 104115 203 104195 523
rect 104179 164 104195 203
rect 104115 163 104195 164
rect 104311 495 104457 563
rect 104601 523 104617 563
rect 104311 489 104511 495
rect 104311 455 104465 489
rect 104311 449 104511 455
rect 104311 163 104457 449
rect 104537 203 104617 523
rect 104601 164 104617 203
rect 104537 163 104617 164
rect 104733 495 104879 563
rect 105023 523 105039 563
rect 104733 489 104933 495
rect 104733 455 104887 489
rect 104733 449 104933 455
rect 104733 163 104879 449
rect 104959 203 105039 523
rect 105023 164 105039 203
rect 104959 163 105039 164
rect 105155 495 105301 563
rect 105445 523 105461 563
rect 105155 489 105355 495
rect 105155 455 105309 489
rect 105155 449 105355 455
rect 105155 163 105301 449
rect 105381 203 105461 523
rect 105445 164 105461 203
rect 105381 163 105461 164
rect 105577 495 105723 563
rect 105867 523 105883 563
rect 105577 489 105777 495
rect 105577 455 105731 489
rect 105577 449 105777 455
rect 105577 163 105723 449
rect 105803 203 105883 523
rect 105867 164 105883 203
rect 105803 163 105883 164
rect 105999 495 106145 563
rect 106289 523 106305 563
rect 105999 489 106199 495
rect 105999 455 106153 489
rect 105999 449 106199 455
rect 105999 163 106145 449
rect 106225 203 106305 523
rect 106289 164 106305 203
rect 106225 163 106305 164
rect 106421 495 106567 563
rect 106711 523 106727 563
rect 106421 489 106621 495
rect 106421 455 106575 489
rect 106421 449 106621 455
rect 106421 163 106567 449
rect 106647 203 106727 523
rect 106711 164 106727 203
rect 106647 163 106727 164
rect 106843 495 106989 563
rect 107133 523 107149 563
rect 106843 489 107043 495
rect 106843 455 106997 489
rect 106843 449 107043 455
rect 106843 163 106989 449
rect 107069 203 107149 523
rect 107133 164 107149 203
rect 107069 163 107149 164
rect 107265 495 107411 563
rect 107555 523 107571 563
rect 107265 489 107465 495
rect 107265 455 107419 489
rect 107265 449 107465 455
rect 107265 163 107411 449
rect 107491 203 107571 523
rect 107555 164 107571 203
rect 107491 163 107571 164
rect 107687 495 107833 563
rect 107977 523 107993 563
rect 107687 489 107887 495
rect 107687 455 107841 489
rect 107687 449 107887 455
rect 107687 163 107833 449
rect 107913 203 107993 523
rect 107977 164 107993 203
rect 107913 163 107993 164
rect 108109 495 108255 563
rect 108399 523 108415 563
rect 108109 489 108309 495
rect 108109 455 108263 489
rect 108109 449 108309 455
rect 108109 163 108255 449
rect 108335 203 108415 523
rect 108399 164 108415 203
rect 108335 163 108415 164
rect 108531 495 108677 563
rect 108821 523 108837 563
rect 108531 489 108731 495
rect 108531 455 108685 489
rect 108531 449 108731 455
rect 108531 163 108677 449
rect 108757 203 108837 523
rect 108821 164 108837 203
rect 108757 163 108837 164
rect 108953 495 109099 563
rect 109243 523 109259 563
rect 108953 489 109153 495
rect 108953 455 109107 489
rect 108953 449 109153 455
rect 108953 163 109099 449
rect 109179 203 109259 523
rect 109243 164 109259 203
rect 109179 163 109259 164
rect 109375 495 109521 563
rect 109665 523 109681 563
rect 109375 489 109575 495
rect 109375 455 109529 489
rect 109375 449 109575 455
rect 109375 163 109521 449
rect 109601 203 109681 523
rect 109665 164 109681 203
rect 109601 163 109681 164
rect 109797 495 109943 563
rect 110087 523 110103 563
rect 109797 489 109997 495
rect 109797 455 109951 489
rect 109797 449 109997 455
rect 109797 163 109943 449
rect 110023 203 110103 523
rect 110087 164 110103 203
rect 110023 163 110103 164
rect 110219 495 110365 563
rect 110509 523 110525 563
rect 110219 489 110419 495
rect 110219 455 110373 489
rect 110219 449 110419 455
rect 110219 163 110365 449
rect 110445 203 110525 523
rect 110509 164 110525 203
rect 110445 163 110525 164
rect 110641 495 110787 563
rect 110931 523 110947 563
rect 110641 489 110841 495
rect 110641 455 110795 489
rect 110641 449 110841 455
rect 110641 163 110787 449
rect 110867 203 110947 523
rect 110931 164 110947 203
rect 110867 163 110947 164
rect 111063 495 111209 563
rect 111353 523 111369 563
rect 111063 489 111263 495
rect 111063 455 111217 489
rect 111063 449 111263 455
rect 111063 163 111209 449
rect 111289 203 111369 523
rect 111353 164 111369 203
rect 111289 163 111369 164
rect 111485 495 111631 563
rect 111775 523 111791 563
rect 111485 489 111685 495
rect 111485 455 111639 489
rect 111485 449 111685 455
rect 111485 163 111631 449
rect 111711 203 111791 523
rect 111775 164 111791 203
rect 111711 163 111791 164
rect 111907 495 112053 563
rect 112197 523 112213 563
rect 111907 489 112107 495
rect 111907 455 112061 489
rect 111907 449 112107 455
rect 111907 163 112053 449
rect 112133 203 112213 523
rect 112197 164 112213 203
rect 112133 163 112213 164
rect 112329 163 112475 563
rect 112619 523 112635 563
rect 112555 203 112635 523
rect 112619 164 112635 203
rect 112555 163 112635 164
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
use hgu_sw_cap  x1[0]
timestamp 1697348449
transform 1 0 111920 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[1]
timestamp 1697348449
transform 1 0 111498 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[2]
timestamp 1697348449
transform 1 0 111076 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[3]
timestamp 1697348449
transform 1 0 110654 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[4]
timestamp 1697348449
transform 1 0 110232 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[5]
timestamp 1697348449
transform 1 0 109810 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[6]
timestamp 1697348449
transform 1 0 109388 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[7]
timestamp 1697348449
transform 1 0 108966 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[8]
timestamp 1697348449
transform 1 0 108544 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[9]
timestamp 1697348449
transform 1 0 108122 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[10]
timestamp 1697348449
transform 1 0 107700 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[11]
timestamp 1697348449
transform 1 0 107278 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[12]
timestamp 1697348449
transform 1 0 106856 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[13]
timestamp 1697348449
transform 1 0 106434 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[14]
timestamp 1697348449
transform 1 0 106012 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[15]
timestamp 1697348449
transform 1 0 105590 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[16]
timestamp 1697348449
transform 1 0 105168 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[17]
timestamp 1697348449
transform 1 0 104746 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[18]
timestamp 1697348449
transform 1 0 104324 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[19]
timestamp 1697348449
transform 1 0 103902 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[20]
timestamp 1697348449
transform 1 0 103480 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[21]
timestamp 1697348449
transform 1 0 103058 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[22]
timestamp 1697348449
transform 1 0 102636 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[23]
timestamp 1697348449
transform 1 0 102214 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[24]
timestamp 1697348449
transform 1 0 101792 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[25]
timestamp 1697348449
transform 1 0 101370 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[26]
timestamp 1697348449
transform 1 0 100948 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[27]
timestamp 1697348449
transform 1 0 100526 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[28]
timestamp 1697348449
transform 1 0 100104 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[29]
timestamp 1697348449
transform 1 0 99682 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[30]
timestamp 1697348449
transform 1 0 99260 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[31]
timestamp 1697348449
transform 1 0 98838 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[32]
timestamp 1697348449
transform 1 0 98416 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[33]
timestamp 1697348449
transform 1 0 97994 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[34]
timestamp 1697348449
transform 1 0 97572 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[35]
timestamp 1697348449
transform 1 0 97150 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[36]
timestamp 1697348449
transform 1 0 96728 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[37]
timestamp 1697348449
transform 1 0 96306 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[38]
timestamp 1697348449
transform 1 0 95884 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[39]
timestamp 1697348449
transform 1 0 95462 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[40]
timestamp 1697348449
transform 1 0 95040 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[41]
timestamp 1697348449
transform 1 0 94618 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[42]
timestamp 1697348449
transform 1 0 94196 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[43]
timestamp 1697348449
transform 1 0 93774 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[44]
timestamp 1697348449
transform 1 0 93352 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[45]
timestamp 1697348449
transform 1 0 92930 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[46]
timestamp 1697348449
transform 1 0 92508 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[47]
timestamp 1697348449
transform 1 0 92086 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[48]
timestamp 1697348449
transform 1 0 91664 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[49]
timestamp 1697348449
transform 1 0 91242 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[50]
timestamp 1697348449
transform 1 0 90820 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[51]
timestamp 1697348449
transform 1 0 90398 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[52]
timestamp 1697348449
transform 1 0 89976 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[53]
timestamp 1697348449
transform 1 0 89554 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[54]
timestamp 1697348449
transform 1 0 89132 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[55]
timestamp 1697348449
transform 1 0 88710 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[56]
timestamp 1697348449
transform 1 0 88288 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[57]
timestamp 1697348449
transform 1 0 87866 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[58]
timestamp 1697348449
transform 1 0 87444 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[59]
timestamp 1697348449
transform 1 0 87022 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[60]
timestamp 1697348449
transform 1 0 86600 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[61]
timestamp 1697348449
transform 1 0 86178 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[62]
timestamp 1697348449
transform 1 0 85756 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[63]
timestamp 1697348449
transform 1 0 85334 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[64]
timestamp 1697348449
transform 1 0 84912 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[65]
timestamp 1697348449
transform 1 0 84490 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[66]
timestamp 1697348449
transform 1 0 84068 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[67]
timestamp 1697348449
transform 1 0 83646 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[68]
timestamp 1697348449
transform 1 0 83224 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[69]
timestamp 1697348449
transform 1 0 82802 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[70]
timestamp 1697348449
transform 1 0 82380 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[71]
timestamp 1697348449
transform 1 0 81958 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[72]
timestamp 1697348449
transform 1 0 81536 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[73]
timestamp 1697348449
transform 1 0 81114 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[74]
timestamp 1697348449
transform 1 0 80692 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[75]
timestamp 1697348449
transform 1 0 80270 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[76]
timestamp 1697348449
transform 1 0 79848 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[77]
timestamp 1697348449
transform 1 0 79426 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[78]
timestamp 1697348449
transform 1 0 79004 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[79]
timestamp 1697348449
transform 1 0 78582 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[80]
timestamp 1697348449
transform 1 0 78160 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[81]
timestamp 1697348449
transform 1 0 77738 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[82]
timestamp 1697348449
transform 1 0 77316 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[83]
timestamp 1697348449
transform 1 0 76894 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[84]
timestamp 1697348449
transform 1 0 76472 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[85]
timestamp 1697348449
transform 1 0 76050 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[86]
timestamp 1697348449
transform 1 0 75628 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[87]
timestamp 1697348449
transform 1 0 75206 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[88]
timestamp 1697348449
transform 1 0 74784 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[89]
timestamp 1697348449
transform 1 0 74362 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[90]
timestamp 1697348449
transform 1 0 73940 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[91]
timestamp 1697348449
transform 1 0 73518 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[92]
timestamp 1697348449
transform 1 0 73096 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[93]
timestamp 1697348449
transform 1 0 72674 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[94]
timestamp 1697348449
transform 1 0 72252 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[95]
timestamp 1697348449
transform 1 0 71830 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[96]
timestamp 1697348449
transform 1 0 71408 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[97]
timestamp 1697348449
transform 1 0 70986 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[98]
timestamp 1697348449
transform 1 0 70564 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[99]
timestamp 1697348449
transform 1 0 70142 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[100]
timestamp 1697348449
transform 1 0 69720 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[101]
timestamp 1697348449
transform 1 0 69298 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[102]
timestamp 1697348449
transform 1 0 68876 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[103]
timestamp 1697348449
transform 1 0 68454 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[104]
timestamp 1697348449
transform 1 0 68032 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[105]
timestamp 1697348449
transform 1 0 67610 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[106]
timestamp 1697348449
transform 1 0 67188 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[107]
timestamp 1697348449
transform 1 0 66766 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[108]
timestamp 1697348449
transform 1 0 66344 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[109]
timestamp 1697348449
transform 1 0 65922 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[110]
timestamp 1697348449
transform 1 0 65500 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[111]
timestamp 1697348449
transform 1 0 65078 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[112]
timestamp 1697348449
transform 1 0 64656 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[113]
timestamp 1697348449
transform 1 0 64234 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[114]
timestamp 1697348449
transform 1 0 63812 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[115]
timestamp 1697348449
transform 1 0 63390 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[116]
timestamp 1697348449
transform 1 0 62968 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[117]
timestamp 1697348449
transform 1 0 62546 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[118]
timestamp 1697348449
transform 1 0 62124 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[119]
timestamp 1697348449
transform 1 0 61702 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[120]
timestamp 1697348449
transform 1 0 61280 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[121]
timestamp 1697348449
transform 1 0 60858 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[122]
timestamp 1697348449
transform 1 0 60436 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[123]
timestamp 1697348449
transform 1 0 60014 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[124]
timestamp 1697348449
transform 1 0 59592 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[125]
timestamp 1697348449
transform 1 0 59170 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[126]
timestamp 1697348449
transform 1 0 58748 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x1[127]
timestamp 1697348449
transform 1 0 58326 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x2
timestamp 1697348449
transform 1 0 4732 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x3[0]
timestamp 1697348449
transform 1 0 5576 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x3[1]
timestamp 1697348449
transform 1 0 5154 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x4[0]
timestamp 1697348449
transform 1 0 7264 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x4[1]
timestamp 1697348449
transform 1 0 6842 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x4[2]
timestamp 1697348449
transform 1 0 6420 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x4[3]
timestamp 1697348449
transform 1 0 5998 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x5[0]
timestamp 1697348449
transform 1 0 10640 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x5[1]
timestamp 1697348449
transform 1 0 10218 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x5[2]
timestamp 1697348449
transform 1 0 9796 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x5[3]
timestamp 1697348449
transform 1 0 9374 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x5[4]
timestamp 1697348449
transform 1 0 8952 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x5[5]
timestamp 1697348449
transform 1 0 8530 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x5[6]
timestamp 1697348449
transform 1 0 8108 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x5[7]
timestamp 1697348449
transform 1 0 7686 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x6[0]
timestamp 1697348449
transform 1 0 17392 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x6[1]
timestamp 1697348449
transform 1 0 16970 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x6[2]
timestamp 1697348449
transform 1 0 16548 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x6[3]
timestamp 1697348449
transform 1 0 16126 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x6[4]
timestamp 1697348449
transform 1 0 15704 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x6[5]
timestamp 1697348449
transform 1 0 15282 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x6[6]
timestamp 1697348449
transform 1 0 14860 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x6[7]
timestamp 1697348449
transform 1 0 14438 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x6[8]
timestamp 1697348449
transform 1 0 14016 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x6[9]
timestamp 1697348449
transform 1 0 13594 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x6[10]
timestamp 1697348449
transform 1 0 13172 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x6[11]
timestamp 1697348449
transform 1 0 12750 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x6[12]
timestamp 1697348449
transform 1 0 12328 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x6[13]
timestamp 1697348449
transform 1 0 11906 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x6[14]
timestamp 1697348449
transform 1 0 11484 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x6[15]
timestamp 1697348449
transform 1 0 11062 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[0]
timestamp 1697348449
transform 1 0 30896 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[1]
timestamp 1697348449
transform 1 0 30474 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[2]
timestamp 1697348449
transform 1 0 30052 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[3]
timestamp 1697348449
transform 1 0 29630 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[4]
timestamp 1697348449
transform 1 0 29208 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[5]
timestamp 1697348449
transform 1 0 28786 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[6]
timestamp 1697348449
transform 1 0 28364 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[7]
timestamp 1697348449
transform 1 0 27942 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[8]
timestamp 1697348449
transform 1 0 27520 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[9]
timestamp 1697348449
transform 1 0 27098 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[10]
timestamp 1697348449
transform 1 0 26676 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[11]
timestamp 1697348449
transform 1 0 26254 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[12]
timestamp 1697348449
transform 1 0 25832 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[13]
timestamp 1697348449
transform 1 0 25410 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[14]
timestamp 1697348449
transform 1 0 24988 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[15]
timestamp 1697348449
transform 1 0 24566 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[16]
timestamp 1697348449
transform 1 0 24144 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[17]
timestamp 1697348449
transform 1 0 23722 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[18]
timestamp 1697348449
transform 1 0 23300 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[19]
timestamp 1697348449
transform 1 0 22878 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[20]
timestamp 1697348449
transform 1 0 22456 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[21]
timestamp 1697348449
transform 1 0 22034 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[22]
timestamp 1697348449
transform 1 0 21612 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[23]
timestamp 1697348449
transform 1 0 21190 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[24]
timestamp 1697348449
transform 1 0 20768 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[25]
timestamp 1697348449
transform 1 0 20346 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[26]
timestamp 1697348449
transform 1 0 19924 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[27]
timestamp 1697348449
transform 1 0 19502 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[28]
timestamp 1697348449
transform 1 0 19080 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[29]
timestamp 1697348449
transform 1 0 18658 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[30]
timestamp 1697348449
transform 1 0 18236 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x7[31]
timestamp 1697348449
transform 1 0 17814 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[0]
timestamp 1697348449
transform 1 0 57904 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[1]
timestamp 1697348449
transform 1 0 57482 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[2]
timestamp 1697348449
transform 1 0 57060 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[3]
timestamp 1697348449
transform 1 0 56638 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[4]
timestamp 1697348449
transform 1 0 56216 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[5]
timestamp 1697348449
transform 1 0 55794 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[6]
timestamp 1697348449
transform 1 0 55372 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[7]
timestamp 1697348449
transform 1 0 54950 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[8]
timestamp 1697348449
transform 1 0 54528 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[9]
timestamp 1697348449
transform 1 0 54106 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[10]
timestamp 1697348449
transform 1 0 53684 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[11]
timestamp 1697348449
transform 1 0 53262 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[12]
timestamp 1697348449
transform 1 0 52840 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[13]
timestamp 1697348449
transform 1 0 52418 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[14]
timestamp 1697348449
transform 1 0 51996 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[15]
timestamp 1697348449
transform 1 0 51574 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[16]
timestamp 1697348449
transform 1 0 51152 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[17]
timestamp 1697348449
transform 1 0 50730 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[18]
timestamp 1697348449
transform 1 0 50308 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[19]
timestamp 1697348449
transform 1 0 49886 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[20]
timestamp 1697348449
transform 1 0 49464 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[21]
timestamp 1697348449
transform 1 0 49042 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[22]
timestamp 1697348449
transform 1 0 48620 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[23]
timestamp 1697348449
transform 1 0 48198 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[24]
timestamp 1697348449
transform 1 0 47776 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[25]
timestamp 1697348449
transform 1 0 47354 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[26]
timestamp 1697348449
transform 1 0 46932 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[27]
timestamp 1697348449
transform 1 0 46510 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[28]
timestamp 1697348449
transform 1 0 46088 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[29]
timestamp 1697348449
transform 1 0 45666 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[30]
timestamp 1697348449
transform 1 0 45244 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[31]
timestamp 1697348449
transform 1 0 44822 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[32]
timestamp 1697348449
transform 1 0 44400 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[33]
timestamp 1697348449
transform 1 0 43978 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[34]
timestamp 1697348449
transform 1 0 43556 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[35]
timestamp 1697348449
transform 1 0 43134 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[36]
timestamp 1697348449
transform 1 0 42712 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[37]
timestamp 1697348449
transform 1 0 42290 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[38]
timestamp 1697348449
transform 1 0 41868 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[39]
timestamp 1697348449
transform 1 0 41446 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[40]
timestamp 1697348449
transform 1 0 41024 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[41]
timestamp 1697348449
transform 1 0 40602 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[42]
timestamp 1697348449
transform 1 0 40180 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[43]
timestamp 1697348449
transform 1 0 39758 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[44]
timestamp 1697348449
transform 1 0 39336 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[45]
timestamp 1697348449
transform 1 0 38914 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[46]
timestamp 1697348449
transform 1 0 38492 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[47]
timestamp 1697348449
transform 1 0 38070 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[48]
timestamp 1697348449
transform 1 0 37648 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[49]
timestamp 1697348449
transform 1 0 37226 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[50]
timestamp 1697348449
transform 1 0 36804 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[51]
timestamp 1697348449
transform 1 0 36382 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[52]
timestamp 1697348449
transform 1 0 35960 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[53]
timestamp 1697348449
transform 1 0 35538 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[54]
timestamp 1697348449
transform 1 0 35116 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[55]
timestamp 1697348449
transform 1 0 34694 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[56]
timestamp 1697348449
transform 1 0 34272 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[57]
timestamp 1697348449
transform 1 0 33850 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[58]
timestamp 1697348449
transform 1 0 33428 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[59]
timestamp 1697348449
transform 1 0 33006 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[60]
timestamp 1697348449
transform 1 0 32584 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[61]
timestamp 1697348449
transform 1 0 32162 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[62]
timestamp 1697348449
transform 1 0 31740 0 1 1776
box -53 -1653 1141 200
use hgu_sw_cap  x8[63]
timestamp 1697348449
transform 1 0 31318 0 1 1776
box -53 -1653 1141 200
use sky130_fd_pr__nfet_01v8_J3KQQP  XM1
timestamp 1697025759
transform 1 0 512 0 1 799
box -565 -252 565 252
use sky130_fd_pr__pfet_01v8_GVE7YE  XM2
timestamp 1697025759
transform 1 0 1370 0 1 793
box -346 -299 346 299
use sky130_fd_pr__nfet_01v8_WENHSZ  XM3
timestamp 1697025759
transform 1 0 2064 0 1 789
box -401 -348 401 348
use sky130_fd_pr__nfet_01v8_L7T3GD  XM4
timestamp 1697025759
transform 1 0 2623 0 1 640
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_XYUFBL  XM5
timestamp 1697025759
transform 1 0 2992 0 1 634
box -211 -299 211 299
use sky130_fd_pr__nfet_01v8_L7T3GD  XM6
timestamp 1697025759
transform 1 0 3361 0 1 534
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_XYUFBL  XM7
timestamp 1697025759
transform 1 0 3730 0 1 528
box -211 -299 211 299
use sky130_fd_pr__nfet_01v8_9NW3WL  XM8
timestamp 1697025759
transform 1 0 4099 0 1 470
box -211 -294 211 294
use sky130_fd_pr__pfet_01v8_XCA4BL  XM9
timestamp 1697025759
transform 1 0 4468 0 1 502
box -211 -379 211 379
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 IN
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 OUT
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 VSS
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE\[0\]}
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE\[1\]}
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE\[2\]}
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE\[3\]}
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 {}
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE\[4\]}
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE\[5\]}
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE\[6\]}
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE\[7\]}
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 {}
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 DELAY_CAP=DELAY_CAP
port 14 nsew
<< end >>
