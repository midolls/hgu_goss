magic
tech sky130A
timestamp 1697616495
<< end >>
