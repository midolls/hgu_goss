magic
tech sky130A
magscale 1 2
timestamp 1699422110
<< error_s >>
rect 13752 4957 13761 4962
rect 13795 4957 13804 4962
rect 13752 4953 13804 4957
rect 13743 4944 13745 4953
rect 13752 4948 13808 4953
rect 13743 4901 13745 4910
rect 13752 4906 13757 4948
rect 13799 4906 13808 4948
rect 13811 4944 13813 4953
rect 13752 4901 13808 4906
rect 13811 4901 13813 4910
rect 13752 4892 13761 4901
rect 13795 4892 13804 4901
<< nwell >>
rect 13332 6954 18192 6996
rect 13332 5670 18192 5724
<< psubdiff >>
rect 13370 7581 13399 7615
rect 13433 7581 13491 7615
rect 13525 7581 13583 7615
rect 13617 7581 13675 7615
rect 13709 7581 13767 7615
rect 13801 7581 13859 7615
rect 13893 7581 13951 7615
rect 13985 7581 14043 7615
rect 14077 7581 14135 7615
rect 14169 7581 14226 7615
rect 14260 7581 14319 7615
rect 14353 7581 14411 7615
rect 14445 7581 14503 7615
rect 14537 7581 14595 7615
rect 14629 7581 14687 7615
rect 14721 7581 14779 7615
rect 14813 7581 14871 7615
rect 14905 7581 14963 7615
rect 14997 7581 15055 7615
rect 15089 7581 15147 7615
rect 15181 7581 15239 7615
rect 15273 7581 15331 7615
rect 15365 7581 15423 7615
rect 15457 7581 15515 7615
rect 15549 7581 15607 7615
rect 15641 7581 15699 7615
rect 15733 7581 15791 7615
rect 15825 7581 15883 7615
rect 15917 7581 15975 7615
rect 16009 7581 16067 7615
rect 16101 7581 16159 7615
rect 16193 7581 16251 7615
rect 16285 7581 16343 7615
rect 16377 7581 16435 7615
rect 16469 7581 16527 7615
rect 16561 7581 16619 7615
rect 16653 7581 16711 7615
rect 16745 7581 16803 7615
rect 16837 7581 16895 7615
rect 16929 7581 16987 7615
rect 17021 7581 17079 7615
rect 17113 7581 17171 7615
rect 17205 7581 17263 7615
rect 17297 7581 17355 7615
rect 17389 7581 17447 7615
rect 17481 7581 17539 7615
rect 17573 7581 17631 7615
rect 17665 7581 17723 7615
rect 17757 7581 17815 7615
rect 17849 7581 17907 7615
rect 17941 7581 17999 7615
rect 18033 7581 18091 7615
rect 18125 7581 18154 7615
rect 13370 6316 13399 6350
rect 13433 6316 13491 6350
rect 13525 6316 13583 6350
rect 13617 6316 13675 6350
rect 13709 6316 13767 6350
rect 13801 6316 13859 6350
rect 13893 6316 13951 6350
rect 13985 6316 14043 6350
rect 14077 6316 14135 6350
rect 14169 6316 14227 6350
rect 14261 6316 14319 6350
rect 14353 6316 14411 6350
rect 14445 6316 14503 6350
rect 14537 6316 14595 6350
rect 14629 6316 14687 6350
rect 14721 6316 14779 6350
rect 14813 6316 14871 6350
rect 14905 6316 14964 6350
rect 14998 6316 15055 6350
rect 15089 6316 15147 6350
rect 15181 6316 15239 6350
rect 15273 6316 15332 6350
rect 15366 6316 15423 6350
rect 15457 6316 15515 6350
rect 15549 6316 15607 6350
rect 15641 6316 15699 6350
rect 15733 6316 15791 6350
rect 15825 6316 15883 6350
rect 15917 6316 15975 6350
rect 16009 6316 16067 6350
rect 16101 6316 16159 6350
rect 16193 6316 16251 6350
rect 16285 6316 16343 6350
rect 16377 6316 16435 6350
rect 16469 6316 16526 6350
rect 16560 6316 16618 6350
rect 16652 6316 16711 6350
rect 16745 6316 16803 6350
rect 16837 6316 16895 6350
rect 16929 6316 16986 6350
rect 17020 6316 17079 6350
rect 17113 6316 17170 6350
rect 17204 6316 17263 6350
rect 17297 6316 17355 6350
rect 17389 6316 17447 6350
rect 17481 6316 17539 6350
rect 17573 6316 17631 6350
rect 17665 6316 17723 6350
rect 17757 6316 17815 6350
rect 17849 6316 17907 6350
rect 17941 6316 17999 6350
rect 18033 6316 18091 6350
rect 18125 6316 18154 6350
rect 13370 5049 13399 5083
rect 13433 5049 13491 5083
rect 13525 5049 13583 5083
rect 13617 5049 13675 5083
rect 13709 5049 13767 5083
rect 13801 5049 13859 5083
rect 13893 5049 13951 5083
rect 13985 5049 14043 5083
rect 14077 5049 14135 5083
rect 14169 5049 14227 5083
rect 14261 5049 14319 5083
rect 14353 5049 14411 5083
rect 14445 5049 14503 5083
rect 14537 5049 14595 5083
rect 14629 5049 14687 5083
rect 14721 5049 14779 5083
rect 14813 5049 14871 5083
rect 14905 5049 14963 5083
rect 14997 5049 15055 5083
rect 15089 5049 15147 5083
rect 15181 5049 15239 5083
rect 15273 5049 15331 5083
rect 15365 5049 15423 5083
rect 15457 5049 15515 5083
rect 15549 5049 15607 5083
rect 15641 5049 15699 5083
rect 15733 5049 15791 5083
rect 15825 5049 15883 5083
rect 15917 5049 15975 5083
rect 16009 5049 16067 5083
rect 16101 5049 16159 5083
rect 16193 5049 16251 5083
rect 16285 5049 16343 5083
rect 16377 5049 16435 5083
rect 16469 5049 16527 5083
rect 16561 5049 16619 5083
rect 16653 5049 16711 5083
rect 16745 5049 16803 5083
rect 16837 5049 16895 5083
rect 16929 5049 16987 5083
rect 17021 5049 17079 5083
rect 17113 5049 17171 5083
rect 17205 5049 17263 5083
rect 17297 5049 17355 5083
rect 17389 5049 17447 5083
rect 17481 5049 17539 5083
rect 17573 5049 17631 5083
rect 17665 5049 17723 5083
rect 17757 5049 17815 5083
rect 17849 5049 17907 5083
rect 17941 5049 17999 5083
rect 18033 5049 18091 5083
rect 18125 5049 18154 5083
<< nsubdiff >>
rect 13370 6955 13400 6989
rect 13434 6955 13491 6989
rect 13525 6955 13584 6989
rect 13618 6955 13675 6989
rect 13709 6955 13766 6989
rect 13800 6955 13860 6989
rect 13894 6955 13951 6989
rect 13985 6955 14044 6989
rect 14078 6955 14135 6989
rect 14169 6955 14227 6989
rect 14261 6955 14318 6989
rect 14352 6955 14411 6989
rect 14445 6955 14504 6989
rect 14538 6955 14595 6989
rect 14629 6955 14687 6989
rect 14721 6955 14779 6989
rect 14813 6955 14871 6989
rect 14905 6955 14963 6989
rect 14997 6955 15055 6989
rect 15089 6955 15147 6989
rect 15181 6955 15240 6989
rect 15274 6955 15330 6989
rect 15364 6955 15423 6989
rect 15457 6955 15516 6989
rect 15550 6955 15608 6989
rect 15642 6955 15699 6989
rect 15733 6955 15792 6989
rect 15826 6955 15884 6989
rect 15918 6955 15976 6989
rect 16010 6955 16068 6989
rect 16102 6955 16160 6989
rect 16194 6955 16252 6989
rect 16286 6955 16343 6989
rect 16377 6955 16434 6989
rect 16468 6955 16527 6989
rect 16561 6955 16620 6989
rect 16654 6955 16712 6989
rect 16746 6955 16803 6989
rect 16837 6955 16897 6989
rect 16931 6955 16987 6989
rect 17021 6955 17078 6989
rect 17112 6955 17171 6989
rect 17205 6955 17264 6989
rect 17298 6955 17356 6989
rect 17390 6955 17447 6989
rect 17481 6955 17539 6989
rect 17573 6955 17631 6989
rect 17665 6955 17722 6989
rect 17756 6955 17814 6989
rect 17848 6955 17907 6989
rect 17941 6955 17999 6989
rect 18033 6955 18091 6989
rect 18125 6955 18154 6989
rect 13370 5674 13402 5708
rect 13436 5674 13492 5708
rect 13526 5674 13585 5708
rect 13619 5674 13675 5708
rect 13709 5674 13766 5708
rect 13800 5674 13860 5708
rect 13894 5674 13951 5708
rect 13985 5674 14043 5708
rect 14077 5674 14135 5708
rect 14169 5674 14228 5708
rect 14262 5674 14319 5708
rect 14353 5674 14411 5708
rect 14445 5674 14503 5708
rect 14537 5674 14595 5708
rect 14629 5674 14688 5708
rect 14722 5674 14779 5708
rect 14813 5674 14870 5708
rect 14904 5674 14963 5708
rect 14997 5674 15056 5708
rect 15090 5674 15147 5708
rect 15181 5674 15239 5708
rect 15273 5674 15331 5708
rect 15365 5674 15423 5708
rect 15457 5674 15516 5708
rect 15550 5674 15606 5708
rect 15640 5674 15699 5708
rect 15733 5674 15791 5708
rect 15825 5674 15884 5708
rect 15918 5674 15978 5708
rect 16012 5674 16067 5708
rect 16101 5674 16159 5708
rect 16193 5674 16251 5708
rect 16285 5674 16343 5708
rect 16377 5674 16435 5708
rect 16469 5674 16527 5708
rect 16561 5674 16619 5708
rect 16653 5674 16711 5708
rect 16745 5674 16803 5708
rect 16837 5674 16895 5708
rect 16929 5674 16987 5708
rect 17021 5674 17079 5708
rect 17113 5674 17171 5708
rect 17205 5674 17263 5708
rect 17297 5674 17355 5708
rect 17389 5674 17447 5708
rect 17481 5674 17539 5708
rect 17573 5674 17631 5708
rect 17665 5674 17723 5708
rect 17757 5674 17815 5708
rect 17849 5674 17907 5708
rect 17941 5674 18000 5708
rect 18034 5674 18091 5708
rect 18125 5674 18154 5708
<< psubdiffcont >>
rect 13399 7581 13433 7615
rect 13491 7581 13525 7615
rect 13583 7581 13617 7615
rect 13675 7581 13709 7615
rect 13767 7581 13801 7615
rect 13859 7581 13893 7615
rect 13951 7581 13985 7615
rect 14043 7581 14077 7615
rect 14135 7581 14169 7615
rect 14226 7581 14260 7615
rect 14319 7581 14353 7615
rect 14411 7581 14445 7615
rect 14503 7581 14537 7615
rect 14595 7581 14629 7615
rect 14687 7581 14721 7615
rect 14779 7581 14813 7615
rect 14871 7581 14905 7615
rect 14963 7581 14997 7615
rect 15055 7581 15089 7615
rect 15147 7581 15181 7615
rect 15239 7581 15273 7615
rect 15331 7581 15365 7615
rect 15423 7581 15457 7615
rect 15515 7581 15549 7615
rect 15607 7581 15641 7615
rect 15699 7581 15733 7615
rect 15791 7581 15825 7615
rect 15883 7581 15917 7615
rect 15975 7581 16009 7615
rect 16067 7581 16101 7615
rect 16159 7581 16193 7615
rect 16251 7581 16285 7615
rect 16343 7581 16377 7615
rect 16435 7581 16469 7615
rect 16527 7581 16561 7615
rect 16619 7581 16653 7615
rect 16711 7581 16745 7615
rect 16803 7581 16837 7615
rect 16895 7581 16929 7615
rect 16987 7581 17021 7615
rect 17079 7581 17113 7615
rect 17171 7581 17205 7615
rect 17263 7581 17297 7615
rect 17355 7581 17389 7615
rect 17447 7581 17481 7615
rect 17539 7581 17573 7615
rect 17631 7581 17665 7615
rect 17723 7581 17757 7615
rect 17815 7581 17849 7615
rect 17907 7581 17941 7615
rect 17999 7581 18033 7615
rect 18091 7581 18125 7615
rect 13399 6316 13433 6350
rect 13491 6316 13525 6350
rect 13583 6316 13617 6350
rect 13675 6316 13709 6350
rect 13767 6316 13801 6350
rect 13859 6316 13893 6350
rect 13951 6316 13985 6350
rect 14043 6316 14077 6350
rect 14135 6316 14169 6350
rect 14227 6316 14261 6350
rect 14319 6316 14353 6350
rect 14411 6316 14445 6350
rect 14503 6316 14537 6350
rect 14595 6316 14629 6350
rect 14687 6316 14721 6350
rect 14779 6316 14813 6350
rect 14871 6316 14905 6350
rect 14964 6316 14998 6350
rect 15055 6316 15089 6350
rect 15147 6316 15181 6350
rect 15239 6316 15273 6350
rect 15332 6316 15366 6350
rect 15423 6316 15457 6350
rect 15515 6316 15549 6350
rect 15607 6316 15641 6350
rect 15699 6316 15733 6350
rect 15791 6316 15825 6350
rect 15883 6316 15917 6350
rect 15975 6316 16009 6350
rect 16067 6316 16101 6350
rect 16159 6316 16193 6350
rect 16251 6316 16285 6350
rect 16343 6316 16377 6350
rect 16435 6316 16469 6350
rect 16526 6316 16560 6350
rect 16618 6316 16652 6350
rect 16711 6316 16745 6350
rect 16803 6316 16837 6350
rect 16895 6316 16929 6350
rect 16986 6316 17020 6350
rect 17079 6316 17113 6350
rect 17170 6316 17204 6350
rect 17263 6316 17297 6350
rect 17355 6316 17389 6350
rect 17447 6316 17481 6350
rect 17539 6316 17573 6350
rect 17631 6316 17665 6350
rect 17723 6316 17757 6350
rect 17815 6316 17849 6350
rect 17907 6316 17941 6350
rect 17999 6316 18033 6350
rect 18091 6316 18125 6350
rect 13399 5049 13433 5083
rect 13491 5049 13525 5083
rect 13583 5049 13617 5083
rect 13675 5049 13709 5083
rect 13767 5049 13801 5083
rect 13859 5049 13893 5083
rect 13951 5049 13985 5083
rect 14043 5049 14077 5083
rect 14135 5049 14169 5083
rect 14227 5049 14261 5083
rect 14319 5049 14353 5083
rect 14411 5049 14445 5083
rect 14503 5049 14537 5083
rect 14595 5049 14629 5083
rect 14687 5049 14721 5083
rect 14779 5049 14813 5083
rect 14871 5049 14905 5083
rect 14963 5049 14997 5083
rect 15055 5049 15089 5083
rect 15147 5049 15181 5083
rect 15239 5049 15273 5083
rect 15331 5049 15365 5083
rect 15423 5049 15457 5083
rect 15515 5049 15549 5083
rect 15607 5049 15641 5083
rect 15699 5049 15733 5083
rect 15791 5049 15825 5083
rect 15883 5049 15917 5083
rect 15975 5049 16009 5083
rect 16067 5049 16101 5083
rect 16159 5049 16193 5083
rect 16251 5049 16285 5083
rect 16343 5049 16377 5083
rect 16435 5049 16469 5083
rect 16527 5049 16561 5083
rect 16619 5049 16653 5083
rect 16711 5049 16745 5083
rect 16803 5049 16837 5083
rect 16895 5049 16929 5083
rect 16987 5049 17021 5083
rect 17079 5049 17113 5083
rect 17171 5049 17205 5083
rect 17263 5049 17297 5083
rect 17355 5049 17389 5083
rect 17447 5049 17481 5083
rect 17539 5049 17573 5083
rect 17631 5049 17665 5083
rect 17723 5049 17757 5083
rect 17815 5049 17849 5083
rect 17907 5049 17941 5083
rect 17999 5049 18033 5083
rect 18091 5049 18125 5083
<< nsubdiffcont >>
rect 13400 6955 13434 6989
rect 13491 6955 13525 6989
rect 13584 6955 13618 6989
rect 13675 6955 13709 6989
rect 13766 6955 13800 6989
rect 13860 6955 13894 6989
rect 13951 6955 13985 6989
rect 14044 6955 14078 6989
rect 14135 6955 14169 6989
rect 14227 6955 14261 6989
rect 14318 6955 14352 6989
rect 14411 6955 14445 6989
rect 14504 6955 14538 6989
rect 14595 6955 14629 6989
rect 14687 6955 14721 6989
rect 14779 6955 14813 6989
rect 14871 6955 14905 6989
rect 14963 6955 14997 6989
rect 15055 6955 15089 6989
rect 15147 6955 15181 6989
rect 15240 6955 15274 6989
rect 15330 6955 15364 6989
rect 15423 6955 15457 6989
rect 15516 6955 15550 6989
rect 15608 6955 15642 6989
rect 15699 6955 15733 6989
rect 15792 6955 15826 6989
rect 15884 6955 15918 6989
rect 15976 6955 16010 6989
rect 16068 6955 16102 6989
rect 16160 6955 16194 6989
rect 16252 6955 16286 6989
rect 16343 6955 16377 6989
rect 16434 6955 16468 6989
rect 16527 6955 16561 6989
rect 16620 6955 16654 6989
rect 16712 6955 16746 6989
rect 16803 6955 16837 6989
rect 16897 6955 16931 6989
rect 16987 6955 17021 6989
rect 17078 6955 17112 6989
rect 17171 6955 17205 6989
rect 17264 6955 17298 6989
rect 17356 6955 17390 6989
rect 17447 6955 17481 6989
rect 17539 6955 17573 6989
rect 17631 6955 17665 6989
rect 17722 6955 17756 6989
rect 17814 6955 17848 6989
rect 17907 6955 17941 6989
rect 17999 6955 18033 6989
rect 18091 6955 18125 6989
rect 13402 5674 13436 5708
rect 13492 5674 13526 5708
rect 13585 5674 13619 5708
rect 13675 5674 13709 5708
rect 13766 5674 13800 5708
rect 13860 5674 13894 5708
rect 13951 5674 13985 5708
rect 14043 5674 14077 5708
rect 14135 5674 14169 5708
rect 14228 5674 14262 5708
rect 14319 5674 14353 5708
rect 14411 5674 14445 5708
rect 14503 5674 14537 5708
rect 14595 5674 14629 5708
rect 14688 5674 14722 5708
rect 14779 5674 14813 5708
rect 14870 5674 14904 5708
rect 14963 5674 14997 5708
rect 15056 5674 15090 5708
rect 15147 5674 15181 5708
rect 15239 5674 15273 5708
rect 15331 5674 15365 5708
rect 15423 5674 15457 5708
rect 15516 5674 15550 5708
rect 15606 5674 15640 5708
rect 15699 5674 15733 5708
rect 15791 5674 15825 5708
rect 15884 5674 15918 5708
rect 15978 5674 16012 5708
rect 16067 5674 16101 5708
rect 16159 5674 16193 5708
rect 16251 5674 16285 5708
rect 16343 5674 16377 5708
rect 16435 5674 16469 5708
rect 16527 5674 16561 5708
rect 16619 5674 16653 5708
rect 16711 5674 16745 5708
rect 16803 5674 16837 5708
rect 16895 5674 16929 5708
rect 16987 5674 17021 5708
rect 17079 5674 17113 5708
rect 17171 5674 17205 5708
rect 17263 5674 17297 5708
rect 17355 5674 17389 5708
rect 17447 5674 17481 5708
rect 17539 5674 17573 5708
rect 17631 5674 17665 5708
rect 17723 5674 17757 5708
rect 17815 5674 17849 5708
rect 17907 5674 17941 5708
rect 18000 5674 18034 5708
rect 18091 5674 18125 5708
<< locali >>
rect 13370 7581 13399 7615
rect 13433 7581 13491 7615
rect 13525 7581 13583 7615
rect 13617 7581 13675 7615
rect 13709 7581 13767 7615
rect 13801 7581 13859 7615
rect 13893 7581 13951 7615
rect 13985 7581 14043 7615
rect 14077 7581 14135 7615
rect 14169 7581 14226 7615
rect 14260 7581 14319 7615
rect 14353 7581 14411 7615
rect 14445 7581 14503 7615
rect 14537 7581 14595 7615
rect 14629 7581 14687 7615
rect 14721 7581 14779 7615
rect 14813 7581 14871 7615
rect 14905 7581 14963 7615
rect 14997 7581 15055 7615
rect 15089 7581 15147 7615
rect 15181 7581 15239 7615
rect 15273 7581 15331 7615
rect 15365 7581 15423 7615
rect 15457 7581 15515 7615
rect 15549 7581 15607 7615
rect 15641 7581 15699 7615
rect 15733 7581 15791 7615
rect 15825 7581 15883 7615
rect 15917 7581 15975 7615
rect 16009 7581 16067 7615
rect 16101 7581 16159 7615
rect 16193 7581 16251 7615
rect 16285 7581 16343 7615
rect 16377 7581 16435 7615
rect 16469 7581 16527 7615
rect 16561 7581 16619 7615
rect 16653 7581 16711 7615
rect 16745 7581 16803 7615
rect 16837 7581 16895 7615
rect 16929 7581 16987 7615
rect 17021 7581 17079 7615
rect 17113 7581 17171 7615
rect 17205 7581 17263 7615
rect 17297 7581 17355 7615
rect 17389 7581 17447 7615
rect 17481 7581 17539 7615
rect 17573 7581 17631 7615
rect 17665 7581 17723 7615
rect 17757 7581 17815 7615
rect 17849 7581 17907 7615
rect 17941 7581 17999 7615
rect 18033 7581 18091 7615
rect 18125 7581 18154 7615
rect 13370 6989 18154 7008
rect 13370 6955 13400 6989
rect 13434 6955 13491 6989
rect 13525 6955 13584 6989
rect 13618 6955 13675 6989
rect 13709 6955 13766 6989
rect 13800 6955 13860 6989
rect 13894 6955 13951 6989
rect 13985 6955 14044 6989
rect 14078 6955 14135 6989
rect 14169 6955 14227 6989
rect 14261 6955 14318 6989
rect 14352 6955 14411 6989
rect 14445 6955 14504 6989
rect 14538 6955 14595 6989
rect 14629 6955 14687 6989
rect 14721 6955 14779 6989
rect 14813 6955 14871 6989
rect 14905 6955 14963 6989
rect 14997 6955 15055 6989
rect 15089 6955 15147 6989
rect 15181 6955 15240 6989
rect 15274 6955 15330 6989
rect 15364 6955 15423 6989
rect 15457 6955 15516 6989
rect 15550 6955 15608 6989
rect 15642 6955 15699 6989
rect 15733 6955 15792 6989
rect 15826 6955 15884 6989
rect 15918 6955 15976 6989
rect 16010 6955 16068 6989
rect 16102 6955 16160 6989
rect 16194 6955 16252 6989
rect 16286 6955 16343 6989
rect 16377 6955 16434 6989
rect 16468 6955 16527 6989
rect 16561 6955 16620 6989
rect 16654 6955 16712 6989
rect 16746 6955 16803 6989
rect 16837 6955 16897 6989
rect 16931 6955 16987 6989
rect 17021 6955 17078 6989
rect 17112 6955 17171 6989
rect 17205 6955 17264 6989
rect 17298 6955 17356 6989
rect 17390 6955 17447 6989
rect 17481 6955 17539 6989
rect 17573 6955 17631 6989
rect 17665 6955 17722 6989
rect 17756 6955 17814 6989
rect 17848 6955 17907 6989
rect 17941 6955 17999 6989
rect 18033 6955 18091 6989
rect 18125 6955 18154 6989
rect 13370 6933 18154 6955
rect 13370 6350 18154 6367
rect 13370 6316 13399 6350
rect 13433 6316 13491 6350
rect 13525 6316 13583 6350
rect 13617 6316 13675 6350
rect 13709 6316 13767 6350
rect 13801 6316 13859 6350
rect 13893 6316 13951 6350
rect 13985 6316 14043 6350
rect 14077 6316 14135 6350
rect 14169 6316 14227 6350
rect 14261 6316 14319 6350
rect 14353 6316 14411 6350
rect 14445 6316 14503 6350
rect 14537 6316 14595 6350
rect 14629 6316 14687 6350
rect 14721 6316 14779 6350
rect 14813 6316 14871 6350
rect 14905 6316 14964 6350
rect 14998 6316 15055 6350
rect 15089 6316 15147 6350
rect 15181 6316 15239 6350
rect 15273 6316 15332 6350
rect 15366 6316 15423 6350
rect 15457 6316 15515 6350
rect 15549 6316 15607 6350
rect 15641 6316 15699 6350
rect 15733 6316 15791 6350
rect 15825 6316 15883 6350
rect 15917 6316 15975 6350
rect 16009 6316 16067 6350
rect 16101 6316 16159 6350
rect 16193 6316 16251 6350
rect 16285 6316 16343 6350
rect 16377 6316 16435 6350
rect 16469 6316 16526 6350
rect 16560 6316 16618 6350
rect 16652 6316 16711 6350
rect 16745 6316 16803 6350
rect 16837 6316 16895 6350
rect 16929 6316 16986 6350
rect 17020 6316 17079 6350
rect 17113 6316 17170 6350
rect 17204 6316 17263 6350
rect 17297 6316 17355 6350
rect 17389 6316 17447 6350
rect 17481 6316 17539 6350
rect 17573 6316 17631 6350
rect 17665 6316 17723 6350
rect 17757 6316 17815 6350
rect 17849 6316 17907 6350
rect 17941 6316 17999 6350
rect 18033 6316 18091 6350
rect 18125 6316 18154 6350
rect 13370 6292 18154 6316
rect 13370 5708 18154 5726
rect 13370 5674 13402 5708
rect 13436 5674 13492 5708
rect 13526 5674 13585 5708
rect 13619 5674 13675 5708
rect 13709 5674 13766 5708
rect 13800 5674 13860 5708
rect 13894 5674 13951 5708
rect 13985 5674 14043 5708
rect 14077 5674 14135 5708
rect 14169 5674 14228 5708
rect 14262 5674 14319 5708
rect 14353 5674 14411 5708
rect 14445 5674 14503 5708
rect 14537 5674 14595 5708
rect 14629 5674 14688 5708
rect 14722 5674 14779 5708
rect 14813 5674 14870 5708
rect 14904 5674 14963 5708
rect 14997 5674 15056 5708
rect 15090 5674 15147 5708
rect 15181 5674 15239 5708
rect 15273 5674 15331 5708
rect 15365 5674 15423 5708
rect 15457 5674 15516 5708
rect 15550 5674 15606 5708
rect 15640 5674 15699 5708
rect 15733 5674 15791 5708
rect 15825 5674 15884 5708
rect 15918 5674 15978 5708
rect 16012 5674 16067 5708
rect 16101 5674 16159 5708
rect 16193 5674 16251 5708
rect 16285 5674 16343 5708
rect 16377 5674 16435 5708
rect 16469 5674 16527 5708
rect 16561 5674 16619 5708
rect 16653 5674 16711 5708
rect 16745 5674 16803 5708
rect 16837 5674 16895 5708
rect 16929 5674 16987 5708
rect 17021 5674 17079 5708
rect 17113 5674 17171 5708
rect 17205 5674 17263 5708
rect 17297 5674 17355 5708
rect 17389 5674 17447 5708
rect 17481 5674 17539 5708
rect 17573 5674 17631 5708
rect 17665 5674 17723 5708
rect 17757 5674 17815 5708
rect 17849 5674 17907 5708
rect 17941 5674 18000 5708
rect 18034 5674 18091 5708
rect 18125 5674 18154 5708
rect 13370 5651 18154 5674
rect 13370 5049 13399 5083
rect 13433 5049 13491 5083
rect 13525 5049 13583 5083
rect 13617 5049 13675 5083
rect 13709 5049 13767 5083
rect 13801 5049 13859 5083
rect 13893 5049 13951 5083
rect 13985 5049 14043 5083
rect 14077 5049 14135 5083
rect 14169 5049 14227 5083
rect 14261 5049 14319 5083
rect 14353 5049 14411 5083
rect 14445 5049 14503 5083
rect 14537 5049 14595 5083
rect 14629 5049 14687 5083
rect 14721 5049 14779 5083
rect 14813 5049 14871 5083
rect 14905 5049 14963 5083
rect 14997 5049 15055 5083
rect 15089 5049 15147 5083
rect 15181 5049 15239 5083
rect 15273 5049 15331 5083
rect 15365 5049 15423 5083
rect 15457 5049 15515 5083
rect 15549 5049 15607 5083
rect 15641 5049 15699 5083
rect 15733 5049 15791 5083
rect 15825 5049 15883 5083
rect 15917 5049 15975 5083
rect 16009 5049 16067 5083
rect 16101 5049 16159 5083
rect 16193 5049 16251 5083
rect 16285 5049 16343 5083
rect 16377 5049 16435 5083
rect 16469 5049 16527 5083
rect 16561 5049 16619 5083
rect 16653 5049 16711 5083
rect 16745 5049 16803 5083
rect 16837 5049 16895 5083
rect 16929 5049 16987 5083
rect 17021 5049 17079 5083
rect 17113 5049 17171 5083
rect 17205 5049 17263 5083
rect 17297 5049 17355 5083
rect 17389 5049 17447 5083
rect 17481 5049 17539 5083
rect 17573 5049 17631 5083
rect 17665 5049 17723 5083
rect 17757 5049 17815 5083
rect 17849 5049 17907 5083
rect 17941 5049 17999 5083
rect 18033 5049 18091 5083
rect 18125 5049 18154 5083
<< viali >>
rect 13416 7294 13450 7328
rect 15805 7276 15839 7310
rect 13417 6625 13451 6659
rect 15806 6628 15840 6662
rect 13419 6011 13453 6045
rect 15803 6011 15837 6045
rect 13415 5336 13449 5370
rect 15804 5325 15838 5359
<< metal1 >>
rect 18424 9269 18495 9315
rect 17602 7984 17899 7991
rect 13338 7918 13937 7946
rect 16645 7890 16703 7963
rect 13338 7862 16703 7890
rect 17501 7834 17560 7954
rect 13338 7806 17560 7834
rect 17602 7778 17934 7984
rect 13285 7750 17934 7778
rect 13285 7612 13339 7750
rect 13409 7655 13415 7707
rect 13467 7695 13473 7707
rect 15803 7695 15809 7707
rect 13467 7667 15809 7695
rect 13467 7655 13473 7667
rect 15803 7655 15809 7667
rect 15861 7695 15867 7707
rect 18467 7695 18495 9269
rect 15861 7667 18495 7695
rect 15861 7655 15867 7667
rect 13285 7516 13400 7612
rect 13491 7581 13525 7615
rect 13583 7581 13617 7615
rect 13675 7581 13709 7615
rect 13767 7581 13801 7615
rect 13859 7581 13893 7615
rect 13951 7581 13985 7615
rect 14043 7581 14077 7615
rect 14135 7581 14169 7615
rect 14226 7581 14260 7615
rect 14319 7581 14353 7615
rect 14411 7581 14445 7615
rect 14503 7581 14537 7615
rect 14595 7581 14629 7615
rect 14687 7581 14721 7615
rect 14779 7581 14813 7615
rect 14871 7581 14905 7615
rect 14963 7581 14997 7615
rect 15055 7581 15089 7615
rect 15147 7581 15181 7615
rect 15239 7581 15273 7615
rect 15331 7581 15365 7615
rect 15423 7581 15457 7615
rect 15515 7581 15549 7615
rect 15607 7581 15641 7615
rect 15699 7581 15733 7615
rect 15791 7581 15825 7615
rect 15883 7581 15917 7615
rect 15975 7581 16009 7615
rect 16067 7581 16101 7615
rect 16159 7581 16193 7615
rect 16251 7581 16285 7615
rect 16343 7581 16377 7615
rect 16435 7581 16469 7615
rect 16527 7581 16561 7615
rect 16619 7581 16653 7615
rect 16711 7581 16745 7615
rect 16803 7581 16837 7615
rect 16895 7581 16929 7615
rect 16987 7581 17021 7615
rect 17079 7581 17113 7615
rect 17171 7581 17205 7615
rect 17263 7581 17297 7615
rect 17355 7581 17389 7615
rect 17447 7581 17481 7615
rect 17539 7581 17573 7615
rect 17631 7581 17665 7615
rect 17723 7581 17757 7615
rect 17815 7581 17849 7615
rect 17907 7581 17941 7615
rect 17999 7581 18033 7615
rect 18091 7581 18125 7615
rect 13406 7337 13458 7343
rect 13406 7279 13458 7285
rect 15798 7322 15850 7328
rect 15798 7264 15850 7270
rect 13491 6954 13525 6988
rect 13584 6955 13618 6989
rect 15792 6954 15826 6988
rect 13407 6669 13459 6675
rect 13407 6611 13459 6617
rect 15797 6673 15849 6679
rect 15797 6615 15849 6621
rect 13399 6315 13433 6349
rect 13491 6316 13525 6350
rect 13583 6316 13617 6350
rect 13675 6316 13709 6350
rect 13767 6316 13801 6350
rect 13859 6316 13893 6350
rect 13951 6316 13985 6350
rect 14043 6316 14077 6350
rect 14135 6316 14169 6350
rect 14227 6316 14261 6350
rect 14319 6316 14353 6350
rect 14411 6316 14445 6350
rect 14503 6316 14537 6350
rect 14595 6316 14629 6350
rect 14687 6316 14721 6350
rect 14779 6316 14813 6350
rect 14871 6316 14905 6350
rect 14964 6316 14998 6350
rect 15055 6316 15089 6350
rect 15147 6316 15181 6350
rect 15239 6316 15273 6350
rect 15332 6316 15366 6350
rect 15423 6316 15457 6350
rect 15515 6316 15549 6350
rect 15607 6316 15641 6350
rect 15699 6316 15733 6350
rect 15791 6316 15825 6350
rect 15883 6316 15917 6350
rect 15975 6316 16009 6350
rect 16067 6316 16101 6350
rect 16159 6316 16193 6350
rect 16251 6316 16285 6350
rect 16343 6316 16377 6350
rect 16435 6316 16469 6350
rect 16526 6316 16560 6350
rect 16618 6316 16652 6350
rect 16711 6316 16745 6350
rect 16803 6316 16837 6350
rect 16895 6316 16929 6350
rect 16986 6316 17020 6350
rect 17079 6316 17113 6350
rect 17170 6316 17204 6350
rect 17263 6316 17297 6350
rect 17355 6316 17389 6350
rect 17447 6316 17481 6350
rect 17539 6316 17573 6350
rect 17631 6316 17665 6350
rect 17723 6316 17757 6350
rect 17815 6316 17849 6350
rect 17907 6316 17941 6350
rect 17999 6316 18033 6350
rect 18091 6316 18125 6350
rect 13409 6056 13461 6062
rect 13409 5998 13461 6004
rect 15796 6057 15848 6063
rect 15796 5999 15848 6005
rect 13404 5381 13456 5387
rect 13404 5323 13456 5329
rect 15797 5370 15849 5376
rect 15797 5312 15849 5318
rect 13399 5049 13433 5083
rect 13491 5049 13525 5083
rect 13583 5049 13617 5083
rect 13675 5049 13709 5083
rect 13767 5049 13801 5083
rect 13859 5049 13893 5083
rect 13951 5049 13985 5083
rect 14043 5049 14077 5083
rect 14135 5049 14169 5083
rect 14227 5049 14261 5083
rect 14319 5049 14353 5083
rect 14411 5049 14445 5083
rect 14503 5049 14537 5083
rect 14595 5049 14629 5083
rect 14687 5049 14721 5083
rect 14779 5049 14813 5083
rect 14871 5049 14905 5083
rect 14963 5049 14997 5083
rect 15055 5049 15089 5083
rect 15147 5049 15181 5083
rect 15239 5049 15273 5083
rect 15331 5049 15365 5083
rect 15423 5049 15457 5083
rect 15515 5049 15549 5083
rect 15607 5049 15641 5083
rect 15699 5049 15733 5083
rect 15791 5049 15825 5083
rect 15883 5049 15917 5083
rect 15975 5049 16009 5083
rect 16067 5049 16101 5083
rect 16159 5049 16193 5083
rect 16251 5049 16285 5083
rect 16343 5049 16377 5083
rect 16435 5049 16469 5083
rect 16527 5049 16561 5083
rect 16619 5049 16653 5083
rect 16711 5049 16745 5083
rect 16803 5049 16837 5083
rect 16895 5049 16929 5083
rect 16987 5049 17021 5083
rect 17079 5049 17113 5083
rect 17171 5049 17205 5083
rect 17263 5049 17297 5083
rect 17355 5049 17389 5083
rect 17447 5049 17481 5083
rect 17539 5049 17573 5083
rect 17631 5049 17665 5083
rect 17723 5049 17757 5083
rect 17815 5049 17849 5083
rect 17907 5049 17941 5083
rect 17999 5049 18033 5083
rect 18091 5049 18125 5083
rect 13745 4901 13752 4953
rect 13804 4901 13811 4953
<< via1 >>
rect 13415 7655 13467 7707
rect 15809 7655 15861 7707
rect 13406 7328 13458 7337
rect 13406 7294 13416 7328
rect 13416 7294 13450 7328
rect 13450 7294 13458 7328
rect 13406 7285 13458 7294
rect 15798 7310 15850 7322
rect 15798 7276 15805 7310
rect 15805 7276 15839 7310
rect 15839 7276 15850 7310
rect 15798 7270 15850 7276
rect 13407 6659 13459 6669
rect 13407 6625 13417 6659
rect 13417 6625 13451 6659
rect 13451 6625 13459 6659
rect 13407 6617 13459 6625
rect 15797 6662 15849 6673
rect 15797 6628 15806 6662
rect 15806 6628 15840 6662
rect 15840 6628 15849 6662
rect 15797 6621 15849 6628
rect 13409 6045 13461 6056
rect 13409 6011 13419 6045
rect 13419 6011 13453 6045
rect 13453 6011 13461 6045
rect 13409 6004 13461 6011
rect 15796 6045 15848 6057
rect 15796 6011 15803 6045
rect 15803 6011 15837 6045
rect 15837 6011 15848 6045
rect 15796 6005 15848 6011
rect 13404 5370 13456 5381
rect 13404 5336 13415 5370
rect 13415 5336 13449 5370
rect 13449 5336 13456 5370
rect 13404 5329 13456 5336
rect 15797 5359 15849 5370
rect 15797 5325 15804 5359
rect 15804 5325 15838 5359
rect 15838 5325 15849 5359
rect 15797 5318 15849 5325
rect 13752 4901 13804 4953
<< metal2 >>
rect 13409 7655 13415 7707
rect 13467 7655 13473 7707
rect 15803 7655 15809 7707
rect 15861 7655 15867 7707
rect 13428 7343 13456 7655
rect 13406 7337 13458 7343
rect 15822 7328 15850 7655
rect 13406 7279 13458 7285
rect 15798 7322 15850 7328
rect 13428 6675 13456 7279
rect 15798 7264 15850 7270
rect 15822 6679 15850 7264
rect 13407 6669 13459 6675
rect 13407 6611 13459 6617
rect 15797 6673 15850 6679
rect 15849 6621 15850 6673
rect 15797 6615 15850 6621
rect 13428 6062 13456 6611
rect 15822 6063 15850 6615
rect 13409 6056 13461 6062
rect 13409 5998 13461 6004
rect 15796 6057 15850 6063
rect 15848 6005 15850 6057
rect 15796 5999 15850 6005
rect 13428 5387 13456 5998
rect 13404 5381 13456 5387
rect 15822 5376 15850 5999
rect 13404 5323 13456 5329
rect 13428 5294 13456 5323
rect 15797 5370 15850 5376
rect 15849 5318 15850 5370
rect 15797 5312 15850 5318
rect 15822 5294 15850 5312
rect 13745 4901 13752 4953
rect 13804 4901 13811 4953
<< via2 >>
rect 13752 4901 13804 4953
<< metal4 >>
rect 11836 10013 12254 10623
rect 18267 10492 19041 10623
rect 18267 10217 18493 10492
rect 18590 10217 19041 10492
rect 18267 9636 19041 10217
rect 11864 7966 12240 9403
rect 11864 7481 18154 7966
rect 12771 6704 13267 7481
rect 18545 7351 19041 9636
rect 13330 6866 19043 7351
rect 12771 6219 18193 6704
rect 12771 5525 13267 6219
rect 18545 6076 19041 6866
rect 13327 5591 19043 6076
rect 12771 5040 18195 5525
use sky130_fd_sc_hd__dfbbp_1  x1[0] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697358018
transform 1 0 13370 0 -1 7564
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x1[1]
timestamp 1697358018
transform 1 0 15762 0 -1 7564
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x1[2]
timestamp 1697358018
transform 1 0 13370 0 1 6380
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x1[3]
timestamp 1697358018
transform 1 0 15762 0 1 6380
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x1[4]
timestamp 1697358018
transform 1 0 13370 0 -1 6284
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x1[5]
timestamp 1697358018
transform 1 0 15762 0 -1 6284
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x1[6]
timestamp 1697358018
transform 1 0 13370 0 1 5100
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x1[7]
timestamp 1697358018
transform 1 0 15762 0 1 5100
box -38 -48 2430 592
use hgu_delay_no_code  x2
timestamp 1699326296
transform 1 0 2492 0 1 7675
box 9238 267 15997 2986
<< labels >>
flabel metal4 11864 7966 12240 9403 0 FreeSans 320 0 0 0 VSS
port 1 nsew
flabel metal4 11836 10013 12254 10623 0 FreeSans 320 0 0 0 VDD
port 2 nsew
<< end >>
