magic
tech sky130A
magscale 1 2
timestamp 1698474146
<< pwell >>
rect 1006 1014 1032 1046
<< metal3 >>
rect 686 1824 1358 1826
rect 686 1760 790 1824
rect 854 1760 870 1824
rect 934 1760 950 1824
rect 1014 1760 1030 1824
rect 1094 1760 1110 1824
rect 1174 1760 1190 1824
rect 1254 1760 1358 1824
rect 686 1758 1358 1760
rect 686 1604 752 1758
rect 686 1540 687 1604
rect 751 1540 752 1604
rect 686 1524 752 1540
rect 686 1460 687 1524
rect 751 1460 752 1524
rect 686 1444 752 1460
rect 686 1380 687 1444
rect 751 1380 752 1444
rect 686 1364 752 1380
rect 686 1300 687 1364
rect 751 1300 752 1364
rect 686 1284 752 1300
rect 686 1220 687 1284
rect 751 1220 752 1284
rect 686 1204 752 1220
rect 686 1140 687 1204
rect 751 1140 752 1204
rect 686 1124 752 1140
rect 686 1060 687 1124
rect 751 1060 752 1124
rect 686 1044 752 1060
rect 686 980 687 1044
rect 751 980 752 1044
rect 686 964 752 980
rect 686 900 687 964
rect 751 900 752 964
rect 686 884 752 900
rect 686 820 687 884
rect 751 820 752 884
rect 686 730 752 820
rect 812 726 872 1758
rect 932 666 992 1696
rect 1052 726 1112 1758
rect 1172 666 1232 1696
rect 1292 1604 1358 1758
rect 1292 1540 1293 1604
rect 1357 1540 1358 1604
rect 1292 1524 1358 1540
rect 1292 1460 1293 1524
rect 1357 1460 1358 1524
rect 1292 1444 1358 1460
rect 1292 1380 1293 1444
rect 1357 1380 1358 1444
rect 1292 1364 1358 1380
rect 1292 1300 1293 1364
rect 1357 1300 1358 1364
rect 1292 1284 1358 1300
rect 1292 1220 1293 1284
rect 1357 1220 1358 1284
rect 1292 1204 1358 1220
rect 1292 1140 1293 1204
rect 1357 1140 1358 1204
rect 1292 1124 1358 1140
rect 1292 1060 1293 1124
rect 1357 1060 1358 1124
rect 1292 1044 1358 1060
rect 1292 980 1293 1044
rect 1357 980 1358 1044
rect 1292 964 1358 980
rect 1292 900 1293 964
rect 1357 900 1358 964
rect 1292 884 1358 900
rect 1292 820 1293 884
rect 1357 820 1358 884
rect 1292 730 1358 820
rect 686 664 1358 666
rect 686 600 790 664
rect 854 600 870 664
rect 934 600 950 664
rect 1014 600 1030 664
rect 1094 600 1110 664
rect 1174 600 1190 664
rect 1254 600 1358 664
rect 686 598 1358 600
<< via3 >>
rect 790 1760 854 1824
rect 870 1760 934 1824
rect 950 1760 1014 1824
rect 1030 1760 1094 1824
rect 1110 1760 1174 1824
rect 1190 1760 1254 1824
rect 687 1540 751 1604
rect 687 1460 751 1524
rect 687 1380 751 1444
rect 687 1300 751 1364
rect 687 1220 751 1284
rect 687 1140 751 1204
rect 687 1060 751 1124
rect 687 980 751 1044
rect 687 900 751 964
rect 687 820 751 884
rect 1293 1540 1357 1604
rect 1293 1460 1357 1524
rect 1293 1380 1357 1444
rect 1293 1300 1357 1364
rect 1293 1220 1357 1284
rect 1293 1140 1357 1204
rect 1293 1060 1357 1124
rect 1293 980 1357 1044
rect 1293 900 1357 964
rect 1293 820 1357 884
rect 790 600 854 664
rect 870 600 934 664
rect 950 600 1014 664
rect 1030 600 1094 664
rect 1110 600 1174 664
rect 1190 600 1254 664
<< metal4 >>
rect 686 1824 1358 1826
rect 686 1760 790 1824
rect 854 1760 870 1824
rect 934 1760 950 1824
rect 1014 1760 1030 1824
rect 1094 1760 1110 1824
rect 1174 1760 1190 1824
rect 1254 1760 1358 1824
rect 686 1758 1358 1760
rect 686 1604 752 1758
rect 686 1540 687 1604
rect 751 1540 752 1604
rect 686 1524 752 1540
rect 686 1460 687 1524
rect 751 1460 752 1524
rect 686 1444 752 1460
rect 686 1380 687 1444
rect 751 1380 752 1444
rect 686 1364 752 1380
rect 686 1300 687 1364
rect 751 1300 752 1364
rect 686 1284 752 1300
rect 686 1220 687 1284
rect 751 1220 752 1284
rect 686 1204 752 1220
rect 686 1140 687 1204
rect 751 1140 752 1204
rect 686 1124 752 1140
rect 686 1060 687 1124
rect 751 1060 752 1124
rect 686 1044 752 1060
rect 686 980 687 1044
rect 751 980 752 1044
rect 686 964 752 980
rect 686 900 687 964
rect 751 900 752 964
rect 686 884 752 900
rect 686 820 687 884
rect 751 820 752 884
rect 686 730 752 820
rect 812 666 872 1696
rect 932 726 992 1758
rect 1052 666 1112 1696
rect 1172 726 1232 1758
rect 1292 1604 1358 1758
rect 1292 1540 1293 1604
rect 1357 1540 1358 1604
rect 1292 1524 1358 1540
rect 1292 1460 1293 1524
rect 1357 1460 1358 1524
rect 1292 1444 1358 1460
rect 1292 1380 1293 1444
rect 1357 1380 1358 1444
rect 1292 1364 1358 1380
rect 1292 1300 1293 1364
rect 1357 1300 1358 1364
rect 1292 1284 1358 1300
rect 1292 1220 1293 1284
rect 1357 1220 1358 1284
rect 1292 1204 1358 1220
rect 1292 1140 1293 1204
rect 1357 1140 1358 1204
rect 1292 1124 1358 1140
rect 1292 1060 1293 1124
rect 1357 1060 1358 1124
rect 1292 1044 1358 1060
rect 1292 980 1293 1044
rect 1357 980 1358 1044
rect 1292 964 1358 980
rect 1292 900 1293 964
rect 1357 900 1358 964
rect 1292 884 1358 900
rect 1292 820 1293 884
rect 1357 820 1358 884
rect 1292 730 1358 820
rect 686 664 1358 666
rect 686 600 790 664
rect 854 600 870 664
rect 934 600 950 664
rect 1014 600 1030 664
rect 1094 600 1110 664
rect 1174 600 1190 664
rect 1254 600 1358 664
rect 686 598 1358 600
<< labels >>
flabel pwell 1006 1014 1032 1046 0 FreeSans 160 0 0 0 SUB
port 9 nsew
flabel metal4 948 1348 974 1380 0 FreeSans 320 0 0 0 CBOT
port 4 nsew
flabel metal4 1066 758 1092 790 0 FreeSans 320 0 0 0 CTOP
port 6 nsew
<< end >>
