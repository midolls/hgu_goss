magic
tech sky130A
timestamp 1697993263
<< pwell >>
rect 45 243 53 251
<< metal1 >>
rect -44 456 198 459
rect -44 430 -18 456
rect 8 430 14 456
rect 40 430 46 456
rect 72 430 78 456
rect 104 430 110 456
rect 136 430 142 456
rect 168 430 198 456
rect -44 427 198 430
rect -44 404 -17 427
rect -44 378 -43 404
rect -44 372 -17 378
rect -44 346 -43 372
rect -44 340 -17 346
rect -44 314 -43 340
rect -44 308 -17 314
rect -44 282 -43 308
rect -44 276 -17 282
rect -44 250 -43 276
rect -44 244 -17 250
rect -44 218 -43 244
rect -44 212 -17 218
rect -44 186 -43 212
rect -44 180 -17 186
rect -44 154 -43 180
rect -44 148 -17 154
rect -44 122 -43 148
rect -44 116 -17 122
rect -44 90 -43 116
rect -44 84 -17 90
rect -44 58 -43 84
rect -44 46 -17 58
rect 0 32 14 413
rect 28 46 42 427
rect 56 32 70 413
rect 84 46 98 427
rect 112 32 126 413
rect 140 46 154 427
rect 171 404 198 427
rect 197 378 198 404
rect 171 372 198 378
rect 197 346 198 372
rect 171 340 198 346
rect 197 314 198 340
rect 171 308 198 314
rect 197 282 198 308
rect 171 276 198 282
rect 197 250 198 276
rect 171 244 198 250
rect 197 218 198 244
rect 171 212 198 218
rect 197 186 198 212
rect 171 180 198 186
rect 197 154 198 180
rect 171 148 198 154
rect 197 122 198 148
rect 171 116 198 122
rect 197 90 198 116
rect 171 84 198 90
rect 197 58 198 84
rect 171 46 198 58
rect 0 29 154 32
rect 0 3 14 29
rect 40 3 46 29
rect 72 3 78 29
rect 104 3 110 29
rect 136 3 154 29
rect 0 0 154 3
<< via1 >>
rect -18 430 8 456
rect 14 430 40 456
rect 46 430 72 456
rect 78 430 104 456
rect 110 430 136 456
rect 142 430 168 456
rect -43 378 -17 404
rect -43 346 -17 372
rect -43 314 -17 340
rect -43 282 -17 308
rect -43 250 -17 276
rect -43 218 -17 244
rect -43 186 -17 212
rect -43 154 -17 180
rect -43 122 -17 148
rect -43 90 -17 116
rect -43 58 -17 84
rect 171 378 197 404
rect 171 346 197 372
rect 171 314 197 340
rect 171 282 197 308
rect 171 250 197 276
rect 171 218 197 244
rect 171 186 197 212
rect 171 154 197 180
rect 171 122 197 148
rect 171 90 197 116
rect 171 58 197 84
rect 14 3 40 29
rect 46 3 72 29
rect 78 3 104 29
rect 110 3 136 29
<< metal2 >>
rect -44 456 198 459
rect -44 430 -18 456
rect 8 430 14 456
rect 40 430 46 456
rect 72 430 78 456
rect 104 430 110 456
rect 136 430 142 456
rect 168 430 198 456
rect -44 427 198 430
rect -44 404 -17 427
rect -44 378 -43 404
rect -44 372 -17 378
rect -44 346 -43 372
rect -44 340 -17 346
rect -44 314 -43 340
rect -44 308 -17 314
rect -44 282 -43 308
rect -44 276 -17 282
rect -44 250 -43 276
rect -44 244 -17 250
rect -44 218 -43 244
rect -44 212 -17 218
rect -44 186 -43 212
rect -44 180 -17 186
rect -44 154 -43 180
rect -44 148 -17 154
rect -44 122 -43 148
rect -44 116 -17 122
rect -44 90 -43 116
rect -44 84 -17 90
rect -44 58 -43 84
rect -44 46 -17 58
rect 0 46 14 427
rect 28 32 42 413
rect 56 46 70 427
rect 84 32 98 413
rect 112 46 126 427
rect 140 32 154 413
rect 171 404 198 427
rect 197 378 198 404
rect 171 372 198 378
rect 197 346 198 372
rect 171 340 198 346
rect 197 314 198 340
rect 171 308 198 314
rect 197 282 198 308
rect 171 276 198 282
rect 197 250 198 276
rect 171 244 198 250
rect 197 218 198 244
rect 171 212 198 218
rect 197 186 198 212
rect 171 180 198 186
rect 197 154 198 180
rect 171 148 198 154
rect 197 122 198 148
rect 171 116 198 122
rect 197 90 198 116
rect 171 84 198 90
rect 197 58 198 84
rect 171 46 198 58
rect 0 29 154 32
rect 0 3 14 29
rect 40 3 46 29
rect 72 3 78 29
rect 104 3 110 29
rect 136 3 154 29
rect 0 0 154 3
<< labels >>
flabel metal2 s 86 55 97 68 0 FreeSans 100 0 0 0 C0
port 1 nsew
flabel metal2 s 58 390 68 403 0 FreeSans 100 0 0 0 C1
port 2 nsew
flabel pwell s 45 243 53 251 0 FreeSans 100 0 0 0 SUB
port 3 nsew
<< properties >>
string device primitive
string GDS_END 4180
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 148
<< end >>
