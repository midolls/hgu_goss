* NGSPICE file created from hgu_delay_flat.ext - technology: sky130A

.subckt hgu_delay_flat out sample_delay_offset in sample_code0[3] sample_code1[3]
+ sample_code2[3] sample_code3[3] sample_code0[0] sample_code0[1] sample_code0[2]
+ sample_code1[2] sample_code1[1] sample_code1[0] sample_code3[0] sample_code3[1]
+ sample_code2[0] sample_code2[1] sample_code2[2] sample_code3[2] VDD VSS
X0 a_7410_3063# x1.IN a_7322_3201# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1 x2.x5.Y sample_delay_offset VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2 VSS x3.IN a_6749_n1239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3 a_7436_1812# x1.IN a_7364_1812# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 x2.x7.delay_signal sample_code2[0] x2.x5[7].x1.CBOT VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X5 a_6465_2476# x4.x7.delay_signal x1.IN VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X6 a_727_1536# in a_655_1674# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X7 a_655_1122# in a_567_1122# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X8 x1.x7.delay_signal sample_code1[1] x1.x3[1].hgu_cdac_unit_psub_0.CBOT VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X9 a_6058_n161# x3.IN a_5970_n161# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X10 VDD sample_code2[3] sample_code2[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X11 a_12767_n299# x2.IN a_12679_n437# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X12 VSS sample_delay_offset x4.x5.Y VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X13 x4.x7.delay_signal sample_code0[0] x4.x5[7].x1.CBOT VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X14 a_12839_n851# x2.IN a_12767_n713# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X15 x2.x3[1].hgu_cdac_unit_psub_0.CBOT sample_code2[1] x2.x7.delay_signal VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X16 x3.x4[3].hgu_cdac_unit_psub_0.CBOT sample_code3[2] x3.x7.delay_signal VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X17 a_6058_n437# x3.IN a_5970_n437# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X18 a_6084_n2102# x3.IN a_5996_n1964# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X19 a_6465_2135# x1.IN VDD VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_6749_n1036# x3.IN VDD VSS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 x4.x7.delay_signal sample_delay_offset x4.x7.hgu_cdac_unit_psub_0.CBOT VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X22 out x3.x7.delay_signal a_40_n1239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X23 x3.x4[3].hgu_cdac_unit_psub_0.CBOT sample_code3[2] x3.x7.delay_signal VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X24 VDD in a_613_3477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X25 a_7436_1260# x1.IN a_7364_1398# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X26 x1.x7.delay_signal sample_delay_offset x1.x7.hgu_cdac_unit_psub_0.CBOT VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X27 a_12793_n2102# x2.IN a_12705_n2240# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X28 a_6084_n2378# x3.IN a_5996_n2240# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X29 x1.x7.delay_signal sample_code1[0] x1.x5[7].x1.CBOT VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X30 x4.x3[1].hgu_cdac_unit_psub_0.CBOT sample_code0[1] x4.x7.delay_signal VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X31 VDD x2.IN a_13174_2135# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X32 x3.x7.delay_signal sample_code3[0] x3.x5[7].x1.CBOT VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X33 x1.x5[7].x1.CBOT sample_code1[0] x1.x7.delay_signal VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X34 x4.x7.delay_signal sample_code0[1] x4.x3[1].hgu_cdac_unit_psub_0.CBOT VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X35 a_7364_2088# x1.IN a_7276_1950# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X36 a_655_1812# in a_567_1674# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X37 a_6058_n851# x3.IN x3.x7.delay_signal VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X38 a_12839_n299# x2.IN a_12767_n299# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X39 x1.x5[7].x1.CBOT sample_code1[0] x1.x7.delay_signal VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X40 a_727_1260# in a_655_1260# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X41 a_13174_2476# x2.IN VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_12793_n1826# x2.IN x2.x7.delay_signal VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X43 x3.x6.x1.CBOT x3.x5.Y x3.x7.delay_signal VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X44 a_727_1536# in a_655_1536# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X45 x3.x7.delay_signal sample_code3[2] x3.x4[3].hgu_cdac_unit_psub_0.CBOT VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X46 sample_code0[0] sample_code0[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X47 x2.x7.delay_signal sample_code2[0] x2.x5[7].x1.CBOT VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X48 x3.x5[7].x1.CBOT sample_code3[0] x3.x7.delay_signal VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X49 a_6130_n575# x3.IN a_6058_n575# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X50 a_7410_3339# x1.IN a_7322_3477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X51 a_6084_n1826# x3.IN a_5996_n1964# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X52 x3.x7.delay_signal sample_code3[2] x3.x4[3].hgu_cdac_unit_psub_0.CBOT VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X53 sample_code1[0] sample_code1[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X54 a_655_1398# in a_567_1398# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X55 x3.x5.Y sample_delay_offset VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X56 x3.x5[7].x1.CBOT sample_code3[0] x3.x7.delay_signal VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X57 a_701_3063# in a_613_3201# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X58 VDD x1.IN a_6465_2135# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X59 x3.x5[7].x1.CBOT sample_code3[0] x3.x7.delay_signal VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X60 x3.IN x2.x7.delay_signal a_6749_n1036# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X61 a_7364_1674# x1.IN a_7276_1674# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X62 x4.x7.delay_signal sample_code0[2] x4.x4[3].hgu_cdac_unit_psub_0.CBOT VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X63 x1.x7.delay_signal x1.IN a_7364_2088# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X64 x4.x5[7].x1.CBOT sample_code0[0] x4.x7.delay_signal VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X65 a_6465_2476# x1.IN VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X66 a_727_1812# in a_655_1950# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X67 VDD x2.x7.delay_signal a_6749_n1239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X68 a_6749_n1239# x3.IN VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X69 x3.x5[7].x1.CBOT sample_code3[0] x3.x7.delay_signal VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X70 VSS sample_code3[3] sample_code3[0] VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X71 x1.x7.delay_signal sample_code1[2] x1.x4[3].hgu_cdac_unit_psub_0.CBOT VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X72 a_12767_n575# x2.IN a_12679_n713# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X73 x2.x4[3].hgu_cdac_unit_psub_0.CBOT sample_code2[2] x2.x7.delay_signal VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X74 a_6058_n713# x3.IN a_5970_n713# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X75 VSS in a_655_1122# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X76 x1.x5[7].x1.CBOT sample_code1[0] x1.x7.delay_signal VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X77 a_12793_n2378# x2.IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X78 a_13174_2476# x1.x7.delay_signal VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X79 VSS x2.IN a_13174_2476# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X80 x2.x4[3].hgu_cdac_unit_psub_0.CBOT sample_code2[2] x2.x7.delay_signal VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X81 a_6130_n299# x3.IN a_6058_n161# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X82 a_7410_3063# x1.IN a_7322_2925# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X83 x1.x4[3].hgu_cdac_unit_psub_0.CBOT sample_code1[2] x1.x7.delay_signal VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X84 VDD sample_delay_offset x1.x5.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X85 x4.x7.delay_signal sample_code0[0] x4.x5[7].x1.CBOT VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X86 a_7436_1536# x1.IN a_7364_1674# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X87 a_6130_n23# x3.IN a_6058_n23# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X88 a_6130_n575# x3.IN a_6058_n437# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X89 a_7410_3339# x1.IN a_7322_3201# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X90 x2.x7.hgu_cdac_unit_psub_0.CBOT sample_delay_offset x2.x7.delay_signal VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X91 x3.x7.delay_signal sample_code3[0] x3.x2.hgu_cdac_unit_psub_0.CBOT VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.43 as=0.122 ps=1.42 w=0.42 l=0.15
X92 a_655_2088# in a_567_1950# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X93 a_7364_1260# x1.IN a_7276_1122# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X94 a_12839_n23# x2.IN a_12767_n23# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X95 a_12839_n575# x2.IN a_12767_n575# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X96 a_7364_1536# x1.IN a_7276_1398# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X97 VDD out a_40_n1036# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X98 a_6058_n299# x3.IN a_5970_n437# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X99 x1.x7.delay_signal sample_code1[0] x1.x5[7].x1.CBOT VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X100 a_40_n1036# out VDD VSS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X101 x1.x7.delay_signal sample_code1[0] x1.x5[7].x1.CBOT VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X102 a_6130_n23# x3.IN a_6058_115# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X103 a_12793_n2102# x2.IN a_12705_n1964# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X104 x3.x3[1].hgu_cdac_unit_psub_0.CBOT sample_code3[1] x3.x7.delay_signal VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X105 x4.x5[7].x1.CBOT sample_code0[0] x4.x7.delay_signal VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X106 a_727_1812# in a_655_1812# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X107 a_12767_n161# x2.IN a_12679_n161# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X108 a_6465_2476# x4.x7.delay_signal VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X109 VSS x1.IN a_6465_2476# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X110 x3.IN x2.x7.delay_signal a_6749_n1239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X111 a_701_3339# in a_613_3477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X112 a_12839_n23# x2.IN a_12767_115# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X113 x2.x7.delay_signal sample_code2[2] x2.x4[3].hgu_cdac_unit_psub_0.CBOT VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X114 x2.x7.delay_signal sample_code2[0] x2.x2.hgu_cdac_unit_psub_0.CBOT VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.43 as=0.122 ps=1.42 w=0.42 l=0.15
X115 x4.x4[3].hgu_cdac_unit_psub_0.CBOT sample_code0[2] x4.x7.delay_signal VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X116 x2.x5[7].x1.CBOT sample_code2[0] x2.x7.delay_signal VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X117 x3.x7.delay_signal sample_code3[0] x3.x5[7].x1.CBOT VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X118 a_6130_n851# x3.IN a_6058_n851# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X119 sample_code1[0] sample_code1[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X120 x2.x6.x1.CBOT x2.x5.Y x2.x7.delay_signal VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X121 a_12767_n437# x2.IN a_12679_n437# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X122 x1.x7.delay_signal x1.IN a_7322_2925# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X123 a_13174_2135# x1.x7.delay_signal x2.IN VSS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X124 x3.x5.Y sample_delay_offset VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X125 a_655_1674# in a_567_1674# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X126 x2.x5[7].x1.CBOT sample_code2[0] x2.x7.delay_signal VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X127 a_7436_1260# x1.IN a_7364_1260# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X128 x2.x5[7].x1.CBOT sample_code2[0] x2.x7.delay_signal VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X129 x3.x7.delay_signal sample_code3[0] x3.x5[7].x1.CBOT VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X130 a_7364_1950# x1.IN a_7276_1950# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X131 a_12793_n2378# x2.IN a_12705_n2240# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X132 x1.x7.delay_signal x1.x5.Y x1.x6.x1.CBOT VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X133 x1.x2.hgu_cdac_unit_psub_0.CBOT sample_code1[0] x1.x7.delay_signal VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X134 a_7436_1536# x1.IN a_7364_1536# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X135 x2.x5.Y sample_delay_offset VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X136 x2.x5[7].x1.CBOT sample_code2[0] x2.x7.delay_signal VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X137 a_12767_n23# x2.IN a_12679_n161# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X138 a_6084_n2102# x3.IN a_5996_n2240# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X139 x3.x7.delay_signal sample_code3[0] x3.x5[7].x1.CBOT VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X140 x1.x3[1].hgu_cdac_unit_psub_0.CBOT sample_code1[1] x1.x7.delay_signal VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X141 a_6058_n23# x3.IN a_5970_n161# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X142 VDD sample_code3[3] sample_code3[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X143 a_727_1260# in a_655_1398# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X144 a_7364_1122# x1.IN a_7276_1122# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X145 a_12767_n851# x2.IN x2.x7.delay_signal VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X146 a_12839_n299# x2.IN a_12767_n161# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X147 VSS x3.x7.delay_signal a_40_n1036# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X148 x4.x5[7].x1.CBOT sample_code0[0] x4.x7.delay_signal VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X149 VSS sample_code2[3] sample_code2[0] VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X150 x2.x7.delay_signal sample_code2[2] x2.x4[3].hgu_cdac_unit_psub_0.CBOT VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X151 VDD x3.IN a_6749_n1036# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X152 x3.x7.delay_signal sample_code3[1] x3.x3[1].hgu_cdac_unit_psub_0.CBOT VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X153 a_12839_n575# x2.IN a_12767_n437# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X154 VSS sample_delay_offset x1.x5.Y VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X155 a_6084_n1826# x3.IN x3.x7.delay_signal VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X156 x3.x7.hgu_cdac_unit_psub_0.CBOT sample_delay_offset x3.x7.delay_signal VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X157 a_6465_2135# x4.x7.delay_signal x1.IN VSS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X158 a_12767_115# x2.IN VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X159 a_701_3063# in a_613_2925# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X160 x1.x4[3].hgu_cdac_unit_psub_0.CBOT sample_code1[2] x1.x7.delay_signal VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X161 VDD sample_delay_offset x4.x5.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X162 a_6058_115# x3.IN VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X163 a_12793_n1826# x2.IN a_12705_n1964# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X164 a_7436_1812# x1.IN a_7364_1950# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X165 x1.x7.delay_signal sample_code1[2] x1.x4[3].hgu_cdac_unit_psub_0.CBOT VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X166 VSS out a_40_n1239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X167 a_701_3339# in a_613_3201# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X168 x4.x2.hgu_cdac_unit_psub_0.CBOT sample_code0[0] x4.x7.delay_signal VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X169 VSS x2.x7.delay_signal a_6749_n1036# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X170 VDD x1.IN a_7322_3477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X171 x1.x5[7].x1.CBOT sample_code1[0] x1.x7.delay_signal VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X172 a_40_n1239# out VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X173 a_6130_n851# x3.IN a_6058_n713# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X174 a_655_1260# in a_567_1122# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X175 x4.x7.delay_signal sample_code0[0] x4.x5[7].x1.CBOT VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X176 a_13174_2135# x1.x7.delay_signal VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X177 a_655_1536# in a_567_1398# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X178 out x3.x7.delay_signal a_40_n1036# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X179 a_7364_1812# x1.IN a_7276_1674# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X180 VSS x1.IN a_7364_1122# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X181 a_12839_n851# x2.IN a_12767_n851# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X182 a_6058_n575# x3.IN a_5970_n713# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X183 x4.x7.delay_signal x4.x5.Y x4.x6.x1.CBOT VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X184 a_13174_2476# x1.x7.delay_signal x2.IN VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X185 x4.x7.delay_signal in a_655_2088# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X186 VDD x3.x7.delay_signal a_40_n1239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X187 x2.x7.delay_signal sample_code2[1] x2.x3[1].hgu_cdac_unit_psub_0.CBOT VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X188 x1.x7.delay_signal sample_code1[0] x1.x5[7].x1.CBOT VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X189 a_12767_n713# x2.IN a_12679_n713# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X190 x4.x7.delay_signal in a_613_2925# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X191 x4.x7.delay_signal sample_code0[2] x4.x4[3].hgu_cdac_unit_psub_0.CBOT VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X192 a_6130_n299# x3.IN a_6058_n299# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X193 x4.x7.delay_signal sample_code0[0] x4.x5[7].x1.CBOT VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X194 x4.x5[7].x1.CBOT sample_code0[0] x4.x7.delay_signal VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X195 a_13174_2135# x2.IN VDD VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X196 a_6084_n2378# x3.IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X197 sample_code0[0] sample_code0[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X198 a_655_1950# in a_567_1950# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X199 x2.x7.delay_signal sample_code2[0] x2.x5[7].x1.CBOT VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X200 x2.x7.delay_signal sample_code2[0] x2.x5[7].x1.CBOT VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X201 x4.x4[3].hgu_cdac_unit_psub_0.CBOT sample_code0[2] x4.x7.delay_signal VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X202 a_6465_2135# x4.x7.delay_signal VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X203 a_7364_1398# x1.IN a_7276_1398# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
.ends

