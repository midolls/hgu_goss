magic
tech sky130A
magscale 1 2
timestamp 1699632744
<< nwell >>
rect -36 2671 2892 3031
rect 4348 2671 7276 3031
rect -42 1526 16670 1890
rect -38 841 16782 1201
rect -38 152 16782 513
<< pwell >>
rect 3 2431 277 2587
rect 279 2431 801 2613
rect 831 2431 2781 2613
rect 4387 2431 4661 2587
rect 4663 2431 5185 2613
rect 5215 2431 7165 2613
rect 33 2393 67 2431
rect 308 2393 342 2431
rect 860 2393 894 2431
rect 4417 2393 4451 2431
rect 4692 2393 4726 2431
rect 5244 2393 5278 2431
rect 1 1425 187 1471
rect 2075 1425 2261 1471
rect 1 1289 781 1425
rect 1481 1289 2261 1425
rect 2393 1425 2579 1471
rect 4467 1425 4653 1471
rect 2393 1289 3173 1425
rect 3873 1289 4653 1425
rect 4785 1425 4971 1471
rect 6857 1425 7043 1471
rect 4785 1289 5565 1425
rect 6263 1289 7043 1425
rect 7177 1425 7363 1471
rect 9251 1425 9437 1471
rect 7177 1289 7957 1425
rect 8657 1289 9437 1425
rect 9569 1425 9755 1471
rect 11643 1425 11829 1471
rect 9569 1289 10349 1425
rect 11049 1289 11829 1425
rect 11961 1425 12147 1471
rect 14033 1425 14219 1471
rect 11961 1289 12741 1425
rect 13439 1289 14219 1425
rect 14353 1425 14539 1471
rect 16427 1425 16613 1471
rect 14353 1289 15133 1425
rect 15833 1289 16613 1425
rect 84 1251 118 1289
rect 2144 1251 2178 1289
rect 2476 1251 2510 1289
rect 4536 1251 4570 1289
rect 4868 1251 4902 1289
rect 6926 1251 6960 1289
rect 7260 1251 7294 1289
rect 9320 1251 9354 1289
rect 9652 1251 9686 1289
rect 11712 1251 11746 1289
rect 12044 1251 12078 1289
rect 14102 1251 14136 1289
rect 14436 1251 14470 1289
rect 16496 1251 16530 1289
rect 1924 781 2391 783
rect 4316 781 4783 783
rect 6708 781 7175 783
rect 9100 781 9567 783
rect 11492 781 11959 783
rect 13884 781 14351 783
rect 16276 781 16743 783
rect 780 737 1235 781
rect 1557 737 2391 781
rect 3172 737 3627 781
rect 3949 737 4783 781
rect 5564 737 6019 781
rect 6341 737 7175 781
rect 7956 737 8411 781
rect 8733 737 9567 781
rect 10348 737 10803 781
rect 11125 737 11959 781
rect 12740 737 13195 781
rect 13517 737 14351 781
rect 15132 737 15587 781
rect 15909 737 16743 781
rect 1 601 2391 737
rect 2393 601 4783 737
rect 4785 601 7175 737
rect 7177 601 9567 737
rect 9569 601 11959 737
rect 11961 601 14351 737
rect 14353 601 16743 737
rect 29 563 63 601
rect 2421 563 2455 601
rect 4813 563 4847 601
rect 7205 563 7239 601
rect 9597 563 9631 601
rect 11989 563 12023 601
rect 14381 563 14415 601
rect 1 92 468 94
rect 2393 92 2860 94
rect 4785 92 5252 94
rect 7177 92 7644 94
rect 9569 92 10036 94
rect 11961 92 12428 94
rect 14353 92 14820 94
rect 1 48 835 92
rect 1157 48 1612 92
rect 2393 48 3227 92
rect 3549 48 4004 92
rect 4785 48 5619 92
rect 5941 48 6396 92
rect 7177 48 8011 92
rect 8333 48 8788 92
rect 9569 48 10403 92
rect 10725 48 11180 92
rect 11961 48 12795 92
rect 13117 48 13572 92
rect 14353 48 15187 92
rect 15509 48 15964 92
rect 1 -88 2391 48
rect 2393 -88 4783 48
rect 4785 -88 7175 48
rect 7177 -88 9567 48
rect 9569 -88 11959 48
rect 11961 -88 14351 48
rect 14353 -88 16743 48
rect 2329 -126 2363 -88
rect 4721 -126 4755 -88
rect 7113 -126 7147 -88
rect 9505 -126 9539 -88
rect 11897 -126 11931 -88
rect 14289 -126 14323 -88
rect 16681 -126 16715 -88
<< scnmos >>
rect 81 2457 111 2561
rect 169 2457 199 2561
rect 357 2457 387 2587
rect 441 2457 471 2587
rect 525 2457 555 2587
rect 609 2457 639 2587
rect 693 2457 723 2587
rect 909 2457 939 2587
rect 993 2457 1023 2587
rect 1077 2457 1107 2587
rect 1161 2457 1191 2587
rect 1245 2457 1275 2587
rect 1329 2457 1359 2587
rect 1413 2457 1443 2587
rect 1497 2457 1527 2587
rect 1581 2457 1611 2587
rect 1665 2457 1695 2587
rect 1749 2457 1779 2587
rect 1833 2457 1863 2587
rect 1917 2457 1947 2587
rect 2001 2457 2031 2587
rect 2085 2457 2115 2587
rect 2169 2457 2199 2587
rect 2253 2457 2283 2587
rect 2337 2457 2367 2587
rect 2421 2457 2451 2587
rect 2505 2457 2535 2587
rect 2589 2457 2619 2587
rect 2673 2457 2703 2587
rect 4465 2457 4495 2561
rect 4553 2457 4583 2561
rect 4741 2457 4771 2587
rect 4825 2457 4855 2587
rect 4909 2457 4939 2587
rect 4993 2457 5023 2587
rect 5077 2457 5107 2587
rect 5293 2457 5323 2587
rect 5377 2457 5407 2587
rect 5461 2457 5491 2587
rect 5545 2457 5575 2587
rect 5629 2457 5659 2587
rect 5713 2457 5743 2587
rect 5797 2457 5827 2587
rect 5881 2457 5911 2587
rect 5965 2457 5995 2587
rect 6049 2457 6079 2587
rect 6133 2457 6163 2587
rect 6217 2457 6247 2587
rect 6301 2457 6331 2587
rect 6385 2457 6415 2587
rect 6469 2457 6499 2587
rect 6553 2457 6583 2587
rect 6637 2457 6667 2587
rect 6721 2457 6751 2587
rect 6805 2457 6835 2587
rect 6889 2457 6919 2587
rect 6973 2457 7003 2587
rect 7057 2457 7087 2587
rect 79 1315 109 1445
rect 188 1315 218 1399
rect 284 1315 314 1399
rect 409 1315 439 1399
rect 505 1315 535 1399
rect 673 1315 703 1399
rect 1559 1315 1589 1399
rect 1727 1315 1757 1399
rect 1823 1315 1853 1399
rect 1948 1315 1978 1399
rect 2044 1315 2074 1399
rect 2153 1315 2183 1445
rect 2471 1315 2501 1445
rect 2580 1315 2610 1399
rect 2676 1315 2706 1399
rect 2801 1315 2831 1399
rect 2897 1315 2927 1399
rect 3065 1315 3095 1399
rect 3951 1315 3981 1399
rect 4119 1315 4149 1399
rect 4215 1315 4245 1399
rect 4340 1315 4370 1399
rect 4436 1315 4466 1399
rect 4545 1315 4575 1445
rect 4863 1315 4893 1445
rect 4972 1315 5002 1399
rect 5068 1315 5098 1399
rect 5193 1315 5223 1399
rect 5289 1315 5319 1399
rect 5457 1315 5487 1399
rect 6341 1315 6371 1399
rect 6509 1315 6539 1399
rect 6605 1315 6635 1399
rect 6730 1315 6760 1399
rect 6826 1315 6856 1399
rect 6935 1315 6965 1445
rect 7255 1315 7285 1445
rect 7364 1315 7394 1399
rect 7460 1315 7490 1399
rect 7585 1315 7615 1399
rect 7681 1315 7711 1399
rect 7849 1315 7879 1399
rect 8735 1315 8765 1399
rect 8903 1315 8933 1399
rect 8999 1315 9029 1399
rect 9124 1315 9154 1399
rect 9220 1315 9250 1399
rect 9329 1315 9359 1445
rect 9647 1315 9677 1445
rect 9756 1315 9786 1399
rect 9852 1315 9882 1399
rect 9977 1315 10007 1399
rect 10073 1315 10103 1399
rect 10241 1315 10271 1399
rect 11127 1315 11157 1399
rect 11295 1315 11325 1399
rect 11391 1315 11421 1399
rect 11516 1315 11546 1399
rect 11612 1315 11642 1399
rect 11721 1315 11751 1445
rect 12039 1315 12069 1445
rect 12148 1315 12178 1399
rect 12244 1315 12274 1399
rect 12369 1315 12399 1399
rect 12465 1315 12495 1399
rect 12633 1315 12663 1399
rect 13517 1315 13547 1399
rect 13685 1315 13715 1399
rect 13781 1315 13811 1399
rect 13906 1315 13936 1399
rect 14002 1315 14032 1399
rect 14111 1315 14141 1445
rect 14431 1315 14461 1445
rect 14540 1315 14570 1399
rect 14636 1315 14666 1399
rect 14761 1315 14791 1399
rect 14857 1315 14887 1399
rect 15025 1315 15055 1399
rect 15911 1315 15941 1399
rect 16079 1315 16109 1399
rect 16175 1315 16205 1399
rect 16300 1315 16330 1399
rect 16396 1315 16426 1399
rect 16505 1315 16535 1445
rect 79 627 109 711
rect 163 627 193 711
rect 351 627 381 711
rect 446 627 476 699
rect 551 627 581 699
rect 647 627 677 711
rect 761 627 791 711
rect 857 627 887 755
rect 941 627 971 755
rect 1129 627 1159 755
rect 1249 627 1279 699
rect 1333 627 1363 699
rect 1428 627 1458 711
rect 1525 627 1555 711
rect 1633 627 1663 755
rect 1717 627 1747 755
rect 1905 627 1935 711
rect 2000 627 2030 757
rect 2188 627 2218 711
rect 2283 627 2313 757
rect 2471 627 2501 711
rect 2555 627 2585 711
rect 2743 627 2773 711
rect 2838 627 2868 699
rect 2943 627 2973 699
rect 3039 627 3069 711
rect 3153 627 3183 711
rect 3249 627 3279 755
rect 3333 627 3363 755
rect 3521 627 3551 755
rect 3641 627 3671 699
rect 3725 627 3755 699
rect 3820 627 3850 711
rect 3917 627 3947 711
rect 4025 627 4055 755
rect 4109 627 4139 755
rect 4297 627 4327 711
rect 4392 627 4422 757
rect 4580 627 4610 711
rect 4675 627 4705 757
rect 4863 627 4893 711
rect 4947 627 4977 711
rect 5135 627 5165 711
rect 5230 627 5260 699
rect 5335 627 5365 699
rect 5431 627 5461 711
rect 5545 627 5575 711
rect 5641 627 5671 755
rect 5725 627 5755 755
rect 5913 627 5943 755
rect 6033 627 6063 699
rect 6117 627 6147 699
rect 6212 627 6242 711
rect 6309 627 6339 711
rect 6417 627 6447 755
rect 6501 627 6531 755
rect 6689 627 6719 711
rect 6784 627 6814 757
rect 6972 627 7002 711
rect 7067 627 7097 757
rect 7255 627 7285 711
rect 7339 627 7369 711
rect 7527 627 7557 711
rect 7622 627 7652 699
rect 7727 627 7757 699
rect 7823 627 7853 711
rect 7937 627 7967 711
rect 8033 627 8063 755
rect 8117 627 8147 755
rect 8305 627 8335 755
rect 8425 627 8455 699
rect 8509 627 8539 699
rect 8604 627 8634 711
rect 8701 627 8731 711
rect 8809 627 8839 755
rect 8893 627 8923 755
rect 9081 627 9111 711
rect 9176 627 9206 757
rect 9364 627 9394 711
rect 9459 627 9489 757
rect 9647 627 9677 711
rect 9731 627 9761 711
rect 9919 627 9949 711
rect 10014 627 10044 699
rect 10119 627 10149 699
rect 10215 627 10245 711
rect 10329 627 10359 711
rect 10425 627 10455 755
rect 10509 627 10539 755
rect 10697 627 10727 755
rect 10817 627 10847 699
rect 10901 627 10931 699
rect 10996 627 11026 711
rect 11093 627 11123 711
rect 11201 627 11231 755
rect 11285 627 11315 755
rect 11473 627 11503 711
rect 11568 627 11598 757
rect 11756 627 11786 711
rect 11851 627 11881 757
rect 12039 627 12069 711
rect 12123 627 12153 711
rect 12311 627 12341 711
rect 12406 627 12436 699
rect 12511 627 12541 699
rect 12607 627 12637 711
rect 12721 627 12751 711
rect 12817 627 12847 755
rect 12901 627 12931 755
rect 13089 627 13119 755
rect 13209 627 13239 699
rect 13293 627 13323 699
rect 13388 627 13418 711
rect 13485 627 13515 711
rect 13593 627 13623 755
rect 13677 627 13707 755
rect 13865 627 13895 711
rect 13960 627 13990 757
rect 14148 627 14178 711
rect 14243 627 14273 757
rect 14431 627 14461 711
rect 14515 627 14545 711
rect 14703 627 14733 711
rect 14798 627 14828 699
rect 14903 627 14933 699
rect 14999 627 15029 711
rect 15113 627 15143 711
rect 15209 627 15239 755
rect 15293 627 15323 755
rect 15481 627 15511 755
rect 15601 627 15631 699
rect 15685 627 15715 699
rect 15780 627 15810 711
rect 15877 627 15907 711
rect 15985 627 16015 755
rect 16069 627 16099 755
rect 16257 627 16287 711
rect 16352 627 16382 757
rect 16540 627 16570 711
rect 16635 627 16665 757
rect 79 -62 109 68
rect 174 -62 204 22
rect 362 -62 392 68
rect 457 -62 487 22
rect 645 -62 675 66
rect 729 -62 759 66
rect 837 -62 867 22
rect 934 -62 964 22
rect 1029 -62 1059 10
rect 1113 -62 1143 10
rect 1233 -62 1263 66
rect 1421 -62 1451 66
rect 1505 -62 1535 66
rect 1601 -62 1631 22
rect 1715 -62 1745 22
rect 1811 -62 1841 10
rect 1916 -62 1946 10
rect 2011 -62 2041 22
rect 2199 -62 2229 22
rect 2283 -62 2313 22
rect 2471 -62 2501 68
rect 2566 -62 2596 22
rect 2754 -62 2784 68
rect 2849 -62 2879 22
rect 3037 -62 3067 66
rect 3121 -62 3151 66
rect 3229 -62 3259 22
rect 3326 -62 3356 22
rect 3421 -62 3451 10
rect 3505 -62 3535 10
rect 3625 -62 3655 66
rect 3813 -62 3843 66
rect 3897 -62 3927 66
rect 3993 -62 4023 22
rect 4107 -62 4137 22
rect 4203 -62 4233 10
rect 4308 -62 4338 10
rect 4403 -62 4433 22
rect 4591 -62 4621 22
rect 4675 -62 4705 22
rect 4863 -62 4893 68
rect 4958 -62 4988 22
rect 5146 -62 5176 68
rect 5241 -62 5271 22
rect 5429 -62 5459 66
rect 5513 -62 5543 66
rect 5621 -62 5651 22
rect 5718 -62 5748 22
rect 5813 -62 5843 10
rect 5897 -62 5927 10
rect 6017 -62 6047 66
rect 6205 -62 6235 66
rect 6289 -62 6319 66
rect 6385 -62 6415 22
rect 6499 -62 6529 22
rect 6595 -62 6625 10
rect 6700 -62 6730 10
rect 6795 -62 6825 22
rect 6983 -62 7013 22
rect 7067 -62 7097 22
rect 7255 -62 7285 68
rect 7350 -62 7380 22
rect 7538 -62 7568 68
rect 7633 -62 7663 22
rect 7821 -62 7851 66
rect 7905 -62 7935 66
rect 8013 -62 8043 22
rect 8110 -62 8140 22
rect 8205 -62 8235 10
rect 8289 -62 8319 10
rect 8409 -62 8439 66
rect 8597 -62 8627 66
rect 8681 -62 8711 66
rect 8777 -62 8807 22
rect 8891 -62 8921 22
rect 8987 -62 9017 10
rect 9092 -62 9122 10
rect 9187 -62 9217 22
rect 9375 -62 9405 22
rect 9459 -62 9489 22
rect 9647 -62 9677 68
rect 9742 -62 9772 22
rect 9930 -62 9960 68
rect 10025 -62 10055 22
rect 10213 -62 10243 66
rect 10297 -62 10327 66
rect 10405 -62 10435 22
rect 10502 -62 10532 22
rect 10597 -62 10627 10
rect 10681 -62 10711 10
rect 10801 -62 10831 66
rect 10989 -62 11019 66
rect 11073 -62 11103 66
rect 11169 -62 11199 22
rect 11283 -62 11313 22
rect 11379 -62 11409 10
rect 11484 -62 11514 10
rect 11579 -62 11609 22
rect 11767 -62 11797 22
rect 11851 -62 11881 22
rect 12039 -62 12069 68
rect 12134 -62 12164 22
rect 12322 -62 12352 68
rect 12417 -62 12447 22
rect 12605 -62 12635 66
rect 12689 -62 12719 66
rect 12797 -62 12827 22
rect 12894 -62 12924 22
rect 12989 -62 13019 10
rect 13073 -62 13103 10
rect 13193 -62 13223 66
rect 13381 -62 13411 66
rect 13465 -62 13495 66
rect 13561 -62 13591 22
rect 13675 -62 13705 22
rect 13771 -62 13801 10
rect 13876 -62 13906 10
rect 13971 -62 14001 22
rect 14159 -62 14189 22
rect 14243 -62 14273 22
rect 14431 -62 14461 68
rect 14526 -62 14556 22
rect 14714 -62 14744 68
rect 14809 -62 14839 22
rect 14997 -62 15027 66
rect 15081 -62 15111 66
rect 15189 -62 15219 22
rect 15286 -62 15316 22
rect 15381 -62 15411 10
rect 15465 -62 15495 10
rect 15585 -62 15615 66
rect 15773 -62 15803 66
rect 15857 -62 15887 66
rect 15953 -62 15983 22
rect 16067 -62 16097 22
rect 16163 -62 16193 10
rect 16268 -62 16298 10
rect 16363 -62 16393 22
rect 16551 -62 16581 22
rect 16635 -62 16665 22
<< scpmoshvt >>
rect 81 2749 111 2907
rect 169 2749 199 2907
rect 357 2707 387 2907
rect 441 2707 471 2907
rect 525 2707 555 2907
rect 609 2707 639 2907
rect 693 2707 723 2907
rect 909 2707 939 2907
rect 993 2707 1023 2907
rect 1077 2707 1107 2907
rect 1161 2707 1191 2907
rect 1245 2707 1275 2907
rect 1329 2707 1359 2907
rect 1413 2707 1443 2907
rect 1497 2707 1527 2907
rect 1581 2707 1611 2907
rect 1665 2707 1695 2907
rect 1749 2707 1779 2907
rect 1833 2707 1863 2907
rect 1917 2707 1947 2907
rect 2001 2707 2031 2907
rect 2085 2707 2115 2907
rect 2169 2707 2199 2907
rect 2253 2707 2283 2907
rect 2337 2707 2367 2907
rect 2421 2707 2451 2907
rect 2505 2707 2535 2907
rect 2589 2707 2619 2907
rect 2673 2707 2703 2907
rect 4465 2749 4495 2907
rect 4553 2749 4583 2907
rect 4741 2707 4771 2907
rect 4825 2707 4855 2907
rect 4909 2707 4939 2907
rect 4993 2707 5023 2907
rect 5077 2707 5107 2907
rect 5293 2707 5323 2907
rect 5377 2707 5407 2907
rect 5461 2707 5491 2907
rect 5545 2707 5575 2907
rect 5629 2707 5659 2907
rect 5713 2707 5743 2907
rect 5797 2707 5827 2907
rect 5881 2707 5911 2907
rect 5965 2707 5995 2907
rect 6049 2707 6079 2907
rect 6133 2707 6163 2907
rect 6217 2707 6247 2907
rect 6301 2707 6331 2907
rect 6385 2707 6415 2907
rect 6469 2707 6499 2907
rect 6553 2707 6583 2907
rect 6637 2707 6667 2907
rect 6721 2707 6751 2907
rect 6805 2707 6835 2907
rect 6889 2707 6919 2907
rect 6973 2707 7003 2907
rect 7057 2707 7087 2907
rect 79 1565 109 1765
rect 188 1642 218 1726
rect 291 1642 321 1726
rect 505 1642 535 1726
rect 577 1642 607 1726
rect 673 1642 703 1726
rect 1559 1642 1589 1726
rect 1655 1642 1685 1726
rect 1727 1642 1757 1726
rect 1941 1642 1971 1726
rect 2044 1642 2074 1726
rect 2153 1565 2183 1765
rect 2471 1565 2501 1765
rect 2580 1642 2610 1726
rect 2683 1642 2713 1726
rect 2897 1642 2927 1726
rect 2969 1642 2999 1726
rect 3065 1642 3095 1726
rect 3951 1642 3981 1726
rect 4047 1642 4077 1726
rect 4119 1642 4149 1726
rect 4333 1642 4363 1726
rect 4436 1642 4466 1726
rect 4545 1565 4575 1765
rect 4863 1565 4893 1765
rect 4972 1642 5002 1726
rect 5075 1642 5105 1726
rect 5289 1642 5319 1726
rect 5361 1642 5391 1726
rect 5457 1642 5487 1726
rect 6341 1642 6371 1726
rect 6437 1642 6467 1726
rect 6509 1642 6539 1726
rect 6723 1642 6753 1726
rect 6826 1642 6856 1726
rect 6935 1565 6965 1765
rect 7255 1565 7285 1765
rect 7364 1642 7394 1726
rect 7467 1642 7497 1726
rect 7681 1642 7711 1726
rect 7753 1642 7783 1726
rect 7849 1642 7879 1726
rect 8735 1642 8765 1726
rect 8831 1642 8861 1726
rect 8903 1642 8933 1726
rect 9117 1642 9147 1726
rect 9220 1642 9250 1726
rect 9329 1565 9359 1765
rect 9647 1565 9677 1765
rect 9756 1642 9786 1726
rect 9859 1642 9889 1726
rect 10073 1642 10103 1726
rect 10145 1642 10175 1726
rect 10241 1642 10271 1726
rect 11127 1642 11157 1726
rect 11223 1642 11253 1726
rect 11295 1642 11325 1726
rect 11509 1642 11539 1726
rect 11612 1642 11642 1726
rect 11721 1565 11751 1765
rect 12039 1565 12069 1765
rect 12148 1642 12178 1726
rect 12251 1642 12281 1726
rect 12465 1642 12495 1726
rect 12537 1642 12567 1726
rect 12633 1642 12663 1726
rect 13517 1642 13547 1726
rect 13613 1642 13643 1726
rect 13685 1642 13715 1726
rect 13899 1642 13929 1726
rect 14002 1642 14032 1726
rect 14111 1565 14141 1765
rect 14431 1565 14461 1765
rect 14540 1642 14570 1726
rect 14643 1642 14673 1726
rect 14857 1642 14887 1726
rect 14929 1642 14959 1726
rect 15025 1642 15055 1726
rect 15911 1642 15941 1726
rect 16007 1642 16037 1726
rect 16079 1642 16109 1726
rect 16293 1642 16323 1726
rect 16396 1642 16426 1726
rect 16505 1565 16535 1765
rect 79 943 109 1071
rect 163 943 193 1071
rect 351 993 381 1077
rect 443 993 473 1077
rect 527 993 557 1077
rect 647 993 677 1077
rect 753 993 783 1077
rect 861 909 891 1077
rect 945 909 975 1077
rect 1082 909 1112 1077
rect 1226 993 1256 1077
rect 1310 993 1340 1077
rect 1415 993 1445 1077
rect 1536 993 1566 1077
rect 1642 909 1672 1077
rect 1714 909 1744 1077
rect 1903 881 1933 1009
rect 2000 877 2030 1077
rect 2188 933 2218 1061
rect 2283 877 2313 1077
rect 2471 943 2501 1071
rect 2555 943 2585 1071
rect 2743 993 2773 1077
rect 2835 993 2865 1077
rect 2919 993 2949 1077
rect 3039 993 3069 1077
rect 3145 993 3175 1077
rect 3253 909 3283 1077
rect 3337 909 3367 1077
rect 3474 909 3504 1077
rect 3618 993 3648 1077
rect 3702 993 3732 1077
rect 3807 993 3837 1077
rect 3928 993 3958 1077
rect 4034 909 4064 1077
rect 4106 909 4136 1077
rect 4295 881 4325 1009
rect 4392 877 4422 1077
rect 4580 933 4610 1061
rect 4675 877 4705 1077
rect 4863 943 4893 1071
rect 4947 943 4977 1071
rect 5135 993 5165 1077
rect 5227 993 5257 1077
rect 5311 993 5341 1077
rect 5431 993 5461 1077
rect 5537 993 5567 1077
rect 5645 909 5675 1077
rect 5729 909 5759 1077
rect 5866 909 5896 1077
rect 6010 993 6040 1077
rect 6094 993 6124 1077
rect 6199 993 6229 1077
rect 6320 993 6350 1077
rect 6426 909 6456 1077
rect 6498 909 6528 1077
rect 6687 881 6717 1009
rect 6784 877 6814 1077
rect 6972 933 7002 1061
rect 7067 877 7097 1077
rect 7255 943 7285 1071
rect 7339 943 7369 1071
rect 7527 993 7557 1077
rect 7619 993 7649 1077
rect 7703 993 7733 1077
rect 7823 993 7853 1077
rect 7929 993 7959 1077
rect 8037 909 8067 1077
rect 8121 909 8151 1077
rect 8258 909 8288 1077
rect 8402 993 8432 1077
rect 8486 993 8516 1077
rect 8591 993 8621 1077
rect 8712 993 8742 1077
rect 8818 909 8848 1077
rect 8890 909 8920 1077
rect 9079 881 9109 1009
rect 9176 877 9206 1077
rect 9364 933 9394 1061
rect 9459 877 9489 1077
rect 9647 943 9677 1071
rect 9731 943 9761 1071
rect 9919 993 9949 1077
rect 10011 993 10041 1077
rect 10095 993 10125 1077
rect 10215 993 10245 1077
rect 10321 993 10351 1077
rect 10429 909 10459 1077
rect 10513 909 10543 1077
rect 10650 909 10680 1077
rect 10794 993 10824 1077
rect 10878 993 10908 1077
rect 10983 993 11013 1077
rect 11104 993 11134 1077
rect 11210 909 11240 1077
rect 11282 909 11312 1077
rect 11471 881 11501 1009
rect 11568 877 11598 1077
rect 11756 933 11786 1061
rect 11851 877 11881 1077
rect 12039 943 12069 1071
rect 12123 943 12153 1071
rect 12311 993 12341 1077
rect 12403 993 12433 1077
rect 12487 993 12517 1077
rect 12607 993 12637 1077
rect 12713 993 12743 1077
rect 12821 909 12851 1077
rect 12905 909 12935 1077
rect 13042 909 13072 1077
rect 13186 993 13216 1077
rect 13270 993 13300 1077
rect 13375 993 13405 1077
rect 13496 993 13526 1077
rect 13602 909 13632 1077
rect 13674 909 13704 1077
rect 13863 881 13893 1009
rect 13960 877 13990 1077
rect 14148 933 14178 1061
rect 14243 877 14273 1077
rect 14431 943 14461 1071
rect 14515 943 14545 1071
rect 14703 993 14733 1077
rect 14795 993 14825 1077
rect 14879 993 14909 1077
rect 14999 993 15029 1077
rect 15105 993 15135 1077
rect 15213 909 15243 1077
rect 15297 909 15327 1077
rect 15434 909 15464 1077
rect 15578 993 15608 1077
rect 15662 993 15692 1077
rect 15767 993 15797 1077
rect 15888 993 15918 1077
rect 15994 909 16024 1077
rect 16066 909 16096 1077
rect 16255 881 16285 1009
rect 16352 877 16382 1077
rect 16540 933 16570 1061
rect 16635 877 16665 1077
rect 79 188 109 388
rect 174 244 204 372
rect 362 188 392 388
rect 459 192 489 320
rect 648 220 678 388
rect 720 220 750 388
rect 826 304 856 388
rect 947 304 977 388
rect 1052 304 1082 388
rect 1136 304 1166 388
rect 1280 220 1310 388
rect 1417 220 1447 388
rect 1501 220 1531 388
rect 1609 304 1639 388
rect 1715 304 1745 388
rect 1835 304 1865 388
rect 1919 304 1949 388
rect 2011 304 2041 388
rect 2199 254 2229 382
rect 2283 254 2313 382
rect 2471 188 2501 388
rect 2566 244 2596 372
rect 2754 188 2784 388
rect 2851 192 2881 320
rect 3040 220 3070 388
rect 3112 220 3142 388
rect 3218 304 3248 388
rect 3339 304 3369 388
rect 3444 304 3474 388
rect 3528 304 3558 388
rect 3672 220 3702 388
rect 3809 220 3839 388
rect 3893 220 3923 388
rect 4001 304 4031 388
rect 4107 304 4137 388
rect 4227 304 4257 388
rect 4311 304 4341 388
rect 4403 304 4433 388
rect 4591 254 4621 382
rect 4675 254 4705 382
rect 4863 188 4893 388
rect 4958 244 4988 372
rect 5146 188 5176 388
rect 5243 192 5273 320
rect 5432 220 5462 388
rect 5504 220 5534 388
rect 5610 304 5640 388
rect 5731 304 5761 388
rect 5836 304 5866 388
rect 5920 304 5950 388
rect 6064 220 6094 388
rect 6201 220 6231 388
rect 6285 220 6315 388
rect 6393 304 6423 388
rect 6499 304 6529 388
rect 6619 304 6649 388
rect 6703 304 6733 388
rect 6795 304 6825 388
rect 6983 254 7013 382
rect 7067 254 7097 382
rect 7255 188 7285 388
rect 7350 244 7380 372
rect 7538 188 7568 388
rect 7635 192 7665 320
rect 7824 220 7854 388
rect 7896 220 7926 388
rect 8002 304 8032 388
rect 8123 304 8153 388
rect 8228 304 8258 388
rect 8312 304 8342 388
rect 8456 220 8486 388
rect 8593 220 8623 388
rect 8677 220 8707 388
rect 8785 304 8815 388
rect 8891 304 8921 388
rect 9011 304 9041 388
rect 9095 304 9125 388
rect 9187 304 9217 388
rect 9375 254 9405 382
rect 9459 254 9489 382
rect 9647 188 9677 388
rect 9742 244 9772 372
rect 9930 188 9960 388
rect 10027 192 10057 320
rect 10216 220 10246 388
rect 10288 220 10318 388
rect 10394 304 10424 388
rect 10515 304 10545 388
rect 10620 304 10650 388
rect 10704 304 10734 388
rect 10848 220 10878 388
rect 10985 220 11015 388
rect 11069 220 11099 388
rect 11177 304 11207 388
rect 11283 304 11313 388
rect 11403 304 11433 388
rect 11487 304 11517 388
rect 11579 304 11609 388
rect 11767 254 11797 382
rect 11851 254 11881 382
rect 12039 188 12069 388
rect 12134 244 12164 372
rect 12322 188 12352 388
rect 12419 192 12449 320
rect 12608 220 12638 388
rect 12680 220 12710 388
rect 12786 304 12816 388
rect 12907 304 12937 388
rect 13012 304 13042 388
rect 13096 304 13126 388
rect 13240 220 13270 388
rect 13377 220 13407 388
rect 13461 220 13491 388
rect 13569 304 13599 388
rect 13675 304 13705 388
rect 13795 304 13825 388
rect 13879 304 13909 388
rect 13971 304 14001 388
rect 14159 254 14189 382
rect 14243 254 14273 382
rect 14431 188 14461 388
rect 14526 244 14556 372
rect 14714 188 14744 388
rect 14811 192 14841 320
rect 15000 220 15030 388
rect 15072 220 15102 388
rect 15178 304 15208 388
rect 15299 304 15329 388
rect 15404 304 15434 388
rect 15488 304 15518 388
rect 15632 220 15662 388
rect 15769 220 15799 388
rect 15853 220 15883 388
rect 15961 304 15991 388
rect 16067 304 16097 388
rect 16187 304 16217 388
rect 16271 304 16301 388
rect 16363 304 16393 388
rect 16551 254 16581 382
rect 16635 254 16665 382
<< ndiff >>
rect 29 2516 81 2561
rect 29 2482 37 2516
rect 71 2482 81 2516
rect 29 2457 81 2482
rect 111 2503 169 2561
rect 111 2469 123 2503
rect 157 2469 169 2503
rect 111 2457 169 2469
rect 199 2533 251 2561
rect 199 2499 209 2533
rect 243 2499 251 2533
rect 199 2457 251 2499
rect 305 2539 357 2587
rect 305 2505 313 2539
rect 347 2505 357 2539
rect 305 2457 357 2505
rect 387 2507 441 2587
rect 387 2473 397 2507
rect 431 2473 441 2507
rect 387 2457 441 2473
rect 471 2539 525 2587
rect 471 2505 481 2539
rect 515 2505 525 2539
rect 471 2457 525 2505
rect 555 2507 609 2587
rect 555 2473 565 2507
rect 599 2473 609 2507
rect 555 2457 609 2473
rect 639 2539 693 2587
rect 639 2505 649 2539
rect 683 2505 693 2539
rect 639 2457 693 2505
rect 723 2571 775 2587
rect 723 2537 733 2571
rect 767 2537 775 2571
rect 723 2503 775 2537
rect 723 2469 733 2503
rect 767 2469 775 2503
rect 723 2457 775 2469
rect 857 2575 909 2587
rect 857 2541 865 2575
rect 899 2541 909 2575
rect 857 2507 909 2541
rect 857 2473 865 2507
rect 899 2473 909 2507
rect 857 2457 909 2473
rect 939 2575 993 2587
rect 939 2541 949 2575
rect 983 2541 993 2575
rect 939 2507 993 2541
rect 939 2473 949 2507
rect 983 2473 993 2507
rect 939 2457 993 2473
rect 1023 2507 1077 2587
rect 1023 2473 1033 2507
rect 1067 2473 1077 2507
rect 1023 2457 1077 2473
rect 1107 2575 1161 2587
rect 1107 2541 1117 2575
rect 1151 2541 1161 2575
rect 1107 2507 1161 2541
rect 1107 2473 1117 2507
rect 1151 2473 1161 2507
rect 1107 2457 1161 2473
rect 1191 2507 1245 2587
rect 1191 2473 1201 2507
rect 1235 2473 1245 2507
rect 1191 2457 1245 2473
rect 1275 2575 1329 2587
rect 1275 2541 1285 2575
rect 1319 2541 1329 2575
rect 1275 2507 1329 2541
rect 1275 2473 1285 2507
rect 1319 2473 1329 2507
rect 1275 2457 1329 2473
rect 1359 2507 1413 2587
rect 1359 2473 1369 2507
rect 1403 2473 1413 2507
rect 1359 2457 1413 2473
rect 1443 2575 1497 2587
rect 1443 2541 1453 2575
rect 1487 2541 1497 2575
rect 1443 2507 1497 2541
rect 1443 2473 1453 2507
rect 1487 2473 1497 2507
rect 1443 2457 1497 2473
rect 1527 2507 1581 2587
rect 1527 2473 1537 2507
rect 1571 2473 1581 2507
rect 1527 2457 1581 2473
rect 1611 2575 1665 2587
rect 1611 2541 1621 2575
rect 1655 2541 1665 2575
rect 1611 2507 1665 2541
rect 1611 2473 1621 2507
rect 1655 2473 1665 2507
rect 1611 2457 1665 2473
rect 1695 2507 1749 2587
rect 1695 2473 1705 2507
rect 1739 2473 1749 2507
rect 1695 2457 1749 2473
rect 1779 2575 1833 2587
rect 1779 2541 1789 2575
rect 1823 2541 1833 2575
rect 1779 2507 1833 2541
rect 1779 2473 1789 2507
rect 1823 2473 1833 2507
rect 1779 2457 1833 2473
rect 1863 2507 1917 2587
rect 1863 2473 1873 2507
rect 1907 2473 1917 2507
rect 1863 2457 1917 2473
rect 1947 2575 2001 2587
rect 1947 2541 1957 2575
rect 1991 2541 2001 2575
rect 1947 2507 2001 2541
rect 1947 2473 1957 2507
rect 1991 2473 2001 2507
rect 1947 2457 2001 2473
rect 2031 2507 2085 2587
rect 2031 2473 2041 2507
rect 2075 2473 2085 2507
rect 2031 2457 2085 2473
rect 2115 2575 2169 2587
rect 2115 2541 2125 2575
rect 2159 2541 2169 2575
rect 2115 2507 2169 2541
rect 2115 2473 2125 2507
rect 2159 2473 2169 2507
rect 2115 2457 2169 2473
rect 2199 2507 2253 2587
rect 2199 2473 2209 2507
rect 2243 2473 2253 2507
rect 2199 2457 2253 2473
rect 2283 2575 2337 2587
rect 2283 2541 2293 2575
rect 2327 2541 2337 2575
rect 2283 2507 2337 2541
rect 2283 2473 2293 2507
rect 2327 2473 2337 2507
rect 2283 2457 2337 2473
rect 2367 2507 2421 2587
rect 2367 2473 2377 2507
rect 2411 2473 2421 2507
rect 2367 2457 2421 2473
rect 2451 2575 2505 2587
rect 2451 2541 2461 2575
rect 2495 2541 2505 2575
rect 2451 2507 2505 2541
rect 2451 2473 2461 2507
rect 2495 2473 2505 2507
rect 2451 2457 2505 2473
rect 2535 2507 2589 2587
rect 2535 2473 2545 2507
rect 2579 2473 2589 2507
rect 2535 2457 2589 2473
rect 2619 2575 2673 2587
rect 2619 2541 2629 2575
rect 2663 2541 2673 2575
rect 2619 2507 2673 2541
rect 2619 2473 2629 2507
rect 2663 2473 2673 2507
rect 2619 2457 2673 2473
rect 2703 2507 2755 2587
rect 2703 2473 2713 2507
rect 2747 2473 2755 2507
rect 2703 2457 2755 2473
rect 4413 2516 4465 2561
rect 4413 2482 4421 2516
rect 4455 2482 4465 2516
rect 4413 2457 4465 2482
rect 4495 2503 4553 2561
rect 4495 2469 4507 2503
rect 4541 2469 4553 2503
rect 4495 2457 4553 2469
rect 4583 2533 4635 2561
rect 4583 2499 4593 2533
rect 4627 2499 4635 2533
rect 4583 2457 4635 2499
rect 4689 2539 4741 2587
rect 4689 2505 4697 2539
rect 4731 2505 4741 2539
rect 4689 2457 4741 2505
rect 4771 2507 4825 2587
rect 4771 2473 4781 2507
rect 4815 2473 4825 2507
rect 4771 2457 4825 2473
rect 4855 2539 4909 2587
rect 4855 2505 4865 2539
rect 4899 2505 4909 2539
rect 4855 2457 4909 2505
rect 4939 2507 4993 2587
rect 4939 2473 4949 2507
rect 4983 2473 4993 2507
rect 4939 2457 4993 2473
rect 5023 2539 5077 2587
rect 5023 2505 5033 2539
rect 5067 2505 5077 2539
rect 5023 2457 5077 2505
rect 5107 2571 5159 2587
rect 5107 2537 5117 2571
rect 5151 2537 5159 2571
rect 5107 2503 5159 2537
rect 5107 2469 5117 2503
rect 5151 2469 5159 2503
rect 5107 2457 5159 2469
rect 5241 2575 5293 2587
rect 5241 2541 5249 2575
rect 5283 2541 5293 2575
rect 5241 2507 5293 2541
rect 5241 2473 5249 2507
rect 5283 2473 5293 2507
rect 5241 2457 5293 2473
rect 5323 2575 5377 2587
rect 5323 2541 5333 2575
rect 5367 2541 5377 2575
rect 5323 2507 5377 2541
rect 5323 2473 5333 2507
rect 5367 2473 5377 2507
rect 5323 2457 5377 2473
rect 5407 2507 5461 2587
rect 5407 2473 5417 2507
rect 5451 2473 5461 2507
rect 5407 2457 5461 2473
rect 5491 2575 5545 2587
rect 5491 2541 5501 2575
rect 5535 2541 5545 2575
rect 5491 2507 5545 2541
rect 5491 2473 5501 2507
rect 5535 2473 5545 2507
rect 5491 2457 5545 2473
rect 5575 2507 5629 2587
rect 5575 2473 5585 2507
rect 5619 2473 5629 2507
rect 5575 2457 5629 2473
rect 5659 2575 5713 2587
rect 5659 2541 5669 2575
rect 5703 2541 5713 2575
rect 5659 2507 5713 2541
rect 5659 2473 5669 2507
rect 5703 2473 5713 2507
rect 5659 2457 5713 2473
rect 5743 2507 5797 2587
rect 5743 2473 5753 2507
rect 5787 2473 5797 2507
rect 5743 2457 5797 2473
rect 5827 2575 5881 2587
rect 5827 2541 5837 2575
rect 5871 2541 5881 2575
rect 5827 2507 5881 2541
rect 5827 2473 5837 2507
rect 5871 2473 5881 2507
rect 5827 2457 5881 2473
rect 5911 2507 5965 2587
rect 5911 2473 5921 2507
rect 5955 2473 5965 2507
rect 5911 2457 5965 2473
rect 5995 2575 6049 2587
rect 5995 2541 6005 2575
rect 6039 2541 6049 2575
rect 5995 2507 6049 2541
rect 5995 2473 6005 2507
rect 6039 2473 6049 2507
rect 5995 2457 6049 2473
rect 6079 2507 6133 2587
rect 6079 2473 6089 2507
rect 6123 2473 6133 2507
rect 6079 2457 6133 2473
rect 6163 2575 6217 2587
rect 6163 2541 6173 2575
rect 6207 2541 6217 2575
rect 6163 2507 6217 2541
rect 6163 2473 6173 2507
rect 6207 2473 6217 2507
rect 6163 2457 6217 2473
rect 6247 2507 6301 2587
rect 6247 2473 6257 2507
rect 6291 2473 6301 2507
rect 6247 2457 6301 2473
rect 6331 2575 6385 2587
rect 6331 2541 6341 2575
rect 6375 2541 6385 2575
rect 6331 2507 6385 2541
rect 6331 2473 6341 2507
rect 6375 2473 6385 2507
rect 6331 2457 6385 2473
rect 6415 2507 6469 2587
rect 6415 2473 6425 2507
rect 6459 2473 6469 2507
rect 6415 2457 6469 2473
rect 6499 2575 6553 2587
rect 6499 2541 6509 2575
rect 6543 2541 6553 2575
rect 6499 2507 6553 2541
rect 6499 2473 6509 2507
rect 6543 2473 6553 2507
rect 6499 2457 6553 2473
rect 6583 2507 6637 2587
rect 6583 2473 6593 2507
rect 6627 2473 6637 2507
rect 6583 2457 6637 2473
rect 6667 2575 6721 2587
rect 6667 2541 6677 2575
rect 6711 2541 6721 2575
rect 6667 2507 6721 2541
rect 6667 2473 6677 2507
rect 6711 2473 6721 2507
rect 6667 2457 6721 2473
rect 6751 2507 6805 2587
rect 6751 2473 6761 2507
rect 6795 2473 6805 2507
rect 6751 2457 6805 2473
rect 6835 2575 6889 2587
rect 6835 2541 6845 2575
rect 6879 2541 6889 2575
rect 6835 2507 6889 2541
rect 6835 2473 6845 2507
rect 6879 2473 6889 2507
rect 6835 2457 6889 2473
rect 6919 2507 6973 2587
rect 6919 2473 6929 2507
rect 6963 2473 6973 2507
rect 6919 2457 6973 2473
rect 7003 2575 7057 2587
rect 7003 2541 7013 2575
rect 7047 2541 7057 2575
rect 7003 2507 7057 2541
rect 7003 2473 7013 2507
rect 7047 2473 7057 2507
rect 7003 2457 7057 2473
rect 7087 2507 7139 2587
rect 7087 2473 7097 2507
rect 7131 2473 7139 2507
rect 7087 2457 7139 2473
rect 27 1380 79 1445
rect 27 1346 35 1380
rect 69 1346 79 1380
rect 27 1315 79 1346
rect 109 1399 161 1445
rect 2101 1399 2153 1445
rect 109 1361 188 1399
rect 109 1327 119 1361
rect 153 1327 188 1361
rect 109 1315 188 1327
rect 218 1315 284 1399
rect 314 1376 409 1399
rect 314 1342 326 1376
rect 360 1342 409 1376
rect 314 1315 409 1342
rect 439 1315 505 1399
rect 535 1376 673 1399
rect 535 1342 561 1376
rect 595 1342 629 1376
rect 663 1342 673 1376
rect 535 1315 673 1342
rect 703 1376 755 1399
rect 703 1342 713 1376
rect 747 1342 755 1376
rect 703 1315 755 1342
rect 1507 1376 1559 1399
rect 1507 1342 1515 1376
rect 1549 1342 1559 1376
rect 1507 1315 1559 1342
rect 1589 1376 1727 1399
rect 1589 1342 1599 1376
rect 1633 1342 1667 1376
rect 1701 1342 1727 1376
rect 1589 1315 1727 1342
rect 1757 1315 1823 1399
rect 1853 1376 1948 1399
rect 1853 1342 1902 1376
rect 1936 1342 1948 1376
rect 1853 1315 1948 1342
rect 1978 1315 2044 1399
rect 2074 1361 2153 1399
rect 2074 1327 2109 1361
rect 2143 1327 2153 1361
rect 2074 1315 2153 1327
rect 2183 1380 2235 1445
rect 2183 1346 2193 1380
rect 2227 1346 2235 1380
rect 2183 1315 2235 1346
rect 2419 1380 2471 1445
rect 2419 1346 2427 1380
rect 2461 1346 2471 1380
rect 2419 1315 2471 1346
rect 2501 1399 2553 1445
rect 4493 1399 4545 1445
rect 2501 1361 2580 1399
rect 2501 1327 2511 1361
rect 2545 1327 2580 1361
rect 2501 1315 2580 1327
rect 2610 1315 2676 1399
rect 2706 1376 2801 1399
rect 2706 1342 2718 1376
rect 2752 1342 2801 1376
rect 2706 1315 2801 1342
rect 2831 1315 2897 1399
rect 2927 1376 3065 1399
rect 2927 1342 2953 1376
rect 2987 1342 3021 1376
rect 3055 1342 3065 1376
rect 2927 1315 3065 1342
rect 3095 1376 3147 1399
rect 3095 1342 3105 1376
rect 3139 1342 3147 1376
rect 3095 1315 3147 1342
rect 3899 1376 3951 1399
rect 3899 1342 3907 1376
rect 3941 1342 3951 1376
rect 3899 1315 3951 1342
rect 3981 1376 4119 1399
rect 3981 1342 3991 1376
rect 4025 1342 4059 1376
rect 4093 1342 4119 1376
rect 3981 1315 4119 1342
rect 4149 1315 4215 1399
rect 4245 1376 4340 1399
rect 4245 1342 4294 1376
rect 4328 1342 4340 1376
rect 4245 1315 4340 1342
rect 4370 1315 4436 1399
rect 4466 1361 4545 1399
rect 4466 1327 4501 1361
rect 4535 1327 4545 1361
rect 4466 1315 4545 1327
rect 4575 1380 4627 1445
rect 4575 1346 4585 1380
rect 4619 1346 4627 1380
rect 4575 1315 4627 1346
rect 4811 1380 4863 1445
rect 4811 1346 4819 1380
rect 4853 1346 4863 1380
rect 4811 1315 4863 1346
rect 4893 1399 4945 1445
rect 6883 1399 6935 1445
rect 4893 1361 4972 1399
rect 4893 1327 4903 1361
rect 4937 1327 4972 1361
rect 4893 1315 4972 1327
rect 5002 1315 5068 1399
rect 5098 1376 5193 1399
rect 5098 1342 5110 1376
rect 5144 1342 5193 1376
rect 5098 1315 5193 1342
rect 5223 1315 5289 1399
rect 5319 1376 5457 1399
rect 5319 1342 5345 1376
rect 5379 1342 5413 1376
rect 5447 1342 5457 1376
rect 5319 1315 5457 1342
rect 5487 1376 5539 1399
rect 5487 1342 5497 1376
rect 5531 1342 5539 1376
rect 5487 1315 5539 1342
rect 6289 1376 6341 1399
rect 6289 1342 6297 1376
rect 6331 1342 6341 1376
rect 6289 1315 6341 1342
rect 6371 1376 6509 1399
rect 6371 1342 6381 1376
rect 6415 1342 6449 1376
rect 6483 1342 6509 1376
rect 6371 1315 6509 1342
rect 6539 1315 6605 1399
rect 6635 1376 6730 1399
rect 6635 1342 6684 1376
rect 6718 1342 6730 1376
rect 6635 1315 6730 1342
rect 6760 1315 6826 1399
rect 6856 1361 6935 1399
rect 6856 1327 6891 1361
rect 6925 1327 6935 1361
rect 6856 1315 6935 1327
rect 6965 1380 7017 1445
rect 6965 1346 6975 1380
rect 7009 1346 7017 1380
rect 6965 1315 7017 1346
rect 7203 1380 7255 1445
rect 7203 1346 7211 1380
rect 7245 1346 7255 1380
rect 7203 1315 7255 1346
rect 7285 1399 7337 1445
rect 9277 1399 9329 1445
rect 7285 1361 7364 1399
rect 7285 1327 7295 1361
rect 7329 1327 7364 1361
rect 7285 1315 7364 1327
rect 7394 1315 7460 1399
rect 7490 1376 7585 1399
rect 7490 1342 7502 1376
rect 7536 1342 7585 1376
rect 7490 1315 7585 1342
rect 7615 1315 7681 1399
rect 7711 1376 7849 1399
rect 7711 1342 7737 1376
rect 7771 1342 7805 1376
rect 7839 1342 7849 1376
rect 7711 1315 7849 1342
rect 7879 1376 7931 1399
rect 7879 1342 7889 1376
rect 7923 1342 7931 1376
rect 7879 1315 7931 1342
rect 8683 1376 8735 1399
rect 8683 1342 8691 1376
rect 8725 1342 8735 1376
rect 8683 1315 8735 1342
rect 8765 1376 8903 1399
rect 8765 1342 8775 1376
rect 8809 1342 8843 1376
rect 8877 1342 8903 1376
rect 8765 1315 8903 1342
rect 8933 1315 8999 1399
rect 9029 1376 9124 1399
rect 9029 1342 9078 1376
rect 9112 1342 9124 1376
rect 9029 1315 9124 1342
rect 9154 1315 9220 1399
rect 9250 1361 9329 1399
rect 9250 1327 9285 1361
rect 9319 1327 9329 1361
rect 9250 1315 9329 1327
rect 9359 1380 9411 1445
rect 9359 1346 9369 1380
rect 9403 1346 9411 1380
rect 9359 1315 9411 1346
rect 9595 1380 9647 1445
rect 9595 1346 9603 1380
rect 9637 1346 9647 1380
rect 9595 1315 9647 1346
rect 9677 1399 9729 1445
rect 11669 1399 11721 1445
rect 9677 1361 9756 1399
rect 9677 1327 9687 1361
rect 9721 1327 9756 1361
rect 9677 1315 9756 1327
rect 9786 1315 9852 1399
rect 9882 1376 9977 1399
rect 9882 1342 9894 1376
rect 9928 1342 9977 1376
rect 9882 1315 9977 1342
rect 10007 1315 10073 1399
rect 10103 1376 10241 1399
rect 10103 1342 10129 1376
rect 10163 1342 10197 1376
rect 10231 1342 10241 1376
rect 10103 1315 10241 1342
rect 10271 1376 10323 1399
rect 10271 1342 10281 1376
rect 10315 1342 10323 1376
rect 10271 1315 10323 1342
rect 11075 1376 11127 1399
rect 11075 1342 11083 1376
rect 11117 1342 11127 1376
rect 11075 1315 11127 1342
rect 11157 1376 11295 1399
rect 11157 1342 11167 1376
rect 11201 1342 11235 1376
rect 11269 1342 11295 1376
rect 11157 1315 11295 1342
rect 11325 1315 11391 1399
rect 11421 1376 11516 1399
rect 11421 1342 11470 1376
rect 11504 1342 11516 1376
rect 11421 1315 11516 1342
rect 11546 1315 11612 1399
rect 11642 1361 11721 1399
rect 11642 1327 11677 1361
rect 11711 1327 11721 1361
rect 11642 1315 11721 1327
rect 11751 1380 11803 1445
rect 11751 1346 11761 1380
rect 11795 1346 11803 1380
rect 11751 1315 11803 1346
rect 11987 1380 12039 1445
rect 11987 1346 11995 1380
rect 12029 1346 12039 1380
rect 11987 1315 12039 1346
rect 12069 1399 12121 1445
rect 14059 1399 14111 1445
rect 12069 1361 12148 1399
rect 12069 1327 12079 1361
rect 12113 1327 12148 1361
rect 12069 1315 12148 1327
rect 12178 1315 12244 1399
rect 12274 1376 12369 1399
rect 12274 1342 12286 1376
rect 12320 1342 12369 1376
rect 12274 1315 12369 1342
rect 12399 1315 12465 1399
rect 12495 1376 12633 1399
rect 12495 1342 12521 1376
rect 12555 1342 12589 1376
rect 12623 1342 12633 1376
rect 12495 1315 12633 1342
rect 12663 1376 12715 1399
rect 12663 1342 12673 1376
rect 12707 1342 12715 1376
rect 12663 1315 12715 1342
rect 13465 1376 13517 1399
rect 13465 1342 13473 1376
rect 13507 1342 13517 1376
rect 13465 1315 13517 1342
rect 13547 1376 13685 1399
rect 13547 1342 13557 1376
rect 13591 1342 13625 1376
rect 13659 1342 13685 1376
rect 13547 1315 13685 1342
rect 13715 1315 13781 1399
rect 13811 1376 13906 1399
rect 13811 1342 13860 1376
rect 13894 1342 13906 1376
rect 13811 1315 13906 1342
rect 13936 1315 14002 1399
rect 14032 1361 14111 1399
rect 14032 1327 14067 1361
rect 14101 1327 14111 1361
rect 14032 1315 14111 1327
rect 14141 1380 14193 1445
rect 14141 1346 14151 1380
rect 14185 1346 14193 1380
rect 14141 1315 14193 1346
rect 14379 1380 14431 1445
rect 14379 1346 14387 1380
rect 14421 1346 14431 1380
rect 14379 1315 14431 1346
rect 14461 1399 14513 1445
rect 16453 1399 16505 1445
rect 14461 1361 14540 1399
rect 14461 1327 14471 1361
rect 14505 1327 14540 1361
rect 14461 1315 14540 1327
rect 14570 1315 14636 1399
rect 14666 1376 14761 1399
rect 14666 1342 14678 1376
rect 14712 1342 14761 1376
rect 14666 1315 14761 1342
rect 14791 1315 14857 1399
rect 14887 1376 15025 1399
rect 14887 1342 14913 1376
rect 14947 1342 14981 1376
rect 15015 1342 15025 1376
rect 14887 1315 15025 1342
rect 15055 1376 15107 1399
rect 15055 1342 15065 1376
rect 15099 1342 15107 1376
rect 15055 1315 15107 1342
rect 15859 1376 15911 1399
rect 15859 1342 15867 1376
rect 15901 1342 15911 1376
rect 15859 1315 15911 1342
rect 15941 1376 16079 1399
rect 15941 1342 15951 1376
rect 15985 1342 16019 1376
rect 16053 1342 16079 1376
rect 15941 1315 16079 1342
rect 16109 1315 16175 1399
rect 16205 1376 16300 1399
rect 16205 1342 16254 1376
rect 16288 1342 16300 1376
rect 16205 1315 16300 1342
rect 16330 1315 16396 1399
rect 16426 1361 16505 1399
rect 16426 1327 16461 1361
rect 16495 1327 16505 1361
rect 16426 1315 16505 1327
rect 16535 1380 16587 1445
rect 16535 1346 16545 1380
rect 16579 1346 16587 1380
rect 16535 1315 16587 1346
rect 27 699 79 711
rect 27 665 35 699
rect 69 665 79 699
rect 27 627 79 665
rect 109 673 163 711
rect 109 639 119 673
rect 153 639 163 673
rect 109 627 163 639
rect 193 699 245 711
rect 193 665 203 699
rect 237 665 245 699
rect 193 627 245 665
rect 299 673 351 711
rect 299 639 307 673
rect 341 639 351 673
rect 299 627 351 639
rect 381 699 431 711
rect 806 711 857 755
rect 596 699 647 711
rect 381 691 446 699
rect 381 657 391 691
rect 425 657 446 691
rect 381 627 446 657
rect 476 673 551 699
rect 476 639 496 673
rect 530 639 551 673
rect 476 627 551 639
rect 581 627 647 699
rect 677 669 761 711
rect 677 635 717 669
rect 751 635 761 669
rect 677 627 761 635
rect 791 675 857 711
rect 791 641 801 675
rect 835 641 857 675
rect 791 627 857 641
rect 887 733 941 755
rect 887 699 897 733
rect 931 699 941 733
rect 887 627 941 699
rect 971 707 1023 755
rect 971 673 981 707
rect 1015 673 1023 707
rect 971 627 1023 673
rect 1077 673 1129 755
rect 1077 639 1085 673
rect 1119 639 1129 673
rect 1077 627 1129 639
rect 1159 699 1209 755
rect 1583 711 1633 755
rect 1378 699 1428 711
rect 1159 627 1249 699
rect 1279 673 1333 699
rect 1279 639 1289 673
rect 1323 639 1333 673
rect 1279 627 1333 639
rect 1363 627 1428 699
rect 1458 669 1525 711
rect 1458 635 1481 669
rect 1515 635 1525 669
rect 1458 627 1525 635
rect 1555 689 1633 711
rect 1555 655 1565 689
rect 1599 655 1633 689
rect 1555 627 1633 655
rect 1663 747 1717 755
rect 1663 713 1673 747
rect 1707 713 1717 747
rect 1663 627 1717 713
rect 1747 681 1799 755
rect 1950 711 2000 757
rect 1747 647 1757 681
rect 1791 647 1799 681
rect 1747 627 1799 647
rect 1853 683 1905 711
rect 1853 649 1861 683
rect 1895 649 1905 683
rect 1853 627 1905 649
rect 1935 673 2000 711
rect 1935 639 1956 673
rect 1990 639 2000 673
rect 1935 627 2000 639
rect 2030 707 2082 757
rect 2233 711 2283 757
rect 2030 673 2040 707
rect 2074 673 2082 707
rect 2030 627 2082 673
rect 2136 699 2188 711
rect 2136 665 2144 699
rect 2178 665 2188 699
rect 2136 627 2188 665
rect 2218 673 2283 711
rect 2218 639 2239 673
rect 2273 639 2283 673
rect 2218 627 2283 639
rect 2313 709 2365 757
rect 2313 675 2323 709
rect 2357 675 2365 709
rect 2313 627 2365 675
rect 2419 699 2471 711
rect 2419 665 2427 699
rect 2461 665 2471 699
rect 2419 627 2471 665
rect 2501 673 2555 711
rect 2501 639 2511 673
rect 2545 639 2555 673
rect 2501 627 2555 639
rect 2585 699 2637 711
rect 2585 665 2595 699
rect 2629 665 2637 699
rect 2585 627 2637 665
rect 2691 673 2743 711
rect 2691 639 2699 673
rect 2733 639 2743 673
rect 2691 627 2743 639
rect 2773 699 2823 711
rect 3198 711 3249 755
rect 2988 699 3039 711
rect 2773 691 2838 699
rect 2773 657 2783 691
rect 2817 657 2838 691
rect 2773 627 2838 657
rect 2868 673 2943 699
rect 2868 639 2888 673
rect 2922 639 2943 673
rect 2868 627 2943 639
rect 2973 627 3039 699
rect 3069 669 3153 711
rect 3069 635 3109 669
rect 3143 635 3153 669
rect 3069 627 3153 635
rect 3183 675 3249 711
rect 3183 641 3193 675
rect 3227 641 3249 675
rect 3183 627 3249 641
rect 3279 733 3333 755
rect 3279 699 3289 733
rect 3323 699 3333 733
rect 3279 627 3333 699
rect 3363 707 3415 755
rect 3363 673 3373 707
rect 3407 673 3415 707
rect 3363 627 3415 673
rect 3469 673 3521 755
rect 3469 639 3477 673
rect 3511 639 3521 673
rect 3469 627 3521 639
rect 3551 699 3601 755
rect 3975 711 4025 755
rect 3770 699 3820 711
rect 3551 627 3641 699
rect 3671 673 3725 699
rect 3671 639 3681 673
rect 3715 639 3725 673
rect 3671 627 3725 639
rect 3755 627 3820 699
rect 3850 669 3917 711
rect 3850 635 3873 669
rect 3907 635 3917 669
rect 3850 627 3917 635
rect 3947 689 4025 711
rect 3947 655 3957 689
rect 3991 655 4025 689
rect 3947 627 4025 655
rect 4055 747 4109 755
rect 4055 713 4065 747
rect 4099 713 4109 747
rect 4055 627 4109 713
rect 4139 681 4191 755
rect 4342 711 4392 757
rect 4139 647 4149 681
rect 4183 647 4191 681
rect 4139 627 4191 647
rect 4245 683 4297 711
rect 4245 649 4253 683
rect 4287 649 4297 683
rect 4245 627 4297 649
rect 4327 673 4392 711
rect 4327 639 4348 673
rect 4382 639 4392 673
rect 4327 627 4392 639
rect 4422 707 4474 757
rect 4625 711 4675 757
rect 4422 673 4432 707
rect 4466 673 4474 707
rect 4422 627 4474 673
rect 4528 699 4580 711
rect 4528 665 4536 699
rect 4570 665 4580 699
rect 4528 627 4580 665
rect 4610 673 4675 711
rect 4610 639 4631 673
rect 4665 639 4675 673
rect 4610 627 4675 639
rect 4705 709 4757 757
rect 4705 675 4715 709
rect 4749 675 4757 709
rect 4705 627 4757 675
rect 4811 699 4863 711
rect 4811 665 4819 699
rect 4853 665 4863 699
rect 4811 627 4863 665
rect 4893 673 4947 711
rect 4893 639 4903 673
rect 4937 639 4947 673
rect 4893 627 4947 639
rect 4977 699 5029 711
rect 4977 665 4987 699
rect 5021 665 5029 699
rect 4977 627 5029 665
rect 5083 673 5135 711
rect 5083 639 5091 673
rect 5125 639 5135 673
rect 5083 627 5135 639
rect 5165 699 5215 711
rect 5590 711 5641 755
rect 5380 699 5431 711
rect 5165 691 5230 699
rect 5165 657 5175 691
rect 5209 657 5230 691
rect 5165 627 5230 657
rect 5260 673 5335 699
rect 5260 639 5280 673
rect 5314 639 5335 673
rect 5260 627 5335 639
rect 5365 627 5431 699
rect 5461 669 5545 711
rect 5461 635 5501 669
rect 5535 635 5545 669
rect 5461 627 5545 635
rect 5575 675 5641 711
rect 5575 641 5585 675
rect 5619 641 5641 675
rect 5575 627 5641 641
rect 5671 733 5725 755
rect 5671 699 5681 733
rect 5715 699 5725 733
rect 5671 627 5725 699
rect 5755 707 5807 755
rect 5755 673 5765 707
rect 5799 673 5807 707
rect 5755 627 5807 673
rect 5861 673 5913 755
rect 5861 639 5869 673
rect 5903 639 5913 673
rect 5861 627 5913 639
rect 5943 699 5993 755
rect 6367 711 6417 755
rect 6162 699 6212 711
rect 5943 627 6033 699
rect 6063 673 6117 699
rect 6063 639 6073 673
rect 6107 639 6117 673
rect 6063 627 6117 639
rect 6147 627 6212 699
rect 6242 669 6309 711
rect 6242 635 6265 669
rect 6299 635 6309 669
rect 6242 627 6309 635
rect 6339 689 6417 711
rect 6339 655 6349 689
rect 6383 655 6417 689
rect 6339 627 6417 655
rect 6447 747 6501 755
rect 6447 713 6457 747
rect 6491 713 6501 747
rect 6447 627 6501 713
rect 6531 681 6583 755
rect 6734 711 6784 757
rect 6531 647 6541 681
rect 6575 647 6583 681
rect 6531 627 6583 647
rect 6637 683 6689 711
rect 6637 649 6645 683
rect 6679 649 6689 683
rect 6637 627 6689 649
rect 6719 673 6784 711
rect 6719 639 6740 673
rect 6774 639 6784 673
rect 6719 627 6784 639
rect 6814 707 6866 757
rect 7017 711 7067 757
rect 6814 673 6824 707
rect 6858 673 6866 707
rect 6814 627 6866 673
rect 6920 699 6972 711
rect 6920 665 6928 699
rect 6962 665 6972 699
rect 6920 627 6972 665
rect 7002 673 7067 711
rect 7002 639 7023 673
rect 7057 639 7067 673
rect 7002 627 7067 639
rect 7097 709 7149 757
rect 7097 675 7107 709
rect 7141 675 7149 709
rect 7097 627 7149 675
rect 7203 699 7255 711
rect 7203 665 7211 699
rect 7245 665 7255 699
rect 7203 627 7255 665
rect 7285 673 7339 711
rect 7285 639 7295 673
rect 7329 639 7339 673
rect 7285 627 7339 639
rect 7369 699 7421 711
rect 7369 665 7379 699
rect 7413 665 7421 699
rect 7369 627 7421 665
rect 7475 673 7527 711
rect 7475 639 7483 673
rect 7517 639 7527 673
rect 7475 627 7527 639
rect 7557 699 7607 711
rect 7982 711 8033 755
rect 7772 699 7823 711
rect 7557 691 7622 699
rect 7557 657 7567 691
rect 7601 657 7622 691
rect 7557 627 7622 657
rect 7652 673 7727 699
rect 7652 639 7672 673
rect 7706 639 7727 673
rect 7652 627 7727 639
rect 7757 627 7823 699
rect 7853 669 7937 711
rect 7853 635 7893 669
rect 7927 635 7937 669
rect 7853 627 7937 635
rect 7967 675 8033 711
rect 7967 641 7977 675
rect 8011 641 8033 675
rect 7967 627 8033 641
rect 8063 733 8117 755
rect 8063 699 8073 733
rect 8107 699 8117 733
rect 8063 627 8117 699
rect 8147 707 8199 755
rect 8147 673 8157 707
rect 8191 673 8199 707
rect 8147 627 8199 673
rect 8253 673 8305 755
rect 8253 639 8261 673
rect 8295 639 8305 673
rect 8253 627 8305 639
rect 8335 699 8385 755
rect 8759 711 8809 755
rect 8554 699 8604 711
rect 8335 627 8425 699
rect 8455 673 8509 699
rect 8455 639 8465 673
rect 8499 639 8509 673
rect 8455 627 8509 639
rect 8539 627 8604 699
rect 8634 669 8701 711
rect 8634 635 8657 669
rect 8691 635 8701 669
rect 8634 627 8701 635
rect 8731 689 8809 711
rect 8731 655 8741 689
rect 8775 655 8809 689
rect 8731 627 8809 655
rect 8839 747 8893 755
rect 8839 713 8849 747
rect 8883 713 8893 747
rect 8839 627 8893 713
rect 8923 681 8975 755
rect 9126 711 9176 757
rect 8923 647 8933 681
rect 8967 647 8975 681
rect 8923 627 8975 647
rect 9029 683 9081 711
rect 9029 649 9037 683
rect 9071 649 9081 683
rect 9029 627 9081 649
rect 9111 673 9176 711
rect 9111 639 9132 673
rect 9166 639 9176 673
rect 9111 627 9176 639
rect 9206 707 9258 757
rect 9409 711 9459 757
rect 9206 673 9216 707
rect 9250 673 9258 707
rect 9206 627 9258 673
rect 9312 699 9364 711
rect 9312 665 9320 699
rect 9354 665 9364 699
rect 9312 627 9364 665
rect 9394 673 9459 711
rect 9394 639 9415 673
rect 9449 639 9459 673
rect 9394 627 9459 639
rect 9489 709 9541 757
rect 9489 675 9499 709
rect 9533 675 9541 709
rect 9489 627 9541 675
rect 9595 699 9647 711
rect 9595 665 9603 699
rect 9637 665 9647 699
rect 9595 627 9647 665
rect 9677 673 9731 711
rect 9677 639 9687 673
rect 9721 639 9731 673
rect 9677 627 9731 639
rect 9761 699 9813 711
rect 9761 665 9771 699
rect 9805 665 9813 699
rect 9761 627 9813 665
rect 9867 673 9919 711
rect 9867 639 9875 673
rect 9909 639 9919 673
rect 9867 627 9919 639
rect 9949 699 9999 711
rect 10374 711 10425 755
rect 10164 699 10215 711
rect 9949 691 10014 699
rect 9949 657 9959 691
rect 9993 657 10014 691
rect 9949 627 10014 657
rect 10044 673 10119 699
rect 10044 639 10064 673
rect 10098 639 10119 673
rect 10044 627 10119 639
rect 10149 627 10215 699
rect 10245 669 10329 711
rect 10245 635 10285 669
rect 10319 635 10329 669
rect 10245 627 10329 635
rect 10359 675 10425 711
rect 10359 641 10369 675
rect 10403 641 10425 675
rect 10359 627 10425 641
rect 10455 733 10509 755
rect 10455 699 10465 733
rect 10499 699 10509 733
rect 10455 627 10509 699
rect 10539 707 10591 755
rect 10539 673 10549 707
rect 10583 673 10591 707
rect 10539 627 10591 673
rect 10645 673 10697 755
rect 10645 639 10653 673
rect 10687 639 10697 673
rect 10645 627 10697 639
rect 10727 699 10777 755
rect 11151 711 11201 755
rect 10946 699 10996 711
rect 10727 627 10817 699
rect 10847 673 10901 699
rect 10847 639 10857 673
rect 10891 639 10901 673
rect 10847 627 10901 639
rect 10931 627 10996 699
rect 11026 669 11093 711
rect 11026 635 11049 669
rect 11083 635 11093 669
rect 11026 627 11093 635
rect 11123 689 11201 711
rect 11123 655 11133 689
rect 11167 655 11201 689
rect 11123 627 11201 655
rect 11231 747 11285 755
rect 11231 713 11241 747
rect 11275 713 11285 747
rect 11231 627 11285 713
rect 11315 681 11367 755
rect 11518 711 11568 757
rect 11315 647 11325 681
rect 11359 647 11367 681
rect 11315 627 11367 647
rect 11421 683 11473 711
rect 11421 649 11429 683
rect 11463 649 11473 683
rect 11421 627 11473 649
rect 11503 673 11568 711
rect 11503 639 11524 673
rect 11558 639 11568 673
rect 11503 627 11568 639
rect 11598 707 11650 757
rect 11801 711 11851 757
rect 11598 673 11608 707
rect 11642 673 11650 707
rect 11598 627 11650 673
rect 11704 699 11756 711
rect 11704 665 11712 699
rect 11746 665 11756 699
rect 11704 627 11756 665
rect 11786 673 11851 711
rect 11786 639 11807 673
rect 11841 639 11851 673
rect 11786 627 11851 639
rect 11881 709 11933 757
rect 11881 675 11891 709
rect 11925 675 11933 709
rect 11881 627 11933 675
rect 11987 699 12039 711
rect 11987 665 11995 699
rect 12029 665 12039 699
rect 11987 627 12039 665
rect 12069 673 12123 711
rect 12069 639 12079 673
rect 12113 639 12123 673
rect 12069 627 12123 639
rect 12153 699 12205 711
rect 12153 665 12163 699
rect 12197 665 12205 699
rect 12153 627 12205 665
rect 12259 673 12311 711
rect 12259 639 12267 673
rect 12301 639 12311 673
rect 12259 627 12311 639
rect 12341 699 12391 711
rect 12766 711 12817 755
rect 12556 699 12607 711
rect 12341 691 12406 699
rect 12341 657 12351 691
rect 12385 657 12406 691
rect 12341 627 12406 657
rect 12436 673 12511 699
rect 12436 639 12456 673
rect 12490 639 12511 673
rect 12436 627 12511 639
rect 12541 627 12607 699
rect 12637 669 12721 711
rect 12637 635 12677 669
rect 12711 635 12721 669
rect 12637 627 12721 635
rect 12751 675 12817 711
rect 12751 641 12761 675
rect 12795 641 12817 675
rect 12751 627 12817 641
rect 12847 733 12901 755
rect 12847 699 12857 733
rect 12891 699 12901 733
rect 12847 627 12901 699
rect 12931 707 12983 755
rect 12931 673 12941 707
rect 12975 673 12983 707
rect 12931 627 12983 673
rect 13037 673 13089 755
rect 13037 639 13045 673
rect 13079 639 13089 673
rect 13037 627 13089 639
rect 13119 699 13169 755
rect 13543 711 13593 755
rect 13338 699 13388 711
rect 13119 627 13209 699
rect 13239 673 13293 699
rect 13239 639 13249 673
rect 13283 639 13293 673
rect 13239 627 13293 639
rect 13323 627 13388 699
rect 13418 669 13485 711
rect 13418 635 13441 669
rect 13475 635 13485 669
rect 13418 627 13485 635
rect 13515 689 13593 711
rect 13515 655 13525 689
rect 13559 655 13593 689
rect 13515 627 13593 655
rect 13623 747 13677 755
rect 13623 713 13633 747
rect 13667 713 13677 747
rect 13623 627 13677 713
rect 13707 681 13759 755
rect 13910 711 13960 757
rect 13707 647 13717 681
rect 13751 647 13759 681
rect 13707 627 13759 647
rect 13813 683 13865 711
rect 13813 649 13821 683
rect 13855 649 13865 683
rect 13813 627 13865 649
rect 13895 673 13960 711
rect 13895 639 13916 673
rect 13950 639 13960 673
rect 13895 627 13960 639
rect 13990 707 14042 757
rect 14193 711 14243 757
rect 13990 673 14000 707
rect 14034 673 14042 707
rect 13990 627 14042 673
rect 14096 699 14148 711
rect 14096 665 14104 699
rect 14138 665 14148 699
rect 14096 627 14148 665
rect 14178 673 14243 711
rect 14178 639 14199 673
rect 14233 639 14243 673
rect 14178 627 14243 639
rect 14273 709 14325 757
rect 14273 675 14283 709
rect 14317 675 14325 709
rect 14273 627 14325 675
rect 14379 699 14431 711
rect 14379 665 14387 699
rect 14421 665 14431 699
rect 14379 627 14431 665
rect 14461 673 14515 711
rect 14461 639 14471 673
rect 14505 639 14515 673
rect 14461 627 14515 639
rect 14545 699 14597 711
rect 14545 665 14555 699
rect 14589 665 14597 699
rect 14545 627 14597 665
rect 14651 673 14703 711
rect 14651 639 14659 673
rect 14693 639 14703 673
rect 14651 627 14703 639
rect 14733 699 14783 711
rect 15158 711 15209 755
rect 14948 699 14999 711
rect 14733 691 14798 699
rect 14733 657 14743 691
rect 14777 657 14798 691
rect 14733 627 14798 657
rect 14828 673 14903 699
rect 14828 639 14848 673
rect 14882 639 14903 673
rect 14828 627 14903 639
rect 14933 627 14999 699
rect 15029 669 15113 711
rect 15029 635 15069 669
rect 15103 635 15113 669
rect 15029 627 15113 635
rect 15143 675 15209 711
rect 15143 641 15153 675
rect 15187 641 15209 675
rect 15143 627 15209 641
rect 15239 733 15293 755
rect 15239 699 15249 733
rect 15283 699 15293 733
rect 15239 627 15293 699
rect 15323 707 15375 755
rect 15323 673 15333 707
rect 15367 673 15375 707
rect 15323 627 15375 673
rect 15429 673 15481 755
rect 15429 639 15437 673
rect 15471 639 15481 673
rect 15429 627 15481 639
rect 15511 699 15561 755
rect 15935 711 15985 755
rect 15730 699 15780 711
rect 15511 627 15601 699
rect 15631 673 15685 699
rect 15631 639 15641 673
rect 15675 639 15685 673
rect 15631 627 15685 639
rect 15715 627 15780 699
rect 15810 669 15877 711
rect 15810 635 15833 669
rect 15867 635 15877 669
rect 15810 627 15877 635
rect 15907 689 15985 711
rect 15907 655 15917 689
rect 15951 655 15985 689
rect 15907 627 15985 655
rect 16015 747 16069 755
rect 16015 713 16025 747
rect 16059 713 16069 747
rect 16015 627 16069 713
rect 16099 681 16151 755
rect 16302 711 16352 757
rect 16099 647 16109 681
rect 16143 647 16151 681
rect 16099 627 16151 647
rect 16205 683 16257 711
rect 16205 649 16213 683
rect 16247 649 16257 683
rect 16205 627 16257 649
rect 16287 673 16352 711
rect 16287 639 16308 673
rect 16342 639 16352 673
rect 16287 627 16352 639
rect 16382 707 16434 757
rect 16585 711 16635 757
rect 16382 673 16392 707
rect 16426 673 16434 707
rect 16382 627 16434 673
rect 16488 699 16540 711
rect 16488 665 16496 699
rect 16530 665 16540 699
rect 16488 627 16540 665
rect 16570 673 16635 711
rect 16570 639 16591 673
rect 16625 639 16635 673
rect 16570 627 16635 639
rect 16665 709 16717 757
rect 16665 675 16675 709
rect 16709 675 16717 709
rect 16665 627 16717 675
rect 27 20 79 68
rect 27 -14 35 20
rect 69 -14 79 20
rect 27 -62 79 -14
rect 109 22 159 68
rect 109 -16 174 22
rect 109 -50 119 -16
rect 153 -50 174 -16
rect 109 -62 174 -50
rect 204 10 256 22
rect 204 -24 214 10
rect 248 -24 256 10
rect 204 -62 256 -24
rect 310 18 362 68
rect 310 -16 318 18
rect 352 -16 362 18
rect 310 -62 362 -16
rect 392 22 442 68
rect 392 -16 457 22
rect 392 -50 402 -16
rect 436 -50 457 -16
rect 392 -62 457 -50
rect 487 -6 539 22
rect 487 -40 497 -6
rect 531 -40 539 -6
rect 487 -62 539 -40
rect 593 -8 645 66
rect 593 -42 601 -8
rect 635 -42 645 -8
rect 593 -62 645 -42
rect 675 58 729 66
rect 675 24 685 58
rect 719 24 729 58
rect 675 -62 729 24
rect 759 22 809 66
rect 759 0 837 22
rect 759 -34 793 0
rect 827 -34 837 0
rect 759 -62 837 -34
rect 867 -20 934 22
rect 867 -54 877 -20
rect 911 -54 934 -20
rect 867 -62 934 -54
rect 964 10 1014 22
rect 1183 10 1233 66
rect 964 -62 1029 10
rect 1059 -16 1113 10
rect 1059 -50 1069 -16
rect 1103 -50 1113 -16
rect 1059 -62 1113 -50
rect 1143 -62 1233 10
rect 1263 -16 1315 66
rect 1263 -50 1273 -16
rect 1307 -50 1315 -16
rect 1263 -62 1315 -50
rect 1369 18 1421 66
rect 1369 -16 1377 18
rect 1411 -16 1421 18
rect 1369 -62 1421 -16
rect 1451 44 1505 66
rect 1451 10 1461 44
rect 1495 10 1505 44
rect 1451 -62 1505 10
rect 1535 22 1586 66
rect 1535 -14 1601 22
rect 1535 -48 1557 -14
rect 1591 -48 1601 -14
rect 1535 -62 1601 -48
rect 1631 -20 1715 22
rect 1631 -54 1641 -20
rect 1675 -54 1715 -20
rect 1631 -62 1715 -54
rect 1745 10 1796 22
rect 1961 10 2011 22
rect 1745 -62 1811 10
rect 1841 -16 1916 10
rect 1841 -50 1862 -16
rect 1896 -50 1916 -16
rect 1841 -62 1916 -50
rect 1946 2 2011 10
rect 1946 -32 1967 2
rect 2001 -32 2011 2
rect 1946 -62 2011 -32
rect 2041 -16 2093 22
rect 2041 -50 2051 -16
rect 2085 -50 2093 -16
rect 2041 -62 2093 -50
rect 2147 10 2199 22
rect 2147 -24 2155 10
rect 2189 -24 2199 10
rect 2147 -62 2199 -24
rect 2229 -16 2283 22
rect 2229 -50 2239 -16
rect 2273 -50 2283 -16
rect 2229 -62 2283 -50
rect 2313 10 2365 22
rect 2313 -24 2323 10
rect 2357 -24 2365 10
rect 2313 -62 2365 -24
rect 2419 20 2471 68
rect 2419 -14 2427 20
rect 2461 -14 2471 20
rect 2419 -62 2471 -14
rect 2501 22 2551 68
rect 2501 -16 2566 22
rect 2501 -50 2511 -16
rect 2545 -50 2566 -16
rect 2501 -62 2566 -50
rect 2596 10 2648 22
rect 2596 -24 2606 10
rect 2640 -24 2648 10
rect 2596 -62 2648 -24
rect 2702 18 2754 68
rect 2702 -16 2710 18
rect 2744 -16 2754 18
rect 2702 -62 2754 -16
rect 2784 22 2834 68
rect 2784 -16 2849 22
rect 2784 -50 2794 -16
rect 2828 -50 2849 -16
rect 2784 -62 2849 -50
rect 2879 -6 2931 22
rect 2879 -40 2889 -6
rect 2923 -40 2931 -6
rect 2879 -62 2931 -40
rect 2985 -8 3037 66
rect 2985 -42 2993 -8
rect 3027 -42 3037 -8
rect 2985 -62 3037 -42
rect 3067 58 3121 66
rect 3067 24 3077 58
rect 3111 24 3121 58
rect 3067 -62 3121 24
rect 3151 22 3201 66
rect 3151 0 3229 22
rect 3151 -34 3185 0
rect 3219 -34 3229 0
rect 3151 -62 3229 -34
rect 3259 -20 3326 22
rect 3259 -54 3269 -20
rect 3303 -54 3326 -20
rect 3259 -62 3326 -54
rect 3356 10 3406 22
rect 3575 10 3625 66
rect 3356 -62 3421 10
rect 3451 -16 3505 10
rect 3451 -50 3461 -16
rect 3495 -50 3505 -16
rect 3451 -62 3505 -50
rect 3535 -62 3625 10
rect 3655 -16 3707 66
rect 3655 -50 3665 -16
rect 3699 -50 3707 -16
rect 3655 -62 3707 -50
rect 3761 18 3813 66
rect 3761 -16 3769 18
rect 3803 -16 3813 18
rect 3761 -62 3813 -16
rect 3843 44 3897 66
rect 3843 10 3853 44
rect 3887 10 3897 44
rect 3843 -62 3897 10
rect 3927 22 3978 66
rect 3927 -14 3993 22
rect 3927 -48 3949 -14
rect 3983 -48 3993 -14
rect 3927 -62 3993 -48
rect 4023 -20 4107 22
rect 4023 -54 4033 -20
rect 4067 -54 4107 -20
rect 4023 -62 4107 -54
rect 4137 10 4188 22
rect 4353 10 4403 22
rect 4137 -62 4203 10
rect 4233 -16 4308 10
rect 4233 -50 4254 -16
rect 4288 -50 4308 -16
rect 4233 -62 4308 -50
rect 4338 2 4403 10
rect 4338 -32 4359 2
rect 4393 -32 4403 2
rect 4338 -62 4403 -32
rect 4433 -16 4485 22
rect 4433 -50 4443 -16
rect 4477 -50 4485 -16
rect 4433 -62 4485 -50
rect 4539 10 4591 22
rect 4539 -24 4547 10
rect 4581 -24 4591 10
rect 4539 -62 4591 -24
rect 4621 -16 4675 22
rect 4621 -50 4631 -16
rect 4665 -50 4675 -16
rect 4621 -62 4675 -50
rect 4705 10 4757 22
rect 4705 -24 4715 10
rect 4749 -24 4757 10
rect 4705 -62 4757 -24
rect 4811 20 4863 68
rect 4811 -14 4819 20
rect 4853 -14 4863 20
rect 4811 -62 4863 -14
rect 4893 22 4943 68
rect 4893 -16 4958 22
rect 4893 -50 4903 -16
rect 4937 -50 4958 -16
rect 4893 -62 4958 -50
rect 4988 10 5040 22
rect 4988 -24 4998 10
rect 5032 -24 5040 10
rect 4988 -62 5040 -24
rect 5094 18 5146 68
rect 5094 -16 5102 18
rect 5136 -16 5146 18
rect 5094 -62 5146 -16
rect 5176 22 5226 68
rect 5176 -16 5241 22
rect 5176 -50 5186 -16
rect 5220 -50 5241 -16
rect 5176 -62 5241 -50
rect 5271 -6 5323 22
rect 5271 -40 5281 -6
rect 5315 -40 5323 -6
rect 5271 -62 5323 -40
rect 5377 -8 5429 66
rect 5377 -42 5385 -8
rect 5419 -42 5429 -8
rect 5377 -62 5429 -42
rect 5459 58 5513 66
rect 5459 24 5469 58
rect 5503 24 5513 58
rect 5459 -62 5513 24
rect 5543 22 5593 66
rect 5543 0 5621 22
rect 5543 -34 5577 0
rect 5611 -34 5621 0
rect 5543 -62 5621 -34
rect 5651 -20 5718 22
rect 5651 -54 5661 -20
rect 5695 -54 5718 -20
rect 5651 -62 5718 -54
rect 5748 10 5798 22
rect 5967 10 6017 66
rect 5748 -62 5813 10
rect 5843 -16 5897 10
rect 5843 -50 5853 -16
rect 5887 -50 5897 -16
rect 5843 -62 5897 -50
rect 5927 -62 6017 10
rect 6047 -16 6099 66
rect 6047 -50 6057 -16
rect 6091 -50 6099 -16
rect 6047 -62 6099 -50
rect 6153 18 6205 66
rect 6153 -16 6161 18
rect 6195 -16 6205 18
rect 6153 -62 6205 -16
rect 6235 44 6289 66
rect 6235 10 6245 44
rect 6279 10 6289 44
rect 6235 -62 6289 10
rect 6319 22 6370 66
rect 6319 -14 6385 22
rect 6319 -48 6341 -14
rect 6375 -48 6385 -14
rect 6319 -62 6385 -48
rect 6415 -20 6499 22
rect 6415 -54 6425 -20
rect 6459 -54 6499 -20
rect 6415 -62 6499 -54
rect 6529 10 6580 22
rect 6745 10 6795 22
rect 6529 -62 6595 10
rect 6625 -16 6700 10
rect 6625 -50 6646 -16
rect 6680 -50 6700 -16
rect 6625 -62 6700 -50
rect 6730 2 6795 10
rect 6730 -32 6751 2
rect 6785 -32 6795 2
rect 6730 -62 6795 -32
rect 6825 -16 6877 22
rect 6825 -50 6835 -16
rect 6869 -50 6877 -16
rect 6825 -62 6877 -50
rect 6931 10 6983 22
rect 6931 -24 6939 10
rect 6973 -24 6983 10
rect 6931 -62 6983 -24
rect 7013 -16 7067 22
rect 7013 -50 7023 -16
rect 7057 -50 7067 -16
rect 7013 -62 7067 -50
rect 7097 10 7149 22
rect 7097 -24 7107 10
rect 7141 -24 7149 10
rect 7097 -62 7149 -24
rect 7203 20 7255 68
rect 7203 -14 7211 20
rect 7245 -14 7255 20
rect 7203 -62 7255 -14
rect 7285 22 7335 68
rect 7285 -16 7350 22
rect 7285 -50 7295 -16
rect 7329 -50 7350 -16
rect 7285 -62 7350 -50
rect 7380 10 7432 22
rect 7380 -24 7390 10
rect 7424 -24 7432 10
rect 7380 -62 7432 -24
rect 7486 18 7538 68
rect 7486 -16 7494 18
rect 7528 -16 7538 18
rect 7486 -62 7538 -16
rect 7568 22 7618 68
rect 7568 -16 7633 22
rect 7568 -50 7578 -16
rect 7612 -50 7633 -16
rect 7568 -62 7633 -50
rect 7663 -6 7715 22
rect 7663 -40 7673 -6
rect 7707 -40 7715 -6
rect 7663 -62 7715 -40
rect 7769 -8 7821 66
rect 7769 -42 7777 -8
rect 7811 -42 7821 -8
rect 7769 -62 7821 -42
rect 7851 58 7905 66
rect 7851 24 7861 58
rect 7895 24 7905 58
rect 7851 -62 7905 24
rect 7935 22 7985 66
rect 7935 0 8013 22
rect 7935 -34 7969 0
rect 8003 -34 8013 0
rect 7935 -62 8013 -34
rect 8043 -20 8110 22
rect 8043 -54 8053 -20
rect 8087 -54 8110 -20
rect 8043 -62 8110 -54
rect 8140 10 8190 22
rect 8359 10 8409 66
rect 8140 -62 8205 10
rect 8235 -16 8289 10
rect 8235 -50 8245 -16
rect 8279 -50 8289 -16
rect 8235 -62 8289 -50
rect 8319 -62 8409 10
rect 8439 -16 8491 66
rect 8439 -50 8449 -16
rect 8483 -50 8491 -16
rect 8439 -62 8491 -50
rect 8545 18 8597 66
rect 8545 -16 8553 18
rect 8587 -16 8597 18
rect 8545 -62 8597 -16
rect 8627 44 8681 66
rect 8627 10 8637 44
rect 8671 10 8681 44
rect 8627 -62 8681 10
rect 8711 22 8762 66
rect 8711 -14 8777 22
rect 8711 -48 8733 -14
rect 8767 -48 8777 -14
rect 8711 -62 8777 -48
rect 8807 -20 8891 22
rect 8807 -54 8817 -20
rect 8851 -54 8891 -20
rect 8807 -62 8891 -54
rect 8921 10 8972 22
rect 9137 10 9187 22
rect 8921 -62 8987 10
rect 9017 -16 9092 10
rect 9017 -50 9038 -16
rect 9072 -50 9092 -16
rect 9017 -62 9092 -50
rect 9122 2 9187 10
rect 9122 -32 9143 2
rect 9177 -32 9187 2
rect 9122 -62 9187 -32
rect 9217 -16 9269 22
rect 9217 -50 9227 -16
rect 9261 -50 9269 -16
rect 9217 -62 9269 -50
rect 9323 10 9375 22
rect 9323 -24 9331 10
rect 9365 -24 9375 10
rect 9323 -62 9375 -24
rect 9405 -16 9459 22
rect 9405 -50 9415 -16
rect 9449 -50 9459 -16
rect 9405 -62 9459 -50
rect 9489 10 9541 22
rect 9489 -24 9499 10
rect 9533 -24 9541 10
rect 9489 -62 9541 -24
rect 9595 20 9647 68
rect 9595 -14 9603 20
rect 9637 -14 9647 20
rect 9595 -62 9647 -14
rect 9677 22 9727 68
rect 9677 -16 9742 22
rect 9677 -50 9687 -16
rect 9721 -50 9742 -16
rect 9677 -62 9742 -50
rect 9772 10 9824 22
rect 9772 -24 9782 10
rect 9816 -24 9824 10
rect 9772 -62 9824 -24
rect 9878 18 9930 68
rect 9878 -16 9886 18
rect 9920 -16 9930 18
rect 9878 -62 9930 -16
rect 9960 22 10010 68
rect 9960 -16 10025 22
rect 9960 -50 9970 -16
rect 10004 -50 10025 -16
rect 9960 -62 10025 -50
rect 10055 -6 10107 22
rect 10055 -40 10065 -6
rect 10099 -40 10107 -6
rect 10055 -62 10107 -40
rect 10161 -8 10213 66
rect 10161 -42 10169 -8
rect 10203 -42 10213 -8
rect 10161 -62 10213 -42
rect 10243 58 10297 66
rect 10243 24 10253 58
rect 10287 24 10297 58
rect 10243 -62 10297 24
rect 10327 22 10377 66
rect 10327 0 10405 22
rect 10327 -34 10361 0
rect 10395 -34 10405 0
rect 10327 -62 10405 -34
rect 10435 -20 10502 22
rect 10435 -54 10445 -20
rect 10479 -54 10502 -20
rect 10435 -62 10502 -54
rect 10532 10 10582 22
rect 10751 10 10801 66
rect 10532 -62 10597 10
rect 10627 -16 10681 10
rect 10627 -50 10637 -16
rect 10671 -50 10681 -16
rect 10627 -62 10681 -50
rect 10711 -62 10801 10
rect 10831 -16 10883 66
rect 10831 -50 10841 -16
rect 10875 -50 10883 -16
rect 10831 -62 10883 -50
rect 10937 18 10989 66
rect 10937 -16 10945 18
rect 10979 -16 10989 18
rect 10937 -62 10989 -16
rect 11019 44 11073 66
rect 11019 10 11029 44
rect 11063 10 11073 44
rect 11019 -62 11073 10
rect 11103 22 11154 66
rect 11103 -14 11169 22
rect 11103 -48 11125 -14
rect 11159 -48 11169 -14
rect 11103 -62 11169 -48
rect 11199 -20 11283 22
rect 11199 -54 11209 -20
rect 11243 -54 11283 -20
rect 11199 -62 11283 -54
rect 11313 10 11364 22
rect 11529 10 11579 22
rect 11313 -62 11379 10
rect 11409 -16 11484 10
rect 11409 -50 11430 -16
rect 11464 -50 11484 -16
rect 11409 -62 11484 -50
rect 11514 2 11579 10
rect 11514 -32 11535 2
rect 11569 -32 11579 2
rect 11514 -62 11579 -32
rect 11609 -16 11661 22
rect 11609 -50 11619 -16
rect 11653 -50 11661 -16
rect 11609 -62 11661 -50
rect 11715 10 11767 22
rect 11715 -24 11723 10
rect 11757 -24 11767 10
rect 11715 -62 11767 -24
rect 11797 -16 11851 22
rect 11797 -50 11807 -16
rect 11841 -50 11851 -16
rect 11797 -62 11851 -50
rect 11881 10 11933 22
rect 11881 -24 11891 10
rect 11925 -24 11933 10
rect 11881 -62 11933 -24
rect 11987 20 12039 68
rect 11987 -14 11995 20
rect 12029 -14 12039 20
rect 11987 -62 12039 -14
rect 12069 22 12119 68
rect 12069 -16 12134 22
rect 12069 -50 12079 -16
rect 12113 -50 12134 -16
rect 12069 -62 12134 -50
rect 12164 10 12216 22
rect 12164 -24 12174 10
rect 12208 -24 12216 10
rect 12164 -62 12216 -24
rect 12270 18 12322 68
rect 12270 -16 12278 18
rect 12312 -16 12322 18
rect 12270 -62 12322 -16
rect 12352 22 12402 68
rect 12352 -16 12417 22
rect 12352 -50 12362 -16
rect 12396 -50 12417 -16
rect 12352 -62 12417 -50
rect 12447 -6 12499 22
rect 12447 -40 12457 -6
rect 12491 -40 12499 -6
rect 12447 -62 12499 -40
rect 12553 -8 12605 66
rect 12553 -42 12561 -8
rect 12595 -42 12605 -8
rect 12553 -62 12605 -42
rect 12635 58 12689 66
rect 12635 24 12645 58
rect 12679 24 12689 58
rect 12635 -62 12689 24
rect 12719 22 12769 66
rect 12719 0 12797 22
rect 12719 -34 12753 0
rect 12787 -34 12797 0
rect 12719 -62 12797 -34
rect 12827 -20 12894 22
rect 12827 -54 12837 -20
rect 12871 -54 12894 -20
rect 12827 -62 12894 -54
rect 12924 10 12974 22
rect 13143 10 13193 66
rect 12924 -62 12989 10
rect 13019 -16 13073 10
rect 13019 -50 13029 -16
rect 13063 -50 13073 -16
rect 13019 -62 13073 -50
rect 13103 -62 13193 10
rect 13223 -16 13275 66
rect 13223 -50 13233 -16
rect 13267 -50 13275 -16
rect 13223 -62 13275 -50
rect 13329 18 13381 66
rect 13329 -16 13337 18
rect 13371 -16 13381 18
rect 13329 -62 13381 -16
rect 13411 44 13465 66
rect 13411 10 13421 44
rect 13455 10 13465 44
rect 13411 -62 13465 10
rect 13495 22 13546 66
rect 13495 -14 13561 22
rect 13495 -48 13517 -14
rect 13551 -48 13561 -14
rect 13495 -62 13561 -48
rect 13591 -20 13675 22
rect 13591 -54 13601 -20
rect 13635 -54 13675 -20
rect 13591 -62 13675 -54
rect 13705 10 13756 22
rect 13921 10 13971 22
rect 13705 -62 13771 10
rect 13801 -16 13876 10
rect 13801 -50 13822 -16
rect 13856 -50 13876 -16
rect 13801 -62 13876 -50
rect 13906 2 13971 10
rect 13906 -32 13927 2
rect 13961 -32 13971 2
rect 13906 -62 13971 -32
rect 14001 -16 14053 22
rect 14001 -50 14011 -16
rect 14045 -50 14053 -16
rect 14001 -62 14053 -50
rect 14107 10 14159 22
rect 14107 -24 14115 10
rect 14149 -24 14159 10
rect 14107 -62 14159 -24
rect 14189 -16 14243 22
rect 14189 -50 14199 -16
rect 14233 -50 14243 -16
rect 14189 -62 14243 -50
rect 14273 10 14325 22
rect 14273 -24 14283 10
rect 14317 -24 14325 10
rect 14273 -62 14325 -24
rect 14379 20 14431 68
rect 14379 -14 14387 20
rect 14421 -14 14431 20
rect 14379 -62 14431 -14
rect 14461 22 14511 68
rect 14461 -16 14526 22
rect 14461 -50 14471 -16
rect 14505 -50 14526 -16
rect 14461 -62 14526 -50
rect 14556 10 14608 22
rect 14556 -24 14566 10
rect 14600 -24 14608 10
rect 14556 -62 14608 -24
rect 14662 18 14714 68
rect 14662 -16 14670 18
rect 14704 -16 14714 18
rect 14662 -62 14714 -16
rect 14744 22 14794 68
rect 14744 -16 14809 22
rect 14744 -50 14754 -16
rect 14788 -50 14809 -16
rect 14744 -62 14809 -50
rect 14839 -6 14891 22
rect 14839 -40 14849 -6
rect 14883 -40 14891 -6
rect 14839 -62 14891 -40
rect 14945 -8 14997 66
rect 14945 -42 14953 -8
rect 14987 -42 14997 -8
rect 14945 -62 14997 -42
rect 15027 58 15081 66
rect 15027 24 15037 58
rect 15071 24 15081 58
rect 15027 -62 15081 24
rect 15111 22 15161 66
rect 15111 0 15189 22
rect 15111 -34 15145 0
rect 15179 -34 15189 0
rect 15111 -62 15189 -34
rect 15219 -20 15286 22
rect 15219 -54 15229 -20
rect 15263 -54 15286 -20
rect 15219 -62 15286 -54
rect 15316 10 15366 22
rect 15535 10 15585 66
rect 15316 -62 15381 10
rect 15411 -16 15465 10
rect 15411 -50 15421 -16
rect 15455 -50 15465 -16
rect 15411 -62 15465 -50
rect 15495 -62 15585 10
rect 15615 -16 15667 66
rect 15615 -50 15625 -16
rect 15659 -50 15667 -16
rect 15615 -62 15667 -50
rect 15721 18 15773 66
rect 15721 -16 15729 18
rect 15763 -16 15773 18
rect 15721 -62 15773 -16
rect 15803 44 15857 66
rect 15803 10 15813 44
rect 15847 10 15857 44
rect 15803 -62 15857 10
rect 15887 22 15938 66
rect 15887 -14 15953 22
rect 15887 -48 15909 -14
rect 15943 -48 15953 -14
rect 15887 -62 15953 -48
rect 15983 -20 16067 22
rect 15983 -54 15993 -20
rect 16027 -54 16067 -20
rect 15983 -62 16067 -54
rect 16097 10 16148 22
rect 16313 10 16363 22
rect 16097 -62 16163 10
rect 16193 -16 16268 10
rect 16193 -50 16214 -16
rect 16248 -50 16268 -16
rect 16193 -62 16268 -50
rect 16298 2 16363 10
rect 16298 -32 16319 2
rect 16353 -32 16363 2
rect 16298 -62 16363 -32
rect 16393 -16 16445 22
rect 16393 -50 16403 -16
rect 16437 -50 16445 -16
rect 16393 -62 16445 -50
rect 16499 10 16551 22
rect 16499 -24 16507 10
rect 16541 -24 16551 10
rect 16499 -62 16551 -24
rect 16581 -16 16635 22
rect 16581 -50 16591 -16
rect 16625 -50 16635 -16
rect 16581 -62 16635 -50
rect 16665 10 16717 22
rect 16665 -24 16675 10
rect 16709 -24 16717 10
rect 16665 -62 16717 -24
<< pdiff >>
rect 29 2887 81 2907
rect 29 2853 37 2887
rect 71 2853 81 2887
rect 29 2819 81 2853
rect 29 2785 37 2819
rect 71 2785 81 2819
rect 29 2749 81 2785
rect 111 2887 169 2907
rect 111 2853 123 2887
rect 157 2853 169 2887
rect 111 2819 169 2853
rect 111 2785 123 2819
rect 157 2785 169 2819
rect 111 2749 169 2785
rect 199 2887 251 2907
rect 199 2853 209 2887
rect 243 2853 251 2887
rect 199 2806 251 2853
rect 199 2772 209 2806
rect 243 2772 251 2806
rect 199 2749 251 2772
rect 305 2889 357 2907
rect 305 2855 313 2889
rect 347 2855 357 2889
rect 305 2821 357 2855
rect 305 2787 313 2821
rect 347 2787 357 2821
rect 305 2753 357 2787
rect 305 2719 313 2753
rect 347 2719 357 2753
rect 305 2707 357 2719
rect 387 2895 441 2907
rect 387 2861 397 2895
rect 431 2861 441 2895
rect 387 2827 441 2861
rect 387 2793 397 2827
rect 431 2793 441 2827
rect 387 2707 441 2793
rect 471 2873 525 2907
rect 471 2839 481 2873
rect 515 2839 525 2873
rect 471 2778 525 2839
rect 471 2744 481 2778
rect 515 2744 525 2778
rect 471 2707 525 2744
rect 555 2895 609 2907
rect 555 2861 565 2895
rect 599 2861 609 2895
rect 555 2827 609 2861
rect 555 2793 565 2827
rect 599 2793 609 2827
rect 555 2707 609 2793
rect 639 2873 693 2907
rect 639 2839 649 2873
rect 683 2839 693 2873
rect 639 2778 693 2839
rect 639 2744 649 2778
rect 683 2744 693 2778
rect 639 2707 693 2744
rect 723 2895 775 2907
rect 723 2861 733 2895
rect 767 2861 775 2895
rect 723 2827 775 2861
rect 723 2793 733 2827
rect 767 2793 775 2827
rect 723 2759 775 2793
rect 723 2725 733 2759
rect 767 2725 775 2759
rect 723 2707 775 2725
rect 857 2895 909 2907
rect 857 2861 865 2895
rect 899 2861 909 2895
rect 857 2827 909 2861
rect 857 2793 865 2827
rect 899 2793 909 2827
rect 857 2759 909 2793
rect 857 2725 865 2759
rect 899 2725 909 2759
rect 857 2707 909 2725
rect 939 2889 993 2907
rect 939 2855 949 2889
rect 983 2855 993 2889
rect 939 2821 993 2855
rect 939 2787 949 2821
rect 983 2787 993 2821
rect 939 2753 993 2787
rect 939 2719 949 2753
rect 983 2719 993 2753
rect 939 2707 993 2719
rect 1023 2895 1077 2907
rect 1023 2861 1033 2895
rect 1067 2861 1077 2895
rect 1023 2827 1077 2861
rect 1023 2793 1033 2827
rect 1067 2793 1077 2827
rect 1023 2707 1077 2793
rect 1107 2889 1161 2907
rect 1107 2855 1117 2889
rect 1151 2855 1161 2889
rect 1107 2821 1161 2855
rect 1107 2787 1117 2821
rect 1151 2787 1161 2821
rect 1107 2753 1161 2787
rect 1107 2719 1117 2753
rect 1151 2719 1161 2753
rect 1107 2707 1161 2719
rect 1191 2895 1245 2907
rect 1191 2861 1201 2895
rect 1235 2861 1245 2895
rect 1191 2827 1245 2861
rect 1191 2793 1201 2827
rect 1235 2793 1245 2827
rect 1191 2707 1245 2793
rect 1275 2889 1329 2907
rect 1275 2855 1285 2889
rect 1319 2855 1329 2889
rect 1275 2821 1329 2855
rect 1275 2787 1285 2821
rect 1319 2787 1329 2821
rect 1275 2753 1329 2787
rect 1275 2719 1285 2753
rect 1319 2719 1329 2753
rect 1275 2707 1329 2719
rect 1359 2895 1413 2907
rect 1359 2861 1369 2895
rect 1403 2861 1413 2895
rect 1359 2827 1413 2861
rect 1359 2793 1369 2827
rect 1403 2793 1413 2827
rect 1359 2707 1413 2793
rect 1443 2889 1497 2907
rect 1443 2855 1453 2889
rect 1487 2855 1497 2889
rect 1443 2821 1497 2855
rect 1443 2787 1453 2821
rect 1487 2787 1497 2821
rect 1443 2753 1497 2787
rect 1443 2719 1453 2753
rect 1487 2719 1497 2753
rect 1443 2707 1497 2719
rect 1527 2895 1581 2907
rect 1527 2861 1537 2895
rect 1571 2861 1581 2895
rect 1527 2827 1581 2861
rect 1527 2793 1537 2827
rect 1571 2793 1581 2827
rect 1527 2707 1581 2793
rect 1611 2889 1665 2907
rect 1611 2855 1621 2889
rect 1655 2855 1665 2889
rect 1611 2821 1665 2855
rect 1611 2787 1621 2821
rect 1655 2787 1665 2821
rect 1611 2753 1665 2787
rect 1611 2719 1621 2753
rect 1655 2719 1665 2753
rect 1611 2707 1665 2719
rect 1695 2895 1749 2907
rect 1695 2861 1705 2895
rect 1739 2861 1749 2895
rect 1695 2827 1749 2861
rect 1695 2793 1705 2827
rect 1739 2793 1749 2827
rect 1695 2707 1749 2793
rect 1779 2889 1833 2907
rect 1779 2855 1789 2889
rect 1823 2855 1833 2889
rect 1779 2821 1833 2855
rect 1779 2787 1789 2821
rect 1823 2787 1833 2821
rect 1779 2753 1833 2787
rect 1779 2719 1789 2753
rect 1823 2719 1833 2753
rect 1779 2707 1833 2719
rect 1863 2895 1917 2907
rect 1863 2861 1873 2895
rect 1907 2861 1917 2895
rect 1863 2827 1917 2861
rect 1863 2793 1873 2827
rect 1907 2793 1917 2827
rect 1863 2707 1917 2793
rect 1947 2889 2001 2907
rect 1947 2855 1957 2889
rect 1991 2855 2001 2889
rect 1947 2821 2001 2855
rect 1947 2787 1957 2821
rect 1991 2787 2001 2821
rect 1947 2753 2001 2787
rect 1947 2719 1957 2753
rect 1991 2719 2001 2753
rect 1947 2707 2001 2719
rect 2031 2895 2085 2907
rect 2031 2861 2041 2895
rect 2075 2861 2085 2895
rect 2031 2827 2085 2861
rect 2031 2793 2041 2827
rect 2075 2793 2085 2827
rect 2031 2707 2085 2793
rect 2115 2889 2169 2907
rect 2115 2855 2125 2889
rect 2159 2855 2169 2889
rect 2115 2821 2169 2855
rect 2115 2787 2125 2821
rect 2159 2787 2169 2821
rect 2115 2753 2169 2787
rect 2115 2719 2125 2753
rect 2159 2719 2169 2753
rect 2115 2707 2169 2719
rect 2199 2895 2253 2907
rect 2199 2861 2209 2895
rect 2243 2861 2253 2895
rect 2199 2827 2253 2861
rect 2199 2793 2209 2827
rect 2243 2793 2253 2827
rect 2199 2707 2253 2793
rect 2283 2889 2337 2907
rect 2283 2855 2293 2889
rect 2327 2855 2337 2889
rect 2283 2821 2337 2855
rect 2283 2787 2293 2821
rect 2327 2787 2337 2821
rect 2283 2753 2337 2787
rect 2283 2719 2293 2753
rect 2327 2719 2337 2753
rect 2283 2707 2337 2719
rect 2367 2895 2421 2907
rect 2367 2861 2377 2895
rect 2411 2861 2421 2895
rect 2367 2827 2421 2861
rect 2367 2793 2377 2827
rect 2411 2793 2421 2827
rect 2367 2707 2421 2793
rect 2451 2889 2505 2907
rect 2451 2855 2461 2889
rect 2495 2855 2505 2889
rect 2451 2821 2505 2855
rect 2451 2787 2461 2821
rect 2495 2787 2505 2821
rect 2451 2753 2505 2787
rect 2451 2719 2461 2753
rect 2495 2719 2505 2753
rect 2451 2707 2505 2719
rect 2535 2895 2589 2907
rect 2535 2861 2545 2895
rect 2579 2861 2589 2895
rect 2535 2827 2589 2861
rect 2535 2793 2545 2827
rect 2579 2793 2589 2827
rect 2535 2707 2589 2793
rect 2619 2889 2673 2907
rect 2619 2855 2629 2889
rect 2663 2855 2673 2889
rect 2619 2821 2673 2855
rect 2619 2787 2629 2821
rect 2663 2787 2673 2821
rect 2619 2753 2673 2787
rect 2619 2719 2629 2753
rect 2663 2719 2673 2753
rect 2619 2707 2673 2719
rect 2703 2895 2755 2907
rect 2703 2861 2713 2895
rect 2747 2861 2755 2895
rect 2703 2827 2755 2861
rect 2703 2793 2713 2827
rect 2747 2793 2755 2827
rect 2703 2707 2755 2793
rect 4413 2887 4465 2907
rect 4413 2853 4421 2887
rect 4455 2853 4465 2887
rect 4413 2819 4465 2853
rect 4413 2785 4421 2819
rect 4455 2785 4465 2819
rect 4413 2749 4465 2785
rect 4495 2887 4553 2907
rect 4495 2853 4507 2887
rect 4541 2853 4553 2887
rect 4495 2819 4553 2853
rect 4495 2785 4507 2819
rect 4541 2785 4553 2819
rect 4495 2749 4553 2785
rect 4583 2887 4635 2907
rect 4583 2853 4593 2887
rect 4627 2853 4635 2887
rect 4583 2806 4635 2853
rect 4583 2772 4593 2806
rect 4627 2772 4635 2806
rect 4583 2749 4635 2772
rect 4689 2889 4741 2907
rect 4689 2855 4697 2889
rect 4731 2855 4741 2889
rect 4689 2821 4741 2855
rect 4689 2787 4697 2821
rect 4731 2787 4741 2821
rect 4689 2753 4741 2787
rect 4689 2719 4697 2753
rect 4731 2719 4741 2753
rect 4689 2707 4741 2719
rect 4771 2895 4825 2907
rect 4771 2861 4781 2895
rect 4815 2861 4825 2895
rect 4771 2827 4825 2861
rect 4771 2793 4781 2827
rect 4815 2793 4825 2827
rect 4771 2707 4825 2793
rect 4855 2873 4909 2907
rect 4855 2839 4865 2873
rect 4899 2839 4909 2873
rect 4855 2778 4909 2839
rect 4855 2744 4865 2778
rect 4899 2744 4909 2778
rect 4855 2707 4909 2744
rect 4939 2895 4993 2907
rect 4939 2861 4949 2895
rect 4983 2861 4993 2895
rect 4939 2827 4993 2861
rect 4939 2793 4949 2827
rect 4983 2793 4993 2827
rect 4939 2707 4993 2793
rect 5023 2873 5077 2907
rect 5023 2839 5033 2873
rect 5067 2839 5077 2873
rect 5023 2778 5077 2839
rect 5023 2744 5033 2778
rect 5067 2744 5077 2778
rect 5023 2707 5077 2744
rect 5107 2895 5159 2907
rect 5107 2861 5117 2895
rect 5151 2861 5159 2895
rect 5107 2827 5159 2861
rect 5107 2793 5117 2827
rect 5151 2793 5159 2827
rect 5107 2759 5159 2793
rect 5107 2725 5117 2759
rect 5151 2725 5159 2759
rect 5107 2707 5159 2725
rect 5241 2895 5293 2907
rect 5241 2861 5249 2895
rect 5283 2861 5293 2895
rect 5241 2827 5293 2861
rect 5241 2793 5249 2827
rect 5283 2793 5293 2827
rect 5241 2759 5293 2793
rect 5241 2725 5249 2759
rect 5283 2725 5293 2759
rect 5241 2707 5293 2725
rect 5323 2889 5377 2907
rect 5323 2855 5333 2889
rect 5367 2855 5377 2889
rect 5323 2821 5377 2855
rect 5323 2787 5333 2821
rect 5367 2787 5377 2821
rect 5323 2753 5377 2787
rect 5323 2719 5333 2753
rect 5367 2719 5377 2753
rect 5323 2707 5377 2719
rect 5407 2895 5461 2907
rect 5407 2861 5417 2895
rect 5451 2861 5461 2895
rect 5407 2827 5461 2861
rect 5407 2793 5417 2827
rect 5451 2793 5461 2827
rect 5407 2707 5461 2793
rect 5491 2889 5545 2907
rect 5491 2855 5501 2889
rect 5535 2855 5545 2889
rect 5491 2821 5545 2855
rect 5491 2787 5501 2821
rect 5535 2787 5545 2821
rect 5491 2753 5545 2787
rect 5491 2719 5501 2753
rect 5535 2719 5545 2753
rect 5491 2707 5545 2719
rect 5575 2895 5629 2907
rect 5575 2861 5585 2895
rect 5619 2861 5629 2895
rect 5575 2827 5629 2861
rect 5575 2793 5585 2827
rect 5619 2793 5629 2827
rect 5575 2707 5629 2793
rect 5659 2889 5713 2907
rect 5659 2855 5669 2889
rect 5703 2855 5713 2889
rect 5659 2821 5713 2855
rect 5659 2787 5669 2821
rect 5703 2787 5713 2821
rect 5659 2753 5713 2787
rect 5659 2719 5669 2753
rect 5703 2719 5713 2753
rect 5659 2707 5713 2719
rect 5743 2895 5797 2907
rect 5743 2861 5753 2895
rect 5787 2861 5797 2895
rect 5743 2827 5797 2861
rect 5743 2793 5753 2827
rect 5787 2793 5797 2827
rect 5743 2707 5797 2793
rect 5827 2889 5881 2907
rect 5827 2855 5837 2889
rect 5871 2855 5881 2889
rect 5827 2821 5881 2855
rect 5827 2787 5837 2821
rect 5871 2787 5881 2821
rect 5827 2753 5881 2787
rect 5827 2719 5837 2753
rect 5871 2719 5881 2753
rect 5827 2707 5881 2719
rect 5911 2895 5965 2907
rect 5911 2861 5921 2895
rect 5955 2861 5965 2895
rect 5911 2827 5965 2861
rect 5911 2793 5921 2827
rect 5955 2793 5965 2827
rect 5911 2707 5965 2793
rect 5995 2889 6049 2907
rect 5995 2855 6005 2889
rect 6039 2855 6049 2889
rect 5995 2821 6049 2855
rect 5995 2787 6005 2821
rect 6039 2787 6049 2821
rect 5995 2753 6049 2787
rect 5995 2719 6005 2753
rect 6039 2719 6049 2753
rect 5995 2707 6049 2719
rect 6079 2895 6133 2907
rect 6079 2861 6089 2895
rect 6123 2861 6133 2895
rect 6079 2827 6133 2861
rect 6079 2793 6089 2827
rect 6123 2793 6133 2827
rect 6079 2707 6133 2793
rect 6163 2889 6217 2907
rect 6163 2855 6173 2889
rect 6207 2855 6217 2889
rect 6163 2821 6217 2855
rect 6163 2787 6173 2821
rect 6207 2787 6217 2821
rect 6163 2753 6217 2787
rect 6163 2719 6173 2753
rect 6207 2719 6217 2753
rect 6163 2707 6217 2719
rect 6247 2895 6301 2907
rect 6247 2861 6257 2895
rect 6291 2861 6301 2895
rect 6247 2827 6301 2861
rect 6247 2793 6257 2827
rect 6291 2793 6301 2827
rect 6247 2707 6301 2793
rect 6331 2889 6385 2907
rect 6331 2855 6341 2889
rect 6375 2855 6385 2889
rect 6331 2821 6385 2855
rect 6331 2787 6341 2821
rect 6375 2787 6385 2821
rect 6331 2753 6385 2787
rect 6331 2719 6341 2753
rect 6375 2719 6385 2753
rect 6331 2707 6385 2719
rect 6415 2895 6469 2907
rect 6415 2861 6425 2895
rect 6459 2861 6469 2895
rect 6415 2827 6469 2861
rect 6415 2793 6425 2827
rect 6459 2793 6469 2827
rect 6415 2707 6469 2793
rect 6499 2889 6553 2907
rect 6499 2855 6509 2889
rect 6543 2855 6553 2889
rect 6499 2821 6553 2855
rect 6499 2787 6509 2821
rect 6543 2787 6553 2821
rect 6499 2753 6553 2787
rect 6499 2719 6509 2753
rect 6543 2719 6553 2753
rect 6499 2707 6553 2719
rect 6583 2895 6637 2907
rect 6583 2861 6593 2895
rect 6627 2861 6637 2895
rect 6583 2827 6637 2861
rect 6583 2793 6593 2827
rect 6627 2793 6637 2827
rect 6583 2707 6637 2793
rect 6667 2889 6721 2907
rect 6667 2855 6677 2889
rect 6711 2855 6721 2889
rect 6667 2821 6721 2855
rect 6667 2787 6677 2821
rect 6711 2787 6721 2821
rect 6667 2753 6721 2787
rect 6667 2719 6677 2753
rect 6711 2719 6721 2753
rect 6667 2707 6721 2719
rect 6751 2895 6805 2907
rect 6751 2861 6761 2895
rect 6795 2861 6805 2895
rect 6751 2827 6805 2861
rect 6751 2793 6761 2827
rect 6795 2793 6805 2827
rect 6751 2707 6805 2793
rect 6835 2889 6889 2907
rect 6835 2855 6845 2889
rect 6879 2855 6889 2889
rect 6835 2821 6889 2855
rect 6835 2787 6845 2821
rect 6879 2787 6889 2821
rect 6835 2753 6889 2787
rect 6835 2719 6845 2753
rect 6879 2719 6889 2753
rect 6835 2707 6889 2719
rect 6919 2895 6973 2907
rect 6919 2861 6929 2895
rect 6963 2861 6973 2895
rect 6919 2827 6973 2861
rect 6919 2793 6929 2827
rect 6963 2793 6973 2827
rect 6919 2707 6973 2793
rect 7003 2889 7057 2907
rect 7003 2855 7013 2889
rect 7047 2855 7057 2889
rect 7003 2821 7057 2855
rect 7003 2787 7013 2821
rect 7047 2787 7057 2821
rect 7003 2753 7057 2787
rect 7003 2719 7013 2753
rect 7047 2719 7057 2753
rect 7003 2707 7057 2719
rect 7087 2895 7139 2907
rect 7087 2861 7097 2895
rect 7131 2861 7139 2895
rect 7087 2827 7139 2861
rect 7087 2793 7097 2827
rect 7131 2793 7139 2827
rect 7087 2707 7139 2793
rect 27 1753 79 1765
rect 27 1719 35 1753
rect 69 1719 79 1753
rect 27 1685 79 1719
rect 27 1651 35 1685
rect 69 1651 79 1685
rect 27 1617 79 1651
rect 27 1583 35 1617
rect 69 1583 79 1617
rect 27 1565 79 1583
rect 109 1753 161 1765
rect 109 1719 119 1753
rect 153 1726 161 1753
rect 2101 1753 2153 1765
rect 2101 1726 2109 1753
rect 153 1719 188 1726
rect 109 1685 188 1719
rect 109 1651 119 1685
rect 153 1651 188 1685
rect 109 1642 188 1651
rect 218 1642 291 1726
rect 321 1693 505 1726
rect 321 1659 355 1693
rect 389 1659 430 1693
rect 464 1659 505 1693
rect 321 1642 505 1659
rect 535 1642 577 1726
rect 607 1693 673 1726
rect 607 1659 627 1693
rect 661 1659 673 1693
rect 607 1642 673 1659
rect 703 1693 759 1726
rect 703 1659 713 1693
rect 747 1659 759 1693
rect 703 1642 759 1659
rect 1503 1693 1559 1726
rect 1503 1659 1515 1693
rect 1549 1659 1559 1693
rect 1503 1642 1559 1659
rect 1589 1693 1655 1726
rect 1589 1659 1601 1693
rect 1635 1659 1655 1693
rect 1589 1642 1655 1659
rect 1685 1642 1727 1726
rect 1757 1693 1941 1726
rect 1757 1659 1798 1693
rect 1832 1659 1873 1693
rect 1907 1659 1941 1693
rect 1757 1642 1941 1659
rect 1971 1642 2044 1726
rect 2074 1719 2109 1726
rect 2143 1719 2153 1753
rect 2074 1685 2153 1719
rect 2074 1651 2109 1685
rect 2143 1651 2153 1685
rect 2074 1642 2153 1651
rect 109 1617 161 1642
rect 109 1583 119 1617
rect 153 1583 161 1617
rect 109 1565 161 1583
rect 2101 1617 2153 1642
rect 2101 1583 2109 1617
rect 2143 1583 2153 1617
rect 2101 1565 2153 1583
rect 2183 1753 2235 1765
rect 2183 1719 2193 1753
rect 2227 1719 2235 1753
rect 2183 1685 2235 1719
rect 2183 1651 2193 1685
rect 2227 1651 2235 1685
rect 2183 1617 2235 1651
rect 2183 1583 2193 1617
rect 2227 1583 2235 1617
rect 2183 1565 2235 1583
rect 2419 1753 2471 1765
rect 2419 1719 2427 1753
rect 2461 1719 2471 1753
rect 2419 1685 2471 1719
rect 2419 1651 2427 1685
rect 2461 1651 2471 1685
rect 2419 1617 2471 1651
rect 2419 1583 2427 1617
rect 2461 1583 2471 1617
rect 2419 1565 2471 1583
rect 2501 1753 2553 1765
rect 2501 1719 2511 1753
rect 2545 1726 2553 1753
rect 4493 1753 4545 1765
rect 4493 1726 4501 1753
rect 2545 1719 2580 1726
rect 2501 1685 2580 1719
rect 2501 1651 2511 1685
rect 2545 1651 2580 1685
rect 2501 1642 2580 1651
rect 2610 1642 2683 1726
rect 2713 1693 2897 1726
rect 2713 1659 2747 1693
rect 2781 1659 2822 1693
rect 2856 1659 2897 1693
rect 2713 1642 2897 1659
rect 2927 1642 2969 1726
rect 2999 1693 3065 1726
rect 2999 1659 3019 1693
rect 3053 1659 3065 1693
rect 2999 1642 3065 1659
rect 3095 1693 3151 1726
rect 3095 1659 3105 1693
rect 3139 1659 3151 1693
rect 3095 1642 3151 1659
rect 3895 1693 3951 1726
rect 3895 1659 3907 1693
rect 3941 1659 3951 1693
rect 3895 1642 3951 1659
rect 3981 1693 4047 1726
rect 3981 1659 3993 1693
rect 4027 1659 4047 1693
rect 3981 1642 4047 1659
rect 4077 1642 4119 1726
rect 4149 1693 4333 1726
rect 4149 1659 4190 1693
rect 4224 1659 4265 1693
rect 4299 1659 4333 1693
rect 4149 1642 4333 1659
rect 4363 1642 4436 1726
rect 4466 1719 4501 1726
rect 4535 1719 4545 1753
rect 4466 1685 4545 1719
rect 4466 1651 4501 1685
rect 4535 1651 4545 1685
rect 4466 1642 4545 1651
rect 2501 1617 2553 1642
rect 2501 1583 2511 1617
rect 2545 1583 2553 1617
rect 2501 1565 2553 1583
rect 4493 1617 4545 1642
rect 4493 1583 4501 1617
rect 4535 1583 4545 1617
rect 4493 1565 4545 1583
rect 4575 1753 4627 1765
rect 4575 1719 4585 1753
rect 4619 1719 4627 1753
rect 4575 1685 4627 1719
rect 4575 1651 4585 1685
rect 4619 1651 4627 1685
rect 4575 1617 4627 1651
rect 4575 1583 4585 1617
rect 4619 1583 4627 1617
rect 4575 1565 4627 1583
rect 4811 1753 4863 1765
rect 4811 1719 4819 1753
rect 4853 1719 4863 1753
rect 4811 1685 4863 1719
rect 4811 1651 4819 1685
rect 4853 1651 4863 1685
rect 4811 1617 4863 1651
rect 4811 1583 4819 1617
rect 4853 1583 4863 1617
rect 4811 1565 4863 1583
rect 4893 1753 4945 1765
rect 4893 1719 4903 1753
rect 4937 1726 4945 1753
rect 6883 1753 6935 1765
rect 6883 1726 6891 1753
rect 4937 1719 4972 1726
rect 4893 1685 4972 1719
rect 4893 1651 4903 1685
rect 4937 1651 4972 1685
rect 4893 1642 4972 1651
rect 5002 1642 5075 1726
rect 5105 1693 5289 1726
rect 5105 1659 5139 1693
rect 5173 1659 5214 1693
rect 5248 1659 5289 1693
rect 5105 1642 5289 1659
rect 5319 1642 5361 1726
rect 5391 1693 5457 1726
rect 5391 1659 5411 1693
rect 5445 1659 5457 1693
rect 5391 1642 5457 1659
rect 5487 1693 5543 1726
rect 5487 1659 5497 1693
rect 5531 1659 5543 1693
rect 5487 1642 5543 1659
rect 6285 1693 6341 1726
rect 6285 1659 6297 1693
rect 6331 1659 6341 1693
rect 6285 1642 6341 1659
rect 6371 1693 6437 1726
rect 6371 1659 6383 1693
rect 6417 1659 6437 1693
rect 6371 1642 6437 1659
rect 6467 1642 6509 1726
rect 6539 1693 6723 1726
rect 6539 1659 6580 1693
rect 6614 1659 6655 1693
rect 6689 1659 6723 1693
rect 6539 1642 6723 1659
rect 6753 1642 6826 1726
rect 6856 1719 6891 1726
rect 6925 1719 6935 1753
rect 6856 1685 6935 1719
rect 6856 1651 6891 1685
rect 6925 1651 6935 1685
rect 6856 1642 6935 1651
rect 4893 1617 4945 1642
rect 4893 1583 4903 1617
rect 4937 1583 4945 1617
rect 4893 1565 4945 1583
rect 6883 1617 6935 1642
rect 6883 1583 6891 1617
rect 6925 1583 6935 1617
rect 6883 1565 6935 1583
rect 6965 1753 7017 1765
rect 6965 1719 6975 1753
rect 7009 1719 7017 1753
rect 6965 1685 7017 1719
rect 6965 1651 6975 1685
rect 7009 1651 7017 1685
rect 6965 1617 7017 1651
rect 6965 1583 6975 1617
rect 7009 1583 7017 1617
rect 6965 1565 7017 1583
rect 7203 1753 7255 1765
rect 7203 1719 7211 1753
rect 7245 1719 7255 1753
rect 7203 1685 7255 1719
rect 7203 1651 7211 1685
rect 7245 1651 7255 1685
rect 7203 1617 7255 1651
rect 7203 1583 7211 1617
rect 7245 1583 7255 1617
rect 7203 1565 7255 1583
rect 7285 1753 7337 1765
rect 7285 1719 7295 1753
rect 7329 1726 7337 1753
rect 9277 1753 9329 1765
rect 9277 1726 9285 1753
rect 7329 1719 7364 1726
rect 7285 1685 7364 1719
rect 7285 1651 7295 1685
rect 7329 1651 7364 1685
rect 7285 1642 7364 1651
rect 7394 1642 7467 1726
rect 7497 1693 7681 1726
rect 7497 1659 7531 1693
rect 7565 1659 7606 1693
rect 7640 1659 7681 1693
rect 7497 1642 7681 1659
rect 7711 1642 7753 1726
rect 7783 1693 7849 1726
rect 7783 1659 7803 1693
rect 7837 1659 7849 1693
rect 7783 1642 7849 1659
rect 7879 1693 7935 1726
rect 7879 1659 7889 1693
rect 7923 1659 7935 1693
rect 7879 1642 7935 1659
rect 8679 1693 8735 1726
rect 8679 1659 8691 1693
rect 8725 1659 8735 1693
rect 8679 1642 8735 1659
rect 8765 1693 8831 1726
rect 8765 1659 8777 1693
rect 8811 1659 8831 1693
rect 8765 1642 8831 1659
rect 8861 1642 8903 1726
rect 8933 1693 9117 1726
rect 8933 1659 8974 1693
rect 9008 1659 9049 1693
rect 9083 1659 9117 1693
rect 8933 1642 9117 1659
rect 9147 1642 9220 1726
rect 9250 1719 9285 1726
rect 9319 1719 9329 1753
rect 9250 1685 9329 1719
rect 9250 1651 9285 1685
rect 9319 1651 9329 1685
rect 9250 1642 9329 1651
rect 7285 1617 7337 1642
rect 7285 1583 7295 1617
rect 7329 1583 7337 1617
rect 7285 1565 7337 1583
rect 9277 1617 9329 1642
rect 9277 1583 9285 1617
rect 9319 1583 9329 1617
rect 9277 1565 9329 1583
rect 9359 1753 9411 1765
rect 9359 1719 9369 1753
rect 9403 1719 9411 1753
rect 9359 1685 9411 1719
rect 9359 1651 9369 1685
rect 9403 1651 9411 1685
rect 9359 1617 9411 1651
rect 9359 1583 9369 1617
rect 9403 1583 9411 1617
rect 9359 1565 9411 1583
rect 9595 1753 9647 1765
rect 9595 1719 9603 1753
rect 9637 1719 9647 1753
rect 9595 1685 9647 1719
rect 9595 1651 9603 1685
rect 9637 1651 9647 1685
rect 9595 1617 9647 1651
rect 9595 1583 9603 1617
rect 9637 1583 9647 1617
rect 9595 1565 9647 1583
rect 9677 1753 9729 1765
rect 9677 1719 9687 1753
rect 9721 1726 9729 1753
rect 11669 1753 11721 1765
rect 11669 1726 11677 1753
rect 9721 1719 9756 1726
rect 9677 1685 9756 1719
rect 9677 1651 9687 1685
rect 9721 1651 9756 1685
rect 9677 1642 9756 1651
rect 9786 1642 9859 1726
rect 9889 1693 10073 1726
rect 9889 1659 9923 1693
rect 9957 1659 9998 1693
rect 10032 1659 10073 1693
rect 9889 1642 10073 1659
rect 10103 1642 10145 1726
rect 10175 1693 10241 1726
rect 10175 1659 10195 1693
rect 10229 1659 10241 1693
rect 10175 1642 10241 1659
rect 10271 1693 10327 1726
rect 10271 1659 10281 1693
rect 10315 1659 10327 1693
rect 10271 1642 10327 1659
rect 11071 1693 11127 1726
rect 11071 1659 11083 1693
rect 11117 1659 11127 1693
rect 11071 1642 11127 1659
rect 11157 1693 11223 1726
rect 11157 1659 11169 1693
rect 11203 1659 11223 1693
rect 11157 1642 11223 1659
rect 11253 1642 11295 1726
rect 11325 1693 11509 1726
rect 11325 1659 11366 1693
rect 11400 1659 11441 1693
rect 11475 1659 11509 1693
rect 11325 1642 11509 1659
rect 11539 1642 11612 1726
rect 11642 1719 11677 1726
rect 11711 1719 11721 1753
rect 11642 1685 11721 1719
rect 11642 1651 11677 1685
rect 11711 1651 11721 1685
rect 11642 1642 11721 1651
rect 9677 1617 9729 1642
rect 9677 1583 9687 1617
rect 9721 1583 9729 1617
rect 9677 1565 9729 1583
rect 11669 1617 11721 1642
rect 11669 1583 11677 1617
rect 11711 1583 11721 1617
rect 11669 1565 11721 1583
rect 11751 1753 11803 1765
rect 11751 1719 11761 1753
rect 11795 1719 11803 1753
rect 11751 1685 11803 1719
rect 11751 1651 11761 1685
rect 11795 1651 11803 1685
rect 11751 1617 11803 1651
rect 11751 1583 11761 1617
rect 11795 1583 11803 1617
rect 11751 1565 11803 1583
rect 11987 1753 12039 1765
rect 11987 1719 11995 1753
rect 12029 1719 12039 1753
rect 11987 1685 12039 1719
rect 11987 1651 11995 1685
rect 12029 1651 12039 1685
rect 11987 1617 12039 1651
rect 11987 1583 11995 1617
rect 12029 1583 12039 1617
rect 11987 1565 12039 1583
rect 12069 1753 12121 1765
rect 12069 1719 12079 1753
rect 12113 1726 12121 1753
rect 14059 1753 14111 1765
rect 14059 1726 14067 1753
rect 12113 1719 12148 1726
rect 12069 1685 12148 1719
rect 12069 1651 12079 1685
rect 12113 1651 12148 1685
rect 12069 1642 12148 1651
rect 12178 1642 12251 1726
rect 12281 1693 12465 1726
rect 12281 1659 12315 1693
rect 12349 1659 12390 1693
rect 12424 1659 12465 1693
rect 12281 1642 12465 1659
rect 12495 1642 12537 1726
rect 12567 1693 12633 1726
rect 12567 1659 12587 1693
rect 12621 1659 12633 1693
rect 12567 1642 12633 1659
rect 12663 1693 12719 1726
rect 12663 1659 12673 1693
rect 12707 1659 12719 1693
rect 12663 1642 12719 1659
rect 13461 1693 13517 1726
rect 13461 1659 13473 1693
rect 13507 1659 13517 1693
rect 13461 1642 13517 1659
rect 13547 1693 13613 1726
rect 13547 1659 13559 1693
rect 13593 1659 13613 1693
rect 13547 1642 13613 1659
rect 13643 1642 13685 1726
rect 13715 1693 13899 1726
rect 13715 1659 13756 1693
rect 13790 1659 13831 1693
rect 13865 1659 13899 1693
rect 13715 1642 13899 1659
rect 13929 1642 14002 1726
rect 14032 1719 14067 1726
rect 14101 1719 14111 1753
rect 14032 1685 14111 1719
rect 14032 1651 14067 1685
rect 14101 1651 14111 1685
rect 14032 1642 14111 1651
rect 12069 1617 12121 1642
rect 12069 1583 12079 1617
rect 12113 1583 12121 1617
rect 12069 1565 12121 1583
rect 14059 1617 14111 1642
rect 14059 1583 14067 1617
rect 14101 1583 14111 1617
rect 14059 1565 14111 1583
rect 14141 1753 14193 1765
rect 14141 1719 14151 1753
rect 14185 1719 14193 1753
rect 14141 1685 14193 1719
rect 14141 1651 14151 1685
rect 14185 1651 14193 1685
rect 14141 1617 14193 1651
rect 14141 1583 14151 1617
rect 14185 1583 14193 1617
rect 14141 1565 14193 1583
rect 14379 1753 14431 1765
rect 14379 1719 14387 1753
rect 14421 1719 14431 1753
rect 14379 1685 14431 1719
rect 14379 1651 14387 1685
rect 14421 1651 14431 1685
rect 14379 1617 14431 1651
rect 14379 1583 14387 1617
rect 14421 1583 14431 1617
rect 14379 1565 14431 1583
rect 14461 1753 14513 1765
rect 14461 1719 14471 1753
rect 14505 1726 14513 1753
rect 16453 1753 16505 1765
rect 16453 1726 16461 1753
rect 14505 1719 14540 1726
rect 14461 1685 14540 1719
rect 14461 1651 14471 1685
rect 14505 1651 14540 1685
rect 14461 1642 14540 1651
rect 14570 1642 14643 1726
rect 14673 1693 14857 1726
rect 14673 1659 14707 1693
rect 14741 1659 14782 1693
rect 14816 1659 14857 1693
rect 14673 1642 14857 1659
rect 14887 1642 14929 1726
rect 14959 1693 15025 1726
rect 14959 1659 14979 1693
rect 15013 1659 15025 1693
rect 14959 1642 15025 1659
rect 15055 1693 15111 1726
rect 15055 1659 15065 1693
rect 15099 1659 15111 1693
rect 15055 1642 15111 1659
rect 15855 1693 15911 1726
rect 15855 1659 15867 1693
rect 15901 1659 15911 1693
rect 15855 1642 15911 1659
rect 15941 1693 16007 1726
rect 15941 1659 15953 1693
rect 15987 1659 16007 1693
rect 15941 1642 16007 1659
rect 16037 1642 16079 1726
rect 16109 1693 16293 1726
rect 16109 1659 16150 1693
rect 16184 1659 16225 1693
rect 16259 1659 16293 1693
rect 16109 1642 16293 1659
rect 16323 1642 16396 1726
rect 16426 1719 16461 1726
rect 16495 1719 16505 1753
rect 16426 1685 16505 1719
rect 16426 1651 16461 1685
rect 16495 1651 16505 1685
rect 16426 1642 16505 1651
rect 14461 1617 14513 1642
rect 14461 1583 14471 1617
rect 14505 1583 14513 1617
rect 14461 1565 14513 1583
rect 16453 1617 16505 1642
rect 16453 1583 16461 1617
rect 16495 1583 16505 1617
rect 16453 1565 16505 1583
rect 16535 1753 16587 1765
rect 16535 1719 16545 1753
rect 16579 1719 16587 1753
rect 16535 1685 16587 1719
rect 16535 1651 16545 1685
rect 16579 1651 16587 1685
rect 16535 1617 16587 1651
rect 16535 1583 16545 1617
rect 16579 1583 16587 1617
rect 16535 1565 16587 1583
rect 27 1057 79 1071
rect 27 1023 35 1057
rect 69 1023 79 1057
rect 27 989 79 1023
rect 27 955 35 989
rect 69 955 79 989
rect 27 943 79 955
rect 109 1041 163 1071
rect 109 1007 119 1041
rect 153 1007 163 1041
rect 109 943 163 1007
rect 193 1057 245 1071
rect 193 1023 203 1057
rect 237 1023 245 1057
rect 193 989 245 1023
rect 299 1041 351 1077
rect 299 1007 307 1041
rect 341 1007 351 1041
rect 299 993 351 1007
rect 381 1057 443 1077
rect 381 1023 391 1057
rect 425 1023 443 1057
rect 381 993 443 1023
rect 473 1064 527 1077
rect 473 1030 483 1064
rect 517 1030 527 1064
rect 473 993 527 1030
rect 557 993 647 1077
rect 677 1055 753 1077
rect 677 1021 697 1055
rect 731 1021 753 1055
rect 677 993 753 1021
rect 783 1039 861 1077
rect 783 1005 817 1039
rect 851 1005 861 1039
rect 783 993 861 1005
rect 193 955 203 989
rect 237 955 245 989
rect 193 943 245 955
rect 799 971 861 993
rect 799 937 817 971
rect 851 937 861 971
rect 799 909 861 937
rect 891 909 945 1077
rect 975 1065 1082 1077
rect 975 1031 991 1065
rect 1025 1031 1082 1065
rect 975 997 1082 1031
rect 975 963 991 997
rect 1025 963 1082 997
rect 975 909 1082 963
rect 1112 993 1226 1077
rect 1256 1064 1310 1077
rect 1256 1030 1266 1064
rect 1300 1030 1310 1064
rect 1256 993 1310 1030
rect 1340 993 1415 1077
rect 1445 1065 1536 1077
rect 1445 1031 1480 1065
rect 1514 1031 1536 1065
rect 1445 993 1536 1031
rect 1566 1039 1642 1077
rect 1566 1005 1588 1039
rect 1622 1005 1642 1039
rect 1566 993 1642 1005
rect 1112 909 1164 993
rect 1592 909 1642 993
rect 1672 909 1714 1077
rect 1744 1065 1796 1077
rect 1744 1031 1754 1065
rect 1788 1031 1796 1065
rect 1744 909 1796 1031
rect 1948 1065 2000 1077
rect 1948 1031 1956 1065
rect 1990 1031 2000 1065
rect 1948 1009 2000 1031
rect 1850 929 1903 1009
rect 1850 895 1858 929
rect 1892 895 1903 929
rect 1850 881 1903 895
rect 1933 881 2000 1009
rect 1950 877 2000 881
rect 2030 1028 2082 1077
rect 2233 1061 2283 1077
rect 2030 994 2040 1028
rect 2074 994 2082 1028
rect 2030 960 2082 994
rect 2030 926 2040 960
rect 2074 926 2082 960
rect 2136 1047 2188 1061
rect 2136 1013 2144 1047
rect 2178 1013 2188 1047
rect 2136 979 2188 1013
rect 2136 945 2144 979
rect 2178 945 2188 979
rect 2136 933 2188 945
rect 2218 1053 2283 1061
rect 2218 1019 2239 1053
rect 2273 1019 2283 1053
rect 2218 985 2283 1019
rect 2218 951 2239 985
rect 2273 951 2283 985
rect 2218 933 2283 951
rect 2030 877 2082 926
rect 2233 877 2283 933
rect 2313 1029 2365 1077
rect 2313 995 2323 1029
rect 2357 995 2365 1029
rect 2313 961 2365 995
rect 2313 927 2323 961
rect 2357 927 2365 961
rect 2419 1057 2471 1071
rect 2419 1023 2427 1057
rect 2461 1023 2471 1057
rect 2419 989 2471 1023
rect 2419 955 2427 989
rect 2461 955 2471 989
rect 2419 943 2471 955
rect 2501 1041 2555 1071
rect 2501 1007 2511 1041
rect 2545 1007 2555 1041
rect 2501 943 2555 1007
rect 2585 1057 2637 1071
rect 2585 1023 2595 1057
rect 2629 1023 2637 1057
rect 2585 989 2637 1023
rect 2691 1041 2743 1077
rect 2691 1007 2699 1041
rect 2733 1007 2743 1041
rect 2691 993 2743 1007
rect 2773 1057 2835 1077
rect 2773 1023 2783 1057
rect 2817 1023 2835 1057
rect 2773 993 2835 1023
rect 2865 1064 2919 1077
rect 2865 1030 2875 1064
rect 2909 1030 2919 1064
rect 2865 993 2919 1030
rect 2949 993 3039 1077
rect 3069 1055 3145 1077
rect 3069 1021 3089 1055
rect 3123 1021 3145 1055
rect 3069 993 3145 1021
rect 3175 1039 3253 1077
rect 3175 1005 3209 1039
rect 3243 1005 3253 1039
rect 3175 993 3253 1005
rect 2585 955 2595 989
rect 2629 955 2637 989
rect 2585 943 2637 955
rect 2313 877 2365 927
rect 3191 971 3253 993
rect 3191 937 3209 971
rect 3243 937 3253 971
rect 3191 909 3253 937
rect 3283 909 3337 1077
rect 3367 1065 3474 1077
rect 3367 1031 3383 1065
rect 3417 1031 3474 1065
rect 3367 997 3474 1031
rect 3367 963 3383 997
rect 3417 963 3474 997
rect 3367 909 3474 963
rect 3504 993 3618 1077
rect 3648 1064 3702 1077
rect 3648 1030 3658 1064
rect 3692 1030 3702 1064
rect 3648 993 3702 1030
rect 3732 993 3807 1077
rect 3837 1065 3928 1077
rect 3837 1031 3872 1065
rect 3906 1031 3928 1065
rect 3837 993 3928 1031
rect 3958 1039 4034 1077
rect 3958 1005 3980 1039
rect 4014 1005 4034 1039
rect 3958 993 4034 1005
rect 3504 909 3556 993
rect 3984 909 4034 993
rect 4064 909 4106 1077
rect 4136 1065 4188 1077
rect 4136 1031 4146 1065
rect 4180 1031 4188 1065
rect 4136 909 4188 1031
rect 4340 1065 4392 1077
rect 4340 1031 4348 1065
rect 4382 1031 4392 1065
rect 4340 1009 4392 1031
rect 4242 929 4295 1009
rect 4242 895 4250 929
rect 4284 895 4295 929
rect 4242 881 4295 895
rect 4325 881 4392 1009
rect 4342 877 4392 881
rect 4422 1028 4474 1077
rect 4625 1061 4675 1077
rect 4422 994 4432 1028
rect 4466 994 4474 1028
rect 4422 960 4474 994
rect 4422 926 4432 960
rect 4466 926 4474 960
rect 4528 1047 4580 1061
rect 4528 1013 4536 1047
rect 4570 1013 4580 1047
rect 4528 979 4580 1013
rect 4528 945 4536 979
rect 4570 945 4580 979
rect 4528 933 4580 945
rect 4610 1053 4675 1061
rect 4610 1019 4631 1053
rect 4665 1019 4675 1053
rect 4610 985 4675 1019
rect 4610 951 4631 985
rect 4665 951 4675 985
rect 4610 933 4675 951
rect 4422 877 4474 926
rect 4625 877 4675 933
rect 4705 1029 4757 1077
rect 4705 995 4715 1029
rect 4749 995 4757 1029
rect 4705 961 4757 995
rect 4705 927 4715 961
rect 4749 927 4757 961
rect 4811 1057 4863 1071
rect 4811 1023 4819 1057
rect 4853 1023 4863 1057
rect 4811 989 4863 1023
rect 4811 955 4819 989
rect 4853 955 4863 989
rect 4811 943 4863 955
rect 4893 1041 4947 1071
rect 4893 1007 4903 1041
rect 4937 1007 4947 1041
rect 4893 943 4947 1007
rect 4977 1057 5029 1071
rect 4977 1023 4987 1057
rect 5021 1023 5029 1057
rect 4977 989 5029 1023
rect 5083 1041 5135 1077
rect 5083 1007 5091 1041
rect 5125 1007 5135 1041
rect 5083 993 5135 1007
rect 5165 1057 5227 1077
rect 5165 1023 5175 1057
rect 5209 1023 5227 1057
rect 5165 993 5227 1023
rect 5257 1064 5311 1077
rect 5257 1030 5267 1064
rect 5301 1030 5311 1064
rect 5257 993 5311 1030
rect 5341 993 5431 1077
rect 5461 1055 5537 1077
rect 5461 1021 5481 1055
rect 5515 1021 5537 1055
rect 5461 993 5537 1021
rect 5567 1039 5645 1077
rect 5567 1005 5601 1039
rect 5635 1005 5645 1039
rect 5567 993 5645 1005
rect 4977 955 4987 989
rect 5021 955 5029 989
rect 4977 943 5029 955
rect 4705 877 4757 927
rect 5583 971 5645 993
rect 5583 937 5601 971
rect 5635 937 5645 971
rect 5583 909 5645 937
rect 5675 909 5729 1077
rect 5759 1065 5866 1077
rect 5759 1031 5775 1065
rect 5809 1031 5866 1065
rect 5759 997 5866 1031
rect 5759 963 5775 997
rect 5809 963 5866 997
rect 5759 909 5866 963
rect 5896 993 6010 1077
rect 6040 1064 6094 1077
rect 6040 1030 6050 1064
rect 6084 1030 6094 1064
rect 6040 993 6094 1030
rect 6124 993 6199 1077
rect 6229 1065 6320 1077
rect 6229 1031 6264 1065
rect 6298 1031 6320 1065
rect 6229 993 6320 1031
rect 6350 1039 6426 1077
rect 6350 1005 6372 1039
rect 6406 1005 6426 1039
rect 6350 993 6426 1005
rect 5896 909 5948 993
rect 6376 909 6426 993
rect 6456 909 6498 1077
rect 6528 1065 6580 1077
rect 6528 1031 6538 1065
rect 6572 1031 6580 1065
rect 6528 909 6580 1031
rect 6732 1065 6784 1077
rect 6732 1031 6740 1065
rect 6774 1031 6784 1065
rect 6732 1009 6784 1031
rect 6634 929 6687 1009
rect 6634 895 6642 929
rect 6676 895 6687 929
rect 6634 881 6687 895
rect 6717 881 6784 1009
rect 6734 877 6784 881
rect 6814 1028 6866 1077
rect 7017 1061 7067 1077
rect 6814 994 6824 1028
rect 6858 994 6866 1028
rect 6814 960 6866 994
rect 6814 926 6824 960
rect 6858 926 6866 960
rect 6920 1047 6972 1061
rect 6920 1013 6928 1047
rect 6962 1013 6972 1047
rect 6920 979 6972 1013
rect 6920 945 6928 979
rect 6962 945 6972 979
rect 6920 933 6972 945
rect 7002 1053 7067 1061
rect 7002 1019 7023 1053
rect 7057 1019 7067 1053
rect 7002 985 7067 1019
rect 7002 951 7023 985
rect 7057 951 7067 985
rect 7002 933 7067 951
rect 6814 877 6866 926
rect 7017 877 7067 933
rect 7097 1029 7149 1077
rect 7097 995 7107 1029
rect 7141 995 7149 1029
rect 7097 961 7149 995
rect 7097 927 7107 961
rect 7141 927 7149 961
rect 7203 1057 7255 1071
rect 7203 1023 7211 1057
rect 7245 1023 7255 1057
rect 7203 989 7255 1023
rect 7203 955 7211 989
rect 7245 955 7255 989
rect 7203 943 7255 955
rect 7285 1041 7339 1071
rect 7285 1007 7295 1041
rect 7329 1007 7339 1041
rect 7285 943 7339 1007
rect 7369 1057 7421 1071
rect 7369 1023 7379 1057
rect 7413 1023 7421 1057
rect 7369 989 7421 1023
rect 7475 1041 7527 1077
rect 7475 1007 7483 1041
rect 7517 1007 7527 1041
rect 7475 993 7527 1007
rect 7557 1057 7619 1077
rect 7557 1023 7567 1057
rect 7601 1023 7619 1057
rect 7557 993 7619 1023
rect 7649 1064 7703 1077
rect 7649 1030 7659 1064
rect 7693 1030 7703 1064
rect 7649 993 7703 1030
rect 7733 993 7823 1077
rect 7853 1055 7929 1077
rect 7853 1021 7873 1055
rect 7907 1021 7929 1055
rect 7853 993 7929 1021
rect 7959 1039 8037 1077
rect 7959 1005 7993 1039
rect 8027 1005 8037 1039
rect 7959 993 8037 1005
rect 7369 955 7379 989
rect 7413 955 7421 989
rect 7369 943 7421 955
rect 7097 877 7149 927
rect 7975 971 8037 993
rect 7975 937 7993 971
rect 8027 937 8037 971
rect 7975 909 8037 937
rect 8067 909 8121 1077
rect 8151 1065 8258 1077
rect 8151 1031 8167 1065
rect 8201 1031 8258 1065
rect 8151 997 8258 1031
rect 8151 963 8167 997
rect 8201 963 8258 997
rect 8151 909 8258 963
rect 8288 993 8402 1077
rect 8432 1064 8486 1077
rect 8432 1030 8442 1064
rect 8476 1030 8486 1064
rect 8432 993 8486 1030
rect 8516 993 8591 1077
rect 8621 1065 8712 1077
rect 8621 1031 8656 1065
rect 8690 1031 8712 1065
rect 8621 993 8712 1031
rect 8742 1039 8818 1077
rect 8742 1005 8764 1039
rect 8798 1005 8818 1039
rect 8742 993 8818 1005
rect 8288 909 8340 993
rect 8768 909 8818 993
rect 8848 909 8890 1077
rect 8920 1065 8972 1077
rect 8920 1031 8930 1065
rect 8964 1031 8972 1065
rect 8920 909 8972 1031
rect 9124 1065 9176 1077
rect 9124 1031 9132 1065
rect 9166 1031 9176 1065
rect 9124 1009 9176 1031
rect 9026 929 9079 1009
rect 9026 895 9034 929
rect 9068 895 9079 929
rect 9026 881 9079 895
rect 9109 881 9176 1009
rect 9126 877 9176 881
rect 9206 1028 9258 1077
rect 9409 1061 9459 1077
rect 9206 994 9216 1028
rect 9250 994 9258 1028
rect 9206 960 9258 994
rect 9206 926 9216 960
rect 9250 926 9258 960
rect 9312 1047 9364 1061
rect 9312 1013 9320 1047
rect 9354 1013 9364 1047
rect 9312 979 9364 1013
rect 9312 945 9320 979
rect 9354 945 9364 979
rect 9312 933 9364 945
rect 9394 1053 9459 1061
rect 9394 1019 9415 1053
rect 9449 1019 9459 1053
rect 9394 985 9459 1019
rect 9394 951 9415 985
rect 9449 951 9459 985
rect 9394 933 9459 951
rect 9206 877 9258 926
rect 9409 877 9459 933
rect 9489 1029 9541 1077
rect 9489 995 9499 1029
rect 9533 995 9541 1029
rect 9489 961 9541 995
rect 9489 927 9499 961
rect 9533 927 9541 961
rect 9595 1057 9647 1071
rect 9595 1023 9603 1057
rect 9637 1023 9647 1057
rect 9595 989 9647 1023
rect 9595 955 9603 989
rect 9637 955 9647 989
rect 9595 943 9647 955
rect 9677 1041 9731 1071
rect 9677 1007 9687 1041
rect 9721 1007 9731 1041
rect 9677 943 9731 1007
rect 9761 1057 9813 1071
rect 9761 1023 9771 1057
rect 9805 1023 9813 1057
rect 9761 989 9813 1023
rect 9867 1041 9919 1077
rect 9867 1007 9875 1041
rect 9909 1007 9919 1041
rect 9867 993 9919 1007
rect 9949 1057 10011 1077
rect 9949 1023 9959 1057
rect 9993 1023 10011 1057
rect 9949 993 10011 1023
rect 10041 1064 10095 1077
rect 10041 1030 10051 1064
rect 10085 1030 10095 1064
rect 10041 993 10095 1030
rect 10125 993 10215 1077
rect 10245 1055 10321 1077
rect 10245 1021 10265 1055
rect 10299 1021 10321 1055
rect 10245 993 10321 1021
rect 10351 1039 10429 1077
rect 10351 1005 10385 1039
rect 10419 1005 10429 1039
rect 10351 993 10429 1005
rect 9761 955 9771 989
rect 9805 955 9813 989
rect 9761 943 9813 955
rect 9489 877 9541 927
rect 10367 971 10429 993
rect 10367 937 10385 971
rect 10419 937 10429 971
rect 10367 909 10429 937
rect 10459 909 10513 1077
rect 10543 1065 10650 1077
rect 10543 1031 10559 1065
rect 10593 1031 10650 1065
rect 10543 997 10650 1031
rect 10543 963 10559 997
rect 10593 963 10650 997
rect 10543 909 10650 963
rect 10680 993 10794 1077
rect 10824 1064 10878 1077
rect 10824 1030 10834 1064
rect 10868 1030 10878 1064
rect 10824 993 10878 1030
rect 10908 993 10983 1077
rect 11013 1065 11104 1077
rect 11013 1031 11048 1065
rect 11082 1031 11104 1065
rect 11013 993 11104 1031
rect 11134 1039 11210 1077
rect 11134 1005 11156 1039
rect 11190 1005 11210 1039
rect 11134 993 11210 1005
rect 10680 909 10732 993
rect 11160 909 11210 993
rect 11240 909 11282 1077
rect 11312 1065 11364 1077
rect 11312 1031 11322 1065
rect 11356 1031 11364 1065
rect 11312 909 11364 1031
rect 11516 1065 11568 1077
rect 11516 1031 11524 1065
rect 11558 1031 11568 1065
rect 11516 1009 11568 1031
rect 11418 929 11471 1009
rect 11418 895 11426 929
rect 11460 895 11471 929
rect 11418 881 11471 895
rect 11501 881 11568 1009
rect 11518 877 11568 881
rect 11598 1028 11650 1077
rect 11801 1061 11851 1077
rect 11598 994 11608 1028
rect 11642 994 11650 1028
rect 11598 960 11650 994
rect 11598 926 11608 960
rect 11642 926 11650 960
rect 11704 1047 11756 1061
rect 11704 1013 11712 1047
rect 11746 1013 11756 1047
rect 11704 979 11756 1013
rect 11704 945 11712 979
rect 11746 945 11756 979
rect 11704 933 11756 945
rect 11786 1053 11851 1061
rect 11786 1019 11807 1053
rect 11841 1019 11851 1053
rect 11786 985 11851 1019
rect 11786 951 11807 985
rect 11841 951 11851 985
rect 11786 933 11851 951
rect 11598 877 11650 926
rect 11801 877 11851 933
rect 11881 1029 11933 1077
rect 11881 995 11891 1029
rect 11925 995 11933 1029
rect 11881 961 11933 995
rect 11881 927 11891 961
rect 11925 927 11933 961
rect 11987 1057 12039 1071
rect 11987 1023 11995 1057
rect 12029 1023 12039 1057
rect 11987 989 12039 1023
rect 11987 955 11995 989
rect 12029 955 12039 989
rect 11987 943 12039 955
rect 12069 1041 12123 1071
rect 12069 1007 12079 1041
rect 12113 1007 12123 1041
rect 12069 943 12123 1007
rect 12153 1057 12205 1071
rect 12153 1023 12163 1057
rect 12197 1023 12205 1057
rect 12153 989 12205 1023
rect 12259 1041 12311 1077
rect 12259 1007 12267 1041
rect 12301 1007 12311 1041
rect 12259 993 12311 1007
rect 12341 1057 12403 1077
rect 12341 1023 12351 1057
rect 12385 1023 12403 1057
rect 12341 993 12403 1023
rect 12433 1064 12487 1077
rect 12433 1030 12443 1064
rect 12477 1030 12487 1064
rect 12433 993 12487 1030
rect 12517 993 12607 1077
rect 12637 1055 12713 1077
rect 12637 1021 12657 1055
rect 12691 1021 12713 1055
rect 12637 993 12713 1021
rect 12743 1039 12821 1077
rect 12743 1005 12777 1039
rect 12811 1005 12821 1039
rect 12743 993 12821 1005
rect 12153 955 12163 989
rect 12197 955 12205 989
rect 12153 943 12205 955
rect 11881 877 11933 927
rect 12759 971 12821 993
rect 12759 937 12777 971
rect 12811 937 12821 971
rect 12759 909 12821 937
rect 12851 909 12905 1077
rect 12935 1065 13042 1077
rect 12935 1031 12951 1065
rect 12985 1031 13042 1065
rect 12935 997 13042 1031
rect 12935 963 12951 997
rect 12985 963 13042 997
rect 12935 909 13042 963
rect 13072 993 13186 1077
rect 13216 1064 13270 1077
rect 13216 1030 13226 1064
rect 13260 1030 13270 1064
rect 13216 993 13270 1030
rect 13300 993 13375 1077
rect 13405 1065 13496 1077
rect 13405 1031 13440 1065
rect 13474 1031 13496 1065
rect 13405 993 13496 1031
rect 13526 1039 13602 1077
rect 13526 1005 13548 1039
rect 13582 1005 13602 1039
rect 13526 993 13602 1005
rect 13072 909 13124 993
rect 13552 909 13602 993
rect 13632 909 13674 1077
rect 13704 1065 13756 1077
rect 13704 1031 13714 1065
rect 13748 1031 13756 1065
rect 13704 909 13756 1031
rect 13908 1065 13960 1077
rect 13908 1031 13916 1065
rect 13950 1031 13960 1065
rect 13908 1009 13960 1031
rect 13810 929 13863 1009
rect 13810 895 13818 929
rect 13852 895 13863 929
rect 13810 881 13863 895
rect 13893 881 13960 1009
rect 13910 877 13960 881
rect 13990 1028 14042 1077
rect 14193 1061 14243 1077
rect 13990 994 14000 1028
rect 14034 994 14042 1028
rect 13990 960 14042 994
rect 13990 926 14000 960
rect 14034 926 14042 960
rect 14096 1047 14148 1061
rect 14096 1013 14104 1047
rect 14138 1013 14148 1047
rect 14096 979 14148 1013
rect 14096 945 14104 979
rect 14138 945 14148 979
rect 14096 933 14148 945
rect 14178 1053 14243 1061
rect 14178 1019 14199 1053
rect 14233 1019 14243 1053
rect 14178 985 14243 1019
rect 14178 951 14199 985
rect 14233 951 14243 985
rect 14178 933 14243 951
rect 13990 877 14042 926
rect 14193 877 14243 933
rect 14273 1029 14325 1077
rect 14273 995 14283 1029
rect 14317 995 14325 1029
rect 14273 961 14325 995
rect 14273 927 14283 961
rect 14317 927 14325 961
rect 14379 1057 14431 1071
rect 14379 1023 14387 1057
rect 14421 1023 14431 1057
rect 14379 989 14431 1023
rect 14379 955 14387 989
rect 14421 955 14431 989
rect 14379 943 14431 955
rect 14461 1041 14515 1071
rect 14461 1007 14471 1041
rect 14505 1007 14515 1041
rect 14461 943 14515 1007
rect 14545 1057 14597 1071
rect 14545 1023 14555 1057
rect 14589 1023 14597 1057
rect 14545 989 14597 1023
rect 14651 1041 14703 1077
rect 14651 1007 14659 1041
rect 14693 1007 14703 1041
rect 14651 993 14703 1007
rect 14733 1057 14795 1077
rect 14733 1023 14743 1057
rect 14777 1023 14795 1057
rect 14733 993 14795 1023
rect 14825 1064 14879 1077
rect 14825 1030 14835 1064
rect 14869 1030 14879 1064
rect 14825 993 14879 1030
rect 14909 993 14999 1077
rect 15029 1055 15105 1077
rect 15029 1021 15049 1055
rect 15083 1021 15105 1055
rect 15029 993 15105 1021
rect 15135 1039 15213 1077
rect 15135 1005 15169 1039
rect 15203 1005 15213 1039
rect 15135 993 15213 1005
rect 14545 955 14555 989
rect 14589 955 14597 989
rect 14545 943 14597 955
rect 14273 877 14325 927
rect 15151 971 15213 993
rect 15151 937 15169 971
rect 15203 937 15213 971
rect 15151 909 15213 937
rect 15243 909 15297 1077
rect 15327 1065 15434 1077
rect 15327 1031 15343 1065
rect 15377 1031 15434 1065
rect 15327 997 15434 1031
rect 15327 963 15343 997
rect 15377 963 15434 997
rect 15327 909 15434 963
rect 15464 993 15578 1077
rect 15608 1064 15662 1077
rect 15608 1030 15618 1064
rect 15652 1030 15662 1064
rect 15608 993 15662 1030
rect 15692 993 15767 1077
rect 15797 1065 15888 1077
rect 15797 1031 15832 1065
rect 15866 1031 15888 1065
rect 15797 993 15888 1031
rect 15918 1039 15994 1077
rect 15918 1005 15940 1039
rect 15974 1005 15994 1039
rect 15918 993 15994 1005
rect 15464 909 15516 993
rect 15944 909 15994 993
rect 16024 909 16066 1077
rect 16096 1065 16148 1077
rect 16096 1031 16106 1065
rect 16140 1031 16148 1065
rect 16096 909 16148 1031
rect 16300 1065 16352 1077
rect 16300 1031 16308 1065
rect 16342 1031 16352 1065
rect 16300 1009 16352 1031
rect 16202 929 16255 1009
rect 16202 895 16210 929
rect 16244 895 16255 929
rect 16202 881 16255 895
rect 16285 881 16352 1009
rect 16302 877 16352 881
rect 16382 1028 16434 1077
rect 16585 1061 16635 1077
rect 16382 994 16392 1028
rect 16426 994 16434 1028
rect 16382 960 16434 994
rect 16382 926 16392 960
rect 16426 926 16434 960
rect 16488 1047 16540 1061
rect 16488 1013 16496 1047
rect 16530 1013 16540 1047
rect 16488 979 16540 1013
rect 16488 945 16496 979
rect 16530 945 16540 979
rect 16488 933 16540 945
rect 16570 1053 16635 1061
rect 16570 1019 16591 1053
rect 16625 1019 16635 1053
rect 16570 985 16635 1019
rect 16570 951 16591 985
rect 16625 951 16635 985
rect 16570 933 16635 951
rect 16382 877 16434 926
rect 16585 877 16635 933
rect 16665 1029 16717 1077
rect 16665 995 16675 1029
rect 16709 995 16717 1029
rect 16665 961 16717 995
rect 16665 927 16675 961
rect 16709 927 16717 961
rect 16665 877 16717 927
rect 27 340 79 388
rect 27 306 35 340
rect 69 306 79 340
rect 27 272 79 306
rect 27 238 35 272
rect 69 238 79 272
rect 27 188 79 238
rect 109 372 159 388
rect 109 364 174 372
rect 109 330 119 364
rect 153 330 174 364
rect 109 296 174 330
rect 109 262 119 296
rect 153 262 174 296
rect 109 244 174 262
rect 204 358 256 372
rect 204 324 214 358
rect 248 324 256 358
rect 204 290 256 324
rect 204 256 214 290
rect 248 256 256 290
rect 204 244 256 256
rect 310 339 362 388
rect 310 305 318 339
rect 352 305 362 339
rect 310 271 362 305
rect 109 188 159 244
rect 310 237 318 271
rect 352 237 362 271
rect 310 188 362 237
rect 392 376 444 388
rect 392 342 402 376
rect 436 342 444 376
rect 596 376 648 388
rect 392 320 444 342
rect 596 342 604 376
rect 638 342 648 376
rect 392 192 459 320
rect 489 240 542 320
rect 489 206 500 240
rect 534 206 542 240
rect 596 220 648 342
rect 678 220 720 388
rect 750 350 826 388
rect 750 316 770 350
rect 804 316 826 350
rect 750 304 826 316
rect 856 376 947 388
rect 856 342 878 376
rect 912 342 947 376
rect 856 304 947 342
rect 977 304 1052 388
rect 1082 375 1136 388
rect 1082 341 1092 375
rect 1126 341 1136 375
rect 1082 304 1136 341
rect 1166 304 1280 388
rect 750 220 800 304
rect 489 192 542 206
rect 392 188 442 192
rect 1228 220 1280 304
rect 1310 376 1417 388
rect 1310 342 1367 376
rect 1401 342 1417 376
rect 1310 308 1417 342
rect 1310 274 1367 308
rect 1401 274 1417 308
rect 1310 220 1417 274
rect 1447 220 1501 388
rect 1531 350 1609 388
rect 1531 316 1541 350
rect 1575 316 1609 350
rect 1531 304 1609 316
rect 1639 366 1715 388
rect 1639 332 1661 366
rect 1695 332 1715 366
rect 1639 304 1715 332
rect 1745 304 1835 388
rect 1865 375 1919 388
rect 1865 341 1875 375
rect 1909 341 1919 375
rect 1865 304 1919 341
rect 1949 368 2011 388
rect 1949 334 1967 368
rect 2001 334 2011 368
rect 1949 304 2011 334
rect 2041 352 2093 388
rect 2041 318 2051 352
rect 2085 318 2093 352
rect 2041 304 2093 318
rect 2147 368 2199 382
rect 2147 334 2155 368
rect 2189 334 2199 368
rect 1531 282 1593 304
rect 1531 248 1541 282
rect 1575 248 1593 282
rect 1531 220 1593 248
rect 2147 300 2199 334
rect 2147 266 2155 300
rect 2189 266 2199 300
rect 2147 254 2199 266
rect 2229 352 2283 382
rect 2229 318 2239 352
rect 2273 318 2283 352
rect 2229 254 2283 318
rect 2313 368 2365 382
rect 2313 334 2323 368
rect 2357 334 2365 368
rect 2313 300 2365 334
rect 2313 266 2323 300
rect 2357 266 2365 300
rect 2313 254 2365 266
rect 2419 340 2471 388
rect 2419 306 2427 340
rect 2461 306 2471 340
rect 2419 272 2471 306
rect 2419 238 2427 272
rect 2461 238 2471 272
rect 2419 188 2471 238
rect 2501 372 2551 388
rect 2501 364 2566 372
rect 2501 330 2511 364
rect 2545 330 2566 364
rect 2501 296 2566 330
rect 2501 262 2511 296
rect 2545 262 2566 296
rect 2501 244 2566 262
rect 2596 358 2648 372
rect 2596 324 2606 358
rect 2640 324 2648 358
rect 2596 290 2648 324
rect 2596 256 2606 290
rect 2640 256 2648 290
rect 2596 244 2648 256
rect 2702 339 2754 388
rect 2702 305 2710 339
rect 2744 305 2754 339
rect 2702 271 2754 305
rect 2501 188 2551 244
rect 2702 237 2710 271
rect 2744 237 2754 271
rect 2702 188 2754 237
rect 2784 376 2836 388
rect 2784 342 2794 376
rect 2828 342 2836 376
rect 2988 376 3040 388
rect 2784 320 2836 342
rect 2988 342 2996 376
rect 3030 342 3040 376
rect 2784 192 2851 320
rect 2881 240 2934 320
rect 2881 206 2892 240
rect 2926 206 2934 240
rect 2988 220 3040 342
rect 3070 220 3112 388
rect 3142 350 3218 388
rect 3142 316 3162 350
rect 3196 316 3218 350
rect 3142 304 3218 316
rect 3248 376 3339 388
rect 3248 342 3270 376
rect 3304 342 3339 376
rect 3248 304 3339 342
rect 3369 304 3444 388
rect 3474 375 3528 388
rect 3474 341 3484 375
rect 3518 341 3528 375
rect 3474 304 3528 341
rect 3558 304 3672 388
rect 3142 220 3192 304
rect 2881 192 2934 206
rect 2784 188 2834 192
rect 3620 220 3672 304
rect 3702 376 3809 388
rect 3702 342 3759 376
rect 3793 342 3809 376
rect 3702 308 3809 342
rect 3702 274 3759 308
rect 3793 274 3809 308
rect 3702 220 3809 274
rect 3839 220 3893 388
rect 3923 350 4001 388
rect 3923 316 3933 350
rect 3967 316 4001 350
rect 3923 304 4001 316
rect 4031 366 4107 388
rect 4031 332 4053 366
rect 4087 332 4107 366
rect 4031 304 4107 332
rect 4137 304 4227 388
rect 4257 375 4311 388
rect 4257 341 4267 375
rect 4301 341 4311 375
rect 4257 304 4311 341
rect 4341 368 4403 388
rect 4341 334 4359 368
rect 4393 334 4403 368
rect 4341 304 4403 334
rect 4433 352 4485 388
rect 4433 318 4443 352
rect 4477 318 4485 352
rect 4433 304 4485 318
rect 4539 368 4591 382
rect 4539 334 4547 368
rect 4581 334 4591 368
rect 3923 282 3985 304
rect 3923 248 3933 282
rect 3967 248 3985 282
rect 3923 220 3985 248
rect 4539 300 4591 334
rect 4539 266 4547 300
rect 4581 266 4591 300
rect 4539 254 4591 266
rect 4621 352 4675 382
rect 4621 318 4631 352
rect 4665 318 4675 352
rect 4621 254 4675 318
rect 4705 368 4757 382
rect 4705 334 4715 368
rect 4749 334 4757 368
rect 4705 300 4757 334
rect 4705 266 4715 300
rect 4749 266 4757 300
rect 4705 254 4757 266
rect 4811 340 4863 388
rect 4811 306 4819 340
rect 4853 306 4863 340
rect 4811 272 4863 306
rect 4811 238 4819 272
rect 4853 238 4863 272
rect 4811 188 4863 238
rect 4893 372 4943 388
rect 4893 364 4958 372
rect 4893 330 4903 364
rect 4937 330 4958 364
rect 4893 296 4958 330
rect 4893 262 4903 296
rect 4937 262 4958 296
rect 4893 244 4958 262
rect 4988 358 5040 372
rect 4988 324 4998 358
rect 5032 324 5040 358
rect 4988 290 5040 324
rect 4988 256 4998 290
rect 5032 256 5040 290
rect 4988 244 5040 256
rect 5094 339 5146 388
rect 5094 305 5102 339
rect 5136 305 5146 339
rect 5094 271 5146 305
rect 4893 188 4943 244
rect 5094 237 5102 271
rect 5136 237 5146 271
rect 5094 188 5146 237
rect 5176 376 5228 388
rect 5176 342 5186 376
rect 5220 342 5228 376
rect 5380 376 5432 388
rect 5176 320 5228 342
rect 5380 342 5388 376
rect 5422 342 5432 376
rect 5176 192 5243 320
rect 5273 240 5326 320
rect 5273 206 5284 240
rect 5318 206 5326 240
rect 5380 220 5432 342
rect 5462 220 5504 388
rect 5534 350 5610 388
rect 5534 316 5554 350
rect 5588 316 5610 350
rect 5534 304 5610 316
rect 5640 376 5731 388
rect 5640 342 5662 376
rect 5696 342 5731 376
rect 5640 304 5731 342
rect 5761 304 5836 388
rect 5866 375 5920 388
rect 5866 341 5876 375
rect 5910 341 5920 375
rect 5866 304 5920 341
rect 5950 304 6064 388
rect 5534 220 5584 304
rect 5273 192 5326 206
rect 5176 188 5226 192
rect 6012 220 6064 304
rect 6094 376 6201 388
rect 6094 342 6151 376
rect 6185 342 6201 376
rect 6094 308 6201 342
rect 6094 274 6151 308
rect 6185 274 6201 308
rect 6094 220 6201 274
rect 6231 220 6285 388
rect 6315 350 6393 388
rect 6315 316 6325 350
rect 6359 316 6393 350
rect 6315 304 6393 316
rect 6423 366 6499 388
rect 6423 332 6445 366
rect 6479 332 6499 366
rect 6423 304 6499 332
rect 6529 304 6619 388
rect 6649 375 6703 388
rect 6649 341 6659 375
rect 6693 341 6703 375
rect 6649 304 6703 341
rect 6733 368 6795 388
rect 6733 334 6751 368
rect 6785 334 6795 368
rect 6733 304 6795 334
rect 6825 352 6877 388
rect 6825 318 6835 352
rect 6869 318 6877 352
rect 6825 304 6877 318
rect 6931 368 6983 382
rect 6931 334 6939 368
rect 6973 334 6983 368
rect 6315 282 6377 304
rect 6315 248 6325 282
rect 6359 248 6377 282
rect 6315 220 6377 248
rect 6931 300 6983 334
rect 6931 266 6939 300
rect 6973 266 6983 300
rect 6931 254 6983 266
rect 7013 352 7067 382
rect 7013 318 7023 352
rect 7057 318 7067 352
rect 7013 254 7067 318
rect 7097 368 7149 382
rect 7097 334 7107 368
rect 7141 334 7149 368
rect 7097 300 7149 334
rect 7097 266 7107 300
rect 7141 266 7149 300
rect 7097 254 7149 266
rect 7203 340 7255 388
rect 7203 306 7211 340
rect 7245 306 7255 340
rect 7203 272 7255 306
rect 7203 238 7211 272
rect 7245 238 7255 272
rect 7203 188 7255 238
rect 7285 372 7335 388
rect 7285 364 7350 372
rect 7285 330 7295 364
rect 7329 330 7350 364
rect 7285 296 7350 330
rect 7285 262 7295 296
rect 7329 262 7350 296
rect 7285 244 7350 262
rect 7380 358 7432 372
rect 7380 324 7390 358
rect 7424 324 7432 358
rect 7380 290 7432 324
rect 7380 256 7390 290
rect 7424 256 7432 290
rect 7380 244 7432 256
rect 7486 339 7538 388
rect 7486 305 7494 339
rect 7528 305 7538 339
rect 7486 271 7538 305
rect 7285 188 7335 244
rect 7486 237 7494 271
rect 7528 237 7538 271
rect 7486 188 7538 237
rect 7568 376 7620 388
rect 7568 342 7578 376
rect 7612 342 7620 376
rect 7772 376 7824 388
rect 7568 320 7620 342
rect 7772 342 7780 376
rect 7814 342 7824 376
rect 7568 192 7635 320
rect 7665 240 7718 320
rect 7665 206 7676 240
rect 7710 206 7718 240
rect 7772 220 7824 342
rect 7854 220 7896 388
rect 7926 350 8002 388
rect 7926 316 7946 350
rect 7980 316 8002 350
rect 7926 304 8002 316
rect 8032 376 8123 388
rect 8032 342 8054 376
rect 8088 342 8123 376
rect 8032 304 8123 342
rect 8153 304 8228 388
rect 8258 375 8312 388
rect 8258 341 8268 375
rect 8302 341 8312 375
rect 8258 304 8312 341
rect 8342 304 8456 388
rect 7926 220 7976 304
rect 7665 192 7718 206
rect 7568 188 7618 192
rect 8404 220 8456 304
rect 8486 376 8593 388
rect 8486 342 8543 376
rect 8577 342 8593 376
rect 8486 308 8593 342
rect 8486 274 8543 308
rect 8577 274 8593 308
rect 8486 220 8593 274
rect 8623 220 8677 388
rect 8707 350 8785 388
rect 8707 316 8717 350
rect 8751 316 8785 350
rect 8707 304 8785 316
rect 8815 366 8891 388
rect 8815 332 8837 366
rect 8871 332 8891 366
rect 8815 304 8891 332
rect 8921 304 9011 388
rect 9041 375 9095 388
rect 9041 341 9051 375
rect 9085 341 9095 375
rect 9041 304 9095 341
rect 9125 368 9187 388
rect 9125 334 9143 368
rect 9177 334 9187 368
rect 9125 304 9187 334
rect 9217 352 9269 388
rect 9217 318 9227 352
rect 9261 318 9269 352
rect 9217 304 9269 318
rect 9323 368 9375 382
rect 9323 334 9331 368
rect 9365 334 9375 368
rect 8707 282 8769 304
rect 8707 248 8717 282
rect 8751 248 8769 282
rect 8707 220 8769 248
rect 9323 300 9375 334
rect 9323 266 9331 300
rect 9365 266 9375 300
rect 9323 254 9375 266
rect 9405 352 9459 382
rect 9405 318 9415 352
rect 9449 318 9459 352
rect 9405 254 9459 318
rect 9489 368 9541 382
rect 9489 334 9499 368
rect 9533 334 9541 368
rect 9489 300 9541 334
rect 9489 266 9499 300
rect 9533 266 9541 300
rect 9489 254 9541 266
rect 9595 340 9647 388
rect 9595 306 9603 340
rect 9637 306 9647 340
rect 9595 272 9647 306
rect 9595 238 9603 272
rect 9637 238 9647 272
rect 9595 188 9647 238
rect 9677 372 9727 388
rect 9677 364 9742 372
rect 9677 330 9687 364
rect 9721 330 9742 364
rect 9677 296 9742 330
rect 9677 262 9687 296
rect 9721 262 9742 296
rect 9677 244 9742 262
rect 9772 358 9824 372
rect 9772 324 9782 358
rect 9816 324 9824 358
rect 9772 290 9824 324
rect 9772 256 9782 290
rect 9816 256 9824 290
rect 9772 244 9824 256
rect 9878 339 9930 388
rect 9878 305 9886 339
rect 9920 305 9930 339
rect 9878 271 9930 305
rect 9677 188 9727 244
rect 9878 237 9886 271
rect 9920 237 9930 271
rect 9878 188 9930 237
rect 9960 376 10012 388
rect 9960 342 9970 376
rect 10004 342 10012 376
rect 10164 376 10216 388
rect 9960 320 10012 342
rect 10164 342 10172 376
rect 10206 342 10216 376
rect 9960 192 10027 320
rect 10057 240 10110 320
rect 10057 206 10068 240
rect 10102 206 10110 240
rect 10164 220 10216 342
rect 10246 220 10288 388
rect 10318 350 10394 388
rect 10318 316 10338 350
rect 10372 316 10394 350
rect 10318 304 10394 316
rect 10424 376 10515 388
rect 10424 342 10446 376
rect 10480 342 10515 376
rect 10424 304 10515 342
rect 10545 304 10620 388
rect 10650 375 10704 388
rect 10650 341 10660 375
rect 10694 341 10704 375
rect 10650 304 10704 341
rect 10734 304 10848 388
rect 10318 220 10368 304
rect 10057 192 10110 206
rect 9960 188 10010 192
rect 10796 220 10848 304
rect 10878 376 10985 388
rect 10878 342 10935 376
rect 10969 342 10985 376
rect 10878 308 10985 342
rect 10878 274 10935 308
rect 10969 274 10985 308
rect 10878 220 10985 274
rect 11015 220 11069 388
rect 11099 350 11177 388
rect 11099 316 11109 350
rect 11143 316 11177 350
rect 11099 304 11177 316
rect 11207 366 11283 388
rect 11207 332 11229 366
rect 11263 332 11283 366
rect 11207 304 11283 332
rect 11313 304 11403 388
rect 11433 375 11487 388
rect 11433 341 11443 375
rect 11477 341 11487 375
rect 11433 304 11487 341
rect 11517 368 11579 388
rect 11517 334 11535 368
rect 11569 334 11579 368
rect 11517 304 11579 334
rect 11609 352 11661 388
rect 11609 318 11619 352
rect 11653 318 11661 352
rect 11609 304 11661 318
rect 11715 368 11767 382
rect 11715 334 11723 368
rect 11757 334 11767 368
rect 11099 282 11161 304
rect 11099 248 11109 282
rect 11143 248 11161 282
rect 11099 220 11161 248
rect 11715 300 11767 334
rect 11715 266 11723 300
rect 11757 266 11767 300
rect 11715 254 11767 266
rect 11797 352 11851 382
rect 11797 318 11807 352
rect 11841 318 11851 352
rect 11797 254 11851 318
rect 11881 368 11933 382
rect 11881 334 11891 368
rect 11925 334 11933 368
rect 11881 300 11933 334
rect 11881 266 11891 300
rect 11925 266 11933 300
rect 11881 254 11933 266
rect 11987 340 12039 388
rect 11987 306 11995 340
rect 12029 306 12039 340
rect 11987 272 12039 306
rect 11987 238 11995 272
rect 12029 238 12039 272
rect 11987 188 12039 238
rect 12069 372 12119 388
rect 12069 364 12134 372
rect 12069 330 12079 364
rect 12113 330 12134 364
rect 12069 296 12134 330
rect 12069 262 12079 296
rect 12113 262 12134 296
rect 12069 244 12134 262
rect 12164 358 12216 372
rect 12164 324 12174 358
rect 12208 324 12216 358
rect 12164 290 12216 324
rect 12164 256 12174 290
rect 12208 256 12216 290
rect 12164 244 12216 256
rect 12270 339 12322 388
rect 12270 305 12278 339
rect 12312 305 12322 339
rect 12270 271 12322 305
rect 12069 188 12119 244
rect 12270 237 12278 271
rect 12312 237 12322 271
rect 12270 188 12322 237
rect 12352 376 12404 388
rect 12352 342 12362 376
rect 12396 342 12404 376
rect 12556 376 12608 388
rect 12352 320 12404 342
rect 12556 342 12564 376
rect 12598 342 12608 376
rect 12352 192 12419 320
rect 12449 240 12502 320
rect 12449 206 12460 240
rect 12494 206 12502 240
rect 12556 220 12608 342
rect 12638 220 12680 388
rect 12710 350 12786 388
rect 12710 316 12730 350
rect 12764 316 12786 350
rect 12710 304 12786 316
rect 12816 376 12907 388
rect 12816 342 12838 376
rect 12872 342 12907 376
rect 12816 304 12907 342
rect 12937 304 13012 388
rect 13042 375 13096 388
rect 13042 341 13052 375
rect 13086 341 13096 375
rect 13042 304 13096 341
rect 13126 304 13240 388
rect 12710 220 12760 304
rect 12449 192 12502 206
rect 12352 188 12402 192
rect 13188 220 13240 304
rect 13270 376 13377 388
rect 13270 342 13327 376
rect 13361 342 13377 376
rect 13270 308 13377 342
rect 13270 274 13327 308
rect 13361 274 13377 308
rect 13270 220 13377 274
rect 13407 220 13461 388
rect 13491 350 13569 388
rect 13491 316 13501 350
rect 13535 316 13569 350
rect 13491 304 13569 316
rect 13599 366 13675 388
rect 13599 332 13621 366
rect 13655 332 13675 366
rect 13599 304 13675 332
rect 13705 304 13795 388
rect 13825 375 13879 388
rect 13825 341 13835 375
rect 13869 341 13879 375
rect 13825 304 13879 341
rect 13909 368 13971 388
rect 13909 334 13927 368
rect 13961 334 13971 368
rect 13909 304 13971 334
rect 14001 352 14053 388
rect 14001 318 14011 352
rect 14045 318 14053 352
rect 14001 304 14053 318
rect 14107 368 14159 382
rect 14107 334 14115 368
rect 14149 334 14159 368
rect 13491 282 13553 304
rect 13491 248 13501 282
rect 13535 248 13553 282
rect 13491 220 13553 248
rect 14107 300 14159 334
rect 14107 266 14115 300
rect 14149 266 14159 300
rect 14107 254 14159 266
rect 14189 352 14243 382
rect 14189 318 14199 352
rect 14233 318 14243 352
rect 14189 254 14243 318
rect 14273 368 14325 382
rect 14273 334 14283 368
rect 14317 334 14325 368
rect 14273 300 14325 334
rect 14273 266 14283 300
rect 14317 266 14325 300
rect 14273 254 14325 266
rect 14379 340 14431 388
rect 14379 306 14387 340
rect 14421 306 14431 340
rect 14379 272 14431 306
rect 14379 238 14387 272
rect 14421 238 14431 272
rect 14379 188 14431 238
rect 14461 372 14511 388
rect 14461 364 14526 372
rect 14461 330 14471 364
rect 14505 330 14526 364
rect 14461 296 14526 330
rect 14461 262 14471 296
rect 14505 262 14526 296
rect 14461 244 14526 262
rect 14556 358 14608 372
rect 14556 324 14566 358
rect 14600 324 14608 358
rect 14556 290 14608 324
rect 14556 256 14566 290
rect 14600 256 14608 290
rect 14556 244 14608 256
rect 14662 339 14714 388
rect 14662 305 14670 339
rect 14704 305 14714 339
rect 14662 271 14714 305
rect 14461 188 14511 244
rect 14662 237 14670 271
rect 14704 237 14714 271
rect 14662 188 14714 237
rect 14744 376 14796 388
rect 14744 342 14754 376
rect 14788 342 14796 376
rect 14948 376 15000 388
rect 14744 320 14796 342
rect 14948 342 14956 376
rect 14990 342 15000 376
rect 14744 192 14811 320
rect 14841 240 14894 320
rect 14841 206 14852 240
rect 14886 206 14894 240
rect 14948 220 15000 342
rect 15030 220 15072 388
rect 15102 350 15178 388
rect 15102 316 15122 350
rect 15156 316 15178 350
rect 15102 304 15178 316
rect 15208 376 15299 388
rect 15208 342 15230 376
rect 15264 342 15299 376
rect 15208 304 15299 342
rect 15329 304 15404 388
rect 15434 375 15488 388
rect 15434 341 15444 375
rect 15478 341 15488 375
rect 15434 304 15488 341
rect 15518 304 15632 388
rect 15102 220 15152 304
rect 14841 192 14894 206
rect 14744 188 14794 192
rect 15580 220 15632 304
rect 15662 376 15769 388
rect 15662 342 15719 376
rect 15753 342 15769 376
rect 15662 308 15769 342
rect 15662 274 15719 308
rect 15753 274 15769 308
rect 15662 220 15769 274
rect 15799 220 15853 388
rect 15883 350 15961 388
rect 15883 316 15893 350
rect 15927 316 15961 350
rect 15883 304 15961 316
rect 15991 366 16067 388
rect 15991 332 16013 366
rect 16047 332 16067 366
rect 15991 304 16067 332
rect 16097 304 16187 388
rect 16217 375 16271 388
rect 16217 341 16227 375
rect 16261 341 16271 375
rect 16217 304 16271 341
rect 16301 368 16363 388
rect 16301 334 16319 368
rect 16353 334 16363 368
rect 16301 304 16363 334
rect 16393 352 16445 388
rect 16393 318 16403 352
rect 16437 318 16445 352
rect 16393 304 16445 318
rect 16499 368 16551 382
rect 16499 334 16507 368
rect 16541 334 16551 368
rect 15883 282 15945 304
rect 15883 248 15893 282
rect 15927 248 15945 282
rect 15883 220 15945 248
rect 16499 300 16551 334
rect 16499 266 16507 300
rect 16541 266 16551 300
rect 16499 254 16551 266
rect 16581 352 16635 382
rect 16581 318 16591 352
rect 16625 318 16635 352
rect 16581 254 16635 318
rect 16665 368 16717 382
rect 16665 334 16675 368
rect 16709 334 16717 368
rect 16665 300 16717 334
rect 16665 266 16675 300
rect 16709 266 16717 300
rect 16665 254 16717 266
<< ndiffc >>
rect 37 2482 71 2516
rect 123 2469 157 2503
rect 209 2499 243 2533
rect 313 2505 347 2539
rect 397 2473 431 2507
rect 481 2505 515 2539
rect 565 2473 599 2507
rect 649 2505 683 2539
rect 733 2537 767 2571
rect 733 2469 767 2503
rect 865 2541 899 2575
rect 865 2473 899 2507
rect 949 2541 983 2575
rect 949 2473 983 2507
rect 1033 2473 1067 2507
rect 1117 2541 1151 2575
rect 1117 2473 1151 2507
rect 1201 2473 1235 2507
rect 1285 2541 1319 2575
rect 1285 2473 1319 2507
rect 1369 2473 1403 2507
rect 1453 2541 1487 2575
rect 1453 2473 1487 2507
rect 1537 2473 1571 2507
rect 1621 2541 1655 2575
rect 1621 2473 1655 2507
rect 1705 2473 1739 2507
rect 1789 2541 1823 2575
rect 1789 2473 1823 2507
rect 1873 2473 1907 2507
rect 1957 2541 1991 2575
rect 1957 2473 1991 2507
rect 2041 2473 2075 2507
rect 2125 2541 2159 2575
rect 2125 2473 2159 2507
rect 2209 2473 2243 2507
rect 2293 2541 2327 2575
rect 2293 2473 2327 2507
rect 2377 2473 2411 2507
rect 2461 2541 2495 2575
rect 2461 2473 2495 2507
rect 2545 2473 2579 2507
rect 2629 2541 2663 2575
rect 2629 2473 2663 2507
rect 2713 2473 2747 2507
rect 4421 2482 4455 2516
rect 4507 2469 4541 2503
rect 4593 2499 4627 2533
rect 4697 2505 4731 2539
rect 4781 2473 4815 2507
rect 4865 2505 4899 2539
rect 4949 2473 4983 2507
rect 5033 2505 5067 2539
rect 5117 2537 5151 2571
rect 5117 2469 5151 2503
rect 5249 2541 5283 2575
rect 5249 2473 5283 2507
rect 5333 2541 5367 2575
rect 5333 2473 5367 2507
rect 5417 2473 5451 2507
rect 5501 2541 5535 2575
rect 5501 2473 5535 2507
rect 5585 2473 5619 2507
rect 5669 2541 5703 2575
rect 5669 2473 5703 2507
rect 5753 2473 5787 2507
rect 5837 2541 5871 2575
rect 5837 2473 5871 2507
rect 5921 2473 5955 2507
rect 6005 2541 6039 2575
rect 6005 2473 6039 2507
rect 6089 2473 6123 2507
rect 6173 2541 6207 2575
rect 6173 2473 6207 2507
rect 6257 2473 6291 2507
rect 6341 2541 6375 2575
rect 6341 2473 6375 2507
rect 6425 2473 6459 2507
rect 6509 2541 6543 2575
rect 6509 2473 6543 2507
rect 6593 2473 6627 2507
rect 6677 2541 6711 2575
rect 6677 2473 6711 2507
rect 6761 2473 6795 2507
rect 6845 2541 6879 2575
rect 6845 2473 6879 2507
rect 6929 2473 6963 2507
rect 7013 2541 7047 2575
rect 7013 2473 7047 2507
rect 7097 2473 7131 2507
rect 35 1346 69 1380
rect 119 1327 153 1361
rect 326 1342 360 1376
rect 561 1342 595 1376
rect 629 1342 663 1376
rect 713 1342 747 1376
rect 1515 1342 1549 1376
rect 1599 1342 1633 1376
rect 1667 1342 1701 1376
rect 1902 1342 1936 1376
rect 2109 1327 2143 1361
rect 2193 1346 2227 1380
rect 2427 1346 2461 1380
rect 2511 1327 2545 1361
rect 2718 1342 2752 1376
rect 2953 1342 2987 1376
rect 3021 1342 3055 1376
rect 3105 1342 3139 1376
rect 3907 1342 3941 1376
rect 3991 1342 4025 1376
rect 4059 1342 4093 1376
rect 4294 1342 4328 1376
rect 4501 1327 4535 1361
rect 4585 1346 4619 1380
rect 4819 1346 4853 1380
rect 4903 1327 4937 1361
rect 5110 1342 5144 1376
rect 5345 1342 5379 1376
rect 5413 1342 5447 1376
rect 5497 1342 5531 1376
rect 6297 1342 6331 1376
rect 6381 1342 6415 1376
rect 6449 1342 6483 1376
rect 6684 1342 6718 1376
rect 6891 1327 6925 1361
rect 6975 1346 7009 1380
rect 7211 1346 7245 1380
rect 7295 1327 7329 1361
rect 7502 1342 7536 1376
rect 7737 1342 7771 1376
rect 7805 1342 7839 1376
rect 7889 1342 7923 1376
rect 8691 1342 8725 1376
rect 8775 1342 8809 1376
rect 8843 1342 8877 1376
rect 9078 1342 9112 1376
rect 9285 1327 9319 1361
rect 9369 1346 9403 1380
rect 9603 1346 9637 1380
rect 9687 1327 9721 1361
rect 9894 1342 9928 1376
rect 10129 1342 10163 1376
rect 10197 1342 10231 1376
rect 10281 1342 10315 1376
rect 11083 1342 11117 1376
rect 11167 1342 11201 1376
rect 11235 1342 11269 1376
rect 11470 1342 11504 1376
rect 11677 1327 11711 1361
rect 11761 1346 11795 1380
rect 11995 1346 12029 1380
rect 12079 1327 12113 1361
rect 12286 1342 12320 1376
rect 12521 1342 12555 1376
rect 12589 1342 12623 1376
rect 12673 1342 12707 1376
rect 13473 1342 13507 1376
rect 13557 1342 13591 1376
rect 13625 1342 13659 1376
rect 13860 1342 13894 1376
rect 14067 1327 14101 1361
rect 14151 1346 14185 1380
rect 14387 1346 14421 1380
rect 14471 1327 14505 1361
rect 14678 1342 14712 1376
rect 14913 1342 14947 1376
rect 14981 1342 15015 1376
rect 15065 1342 15099 1376
rect 15867 1342 15901 1376
rect 15951 1342 15985 1376
rect 16019 1342 16053 1376
rect 16254 1342 16288 1376
rect 16461 1327 16495 1361
rect 16545 1346 16579 1380
rect 35 665 69 699
rect 119 639 153 673
rect 203 665 237 699
rect 307 639 341 673
rect 391 657 425 691
rect 496 639 530 673
rect 717 635 751 669
rect 801 641 835 675
rect 897 699 931 733
rect 981 673 1015 707
rect 1085 639 1119 673
rect 1289 639 1323 673
rect 1481 635 1515 669
rect 1565 655 1599 689
rect 1673 713 1707 747
rect 1757 647 1791 681
rect 1861 649 1895 683
rect 1956 639 1990 673
rect 2040 673 2074 707
rect 2144 665 2178 699
rect 2239 639 2273 673
rect 2323 675 2357 709
rect 2427 665 2461 699
rect 2511 639 2545 673
rect 2595 665 2629 699
rect 2699 639 2733 673
rect 2783 657 2817 691
rect 2888 639 2922 673
rect 3109 635 3143 669
rect 3193 641 3227 675
rect 3289 699 3323 733
rect 3373 673 3407 707
rect 3477 639 3511 673
rect 3681 639 3715 673
rect 3873 635 3907 669
rect 3957 655 3991 689
rect 4065 713 4099 747
rect 4149 647 4183 681
rect 4253 649 4287 683
rect 4348 639 4382 673
rect 4432 673 4466 707
rect 4536 665 4570 699
rect 4631 639 4665 673
rect 4715 675 4749 709
rect 4819 665 4853 699
rect 4903 639 4937 673
rect 4987 665 5021 699
rect 5091 639 5125 673
rect 5175 657 5209 691
rect 5280 639 5314 673
rect 5501 635 5535 669
rect 5585 641 5619 675
rect 5681 699 5715 733
rect 5765 673 5799 707
rect 5869 639 5903 673
rect 6073 639 6107 673
rect 6265 635 6299 669
rect 6349 655 6383 689
rect 6457 713 6491 747
rect 6541 647 6575 681
rect 6645 649 6679 683
rect 6740 639 6774 673
rect 6824 673 6858 707
rect 6928 665 6962 699
rect 7023 639 7057 673
rect 7107 675 7141 709
rect 7211 665 7245 699
rect 7295 639 7329 673
rect 7379 665 7413 699
rect 7483 639 7517 673
rect 7567 657 7601 691
rect 7672 639 7706 673
rect 7893 635 7927 669
rect 7977 641 8011 675
rect 8073 699 8107 733
rect 8157 673 8191 707
rect 8261 639 8295 673
rect 8465 639 8499 673
rect 8657 635 8691 669
rect 8741 655 8775 689
rect 8849 713 8883 747
rect 8933 647 8967 681
rect 9037 649 9071 683
rect 9132 639 9166 673
rect 9216 673 9250 707
rect 9320 665 9354 699
rect 9415 639 9449 673
rect 9499 675 9533 709
rect 9603 665 9637 699
rect 9687 639 9721 673
rect 9771 665 9805 699
rect 9875 639 9909 673
rect 9959 657 9993 691
rect 10064 639 10098 673
rect 10285 635 10319 669
rect 10369 641 10403 675
rect 10465 699 10499 733
rect 10549 673 10583 707
rect 10653 639 10687 673
rect 10857 639 10891 673
rect 11049 635 11083 669
rect 11133 655 11167 689
rect 11241 713 11275 747
rect 11325 647 11359 681
rect 11429 649 11463 683
rect 11524 639 11558 673
rect 11608 673 11642 707
rect 11712 665 11746 699
rect 11807 639 11841 673
rect 11891 675 11925 709
rect 11995 665 12029 699
rect 12079 639 12113 673
rect 12163 665 12197 699
rect 12267 639 12301 673
rect 12351 657 12385 691
rect 12456 639 12490 673
rect 12677 635 12711 669
rect 12761 641 12795 675
rect 12857 699 12891 733
rect 12941 673 12975 707
rect 13045 639 13079 673
rect 13249 639 13283 673
rect 13441 635 13475 669
rect 13525 655 13559 689
rect 13633 713 13667 747
rect 13717 647 13751 681
rect 13821 649 13855 683
rect 13916 639 13950 673
rect 14000 673 14034 707
rect 14104 665 14138 699
rect 14199 639 14233 673
rect 14283 675 14317 709
rect 14387 665 14421 699
rect 14471 639 14505 673
rect 14555 665 14589 699
rect 14659 639 14693 673
rect 14743 657 14777 691
rect 14848 639 14882 673
rect 15069 635 15103 669
rect 15153 641 15187 675
rect 15249 699 15283 733
rect 15333 673 15367 707
rect 15437 639 15471 673
rect 15641 639 15675 673
rect 15833 635 15867 669
rect 15917 655 15951 689
rect 16025 713 16059 747
rect 16109 647 16143 681
rect 16213 649 16247 683
rect 16308 639 16342 673
rect 16392 673 16426 707
rect 16496 665 16530 699
rect 16591 639 16625 673
rect 16675 675 16709 709
rect 35 -14 69 20
rect 119 -50 153 -16
rect 214 -24 248 10
rect 318 -16 352 18
rect 402 -50 436 -16
rect 497 -40 531 -6
rect 601 -42 635 -8
rect 685 24 719 58
rect 793 -34 827 0
rect 877 -54 911 -20
rect 1069 -50 1103 -16
rect 1273 -50 1307 -16
rect 1377 -16 1411 18
rect 1461 10 1495 44
rect 1557 -48 1591 -14
rect 1641 -54 1675 -20
rect 1862 -50 1896 -16
rect 1967 -32 2001 2
rect 2051 -50 2085 -16
rect 2155 -24 2189 10
rect 2239 -50 2273 -16
rect 2323 -24 2357 10
rect 2427 -14 2461 20
rect 2511 -50 2545 -16
rect 2606 -24 2640 10
rect 2710 -16 2744 18
rect 2794 -50 2828 -16
rect 2889 -40 2923 -6
rect 2993 -42 3027 -8
rect 3077 24 3111 58
rect 3185 -34 3219 0
rect 3269 -54 3303 -20
rect 3461 -50 3495 -16
rect 3665 -50 3699 -16
rect 3769 -16 3803 18
rect 3853 10 3887 44
rect 3949 -48 3983 -14
rect 4033 -54 4067 -20
rect 4254 -50 4288 -16
rect 4359 -32 4393 2
rect 4443 -50 4477 -16
rect 4547 -24 4581 10
rect 4631 -50 4665 -16
rect 4715 -24 4749 10
rect 4819 -14 4853 20
rect 4903 -50 4937 -16
rect 4998 -24 5032 10
rect 5102 -16 5136 18
rect 5186 -50 5220 -16
rect 5281 -40 5315 -6
rect 5385 -42 5419 -8
rect 5469 24 5503 58
rect 5577 -34 5611 0
rect 5661 -54 5695 -20
rect 5853 -50 5887 -16
rect 6057 -50 6091 -16
rect 6161 -16 6195 18
rect 6245 10 6279 44
rect 6341 -48 6375 -14
rect 6425 -54 6459 -20
rect 6646 -50 6680 -16
rect 6751 -32 6785 2
rect 6835 -50 6869 -16
rect 6939 -24 6973 10
rect 7023 -50 7057 -16
rect 7107 -24 7141 10
rect 7211 -14 7245 20
rect 7295 -50 7329 -16
rect 7390 -24 7424 10
rect 7494 -16 7528 18
rect 7578 -50 7612 -16
rect 7673 -40 7707 -6
rect 7777 -42 7811 -8
rect 7861 24 7895 58
rect 7969 -34 8003 0
rect 8053 -54 8087 -20
rect 8245 -50 8279 -16
rect 8449 -50 8483 -16
rect 8553 -16 8587 18
rect 8637 10 8671 44
rect 8733 -48 8767 -14
rect 8817 -54 8851 -20
rect 9038 -50 9072 -16
rect 9143 -32 9177 2
rect 9227 -50 9261 -16
rect 9331 -24 9365 10
rect 9415 -50 9449 -16
rect 9499 -24 9533 10
rect 9603 -14 9637 20
rect 9687 -50 9721 -16
rect 9782 -24 9816 10
rect 9886 -16 9920 18
rect 9970 -50 10004 -16
rect 10065 -40 10099 -6
rect 10169 -42 10203 -8
rect 10253 24 10287 58
rect 10361 -34 10395 0
rect 10445 -54 10479 -20
rect 10637 -50 10671 -16
rect 10841 -50 10875 -16
rect 10945 -16 10979 18
rect 11029 10 11063 44
rect 11125 -48 11159 -14
rect 11209 -54 11243 -20
rect 11430 -50 11464 -16
rect 11535 -32 11569 2
rect 11619 -50 11653 -16
rect 11723 -24 11757 10
rect 11807 -50 11841 -16
rect 11891 -24 11925 10
rect 11995 -14 12029 20
rect 12079 -50 12113 -16
rect 12174 -24 12208 10
rect 12278 -16 12312 18
rect 12362 -50 12396 -16
rect 12457 -40 12491 -6
rect 12561 -42 12595 -8
rect 12645 24 12679 58
rect 12753 -34 12787 0
rect 12837 -54 12871 -20
rect 13029 -50 13063 -16
rect 13233 -50 13267 -16
rect 13337 -16 13371 18
rect 13421 10 13455 44
rect 13517 -48 13551 -14
rect 13601 -54 13635 -20
rect 13822 -50 13856 -16
rect 13927 -32 13961 2
rect 14011 -50 14045 -16
rect 14115 -24 14149 10
rect 14199 -50 14233 -16
rect 14283 -24 14317 10
rect 14387 -14 14421 20
rect 14471 -50 14505 -16
rect 14566 -24 14600 10
rect 14670 -16 14704 18
rect 14754 -50 14788 -16
rect 14849 -40 14883 -6
rect 14953 -42 14987 -8
rect 15037 24 15071 58
rect 15145 -34 15179 0
rect 15229 -54 15263 -20
rect 15421 -50 15455 -16
rect 15625 -50 15659 -16
rect 15729 -16 15763 18
rect 15813 10 15847 44
rect 15909 -48 15943 -14
rect 15993 -54 16027 -20
rect 16214 -50 16248 -16
rect 16319 -32 16353 2
rect 16403 -50 16437 -16
rect 16507 -24 16541 10
rect 16591 -50 16625 -16
rect 16675 -24 16709 10
<< pdiffc >>
rect 37 2853 71 2887
rect 37 2785 71 2819
rect 123 2853 157 2887
rect 123 2785 157 2819
rect 209 2853 243 2887
rect 209 2772 243 2806
rect 313 2855 347 2889
rect 313 2787 347 2821
rect 313 2719 347 2753
rect 397 2861 431 2895
rect 397 2793 431 2827
rect 481 2839 515 2873
rect 481 2744 515 2778
rect 565 2861 599 2895
rect 565 2793 599 2827
rect 649 2839 683 2873
rect 649 2744 683 2778
rect 733 2861 767 2895
rect 733 2793 767 2827
rect 733 2725 767 2759
rect 865 2861 899 2895
rect 865 2793 899 2827
rect 865 2725 899 2759
rect 949 2855 983 2889
rect 949 2787 983 2821
rect 949 2719 983 2753
rect 1033 2861 1067 2895
rect 1033 2793 1067 2827
rect 1117 2855 1151 2889
rect 1117 2787 1151 2821
rect 1117 2719 1151 2753
rect 1201 2861 1235 2895
rect 1201 2793 1235 2827
rect 1285 2855 1319 2889
rect 1285 2787 1319 2821
rect 1285 2719 1319 2753
rect 1369 2861 1403 2895
rect 1369 2793 1403 2827
rect 1453 2855 1487 2889
rect 1453 2787 1487 2821
rect 1453 2719 1487 2753
rect 1537 2861 1571 2895
rect 1537 2793 1571 2827
rect 1621 2855 1655 2889
rect 1621 2787 1655 2821
rect 1621 2719 1655 2753
rect 1705 2861 1739 2895
rect 1705 2793 1739 2827
rect 1789 2855 1823 2889
rect 1789 2787 1823 2821
rect 1789 2719 1823 2753
rect 1873 2861 1907 2895
rect 1873 2793 1907 2827
rect 1957 2855 1991 2889
rect 1957 2787 1991 2821
rect 1957 2719 1991 2753
rect 2041 2861 2075 2895
rect 2041 2793 2075 2827
rect 2125 2855 2159 2889
rect 2125 2787 2159 2821
rect 2125 2719 2159 2753
rect 2209 2861 2243 2895
rect 2209 2793 2243 2827
rect 2293 2855 2327 2889
rect 2293 2787 2327 2821
rect 2293 2719 2327 2753
rect 2377 2861 2411 2895
rect 2377 2793 2411 2827
rect 2461 2855 2495 2889
rect 2461 2787 2495 2821
rect 2461 2719 2495 2753
rect 2545 2861 2579 2895
rect 2545 2793 2579 2827
rect 2629 2855 2663 2889
rect 2629 2787 2663 2821
rect 2629 2719 2663 2753
rect 2713 2861 2747 2895
rect 2713 2793 2747 2827
rect 4421 2853 4455 2887
rect 4421 2785 4455 2819
rect 4507 2853 4541 2887
rect 4507 2785 4541 2819
rect 4593 2853 4627 2887
rect 4593 2772 4627 2806
rect 4697 2855 4731 2889
rect 4697 2787 4731 2821
rect 4697 2719 4731 2753
rect 4781 2861 4815 2895
rect 4781 2793 4815 2827
rect 4865 2839 4899 2873
rect 4865 2744 4899 2778
rect 4949 2861 4983 2895
rect 4949 2793 4983 2827
rect 5033 2839 5067 2873
rect 5033 2744 5067 2778
rect 5117 2861 5151 2895
rect 5117 2793 5151 2827
rect 5117 2725 5151 2759
rect 5249 2861 5283 2895
rect 5249 2793 5283 2827
rect 5249 2725 5283 2759
rect 5333 2855 5367 2889
rect 5333 2787 5367 2821
rect 5333 2719 5367 2753
rect 5417 2861 5451 2895
rect 5417 2793 5451 2827
rect 5501 2855 5535 2889
rect 5501 2787 5535 2821
rect 5501 2719 5535 2753
rect 5585 2861 5619 2895
rect 5585 2793 5619 2827
rect 5669 2855 5703 2889
rect 5669 2787 5703 2821
rect 5669 2719 5703 2753
rect 5753 2861 5787 2895
rect 5753 2793 5787 2827
rect 5837 2855 5871 2889
rect 5837 2787 5871 2821
rect 5837 2719 5871 2753
rect 5921 2861 5955 2895
rect 5921 2793 5955 2827
rect 6005 2855 6039 2889
rect 6005 2787 6039 2821
rect 6005 2719 6039 2753
rect 6089 2861 6123 2895
rect 6089 2793 6123 2827
rect 6173 2855 6207 2889
rect 6173 2787 6207 2821
rect 6173 2719 6207 2753
rect 6257 2861 6291 2895
rect 6257 2793 6291 2827
rect 6341 2855 6375 2889
rect 6341 2787 6375 2821
rect 6341 2719 6375 2753
rect 6425 2861 6459 2895
rect 6425 2793 6459 2827
rect 6509 2855 6543 2889
rect 6509 2787 6543 2821
rect 6509 2719 6543 2753
rect 6593 2861 6627 2895
rect 6593 2793 6627 2827
rect 6677 2855 6711 2889
rect 6677 2787 6711 2821
rect 6677 2719 6711 2753
rect 6761 2861 6795 2895
rect 6761 2793 6795 2827
rect 6845 2855 6879 2889
rect 6845 2787 6879 2821
rect 6845 2719 6879 2753
rect 6929 2861 6963 2895
rect 6929 2793 6963 2827
rect 7013 2855 7047 2889
rect 7013 2787 7047 2821
rect 7013 2719 7047 2753
rect 7097 2861 7131 2895
rect 7097 2793 7131 2827
rect 35 1719 69 1753
rect 35 1651 69 1685
rect 35 1583 69 1617
rect 119 1719 153 1753
rect 119 1651 153 1685
rect 355 1659 389 1693
rect 430 1659 464 1693
rect 627 1659 661 1693
rect 713 1659 747 1693
rect 1515 1659 1549 1693
rect 1601 1659 1635 1693
rect 1798 1659 1832 1693
rect 1873 1659 1907 1693
rect 2109 1719 2143 1753
rect 2109 1651 2143 1685
rect 119 1583 153 1617
rect 2109 1583 2143 1617
rect 2193 1719 2227 1753
rect 2193 1651 2227 1685
rect 2193 1583 2227 1617
rect 2427 1719 2461 1753
rect 2427 1651 2461 1685
rect 2427 1583 2461 1617
rect 2511 1719 2545 1753
rect 2511 1651 2545 1685
rect 2747 1659 2781 1693
rect 2822 1659 2856 1693
rect 3019 1659 3053 1693
rect 3105 1659 3139 1693
rect 3907 1659 3941 1693
rect 3993 1659 4027 1693
rect 4190 1659 4224 1693
rect 4265 1659 4299 1693
rect 4501 1719 4535 1753
rect 4501 1651 4535 1685
rect 2511 1583 2545 1617
rect 4501 1583 4535 1617
rect 4585 1719 4619 1753
rect 4585 1651 4619 1685
rect 4585 1583 4619 1617
rect 4819 1719 4853 1753
rect 4819 1651 4853 1685
rect 4819 1583 4853 1617
rect 4903 1719 4937 1753
rect 4903 1651 4937 1685
rect 5139 1659 5173 1693
rect 5214 1659 5248 1693
rect 5411 1659 5445 1693
rect 5497 1659 5531 1693
rect 6297 1659 6331 1693
rect 6383 1659 6417 1693
rect 6580 1659 6614 1693
rect 6655 1659 6689 1693
rect 6891 1719 6925 1753
rect 6891 1651 6925 1685
rect 4903 1583 4937 1617
rect 6891 1583 6925 1617
rect 6975 1719 7009 1753
rect 6975 1651 7009 1685
rect 6975 1583 7009 1617
rect 7211 1719 7245 1753
rect 7211 1651 7245 1685
rect 7211 1583 7245 1617
rect 7295 1719 7329 1753
rect 7295 1651 7329 1685
rect 7531 1659 7565 1693
rect 7606 1659 7640 1693
rect 7803 1659 7837 1693
rect 7889 1659 7923 1693
rect 8691 1659 8725 1693
rect 8777 1659 8811 1693
rect 8974 1659 9008 1693
rect 9049 1659 9083 1693
rect 9285 1719 9319 1753
rect 9285 1651 9319 1685
rect 7295 1583 7329 1617
rect 9285 1583 9319 1617
rect 9369 1719 9403 1753
rect 9369 1651 9403 1685
rect 9369 1583 9403 1617
rect 9603 1719 9637 1753
rect 9603 1651 9637 1685
rect 9603 1583 9637 1617
rect 9687 1719 9721 1753
rect 9687 1651 9721 1685
rect 9923 1659 9957 1693
rect 9998 1659 10032 1693
rect 10195 1659 10229 1693
rect 10281 1659 10315 1693
rect 11083 1659 11117 1693
rect 11169 1659 11203 1693
rect 11366 1659 11400 1693
rect 11441 1659 11475 1693
rect 11677 1719 11711 1753
rect 11677 1651 11711 1685
rect 9687 1583 9721 1617
rect 11677 1583 11711 1617
rect 11761 1719 11795 1753
rect 11761 1651 11795 1685
rect 11761 1583 11795 1617
rect 11995 1719 12029 1753
rect 11995 1651 12029 1685
rect 11995 1583 12029 1617
rect 12079 1719 12113 1753
rect 12079 1651 12113 1685
rect 12315 1659 12349 1693
rect 12390 1659 12424 1693
rect 12587 1659 12621 1693
rect 12673 1659 12707 1693
rect 13473 1659 13507 1693
rect 13559 1659 13593 1693
rect 13756 1659 13790 1693
rect 13831 1659 13865 1693
rect 14067 1719 14101 1753
rect 14067 1651 14101 1685
rect 12079 1583 12113 1617
rect 14067 1583 14101 1617
rect 14151 1719 14185 1753
rect 14151 1651 14185 1685
rect 14151 1583 14185 1617
rect 14387 1719 14421 1753
rect 14387 1651 14421 1685
rect 14387 1583 14421 1617
rect 14471 1719 14505 1753
rect 14471 1651 14505 1685
rect 14707 1659 14741 1693
rect 14782 1659 14816 1693
rect 14979 1659 15013 1693
rect 15065 1659 15099 1693
rect 15867 1659 15901 1693
rect 15953 1659 15987 1693
rect 16150 1659 16184 1693
rect 16225 1659 16259 1693
rect 16461 1719 16495 1753
rect 16461 1651 16495 1685
rect 14471 1583 14505 1617
rect 16461 1583 16495 1617
rect 16545 1719 16579 1753
rect 16545 1651 16579 1685
rect 16545 1583 16579 1617
rect 35 1023 69 1057
rect 35 955 69 989
rect 119 1007 153 1041
rect 203 1023 237 1057
rect 307 1007 341 1041
rect 391 1023 425 1057
rect 483 1030 517 1064
rect 697 1021 731 1055
rect 817 1005 851 1039
rect 203 955 237 989
rect 817 937 851 971
rect 991 1031 1025 1065
rect 991 963 1025 997
rect 1266 1030 1300 1064
rect 1480 1031 1514 1065
rect 1588 1005 1622 1039
rect 1754 1031 1788 1065
rect 1956 1031 1990 1065
rect 1858 895 1892 929
rect 2040 994 2074 1028
rect 2040 926 2074 960
rect 2144 1013 2178 1047
rect 2144 945 2178 979
rect 2239 1019 2273 1053
rect 2239 951 2273 985
rect 2323 995 2357 1029
rect 2323 927 2357 961
rect 2427 1023 2461 1057
rect 2427 955 2461 989
rect 2511 1007 2545 1041
rect 2595 1023 2629 1057
rect 2699 1007 2733 1041
rect 2783 1023 2817 1057
rect 2875 1030 2909 1064
rect 3089 1021 3123 1055
rect 3209 1005 3243 1039
rect 2595 955 2629 989
rect 3209 937 3243 971
rect 3383 1031 3417 1065
rect 3383 963 3417 997
rect 3658 1030 3692 1064
rect 3872 1031 3906 1065
rect 3980 1005 4014 1039
rect 4146 1031 4180 1065
rect 4348 1031 4382 1065
rect 4250 895 4284 929
rect 4432 994 4466 1028
rect 4432 926 4466 960
rect 4536 1013 4570 1047
rect 4536 945 4570 979
rect 4631 1019 4665 1053
rect 4631 951 4665 985
rect 4715 995 4749 1029
rect 4715 927 4749 961
rect 4819 1023 4853 1057
rect 4819 955 4853 989
rect 4903 1007 4937 1041
rect 4987 1023 5021 1057
rect 5091 1007 5125 1041
rect 5175 1023 5209 1057
rect 5267 1030 5301 1064
rect 5481 1021 5515 1055
rect 5601 1005 5635 1039
rect 4987 955 5021 989
rect 5601 937 5635 971
rect 5775 1031 5809 1065
rect 5775 963 5809 997
rect 6050 1030 6084 1064
rect 6264 1031 6298 1065
rect 6372 1005 6406 1039
rect 6538 1031 6572 1065
rect 6740 1031 6774 1065
rect 6642 895 6676 929
rect 6824 994 6858 1028
rect 6824 926 6858 960
rect 6928 1013 6962 1047
rect 6928 945 6962 979
rect 7023 1019 7057 1053
rect 7023 951 7057 985
rect 7107 995 7141 1029
rect 7107 927 7141 961
rect 7211 1023 7245 1057
rect 7211 955 7245 989
rect 7295 1007 7329 1041
rect 7379 1023 7413 1057
rect 7483 1007 7517 1041
rect 7567 1023 7601 1057
rect 7659 1030 7693 1064
rect 7873 1021 7907 1055
rect 7993 1005 8027 1039
rect 7379 955 7413 989
rect 7993 937 8027 971
rect 8167 1031 8201 1065
rect 8167 963 8201 997
rect 8442 1030 8476 1064
rect 8656 1031 8690 1065
rect 8764 1005 8798 1039
rect 8930 1031 8964 1065
rect 9132 1031 9166 1065
rect 9034 895 9068 929
rect 9216 994 9250 1028
rect 9216 926 9250 960
rect 9320 1013 9354 1047
rect 9320 945 9354 979
rect 9415 1019 9449 1053
rect 9415 951 9449 985
rect 9499 995 9533 1029
rect 9499 927 9533 961
rect 9603 1023 9637 1057
rect 9603 955 9637 989
rect 9687 1007 9721 1041
rect 9771 1023 9805 1057
rect 9875 1007 9909 1041
rect 9959 1023 9993 1057
rect 10051 1030 10085 1064
rect 10265 1021 10299 1055
rect 10385 1005 10419 1039
rect 9771 955 9805 989
rect 10385 937 10419 971
rect 10559 1031 10593 1065
rect 10559 963 10593 997
rect 10834 1030 10868 1064
rect 11048 1031 11082 1065
rect 11156 1005 11190 1039
rect 11322 1031 11356 1065
rect 11524 1031 11558 1065
rect 11426 895 11460 929
rect 11608 994 11642 1028
rect 11608 926 11642 960
rect 11712 1013 11746 1047
rect 11712 945 11746 979
rect 11807 1019 11841 1053
rect 11807 951 11841 985
rect 11891 995 11925 1029
rect 11891 927 11925 961
rect 11995 1023 12029 1057
rect 11995 955 12029 989
rect 12079 1007 12113 1041
rect 12163 1023 12197 1057
rect 12267 1007 12301 1041
rect 12351 1023 12385 1057
rect 12443 1030 12477 1064
rect 12657 1021 12691 1055
rect 12777 1005 12811 1039
rect 12163 955 12197 989
rect 12777 937 12811 971
rect 12951 1031 12985 1065
rect 12951 963 12985 997
rect 13226 1030 13260 1064
rect 13440 1031 13474 1065
rect 13548 1005 13582 1039
rect 13714 1031 13748 1065
rect 13916 1031 13950 1065
rect 13818 895 13852 929
rect 14000 994 14034 1028
rect 14000 926 14034 960
rect 14104 1013 14138 1047
rect 14104 945 14138 979
rect 14199 1019 14233 1053
rect 14199 951 14233 985
rect 14283 995 14317 1029
rect 14283 927 14317 961
rect 14387 1023 14421 1057
rect 14387 955 14421 989
rect 14471 1007 14505 1041
rect 14555 1023 14589 1057
rect 14659 1007 14693 1041
rect 14743 1023 14777 1057
rect 14835 1030 14869 1064
rect 15049 1021 15083 1055
rect 15169 1005 15203 1039
rect 14555 955 14589 989
rect 15169 937 15203 971
rect 15343 1031 15377 1065
rect 15343 963 15377 997
rect 15618 1030 15652 1064
rect 15832 1031 15866 1065
rect 15940 1005 15974 1039
rect 16106 1031 16140 1065
rect 16308 1031 16342 1065
rect 16210 895 16244 929
rect 16392 994 16426 1028
rect 16392 926 16426 960
rect 16496 1013 16530 1047
rect 16496 945 16530 979
rect 16591 1019 16625 1053
rect 16591 951 16625 985
rect 16675 995 16709 1029
rect 16675 927 16709 961
rect 35 306 69 340
rect 35 238 69 272
rect 119 330 153 364
rect 119 262 153 296
rect 214 324 248 358
rect 214 256 248 290
rect 318 305 352 339
rect 318 237 352 271
rect 402 342 436 376
rect 604 342 638 376
rect 500 206 534 240
rect 770 316 804 350
rect 878 342 912 376
rect 1092 341 1126 375
rect 1367 342 1401 376
rect 1367 274 1401 308
rect 1541 316 1575 350
rect 1661 332 1695 366
rect 1875 341 1909 375
rect 1967 334 2001 368
rect 2051 318 2085 352
rect 2155 334 2189 368
rect 1541 248 1575 282
rect 2155 266 2189 300
rect 2239 318 2273 352
rect 2323 334 2357 368
rect 2323 266 2357 300
rect 2427 306 2461 340
rect 2427 238 2461 272
rect 2511 330 2545 364
rect 2511 262 2545 296
rect 2606 324 2640 358
rect 2606 256 2640 290
rect 2710 305 2744 339
rect 2710 237 2744 271
rect 2794 342 2828 376
rect 2996 342 3030 376
rect 2892 206 2926 240
rect 3162 316 3196 350
rect 3270 342 3304 376
rect 3484 341 3518 375
rect 3759 342 3793 376
rect 3759 274 3793 308
rect 3933 316 3967 350
rect 4053 332 4087 366
rect 4267 341 4301 375
rect 4359 334 4393 368
rect 4443 318 4477 352
rect 4547 334 4581 368
rect 3933 248 3967 282
rect 4547 266 4581 300
rect 4631 318 4665 352
rect 4715 334 4749 368
rect 4715 266 4749 300
rect 4819 306 4853 340
rect 4819 238 4853 272
rect 4903 330 4937 364
rect 4903 262 4937 296
rect 4998 324 5032 358
rect 4998 256 5032 290
rect 5102 305 5136 339
rect 5102 237 5136 271
rect 5186 342 5220 376
rect 5388 342 5422 376
rect 5284 206 5318 240
rect 5554 316 5588 350
rect 5662 342 5696 376
rect 5876 341 5910 375
rect 6151 342 6185 376
rect 6151 274 6185 308
rect 6325 316 6359 350
rect 6445 332 6479 366
rect 6659 341 6693 375
rect 6751 334 6785 368
rect 6835 318 6869 352
rect 6939 334 6973 368
rect 6325 248 6359 282
rect 6939 266 6973 300
rect 7023 318 7057 352
rect 7107 334 7141 368
rect 7107 266 7141 300
rect 7211 306 7245 340
rect 7211 238 7245 272
rect 7295 330 7329 364
rect 7295 262 7329 296
rect 7390 324 7424 358
rect 7390 256 7424 290
rect 7494 305 7528 339
rect 7494 237 7528 271
rect 7578 342 7612 376
rect 7780 342 7814 376
rect 7676 206 7710 240
rect 7946 316 7980 350
rect 8054 342 8088 376
rect 8268 341 8302 375
rect 8543 342 8577 376
rect 8543 274 8577 308
rect 8717 316 8751 350
rect 8837 332 8871 366
rect 9051 341 9085 375
rect 9143 334 9177 368
rect 9227 318 9261 352
rect 9331 334 9365 368
rect 8717 248 8751 282
rect 9331 266 9365 300
rect 9415 318 9449 352
rect 9499 334 9533 368
rect 9499 266 9533 300
rect 9603 306 9637 340
rect 9603 238 9637 272
rect 9687 330 9721 364
rect 9687 262 9721 296
rect 9782 324 9816 358
rect 9782 256 9816 290
rect 9886 305 9920 339
rect 9886 237 9920 271
rect 9970 342 10004 376
rect 10172 342 10206 376
rect 10068 206 10102 240
rect 10338 316 10372 350
rect 10446 342 10480 376
rect 10660 341 10694 375
rect 10935 342 10969 376
rect 10935 274 10969 308
rect 11109 316 11143 350
rect 11229 332 11263 366
rect 11443 341 11477 375
rect 11535 334 11569 368
rect 11619 318 11653 352
rect 11723 334 11757 368
rect 11109 248 11143 282
rect 11723 266 11757 300
rect 11807 318 11841 352
rect 11891 334 11925 368
rect 11891 266 11925 300
rect 11995 306 12029 340
rect 11995 238 12029 272
rect 12079 330 12113 364
rect 12079 262 12113 296
rect 12174 324 12208 358
rect 12174 256 12208 290
rect 12278 305 12312 339
rect 12278 237 12312 271
rect 12362 342 12396 376
rect 12564 342 12598 376
rect 12460 206 12494 240
rect 12730 316 12764 350
rect 12838 342 12872 376
rect 13052 341 13086 375
rect 13327 342 13361 376
rect 13327 274 13361 308
rect 13501 316 13535 350
rect 13621 332 13655 366
rect 13835 341 13869 375
rect 13927 334 13961 368
rect 14011 318 14045 352
rect 14115 334 14149 368
rect 13501 248 13535 282
rect 14115 266 14149 300
rect 14199 318 14233 352
rect 14283 334 14317 368
rect 14283 266 14317 300
rect 14387 306 14421 340
rect 14387 238 14421 272
rect 14471 330 14505 364
rect 14471 262 14505 296
rect 14566 324 14600 358
rect 14566 256 14600 290
rect 14670 305 14704 339
rect 14670 237 14704 271
rect 14754 342 14788 376
rect 14956 342 14990 376
rect 14852 206 14886 240
rect 15122 316 15156 350
rect 15230 342 15264 376
rect 15444 341 15478 375
rect 15719 342 15753 376
rect 15719 274 15753 308
rect 15893 316 15927 350
rect 16013 332 16047 366
rect 16227 341 16261 375
rect 16319 334 16353 368
rect 16403 318 16437 352
rect 16507 334 16541 368
rect 15893 248 15927 282
rect 16507 266 16541 300
rect 16591 318 16625 352
rect 16675 334 16709 368
rect 16675 266 16709 300
<< psubdiff >>
rect 2 2369 31 2403
rect 65 2369 123 2403
rect 157 2369 215 2403
rect 249 2369 307 2403
rect 341 2369 399 2403
rect 433 2369 491 2403
rect 525 2369 583 2403
rect 617 2369 675 2403
rect 709 2369 767 2403
rect 801 2369 859 2403
rect 893 2369 951 2403
rect 985 2369 1043 2403
rect 1077 2369 1135 2403
rect 1169 2369 1227 2403
rect 1261 2369 1319 2403
rect 1353 2369 1411 2403
rect 1445 2369 1503 2403
rect 1537 2369 1595 2403
rect 1629 2369 1687 2403
rect 1721 2369 1779 2403
rect 1813 2369 1871 2403
rect 1905 2369 1963 2403
rect 1997 2369 2055 2403
rect 2089 2369 2147 2403
rect 2181 2369 2239 2403
rect 2273 2369 2331 2403
rect 2365 2369 2423 2403
rect 2457 2369 2515 2403
rect 2549 2369 2607 2403
rect 2641 2369 2699 2403
rect 2733 2369 2791 2403
rect 2825 2369 2854 2403
rect 4386 2369 4415 2403
rect 4449 2369 4507 2403
rect 4541 2369 4599 2403
rect 4633 2369 4691 2403
rect 4725 2369 4783 2403
rect 4817 2369 4875 2403
rect 4909 2369 4967 2403
rect 5001 2369 5059 2403
rect 5093 2369 5151 2403
rect 5185 2369 5243 2403
rect 5277 2369 5335 2403
rect 5369 2369 5427 2403
rect 5461 2369 5519 2403
rect 5553 2369 5611 2403
rect 5645 2369 5703 2403
rect 5737 2369 5795 2403
rect 5829 2369 5887 2403
rect 5921 2369 5979 2403
rect 6013 2369 6071 2403
rect 6105 2369 6163 2403
rect 6197 2369 6255 2403
rect 6289 2369 6347 2403
rect 6381 2369 6439 2403
rect 6473 2369 6531 2403
rect 6565 2369 6623 2403
rect 6657 2369 6715 2403
rect 6749 2369 6807 2403
rect 6841 2369 6899 2403
rect 6933 2369 6991 2403
rect 7025 2369 7083 2403
rect 7117 2369 7175 2403
rect 7209 2369 7238 2403
rect 0 1227 29 1261
rect 63 1227 121 1261
rect 155 1227 213 1261
rect 247 1227 305 1261
rect 339 1227 397 1261
rect 431 1227 489 1261
rect 523 1227 581 1261
rect 615 1227 673 1261
rect 707 1227 765 1261
rect 799 1227 857 1261
rect 891 1227 949 1261
rect 983 1227 1041 1261
rect 1075 1227 1133 1261
rect 1167 1227 1225 1261
rect 1259 1227 1317 1261
rect 1351 1227 1409 1261
rect 1443 1227 1501 1261
rect 1535 1227 1593 1261
rect 1627 1227 1685 1261
rect 1719 1227 1777 1261
rect 1811 1227 1869 1261
rect 1903 1227 1961 1261
rect 1995 1227 2053 1261
rect 2087 1227 2145 1261
rect 2179 1227 2237 1261
rect 2271 1227 2329 1261
rect 2363 1227 2421 1261
rect 2455 1227 2513 1261
rect 2547 1227 2605 1261
rect 2639 1227 2697 1261
rect 2731 1227 2789 1261
rect 2823 1227 2881 1261
rect 2915 1227 2973 1261
rect 3007 1227 3065 1261
rect 3099 1227 3157 1261
rect 3191 1227 3249 1261
rect 3283 1227 3341 1261
rect 3375 1227 3433 1261
rect 3467 1227 3525 1261
rect 3559 1227 3617 1261
rect 3651 1227 3709 1261
rect 3743 1227 3801 1261
rect 3835 1227 3893 1261
rect 3927 1227 3985 1261
rect 4019 1227 4077 1261
rect 4111 1227 4169 1261
rect 4203 1227 4261 1261
rect 4295 1227 4353 1261
rect 4387 1227 4445 1261
rect 4479 1227 4537 1261
rect 4571 1227 4629 1261
rect 4663 1227 4721 1261
rect 4755 1227 4813 1261
rect 4847 1227 4905 1261
rect 4939 1227 4997 1261
rect 5031 1227 5089 1261
rect 5123 1227 5181 1261
rect 5215 1227 5273 1261
rect 5307 1227 5365 1261
rect 5399 1227 5457 1261
rect 5491 1227 5549 1261
rect 5583 1227 5641 1261
rect 5675 1231 6245 1261
rect 5675 1227 5704 1231
rect 6216 1227 6245 1231
rect 6279 1227 6337 1261
rect 6371 1227 6429 1261
rect 6463 1227 6521 1261
rect 6555 1227 6613 1261
rect 6647 1227 6705 1261
rect 6739 1227 6797 1261
rect 6831 1227 6889 1261
rect 6923 1227 6981 1261
rect 7015 1227 7073 1261
rect 7107 1227 7165 1261
rect 7199 1227 7257 1261
rect 7291 1227 7349 1261
rect 7383 1227 7441 1261
rect 7475 1227 7533 1261
rect 7567 1227 7625 1261
rect 7659 1227 7717 1261
rect 7751 1227 7809 1261
rect 7843 1227 7901 1261
rect 7935 1227 7993 1261
rect 8027 1227 8085 1261
rect 8119 1227 8177 1261
rect 8211 1227 8269 1261
rect 8303 1227 8361 1261
rect 8395 1227 8453 1261
rect 8487 1227 8545 1261
rect 8579 1227 8637 1261
rect 8671 1227 8729 1261
rect 8763 1227 8821 1261
rect 8855 1227 8913 1261
rect 8947 1227 9005 1261
rect 9039 1227 9097 1261
rect 9131 1227 9189 1261
rect 9223 1227 9281 1261
rect 9315 1227 9373 1261
rect 9407 1227 9465 1261
rect 9499 1227 9557 1261
rect 9591 1227 9649 1261
rect 9683 1227 9741 1261
rect 9775 1227 9833 1261
rect 9867 1227 9925 1261
rect 9959 1227 10017 1261
rect 10051 1227 10109 1261
rect 10143 1227 10201 1261
rect 10235 1227 10293 1261
rect 10327 1227 10385 1261
rect 10419 1227 10477 1261
rect 10511 1227 10569 1261
rect 10603 1227 10661 1261
rect 10695 1227 10753 1261
rect 10787 1227 10845 1261
rect 10879 1227 10937 1261
rect 10971 1227 11029 1261
rect 11063 1227 11121 1261
rect 11155 1227 11213 1261
rect 11247 1227 11305 1261
rect 11339 1227 11397 1261
rect 11431 1227 11489 1261
rect 11523 1227 11581 1261
rect 11615 1227 11673 1261
rect 11707 1227 11765 1261
rect 11799 1227 11857 1261
rect 11891 1231 12011 1261
rect 11891 1227 11920 1231
rect 11982 1227 12011 1231
rect 12045 1227 12103 1261
rect 12137 1227 12195 1261
rect 12229 1227 12287 1261
rect 12321 1227 12379 1261
rect 12413 1227 12471 1261
rect 12505 1227 12563 1261
rect 12597 1227 12655 1261
rect 12689 1227 12747 1261
rect 12781 1227 12839 1261
rect 12873 1227 12931 1261
rect 12965 1227 13023 1261
rect 13057 1227 13115 1261
rect 13149 1227 13207 1261
rect 13241 1227 13299 1261
rect 13333 1227 13391 1261
rect 13425 1227 13483 1261
rect 13517 1227 13575 1261
rect 13609 1227 13667 1261
rect 13701 1227 13759 1261
rect 13793 1227 13851 1261
rect 13885 1227 13943 1261
rect 13977 1227 14035 1261
rect 14069 1227 14127 1261
rect 14161 1227 14219 1261
rect 14253 1227 14311 1261
rect 14345 1227 14403 1261
rect 14437 1227 14495 1261
rect 14529 1227 14587 1261
rect 14621 1227 14679 1261
rect 14713 1227 14771 1261
rect 14805 1227 14863 1261
rect 14897 1227 14955 1261
rect 14989 1227 15047 1261
rect 15081 1227 15139 1261
rect 15173 1227 15231 1261
rect 15265 1227 15323 1261
rect 15357 1227 15415 1261
rect 15449 1227 15507 1261
rect 15541 1227 15599 1261
rect 15633 1227 15691 1261
rect 15725 1227 15783 1261
rect 15817 1227 15875 1261
rect 15909 1227 15967 1261
rect 16001 1227 16059 1261
rect 16093 1227 16151 1261
rect 16185 1227 16243 1261
rect 16277 1227 16335 1261
rect 16369 1227 16427 1261
rect 16461 1227 16519 1261
rect 16553 1231 16614 1261
rect 16553 1227 16582 1231
rect -1 543 29 573
rect 0 539 29 543
rect 63 539 121 573
rect 155 539 213 573
rect 247 539 305 573
rect 339 539 397 573
rect 431 539 489 573
rect 523 539 581 573
rect 615 539 673 573
rect 707 539 765 573
rect 799 539 857 573
rect 891 539 949 573
rect 983 539 1041 573
rect 1075 539 1133 573
rect 1167 539 1225 573
rect 1259 539 1317 573
rect 1351 539 1409 573
rect 1443 539 1501 573
rect 1535 539 1593 573
rect 1627 539 1685 573
rect 1719 539 1777 573
rect 1811 539 1869 573
rect 1903 539 1961 573
rect 1995 539 2053 573
rect 2087 539 2145 573
rect 2179 539 2237 573
rect 2271 539 2329 573
rect 2363 539 2421 573
rect 2455 539 2513 573
rect 2547 539 2605 573
rect 2639 539 2697 573
rect 2731 539 2789 573
rect 2823 539 2881 573
rect 2915 539 2973 573
rect 3007 539 3065 573
rect 3099 539 3157 573
rect 3191 539 3249 573
rect 3283 539 3341 573
rect 3375 539 3433 573
rect 3467 539 3525 573
rect 3559 539 3617 573
rect 3651 539 3709 573
rect 3743 539 3801 573
rect 3835 539 3893 573
rect 3927 539 3985 573
rect 4019 539 4077 573
rect 4111 539 4169 573
rect 4203 539 4261 573
rect 4295 539 4353 573
rect 4387 539 4445 573
rect 4479 539 4537 573
rect 4571 539 4629 573
rect 4663 539 4721 573
rect 4755 539 4813 573
rect 4847 539 4905 573
rect 4939 539 4997 573
rect 5031 539 5089 573
rect 5123 539 5181 573
rect 5215 539 5273 573
rect 5307 539 5365 573
rect 5399 539 5457 573
rect 5491 539 5549 573
rect 5583 539 5641 573
rect 5675 539 5733 573
rect 5767 539 5825 573
rect 5859 539 5917 573
rect 5951 539 6009 573
rect 6043 539 6101 573
rect 6135 539 6193 573
rect 6227 539 6285 573
rect 6319 539 6377 573
rect 6411 539 6469 573
rect 6503 539 6561 573
rect 6595 539 6653 573
rect 6687 539 6745 573
rect 6779 539 6837 573
rect 6871 539 6929 573
rect 6963 539 7021 573
rect 7055 539 7113 573
rect 7147 539 7205 573
rect 7239 539 7297 573
rect 7331 539 7389 573
rect 7423 539 7481 573
rect 7515 539 7573 573
rect 7607 539 7665 573
rect 7699 539 7757 573
rect 7791 539 7849 573
rect 7883 539 7941 573
rect 7975 539 8033 573
rect 8067 539 8125 573
rect 8159 539 8217 573
rect 8251 539 8309 573
rect 8343 539 8401 573
rect 8435 539 8493 573
rect 8527 539 8585 573
rect 8619 539 8677 573
rect 8711 539 8769 573
rect 8803 539 8861 573
rect 8895 539 8953 573
rect 8987 539 9045 573
rect 9079 539 9137 573
rect 9171 539 9229 573
rect 9263 539 9321 573
rect 9355 539 9413 573
rect 9447 539 9505 573
rect 9539 539 9597 573
rect 9631 539 9689 573
rect 9723 539 9781 573
rect 9815 539 9873 573
rect 9907 539 9965 573
rect 9999 539 10057 573
rect 10091 539 10149 573
rect 10183 539 10241 573
rect 10275 539 10333 573
rect 10367 539 10425 573
rect 10459 539 10517 573
rect 10551 539 10609 573
rect 10643 539 10701 573
rect 10735 539 10793 573
rect 10827 539 10885 573
rect 10919 539 10977 573
rect 11011 539 11069 573
rect 11103 539 11161 573
rect 11195 539 11253 573
rect 11287 539 11345 573
rect 11379 539 11437 573
rect 11471 539 11529 573
rect 11563 539 11621 573
rect 11655 539 11713 573
rect 11747 539 11805 573
rect 11839 539 11897 573
rect 11931 539 11989 573
rect 12023 539 12081 573
rect 12115 539 12173 573
rect 12207 539 12265 573
rect 12299 539 12357 573
rect 12391 539 12449 573
rect 12483 539 12541 573
rect 12575 539 12633 573
rect 12667 539 12725 573
rect 12759 539 12817 573
rect 12851 539 12909 573
rect 12943 539 13001 573
rect 13035 539 13093 573
rect 13127 539 13185 573
rect 13219 539 13277 573
rect 13311 539 13369 573
rect 13403 539 13461 573
rect 13495 539 13553 573
rect 13587 539 13645 573
rect 13679 539 13737 573
rect 13771 539 13829 573
rect 13863 539 13921 573
rect 13955 539 14013 573
rect 14047 539 14105 573
rect 14139 539 14197 573
rect 14231 539 14289 573
rect 14323 539 14381 573
rect 14415 539 14473 573
rect 14507 539 14565 573
rect 14599 539 14657 573
rect 14691 539 14749 573
rect 14783 539 14841 573
rect 14875 539 14933 573
rect 14967 539 15025 573
rect 15059 539 15117 573
rect 15151 539 15209 573
rect 15243 539 15301 573
rect 15335 539 15393 573
rect 15427 539 15485 573
rect 15519 539 15577 573
rect 15611 539 15669 573
rect 15703 539 15761 573
rect 15795 539 15853 573
rect 15887 539 15945 573
rect 15979 539 16037 573
rect 16071 539 16129 573
rect 16163 539 16221 573
rect 16255 539 16313 573
rect 16347 539 16405 573
rect 16439 539 16497 573
rect 16531 539 16589 573
rect 16623 539 16681 573
rect 16715 539 16744 573
rect 0 -150 29 -116
rect 63 -150 121 -116
rect 155 -150 213 -116
rect 247 -150 305 -116
rect 339 -150 397 -116
rect 431 -150 489 -116
rect 523 -150 581 -116
rect 615 -150 673 -116
rect 707 -150 765 -116
rect 799 -150 857 -116
rect 891 -150 949 -116
rect 983 -150 1041 -116
rect 1075 -150 1133 -116
rect 1167 -150 1225 -116
rect 1259 -150 1317 -116
rect 1351 -150 1409 -116
rect 1443 -150 1501 -116
rect 1535 -150 1593 -116
rect 1627 -150 1685 -116
rect 1719 -150 1777 -116
rect 1811 -150 1869 -116
rect 1903 -150 1961 -116
rect 1995 -150 2053 -116
rect 2087 -150 2145 -116
rect 2179 -150 2237 -116
rect 2271 -150 2329 -116
rect 2363 -150 2421 -116
rect 2455 -150 2513 -116
rect 2547 -150 2605 -116
rect 2639 -150 2697 -116
rect 2731 -150 2789 -116
rect 2823 -150 2881 -116
rect 2915 -150 2973 -116
rect 3007 -150 3065 -116
rect 3099 -150 3157 -116
rect 3191 -150 3249 -116
rect 3283 -150 3341 -116
rect 3375 -150 3433 -116
rect 3467 -150 3525 -116
rect 3559 -150 3617 -116
rect 3651 -150 3709 -116
rect 3743 -150 3801 -116
rect 3835 -150 3893 -116
rect 3927 -150 3985 -116
rect 4019 -150 4077 -116
rect 4111 -150 4169 -116
rect 4203 -150 4261 -116
rect 4295 -150 4353 -116
rect 4387 -150 4445 -116
rect 4479 -150 4537 -116
rect 4571 -150 4629 -116
rect 4663 -150 4721 -116
rect 4755 -150 4813 -116
rect 4847 -150 4905 -116
rect 4939 -150 4997 -116
rect 5031 -150 5089 -116
rect 5123 -150 5181 -116
rect 5215 -150 5273 -116
rect 5307 -150 5365 -116
rect 5399 -150 5457 -116
rect 5491 -150 5549 -116
rect 5583 -150 5641 -116
rect 5675 -150 5733 -116
rect 5767 -150 5825 -116
rect 5859 -150 5917 -116
rect 5951 -150 6009 -116
rect 6043 -150 6101 -116
rect 6135 -150 6193 -116
rect 6227 -150 6285 -116
rect 6319 -150 6377 -116
rect 6411 -150 6469 -116
rect 6503 -150 6561 -116
rect 6595 -150 6653 -116
rect 6687 -150 6745 -116
rect 6779 -150 6837 -116
rect 6871 -150 6929 -116
rect 6963 -150 7021 -116
rect 7055 -150 7113 -116
rect 7147 -150 7205 -116
rect 7239 -150 7297 -116
rect 7331 -150 7389 -116
rect 7423 -150 7481 -116
rect 7515 -150 7573 -116
rect 7607 -150 7665 -116
rect 7699 -150 7757 -116
rect 7791 -150 7849 -116
rect 7883 -150 7941 -116
rect 7975 -150 8033 -116
rect 8067 -150 8125 -116
rect 8159 -150 8217 -116
rect 8251 -150 8309 -116
rect 8343 -150 8401 -116
rect 8435 -150 8493 -116
rect 8527 -150 8585 -116
rect 8619 -150 8677 -116
rect 8711 -150 8769 -116
rect 8803 -150 8861 -116
rect 8895 -150 8953 -116
rect 8987 -150 9045 -116
rect 9079 -150 9137 -116
rect 9171 -150 9229 -116
rect 9263 -150 9321 -116
rect 9355 -150 9413 -116
rect 9447 -150 9505 -116
rect 9539 -150 9597 -116
rect 9631 -150 9689 -116
rect 9723 -150 9781 -116
rect 9815 -150 9873 -116
rect 9907 -150 9965 -116
rect 9999 -150 10057 -116
rect 10091 -150 10149 -116
rect 10183 -150 10241 -116
rect 10275 -150 10333 -116
rect 10367 -150 10425 -116
rect 10459 -150 10517 -116
rect 10551 -150 10609 -116
rect 10643 -150 10701 -116
rect 10735 -150 10793 -116
rect 10827 -150 10885 -116
rect 10919 -150 10977 -116
rect 11011 -150 11069 -116
rect 11103 -150 11161 -116
rect 11195 -150 11253 -116
rect 11287 -150 11345 -116
rect 11379 -150 11437 -116
rect 11471 -150 11529 -116
rect 11563 -150 11621 -116
rect 11655 -150 11713 -116
rect 11747 -150 11805 -116
rect 11839 -150 11897 -116
rect 11931 -150 11989 -116
rect 12023 -150 12081 -116
rect 12115 -150 12173 -116
rect 12207 -150 12265 -116
rect 12299 -150 12357 -116
rect 12391 -150 12449 -116
rect 12483 -150 12541 -116
rect 12575 -150 12633 -116
rect 12667 -150 12725 -116
rect 12759 -150 12817 -116
rect 12851 -150 12909 -116
rect 12943 -150 13001 -116
rect 13035 -150 13093 -116
rect 13127 -150 13185 -116
rect 13219 -150 13277 -116
rect 13311 -150 13369 -116
rect 13403 -150 13461 -116
rect 13495 -150 13553 -116
rect 13587 -150 13645 -116
rect 13679 -150 13737 -116
rect 13771 -150 13829 -116
rect 13863 -150 13921 -116
rect 13955 -150 14013 -116
rect 14047 -150 14105 -116
rect 14139 -150 14197 -116
rect 14231 -150 14289 -116
rect 14323 -150 14381 -116
rect 14415 -150 14473 -116
rect 14507 -150 14565 -116
rect 14599 -150 14657 -116
rect 14691 -150 14749 -116
rect 14783 -150 14841 -116
rect 14875 -150 14933 -116
rect 14967 -150 15025 -116
rect 15059 -150 15117 -116
rect 15151 -150 15209 -116
rect 15243 -150 15301 -116
rect 15335 -150 15393 -116
rect 15427 -150 15485 -116
rect 15519 -150 15577 -116
rect 15611 -150 15669 -116
rect 15703 -150 15761 -116
rect 15795 -150 15853 -116
rect 15887 -150 15945 -116
rect 15979 -150 16037 -116
rect 16071 -150 16129 -116
rect 16163 -150 16221 -116
rect 16255 -150 16313 -116
rect 16347 -150 16405 -116
rect 16439 -150 16497 -116
rect 16531 -150 16589 -116
rect 16623 -150 16681 -116
rect 16715 -150 16744 -116
<< nsubdiff >>
rect 2 2961 31 2995
rect 65 2961 123 2995
rect 157 2961 215 2995
rect 249 2961 307 2995
rect 341 2961 399 2995
rect 433 2961 491 2995
rect 525 2961 583 2995
rect 617 2961 675 2995
rect 709 2961 767 2995
rect 801 2961 859 2995
rect 893 2961 951 2995
rect 985 2961 1043 2995
rect 1077 2961 1135 2995
rect 1169 2961 1227 2995
rect 1261 2961 1319 2995
rect 1353 2961 1411 2995
rect 1445 2961 1503 2995
rect 1537 2961 1595 2995
rect 1629 2961 1687 2995
rect 1721 2961 1779 2995
rect 1813 2961 1871 2995
rect 1905 2961 1963 2995
rect 1997 2961 2055 2995
rect 2089 2961 2147 2995
rect 2181 2961 2239 2995
rect 2273 2961 2331 2995
rect 2365 2961 2423 2995
rect 2457 2961 2515 2995
rect 2549 2961 2607 2995
rect 2641 2961 2699 2995
rect 2733 2961 2791 2995
rect 2825 2961 2854 2995
rect 4386 2961 4415 2995
rect 4449 2961 4507 2995
rect 4541 2961 4599 2995
rect 4633 2961 4691 2995
rect 4725 2961 4783 2995
rect 4817 2961 4875 2995
rect 4909 2961 4967 2995
rect 5001 2961 5059 2995
rect 5093 2961 5151 2995
rect 5185 2961 5243 2995
rect 5277 2961 5335 2995
rect 5369 2961 5427 2995
rect 5461 2961 5519 2995
rect 5553 2961 5611 2995
rect 5645 2961 5703 2995
rect 5737 2961 5795 2995
rect 5829 2961 5887 2995
rect 5921 2961 5979 2995
rect 6013 2961 6071 2995
rect 6105 2961 6163 2995
rect 6197 2961 6255 2995
rect 6289 2961 6347 2995
rect 6381 2961 6439 2995
rect 6473 2961 6531 2995
rect 6565 2961 6623 2995
rect 6657 2961 6715 2995
rect 6749 2961 6807 2995
rect 6841 2961 6899 2995
rect 6933 2961 6991 2995
rect 7025 2961 7083 2995
rect 7117 2961 7175 2995
rect 7209 2961 7238 2995
rect 0 1819 29 1853
rect 63 1819 121 1853
rect 155 1819 213 1853
rect 247 1819 305 1853
rect 339 1819 397 1853
rect 431 1819 489 1853
rect 523 1819 581 1853
rect 615 1819 673 1853
rect 707 1819 765 1853
rect 799 1819 857 1853
rect 891 1819 949 1853
rect 983 1819 1041 1853
rect 1075 1819 1133 1853
rect 1167 1819 1225 1853
rect 1259 1819 1317 1853
rect 1351 1819 1409 1853
rect 1443 1819 1501 1853
rect 1535 1819 1593 1853
rect 1627 1819 1685 1853
rect 1719 1819 1777 1853
rect 1811 1819 1869 1853
rect 1903 1819 1961 1853
rect 1995 1819 2053 1853
rect 2087 1819 2145 1853
rect 2179 1819 2237 1853
rect 2271 1819 2329 1853
rect 2363 1819 2421 1853
rect 2455 1819 2513 1853
rect 2547 1819 2605 1853
rect 2639 1819 2697 1853
rect 2731 1819 2789 1853
rect 2823 1819 2881 1853
rect 2915 1819 2973 1853
rect 3007 1819 3065 1853
rect 3099 1819 3157 1853
rect 3191 1819 3249 1853
rect 3283 1819 3341 1853
rect 3375 1819 3433 1853
rect 3467 1819 3525 1853
rect 3559 1819 3617 1853
rect 3651 1819 3709 1853
rect 3743 1819 3801 1853
rect 3835 1819 3893 1853
rect 3927 1819 3985 1853
rect 4019 1819 4077 1853
rect 4111 1819 4169 1853
rect 4203 1819 4261 1853
rect 4295 1819 4353 1853
rect 4387 1819 4445 1853
rect 4479 1819 4537 1853
rect 4571 1819 4629 1853
rect 4663 1819 4721 1853
rect 4755 1819 4813 1853
rect 4847 1819 4905 1853
rect 4939 1819 4997 1853
rect 5031 1819 5089 1853
rect 5123 1819 5181 1853
rect 5215 1819 5273 1853
rect 5307 1819 5365 1853
rect 5399 1819 5457 1853
rect 5491 1819 5549 1853
rect 5583 1819 5641 1853
rect 5675 1849 5704 1853
rect 6216 1849 6245 1853
rect 5675 1819 6245 1849
rect 6279 1819 6337 1853
rect 6371 1819 6429 1853
rect 6463 1819 6521 1853
rect 6555 1819 6613 1853
rect 6647 1819 6705 1853
rect 6739 1819 6797 1853
rect 6831 1819 6889 1853
rect 6923 1819 6981 1853
rect 7015 1819 7073 1853
rect 7107 1819 7165 1853
rect 7199 1819 7257 1853
rect 7291 1819 7349 1853
rect 7383 1819 7441 1853
rect 7475 1819 7533 1853
rect 7567 1819 7625 1853
rect 7659 1819 7717 1853
rect 7751 1819 7809 1853
rect 7843 1819 7901 1853
rect 7935 1819 7993 1853
rect 8027 1819 8085 1853
rect 8119 1819 8177 1853
rect 8211 1819 8269 1853
rect 8303 1819 8361 1853
rect 8395 1819 8453 1853
rect 8487 1819 8545 1853
rect 8579 1819 8637 1853
rect 8671 1819 8729 1853
rect 8763 1819 8821 1853
rect 8855 1819 8913 1853
rect 8947 1819 9005 1853
rect 9039 1819 9097 1853
rect 9131 1819 9189 1853
rect 9223 1819 9281 1853
rect 9315 1819 9373 1853
rect 9407 1819 9465 1853
rect 9499 1819 9557 1853
rect 9591 1819 9649 1853
rect 9683 1819 9741 1853
rect 9775 1819 9833 1853
rect 9867 1819 9925 1853
rect 9959 1819 10017 1853
rect 10051 1819 10109 1853
rect 10143 1819 10201 1853
rect 10235 1819 10293 1853
rect 10327 1819 10385 1853
rect 10419 1819 10477 1853
rect 10511 1819 10569 1853
rect 10603 1819 10661 1853
rect 10695 1819 10753 1853
rect 10787 1819 10845 1853
rect 10879 1819 10937 1853
rect 10971 1819 11029 1853
rect 11063 1819 11121 1853
rect 11155 1819 11213 1853
rect 11247 1819 11305 1853
rect 11339 1819 11397 1853
rect 11431 1819 11489 1853
rect 11523 1819 11581 1853
rect 11615 1819 11673 1853
rect 11707 1819 11765 1853
rect 11799 1819 11857 1853
rect 11891 1849 11920 1853
rect 11982 1849 12011 1853
rect 11891 1819 12011 1849
rect 12045 1819 12103 1853
rect 12137 1819 12195 1853
rect 12229 1819 12287 1853
rect 12321 1819 12379 1853
rect 12413 1819 12471 1853
rect 12505 1819 12563 1853
rect 12597 1819 12655 1853
rect 12689 1819 12747 1853
rect 12781 1819 12839 1853
rect 12873 1819 12931 1853
rect 12965 1819 13023 1853
rect 13057 1819 13115 1853
rect 13149 1819 13207 1853
rect 13241 1819 13299 1853
rect 13333 1819 13391 1853
rect 13425 1819 13483 1853
rect 13517 1819 13575 1853
rect 13609 1819 13667 1853
rect 13701 1819 13759 1853
rect 13793 1819 13851 1853
rect 13885 1819 13943 1853
rect 13977 1819 14035 1853
rect 14069 1819 14127 1853
rect 14161 1819 14219 1853
rect 14253 1819 14311 1853
rect 14345 1819 14403 1853
rect 14437 1819 14495 1853
rect 14529 1819 14587 1853
rect 14621 1819 14679 1853
rect 14713 1819 14771 1853
rect 14805 1819 14863 1853
rect 14897 1819 14955 1853
rect 14989 1819 15047 1853
rect 15081 1819 15139 1853
rect 15173 1819 15231 1853
rect 15265 1819 15323 1853
rect 15357 1819 15415 1853
rect 15449 1819 15507 1853
rect 15541 1819 15599 1853
rect 15633 1819 15691 1853
rect 15725 1819 15783 1853
rect 15817 1819 15875 1853
rect 15909 1819 15967 1853
rect 16001 1819 16059 1853
rect 16093 1819 16151 1853
rect 16185 1819 16243 1853
rect 16277 1819 16335 1853
rect 16369 1819 16427 1853
rect 16461 1819 16519 1853
rect 16553 1849 16582 1853
rect 16553 1819 16614 1849
rect 3704 1804 3757 1819
rect 1 1161 29 1165
rect -1 1131 29 1161
rect 63 1131 121 1165
rect 155 1131 213 1165
rect 247 1131 305 1165
rect 339 1131 397 1165
rect 431 1131 489 1165
rect 523 1131 581 1165
rect 615 1131 673 1165
rect 707 1131 765 1165
rect 799 1131 857 1165
rect 891 1131 949 1165
rect 983 1131 1041 1165
rect 1075 1131 1133 1165
rect 1167 1131 1225 1165
rect 1259 1131 1317 1165
rect 1351 1131 1409 1165
rect 1443 1131 1501 1165
rect 1535 1131 1593 1165
rect 1627 1131 1685 1165
rect 1719 1131 1777 1165
rect 1811 1161 1835 1165
rect 1811 1131 1843 1161
rect 2029 1161 2053 1165
rect 1995 1131 2053 1161
rect 2087 1131 2145 1165
rect 2179 1131 2237 1165
rect 2271 1131 2329 1165
rect 2363 1131 2421 1165
rect 2455 1131 2513 1165
rect 2547 1131 2605 1165
rect 2639 1131 2697 1165
rect 2731 1131 2789 1165
rect 2823 1131 2881 1165
rect 2915 1131 2973 1165
rect 3007 1131 3065 1165
rect 3099 1131 3157 1165
rect 3191 1131 3249 1165
rect 3283 1131 3341 1165
rect 3375 1131 3433 1165
rect 3467 1131 3525 1165
rect 3559 1131 3617 1165
rect 3651 1131 3709 1165
rect 3743 1131 3801 1165
rect 3835 1131 3893 1165
rect 3927 1131 3985 1165
rect 4019 1131 4077 1165
rect 4111 1131 4169 1165
rect 4203 1161 4227 1165
rect 4203 1131 4254 1161
rect 4421 1161 4445 1165
rect 4387 1131 4445 1161
rect 4479 1131 4537 1165
rect 4571 1131 4629 1165
rect 4663 1131 4721 1165
rect 4755 1131 4813 1165
rect 4847 1131 4905 1165
rect 4939 1131 4997 1165
rect 5031 1131 5089 1165
rect 5123 1131 5181 1165
rect 5215 1131 5273 1165
rect 5307 1131 5365 1165
rect 5399 1131 5457 1165
rect 5491 1131 5549 1165
rect 5583 1131 5641 1165
rect 5675 1131 5733 1165
rect 5767 1131 5825 1165
rect 5859 1131 5917 1165
rect 5951 1131 6009 1165
rect 6043 1131 6101 1165
rect 6135 1131 6193 1165
rect 6227 1131 6285 1165
rect 6319 1131 6377 1165
rect 6411 1131 6469 1165
rect 6503 1131 6561 1165
rect 6595 1161 6619 1165
rect 6595 1131 6643 1161
rect 6813 1161 6837 1165
rect 6779 1131 6837 1161
rect 6871 1131 6929 1165
rect 6963 1131 7021 1165
rect 7055 1131 7113 1165
rect 7147 1131 7205 1165
rect 7239 1131 7297 1165
rect 7331 1131 7389 1165
rect 7423 1131 7481 1165
rect 7515 1131 7573 1165
rect 7607 1131 7665 1165
rect 7699 1131 7757 1165
rect 7791 1131 7849 1165
rect 7883 1131 7941 1165
rect 7975 1131 8033 1165
rect 8067 1131 8125 1165
rect 8159 1131 8217 1165
rect 8251 1131 8309 1165
rect 8343 1131 8401 1165
rect 8435 1131 8493 1165
rect 8527 1131 8585 1165
rect 8619 1131 8677 1165
rect 8711 1131 8769 1165
rect 8803 1131 8861 1165
rect 8895 1131 8953 1165
rect 8987 1161 9011 1165
rect 8987 1131 9037 1161
rect 9205 1161 9229 1165
rect 9171 1131 9229 1161
rect 9263 1131 9321 1165
rect 9355 1131 9413 1165
rect 9447 1131 9505 1165
rect 9539 1131 9597 1165
rect 9631 1131 9689 1165
rect 9723 1131 9781 1165
rect 9815 1131 9873 1165
rect 9907 1131 9965 1165
rect 9999 1131 10057 1165
rect 10091 1131 10149 1165
rect 10183 1131 10241 1165
rect 10275 1131 10333 1165
rect 10367 1131 10425 1165
rect 10459 1131 10517 1165
rect 10551 1131 10609 1165
rect 10643 1131 10701 1165
rect 10735 1131 10793 1165
rect 10827 1131 10885 1165
rect 10919 1131 10977 1165
rect 11011 1131 11069 1165
rect 11103 1131 11161 1165
rect 11195 1131 11253 1165
rect 11287 1131 11345 1165
rect 11379 1161 11403 1165
rect 11379 1131 11427 1161
rect 11597 1161 11621 1165
rect 11563 1131 11621 1161
rect 11655 1131 11713 1165
rect 11747 1131 11805 1165
rect 11839 1131 11897 1165
rect 11931 1131 11989 1165
rect 12023 1131 12081 1165
rect 12115 1131 12173 1165
rect 12207 1131 12265 1165
rect 12299 1131 12357 1165
rect 12391 1131 12449 1165
rect 12483 1131 12541 1165
rect 12575 1131 12633 1165
rect 12667 1131 12725 1165
rect 12759 1131 12817 1165
rect 12851 1131 12909 1165
rect 12943 1131 13001 1165
rect 13035 1131 13093 1165
rect 13127 1131 13185 1165
rect 13219 1131 13277 1165
rect 13311 1131 13369 1165
rect 13403 1131 13461 1165
rect 13495 1131 13553 1165
rect 13587 1131 13645 1165
rect 13679 1131 13737 1165
rect 13771 1161 13795 1165
rect 13771 1131 13819 1161
rect 13989 1161 14013 1165
rect 13955 1131 14013 1161
rect 14047 1131 14105 1165
rect 14139 1131 14197 1165
rect 14231 1131 14289 1165
rect 14323 1131 14381 1165
rect 14415 1131 14473 1165
rect 14507 1131 14565 1165
rect 14599 1131 14657 1165
rect 14691 1131 14749 1165
rect 14783 1131 14841 1165
rect 14875 1131 14933 1165
rect 14967 1131 15025 1165
rect 15059 1131 15117 1165
rect 15151 1131 15209 1165
rect 15243 1131 15301 1165
rect 15335 1131 15393 1165
rect 15427 1131 15485 1165
rect 15519 1131 15577 1165
rect 15611 1131 15669 1165
rect 15703 1131 15761 1165
rect 15795 1131 15853 1165
rect 15887 1131 15945 1165
rect 15979 1131 16037 1165
rect 16071 1131 16129 1165
rect 16163 1161 16187 1165
rect 16163 1131 16211 1161
rect 16381 1161 16405 1165
rect 16347 1131 16405 1161
rect 16439 1131 16497 1165
rect 16531 1131 16589 1165
rect 16623 1131 16681 1165
rect 16715 1131 16744 1165
rect 0 476 571 477
rect 0 442 29 476
rect 63 442 121 476
rect 155 442 213 476
rect 247 442 305 476
rect 339 442 394 476
rect 428 442 496 476
rect 530 442 581 476
rect 615 442 673 476
rect 707 442 765 476
rect 799 442 857 476
rect 891 442 949 476
rect 983 442 1041 476
rect 1075 442 1133 476
rect 1167 442 1225 476
rect 1259 442 1317 476
rect 1351 442 1409 476
rect 1443 442 1501 476
rect 1535 442 1559 476
rect 1753 442 1777 476
rect 1811 442 1869 476
rect 1903 442 1961 476
rect 1995 442 2053 476
rect 2087 442 2145 476
rect 2179 442 2237 476
rect 2271 442 2329 476
rect 2363 442 2421 476
rect 2455 442 2513 476
rect 2547 442 2605 476
rect 2639 442 2697 476
rect 2731 442 2791 476
rect 2825 442 2882 476
rect 2916 442 2973 476
rect 3007 442 3065 476
rect 3099 442 3157 476
rect 3191 442 3249 476
rect 3283 442 3341 476
rect 3375 442 3433 476
rect 3467 442 3525 476
rect 3559 442 3617 476
rect 3651 442 3709 476
rect 3743 442 3801 476
rect 3835 442 3893 476
rect 3927 442 3955 476
rect 4145 442 4169 476
rect 4203 442 4261 476
rect 4295 442 4353 476
rect 4387 442 4445 476
rect 4479 442 4537 476
rect 4571 442 4629 476
rect 4663 442 4721 476
rect 4755 442 4813 476
rect 4847 442 4905 476
rect 4939 442 4997 476
rect 5031 442 5089 476
rect 5123 442 5179 476
rect 5213 442 5273 476
rect 5307 442 5365 476
rect 5399 442 5457 476
rect 5491 442 5549 476
rect 5583 442 5641 476
rect 5675 442 5733 476
rect 5767 442 5825 476
rect 5859 442 5917 476
rect 5951 442 6009 476
rect 6043 442 6101 476
rect 6135 442 6193 476
rect 6227 442 6285 476
rect 6319 442 6353 476
rect 6518 442 6561 476
rect 6595 442 6653 476
rect 6687 442 6745 476
rect 6779 442 6837 476
rect 6871 442 6929 476
rect 6963 442 7021 476
rect 7055 442 7113 476
rect 7147 442 7205 476
rect 7239 442 7297 476
rect 7331 442 7389 476
rect 7423 442 7481 476
rect 7515 442 7574 476
rect 7608 442 7665 476
rect 7699 442 7757 476
rect 7791 442 7849 476
rect 7883 442 7941 476
rect 7975 442 8033 476
rect 8067 442 8125 476
rect 8159 442 8217 476
rect 8251 442 8309 476
rect 8343 442 8401 476
rect 8435 442 8493 476
rect 8527 442 8585 476
rect 8619 442 8677 476
rect 8711 442 8745 476
rect 8929 442 8953 476
rect 8987 442 9045 476
rect 9079 442 9137 476
rect 9171 442 9229 476
rect 9263 442 9321 476
rect 9355 442 9413 476
rect 9447 442 9505 476
rect 9539 442 9597 476
rect 9631 442 9689 476
rect 9723 442 9781 476
rect 9815 442 9873 476
rect 9907 442 9963 476
rect 9997 442 10058 476
rect 10092 442 10149 476
rect 10183 442 10241 476
rect 10275 442 10333 476
rect 10367 442 10425 476
rect 10459 442 10517 476
rect 10551 442 10609 476
rect 10643 442 10701 476
rect 10735 442 10793 476
rect 10827 442 10885 476
rect 10919 442 10977 476
rect 11011 442 11069 476
rect 11103 442 11127 476
rect 11315 442 11345 476
rect 11379 442 11437 476
rect 11471 442 11529 476
rect 11563 442 11621 476
rect 11655 442 11713 476
rect 11747 442 11805 476
rect 11839 442 11897 476
rect 11931 442 11989 476
rect 12023 442 12081 476
rect 12115 442 12173 476
rect 12207 442 12265 476
rect 12299 442 12357 476
rect 12391 442 12448 476
rect 12482 442 12541 476
rect 12575 442 12633 476
rect 12667 442 12725 476
rect 12759 442 12817 476
rect 12851 442 12909 476
rect 12943 442 13001 476
rect 13035 442 13093 476
rect 13127 442 13185 476
rect 13219 442 13277 476
rect 13311 442 13369 476
rect 13403 442 13461 476
rect 13495 442 13519 476
rect 13639 442 13737 476
rect 13771 442 13829 476
rect 13863 442 13921 476
rect 13955 442 14013 476
rect 14047 442 14105 476
rect 14139 442 14197 476
rect 14231 442 14289 476
rect 14323 442 14381 476
rect 14415 442 14473 476
rect 14507 442 14565 476
rect 14599 442 14657 476
rect 14691 442 14748 476
rect 14782 442 14842 476
rect 14876 442 14933 476
rect 14967 442 15025 476
rect 15059 442 15117 476
rect 15151 442 15209 476
rect 15243 442 15301 476
rect 15335 442 15393 476
rect 15427 442 15485 476
rect 15519 442 15577 476
rect 15611 442 15669 476
rect 15703 442 15761 476
rect 15795 442 15853 476
rect 15887 442 15921 476
rect 16031 442 16129 476
rect 16163 442 16221 476
rect 16255 442 16313 476
rect 16347 442 16405 476
rect 16439 442 16497 476
rect 16531 442 16589 476
rect 16623 442 16681 476
rect 16715 442 16744 476
<< psubdiffcont >>
rect 31 2369 65 2403
rect 123 2369 157 2403
rect 215 2369 249 2403
rect 307 2369 341 2403
rect 399 2369 433 2403
rect 491 2369 525 2403
rect 583 2369 617 2403
rect 675 2369 709 2403
rect 767 2369 801 2403
rect 859 2369 893 2403
rect 951 2369 985 2403
rect 1043 2369 1077 2403
rect 1135 2369 1169 2403
rect 1227 2369 1261 2403
rect 1319 2369 1353 2403
rect 1411 2369 1445 2403
rect 1503 2369 1537 2403
rect 1595 2369 1629 2403
rect 1687 2369 1721 2403
rect 1779 2369 1813 2403
rect 1871 2369 1905 2403
rect 1963 2369 1997 2403
rect 2055 2369 2089 2403
rect 2147 2369 2181 2403
rect 2239 2369 2273 2403
rect 2331 2369 2365 2403
rect 2423 2369 2457 2403
rect 2515 2369 2549 2403
rect 2607 2369 2641 2403
rect 2699 2369 2733 2403
rect 2791 2369 2825 2403
rect 4415 2369 4449 2403
rect 4507 2369 4541 2403
rect 4599 2369 4633 2403
rect 4691 2369 4725 2403
rect 4783 2369 4817 2403
rect 4875 2369 4909 2403
rect 4967 2369 5001 2403
rect 5059 2369 5093 2403
rect 5151 2369 5185 2403
rect 5243 2369 5277 2403
rect 5335 2369 5369 2403
rect 5427 2369 5461 2403
rect 5519 2369 5553 2403
rect 5611 2369 5645 2403
rect 5703 2369 5737 2403
rect 5795 2369 5829 2403
rect 5887 2369 5921 2403
rect 5979 2369 6013 2403
rect 6071 2369 6105 2403
rect 6163 2369 6197 2403
rect 6255 2369 6289 2403
rect 6347 2369 6381 2403
rect 6439 2369 6473 2403
rect 6531 2369 6565 2403
rect 6623 2369 6657 2403
rect 6715 2369 6749 2403
rect 6807 2369 6841 2403
rect 6899 2369 6933 2403
rect 6991 2369 7025 2403
rect 7083 2369 7117 2403
rect 7175 2369 7209 2403
rect 29 1227 63 1261
rect 121 1227 155 1261
rect 213 1227 247 1261
rect 305 1227 339 1261
rect 397 1227 431 1261
rect 489 1227 523 1261
rect 581 1227 615 1261
rect 673 1227 707 1261
rect 765 1227 799 1261
rect 857 1227 891 1261
rect 949 1227 983 1261
rect 1041 1227 1075 1261
rect 1133 1227 1167 1261
rect 1225 1227 1259 1261
rect 1317 1227 1351 1261
rect 1409 1227 1443 1261
rect 1501 1227 1535 1261
rect 1593 1227 1627 1261
rect 1685 1227 1719 1261
rect 1777 1227 1811 1261
rect 1869 1227 1903 1261
rect 1961 1227 1995 1261
rect 2053 1227 2087 1261
rect 2145 1227 2179 1261
rect 2237 1227 2271 1261
rect 2329 1227 2363 1261
rect 2421 1227 2455 1261
rect 2513 1227 2547 1261
rect 2605 1227 2639 1261
rect 2697 1227 2731 1261
rect 2789 1227 2823 1261
rect 2881 1227 2915 1261
rect 2973 1227 3007 1261
rect 3065 1227 3099 1261
rect 3157 1227 3191 1261
rect 3249 1227 3283 1261
rect 3341 1227 3375 1261
rect 3433 1227 3467 1261
rect 3525 1227 3559 1261
rect 3617 1227 3651 1261
rect 3709 1227 3743 1261
rect 3801 1227 3835 1261
rect 3893 1227 3927 1261
rect 3985 1227 4019 1261
rect 4077 1227 4111 1261
rect 4169 1227 4203 1261
rect 4261 1227 4295 1261
rect 4353 1227 4387 1261
rect 4445 1227 4479 1261
rect 4537 1227 4571 1261
rect 4629 1227 4663 1261
rect 4721 1227 4755 1261
rect 4813 1227 4847 1261
rect 4905 1227 4939 1261
rect 4997 1227 5031 1261
rect 5089 1227 5123 1261
rect 5181 1227 5215 1261
rect 5273 1227 5307 1261
rect 5365 1227 5399 1261
rect 5457 1227 5491 1261
rect 5549 1227 5583 1261
rect 5641 1227 5675 1261
rect 6245 1227 6279 1261
rect 6337 1227 6371 1261
rect 6429 1227 6463 1261
rect 6521 1227 6555 1261
rect 6613 1227 6647 1261
rect 6705 1227 6739 1261
rect 6797 1227 6831 1261
rect 6889 1227 6923 1261
rect 6981 1227 7015 1261
rect 7073 1227 7107 1261
rect 7165 1227 7199 1261
rect 7257 1227 7291 1261
rect 7349 1227 7383 1261
rect 7441 1227 7475 1261
rect 7533 1227 7567 1261
rect 7625 1227 7659 1261
rect 7717 1227 7751 1261
rect 7809 1227 7843 1261
rect 7901 1227 7935 1261
rect 7993 1227 8027 1261
rect 8085 1227 8119 1261
rect 8177 1227 8211 1261
rect 8269 1227 8303 1261
rect 8361 1227 8395 1261
rect 8453 1227 8487 1261
rect 8545 1227 8579 1261
rect 8637 1227 8671 1261
rect 8729 1227 8763 1261
rect 8821 1227 8855 1261
rect 8913 1227 8947 1261
rect 9005 1227 9039 1261
rect 9097 1227 9131 1261
rect 9189 1227 9223 1261
rect 9281 1227 9315 1261
rect 9373 1227 9407 1261
rect 9465 1227 9499 1261
rect 9557 1227 9591 1261
rect 9649 1227 9683 1261
rect 9741 1227 9775 1261
rect 9833 1227 9867 1261
rect 9925 1227 9959 1261
rect 10017 1227 10051 1261
rect 10109 1227 10143 1261
rect 10201 1227 10235 1261
rect 10293 1227 10327 1261
rect 10385 1227 10419 1261
rect 10477 1227 10511 1261
rect 10569 1227 10603 1261
rect 10661 1227 10695 1261
rect 10753 1227 10787 1261
rect 10845 1227 10879 1261
rect 10937 1227 10971 1261
rect 11029 1227 11063 1261
rect 11121 1227 11155 1261
rect 11213 1227 11247 1261
rect 11305 1227 11339 1261
rect 11397 1227 11431 1261
rect 11489 1227 11523 1261
rect 11581 1227 11615 1261
rect 11673 1227 11707 1261
rect 11765 1227 11799 1261
rect 11857 1227 11891 1261
rect 12011 1227 12045 1261
rect 12103 1227 12137 1261
rect 12195 1227 12229 1261
rect 12287 1227 12321 1261
rect 12379 1227 12413 1261
rect 12471 1227 12505 1261
rect 12563 1227 12597 1261
rect 12655 1227 12689 1261
rect 12747 1227 12781 1261
rect 12839 1227 12873 1261
rect 12931 1227 12965 1261
rect 13023 1227 13057 1261
rect 13115 1227 13149 1261
rect 13207 1227 13241 1261
rect 13299 1227 13333 1261
rect 13391 1227 13425 1261
rect 13483 1227 13517 1261
rect 13575 1227 13609 1261
rect 13667 1227 13701 1261
rect 13759 1227 13793 1261
rect 13851 1227 13885 1261
rect 13943 1227 13977 1261
rect 14035 1227 14069 1261
rect 14127 1227 14161 1261
rect 14219 1227 14253 1261
rect 14311 1227 14345 1261
rect 14403 1227 14437 1261
rect 14495 1227 14529 1261
rect 14587 1227 14621 1261
rect 14679 1227 14713 1261
rect 14771 1227 14805 1261
rect 14863 1227 14897 1261
rect 14955 1227 14989 1261
rect 15047 1227 15081 1261
rect 15139 1227 15173 1261
rect 15231 1227 15265 1261
rect 15323 1227 15357 1261
rect 15415 1227 15449 1261
rect 15507 1227 15541 1261
rect 15599 1227 15633 1261
rect 15691 1227 15725 1261
rect 15783 1227 15817 1261
rect 15875 1227 15909 1261
rect 15967 1227 16001 1261
rect 16059 1227 16093 1261
rect 16151 1227 16185 1261
rect 16243 1227 16277 1261
rect 16335 1227 16369 1261
rect 16427 1227 16461 1261
rect 16519 1227 16553 1261
rect 29 539 63 573
rect 121 539 155 573
rect 213 539 247 573
rect 305 539 339 573
rect 397 539 431 573
rect 489 539 523 573
rect 581 539 615 573
rect 673 539 707 573
rect 765 539 799 573
rect 857 539 891 573
rect 949 539 983 573
rect 1041 539 1075 573
rect 1133 539 1167 573
rect 1225 539 1259 573
rect 1317 539 1351 573
rect 1409 539 1443 573
rect 1501 539 1535 573
rect 1593 539 1627 573
rect 1685 539 1719 573
rect 1777 539 1811 573
rect 1869 539 1903 573
rect 1961 539 1995 573
rect 2053 539 2087 573
rect 2145 539 2179 573
rect 2237 539 2271 573
rect 2329 539 2363 573
rect 2421 539 2455 573
rect 2513 539 2547 573
rect 2605 539 2639 573
rect 2697 539 2731 573
rect 2789 539 2823 573
rect 2881 539 2915 573
rect 2973 539 3007 573
rect 3065 539 3099 573
rect 3157 539 3191 573
rect 3249 539 3283 573
rect 3341 539 3375 573
rect 3433 539 3467 573
rect 3525 539 3559 573
rect 3617 539 3651 573
rect 3709 539 3743 573
rect 3801 539 3835 573
rect 3893 539 3927 573
rect 3985 539 4019 573
rect 4077 539 4111 573
rect 4169 539 4203 573
rect 4261 539 4295 573
rect 4353 539 4387 573
rect 4445 539 4479 573
rect 4537 539 4571 573
rect 4629 539 4663 573
rect 4721 539 4755 573
rect 4813 539 4847 573
rect 4905 539 4939 573
rect 4997 539 5031 573
rect 5089 539 5123 573
rect 5181 539 5215 573
rect 5273 539 5307 573
rect 5365 539 5399 573
rect 5457 539 5491 573
rect 5549 539 5583 573
rect 5641 539 5675 573
rect 5733 539 5767 573
rect 5825 539 5859 573
rect 5917 539 5951 573
rect 6009 539 6043 573
rect 6101 539 6135 573
rect 6193 539 6227 573
rect 6285 539 6319 573
rect 6377 539 6411 573
rect 6469 539 6503 573
rect 6561 539 6595 573
rect 6653 539 6687 573
rect 6745 539 6779 573
rect 6837 539 6871 573
rect 6929 539 6963 573
rect 7021 539 7055 573
rect 7113 539 7147 573
rect 7205 539 7239 573
rect 7297 539 7331 573
rect 7389 539 7423 573
rect 7481 539 7515 573
rect 7573 539 7607 573
rect 7665 539 7699 573
rect 7757 539 7791 573
rect 7849 539 7883 573
rect 7941 539 7975 573
rect 8033 539 8067 573
rect 8125 539 8159 573
rect 8217 539 8251 573
rect 8309 539 8343 573
rect 8401 539 8435 573
rect 8493 539 8527 573
rect 8585 539 8619 573
rect 8677 539 8711 573
rect 8769 539 8803 573
rect 8861 539 8895 573
rect 8953 539 8987 573
rect 9045 539 9079 573
rect 9137 539 9171 573
rect 9229 539 9263 573
rect 9321 539 9355 573
rect 9413 539 9447 573
rect 9505 539 9539 573
rect 9597 539 9631 573
rect 9689 539 9723 573
rect 9781 539 9815 573
rect 9873 539 9907 573
rect 9965 539 9999 573
rect 10057 539 10091 573
rect 10149 539 10183 573
rect 10241 539 10275 573
rect 10333 539 10367 573
rect 10425 539 10459 573
rect 10517 539 10551 573
rect 10609 539 10643 573
rect 10701 539 10735 573
rect 10793 539 10827 573
rect 10885 539 10919 573
rect 10977 539 11011 573
rect 11069 539 11103 573
rect 11161 539 11195 573
rect 11253 539 11287 573
rect 11345 539 11379 573
rect 11437 539 11471 573
rect 11529 539 11563 573
rect 11621 539 11655 573
rect 11713 539 11747 573
rect 11805 539 11839 573
rect 11897 539 11931 573
rect 11989 539 12023 573
rect 12081 539 12115 573
rect 12173 539 12207 573
rect 12265 539 12299 573
rect 12357 539 12391 573
rect 12449 539 12483 573
rect 12541 539 12575 573
rect 12633 539 12667 573
rect 12725 539 12759 573
rect 12817 539 12851 573
rect 12909 539 12943 573
rect 13001 539 13035 573
rect 13093 539 13127 573
rect 13185 539 13219 573
rect 13277 539 13311 573
rect 13369 539 13403 573
rect 13461 539 13495 573
rect 13553 539 13587 573
rect 13645 539 13679 573
rect 13737 539 13771 573
rect 13829 539 13863 573
rect 13921 539 13955 573
rect 14013 539 14047 573
rect 14105 539 14139 573
rect 14197 539 14231 573
rect 14289 539 14323 573
rect 14381 539 14415 573
rect 14473 539 14507 573
rect 14565 539 14599 573
rect 14657 539 14691 573
rect 14749 539 14783 573
rect 14841 539 14875 573
rect 14933 539 14967 573
rect 15025 539 15059 573
rect 15117 539 15151 573
rect 15209 539 15243 573
rect 15301 539 15335 573
rect 15393 539 15427 573
rect 15485 539 15519 573
rect 15577 539 15611 573
rect 15669 539 15703 573
rect 15761 539 15795 573
rect 15853 539 15887 573
rect 15945 539 15979 573
rect 16037 539 16071 573
rect 16129 539 16163 573
rect 16221 539 16255 573
rect 16313 539 16347 573
rect 16405 539 16439 573
rect 16497 539 16531 573
rect 16589 539 16623 573
rect 16681 539 16715 573
rect 29 -150 63 -116
rect 121 -150 155 -116
rect 213 -150 247 -116
rect 305 -150 339 -116
rect 397 -150 431 -116
rect 489 -150 523 -116
rect 581 -150 615 -116
rect 673 -150 707 -116
rect 765 -150 799 -116
rect 857 -150 891 -116
rect 949 -150 983 -116
rect 1041 -150 1075 -116
rect 1133 -150 1167 -116
rect 1225 -150 1259 -116
rect 1317 -150 1351 -116
rect 1409 -150 1443 -116
rect 1501 -150 1535 -116
rect 1593 -150 1627 -116
rect 1685 -150 1719 -116
rect 1777 -150 1811 -116
rect 1869 -150 1903 -116
rect 1961 -150 1995 -116
rect 2053 -150 2087 -116
rect 2145 -150 2179 -116
rect 2237 -150 2271 -116
rect 2329 -150 2363 -116
rect 2421 -150 2455 -116
rect 2513 -150 2547 -116
rect 2605 -150 2639 -116
rect 2697 -150 2731 -116
rect 2789 -150 2823 -116
rect 2881 -150 2915 -116
rect 2973 -150 3007 -116
rect 3065 -150 3099 -116
rect 3157 -150 3191 -116
rect 3249 -150 3283 -116
rect 3341 -150 3375 -116
rect 3433 -150 3467 -116
rect 3525 -150 3559 -116
rect 3617 -150 3651 -116
rect 3709 -150 3743 -116
rect 3801 -150 3835 -116
rect 3893 -150 3927 -116
rect 3985 -150 4019 -116
rect 4077 -150 4111 -116
rect 4169 -150 4203 -116
rect 4261 -150 4295 -116
rect 4353 -150 4387 -116
rect 4445 -150 4479 -116
rect 4537 -150 4571 -116
rect 4629 -150 4663 -116
rect 4721 -150 4755 -116
rect 4813 -150 4847 -116
rect 4905 -150 4939 -116
rect 4997 -150 5031 -116
rect 5089 -150 5123 -116
rect 5181 -150 5215 -116
rect 5273 -150 5307 -116
rect 5365 -150 5399 -116
rect 5457 -150 5491 -116
rect 5549 -150 5583 -116
rect 5641 -150 5675 -116
rect 5733 -150 5767 -116
rect 5825 -150 5859 -116
rect 5917 -150 5951 -116
rect 6009 -150 6043 -116
rect 6101 -150 6135 -116
rect 6193 -150 6227 -116
rect 6285 -150 6319 -116
rect 6377 -150 6411 -116
rect 6469 -150 6503 -116
rect 6561 -150 6595 -116
rect 6653 -150 6687 -116
rect 6745 -150 6779 -116
rect 6837 -150 6871 -116
rect 6929 -150 6963 -116
rect 7021 -150 7055 -116
rect 7113 -150 7147 -116
rect 7205 -150 7239 -116
rect 7297 -150 7331 -116
rect 7389 -150 7423 -116
rect 7481 -150 7515 -116
rect 7573 -150 7607 -116
rect 7665 -150 7699 -116
rect 7757 -150 7791 -116
rect 7849 -150 7883 -116
rect 7941 -150 7975 -116
rect 8033 -150 8067 -116
rect 8125 -150 8159 -116
rect 8217 -150 8251 -116
rect 8309 -150 8343 -116
rect 8401 -150 8435 -116
rect 8493 -150 8527 -116
rect 8585 -150 8619 -116
rect 8677 -150 8711 -116
rect 8769 -150 8803 -116
rect 8861 -150 8895 -116
rect 8953 -150 8987 -116
rect 9045 -150 9079 -116
rect 9137 -150 9171 -116
rect 9229 -150 9263 -116
rect 9321 -150 9355 -116
rect 9413 -150 9447 -116
rect 9505 -150 9539 -116
rect 9597 -150 9631 -116
rect 9689 -150 9723 -116
rect 9781 -150 9815 -116
rect 9873 -150 9907 -116
rect 9965 -150 9999 -116
rect 10057 -150 10091 -116
rect 10149 -150 10183 -116
rect 10241 -150 10275 -116
rect 10333 -150 10367 -116
rect 10425 -150 10459 -116
rect 10517 -150 10551 -116
rect 10609 -150 10643 -116
rect 10701 -150 10735 -116
rect 10793 -150 10827 -116
rect 10885 -150 10919 -116
rect 10977 -150 11011 -116
rect 11069 -150 11103 -116
rect 11161 -150 11195 -116
rect 11253 -150 11287 -116
rect 11345 -150 11379 -116
rect 11437 -150 11471 -116
rect 11529 -150 11563 -116
rect 11621 -150 11655 -116
rect 11713 -150 11747 -116
rect 11805 -150 11839 -116
rect 11897 -150 11931 -116
rect 11989 -150 12023 -116
rect 12081 -150 12115 -116
rect 12173 -150 12207 -116
rect 12265 -150 12299 -116
rect 12357 -150 12391 -116
rect 12449 -150 12483 -116
rect 12541 -150 12575 -116
rect 12633 -150 12667 -116
rect 12725 -150 12759 -116
rect 12817 -150 12851 -116
rect 12909 -150 12943 -116
rect 13001 -150 13035 -116
rect 13093 -150 13127 -116
rect 13185 -150 13219 -116
rect 13277 -150 13311 -116
rect 13369 -150 13403 -116
rect 13461 -150 13495 -116
rect 13553 -150 13587 -116
rect 13645 -150 13679 -116
rect 13737 -150 13771 -116
rect 13829 -150 13863 -116
rect 13921 -150 13955 -116
rect 14013 -150 14047 -116
rect 14105 -150 14139 -116
rect 14197 -150 14231 -116
rect 14289 -150 14323 -116
rect 14381 -150 14415 -116
rect 14473 -150 14507 -116
rect 14565 -150 14599 -116
rect 14657 -150 14691 -116
rect 14749 -150 14783 -116
rect 14841 -150 14875 -116
rect 14933 -150 14967 -116
rect 15025 -150 15059 -116
rect 15117 -150 15151 -116
rect 15209 -150 15243 -116
rect 15301 -150 15335 -116
rect 15393 -150 15427 -116
rect 15485 -150 15519 -116
rect 15577 -150 15611 -116
rect 15669 -150 15703 -116
rect 15761 -150 15795 -116
rect 15853 -150 15887 -116
rect 15945 -150 15979 -116
rect 16037 -150 16071 -116
rect 16129 -150 16163 -116
rect 16221 -150 16255 -116
rect 16313 -150 16347 -116
rect 16405 -150 16439 -116
rect 16497 -150 16531 -116
rect 16589 -150 16623 -116
rect 16681 -150 16715 -116
<< nsubdiffcont >>
rect 31 2961 65 2995
rect 123 2961 157 2995
rect 215 2961 249 2995
rect 307 2961 341 2995
rect 399 2961 433 2995
rect 491 2961 525 2995
rect 583 2961 617 2995
rect 675 2961 709 2995
rect 767 2961 801 2995
rect 859 2961 893 2995
rect 951 2961 985 2995
rect 1043 2961 1077 2995
rect 1135 2961 1169 2995
rect 1227 2961 1261 2995
rect 1319 2961 1353 2995
rect 1411 2961 1445 2995
rect 1503 2961 1537 2995
rect 1595 2961 1629 2995
rect 1687 2961 1721 2995
rect 1779 2961 1813 2995
rect 1871 2961 1905 2995
rect 1963 2961 1997 2995
rect 2055 2961 2089 2995
rect 2147 2961 2181 2995
rect 2239 2961 2273 2995
rect 2331 2961 2365 2995
rect 2423 2961 2457 2995
rect 2515 2961 2549 2995
rect 2607 2961 2641 2995
rect 2699 2961 2733 2995
rect 2791 2961 2825 2995
rect 4415 2961 4449 2995
rect 4507 2961 4541 2995
rect 4599 2961 4633 2995
rect 4691 2961 4725 2995
rect 4783 2961 4817 2995
rect 4875 2961 4909 2995
rect 4967 2961 5001 2995
rect 5059 2961 5093 2995
rect 5151 2961 5185 2995
rect 5243 2961 5277 2995
rect 5335 2961 5369 2995
rect 5427 2961 5461 2995
rect 5519 2961 5553 2995
rect 5611 2961 5645 2995
rect 5703 2961 5737 2995
rect 5795 2961 5829 2995
rect 5887 2961 5921 2995
rect 5979 2961 6013 2995
rect 6071 2961 6105 2995
rect 6163 2961 6197 2995
rect 6255 2961 6289 2995
rect 6347 2961 6381 2995
rect 6439 2961 6473 2995
rect 6531 2961 6565 2995
rect 6623 2961 6657 2995
rect 6715 2961 6749 2995
rect 6807 2961 6841 2995
rect 6899 2961 6933 2995
rect 6991 2961 7025 2995
rect 7083 2961 7117 2995
rect 7175 2961 7209 2995
rect 29 1819 63 1853
rect 121 1819 155 1853
rect 213 1819 247 1853
rect 305 1819 339 1853
rect 397 1819 431 1853
rect 489 1819 523 1853
rect 581 1819 615 1853
rect 673 1819 707 1853
rect 765 1819 799 1853
rect 857 1819 891 1853
rect 949 1819 983 1853
rect 1041 1819 1075 1853
rect 1133 1819 1167 1853
rect 1225 1819 1259 1853
rect 1317 1819 1351 1853
rect 1409 1819 1443 1853
rect 1501 1819 1535 1853
rect 1593 1819 1627 1853
rect 1685 1819 1719 1853
rect 1777 1819 1811 1853
rect 1869 1819 1903 1853
rect 1961 1819 1995 1853
rect 2053 1819 2087 1853
rect 2145 1819 2179 1853
rect 2237 1819 2271 1853
rect 2329 1819 2363 1853
rect 2421 1819 2455 1853
rect 2513 1819 2547 1853
rect 2605 1819 2639 1853
rect 2697 1819 2731 1853
rect 2789 1819 2823 1853
rect 2881 1819 2915 1853
rect 2973 1819 3007 1853
rect 3065 1819 3099 1853
rect 3157 1819 3191 1853
rect 3249 1819 3283 1853
rect 3341 1819 3375 1853
rect 3433 1819 3467 1853
rect 3525 1819 3559 1853
rect 3617 1819 3651 1853
rect 3709 1819 3743 1853
rect 3801 1819 3835 1853
rect 3893 1819 3927 1853
rect 3985 1819 4019 1853
rect 4077 1819 4111 1853
rect 4169 1819 4203 1853
rect 4261 1819 4295 1853
rect 4353 1819 4387 1853
rect 4445 1819 4479 1853
rect 4537 1819 4571 1853
rect 4629 1819 4663 1853
rect 4721 1819 4755 1853
rect 4813 1819 4847 1853
rect 4905 1819 4939 1853
rect 4997 1819 5031 1853
rect 5089 1819 5123 1853
rect 5181 1819 5215 1853
rect 5273 1819 5307 1853
rect 5365 1819 5399 1853
rect 5457 1819 5491 1853
rect 5549 1819 5583 1853
rect 5641 1819 5675 1853
rect 6245 1819 6279 1853
rect 6337 1819 6371 1853
rect 6429 1819 6463 1853
rect 6521 1819 6555 1853
rect 6613 1819 6647 1853
rect 6705 1819 6739 1853
rect 6797 1819 6831 1853
rect 6889 1819 6923 1853
rect 6981 1819 7015 1853
rect 7073 1819 7107 1853
rect 7165 1819 7199 1853
rect 7257 1819 7291 1853
rect 7349 1819 7383 1853
rect 7441 1819 7475 1853
rect 7533 1819 7567 1853
rect 7625 1819 7659 1853
rect 7717 1819 7751 1853
rect 7809 1819 7843 1853
rect 7901 1819 7935 1853
rect 7993 1819 8027 1853
rect 8085 1819 8119 1853
rect 8177 1819 8211 1853
rect 8269 1819 8303 1853
rect 8361 1819 8395 1853
rect 8453 1819 8487 1853
rect 8545 1819 8579 1853
rect 8637 1819 8671 1853
rect 8729 1819 8763 1853
rect 8821 1819 8855 1853
rect 8913 1819 8947 1853
rect 9005 1819 9039 1853
rect 9097 1819 9131 1853
rect 9189 1819 9223 1853
rect 9281 1819 9315 1853
rect 9373 1819 9407 1853
rect 9465 1819 9499 1853
rect 9557 1819 9591 1853
rect 9649 1819 9683 1853
rect 9741 1819 9775 1853
rect 9833 1819 9867 1853
rect 9925 1819 9959 1853
rect 10017 1819 10051 1853
rect 10109 1819 10143 1853
rect 10201 1819 10235 1853
rect 10293 1819 10327 1853
rect 10385 1819 10419 1853
rect 10477 1819 10511 1853
rect 10569 1819 10603 1853
rect 10661 1819 10695 1853
rect 10753 1819 10787 1853
rect 10845 1819 10879 1853
rect 10937 1819 10971 1853
rect 11029 1819 11063 1853
rect 11121 1819 11155 1853
rect 11213 1819 11247 1853
rect 11305 1819 11339 1853
rect 11397 1819 11431 1853
rect 11489 1819 11523 1853
rect 11581 1819 11615 1853
rect 11673 1819 11707 1853
rect 11765 1819 11799 1853
rect 11857 1819 11891 1853
rect 12011 1819 12045 1853
rect 12103 1819 12137 1853
rect 12195 1819 12229 1853
rect 12287 1819 12321 1853
rect 12379 1819 12413 1853
rect 12471 1819 12505 1853
rect 12563 1819 12597 1853
rect 12655 1819 12689 1853
rect 12747 1819 12781 1853
rect 12839 1819 12873 1853
rect 12931 1819 12965 1853
rect 13023 1819 13057 1853
rect 13115 1819 13149 1853
rect 13207 1819 13241 1853
rect 13299 1819 13333 1853
rect 13391 1819 13425 1853
rect 13483 1819 13517 1853
rect 13575 1819 13609 1853
rect 13667 1819 13701 1853
rect 13759 1819 13793 1853
rect 13851 1819 13885 1853
rect 13943 1819 13977 1853
rect 14035 1819 14069 1853
rect 14127 1819 14161 1853
rect 14219 1819 14253 1853
rect 14311 1819 14345 1853
rect 14403 1819 14437 1853
rect 14495 1819 14529 1853
rect 14587 1819 14621 1853
rect 14679 1819 14713 1853
rect 14771 1819 14805 1853
rect 14863 1819 14897 1853
rect 14955 1819 14989 1853
rect 15047 1819 15081 1853
rect 15139 1819 15173 1853
rect 15231 1819 15265 1853
rect 15323 1819 15357 1853
rect 15415 1819 15449 1853
rect 15507 1819 15541 1853
rect 15599 1819 15633 1853
rect 15691 1819 15725 1853
rect 15783 1819 15817 1853
rect 15875 1819 15909 1853
rect 15967 1819 16001 1853
rect 16059 1819 16093 1853
rect 16151 1819 16185 1853
rect 16243 1819 16277 1853
rect 16335 1819 16369 1853
rect 16427 1819 16461 1853
rect 16519 1819 16553 1853
rect 29 1131 63 1165
rect 121 1131 155 1165
rect 213 1131 247 1165
rect 305 1131 339 1165
rect 397 1131 431 1165
rect 489 1131 523 1165
rect 581 1131 615 1165
rect 673 1131 707 1165
rect 765 1131 799 1165
rect 857 1131 891 1165
rect 949 1131 983 1165
rect 1041 1131 1075 1165
rect 1133 1131 1167 1165
rect 1225 1131 1259 1165
rect 1317 1131 1351 1165
rect 1409 1131 1443 1165
rect 1501 1131 1535 1165
rect 1593 1131 1627 1165
rect 1685 1131 1719 1165
rect 1777 1131 1811 1165
rect 2053 1131 2087 1165
rect 2145 1131 2179 1165
rect 2237 1131 2271 1165
rect 2329 1131 2363 1165
rect 2421 1131 2455 1165
rect 2513 1131 2547 1165
rect 2605 1131 2639 1165
rect 2697 1131 2731 1165
rect 2789 1131 2823 1165
rect 2881 1131 2915 1165
rect 2973 1131 3007 1165
rect 3065 1131 3099 1165
rect 3157 1131 3191 1165
rect 3249 1131 3283 1165
rect 3341 1131 3375 1165
rect 3433 1131 3467 1165
rect 3525 1131 3559 1165
rect 3617 1131 3651 1165
rect 3709 1131 3743 1165
rect 3801 1131 3835 1165
rect 3893 1131 3927 1165
rect 3985 1131 4019 1165
rect 4077 1131 4111 1165
rect 4169 1131 4203 1165
rect 4445 1131 4479 1165
rect 4537 1131 4571 1165
rect 4629 1131 4663 1165
rect 4721 1131 4755 1165
rect 4813 1131 4847 1165
rect 4905 1131 4939 1165
rect 4997 1131 5031 1165
rect 5089 1131 5123 1165
rect 5181 1131 5215 1165
rect 5273 1131 5307 1165
rect 5365 1131 5399 1165
rect 5457 1131 5491 1165
rect 5549 1131 5583 1165
rect 5641 1131 5675 1165
rect 5733 1131 5767 1165
rect 5825 1131 5859 1165
rect 5917 1131 5951 1165
rect 6009 1131 6043 1165
rect 6101 1131 6135 1165
rect 6193 1131 6227 1165
rect 6285 1131 6319 1165
rect 6377 1131 6411 1165
rect 6469 1131 6503 1165
rect 6561 1131 6595 1165
rect 6837 1131 6871 1165
rect 6929 1131 6963 1165
rect 7021 1131 7055 1165
rect 7113 1131 7147 1165
rect 7205 1131 7239 1165
rect 7297 1131 7331 1165
rect 7389 1131 7423 1165
rect 7481 1131 7515 1165
rect 7573 1131 7607 1165
rect 7665 1131 7699 1165
rect 7757 1131 7791 1165
rect 7849 1131 7883 1165
rect 7941 1131 7975 1165
rect 8033 1131 8067 1165
rect 8125 1131 8159 1165
rect 8217 1131 8251 1165
rect 8309 1131 8343 1165
rect 8401 1131 8435 1165
rect 8493 1131 8527 1165
rect 8585 1131 8619 1165
rect 8677 1131 8711 1165
rect 8769 1131 8803 1165
rect 8861 1131 8895 1165
rect 8953 1131 8987 1165
rect 9229 1131 9263 1165
rect 9321 1131 9355 1165
rect 9413 1131 9447 1165
rect 9505 1131 9539 1165
rect 9597 1131 9631 1165
rect 9689 1131 9723 1165
rect 9781 1131 9815 1165
rect 9873 1131 9907 1165
rect 9965 1131 9999 1165
rect 10057 1131 10091 1165
rect 10149 1131 10183 1165
rect 10241 1131 10275 1165
rect 10333 1131 10367 1165
rect 10425 1131 10459 1165
rect 10517 1131 10551 1165
rect 10609 1131 10643 1165
rect 10701 1131 10735 1165
rect 10793 1131 10827 1165
rect 10885 1131 10919 1165
rect 10977 1131 11011 1165
rect 11069 1131 11103 1165
rect 11161 1131 11195 1165
rect 11253 1131 11287 1165
rect 11345 1131 11379 1165
rect 11621 1131 11655 1165
rect 11713 1131 11747 1165
rect 11805 1131 11839 1165
rect 11897 1131 11931 1165
rect 11989 1131 12023 1165
rect 12081 1131 12115 1165
rect 12173 1131 12207 1165
rect 12265 1131 12299 1165
rect 12357 1131 12391 1165
rect 12449 1131 12483 1165
rect 12541 1131 12575 1165
rect 12633 1131 12667 1165
rect 12725 1131 12759 1165
rect 12817 1131 12851 1165
rect 12909 1131 12943 1165
rect 13001 1131 13035 1165
rect 13093 1131 13127 1165
rect 13185 1131 13219 1165
rect 13277 1131 13311 1165
rect 13369 1131 13403 1165
rect 13461 1131 13495 1165
rect 13553 1131 13587 1165
rect 13645 1131 13679 1165
rect 13737 1131 13771 1165
rect 14013 1131 14047 1165
rect 14105 1131 14139 1165
rect 14197 1131 14231 1165
rect 14289 1131 14323 1165
rect 14381 1131 14415 1165
rect 14473 1131 14507 1165
rect 14565 1131 14599 1165
rect 14657 1131 14691 1165
rect 14749 1131 14783 1165
rect 14841 1131 14875 1165
rect 14933 1131 14967 1165
rect 15025 1131 15059 1165
rect 15117 1131 15151 1165
rect 15209 1131 15243 1165
rect 15301 1131 15335 1165
rect 15393 1131 15427 1165
rect 15485 1131 15519 1165
rect 15577 1131 15611 1165
rect 15669 1131 15703 1165
rect 15761 1131 15795 1165
rect 15853 1131 15887 1165
rect 15945 1131 15979 1165
rect 16037 1131 16071 1165
rect 16129 1131 16163 1165
rect 16405 1131 16439 1165
rect 16497 1131 16531 1165
rect 16589 1131 16623 1165
rect 16681 1131 16715 1165
rect 29 442 63 476
rect 121 442 155 476
rect 213 442 247 476
rect 305 442 339 476
rect 394 442 428 476
rect 496 442 530 476
rect 581 442 615 476
rect 673 442 707 476
rect 765 442 799 476
rect 857 442 891 476
rect 949 442 983 476
rect 1041 442 1075 476
rect 1133 442 1167 476
rect 1225 442 1259 476
rect 1317 442 1351 476
rect 1409 442 1443 476
rect 1501 442 1535 476
rect 1777 442 1811 476
rect 1869 442 1903 476
rect 1961 442 1995 476
rect 2053 442 2087 476
rect 2145 442 2179 476
rect 2237 442 2271 476
rect 2329 442 2363 476
rect 2421 442 2455 476
rect 2513 442 2547 476
rect 2605 442 2639 476
rect 2697 442 2731 476
rect 2791 442 2825 476
rect 2882 442 2916 476
rect 2973 442 3007 476
rect 3065 442 3099 476
rect 3157 442 3191 476
rect 3249 442 3283 476
rect 3341 442 3375 476
rect 3433 442 3467 476
rect 3525 442 3559 476
rect 3617 442 3651 476
rect 3709 442 3743 476
rect 3801 442 3835 476
rect 3893 442 3927 476
rect 4169 442 4203 476
rect 4261 442 4295 476
rect 4353 442 4387 476
rect 4445 442 4479 476
rect 4537 442 4571 476
rect 4629 442 4663 476
rect 4721 442 4755 476
rect 4813 442 4847 476
rect 4905 442 4939 476
rect 4997 442 5031 476
rect 5089 442 5123 476
rect 5179 442 5213 476
rect 5273 442 5307 476
rect 5365 442 5399 476
rect 5457 442 5491 476
rect 5549 442 5583 476
rect 5641 442 5675 476
rect 5733 442 5767 476
rect 5825 442 5859 476
rect 5917 442 5951 476
rect 6009 442 6043 476
rect 6101 442 6135 476
rect 6193 442 6227 476
rect 6285 442 6319 476
rect 6561 442 6595 476
rect 6653 442 6687 476
rect 6745 442 6779 476
rect 6837 442 6871 476
rect 6929 442 6963 476
rect 7021 442 7055 476
rect 7113 442 7147 476
rect 7205 442 7239 476
rect 7297 442 7331 476
rect 7389 442 7423 476
rect 7481 442 7515 476
rect 7574 442 7608 476
rect 7665 442 7699 476
rect 7757 442 7791 476
rect 7849 442 7883 476
rect 7941 442 7975 476
rect 8033 442 8067 476
rect 8125 442 8159 476
rect 8217 442 8251 476
rect 8309 442 8343 476
rect 8401 442 8435 476
rect 8493 442 8527 476
rect 8585 442 8619 476
rect 8677 442 8711 476
rect 8953 442 8987 476
rect 9045 442 9079 476
rect 9137 442 9171 476
rect 9229 442 9263 476
rect 9321 442 9355 476
rect 9413 442 9447 476
rect 9505 442 9539 476
rect 9597 442 9631 476
rect 9689 442 9723 476
rect 9781 442 9815 476
rect 9873 442 9907 476
rect 9963 442 9997 476
rect 10058 442 10092 476
rect 10149 442 10183 476
rect 10241 442 10275 476
rect 10333 442 10367 476
rect 10425 442 10459 476
rect 10517 442 10551 476
rect 10609 442 10643 476
rect 10701 442 10735 476
rect 10793 442 10827 476
rect 10885 442 10919 476
rect 10977 442 11011 476
rect 11069 442 11103 476
rect 11345 442 11379 476
rect 11437 442 11471 476
rect 11529 442 11563 476
rect 11621 442 11655 476
rect 11713 442 11747 476
rect 11805 442 11839 476
rect 11897 442 11931 476
rect 11989 442 12023 476
rect 12081 442 12115 476
rect 12173 442 12207 476
rect 12265 442 12299 476
rect 12357 442 12391 476
rect 12448 442 12482 476
rect 12541 442 12575 476
rect 12633 442 12667 476
rect 12725 442 12759 476
rect 12817 442 12851 476
rect 12909 442 12943 476
rect 13001 442 13035 476
rect 13093 442 13127 476
rect 13185 442 13219 476
rect 13277 442 13311 476
rect 13369 442 13403 476
rect 13461 442 13495 476
rect 13737 442 13771 476
rect 13829 442 13863 476
rect 13921 442 13955 476
rect 14013 442 14047 476
rect 14105 442 14139 476
rect 14197 442 14231 476
rect 14289 442 14323 476
rect 14381 442 14415 476
rect 14473 442 14507 476
rect 14565 442 14599 476
rect 14657 442 14691 476
rect 14748 442 14782 476
rect 14842 442 14876 476
rect 14933 442 14967 476
rect 15025 442 15059 476
rect 15117 442 15151 476
rect 15209 442 15243 476
rect 15301 442 15335 476
rect 15393 442 15427 476
rect 15485 442 15519 476
rect 15577 442 15611 476
rect 15669 442 15703 476
rect 15761 442 15795 476
rect 15853 442 15887 476
rect 16129 442 16163 476
rect 16221 442 16255 476
rect 16313 442 16347 476
rect 16405 442 16439 476
rect 16497 442 16531 476
rect 16589 442 16623 476
rect 16681 442 16715 476
<< poly >>
rect 81 2907 111 2933
rect 169 2907 199 2933
rect 357 2907 387 2933
rect 441 2907 471 2933
rect 525 2907 555 2933
rect 609 2907 639 2933
rect 693 2907 723 2933
rect 909 2907 939 2933
rect 993 2907 1023 2933
rect 1077 2907 1107 2933
rect 1161 2907 1191 2933
rect 1245 2907 1275 2933
rect 1329 2907 1359 2933
rect 1413 2907 1443 2933
rect 1497 2907 1527 2933
rect 1581 2907 1611 2933
rect 1665 2907 1695 2933
rect 1749 2907 1779 2933
rect 1833 2907 1863 2933
rect 1917 2907 1947 2933
rect 2001 2907 2031 2933
rect 2085 2907 2115 2933
rect 2169 2907 2199 2933
rect 2253 2907 2283 2933
rect 2337 2907 2367 2933
rect 2421 2907 2451 2933
rect 2505 2907 2535 2933
rect 2589 2907 2619 2933
rect 2673 2907 2703 2933
rect 4465 2907 4495 2933
rect 4553 2907 4583 2933
rect 4741 2907 4771 2933
rect 4825 2907 4855 2933
rect 4909 2907 4939 2933
rect 4993 2907 5023 2933
rect 5077 2907 5107 2933
rect 5293 2907 5323 2933
rect 5377 2907 5407 2933
rect 5461 2907 5491 2933
rect 5545 2907 5575 2933
rect 5629 2907 5659 2933
rect 5713 2907 5743 2933
rect 5797 2907 5827 2933
rect 5881 2907 5911 2933
rect 5965 2907 5995 2933
rect 6049 2907 6079 2933
rect 6133 2907 6163 2933
rect 6217 2907 6247 2933
rect 6301 2907 6331 2933
rect 6385 2907 6415 2933
rect 6469 2907 6499 2933
rect 6553 2907 6583 2933
rect 6637 2907 6667 2933
rect 6721 2907 6751 2933
rect 6805 2907 6835 2933
rect 6889 2907 6919 2933
rect 6973 2907 7003 2933
rect 7057 2907 7087 2933
rect 81 2734 111 2749
rect 75 2710 111 2734
rect 75 2675 105 2710
rect 169 2688 199 2749
rect 4465 2734 4495 2749
rect 4459 2710 4495 2734
rect 29 2659 105 2675
rect 29 2625 39 2659
rect 73 2625 105 2659
rect 29 2609 105 2625
rect 147 2672 201 2688
rect 147 2638 157 2672
rect 191 2638 201 2672
rect 357 2671 387 2707
rect 147 2622 201 2638
rect 306 2659 387 2671
rect 441 2669 471 2707
rect 525 2669 555 2707
rect 609 2669 639 2707
rect 693 2669 723 2707
rect 306 2625 322 2659
rect 356 2625 387 2659
rect 75 2600 105 2609
rect 75 2576 111 2600
rect 81 2561 111 2576
rect 169 2561 199 2622
rect 306 2613 387 2625
rect 440 2659 723 2669
rect 440 2625 456 2659
rect 490 2625 723 2659
rect 440 2615 723 2625
rect 357 2587 387 2613
rect 441 2587 471 2615
rect 525 2587 555 2615
rect 609 2587 639 2615
rect 693 2587 723 2615
rect 909 2669 939 2707
rect 993 2669 1023 2707
rect 1077 2669 1107 2707
rect 1161 2669 1191 2707
rect 1245 2669 1275 2707
rect 1329 2669 1359 2707
rect 909 2659 1359 2669
rect 909 2625 933 2659
rect 967 2625 1001 2659
rect 1035 2625 1069 2659
rect 1103 2625 1137 2659
rect 1171 2625 1205 2659
rect 1239 2625 1273 2659
rect 1307 2625 1359 2659
rect 909 2615 1359 2625
rect 909 2587 939 2615
rect 993 2587 1023 2615
rect 1077 2587 1107 2615
rect 1161 2587 1191 2615
rect 1245 2587 1275 2615
rect 1329 2587 1359 2615
rect 1413 2669 1443 2707
rect 1497 2669 1527 2707
rect 1581 2669 1611 2707
rect 1665 2669 1695 2707
rect 1749 2669 1779 2707
rect 1833 2669 1863 2707
rect 1917 2669 1947 2707
rect 2001 2669 2031 2707
rect 2085 2669 2115 2707
rect 2169 2669 2199 2707
rect 2253 2669 2283 2707
rect 2337 2669 2367 2707
rect 2421 2669 2451 2707
rect 2505 2669 2535 2707
rect 2589 2669 2619 2707
rect 2673 2669 2703 2707
rect 4459 2675 4489 2710
rect 4553 2688 4583 2749
rect 1413 2659 2707 2669
rect 1413 2625 1433 2659
rect 1467 2625 1501 2659
rect 1535 2625 1569 2659
rect 1603 2625 1637 2659
rect 1671 2625 1705 2659
rect 1739 2625 1773 2659
rect 1807 2625 1841 2659
rect 1875 2625 1909 2659
rect 1943 2625 1977 2659
rect 2011 2625 2045 2659
rect 2079 2625 2113 2659
rect 2147 2625 2181 2659
rect 2215 2625 2249 2659
rect 2283 2625 2317 2659
rect 2351 2625 2385 2659
rect 2419 2625 2453 2659
rect 2487 2625 2521 2659
rect 2555 2625 2589 2659
rect 2623 2625 2657 2659
rect 2691 2625 2707 2659
rect 1413 2615 2707 2625
rect 4413 2659 4489 2675
rect 4413 2625 4423 2659
rect 4457 2625 4489 2659
rect 1413 2587 1443 2615
rect 1497 2587 1527 2615
rect 1581 2587 1611 2615
rect 1665 2587 1695 2615
rect 1749 2587 1779 2615
rect 1833 2587 1863 2615
rect 1917 2587 1947 2615
rect 2001 2587 2031 2615
rect 2085 2587 2115 2615
rect 2169 2587 2199 2615
rect 2253 2587 2283 2615
rect 2337 2587 2367 2615
rect 2421 2587 2451 2615
rect 2505 2587 2535 2615
rect 2589 2587 2619 2615
rect 2673 2587 2703 2615
rect 4413 2609 4489 2625
rect 4531 2672 4585 2688
rect 4531 2638 4541 2672
rect 4575 2638 4585 2672
rect 4741 2671 4771 2707
rect 4531 2622 4585 2638
rect 4690 2659 4771 2671
rect 4825 2669 4855 2707
rect 4909 2669 4939 2707
rect 4993 2669 5023 2707
rect 5077 2669 5107 2707
rect 4690 2625 4706 2659
rect 4740 2625 4771 2659
rect 4459 2600 4489 2609
rect 4459 2576 4495 2600
rect 4465 2561 4495 2576
rect 4553 2561 4583 2622
rect 4690 2613 4771 2625
rect 4824 2659 5107 2669
rect 4824 2625 4840 2659
rect 4874 2625 5107 2659
rect 4824 2615 5107 2625
rect 4741 2587 4771 2613
rect 4825 2587 4855 2615
rect 4909 2587 4939 2615
rect 4993 2587 5023 2615
rect 5077 2587 5107 2615
rect 5293 2669 5323 2707
rect 5377 2669 5407 2707
rect 5461 2669 5491 2707
rect 5545 2669 5575 2707
rect 5629 2669 5659 2707
rect 5713 2669 5743 2707
rect 5293 2659 5743 2669
rect 5293 2625 5317 2659
rect 5351 2625 5385 2659
rect 5419 2625 5453 2659
rect 5487 2625 5521 2659
rect 5555 2625 5589 2659
rect 5623 2625 5657 2659
rect 5691 2625 5743 2659
rect 5293 2615 5743 2625
rect 5293 2587 5323 2615
rect 5377 2587 5407 2615
rect 5461 2587 5491 2615
rect 5545 2587 5575 2615
rect 5629 2587 5659 2615
rect 5713 2587 5743 2615
rect 5797 2669 5827 2707
rect 5881 2669 5911 2707
rect 5965 2669 5995 2707
rect 6049 2669 6079 2707
rect 6133 2669 6163 2707
rect 6217 2669 6247 2707
rect 6301 2669 6331 2707
rect 6385 2669 6415 2707
rect 6469 2669 6499 2707
rect 6553 2669 6583 2707
rect 6637 2669 6667 2707
rect 6721 2669 6751 2707
rect 6805 2669 6835 2707
rect 6889 2669 6919 2707
rect 6973 2669 7003 2707
rect 7057 2669 7087 2707
rect 5797 2659 7091 2669
rect 5797 2625 5817 2659
rect 5851 2625 5885 2659
rect 5919 2625 5953 2659
rect 5987 2625 6021 2659
rect 6055 2625 6089 2659
rect 6123 2625 6157 2659
rect 6191 2625 6225 2659
rect 6259 2625 6293 2659
rect 6327 2625 6361 2659
rect 6395 2625 6429 2659
rect 6463 2625 6497 2659
rect 6531 2625 6565 2659
rect 6599 2625 6633 2659
rect 6667 2625 6701 2659
rect 6735 2625 6769 2659
rect 6803 2625 6837 2659
rect 6871 2625 6905 2659
rect 6939 2625 6973 2659
rect 7007 2625 7041 2659
rect 7075 2625 7091 2659
rect 5797 2615 7091 2625
rect 5797 2587 5827 2615
rect 5881 2587 5911 2615
rect 5965 2587 5995 2615
rect 6049 2587 6079 2615
rect 6133 2587 6163 2615
rect 6217 2587 6247 2615
rect 6301 2587 6331 2615
rect 6385 2587 6415 2615
rect 6469 2587 6499 2615
rect 6553 2587 6583 2615
rect 6637 2587 6667 2615
rect 6721 2587 6751 2615
rect 6805 2587 6835 2615
rect 6889 2587 6919 2615
rect 6973 2587 7003 2615
rect 7057 2587 7087 2615
rect 81 2431 111 2457
rect 169 2431 199 2457
rect 357 2431 387 2457
rect 441 2431 471 2457
rect 525 2431 555 2457
rect 609 2431 639 2457
rect 693 2431 723 2457
rect 909 2431 939 2457
rect 993 2431 1023 2457
rect 1077 2431 1107 2457
rect 1161 2431 1191 2457
rect 1245 2431 1275 2457
rect 1329 2431 1359 2457
rect 1413 2431 1443 2457
rect 1497 2431 1527 2457
rect 1581 2431 1611 2457
rect 1665 2431 1695 2457
rect 1749 2431 1779 2457
rect 1833 2431 1863 2457
rect 1917 2431 1947 2457
rect 2001 2431 2031 2457
rect 2085 2431 2115 2457
rect 2169 2431 2199 2457
rect 2253 2431 2283 2457
rect 2337 2431 2367 2457
rect 2421 2431 2451 2457
rect 2505 2431 2535 2457
rect 2589 2431 2619 2457
rect 2673 2431 2703 2457
rect 4465 2431 4495 2457
rect 4553 2431 4583 2457
rect 4741 2431 4771 2457
rect 4825 2431 4855 2457
rect 4909 2431 4939 2457
rect 4993 2431 5023 2457
rect 5077 2431 5107 2457
rect 5293 2431 5323 2457
rect 5377 2431 5407 2457
rect 5461 2431 5491 2457
rect 5545 2431 5575 2457
rect 5629 2431 5659 2457
rect 5713 2431 5743 2457
rect 5797 2431 5827 2457
rect 5881 2431 5911 2457
rect 5965 2431 5995 2457
rect 6049 2431 6079 2457
rect 6133 2431 6163 2457
rect 6217 2431 6247 2457
rect 6301 2431 6331 2457
rect 6385 2431 6415 2457
rect 6469 2431 6499 2457
rect 6553 2431 6583 2457
rect 6637 2431 6667 2457
rect 6721 2431 6751 2457
rect 6805 2431 6835 2457
rect 6889 2431 6919 2457
rect 6973 2431 7003 2457
rect 7057 2431 7087 2457
rect 79 1765 109 1791
rect 2153 1765 2183 1791
rect 2471 1765 2501 1791
rect 4545 1765 4575 1791
rect 4863 1765 4893 1791
rect 6935 1765 6965 1791
rect 7255 1765 7285 1791
rect 9329 1765 9359 1791
rect 9647 1765 9677 1791
rect 11721 1765 11751 1791
rect 12039 1765 12069 1791
rect 14111 1765 14141 1791
rect 14431 1765 14461 1791
rect 16505 1765 16535 1791
rect 188 1726 218 1752
rect 291 1726 321 1752
rect 505 1726 535 1752
rect 577 1726 607 1752
rect 673 1726 703 1752
rect 1559 1726 1589 1752
rect 1655 1726 1685 1752
rect 1727 1726 1757 1752
rect 1941 1726 1971 1752
rect 2044 1726 2074 1752
rect 79 1533 109 1565
rect 188 1533 218 1642
rect 291 1627 321 1642
rect 291 1597 439 1627
rect 505 1610 535 1642
rect 76 1517 130 1533
rect 76 1483 86 1517
rect 120 1483 130 1517
rect 76 1467 130 1483
rect 172 1517 226 1533
rect 172 1483 182 1517
rect 216 1483 226 1517
rect 409 1497 439 1597
rect 481 1594 535 1610
rect 481 1560 491 1594
rect 525 1560 535 1594
rect 481 1544 535 1560
rect 172 1467 226 1483
rect 284 1481 367 1497
rect 79 1445 109 1467
rect 188 1399 218 1467
rect 284 1447 323 1481
rect 357 1447 367 1481
rect 284 1431 367 1447
rect 409 1481 463 1497
rect 577 1491 607 1642
rect 673 1610 703 1642
rect 649 1594 703 1610
rect 649 1560 659 1594
rect 693 1560 703 1594
rect 649 1544 703 1560
rect 409 1447 419 1481
rect 453 1447 463 1481
rect 565 1481 631 1491
rect 565 1467 581 1481
rect 409 1431 463 1447
rect 505 1447 581 1467
rect 615 1447 631 1481
rect 505 1437 631 1447
rect 284 1399 314 1431
rect 409 1399 439 1431
rect 505 1399 535 1437
rect 673 1399 703 1544
rect 1559 1610 1589 1642
rect 1559 1594 1613 1610
rect 1559 1560 1569 1594
rect 1603 1560 1613 1594
rect 1559 1544 1613 1560
rect 1559 1399 1589 1544
rect 1655 1491 1685 1642
rect 1727 1610 1757 1642
rect 1941 1627 1971 1642
rect 1727 1594 1781 1610
rect 1727 1560 1737 1594
rect 1771 1560 1781 1594
rect 1727 1544 1781 1560
rect 1823 1597 1971 1627
rect 1823 1497 1853 1597
rect 2044 1533 2074 1642
rect 2580 1726 2610 1752
rect 2683 1726 2713 1752
rect 2897 1726 2927 1752
rect 2969 1726 2999 1752
rect 3065 1726 3095 1752
rect 3951 1726 3981 1752
rect 4047 1726 4077 1752
rect 4119 1726 4149 1752
rect 4333 1726 4363 1752
rect 4436 1726 4466 1752
rect 2153 1533 2183 1565
rect 2471 1533 2501 1565
rect 2580 1533 2610 1642
rect 2683 1627 2713 1642
rect 2683 1597 2831 1627
rect 2897 1610 2927 1642
rect 2036 1517 2090 1533
rect 1631 1481 1697 1491
rect 1631 1447 1647 1481
rect 1681 1467 1697 1481
rect 1799 1481 1853 1497
rect 1681 1447 1757 1467
rect 1631 1437 1757 1447
rect 1727 1399 1757 1437
rect 1799 1447 1809 1481
rect 1843 1447 1853 1481
rect 1799 1431 1853 1447
rect 1895 1481 1978 1497
rect 1895 1447 1905 1481
rect 1939 1447 1978 1481
rect 2036 1483 2046 1517
rect 2080 1483 2090 1517
rect 2036 1467 2090 1483
rect 2132 1517 2186 1533
rect 2132 1483 2142 1517
rect 2176 1483 2186 1517
rect 2132 1467 2186 1483
rect 2468 1517 2522 1533
rect 2468 1483 2478 1517
rect 2512 1483 2522 1517
rect 2468 1467 2522 1483
rect 2564 1517 2618 1533
rect 2564 1483 2574 1517
rect 2608 1483 2618 1517
rect 2801 1497 2831 1597
rect 2873 1594 2927 1610
rect 2873 1560 2883 1594
rect 2917 1560 2927 1594
rect 2873 1544 2927 1560
rect 2564 1467 2618 1483
rect 2676 1481 2759 1497
rect 1895 1431 1978 1447
rect 1823 1399 1853 1431
rect 1948 1399 1978 1431
rect 2044 1399 2074 1467
rect 2153 1445 2183 1467
rect 2471 1445 2501 1467
rect 2580 1399 2610 1467
rect 2676 1447 2715 1481
rect 2749 1447 2759 1481
rect 2676 1431 2759 1447
rect 2801 1481 2855 1497
rect 2969 1491 2999 1642
rect 3065 1610 3095 1642
rect 3041 1594 3095 1610
rect 3041 1560 3051 1594
rect 3085 1560 3095 1594
rect 3041 1544 3095 1560
rect 2801 1447 2811 1481
rect 2845 1447 2855 1481
rect 2957 1481 3023 1491
rect 2957 1467 2973 1481
rect 2801 1431 2855 1447
rect 2897 1447 2973 1467
rect 3007 1447 3023 1481
rect 2897 1437 3023 1447
rect 2676 1399 2706 1431
rect 2801 1399 2831 1431
rect 2897 1399 2927 1437
rect 3065 1399 3095 1544
rect 3951 1610 3981 1642
rect 3951 1594 4005 1610
rect 3951 1560 3961 1594
rect 3995 1560 4005 1594
rect 3951 1544 4005 1560
rect 3951 1399 3981 1544
rect 4047 1491 4077 1642
rect 4119 1610 4149 1642
rect 4333 1627 4363 1642
rect 4119 1594 4173 1610
rect 4119 1560 4129 1594
rect 4163 1560 4173 1594
rect 4119 1544 4173 1560
rect 4215 1597 4363 1627
rect 4215 1497 4245 1597
rect 4436 1533 4466 1642
rect 4972 1726 5002 1752
rect 5075 1726 5105 1752
rect 5289 1726 5319 1752
rect 5361 1726 5391 1752
rect 5457 1726 5487 1752
rect 6341 1726 6371 1752
rect 6437 1726 6467 1752
rect 6509 1726 6539 1752
rect 6723 1726 6753 1752
rect 6826 1726 6856 1752
rect 4545 1533 4575 1565
rect 4863 1533 4893 1565
rect 4972 1533 5002 1642
rect 5075 1627 5105 1642
rect 5075 1597 5223 1627
rect 5289 1610 5319 1642
rect 4428 1517 4482 1533
rect 4023 1481 4089 1491
rect 4023 1447 4039 1481
rect 4073 1467 4089 1481
rect 4191 1481 4245 1497
rect 4073 1447 4149 1467
rect 4023 1437 4149 1447
rect 4119 1399 4149 1437
rect 4191 1447 4201 1481
rect 4235 1447 4245 1481
rect 4191 1431 4245 1447
rect 4287 1481 4370 1497
rect 4287 1447 4297 1481
rect 4331 1447 4370 1481
rect 4428 1483 4438 1517
rect 4472 1483 4482 1517
rect 4428 1467 4482 1483
rect 4524 1517 4578 1533
rect 4524 1483 4534 1517
rect 4568 1483 4578 1517
rect 4524 1467 4578 1483
rect 4860 1517 4914 1533
rect 4860 1483 4870 1517
rect 4904 1483 4914 1517
rect 4860 1467 4914 1483
rect 4956 1517 5010 1533
rect 4956 1483 4966 1517
rect 5000 1483 5010 1517
rect 5193 1497 5223 1597
rect 5265 1594 5319 1610
rect 5265 1560 5275 1594
rect 5309 1560 5319 1594
rect 5265 1544 5319 1560
rect 4956 1467 5010 1483
rect 5068 1481 5151 1497
rect 4287 1431 4370 1447
rect 4215 1399 4245 1431
rect 4340 1399 4370 1431
rect 4436 1399 4466 1467
rect 4545 1445 4575 1467
rect 4863 1445 4893 1467
rect 4972 1399 5002 1467
rect 5068 1447 5107 1481
rect 5141 1447 5151 1481
rect 5068 1431 5151 1447
rect 5193 1481 5247 1497
rect 5361 1491 5391 1642
rect 5457 1610 5487 1642
rect 5433 1594 5487 1610
rect 5433 1560 5443 1594
rect 5477 1560 5487 1594
rect 5433 1544 5487 1560
rect 5193 1447 5203 1481
rect 5237 1447 5247 1481
rect 5349 1481 5415 1491
rect 5349 1467 5365 1481
rect 5193 1431 5247 1447
rect 5289 1447 5365 1467
rect 5399 1447 5415 1481
rect 5289 1437 5415 1447
rect 5068 1399 5098 1431
rect 5193 1399 5223 1431
rect 5289 1399 5319 1437
rect 5457 1399 5487 1544
rect 6341 1610 6371 1642
rect 6341 1594 6395 1610
rect 6341 1560 6351 1594
rect 6385 1560 6395 1594
rect 6341 1544 6395 1560
rect 6341 1399 6371 1544
rect 6437 1491 6467 1642
rect 6509 1610 6539 1642
rect 6723 1627 6753 1642
rect 6509 1594 6563 1610
rect 6509 1560 6519 1594
rect 6553 1560 6563 1594
rect 6509 1544 6563 1560
rect 6605 1597 6753 1627
rect 6605 1497 6635 1597
rect 6826 1533 6856 1642
rect 7364 1726 7394 1752
rect 7467 1726 7497 1752
rect 7681 1726 7711 1752
rect 7753 1726 7783 1752
rect 7849 1726 7879 1752
rect 8735 1726 8765 1752
rect 8831 1726 8861 1752
rect 8903 1726 8933 1752
rect 9117 1726 9147 1752
rect 9220 1726 9250 1752
rect 6935 1533 6965 1565
rect 7255 1533 7285 1565
rect 7364 1533 7394 1642
rect 7467 1627 7497 1642
rect 7467 1597 7615 1627
rect 7681 1610 7711 1642
rect 6818 1517 6872 1533
rect 6413 1481 6479 1491
rect 6413 1447 6429 1481
rect 6463 1467 6479 1481
rect 6581 1481 6635 1497
rect 6463 1447 6539 1467
rect 6413 1437 6539 1447
rect 6509 1399 6539 1437
rect 6581 1447 6591 1481
rect 6625 1447 6635 1481
rect 6581 1431 6635 1447
rect 6677 1481 6760 1497
rect 6677 1447 6687 1481
rect 6721 1447 6760 1481
rect 6818 1483 6828 1517
rect 6862 1483 6872 1517
rect 6818 1467 6872 1483
rect 6914 1517 6968 1533
rect 6914 1483 6924 1517
rect 6958 1483 6968 1517
rect 6914 1467 6968 1483
rect 7252 1517 7306 1533
rect 7252 1483 7262 1517
rect 7296 1483 7306 1517
rect 7252 1467 7306 1483
rect 7348 1517 7402 1533
rect 7348 1483 7358 1517
rect 7392 1483 7402 1517
rect 7585 1497 7615 1597
rect 7657 1594 7711 1610
rect 7657 1560 7667 1594
rect 7701 1560 7711 1594
rect 7657 1544 7711 1560
rect 7348 1467 7402 1483
rect 7460 1481 7543 1497
rect 6677 1431 6760 1447
rect 6605 1399 6635 1431
rect 6730 1399 6760 1431
rect 6826 1399 6856 1467
rect 6935 1445 6965 1467
rect 7255 1445 7285 1467
rect 7364 1399 7394 1467
rect 7460 1447 7499 1481
rect 7533 1447 7543 1481
rect 7460 1431 7543 1447
rect 7585 1481 7639 1497
rect 7753 1491 7783 1642
rect 7849 1610 7879 1642
rect 7825 1594 7879 1610
rect 7825 1560 7835 1594
rect 7869 1560 7879 1594
rect 7825 1544 7879 1560
rect 7585 1447 7595 1481
rect 7629 1447 7639 1481
rect 7741 1481 7807 1491
rect 7741 1467 7757 1481
rect 7585 1431 7639 1447
rect 7681 1447 7757 1467
rect 7791 1447 7807 1481
rect 7681 1437 7807 1447
rect 7460 1399 7490 1431
rect 7585 1399 7615 1431
rect 7681 1399 7711 1437
rect 7849 1399 7879 1544
rect 8735 1610 8765 1642
rect 8735 1594 8789 1610
rect 8735 1560 8745 1594
rect 8779 1560 8789 1594
rect 8735 1544 8789 1560
rect 8735 1399 8765 1544
rect 8831 1491 8861 1642
rect 8903 1610 8933 1642
rect 9117 1627 9147 1642
rect 8903 1594 8957 1610
rect 8903 1560 8913 1594
rect 8947 1560 8957 1594
rect 8903 1544 8957 1560
rect 8999 1597 9147 1627
rect 8999 1497 9029 1597
rect 9220 1533 9250 1642
rect 9756 1726 9786 1752
rect 9859 1726 9889 1752
rect 10073 1726 10103 1752
rect 10145 1726 10175 1752
rect 10241 1726 10271 1752
rect 11127 1726 11157 1752
rect 11223 1726 11253 1752
rect 11295 1726 11325 1752
rect 11509 1726 11539 1752
rect 11612 1726 11642 1752
rect 9329 1533 9359 1565
rect 9647 1533 9677 1565
rect 9756 1533 9786 1642
rect 9859 1627 9889 1642
rect 9859 1597 10007 1627
rect 10073 1610 10103 1642
rect 9212 1517 9266 1533
rect 8807 1481 8873 1491
rect 8807 1447 8823 1481
rect 8857 1467 8873 1481
rect 8975 1481 9029 1497
rect 8857 1447 8933 1467
rect 8807 1437 8933 1447
rect 8903 1399 8933 1437
rect 8975 1447 8985 1481
rect 9019 1447 9029 1481
rect 8975 1431 9029 1447
rect 9071 1481 9154 1497
rect 9071 1447 9081 1481
rect 9115 1447 9154 1481
rect 9212 1483 9222 1517
rect 9256 1483 9266 1517
rect 9212 1467 9266 1483
rect 9308 1517 9362 1533
rect 9308 1483 9318 1517
rect 9352 1483 9362 1517
rect 9308 1467 9362 1483
rect 9644 1517 9698 1533
rect 9644 1483 9654 1517
rect 9688 1483 9698 1517
rect 9644 1467 9698 1483
rect 9740 1517 9794 1533
rect 9740 1483 9750 1517
rect 9784 1483 9794 1517
rect 9977 1497 10007 1597
rect 10049 1594 10103 1610
rect 10049 1560 10059 1594
rect 10093 1560 10103 1594
rect 10049 1544 10103 1560
rect 9740 1467 9794 1483
rect 9852 1481 9935 1497
rect 9071 1431 9154 1447
rect 8999 1399 9029 1431
rect 9124 1399 9154 1431
rect 9220 1399 9250 1467
rect 9329 1445 9359 1467
rect 9647 1445 9677 1467
rect 9756 1399 9786 1467
rect 9852 1447 9891 1481
rect 9925 1447 9935 1481
rect 9852 1431 9935 1447
rect 9977 1481 10031 1497
rect 10145 1491 10175 1642
rect 10241 1610 10271 1642
rect 10217 1594 10271 1610
rect 10217 1560 10227 1594
rect 10261 1560 10271 1594
rect 10217 1544 10271 1560
rect 9977 1447 9987 1481
rect 10021 1447 10031 1481
rect 10133 1481 10199 1491
rect 10133 1467 10149 1481
rect 9977 1431 10031 1447
rect 10073 1447 10149 1467
rect 10183 1447 10199 1481
rect 10073 1437 10199 1447
rect 9852 1399 9882 1431
rect 9977 1399 10007 1431
rect 10073 1399 10103 1437
rect 10241 1399 10271 1544
rect 11127 1610 11157 1642
rect 11127 1594 11181 1610
rect 11127 1560 11137 1594
rect 11171 1560 11181 1594
rect 11127 1544 11181 1560
rect 11127 1399 11157 1544
rect 11223 1491 11253 1642
rect 11295 1610 11325 1642
rect 11509 1627 11539 1642
rect 11295 1594 11349 1610
rect 11295 1560 11305 1594
rect 11339 1560 11349 1594
rect 11295 1544 11349 1560
rect 11391 1597 11539 1627
rect 11391 1497 11421 1597
rect 11612 1533 11642 1642
rect 12148 1726 12178 1752
rect 12251 1726 12281 1752
rect 12465 1726 12495 1752
rect 12537 1726 12567 1752
rect 12633 1726 12663 1752
rect 13517 1726 13547 1752
rect 13613 1726 13643 1752
rect 13685 1726 13715 1752
rect 13899 1726 13929 1752
rect 14002 1726 14032 1752
rect 11721 1533 11751 1565
rect 12039 1533 12069 1565
rect 12148 1533 12178 1642
rect 12251 1627 12281 1642
rect 12251 1597 12399 1627
rect 12465 1610 12495 1642
rect 11604 1517 11658 1533
rect 11199 1481 11265 1491
rect 11199 1447 11215 1481
rect 11249 1467 11265 1481
rect 11367 1481 11421 1497
rect 11249 1447 11325 1467
rect 11199 1437 11325 1447
rect 11295 1399 11325 1437
rect 11367 1447 11377 1481
rect 11411 1447 11421 1481
rect 11367 1431 11421 1447
rect 11463 1481 11546 1497
rect 11463 1447 11473 1481
rect 11507 1447 11546 1481
rect 11604 1483 11614 1517
rect 11648 1483 11658 1517
rect 11604 1467 11658 1483
rect 11700 1517 11754 1533
rect 11700 1483 11710 1517
rect 11744 1483 11754 1517
rect 11700 1467 11754 1483
rect 12036 1517 12090 1533
rect 12036 1483 12046 1517
rect 12080 1483 12090 1517
rect 12036 1467 12090 1483
rect 12132 1517 12186 1533
rect 12132 1483 12142 1517
rect 12176 1483 12186 1517
rect 12369 1497 12399 1597
rect 12441 1594 12495 1610
rect 12441 1560 12451 1594
rect 12485 1560 12495 1594
rect 12441 1544 12495 1560
rect 12132 1467 12186 1483
rect 12244 1481 12327 1497
rect 11463 1431 11546 1447
rect 11391 1399 11421 1431
rect 11516 1399 11546 1431
rect 11612 1399 11642 1467
rect 11721 1445 11751 1467
rect 12039 1445 12069 1467
rect 12148 1399 12178 1467
rect 12244 1447 12283 1481
rect 12317 1447 12327 1481
rect 12244 1431 12327 1447
rect 12369 1481 12423 1497
rect 12537 1491 12567 1642
rect 12633 1610 12663 1642
rect 12609 1594 12663 1610
rect 12609 1560 12619 1594
rect 12653 1560 12663 1594
rect 12609 1544 12663 1560
rect 12369 1447 12379 1481
rect 12413 1447 12423 1481
rect 12525 1481 12591 1491
rect 12525 1467 12541 1481
rect 12369 1431 12423 1447
rect 12465 1447 12541 1467
rect 12575 1447 12591 1481
rect 12465 1437 12591 1447
rect 12244 1399 12274 1431
rect 12369 1399 12399 1431
rect 12465 1399 12495 1437
rect 12633 1399 12663 1544
rect 13517 1610 13547 1642
rect 13517 1594 13571 1610
rect 13517 1560 13527 1594
rect 13561 1560 13571 1594
rect 13517 1544 13571 1560
rect 13517 1399 13547 1544
rect 13613 1491 13643 1642
rect 13685 1610 13715 1642
rect 13899 1627 13929 1642
rect 13685 1594 13739 1610
rect 13685 1560 13695 1594
rect 13729 1560 13739 1594
rect 13685 1544 13739 1560
rect 13781 1597 13929 1627
rect 13781 1497 13811 1597
rect 14002 1533 14032 1642
rect 14540 1726 14570 1752
rect 14643 1726 14673 1752
rect 14857 1726 14887 1752
rect 14929 1726 14959 1752
rect 15025 1726 15055 1752
rect 15911 1726 15941 1752
rect 16007 1726 16037 1752
rect 16079 1726 16109 1752
rect 16293 1726 16323 1752
rect 16396 1726 16426 1752
rect 14111 1533 14141 1565
rect 14431 1533 14461 1565
rect 14540 1533 14570 1642
rect 14643 1627 14673 1642
rect 14643 1597 14791 1627
rect 14857 1610 14887 1642
rect 13994 1517 14048 1533
rect 13589 1481 13655 1491
rect 13589 1447 13605 1481
rect 13639 1467 13655 1481
rect 13757 1481 13811 1497
rect 13639 1447 13715 1467
rect 13589 1437 13715 1447
rect 13685 1399 13715 1437
rect 13757 1447 13767 1481
rect 13801 1447 13811 1481
rect 13757 1431 13811 1447
rect 13853 1481 13936 1497
rect 13853 1447 13863 1481
rect 13897 1447 13936 1481
rect 13994 1483 14004 1517
rect 14038 1483 14048 1517
rect 13994 1467 14048 1483
rect 14090 1517 14144 1533
rect 14090 1483 14100 1517
rect 14134 1483 14144 1517
rect 14090 1467 14144 1483
rect 14428 1517 14482 1533
rect 14428 1483 14438 1517
rect 14472 1483 14482 1517
rect 14428 1467 14482 1483
rect 14524 1517 14578 1533
rect 14524 1483 14534 1517
rect 14568 1483 14578 1517
rect 14761 1497 14791 1597
rect 14833 1594 14887 1610
rect 14833 1560 14843 1594
rect 14877 1560 14887 1594
rect 14833 1544 14887 1560
rect 14524 1467 14578 1483
rect 14636 1481 14719 1497
rect 13853 1431 13936 1447
rect 13781 1399 13811 1431
rect 13906 1399 13936 1431
rect 14002 1399 14032 1467
rect 14111 1445 14141 1467
rect 14431 1445 14461 1467
rect 14540 1399 14570 1467
rect 14636 1447 14675 1481
rect 14709 1447 14719 1481
rect 14636 1431 14719 1447
rect 14761 1481 14815 1497
rect 14929 1491 14959 1642
rect 15025 1610 15055 1642
rect 15001 1594 15055 1610
rect 15001 1560 15011 1594
rect 15045 1560 15055 1594
rect 15001 1544 15055 1560
rect 14761 1447 14771 1481
rect 14805 1447 14815 1481
rect 14917 1481 14983 1491
rect 14917 1467 14933 1481
rect 14761 1431 14815 1447
rect 14857 1447 14933 1467
rect 14967 1447 14983 1481
rect 14857 1437 14983 1447
rect 14636 1399 14666 1431
rect 14761 1399 14791 1431
rect 14857 1399 14887 1437
rect 15025 1399 15055 1544
rect 15911 1610 15941 1642
rect 15911 1594 15965 1610
rect 15911 1560 15921 1594
rect 15955 1560 15965 1594
rect 15911 1544 15965 1560
rect 15911 1399 15941 1544
rect 16007 1491 16037 1642
rect 16079 1610 16109 1642
rect 16293 1627 16323 1642
rect 16079 1594 16133 1610
rect 16079 1560 16089 1594
rect 16123 1560 16133 1594
rect 16079 1544 16133 1560
rect 16175 1597 16323 1627
rect 16175 1497 16205 1597
rect 16396 1533 16426 1642
rect 16505 1533 16535 1565
rect 16388 1517 16442 1533
rect 15983 1481 16049 1491
rect 15983 1447 15999 1481
rect 16033 1467 16049 1481
rect 16151 1481 16205 1497
rect 16033 1447 16109 1467
rect 15983 1437 16109 1447
rect 16079 1399 16109 1437
rect 16151 1447 16161 1481
rect 16195 1447 16205 1481
rect 16151 1431 16205 1447
rect 16247 1481 16330 1497
rect 16247 1447 16257 1481
rect 16291 1447 16330 1481
rect 16388 1483 16398 1517
rect 16432 1483 16442 1517
rect 16388 1467 16442 1483
rect 16484 1517 16538 1533
rect 16484 1483 16494 1517
rect 16528 1483 16538 1517
rect 16484 1467 16538 1483
rect 16247 1431 16330 1447
rect 16175 1399 16205 1431
rect 16300 1399 16330 1431
rect 16396 1399 16426 1467
rect 16505 1445 16535 1467
rect 79 1289 109 1315
rect 188 1289 218 1315
rect 284 1289 314 1315
rect 409 1289 439 1315
rect 505 1289 535 1315
rect 673 1289 703 1315
rect 1559 1289 1589 1315
rect 1727 1289 1757 1315
rect 1823 1289 1853 1315
rect 1948 1289 1978 1315
rect 2044 1289 2074 1315
rect 2153 1289 2183 1315
rect 2471 1289 2501 1315
rect 2580 1289 2610 1315
rect 2676 1289 2706 1315
rect 2801 1289 2831 1315
rect 2897 1289 2927 1315
rect 3065 1289 3095 1315
rect 3951 1289 3981 1315
rect 4119 1289 4149 1315
rect 4215 1289 4245 1315
rect 4340 1289 4370 1315
rect 4436 1289 4466 1315
rect 4545 1289 4575 1315
rect 4863 1289 4893 1315
rect 4972 1289 5002 1315
rect 5068 1289 5098 1315
rect 5193 1289 5223 1315
rect 5289 1289 5319 1315
rect 5457 1289 5487 1315
rect 6341 1289 6371 1315
rect 6509 1289 6539 1315
rect 6605 1289 6635 1315
rect 6730 1289 6760 1315
rect 6826 1289 6856 1315
rect 6935 1289 6965 1315
rect 7255 1289 7285 1315
rect 7364 1289 7394 1315
rect 7460 1289 7490 1315
rect 7585 1289 7615 1315
rect 7681 1289 7711 1315
rect 7849 1289 7879 1315
rect 8735 1289 8765 1315
rect 8903 1289 8933 1315
rect 8999 1289 9029 1315
rect 9124 1289 9154 1315
rect 9220 1289 9250 1315
rect 9329 1289 9359 1315
rect 9647 1289 9677 1315
rect 9756 1289 9786 1315
rect 9852 1289 9882 1315
rect 9977 1289 10007 1315
rect 10073 1289 10103 1315
rect 10241 1289 10271 1315
rect 11127 1289 11157 1315
rect 11295 1289 11325 1315
rect 11391 1289 11421 1315
rect 11516 1289 11546 1315
rect 11612 1289 11642 1315
rect 11721 1289 11751 1315
rect 12039 1289 12069 1315
rect 12148 1289 12178 1315
rect 12244 1289 12274 1315
rect 12369 1289 12399 1315
rect 12465 1289 12495 1315
rect 12633 1289 12663 1315
rect 13517 1289 13547 1315
rect 13685 1289 13715 1315
rect 13781 1289 13811 1315
rect 13906 1289 13936 1315
rect 14002 1289 14032 1315
rect 14111 1289 14141 1315
rect 14431 1289 14461 1315
rect 14540 1289 14570 1315
rect 14636 1289 14666 1315
rect 14761 1289 14791 1315
rect 14857 1289 14887 1315
rect 15025 1289 15055 1315
rect 15911 1289 15941 1315
rect 16079 1289 16109 1315
rect 16175 1289 16205 1315
rect 16300 1289 16330 1315
rect 16396 1289 16426 1315
rect 16505 1289 16535 1315
rect 1885 1158 1951 1174
rect 1885 1124 1901 1158
rect 1935 1124 1951 1158
rect 4277 1157 4343 1173
rect 1885 1108 1951 1124
rect 4277 1123 4293 1157
rect 4327 1123 4343 1157
rect 6669 1157 6735 1173
rect 79 1071 109 1097
rect 163 1071 193 1097
rect 351 1077 381 1103
rect 443 1077 473 1103
rect 527 1077 557 1103
rect 647 1077 677 1103
rect 753 1077 783 1103
rect 861 1077 891 1103
rect 945 1077 975 1103
rect 1082 1077 1112 1103
rect 1226 1077 1256 1103
rect 1310 1077 1340 1103
rect 1415 1077 1445 1103
rect 1536 1077 1566 1103
rect 1642 1077 1672 1103
rect 1714 1077 1744 1103
rect 79 928 109 943
rect 45 898 109 928
rect 45 860 75 898
rect 21 844 75 860
rect 163 854 193 943
rect 21 810 31 844
rect 65 810 75 844
rect 21 794 75 810
rect 117 844 193 854
rect 351 847 381 993
rect 443 859 473 993
rect 527 955 557 993
rect 647 961 677 993
rect 515 945 581 955
rect 515 911 531 945
rect 565 911 581 945
rect 515 901 581 911
rect 647 945 711 961
rect 647 911 667 945
rect 701 911 711 945
rect 647 895 711 911
rect 117 810 133 844
rect 167 810 193 844
rect 117 800 193 810
rect 45 756 75 794
rect 45 726 109 756
rect 79 711 109 726
rect 163 711 193 800
rect 339 831 393 847
rect 339 797 349 831
rect 383 797 393 831
rect 443 829 581 859
rect 339 781 393 797
rect 551 799 581 829
rect 351 711 381 781
rect 446 771 509 787
rect 446 737 465 771
rect 499 737 509 771
rect 446 721 509 737
rect 551 783 605 799
rect 551 749 561 783
rect 595 749 605 783
rect 551 733 605 749
rect 446 699 476 721
rect 551 699 581 733
rect 647 711 677 895
rect 753 809 783 993
rect 1226 961 1256 993
rect 1202 945 1256 961
rect 1310 955 1340 993
rect 1415 961 1445 993
rect 1202 911 1212 945
rect 1246 911 1256 945
rect 861 877 891 909
rect 945 877 975 909
rect 825 861 891 877
rect 825 827 835 861
rect 869 827 891 861
rect 825 811 891 827
rect 941 861 1031 877
rect 941 827 987 861
rect 1021 827 1031 861
rect 941 811 1031 827
rect 1082 843 1112 909
rect 1202 895 1256 911
rect 1298 945 1364 955
rect 1298 911 1314 945
rect 1348 911 1364 945
rect 1298 901 1364 911
rect 1415 945 1494 961
rect 1415 911 1450 945
rect 1484 911 1494 945
rect 1415 895 1494 911
rect 1226 859 1256 895
rect 1082 827 1159 843
rect 1226 829 1363 859
rect 1082 813 1115 827
rect 723 793 783 809
rect 723 759 733 793
rect 767 773 783 793
rect 767 759 791 773
rect 723 743 791 759
rect 857 755 887 811
rect 941 755 971 811
rect 1105 793 1115 813
rect 1149 793 1159 827
rect 1105 777 1159 793
rect 1129 755 1159 777
rect 1237 771 1291 787
rect 761 711 791 743
rect 1237 737 1247 771
rect 1281 737 1291 771
rect 1237 721 1291 737
rect 1249 699 1279 721
rect 1333 699 1363 829
rect 1428 711 1458 895
rect 1536 816 1566 993
rect 1903 1009 1933 1108
rect 4277 1107 4343 1123
rect 6669 1123 6685 1157
rect 6719 1123 6735 1157
rect 9061 1158 9127 1174
rect 6669 1107 6735 1123
rect 9061 1124 9077 1158
rect 9111 1124 9127 1158
rect 11453 1158 11519 1174
rect 9061 1108 9127 1124
rect 11453 1124 11469 1158
rect 11503 1124 11519 1158
rect 13845 1157 13911 1173
rect 11453 1108 11519 1124
rect 13845 1123 13861 1157
rect 13895 1123 13911 1157
rect 16237 1157 16303 1173
rect 2000 1077 2030 1103
rect 1642 861 1672 909
rect 1501 793 1566 816
rect 1608 845 1672 861
rect 1608 811 1618 845
rect 1652 811 1672 845
rect 1714 877 1744 909
rect 1714 861 1798 877
rect 1714 827 1754 861
rect 1788 827 1798 861
rect 1903 849 1933 881
rect 2188 1061 2218 1087
rect 2283 1077 2313 1103
rect 2188 917 2218 933
rect 2163 887 2218 917
rect 1714 811 1798 827
rect 1853 833 1935 849
rect 2000 845 2030 877
rect 1608 795 1672 811
rect 1501 759 1511 793
rect 1545 786 1566 793
rect 1545 759 1555 786
rect 1501 743 1555 759
rect 1633 755 1663 795
rect 1717 755 1747 811
rect 1853 799 1863 833
rect 1897 799 1935 833
rect 1853 783 1935 799
rect 1525 711 1555 743
rect 1905 711 1935 783
rect 1981 839 2035 845
rect 2163 839 2193 887
rect 2471 1071 2501 1097
rect 2555 1071 2585 1097
rect 2743 1077 2773 1103
rect 2835 1077 2865 1103
rect 2919 1077 2949 1103
rect 3039 1077 3069 1103
rect 3145 1077 3175 1103
rect 3253 1077 3283 1103
rect 3337 1077 3367 1103
rect 3474 1077 3504 1103
rect 3618 1077 3648 1103
rect 3702 1077 3732 1103
rect 3807 1077 3837 1103
rect 3928 1077 3958 1103
rect 4034 1077 4064 1103
rect 4106 1077 4136 1103
rect 2471 928 2501 943
rect 2437 898 2501 928
rect 2283 845 2313 877
rect 2437 860 2467 898
rect 1981 829 2193 839
rect 1981 795 1991 829
rect 2025 795 2193 829
rect 1981 785 2193 795
rect 1981 779 2030 785
rect 2000 757 2030 779
rect 2163 756 2193 785
rect 2255 829 2314 845
rect 2255 795 2265 829
rect 2299 795 2314 829
rect 2255 779 2314 795
rect 2413 844 2467 860
rect 2555 854 2585 943
rect 2413 810 2423 844
rect 2457 810 2467 844
rect 2413 794 2467 810
rect 2509 844 2585 854
rect 2743 847 2773 993
rect 2835 859 2865 993
rect 2919 955 2949 993
rect 3039 961 3069 993
rect 2907 945 2973 955
rect 2907 911 2923 945
rect 2957 911 2973 945
rect 2907 901 2973 911
rect 3039 945 3103 961
rect 3039 911 3059 945
rect 3093 911 3103 945
rect 3039 895 3103 911
rect 2509 810 2525 844
rect 2559 810 2585 844
rect 2509 800 2585 810
rect 2283 757 2313 779
rect 2163 726 2218 756
rect 2188 711 2218 726
rect 2437 756 2467 794
rect 2437 726 2501 756
rect 2471 711 2501 726
rect 2555 711 2585 800
rect 2731 831 2785 847
rect 2731 797 2741 831
rect 2775 797 2785 831
rect 2835 829 2973 859
rect 2731 781 2785 797
rect 2943 799 2973 829
rect 2743 711 2773 781
rect 2838 771 2901 787
rect 2838 737 2857 771
rect 2891 737 2901 771
rect 2838 721 2901 737
rect 2943 783 2997 799
rect 2943 749 2953 783
rect 2987 749 2997 783
rect 2943 733 2997 749
rect 2838 699 2868 721
rect 2943 699 2973 733
rect 3039 711 3069 895
rect 3145 809 3175 993
rect 3618 961 3648 993
rect 3594 945 3648 961
rect 3702 955 3732 993
rect 3807 961 3837 993
rect 3594 911 3604 945
rect 3638 911 3648 945
rect 3253 877 3283 909
rect 3337 877 3367 909
rect 3217 861 3283 877
rect 3217 827 3227 861
rect 3261 827 3283 861
rect 3217 811 3283 827
rect 3333 861 3423 877
rect 3333 827 3379 861
rect 3413 827 3423 861
rect 3333 811 3423 827
rect 3474 843 3504 909
rect 3594 895 3648 911
rect 3690 945 3756 955
rect 3690 911 3706 945
rect 3740 911 3756 945
rect 3690 901 3756 911
rect 3807 945 3886 961
rect 3807 911 3842 945
rect 3876 911 3886 945
rect 3807 895 3886 911
rect 3618 859 3648 895
rect 3474 827 3551 843
rect 3618 829 3755 859
rect 3474 813 3507 827
rect 3115 793 3175 809
rect 3115 759 3125 793
rect 3159 773 3175 793
rect 3159 759 3183 773
rect 3115 743 3183 759
rect 3249 755 3279 811
rect 3333 755 3363 811
rect 3497 793 3507 813
rect 3541 793 3551 827
rect 3497 777 3551 793
rect 3521 755 3551 777
rect 3629 771 3683 787
rect 3153 711 3183 743
rect 3629 737 3639 771
rect 3673 737 3683 771
rect 3629 721 3683 737
rect 3641 699 3671 721
rect 3725 699 3755 829
rect 3820 711 3850 895
rect 3928 816 3958 993
rect 4295 1009 4325 1107
rect 4392 1077 4422 1103
rect 4034 861 4064 909
rect 3893 793 3958 816
rect 4000 845 4064 861
rect 4000 811 4010 845
rect 4044 811 4064 845
rect 4106 877 4136 909
rect 4106 861 4190 877
rect 4106 827 4146 861
rect 4180 827 4190 861
rect 4295 849 4325 881
rect 4580 1061 4610 1087
rect 4675 1077 4705 1103
rect 4580 917 4610 933
rect 4555 887 4610 917
rect 4106 811 4190 827
rect 4245 833 4327 849
rect 4392 845 4422 877
rect 4000 795 4064 811
rect 3893 759 3903 793
rect 3937 786 3958 793
rect 3937 759 3947 786
rect 3893 743 3947 759
rect 4025 755 4055 795
rect 4109 755 4139 811
rect 4245 799 4255 833
rect 4289 799 4327 833
rect 4245 783 4327 799
rect 3917 711 3947 743
rect 4297 711 4327 783
rect 4373 839 4427 845
rect 4555 839 4585 887
rect 4863 1071 4893 1097
rect 4947 1071 4977 1097
rect 5135 1077 5165 1103
rect 5227 1077 5257 1103
rect 5311 1077 5341 1103
rect 5431 1077 5461 1103
rect 5537 1077 5567 1103
rect 5645 1077 5675 1103
rect 5729 1077 5759 1103
rect 5866 1077 5896 1103
rect 6010 1077 6040 1103
rect 6094 1077 6124 1103
rect 6199 1077 6229 1103
rect 6320 1077 6350 1103
rect 6426 1077 6456 1103
rect 6498 1077 6528 1103
rect 4863 928 4893 943
rect 4829 898 4893 928
rect 4675 845 4705 877
rect 4829 860 4859 898
rect 4373 829 4585 839
rect 4373 795 4383 829
rect 4417 795 4585 829
rect 4373 785 4585 795
rect 4373 779 4422 785
rect 4392 757 4422 779
rect 4555 756 4585 785
rect 4647 829 4706 845
rect 4647 795 4657 829
rect 4691 795 4706 829
rect 4647 779 4706 795
rect 4805 844 4859 860
rect 4947 854 4977 943
rect 4805 810 4815 844
rect 4849 810 4859 844
rect 4805 794 4859 810
rect 4901 844 4977 854
rect 5135 847 5165 993
rect 5227 859 5257 993
rect 5311 955 5341 993
rect 5431 961 5461 993
rect 5299 945 5365 955
rect 5299 911 5315 945
rect 5349 911 5365 945
rect 5299 901 5365 911
rect 5431 945 5495 961
rect 5431 911 5451 945
rect 5485 911 5495 945
rect 5431 895 5495 911
rect 4901 810 4917 844
rect 4951 810 4977 844
rect 4901 800 4977 810
rect 4675 757 4705 779
rect 4555 726 4610 756
rect 4580 711 4610 726
rect 4829 756 4859 794
rect 4829 726 4893 756
rect 4863 711 4893 726
rect 4947 711 4977 800
rect 5123 831 5177 847
rect 5123 797 5133 831
rect 5167 797 5177 831
rect 5227 829 5365 859
rect 5123 781 5177 797
rect 5335 799 5365 829
rect 5135 711 5165 781
rect 5230 771 5293 787
rect 5230 737 5249 771
rect 5283 737 5293 771
rect 5230 721 5293 737
rect 5335 783 5389 799
rect 5335 749 5345 783
rect 5379 749 5389 783
rect 5335 733 5389 749
rect 5230 699 5260 721
rect 5335 699 5365 733
rect 5431 711 5461 895
rect 5537 809 5567 993
rect 6010 961 6040 993
rect 5986 945 6040 961
rect 6094 955 6124 993
rect 6199 961 6229 993
rect 5986 911 5996 945
rect 6030 911 6040 945
rect 5645 877 5675 909
rect 5729 877 5759 909
rect 5609 861 5675 877
rect 5609 827 5619 861
rect 5653 827 5675 861
rect 5609 811 5675 827
rect 5725 861 5815 877
rect 5725 827 5771 861
rect 5805 827 5815 861
rect 5725 811 5815 827
rect 5866 843 5896 909
rect 5986 895 6040 911
rect 6082 945 6148 955
rect 6082 911 6098 945
rect 6132 911 6148 945
rect 6082 901 6148 911
rect 6199 945 6278 961
rect 6199 911 6234 945
rect 6268 911 6278 945
rect 6199 895 6278 911
rect 6010 859 6040 895
rect 5866 827 5943 843
rect 6010 829 6147 859
rect 5866 813 5899 827
rect 5507 793 5567 809
rect 5507 759 5517 793
rect 5551 773 5567 793
rect 5551 759 5575 773
rect 5507 743 5575 759
rect 5641 755 5671 811
rect 5725 755 5755 811
rect 5889 793 5899 813
rect 5933 793 5943 827
rect 5889 777 5943 793
rect 5913 755 5943 777
rect 6021 771 6075 787
rect 5545 711 5575 743
rect 6021 737 6031 771
rect 6065 737 6075 771
rect 6021 721 6075 737
rect 6033 699 6063 721
rect 6117 699 6147 829
rect 6212 711 6242 895
rect 6320 816 6350 993
rect 6687 1009 6717 1107
rect 6784 1077 6814 1103
rect 6426 861 6456 909
rect 6285 793 6350 816
rect 6392 845 6456 861
rect 6392 811 6402 845
rect 6436 811 6456 845
rect 6498 877 6528 909
rect 6498 861 6582 877
rect 6498 827 6538 861
rect 6572 827 6582 861
rect 6687 849 6717 881
rect 6972 1061 7002 1087
rect 7067 1077 7097 1103
rect 6972 917 7002 933
rect 6947 887 7002 917
rect 6498 811 6582 827
rect 6637 833 6719 849
rect 6784 845 6814 877
rect 6392 795 6456 811
rect 6285 759 6295 793
rect 6329 786 6350 793
rect 6329 759 6339 786
rect 6285 743 6339 759
rect 6417 755 6447 795
rect 6501 755 6531 811
rect 6637 799 6647 833
rect 6681 799 6719 833
rect 6637 783 6719 799
rect 6309 711 6339 743
rect 6689 711 6719 783
rect 6765 839 6819 845
rect 6947 839 6977 887
rect 7255 1071 7285 1097
rect 7339 1071 7369 1097
rect 7527 1077 7557 1103
rect 7619 1077 7649 1103
rect 7703 1077 7733 1103
rect 7823 1077 7853 1103
rect 7929 1077 7959 1103
rect 8037 1077 8067 1103
rect 8121 1077 8151 1103
rect 8258 1077 8288 1103
rect 8402 1077 8432 1103
rect 8486 1077 8516 1103
rect 8591 1077 8621 1103
rect 8712 1077 8742 1103
rect 8818 1077 8848 1103
rect 8890 1077 8920 1103
rect 7255 928 7285 943
rect 7221 898 7285 928
rect 7067 845 7097 877
rect 7221 860 7251 898
rect 6765 829 6977 839
rect 6765 795 6775 829
rect 6809 795 6977 829
rect 6765 785 6977 795
rect 6765 779 6814 785
rect 6784 757 6814 779
rect 6947 756 6977 785
rect 7039 829 7098 845
rect 7039 795 7049 829
rect 7083 795 7098 829
rect 7039 779 7098 795
rect 7197 844 7251 860
rect 7339 854 7369 943
rect 7197 810 7207 844
rect 7241 810 7251 844
rect 7197 794 7251 810
rect 7293 844 7369 854
rect 7527 847 7557 993
rect 7619 859 7649 993
rect 7703 955 7733 993
rect 7823 961 7853 993
rect 7691 945 7757 955
rect 7691 911 7707 945
rect 7741 911 7757 945
rect 7691 901 7757 911
rect 7823 945 7887 961
rect 7823 911 7843 945
rect 7877 911 7887 945
rect 7823 895 7887 911
rect 7293 810 7309 844
rect 7343 810 7369 844
rect 7293 800 7369 810
rect 7067 757 7097 779
rect 6947 726 7002 756
rect 6972 711 7002 726
rect 7221 756 7251 794
rect 7221 726 7285 756
rect 7255 711 7285 726
rect 7339 711 7369 800
rect 7515 831 7569 847
rect 7515 797 7525 831
rect 7559 797 7569 831
rect 7619 829 7757 859
rect 7515 781 7569 797
rect 7727 799 7757 829
rect 7527 711 7557 781
rect 7622 771 7685 787
rect 7622 737 7641 771
rect 7675 737 7685 771
rect 7622 721 7685 737
rect 7727 783 7781 799
rect 7727 749 7737 783
rect 7771 749 7781 783
rect 7727 733 7781 749
rect 7622 699 7652 721
rect 7727 699 7757 733
rect 7823 711 7853 895
rect 7929 809 7959 993
rect 8402 961 8432 993
rect 8378 945 8432 961
rect 8486 955 8516 993
rect 8591 961 8621 993
rect 8378 911 8388 945
rect 8422 911 8432 945
rect 8037 877 8067 909
rect 8121 877 8151 909
rect 8001 861 8067 877
rect 8001 827 8011 861
rect 8045 827 8067 861
rect 8001 811 8067 827
rect 8117 861 8207 877
rect 8117 827 8163 861
rect 8197 827 8207 861
rect 8117 811 8207 827
rect 8258 843 8288 909
rect 8378 895 8432 911
rect 8474 945 8540 955
rect 8474 911 8490 945
rect 8524 911 8540 945
rect 8474 901 8540 911
rect 8591 945 8670 961
rect 8591 911 8626 945
rect 8660 911 8670 945
rect 8591 895 8670 911
rect 8402 859 8432 895
rect 8258 827 8335 843
rect 8402 829 8539 859
rect 8258 813 8291 827
rect 7899 793 7959 809
rect 7899 759 7909 793
rect 7943 773 7959 793
rect 7943 759 7967 773
rect 7899 743 7967 759
rect 8033 755 8063 811
rect 8117 755 8147 811
rect 8281 793 8291 813
rect 8325 793 8335 827
rect 8281 777 8335 793
rect 8305 755 8335 777
rect 8413 771 8467 787
rect 7937 711 7967 743
rect 8413 737 8423 771
rect 8457 737 8467 771
rect 8413 721 8467 737
rect 8425 699 8455 721
rect 8509 699 8539 829
rect 8604 711 8634 895
rect 8712 816 8742 993
rect 9079 1009 9109 1108
rect 9176 1077 9206 1103
rect 8818 861 8848 909
rect 8677 793 8742 816
rect 8784 845 8848 861
rect 8784 811 8794 845
rect 8828 811 8848 845
rect 8890 877 8920 909
rect 8890 861 8974 877
rect 8890 827 8930 861
rect 8964 827 8974 861
rect 9079 849 9109 881
rect 9364 1061 9394 1087
rect 9459 1077 9489 1103
rect 9364 917 9394 933
rect 9339 887 9394 917
rect 8890 811 8974 827
rect 9029 833 9111 849
rect 9176 845 9206 877
rect 8784 795 8848 811
rect 8677 759 8687 793
rect 8721 786 8742 793
rect 8721 759 8731 786
rect 8677 743 8731 759
rect 8809 755 8839 795
rect 8893 755 8923 811
rect 9029 799 9039 833
rect 9073 799 9111 833
rect 9029 783 9111 799
rect 8701 711 8731 743
rect 9081 711 9111 783
rect 9157 839 9211 845
rect 9339 839 9369 887
rect 9647 1071 9677 1097
rect 9731 1071 9761 1097
rect 9919 1077 9949 1103
rect 10011 1077 10041 1103
rect 10095 1077 10125 1103
rect 10215 1077 10245 1103
rect 10321 1077 10351 1103
rect 10429 1077 10459 1103
rect 10513 1077 10543 1103
rect 10650 1077 10680 1103
rect 10794 1077 10824 1103
rect 10878 1077 10908 1103
rect 10983 1077 11013 1103
rect 11104 1077 11134 1103
rect 11210 1077 11240 1103
rect 11282 1077 11312 1103
rect 9647 928 9677 943
rect 9613 898 9677 928
rect 9459 845 9489 877
rect 9613 860 9643 898
rect 9157 829 9369 839
rect 9157 795 9167 829
rect 9201 795 9369 829
rect 9157 785 9369 795
rect 9157 779 9206 785
rect 9176 757 9206 779
rect 9339 756 9369 785
rect 9431 829 9490 845
rect 9431 795 9441 829
rect 9475 795 9490 829
rect 9431 779 9490 795
rect 9589 844 9643 860
rect 9731 854 9761 943
rect 9589 810 9599 844
rect 9633 810 9643 844
rect 9589 794 9643 810
rect 9685 844 9761 854
rect 9919 847 9949 993
rect 10011 859 10041 993
rect 10095 955 10125 993
rect 10215 961 10245 993
rect 10083 945 10149 955
rect 10083 911 10099 945
rect 10133 911 10149 945
rect 10083 901 10149 911
rect 10215 945 10279 961
rect 10215 911 10235 945
rect 10269 911 10279 945
rect 10215 895 10279 911
rect 9685 810 9701 844
rect 9735 810 9761 844
rect 9685 800 9761 810
rect 9459 757 9489 779
rect 9339 726 9394 756
rect 9364 711 9394 726
rect 9613 756 9643 794
rect 9613 726 9677 756
rect 9647 711 9677 726
rect 9731 711 9761 800
rect 9907 831 9961 847
rect 9907 797 9917 831
rect 9951 797 9961 831
rect 10011 829 10149 859
rect 9907 781 9961 797
rect 10119 799 10149 829
rect 9919 711 9949 781
rect 10014 771 10077 787
rect 10014 737 10033 771
rect 10067 737 10077 771
rect 10014 721 10077 737
rect 10119 783 10173 799
rect 10119 749 10129 783
rect 10163 749 10173 783
rect 10119 733 10173 749
rect 10014 699 10044 721
rect 10119 699 10149 733
rect 10215 711 10245 895
rect 10321 809 10351 993
rect 10794 961 10824 993
rect 10770 945 10824 961
rect 10878 955 10908 993
rect 10983 961 11013 993
rect 10770 911 10780 945
rect 10814 911 10824 945
rect 10429 877 10459 909
rect 10513 877 10543 909
rect 10393 861 10459 877
rect 10393 827 10403 861
rect 10437 827 10459 861
rect 10393 811 10459 827
rect 10509 861 10599 877
rect 10509 827 10555 861
rect 10589 827 10599 861
rect 10509 811 10599 827
rect 10650 843 10680 909
rect 10770 895 10824 911
rect 10866 945 10932 955
rect 10866 911 10882 945
rect 10916 911 10932 945
rect 10866 901 10932 911
rect 10983 945 11062 961
rect 10983 911 11018 945
rect 11052 911 11062 945
rect 10983 895 11062 911
rect 10794 859 10824 895
rect 10650 827 10727 843
rect 10794 829 10931 859
rect 10650 813 10683 827
rect 10291 793 10351 809
rect 10291 759 10301 793
rect 10335 773 10351 793
rect 10335 759 10359 773
rect 10291 743 10359 759
rect 10425 755 10455 811
rect 10509 755 10539 811
rect 10673 793 10683 813
rect 10717 793 10727 827
rect 10673 777 10727 793
rect 10697 755 10727 777
rect 10805 771 10859 787
rect 10329 711 10359 743
rect 10805 737 10815 771
rect 10849 737 10859 771
rect 10805 721 10859 737
rect 10817 699 10847 721
rect 10901 699 10931 829
rect 10996 711 11026 895
rect 11104 816 11134 993
rect 11471 1009 11501 1108
rect 13845 1107 13911 1123
rect 16237 1123 16253 1157
rect 16287 1123 16303 1157
rect 16237 1107 16303 1123
rect 11568 1077 11598 1103
rect 11210 861 11240 909
rect 11069 793 11134 816
rect 11176 845 11240 861
rect 11176 811 11186 845
rect 11220 811 11240 845
rect 11282 877 11312 909
rect 11282 861 11366 877
rect 11282 827 11322 861
rect 11356 827 11366 861
rect 11471 849 11501 881
rect 11756 1061 11786 1087
rect 11851 1077 11881 1103
rect 11756 917 11786 933
rect 11731 887 11786 917
rect 11282 811 11366 827
rect 11421 833 11503 849
rect 11568 845 11598 877
rect 11176 795 11240 811
rect 11069 759 11079 793
rect 11113 786 11134 793
rect 11113 759 11123 786
rect 11069 743 11123 759
rect 11201 755 11231 795
rect 11285 755 11315 811
rect 11421 799 11431 833
rect 11465 799 11503 833
rect 11421 783 11503 799
rect 11093 711 11123 743
rect 11473 711 11503 783
rect 11549 839 11603 845
rect 11731 839 11761 887
rect 12039 1071 12069 1097
rect 12123 1071 12153 1097
rect 12311 1077 12341 1103
rect 12403 1077 12433 1103
rect 12487 1077 12517 1103
rect 12607 1077 12637 1103
rect 12713 1077 12743 1103
rect 12821 1077 12851 1103
rect 12905 1077 12935 1103
rect 13042 1077 13072 1103
rect 13186 1077 13216 1103
rect 13270 1077 13300 1103
rect 13375 1077 13405 1103
rect 13496 1077 13526 1103
rect 13602 1077 13632 1103
rect 13674 1077 13704 1103
rect 12039 928 12069 943
rect 12005 898 12069 928
rect 11851 845 11881 877
rect 12005 860 12035 898
rect 11549 829 11761 839
rect 11549 795 11559 829
rect 11593 795 11761 829
rect 11549 785 11761 795
rect 11549 779 11598 785
rect 11568 757 11598 779
rect 11731 756 11761 785
rect 11823 829 11882 845
rect 11823 795 11833 829
rect 11867 795 11882 829
rect 11823 779 11882 795
rect 11981 844 12035 860
rect 12123 854 12153 943
rect 11981 810 11991 844
rect 12025 810 12035 844
rect 11981 794 12035 810
rect 12077 844 12153 854
rect 12311 847 12341 993
rect 12403 859 12433 993
rect 12487 955 12517 993
rect 12607 961 12637 993
rect 12475 945 12541 955
rect 12475 911 12491 945
rect 12525 911 12541 945
rect 12475 901 12541 911
rect 12607 945 12671 961
rect 12607 911 12627 945
rect 12661 911 12671 945
rect 12607 895 12671 911
rect 12077 810 12093 844
rect 12127 810 12153 844
rect 12077 800 12153 810
rect 11851 757 11881 779
rect 11731 726 11786 756
rect 11756 711 11786 726
rect 12005 756 12035 794
rect 12005 726 12069 756
rect 12039 711 12069 726
rect 12123 711 12153 800
rect 12299 831 12353 847
rect 12299 797 12309 831
rect 12343 797 12353 831
rect 12403 829 12541 859
rect 12299 781 12353 797
rect 12511 799 12541 829
rect 12311 711 12341 781
rect 12406 771 12469 787
rect 12406 737 12425 771
rect 12459 737 12469 771
rect 12406 721 12469 737
rect 12511 783 12565 799
rect 12511 749 12521 783
rect 12555 749 12565 783
rect 12511 733 12565 749
rect 12406 699 12436 721
rect 12511 699 12541 733
rect 12607 711 12637 895
rect 12713 809 12743 993
rect 13186 961 13216 993
rect 13162 945 13216 961
rect 13270 955 13300 993
rect 13375 961 13405 993
rect 13162 911 13172 945
rect 13206 911 13216 945
rect 12821 877 12851 909
rect 12905 877 12935 909
rect 12785 861 12851 877
rect 12785 827 12795 861
rect 12829 827 12851 861
rect 12785 811 12851 827
rect 12901 861 12991 877
rect 12901 827 12947 861
rect 12981 827 12991 861
rect 12901 811 12991 827
rect 13042 843 13072 909
rect 13162 895 13216 911
rect 13258 945 13324 955
rect 13258 911 13274 945
rect 13308 911 13324 945
rect 13258 901 13324 911
rect 13375 945 13454 961
rect 13375 911 13410 945
rect 13444 911 13454 945
rect 13375 895 13454 911
rect 13186 859 13216 895
rect 13042 827 13119 843
rect 13186 829 13323 859
rect 13042 813 13075 827
rect 12683 793 12743 809
rect 12683 759 12693 793
rect 12727 773 12743 793
rect 12727 759 12751 773
rect 12683 743 12751 759
rect 12817 755 12847 811
rect 12901 755 12931 811
rect 13065 793 13075 813
rect 13109 793 13119 827
rect 13065 777 13119 793
rect 13089 755 13119 777
rect 13197 771 13251 787
rect 12721 711 12751 743
rect 13197 737 13207 771
rect 13241 737 13251 771
rect 13197 721 13251 737
rect 13209 699 13239 721
rect 13293 699 13323 829
rect 13388 711 13418 895
rect 13496 816 13526 993
rect 13863 1009 13893 1107
rect 13960 1077 13990 1103
rect 13602 861 13632 909
rect 13461 793 13526 816
rect 13568 845 13632 861
rect 13568 811 13578 845
rect 13612 811 13632 845
rect 13674 877 13704 909
rect 13674 861 13758 877
rect 13674 827 13714 861
rect 13748 827 13758 861
rect 13863 849 13893 881
rect 14148 1061 14178 1087
rect 14243 1077 14273 1103
rect 14148 917 14178 933
rect 14123 887 14178 917
rect 13674 811 13758 827
rect 13813 833 13895 849
rect 13960 845 13990 877
rect 13568 795 13632 811
rect 13461 759 13471 793
rect 13505 786 13526 793
rect 13505 759 13515 786
rect 13461 743 13515 759
rect 13593 755 13623 795
rect 13677 755 13707 811
rect 13813 799 13823 833
rect 13857 799 13895 833
rect 13813 783 13895 799
rect 13485 711 13515 743
rect 13865 711 13895 783
rect 13941 839 13995 845
rect 14123 839 14153 887
rect 14431 1071 14461 1097
rect 14515 1071 14545 1097
rect 14703 1077 14733 1103
rect 14795 1077 14825 1103
rect 14879 1077 14909 1103
rect 14999 1077 15029 1103
rect 15105 1077 15135 1103
rect 15213 1077 15243 1103
rect 15297 1077 15327 1103
rect 15434 1077 15464 1103
rect 15578 1077 15608 1103
rect 15662 1077 15692 1103
rect 15767 1077 15797 1103
rect 15888 1077 15918 1103
rect 15994 1077 16024 1103
rect 16066 1077 16096 1103
rect 14431 928 14461 943
rect 14397 898 14461 928
rect 14243 845 14273 877
rect 14397 860 14427 898
rect 13941 829 14153 839
rect 13941 795 13951 829
rect 13985 795 14153 829
rect 13941 785 14153 795
rect 13941 779 13990 785
rect 13960 757 13990 779
rect 14123 756 14153 785
rect 14215 829 14274 845
rect 14215 795 14225 829
rect 14259 795 14274 829
rect 14215 779 14274 795
rect 14373 844 14427 860
rect 14515 854 14545 943
rect 14373 810 14383 844
rect 14417 810 14427 844
rect 14373 794 14427 810
rect 14469 844 14545 854
rect 14703 847 14733 993
rect 14795 859 14825 993
rect 14879 955 14909 993
rect 14999 961 15029 993
rect 14867 945 14933 955
rect 14867 911 14883 945
rect 14917 911 14933 945
rect 14867 901 14933 911
rect 14999 945 15063 961
rect 14999 911 15019 945
rect 15053 911 15063 945
rect 14999 895 15063 911
rect 14469 810 14485 844
rect 14519 810 14545 844
rect 14469 800 14545 810
rect 14243 757 14273 779
rect 14123 726 14178 756
rect 14148 711 14178 726
rect 14397 756 14427 794
rect 14397 726 14461 756
rect 14431 711 14461 726
rect 14515 711 14545 800
rect 14691 831 14745 847
rect 14691 797 14701 831
rect 14735 797 14745 831
rect 14795 829 14933 859
rect 14691 781 14745 797
rect 14903 799 14933 829
rect 14703 711 14733 781
rect 14798 771 14861 787
rect 14798 737 14817 771
rect 14851 737 14861 771
rect 14798 721 14861 737
rect 14903 783 14957 799
rect 14903 749 14913 783
rect 14947 749 14957 783
rect 14903 733 14957 749
rect 14798 699 14828 721
rect 14903 699 14933 733
rect 14999 711 15029 895
rect 15105 809 15135 993
rect 15578 961 15608 993
rect 15554 945 15608 961
rect 15662 955 15692 993
rect 15767 961 15797 993
rect 15554 911 15564 945
rect 15598 911 15608 945
rect 15213 877 15243 909
rect 15297 877 15327 909
rect 15177 861 15243 877
rect 15177 827 15187 861
rect 15221 827 15243 861
rect 15177 811 15243 827
rect 15293 861 15383 877
rect 15293 827 15339 861
rect 15373 827 15383 861
rect 15293 811 15383 827
rect 15434 843 15464 909
rect 15554 895 15608 911
rect 15650 945 15716 955
rect 15650 911 15666 945
rect 15700 911 15716 945
rect 15650 901 15716 911
rect 15767 945 15846 961
rect 15767 911 15802 945
rect 15836 911 15846 945
rect 15767 895 15846 911
rect 15578 859 15608 895
rect 15434 827 15511 843
rect 15578 829 15715 859
rect 15434 813 15467 827
rect 15075 793 15135 809
rect 15075 759 15085 793
rect 15119 773 15135 793
rect 15119 759 15143 773
rect 15075 743 15143 759
rect 15209 755 15239 811
rect 15293 755 15323 811
rect 15457 793 15467 813
rect 15501 793 15511 827
rect 15457 777 15511 793
rect 15481 755 15511 777
rect 15589 771 15643 787
rect 15113 711 15143 743
rect 15589 737 15599 771
rect 15633 737 15643 771
rect 15589 721 15643 737
rect 15601 699 15631 721
rect 15685 699 15715 829
rect 15780 711 15810 895
rect 15888 816 15918 993
rect 16255 1009 16285 1107
rect 16352 1077 16382 1103
rect 15994 861 16024 909
rect 15853 793 15918 816
rect 15960 845 16024 861
rect 15960 811 15970 845
rect 16004 811 16024 845
rect 16066 877 16096 909
rect 16066 861 16150 877
rect 16066 827 16106 861
rect 16140 827 16150 861
rect 16255 849 16285 881
rect 16540 1061 16570 1087
rect 16635 1077 16665 1103
rect 16540 917 16570 933
rect 16515 887 16570 917
rect 16066 811 16150 827
rect 16205 833 16287 849
rect 16352 845 16382 877
rect 15960 795 16024 811
rect 15853 759 15863 793
rect 15897 786 15918 793
rect 15897 759 15907 786
rect 15853 743 15907 759
rect 15985 755 16015 795
rect 16069 755 16099 811
rect 16205 799 16215 833
rect 16249 799 16287 833
rect 16205 783 16287 799
rect 15877 711 15907 743
rect 16257 711 16287 783
rect 16333 839 16387 845
rect 16515 839 16545 887
rect 16635 845 16665 877
rect 16333 829 16545 839
rect 16333 795 16343 829
rect 16377 795 16545 829
rect 16333 785 16545 795
rect 16333 779 16382 785
rect 16352 757 16382 779
rect 16515 756 16545 785
rect 16607 829 16666 845
rect 16607 795 16617 829
rect 16651 795 16666 829
rect 16607 779 16666 795
rect 16635 757 16665 779
rect 16515 726 16570 756
rect 16540 711 16570 726
rect 79 601 109 627
rect 163 601 193 627
rect 351 601 381 627
rect 446 601 476 627
rect 551 601 581 627
rect 647 601 677 627
rect 761 601 791 627
rect 857 601 887 627
rect 941 601 971 627
rect 1129 601 1159 627
rect 1249 601 1279 627
rect 1333 601 1363 627
rect 1428 601 1458 627
rect 1525 601 1555 627
rect 1633 601 1663 627
rect 1717 601 1747 627
rect 1905 601 1935 627
rect 2000 601 2030 627
rect 2188 601 2218 627
rect 2283 601 2313 627
rect 2471 601 2501 627
rect 2555 601 2585 627
rect 2743 601 2773 627
rect 2838 601 2868 627
rect 2943 601 2973 627
rect 3039 601 3069 627
rect 3153 601 3183 627
rect 3249 601 3279 627
rect 3333 601 3363 627
rect 3521 601 3551 627
rect 3641 601 3671 627
rect 3725 601 3755 627
rect 3820 601 3850 627
rect 3917 601 3947 627
rect 4025 601 4055 627
rect 4109 601 4139 627
rect 4297 601 4327 627
rect 4392 601 4422 627
rect 4580 601 4610 627
rect 4675 601 4705 627
rect 4863 601 4893 627
rect 4947 601 4977 627
rect 5135 601 5165 627
rect 5230 601 5260 627
rect 5335 601 5365 627
rect 5431 601 5461 627
rect 5545 601 5575 627
rect 5641 601 5671 627
rect 5725 601 5755 627
rect 5913 601 5943 627
rect 6033 601 6063 627
rect 6117 601 6147 627
rect 6212 601 6242 627
rect 6309 601 6339 627
rect 6417 601 6447 627
rect 6501 601 6531 627
rect 6689 601 6719 627
rect 6784 601 6814 627
rect 6972 601 7002 627
rect 7067 601 7097 627
rect 7255 601 7285 627
rect 7339 601 7369 627
rect 7527 601 7557 627
rect 7622 601 7652 627
rect 7727 601 7757 627
rect 7823 601 7853 627
rect 7937 601 7967 627
rect 8033 601 8063 627
rect 8117 601 8147 627
rect 8305 601 8335 627
rect 8425 601 8455 627
rect 8509 601 8539 627
rect 8604 601 8634 627
rect 8701 601 8731 627
rect 8809 601 8839 627
rect 8893 601 8923 627
rect 9081 601 9111 627
rect 9176 601 9206 627
rect 9364 601 9394 627
rect 9459 601 9489 627
rect 9647 601 9677 627
rect 9731 601 9761 627
rect 9919 601 9949 627
rect 10014 601 10044 627
rect 10119 601 10149 627
rect 10215 601 10245 627
rect 10329 601 10359 627
rect 10425 601 10455 627
rect 10509 601 10539 627
rect 10697 601 10727 627
rect 10817 601 10847 627
rect 10901 601 10931 627
rect 10996 601 11026 627
rect 11093 601 11123 627
rect 11201 601 11231 627
rect 11285 601 11315 627
rect 11473 601 11503 627
rect 11568 601 11598 627
rect 11756 601 11786 627
rect 11851 601 11881 627
rect 12039 601 12069 627
rect 12123 601 12153 627
rect 12311 601 12341 627
rect 12406 601 12436 627
rect 12511 601 12541 627
rect 12607 601 12637 627
rect 12721 601 12751 627
rect 12817 601 12847 627
rect 12901 601 12931 627
rect 13089 601 13119 627
rect 13209 601 13239 627
rect 13293 601 13323 627
rect 13388 601 13418 627
rect 13485 601 13515 627
rect 13593 601 13623 627
rect 13677 601 13707 627
rect 13865 601 13895 627
rect 13960 601 13990 627
rect 14148 601 14178 627
rect 14243 601 14273 627
rect 14431 601 14461 627
rect 14515 601 14545 627
rect 14703 601 14733 627
rect 14798 601 14828 627
rect 14903 601 14933 627
rect 14999 601 15029 627
rect 15113 601 15143 627
rect 15209 601 15239 627
rect 15293 601 15323 627
rect 15481 601 15511 627
rect 15601 601 15631 627
rect 15685 601 15715 627
rect 15780 601 15810 627
rect 15877 601 15907 627
rect 15985 601 16015 627
rect 16069 601 16099 627
rect 16257 601 16287 627
rect 16352 601 16382 627
rect 16540 601 16570 627
rect 16635 601 16665 627
rect 1591 472 1657 488
rect 1591 438 1607 472
rect 1641 438 1657 472
rect 3983 472 4049 488
rect 1591 422 1657 438
rect 3983 438 3999 472
rect 4033 438 4049 472
rect 6375 472 6441 488
rect 3983 422 4049 438
rect 6375 438 6391 472
rect 6425 438 6441 472
rect 8767 472 8833 488
rect 6375 422 6441 438
rect 8767 438 8783 472
rect 8817 438 8833 472
rect 11159 472 11225 488
rect 8767 422 8833 438
rect 11159 438 11175 472
rect 11209 438 11225 472
rect 13551 472 13617 488
rect 11159 422 11225 438
rect 13551 438 13567 472
rect 13601 438 13617 472
rect 15943 469 16009 485
rect 13551 422 13617 438
rect 15943 435 15959 469
rect 15993 435 16009 469
rect 79 388 109 414
rect 174 372 204 398
rect 362 388 392 414
rect 648 388 678 414
rect 720 388 750 414
rect 826 388 856 414
rect 947 388 977 414
rect 1052 388 1082 414
rect 1136 388 1166 414
rect 1280 388 1310 414
rect 1417 388 1447 414
rect 1501 388 1531 414
rect 1609 388 1639 422
rect 1715 388 1745 414
rect 1835 388 1865 414
rect 1919 388 1949 414
rect 2011 388 2041 414
rect 174 228 204 244
rect 174 198 229 228
rect 79 156 109 188
rect 78 140 137 156
rect 78 106 93 140
rect 127 106 137 140
rect 78 90 137 106
rect 199 150 229 198
rect 459 320 489 346
rect 362 156 392 188
rect 459 160 489 192
rect 648 188 678 220
rect 594 172 678 188
rect 357 150 411 156
rect 199 140 411 150
rect 199 106 367 140
rect 401 106 411 140
rect 199 96 411 106
rect 79 68 109 90
rect 199 67 229 96
rect 362 90 411 96
rect 457 144 539 160
rect 457 110 495 144
rect 529 110 539 144
rect 594 138 604 172
rect 638 138 678 172
rect 594 122 678 138
rect 720 172 750 220
rect 720 156 784 172
rect 720 122 740 156
rect 774 122 784 156
rect 457 94 539 110
rect 362 68 392 90
rect 174 37 229 67
rect 174 22 204 37
rect 457 22 487 94
rect 645 66 675 122
rect 720 106 784 122
rect 826 127 856 304
rect 947 272 977 304
rect 898 256 977 272
rect 1052 266 1082 304
rect 1136 272 1166 304
rect 898 222 908 256
rect 942 222 977 256
rect 898 206 977 222
rect 1028 256 1094 266
rect 1028 222 1044 256
rect 1078 222 1094 256
rect 1028 212 1094 222
rect 1136 256 1190 272
rect 1136 222 1146 256
rect 1180 222 1190 256
rect 1136 206 1190 222
rect 2199 382 2229 408
rect 2283 382 2313 408
rect 2471 388 2501 414
rect 729 66 759 106
rect 826 104 891 127
rect 826 97 847 104
rect 837 70 847 97
rect 881 70 891 104
rect 837 54 891 70
rect 837 22 867 54
rect 934 22 964 206
rect 1136 170 1166 206
rect 1029 140 1166 170
rect 1280 154 1310 220
rect 1417 188 1447 220
rect 1501 188 1531 220
rect 1029 10 1059 140
rect 1233 138 1310 154
rect 1233 104 1243 138
rect 1277 124 1310 138
rect 1361 172 1451 188
rect 1361 138 1371 172
rect 1405 138 1451 172
rect 1277 104 1287 124
rect 1361 122 1451 138
rect 1501 172 1567 188
rect 1501 138 1523 172
rect 1557 138 1567 172
rect 1501 122 1567 138
rect 1101 82 1155 98
rect 1101 48 1111 82
rect 1145 48 1155 82
rect 1233 88 1287 104
rect 1233 66 1263 88
rect 1421 66 1451 122
rect 1505 66 1535 122
rect 1609 120 1639 304
rect 1715 272 1745 304
rect 1681 256 1745 272
rect 1835 266 1865 304
rect 1681 222 1691 256
rect 1725 222 1745 256
rect 1681 206 1745 222
rect 1811 256 1877 266
rect 1811 222 1827 256
rect 1861 222 1877 256
rect 1811 212 1877 222
rect 1609 104 1669 120
rect 1609 84 1625 104
rect 1601 70 1625 84
rect 1659 70 1669 104
rect 1101 32 1155 48
rect 1113 10 1143 32
rect 1601 54 1669 70
rect 1601 22 1631 54
rect 1715 22 1745 206
rect 1919 170 1949 304
rect 1811 140 1949 170
rect 2011 158 2041 304
rect 2199 165 2229 254
rect 2283 239 2313 254
rect 2283 209 2347 239
rect 2317 171 2347 209
rect 2566 372 2596 398
rect 2754 388 2784 414
rect 3040 388 3070 414
rect 3112 388 3142 414
rect 3218 388 3248 414
rect 3339 388 3369 414
rect 3444 388 3474 414
rect 3528 388 3558 414
rect 3672 388 3702 414
rect 3809 388 3839 414
rect 3893 388 3923 414
rect 4001 388 4031 422
rect 4107 388 4137 414
rect 4227 388 4257 414
rect 4311 388 4341 414
rect 4403 388 4433 414
rect 2566 228 2596 244
rect 2566 198 2621 228
rect 1999 142 2053 158
rect 1811 110 1841 140
rect 1787 94 1841 110
rect 1999 108 2009 142
rect 2043 108 2053 142
rect 1787 60 1797 94
rect 1831 60 1841 94
rect 1787 44 1841 60
rect 1811 10 1841 44
rect 1883 82 1946 98
rect 1999 92 2053 108
rect 2199 155 2275 165
rect 2199 121 2225 155
rect 2259 121 2275 155
rect 2199 111 2275 121
rect 2317 155 2371 171
rect 2471 156 2501 188
rect 2317 121 2327 155
rect 2361 121 2371 155
rect 1883 48 1893 82
rect 1927 48 1946 82
rect 1883 32 1946 48
rect 1916 10 1946 32
rect 2011 22 2041 92
rect 2199 22 2229 111
rect 2317 105 2371 121
rect 2470 140 2529 156
rect 2470 106 2485 140
rect 2519 106 2529 140
rect 2317 67 2347 105
rect 2470 90 2529 106
rect 2591 150 2621 198
rect 2851 320 2881 346
rect 2754 156 2784 188
rect 2851 160 2881 192
rect 3040 188 3070 220
rect 2986 172 3070 188
rect 2749 150 2803 156
rect 2591 140 2803 150
rect 2591 106 2759 140
rect 2793 106 2803 140
rect 2591 96 2803 106
rect 2471 68 2501 90
rect 2283 37 2347 67
rect 2283 22 2313 37
rect 2591 67 2621 96
rect 2754 90 2803 96
rect 2849 144 2931 160
rect 2849 110 2887 144
rect 2921 110 2931 144
rect 2986 138 2996 172
rect 3030 138 3070 172
rect 2986 122 3070 138
rect 3112 172 3142 220
rect 3112 156 3176 172
rect 3112 122 3132 156
rect 3166 122 3176 156
rect 2849 94 2931 110
rect 2754 68 2784 90
rect 2566 37 2621 67
rect 2566 22 2596 37
rect 2849 22 2879 94
rect 3037 66 3067 122
rect 3112 106 3176 122
rect 3218 127 3248 304
rect 3339 272 3369 304
rect 3290 256 3369 272
rect 3444 266 3474 304
rect 3528 272 3558 304
rect 3290 222 3300 256
rect 3334 222 3369 256
rect 3290 206 3369 222
rect 3420 256 3486 266
rect 3420 222 3436 256
rect 3470 222 3486 256
rect 3420 212 3486 222
rect 3528 256 3582 272
rect 3528 222 3538 256
rect 3572 222 3582 256
rect 3528 206 3582 222
rect 4591 382 4621 408
rect 4675 382 4705 408
rect 4863 388 4893 414
rect 3121 66 3151 106
rect 3218 104 3283 127
rect 3218 97 3239 104
rect 3229 70 3239 97
rect 3273 70 3283 104
rect 3229 54 3283 70
rect 3229 22 3259 54
rect 3326 22 3356 206
rect 3528 170 3558 206
rect 3421 140 3558 170
rect 3672 154 3702 220
rect 3809 188 3839 220
rect 3893 188 3923 220
rect 3421 10 3451 140
rect 3625 138 3702 154
rect 3625 104 3635 138
rect 3669 124 3702 138
rect 3753 172 3843 188
rect 3753 138 3763 172
rect 3797 138 3843 172
rect 3669 104 3679 124
rect 3753 122 3843 138
rect 3893 172 3959 188
rect 3893 138 3915 172
rect 3949 138 3959 172
rect 3893 122 3959 138
rect 3493 82 3547 98
rect 3493 48 3503 82
rect 3537 48 3547 82
rect 3625 88 3679 104
rect 3625 66 3655 88
rect 3813 66 3843 122
rect 3897 66 3927 122
rect 4001 120 4031 304
rect 4107 272 4137 304
rect 4073 256 4137 272
rect 4227 266 4257 304
rect 4073 222 4083 256
rect 4117 222 4137 256
rect 4073 206 4137 222
rect 4203 256 4269 266
rect 4203 222 4219 256
rect 4253 222 4269 256
rect 4203 212 4269 222
rect 4001 104 4061 120
rect 4001 84 4017 104
rect 3993 70 4017 84
rect 4051 70 4061 104
rect 3493 32 3547 48
rect 3505 10 3535 32
rect 3993 54 4061 70
rect 3993 22 4023 54
rect 4107 22 4137 206
rect 4311 170 4341 304
rect 4203 140 4341 170
rect 4403 158 4433 304
rect 4591 165 4621 254
rect 4675 239 4705 254
rect 4675 209 4739 239
rect 4709 171 4739 209
rect 4958 372 4988 398
rect 5146 388 5176 414
rect 5432 388 5462 414
rect 5504 388 5534 414
rect 5610 388 5640 414
rect 5731 388 5761 414
rect 5836 388 5866 414
rect 5920 388 5950 414
rect 6064 388 6094 414
rect 6201 388 6231 414
rect 6285 388 6315 414
rect 6393 388 6423 422
rect 6499 388 6529 414
rect 6619 388 6649 414
rect 6703 388 6733 414
rect 6795 388 6825 414
rect 4958 228 4988 244
rect 4958 198 5013 228
rect 4391 142 4445 158
rect 4203 110 4233 140
rect 4179 94 4233 110
rect 4391 108 4401 142
rect 4435 108 4445 142
rect 4179 60 4189 94
rect 4223 60 4233 94
rect 4179 44 4233 60
rect 4203 10 4233 44
rect 4275 82 4338 98
rect 4391 92 4445 108
rect 4591 155 4667 165
rect 4591 121 4617 155
rect 4651 121 4667 155
rect 4591 111 4667 121
rect 4709 155 4763 171
rect 4863 156 4893 188
rect 4709 121 4719 155
rect 4753 121 4763 155
rect 4275 48 4285 82
rect 4319 48 4338 82
rect 4275 32 4338 48
rect 4308 10 4338 32
rect 4403 22 4433 92
rect 4591 22 4621 111
rect 4709 105 4763 121
rect 4862 140 4921 156
rect 4862 106 4877 140
rect 4911 106 4921 140
rect 4709 67 4739 105
rect 4862 90 4921 106
rect 4983 150 5013 198
rect 5243 320 5273 346
rect 5146 156 5176 188
rect 5243 160 5273 192
rect 5432 188 5462 220
rect 5378 172 5462 188
rect 5141 150 5195 156
rect 4983 140 5195 150
rect 4983 106 5151 140
rect 5185 106 5195 140
rect 4983 96 5195 106
rect 4863 68 4893 90
rect 4675 37 4739 67
rect 4675 22 4705 37
rect 4983 67 5013 96
rect 5146 90 5195 96
rect 5241 144 5323 160
rect 5241 110 5279 144
rect 5313 110 5323 144
rect 5378 138 5388 172
rect 5422 138 5462 172
rect 5378 122 5462 138
rect 5504 172 5534 220
rect 5504 156 5568 172
rect 5504 122 5524 156
rect 5558 122 5568 156
rect 5241 94 5323 110
rect 5146 68 5176 90
rect 4958 37 5013 67
rect 4958 22 4988 37
rect 5241 22 5271 94
rect 5429 66 5459 122
rect 5504 106 5568 122
rect 5610 127 5640 304
rect 5731 272 5761 304
rect 5682 256 5761 272
rect 5836 266 5866 304
rect 5920 272 5950 304
rect 5682 222 5692 256
rect 5726 222 5761 256
rect 5682 206 5761 222
rect 5812 256 5878 266
rect 5812 222 5828 256
rect 5862 222 5878 256
rect 5812 212 5878 222
rect 5920 256 5974 272
rect 5920 222 5930 256
rect 5964 222 5974 256
rect 5920 206 5974 222
rect 6983 382 7013 408
rect 7067 382 7097 408
rect 7255 388 7285 414
rect 5513 66 5543 106
rect 5610 104 5675 127
rect 5610 97 5631 104
rect 5621 70 5631 97
rect 5665 70 5675 104
rect 5621 54 5675 70
rect 5621 22 5651 54
rect 5718 22 5748 206
rect 5920 170 5950 206
rect 5813 140 5950 170
rect 6064 154 6094 220
rect 6201 188 6231 220
rect 6285 188 6315 220
rect 5813 10 5843 140
rect 6017 138 6094 154
rect 6017 104 6027 138
rect 6061 124 6094 138
rect 6145 172 6235 188
rect 6145 138 6155 172
rect 6189 138 6235 172
rect 6061 104 6071 124
rect 6145 122 6235 138
rect 6285 172 6351 188
rect 6285 138 6307 172
rect 6341 138 6351 172
rect 6285 122 6351 138
rect 5885 82 5939 98
rect 5885 48 5895 82
rect 5929 48 5939 82
rect 6017 88 6071 104
rect 6017 66 6047 88
rect 6205 66 6235 122
rect 6289 66 6319 122
rect 6393 120 6423 304
rect 6499 272 6529 304
rect 6465 256 6529 272
rect 6619 266 6649 304
rect 6465 222 6475 256
rect 6509 222 6529 256
rect 6465 206 6529 222
rect 6595 256 6661 266
rect 6595 222 6611 256
rect 6645 222 6661 256
rect 6595 212 6661 222
rect 6393 104 6453 120
rect 6393 84 6409 104
rect 6385 70 6409 84
rect 6443 70 6453 104
rect 5885 32 5939 48
rect 5897 10 5927 32
rect 6385 54 6453 70
rect 6385 22 6415 54
rect 6499 22 6529 206
rect 6703 170 6733 304
rect 6595 140 6733 170
rect 6795 158 6825 304
rect 6983 165 7013 254
rect 7067 239 7097 254
rect 7067 209 7131 239
rect 7101 171 7131 209
rect 7350 372 7380 398
rect 7538 388 7568 414
rect 7824 388 7854 414
rect 7896 388 7926 414
rect 8002 388 8032 414
rect 8123 388 8153 414
rect 8228 388 8258 414
rect 8312 388 8342 414
rect 8456 388 8486 414
rect 8593 388 8623 414
rect 8677 388 8707 414
rect 8785 388 8815 422
rect 8891 388 8921 414
rect 9011 388 9041 414
rect 9095 388 9125 414
rect 9187 388 9217 414
rect 7350 228 7380 244
rect 7350 198 7405 228
rect 6783 142 6837 158
rect 6595 110 6625 140
rect 6571 94 6625 110
rect 6783 108 6793 142
rect 6827 108 6837 142
rect 6571 60 6581 94
rect 6615 60 6625 94
rect 6571 44 6625 60
rect 6595 10 6625 44
rect 6667 82 6730 98
rect 6783 92 6837 108
rect 6983 155 7059 165
rect 6983 121 7009 155
rect 7043 121 7059 155
rect 6983 111 7059 121
rect 7101 155 7155 171
rect 7255 156 7285 188
rect 7101 121 7111 155
rect 7145 121 7155 155
rect 6667 48 6677 82
rect 6711 48 6730 82
rect 6667 32 6730 48
rect 6700 10 6730 32
rect 6795 22 6825 92
rect 6983 22 7013 111
rect 7101 105 7155 121
rect 7254 140 7313 156
rect 7254 106 7269 140
rect 7303 106 7313 140
rect 7101 67 7131 105
rect 7254 90 7313 106
rect 7375 150 7405 198
rect 7635 320 7665 346
rect 7538 156 7568 188
rect 7635 160 7665 192
rect 7824 188 7854 220
rect 7770 172 7854 188
rect 7533 150 7587 156
rect 7375 140 7587 150
rect 7375 106 7543 140
rect 7577 106 7587 140
rect 7375 96 7587 106
rect 7255 68 7285 90
rect 7067 37 7131 67
rect 7067 22 7097 37
rect 7375 67 7405 96
rect 7538 90 7587 96
rect 7633 144 7715 160
rect 7633 110 7671 144
rect 7705 110 7715 144
rect 7770 138 7780 172
rect 7814 138 7854 172
rect 7770 122 7854 138
rect 7896 172 7926 220
rect 7896 156 7960 172
rect 7896 122 7916 156
rect 7950 122 7960 156
rect 7633 94 7715 110
rect 7538 68 7568 90
rect 7350 37 7405 67
rect 7350 22 7380 37
rect 7633 22 7663 94
rect 7821 66 7851 122
rect 7896 106 7960 122
rect 8002 127 8032 304
rect 8123 272 8153 304
rect 8074 256 8153 272
rect 8228 266 8258 304
rect 8312 272 8342 304
rect 8074 222 8084 256
rect 8118 222 8153 256
rect 8074 206 8153 222
rect 8204 256 8270 266
rect 8204 222 8220 256
rect 8254 222 8270 256
rect 8204 212 8270 222
rect 8312 256 8366 272
rect 8312 222 8322 256
rect 8356 222 8366 256
rect 8312 206 8366 222
rect 9375 382 9405 408
rect 9459 382 9489 408
rect 9647 388 9677 414
rect 7905 66 7935 106
rect 8002 104 8067 127
rect 8002 97 8023 104
rect 8013 70 8023 97
rect 8057 70 8067 104
rect 8013 54 8067 70
rect 8013 22 8043 54
rect 8110 22 8140 206
rect 8312 170 8342 206
rect 8205 140 8342 170
rect 8456 154 8486 220
rect 8593 188 8623 220
rect 8677 188 8707 220
rect 8205 10 8235 140
rect 8409 138 8486 154
rect 8409 104 8419 138
rect 8453 124 8486 138
rect 8537 172 8627 188
rect 8537 138 8547 172
rect 8581 138 8627 172
rect 8453 104 8463 124
rect 8537 122 8627 138
rect 8677 172 8743 188
rect 8677 138 8699 172
rect 8733 138 8743 172
rect 8677 122 8743 138
rect 8277 82 8331 98
rect 8277 48 8287 82
rect 8321 48 8331 82
rect 8409 88 8463 104
rect 8409 66 8439 88
rect 8597 66 8627 122
rect 8681 66 8711 122
rect 8785 120 8815 304
rect 8891 272 8921 304
rect 8857 256 8921 272
rect 9011 266 9041 304
rect 8857 222 8867 256
rect 8901 222 8921 256
rect 8857 206 8921 222
rect 8987 256 9053 266
rect 8987 222 9003 256
rect 9037 222 9053 256
rect 8987 212 9053 222
rect 8785 104 8845 120
rect 8785 84 8801 104
rect 8777 70 8801 84
rect 8835 70 8845 104
rect 8277 32 8331 48
rect 8289 10 8319 32
rect 8777 54 8845 70
rect 8777 22 8807 54
rect 8891 22 8921 206
rect 9095 170 9125 304
rect 8987 140 9125 170
rect 9187 158 9217 304
rect 9375 165 9405 254
rect 9459 239 9489 254
rect 9459 209 9523 239
rect 9493 171 9523 209
rect 9742 372 9772 398
rect 9930 388 9960 414
rect 10216 388 10246 414
rect 10288 388 10318 414
rect 10394 388 10424 414
rect 10515 388 10545 414
rect 10620 388 10650 414
rect 10704 388 10734 414
rect 10848 388 10878 414
rect 10985 388 11015 414
rect 11069 388 11099 414
rect 11177 388 11207 422
rect 11283 388 11313 414
rect 11403 388 11433 414
rect 11487 388 11517 414
rect 11579 388 11609 414
rect 9742 228 9772 244
rect 9742 198 9797 228
rect 9175 142 9229 158
rect 8987 110 9017 140
rect 8963 94 9017 110
rect 9175 108 9185 142
rect 9219 108 9229 142
rect 8963 60 8973 94
rect 9007 60 9017 94
rect 8963 44 9017 60
rect 8987 10 9017 44
rect 9059 82 9122 98
rect 9175 92 9229 108
rect 9375 155 9451 165
rect 9375 121 9401 155
rect 9435 121 9451 155
rect 9375 111 9451 121
rect 9493 155 9547 171
rect 9647 156 9677 188
rect 9493 121 9503 155
rect 9537 121 9547 155
rect 9059 48 9069 82
rect 9103 48 9122 82
rect 9059 32 9122 48
rect 9092 10 9122 32
rect 9187 22 9217 92
rect 9375 22 9405 111
rect 9493 105 9547 121
rect 9646 140 9705 156
rect 9646 106 9661 140
rect 9695 106 9705 140
rect 9493 67 9523 105
rect 9646 90 9705 106
rect 9767 150 9797 198
rect 10027 320 10057 346
rect 9930 156 9960 188
rect 10027 160 10057 192
rect 10216 188 10246 220
rect 10162 172 10246 188
rect 9925 150 9979 156
rect 9767 140 9979 150
rect 9767 106 9935 140
rect 9969 106 9979 140
rect 9767 96 9979 106
rect 9647 68 9677 90
rect 9459 37 9523 67
rect 9459 22 9489 37
rect 9767 67 9797 96
rect 9930 90 9979 96
rect 10025 144 10107 160
rect 10025 110 10063 144
rect 10097 110 10107 144
rect 10162 138 10172 172
rect 10206 138 10246 172
rect 10162 122 10246 138
rect 10288 172 10318 220
rect 10288 156 10352 172
rect 10288 122 10308 156
rect 10342 122 10352 156
rect 10025 94 10107 110
rect 9930 68 9960 90
rect 9742 37 9797 67
rect 9742 22 9772 37
rect 10025 22 10055 94
rect 10213 66 10243 122
rect 10288 106 10352 122
rect 10394 127 10424 304
rect 10515 272 10545 304
rect 10466 256 10545 272
rect 10620 266 10650 304
rect 10704 272 10734 304
rect 10466 222 10476 256
rect 10510 222 10545 256
rect 10466 206 10545 222
rect 10596 256 10662 266
rect 10596 222 10612 256
rect 10646 222 10662 256
rect 10596 212 10662 222
rect 10704 256 10758 272
rect 10704 222 10714 256
rect 10748 222 10758 256
rect 10704 206 10758 222
rect 11767 382 11797 408
rect 11851 382 11881 408
rect 12039 388 12069 414
rect 10297 66 10327 106
rect 10394 104 10459 127
rect 10394 97 10415 104
rect 10405 70 10415 97
rect 10449 70 10459 104
rect 10405 54 10459 70
rect 10405 22 10435 54
rect 10502 22 10532 206
rect 10704 170 10734 206
rect 10597 140 10734 170
rect 10848 154 10878 220
rect 10985 188 11015 220
rect 11069 188 11099 220
rect 10597 10 10627 140
rect 10801 138 10878 154
rect 10801 104 10811 138
rect 10845 124 10878 138
rect 10929 172 11019 188
rect 10929 138 10939 172
rect 10973 138 11019 172
rect 10845 104 10855 124
rect 10929 122 11019 138
rect 11069 172 11135 188
rect 11069 138 11091 172
rect 11125 138 11135 172
rect 11069 122 11135 138
rect 10669 82 10723 98
rect 10669 48 10679 82
rect 10713 48 10723 82
rect 10801 88 10855 104
rect 10801 66 10831 88
rect 10989 66 11019 122
rect 11073 66 11103 122
rect 11177 120 11207 304
rect 11283 272 11313 304
rect 11249 256 11313 272
rect 11403 266 11433 304
rect 11249 222 11259 256
rect 11293 222 11313 256
rect 11249 206 11313 222
rect 11379 256 11445 266
rect 11379 222 11395 256
rect 11429 222 11445 256
rect 11379 212 11445 222
rect 11177 104 11237 120
rect 11177 84 11193 104
rect 11169 70 11193 84
rect 11227 70 11237 104
rect 10669 32 10723 48
rect 10681 10 10711 32
rect 11169 54 11237 70
rect 11169 22 11199 54
rect 11283 22 11313 206
rect 11487 170 11517 304
rect 11379 140 11517 170
rect 11579 158 11609 304
rect 11767 165 11797 254
rect 11851 239 11881 254
rect 11851 209 11915 239
rect 11885 171 11915 209
rect 12134 372 12164 398
rect 12322 388 12352 414
rect 12608 388 12638 414
rect 12680 388 12710 414
rect 12786 388 12816 414
rect 12907 388 12937 414
rect 13012 388 13042 414
rect 13096 388 13126 414
rect 13240 388 13270 414
rect 13377 388 13407 414
rect 13461 388 13491 414
rect 13569 388 13599 422
rect 15943 419 16009 435
rect 13675 388 13705 414
rect 13795 388 13825 414
rect 13879 388 13909 414
rect 13971 388 14001 414
rect 12134 228 12164 244
rect 12134 198 12189 228
rect 11567 142 11621 158
rect 11379 110 11409 140
rect 11355 94 11409 110
rect 11567 108 11577 142
rect 11611 108 11621 142
rect 11355 60 11365 94
rect 11399 60 11409 94
rect 11355 44 11409 60
rect 11379 10 11409 44
rect 11451 82 11514 98
rect 11567 92 11621 108
rect 11767 155 11843 165
rect 11767 121 11793 155
rect 11827 121 11843 155
rect 11767 111 11843 121
rect 11885 155 11939 171
rect 12039 156 12069 188
rect 11885 121 11895 155
rect 11929 121 11939 155
rect 11451 48 11461 82
rect 11495 48 11514 82
rect 11451 32 11514 48
rect 11484 10 11514 32
rect 11579 22 11609 92
rect 11767 22 11797 111
rect 11885 105 11939 121
rect 12038 140 12097 156
rect 12038 106 12053 140
rect 12087 106 12097 140
rect 11885 67 11915 105
rect 12038 90 12097 106
rect 12159 150 12189 198
rect 12419 320 12449 346
rect 12322 156 12352 188
rect 12419 160 12449 192
rect 12608 188 12638 220
rect 12554 172 12638 188
rect 12317 150 12371 156
rect 12159 140 12371 150
rect 12159 106 12327 140
rect 12361 106 12371 140
rect 12159 96 12371 106
rect 12039 68 12069 90
rect 11851 37 11915 67
rect 11851 22 11881 37
rect 12159 67 12189 96
rect 12322 90 12371 96
rect 12417 144 12499 160
rect 12417 110 12455 144
rect 12489 110 12499 144
rect 12554 138 12564 172
rect 12598 138 12638 172
rect 12554 122 12638 138
rect 12680 172 12710 220
rect 12680 156 12744 172
rect 12680 122 12700 156
rect 12734 122 12744 156
rect 12417 94 12499 110
rect 12322 68 12352 90
rect 12134 37 12189 67
rect 12134 22 12164 37
rect 12417 22 12447 94
rect 12605 66 12635 122
rect 12680 106 12744 122
rect 12786 127 12816 304
rect 12907 272 12937 304
rect 12858 256 12937 272
rect 13012 266 13042 304
rect 13096 272 13126 304
rect 12858 222 12868 256
rect 12902 222 12937 256
rect 12858 206 12937 222
rect 12988 256 13054 266
rect 12988 222 13004 256
rect 13038 222 13054 256
rect 12988 212 13054 222
rect 13096 256 13150 272
rect 13096 222 13106 256
rect 13140 222 13150 256
rect 13096 206 13150 222
rect 14159 382 14189 408
rect 14243 382 14273 408
rect 14431 388 14461 414
rect 12689 66 12719 106
rect 12786 104 12851 127
rect 12786 97 12807 104
rect 12797 70 12807 97
rect 12841 70 12851 104
rect 12797 54 12851 70
rect 12797 22 12827 54
rect 12894 22 12924 206
rect 13096 170 13126 206
rect 12989 140 13126 170
rect 13240 154 13270 220
rect 13377 188 13407 220
rect 13461 188 13491 220
rect 12989 10 13019 140
rect 13193 138 13270 154
rect 13193 104 13203 138
rect 13237 124 13270 138
rect 13321 172 13411 188
rect 13321 138 13331 172
rect 13365 138 13411 172
rect 13237 104 13247 124
rect 13321 122 13411 138
rect 13461 172 13527 188
rect 13461 138 13483 172
rect 13517 138 13527 172
rect 13461 122 13527 138
rect 13061 82 13115 98
rect 13061 48 13071 82
rect 13105 48 13115 82
rect 13193 88 13247 104
rect 13193 66 13223 88
rect 13381 66 13411 122
rect 13465 66 13495 122
rect 13569 120 13599 304
rect 13675 272 13705 304
rect 13641 256 13705 272
rect 13795 266 13825 304
rect 13641 222 13651 256
rect 13685 222 13705 256
rect 13641 206 13705 222
rect 13771 256 13837 266
rect 13771 222 13787 256
rect 13821 222 13837 256
rect 13771 212 13837 222
rect 13569 104 13629 120
rect 13569 84 13585 104
rect 13561 70 13585 84
rect 13619 70 13629 104
rect 13061 32 13115 48
rect 13073 10 13103 32
rect 13561 54 13629 70
rect 13561 22 13591 54
rect 13675 22 13705 206
rect 13879 170 13909 304
rect 13771 140 13909 170
rect 13971 158 14001 304
rect 14159 165 14189 254
rect 14243 239 14273 254
rect 14243 209 14307 239
rect 14277 171 14307 209
rect 14526 372 14556 398
rect 14714 388 14744 414
rect 15000 388 15030 414
rect 15072 388 15102 414
rect 15178 388 15208 414
rect 15299 388 15329 414
rect 15404 388 15434 414
rect 15488 388 15518 414
rect 15632 388 15662 414
rect 15769 388 15799 414
rect 15853 388 15883 414
rect 15961 388 15991 419
rect 16067 388 16097 414
rect 16187 388 16217 414
rect 16271 388 16301 414
rect 16363 388 16393 414
rect 14526 228 14556 244
rect 14526 198 14581 228
rect 13959 142 14013 158
rect 13771 110 13801 140
rect 13747 94 13801 110
rect 13959 108 13969 142
rect 14003 108 14013 142
rect 13747 60 13757 94
rect 13791 60 13801 94
rect 13747 44 13801 60
rect 13771 10 13801 44
rect 13843 82 13906 98
rect 13959 92 14013 108
rect 14159 155 14235 165
rect 14159 121 14185 155
rect 14219 121 14235 155
rect 14159 111 14235 121
rect 14277 155 14331 171
rect 14431 156 14461 188
rect 14277 121 14287 155
rect 14321 121 14331 155
rect 13843 48 13853 82
rect 13887 48 13906 82
rect 13843 32 13906 48
rect 13876 10 13906 32
rect 13971 22 14001 92
rect 14159 22 14189 111
rect 14277 105 14331 121
rect 14430 140 14489 156
rect 14430 106 14445 140
rect 14479 106 14489 140
rect 14277 67 14307 105
rect 14430 90 14489 106
rect 14551 150 14581 198
rect 14811 320 14841 346
rect 14714 156 14744 188
rect 14811 160 14841 192
rect 15000 188 15030 220
rect 14946 172 15030 188
rect 14709 150 14763 156
rect 14551 140 14763 150
rect 14551 106 14719 140
rect 14753 106 14763 140
rect 14551 96 14763 106
rect 14431 68 14461 90
rect 14243 37 14307 67
rect 14243 22 14273 37
rect 14551 67 14581 96
rect 14714 90 14763 96
rect 14809 144 14891 160
rect 14809 110 14847 144
rect 14881 110 14891 144
rect 14946 138 14956 172
rect 14990 138 15030 172
rect 14946 122 15030 138
rect 15072 172 15102 220
rect 15072 156 15136 172
rect 15072 122 15092 156
rect 15126 122 15136 156
rect 14809 94 14891 110
rect 14714 68 14744 90
rect 14526 37 14581 67
rect 14526 22 14556 37
rect 14809 22 14839 94
rect 14997 66 15027 122
rect 15072 106 15136 122
rect 15178 127 15208 304
rect 15299 272 15329 304
rect 15250 256 15329 272
rect 15404 266 15434 304
rect 15488 272 15518 304
rect 15250 222 15260 256
rect 15294 222 15329 256
rect 15250 206 15329 222
rect 15380 256 15446 266
rect 15380 222 15396 256
rect 15430 222 15446 256
rect 15380 212 15446 222
rect 15488 256 15542 272
rect 15488 222 15498 256
rect 15532 222 15542 256
rect 15488 206 15542 222
rect 16551 382 16581 408
rect 16635 382 16665 408
rect 15081 66 15111 106
rect 15178 104 15243 127
rect 15178 97 15199 104
rect 15189 70 15199 97
rect 15233 70 15243 104
rect 15189 54 15243 70
rect 15189 22 15219 54
rect 15286 22 15316 206
rect 15488 170 15518 206
rect 15381 140 15518 170
rect 15632 154 15662 220
rect 15769 188 15799 220
rect 15853 188 15883 220
rect 15381 10 15411 140
rect 15585 138 15662 154
rect 15585 104 15595 138
rect 15629 124 15662 138
rect 15713 172 15803 188
rect 15713 138 15723 172
rect 15757 138 15803 172
rect 15629 104 15639 124
rect 15713 122 15803 138
rect 15853 172 15919 188
rect 15853 138 15875 172
rect 15909 138 15919 172
rect 15853 122 15919 138
rect 15453 82 15507 98
rect 15453 48 15463 82
rect 15497 48 15507 82
rect 15585 88 15639 104
rect 15585 66 15615 88
rect 15773 66 15803 122
rect 15857 66 15887 122
rect 15961 120 15991 304
rect 16067 272 16097 304
rect 16033 256 16097 272
rect 16187 266 16217 304
rect 16033 222 16043 256
rect 16077 222 16097 256
rect 16033 206 16097 222
rect 16163 256 16229 266
rect 16163 222 16179 256
rect 16213 222 16229 256
rect 16163 212 16229 222
rect 15961 104 16021 120
rect 15961 84 15977 104
rect 15953 70 15977 84
rect 16011 70 16021 104
rect 15453 32 15507 48
rect 15465 10 15495 32
rect 15953 54 16021 70
rect 15953 22 15983 54
rect 16067 22 16097 206
rect 16271 170 16301 304
rect 16163 140 16301 170
rect 16363 158 16393 304
rect 16551 165 16581 254
rect 16635 239 16665 254
rect 16635 209 16699 239
rect 16669 171 16699 209
rect 16351 142 16405 158
rect 16163 110 16193 140
rect 16139 94 16193 110
rect 16351 108 16361 142
rect 16395 108 16405 142
rect 16139 60 16149 94
rect 16183 60 16193 94
rect 16139 44 16193 60
rect 16163 10 16193 44
rect 16235 82 16298 98
rect 16351 92 16405 108
rect 16551 155 16627 165
rect 16551 121 16577 155
rect 16611 121 16627 155
rect 16551 111 16627 121
rect 16669 155 16723 171
rect 16669 121 16679 155
rect 16713 121 16723 155
rect 16235 48 16245 82
rect 16279 48 16298 82
rect 16235 32 16298 48
rect 16268 10 16298 32
rect 16363 22 16393 92
rect 16551 22 16581 111
rect 16669 105 16723 121
rect 16669 67 16699 105
rect 16635 37 16699 67
rect 16635 22 16665 37
rect 79 -88 109 -62
rect 174 -88 204 -62
rect 362 -88 392 -62
rect 457 -88 487 -62
rect 645 -88 675 -62
rect 729 -88 759 -62
rect 837 -88 867 -62
rect 934 -88 964 -62
rect 1029 -88 1059 -62
rect 1113 -88 1143 -62
rect 1233 -88 1263 -62
rect 1421 -88 1451 -62
rect 1505 -88 1535 -62
rect 1601 -88 1631 -62
rect 1715 -88 1745 -62
rect 1811 -88 1841 -62
rect 1916 -88 1946 -62
rect 2011 -88 2041 -62
rect 2199 -88 2229 -62
rect 2283 -88 2313 -62
rect 2471 -88 2501 -62
rect 2566 -88 2596 -62
rect 2754 -88 2784 -62
rect 2849 -88 2879 -62
rect 3037 -88 3067 -62
rect 3121 -88 3151 -62
rect 3229 -88 3259 -62
rect 3326 -88 3356 -62
rect 3421 -88 3451 -62
rect 3505 -88 3535 -62
rect 3625 -88 3655 -62
rect 3813 -88 3843 -62
rect 3897 -88 3927 -62
rect 3993 -88 4023 -62
rect 4107 -88 4137 -62
rect 4203 -88 4233 -62
rect 4308 -88 4338 -62
rect 4403 -88 4433 -62
rect 4591 -88 4621 -62
rect 4675 -88 4705 -62
rect 4863 -88 4893 -62
rect 4958 -88 4988 -62
rect 5146 -88 5176 -62
rect 5241 -88 5271 -62
rect 5429 -88 5459 -62
rect 5513 -88 5543 -62
rect 5621 -88 5651 -62
rect 5718 -88 5748 -62
rect 5813 -88 5843 -62
rect 5897 -88 5927 -62
rect 6017 -88 6047 -62
rect 6205 -88 6235 -62
rect 6289 -88 6319 -62
rect 6385 -88 6415 -62
rect 6499 -88 6529 -62
rect 6595 -88 6625 -62
rect 6700 -88 6730 -62
rect 6795 -88 6825 -62
rect 6983 -88 7013 -62
rect 7067 -88 7097 -62
rect 7255 -88 7285 -62
rect 7350 -88 7380 -62
rect 7538 -88 7568 -62
rect 7633 -88 7663 -62
rect 7821 -88 7851 -62
rect 7905 -88 7935 -62
rect 8013 -88 8043 -62
rect 8110 -88 8140 -62
rect 8205 -88 8235 -62
rect 8289 -88 8319 -62
rect 8409 -88 8439 -62
rect 8597 -88 8627 -62
rect 8681 -88 8711 -62
rect 8777 -88 8807 -62
rect 8891 -88 8921 -62
rect 8987 -88 9017 -62
rect 9092 -88 9122 -62
rect 9187 -88 9217 -62
rect 9375 -88 9405 -62
rect 9459 -88 9489 -62
rect 9647 -88 9677 -62
rect 9742 -88 9772 -62
rect 9930 -88 9960 -62
rect 10025 -88 10055 -62
rect 10213 -88 10243 -62
rect 10297 -88 10327 -62
rect 10405 -88 10435 -62
rect 10502 -88 10532 -62
rect 10597 -88 10627 -62
rect 10681 -88 10711 -62
rect 10801 -88 10831 -62
rect 10989 -88 11019 -62
rect 11073 -88 11103 -62
rect 11169 -88 11199 -62
rect 11283 -88 11313 -62
rect 11379 -88 11409 -62
rect 11484 -88 11514 -62
rect 11579 -88 11609 -62
rect 11767 -88 11797 -62
rect 11851 -88 11881 -62
rect 12039 -88 12069 -62
rect 12134 -88 12164 -62
rect 12322 -88 12352 -62
rect 12417 -88 12447 -62
rect 12605 -88 12635 -62
rect 12689 -88 12719 -62
rect 12797 -88 12827 -62
rect 12894 -88 12924 -62
rect 12989 -88 13019 -62
rect 13073 -88 13103 -62
rect 13193 -88 13223 -62
rect 13381 -88 13411 -62
rect 13465 -88 13495 -62
rect 13561 -88 13591 -62
rect 13675 -88 13705 -62
rect 13771 -88 13801 -62
rect 13876 -88 13906 -62
rect 13971 -88 14001 -62
rect 14159 -88 14189 -62
rect 14243 -88 14273 -62
rect 14431 -88 14461 -62
rect 14526 -88 14556 -62
rect 14714 -88 14744 -62
rect 14809 -88 14839 -62
rect 14997 -88 15027 -62
rect 15081 -88 15111 -62
rect 15189 -88 15219 -62
rect 15286 -88 15316 -62
rect 15381 -88 15411 -62
rect 15465 -88 15495 -62
rect 15585 -88 15615 -62
rect 15773 -88 15803 -62
rect 15857 -88 15887 -62
rect 15953 -88 15983 -62
rect 16067 -88 16097 -62
rect 16163 -88 16193 -62
rect 16268 -88 16298 -62
rect 16363 -88 16393 -62
rect 16551 -88 16581 -62
rect 16635 -88 16665 -62
<< polycont >>
rect 39 2625 73 2659
rect 157 2638 191 2672
rect 322 2625 356 2659
rect 456 2625 490 2659
rect 933 2625 967 2659
rect 1001 2625 1035 2659
rect 1069 2625 1103 2659
rect 1137 2625 1171 2659
rect 1205 2625 1239 2659
rect 1273 2625 1307 2659
rect 1433 2625 1467 2659
rect 1501 2625 1535 2659
rect 1569 2625 1603 2659
rect 1637 2625 1671 2659
rect 1705 2625 1739 2659
rect 1773 2625 1807 2659
rect 1841 2625 1875 2659
rect 1909 2625 1943 2659
rect 1977 2625 2011 2659
rect 2045 2625 2079 2659
rect 2113 2625 2147 2659
rect 2181 2625 2215 2659
rect 2249 2625 2283 2659
rect 2317 2625 2351 2659
rect 2385 2625 2419 2659
rect 2453 2625 2487 2659
rect 2521 2625 2555 2659
rect 2589 2625 2623 2659
rect 2657 2625 2691 2659
rect 4423 2625 4457 2659
rect 4541 2638 4575 2672
rect 4706 2625 4740 2659
rect 4840 2625 4874 2659
rect 5317 2625 5351 2659
rect 5385 2625 5419 2659
rect 5453 2625 5487 2659
rect 5521 2625 5555 2659
rect 5589 2625 5623 2659
rect 5657 2625 5691 2659
rect 5817 2625 5851 2659
rect 5885 2625 5919 2659
rect 5953 2625 5987 2659
rect 6021 2625 6055 2659
rect 6089 2625 6123 2659
rect 6157 2625 6191 2659
rect 6225 2625 6259 2659
rect 6293 2625 6327 2659
rect 6361 2625 6395 2659
rect 6429 2625 6463 2659
rect 6497 2625 6531 2659
rect 6565 2625 6599 2659
rect 6633 2625 6667 2659
rect 6701 2625 6735 2659
rect 6769 2625 6803 2659
rect 6837 2625 6871 2659
rect 6905 2625 6939 2659
rect 6973 2625 7007 2659
rect 7041 2625 7075 2659
rect 86 1483 120 1517
rect 182 1483 216 1517
rect 491 1560 525 1594
rect 323 1447 357 1481
rect 659 1560 693 1594
rect 419 1447 453 1481
rect 581 1447 615 1481
rect 1569 1560 1603 1594
rect 1737 1560 1771 1594
rect 1647 1447 1681 1481
rect 1809 1447 1843 1481
rect 1905 1447 1939 1481
rect 2046 1483 2080 1517
rect 2142 1483 2176 1517
rect 2478 1483 2512 1517
rect 2574 1483 2608 1517
rect 2883 1560 2917 1594
rect 2715 1447 2749 1481
rect 3051 1560 3085 1594
rect 2811 1447 2845 1481
rect 2973 1447 3007 1481
rect 3961 1560 3995 1594
rect 4129 1560 4163 1594
rect 4039 1447 4073 1481
rect 4201 1447 4235 1481
rect 4297 1447 4331 1481
rect 4438 1483 4472 1517
rect 4534 1483 4568 1517
rect 4870 1483 4904 1517
rect 4966 1483 5000 1517
rect 5275 1560 5309 1594
rect 5107 1447 5141 1481
rect 5443 1560 5477 1594
rect 5203 1447 5237 1481
rect 5365 1447 5399 1481
rect 6351 1560 6385 1594
rect 6519 1560 6553 1594
rect 6429 1447 6463 1481
rect 6591 1447 6625 1481
rect 6687 1447 6721 1481
rect 6828 1483 6862 1517
rect 6924 1483 6958 1517
rect 7262 1483 7296 1517
rect 7358 1483 7392 1517
rect 7667 1560 7701 1594
rect 7499 1447 7533 1481
rect 7835 1560 7869 1594
rect 7595 1447 7629 1481
rect 7757 1447 7791 1481
rect 8745 1560 8779 1594
rect 8913 1560 8947 1594
rect 8823 1447 8857 1481
rect 8985 1447 9019 1481
rect 9081 1447 9115 1481
rect 9222 1483 9256 1517
rect 9318 1483 9352 1517
rect 9654 1483 9688 1517
rect 9750 1483 9784 1517
rect 10059 1560 10093 1594
rect 9891 1447 9925 1481
rect 10227 1560 10261 1594
rect 9987 1447 10021 1481
rect 10149 1447 10183 1481
rect 11137 1560 11171 1594
rect 11305 1560 11339 1594
rect 11215 1447 11249 1481
rect 11377 1447 11411 1481
rect 11473 1447 11507 1481
rect 11614 1483 11648 1517
rect 11710 1483 11744 1517
rect 12046 1483 12080 1517
rect 12142 1483 12176 1517
rect 12451 1560 12485 1594
rect 12283 1447 12317 1481
rect 12619 1560 12653 1594
rect 12379 1447 12413 1481
rect 12541 1447 12575 1481
rect 13527 1560 13561 1594
rect 13695 1560 13729 1594
rect 13605 1447 13639 1481
rect 13767 1447 13801 1481
rect 13863 1447 13897 1481
rect 14004 1483 14038 1517
rect 14100 1483 14134 1517
rect 14438 1483 14472 1517
rect 14534 1483 14568 1517
rect 14843 1560 14877 1594
rect 14675 1447 14709 1481
rect 15011 1560 15045 1594
rect 14771 1447 14805 1481
rect 14933 1447 14967 1481
rect 15921 1560 15955 1594
rect 16089 1560 16123 1594
rect 15999 1447 16033 1481
rect 16161 1447 16195 1481
rect 16257 1447 16291 1481
rect 16398 1483 16432 1517
rect 16494 1483 16528 1517
rect 1901 1124 1935 1158
rect 4293 1123 4327 1157
rect 31 810 65 844
rect 531 911 565 945
rect 667 911 701 945
rect 133 810 167 844
rect 349 797 383 831
rect 465 737 499 771
rect 561 749 595 783
rect 1212 911 1246 945
rect 835 827 869 861
rect 987 827 1021 861
rect 1314 911 1348 945
rect 1450 911 1484 945
rect 733 759 767 793
rect 1115 793 1149 827
rect 1247 737 1281 771
rect 6685 1123 6719 1157
rect 9077 1124 9111 1158
rect 11469 1124 11503 1158
rect 13861 1123 13895 1157
rect 1618 811 1652 845
rect 1754 827 1788 861
rect 1511 759 1545 793
rect 1863 799 1897 833
rect 1991 795 2025 829
rect 2265 795 2299 829
rect 2423 810 2457 844
rect 2923 911 2957 945
rect 3059 911 3093 945
rect 2525 810 2559 844
rect 2741 797 2775 831
rect 2857 737 2891 771
rect 2953 749 2987 783
rect 3604 911 3638 945
rect 3227 827 3261 861
rect 3379 827 3413 861
rect 3706 911 3740 945
rect 3842 911 3876 945
rect 3125 759 3159 793
rect 3507 793 3541 827
rect 3639 737 3673 771
rect 4010 811 4044 845
rect 4146 827 4180 861
rect 3903 759 3937 793
rect 4255 799 4289 833
rect 4383 795 4417 829
rect 4657 795 4691 829
rect 4815 810 4849 844
rect 5315 911 5349 945
rect 5451 911 5485 945
rect 4917 810 4951 844
rect 5133 797 5167 831
rect 5249 737 5283 771
rect 5345 749 5379 783
rect 5996 911 6030 945
rect 5619 827 5653 861
rect 5771 827 5805 861
rect 6098 911 6132 945
rect 6234 911 6268 945
rect 5517 759 5551 793
rect 5899 793 5933 827
rect 6031 737 6065 771
rect 6402 811 6436 845
rect 6538 827 6572 861
rect 6295 759 6329 793
rect 6647 799 6681 833
rect 6775 795 6809 829
rect 7049 795 7083 829
rect 7207 810 7241 844
rect 7707 911 7741 945
rect 7843 911 7877 945
rect 7309 810 7343 844
rect 7525 797 7559 831
rect 7641 737 7675 771
rect 7737 749 7771 783
rect 8388 911 8422 945
rect 8011 827 8045 861
rect 8163 827 8197 861
rect 8490 911 8524 945
rect 8626 911 8660 945
rect 7909 759 7943 793
rect 8291 793 8325 827
rect 8423 737 8457 771
rect 8794 811 8828 845
rect 8930 827 8964 861
rect 8687 759 8721 793
rect 9039 799 9073 833
rect 9167 795 9201 829
rect 9441 795 9475 829
rect 9599 810 9633 844
rect 10099 911 10133 945
rect 10235 911 10269 945
rect 9701 810 9735 844
rect 9917 797 9951 831
rect 10033 737 10067 771
rect 10129 749 10163 783
rect 10780 911 10814 945
rect 10403 827 10437 861
rect 10555 827 10589 861
rect 10882 911 10916 945
rect 11018 911 11052 945
rect 10301 759 10335 793
rect 10683 793 10717 827
rect 10815 737 10849 771
rect 16253 1123 16287 1157
rect 11186 811 11220 845
rect 11322 827 11356 861
rect 11079 759 11113 793
rect 11431 799 11465 833
rect 11559 795 11593 829
rect 11833 795 11867 829
rect 11991 810 12025 844
rect 12491 911 12525 945
rect 12627 911 12661 945
rect 12093 810 12127 844
rect 12309 797 12343 831
rect 12425 737 12459 771
rect 12521 749 12555 783
rect 13172 911 13206 945
rect 12795 827 12829 861
rect 12947 827 12981 861
rect 13274 911 13308 945
rect 13410 911 13444 945
rect 12693 759 12727 793
rect 13075 793 13109 827
rect 13207 737 13241 771
rect 13578 811 13612 845
rect 13714 827 13748 861
rect 13471 759 13505 793
rect 13823 799 13857 833
rect 13951 795 13985 829
rect 14225 795 14259 829
rect 14383 810 14417 844
rect 14883 911 14917 945
rect 15019 911 15053 945
rect 14485 810 14519 844
rect 14701 797 14735 831
rect 14817 737 14851 771
rect 14913 749 14947 783
rect 15564 911 15598 945
rect 15187 827 15221 861
rect 15339 827 15373 861
rect 15666 911 15700 945
rect 15802 911 15836 945
rect 15085 759 15119 793
rect 15467 793 15501 827
rect 15599 737 15633 771
rect 15970 811 16004 845
rect 16106 827 16140 861
rect 15863 759 15897 793
rect 16215 799 16249 833
rect 16343 795 16377 829
rect 16617 795 16651 829
rect 1607 438 1641 472
rect 3999 438 4033 472
rect 6391 438 6425 472
rect 8783 438 8817 472
rect 11175 438 11209 472
rect 13567 438 13601 472
rect 15959 435 15993 469
rect 93 106 127 140
rect 367 106 401 140
rect 495 110 529 144
rect 604 138 638 172
rect 740 122 774 156
rect 908 222 942 256
rect 1044 222 1078 256
rect 1146 222 1180 256
rect 847 70 881 104
rect 1243 104 1277 138
rect 1371 138 1405 172
rect 1523 138 1557 172
rect 1111 48 1145 82
rect 1691 222 1725 256
rect 1827 222 1861 256
rect 1625 70 1659 104
rect 2009 108 2043 142
rect 1797 60 1831 94
rect 2225 121 2259 155
rect 2327 121 2361 155
rect 1893 48 1927 82
rect 2485 106 2519 140
rect 2759 106 2793 140
rect 2887 110 2921 144
rect 2996 138 3030 172
rect 3132 122 3166 156
rect 3300 222 3334 256
rect 3436 222 3470 256
rect 3538 222 3572 256
rect 3239 70 3273 104
rect 3635 104 3669 138
rect 3763 138 3797 172
rect 3915 138 3949 172
rect 3503 48 3537 82
rect 4083 222 4117 256
rect 4219 222 4253 256
rect 4017 70 4051 104
rect 4401 108 4435 142
rect 4189 60 4223 94
rect 4617 121 4651 155
rect 4719 121 4753 155
rect 4285 48 4319 82
rect 4877 106 4911 140
rect 5151 106 5185 140
rect 5279 110 5313 144
rect 5388 138 5422 172
rect 5524 122 5558 156
rect 5692 222 5726 256
rect 5828 222 5862 256
rect 5930 222 5964 256
rect 5631 70 5665 104
rect 6027 104 6061 138
rect 6155 138 6189 172
rect 6307 138 6341 172
rect 5895 48 5929 82
rect 6475 222 6509 256
rect 6611 222 6645 256
rect 6409 70 6443 104
rect 6793 108 6827 142
rect 6581 60 6615 94
rect 7009 121 7043 155
rect 7111 121 7145 155
rect 6677 48 6711 82
rect 7269 106 7303 140
rect 7543 106 7577 140
rect 7671 110 7705 144
rect 7780 138 7814 172
rect 7916 122 7950 156
rect 8084 222 8118 256
rect 8220 222 8254 256
rect 8322 222 8356 256
rect 8023 70 8057 104
rect 8419 104 8453 138
rect 8547 138 8581 172
rect 8699 138 8733 172
rect 8287 48 8321 82
rect 8867 222 8901 256
rect 9003 222 9037 256
rect 8801 70 8835 104
rect 9185 108 9219 142
rect 8973 60 9007 94
rect 9401 121 9435 155
rect 9503 121 9537 155
rect 9069 48 9103 82
rect 9661 106 9695 140
rect 9935 106 9969 140
rect 10063 110 10097 144
rect 10172 138 10206 172
rect 10308 122 10342 156
rect 10476 222 10510 256
rect 10612 222 10646 256
rect 10714 222 10748 256
rect 10415 70 10449 104
rect 10811 104 10845 138
rect 10939 138 10973 172
rect 11091 138 11125 172
rect 10679 48 10713 82
rect 11259 222 11293 256
rect 11395 222 11429 256
rect 11193 70 11227 104
rect 11577 108 11611 142
rect 11365 60 11399 94
rect 11793 121 11827 155
rect 11895 121 11929 155
rect 11461 48 11495 82
rect 12053 106 12087 140
rect 12327 106 12361 140
rect 12455 110 12489 144
rect 12564 138 12598 172
rect 12700 122 12734 156
rect 12868 222 12902 256
rect 13004 222 13038 256
rect 13106 222 13140 256
rect 12807 70 12841 104
rect 13203 104 13237 138
rect 13331 138 13365 172
rect 13483 138 13517 172
rect 13071 48 13105 82
rect 13651 222 13685 256
rect 13787 222 13821 256
rect 13585 70 13619 104
rect 13969 108 14003 142
rect 13757 60 13791 94
rect 14185 121 14219 155
rect 14287 121 14321 155
rect 13853 48 13887 82
rect 14445 106 14479 140
rect 14719 106 14753 140
rect 14847 110 14881 144
rect 14956 138 14990 172
rect 15092 122 15126 156
rect 15260 222 15294 256
rect 15396 222 15430 256
rect 15498 222 15532 256
rect 15199 70 15233 104
rect 15595 104 15629 138
rect 15723 138 15757 172
rect 15875 138 15909 172
rect 15463 48 15497 82
rect 16043 222 16077 256
rect 16179 222 16213 256
rect 15977 70 16011 104
rect 16361 108 16395 142
rect 16149 60 16183 94
rect 16577 121 16611 155
rect 16679 121 16713 155
rect 16245 48 16279 82
<< locali >>
rect 2 2937 31 2995
rect 65 2937 123 2995
rect 157 2937 215 2995
rect 249 2937 307 2995
rect 341 2937 399 2995
rect 433 2937 491 2995
rect 525 2937 583 2995
rect 617 2937 675 2995
rect 709 2937 767 2995
rect 801 2937 859 2995
rect 893 2937 951 2995
rect 985 2937 1043 2995
rect 1077 2937 1135 2995
rect 1169 2937 1227 2995
rect 1261 2937 1319 2995
rect 1353 2937 1411 2995
rect 1445 2937 1503 2995
rect 1537 2937 1595 2995
rect 1629 2937 1687 2995
rect 1721 2937 1779 2995
rect 1813 2937 1871 2995
rect 1905 2937 1963 2995
rect 1997 2937 2055 2995
rect 2089 2937 2147 2995
rect 2181 2937 2239 2995
rect 2273 2937 2331 2995
rect 2365 2937 2423 2995
rect 2457 2937 2515 2995
rect 2549 2937 2607 2995
rect 2641 2937 2699 2995
rect 2733 2937 2791 2995
rect 2825 2937 2854 2995
rect 4386 2937 4415 2995
rect 4449 2937 4507 2995
rect 4541 2937 4599 2995
rect 4633 2937 4691 2995
rect 4725 2937 4783 2995
rect 4817 2937 4875 2995
rect 4909 2937 4967 2995
rect 5001 2937 5059 2995
rect 5093 2937 5151 2995
rect 5185 2937 5243 2995
rect 5277 2937 5335 2995
rect 5369 2937 5427 2995
rect 5461 2937 5519 2995
rect 5553 2937 5611 2995
rect 5645 2937 5703 2995
rect 5737 2937 5795 2995
rect 5829 2937 5887 2995
rect 5921 2937 5979 2995
rect 6013 2937 6071 2995
rect 6105 2937 6163 2995
rect 6197 2937 6255 2995
rect 6289 2937 6347 2995
rect 6381 2937 6439 2995
rect 6473 2937 6531 2995
rect 6565 2937 6623 2995
rect 6657 2937 6715 2995
rect 6749 2937 6807 2995
rect 6841 2937 6899 2995
rect 6933 2937 6991 2995
rect 7025 2937 7083 2995
rect 7117 2937 7175 2995
rect 7209 2937 7238 2995
rect 35 2887 71 2903
rect 35 2853 37 2887
rect 35 2819 71 2853
rect 35 2785 37 2819
rect 107 2887 173 2937
rect 107 2853 123 2887
rect 157 2853 173 2887
rect 107 2819 173 2853
rect 107 2785 123 2819
rect 157 2785 173 2819
rect 207 2887 261 2903
rect 207 2853 209 2887
rect 243 2853 261 2887
rect 207 2806 261 2853
rect 35 2751 71 2785
rect 207 2772 209 2806
rect 243 2772 261 2806
rect 35 2717 170 2751
rect 207 2722 261 2772
rect 136 2688 170 2717
rect 23 2675 91 2681
rect 23 2625 39 2675
rect 73 2625 91 2675
rect 23 2607 91 2625
rect 136 2672 191 2688
rect 136 2638 157 2672
rect 136 2622 191 2638
rect 225 2670 261 2722
rect 297 2889 363 2903
rect 297 2855 313 2889
rect 347 2855 363 2889
rect 297 2821 363 2855
rect 297 2787 313 2821
rect 347 2787 363 2821
rect 297 2753 363 2787
rect 397 2895 445 2937
rect 431 2861 445 2895
rect 397 2827 445 2861
rect 431 2793 445 2827
rect 397 2777 445 2793
rect 481 2873 515 2903
rect 481 2778 515 2839
rect 297 2719 313 2753
rect 347 2741 363 2753
rect 549 2895 615 2937
rect 549 2861 565 2895
rect 599 2861 615 2895
rect 549 2827 615 2861
rect 549 2793 565 2827
rect 599 2793 615 2827
rect 549 2777 615 2793
rect 649 2873 683 2903
rect 649 2778 683 2839
rect 347 2719 440 2741
rect 297 2707 440 2719
rect 296 2670 372 2673
rect 225 2659 372 2670
rect 225 2626 322 2659
rect 136 2571 170 2622
rect 37 2537 170 2571
rect 225 2562 261 2626
rect 296 2625 322 2626
rect 356 2625 372 2659
rect 406 2659 440 2707
rect 481 2733 515 2744
rect 649 2733 683 2744
rect 481 2699 683 2733
rect 717 2895 783 2937
rect 717 2861 733 2895
rect 767 2861 783 2895
rect 717 2827 783 2861
rect 717 2793 733 2827
rect 767 2793 783 2827
rect 717 2759 783 2793
rect 717 2725 733 2759
rect 767 2725 783 2759
rect 717 2707 783 2725
rect 865 2895 899 2937
rect 865 2827 899 2861
rect 865 2759 899 2793
rect 865 2699 899 2725
rect 933 2889 999 2903
rect 933 2855 949 2889
rect 983 2855 999 2889
rect 933 2821 999 2855
rect 933 2787 949 2821
rect 983 2787 999 2821
rect 933 2753 999 2787
rect 1033 2895 1067 2937
rect 1033 2827 1067 2861
rect 1033 2777 1067 2793
rect 1101 2889 1167 2903
rect 1101 2855 1117 2889
rect 1151 2855 1167 2889
rect 1101 2821 1167 2855
rect 1101 2787 1117 2821
rect 1151 2787 1167 2821
rect 933 2719 949 2753
rect 983 2733 999 2753
rect 1101 2753 1167 2787
rect 1201 2895 1235 2937
rect 1201 2827 1235 2861
rect 1201 2777 1235 2793
rect 1269 2889 1335 2903
rect 1269 2855 1285 2889
rect 1319 2855 1335 2889
rect 1269 2821 1335 2855
rect 1269 2787 1285 2821
rect 1319 2787 1335 2821
rect 1101 2733 1117 2753
rect 983 2719 1117 2733
rect 1151 2733 1167 2753
rect 1269 2753 1335 2787
rect 1369 2895 1403 2937
rect 1369 2827 1403 2861
rect 1369 2777 1403 2793
rect 1437 2889 1503 2903
rect 1437 2855 1453 2889
rect 1487 2855 1503 2889
rect 1437 2821 1503 2855
rect 1437 2787 1453 2821
rect 1487 2787 1503 2821
rect 1269 2733 1285 2753
rect 1151 2719 1285 2733
rect 1319 2733 1335 2753
rect 1437 2753 1503 2787
rect 1537 2895 1571 2937
rect 1537 2827 1571 2861
rect 1537 2777 1571 2793
rect 1605 2889 1671 2903
rect 1605 2855 1621 2889
rect 1655 2855 1671 2889
rect 1605 2821 1671 2855
rect 1605 2787 1621 2821
rect 1655 2787 1671 2821
rect 1319 2719 1403 2733
rect 933 2699 1403 2719
rect 1437 2719 1453 2753
rect 1487 2733 1503 2753
rect 1605 2753 1671 2787
rect 1705 2895 1739 2937
rect 1705 2827 1739 2861
rect 1705 2777 1739 2793
rect 1773 2889 1839 2903
rect 1773 2855 1789 2889
rect 1823 2855 1839 2889
rect 1773 2821 1839 2855
rect 1773 2787 1789 2821
rect 1823 2787 1839 2821
rect 1605 2733 1621 2753
rect 1487 2719 1621 2733
rect 1655 2733 1671 2753
rect 1773 2753 1839 2787
rect 1873 2895 1907 2937
rect 1873 2827 1907 2861
rect 1873 2777 1907 2793
rect 1941 2889 2007 2903
rect 1941 2855 1957 2889
rect 1991 2855 2007 2889
rect 1941 2821 2007 2855
rect 1941 2787 1957 2821
rect 1991 2787 2007 2821
rect 1773 2733 1789 2753
rect 1655 2719 1789 2733
rect 1823 2733 1839 2753
rect 1941 2753 2007 2787
rect 2041 2895 2075 2937
rect 2041 2827 2075 2861
rect 2041 2777 2075 2793
rect 2109 2889 2175 2903
rect 2109 2855 2125 2889
rect 2159 2855 2175 2889
rect 2109 2821 2175 2855
rect 2109 2787 2125 2821
rect 2159 2787 2175 2821
rect 1941 2733 1957 2753
rect 1823 2719 1957 2733
rect 1991 2733 2007 2753
rect 2109 2753 2175 2787
rect 2209 2895 2243 2937
rect 2209 2827 2243 2861
rect 2209 2777 2243 2793
rect 2277 2889 2343 2903
rect 2277 2855 2293 2889
rect 2327 2855 2343 2889
rect 2277 2821 2343 2855
rect 2277 2787 2293 2821
rect 2327 2787 2343 2821
rect 2109 2733 2125 2753
rect 1991 2719 2125 2733
rect 2159 2733 2175 2753
rect 2277 2753 2343 2787
rect 2377 2895 2411 2937
rect 2377 2827 2411 2861
rect 2377 2777 2411 2793
rect 2445 2889 2511 2903
rect 2445 2855 2461 2889
rect 2495 2855 2511 2889
rect 2445 2821 2511 2855
rect 2445 2787 2461 2821
rect 2495 2787 2511 2821
rect 2277 2733 2293 2753
rect 2159 2719 2293 2733
rect 2327 2733 2343 2753
rect 2445 2753 2511 2787
rect 2545 2895 2579 2937
rect 2545 2827 2579 2861
rect 2545 2777 2579 2793
rect 2613 2889 2679 2903
rect 2613 2855 2629 2889
rect 2663 2855 2679 2889
rect 2613 2821 2679 2855
rect 2613 2787 2629 2821
rect 2663 2787 2679 2821
rect 2445 2733 2461 2753
rect 2327 2719 2461 2733
rect 2495 2733 2511 2753
rect 2613 2753 2679 2787
rect 2713 2895 2747 2937
rect 4419 2887 4455 2903
rect 2713 2827 2747 2861
rect 2713 2777 2747 2793
rect 2613 2733 2629 2753
rect 2495 2719 2629 2733
rect 2663 2733 2679 2753
rect 2782 2733 2837 2882
rect 2663 2719 2837 2733
rect 1437 2699 2837 2719
rect 4419 2853 4421 2887
rect 4419 2819 4455 2853
rect 4419 2785 4421 2819
rect 4491 2887 4557 2937
rect 4491 2853 4507 2887
rect 4541 2853 4557 2887
rect 4491 2819 4557 2853
rect 4491 2785 4507 2819
rect 4541 2785 4557 2819
rect 4591 2887 4645 2903
rect 4591 2853 4593 2887
rect 4627 2853 4645 2887
rect 4591 2806 4645 2853
rect 4419 2751 4455 2785
rect 4591 2772 4593 2806
rect 4627 2772 4645 2806
rect 4419 2717 4554 2751
rect 4591 2722 4645 2772
rect 584 2664 683 2699
rect 1368 2665 1403 2699
rect 2761 2665 2837 2699
rect 4520 2688 4554 2717
rect 847 2664 1327 2665
rect 584 2659 1327 2664
rect 406 2625 456 2659
rect 490 2625 506 2659
rect 584 2626 933 2659
rect 406 2591 440 2625
rect 584 2591 683 2626
rect 847 2625 933 2626
rect 967 2625 1001 2659
rect 1035 2625 1069 2659
rect 1103 2625 1137 2659
rect 1171 2625 1205 2659
rect 1239 2625 1273 2659
rect 1307 2625 1327 2659
rect 1368 2659 2712 2665
rect 1368 2625 1433 2659
rect 1467 2625 1501 2659
rect 1535 2625 1569 2659
rect 1603 2625 1637 2659
rect 1671 2625 1705 2659
rect 1739 2625 1773 2659
rect 1807 2625 1841 2659
rect 1875 2625 1909 2659
rect 1943 2625 1977 2659
rect 2011 2625 2045 2659
rect 2079 2625 2113 2659
rect 2147 2625 2181 2659
rect 2215 2625 2249 2659
rect 2283 2625 2317 2659
rect 2351 2625 2385 2659
rect 2419 2625 2453 2659
rect 2487 2625 2521 2659
rect 2555 2625 2589 2659
rect 2623 2625 2657 2659
rect 2691 2625 2712 2659
rect 2761 2664 2915 2665
rect 2761 2630 2876 2664
rect 2910 2630 2915 2664
rect 2761 2629 2915 2630
rect 4407 2659 4475 2681
rect 1368 2591 1403 2625
rect 2761 2591 2837 2629
rect 4407 2624 4423 2659
rect 4457 2624 4475 2659
rect 4407 2607 4475 2624
rect 4520 2672 4575 2688
rect 4520 2638 4541 2672
rect 4520 2622 4575 2638
rect 4609 2672 4645 2722
rect 4681 2889 4747 2903
rect 4681 2855 4697 2889
rect 4731 2855 4747 2889
rect 4681 2821 4747 2855
rect 4681 2787 4697 2821
rect 4731 2787 4747 2821
rect 4681 2753 4747 2787
rect 4781 2895 4829 2937
rect 4815 2861 4829 2895
rect 4781 2827 4829 2861
rect 4815 2793 4829 2827
rect 4781 2777 4829 2793
rect 4865 2873 4899 2903
rect 4865 2778 4899 2839
rect 4681 2719 4697 2753
rect 4731 2741 4747 2753
rect 4933 2895 4999 2937
rect 4933 2861 4949 2895
rect 4983 2861 4999 2895
rect 4933 2827 4999 2861
rect 4933 2793 4949 2827
rect 4983 2793 4999 2827
rect 4933 2777 4999 2793
rect 5033 2873 5067 2903
rect 5033 2778 5067 2839
rect 4731 2719 4824 2741
rect 4681 2707 4824 2719
rect 4680 2672 4756 2673
rect 4609 2659 4756 2672
rect 4609 2626 4706 2659
rect 37 2516 71 2537
rect 209 2533 261 2562
rect 37 2461 71 2482
rect 107 2469 123 2503
rect 157 2469 173 2503
rect 107 2427 173 2469
rect 243 2499 261 2533
rect 209 2461 261 2499
rect 313 2557 440 2591
rect 481 2557 683 2591
rect 313 2539 347 2557
rect 481 2539 515 2557
rect 313 2461 347 2505
rect 383 2507 431 2523
rect 383 2473 397 2507
rect 383 2427 431 2473
rect 649 2539 683 2557
rect 481 2461 515 2505
rect 549 2507 615 2523
rect 549 2473 565 2507
rect 599 2473 615 2507
rect 549 2427 615 2473
rect 649 2461 683 2505
rect 717 2571 783 2587
rect 717 2537 733 2571
rect 767 2537 783 2571
rect 717 2503 783 2537
rect 717 2469 733 2503
rect 767 2469 783 2503
rect 717 2427 783 2469
rect 865 2575 899 2591
rect 865 2507 899 2541
rect 865 2427 899 2473
rect 933 2575 1403 2591
rect 933 2541 949 2575
rect 983 2557 1117 2575
rect 983 2541 999 2557
rect 933 2507 999 2541
rect 1101 2541 1117 2557
rect 1151 2557 1285 2575
rect 1151 2541 1167 2557
rect 933 2473 949 2507
rect 983 2473 999 2507
rect 933 2462 999 2473
rect 1033 2507 1067 2523
rect 1033 2427 1067 2473
rect 1101 2507 1167 2541
rect 1269 2541 1285 2557
rect 1319 2557 1403 2575
rect 1437 2575 2837 2591
rect 1319 2541 1335 2557
rect 1101 2473 1117 2507
rect 1151 2473 1167 2507
rect 1101 2462 1167 2473
rect 1201 2507 1235 2523
rect 1201 2427 1235 2473
rect 1269 2507 1335 2541
rect 1437 2541 1453 2575
rect 1487 2557 1621 2575
rect 1487 2541 1503 2557
rect 1269 2473 1285 2507
rect 1319 2473 1335 2507
rect 1269 2462 1335 2473
rect 1369 2507 1403 2523
rect 1369 2427 1403 2473
rect 1437 2507 1503 2541
rect 1605 2541 1621 2557
rect 1655 2557 1789 2575
rect 1655 2541 1671 2557
rect 1437 2473 1453 2507
rect 1487 2473 1503 2507
rect 1437 2462 1503 2473
rect 1537 2507 1571 2523
rect 1437 2461 1487 2462
rect 1537 2427 1571 2473
rect 1605 2507 1671 2541
rect 1773 2541 1789 2557
rect 1823 2557 1957 2575
rect 1823 2541 1839 2557
rect 1605 2473 1621 2507
rect 1655 2473 1671 2507
rect 1605 2462 1671 2473
rect 1705 2507 1739 2523
rect 1621 2461 1655 2462
rect 1705 2427 1739 2473
rect 1773 2507 1839 2541
rect 1941 2541 1957 2557
rect 1991 2557 2125 2575
rect 1991 2541 2007 2557
rect 1773 2473 1789 2507
rect 1823 2473 1839 2507
rect 1773 2462 1839 2473
rect 1873 2507 1907 2523
rect 1789 2461 1823 2462
rect 1873 2427 1907 2473
rect 1941 2507 2007 2541
rect 2109 2541 2125 2557
rect 2159 2557 2293 2575
rect 2159 2541 2175 2557
rect 1941 2473 1957 2507
rect 1991 2473 2007 2507
rect 1941 2462 2007 2473
rect 2041 2507 2075 2523
rect 2041 2427 2075 2473
rect 2109 2507 2175 2541
rect 2277 2541 2293 2557
rect 2327 2557 2461 2575
rect 2327 2541 2343 2557
rect 2109 2473 2125 2507
rect 2159 2473 2175 2507
rect 2109 2462 2175 2473
rect 2209 2507 2243 2523
rect 2209 2427 2243 2473
rect 2277 2507 2343 2541
rect 2445 2541 2461 2557
rect 2495 2557 2629 2575
rect 2495 2541 2511 2557
rect 2277 2473 2293 2507
rect 2327 2473 2343 2507
rect 2277 2462 2343 2473
rect 2377 2507 2411 2523
rect 2377 2427 2411 2473
rect 2445 2507 2511 2541
rect 2613 2541 2629 2557
rect 2663 2557 2837 2575
rect 4520 2571 4554 2622
rect 2663 2541 2679 2557
rect 2445 2473 2461 2507
rect 2495 2473 2511 2507
rect 2445 2462 2511 2473
rect 2545 2507 2579 2523
rect 2545 2427 2579 2473
rect 2613 2507 2679 2541
rect 2613 2473 2629 2507
rect 2663 2473 2679 2507
rect 2613 2462 2679 2473
rect 2713 2507 2747 2523
rect 2782 2483 2837 2557
rect 4421 2537 4554 2571
rect 4609 2562 4645 2626
rect 4680 2625 4706 2626
rect 4740 2625 4756 2659
rect 4790 2659 4824 2707
rect 4865 2733 4899 2744
rect 5033 2733 5067 2744
rect 4865 2699 5067 2733
rect 5101 2895 5167 2937
rect 5101 2861 5117 2895
rect 5151 2861 5167 2895
rect 5101 2827 5167 2861
rect 5101 2793 5117 2827
rect 5151 2793 5167 2827
rect 5101 2759 5167 2793
rect 5101 2725 5117 2759
rect 5151 2725 5167 2759
rect 5101 2707 5167 2725
rect 5249 2895 5283 2937
rect 5249 2827 5283 2861
rect 5249 2759 5283 2793
rect 5249 2699 5283 2725
rect 5317 2889 5383 2903
rect 5317 2855 5333 2889
rect 5367 2855 5383 2889
rect 5317 2821 5383 2855
rect 5317 2787 5333 2821
rect 5367 2787 5383 2821
rect 5317 2753 5383 2787
rect 5417 2895 5451 2937
rect 5417 2827 5451 2861
rect 5417 2777 5451 2793
rect 5485 2889 5551 2903
rect 5485 2855 5501 2889
rect 5535 2855 5551 2889
rect 5485 2821 5551 2855
rect 5485 2787 5501 2821
rect 5535 2787 5551 2821
rect 5317 2719 5333 2753
rect 5367 2733 5383 2753
rect 5485 2753 5551 2787
rect 5585 2895 5619 2937
rect 5585 2827 5619 2861
rect 5585 2777 5619 2793
rect 5653 2889 5719 2903
rect 5653 2855 5669 2889
rect 5703 2855 5719 2889
rect 5653 2821 5719 2855
rect 5653 2787 5669 2821
rect 5703 2787 5719 2821
rect 5485 2733 5501 2753
rect 5367 2719 5501 2733
rect 5535 2733 5551 2753
rect 5653 2753 5719 2787
rect 5753 2895 5787 2937
rect 5753 2827 5787 2861
rect 5753 2777 5787 2793
rect 5821 2889 5887 2903
rect 5821 2855 5837 2889
rect 5871 2855 5887 2889
rect 5821 2821 5887 2855
rect 5821 2787 5837 2821
rect 5871 2787 5887 2821
rect 5653 2733 5669 2753
rect 5535 2719 5669 2733
rect 5703 2733 5719 2753
rect 5821 2753 5887 2787
rect 5921 2895 5955 2937
rect 5921 2827 5955 2861
rect 5921 2777 5955 2793
rect 5989 2889 6055 2903
rect 5989 2855 6005 2889
rect 6039 2855 6055 2889
rect 5989 2821 6055 2855
rect 5989 2787 6005 2821
rect 6039 2787 6055 2821
rect 5703 2719 5787 2733
rect 5317 2699 5787 2719
rect 5821 2719 5837 2753
rect 5871 2733 5887 2753
rect 5989 2753 6055 2787
rect 6089 2895 6123 2937
rect 6089 2827 6123 2861
rect 6089 2777 6123 2793
rect 6157 2889 6223 2903
rect 6157 2855 6173 2889
rect 6207 2855 6223 2889
rect 6157 2821 6223 2855
rect 6157 2787 6173 2821
rect 6207 2787 6223 2821
rect 5989 2733 6005 2753
rect 5871 2719 6005 2733
rect 6039 2733 6055 2753
rect 6157 2753 6223 2787
rect 6257 2895 6291 2937
rect 6257 2827 6291 2861
rect 6257 2777 6291 2793
rect 6325 2889 6391 2903
rect 6325 2855 6341 2889
rect 6375 2855 6391 2889
rect 6325 2821 6391 2855
rect 6325 2787 6341 2821
rect 6375 2787 6391 2821
rect 6157 2733 6173 2753
rect 6039 2719 6173 2733
rect 6207 2733 6223 2753
rect 6325 2753 6391 2787
rect 6425 2895 6459 2937
rect 6425 2827 6459 2861
rect 6425 2777 6459 2793
rect 6493 2889 6559 2903
rect 6493 2855 6509 2889
rect 6543 2855 6559 2889
rect 6493 2821 6559 2855
rect 6493 2787 6509 2821
rect 6543 2787 6559 2821
rect 6325 2733 6341 2753
rect 6207 2719 6341 2733
rect 6375 2733 6391 2753
rect 6493 2753 6559 2787
rect 6593 2895 6627 2937
rect 6593 2827 6627 2861
rect 6593 2777 6627 2793
rect 6661 2889 6727 2903
rect 6661 2855 6677 2889
rect 6711 2855 6727 2889
rect 6661 2821 6727 2855
rect 6661 2787 6677 2821
rect 6711 2787 6727 2821
rect 6493 2733 6509 2753
rect 6375 2719 6509 2733
rect 6543 2733 6559 2753
rect 6661 2753 6727 2787
rect 6761 2895 6795 2937
rect 6761 2827 6795 2861
rect 6761 2777 6795 2793
rect 6829 2889 6895 2903
rect 6829 2855 6845 2889
rect 6879 2855 6895 2889
rect 6829 2821 6895 2855
rect 6829 2787 6845 2821
rect 6879 2787 6895 2821
rect 6661 2733 6677 2753
rect 6543 2719 6677 2733
rect 6711 2733 6727 2753
rect 6829 2753 6895 2787
rect 6929 2895 6963 2937
rect 6929 2827 6963 2861
rect 6929 2777 6963 2793
rect 6997 2889 7063 2903
rect 6997 2855 7013 2889
rect 7047 2855 7063 2889
rect 6997 2821 7063 2855
rect 6997 2787 7013 2821
rect 7047 2787 7063 2821
rect 6829 2733 6845 2753
rect 6711 2719 6845 2733
rect 6879 2733 6895 2753
rect 6997 2753 7063 2787
rect 7097 2895 7131 2937
rect 7097 2827 7131 2861
rect 7097 2777 7131 2793
rect 6997 2733 7013 2753
rect 6879 2719 7013 2733
rect 7047 2733 7063 2753
rect 7166 2733 7221 2882
rect 7047 2719 7221 2733
rect 5821 2699 7221 2719
rect 4968 2666 5067 2699
rect 4968 2665 5238 2666
rect 5752 2665 5787 2699
rect 7145 2666 7221 2699
rect 4968 2659 5711 2665
rect 4790 2625 4840 2659
rect 4874 2625 4890 2659
rect 4968 2626 5317 2659
rect 4790 2591 4824 2625
rect 4968 2591 5067 2626
rect 5231 2625 5317 2626
rect 5351 2625 5385 2659
rect 5419 2625 5453 2659
rect 5487 2625 5521 2659
rect 5555 2625 5589 2659
rect 5623 2625 5657 2659
rect 5691 2625 5711 2659
rect 5752 2659 7096 2665
rect 5752 2625 5817 2659
rect 5851 2625 5885 2659
rect 5919 2625 5953 2659
rect 5987 2625 6021 2659
rect 6055 2625 6089 2659
rect 6123 2625 6157 2659
rect 6191 2625 6225 2659
rect 6259 2625 6293 2659
rect 6327 2625 6361 2659
rect 6395 2625 6429 2659
rect 6463 2625 6497 2659
rect 6531 2625 6565 2659
rect 6599 2625 6633 2659
rect 6667 2625 6701 2659
rect 6735 2625 6769 2659
rect 6803 2625 6837 2659
rect 6871 2625 6905 2659
rect 6939 2625 6973 2659
rect 7007 2625 7041 2659
rect 7075 2625 7096 2659
rect 7145 2632 7176 2666
rect 7210 2632 7221 2666
rect 5752 2591 5787 2625
rect 7145 2591 7221 2632
rect 4421 2516 4455 2537
rect 2713 2427 2747 2473
rect 4593 2533 4645 2562
rect 4421 2461 4455 2482
rect 4491 2469 4507 2503
rect 4541 2469 4557 2503
rect 4491 2427 4557 2469
rect 4627 2499 4645 2533
rect 4593 2461 4645 2499
rect 4697 2557 4824 2591
rect 4865 2557 5067 2591
rect 4697 2539 4731 2557
rect 4865 2539 4899 2557
rect 4697 2461 4731 2505
rect 4767 2507 4815 2523
rect 4767 2473 4781 2507
rect 4767 2427 4815 2473
rect 5033 2539 5067 2557
rect 4865 2461 4899 2505
rect 4933 2507 4999 2523
rect 4933 2473 4949 2507
rect 4983 2473 4999 2507
rect 4933 2427 4999 2473
rect 5033 2461 5067 2505
rect 5101 2571 5167 2587
rect 5101 2537 5117 2571
rect 5151 2537 5167 2571
rect 5101 2503 5167 2537
rect 5101 2469 5117 2503
rect 5151 2469 5167 2503
rect 5101 2427 5167 2469
rect 5249 2575 5283 2591
rect 5249 2507 5283 2541
rect 5249 2427 5283 2473
rect 5317 2575 5787 2591
rect 5317 2541 5333 2575
rect 5367 2557 5501 2575
rect 5367 2541 5383 2557
rect 5317 2507 5383 2541
rect 5485 2541 5501 2557
rect 5535 2557 5669 2575
rect 5535 2541 5551 2557
rect 5317 2473 5333 2507
rect 5367 2473 5383 2507
rect 5317 2462 5383 2473
rect 5417 2507 5451 2523
rect 5417 2427 5451 2473
rect 5485 2507 5551 2541
rect 5653 2541 5669 2557
rect 5703 2557 5787 2575
rect 5821 2575 7221 2591
rect 5703 2541 5719 2557
rect 5485 2473 5501 2507
rect 5535 2473 5551 2507
rect 5485 2462 5551 2473
rect 5585 2507 5619 2523
rect 5585 2427 5619 2473
rect 5653 2507 5719 2541
rect 5821 2541 5837 2575
rect 5871 2557 6005 2575
rect 5871 2541 5887 2557
rect 5653 2473 5669 2507
rect 5703 2473 5719 2507
rect 5653 2462 5719 2473
rect 5753 2507 5787 2523
rect 5753 2427 5787 2473
rect 5821 2507 5887 2541
rect 5989 2541 6005 2557
rect 6039 2557 6173 2575
rect 6039 2541 6055 2557
rect 5821 2473 5837 2507
rect 5871 2473 5887 2507
rect 5821 2462 5887 2473
rect 5921 2507 5955 2523
rect 5821 2461 5871 2462
rect 5921 2427 5955 2473
rect 5989 2507 6055 2541
rect 6157 2541 6173 2557
rect 6207 2557 6341 2575
rect 6207 2541 6223 2557
rect 5989 2473 6005 2507
rect 6039 2473 6055 2507
rect 5989 2462 6055 2473
rect 6089 2507 6123 2523
rect 6005 2461 6039 2462
rect 6089 2427 6123 2473
rect 6157 2507 6223 2541
rect 6325 2541 6341 2557
rect 6375 2557 6509 2575
rect 6375 2541 6391 2557
rect 6157 2473 6173 2507
rect 6207 2473 6223 2507
rect 6157 2462 6223 2473
rect 6257 2507 6291 2523
rect 6173 2461 6207 2462
rect 6257 2427 6291 2473
rect 6325 2507 6391 2541
rect 6493 2541 6509 2557
rect 6543 2557 6677 2575
rect 6543 2541 6559 2557
rect 6325 2473 6341 2507
rect 6375 2473 6391 2507
rect 6325 2462 6391 2473
rect 6425 2507 6459 2523
rect 6425 2427 6459 2473
rect 6493 2507 6559 2541
rect 6661 2541 6677 2557
rect 6711 2557 6845 2575
rect 6711 2541 6727 2557
rect 6493 2473 6509 2507
rect 6543 2473 6559 2507
rect 6493 2462 6559 2473
rect 6593 2507 6627 2523
rect 6593 2427 6627 2473
rect 6661 2507 6727 2541
rect 6829 2541 6845 2557
rect 6879 2557 7013 2575
rect 6879 2541 6895 2557
rect 6661 2473 6677 2507
rect 6711 2473 6727 2507
rect 6661 2462 6727 2473
rect 6761 2507 6795 2523
rect 6761 2427 6795 2473
rect 6829 2507 6895 2541
rect 6997 2541 7013 2557
rect 7047 2557 7221 2575
rect 7047 2541 7063 2557
rect 6829 2473 6845 2507
rect 6879 2473 6895 2507
rect 6829 2462 6895 2473
rect 6929 2507 6963 2523
rect 6929 2427 6963 2473
rect 6997 2507 7063 2541
rect 6997 2473 7013 2507
rect 7047 2473 7063 2507
rect 6997 2462 7063 2473
rect 7097 2507 7131 2523
rect 7166 2483 7221 2557
rect 7097 2427 7131 2473
rect 2 2369 31 2427
rect 65 2369 123 2427
rect 157 2369 215 2427
rect 249 2369 307 2427
rect 341 2369 399 2427
rect 433 2369 491 2427
rect 525 2369 583 2427
rect 617 2369 675 2427
rect 709 2369 767 2427
rect 801 2369 859 2427
rect 893 2369 951 2427
rect 985 2369 1043 2427
rect 1077 2369 1135 2427
rect 1169 2369 1227 2427
rect 1261 2369 1319 2427
rect 1353 2369 1411 2427
rect 1445 2369 1503 2427
rect 1537 2369 1595 2427
rect 1629 2369 1687 2427
rect 1721 2369 1779 2427
rect 1813 2369 1871 2427
rect 1905 2369 1963 2427
rect 1997 2369 2055 2427
rect 2089 2369 2147 2427
rect 2181 2369 2239 2427
rect 2273 2369 2331 2427
rect 2365 2369 2423 2427
rect 2457 2369 2515 2427
rect 2549 2369 2607 2427
rect 2641 2369 2699 2427
rect 2733 2369 2791 2427
rect 2825 2369 2854 2427
rect 4386 2369 4415 2427
rect 4449 2369 4507 2427
rect 4541 2369 4599 2427
rect 4633 2369 4691 2427
rect 4725 2369 4783 2427
rect 4817 2369 4875 2427
rect 4909 2369 4967 2427
rect 5001 2369 5059 2427
rect 5093 2369 5151 2427
rect 5185 2369 5243 2427
rect 5277 2369 5335 2427
rect 5369 2369 5427 2427
rect 5461 2369 5519 2427
rect 5553 2369 5611 2427
rect 5645 2369 5703 2427
rect 5737 2369 5795 2427
rect 5829 2369 5887 2427
rect 5921 2369 5979 2427
rect 6013 2369 6071 2427
rect 6105 2369 6163 2427
rect 6197 2369 6255 2427
rect 6289 2369 6347 2427
rect 6381 2369 6439 2427
rect 6473 2369 6531 2427
rect 6565 2369 6623 2427
rect 6657 2369 6715 2427
rect 6749 2369 6807 2427
rect 6841 2369 6899 2427
rect 6933 2369 6991 2427
rect 7025 2369 7083 2427
rect 7117 2369 7175 2427
rect 7209 2369 7238 2427
rect 0 1795 29 1853
rect 63 1795 121 1853
rect 155 1795 213 1853
rect 247 1795 305 1853
rect 339 1795 397 1853
rect 431 1795 489 1853
rect 523 1795 581 1853
rect 615 1795 673 1853
rect 707 1795 765 1853
rect 799 1819 857 1853
rect 891 1819 949 1853
rect 983 1819 1041 1853
rect 1075 1819 1133 1853
rect 1167 1819 1225 1853
rect 1259 1819 1317 1853
rect 1351 1819 1409 1853
rect 1443 1829 1501 1853
rect 1443 1819 1463 1829
rect 799 1804 1463 1819
rect 799 1795 828 1804
rect 1434 1795 1463 1804
rect 1497 1819 1501 1829
rect 1535 1829 1593 1853
rect 1535 1819 1555 1829
rect 1497 1795 1555 1819
rect 1589 1819 1593 1829
rect 1627 1829 1685 1853
rect 1627 1819 1647 1829
rect 1589 1795 1647 1819
rect 1681 1819 1685 1829
rect 1719 1829 1777 1853
rect 1719 1819 1739 1829
rect 1681 1795 1739 1819
rect 1773 1819 1777 1829
rect 1811 1829 1869 1853
rect 1811 1819 1831 1829
rect 1773 1795 1831 1819
rect 1865 1819 1869 1829
rect 1903 1829 1961 1853
rect 1903 1819 1923 1829
rect 1865 1795 1923 1819
rect 1957 1819 1961 1829
rect 1995 1829 2053 1853
rect 1995 1819 2015 1829
rect 1957 1795 2015 1819
rect 2049 1819 2053 1829
rect 2087 1829 2145 1853
rect 2087 1819 2107 1829
rect 2049 1795 2107 1819
rect 2141 1819 2145 1829
rect 2179 1829 2237 1853
rect 2179 1819 2199 1829
rect 2141 1795 2199 1819
rect 2233 1819 2237 1829
rect 2271 1819 2329 1853
rect 2363 1819 2421 1853
rect 2233 1804 2421 1819
rect 2233 1795 2262 1804
rect 2392 1795 2421 1804
rect 2455 1795 2513 1853
rect 2547 1795 2605 1853
rect 2639 1795 2697 1853
rect 2731 1795 2789 1853
rect 2823 1795 2881 1853
rect 2915 1795 2973 1853
rect 3007 1795 3065 1853
rect 3099 1795 3157 1853
rect 3191 1819 3249 1853
rect 3283 1819 3341 1853
rect 3375 1819 3433 1853
rect 3467 1819 3525 1853
rect 3559 1819 3617 1853
rect 3651 1819 3709 1853
rect 3743 1819 3801 1853
rect 3835 1829 3893 1853
rect 3835 1819 3855 1829
rect 3191 1804 3855 1819
rect 3191 1795 3220 1804
rect 3826 1795 3855 1804
rect 3889 1819 3893 1829
rect 3927 1829 3985 1853
rect 3927 1819 3947 1829
rect 3889 1795 3947 1819
rect 3981 1819 3985 1829
rect 4019 1829 4077 1853
rect 4019 1819 4039 1829
rect 3981 1795 4039 1819
rect 4073 1819 4077 1829
rect 4111 1829 4169 1853
rect 4111 1819 4131 1829
rect 4073 1795 4131 1819
rect 4165 1819 4169 1829
rect 4203 1829 4261 1853
rect 4203 1819 4223 1829
rect 4165 1795 4223 1819
rect 4257 1819 4261 1829
rect 4295 1829 4353 1853
rect 4295 1819 4315 1829
rect 4257 1795 4315 1819
rect 4349 1819 4353 1829
rect 4387 1829 4445 1853
rect 4387 1819 4407 1829
rect 4349 1795 4407 1819
rect 4441 1819 4445 1829
rect 4479 1829 4537 1853
rect 4479 1819 4499 1829
rect 4441 1795 4499 1819
rect 4533 1819 4537 1829
rect 4571 1829 4629 1853
rect 4571 1819 4591 1829
rect 4533 1795 4591 1819
rect 4625 1819 4629 1829
rect 4663 1819 4721 1853
rect 4755 1819 4813 1853
rect 4625 1804 4813 1819
rect 4625 1795 4654 1804
rect 4784 1795 4813 1804
rect 4847 1795 4905 1853
rect 4939 1795 4997 1853
rect 5031 1795 5089 1853
rect 5123 1795 5181 1853
rect 5215 1795 5273 1853
rect 5307 1795 5365 1853
rect 5399 1795 5457 1853
rect 5491 1795 5549 1853
rect 5583 1819 5641 1853
rect 5675 1819 6245 1853
rect 5583 1804 6245 1819
rect 5583 1795 5612 1804
rect 6216 1795 6245 1804
rect 6279 1795 6337 1853
rect 6371 1795 6429 1853
rect 6463 1795 6521 1853
rect 6555 1795 6613 1853
rect 6647 1795 6705 1853
rect 6739 1795 6797 1853
rect 6831 1795 6889 1853
rect 6923 1795 6981 1853
rect 7015 1819 7073 1853
rect 7107 1819 7165 1853
rect 7199 1829 7257 1853
rect 7199 1819 7205 1829
rect 7015 1804 7205 1819
rect 7015 1795 7044 1804
rect 7176 1795 7205 1804
rect 7239 1819 7257 1829
rect 7291 1829 7349 1853
rect 7291 1819 7297 1829
rect 7239 1795 7297 1819
rect 7331 1819 7349 1829
rect 7383 1829 7441 1853
rect 7383 1819 7389 1829
rect 7331 1795 7389 1819
rect 7423 1819 7441 1829
rect 7475 1829 7533 1853
rect 7475 1819 7481 1829
rect 7423 1795 7481 1819
rect 7515 1819 7533 1829
rect 7567 1829 7625 1853
rect 7567 1819 7573 1829
rect 7515 1795 7573 1819
rect 7607 1819 7625 1829
rect 7659 1829 7717 1853
rect 7659 1819 7665 1829
rect 7607 1795 7665 1819
rect 7699 1819 7717 1829
rect 7751 1829 7809 1853
rect 7751 1819 7757 1829
rect 7699 1795 7757 1819
rect 7791 1819 7809 1829
rect 7843 1829 7901 1853
rect 7843 1819 7849 1829
rect 7791 1795 7849 1819
rect 7883 1819 7901 1829
rect 7935 1829 7993 1853
rect 7935 1819 7941 1829
rect 7883 1795 7941 1819
rect 7975 1819 7993 1829
rect 8027 1819 8085 1853
rect 8119 1819 8177 1853
rect 8211 1819 8269 1853
rect 8303 1819 8361 1853
rect 8395 1819 8453 1853
rect 8487 1819 8545 1853
rect 8579 1819 8637 1853
rect 8671 1829 8729 1853
rect 8763 1829 8821 1853
rect 8855 1829 8913 1853
rect 8947 1829 9005 1853
rect 9039 1829 9097 1853
rect 9131 1829 9189 1853
rect 9223 1829 9281 1853
rect 9315 1829 9373 1853
rect 9407 1829 9465 1853
rect 8673 1819 8729 1829
rect 8765 1819 8821 1829
rect 8857 1819 8913 1829
rect 8949 1819 9005 1829
rect 9041 1819 9097 1829
rect 9133 1819 9189 1829
rect 9225 1819 9281 1829
rect 9317 1819 9373 1829
rect 9409 1819 9465 1829
rect 9499 1819 9557 1853
rect 9591 1829 9649 1853
rect 9591 1819 9597 1829
rect 7975 1804 8639 1819
rect 7975 1795 8004 1804
rect 8610 1795 8639 1804
rect 8673 1795 8731 1819
rect 8765 1795 8823 1819
rect 8857 1795 8915 1819
rect 8949 1795 9007 1819
rect 9041 1795 9099 1819
rect 9133 1795 9191 1819
rect 9225 1795 9283 1819
rect 9317 1795 9375 1819
rect 9409 1804 9597 1819
rect 9409 1795 9438 1804
rect 9568 1795 9597 1804
rect 9631 1819 9649 1829
rect 9683 1829 9741 1853
rect 9683 1819 9689 1829
rect 9631 1795 9689 1819
rect 9723 1819 9741 1829
rect 9775 1829 9833 1853
rect 9775 1819 9781 1829
rect 9723 1795 9781 1819
rect 9815 1819 9833 1829
rect 9867 1829 9925 1853
rect 9867 1819 9873 1829
rect 9815 1795 9873 1819
rect 9907 1819 9925 1829
rect 9959 1829 10017 1853
rect 9959 1819 9965 1829
rect 9907 1795 9965 1819
rect 9999 1819 10017 1829
rect 10051 1829 10109 1853
rect 10051 1819 10057 1829
rect 9999 1795 10057 1819
rect 10091 1819 10109 1829
rect 10143 1829 10201 1853
rect 10143 1819 10149 1829
rect 10091 1795 10149 1819
rect 10183 1819 10201 1829
rect 10235 1829 10293 1853
rect 10235 1819 10241 1829
rect 10183 1795 10241 1819
rect 10275 1819 10293 1829
rect 10327 1829 10385 1853
rect 10327 1819 10333 1829
rect 10275 1795 10333 1819
rect 10367 1819 10385 1829
rect 10419 1819 10477 1853
rect 10511 1819 10569 1853
rect 10603 1819 10661 1853
rect 10695 1819 10753 1853
rect 10787 1819 10845 1853
rect 10879 1819 10937 1853
rect 10971 1819 11029 1853
rect 11063 1829 11121 1853
rect 11155 1829 11213 1853
rect 11247 1829 11305 1853
rect 11339 1829 11397 1853
rect 11431 1829 11489 1853
rect 11523 1829 11581 1853
rect 11615 1829 11673 1853
rect 11707 1829 11765 1853
rect 11799 1829 11857 1853
rect 11065 1819 11121 1829
rect 11157 1819 11213 1829
rect 11249 1819 11305 1829
rect 11341 1819 11397 1829
rect 11433 1819 11489 1829
rect 11525 1819 11581 1829
rect 11617 1819 11673 1829
rect 11709 1819 11765 1829
rect 11801 1819 11857 1829
rect 11891 1829 12011 1853
rect 12045 1829 12103 1853
rect 12137 1829 12195 1853
rect 12229 1829 12287 1853
rect 12321 1829 12379 1853
rect 12413 1829 12471 1853
rect 12505 1829 12563 1853
rect 12597 1829 12655 1853
rect 12689 1829 12747 1853
rect 11891 1819 11989 1829
rect 12045 1819 12081 1829
rect 12137 1819 12173 1829
rect 12229 1819 12265 1829
rect 12321 1819 12357 1829
rect 12413 1819 12449 1829
rect 12505 1819 12541 1829
rect 12597 1819 12633 1829
rect 12689 1819 12725 1829
rect 12781 1819 12839 1853
rect 12873 1819 12931 1853
rect 12965 1819 13023 1853
rect 13057 1819 13115 1853
rect 13149 1819 13207 1853
rect 13241 1819 13299 1853
rect 13333 1819 13391 1853
rect 13425 1829 13483 1853
rect 13517 1829 13575 1853
rect 13609 1829 13667 1853
rect 13701 1829 13759 1853
rect 13793 1829 13851 1853
rect 13885 1829 13943 1853
rect 13977 1829 14035 1853
rect 14069 1829 14127 1853
rect 14161 1829 14219 1853
rect 13455 1819 13483 1829
rect 13547 1819 13575 1829
rect 13639 1819 13667 1829
rect 13731 1819 13759 1829
rect 13823 1819 13851 1829
rect 13915 1819 13943 1829
rect 14007 1819 14035 1829
rect 14099 1819 14127 1829
rect 14191 1819 14219 1829
rect 14253 1819 14311 1853
rect 14345 1829 14403 1853
rect 14437 1829 14495 1853
rect 14529 1829 14587 1853
rect 14621 1829 14679 1853
rect 14713 1829 14771 1853
rect 14805 1829 14863 1853
rect 14897 1829 14955 1853
rect 14989 1829 15047 1853
rect 15081 1829 15139 1853
rect 14345 1819 14381 1829
rect 14437 1819 14473 1829
rect 14529 1819 14565 1829
rect 14621 1819 14657 1829
rect 14713 1819 14749 1829
rect 14805 1819 14841 1829
rect 14897 1819 14933 1829
rect 14989 1819 15025 1829
rect 15081 1819 15117 1829
rect 15173 1819 15231 1853
rect 15265 1819 15323 1853
rect 15357 1819 15415 1853
rect 15449 1819 15507 1853
rect 15541 1819 15599 1853
rect 15633 1819 15691 1853
rect 15725 1819 15783 1853
rect 15817 1829 15875 1853
rect 15909 1829 15967 1853
rect 16001 1829 16059 1853
rect 16093 1829 16151 1853
rect 16185 1829 16243 1853
rect 16277 1829 16335 1853
rect 16369 1829 16427 1853
rect 16461 1829 16519 1853
rect 16553 1829 16614 1853
rect 15849 1819 15875 1829
rect 15941 1819 15967 1829
rect 16033 1819 16059 1829
rect 16125 1819 16151 1829
rect 16217 1819 16243 1829
rect 16309 1819 16335 1829
rect 16401 1819 16427 1829
rect 16493 1819 16519 1829
rect 10367 1804 11031 1819
rect 10367 1795 10396 1804
rect 11002 1795 11031 1804
rect 11065 1795 11123 1819
rect 11157 1795 11215 1819
rect 11249 1795 11307 1819
rect 11341 1795 11399 1819
rect 11433 1795 11491 1819
rect 11525 1795 11583 1819
rect 11617 1795 11675 1819
rect 11709 1795 11767 1819
rect 11801 1804 11989 1819
rect 11801 1795 11830 1804
rect 11960 1795 11989 1804
rect 12023 1795 12081 1819
rect 12115 1795 12173 1819
rect 12207 1795 12265 1819
rect 12299 1795 12357 1819
rect 12391 1795 12449 1819
rect 12483 1795 12541 1819
rect 12575 1795 12633 1819
rect 12667 1795 12725 1819
rect 12759 1804 13421 1819
rect 12759 1795 12788 1804
rect 13392 1795 13421 1804
rect 13455 1795 13513 1819
rect 13547 1795 13605 1819
rect 13639 1795 13697 1819
rect 13731 1795 13789 1819
rect 13823 1795 13881 1819
rect 13915 1795 13973 1819
rect 14007 1795 14065 1819
rect 14099 1795 14157 1819
rect 14191 1804 14381 1819
rect 14191 1795 14220 1804
rect 14352 1795 14381 1804
rect 14415 1795 14473 1819
rect 14507 1795 14565 1819
rect 14599 1795 14657 1819
rect 14691 1795 14749 1819
rect 14783 1795 14841 1819
rect 14875 1795 14933 1819
rect 14967 1795 15025 1819
rect 15059 1795 15117 1819
rect 15151 1804 15815 1819
rect 15151 1795 15180 1804
rect 15786 1795 15815 1804
rect 15849 1795 15907 1819
rect 15941 1795 15999 1819
rect 16033 1795 16091 1819
rect 16125 1795 16183 1819
rect 16217 1795 16275 1819
rect 16309 1795 16367 1819
rect 16401 1795 16459 1819
rect 16493 1795 16551 1819
rect 16585 1795 16614 1829
rect 18 1753 85 1761
rect 18 1719 35 1753
rect 69 1719 85 1753
rect 18 1685 85 1719
rect 18 1651 35 1685
rect 69 1651 85 1685
rect 18 1617 85 1651
rect 18 1583 35 1617
rect 69 1583 85 1617
rect 18 1567 85 1583
rect 119 1753 153 1795
rect 119 1685 153 1719
rect 119 1617 153 1651
rect 119 1567 153 1583
rect 187 1727 593 1761
rect 18 1433 52 1567
rect 187 1533 221 1727
rect 86 1517 137 1533
rect 120 1483 137 1517
rect 86 1467 137 1483
rect 182 1517 221 1533
rect 216 1483 221 1517
rect 182 1467 221 1483
rect 255 1659 355 1693
rect 389 1659 430 1693
rect 464 1659 480 1693
rect 103 1433 137 1467
rect 255 1433 289 1659
rect 18 1406 69 1433
rect 18 1372 28 1406
rect 62 1380 69 1406
rect 103 1399 289 1433
rect 323 1607 525 1625
rect 323 1591 484 1607
rect 518 1594 525 1607
rect 323 1481 357 1591
rect 487 1560 491 1573
rect 323 1431 357 1447
rect 398 1481 453 1551
rect 398 1447 419 1481
rect 18 1346 35 1372
rect 254 1392 289 1399
rect 254 1376 360 1392
rect 18 1319 69 1346
rect 103 1361 169 1365
rect 103 1327 119 1361
rect 153 1327 169 1361
rect 103 1285 169 1327
rect 254 1342 326 1376
rect 254 1319 360 1342
rect 398 1285 453 1447
rect 487 1319 525 1560
rect 559 1594 593 1727
rect 627 1693 661 1795
rect 627 1643 661 1659
rect 708 1693 811 1725
rect 708 1659 713 1693
rect 747 1659 811 1693
rect 708 1643 811 1659
rect 559 1591 659 1594
rect 559 1557 656 1591
rect 693 1560 709 1594
rect 690 1557 709 1560
rect 559 1556 709 1557
rect 743 1481 811 1643
rect 565 1447 581 1481
rect 615 1447 811 1481
rect 1451 1693 1554 1725
rect 1451 1659 1515 1693
rect 1549 1659 1554 1693
rect 1451 1643 1554 1659
rect 1601 1693 1635 1795
rect 1601 1643 1635 1659
rect 1669 1727 2075 1761
rect 1451 1481 1519 1643
rect 1669 1594 1703 1727
rect 1782 1659 1798 1693
rect 1832 1659 1873 1693
rect 1907 1659 2007 1693
rect 1553 1592 1569 1594
rect 1553 1558 1566 1592
rect 1603 1560 1703 1594
rect 1600 1558 1703 1560
rect 1553 1556 1703 1558
rect 1737 1607 1939 1625
rect 1737 1594 1746 1607
rect 1780 1591 1939 1607
rect 1771 1560 1775 1573
rect 1451 1447 1647 1481
rect 1681 1447 1697 1481
rect 561 1376 663 1392
rect 595 1342 629 1376
rect 561 1285 663 1342
rect 707 1376 756 1447
rect 707 1342 713 1376
rect 747 1342 756 1376
rect 707 1326 756 1342
rect 1506 1376 1555 1447
rect 1506 1342 1515 1376
rect 1549 1342 1555 1376
rect 1506 1326 1555 1342
rect 1599 1376 1701 1392
rect 1633 1342 1667 1376
rect 1599 1285 1701 1342
rect 1737 1319 1775 1560
rect 1809 1481 1864 1551
rect 1843 1447 1864 1481
rect 1809 1285 1864 1447
rect 1905 1481 1939 1591
rect 1905 1431 1939 1447
rect 1973 1433 2007 1659
rect 2041 1533 2075 1727
rect 2109 1753 2143 1795
rect 2109 1685 2143 1719
rect 2109 1617 2143 1651
rect 2109 1567 2143 1583
rect 2177 1753 2244 1761
rect 2177 1719 2193 1753
rect 2227 1719 2244 1753
rect 2177 1685 2244 1719
rect 2177 1651 2193 1685
rect 2227 1651 2244 1685
rect 2177 1617 2244 1651
rect 2177 1583 2193 1617
rect 2227 1583 2244 1617
rect 2177 1567 2244 1583
rect 2041 1517 2080 1533
rect 2041 1483 2046 1517
rect 2041 1467 2080 1483
rect 2125 1517 2176 1533
rect 2125 1483 2142 1517
rect 2125 1467 2176 1483
rect 2125 1433 2159 1467
rect 2210 1433 2244 1567
rect 1973 1399 2159 1433
rect 2193 1404 2244 1433
rect 1973 1392 2008 1399
rect 1902 1376 2008 1392
rect 1936 1342 2008 1376
rect 2193 1380 2204 1404
rect 2238 1370 2244 1404
rect 1902 1319 2008 1342
rect 2093 1361 2159 1365
rect 2093 1327 2109 1361
rect 2143 1327 2159 1361
rect 2093 1285 2159 1327
rect 2227 1346 2244 1370
rect 2193 1319 2244 1346
rect 2410 1753 2477 1761
rect 2410 1719 2427 1753
rect 2461 1719 2477 1753
rect 2410 1685 2477 1719
rect 2410 1651 2427 1685
rect 2461 1651 2477 1685
rect 2410 1617 2477 1651
rect 2410 1583 2427 1617
rect 2461 1583 2477 1617
rect 2410 1567 2477 1583
rect 2511 1753 2545 1795
rect 2511 1685 2545 1719
rect 2511 1617 2545 1651
rect 2511 1567 2545 1583
rect 2579 1727 2985 1761
rect 2410 1433 2444 1567
rect 2579 1533 2613 1727
rect 2478 1517 2529 1533
rect 2512 1483 2529 1517
rect 2478 1467 2529 1483
rect 2574 1517 2613 1533
rect 2608 1483 2613 1517
rect 2574 1467 2613 1483
rect 2647 1659 2747 1693
rect 2781 1659 2822 1693
rect 2856 1659 2872 1693
rect 2495 1433 2529 1467
rect 2647 1433 2681 1659
rect 2410 1406 2461 1433
rect 2410 1372 2420 1406
rect 2454 1380 2461 1406
rect 2495 1399 2681 1433
rect 2715 1606 2917 1625
rect 2715 1591 2877 1606
rect 2911 1594 2917 1606
rect 2715 1481 2749 1591
rect 2879 1560 2883 1572
rect 2715 1431 2749 1447
rect 2790 1481 2845 1551
rect 2790 1447 2811 1481
rect 2410 1346 2427 1372
rect 2646 1392 2681 1399
rect 2646 1376 2752 1392
rect 2410 1319 2461 1346
rect 2495 1361 2561 1365
rect 2495 1327 2511 1361
rect 2545 1327 2561 1361
rect 2495 1285 2561 1327
rect 2646 1342 2718 1376
rect 2646 1319 2752 1342
rect 2790 1285 2845 1447
rect 2879 1319 2917 1560
rect 2951 1594 2985 1727
rect 3019 1693 3053 1795
rect 3019 1643 3053 1659
rect 3100 1693 3203 1725
rect 3100 1659 3105 1693
rect 3139 1659 3203 1693
rect 3100 1643 3203 1659
rect 2951 1590 3051 1594
rect 2951 1556 3048 1590
rect 3085 1560 3101 1594
rect 3082 1556 3101 1560
rect 3135 1481 3203 1643
rect 2957 1447 2973 1481
rect 3007 1447 3203 1481
rect 3843 1693 3946 1725
rect 3843 1659 3907 1693
rect 3941 1659 3946 1693
rect 3843 1643 3946 1659
rect 3993 1693 4027 1795
rect 3993 1643 4027 1659
rect 4061 1727 4467 1761
rect 3843 1481 3911 1643
rect 4061 1594 4095 1727
rect 4174 1659 4190 1693
rect 4224 1659 4265 1693
rect 4299 1659 4399 1693
rect 3945 1591 3961 1594
rect 3945 1557 3958 1591
rect 3995 1560 4095 1594
rect 3992 1557 4095 1560
rect 3945 1556 4095 1557
rect 4129 1607 4331 1625
rect 4129 1594 4138 1607
rect 4172 1591 4331 1607
rect 4163 1560 4167 1573
rect 3843 1447 4039 1481
rect 4073 1447 4089 1481
rect 2953 1376 3055 1392
rect 2987 1342 3021 1376
rect 2953 1285 3055 1342
rect 3099 1376 3148 1447
rect 3099 1342 3105 1376
rect 3139 1342 3148 1376
rect 3099 1326 3148 1342
rect 3898 1376 3947 1447
rect 3898 1342 3907 1376
rect 3941 1342 3947 1376
rect 3898 1326 3947 1342
rect 3991 1376 4093 1392
rect 4025 1342 4059 1376
rect 3991 1285 4093 1342
rect 4129 1319 4167 1560
rect 4201 1481 4256 1551
rect 4235 1447 4256 1481
rect 4201 1285 4256 1447
rect 4297 1481 4331 1591
rect 4297 1431 4331 1447
rect 4365 1433 4399 1659
rect 4433 1533 4467 1727
rect 4501 1753 4535 1795
rect 4501 1685 4535 1719
rect 4501 1617 4535 1651
rect 4501 1567 4535 1583
rect 4569 1753 4636 1761
rect 4569 1719 4585 1753
rect 4619 1719 4636 1753
rect 4569 1685 4636 1719
rect 4569 1651 4585 1685
rect 4619 1651 4636 1685
rect 4569 1617 4636 1651
rect 4569 1583 4585 1617
rect 4619 1583 4636 1617
rect 4569 1567 4636 1583
rect 4433 1517 4472 1533
rect 4433 1483 4438 1517
rect 4433 1467 4472 1483
rect 4517 1517 4568 1533
rect 4517 1483 4534 1517
rect 4517 1467 4568 1483
rect 4517 1433 4551 1467
rect 4602 1433 4636 1567
rect 4365 1399 4551 1433
rect 4585 1404 4636 1433
rect 4365 1392 4400 1399
rect 4294 1376 4400 1392
rect 4328 1342 4400 1376
rect 4585 1380 4598 1404
rect 4632 1370 4636 1404
rect 4294 1319 4400 1342
rect 4485 1361 4551 1365
rect 4485 1327 4501 1361
rect 4535 1327 4551 1361
rect 4485 1285 4551 1327
rect 4619 1346 4636 1370
rect 4585 1319 4636 1346
rect 4802 1753 4869 1761
rect 4802 1719 4819 1753
rect 4853 1719 4869 1753
rect 4802 1685 4869 1719
rect 4802 1651 4819 1685
rect 4853 1651 4869 1685
rect 4802 1617 4869 1651
rect 4802 1583 4819 1617
rect 4853 1583 4869 1617
rect 4802 1567 4869 1583
rect 4903 1753 4937 1795
rect 4903 1685 4937 1719
rect 4903 1617 4937 1651
rect 4903 1567 4937 1583
rect 4971 1727 5377 1761
rect 4802 1433 4836 1567
rect 4971 1533 5005 1727
rect 4870 1517 4921 1533
rect 4904 1483 4921 1517
rect 4870 1467 4921 1483
rect 4966 1517 5005 1533
rect 5000 1483 5005 1517
rect 4966 1467 5005 1483
rect 5039 1659 5139 1693
rect 5173 1659 5214 1693
rect 5248 1659 5264 1693
rect 4887 1433 4921 1467
rect 5039 1433 5073 1659
rect 4802 1406 4853 1433
rect 4802 1372 4812 1406
rect 4846 1380 4853 1406
rect 4887 1399 5073 1433
rect 5107 1606 5309 1625
rect 5107 1591 5269 1606
rect 5303 1594 5309 1606
rect 5107 1481 5141 1591
rect 5271 1560 5275 1572
rect 5107 1431 5141 1447
rect 5182 1481 5237 1551
rect 5182 1447 5203 1481
rect 4802 1346 4819 1372
rect 5038 1392 5073 1399
rect 5038 1376 5144 1392
rect 4802 1319 4853 1346
rect 4887 1361 4953 1365
rect 4887 1327 4903 1361
rect 4937 1327 4953 1361
rect 4887 1285 4953 1327
rect 5038 1342 5110 1376
rect 5038 1319 5144 1342
rect 5182 1285 5237 1447
rect 5271 1319 5309 1560
rect 5343 1594 5377 1727
rect 5411 1693 5445 1795
rect 5411 1643 5445 1659
rect 5492 1693 5595 1725
rect 5492 1659 5497 1693
rect 5531 1659 5595 1693
rect 5492 1643 5595 1659
rect 5343 1591 5443 1594
rect 5343 1557 5439 1591
rect 5477 1560 5493 1594
rect 5473 1557 5493 1560
rect 5343 1556 5493 1557
rect 5527 1481 5595 1643
rect 5349 1447 5365 1481
rect 5399 1447 5595 1481
rect 6233 1693 6336 1725
rect 6233 1659 6297 1693
rect 6331 1659 6336 1693
rect 6233 1643 6336 1659
rect 6383 1693 6417 1795
rect 6383 1643 6417 1659
rect 6451 1727 6857 1761
rect 6233 1481 6301 1643
rect 6451 1594 6485 1727
rect 6564 1659 6580 1693
rect 6614 1659 6655 1693
rect 6689 1659 6789 1693
rect 6335 1591 6351 1594
rect 6335 1557 6348 1591
rect 6385 1560 6485 1594
rect 6382 1557 6485 1560
rect 6335 1556 6485 1557
rect 6519 1608 6721 1625
rect 6519 1594 6529 1608
rect 6563 1591 6721 1608
rect 6553 1560 6557 1574
rect 6233 1447 6429 1481
rect 6463 1447 6479 1481
rect 5345 1376 5447 1392
rect 5379 1342 5413 1376
rect 5345 1285 5447 1342
rect 5491 1376 5540 1447
rect 5491 1342 5497 1376
rect 5531 1342 5540 1376
rect 5491 1326 5540 1342
rect 6288 1376 6337 1447
rect 6288 1342 6297 1376
rect 6331 1342 6337 1376
rect 6288 1326 6337 1342
rect 6381 1376 6483 1392
rect 6415 1342 6449 1376
rect 6381 1285 6483 1342
rect 6519 1319 6557 1560
rect 6591 1481 6646 1551
rect 6625 1447 6646 1481
rect 6591 1285 6646 1447
rect 6687 1481 6721 1591
rect 6687 1431 6721 1447
rect 6755 1433 6789 1659
rect 6823 1533 6857 1727
rect 6891 1753 6925 1795
rect 6891 1685 6925 1719
rect 6891 1617 6925 1651
rect 6891 1567 6925 1583
rect 6959 1753 7026 1761
rect 6959 1719 6975 1753
rect 7009 1719 7026 1753
rect 6959 1685 7026 1719
rect 6959 1651 6975 1685
rect 7009 1651 7026 1685
rect 6959 1617 7026 1651
rect 6959 1583 6975 1617
rect 7009 1583 7026 1617
rect 6959 1567 7026 1583
rect 6823 1517 6862 1533
rect 6823 1483 6828 1517
rect 6823 1467 6862 1483
rect 6907 1517 6958 1533
rect 6907 1483 6924 1517
rect 6907 1467 6958 1483
rect 6907 1433 6941 1467
rect 6992 1433 7026 1567
rect 6755 1399 6941 1433
rect 6975 1406 7026 1433
rect 6755 1392 6790 1399
rect 6684 1376 6790 1392
rect 6718 1342 6790 1376
rect 6975 1380 6988 1406
rect 7022 1372 7026 1406
rect 6684 1319 6790 1342
rect 6875 1361 6941 1365
rect 6875 1327 6891 1361
rect 6925 1327 6941 1361
rect 6875 1285 6941 1327
rect 7009 1346 7026 1372
rect 6975 1319 7026 1346
rect 7194 1753 7261 1761
rect 7194 1719 7211 1753
rect 7245 1719 7261 1753
rect 7194 1685 7261 1719
rect 7194 1651 7211 1685
rect 7245 1651 7261 1685
rect 7194 1617 7261 1651
rect 7194 1583 7211 1617
rect 7245 1583 7261 1617
rect 7194 1567 7261 1583
rect 7295 1753 7329 1795
rect 7295 1685 7329 1719
rect 7295 1617 7329 1651
rect 7295 1567 7329 1583
rect 7363 1727 7769 1761
rect 7194 1433 7228 1567
rect 7363 1533 7397 1727
rect 7262 1517 7313 1533
rect 7296 1483 7313 1517
rect 7262 1467 7313 1483
rect 7358 1517 7397 1533
rect 7392 1483 7397 1517
rect 7358 1467 7397 1483
rect 7431 1659 7531 1693
rect 7565 1659 7606 1693
rect 7640 1659 7656 1693
rect 7279 1433 7313 1467
rect 7431 1433 7465 1659
rect 7194 1406 7245 1433
rect 7194 1372 7204 1406
rect 7238 1380 7245 1406
rect 7279 1399 7465 1433
rect 7499 1607 7701 1625
rect 7499 1591 7661 1607
rect 7695 1594 7701 1607
rect 7499 1481 7533 1591
rect 7663 1560 7667 1573
rect 7499 1431 7533 1447
rect 7574 1481 7629 1551
rect 7574 1447 7595 1481
rect 7194 1346 7211 1372
rect 7430 1392 7465 1399
rect 7430 1376 7536 1392
rect 7194 1319 7245 1346
rect 7279 1361 7345 1365
rect 7279 1327 7295 1361
rect 7329 1327 7345 1361
rect 7279 1285 7345 1327
rect 7430 1342 7502 1376
rect 7430 1319 7536 1342
rect 7574 1285 7629 1447
rect 7663 1319 7701 1560
rect 7735 1594 7769 1727
rect 7803 1693 7837 1795
rect 7803 1643 7837 1659
rect 7884 1693 7987 1725
rect 7884 1659 7889 1693
rect 7923 1659 7987 1693
rect 7884 1643 7987 1659
rect 7735 1591 7835 1594
rect 7735 1557 7832 1591
rect 7869 1560 7885 1594
rect 7866 1557 7885 1560
rect 7735 1556 7885 1557
rect 7919 1481 7987 1643
rect 7741 1447 7757 1481
rect 7791 1447 7987 1481
rect 8627 1693 8730 1725
rect 8627 1659 8691 1693
rect 8725 1659 8730 1693
rect 8627 1643 8730 1659
rect 8777 1693 8811 1795
rect 8777 1643 8811 1659
rect 8845 1727 9251 1761
rect 8627 1481 8695 1643
rect 8845 1594 8879 1727
rect 8958 1659 8974 1693
rect 9008 1659 9049 1693
rect 9083 1659 9183 1693
rect 8729 1592 8745 1594
rect 8729 1558 8742 1592
rect 8779 1560 8879 1594
rect 8776 1558 8879 1560
rect 8729 1556 8879 1558
rect 8913 1608 9115 1625
rect 8913 1594 8922 1608
rect 8956 1591 9115 1608
rect 8947 1560 8951 1574
rect 8627 1447 8823 1481
rect 8857 1447 8873 1481
rect 7737 1376 7839 1392
rect 7771 1342 7805 1376
rect 7737 1285 7839 1342
rect 7883 1376 7932 1447
rect 7883 1342 7889 1376
rect 7923 1342 7932 1376
rect 7883 1326 7932 1342
rect 8682 1376 8731 1447
rect 8682 1342 8691 1376
rect 8725 1342 8731 1376
rect 8682 1326 8731 1342
rect 8775 1376 8877 1392
rect 8809 1342 8843 1376
rect 8775 1285 8877 1342
rect 8913 1319 8951 1560
rect 8985 1481 9040 1551
rect 9019 1447 9040 1481
rect 8985 1285 9040 1447
rect 9081 1481 9115 1591
rect 9081 1431 9115 1447
rect 9149 1433 9183 1659
rect 9217 1533 9251 1727
rect 9285 1753 9319 1795
rect 9285 1685 9319 1719
rect 9285 1617 9319 1651
rect 9285 1567 9319 1583
rect 9353 1753 9420 1761
rect 9353 1719 9369 1753
rect 9403 1719 9420 1753
rect 9353 1685 9420 1719
rect 9353 1651 9369 1685
rect 9403 1651 9420 1685
rect 9353 1617 9420 1651
rect 9353 1583 9369 1617
rect 9403 1583 9420 1617
rect 9353 1567 9420 1583
rect 9217 1517 9256 1533
rect 9217 1483 9222 1517
rect 9217 1467 9256 1483
rect 9301 1517 9352 1533
rect 9301 1483 9318 1517
rect 9301 1467 9352 1483
rect 9301 1433 9335 1467
rect 9386 1433 9420 1567
rect 9149 1399 9335 1433
rect 9369 1404 9420 1433
rect 9149 1392 9184 1399
rect 9078 1376 9184 1392
rect 9112 1342 9184 1376
rect 9369 1380 9380 1404
rect 9414 1370 9420 1404
rect 9078 1319 9184 1342
rect 9269 1361 9335 1365
rect 9269 1327 9285 1361
rect 9319 1327 9335 1361
rect 9269 1285 9335 1327
rect 9403 1346 9420 1370
rect 9369 1319 9420 1346
rect 9586 1753 9653 1761
rect 9586 1719 9603 1753
rect 9637 1719 9653 1753
rect 9586 1685 9653 1719
rect 9586 1651 9603 1685
rect 9637 1651 9653 1685
rect 9586 1617 9653 1651
rect 9586 1583 9603 1617
rect 9637 1583 9653 1617
rect 9586 1567 9653 1583
rect 9687 1753 9721 1795
rect 9687 1685 9721 1719
rect 9687 1617 9721 1651
rect 9687 1567 9721 1583
rect 9755 1727 10161 1761
rect 9586 1433 9620 1567
rect 9755 1533 9789 1727
rect 9654 1517 9705 1533
rect 9688 1483 9705 1517
rect 9654 1467 9705 1483
rect 9750 1517 9789 1533
rect 9784 1483 9789 1517
rect 9750 1467 9789 1483
rect 9823 1659 9923 1693
rect 9957 1659 9998 1693
rect 10032 1659 10048 1693
rect 9671 1433 9705 1467
rect 9823 1433 9857 1659
rect 9586 1407 9637 1433
rect 9586 1373 9595 1407
rect 9629 1380 9637 1407
rect 9671 1399 9857 1433
rect 9891 1606 10093 1625
rect 9891 1591 10052 1606
rect 10086 1594 10093 1606
rect 9891 1481 9925 1591
rect 10055 1560 10059 1572
rect 9891 1431 9925 1447
rect 9966 1481 10021 1551
rect 9966 1447 9987 1481
rect 9586 1346 9603 1373
rect 9822 1392 9857 1399
rect 9822 1376 9928 1392
rect 9586 1319 9637 1346
rect 9671 1361 9737 1365
rect 9671 1327 9687 1361
rect 9721 1327 9737 1361
rect 9671 1285 9737 1327
rect 9822 1342 9894 1376
rect 9822 1319 9928 1342
rect 9966 1285 10021 1447
rect 10055 1319 10093 1560
rect 10127 1594 10161 1727
rect 10195 1693 10229 1795
rect 10195 1643 10229 1659
rect 10276 1693 10379 1725
rect 10276 1659 10281 1693
rect 10315 1659 10379 1693
rect 10276 1643 10379 1659
rect 10127 1592 10227 1594
rect 10127 1558 10223 1592
rect 10261 1560 10277 1594
rect 10257 1558 10277 1560
rect 10127 1556 10277 1558
rect 10311 1481 10379 1643
rect 10133 1447 10149 1481
rect 10183 1447 10379 1481
rect 11019 1693 11122 1725
rect 11019 1659 11083 1693
rect 11117 1659 11122 1693
rect 11019 1643 11122 1659
rect 11169 1693 11203 1795
rect 11169 1643 11203 1659
rect 11237 1727 11643 1761
rect 11019 1481 11087 1643
rect 11237 1594 11271 1727
rect 11350 1659 11366 1693
rect 11400 1659 11441 1693
rect 11475 1659 11575 1693
rect 11121 1591 11137 1594
rect 11121 1557 11134 1591
rect 11171 1560 11271 1594
rect 11168 1557 11271 1560
rect 11121 1556 11271 1557
rect 11305 1608 11507 1625
rect 11305 1594 11315 1608
rect 11349 1591 11507 1608
rect 11339 1560 11343 1574
rect 11019 1447 11215 1481
rect 11249 1447 11265 1481
rect 10129 1376 10231 1392
rect 10163 1342 10197 1376
rect 10129 1285 10231 1342
rect 10275 1376 10324 1447
rect 10275 1342 10281 1376
rect 10315 1342 10324 1376
rect 10275 1326 10324 1342
rect 11074 1376 11123 1447
rect 11074 1342 11083 1376
rect 11117 1342 11123 1376
rect 11074 1326 11123 1342
rect 11167 1376 11269 1392
rect 11201 1342 11235 1376
rect 11167 1285 11269 1342
rect 11305 1319 11343 1560
rect 11377 1481 11432 1551
rect 11411 1447 11432 1481
rect 11377 1285 11432 1447
rect 11473 1481 11507 1591
rect 11473 1431 11507 1447
rect 11541 1433 11575 1659
rect 11609 1533 11643 1727
rect 11677 1753 11711 1795
rect 11677 1685 11711 1719
rect 11677 1617 11711 1651
rect 11677 1567 11711 1583
rect 11745 1753 11812 1761
rect 11745 1719 11761 1753
rect 11795 1719 11812 1753
rect 11745 1685 11812 1719
rect 11745 1651 11761 1685
rect 11795 1651 11812 1685
rect 11745 1617 11812 1651
rect 11745 1583 11761 1617
rect 11795 1583 11812 1617
rect 11745 1567 11812 1583
rect 11609 1517 11648 1533
rect 11609 1483 11614 1517
rect 11609 1467 11648 1483
rect 11693 1517 11744 1533
rect 11693 1483 11710 1517
rect 11693 1467 11744 1483
rect 11693 1433 11727 1467
rect 11778 1433 11812 1567
rect 11541 1399 11727 1433
rect 11761 1406 11812 1433
rect 11541 1392 11576 1399
rect 11470 1376 11576 1392
rect 11504 1342 11576 1376
rect 11761 1380 11772 1406
rect 11806 1372 11812 1406
rect 11470 1319 11576 1342
rect 11661 1361 11727 1365
rect 11661 1327 11677 1361
rect 11711 1327 11727 1361
rect 11661 1285 11727 1327
rect 11795 1346 11812 1372
rect 11761 1319 11812 1346
rect 11978 1753 12045 1761
rect 11978 1719 11995 1753
rect 12029 1719 12045 1753
rect 11978 1685 12045 1719
rect 11978 1651 11995 1685
rect 12029 1651 12045 1685
rect 11978 1617 12045 1651
rect 11978 1583 11995 1617
rect 12029 1583 12045 1617
rect 11978 1567 12045 1583
rect 12079 1753 12113 1795
rect 12079 1685 12113 1719
rect 12079 1617 12113 1651
rect 12079 1567 12113 1583
rect 12147 1727 12553 1761
rect 11978 1433 12012 1567
rect 12147 1533 12181 1727
rect 12046 1517 12097 1533
rect 12080 1483 12097 1517
rect 12046 1467 12097 1483
rect 12142 1517 12181 1533
rect 12176 1483 12181 1517
rect 12142 1467 12181 1483
rect 12215 1659 12315 1693
rect 12349 1659 12390 1693
rect 12424 1659 12440 1693
rect 12063 1433 12097 1467
rect 12215 1433 12249 1659
rect 11978 1406 12029 1433
rect 11978 1372 11987 1406
rect 12021 1380 12029 1406
rect 12063 1399 12249 1433
rect 12283 1605 12485 1625
rect 12283 1591 12444 1605
rect 12478 1594 12485 1605
rect 12283 1481 12317 1591
rect 12447 1560 12451 1571
rect 12283 1431 12317 1447
rect 12358 1481 12413 1551
rect 12358 1447 12379 1481
rect 11978 1346 11995 1372
rect 12214 1392 12249 1399
rect 12214 1376 12320 1392
rect 11978 1319 12029 1346
rect 12063 1361 12129 1365
rect 12063 1327 12079 1361
rect 12113 1327 12129 1361
rect 12063 1285 12129 1327
rect 12214 1342 12286 1376
rect 12214 1319 12320 1342
rect 12358 1285 12413 1447
rect 12447 1319 12485 1560
rect 12519 1594 12553 1727
rect 12587 1693 12621 1795
rect 12587 1643 12621 1659
rect 12668 1693 12771 1725
rect 12668 1659 12673 1693
rect 12707 1659 12771 1693
rect 12668 1643 12771 1659
rect 12519 1592 12619 1594
rect 12519 1558 12615 1592
rect 12653 1560 12669 1594
rect 12649 1558 12669 1560
rect 12519 1556 12669 1558
rect 12703 1481 12771 1643
rect 12525 1447 12541 1481
rect 12575 1447 12771 1481
rect 13409 1693 13512 1725
rect 13409 1659 13473 1693
rect 13507 1659 13512 1693
rect 13409 1643 13512 1659
rect 13559 1693 13593 1795
rect 13559 1643 13593 1659
rect 13627 1727 14033 1761
rect 13409 1481 13477 1643
rect 13627 1594 13661 1727
rect 13740 1659 13756 1693
rect 13790 1659 13831 1693
rect 13865 1659 13965 1693
rect 13511 1591 13527 1594
rect 13511 1557 13523 1591
rect 13561 1560 13661 1594
rect 13557 1557 13661 1560
rect 13511 1556 13661 1557
rect 13695 1608 13897 1625
rect 13695 1594 13704 1608
rect 13738 1591 13897 1608
rect 13729 1560 13733 1574
rect 13409 1447 13605 1481
rect 13639 1447 13655 1481
rect 12521 1376 12623 1392
rect 12555 1342 12589 1376
rect 12521 1285 12623 1342
rect 12667 1376 12716 1447
rect 12667 1342 12673 1376
rect 12707 1342 12716 1376
rect 12667 1326 12716 1342
rect 13464 1376 13513 1447
rect 13464 1342 13473 1376
rect 13507 1342 13513 1376
rect 13464 1326 13513 1342
rect 13557 1376 13659 1392
rect 13591 1342 13625 1376
rect 13557 1285 13659 1342
rect 13695 1319 13733 1560
rect 13767 1481 13822 1551
rect 13801 1447 13822 1481
rect 13767 1285 13822 1447
rect 13863 1481 13897 1591
rect 13863 1431 13897 1447
rect 13931 1433 13965 1659
rect 13999 1533 14033 1727
rect 14067 1753 14101 1795
rect 14067 1685 14101 1719
rect 14067 1617 14101 1651
rect 14067 1567 14101 1583
rect 14135 1753 14202 1761
rect 14135 1719 14151 1753
rect 14185 1719 14202 1753
rect 14135 1685 14202 1719
rect 14135 1651 14151 1685
rect 14185 1651 14202 1685
rect 14135 1617 14202 1651
rect 14135 1583 14151 1617
rect 14185 1583 14202 1617
rect 14135 1567 14202 1583
rect 13999 1517 14038 1533
rect 13999 1483 14004 1517
rect 13999 1467 14038 1483
rect 14083 1517 14134 1533
rect 14083 1483 14100 1517
rect 14083 1467 14134 1483
rect 14083 1433 14117 1467
rect 14168 1433 14202 1567
rect 13931 1399 14117 1433
rect 14151 1404 14202 1433
rect 13931 1392 13966 1399
rect 13860 1376 13966 1392
rect 13894 1342 13966 1376
rect 14151 1380 14164 1404
rect 14198 1370 14202 1404
rect 13860 1319 13966 1342
rect 14051 1361 14117 1365
rect 14051 1327 14067 1361
rect 14101 1327 14117 1361
rect 14051 1285 14117 1327
rect 14185 1346 14202 1370
rect 14151 1319 14202 1346
rect 14370 1753 14437 1761
rect 14370 1719 14387 1753
rect 14421 1719 14437 1753
rect 14370 1685 14437 1719
rect 14370 1651 14387 1685
rect 14421 1651 14437 1685
rect 14370 1617 14437 1651
rect 14370 1583 14387 1617
rect 14421 1583 14437 1617
rect 14370 1567 14437 1583
rect 14471 1753 14505 1795
rect 14471 1685 14505 1719
rect 14471 1617 14505 1651
rect 14471 1567 14505 1583
rect 14539 1727 14945 1761
rect 14370 1433 14404 1567
rect 14539 1533 14573 1727
rect 14438 1517 14489 1533
rect 14472 1483 14489 1517
rect 14438 1467 14489 1483
rect 14534 1517 14573 1533
rect 14568 1483 14573 1517
rect 14534 1467 14573 1483
rect 14607 1659 14707 1693
rect 14741 1659 14782 1693
rect 14816 1659 14832 1693
rect 14455 1433 14489 1467
rect 14607 1433 14641 1659
rect 14370 1407 14421 1433
rect 14370 1373 14380 1407
rect 14414 1380 14421 1407
rect 14455 1399 14641 1433
rect 14675 1606 14877 1625
rect 14675 1591 14836 1606
rect 14870 1594 14877 1606
rect 14675 1481 14709 1591
rect 14839 1560 14843 1572
rect 14675 1431 14709 1447
rect 14750 1481 14805 1551
rect 14750 1447 14771 1481
rect 14370 1346 14387 1373
rect 14606 1392 14641 1399
rect 14606 1376 14712 1392
rect 14370 1319 14421 1346
rect 14455 1361 14521 1365
rect 14455 1327 14471 1361
rect 14505 1327 14521 1361
rect 14455 1285 14521 1327
rect 14606 1342 14678 1376
rect 14606 1319 14712 1342
rect 14750 1285 14805 1447
rect 14839 1319 14877 1560
rect 14911 1594 14945 1727
rect 14979 1693 15013 1795
rect 14979 1643 15013 1659
rect 15060 1693 15163 1725
rect 15060 1659 15065 1693
rect 15099 1659 15163 1693
rect 15060 1643 15163 1659
rect 14911 1592 15011 1594
rect 14911 1558 15008 1592
rect 15045 1560 15061 1594
rect 15042 1558 15061 1560
rect 14911 1556 15061 1558
rect 15095 1481 15163 1643
rect 14917 1447 14933 1481
rect 14967 1447 15163 1481
rect 15803 1693 15906 1725
rect 15803 1659 15867 1693
rect 15901 1659 15906 1693
rect 15803 1643 15906 1659
rect 15953 1693 15987 1795
rect 15953 1643 15987 1659
rect 16021 1727 16427 1761
rect 15803 1481 15871 1643
rect 16021 1594 16055 1727
rect 16134 1659 16150 1693
rect 16184 1659 16225 1693
rect 16259 1659 16359 1693
rect 15905 1592 15921 1594
rect 15905 1558 15918 1592
rect 15955 1560 16055 1594
rect 15952 1558 16055 1560
rect 15905 1556 16055 1558
rect 16089 1608 16291 1625
rect 16089 1594 16099 1608
rect 16133 1591 16291 1608
rect 16123 1560 16127 1574
rect 15803 1447 15999 1481
rect 16033 1447 16049 1481
rect 14913 1376 15015 1392
rect 14947 1342 14981 1376
rect 14913 1285 15015 1342
rect 15059 1376 15108 1447
rect 15059 1342 15065 1376
rect 15099 1342 15108 1376
rect 15059 1326 15108 1342
rect 15858 1376 15907 1447
rect 15858 1342 15867 1376
rect 15901 1342 15907 1376
rect 15858 1326 15907 1342
rect 15951 1376 16053 1392
rect 15985 1342 16019 1376
rect 15951 1285 16053 1342
rect 16089 1319 16127 1560
rect 16161 1481 16216 1551
rect 16195 1447 16216 1481
rect 16161 1285 16216 1447
rect 16257 1481 16291 1591
rect 16257 1431 16291 1447
rect 16325 1433 16359 1659
rect 16393 1533 16427 1727
rect 16461 1753 16495 1795
rect 16461 1685 16495 1719
rect 16461 1617 16495 1651
rect 16461 1567 16495 1583
rect 16529 1753 16596 1761
rect 16529 1719 16545 1753
rect 16579 1719 16596 1753
rect 16529 1685 16596 1719
rect 16529 1651 16545 1685
rect 16579 1651 16596 1685
rect 16529 1617 16596 1651
rect 16529 1583 16545 1617
rect 16579 1583 16596 1617
rect 16529 1567 16596 1583
rect 16393 1517 16432 1533
rect 16393 1483 16398 1517
rect 16393 1467 16432 1483
rect 16477 1517 16528 1533
rect 16477 1483 16494 1517
rect 16477 1467 16528 1483
rect 16477 1433 16511 1467
rect 16562 1433 16596 1567
rect 16325 1399 16511 1433
rect 16545 1406 16596 1433
rect 16325 1392 16360 1399
rect 16254 1376 16360 1392
rect 16288 1342 16360 1376
rect 16545 1380 16556 1406
rect 16590 1372 16596 1406
rect 16254 1319 16360 1342
rect 16445 1361 16511 1365
rect 16445 1327 16461 1361
rect 16495 1327 16511 1361
rect 16445 1285 16511 1327
rect 16579 1346 16596 1372
rect 16545 1319 16596 1346
rect 0 1227 29 1285
rect 63 1227 121 1285
rect 155 1227 213 1285
rect 247 1227 305 1285
rect 339 1227 397 1285
rect 431 1227 489 1285
rect 523 1227 581 1285
rect 615 1227 673 1285
rect 707 1227 765 1285
rect 799 1276 828 1285
rect 1434 1276 1463 1285
rect 799 1261 1463 1276
rect 799 1227 857 1261
rect 891 1227 949 1261
rect 983 1227 1041 1261
rect 1075 1227 1133 1261
rect 1167 1227 1225 1261
rect 1259 1227 1317 1261
rect 1351 1227 1409 1261
rect 1443 1251 1463 1261
rect 1497 1261 1555 1285
rect 1497 1251 1501 1261
rect 1443 1227 1501 1251
rect 1535 1251 1555 1261
rect 1589 1261 1647 1285
rect 1589 1251 1593 1261
rect 1535 1227 1593 1251
rect 1627 1251 1647 1261
rect 1681 1261 1739 1285
rect 1681 1251 1685 1261
rect 1627 1227 1685 1251
rect 1719 1251 1739 1261
rect 1773 1261 1831 1285
rect 1773 1251 1777 1261
rect 1719 1227 1777 1251
rect 1811 1251 1831 1261
rect 1865 1261 1923 1285
rect 1865 1251 1869 1261
rect 1811 1227 1869 1251
rect 1903 1251 1923 1261
rect 1957 1261 2015 1285
rect 1957 1251 1961 1261
rect 1903 1227 1961 1251
rect 1995 1251 2015 1261
rect 2049 1261 2107 1285
rect 2049 1251 2053 1261
rect 1995 1227 2053 1251
rect 2087 1251 2107 1261
rect 2141 1261 2199 1285
rect 2141 1251 2145 1261
rect 2087 1227 2145 1251
rect 2179 1251 2199 1261
rect 2233 1276 2262 1285
rect 2392 1276 2421 1285
rect 2233 1261 2421 1276
rect 2233 1251 2237 1261
rect 2179 1227 2237 1251
rect 2271 1227 2329 1261
rect 2363 1227 2421 1261
rect 2455 1227 2513 1285
rect 2547 1227 2605 1285
rect 2639 1227 2697 1285
rect 2731 1227 2789 1285
rect 2823 1227 2881 1285
rect 2915 1227 2973 1285
rect 3007 1227 3065 1285
rect 3099 1227 3157 1285
rect 3191 1276 3220 1285
rect 3826 1276 3855 1285
rect 3191 1261 3855 1276
rect 3191 1227 3249 1261
rect 3283 1227 3341 1261
rect 3375 1227 3433 1261
rect 3467 1227 3525 1261
rect 3559 1227 3617 1261
rect 3651 1227 3709 1261
rect 3743 1227 3801 1261
rect 3835 1251 3855 1261
rect 3889 1261 3947 1285
rect 3889 1251 3893 1261
rect 3835 1227 3893 1251
rect 3927 1251 3947 1261
rect 3981 1261 4039 1285
rect 3981 1251 3985 1261
rect 3927 1227 3985 1251
rect 4019 1251 4039 1261
rect 4073 1261 4131 1285
rect 4073 1251 4077 1261
rect 4019 1227 4077 1251
rect 4111 1251 4131 1261
rect 4165 1261 4223 1285
rect 4165 1251 4169 1261
rect 4111 1227 4169 1251
rect 4203 1251 4223 1261
rect 4257 1261 4315 1285
rect 4257 1251 4261 1261
rect 4203 1227 4261 1251
rect 4295 1251 4315 1261
rect 4349 1261 4407 1285
rect 4349 1251 4353 1261
rect 4295 1227 4353 1251
rect 4387 1251 4407 1261
rect 4441 1261 4499 1285
rect 4441 1251 4445 1261
rect 4387 1227 4445 1251
rect 4479 1251 4499 1261
rect 4533 1261 4591 1285
rect 4533 1251 4537 1261
rect 4479 1227 4537 1251
rect 4571 1251 4591 1261
rect 4625 1276 4654 1285
rect 4784 1276 4813 1285
rect 4625 1261 4813 1276
rect 4625 1251 4629 1261
rect 4571 1227 4629 1251
rect 4663 1227 4721 1261
rect 4755 1227 4813 1261
rect 4847 1227 4905 1285
rect 4939 1227 4997 1285
rect 5031 1227 5089 1285
rect 5123 1227 5181 1285
rect 5215 1227 5273 1285
rect 5307 1227 5365 1285
rect 5399 1227 5457 1285
rect 5491 1227 5549 1285
rect 5583 1276 5612 1285
rect 6216 1276 6245 1285
rect 5583 1261 6245 1276
rect 5583 1227 5641 1261
rect 5675 1227 6245 1261
rect 6279 1227 6337 1285
rect 6371 1227 6429 1285
rect 6463 1227 6521 1285
rect 6555 1227 6613 1285
rect 6647 1227 6705 1285
rect 6739 1227 6797 1285
rect 6831 1227 6889 1285
rect 6923 1227 6981 1285
rect 7015 1276 7044 1285
rect 7176 1276 7205 1285
rect 7015 1261 7205 1276
rect 7015 1227 7073 1261
rect 7107 1227 7165 1261
rect 7199 1251 7205 1261
rect 7239 1261 7297 1285
rect 7239 1251 7257 1261
rect 7199 1227 7257 1251
rect 7291 1251 7297 1261
rect 7331 1261 7389 1285
rect 7331 1251 7349 1261
rect 7291 1227 7349 1251
rect 7383 1251 7389 1261
rect 7423 1261 7481 1285
rect 7423 1251 7441 1261
rect 7383 1227 7441 1251
rect 7475 1251 7481 1261
rect 7515 1261 7573 1285
rect 7515 1251 7533 1261
rect 7475 1227 7533 1251
rect 7567 1251 7573 1261
rect 7607 1261 7665 1285
rect 7607 1251 7625 1261
rect 7567 1227 7625 1251
rect 7659 1251 7665 1261
rect 7699 1261 7757 1285
rect 7699 1251 7717 1261
rect 7659 1227 7717 1251
rect 7751 1251 7757 1261
rect 7791 1261 7849 1285
rect 7791 1251 7809 1261
rect 7751 1227 7809 1251
rect 7843 1251 7849 1261
rect 7883 1261 7941 1285
rect 7883 1251 7901 1261
rect 7843 1227 7901 1251
rect 7935 1251 7941 1261
rect 7975 1276 8004 1285
rect 8610 1276 8639 1285
rect 7975 1261 8639 1276
rect 8673 1261 8731 1285
rect 8765 1261 8823 1285
rect 8857 1261 8915 1285
rect 8949 1261 9007 1285
rect 9041 1261 9099 1285
rect 9133 1261 9191 1285
rect 9225 1261 9283 1285
rect 9317 1261 9375 1285
rect 9409 1276 9438 1285
rect 9568 1276 9597 1285
rect 9409 1261 9597 1276
rect 7975 1251 7993 1261
rect 7935 1227 7993 1251
rect 8027 1227 8085 1261
rect 8119 1227 8177 1261
rect 8211 1227 8269 1261
rect 8303 1227 8361 1261
rect 8395 1227 8453 1261
rect 8487 1227 8545 1261
rect 8579 1227 8637 1261
rect 8673 1251 8729 1261
rect 8765 1251 8821 1261
rect 8857 1251 8913 1261
rect 8949 1251 9005 1261
rect 9041 1251 9097 1261
rect 9133 1251 9189 1261
rect 9225 1251 9281 1261
rect 9317 1251 9373 1261
rect 9409 1251 9465 1261
rect 8671 1227 8729 1251
rect 8763 1227 8821 1251
rect 8855 1227 8913 1251
rect 8947 1227 9005 1251
rect 9039 1227 9097 1251
rect 9131 1227 9189 1251
rect 9223 1227 9281 1251
rect 9315 1227 9373 1251
rect 9407 1227 9465 1251
rect 9499 1227 9557 1261
rect 9591 1251 9597 1261
rect 9631 1261 9689 1285
rect 9631 1251 9649 1261
rect 9591 1227 9649 1251
rect 9683 1251 9689 1261
rect 9723 1261 9781 1285
rect 9723 1251 9741 1261
rect 9683 1227 9741 1251
rect 9775 1251 9781 1261
rect 9815 1261 9873 1285
rect 9815 1251 9833 1261
rect 9775 1227 9833 1251
rect 9867 1251 9873 1261
rect 9907 1261 9965 1285
rect 9907 1251 9925 1261
rect 9867 1227 9925 1251
rect 9959 1251 9965 1261
rect 9999 1261 10057 1285
rect 9999 1251 10017 1261
rect 9959 1227 10017 1251
rect 10051 1251 10057 1261
rect 10091 1261 10149 1285
rect 10091 1251 10109 1261
rect 10051 1227 10109 1251
rect 10143 1251 10149 1261
rect 10183 1261 10241 1285
rect 10183 1251 10201 1261
rect 10143 1227 10201 1251
rect 10235 1251 10241 1261
rect 10275 1261 10333 1285
rect 10275 1251 10293 1261
rect 10235 1227 10293 1251
rect 10327 1251 10333 1261
rect 10367 1276 10396 1285
rect 11002 1276 11031 1285
rect 10367 1261 11031 1276
rect 11065 1261 11123 1285
rect 11157 1261 11215 1285
rect 11249 1261 11307 1285
rect 11341 1261 11399 1285
rect 11433 1261 11491 1285
rect 11525 1261 11583 1285
rect 11617 1261 11675 1285
rect 11709 1261 11767 1285
rect 11801 1276 11830 1285
rect 11960 1276 11989 1285
rect 11801 1261 11989 1276
rect 12023 1261 12081 1285
rect 12115 1261 12173 1285
rect 12207 1261 12265 1285
rect 12299 1261 12357 1285
rect 12391 1261 12449 1285
rect 12483 1261 12541 1285
rect 12575 1261 12633 1285
rect 12667 1261 12725 1285
rect 12759 1276 12788 1285
rect 13392 1276 13421 1285
rect 12759 1261 13421 1276
rect 13455 1261 13513 1285
rect 13547 1261 13605 1285
rect 13639 1261 13697 1285
rect 13731 1261 13789 1285
rect 13823 1261 13881 1285
rect 13915 1261 13973 1285
rect 14007 1261 14065 1285
rect 14099 1261 14157 1285
rect 14191 1276 14220 1285
rect 14352 1276 14381 1285
rect 14191 1261 14381 1276
rect 14415 1261 14473 1285
rect 14507 1261 14565 1285
rect 14599 1261 14657 1285
rect 14691 1261 14749 1285
rect 14783 1261 14841 1285
rect 14875 1261 14933 1285
rect 14967 1261 15025 1285
rect 15059 1261 15117 1285
rect 15151 1276 15180 1285
rect 15786 1276 15815 1285
rect 15151 1261 15815 1276
rect 15849 1261 15907 1285
rect 15941 1261 15999 1285
rect 16033 1261 16091 1285
rect 16125 1261 16183 1285
rect 16217 1261 16275 1285
rect 16309 1261 16367 1285
rect 16401 1261 16459 1285
rect 16493 1261 16551 1285
rect 10367 1251 10385 1261
rect 10327 1227 10385 1251
rect 10419 1227 10477 1261
rect 10511 1227 10569 1261
rect 10603 1227 10661 1261
rect 10695 1227 10753 1261
rect 10787 1227 10845 1261
rect 10879 1227 10937 1261
rect 10971 1227 11029 1261
rect 11065 1251 11121 1261
rect 11157 1251 11213 1261
rect 11249 1251 11305 1261
rect 11341 1251 11397 1261
rect 11433 1251 11489 1261
rect 11525 1251 11581 1261
rect 11617 1251 11673 1261
rect 11709 1251 11765 1261
rect 11801 1251 11857 1261
rect 11063 1227 11121 1251
rect 11155 1227 11213 1251
rect 11247 1227 11305 1251
rect 11339 1227 11397 1251
rect 11431 1227 11489 1251
rect 11523 1227 11581 1251
rect 11615 1227 11673 1251
rect 11707 1227 11765 1251
rect 11799 1227 11857 1251
rect 11891 1251 11989 1261
rect 12045 1251 12081 1261
rect 12137 1251 12173 1261
rect 12229 1251 12265 1261
rect 12321 1251 12357 1261
rect 12413 1251 12449 1261
rect 12505 1251 12541 1261
rect 12597 1251 12633 1261
rect 12689 1251 12725 1261
rect 11891 1227 12011 1251
rect 12045 1227 12103 1251
rect 12137 1227 12195 1251
rect 12229 1227 12287 1251
rect 12321 1227 12379 1251
rect 12413 1227 12471 1251
rect 12505 1227 12563 1251
rect 12597 1227 12655 1251
rect 12689 1227 12747 1251
rect 12781 1227 12839 1261
rect 12873 1227 12931 1261
rect 12965 1227 13023 1261
rect 13057 1227 13115 1261
rect 13149 1227 13207 1261
rect 13241 1227 13299 1261
rect 13333 1227 13391 1261
rect 13455 1251 13483 1261
rect 13547 1251 13575 1261
rect 13639 1251 13667 1261
rect 13731 1251 13759 1261
rect 13823 1251 13851 1261
rect 13915 1251 13943 1261
rect 14007 1251 14035 1261
rect 14099 1251 14127 1261
rect 14191 1251 14219 1261
rect 13425 1227 13483 1251
rect 13517 1227 13575 1251
rect 13609 1227 13667 1251
rect 13701 1227 13759 1251
rect 13793 1227 13851 1251
rect 13885 1227 13943 1251
rect 13977 1227 14035 1251
rect 14069 1227 14127 1251
rect 14161 1227 14219 1251
rect 14253 1227 14311 1261
rect 14345 1251 14381 1261
rect 14437 1251 14473 1261
rect 14529 1251 14565 1261
rect 14621 1251 14657 1261
rect 14713 1251 14749 1261
rect 14805 1251 14841 1261
rect 14897 1251 14933 1261
rect 14989 1251 15025 1261
rect 15081 1251 15117 1261
rect 14345 1227 14403 1251
rect 14437 1227 14495 1251
rect 14529 1227 14587 1251
rect 14621 1227 14679 1251
rect 14713 1227 14771 1251
rect 14805 1227 14863 1251
rect 14897 1227 14955 1251
rect 14989 1227 15047 1251
rect 15081 1227 15139 1251
rect 15173 1227 15231 1261
rect 15265 1227 15323 1261
rect 15357 1227 15415 1261
rect 15449 1227 15507 1261
rect 15541 1227 15599 1261
rect 15633 1227 15691 1261
rect 15725 1227 15783 1261
rect 15849 1251 15875 1261
rect 15941 1251 15967 1261
rect 16033 1251 16059 1261
rect 16125 1251 16151 1261
rect 16217 1251 16243 1261
rect 16309 1251 16335 1261
rect 16401 1251 16427 1261
rect 16493 1251 16519 1261
rect 16585 1251 16614 1285
rect 15817 1227 15875 1251
rect 15909 1227 15967 1251
rect 16001 1227 16059 1251
rect 16093 1227 16151 1251
rect 16185 1227 16243 1251
rect 16277 1227 16335 1251
rect 16369 1227 16427 1251
rect 16461 1227 16519 1251
rect 16553 1227 16614 1251
rect 16237 1165 16303 1173
rect 0 1107 29 1165
rect 63 1107 121 1165
rect 155 1107 213 1165
rect 247 1107 305 1165
rect 339 1107 397 1165
rect 431 1107 489 1165
rect 523 1107 581 1165
rect 615 1107 673 1165
rect 707 1107 765 1165
rect 799 1107 857 1165
rect 891 1107 949 1165
rect 983 1107 1041 1165
rect 1075 1107 1133 1165
rect 1167 1107 1225 1165
rect 1259 1107 1317 1165
rect 1351 1107 1409 1165
rect 1443 1107 1501 1165
rect 1535 1107 1593 1165
rect 1627 1107 1685 1165
rect 1719 1107 1777 1165
rect 1811 1158 2053 1165
rect 1811 1141 1901 1158
rect 1935 1141 2053 1158
rect 1811 1107 1869 1141
rect 1935 1124 1961 1141
rect 1903 1107 1961 1124
rect 1995 1107 2053 1141
rect 2087 1107 2145 1165
rect 2179 1107 2237 1165
rect 2271 1107 2329 1165
rect 2363 1107 2421 1165
rect 2455 1107 2513 1165
rect 2547 1107 2605 1165
rect 2639 1107 2697 1165
rect 2731 1107 2789 1165
rect 2823 1107 2881 1165
rect 2915 1107 2973 1165
rect 3007 1107 3065 1165
rect 3099 1107 3157 1165
rect 3191 1107 3249 1165
rect 3283 1107 3341 1165
rect 3375 1107 3433 1165
rect 3467 1107 3525 1165
rect 3559 1107 3617 1165
rect 3651 1107 3709 1165
rect 3743 1107 3801 1165
rect 3835 1107 3893 1165
rect 3927 1107 3985 1165
rect 4019 1107 4077 1165
rect 4111 1107 4169 1165
rect 4203 1157 4445 1165
rect 4203 1141 4293 1157
rect 4327 1141 4445 1157
rect 4203 1107 4261 1141
rect 4327 1123 4353 1141
rect 4295 1107 4353 1123
rect 4387 1107 4445 1141
rect 4479 1107 4537 1165
rect 4571 1107 4629 1165
rect 4663 1107 4721 1165
rect 4755 1107 4813 1165
rect 4847 1107 4905 1165
rect 4939 1107 4997 1165
rect 5031 1107 5089 1165
rect 5123 1107 5181 1165
rect 5215 1107 5273 1165
rect 5307 1107 5365 1165
rect 5399 1107 5457 1165
rect 5491 1107 5549 1165
rect 5583 1107 5641 1165
rect 5675 1107 5733 1165
rect 5767 1107 5825 1165
rect 5859 1107 5917 1165
rect 5951 1107 6009 1165
rect 6043 1107 6101 1165
rect 6135 1107 6193 1165
rect 6227 1107 6285 1165
rect 6319 1107 6377 1165
rect 6411 1107 6469 1165
rect 6503 1107 6561 1165
rect 6595 1157 6837 1165
rect 6595 1141 6685 1157
rect 6719 1141 6837 1157
rect 6595 1107 6653 1141
rect 6719 1123 6745 1141
rect 6687 1107 6745 1123
rect 6779 1107 6837 1141
rect 6871 1107 6929 1165
rect 6963 1107 7021 1165
rect 7055 1107 7113 1165
rect 7147 1107 7205 1165
rect 7239 1107 7297 1165
rect 7331 1107 7389 1165
rect 7423 1107 7481 1165
rect 7515 1107 7573 1165
rect 7607 1107 7665 1165
rect 7699 1107 7757 1165
rect 7791 1107 7849 1165
rect 7883 1107 7941 1165
rect 7975 1107 8033 1165
rect 8067 1107 8125 1165
rect 8159 1107 8217 1165
rect 8251 1107 8309 1165
rect 8343 1107 8401 1165
rect 8435 1107 8493 1165
rect 8527 1107 8585 1165
rect 8619 1107 8677 1165
rect 8711 1107 8769 1165
rect 8803 1107 8861 1165
rect 8895 1107 8953 1165
rect 8987 1158 9229 1165
rect 8987 1141 9077 1158
rect 9111 1141 9229 1158
rect 8987 1107 9045 1141
rect 9111 1124 9137 1141
rect 9079 1107 9137 1124
rect 9171 1107 9229 1141
rect 9263 1107 9321 1165
rect 9355 1107 9413 1165
rect 9447 1107 9505 1165
rect 9539 1107 9597 1165
rect 9631 1107 9689 1165
rect 9723 1107 9781 1165
rect 9815 1107 9873 1165
rect 9907 1107 9965 1165
rect 9999 1107 10057 1165
rect 10091 1107 10149 1165
rect 10183 1107 10241 1165
rect 10275 1107 10333 1165
rect 10367 1107 10425 1165
rect 10459 1107 10517 1165
rect 10551 1107 10609 1165
rect 10643 1107 10701 1165
rect 10735 1107 10793 1165
rect 10827 1107 10885 1165
rect 10919 1107 10977 1165
rect 11011 1107 11069 1165
rect 11103 1107 11161 1165
rect 11195 1107 11253 1165
rect 11287 1107 11345 1165
rect 11379 1158 11621 1165
rect 11379 1141 11469 1158
rect 11503 1141 11621 1158
rect 11379 1107 11437 1141
rect 11503 1124 11529 1141
rect 11471 1107 11529 1124
rect 11563 1107 11621 1141
rect 11655 1107 11713 1165
rect 11747 1107 11805 1165
rect 11839 1107 11897 1165
rect 11931 1107 11989 1165
rect 12023 1107 12081 1165
rect 12115 1107 12173 1165
rect 12207 1107 12265 1165
rect 12299 1107 12357 1165
rect 12391 1107 12449 1165
rect 12483 1107 12541 1165
rect 12575 1107 12633 1165
rect 12667 1107 12725 1165
rect 12759 1107 12817 1165
rect 12851 1107 12909 1165
rect 12943 1107 13001 1165
rect 13035 1107 13093 1165
rect 13127 1107 13185 1165
rect 13219 1107 13277 1165
rect 13311 1107 13369 1165
rect 13403 1107 13461 1165
rect 13495 1107 13553 1165
rect 13587 1107 13645 1165
rect 13679 1107 13737 1165
rect 13771 1157 14013 1165
rect 13771 1141 13861 1157
rect 13895 1141 14013 1157
rect 13771 1107 13829 1141
rect 13895 1123 13921 1141
rect 13863 1107 13921 1123
rect 13955 1107 14013 1141
rect 14047 1107 14105 1165
rect 14139 1107 14197 1165
rect 14231 1107 14289 1165
rect 14323 1107 14381 1165
rect 14415 1107 14473 1165
rect 14507 1107 14565 1165
rect 14599 1107 14657 1165
rect 14691 1107 14749 1165
rect 14783 1107 14841 1165
rect 14875 1107 14933 1165
rect 14967 1107 15025 1165
rect 15059 1107 15117 1165
rect 15151 1107 15209 1165
rect 15243 1107 15301 1165
rect 15335 1107 15393 1165
rect 15427 1107 15485 1165
rect 15519 1107 15577 1165
rect 15611 1107 15669 1165
rect 15703 1107 15761 1165
rect 15795 1107 15853 1165
rect 15887 1107 15945 1165
rect 15979 1107 16037 1165
rect 16071 1107 16129 1165
rect 16163 1157 16405 1165
rect 16163 1141 16253 1157
rect 16287 1141 16405 1157
rect 16163 1107 16221 1141
rect 16287 1123 16313 1141
rect 16255 1107 16313 1123
rect 16347 1107 16405 1141
rect 16439 1107 16497 1165
rect 16531 1107 16589 1165
rect 16623 1107 16681 1165
rect 16715 1107 16744 1165
rect 35 1057 69 1073
rect 35 989 69 1023
rect 103 1041 169 1107
rect 103 1007 119 1041
rect 153 1007 169 1041
rect 203 1057 247 1073
rect 237 1023 247 1057
rect 203 989 247 1023
rect 286 1041 357 1107
rect 286 1007 307 1041
rect 341 1007 357 1041
rect 391 1057 425 1073
rect 467 1030 483 1064
rect 517 1030 633 1064
rect 69 955 168 973
rect 35 939 168 955
rect 17 859 87 905
rect 17 825 26 859
rect 60 844 87 859
rect 17 810 31 825
rect 65 810 87 844
rect 17 775 87 810
rect 122 844 168 939
rect 122 810 133 844
rect 167 810 168 844
rect 122 767 168 810
rect 35 733 122 741
rect 156 733 168 767
rect 35 707 168 733
rect 237 971 247 989
rect 391 973 425 1023
rect 203 937 213 955
rect 35 699 69 707
rect 203 699 247 937
rect 281 939 425 973
rect 281 745 315 939
rect 465 937 489 971
rect 523 945 565 971
rect 523 937 531 945
rect 465 911 531 937
rect 349 883 431 905
rect 349 849 366 883
rect 400 849 431 883
rect 349 831 431 849
rect 383 797 431 831
rect 349 781 431 797
rect 465 895 565 911
rect 465 771 509 895
rect 599 861 633 1030
rect 681 1055 757 1107
rect 975 1065 1041 1107
rect 681 1021 697 1055
rect 731 1021 757 1055
rect 817 1039 851 1055
rect 817 987 851 1005
rect 975 1031 991 1065
rect 1025 1031 1041 1065
rect 1464 1065 1540 1107
rect 975 997 1041 1031
rect 1250 1030 1266 1064
rect 1300 1030 1416 1064
rect 1464 1031 1480 1065
rect 1514 1031 1540 1065
rect 1728 1065 2006 1107
rect 1588 1039 1622 1055
rect 667 971 937 987
rect 667 945 817 971
rect 701 937 817 945
rect 851 937 937 971
rect 975 963 991 997
rect 1025 963 1041 997
rect 1212 971 1259 977
rect 701 911 717 937
rect 667 895 717 911
rect 819 861 869 877
rect 599 827 835 861
rect 599 819 683 827
rect 281 707 425 745
rect 499 737 509 771
rect 465 721 509 737
rect 545 749 561 783
rect 595 767 615 783
rect 545 733 581 749
rect 545 709 615 733
rect 35 649 69 665
rect 103 639 119 673
rect 153 639 169 673
rect 237 665 247 699
rect 391 691 425 707
rect 203 649 247 665
rect 103 597 169 639
rect 286 639 307 673
rect 341 639 357 673
rect 649 673 683 819
rect 825 811 869 827
rect 903 793 937 937
rect 1212 945 1225 971
rect 1246 911 1259 937
rect 971 903 1172 911
rect 971 869 1133 903
rect 1167 869 1172 903
rect 1212 895 1259 911
rect 1307 945 1348 961
rect 1307 911 1314 945
rect 971 863 1172 869
rect 971 861 1037 863
rect 971 827 987 861
rect 1021 827 1037 861
rect 1307 841 1348 911
rect 1213 835 1348 841
rect 1099 793 1115 827
rect 1149 793 1165 827
rect 717 759 733 793
rect 767 773 783 793
rect 767 767 799 773
rect 717 733 765 759
rect 903 759 1165 793
rect 1213 801 1225 835
rect 1259 805 1348 835
rect 1382 861 1416 1030
rect 1728 1031 1754 1065
rect 1788 1031 1956 1065
rect 1990 1031 2006 1065
rect 1588 997 1622 1005
rect 2040 1028 2097 1073
rect 1450 963 2006 997
rect 1450 945 1500 963
rect 1484 911 1500 945
rect 1450 895 1500 911
rect 1382 845 1652 861
rect 1382 827 1618 845
rect 1259 801 1281 805
rect 1213 792 1281 801
rect 1237 771 1281 792
rect 903 733 947 759
rect 717 727 799 733
rect 881 699 897 733
rect 931 699 947 733
rect 1237 737 1247 771
rect 981 707 1015 723
rect 1237 721 1281 737
rect 391 641 425 657
rect 286 597 357 639
rect 480 639 496 673
rect 530 639 683 673
rect 480 633 683 639
rect 717 669 751 685
rect 717 597 751 635
rect 785 675 851 681
rect 785 641 801 675
rect 835 665 851 675
rect 1382 673 1416 827
rect 1608 811 1618 827
rect 1608 795 1652 811
rect 1456 759 1511 793
rect 1545 767 1565 793
rect 1456 733 1515 759
rect 1549 733 1565 767
rect 1686 748 1720 963
rect 1754 903 1858 929
rect 1754 869 1771 903
rect 1805 895 1858 903
rect 1892 895 1911 929
rect 1805 869 1811 895
rect 1754 861 1811 869
rect 1788 827 1811 861
rect 1972 845 2006 963
rect 2074 994 2097 1028
rect 2040 960 2097 994
rect 2074 955 2097 960
rect 2040 921 2051 926
rect 2085 921 2097 955
rect 2040 906 2097 921
rect 1754 802 1811 827
rect 1767 765 1811 802
rect 1847 833 1938 845
rect 1847 799 1863 833
rect 1897 799 1938 833
rect 1972 829 2025 845
rect 1972 795 1991 829
rect 1972 779 2025 795
rect 1686 747 1723 748
rect 1456 727 1565 733
rect 1643 713 1673 747
rect 1707 713 1723 747
rect 1767 731 1895 765
rect 981 665 1015 673
rect 835 641 1015 665
rect 785 631 1015 641
rect 1065 639 1085 673
rect 1119 639 1135 673
rect 1065 597 1135 639
rect 1260 639 1289 673
rect 1323 639 1416 673
rect 1260 633 1416 639
rect 1450 669 1515 685
rect 1450 635 1481 669
rect 1450 597 1515 635
rect 1549 655 1565 689
rect 1599 665 1615 689
rect 1757 681 1791 697
rect 1599 655 1757 665
rect 1549 647 1757 655
rect 1549 631 1791 647
rect 1853 683 1895 731
rect 1853 649 1861 683
rect 1853 633 1895 649
rect 1945 673 2006 741
rect 2061 723 2097 906
rect 1945 639 1956 673
rect 1990 639 2006 673
rect 1945 597 2006 639
rect 2040 707 2097 723
rect 2074 673 2097 707
rect 2040 631 2097 673
rect 2132 1047 2195 1063
rect 2132 1013 2144 1047
rect 2178 1013 2195 1047
rect 2132 979 2195 1013
rect 2132 945 2144 979
rect 2178 945 2195 979
rect 2132 845 2195 945
rect 2231 1053 2289 1107
rect 2231 1019 2239 1053
rect 2273 1019 2289 1053
rect 2231 985 2289 1019
rect 2231 951 2239 985
rect 2273 951 2289 985
rect 2231 933 2289 951
rect 2323 1034 2375 1073
rect 2323 1029 2334 1034
rect 2368 1000 2375 1034
rect 2357 995 2375 1000
rect 2323 961 2375 995
rect 2357 927 2375 961
rect 2427 1057 2461 1073
rect 2427 989 2461 1023
rect 2495 1041 2561 1107
rect 2495 1007 2511 1041
rect 2545 1007 2561 1041
rect 2595 1057 2639 1073
rect 2629 1023 2639 1057
rect 2595 989 2639 1023
rect 2678 1041 2749 1107
rect 2678 1007 2699 1041
rect 2733 1007 2749 1041
rect 2783 1057 2817 1073
rect 2859 1030 2875 1064
rect 2909 1030 3025 1064
rect 2461 955 2560 973
rect 2427 939 2560 955
rect 2323 871 2375 927
rect 2132 829 2299 845
rect 2132 795 2265 829
rect 2132 779 2299 795
rect 2132 699 2195 779
rect 2333 745 2375 871
rect 2409 859 2479 905
rect 2409 825 2418 859
rect 2452 844 2479 859
rect 2409 810 2423 825
rect 2457 810 2479 844
rect 2409 775 2479 810
rect 2514 844 2560 939
rect 2514 810 2525 844
rect 2559 810 2560 844
rect 2132 665 2144 699
rect 2178 665 2195 699
rect 2323 709 2375 745
rect 2514 767 2560 810
rect 2132 631 2195 665
rect 2230 673 2289 689
rect 2230 639 2239 673
rect 2273 639 2289 673
rect 2230 597 2289 639
rect 2357 675 2375 709
rect 2323 631 2375 675
rect 2427 733 2514 741
rect 2548 733 2560 767
rect 2427 707 2560 733
rect 2629 971 2639 989
rect 2783 973 2817 1023
rect 2595 937 2605 955
rect 2427 699 2461 707
rect 2595 699 2639 937
rect 2673 939 2817 973
rect 2673 745 2707 939
rect 2857 937 2881 971
rect 2915 945 2957 971
rect 2915 937 2923 945
rect 2857 911 2923 937
rect 2741 883 2823 905
rect 2741 849 2758 883
rect 2792 849 2823 883
rect 2741 831 2823 849
rect 2775 797 2823 831
rect 2741 781 2823 797
rect 2857 895 2957 911
rect 2857 771 2901 895
rect 2991 861 3025 1030
rect 3073 1055 3149 1107
rect 3367 1065 3433 1107
rect 3073 1021 3089 1055
rect 3123 1021 3149 1055
rect 3209 1039 3243 1055
rect 3209 987 3243 1005
rect 3367 1031 3383 1065
rect 3417 1031 3433 1065
rect 3856 1065 3932 1107
rect 3367 997 3433 1031
rect 3642 1030 3658 1064
rect 3692 1030 3808 1064
rect 3856 1031 3872 1065
rect 3906 1031 3932 1065
rect 4120 1065 4398 1107
rect 3980 1039 4014 1055
rect 3059 971 3329 987
rect 3059 945 3209 971
rect 3093 937 3209 945
rect 3243 937 3329 971
rect 3367 963 3383 997
rect 3417 963 3433 997
rect 3604 971 3651 977
rect 3093 911 3109 937
rect 3059 895 3109 911
rect 3211 861 3261 877
rect 2991 827 3227 861
rect 2991 819 3075 827
rect 2673 707 2817 745
rect 2891 737 2901 771
rect 2857 721 2901 737
rect 2937 749 2953 783
rect 2987 767 3007 783
rect 2937 733 2973 749
rect 2937 709 3007 733
rect 2427 649 2461 665
rect 2495 639 2511 673
rect 2545 639 2561 673
rect 2629 665 2639 699
rect 2783 691 2817 707
rect 2595 649 2639 665
rect 2495 597 2561 639
rect 2678 639 2699 673
rect 2733 639 2749 673
rect 3041 673 3075 819
rect 3217 811 3261 827
rect 3295 793 3329 937
rect 3604 945 3617 971
rect 3638 911 3651 937
rect 3363 903 3564 911
rect 3363 869 3525 903
rect 3559 869 3564 903
rect 3604 895 3651 911
rect 3699 945 3740 961
rect 3699 911 3706 945
rect 3363 863 3564 869
rect 3363 861 3429 863
rect 3363 827 3379 861
rect 3413 827 3429 861
rect 3699 841 3740 911
rect 3605 835 3740 841
rect 3491 793 3507 827
rect 3541 793 3557 827
rect 3109 759 3125 793
rect 3159 773 3175 793
rect 3159 767 3191 773
rect 3109 733 3157 759
rect 3295 759 3557 793
rect 3605 801 3617 835
rect 3651 805 3740 835
rect 3774 861 3808 1030
rect 4120 1031 4146 1065
rect 4180 1031 4348 1065
rect 4382 1031 4398 1065
rect 3980 997 4014 1005
rect 4432 1028 4489 1073
rect 3842 963 4398 997
rect 3842 945 3892 963
rect 3876 911 3892 945
rect 3842 895 3892 911
rect 3774 845 4044 861
rect 3774 827 4010 845
rect 3651 801 3673 805
rect 3605 792 3673 801
rect 3629 771 3673 792
rect 3295 733 3339 759
rect 3109 727 3191 733
rect 3273 699 3289 733
rect 3323 699 3339 733
rect 3629 737 3639 771
rect 3373 707 3407 723
rect 3629 721 3673 737
rect 2783 641 2817 657
rect 2678 597 2749 639
rect 2872 639 2888 673
rect 2922 639 3075 673
rect 2872 633 3075 639
rect 3109 669 3143 685
rect 3109 597 3143 635
rect 3177 675 3243 681
rect 3177 641 3193 675
rect 3227 665 3243 675
rect 3774 673 3808 827
rect 4000 811 4010 827
rect 4000 795 4044 811
rect 3848 759 3903 793
rect 3937 767 3957 793
rect 3848 733 3907 759
rect 3941 733 3957 767
rect 4078 748 4112 963
rect 4146 903 4250 929
rect 4146 869 4163 903
rect 4197 895 4250 903
rect 4284 895 4303 929
rect 4197 869 4203 895
rect 4146 861 4203 869
rect 4180 827 4203 861
rect 4364 845 4398 963
rect 4466 994 4489 1028
rect 4432 960 4489 994
rect 4466 956 4489 960
rect 4432 922 4443 926
rect 4477 922 4489 956
rect 4432 906 4489 922
rect 4146 802 4203 827
rect 4159 765 4203 802
rect 4239 833 4330 845
rect 4239 799 4255 833
rect 4289 799 4330 833
rect 4364 829 4417 845
rect 4364 795 4383 829
rect 4364 779 4417 795
rect 4078 747 4115 748
rect 3848 727 3957 733
rect 4035 713 4065 747
rect 4099 713 4115 747
rect 4159 731 4287 765
rect 3373 665 3407 673
rect 3227 641 3407 665
rect 3177 631 3407 641
rect 3457 639 3477 673
rect 3511 639 3527 673
rect 3457 597 3527 639
rect 3652 639 3681 673
rect 3715 639 3808 673
rect 3652 633 3808 639
rect 3842 669 3907 685
rect 3842 635 3873 669
rect 3842 597 3907 635
rect 3941 655 3957 689
rect 3991 665 4007 689
rect 4149 681 4183 697
rect 3991 655 4149 665
rect 3941 647 4149 655
rect 3941 631 4183 647
rect 4245 683 4287 731
rect 4245 649 4253 683
rect 4245 633 4287 649
rect 4337 673 4398 741
rect 4453 723 4489 906
rect 4337 639 4348 673
rect 4382 639 4398 673
rect 4337 597 4398 639
rect 4432 707 4489 723
rect 4466 673 4489 707
rect 4432 631 4489 673
rect 4524 1047 4587 1063
rect 4524 1013 4536 1047
rect 4570 1013 4587 1047
rect 4524 979 4587 1013
rect 4524 945 4536 979
rect 4570 945 4587 979
rect 4524 845 4587 945
rect 4623 1053 4681 1107
rect 4623 1019 4631 1053
rect 4665 1019 4681 1053
rect 4623 985 4681 1019
rect 4623 951 4631 985
rect 4665 951 4681 985
rect 4623 933 4681 951
rect 4715 1034 4767 1073
rect 4715 1029 4726 1034
rect 4760 1000 4767 1034
rect 4749 995 4767 1000
rect 4715 961 4767 995
rect 4749 927 4767 961
rect 4819 1057 4853 1073
rect 4819 989 4853 1023
rect 4887 1041 4953 1107
rect 4887 1007 4903 1041
rect 4937 1007 4953 1041
rect 4987 1057 5031 1073
rect 5021 1023 5031 1057
rect 4987 989 5031 1023
rect 5070 1041 5141 1107
rect 5070 1007 5091 1041
rect 5125 1007 5141 1041
rect 5175 1057 5209 1073
rect 5251 1030 5267 1064
rect 5301 1030 5417 1064
rect 4853 955 4952 973
rect 4819 939 4952 955
rect 4715 871 4767 927
rect 4524 829 4691 845
rect 4524 795 4657 829
rect 4524 779 4691 795
rect 4524 699 4587 779
rect 4725 745 4767 871
rect 4801 859 4871 905
rect 4801 825 4810 859
rect 4844 844 4871 859
rect 4801 810 4815 825
rect 4849 810 4871 844
rect 4801 775 4871 810
rect 4906 844 4952 939
rect 4906 810 4917 844
rect 4951 810 4952 844
rect 4524 665 4536 699
rect 4570 665 4587 699
rect 4715 709 4767 745
rect 4906 767 4952 810
rect 4524 631 4587 665
rect 4622 673 4681 689
rect 4622 639 4631 673
rect 4665 639 4681 673
rect 4622 597 4681 639
rect 4749 675 4767 709
rect 4715 631 4767 675
rect 4819 733 4906 741
rect 4940 733 4952 767
rect 4819 707 4952 733
rect 5021 971 5031 989
rect 5175 973 5209 1023
rect 4987 937 4997 955
rect 4819 699 4853 707
rect 4987 699 5031 937
rect 5065 939 5209 973
rect 5065 745 5099 939
rect 5249 937 5273 971
rect 5307 945 5349 971
rect 5307 937 5315 945
rect 5249 911 5315 937
rect 5133 884 5215 905
rect 5133 850 5150 884
rect 5184 850 5215 884
rect 5133 831 5215 850
rect 5167 797 5215 831
rect 5133 781 5215 797
rect 5249 895 5349 911
rect 5249 771 5293 895
rect 5383 861 5417 1030
rect 5465 1055 5541 1107
rect 5759 1065 5825 1107
rect 5465 1021 5481 1055
rect 5515 1021 5541 1055
rect 5601 1039 5635 1055
rect 5601 987 5635 1005
rect 5759 1031 5775 1065
rect 5809 1031 5825 1065
rect 6248 1065 6324 1107
rect 5759 997 5825 1031
rect 6034 1030 6050 1064
rect 6084 1030 6200 1064
rect 6248 1031 6264 1065
rect 6298 1031 6324 1065
rect 6512 1065 6790 1107
rect 6372 1039 6406 1055
rect 5451 971 5721 987
rect 5451 945 5601 971
rect 5485 937 5601 945
rect 5635 937 5721 971
rect 5759 963 5775 997
rect 5809 963 5825 997
rect 5996 971 6043 977
rect 5485 911 5501 937
rect 5451 895 5501 911
rect 5603 861 5653 877
rect 5383 827 5619 861
rect 5383 819 5467 827
rect 5065 707 5209 745
rect 5283 737 5293 771
rect 5249 721 5293 737
rect 5329 749 5345 783
rect 5379 767 5399 783
rect 5329 733 5365 749
rect 5329 709 5399 733
rect 4819 649 4853 665
rect 4887 639 4903 673
rect 4937 639 4953 673
rect 5021 665 5031 699
rect 5175 691 5209 707
rect 4987 649 5031 665
rect 4887 597 4953 639
rect 5070 639 5091 673
rect 5125 639 5141 673
rect 5433 673 5467 819
rect 5609 811 5653 827
rect 5687 793 5721 937
rect 5996 945 6009 971
rect 6030 911 6043 937
rect 5755 903 5956 911
rect 5755 869 5917 903
rect 5951 869 5956 903
rect 5996 895 6043 911
rect 6091 945 6132 961
rect 6091 911 6098 945
rect 5755 863 5956 869
rect 5755 861 5821 863
rect 5755 827 5771 861
rect 5805 827 5821 861
rect 6091 841 6132 911
rect 5997 835 6132 841
rect 5883 793 5899 827
rect 5933 793 5949 827
rect 5501 759 5517 793
rect 5551 773 5567 793
rect 5551 767 5583 773
rect 5501 733 5549 759
rect 5687 759 5949 793
rect 5997 801 6009 835
rect 6043 805 6132 835
rect 6166 861 6200 1030
rect 6512 1031 6538 1065
rect 6572 1031 6740 1065
rect 6774 1031 6790 1065
rect 6372 997 6406 1005
rect 6824 1028 6881 1073
rect 6234 963 6790 997
rect 6234 945 6284 963
rect 6268 911 6284 945
rect 6234 895 6284 911
rect 6166 845 6436 861
rect 6166 827 6402 845
rect 6043 801 6065 805
rect 5997 792 6065 801
rect 6021 771 6065 792
rect 5687 733 5731 759
rect 5501 727 5583 733
rect 5665 699 5681 733
rect 5715 699 5731 733
rect 6021 737 6031 771
rect 5765 707 5799 723
rect 6021 721 6065 737
rect 5175 641 5209 657
rect 5070 597 5141 639
rect 5264 639 5280 673
rect 5314 639 5467 673
rect 5264 633 5467 639
rect 5501 669 5535 685
rect 5501 597 5535 635
rect 5569 675 5635 681
rect 5569 641 5585 675
rect 5619 665 5635 675
rect 6166 673 6200 827
rect 6392 811 6402 827
rect 6392 795 6436 811
rect 6240 759 6295 793
rect 6329 767 6349 793
rect 6240 733 6299 759
rect 6333 733 6349 767
rect 6470 748 6504 963
rect 6538 903 6642 929
rect 6538 869 6555 903
rect 6589 895 6642 903
rect 6676 895 6695 929
rect 6589 869 6595 895
rect 6538 861 6595 869
rect 6572 827 6595 861
rect 6756 845 6790 963
rect 6858 994 6881 1028
rect 6824 960 6881 994
rect 6858 956 6881 960
rect 6824 922 6834 926
rect 6868 922 6881 956
rect 6824 906 6881 922
rect 6538 802 6595 827
rect 6551 765 6595 802
rect 6631 833 6722 845
rect 6631 799 6647 833
rect 6681 799 6722 833
rect 6756 829 6809 845
rect 6756 795 6775 829
rect 6756 779 6809 795
rect 6470 747 6507 748
rect 6240 727 6349 733
rect 6427 713 6457 747
rect 6491 713 6507 747
rect 6551 731 6679 765
rect 5765 665 5799 673
rect 5619 641 5799 665
rect 5569 631 5799 641
rect 5849 639 5869 673
rect 5903 639 5919 673
rect 5849 597 5919 639
rect 6044 639 6073 673
rect 6107 639 6200 673
rect 6044 633 6200 639
rect 6234 669 6299 685
rect 6234 635 6265 669
rect 6234 597 6299 635
rect 6333 655 6349 689
rect 6383 665 6399 689
rect 6541 681 6575 697
rect 6383 655 6541 665
rect 6333 647 6541 655
rect 6333 631 6575 647
rect 6637 683 6679 731
rect 6637 649 6645 683
rect 6637 633 6679 649
rect 6729 673 6790 741
rect 6845 723 6881 906
rect 6729 639 6740 673
rect 6774 639 6790 673
rect 6729 597 6790 639
rect 6824 707 6881 723
rect 6858 673 6881 707
rect 6824 631 6881 673
rect 6916 1047 6979 1063
rect 6916 1013 6928 1047
rect 6962 1013 6979 1047
rect 6916 979 6979 1013
rect 6916 945 6928 979
rect 6962 945 6979 979
rect 6916 845 6979 945
rect 7015 1053 7073 1107
rect 7015 1019 7023 1053
rect 7057 1019 7073 1053
rect 7015 985 7073 1019
rect 7015 951 7023 985
rect 7057 951 7073 985
rect 7015 933 7073 951
rect 7107 1034 7159 1073
rect 7107 1029 7118 1034
rect 7152 1000 7159 1034
rect 7141 995 7159 1000
rect 7107 961 7159 995
rect 7141 927 7159 961
rect 7211 1057 7245 1073
rect 7211 989 7245 1023
rect 7279 1041 7345 1107
rect 7279 1007 7295 1041
rect 7329 1007 7345 1041
rect 7379 1057 7423 1073
rect 7413 1023 7423 1057
rect 7379 989 7423 1023
rect 7462 1041 7533 1107
rect 7462 1007 7483 1041
rect 7517 1007 7533 1041
rect 7567 1057 7601 1073
rect 7643 1030 7659 1064
rect 7693 1030 7809 1064
rect 7245 955 7344 973
rect 7211 939 7344 955
rect 7107 871 7159 927
rect 6916 829 7083 845
rect 6916 795 7049 829
rect 6916 779 7083 795
rect 6916 699 6979 779
rect 7117 745 7159 871
rect 7193 859 7263 905
rect 7193 825 7202 859
rect 7236 844 7263 859
rect 7193 810 7207 825
rect 7241 810 7263 844
rect 7193 775 7263 810
rect 7298 844 7344 939
rect 7298 810 7309 844
rect 7343 810 7344 844
rect 6916 665 6928 699
rect 6962 665 6979 699
rect 7107 709 7159 745
rect 7298 767 7344 810
rect 6916 631 6979 665
rect 7014 673 7073 689
rect 7014 639 7023 673
rect 7057 639 7073 673
rect 7014 597 7073 639
rect 7141 675 7159 709
rect 7107 631 7159 675
rect 7211 733 7298 741
rect 7332 733 7344 767
rect 7211 707 7344 733
rect 7413 971 7423 989
rect 7567 973 7601 1023
rect 7379 937 7389 955
rect 7211 699 7245 707
rect 7379 699 7423 937
rect 7457 939 7601 973
rect 7457 745 7491 939
rect 7641 937 7665 971
rect 7699 945 7741 971
rect 7699 937 7707 945
rect 7641 911 7707 937
rect 7525 884 7607 905
rect 7525 850 7542 884
rect 7576 850 7607 884
rect 7525 831 7607 850
rect 7559 797 7607 831
rect 7525 781 7607 797
rect 7641 895 7741 911
rect 7641 771 7685 895
rect 7775 861 7809 1030
rect 7857 1055 7933 1107
rect 8151 1065 8217 1107
rect 7857 1021 7873 1055
rect 7907 1021 7933 1055
rect 7993 1039 8027 1055
rect 7993 987 8027 1005
rect 8151 1031 8167 1065
rect 8201 1031 8217 1065
rect 8640 1065 8716 1107
rect 8151 997 8217 1031
rect 8426 1030 8442 1064
rect 8476 1030 8592 1064
rect 8640 1031 8656 1065
rect 8690 1031 8716 1065
rect 8904 1065 9182 1107
rect 8764 1039 8798 1055
rect 7843 971 8113 987
rect 7843 945 7993 971
rect 7877 937 7993 945
rect 8027 937 8113 971
rect 8151 963 8167 997
rect 8201 963 8217 997
rect 8388 971 8435 977
rect 7877 911 7893 937
rect 7843 895 7893 911
rect 7995 861 8045 877
rect 7775 827 8011 861
rect 7775 819 7859 827
rect 7457 707 7601 745
rect 7675 737 7685 771
rect 7641 721 7685 737
rect 7721 749 7737 783
rect 7771 767 7791 783
rect 7721 733 7757 749
rect 7721 709 7791 733
rect 7211 649 7245 665
rect 7279 639 7295 673
rect 7329 639 7345 673
rect 7413 665 7423 699
rect 7567 691 7601 707
rect 7379 649 7423 665
rect 7279 597 7345 639
rect 7462 639 7483 673
rect 7517 639 7533 673
rect 7825 673 7859 819
rect 8001 811 8045 827
rect 8079 793 8113 937
rect 8388 945 8401 971
rect 8422 911 8435 937
rect 8147 903 8348 911
rect 8147 869 8309 903
rect 8343 869 8348 903
rect 8388 895 8435 911
rect 8483 945 8524 961
rect 8483 911 8490 945
rect 8147 863 8348 869
rect 8147 861 8213 863
rect 8147 827 8163 861
rect 8197 827 8213 861
rect 8483 841 8524 911
rect 8389 835 8524 841
rect 8275 793 8291 827
rect 8325 793 8341 827
rect 7893 759 7909 793
rect 7943 773 7959 793
rect 7943 767 7975 773
rect 7893 733 7941 759
rect 8079 759 8341 793
rect 8389 801 8401 835
rect 8435 805 8524 835
rect 8558 861 8592 1030
rect 8904 1031 8930 1065
rect 8964 1031 9132 1065
rect 9166 1031 9182 1065
rect 8764 997 8798 1005
rect 9216 1028 9273 1073
rect 8626 963 9182 997
rect 8626 945 8676 963
rect 8660 911 8676 945
rect 8626 895 8676 911
rect 8558 845 8828 861
rect 8558 827 8794 845
rect 8435 801 8457 805
rect 8389 792 8457 801
rect 8413 771 8457 792
rect 8079 733 8123 759
rect 7893 727 7975 733
rect 8057 699 8073 733
rect 8107 699 8123 733
rect 8413 737 8423 771
rect 8157 707 8191 723
rect 8413 721 8457 737
rect 7567 641 7601 657
rect 7462 597 7533 639
rect 7656 639 7672 673
rect 7706 639 7859 673
rect 7656 633 7859 639
rect 7893 669 7927 685
rect 7893 597 7927 635
rect 7961 675 8027 681
rect 7961 641 7977 675
rect 8011 665 8027 675
rect 8558 673 8592 827
rect 8784 811 8794 827
rect 8784 795 8828 811
rect 8632 759 8687 793
rect 8721 767 8741 793
rect 8632 733 8691 759
rect 8725 733 8741 767
rect 8862 748 8896 963
rect 8930 903 9034 929
rect 8930 869 8947 903
rect 8981 895 9034 903
rect 9068 895 9087 929
rect 8981 869 8987 895
rect 8930 861 8987 869
rect 8964 827 8987 861
rect 9148 845 9182 963
rect 9250 994 9273 1028
rect 9216 960 9273 994
rect 9250 957 9273 960
rect 9216 923 9227 926
rect 9261 923 9273 957
rect 9216 906 9273 923
rect 8930 802 8987 827
rect 8943 765 8987 802
rect 9023 833 9114 845
rect 9023 799 9039 833
rect 9073 799 9114 833
rect 9148 829 9201 845
rect 9148 795 9167 829
rect 9148 779 9201 795
rect 8862 747 8899 748
rect 8632 727 8741 733
rect 8819 713 8849 747
rect 8883 713 8899 747
rect 8943 731 9071 765
rect 8157 665 8191 673
rect 8011 641 8191 665
rect 7961 631 8191 641
rect 8241 639 8261 673
rect 8295 639 8311 673
rect 8241 597 8311 639
rect 8436 639 8465 673
rect 8499 639 8592 673
rect 8436 633 8592 639
rect 8626 669 8691 685
rect 8626 635 8657 669
rect 8626 597 8691 635
rect 8725 655 8741 689
rect 8775 665 8791 689
rect 8933 681 8967 697
rect 8775 655 8933 665
rect 8725 647 8933 655
rect 8725 631 8967 647
rect 9029 683 9071 731
rect 9029 649 9037 683
rect 9029 633 9071 649
rect 9121 673 9182 741
rect 9237 723 9273 906
rect 9121 639 9132 673
rect 9166 639 9182 673
rect 9121 597 9182 639
rect 9216 707 9273 723
rect 9250 673 9273 707
rect 9216 631 9273 673
rect 9308 1047 9371 1063
rect 9308 1013 9320 1047
rect 9354 1013 9371 1047
rect 9308 979 9371 1013
rect 9308 945 9320 979
rect 9354 945 9371 979
rect 9308 845 9371 945
rect 9407 1053 9465 1107
rect 9407 1019 9415 1053
rect 9449 1019 9465 1053
rect 9407 985 9465 1019
rect 9407 951 9415 985
rect 9449 951 9465 985
rect 9407 933 9465 951
rect 9499 1034 9551 1073
rect 9499 1029 9510 1034
rect 9544 1000 9551 1034
rect 9533 995 9551 1000
rect 9499 961 9551 995
rect 9533 927 9551 961
rect 9603 1057 9637 1073
rect 9603 989 9637 1023
rect 9671 1041 9737 1107
rect 9671 1007 9687 1041
rect 9721 1007 9737 1041
rect 9771 1057 9815 1073
rect 9805 1023 9815 1057
rect 9771 989 9815 1023
rect 9854 1041 9925 1107
rect 9854 1007 9875 1041
rect 9909 1007 9925 1041
rect 9959 1057 9993 1073
rect 10035 1030 10051 1064
rect 10085 1030 10201 1064
rect 9637 955 9736 973
rect 9603 939 9736 955
rect 9499 871 9551 927
rect 9308 829 9475 845
rect 9308 795 9441 829
rect 9308 779 9475 795
rect 9308 699 9371 779
rect 9509 745 9551 871
rect 9585 860 9655 905
rect 9585 826 9593 860
rect 9627 844 9655 860
rect 9585 810 9599 826
rect 9633 810 9655 844
rect 9585 775 9655 810
rect 9690 844 9736 939
rect 9690 810 9701 844
rect 9735 810 9736 844
rect 9308 665 9320 699
rect 9354 665 9371 699
rect 9499 709 9551 745
rect 9690 767 9736 810
rect 9308 631 9371 665
rect 9406 673 9465 689
rect 9406 639 9415 673
rect 9449 639 9465 673
rect 9406 597 9465 639
rect 9533 675 9551 709
rect 9499 631 9551 675
rect 9603 733 9690 741
rect 9724 733 9736 767
rect 9603 707 9736 733
rect 9805 971 9815 989
rect 9959 973 9993 1023
rect 9771 937 9781 955
rect 9603 699 9637 707
rect 9771 699 9815 937
rect 9849 939 9993 973
rect 9849 745 9883 939
rect 10033 937 10057 971
rect 10091 945 10133 971
rect 10091 937 10099 945
rect 10033 911 10099 937
rect 9917 883 9999 905
rect 9917 849 9934 883
rect 9968 849 9999 883
rect 9917 831 9999 849
rect 9951 797 9999 831
rect 9917 781 9999 797
rect 10033 895 10133 911
rect 10033 771 10077 895
rect 10167 861 10201 1030
rect 10249 1055 10325 1107
rect 10543 1065 10609 1107
rect 10249 1021 10265 1055
rect 10299 1021 10325 1055
rect 10385 1039 10419 1055
rect 10385 987 10419 1005
rect 10543 1031 10559 1065
rect 10593 1031 10609 1065
rect 11032 1065 11108 1107
rect 10543 997 10609 1031
rect 10818 1030 10834 1064
rect 10868 1030 10984 1064
rect 11032 1031 11048 1065
rect 11082 1031 11108 1065
rect 11296 1065 11574 1107
rect 11156 1039 11190 1055
rect 10235 971 10505 987
rect 10235 945 10385 971
rect 10269 937 10385 945
rect 10419 937 10505 971
rect 10543 963 10559 997
rect 10593 963 10609 997
rect 10780 971 10827 977
rect 10269 911 10285 937
rect 10235 895 10285 911
rect 10387 861 10437 877
rect 10167 827 10403 861
rect 10167 819 10251 827
rect 9849 707 9993 745
rect 10067 737 10077 771
rect 10033 721 10077 737
rect 10113 749 10129 783
rect 10163 767 10183 783
rect 10113 733 10149 749
rect 10113 709 10183 733
rect 9603 649 9637 665
rect 9671 639 9687 673
rect 9721 639 9737 673
rect 9805 665 9815 699
rect 9959 691 9993 707
rect 9771 649 9815 665
rect 9671 597 9737 639
rect 9854 639 9875 673
rect 9909 639 9925 673
rect 10217 673 10251 819
rect 10393 811 10437 827
rect 10471 793 10505 937
rect 10780 945 10793 971
rect 10814 911 10827 937
rect 10539 903 10740 911
rect 10539 869 10701 903
rect 10735 869 10740 903
rect 10780 895 10827 911
rect 10875 945 10916 961
rect 10875 911 10882 945
rect 10539 863 10740 869
rect 10539 861 10605 863
rect 10539 827 10555 861
rect 10589 827 10605 861
rect 10875 841 10916 911
rect 10781 835 10916 841
rect 10667 793 10683 827
rect 10717 793 10733 827
rect 10285 759 10301 793
rect 10335 773 10351 793
rect 10335 767 10367 773
rect 10285 733 10333 759
rect 10471 759 10733 793
rect 10781 801 10793 835
rect 10827 805 10916 835
rect 10950 861 10984 1030
rect 11296 1031 11322 1065
rect 11356 1031 11524 1065
rect 11558 1031 11574 1065
rect 11156 997 11190 1005
rect 11608 1028 11665 1073
rect 11018 963 11574 997
rect 11018 945 11068 963
rect 11052 911 11068 945
rect 11018 895 11068 911
rect 10950 845 11220 861
rect 10950 827 11186 845
rect 10827 801 10849 805
rect 10781 792 10849 801
rect 10805 771 10849 792
rect 10471 733 10515 759
rect 10285 727 10367 733
rect 10449 699 10465 733
rect 10499 699 10515 733
rect 10805 737 10815 771
rect 10549 707 10583 723
rect 10805 721 10849 737
rect 9959 641 9993 657
rect 9854 597 9925 639
rect 10048 639 10064 673
rect 10098 639 10251 673
rect 10048 633 10251 639
rect 10285 669 10319 685
rect 10285 597 10319 635
rect 10353 675 10419 681
rect 10353 641 10369 675
rect 10403 665 10419 675
rect 10950 673 10984 827
rect 11176 811 11186 827
rect 11176 795 11220 811
rect 11024 759 11079 793
rect 11113 767 11133 793
rect 11024 733 11083 759
rect 11117 733 11133 767
rect 11254 748 11288 963
rect 11322 903 11426 929
rect 11322 869 11339 903
rect 11373 895 11426 903
rect 11460 895 11479 929
rect 11373 869 11379 895
rect 11322 861 11379 869
rect 11356 827 11379 861
rect 11540 845 11574 963
rect 11642 994 11665 1028
rect 11608 960 11665 994
rect 11642 956 11665 960
rect 11608 922 11618 926
rect 11652 922 11665 956
rect 11608 906 11665 922
rect 11322 802 11379 827
rect 11335 765 11379 802
rect 11415 833 11506 845
rect 11415 799 11431 833
rect 11465 799 11506 833
rect 11540 829 11593 845
rect 11540 795 11559 829
rect 11540 779 11593 795
rect 11254 747 11291 748
rect 11024 727 11133 733
rect 11211 713 11241 747
rect 11275 713 11291 747
rect 11335 731 11463 765
rect 10549 665 10583 673
rect 10403 641 10583 665
rect 10353 631 10583 641
rect 10633 639 10653 673
rect 10687 639 10703 673
rect 10633 597 10703 639
rect 10828 639 10857 673
rect 10891 639 10984 673
rect 10828 633 10984 639
rect 11018 669 11083 685
rect 11018 635 11049 669
rect 11018 597 11083 635
rect 11117 655 11133 689
rect 11167 665 11183 689
rect 11325 681 11359 697
rect 11167 655 11325 665
rect 11117 647 11325 655
rect 11117 631 11359 647
rect 11421 683 11463 731
rect 11421 649 11429 683
rect 11421 633 11463 649
rect 11513 673 11574 741
rect 11629 723 11665 906
rect 11513 639 11524 673
rect 11558 639 11574 673
rect 11513 597 11574 639
rect 11608 707 11665 723
rect 11642 673 11665 707
rect 11608 631 11665 673
rect 11700 1047 11763 1063
rect 11700 1013 11712 1047
rect 11746 1013 11763 1047
rect 11700 979 11763 1013
rect 11700 945 11712 979
rect 11746 945 11763 979
rect 11700 845 11763 945
rect 11799 1053 11857 1107
rect 11799 1019 11807 1053
rect 11841 1019 11857 1053
rect 11799 985 11857 1019
rect 11799 951 11807 985
rect 11841 951 11857 985
rect 11799 933 11857 951
rect 11891 1034 11943 1073
rect 11891 1029 11902 1034
rect 11936 1000 11943 1034
rect 11925 995 11943 1000
rect 11891 961 11943 995
rect 11925 927 11943 961
rect 11995 1057 12029 1073
rect 11995 989 12029 1023
rect 12063 1041 12129 1107
rect 12063 1007 12079 1041
rect 12113 1007 12129 1041
rect 12163 1057 12207 1073
rect 12197 1023 12207 1057
rect 12163 989 12207 1023
rect 12246 1041 12317 1107
rect 12246 1007 12267 1041
rect 12301 1007 12317 1041
rect 12351 1057 12385 1073
rect 12427 1030 12443 1064
rect 12477 1030 12593 1064
rect 12029 955 12128 973
rect 11995 939 12128 955
rect 11891 871 11943 927
rect 11700 829 11867 845
rect 11700 795 11833 829
rect 11700 779 11867 795
rect 11700 699 11763 779
rect 11901 745 11943 871
rect 11977 859 12047 905
rect 11977 825 11985 859
rect 12019 844 12047 859
rect 11977 810 11991 825
rect 12025 810 12047 844
rect 11977 775 12047 810
rect 12082 844 12128 939
rect 12082 810 12093 844
rect 12127 810 12128 844
rect 11700 665 11712 699
rect 11746 665 11763 699
rect 11891 709 11943 745
rect 12082 767 12128 810
rect 11700 631 11763 665
rect 11798 673 11857 689
rect 11798 639 11807 673
rect 11841 639 11857 673
rect 11798 597 11857 639
rect 11925 675 11943 709
rect 11891 631 11943 675
rect 11995 733 12082 741
rect 12116 733 12128 767
rect 11995 707 12128 733
rect 12197 971 12207 989
rect 12351 973 12385 1023
rect 12163 937 12173 955
rect 11995 699 12029 707
rect 12163 699 12207 937
rect 12241 939 12385 973
rect 12241 745 12275 939
rect 12425 937 12449 971
rect 12483 945 12525 971
rect 12483 937 12491 945
rect 12425 911 12491 937
rect 12309 884 12391 905
rect 12309 850 12326 884
rect 12360 850 12391 884
rect 12309 831 12391 850
rect 12343 797 12391 831
rect 12309 781 12391 797
rect 12425 895 12525 911
rect 12425 771 12469 895
rect 12559 861 12593 1030
rect 12641 1055 12717 1107
rect 12935 1065 13001 1107
rect 12641 1021 12657 1055
rect 12691 1021 12717 1055
rect 12777 1039 12811 1055
rect 12777 987 12811 1005
rect 12935 1031 12951 1065
rect 12985 1031 13001 1065
rect 13424 1065 13500 1107
rect 12935 997 13001 1031
rect 13210 1030 13226 1064
rect 13260 1030 13376 1064
rect 13424 1031 13440 1065
rect 13474 1031 13500 1065
rect 13688 1065 13966 1107
rect 13548 1039 13582 1055
rect 12627 971 12897 987
rect 12627 945 12777 971
rect 12661 937 12777 945
rect 12811 937 12897 971
rect 12935 963 12951 997
rect 12985 963 13001 997
rect 13172 971 13219 977
rect 12661 911 12677 937
rect 12627 895 12677 911
rect 12779 861 12829 877
rect 12559 827 12795 861
rect 12559 819 12643 827
rect 12241 707 12385 745
rect 12459 737 12469 771
rect 12425 721 12469 737
rect 12505 749 12521 783
rect 12555 767 12575 783
rect 12505 733 12541 749
rect 12505 709 12575 733
rect 11995 649 12029 665
rect 12063 639 12079 673
rect 12113 639 12129 673
rect 12197 665 12207 699
rect 12351 691 12385 707
rect 12163 649 12207 665
rect 12063 597 12129 639
rect 12246 639 12267 673
rect 12301 639 12317 673
rect 12609 673 12643 819
rect 12785 811 12829 827
rect 12863 793 12897 937
rect 13172 945 13185 971
rect 13206 911 13219 937
rect 12931 903 13132 911
rect 12931 869 13093 903
rect 13127 869 13132 903
rect 13172 895 13219 911
rect 13267 945 13308 961
rect 13267 911 13274 945
rect 12931 863 13132 869
rect 12931 861 12997 863
rect 12931 827 12947 861
rect 12981 827 12997 861
rect 13267 841 13308 911
rect 13173 835 13308 841
rect 13059 793 13075 827
rect 13109 793 13125 827
rect 12677 759 12693 793
rect 12727 773 12743 793
rect 12727 767 12759 773
rect 12677 733 12725 759
rect 12863 759 13125 793
rect 13173 801 13185 835
rect 13219 805 13308 835
rect 13342 861 13376 1030
rect 13688 1031 13714 1065
rect 13748 1031 13916 1065
rect 13950 1031 13966 1065
rect 13548 997 13582 1005
rect 14000 1028 14057 1073
rect 13410 963 13966 997
rect 13410 945 13460 963
rect 13444 911 13460 945
rect 13410 895 13460 911
rect 13342 845 13612 861
rect 13342 827 13578 845
rect 13219 801 13241 805
rect 13173 792 13241 801
rect 13197 771 13241 792
rect 12863 733 12907 759
rect 12677 727 12759 733
rect 12841 699 12857 733
rect 12891 699 12907 733
rect 13197 737 13207 771
rect 12941 707 12975 723
rect 13197 721 13241 737
rect 12351 641 12385 657
rect 12246 597 12317 639
rect 12440 639 12456 673
rect 12490 639 12643 673
rect 12440 633 12643 639
rect 12677 669 12711 685
rect 12677 597 12711 635
rect 12745 675 12811 681
rect 12745 641 12761 675
rect 12795 665 12811 675
rect 13342 673 13376 827
rect 13568 811 13578 827
rect 13568 795 13612 811
rect 13416 759 13471 793
rect 13505 767 13525 793
rect 13416 733 13475 759
rect 13509 733 13525 767
rect 13646 748 13680 963
rect 13714 903 13818 929
rect 13714 869 13731 903
rect 13765 895 13818 903
rect 13852 895 13871 929
rect 13765 869 13771 895
rect 13714 861 13771 869
rect 13748 827 13771 861
rect 13932 845 13966 963
rect 14034 994 14057 1028
rect 14000 960 14057 994
rect 14034 955 14057 960
rect 14000 921 14011 926
rect 14045 921 14057 955
rect 14000 906 14057 921
rect 13714 802 13771 827
rect 13727 765 13771 802
rect 13807 833 13898 845
rect 13807 799 13823 833
rect 13857 799 13898 833
rect 13932 829 13985 845
rect 13932 795 13951 829
rect 13932 779 13985 795
rect 13646 747 13683 748
rect 13416 727 13525 733
rect 13603 713 13633 747
rect 13667 713 13683 747
rect 13727 731 13855 765
rect 12941 665 12975 673
rect 12795 641 12975 665
rect 12745 631 12975 641
rect 13025 639 13045 673
rect 13079 639 13095 673
rect 13025 597 13095 639
rect 13220 639 13249 673
rect 13283 639 13376 673
rect 13220 633 13376 639
rect 13410 669 13475 685
rect 13410 635 13441 669
rect 13410 597 13475 635
rect 13509 655 13525 689
rect 13559 665 13575 689
rect 13717 681 13751 697
rect 13559 655 13717 665
rect 13509 647 13717 655
rect 13509 631 13751 647
rect 13813 683 13855 731
rect 13813 649 13821 683
rect 13813 633 13855 649
rect 13905 673 13966 741
rect 14021 723 14057 906
rect 13905 639 13916 673
rect 13950 639 13966 673
rect 13905 597 13966 639
rect 14000 707 14057 723
rect 14034 673 14057 707
rect 14000 631 14057 673
rect 14092 1047 14155 1063
rect 14092 1013 14104 1047
rect 14138 1013 14155 1047
rect 14092 979 14155 1013
rect 14092 945 14104 979
rect 14138 945 14155 979
rect 14092 845 14155 945
rect 14191 1053 14249 1107
rect 14191 1019 14199 1053
rect 14233 1019 14249 1053
rect 14191 985 14249 1019
rect 14191 951 14199 985
rect 14233 951 14249 985
rect 14191 933 14249 951
rect 14283 1034 14335 1073
rect 14283 1029 14294 1034
rect 14328 1000 14335 1034
rect 14317 995 14335 1000
rect 14283 961 14335 995
rect 14317 927 14335 961
rect 14387 1057 14421 1073
rect 14387 989 14421 1023
rect 14455 1041 14521 1107
rect 14455 1007 14471 1041
rect 14505 1007 14521 1041
rect 14555 1057 14599 1073
rect 14589 1023 14599 1057
rect 14555 989 14599 1023
rect 14638 1041 14709 1107
rect 14638 1007 14659 1041
rect 14693 1007 14709 1041
rect 14743 1057 14777 1073
rect 14819 1030 14835 1064
rect 14869 1030 14985 1064
rect 14421 955 14520 973
rect 14387 939 14520 955
rect 14283 871 14335 927
rect 14092 829 14259 845
rect 14092 795 14225 829
rect 14092 779 14259 795
rect 14092 699 14155 779
rect 14293 745 14335 871
rect 14369 860 14439 905
rect 14369 826 14378 860
rect 14412 844 14439 860
rect 14369 810 14383 826
rect 14417 810 14439 844
rect 14369 775 14439 810
rect 14474 844 14520 939
rect 14474 810 14485 844
rect 14519 810 14520 844
rect 14092 665 14104 699
rect 14138 665 14155 699
rect 14283 709 14335 745
rect 14474 767 14520 810
rect 14092 631 14155 665
rect 14190 673 14249 689
rect 14190 639 14199 673
rect 14233 639 14249 673
rect 14190 597 14249 639
rect 14317 675 14335 709
rect 14283 631 14335 675
rect 14387 733 14474 741
rect 14508 733 14520 767
rect 14387 707 14520 733
rect 14589 971 14599 989
rect 14743 973 14777 1023
rect 14555 937 14565 955
rect 14387 699 14421 707
rect 14555 699 14599 937
rect 14633 939 14777 973
rect 14633 745 14667 939
rect 14817 937 14841 971
rect 14875 945 14917 971
rect 14875 937 14883 945
rect 14817 911 14883 937
rect 14701 883 14783 905
rect 14701 849 14719 883
rect 14753 849 14783 883
rect 14701 831 14783 849
rect 14735 797 14783 831
rect 14701 781 14783 797
rect 14817 895 14917 911
rect 14817 771 14861 895
rect 14951 861 14985 1030
rect 15033 1055 15109 1107
rect 15327 1065 15393 1107
rect 15033 1021 15049 1055
rect 15083 1021 15109 1055
rect 15169 1039 15203 1055
rect 15169 987 15203 1005
rect 15327 1031 15343 1065
rect 15377 1031 15393 1065
rect 15816 1065 15892 1107
rect 15327 997 15393 1031
rect 15602 1030 15618 1064
rect 15652 1030 15768 1064
rect 15816 1031 15832 1065
rect 15866 1031 15892 1065
rect 16080 1065 16358 1107
rect 15940 1039 15974 1055
rect 15019 971 15289 987
rect 15019 945 15169 971
rect 15053 937 15169 945
rect 15203 937 15289 971
rect 15327 963 15343 997
rect 15377 963 15393 997
rect 15564 971 15611 977
rect 15053 911 15069 937
rect 15019 895 15069 911
rect 15171 861 15221 877
rect 14951 827 15187 861
rect 14951 819 15035 827
rect 14633 707 14777 745
rect 14851 737 14861 771
rect 14817 721 14861 737
rect 14897 749 14913 783
rect 14947 767 14967 783
rect 14897 733 14933 749
rect 14897 709 14967 733
rect 14387 649 14421 665
rect 14455 639 14471 673
rect 14505 639 14521 673
rect 14589 665 14599 699
rect 14743 691 14777 707
rect 14555 649 14599 665
rect 14455 597 14521 639
rect 14638 639 14659 673
rect 14693 639 14709 673
rect 15001 673 15035 819
rect 15177 811 15221 827
rect 15255 793 15289 937
rect 15564 945 15577 971
rect 15598 911 15611 937
rect 15323 903 15524 911
rect 15323 869 15485 903
rect 15519 869 15524 903
rect 15564 895 15611 911
rect 15659 945 15700 961
rect 15659 911 15666 945
rect 15323 863 15524 869
rect 15323 861 15389 863
rect 15323 827 15339 861
rect 15373 827 15389 861
rect 15659 841 15700 911
rect 15565 835 15700 841
rect 15451 793 15467 827
rect 15501 793 15517 827
rect 15069 759 15085 793
rect 15119 773 15135 793
rect 15119 767 15151 773
rect 15069 733 15117 759
rect 15255 759 15517 793
rect 15565 801 15577 835
rect 15611 805 15700 835
rect 15734 861 15768 1030
rect 16080 1031 16106 1065
rect 16140 1031 16308 1065
rect 16342 1031 16358 1065
rect 15940 997 15974 1005
rect 16392 1028 16449 1073
rect 15802 963 16358 997
rect 15802 945 15852 963
rect 15836 911 15852 945
rect 15802 895 15852 911
rect 15734 845 16004 861
rect 15734 827 15970 845
rect 15611 801 15633 805
rect 15565 792 15633 801
rect 15589 771 15633 792
rect 15255 733 15299 759
rect 15069 727 15151 733
rect 15233 699 15249 733
rect 15283 699 15299 733
rect 15589 737 15599 771
rect 15333 707 15367 723
rect 15589 721 15633 737
rect 14743 641 14777 657
rect 14638 597 14709 639
rect 14832 639 14848 673
rect 14882 639 15035 673
rect 14832 633 15035 639
rect 15069 669 15103 685
rect 15069 597 15103 635
rect 15137 675 15203 681
rect 15137 641 15153 675
rect 15187 665 15203 675
rect 15734 673 15768 827
rect 15960 811 15970 827
rect 15960 795 16004 811
rect 15808 759 15863 793
rect 15897 767 15917 793
rect 15808 733 15867 759
rect 15901 733 15917 767
rect 16038 748 16072 963
rect 16106 903 16210 929
rect 16106 869 16123 903
rect 16157 895 16210 903
rect 16244 895 16263 929
rect 16157 869 16163 895
rect 16106 861 16163 869
rect 16140 827 16163 861
rect 16324 845 16358 963
rect 16426 994 16449 1028
rect 16392 960 16449 994
rect 16426 957 16449 960
rect 16392 923 16404 926
rect 16438 923 16449 957
rect 16392 906 16449 923
rect 16106 802 16163 827
rect 16119 765 16163 802
rect 16199 833 16290 845
rect 16199 799 16215 833
rect 16249 799 16290 833
rect 16324 829 16377 845
rect 16324 795 16343 829
rect 16324 779 16377 795
rect 16038 747 16075 748
rect 15808 727 15917 733
rect 15995 713 16025 747
rect 16059 713 16075 747
rect 16119 731 16247 765
rect 15333 665 15367 673
rect 15187 641 15367 665
rect 15137 631 15367 641
rect 15417 639 15437 673
rect 15471 639 15487 673
rect 15417 597 15487 639
rect 15612 639 15641 673
rect 15675 639 15768 673
rect 15612 633 15768 639
rect 15802 669 15867 685
rect 15802 635 15833 669
rect 15802 597 15867 635
rect 15901 655 15917 689
rect 15951 665 15967 689
rect 16109 681 16143 697
rect 15951 655 16109 665
rect 15901 647 16109 655
rect 15901 631 16143 647
rect 16205 683 16247 731
rect 16205 649 16213 683
rect 16205 633 16247 649
rect 16297 673 16358 741
rect 16413 723 16449 906
rect 16297 639 16308 673
rect 16342 639 16358 673
rect 16297 597 16358 639
rect 16392 707 16449 723
rect 16426 673 16449 707
rect 16392 631 16449 673
rect 16484 1047 16547 1063
rect 16484 1013 16496 1047
rect 16530 1013 16547 1047
rect 16484 979 16547 1013
rect 16484 945 16496 979
rect 16530 945 16547 979
rect 16484 845 16547 945
rect 16583 1053 16641 1107
rect 16583 1019 16591 1053
rect 16625 1019 16641 1053
rect 16583 985 16641 1019
rect 16583 951 16591 985
rect 16625 951 16641 985
rect 16583 933 16641 951
rect 16675 1034 16727 1073
rect 16675 1029 16686 1034
rect 16720 1000 16727 1034
rect 16709 995 16727 1000
rect 16675 961 16727 995
rect 16709 927 16727 961
rect 16675 871 16727 927
rect 16484 829 16651 845
rect 16484 795 16617 829
rect 16484 779 16651 795
rect 16484 699 16547 779
rect 16685 745 16727 871
rect 16484 665 16496 699
rect 16530 665 16547 699
rect 16675 709 16727 745
rect 16484 631 16547 665
rect 16582 673 16641 689
rect 16582 639 16591 673
rect 16625 639 16641 673
rect 16582 597 16641 639
rect 16709 675 16727 709
rect 16675 631 16727 675
rect 0 539 29 597
rect 63 539 121 597
rect 155 539 213 597
rect 247 539 305 597
rect 339 539 397 597
rect 431 539 489 597
rect 523 539 581 597
rect 615 539 673 597
rect 707 539 765 597
rect 799 539 857 597
rect 891 539 949 597
rect 983 539 1041 597
rect 1075 539 1133 597
rect 1167 539 1225 597
rect 1259 539 1317 597
rect 1351 539 1409 597
rect 1443 539 1501 597
rect 1535 539 1593 597
rect 1627 539 1685 597
rect 1719 539 1777 597
rect 1811 539 1869 597
rect 1903 539 1961 597
rect 1995 539 2053 597
rect 2087 539 2145 597
rect 2179 539 2237 597
rect 2271 539 2329 597
rect 2363 539 2421 597
rect 2455 539 2513 597
rect 2547 539 2605 597
rect 2639 539 2697 597
rect 2731 539 2789 597
rect 2823 539 2881 597
rect 2915 539 2973 597
rect 3007 539 3065 597
rect 3099 539 3157 597
rect 3191 539 3249 597
rect 3283 539 3341 597
rect 3375 539 3433 597
rect 3467 539 3525 597
rect 3559 539 3617 597
rect 3651 539 3709 597
rect 3743 539 3801 597
rect 3835 539 3893 597
rect 3927 539 3985 597
rect 4019 539 4077 597
rect 4111 539 4169 597
rect 4203 539 4261 597
rect 4295 539 4353 597
rect 4387 539 4445 597
rect 4479 539 4537 597
rect 4571 539 4629 597
rect 4663 539 4721 597
rect 4755 539 4813 597
rect 4847 539 4905 597
rect 4939 539 4997 597
rect 5031 539 5089 597
rect 5123 539 5181 597
rect 5215 539 5273 597
rect 5307 539 5365 597
rect 5399 539 5457 597
rect 5491 539 5549 597
rect 5583 539 5641 597
rect 5675 539 5733 597
rect 5767 539 5825 597
rect 5859 539 5917 597
rect 5951 539 6009 597
rect 6043 539 6101 597
rect 6135 539 6193 597
rect 6227 539 6285 597
rect 6319 539 6377 597
rect 6411 539 6469 597
rect 6503 539 6561 597
rect 6595 539 6653 597
rect 6687 539 6745 597
rect 6779 539 6837 597
rect 6871 539 6929 597
rect 6963 539 7021 597
rect 7055 539 7113 597
rect 7147 539 7205 597
rect 7239 539 7297 597
rect 7331 539 7389 597
rect 7423 539 7481 597
rect 7515 539 7573 597
rect 7607 539 7665 597
rect 7699 539 7757 597
rect 7791 539 7849 597
rect 7883 539 7941 597
rect 7975 539 8033 597
rect 8067 539 8125 597
rect 8159 539 8217 597
rect 8251 539 8309 597
rect 8343 539 8401 597
rect 8435 539 8493 597
rect 8527 539 8585 597
rect 8619 539 8677 597
rect 8711 539 8769 597
rect 8803 539 8861 597
rect 8895 539 8953 597
rect 8987 539 9045 597
rect 9079 539 9137 597
rect 9171 539 9229 597
rect 9263 539 9321 597
rect 9355 539 9413 597
rect 9447 539 9505 597
rect 9539 539 9597 597
rect 9631 539 9689 597
rect 9723 539 9781 597
rect 9815 539 9873 597
rect 9907 539 9965 597
rect 9999 539 10057 597
rect 10091 539 10149 597
rect 10183 539 10241 597
rect 10275 539 10333 597
rect 10367 539 10425 597
rect 10459 539 10517 597
rect 10551 539 10609 597
rect 10643 539 10701 597
rect 10735 539 10793 597
rect 10827 539 10885 597
rect 10919 539 10977 597
rect 11011 539 11069 597
rect 11103 539 11161 597
rect 11195 539 11253 597
rect 11287 539 11345 597
rect 11379 539 11437 597
rect 11471 539 11529 597
rect 11563 539 11621 597
rect 11655 539 11713 597
rect 11747 539 11805 597
rect 11839 539 11897 597
rect 11931 539 11989 597
rect 12023 539 12081 597
rect 12115 539 12173 597
rect 12207 539 12265 597
rect 12299 539 12357 597
rect 12391 539 12449 597
rect 12483 539 12541 597
rect 12575 539 12633 597
rect 12667 539 12725 597
rect 12759 539 12817 597
rect 12851 539 12909 597
rect 12943 539 13001 597
rect 13035 539 13093 597
rect 13127 539 13185 597
rect 13219 539 13277 597
rect 13311 539 13369 597
rect 13403 539 13461 597
rect 13495 539 13553 597
rect 13587 539 13645 597
rect 13679 539 13737 597
rect 13771 539 13829 597
rect 13863 539 13921 597
rect 13955 539 14013 597
rect 14047 539 14105 597
rect 14139 539 14197 597
rect 14231 539 14289 597
rect 14323 539 14381 597
rect 14415 539 14473 597
rect 14507 539 14565 597
rect 14599 539 14657 597
rect 14691 539 14749 597
rect 14783 539 14841 597
rect 14875 539 14933 597
rect 14967 539 15025 597
rect 15059 539 15117 597
rect 15151 539 15209 597
rect 15243 539 15301 597
rect 15335 539 15393 597
rect 15427 539 15485 597
rect 15519 539 15577 597
rect 15611 539 15669 597
rect 15703 539 15761 597
rect 15795 539 15853 597
rect 15887 539 15945 597
rect 15979 539 16037 597
rect 16071 539 16129 597
rect 16163 539 16221 597
rect 16255 539 16313 597
rect 16347 539 16405 597
rect 16439 539 16497 597
rect 16531 539 16589 597
rect 16623 539 16681 597
rect 16715 539 16744 597
rect 0 476 571 477
rect 0 418 29 476
rect 63 418 121 476
rect 155 418 213 476
rect 247 418 305 476
rect 339 442 394 476
rect 428 452 496 476
rect 339 418 397 442
rect 431 418 489 452
rect 530 442 581 476
rect 523 418 581 442
rect 615 418 673 476
rect 707 418 765 476
rect 799 418 857 476
rect 891 418 949 476
rect 983 418 1041 476
rect 1075 418 1133 476
rect 1167 418 1225 476
rect 1259 418 1317 476
rect 1351 418 1409 476
rect 1443 418 1501 476
rect 1535 472 1777 476
rect 1535 452 1607 472
rect 1641 452 1777 472
rect 1535 418 1593 452
rect 1641 438 1685 452
rect 1627 418 1685 438
rect 1719 418 1777 452
rect 1811 418 1869 476
rect 1903 418 1961 476
rect 1995 418 2053 476
rect 2087 418 2145 476
rect 2179 418 2237 476
rect 2271 418 2329 476
rect 2363 418 2421 476
rect 2455 418 2513 476
rect 2547 418 2605 476
rect 2639 418 2697 476
rect 2731 452 2791 476
rect 2825 452 2882 476
rect 2731 418 2789 452
rect 2825 442 2881 452
rect 2916 442 2973 476
rect 2823 418 2881 442
rect 2915 418 2973 442
rect 3007 418 3065 476
rect 3099 418 3157 476
rect 3191 418 3249 476
rect 3283 418 3341 476
rect 3375 418 3433 476
rect 3467 418 3525 476
rect 3559 418 3617 476
rect 3651 418 3709 476
rect 3743 418 3801 476
rect 3835 418 3893 476
rect 3927 472 4169 476
rect 3927 452 3999 472
rect 4033 452 4169 472
rect 3927 418 3985 452
rect 4033 438 4077 452
rect 4019 418 4077 438
rect 4111 418 4169 452
rect 4203 418 4261 476
rect 4295 418 4353 476
rect 4387 418 4445 476
rect 4479 418 4537 476
rect 4571 418 4629 476
rect 4663 418 4721 476
rect 4755 418 4813 476
rect 4847 418 4905 476
rect 4939 418 4997 476
rect 5031 418 5089 476
rect 5123 442 5179 476
rect 5213 452 5273 476
rect 5123 418 5181 442
rect 5215 418 5273 452
rect 5307 418 5365 476
rect 5399 418 5457 476
rect 5491 418 5549 476
rect 5583 418 5641 476
rect 5675 418 5733 476
rect 5767 418 5825 476
rect 5859 418 5917 476
rect 5951 418 6009 476
rect 6043 418 6101 476
rect 6135 418 6193 476
rect 6227 418 6285 476
rect 6319 472 6561 476
rect 6319 452 6391 472
rect 6425 452 6561 472
rect 6319 418 6377 452
rect 6425 438 6469 452
rect 6411 418 6469 438
rect 6503 418 6561 452
rect 6595 418 6653 476
rect 6687 418 6745 476
rect 6779 418 6837 476
rect 6871 418 6929 476
rect 6963 418 7021 476
rect 7055 418 7113 476
rect 7147 418 7205 476
rect 7239 418 7297 476
rect 7331 418 7389 476
rect 7423 418 7481 476
rect 7515 452 7574 476
rect 7515 418 7573 452
rect 7608 442 7665 476
rect 7607 418 7665 442
rect 7699 418 7757 476
rect 7791 418 7849 476
rect 7883 418 7941 476
rect 7975 418 8033 476
rect 8067 418 8125 476
rect 8159 418 8217 476
rect 8251 418 8309 476
rect 8343 418 8401 476
rect 8435 418 8493 476
rect 8527 418 8585 476
rect 8619 418 8677 476
rect 8711 472 8953 476
rect 8711 452 8783 472
rect 8817 452 8953 472
rect 8711 418 8769 452
rect 8817 438 8861 452
rect 8803 418 8861 438
rect 8895 418 8953 452
rect 8987 418 9045 476
rect 9079 418 9137 476
rect 9171 418 9229 476
rect 9263 418 9321 476
rect 9355 418 9413 476
rect 9447 418 9505 476
rect 9539 418 9597 476
rect 9631 418 9689 476
rect 9723 418 9781 476
rect 9815 418 9873 476
rect 9907 442 9963 476
rect 9997 452 10058 476
rect 9907 418 9965 442
rect 9999 418 10057 452
rect 10092 442 10149 476
rect 10091 418 10149 442
rect 10183 418 10241 476
rect 10275 418 10333 476
rect 10367 418 10425 476
rect 10459 418 10517 476
rect 10551 418 10609 476
rect 10643 418 10701 476
rect 10735 418 10793 476
rect 10827 418 10885 476
rect 10919 418 10977 476
rect 11011 418 11069 476
rect 11103 472 11345 476
rect 11103 452 11175 472
rect 11209 452 11345 472
rect 11103 418 11161 452
rect 11209 438 11253 452
rect 11195 418 11253 438
rect 11287 418 11345 452
rect 11379 418 11437 476
rect 11471 418 11529 476
rect 11563 418 11621 476
rect 11655 418 11713 476
rect 11747 418 11805 476
rect 11839 418 11897 476
rect 11931 418 11989 476
rect 12023 418 12081 476
rect 12115 418 12173 476
rect 12207 418 12265 476
rect 12299 418 12357 476
rect 12391 442 12448 476
rect 12482 452 12541 476
rect 12391 418 12449 442
rect 12483 418 12541 452
rect 12575 418 12633 476
rect 12667 418 12725 476
rect 12759 418 12817 476
rect 12851 418 12909 476
rect 12943 418 13001 476
rect 13035 418 13093 476
rect 13127 418 13185 476
rect 13219 418 13277 476
rect 13311 418 13369 476
rect 13403 418 13461 476
rect 13495 472 13737 476
rect 13495 452 13567 472
rect 13601 452 13737 472
rect 13495 418 13553 452
rect 13601 438 13645 452
rect 13587 418 13645 438
rect 13679 418 13737 452
rect 13771 418 13829 476
rect 13863 418 13921 476
rect 13955 418 14013 476
rect 14047 418 14105 476
rect 14139 418 14197 476
rect 14231 418 14289 476
rect 14323 418 14381 476
rect 14415 418 14473 476
rect 14507 418 14565 476
rect 14599 418 14657 476
rect 14691 442 14748 476
rect 14782 452 14842 476
rect 14691 418 14749 442
rect 14783 418 14841 452
rect 14876 442 14933 476
rect 14875 418 14933 442
rect 14967 418 15025 476
rect 15059 418 15117 476
rect 15151 418 15209 476
rect 15243 418 15301 476
rect 15335 418 15393 476
rect 15427 418 15485 476
rect 15519 418 15577 476
rect 15611 418 15669 476
rect 15703 418 15761 476
rect 15795 418 15853 476
rect 15887 469 16129 476
rect 15887 452 15959 469
rect 15993 452 16129 469
rect 15887 418 15945 452
rect 15993 435 16037 452
rect 15979 418 16037 435
rect 16071 418 16129 452
rect 16163 418 16221 476
rect 16255 418 16313 476
rect 16347 418 16405 476
rect 16439 418 16497 476
rect 16531 418 16589 476
rect 16623 418 16681 476
rect 16715 418 16744 476
rect 17 342 69 384
rect 17 308 26 342
rect 60 340 69 342
rect 17 306 35 308
rect 17 272 69 306
rect 17 238 35 272
rect 103 364 161 418
rect 103 330 119 364
rect 153 330 161 364
rect 103 296 161 330
rect 103 262 119 296
rect 153 262 161 296
rect 103 244 161 262
rect 197 358 260 374
rect 197 324 214 358
rect 248 324 260 358
rect 197 290 260 324
rect 197 256 214 290
rect 248 256 260 290
rect 17 182 69 238
rect 17 56 59 182
rect 197 156 260 256
rect 93 140 260 156
rect 127 106 260 140
rect 93 90 260 106
rect 17 20 69 56
rect 17 -14 35 20
rect 197 10 260 90
rect 17 -58 69 -14
rect 103 -16 162 0
rect 103 -50 119 -16
rect 153 -50 162 -16
rect 103 -92 162 -50
rect 197 -24 214 10
rect 248 -24 260 10
rect 197 -58 260 -24
rect 295 339 352 384
rect 386 376 664 418
rect 386 342 402 376
rect 436 342 604 376
rect 638 342 664 376
rect 852 376 928 418
rect 770 350 804 366
rect 295 305 318 339
rect 852 342 878 376
rect 912 342 928 376
rect 1351 376 1417 418
rect 770 308 804 316
rect 976 341 1092 375
rect 1126 341 1142 375
rect 1351 342 1367 376
rect 1401 342 1417 376
rect 1635 366 1711 418
rect 295 276 352 305
rect 295 242 306 276
rect 340 271 352 276
rect 295 237 318 242
rect 295 217 352 237
rect 386 274 942 308
rect 295 34 331 217
rect 386 156 420 274
rect 481 206 500 240
rect 534 214 638 240
rect 534 206 587 214
rect 581 180 587 206
rect 621 180 638 214
rect 581 172 638 180
rect 367 140 420 156
rect 401 106 420 140
rect 454 148 545 156
rect 454 144 502 148
rect 454 110 495 144
rect 536 114 545 148
rect 529 110 545 114
rect 581 138 604 172
rect 581 113 638 138
rect 367 90 420 106
rect 581 76 625 113
rect 295 18 352 34
rect 295 -16 318 18
rect 295 -58 352 -16
rect 386 -16 447 52
rect 386 -50 402 -16
rect 436 -50 447 -16
rect 386 -92 447 -50
rect 497 42 625 76
rect 672 59 706 274
rect 892 256 942 274
rect 892 222 908 256
rect 892 206 942 222
rect 976 172 1010 341
rect 1351 308 1417 342
rect 1133 282 1180 288
rect 740 156 1010 172
rect 774 138 1010 156
rect 774 122 784 138
rect 740 106 784 122
rect 669 58 706 59
rect 827 78 847 104
rect 497 -6 539 42
rect 669 24 685 58
rect 719 24 749 58
rect 827 44 843 78
rect 881 70 936 104
rect 877 44 936 70
rect 827 38 936 44
rect 531 -40 539 -6
rect 497 -56 539 -40
rect 601 -8 635 8
rect 777 -24 793 0
rect 635 -34 793 -24
rect 827 -34 843 0
rect 635 -42 843 -34
rect 601 -58 843 -42
rect 877 -20 942 -4
rect 911 -54 942 -20
rect 877 -92 942 -54
rect 976 -16 1010 138
rect 1044 256 1085 272
rect 1078 222 1085 256
rect 1044 152 1085 222
rect 1167 256 1180 282
rect 1351 274 1367 308
rect 1401 274 1417 308
rect 1541 350 1575 366
rect 1635 332 1661 366
rect 1695 332 1711 366
rect 1759 341 1875 375
rect 1909 341 1925 375
rect 1967 368 2001 384
rect 1541 298 1575 316
rect 1455 282 1725 298
rect 1133 222 1146 248
rect 1455 248 1541 282
rect 1575 256 1725 282
rect 1575 248 1691 256
rect 1133 206 1180 222
rect 1220 214 1421 222
rect 1220 180 1225 214
rect 1259 180 1421 214
rect 1220 174 1421 180
rect 1355 172 1421 174
rect 1044 146 1179 152
rect 1044 116 1133 146
rect 1111 112 1133 116
rect 1167 112 1179 146
rect 1355 138 1371 172
rect 1405 138 1421 172
rect 1111 103 1179 112
rect 1227 104 1243 138
rect 1277 104 1293 138
rect 1455 104 1489 248
rect 1675 222 1691 248
rect 1675 206 1725 222
rect 1523 172 1573 188
rect 1759 172 1793 341
rect 1967 284 2001 334
rect 2035 352 2106 418
rect 2035 318 2051 352
rect 2085 318 2106 352
rect 2145 368 2189 384
rect 2145 334 2155 368
rect 2145 300 2189 334
rect 2223 352 2289 418
rect 2223 318 2239 352
rect 2273 318 2289 352
rect 2323 368 2357 384
rect 1827 256 1869 282
rect 1861 248 1869 256
rect 1903 248 1927 282
rect 1967 250 2111 284
rect 1861 222 1927 248
rect 1827 206 1927 222
rect 1557 138 1793 172
rect 1523 122 1567 138
rect 1709 130 1793 138
rect 1111 82 1155 103
rect 1145 48 1155 82
rect 1227 70 1489 104
rect 1609 84 1625 104
rect 1111 32 1155 48
rect 1445 44 1489 70
rect 1593 78 1625 84
rect 1659 70 1675 104
rect 1627 44 1675 70
rect 1377 18 1411 34
rect 1445 10 1461 44
rect 1495 10 1511 44
rect 1593 38 1675 44
rect 976 -50 1069 -16
rect 1103 -50 1132 -16
rect 976 -56 1132 -50
rect 1257 -50 1273 -16
rect 1307 -50 1327 -16
rect 1257 -92 1327 -50
rect 1377 -24 1411 -16
rect 1541 -14 1607 -8
rect 1541 -24 1557 -14
rect 1377 -48 1557 -24
rect 1591 -48 1607 -14
rect 1377 -58 1607 -48
rect 1641 -20 1675 -4
rect 1641 -92 1675 -54
rect 1709 -16 1743 130
rect 1777 78 1797 94
rect 1831 60 1847 94
rect 1811 44 1847 60
rect 1777 20 1847 44
rect 1883 82 1927 206
rect 1961 149 2043 216
rect 1961 115 1968 149
rect 2002 142 2043 149
rect 2002 115 2009 142
rect 1961 108 2009 115
rect 1961 92 2043 108
rect 1883 48 1893 82
rect 2077 56 2111 250
rect 1883 32 1927 48
rect 1967 18 2111 56
rect 2145 282 2155 300
rect 2323 300 2357 334
rect 2179 248 2189 266
rect 1967 2 2001 18
rect 1709 -50 1862 -16
rect 1896 -50 1912 -16
rect 2145 10 2189 248
rect 2224 266 2323 284
rect 2224 250 2357 266
rect 2409 342 2461 384
rect 2409 308 2418 342
rect 2452 340 2461 342
rect 2409 306 2427 308
rect 2409 272 2461 306
rect 2224 155 2270 250
rect 2409 238 2427 272
rect 2495 364 2553 418
rect 2495 330 2511 364
rect 2545 330 2553 364
rect 2495 296 2553 330
rect 2495 262 2511 296
rect 2545 262 2553 296
rect 2495 244 2553 262
rect 2589 358 2652 374
rect 2589 324 2606 358
rect 2640 324 2652 358
rect 2589 290 2652 324
rect 2589 256 2606 290
rect 2640 256 2652 290
rect 2224 121 2225 155
rect 2259 121 2270 155
rect 2224 78 2270 121
rect 2305 205 2375 216
rect 2305 171 2314 205
rect 2348 171 2375 205
rect 2305 155 2375 171
rect 2305 121 2327 155
rect 2361 121 2375 155
rect 2305 86 2375 121
rect 2409 182 2461 238
rect 2224 44 2236 78
rect 2409 56 2451 182
rect 2589 156 2652 256
rect 2485 140 2652 156
rect 2519 106 2652 140
rect 2485 90 2652 106
rect 2270 44 2357 52
rect 2224 18 2357 44
rect 1967 -48 2001 -32
rect 1709 -56 1912 -50
rect 2035 -50 2051 -16
rect 2085 -50 2106 -16
rect 2145 -24 2155 10
rect 2323 10 2357 18
rect 2145 -40 2189 -24
rect 2035 -92 2106 -50
rect 2223 -50 2239 -16
rect 2273 -50 2289 -16
rect 2323 -40 2357 -24
rect 2409 20 2461 56
rect 2409 -14 2427 20
rect 2589 10 2652 90
rect 2223 -92 2289 -50
rect 2409 -58 2461 -14
rect 2495 -16 2554 0
rect 2495 -50 2511 -16
rect 2545 -50 2554 -16
rect 2495 -92 2554 -50
rect 2589 -24 2606 10
rect 2640 -24 2652 10
rect 2589 -58 2652 -24
rect 2687 339 2744 384
rect 2778 376 3056 418
rect 2778 342 2794 376
rect 2828 342 2996 376
rect 3030 342 3056 376
rect 3244 376 3320 418
rect 3162 350 3196 366
rect 2687 305 2710 339
rect 3244 342 3270 376
rect 3304 342 3320 376
rect 3743 376 3809 418
rect 3162 308 3196 316
rect 3368 341 3484 375
rect 3518 341 3534 375
rect 3743 342 3759 376
rect 3793 342 3809 376
rect 4027 366 4103 418
rect 2687 276 2744 305
rect 2687 242 2698 276
rect 2732 271 2744 276
rect 2687 237 2710 242
rect 2687 217 2744 237
rect 2778 274 3334 308
rect 2687 34 2723 217
rect 2778 156 2812 274
rect 2873 206 2892 240
rect 2926 214 3030 240
rect 2926 206 2979 214
rect 2973 180 2979 206
rect 3013 180 3030 214
rect 2973 172 3030 180
rect 2759 140 2812 156
rect 2793 106 2812 140
rect 2846 150 2937 156
rect 2846 144 2891 150
rect 2846 110 2887 144
rect 2925 116 2937 150
rect 2921 110 2937 116
rect 2973 138 2996 172
rect 2973 113 3030 138
rect 2759 90 2812 106
rect 2973 76 3017 113
rect 2687 18 2744 34
rect 2687 -16 2710 18
rect 2687 -58 2744 -16
rect 2778 -16 2839 52
rect 2778 -50 2794 -16
rect 2828 -50 2839 -16
rect 2778 -92 2839 -50
rect 2889 42 3017 76
rect 3064 59 3098 274
rect 3284 256 3334 274
rect 3284 222 3300 256
rect 3284 206 3334 222
rect 3368 172 3402 341
rect 3743 308 3809 342
rect 3525 282 3572 288
rect 3132 156 3402 172
rect 3166 138 3402 156
rect 3166 122 3176 138
rect 3132 106 3176 122
rect 3061 58 3098 59
rect 3219 78 3239 104
rect 2889 -6 2931 42
rect 3061 24 3077 58
rect 3111 24 3141 58
rect 3219 44 3235 78
rect 3273 70 3328 104
rect 3269 44 3328 70
rect 3219 38 3328 44
rect 2923 -40 2931 -6
rect 2889 -56 2931 -40
rect 2993 -8 3027 8
rect 3169 -24 3185 0
rect 3027 -34 3185 -24
rect 3219 -34 3235 0
rect 3027 -42 3235 -34
rect 2993 -58 3235 -42
rect 3269 -20 3334 -4
rect 3303 -54 3334 -20
rect 3269 -92 3334 -54
rect 3368 -16 3402 138
rect 3436 256 3477 272
rect 3470 222 3477 256
rect 3436 152 3477 222
rect 3559 256 3572 282
rect 3743 274 3759 308
rect 3793 274 3809 308
rect 3933 350 3967 366
rect 4027 332 4053 366
rect 4087 332 4103 366
rect 4151 341 4267 375
rect 4301 341 4317 375
rect 4359 368 4393 384
rect 3933 298 3967 316
rect 3847 282 4117 298
rect 3525 222 3538 248
rect 3847 248 3933 282
rect 3967 256 4117 282
rect 3967 248 4083 256
rect 3525 206 3572 222
rect 3612 214 3813 222
rect 3612 180 3617 214
rect 3651 180 3813 214
rect 3612 174 3813 180
rect 3747 172 3813 174
rect 3436 146 3571 152
rect 3436 116 3525 146
rect 3503 112 3525 116
rect 3559 112 3571 146
rect 3747 138 3763 172
rect 3797 138 3813 172
rect 3503 103 3571 112
rect 3619 104 3635 138
rect 3669 104 3685 138
rect 3847 104 3881 248
rect 4067 222 4083 248
rect 4067 206 4117 222
rect 3915 172 3965 188
rect 4151 172 4185 341
rect 4359 284 4393 334
rect 4427 352 4498 418
rect 4427 318 4443 352
rect 4477 318 4498 352
rect 4537 368 4581 384
rect 4537 334 4547 368
rect 4537 300 4581 334
rect 4615 352 4681 418
rect 4615 318 4631 352
rect 4665 318 4681 352
rect 4715 368 4749 384
rect 4219 256 4261 282
rect 4253 248 4261 256
rect 4295 248 4319 282
rect 4359 250 4503 284
rect 4253 222 4319 248
rect 4219 206 4319 222
rect 3949 138 4185 172
rect 3915 122 3959 138
rect 4101 130 4185 138
rect 3503 82 3547 103
rect 3537 48 3547 82
rect 3619 70 3881 104
rect 4001 84 4017 104
rect 3503 32 3547 48
rect 3837 44 3881 70
rect 3985 78 4017 84
rect 4051 70 4067 104
rect 4019 44 4067 70
rect 3769 18 3803 34
rect 3837 10 3853 44
rect 3887 10 3903 44
rect 3985 38 4067 44
rect 3368 -50 3461 -16
rect 3495 -50 3524 -16
rect 3368 -56 3524 -50
rect 3649 -50 3665 -16
rect 3699 -50 3719 -16
rect 3649 -92 3719 -50
rect 3769 -24 3803 -16
rect 3933 -14 3999 -8
rect 3933 -24 3949 -14
rect 3769 -48 3949 -24
rect 3983 -48 3999 -14
rect 3769 -58 3999 -48
rect 4033 -20 4067 -4
rect 4033 -92 4067 -54
rect 4101 -16 4135 130
rect 4169 78 4189 94
rect 4223 60 4239 94
rect 4203 44 4239 60
rect 4169 20 4239 44
rect 4275 82 4319 206
rect 4353 149 4435 216
rect 4353 115 4360 149
rect 4394 142 4435 149
rect 4394 115 4401 142
rect 4353 108 4401 115
rect 4353 92 4435 108
rect 4275 48 4285 82
rect 4469 56 4503 250
rect 4275 32 4319 48
rect 4359 18 4503 56
rect 4537 282 4547 300
rect 4715 300 4749 334
rect 4571 248 4581 266
rect 4359 2 4393 18
rect 4101 -50 4254 -16
rect 4288 -50 4304 -16
rect 4537 10 4581 248
rect 4616 266 4715 284
rect 4616 250 4749 266
rect 4801 342 4853 384
rect 4801 308 4811 342
rect 4845 340 4853 342
rect 4801 306 4819 308
rect 4801 272 4853 306
rect 4616 155 4662 250
rect 4801 238 4819 272
rect 4887 364 4945 418
rect 4887 330 4903 364
rect 4937 330 4945 364
rect 4887 296 4945 330
rect 4887 262 4903 296
rect 4937 262 4945 296
rect 4887 244 4945 262
rect 4981 358 5044 374
rect 4981 324 4998 358
rect 5032 324 5044 358
rect 4981 290 5044 324
rect 4981 256 4998 290
rect 5032 256 5044 290
rect 4616 121 4617 155
rect 4651 121 4662 155
rect 4616 78 4662 121
rect 4697 205 4767 216
rect 4697 171 4708 205
rect 4742 171 4767 205
rect 4697 155 4767 171
rect 4697 121 4719 155
rect 4753 121 4767 155
rect 4697 86 4767 121
rect 4801 182 4853 238
rect 4616 44 4628 78
rect 4801 56 4843 182
rect 4981 156 5044 256
rect 4877 140 5044 156
rect 4911 106 5044 140
rect 4877 90 5044 106
rect 4662 44 4749 52
rect 4616 18 4749 44
rect 4359 -48 4393 -32
rect 4101 -56 4304 -50
rect 4427 -50 4443 -16
rect 4477 -50 4498 -16
rect 4537 -24 4547 10
rect 4715 10 4749 18
rect 4537 -40 4581 -24
rect 4427 -92 4498 -50
rect 4615 -50 4631 -16
rect 4665 -50 4681 -16
rect 4715 -40 4749 -24
rect 4801 20 4853 56
rect 4801 -14 4819 20
rect 4981 10 5044 90
rect 4615 -92 4681 -50
rect 4801 -58 4853 -14
rect 4887 -16 4946 0
rect 4887 -50 4903 -16
rect 4937 -50 4946 -16
rect 4887 -92 4946 -50
rect 4981 -24 4998 10
rect 5032 -24 5044 10
rect 4981 -58 5044 -24
rect 5079 339 5136 384
rect 5170 376 5448 418
rect 5170 342 5186 376
rect 5220 342 5388 376
rect 5422 342 5448 376
rect 5636 376 5712 418
rect 5554 350 5588 366
rect 5079 305 5102 339
rect 5636 342 5662 376
rect 5696 342 5712 376
rect 6135 376 6201 418
rect 5554 308 5588 316
rect 5760 341 5876 375
rect 5910 341 5926 375
rect 6135 342 6151 376
rect 6185 342 6201 376
rect 6419 366 6495 418
rect 5079 276 5136 305
rect 5079 242 5089 276
rect 5123 271 5136 276
rect 5079 237 5102 242
rect 5079 217 5136 237
rect 5170 274 5726 308
rect 5079 34 5115 217
rect 5170 156 5204 274
rect 5265 206 5284 240
rect 5318 214 5422 240
rect 5318 206 5371 214
rect 5365 180 5371 206
rect 5405 180 5422 214
rect 5365 172 5422 180
rect 5151 140 5204 156
rect 5185 106 5204 140
rect 5238 150 5329 156
rect 5238 144 5284 150
rect 5238 110 5279 144
rect 5318 116 5329 150
rect 5313 110 5329 116
rect 5365 138 5388 172
rect 5365 113 5422 138
rect 5151 90 5204 106
rect 5365 76 5409 113
rect 5079 18 5136 34
rect 5079 -16 5102 18
rect 5079 -58 5136 -16
rect 5170 -16 5231 52
rect 5170 -50 5186 -16
rect 5220 -50 5231 -16
rect 5170 -92 5231 -50
rect 5281 42 5409 76
rect 5456 59 5490 274
rect 5676 256 5726 274
rect 5676 222 5692 256
rect 5676 206 5726 222
rect 5760 172 5794 341
rect 6135 308 6201 342
rect 5917 282 5964 288
rect 5524 156 5794 172
rect 5558 138 5794 156
rect 5558 122 5568 138
rect 5524 106 5568 122
rect 5453 58 5490 59
rect 5611 78 5631 104
rect 5281 -6 5323 42
rect 5453 24 5469 58
rect 5503 24 5533 58
rect 5611 44 5627 78
rect 5665 70 5720 104
rect 5661 44 5720 70
rect 5611 38 5720 44
rect 5315 -40 5323 -6
rect 5281 -56 5323 -40
rect 5385 -8 5419 8
rect 5561 -24 5577 0
rect 5419 -34 5577 -24
rect 5611 -34 5627 0
rect 5419 -42 5627 -34
rect 5385 -58 5627 -42
rect 5661 -20 5726 -4
rect 5695 -54 5726 -20
rect 5661 -92 5726 -54
rect 5760 -16 5794 138
rect 5828 256 5869 272
rect 5862 222 5869 256
rect 5828 152 5869 222
rect 5951 256 5964 282
rect 6135 274 6151 308
rect 6185 274 6201 308
rect 6325 350 6359 366
rect 6419 332 6445 366
rect 6479 332 6495 366
rect 6543 341 6659 375
rect 6693 341 6709 375
rect 6751 368 6785 384
rect 6325 298 6359 316
rect 6239 282 6509 298
rect 5917 222 5930 248
rect 6239 248 6325 282
rect 6359 256 6509 282
rect 6359 248 6475 256
rect 5917 206 5964 222
rect 6004 214 6205 222
rect 6004 180 6009 214
rect 6043 180 6205 214
rect 6004 174 6205 180
rect 6139 172 6205 174
rect 5828 146 5963 152
rect 5828 116 5917 146
rect 5895 112 5917 116
rect 5951 112 5963 146
rect 6139 138 6155 172
rect 6189 138 6205 172
rect 5895 103 5963 112
rect 6011 104 6027 138
rect 6061 104 6077 138
rect 6239 104 6273 248
rect 6459 222 6475 248
rect 6459 206 6509 222
rect 6307 172 6357 188
rect 6543 172 6577 341
rect 6751 284 6785 334
rect 6819 352 6890 418
rect 6819 318 6835 352
rect 6869 318 6890 352
rect 6929 368 6973 384
rect 6929 334 6939 368
rect 6929 300 6973 334
rect 7007 352 7073 418
rect 7007 318 7023 352
rect 7057 318 7073 352
rect 7107 368 7141 384
rect 6611 256 6653 282
rect 6645 248 6653 256
rect 6687 248 6711 282
rect 6751 250 6895 284
rect 6645 222 6711 248
rect 6611 206 6711 222
rect 6341 138 6577 172
rect 6307 122 6351 138
rect 6493 130 6577 138
rect 5895 82 5939 103
rect 5929 48 5939 82
rect 6011 70 6273 104
rect 6393 84 6409 104
rect 5895 32 5939 48
rect 6229 44 6273 70
rect 6377 78 6409 84
rect 6443 70 6459 104
rect 6411 44 6459 70
rect 6161 18 6195 34
rect 6229 10 6245 44
rect 6279 10 6295 44
rect 6377 38 6459 44
rect 5760 -50 5853 -16
rect 5887 -50 5916 -16
rect 5760 -56 5916 -50
rect 6041 -50 6057 -16
rect 6091 -50 6111 -16
rect 6041 -92 6111 -50
rect 6161 -24 6195 -16
rect 6325 -14 6391 -8
rect 6325 -24 6341 -14
rect 6161 -48 6341 -24
rect 6375 -48 6391 -14
rect 6161 -58 6391 -48
rect 6425 -20 6459 -4
rect 6425 -92 6459 -54
rect 6493 -16 6527 130
rect 6561 78 6581 94
rect 6615 60 6631 94
rect 6595 44 6631 60
rect 6561 20 6631 44
rect 6667 82 6711 206
rect 6745 150 6827 216
rect 6745 116 6751 150
rect 6785 142 6827 150
rect 6785 116 6793 142
rect 6745 108 6793 116
rect 6745 92 6827 108
rect 6667 48 6677 82
rect 6861 56 6895 250
rect 6667 32 6711 48
rect 6751 18 6895 56
rect 6929 282 6939 300
rect 7107 300 7141 334
rect 6963 248 6973 266
rect 6751 2 6785 18
rect 6493 -50 6646 -16
rect 6680 -50 6696 -16
rect 6929 10 6973 248
rect 7008 266 7107 284
rect 7008 250 7141 266
rect 7193 342 7245 384
rect 7193 308 7202 342
rect 7236 340 7245 342
rect 7193 306 7211 308
rect 7193 272 7245 306
rect 7008 155 7054 250
rect 7193 238 7211 272
rect 7279 364 7337 418
rect 7279 330 7295 364
rect 7329 330 7337 364
rect 7279 296 7337 330
rect 7279 262 7295 296
rect 7329 262 7337 296
rect 7279 244 7337 262
rect 7373 358 7436 374
rect 7373 324 7390 358
rect 7424 324 7436 358
rect 7373 290 7436 324
rect 7373 256 7390 290
rect 7424 256 7436 290
rect 7008 121 7009 155
rect 7043 121 7054 155
rect 7008 78 7054 121
rect 7089 207 7159 216
rect 7089 173 7098 207
rect 7132 173 7159 207
rect 7089 155 7159 173
rect 7089 121 7111 155
rect 7145 121 7159 155
rect 7089 86 7159 121
rect 7193 182 7245 238
rect 7008 44 7020 78
rect 7193 56 7235 182
rect 7373 156 7436 256
rect 7269 140 7436 156
rect 7303 106 7436 140
rect 7269 90 7436 106
rect 7054 44 7141 52
rect 7008 18 7141 44
rect 6751 -48 6785 -32
rect 6493 -56 6696 -50
rect 6819 -50 6835 -16
rect 6869 -50 6890 -16
rect 6929 -24 6939 10
rect 7107 10 7141 18
rect 6929 -40 6973 -24
rect 6819 -92 6890 -50
rect 7007 -50 7023 -16
rect 7057 -50 7073 -16
rect 7107 -40 7141 -24
rect 7193 20 7245 56
rect 7193 -14 7211 20
rect 7373 10 7436 90
rect 7007 -92 7073 -50
rect 7193 -58 7245 -14
rect 7279 -16 7338 0
rect 7279 -50 7295 -16
rect 7329 -50 7338 -16
rect 7279 -92 7338 -50
rect 7373 -24 7390 10
rect 7424 -24 7436 10
rect 7373 -58 7436 -24
rect 7471 339 7528 384
rect 7562 376 7840 418
rect 7562 342 7578 376
rect 7612 342 7780 376
rect 7814 342 7840 376
rect 8028 376 8104 418
rect 7946 350 7980 366
rect 7471 305 7494 339
rect 8028 342 8054 376
rect 8088 342 8104 376
rect 8527 376 8593 418
rect 7946 308 7980 316
rect 8152 341 8268 375
rect 8302 341 8318 375
rect 8527 342 8543 376
rect 8577 342 8593 376
rect 8811 366 8887 418
rect 7471 276 7528 305
rect 7471 242 7482 276
rect 7516 271 7528 276
rect 7471 237 7494 242
rect 7471 217 7528 237
rect 7562 274 8118 308
rect 7471 34 7507 217
rect 7562 156 7596 274
rect 7657 206 7676 240
rect 7710 214 7814 240
rect 7710 206 7763 214
rect 7757 180 7763 206
rect 7797 180 7814 214
rect 7757 172 7814 180
rect 7543 140 7596 156
rect 7577 106 7596 140
rect 7630 150 7721 156
rect 7630 144 7677 150
rect 7630 110 7671 144
rect 7711 116 7721 150
rect 7705 110 7721 116
rect 7757 138 7780 172
rect 7757 113 7814 138
rect 7543 90 7596 106
rect 7757 76 7801 113
rect 7471 18 7528 34
rect 7471 -16 7494 18
rect 7471 -58 7528 -16
rect 7562 -16 7623 52
rect 7562 -50 7578 -16
rect 7612 -50 7623 -16
rect 7562 -92 7623 -50
rect 7673 42 7801 76
rect 7848 59 7882 274
rect 8068 256 8118 274
rect 8068 222 8084 256
rect 8068 206 8118 222
rect 8152 172 8186 341
rect 8527 308 8593 342
rect 8309 282 8356 288
rect 7916 156 8186 172
rect 7950 138 8186 156
rect 7950 122 7960 138
rect 7916 106 7960 122
rect 7845 58 7882 59
rect 8003 78 8023 104
rect 7673 -6 7715 42
rect 7845 24 7861 58
rect 7895 24 7925 58
rect 8003 44 8019 78
rect 8057 70 8112 104
rect 8053 44 8112 70
rect 8003 38 8112 44
rect 7707 -40 7715 -6
rect 7673 -56 7715 -40
rect 7777 -8 7811 8
rect 7953 -24 7969 0
rect 7811 -34 7969 -24
rect 8003 -34 8019 0
rect 7811 -42 8019 -34
rect 7777 -58 8019 -42
rect 8053 -20 8118 -4
rect 8087 -54 8118 -20
rect 8053 -92 8118 -54
rect 8152 -16 8186 138
rect 8220 256 8261 272
rect 8254 222 8261 256
rect 8220 152 8261 222
rect 8343 256 8356 282
rect 8527 274 8543 308
rect 8577 274 8593 308
rect 8717 350 8751 366
rect 8811 332 8837 366
rect 8871 332 8887 366
rect 8935 341 9051 375
rect 9085 341 9101 375
rect 9143 368 9177 384
rect 8717 298 8751 316
rect 8631 282 8901 298
rect 8309 222 8322 248
rect 8631 248 8717 282
rect 8751 256 8901 282
rect 8751 248 8867 256
rect 8309 206 8356 222
rect 8396 214 8597 222
rect 8396 180 8401 214
rect 8435 180 8597 214
rect 8396 174 8597 180
rect 8531 172 8597 174
rect 8220 146 8355 152
rect 8220 116 8309 146
rect 8287 112 8309 116
rect 8343 112 8355 146
rect 8531 138 8547 172
rect 8581 138 8597 172
rect 8287 103 8355 112
rect 8403 104 8419 138
rect 8453 104 8469 138
rect 8631 104 8665 248
rect 8851 222 8867 248
rect 8851 206 8901 222
rect 8699 172 8749 188
rect 8935 172 8969 341
rect 9143 284 9177 334
rect 9211 352 9282 418
rect 9211 318 9227 352
rect 9261 318 9282 352
rect 9321 368 9365 384
rect 9321 334 9331 368
rect 9321 300 9365 334
rect 9399 352 9465 418
rect 9399 318 9415 352
rect 9449 318 9465 352
rect 9499 368 9533 384
rect 9003 256 9045 282
rect 9037 248 9045 256
rect 9079 248 9103 282
rect 9143 250 9287 284
rect 9037 222 9103 248
rect 9003 206 9103 222
rect 8733 138 8969 172
rect 8699 122 8743 138
rect 8885 130 8969 138
rect 8287 82 8331 103
rect 8321 48 8331 82
rect 8403 70 8665 104
rect 8785 84 8801 104
rect 8287 32 8331 48
rect 8621 44 8665 70
rect 8769 78 8801 84
rect 8835 70 8851 104
rect 8803 44 8851 70
rect 8553 18 8587 34
rect 8621 10 8637 44
rect 8671 10 8687 44
rect 8769 38 8851 44
rect 8152 -50 8245 -16
rect 8279 -50 8308 -16
rect 8152 -56 8308 -50
rect 8433 -50 8449 -16
rect 8483 -50 8503 -16
rect 8433 -92 8503 -50
rect 8553 -24 8587 -16
rect 8717 -14 8783 -8
rect 8717 -24 8733 -14
rect 8553 -48 8733 -24
rect 8767 -48 8783 -14
rect 8553 -58 8783 -48
rect 8817 -20 8851 -4
rect 8817 -92 8851 -54
rect 8885 -16 8919 130
rect 8953 78 8973 94
rect 9007 60 9023 94
rect 8987 44 9023 60
rect 8953 20 9023 44
rect 9059 82 9103 206
rect 9137 149 9219 216
rect 9137 115 9144 149
rect 9178 142 9219 149
rect 9178 115 9185 142
rect 9137 108 9185 115
rect 9137 92 9219 108
rect 9059 48 9069 82
rect 9253 56 9287 250
rect 9059 32 9103 48
rect 9143 18 9287 56
rect 9321 282 9331 300
rect 9499 300 9533 334
rect 9355 248 9365 266
rect 9143 2 9177 18
rect 8885 -50 9038 -16
rect 9072 -50 9088 -16
rect 9321 10 9365 248
rect 9400 266 9499 284
rect 9400 250 9533 266
rect 9585 341 9637 384
rect 9585 307 9594 341
rect 9628 340 9637 341
rect 9585 306 9603 307
rect 9585 272 9637 306
rect 9400 155 9446 250
rect 9585 238 9603 272
rect 9671 364 9729 418
rect 9671 330 9687 364
rect 9721 330 9729 364
rect 9671 296 9729 330
rect 9671 262 9687 296
rect 9721 262 9729 296
rect 9671 244 9729 262
rect 9765 358 9828 374
rect 9765 324 9782 358
rect 9816 324 9828 358
rect 9765 290 9828 324
rect 9765 256 9782 290
rect 9816 256 9828 290
rect 9400 121 9401 155
rect 9435 121 9446 155
rect 9400 78 9446 121
rect 9481 205 9551 216
rect 9481 171 9490 205
rect 9524 171 9551 205
rect 9481 155 9551 171
rect 9481 121 9503 155
rect 9537 121 9551 155
rect 9481 86 9551 121
rect 9585 182 9637 238
rect 9400 44 9412 78
rect 9585 56 9627 182
rect 9765 156 9828 256
rect 9661 140 9828 156
rect 9695 106 9828 140
rect 9661 90 9828 106
rect 9446 44 9533 52
rect 9400 18 9533 44
rect 9143 -48 9177 -32
rect 8885 -56 9088 -50
rect 9211 -50 9227 -16
rect 9261 -50 9282 -16
rect 9321 -24 9331 10
rect 9499 10 9533 18
rect 9321 -40 9365 -24
rect 9211 -92 9282 -50
rect 9399 -50 9415 -16
rect 9449 -50 9465 -16
rect 9499 -40 9533 -24
rect 9585 20 9637 56
rect 9585 -14 9603 20
rect 9765 10 9828 90
rect 9399 -92 9465 -50
rect 9585 -58 9637 -14
rect 9671 -16 9730 0
rect 9671 -50 9687 -16
rect 9721 -50 9730 -16
rect 9671 -92 9730 -50
rect 9765 -24 9782 10
rect 9816 -24 9828 10
rect 9765 -58 9828 -24
rect 9863 339 9920 384
rect 9954 376 10232 418
rect 9954 342 9970 376
rect 10004 342 10172 376
rect 10206 342 10232 376
rect 10420 376 10496 418
rect 10338 350 10372 366
rect 9863 305 9886 339
rect 10420 342 10446 376
rect 10480 342 10496 376
rect 10919 376 10985 418
rect 10338 308 10372 316
rect 10544 341 10660 375
rect 10694 341 10710 375
rect 10919 342 10935 376
rect 10969 342 10985 376
rect 11203 366 11279 418
rect 9863 276 9920 305
rect 9863 242 9874 276
rect 9908 271 9920 276
rect 9863 237 9886 242
rect 9863 217 9920 237
rect 9954 274 10510 308
rect 9863 34 9899 217
rect 9954 156 9988 274
rect 10049 206 10068 240
rect 10102 214 10206 240
rect 10102 206 10155 214
rect 10149 180 10155 206
rect 10189 180 10206 214
rect 10149 172 10206 180
rect 9935 140 9988 156
rect 9969 106 9988 140
rect 10022 150 10113 156
rect 10022 144 10068 150
rect 10022 110 10063 144
rect 10102 116 10113 150
rect 10097 110 10113 116
rect 10149 138 10172 172
rect 10149 113 10206 138
rect 9935 90 9988 106
rect 10149 76 10193 113
rect 9863 18 9920 34
rect 9863 -16 9886 18
rect 9863 -58 9920 -16
rect 9954 -16 10015 52
rect 9954 -50 9970 -16
rect 10004 -50 10015 -16
rect 9954 -92 10015 -50
rect 10065 42 10193 76
rect 10240 59 10274 274
rect 10460 256 10510 274
rect 10460 222 10476 256
rect 10460 206 10510 222
rect 10544 172 10578 341
rect 10919 308 10985 342
rect 10701 282 10748 288
rect 10308 156 10578 172
rect 10342 138 10578 156
rect 10342 122 10352 138
rect 10308 106 10352 122
rect 10237 58 10274 59
rect 10395 78 10415 104
rect 10065 -6 10107 42
rect 10237 24 10253 58
rect 10287 24 10317 58
rect 10395 44 10411 78
rect 10449 70 10504 104
rect 10445 44 10504 70
rect 10395 38 10504 44
rect 10099 -40 10107 -6
rect 10065 -56 10107 -40
rect 10169 -8 10203 8
rect 10345 -24 10361 0
rect 10203 -34 10361 -24
rect 10395 -34 10411 0
rect 10203 -42 10411 -34
rect 10169 -58 10411 -42
rect 10445 -20 10510 -4
rect 10479 -54 10510 -20
rect 10445 -92 10510 -54
rect 10544 -16 10578 138
rect 10612 256 10653 272
rect 10646 222 10653 256
rect 10612 152 10653 222
rect 10735 256 10748 282
rect 10919 274 10935 308
rect 10969 274 10985 308
rect 11109 350 11143 366
rect 11203 332 11229 366
rect 11263 332 11279 366
rect 11327 341 11443 375
rect 11477 341 11493 375
rect 11535 368 11569 384
rect 11109 298 11143 316
rect 11023 282 11293 298
rect 10701 222 10714 248
rect 11023 248 11109 282
rect 11143 256 11293 282
rect 11143 248 11259 256
rect 10701 206 10748 222
rect 10788 214 10989 222
rect 10788 180 10793 214
rect 10827 180 10989 214
rect 10788 174 10989 180
rect 10923 172 10989 174
rect 10612 146 10747 152
rect 10612 116 10701 146
rect 10679 112 10701 116
rect 10735 112 10747 146
rect 10923 138 10939 172
rect 10973 138 10989 172
rect 10679 103 10747 112
rect 10795 104 10811 138
rect 10845 104 10861 138
rect 11023 104 11057 248
rect 11243 222 11259 248
rect 11243 206 11293 222
rect 11091 172 11141 188
rect 11327 172 11361 341
rect 11535 284 11569 334
rect 11603 352 11674 418
rect 11603 318 11619 352
rect 11653 318 11674 352
rect 11713 368 11757 384
rect 11713 334 11723 368
rect 11713 300 11757 334
rect 11791 352 11857 418
rect 11791 318 11807 352
rect 11841 318 11857 352
rect 11891 368 11925 384
rect 11395 256 11437 282
rect 11429 248 11437 256
rect 11471 248 11495 282
rect 11535 250 11679 284
rect 11429 222 11495 248
rect 11395 206 11495 222
rect 11125 138 11361 172
rect 11091 122 11135 138
rect 11277 130 11361 138
rect 10679 82 10723 103
rect 10713 48 10723 82
rect 10795 70 11057 104
rect 11177 84 11193 104
rect 10679 32 10723 48
rect 11013 44 11057 70
rect 11161 78 11193 84
rect 11227 70 11243 104
rect 11195 44 11243 70
rect 10945 18 10979 34
rect 11013 10 11029 44
rect 11063 10 11079 44
rect 11161 38 11243 44
rect 10544 -50 10637 -16
rect 10671 -50 10700 -16
rect 10544 -56 10700 -50
rect 10825 -50 10841 -16
rect 10875 -50 10895 -16
rect 10825 -92 10895 -50
rect 10945 -24 10979 -16
rect 11109 -14 11175 -8
rect 11109 -24 11125 -14
rect 10945 -48 11125 -24
rect 11159 -48 11175 -14
rect 10945 -58 11175 -48
rect 11209 -20 11243 -4
rect 11209 -92 11243 -54
rect 11277 -16 11311 130
rect 11345 78 11365 94
rect 11399 60 11415 94
rect 11379 44 11415 60
rect 11345 20 11415 44
rect 11451 82 11495 206
rect 11529 149 11611 216
rect 11529 115 11535 149
rect 11569 142 11611 149
rect 11569 115 11577 142
rect 11529 108 11577 115
rect 11529 92 11611 108
rect 11451 48 11461 82
rect 11645 56 11679 250
rect 11451 32 11495 48
rect 11535 18 11679 56
rect 11713 282 11723 300
rect 11891 300 11925 334
rect 11747 248 11757 266
rect 11535 2 11569 18
rect 11277 -50 11430 -16
rect 11464 -50 11480 -16
rect 11713 10 11757 248
rect 11792 266 11891 284
rect 11792 250 11925 266
rect 11977 343 12029 384
rect 11977 309 11987 343
rect 12021 340 12029 343
rect 11977 306 11995 309
rect 11977 272 12029 306
rect 11792 155 11838 250
rect 11977 238 11995 272
rect 12063 364 12121 418
rect 12063 330 12079 364
rect 12113 330 12121 364
rect 12063 296 12121 330
rect 12063 262 12079 296
rect 12113 262 12121 296
rect 12063 244 12121 262
rect 12157 358 12220 374
rect 12157 324 12174 358
rect 12208 324 12220 358
rect 12157 290 12220 324
rect 12157 256 12174 290
rect 12208 256 12220 290
rect 11792 121 11793 155
rect 11827 121 11838 155
rect 11792 78 11838 121
rect 11873 207 11943 216
rect 11873 173 11882 207
rect 11916 173 11943 207
rect 11873 155 11943 173
rect 11873 121 11895 155
rect 11929 121 11943 155
rect 11873 86 11943 121
rect 11977 182 12029 238
rect 11792 44 11804 78
rect 11977 56 12019 182
rect 12157 156 12220 256
rect 12053 140 12220 156
rect 12087 106 12220 140
rect 12053 90 12220 106
rect 11838 44 11925 52
rect 11792 18 11925 44
rect 11535 -48 11569 -32
rect 11277 -56 11480 -50
rect 11603 -50 11619 -16
rect 11653 -50 11674 -16
rect 11713 -24 11723 10
rect 11891 10 11925 18
rect 11713 -40 11757 -24
rect 11603 -92 11674 -50
rect 11791 -50 11807 -16
rect 11841 -50 11857 -16
rect 11891 -40 11925 -24
rect 11977 20 12029 56
rect 11977 -14 11995 20
rect 12157 10 12220 90
rect 11791 -92 11857 -50
rect 11977 -58 12029 -14
rect 12063 -16 12122 0
rect 12063 -50 12079 -16
rect 12113 -50 12122 -16
rect 12063 -92 12122 -50
rect 12157 -24 12174 10
rect 12208 -24 12220 10
rect 12157 -58 12220 -24
rect 12255 339 12312 384
rect 12346 376 12624 418
rect 12346 342 12362 376
rect 12396 342 12564 376
rect 12598 342 12624 376
rect 12812 376 12888 418
rect 12730 350 12764 366
rect 12255 305 12278 339
rect 12812 342 12838 376
rect 12872 342 12888 376
rect 13311 376 13377 418
rect 12730 308 12764 316
rect 12936 341 13052 375
rect 13086 341 13102 375
rect 13311 342 13327 376
rect 13361 342 13377 376
rect 13595 366 13671 418
rect 12255 277 12312 305
rect 12255 243 12265 277
rect 12299 271 12312 277
rect 12255 237 12278 243
rect 12255 217 12312 237
rect 12346 274 12902 308
rect 12255 34 12291 217
rect 12346 156 12380 274
rect 12441 206 12460 240
rect 12494 214 12598 240
rect 12494 206 12547 214
rect 12541 180 12547 206
rect 12581 180 12598 214
rect 12541 172 12598 180
rect 12327 140 12380 156
rect 12361 106 12380 140
rect 12414 150 12505 156
rect 12414 144 12461 150
rect 12414 110 12455 144
rect 12495 116 12505 150
rect 12489 110 12505 116
rect 12541 138 12564 172
rect 12541 113 12598 138
rect 12327 90 12380 106
rect 12541 76 12585 113
rect 12255 18 12312 34
rect 12255 -16 12278 18
rect 12255 -58 12312 -16
rect 12346 -16 12407 52
rect 12346 -50 12362 -16
rect 12396 -50 12407 -16
rect 12346 -92 12407 -50
rect 12457 42 12585 76
rect 12632 59 12666 274
rect 12852 256 12902 274
rect 12852 222 12868 256
rect 12852 206 12902 222
rect 12936 172 12970 341
rect 13311 308 13377 342
rect 13093 282 13140 288
rect 12700 156 12970 172
rect 12734 138 12970 156
rect 12734 122 12744 138
rect 12700 106 12744 122
rect 12629 58 12666 59
rect 12787 78 12807 104
rect 12457 -6 12499 42
rect 12629 24 12645 58
rect 12679 24 12709 58
rect 12787 44 12803 78
rect 12841 70 12896 104
rect 12837 44 12896 70
rect 12787 38 12896 44
rect 12491 -40 12499 -6
rect 12457 -56 12499 -40
rect 12561 -8 12595 8
rect 12737 -24 12753 0
rect 12595 -34 12753 -24
rect 12787 -34 12803 0
rect 12595 -42 12803 -34
rect 12561 -58 12803 -42
rect 12837 -20 12902 -4
rect 12871 -54 12902 -20
rect 12837 -92 12902 -54
rect 12936 -16 12970 138
rect 13004 256 13045 272
rect 13038 222 13045 256
rect 13004 152 13045 222
rect 13127 256 13140 282
rect 13311 274 13327 308
rect 13361 274 13377 308
rect 13501 350 13535 366
rect 13595 332 13621 366
rect 13655 332 13671 366
rect 13719 341 13835 375
rect 13869 341 13885 375
rect 13927 368 13961 384
rect 13501 298 13535 316
rect 13415 282 13685 298
rect 13093 222 13106 248
rect 13415 248 13501 282
rect 13535 256 13685 282
rect 13535 248 13651 256
rect 13093 206 13140 222
rect 13180 214 13381 222
rect 13180 180 13185 214
rect 13219 180 13381 214
rect 13180 174 13381 180
rect 13315 172 13381 174
rect 13004 146 13139 152
rect 13004 116 13093 146
rect 13071 112 13093 116
rect 13127 112 13139 146
rect 13315 138 13331 172
rect 13365 138 13381 172
rect 13071 103 13139 112
rect 13187 104 13203 138
rect 13237 104 13253 138
rect 13415 104 13449 248
rect 13635 222 13651 248
rect 13635 206 13685 222
rect 13483 172 13533 188
rect 13719 172 13753 341
rect 13927 284 13961 334
rect 13995 352 14066 418
rect 13995 318 14011 352
rect 14045 318 14066 352
rect 14105 368 14149 384
rect 14105 334 14115 368
rect 14105 300 14149 334
rect 14183 352 14249 418
rect 14183 318 14199 352
rect 14233 318 14249 352
rect 14283 368 14317 384
rect 13787 256 13829 282
rect 13821 248 13829 256
rect 13863 248 13887 282
rect 13927 250 14071 284
rect 13821 222 13887 248
rect 13787 206 13887 222
rect 13517 138 13753 172
rect 13483 122 13527 138
rect 13669 130 13753 138
rect 13071 82 13115 103
rect 13105 48 13115 82
rect 13187 70 13449 104
rect 13569 84 13585 104
rect 13071 32 13115 48
rect 13405 44 13449 70
rect 13553 78 13585 84
rect 13619 70 13635 104
rect 13587 44 13635 70
rect 13337 18 13371 34
rect 13405 10 13421 44
rect 13455 10 13471 44
rect 13553 38 13635 44
rect 12936 -50 13029 -16
rect 13063 -50 13092 -16
rect 12936 -56 13092 -50
rect 13217 -50 13233 -16
rect 13267 -50 13287 -16
rect 13217 -92 13287 -50
rect 13337 -24 13371 -16
rect 13501 -14 13567 -8
rect 13501 -24 13517 -14
rect 13337 -48 13517 -24
rect 13551 -48 13567 -14
rect 13337 -58 13567 -48
rect 13601 -20 13635 -4
rect 13601 -92 13635 -54
rect 13669 -16 13703 130
rect 13737 78 13757 94
rect 13791 60 13807 94
rect 13771 44 13807 60
rect 13737 20 13807 44
rect 13843 82 13887 206
rect 13921 149 14003 216
rect 13921 115 13928 149
rect 13962 142 14003 149
rect 13962 115 13969 142
rect 13921 108 13969 115
rect 13921 92 14003 108
rect 13843 48 13853 82
rect 14037 56 14071 250
rect 13843 32 13887 48
rect 13927 18 14071 56
rect 14105 282 14115 300
rect 14283 300 14317 334
rect 14139 248 14149 266
rect 13927 2 13961 18
rect 13669 -50 13822 -16
rect 13856 -50 13872 -16
rect 14105 10 14149 248
rect 14184 266 14283 284
rect 14184 250 14317 266
rect 14369 343 14421 384
rect 14369 309 14378 343
rect 14412 340 14421 343
rect 14369 306 14387 309
rect 14369 272 14421 306
rect 14184 155 14230 250
rect 14369 238 14387 272
rect 14455 364 14513 418
rect 14455 330 14471 364
rect 14505 330 14513 364
rect 14455 296 14513 330
rect 14455 262 14471 296
rect 14505 262 14513 296
rect 14455 244 14513 262
rect 14549 358 14612 374
rect 14549 324 14566 358
rect 14600 324 14612 358
rect 14549 290 14612 324
rect 14549 256 14566 290
rect 14600 256 14612 290
rect 14184 121 14185 155
rect 14219 121 14230 155
rect 14184 78 14230 121
rect 14265 205 14335 216
rect 14265 171 14274 205
rect 14308 171 14335 205
rect 14265 155 14335 171
rect 14265 121 14287 155
rect 14321 121 14335 155
rect 14265 86 14335 121
rect 14369 182 14421 238
rect 14184 44 14196 78
rect 14369 56 14411 182
rect 14549 156 14612 256
rect 14445 140 14612 156
rect 14479 106 14612 140
rect 14445 90 14612 106
rect 14230 44 14317 52
rect 14184 18 14317 44
rect 13927 -48 13961 -32
rect 13669 -56 13872 -50
rect 13995 -50 14011 -16
rect 14045 -50 14066 -16
rect 14105 -24 14115 10
rect 14283 10 14317 18
rect 14105 -40 14149 -24
rect 13995 -92 14066 -50
rect 14183 -50 14199 -16
rect 14233 -50 14249 -16
rect 14283 -40 14317 -24
rect 14369 20 14421 56
rect 14369 -14 14387 20
rect 14549 10 14612 90
rect 14183 -92 14249 -50
rect 14369 -58 14421 -14
rect 14455 -16 14514 0
rect 14455 -50 14471 -16
rect 14505 -50 14514 -16
rect 14455 -92 14514 -50
rect 14549 -24 14566 10
rect 14600 -24 14612 10
rect 14549 -58 14612 -24
rect 14647 339 14704 384
rect 14738 376 15016 418
rect 14738 342 14754 376
rect 14788 342 14956 376
rect 14990 342 15016 376
rect 15204 376 15280 418
rect 15122 350 15156 366
rect 14647 305 14670 339
rect 15204 342 15230 376
rect 15264 342 15280 376
rect 15703 376 15769 418
rect 15122 308 15156 316
rect 15328 341 15444 375
rect 15478 341 15494 375
rect 15703 342 15719 376
rect 15753 342 15769 376
rect 15987 366 16063 418
rect 14647 276 14704 305
rect 14647 242 14658 276
rect 14692 271 14704 276
rect 14647 237 14670 242
rect 14647 217 14704 237
rect 14738 274 15294 308
rect 14647 34 14683 217
rect 14738 156 14772 274
rect 14833 206 14852 240
rect 14886 214 14990 240
rect 14886 206 14939 214
rect 14933 180 14939 206
rect 14973 180 14990 214
rect 14933 172 14990 180
rect 14719 140 14772 156
rect 14753 106 14772 140
rect 14806 150 14897 156
rect 14806 144 14852 150
rect 14806 110 14847 144
rect 14886 116 14897 150
rect 14881 110 14897 116
rect 14933 138 14956 172
rect 14933 113 14990 138
rect 14719 90 14772 106
rect 14933 76 14977 113
rect 14647 18 14704 34
rect 14647 -16 14670 18
rect 14647 -58 14704 -16
rect 14738 -16 14799 52
rect 14738 -50 14754 -16
rect 14788 -50 14799 -16
rect 14738 -92 14799 -50
rect 14849 42 14977 76
rect 15024 59 15058 274
rect 15244 256 15294 274
rect 15244 222 15260 256
rect 15244 206 15294 222
rect 15328 172 15362 341
rect 15703 308 15769 342
rect 15485 282 15532 288
rect 15092 156 15362 172
rect 15126 138 15362 156
rect 15126 122 15136 138
rect 15092 106 15136 122
rect 15021 58 15058 59
rect 15179 78 15199 104
rect 14849 -6 14891 42
rect 15021 24 15037 58
rect 15071 24 15101 58
rect 15179 44 15195 78
rect 15233 70 15288 104
rect 15229 44 15288 70
rect 15179 38 15288 44
rect 14883 -40 14891 -6
rect 14849 -56 14891 -40
rect 14953 -8 14987 8
rect 15129 -24 15145 0
rect 14987 -34 15145 -24
rect 15179 -34 15195 0
rect 14987 -42 15195 -34
rect 14953 -58 15195 -42
rect 15229 -20 15294 -4
rect 15263 -54 15294 -20
rect 15229 -92 15294 -54
rect 15328 -16 15362 138
rect 15396 256 15437 272
rect 15430 222 15437 256
rect 15396 152 15437 222
rect 15519 256 15532 282
rect 15703 274 15719 308
rect 15753 274 15769 308
rect 15893 350 15927 366
rect 15987 332 16013 366
rect 16047 332 16063 366
rect 16111 341 16227 375
rect 16261 341 16277 375
rect 16319 368 16353 384
rect 15893 298 15927 316
rect 15807 282 16077 298
rect 15485 222 15498 248
rect 15807 248 15893 282
rect 15927 256 16077 282
rect 15927 248 16043 256
rect 15485 206 15532 222
rect 15572 214 15773 222
rect 15572 180 15577 214
rect 15611 180 15773 214
rect 15572 174 15773 180
rect 15707 172 15773 174
rect 15396 146 15531 152
rect 15396 116 15485 146
rect 15463 112 15485 116
rect 15519 112 15531 146
rect 15707 138 15723 172
rect 15757 138 15773 172
rect 15463 103 15531 112
rect 15579 104 15595 138
rect 15629 104 15645 138
rect 15807 104 15841 248
rect 16027 222 16043 248
rect 16027 206 16077 222
rect 15875 172 15925 188
rect 16111 172 16145 341
rect 16319 284 16353 334
rect 16387 352 16458 418
rect 16387 318 16403 352
rect 16437 318 16458 352
rect 16497 368 16541 384
rect 16497 334 16507 368
rect 16497 300 16541 334
rect 16575 352 16641 418
rect 16575 318 16591 352
rect 16625 318 16641 352
rect 16675 368 16709 384
rect 16179 256 16221 282
rect 16213 248 16221 256
rect 16255 248 16279 282
rect 16319 250 16463 284
rect 16213 222 16279 248
rect 16179 206 16279 222
rect 15909 138 16145 172
rect 15875 122 15919 138
rect 16061 130 16145 138
rect 15463 82 15507 103
rect 15497 48 15507 82
rect 15579 70 15841 104
rect 15961 84 15977 104
rect 15463 32 15507 48
rect 15797 44 15841 70
rect 15945 78 15977 84
rect 16011 70 16027 104
rect 15979 44 16027 70
rect 15729 18 15763 34
rect 15797 10 15813 44
rect 15847 10 15863 44
rect 15945 38 16027 44
rect 15328 -50 15421 -16
rect 15455 -50 15484 -16
rect 15328 -56 15484 -50
rect 15609 -50 15625 -16
rect 15659 -50 15679 -16
rect 15609 -92 15679 -50
rect 15729 -24 15763 -16
rect 15893 -14 15959 -8
rect 15893 -24 15909 -14
rect 15729 -48 15909 -24
rect 15943 -48 15959 -14
rect 15729 -58 15959 -48
rect 15993 -20 16027 -4
rect 15993 -92 16027 -54
rect 16061 -16 16095 130
rect 16129 78 16149 94
rect 16183 60 16199 94
rect 16163 44 16199 60
rect 16129 20 16199 44
rect 16235 82 16279 206
rect 16313 149 16395 216
rect 16313 115 16321 149
rect 16355 142 16395 149
rect 16355 115 16361 142
rect 16313 108 16361 115
rect 16313 92 16395 108
rect 16235 48 16245 82
rect 16429 56 16463 250
rect 16235 32 16279 48
rect 16319 18 16463 56
rect 16497 282 16507 300
rect 16675 300 16709 334
rect 16531 248 16541 266
rect 16319 2 16353 18
rect 16061 -50 16214 -16
rect 16248 -50 16264 -16
rect 16497 10 16541 248
rect 16576 266 16675 284
rect 16576 250 16709 266
rect 16576 155 16622 250
rect 16576 121 16577 155
rect 16611 121 16622 155
rect 16576 78 16622 121
rect 16657 207 16727 216
rect 16657 173 16666 207
rect 16700 173 16727 207
rect 16657 155 16727 173
rect 16657 121 16679 155
rect 16713 121 16727 155
rect 16657 86 16727 121
rect 16576 44 16588 78
rect 16622 44 16709 52
rect 16576 18 16709 44
rect 16319 -48 16353 -32
rect 16061 -56 16264 -50
rect 16387 -50 16403 -16
rect 16437 -50 16458 -16
rect 16497 -24 16507 10
rect 16675 10 16709 18
rect 16497 -40 16541 -24
rect 16387 -92 16458 -50
rect 16575 -50 16591 -16
rect 16625 -50 16641 -16
rect 16675 -40 16709 -24
rect 16575 -92 16641 -50
rect 0 -150 29 -92
rect 63 -150 121 -92
rect 155 -150 213 -92
rect 247 -150 305 -92
rect 339 -150 397 -92
rect 431 -150 489 -92
rect 523 -150 581 -92
rect 615 -150 673 -92
rect 707 -150 765 -92
rect 799 -150 857 -92
rect 891 -150 949 -92
rect 983 -150 1041 -92
rect 1075 -150 1133 -92
rect 1167 -150 1225 -92
rect 1259 -150 1317 -92
rect 1351 -150 1409 -92
rect 1443 -150 1501 -92
rect 1535 -150 1593 -92
rect 1627 -150 1685 -92
rect 1719 -150 1777 -92
rect 1811 -150 1869 -92
rect 1903 -150 1961 -92
rect 1995 -150 2053 -92
rect 2087 -150 2145 -92
rect 2179 -150 2237 -92
rect 2271 -150 2329 -92
rect 2363 -150 2421 -92
rect 2455 -150 2513 -92
rect 2547 -150 2605 -92
rect 2639 -150 2697 -92
rect 2731 -150 2789 -92
rect 2823 -150 2881 -92
rect 2915 -150 2973 -92
rect 3007 -150 3065 -92
rect 3099 -150 3157 -92
rect 3191 -150 3249 -92
rect 3283 -150 3341 -92
rect 3375 -150 3433 -92
rect 3467 -150 3525 -92
rect 3559 -150 3617 -92
rect 3651 -150 3709 -92
rect 3743 -150 3801 -92
rect 3835 -150 3893 -92
rect 3927 -150 3985 -92
rect 4019 -150 4077 -92
rect 4111 -150 4169 -92
rect 4203 -150 4261 -92
rect 4295 -150 4353 -92
rect 4387 -150 4445 -92
rect 4479 -150 4537 -92
rect 4571 -150 4629 -92
rect 4663 -150 4721 -92
rect 4755 -150 4813 -92
rect 4847 -150 4905 -92
rect 4939 -150 4997 -92
rect 5031 -150 5089 -92
rect 5123 -150 5181 -92
rect 5215 -150 5273 -92
rect 5307 -150 5365 -92
rect 5399 -150 5457 -92
rect 5491 -150 5549 -92
rect 5583 -150 5641 -92
rect 5675 -150 5733 -92
rect 5767 -150 5825 -92
rect 5859 -150 5917 -92
rect 5951 -150 6009 -92
rect 6043 -150 6101 -92
rect 6135 -150 6193 -92
rect 6227 -150 6285 -92
rect 6319 -150 6377 -92
rect 6411 -150 6469 -92
rect 6503 -150 6561 -92
rect 6595 -150 6653 -92
rect 6687 -150 6745 -92
rect 6779 -150 6837 -92
rect 6871 -150 6929 -92
rect 6963 -150 7021 -92
rect 7055 -150 7113 -92
rect 7147 -150 7205 -92
rect 7239 -150 7297 -92
rect 7331 -150 7389 -92
rect 7423 -150 7481 -92
rect 7515 -150 7573 -92
rect 7607 -150 7665 -92
rect 7699 -150 7757 -92
rect 7791 -150 7849 -92
rect 7883 -150 7941 -92
rect 7975 -150 8033 -92
rect 8067 -150 8125 -92
rect 8159 -150 8217 -92
rect 8251 -150 8309 -92
rect 8343 -150 8401 -92
rect 8435 -150 8493 -92
rect 8527 -150 8585 -92
rect 8619 -150 8677 -92
rect 8711 -150 8769 -92
rect 8803 -150 8861 -92
rect 8895 -150 8953 -92
rect 8987 -150 9045 -92
rect 9079 -150 9137 -92
rect 9171 -150 9229 -92
rect 9263 -150 9321 -92
rect 9355 -150 9413 -92
rect 9447 -150 9505 -92
rect 9539 -150 9597 -92
rect 9631 -150 9689 -92
rect 9723 -150 9781 -92
rect 9815 -150 9873 -92
rect 9907 -150 9965 -92
rect 9999 -150 10057 -92
rect 10091 -150 10149 -92
rect 10183 -150 10241 -92
rect 10275 -150 10333 -92
rect 10367 -150 10425 -92
rect 10459 -150 10517 -92
rect 10551 -150 10609 -92
rect 10643 -150 10701 -92
rect 10735 -150 10793 -92
rect 10827 -150 10885 -92
rect 10919 -150 10977 -92
rect 11011 -150 11069 -92
rect 11103 -150 11161 -92
rect 11195 -150 11253 -92
rect 11287 -150 11345 -92
rect 11379 -150 11437 -92
rect 11471 -150 11529 -92
rect 11563 -150 11621 -92
rect 11655 -150 11713 -92
rect 11747 -150 11805 -92
rect 11839 -150 11897 -92
rect 11931 -150 11989 -92
rect 12023 -150 12081 -92
rect 12115 -150 12173 -92
rect 12207 -150 12265 -92
rect 12299 -150 12357 -92
rect 12391 -150 12449 -92
rect 12483 -150 12541 -92
rect 12575 -150 12633 -92
rect 12667 -150 12725 -92
rect 12759 -150 12817 -92
rect 12851 -150 12909 -92
rect 12943 -150 13001 -92
rect 13035 -150 13093 -92
rect 13127 -150 13185 -92
rect 13219 -150 13277 -92
rect 13311 -150 13369 -92
rect 13403 -150 13461 -92
rect 13495 -150 13553 -92
rect 13587 -150 13645 -92
rect 13679 -150 13737 -92
rect 13771 -150 13829 -92
rect 13863 -150 13921 -92
rect 13955 -150 14013 -92
rect 14047 -150 14105 -92
rect 14139 -150 14197 -92
rect 14231 -150 14289 -92
rect 14323 -150 14381 -92
rect 14415 -150 14473 -92
rect 14507 -150 14565 -92
rect 14599 -150 14657 -92
rect 14691 -150 14749 -92
rect 14783 -150 14841 -92
rect 14875 -150 14933 -92
rect 14967 -150 15025 -92
rect 15059 -150 15117 -92
rect 15151 -150 15209 -92
rect 15243 -150 15301 -92
rect 15335 -150 15393 -92
rect 15427 -150 15485 -92
rect 15519 -150 15577 -92
rect 15611 -150 15669 -92
rect 15703 -150 15761 -92
rect 15795 -150 15853 -92
rect 15887 -150 15945 -92
rect 15979 -150 16037 -92
rect 16071 -150 16129 -92
rect 16163 -150 16221 -92
rect 16255 -150 16313 -92
rect 16347 -150 16405 -92
rect 16439 -150 16497 -92
rect 16531 -150 16589 -92
rect 16623 -150 16681 -92
rect 16715 -150 16744 -92
<< viali >>
rect 31 2961 65 2971
rect 31 2937 65 2961
rect 123 2961 157 2971
rect 123 2937 157 2961
rect 215 2961 249 2971
rect 215 2937 249 2961
rect 307 2961 341 2971
rect 307 2937 341 2961
rect 399 2961 433 2971
rect 399 2937 433 2961
rect 491 2961 525 2971
rect 491 2937 525 2961
rect 583 2961 617 2971
rect 583 2937 617 2961
rect 675 2961 709 2971
rect 675 2937 709 2961
rect 767 2961 801 2971
rect 767 2937 801 2961
rect 859 2961 893 2971
rect 859 2937 893 2961
rect 951 2961 985 2971
rect 951 2937 985 2961
rect 1043 2961 1077 2971
rect 1043 2937 1077 2961
rect 1135 2961 1169 2971
rect 1135 2937 1169 2961
rect 1227 2961 1261 2971
rect 1227 2937 1261 2961
rect 1319 2961 1353 2971
rect 1319 2937 1353 2961
rect 1411 2961 1445 2971
rect 1411 2937 1445 2961
rect 1503 2961 1537 2971
rect 1503 2937 1537 2961
rect 1595 2961 1629 2971
rect 1595 2937 1629 2961
rect 1687 2961 1721 2971
rect 1687 2937 1721 2961
rect 1779 2961 1813 2971
rect 1779 2937 1813 2961
rect 1871 2961 1905 2971
rect 1871 2937 1905 2961
rect 1963 2961 1997 2971
rect 1963 2937 1997 2961
rect 2055 2961 2089 2971
rect 2055 2937 2089 2961
rect 2147 2961 2181 2971
rect 2147 2937 2181 2961
rect 2239 2961 2273 2971
rect 2239 2937 2273 2961
rect 2331 2961 2365 2971
rect 2331 2937 2365 2961
rect 2423 2961 2457 2971
rect 2423 2937 2457 2961
rect 2515 2961 2549 2971
rect 2515 2937 2549 2961
rect 2607 2961 2641 2971
rect 2607 2937 2641 2961
rect 2699 2961 2733 2971
rect 2699 2937 2733 2961
rect 2791 2961 2825 2971
rect 2791 2937 2825 2961
rect 4415 2961 4449 2971
rect 4415 2937 4449 2961
rect 4507 2961 4541 2971
rect 4507 2937 4541 2961
rect 4599 2961 4633 2971
rect 4599 2937 4633 2961
rect 4691 2961 4725 2971
rect 4691 2937 4725 2961
rect 4783 2961 4817 2971
rect 4783 2937 4817 2961
rect 4875 2961 4909 2971
rect 4875 2937 4909 2961
rect 4967 2961 5001 2971
rect 4967 2937 5001 2961
rect 5059 2961 5093 2971
rect 5059 2937 5093 2961
rect 5151 2961 5185 2971
rect 5151 2937 5185 2961
rect 5243 2961 5277 2971
rect 5243 2937 5277 2961
rect 5335 2961 5369 2971
rect 5335 2937 5369 2961
rect 5427 2961 5461 2971
rect 5427 2937 5461 2961
rect 5519 2961 5553 2971
rect 5519 2937 5553 2961
rect 5611 2961 5645 2971
rect 5611 2937 5645 2961
rect 5703 2961 5737 2971
rect 5703 2937 5737 2961
rect 5795 2961 5829 2971
rect 5795 2937 5829 2961
rect 5887 2961 5921 2971
rect 5887 2937 5921 2961
rect 5979 2961 6013 2971
rect 5979 2937 6013 2961
rect 6071 2961 6105 2971
rect 6071 2937 6105 2961
rect 6163 2961 6197 2971
rect 6163 2937 6197 2961
rect 6255 2961 6289 2971
rect 6255 2937 6289 2961
rect 6347 2961 6381 2971
rect 6347 2937 6381 2961
rect 6439 2961 6473 2971
rect 6439 2937 6473 2961
rect 6531 2961 6565 2971
rect 6531 2937 6565 2961
rect 6623 2961 6657 2971
rect 6623 2937 6657 2961
rect 6715 2961 6749 2971
rect 6715 2937 6749 2961
rect 6807 2961 6841 2971
rect 6807 2937 6841 2961
rect 6899 2961 6933 2971
rect 6899 2937 6933 2961
rect 6991 2961 7025 2971
rect 6991 2937 7025 2961
rect 7083 2961 7117 2971
rect 7083 2937 7117 2961
rect 7175 2961 7209 2971
rect 7175 2937 7209 2961
rect 39 2659 73 2675
rect 39 2641 73 2659
rect 2876 2630 2910 2664
rect 4423 2625 4457 2658
rect 4423 2624 4457 2625
rect 7176 2632 7210 2666
rect 31 2403 65 2427
rect 31 2393 65 2403
rect 123 2403 157 2427
rect 123 2393 157 2403
rect 215 2403 249 2427
rect 215 2393 249 2403
rect 307 2403 341 2427
rect 307 2393 341 2403
rect 399 2403 433 2427
rect 399 2393 433 2403
rect 491 2403 525 2427
rect 491 2393 525 2403
rect 583 2403 617 2427
rect 583 2393 617 2403
rect 675 2403 709 2427
rect 675 2393 709 2403
rect 767 2403 801 2427
rect 767 2393 801 2403
rect 859 2403 893 2427
rect 859 2393 893 2403
rect 951 2403 985 2427
rect 951 2393 985 2403
rect 1043 2403 1077 2427
rect 1043 2393 1077 2403
rect 1135 2403 1169 2427
rect 1135 2393 1169 2403
rect 1227 2403 1261 2427
rect 1227 2393 1261 2403
rect 1319 2403 1353 2427
rect 1319 2393 1353 2403
rect 1411 2403 1445 2427
rect 1411 2393 1445 2403
rect 1503 2403 1537 2427
rect 1503 2393 1537 2403
rect 1595 2403 1629 2427
rect 1595 2393 1629 2403
rect 1687 2403 1721 2427
rect 1687 2393 1721 2403
rect 1779 2403 1813 2427
rect 1779 2393 1813 2403
rect 1871 2403 1905 2427
rect 1871 2393 1905 2403
rect 1963 2403 1997 2427
rect 1963 2393 1997 2403
rect 2055 2403 2089 2427
rect 2055 2393 2089 2403
rect 2147 2403 2181 2427
rect 2147 2393 2181 2403
rect 2239 2403 2273 2427
rect 2239 2393 2273 2403
rect 2331 2403 2365 2427
rect 2331 2393 2365 2403
rect 2423 2403 2457 2427
rect 2423 2393 2457 2403
rect 2515 2403 2549 2427
rect 2515 2393 2549 2403
rect 2607 2403 2641 2427
rect 2607 2393 2641 2403
rect 2699 2403 2733 2427
rect 2699 2393 2733 2403
rect 2791 2403 2825 2427
rect 2791 2393 2825 2403
rect 4415 2403 4449 2427
rect 4415 2393 4449 2403
rect 4507 2403 4541 2427
rect 4507 2393 4541 2403
rect 4599 2403 4633 2427
rect 4599 2393 4633 2403
rect 4691 2403 4725 2427
rect 4691 2393 4725 2403
rect 4783 2403 4817 2427
rect 4783 2393 4817 2403
rect 4875 2403 4909 2427
rect 4875 2393 4909 2403
rect 4967 2403 5001 2427
rect 4967 2393 5001 2403
rect 5059 2403 5093 2427
rect 5059 2393 5093 2403
rect 5151 2403 5185 2427
rect 5151 2393 5185 2403
rect 5243 2403 5277 2427
rect 5243 2393 5277 2403
rect 5335 2403 5369 2427
rect 5335 2393 5369 2403
rect 5427 2403 5461 2427
rect 5427 2393 5461 2403
rect 5519 2403 5553 2427
rect 5519 2393 5553 2403
rect 5611 2403 5645 2427
rect 5611 2393 5645 2403
rect 5703 2403 5737 2427
rect 5703 2393 5737 2403
rect 5795 2403 5829 2427
rect 5795 2393 5829 2403
rect 5887 2403 5921 2427
rect 5887 2393 5921 2403
rect 5979 2403 6013 2427
rect 5979 2393 6013 2403
rect 6071 2403 6105 2427
rect 6071 2393 6105 2403
rect 6163 2403 6197 2427
rect 6163 2393 6197 2403
rect 6255 2403 6289 2427
rect 6255 2393 6289 2403
rect 6347 2403 6381 2427
rect 6347 2393 6381 2403
rect 6439 2403 6473 2427
rect 6439 2393 6473 2403
rect 6531 2403 6565 2427
rect 6531 2393 6565 2403
rect 6623 2403 6657 2427
rect 6623 2393 6657 2403
rect 6715 2403 6749 2427
rect 6715 2393 6749 2403
rect 6807 2403 6841 2427
rect 6807 2393 6841 2403
rect 6899 2403 6933 2427
rect 6899 2393 6933 2403
rect 6991 2403 7025 2427
rect 6991 2393 7025 2403
rect 7083 2403 7117 2427
rect 7083 2393 7117 2403
rect 7175 2403 7209 2427
rect 7175 2393 7209 2403
rect 29 1819 63 1829
rect 29 1795 63 1819
rect 121 1819 155 1829
rect 121 1795 155 1819
rect 213 1819 247 1829
rect 213 1795 247 1819
rect 305 1819 339 1829
rect 305 1795 339 1819
rect 397 1819 431 1829
rect 397 1795 431 1819
rect 489 1819 523 1829
rect 489 1795 523 1819
rect 581 1819 615 1829
rect 581 1795 615 1819
rect 673 1819 707 1829
rect 673 1795 707 1819
rect 765 1819 799 1829
rect 765 1795 799 1819
rect 1463 1795 1497 1829
rect 1555 1795 1589 1829
rect 1647 1795 1681 1829
rect 1739 1795 1773 1829
rect 1831 1795 1865 1829
rect 1923 1795 1957 1829
rect 2015 1795 2049 1829
rect 2107 1795 2141 1829
rect 2199 1795 2233 1829
rect 2421 1819 2455 1829
rect 2421 1795 2455 1819
rect 2513 1819 2547 1829
rect 2513 1795 2547 1819
rect 2605 1819 2639 1829
rect 2605 1795 2639 1819
rect 2697 1819 2731 1829
rect 2697 1795 2731 1819
rect 2789 1819 2823 1829
rect 2789 1795 2823 1819
rect 2881 1819 2915 1829
rect 2881 1795 2915 1819
rect 2973 1819 3007 1829
rect 2973 1795 3007 1819
rect 3065 1819 3099 1829
rect 3065 1795 3099 1819
rect 3157 1819 3191 1829
rect 3157 1795 3191 1819
rect 3855 1795 3889 1829
rect 3947 1795 3981 1829
rect 4039 1795 4073 1829
rect 4131 1795 4165 1829
rect 4223 1795 4257 1829
rect 4315 1795 4349 1829
rect 4407 1795 4441 1829
rect 4499 1795 4533 1829
rect 4591 1795 4625 1829
rect 4813 1819 4847 1829
rect 4813 1795 4847 1819
rect 4905 1819 4939 1829
rect 4905 1795 4939 1819
rect 4997 1819 5031 1829
rect 4997 1795 5031 1819
rect 5089 1819 5123 1829
rect 5089 1795 5123 1819
rect 5181 1819 5215 1829
rect 5181 1795 5215 1819
rect 5273 1819 5307 1829
rect 5273 1795 5307 1819
rect 5365 1819 5399 1829
rect 5365 1795 5399 1819
rect 5457 1819 5491 1829
rect 5457 1795 5491 1819
rect 5549 1819 5583 1829
rect 6245 1819 6279 1829
rect 5549 1795 5583 1819
rect 6245 1795 6279 1819
rect 6337 1819 6371 1829
rect 6337 1795 6371 1819
rect 6429 1819 6463 1829
rect 6429 1795 6463 1819
rect 6521 1819 6555 1829
rect 6521 1795 6555 1819
rect 6613 1819 6647 1829
rect 6613 1795 6647 1819
rect 6705 1819 6739 1829
rect 6705 1795 6739 1819
rect 6797 1819 6831 1829
rect 6797 1795 6831 1819
rect 6889 1819 6923 1829
rect 6889 1795 6923 1819
rect 6981 1819 7015 1829
rect 6981 1795 7015 1819
rect 7205 1795 7239 1829
rect 7297 1795 7331 1829
rect 7389 1795 7423 1829
rect 7481 1795 7515 1829
rect 7573 1795 7607 1829
rect 7665 1795 7699 1829
rect 7757 1795 7791 1829
rect 7849 1795 7883 1829
rect 7941 1795 7975 1829
rect 8639 1819 8671 1829
rect 8671 1819 8673 1829
rect 8731 1819 8763 1829
rect 8763 1819 8765 1829
rect 8823 1819 8855 1829
rect 8855 1819 8857 1829
rect 8915 1819 8947 1829
rect 8947 1819 8949 1829
rect 9007 1819 9039 1829
rect 9039 1819 9041 1829
rect 9099 1819 9131 1829
rect 9131 1819 9133 1829
rect 9191 1819 9223 1829
rect 9223 1819 9225 1829
rect 9283 1819 9315 1829
rect 9315 1819 9317 1829
rect 9375 1819 9407 1829
rect 9407 1819 9409 1829
rect 8639 1795 8673 1819
rect 8731 1795 8765 1819
rect 8823 1795 8857 1819
rect 8915 1795 8949 1819
rect 9007 1795 9041 1819
rect 9099 1795 9133 1819
rect 9191 1795 9225 1819
rect 9283 1795 9317 1819
rect 9375 1795 9409 1819
rect 9597 1795 9631 1829
rect 9689 1795 9723 1829
rect 9781 1795 9815 1829
rect 9873 1795 9907 1829
rect 9965 1795 9999 1829
rect 10057 1795 10091 1829
rect 10149 1795 10183 1829
rect 10241 1795 10275 1829
rect 10333 1795 10367 1829
rect 11031 1819 11063 1829
rect 11063 1819 11065 1829
rect 11123 1819 11155 1829
rect 11155 1819 11157 1829
rect 11215 1819 11247 1829
rect 11247 1819 11249 1829
rect 11307 1819 11339 1829
rect 11339 1819 11341 1829
rect 11399 1819 11431 1829
rect 11431 1819 11433 1829
rect 11491 1819 11523 1829
rect 11523 1819 11525 1829
rect 11583 1819 11615 1829
rect 11615 1819 11617 1829
rect 11675 1819 11707 1829
rect 11707 1819 11709 1829
rect 11767 1819 11799 1829
rect 11799 1819 11801 1829
rect 11989 1819 12011 1829
rect 12011 1819 12023 1829
rect 12081 1819 12103 1829
rect 12103 1819 12115 1829
rect 12173 1819 12195 1829
rect 12195 1819 12207 1829
rect 12265 1819 12287 1829
rect 12287 1819 12299 1829
rect 12357 1819 12379 1829
rect 12379 1819 12391 1829
rect 12449 1819 12471 1829
rect 12471 1819 12483 1829
rect 12541 1819 12563 1829
rect 12563 1819 12575 1829
rect 12633 1819 12655 1829
rect 12655 1819 12667 1829
rect 12725 1819 12747 1829
rect 12747 1819 12759 1829
rect 13421 1819 13425 1829
rect 13425 1819 13455 1829
rect 13513 1819 13517 1829
rect 13517 1819 13547 1829
rect 13605 1819 13609 1829
rect 13609 1819 13639 1829
rect 13697 1819 13701 1829
rect 13701 1819 13731 1829
rect 13789 1819 13793 1829
rect 13793 1819 13823 1829
rect 13881 1819 13885 1829
rect 13885 1819 13915 1829
rect 13973 1819 13977 1829
rect 13977 1819 14007 1829
rect 14065 1819 14069 1829
rect 14069 1819 14099 1829
rect 14157 1819 14161 1829
rect 14161 1819 14191 1829
rect 14381 1819 14403 1829
rect 14403 1819 14415 1829
rect 14473 1819 14495 1829
rect 14495 1819 14507 1829
rect 14565 1819 14587 1829
rect 14587 1819 14599 1829
rect 14657 1819 14679 1829
rect 14679 1819 14691 1829
rect 14749 1819 14771 1829
rect 14771 1819 14783 1829
rect 14841 1819 14863 1829
rect 14863 1819 14875 1829
rect 14933 1819 14955 1829
rect 14955 1819 14967 1829
rect 15025 1819 15047 1829
rect 15047 1819 15059 1829
rect 15117 1819 15139 1829
rect 15139 1819 15151 1829
rect 15815 1819 15817 1829
rect 15817 1819 15849 1829
rect 15907 1819 15909 1829
rect 15909 1819 15941 1829
rect 15999 1819 16001 1829
rect 16001 1819 16033 1829
rect 16091 1819 16093 1829
rect 16093 1819 16125 1829
rect 16183 1819 16185 1829
rect 16185 1819 16217 1829
rect 16275 1819 16277 1829
rect 16277 1819 16309 1829
rect 16367 1819 16369 1829
rect 16369 1819 16401 1829
rect 16459 1819 16461 1829
rect 16461 1819 16493 1829
rect 16551 1819 16553 1829
rect 16553 1819 16585 1829
rect 11031 1795 11065 1819
rect 11123 1795 11157 1819
rect 11215 1795 11249 1819
rect 11307 1795 11341 1819
rect 11399 1795 11433 1819
rect 11491 1795 11525 1819
rect 11583 1795 11617 1819
rect 11675 1795 11709 1819
rect 11767 1795 11801 1819
rect 11989 1795 12023 1819
rect 12081 1795 12115 1819
rect 12173 1795 12207 1819
rect 12265 1795 12299 1819
rect 12357 1795 12391 1819
rect 12449 1795 12483 1819
rect 12541 1795 12575 1819
rect 12633 1795 12667 1819
rect 12725 1795 12759 1819
rect 13421 1795 13455 1819
rect 13513 1795 13547 1819
rect 13605 1795 13639 1819
rect 13697 1795 13731 1819
rect 13789 1795 13823 1819
rect 13881 1795 13915 1819
rect 13973 1795 14007 1819
rect 14065 1795 14099 1819
rect 14157 1795 14191 1819
rect 14381 1795 14415 1819
rect 14473 1795 14507 1819
rect 14565 1795 14599 1819
rect 14657 1795 14691 1819
rect 14749 1795 14783 1819
rect 14841 1795 14875 1819
rect 14933 1795 14967 1819
rect 15025 1795 15059 1819
rect 15117 1795 15151 1819
rect 15815 1795 15849 1819
rect 15907 1795 15941 1819
rect 15999 1795 16033 1819
rect 16091 1795 16125 1819
rect 16183 1795 16217 1819
rect 16275 1795 16309 1819
rect 16367 1795 16401 1819
rect 16459 1795 16493 1819
rect 16551 1795 16585 1819
rect 28 1380 62 1406
rect 484 1594 518 1607
rect 484 1573 491 1594
rect 491 1573 518 1594
rect 28 1372 35 1380
rect 35 1372 62 1380
rect 656 1560 659 1591
rect 659 1560 690 1591
rect 656 1557 690 1560
rect 1566 1560 1569 1592
rect 1569 1560 1600 1592
rect 1566 1558 1600 1560
rect 1746 1594 1780 1607
rect 1746 1573 1771 1594
rect 1771 1573 1780 1594
rect 2204 1380 2238 1404
rect 2204 1370 2227 1380
rect 2227 1370 2238 1380
rect 2420 1380 2454 1406
rect 2877 1594 2911 1606
rect 2877 1572 2883 1594
rect 2883 1572 2911 1594
rect 2420 1372 2427 1380
rect 2427 1372 2454 1380
rect 3048 1560 3051 1590
rect 3051 1560 3082 1590
rect 3048 1556 3082 1560
rect 3958 1560 3961 1591
rect 3961 1560 3992 1591
rect 3958 1557 3992 1560
rect 4138 1594 4172 1607
rect 4138 1573 4163 1594
rect 4163 1573 4172 1594
rect 4598 1380 4632 1404
rect 4598 1370 4619 1380
rect 4619 1370 4632 1380
rect 4812 1380 4846 1406
rect 5269 1594 5303 1606
rect 5269 1572 5275 1594
rect 5275 1572 5303 1594
rect 4812 1372 4819 1380
rect 4819 1372 4846 1380
rect 5439 1560 5443 1591
rect 5443 1560 5473 1591
rect 5439 1557 5473 1560
rect 6348 1560 6351 1591
rect 6351 1560 6382 1591
rect 6348 1557 6382 1560
rect 6529 1594 6563 1608
rect 6529 1574 6553 1594
rect 6553 1574 6563 1594
rect 6988 1380 7022 1406
rect 6988 1372 7009 1380
rect 7009 1372 7022 1380
rect 7204 1380 7238 1406
rect 7661 1594 7695 1607
rect 7661 1573 7667 1594
rect 7667 1573 7695 1594
rect 7204 1372 7211 1380
rect 7211 1372 7238 1380
rect 7832 1560 7835 1591
rect 7835 1560 7866 1591
rect 7832 1557 7866 1560
rect 8742 1560 8745 1592
rect 8745 1560 8776 1592
rect 8742 1558 8776 1560
rect 8922 1594 8956 1608
rect 8922 1574 8947 1594
rect 8947 1574 8956 1594
rect 9380 1380 9414 1404
rect 9380 1370 9403 1380
rect 9403 1370 9414 1380
rect 9595 1380 9629 1407
rect 10052 1594 10086 1606
rect 10052 1572 10059 1594
rect 10059 1572 10086 1594
rect 9595 1373 9603 1380
rect 9603 1373 9629 1380
rect 10223 1560 10227 1592
rect 10227 1560 10257 1592
rect 10223 1558 10257 1560
rect 11134 1560 11137 1591
rect 11137 1560 11168 1591
rect 11134 1557 11168 1560
rect 11315 1594 11349 1608
rect 11315 1574 11339 1594
rect 11339 1574 11349 1594
rect 11772 1380 11806 1406
rect 11772 1372 11795 1380
rect 11795 1372 11806 1380
rect 11987 1380 12021 1406
rect 12444 1594 12478 1605
rect 12444 1571 12451 1594
rect 12451 1571 12478 1594
rect 11987 1372 11995 1380
rect 11995 1372 12021 1380
rect 12615 1560 12619 1592
rect 12619 1560 12649 1592
rect 12615 1558 12649 1560
rect 13523 1560 13527 1591
rect 13527 1560 13557 1591
rect 13523 1557 13557 1560
rect 13704 1594 13738 1608
rect 13704 1574 13729 1594
rect 13729 1574 13738 1594
rect 14164 1380 14198 1404
rect 14164 1370 14185 1380
rect 14185 1370 14198 1380
rect 14380 1380 14414 1407
rect 14836 1594 14870 1606
rect 14836 1572 14843 1594
rect 14843 1572 14870 1594
rect 14380 1373 14387 1380
rect 14387 1373 14414 1380
rect 15008 1560 15011 1592
rect 15011 1560 15042 1592
rect 15008 1558 15042 1560
rect 15918 1560 15921 1592
rect 15921 1560 15952 1592
rect 15918 1558 15952 1560
rect 16099 1594 16133 1608
rect 16099 1574 16123 1594
rect 16123 1574 16133 1594
rect 16556 1380 16590 1406
rect 16556 1372 16579 1380
rect 16579 1372 16590 1380
rect 29 1261 63 1285
rect 29 1251 63 1261
rect 121 1261 155 1285
rect 121 1251 155 1261
rect 213 1261 247 1285
rect 213 1251 247 1261
rect 305 1261 339 1285
rect 305 1251 339 1261
rect 397 1261 431 1285
rect 397 1251 431 1261
rect 489 1261 523 1285
rect 489 1251 523 1261
rect 581 1261 615 1285
rect 581 1251 615 1261
rect 673 1261 707 1285
rect 673 1251 707 1261
rect 765 1261 799 1285
rect 765 1251 799 1261
rect 1463 1251 1497 1285
rect 1555 1251 1589 1285
rect 1647 1251 1681 1285
rect 1739 1251 1773 1285
rect 1831 1251 1865 1285
rect 1923 1251 1957 1285
rect 2015 1251 2049 1285
rect 2107 1251 2141 1285
rect 2199 1251 2233 1285
rect 2421 1261 2455 1285
rect 2421 1251 2455 1261
rect 2513 1261 2547 1285
rect 2513 1251 2547 1261
rect 2605 1261 2639 1285
rect 2605 1251 2639 1261
rect 2697 1261 2731 1285
rect 2697 1251 2731 1261
rect 2789 1261 2823 1285
rect 2789 1251 2823 1261
rect 2881 1261 2915 1285
rect 2881 1251 2915 1261
rect 2973 1261 3007 1285
rect 2973 1251 3007 1261
rect 3065 1261 3099 1285
rect 3065 1251 3099 1261
rect 3157 1261 3191 1285
rect 3157 1251 3191 1261
rect 3855 1251 3889 1285
rect 3947 1251 3981 1285
rect 4039 1251 4073 1285
rect 4131 1251 4165 1285
rect 4223 1251 4257 1285
rect 4315 1251 4349 1285
rect 4407 1251 4441 1285
rect 4499 1251 4533 1285
rect 4591 1251 4625 1285
rect 4813 1261 4847 1285
rect 4813 1251 4847 1261
rect 4905 1261 4939 1285
rect 4905 1251 4939 1261
rect 4997 1261 5031 1285
rect 4997 1251 5031 1261
rect 5089 1261 5123 1285
rect 5089 1251 5123 1261
rect 5181 1261 5215 1285
rect 5181 1251 5215 1261
rect 5273 1261 5307 1285
rect 5273 1251 5307 1261
rect 5365 1261 5399 1285
rect 5365 1251 5399 1261
rect 5457 1261 5491 1285
rect 5457 1251 5491 1261
rect 5549 1261 5583 1285
rect 6245 1261 6279 1285
rect 5549 1251 5583 1261
rect 6245 1251 6279 1261
rect 6337 1261 6371 1285
rect 6337 1251 6371 1261
rect 6429 1261 6463 1285
rect 6429 1251 6463 1261
rect 6521 1261 6555 1285
rect 6521 1251 6555 1261
rect 6613 1261 6647 1285
rect 6613 1251 6647 1261
rect 6705 1261 6739 1285
rect 6705 1251 6739 1261
rect 6797 1261 6831 1285
rect 6797 1251 6831 1261
rect 6889 1261 6923 1285
rect 6889 1251 6923 1261
rect 6981 1261 7015 1285
rect 6981 1251 7015 1261
rect 7205 1251 7239 1285
rect 7297 1251 7331 1285
rect 7389 1251 7423 1285
rect 7481 1251 7515 1285
rect 7573 1251 7607 1285
rect 7665 1251 7699 1285
rect 7757 1251 7791 1285
rect 7849 1251 7883 1285
rect 7941 1251 7975 1285
rect 8639 1261 8673 1285
rect 8731 1261 8765 1285
rect 8823 1261 8857 1285
rect 8915 1261 8949 1285
rect 9007 1261 9041 1285
rect 9099 1261 9133 1285
rect 9191 1261 9225 1285
rect 9283 1261 9317 1285
rect 9375 1261 9409 1285
rect 8639 1251 8671 1261
rect 8671 1251 8673 1261
rect 8731 1251 8763 1261
rect 8763 1251 8765 1261
rect 8823 1251 8855 1261
rect 8855 1251 8857 1261
rect 8915 1251 8947 1261
rect 8947 1251 8949 1261
rect 9007 1251 9039 1261
rect 9039 1251 9041 1261
rect 9099 1251 9131 1261
rect 9131 1251 9133 1261
rect 9191 1251 9223 1261
rect 9223 1251 9225 1261
rect 9283 1251 9315 1261
rect 9315 1251 9317 1261
rect 9375 1251 9407 1261
rect 9407 1251 9409 1261
rect 9597 1251 9631 1285
rect 9689 1251 9723 1285
rect 9781 1251 9815 1285
rect 9873 1251 9907 1285
rect 9965 1251 9999 1285
rect 10057 1251 10091 1285
rect 10149 1251 10183 1285
rect 10241 1251 10275 1285
rect 10333 1251 10367 1285
rect 11031 1261 11065 1285
rect 11123 1261 11157 1285
rect 11215 1261 11249 1285
rect 11307 1261 11341 1285
rect 11399 1261 11433 1285
rect 11491 1261 11525 1285
rect 11583 1261 11617 1285
rect 11675 1261 11709 1285
rect 11767 1261 11801 1285
rect 11989 1261 12023 1285
rect 12081 1261 12115 1285
rect 12173 1261 12207 1285
rect 12265 1261 12299 1285
rect 12357 1261 12391 1285
rect 12449 1261 12483 1285
rect 12541 1261 12575 1285
rect 12633 1261 12667 1285
rect 12725 1261 12759 1285
rect 13421 1261 13455 1285
rect 13513 1261 13547 1285
rect 13605 1261 13639 1285
rect 13697 1261 13731 1285
rect 13789 1261 13823 1285
rect 13881 1261 13915 1285
rect 13973 1261 14007 1285
rect 14065 1261 14099 1285
rect 14157 1261 14191 1285
rect 14381 1261 14415 1285
rect 14473 1261 14507 1285
rect 14565 1261 14599 1285
rect 14657 1261 14691 1285
rect 14749 1261 14783 1285
rect 14841 1261 14875 1285
rect 14933 1261 14967 1285
rect 15025 1261 15059 1285
rect 15117 1261 15151 1285
rect 15815 1261 15849 1285
rect 15907 1261 15941 1285
rect 15999 1261 16033 1285
rect 16091 1261 16125 1285
rect 16183 1261 16217 1285
rect 16275 1261 16309 1285
rect 16367 1261 16401 1285
rect 16459 1261 16493 1285
rect 16551 1261 16585 1285
rect 11031 1251 11063 1261
rect 11063 1251 11065 1261
rect 11123 1251 11155 1261
rect 11155 1251 11157 1261
rect 11215 1251 11247 1261
rect 11247 1251 11249 1261
rect 11307 1251 11339 1261
rect 11339 1251 11341 1261
rect 11399 1251 11431 1261
rect 11431 1251 11433 1261
rect 11491 1251 11523 1261
rect 11523 1251 11525 1261
rect 11583 1251 11615 1261
rect 11615 1251 11617 1261
rect 11675 1251 11707 1261
rect 11707 1251 11709 1261
rect 11767 1251 11799 1261
rect 11799 1251 11801 1261
rect 11989 1251 12011 1261
rect 12011 1251 12023 1261
rect 12081 1251 12103 1261
rect 12103 1251 12115 1261
rect 12173 1251 12195 1261
rect 12195 1251 12207 1261
rect 12265 1251 12287 1261
rect 12287 1251 12299 1261
rect 12357 1251 12379 1261
rect 12379 1251 12391 1261
rect 12449 1251 12471 1261
rect 12471 1251 12483 1261
rect 12541 1251 12563 1261
rect 12563 1251 12575 1261
rect 12633 1251 12655 1261
rect 12655 1251 12667 1261
rect 12725 1251 12747 1261
rect 12747 1251 12759 1261
rect 13421 1251 13425 1261
rect 13425 1251 13455 1261
rect 13513 1251 13517 1261
rect 13517 1251 13547 1261
rect 13605 1251 13609 1261
rect 13609 1251 13639 1261
rect 13697 1251 13701 1261
rect 13701 1251 13731 1261
rect 13789 1251 13793 1261
rect 13793 1251 13823 1261
rect 13881 1251 13885 1261
rect 13885 1251 13915 1261
rect 13973 1251 13977 1261
rect 13977 1251 14007 1261
rect 14065 1251 14069 1261
rect 14069 1251 14099 1261
rect 14157 1251 14161 1261
rect 14161 1251 14191 1261
rect 14381 1251 14403 1261
rect 14403 1251 14415 1261
rect 14473 1251 14495 1261
rect 14495 1251 14507 1261
rect 14565 1251 14587 1261
rect 14587 1251 14599 1261
rect 14657 1251 14679 1261
rect 14679 1251 14691 1261
rect 14749 1251 14771 1261
rect 14771 1251 14783 1261
rect 14841 1251 14863 1261
rect 14863 1251 14875 1261
rect 14933 1251 14955 1261
rect 14955 1251 14967 1261
rect 15025 1251 15047 1261
rect 15047 1251 15059 1261
rect 15117 1251 15139 1261
rect 15139 1251 15151 1261
rect 15815 1251 15817 1261
rect 15817 1251 15849 1261
rect 15907 1251 15909 1261
rect 15909 1251 15941 1261
rect 15999 1251 16001 1261
rect 16001 1251 16033 1261
rect 16091 1251 16093 1261
rect 16093 1251 16125 1261
rect 16183 1251 16185 1261
rect 16185 1251 16217 1261
rect 16275 1251 16277 1261
rect 16277 1251 16309 1261
rect 16367 1251 16369 1261
rect 16369 1251 16401 1261
rect 16459 1251 16461 1261
rect 16461 1251 16493 1261
rect 16551 1251 16553 1261
rect 16553 1251 16585 1261
rect 29 1131 63 1141
rect 29 1107 63 1131
rect 121 1131 155 1141
rect 121 1107 155 1131
rect 213 1131 247 1141
rect 213 1107 247 1131
rect 305 1131 339 1141
rect 305 1107 339 1131
rect 397 1131 431 1141
rect 397 1107 431 1131
rect 489 1131 523 1141
rect 489 1107 523 1131
rect 581 1131 615 1141
rect 581 1107 615 1131
rect 673 1131 707 1141
rect 673 1107 707 1131
rect 765 1131 799 1141
rect 765 1107 799 1131
rect 857 1131 891 1141
rect 857 1107 891 1131
rect 949 1131 983 1141
rect 949 1107 983 1131
rect 1041 1131 1075 1141
rect 1041 1107 1075 1131
rect 1133 1131 1167 1141
rect 1133 1107 1167 1131
rect 1225 1131 1259 1141
rect 1225 1107 1259 1131
rect 1317 1131 1351 1141
rect 1317 1107 1351 1131
rect 1409 1131 1443 1141
rect 1409 1107 1443 1131
rect 1501 1131 1535 1141
rect 1501 1107 1535 1131
rect 1593 1131 1627 1141
rect 1593 1107 1627 1131
rect 1685 1131 1719 1141
rect 1685 1107 1719 1131
rect 1777 1131 1811 1141
rect 1777 1107 1811 1131
rect 1869 1124 1901 1141
rect 1901 1124 1903 1141
rect 1869 1107 1903 1124
rect 1961 1107 1995 1141
rect 2053 1131 2087 1141
rect 2053 1107 2087 1131
rect 2145 1131 2179 1141
rect 2145 1107 2179 1131
rect 2237 1131 2271 1141
rect 2237 1107 2271 1131
rect 2329 1131 2363 1141
rect 2329 1107 2363 1131
rect 2421 1131 2455 1141
rect 2421 1107 2455 1131
rect 2513 1131 2547 1141
rect 2513 1107 2547 1131
rect 2605 1131 2639 1141
rect 2605 1107 2639 1131
rect 2697 1131 2731 1141
rect 2697 1107 2731 1131
rect 2789 1131 2823 1141
rect 2789 1107 2823 1131
rect 2881 1131 2915 1141
rect 2881 1107 2915 1131
rect 2973 1131 3007 1141
rect 2973 1107 3007 1131
rect 3065 1131 3099 1141
rect 3065 1107 3099 1131
rect 3157 1131 3191 1141
rect 3157 1107 3191 1131
rect 3249 1131 3283 1141
rect 3249 1107 3283 1131
rect 3341 1131 3375 1141
rect 3341 1107 3375 1131
rect 3433 1131 3467 1141
rect 3433 1107 3467 1131
rect 3525 1131 3559 1141
rect 3525 1107 3559 1131
rect 3617 1131 3651 1141
rect 3617 1107 3651 1131
rect 3709 1131 3743 1141
rect 3709 1107 3743 1131
rect 3801 1131 3835 1141
rect 3801 1107 3835 1131
rect 3893 1131 3927 1141
rect 3893 1107 3927 1131
rect 3985 1131 4019 1141
rect 3985 1107 4019 1131
rect 4077 1131 4111 1141
rect 4077 1107 4111 1131
rect 4169 1131 4203 1141
rect 4169 1107 4203 1131
rect 4261 1123 4293 1141
rect 4293 1123 4295 1141
rect 4261 1107 4295 1123
rect 4353 1107 4387 1141
rect 4445 1131 4479 1141
rect 4445 1107 4479 1131
rect 4537 1131 4571 1141
rect 4537 1107 4571 1131
rect 4629 1131 4663 1141
rect 4629 1107 4663 1131
rect 4721 1131 4755 1141
rect 4721 1107 4755 1131
rect 4813 1131 4847 1141
rect 4813 1107 4847 1131
rect 4905 1131 4939 1141
rect 4905 1107 4939 1131
rect 4997 1131 5031 1141
rect 4997 1107 5031 1131
rect 5089 1131 5123 1141
rect 5089 1107 5123 1131
rect 5181 1131 5215 1141
rect 5181 1107 5215 1131
rect 5273 1131 5307 1141
rect 5273 1107 5307 1131
rect 5365 1131 5399 1141
rect 5365 1107 5399 1131
rect 5457 1131 5491 1141
rect 5457 1107 5491 1131
rect 5549 1131 5583 1141
rect 5549 1107 5583 1131
rect 5641 1131 5675 1141
rect 5641 1107 5675 1131
rect 5733 1131 5767 1141
rect 5733 1107 5767 1131
rect 5825 1131 5859 1141
rect 5825 1107 5859 1131
rect 5917 1131 5951 1141
rect 5917 1107 5951 1131
rect 6009 1131 6043 1141
rect 6009 1107 6043 1131
rect 6101 1131 6135 1141
rect 6101 1107 6135 1131
rect 6193 1131 6227 1141
rect 6193 1107 6227 1131
rect 6285 1131 6319 1141
rect 6285 1107 6319 1131
rect 6377 1131 6411 1141
rect 6377 1107 6411 1131
rect 6469 1131 6503 1141
rect 6469 1107 6503 1131
rect 6561 1131 6595 1141
rect 6561 1107 6595 1131
rect 6653 1123 6685 1141
rect 6685 1123 6687 1141
rect 6653 1107 6687 1123
rect 6745 1107 6779 1141
rect 6837 1131 6871 1141
rect 6837 1107 6871 1131
rect 6929 1131 6963 1141
rect 6929 1107 6963 1131
rect 7021 1131 7055 1141
rect 7021 1107 7055 1131
rect 7113 1131 7147 1141
rect 7113 1107 7147 1131
rect 7205 1131 7239 1141
rect 7205 1107 7239 1131
rect 7297 1131 7331 1141
rect 7297 1107 7331 1131
rect 7389 1131 7423 1141
rect 7389 1107 7423 1131
rect 7481 1131 7515 1141
rect 7481 1107 7515 1131
rect 7573 1131 7607 1141
rect 7573 1107 7607 1131
rect 7665 1131 7699 1141
rect 7665 1107 7699 1131
rect 7757 1131 7791 1141
rect 7757 1107 7791 1131
rect 7849 1131 7883 1141
rect 7849 1107 7883 1131
rect 7941 1131 7975 1141
rect 7941 1107 7975 1131
rect 8033 1131 8067 1141
rect 8033 1107 8067 1131
rect 8125 1131 8159 1141
rect 8125 1107 8159 1131
rect 8217 1131 8251 1141
rect 8217 1107 8251 1131
rect 8309 1131 8343 1141
rect 8309 1107 8343 1131
rect 8401 1131 8435 1141
rect 8401 1107 8435 1131
rect 8493 1131 8527 1141
rect 8493 1107 8527 1131
rect 8585 1131 8619 1141
rect 8585 1107 8619 1131
rect 8677 1131 8711 1141
rect 8677 1107 8711 1131
rect 8769 1131 8803 1141
rect 8769 1107 8803 1131
rect 8861 1131 8895 1141
rect 8861 1107 8895 1131
rect 8953 1131 8987 1141
rect 8953 1107 8987 1131
rect 9045 1124 9077 1141
rect 9077 1124 9079 1141
rect 9045 1107 9079 1124
rect 9137 1107 9171 1141
rect 9229 1131 9263 1141
rect 9229 1107 9263 1131
rect 9321 1131 9355 1141
rect 9321 1107 9355 1131
rect 9413 1131 9447 1141
rect 9413 1107 9447 1131
rect 9505 1131 9539 1141
rect 9505 1107 9539 1131
rect 9597 1131 9631 1141
rect 9597 1107 9631 1131
rect 9689 1131 9723 1141
rect 9689 1107 9723 1131
rect 9781 1131 9815 1141
rect 9781 1107 9815 1131
rect 9873 1131 9907 1141
rect 9873 1107 9907 1131
rect 9965 1131 9999 1141
rect 9965 1107 9999 1131
rect 10057 1131 10091 1141
rect 10057 1107 10091 1131
rect 10149 1131 10183 1141
rect 10149 1107 10183 1131
rect 10241 1131 10275 1141
rect 10241 1107 10275 1131
rect 10333 1131 10367 1141
rect 10333 1107 10367 1131
rect 10425 1131 10459 1141
rect 10425 1107 10459 1131
rect 10517 1131 10551 1141
rect 10517 1107 10551 1131
rect 10609 1131 10643 1141
rect 10609 1107 10643 1131
rect 10701 1131 10735 1141
rect 10701 1107 10735 1131
rect 10793 1131 10827 1141
rect 10793 1107 10827 1131
rect 10885 1131 10919 1141
rect 10885 1107 10919 1131
rect 10977 1131 11011 1141
rect 10977 1107 11011 1131
rect 11069 1131 11103 1141
rect 11069 1107 11103 1131
rect 11161 1131 11195 1141
rect 11161 1107 11195 1131
rect 11253 1131 11287 1141
rect 11253 1107 11287 1131
rect 11345 1131 11379 1141
rect 11345 1107 11379 1131
rect 11437 1124 11469 1141
rect 11469 1124 11471 1141
rect 11437 1107 11471 1124
rect 11529 1107 11563 1141
rect 11621 1131 11655 1141
rect 11621 1107 11655 1131
rect 11713 1131 11747 1141
rect 11713 1107 11747 1131
rect 11805 1131 11839 1141
rect 11805 1107 11839 1131
rect 11897 1131 11931 1141
rect 11897 1107 11931 1131
rect 11989 1131 12023 1141
rect 11989 1107 12023 1131
rect 12081 1131 12115 1141
rect 12081 1107 12115 1131
rect 12173 1131 12207 1141
rect 12173 1107 12207 1131
rect 12265 1131 12299 1141
rect 12265 1107 12299 1131
rect 12357 1131 12391 1141
rect 12357 1107 12391 1131
rect 12449 1131 12483 1141
rect 12449 1107 12483 1131
rect 12541 1131 12575 1141
rect 12541 1107 12575 1131
rect 12633 1131 12667 1141
rect 12633 1107 12667 1131
rect 12725 1131 12759 1141
rect 12725 1107 12759 1131
rect 12817 1131 12851 1141
rect 12817 1107 12851 1131
rect 12909 1131 12943 1141
rect 12909 1107 12943 1131
rect 13001 1131 13035 1141
rect 13001 1107 13035 1131
rect 13093 1131 13127 1141
rect 13093 1107 13127 1131
rect 13185 1131 13219 1141
rect 13185 1107 13219 1131
rect 13277 1131 13311 1141
rect 13277 1107 13311 1131
rect 13369 1131 13403 1141
rect 13369 1107 13403 1131
rect 13461 1131 13495 1141
rect 13461 1107 13495 1131
rect 13553 1131 13587 1141
rect 13553 1107 13587 1131
rect 13645 1131 13679 1141
rect 13645 1107 13679 1131
rect 13737 1131 13771 1141
rect 13737 1107 13771 1131
rect 13829 1123 13861 1141
rect 13861 1123 13863 1141
rect 13829 1107 13863 1123
rect 13921 1107 13955 1141
rect 14013 1131 14047 1141
rect 14013 1107 14047 1131
rect 14105 1131 14139 1141
rect 14105 1107 14139 1131
rect 14197 1131 14231 1141
rect 14197 1107 14231 1131
rect 14289 1131 14323 1141
rect 14289 1107 14323 1131
rect 14381 1131 14415 1141
rect 14381 1107 14415 1131
rect 14473 1131 14507 1141
rect 14473 1107 14507 1131
rect 14565 1131 14599 1141
rect 14565 1107 14599 1131
rect 14657 1131 14691 1141
rect 14657 1107 14691 1131
rect 14749 1131 14783 1141
rect 14749 1107 14783 1131
rect 14841 1131 14875 1141
rect 14841 1107 14875 1131
rect 14933 1131 14967 1141
rect 14933 1107 14967 1131
rect 15025 1131 15059 1141
rect 15025 1107 15059 1131
rect 15117 1131 15151 1141
rect 15117 1107 15151 1131
rect 15209 1131 15243 1141
rect 15209 1107 15243 1131
rect 15301 1131 15335 1141
rect 15301 1107 15335 1131
rect 15393 1131 15427 1141
rect 15393 1107 15427 1131
rect 15485 1131 15519 1141
rect 15485 1107 15519 1131
rect 15577 1131 15611 1141
rect 15577 1107 15611 1131
rect 15669 1131 15703 1141
rect 15669 1107 15703 1131
rect 15761 1131 15795 1141
rect 15761 1107 15795 1131
rect 15853 1131 15887 1141
rect 15853 1107 15887 1131
rect 15945 1131 15979 1141
rect 15945 1107 15979 1131
rect 16037 1131 16071 1141
rect 16037 1107 16071 1131
rect 16129 1131 16163 1141
rect 16129 1107 16163 1131
rect 16221 1123 16253 1141
rect 16253 1123 16255 1141
rect 16221 1107 16255 1123
rect 16313 1107 16347 1141
rect 16405 1131 16439 1141
rect 16405 1107 16439 1131
rect 16497 1131 16531 1141
rect 16497 1107 16531 1131
rect 16589 1131 16623 1141
rect 16589 1107 16623 1131
rect 16681 1131 16715 1141
rect 16681 1107 16715 1131
rect 26 844 60 859
rect 26 825 31 844
rect 31 825 60 844
rect 122 733 156 767
rect 213 955 237 971
rect 237 955 247 971
rect 213 937 247 955
rect 489 937 523 971
rect 366 849 400 883
rect 581 749 595 767
rect 595 749 615 767
rect 581 733 615 749
rect 1225 945 1259 971
rect 1225 937 1246 945
rect 1246 937 1259 945
rect 1133 869 1167 903
rect 765 759 767 767
rect 767 759 799 767
rect 765 733 799 759
rect 1225 801 1259 835
rect 1515 759 1545 767
rect 1545 759 1549 767
rect 1515 733 1549 759
rect 1771 869 1805 903
rect 2051 926 2074 955
rect 2074 926 2085 955
rect 2051 921 2085 926
rect 2334 1029 2368 1034
rect 2334 1000 2357 1029
rect 2357 1000 2368 1029
rect 2418 844 2452 859
rect 2418 825 2423 844
rect 2423 825 2452 844
rect 2514 733 2548 767
rect 2605 955 2629 971
rect 2629 955 2639 971
rect 2605 937 2639 955
rect 2881 937 2915 971
rect 2758 849 2792 883
rect 2973 749 2987 767
rect 2987 749 3007 767
rect 2973 733 3007 749
rect 3617 945 3651 971
rect 3617 937 3638 945
rect 3638 937 3651 945
rect 3525 869 3559 903
rect 3157 759 3159 767
rect 3159 759 3191 767
rect 3157 733 3191 759
rect 3617 801 3651 835
rect 3907 759 3937 767
rect 3937 759 3941 767
rect 3907 733 3941 759
rect 4163 869 4197 903
rect 4443 926 4466 956
rect 4466 926 4477 956
rect 4443 922 4477 926
rect 4726 1029 4760 1034
rect 4726 1000 4749 1029
rect 4749 1000 4760 1029
rect 4810 844 4844 859
rect 4810 825 4815 844
rect 4815 825 4844 844
rect 4906 733 4940 767
rect 4997 955 5021 971
rect 5021 955 5031 971
rect 4997 937 5031 955
rect 5273 937 5307 971
rect 5150 850 5184 884
rect 5365 749 5379 767
rect 5379 749 5399 767
rect 5365 733 5399 749
rect 6009 945 6043 971
rect 6009 937 6030 945
rect 6030 937 6043 945
rect 5917 869 5951 903
rect 5549 759 5551 767
rect 5551 759 5583 767
rect 5549 733 5583 759
rect 6009 801 6043 835
rect 6299 759 6329 767
rect 6329 759 6333 767
rect 6299 733 6333 759
rect 6555 869 6589 903
rect 6834 926 6858 956
rect 6858 926 6868 956
rect 6834 922 6868 926
rect 7118 1029 7152 1034
rect 7118 1000 7141 1029
rect 7141 1000 7152 1029
rect 7202 844 7236 859
rect 7202 825 7207 844
rect 7207 825 7236 844
rect 7298 733 7332 767
rect 7389 955 7413 971
rect 7413 955 7423 971
rect 7389 937 7423 955
rect 7665 937 7699 971
rect 7542 850 7576 884
rect 7757 749 7771 767
rect 7771 749 7791 767
rect 7757 733 7791 749
rect 8401 945 8435 971
rect 8401 937 8422 945
rect 8422 937 8435 945
rect 8309 869 8343 903
rect 7941 759 7943 767
rect 7943 759 7975 767
rect 7941 733 7975 759
rect 8401 801 8435 835
rect 8691 759 8721 767
rect 8721 759 8725 767
rect 8691 733 8725 759
rect 8947 869 8981 903
rect 9227 926 9250 957
rect 9250 926 9261 957
rect 9227 923 9261 926
rect 9510 1029 9544 1034
rect 9510 1000 9533 1029
rect 9533 1000 9544 1029
rect 9593 844 9627 860
rect 9593 826 9599 844
rect 9599 826 9627 844
rect 9690 733 9724 767
rect 9781 955 9805 971
rect 9805 955 9815 971
rect 9781 937 9815 955
rect 10057 937 10091 971
rect 9934 849 9968 883
rect 10149 749 10163 767
rect 10163 749 10183 767
rect 10149 733 10183 749
rect 10793 945 10827 971
rect 10793 937 10814 945
rect 10814 937 10827 945
rect 10701 869 10735 903
rect 10333 759 10335 767
rect 10335 759 10367 767
rect 10333 733 10367 759
rect 10793 801 10827 835
rect 11083 759 11113 767
rect 11113 759 11117 767
rect 11083 733 11117 759
rect 11339 869 11373 903
rect 11618 926 11642 956
rect 11642 926 11652 956
rect 11618 922 11652 926
rect 11902 1029 11936 1034
rect 11902 1000 11925 1029
rect 11925 1000 11936 1029
rect 11985 844 12019 859
rect 11985 825 11991 844
rect 11991 825 12019 844
rect 12082 733 12116 767
rect 12173 955 12197 971
rect 12197 955 12207 971
rect 12173 937 12207 955
rect 12449 937 12483 971
rect 12326 850 12360 884
rect 12541 749 12555 767
rect 12555 749 12575 767
rect 12541 733 12575 749
rect 13185 945 13219 971
rect 13185 937 13206 945
rect 13206 937 13219 945
rect 13093 869 13127 903
rect 12725 759 12727 767
rect 12727 759 12759 767
rect 12725 733 12759 759
rect 13185 801 13219 835
rect 13475 759 13505 767
rect 13505 759 13509 767
rect 13475 733 13509 759
rect 13731 869 13765 903
rect 14011 926 14034 955
rect 14034 926 14045 955
rect 14011 921 14045 926
rect 14294 1029 14328 1034
rect 14294 1000 14317 1029
rect 14317 1000 14328 1029
rect 14378 844 14412 860
rect 14378 826 14383 844
rect 14383 826 14412 844
rect 14474 733 14508 767
rect 14565 955 14589 971
rect 14589 955 14599 971
rect 14565 937 14599 955
rect 14841 937 14875 971
rect 14719 849 14753 883
rect 14933 749 14947 767
rect 14947 749 14967 767
rect 14933 733 14967 749
rect 15577 945 15611 971
rect 15577 937 15598 945
rect 15598 937 15611 945
rect 15485 869 15519 903
rect 15117 759 15119 767
rect 15119 759 15151 767
rect 15117 733 15151 759
rect 15577 801 15611 835
rect 15867 759 15897 767
rect 15897 759 15901 767
rect 15867 733 15901 759
rect 16123 869 16157 903
rect 16404 926 16426 957
rect 16426 926 16438 957
rect 16404 923 16438 926
rect 16686 1029 16720 1034
rect 16686 1000 16709 1029
rect 16709 1000 16720 1029
rect 29 573 63 597
rect 29 563 63 573
rect 121 573 155 597
rect 121 563 155 573
rect 213 573 247 597
rect 213 563 247 573
rect 305 573 339 597
rect 305 563 339 573
rect 397 573 431 597
rect 397 563 431 573
rect 489 573 523 597
rect 489 563 523 573
rect 581 573 615 597
rect 581 563 615 573
rect 673 573 707 597
rect 673 563 707 573
rect 765 573 799 597
rect 765 563 799 573
rect 857 573 891 597
rect 857 563 891 573
rect 949 573 983 597
rect 949 563 983 573
rect 1041 573 1075 597
rect 1041 563 1075 573
rect 1133 573 1167 597
rect 1133 563 1167 573
rect 1225 573 1259 597
rect 1225 563 1259 573
rect 1317 573 1351 597
rect 1317 563 1351 573
rect 1409 573 1443 597
rect 1409 563 1443 573
rect 1501 573 1535 597
rect 1501 563 1535 573
rect 1593 573 1627 597
rect 1593 563 1627 573
rect 1685 573 1719 597
rect 1685 563 1719 573
rect 1777 573 1811 597
rect 1777 563 1811 573
rect 1869 573 1903 597
rect 1869 563 1903 573
rect 1961 573 1995 597
rect 1961 563 1995 573
rect 2053 573 2087 597
rect 2053 563 2087 573
rect 2145 573 2179 597
rect 2145 563 2179 573
rect 2237 573 2271 597
rect 2237 563 2271 573
rect 2329 573 2363 597
rect 2329 563 2363 573
rect 2421 573 2455 597
rect 2421 563 2455 573
rect 2513 573 2547 597
rect 2513 563 2547 573
rect 2605 573 2639 597
rect 2605 563 2639 573
rect 2697 573 2731 597
rect 2697 563 2731 573
rect 2789 573 2823 597
rect 2789 563 2823 573
rect 2881 573 2915 597
rect 2881 563 2915 573
rect 2973 573 3007 597
rect 2973 563 3007 573
rect 3065 573 3099 597
rect 3065 563 3099 573
rect 3157 573 3191 597
rect 3157 563 3191 573
rect 3249 573 3283 597
rect 3249 563 3283 573
rect 3341 573 3375 597
rect 3341 563 3375 573
rect 3433 573 3467 597
rect 3433 563 3467 573
rect 3525 573 3559 597
rect 3525 563 3559 573
rect 3617 573 3651 597
rect 3617 563 3651 573
rect 3709 573 3743 597
rect 3709 563 3743 573
rect 3801 573 3835 597
rect 3801 563 3835 573
rect 3893 573 3927 597
rect 3893 563 3927 573
rect 3985 573 4019 597
rect 3985 563 4019 573
rect 4077 573 4111 597
rect 4077 563 4111 573
rect 4169 573 4203 597
rect 4169 563 4203 573
rect 4261 573 4295 597
rect 4261 563 4295 573
rect 4353 573 4387 597
rect 4353 563 4387 573
rect 4445 573 4479 597
rect 4445 563 4479 573
rect 4537 573 4571 597
rect 4537 563 4571 573
rect 4629 573 4663 597
rect 4629 563 4663 573
rect 4721 573 4755 597
rect 4721 563 4755 573
rect 4813 573 4847 597
rect 4813 563 4847 573
rect 4905 573 4939 597
rect 4905 563 4939 573
rect 4997 573 5031 597
rect 4997 563 5031 573
rect 5089 573 5123 597
rect 5089 563 5123 573
rect 5181 573 5215 597
rect 5181 563 5215 573
rect 5273 573 5307 597
rect 5273 563 5307 573
rect 5365 573 5399 597
rect 5365 563 5399 573
rect 5457 573 5491 597
rect 5457 563 5491 573
rect 5549 573 5583 597
rect 5549 563 5583 573
rect 5641 573 5675 597
rect 5641 563 5675 573
rect 5733 573 5767 597
rect 5733 563 5767 573
rect 5825 573 5859 597
rect 5825 563 5859 573
rect 5917 573 5951 597
rect 5917 563 5951 573
rect 6009 573 6043 597
rect 6009 563 6043 573
rect 6101 573 6135 597
rect 6101 563 6135 573
rect 6193 573 6227 597
rect 6193 563 6227 573
rect 6285 573 6319 597
rect 6285 563 6319 573
rect 6377 573 6411 597
rect 6377 563 6411 573
rect 6469 573 6503 597
rect 6469 563 6503 573
rect 6561 573 6595 597
rect 6561 563 6595 573
rect 6653 573 6687 597
rect 6653 563 6687 573
rect 6745 573 6779 597
rect 6745 563 6779 573
rect 6837 573 6871 597
rect 6837 563 6871 573
rect 6929 573 6963 597
rect 6929 563 6963 573
rect 7021 573 7055 597
rect 7021 563 7055 573
rect 7113 573 7147 597
rect 7113 563 7147 573
rect 7205 573 7239 597
rect 7205 563 7239 573
rect 7297 573 7331 597
rect 7297 563 7331 573
rect 7389 573 7423 597
rect 7389 563 7423 573
rect 7481 573 7515 597
rect 7481 563 7515 573
rect 7573 573 7607 597
rect 7573 563 7607 573
rect 7665 573 7699 597
rect 7665 563 7699 573
rect 7757 573 7791 597
rect 7757 563 7791 573
rect 7849 573 7883 597
rect 7849 563 7883 573
rect 7941 573 7975 597
rect 7941 563 7975 573
rect 8033 573 8067 597
rect 8033 563 8067 573
rect 8125 573 8159 597
rect 8125 563 8159 573
rect 8217 573 8251 597
rect 8217 563 8251 573
rect 8309 573 8343 597
rect 8309 563 8343 573
rect 8401 573 8435 597
rect 8401 563 8435 573
rect 8493 573 8527 597
rect 8493 563 8527 573
rect 8585 573 8619 597
rect 8585 563 8619 573
rect 8677 573 8711 597
rect 8677 563 8711 573
rect 8769 573 8803 597
rect 8769 563 8803 573
rect 8861 573 8895 597
rect 8861 563 8895 573
rect 8953 573 8987 597
rect 8953 563 8987 573
rect 9045 573 9079 597
rect 9045 563 9079 573
rect 9137 573 9171 597
rect 9137 563 9171 573
rect 9229 573 9263 597
rect 9229 563 9263 573
rect 9321 573 9355 597
rect 9321 563 9355 573
rect 9413 573 9447 597
rect 9413 563 9447 573
rect 9505 573 9539 597
rect 9505 563 9539 573
rect 9597 573 9631 597
rect 9597 563 9631 573
rect 9689 573 9723 597
rect 9689 563 9723 573
rect 9781 573 9815 597
rect 9781 563 9815 573
rect 9873 573 9907 597
rect 9873 563 9907 573
rect 9965 573 9999 597
rect 9965 563 9999 573
rect 10057 573 10091 597
rect 10057 563 10091 573
rect 10149 573 10183 597
rect 10149 563 10183 573
rect 10241 573 10275 597
rect 10241 563 10275 573
rect 10333 573 10367 597
rect 10333 563 10367 573
rect 10425 573 10459 597
rect 10425 563 10459 573
rect 10517 573 10551 597
rect 10517 563 10551 573
rect 10609 573 10643 597
rect 10609 563 10643 573
rect 10701 573 10735 597
rect 10701 563 10735 573
rect 10793 573 10827 597
rect 10793 563 10827 573
rect 10885 573 10919 597
rect 10885 563 10919 573
rect 10977 573 11011 597
rect 10977 563 11011 573
rect 11069 573 11103 597
rect 11069 563 11103 573
rect 11161 573 11195 597
rect 11161 563 11195 573
rect 11253 573 11287 597
rect 11253 563 11287 573
rect 11345 573 11379 597
rect 11345 563 11379 573
rect 11437 573 11471 597
rect 11437 563 11471 573
rect 11529 573 11563 597
rect 11529 563 11563 573
rect 11621 573 11655 597
rect 11621 563 11655 573
rect 11713 573 11747 597
rect 11713 563 11747 573
rect 11805 573 11839 597
rect 11805 563 11839 573
rect 11897 573 11931 597
rect 11897 563 11931 573
rect 11989 573 12023 597
rect 11989 563 12023 573
rect 12081 573 12115 597
rect 12081 563 12115 573
rect 12173 573 12207 597
rect 12173 563 12207 573
rect 12265 573 12299 597
rect 12265 563 12299 573
rect 12357 573 12391 597
rect 12357 563 12391 573
rect 12449 573 12483 597
rect 12449 563 12483 573
rect 12541 573 12575 597
rect 12541 563 12575 573
rect 12633 573 12667 597
rect 12633 563 12667 573
rect 12725 573 12759 597
rect 12725 563 12759 573
rect 12817 573 12851 597
rect 12817 563 12851 573
rect 12909 573 12943 597
rect 12909 563 12943 573
rect 13001 573 13035 597
rect 13001 563 13035 573
rect 13093 573 13127 597
rect 13093 563 13127 573
rect 13185 573 13219 597
rect 13185 563 13219 573
rect 13277 573 13311 597
rect 13277 563 13311 573
rect 13369 573 13403 597
rect 13369 563 13403 573
rect 13461 573 13495 597
rect 13461 563 13495 573
rect 13553 573 13587 597
rect 13553 563 13587 573
rect 13645 573 13679 597
rect 13645 563 13679 573
rect 13737 573 13771 597
rect 13737 563 13771 573
rect 13829 573 13863 597
rect 13829 563 13863 573
rect 13921 573 13955 597
rect 13921 563 13955 573
rect 14013 573 14047 597
rect 14013 563 14047 573
rect 14105 573 14139 597
rect 14105 563 14139 573
rect 14197 573 14231 597
rect 14197 563 14231 573
rect 14289 573 14323 597
rect 14289 563 14323 573
rect 14381 573 14415 597
rect 14381 563 14415 573
rect 14473 573 14507 597
rect 14473 563 14507 573
rect 14565 573 14599 597
rect 14565 563 14599 573
rect 14657 573 14691 597
rect 14657 563 14691 573
rect 14749 573 14783 597
rect 14749 563 14783 573
rect 14841 573 14875 597
rect 14841 563 14875 573
rect 14933 573 14967 597
rect 14933 563 14967 573
rect 15025 573 15059 597
rect 15025 563 15059 573
rect 15117 573 15151 597
rect 15117 563 15151 573
rect 15209 573 15243 597
rect 15209 563 15243 573
rect 15301 573 15335 597
rect 15301 563 15335 573
rect 15393 573 15427 597
rect 15393 563 15427 573
rect 15485 573 15519 597
rect 15485 563 15519 573
rect 15577 573 15611 597
rect 15577 563 15611 573
rect 15669 573 15703 597
rect 15669 563 15703 573
rect 15761 573 15795 597
rect 15761 563 15795 573
rect 15853 573 15887 597
rect 15853 563 15887 573
rect 15945 573 15979 597
rect 15945 563 15979 573
rect 16037 573 16071 597
rect 16037 563 16071 573
rect 16129 573 16163 597
rect 16129 563 16163 573
rect 16221 573 16255 597
rect 16221 563 16255 573
rect 16313 573 16347 597
rect 16313 563 16347 573
rect 16405 573 16439 597
rect 16405 563 16439 573
rect 16497 573 16531 597
rect 16497 563 16531 573
rect 16589 573 16623 597
rect 16589 563 16623 573
rect 16681 573 16715 597
rect 16681 563 16715 573
rect 29 442 63 452
rect 29 418 63 442
rect 121 442 155 452
rect 121 418 155 442
rect 213 442 247 452
rect 213 418 247 442
rect 305 442 339 452
rect 397 442 428 452
rect 428 442 431 452
rect 305 418 339 442
rect 397 418 431 442
rect 489 442 496 452
rect 496 442 523 452
rect 581 442 615 452
rect 489 418 523 442
rect 581 418 615 442
rect 673 442 707 452
rect 673 418 707 442
rect 765 442 799 452
rect 765 418 799 442
rect 857 442 891 452
rect 857 418 891 442
rect 949 442 983 452
rect 949 418 983 442
rect 1041 442 1075 452
rect 1041 418 1075 442
rect 1133 442 1167 452
rect 1133 418 1167 442
rect 1225 442 1259 452
rect 1225 418 1259 442
rect 1317 442 1351 452
rect 1317 418 1351 442
rect 1409 442 1443 452
rect 1409 418 1443 442
rect 1501 442 1535 452
rect 1501 418 1535 442
rect 1593 438 1607 452
rect 1607 438 1627 452
rect 1593 418 1627 438
rect 1685 418 1719 452
rect 1777 442 1811 452
rect 1777 418 1811 442
rect 1869 442 1903 452
rect 1869 418 1903 442
rect 1961 442 1995 452
rect 1961 418 1995 442
rect 2053 442 2087 452
rect 2053 418 2087 442
rect 2145 442 2179 452
rect 2145 418 2179 442
rect 2237 442 2271 452
rect 2237 418 2271 442
rect 2329 442 2363 452
rect 2329 418 2363 442
rect 2421 442 2455 452
rect 2421 418 2455 442
rect 2513 442 2547 452
rect 2513 418 2547 442
rect 2605 442 2639 452
rect 2605 418 2639 442
rect 2697 442 2731 452
rect 2697 418 2731 442
rect 2789 442 2791 452
rect 2791 442 2823 452
rect 2881 442 2882 452
rect 2882 442 2915 452
rect 2973 442 3007 452
rect 2789 418 2823 442
rect 2881 418 2915 442
rect 2973 418 3007 442
rect 3065 442 3099 452
rect 3065 418 3099 442
rect 3157 442 3191 452
rect 3157 418 3191 442
rect 3249 442 3283 452
rect 3249 418 3283 442
rect 3341 442 3375 452
rect 3341 418 3375 442
rect 3433 442 3467 452
rect 3433 418 3467 442
rect 3525 442 3559 452
rect 3525 418 3559 442
rect 3617 442 3651 452
rect 3617 418 3651 442
rect 3709 442 3743 452
rect 3709 418 3743 442
rect 3801 442 3835 452
rect 3801 418 3835 442
rect 3893 442 3927 452
rect 3893 418 3927 442
rect 3985 438 3999 452
rect 3999 438 4019 452
rect 3985 418 4019 438
rect 4077 418 4111 452
rect 4169 442 4203 452
rect 4169 418 4203 442
rect 4261 442 4295 452
rect 4261 418 4295 442
rect 4353 442 4387 452
rect 4353 418 4387 442
rect 4445 442 4479 452
rect 4445 418 4479 442
rect 4537 442 4571 452
rect 4537 418 4571 442
rect 4629 442 4663 452
rect 4629 418 4663 442
rect 4721 442 4755 452
rect 4721 418 4755 442
rect 4813 442 4847 452
rect 4813 418 4847 442
rect 4905 442 4939 452
rect 4905 418 4939 442
rect 4997 442 5031 452
rect 4997 418 5031 442
rect 5089 442 5123 452
rect 5181 442 5213 452
rect 5213 442 5215 452
rect 5089 418 5123 442
rect 5181 418 5215 442
rect 5273 442 5307 452
rect 5273 418 5307 442
rect 5365 442 5399 452
rect 5365 418 5399 442
rect 5457 442 5491 452
rect 5457 418 5491 442
rect 5549 442 5583 452
rect 5549 418 5583 442
rect 5641 442 5675 452
rect 5641 418 5675 442
rect 5733 442 5767 452
rect 5733 418 5767 442
rect 5825 442 5859 452
rect 5825 418 5859 442
rect 5917 442 5951 452
rect 5917 418 5951 442
rect 6009 442 6043 452
rect 6009 418 6043 442
rect 6101 442 6135 452
rect 6101 418 6135 442
rect 6193 442 6227 452
rect 6193 418 6227 442
rect 6285 442 6319 452
rect 6285 418 6319 442
rect 6377 438 6391 452
rect 6391 438 6411 452
rect 6377 418 6411 438
rect 6469 418 6503 452
rect 6561 442 6595 452
rect 6561 418 6595 442
rect 6653 442 6687 452
rect 6653 418 6687 442
rect 6745 442 6779 452
rect 6745 418 6779 442
rect 6837 442 6871 452
rect 6837 418 6871 442
rect 6929 442 6963 452
rect 6929 418 6963 442
rect 7021 442 7055 452
rect 7021 418 7055 442
rect 7113 442 7147 452
rect 7113 418 7147 442
rect 7205 442 7239 452
rect 7205 418 7239 442
rect 7297 442 7331 452
rect 7297 418 7331 442
rect 7389 442 7423 452
rect 7389 418 7423 442
rect 7481 442 7515 452
rect 7481 418 7515 442
rect 7573 442 7574 452
rect 7574 442 7607 452
rect 7665 442 7699 452
rect 7573 418 7607 442
rect 7665 418 7699 442
rect 7757 442 7791 452
rect 7757 418 7791 442
rect 7849 442 7883 452
rect 7849 418 7883 442
rect 7941 442 7975 452
rect 7941 418 7975 442
rect 8033 442 8067 452
rect 8033 418 8067 442
rect 8125 442 8159 452
rect 8125 418 8159 442
rect 8217 442 8251 452
rect 8217 418 8251 442
rect 8309 442 8343 452
rect 8309 418 8343 442
rect 8401 442 8435 452
rect 8401 418 8435 442
rect 8493 442 8527 452
rect 8493 418 8527 442
rect 8585 442 8619 452
rect 8585 418 8619 442
rect 8677 442 8711 452
rect 8677 418 8711 442
rect 8769 438 8783 452
rect 8783 438 8803 452
rect 8769 418 8803 438
rect 8861 418 8895 452
rect 8953 442 8987 452
rect 8953 418 8987 442
rect 9045 442 9079 452
rect 9045 418 9079 442
rect 9137 442 9171 452
rect 9137 418 9171 442
rect 9229 442 9263 452
rect 9229 418 9263 442
rect 9321 442 9355 452
rect 9321 418 9355 442
rect 9413 442 9447 452
rect 9413 418 9447 442
rect 9505 442 9539 452
rect 9505 418 9539 442
rect 9597 442 9631 452
rect 9597 418 9631 442
rect 9689 442 9723 452
rect 9689 418 9723 442
rect 9781 442 9815 452
rect 9781 418 9815 442
rect 9873 442 9907 452
rect 9965 442 9997 452
rect 9997 442 9999 452
rect 9873 418 9907 442
rect 9965 418 9999 442
rect 10057 442 10058 452
rect 10058 442 10091 452
rect 10149 442 10183 452
rect 10057 418 10091 442
rect 10149 418 10183 442
rect 10241 442 10275 452
rect 10241 418 10275 442
rect 10333 442 10367 452
rect 10333 418 10367 442
rect 10425 442 10459 452
rect 10425 418 10459 442
rect 10517 442 10551 452
rect 10517 418 10551 442
rect 10609 442 10643 452
rect 10609 418 10643 442
rect 10701 442 10735 452
rect 10701 418 10735 442
rect 10793 442 10827 452
rect 10793 418 10827 442
rect 10885 442 10919 452
rect 10885 418 10919 442
rect 10977 442 11011 452
rect 10977 418 11011 442
rect 11069 442 11103 452
rect 11069 418 11103 442
rect 11161 438 11175 452
rect 11175 438 11195 452
rect 11161 418 11195 438
rect 11253 418 11287 452
rect 11345 442 11379 452
rect 11345 418 11379 442
rect 11437 442 11471 452
rect 11437 418 11471 442
rect 11529 442 11563 452
rect 11529 418 11563 442
rect 11621 442 11655 452
rect 11621 418 11655 442
rect 11713 442 11747 452
rect 11713 418 11747 442
rect 11805 442 11839 452
rect 11805 418 11839 442
rect 11897 442 11931 452
rect 11897 418 11931 442
rect 11989 442 12023 452
rect 11989 418 12023 442
rect 12081 442 12115 452
rect 12081 418 12115 442
rect 12173 442 12207 452
rect 12173 418 12207 442
rect 12265 442 12299 452
rect 12265 418 12299 442
rect 12357 442 12391 452
rect 12449 442 12482 452
rect 12482 442 12483 452
rect 12357 418 12391 442
rect 12449 418 12483 442
rect 12541 442 12575 452
rect 12541 418 12575 442
rect 12633 442 12667 452
rect 12633 418 12667 442
rect 12725 442 12759 452
rect 12725 418 12759 442
rect 12817 442 12851 452
rect 12817 418 12851 442
rect 12909 442 12943 452
rect 12909 418 12943 442
rect 13001 442 13035 452
rect 13001 418 13035 442
rect 13093 442 13127 452
rect 13093 418 13127 442
rect 13185 442 13219 452
rect 13185 418 13219 442
rect 13277 442 13311 452
rect 13277 418 13311 442
rect 13369 442 13403 452
rect 13369 418 13403 442
rect 13461 442 13495 452
rect 13461 418 13495 442
rect 13553 438 13567 452
rect 13567 438 13587 452
rect 13553 418 13587 438
rect 13645 418 13679 452
rect 13737 442 13771 452
rect 13737 418 13771 442
rect 13829 442 13863 452
rect 13829 418 13863 442
rect 13921 442 13955 452
rect 13921 418 13955 442
rect 14013 442 14047 452
rect 14013 418 14047 442
rect 14105 442 14139 452
rect 14105 418 14139 442
rect 14197 442 14231 452
rect 14197 418 14231 442
rect 14289 442 14323 452
rect 14289 418 14323 442
rect 14381 442 14415 452
rect 14381 418 14415 442
rect 14473 442 14507 452
rect 14473 418 14507 442
rect 14565 442 14599 452
rect 14565 418 14599 442
rect 14657 442 14691 452
rect 14749 442 14782 452
rect 14782 442 14783 452
rect 14657 418 14691 442
rect 14749 418 14783 442
rect 14841 442 14842 452
rect 14842 442 14875 452
rect 14933 442 14967 452
rect 14841 418 14875 442
rect 14933 418 14967 442
rect 15025 442 15059 452
rect 15025 418 15059 442
rect 15117 442 15151 452
rect 15117 418 15151 442
rect 15209 442 15243 452
rect 15209 418 15243 442
rect 15301 442 15335 452
rect 15301 418 15335 442
rect 15393 442 15427 452
rect 15393 418 15427 442
rect 15485 442 15519 452
rect 15485 418 15519 442
rect 15577 442 15611 452
rect 15577 418 15611 442
rect 15669 442 15703 452
rect 15669 418 15703 442
rect 15761 442 15795 452
rect 15761 418 15795 442
rect 15853 442 15887 452
rect 15853 418 15887 442
rect 15945 435 15959 452
rect 15959 435 15979 452
rect 15945 418 15979 435
rect 16037 418 16071 452
rect 16129 442 16163 452
rect 16129 418 16163 442
rect 16221 442 16255 452
rect 16221 418 16255 442
rect 16313 442 16347 452
rect 16313 418 16347 442
rect 16405 442 16439 452
rect 16405 418 16439 442
rect 16497 442 16531 452
rect 16497 418 16531 442
rect 16589 442 16623 452
rect 16589 418 16623 442
rect 16681 442 16715 452
rect 16681 418 16715 442
rect 26 340 60 342
rect 26 308 35 340
rect 35 308 60 340
rect 306 271 340 276
rect 306 242 318 271
rect 318 242 340 271
rect 587 180 621 214
rect 502 144 536 148
rect 502 114 529 144
rect 529 114 536 144
rect 843 70 847 78
rect 847 70 877 78
rect 843 44 877 70
rect 1133 256 1167 282
rect 1133 248 1146 256
rect 1146 248 1167 256
rect 1225 180 1259 214
rect 1133 112 1167 146
rect 1869 248 1903 282
rect 1593 70 1625 78
rect 1625 70 1627 78
rect 1593 44 1627 70
rect 1777 60 1797 78
rect 1797 60 1811 78
rect 1777 44 1811 60
rect 1968 115 2002 149
rect 2145 266 2155 282
rect 2155 266 2179 282
rect 2145 248 2179 266
rect 2418 340 2452 342
rect 2418 308 2427 340
rect 2427 308 2452 340
rect 2314 171 2348 205
rect 2236 44 2270 78
rect 2698 271 2732 276
rect 2698 242 2710 271
rect 2710 242 2732 271
rect 2979 180 3013 214
rect 2891 144 2925 150
rect 2891 116 2921 144
rect 2921 116 2925 144
rect 3235 70 3239 78
rect 3239 70 3269 78
rect 3235 44 3269 70
rect 3525 256 3559 282
rect 3525 248 3538 256
rect 3538 248 3559 256
rect 3617 180 3651 214
rect 3525 112 3559 146
rect 4261 248 4295 282
rect 3985 70 4017 78
rect 4017 70 4019 78
rect 3985 44 4019 70
rect 4169 60 4189 78
rect 4189 60 4203 78
rect 4169 44 4203 60
rect 4360 115 4394 149
rect 4537 266 4547 282
rect 4547 266 4571 282
rect 4537 248 4571 266
rect 4811 340 4845 342
rect 4811 308 4819 340
rect 4819 308 4845 340
rect 4708 171 4742 205
rect 4628 44 4662 78
rect 5089 271 5123 276
rect 5089 242 5102 271
rect 5102 242 5123 271
rect 5371 180 5405 214
rect 5284 144 5318 150
rect 5284 116 5313 144
rect 5313 116 5318 144
rect 5627 70 5631 78
rect 5631 70 5661 78
rect 5627 44 5661 70
rect 5917 256 5951 282
rect 5917 248 5930 256
rect 5930 248 5951 256
rect 6009 180 6043 214
rect 5917 112 5951 146
rect 6653 248 6687 282
rect 6377 70 6409 78
rect 6409 70 6411 78
rect 6377 44 6411 70
rect 6561 60 6581 78
rect 6581 60 6595 78
rect 6561 44 6595 60
rect 6751 116 6785 150
rect 6929 266 6939 282
rect 6939 266 6963 282
rect 6929 248 6963 266
rect 7202 340 7236 342
rect 7202 308 7211 340
rect 7211 308 7236 340
rect 7098 173 7132 207
rect 7020 44 7054 78
rect 7482 271 7516 276
rect 7482 242 7494 271
rect 7494 242 7516 271
rect 7763 180 7797 214
rect 7677 144 7711 150
rect 7677 116 7705 144
rect 7705 116 7711 144
rect 8019 70 8023 78
rect 8023 70 8053 78
rect 8019 44 8053 70
rect 8309 256 8343 282
rect 8309 248 8322 256
rect 8322 248 8343 256
rect 8401 180 8435 214
rect 8309 112 8343 146
rect 9045 248 9079 282
rect 8769 70 8801 78
rect 8801 70 8803 78
rect 8769 44 8803 70
rect 8953 60 8973 78
rect 8973 60 8987 78
rect 8953 44 8987 60
rect 9144 115 9178 149
rect 9321 266 9331 282
rect 9331 266 9355 282
rect 9321 248 9355 266
rect 9594 340 9628 341
rect 9594 307 9603 340
rect 9603 307 9628 340
rect 9490 171 9524 205
rect 9412 44 9446 78
rect 9874 271 9908 276
rect 9874 242 9886 271
rect 9886 242 9908 271
rect 10155 180 10189 214
rect 10068 144 10102 150
rect 10068 116 10097 144
rect 10097 116 10102 144
rect 10411 70 10415 78
rect 10415 70 10445 78
rect 10411 44 10445 70
rect 10701 256 10735 282
rect 10701 248 10714 256
rect 10714 248 10735 256
rect 10793 180 10827 214
rect 10701 112 10735 146
rect 11437 248 11471 282
rect 11161 70 11193 78
rect 11193 70 11195 78
rect 11161 44 11195 70
rect 11345 60 11365 78
rect 11365 60 11379 78
rect 11345 44 11379 60
rect 11535 115 11569 149
rect 11713 266 11723 282
rect 11723 266 11747 282
rect 11713 248 11747 266
rect 11987 340 12021 343
rect 11987 309 11995 340
rect 11995 309 12021 340
rect 11882 173 11916 207
rect 11804 44 11838 78
rect 12265 271 12299 277
rect 12265 243 12278 271
rect 12278 243 12299 271
rect 12547 180 12581 214
rect 12461 144 12495 150
rect 12461 116 12489 144
rect 12489 116 12495 144
rect 12803 70 12807 78
rect 12807 70 12837 78
rect 12803 44 12837 70
rect 13093 256 13127 282
rect 13093 248 13106 256
rect 13106 248 13127 256
rect 13185 180 13219 214
rect 13093 112 13127 146
rect 13829 248 13863 282
rect 13553 70 13585 78
rect 13585 70 13587 78
rect 13553 44 13587 70
rect 13737 60 13757 78
rect 13757 60 13771 78
rect 13737 44 13771 60
rect 13928 115 13962 149
rect 14105 266 14115 282
rect 14115 266 14139 282
rect 14105 248 14139 266
rect 14378 340 14412 343
rect 14378 309 14387 340
rect 14387 309 14412 340
rect 14274 171 14308 205
rect 14196 44 14230 78
rect 14658 271 14692 276
rect 14658 242 14670 271
rect 14670 242 14692 271
rect 14939 180 14973 214
rect 14852 144 14886 150
rect 14852 116 14881 144
rect 14881 116 14886 144
rect 15195 70 15199 78
rect 15199 70 15229 78
rect 15195 44 15229 70
rect 15485 256 15519 282
rect 15485 248 15498 256
rect 15498 248 15519 256
rect 15577 180 15611 214
rect 15485 112 15519 146
rect 16221 248 16255 282
rect 15945 70 15977 78
rect 15977 70 15979 78
rect 15945 44 15979 70
rect 16129 60 16149 78
rect 16149 60 16163 78
rect 16129 44 16163 60
rect 16321 115 16355 149
rect 16497 266 16507 282
rect 16507 266 16531 282
rect 16497 248 16531 266
rect 16666 173 16700 207
rect 16588 44 16622 78
rect 29 -116 63 -92
rect 29 -126 63 -116
rect 121 -116 155 -92
rect 121 -126 155 -116
rect 213 -116 247 -92
rect 213 -126 247 -116
rect 305 -116 339 -92
rect 305 -126 339 -116
rect 397 -116 431 -92
rect 397 -126 431 -116
rect 489 -116 523 -92
rect 489 -126 523 -116
rect 581 -116 615 -92
rect 581 -126 615 -116
rect 673 -116 707 -92
rect 673 -126 707 -116
rect 765 -116 799 -92
rect 765 -126 799 -116
rect 857 -116 891 -92
rect 857 -126 891 -116
rect 949 -116 983 -92
rect 949 -126 983 -116
rect 1041 -116 1075 -92
rect 1041 -126 1075 -116
rect 1133 -116 1167 -92
rect 1133 -126 1167 -116
rect 1225 -116 1259 -92
rect 1225 -126 1259 -116
rect 1317 -116 1351 -92
rect 1317 -126 1351 -116
rect 1409 -116 1443 -92
rect 1409 -126 1443 -116
rect 1501 -116 1535 -92
rect 1501 -126 1535 -116
rect 1593 -116 1627 -92
rect 1593 -126 1627 -116
rect 1685 -116 1719 -92
rect 1685 -126 1719 -116
rect 1777 -116 1811 -92
rect 1777 -126 1811 -116
rect 1869 -116 1903 -92
rect 1869 -126 1903 -116
rect 1961 -116 1995 -92
rect 1961 -126 1995 -116
rect 2053 -116 2087 -92
rect 2053 -126 2087 -116
rect 2145 -116 2179 -92
rect 2145 -126 2179 -116
rect 2237 -116 2271 -92
rect 2237 -126 2271 -116
rect 2329 -116 2363 -92
rect 2329 -126 2363 -116
rect 2421 -116 2455 -92
rect 2421 -126 2455 -116
rect 2513 -116 2547 -92
rect 2513 -126 2547 -116
rect 2605 -116 2639 -92
rect 2605 -126 2639 -116
rect 2697 -116 2731 -92
rect 2697 -126 2731 -116
rect 2789 -116 2823 -92
rect 2789 -126 2823 -116
rect 2881 -116 2915 -92
rect 2881 -126 2915 -116
rect 2973 -116 3007 -92
rect 2973 -126 3007 -116
rect 3065 -116 3099 -92
rect 3065 -126 3099 -116
rect 3157 -116 3191 -92
rect 3157 -126 3191 -116
rect 3249 -116 3283 -92
rect 3249 -126 3283 -116
rect 3341 -116 3375 -92
rect 3341 -126 3375 -116
rect 3433 -116 3467 -92
rect 3433 -126 3467 -116
rect 3525 -116 3559 -92
rect 3525 -126 3559 -116
rect 3617 -116 3651 -92
rect 3617 -126 3651 -116
rect 3709 -116 3743 -92
rect 3709 -126 3743 -116
rect 3801 -116 3835 -92
rect 3801 -126 3835 -116
rect 3893 -116 3927 -92
rect 3893 -126 3927 -116
rect 3985 -116 4019 -92
rect 3985 -126 4019 -116
rect 4077 -116 4111 -92
rect 4077 -126 4111 -116
rect 4169 -116 4203 -92
rect 4169 -126 4203 -116
rect 4261 -116 4295 -92
rect 4261 -126 4295 -116
rect 4353 -116 4387 -92
rect 4353 -126 4387 -116
rect 4445 -116 4479 -92
rect 4445 -126 4479 -116
rect 4537 -116 4571 -92
rect 4537 -126 4571 -116
rect 4629 -116 4663 -92
rect 4629 -126 4663 -116
rect 4721 -116 4755 -92
rect 4721 -126 4755 -116
rect 4813 -116 4847 -92
rect 4813 -126 4847 -116
rect 4905 -116 4939 -92
rect 4905 -126 4939 -116
rect 4997 -116 5031 -92
rect 4997 -126 5031 -116
rect 5089 -116 5123 -92
rect 5089 -126 5123 -116
rect 5181 -116 5215 -92
rect 5181 -126 5215 -116
rect 5273 -116 5307 -92
rect 5273 -126 5307 -116
rect 5365 -116 5399 -92
rect 5365 -126 5399 -116
rect 5457 -116 5491 -92
rect 5457 -126 5491 -116
rect 5549 -116 5583 -92
rect 5549 -126 5583 -116
rect 5641 -116 5675 -92
rect 5641 -126 5675 -116
rect 5733 -116 5767 -92
rect 5733 -126 5767 -116
rect 5825 -116 5859 -92
rect 5825 -126 5859 -116
rect 5917 -116 5951 -92
rect 5917 -126 5951 -116
rect 6009 -116 6043 -92
rect 6009 -126 6043 -116
rect 6101 -116 6135 -92
rect 6101 -126 6135 -116
rect 6193 -116 6227 -92
rect 6193 -126 6227 -116
rect 6285 -116 6319 -92
rect 6285 -126 6319 -116
rect 6377 -116 6411 -92
rect 6377 -126 6411 -116
rect 6469 -116 6503 -92
rect 6469 -126 6503 -116
rect 6561 -116 6595 -92
rect 6561 -126 6595 -116
rect 6653 -116 6687 -92
rect 6653 -126 6687 -116
rect 6745 -116 6779 -92
rect 6745 -126 6779 -116
rect 6837 -116 6871 -92
rect 6837 -126 6871 -116
rect 6929 -116 6963 -92
rect 6929 -126 6963 -116
rect 7021 -116 7055 -92
rect 7021 -126 7055 -116
rect 7113 -116 7147 -92
rect 7113 -126 7147 -116
rect 7205 -116 7239 -92
rect 7205 -126 7239 -116
rect 7297 -116 7331 -92
rect 7297 -126 7331 -116
rect 7389 -116 7423 -92
rect 7389 -126 7423 -116
rect 7481 -116 7515 -92
rect 7481 -126 7515 -116
rect 7573 -116 7607 -92
rect 7573 -126 7607 -116
rect 7665 -116 7699 -92
rect 7665 -126 7699 -116
rect 7757 -116 7791 -92
rect 7757 -126 7791 -116
rect 7849 -116 7883 -92
rect 7849 -126 7883 -116
rect 7941 -116 7975 -92
rect 7941 -126 7975 -116
rect 8033 -116 8067 -92
rect 8033 -126 8067 -116
rect 8125 -116 8159 -92
rect 8125 -126 8159 -116
rect 8217 -116 8251 -92
rect 8217 -126 8251 -116
rect 8309 -116 8343 -92
rect 8309 -126 8343 -116
rect 8401 -116 8435 -92
rect 8401 -126 8435 -116
rect 8493 -116 8527 -92
rect 8493 -126 8527 -116
rect 8585 -116 8619 -92
rect 8585 -126 8619 -116
rect 8677 -116 8711 -92
rect 8677 -126 8711 -116
rect 8769 -116 8803 -92
rect 8769 -126 8803 -116
rect 8861 -116 8895 -92
rect 8861 -126 8895 -116
rect 8953 -116 8987 -92
rect 8953 -126 8987 -116
rect 9045 -116 9079 -92
rect 9045 -126 9079 -116
rect 9137 -116 9171 -92
rect 9137 -126 9171 -116
rect 9229 -116 9263 -92
rect 9229 -126 9263 -116
rect 9321 -116 9355 -92
rect 9321 -126 9355 -116
rect 9413 -116 9447 -92
rect 9413 -126 9447 -116
rect 9505 -116 9539 -92
rect 9505 -126 9539 -116
rect 9597 -116 9631 -92
rect 9597 -126 9631 -116
rect 9689 -116 9723 -92
rect 9689 -126 9723 -116
rect 9781 -116 9815 -92
rect 9781 -126 9815 -116
rect 9873 -116 9907 -92
rect 9873 -126 9907 -116
rect 9965 -116 9999 -92
rect 9965 -126 9999 -116
rect 10057 -116 10091 -92
rect 10057 -126 10091 -116
rect 10149 -116 10183 -92
rect 10149 -126 10183 -116
rect 10241 -116 10275 -92
rect 10241 -126 10275 -116
rect 10333 -116 10367 -92
rect 10333 -126 10367 -116
rect 10425 -116 10459 -92
rect 10425 -126 10459 -116
rect 10517 -116 10551 -92
rect 10517 -126 10551 -116
rect 10609 -116 10643 -92
rect 10609 -126 10643 -116
rect 10701 -116 10735 -92
rect 10701 -126 10735 -116
rect 10793 -116 10827 -92
rect 10793 -126 10827 -116
rect 10885 -116 10919 -92
rect 10885 -126 10919 -116
rect 10977 -116 11011 -92
rect 10977 -126 11011 -116
rect 11069 -116 11103 -92
rect 11069 -126 11103 -116
rect 11161 -116 11195 -92
rect 11161 -126 11195 -116
rect 11253 -116 11287 -92
rect 11253 -126 11287 -116
rect 11345 -116 11379 -92
rect 11345 -126 11379 -116
rect 11437 -116 11471 -92
rect 11437 -126 11471 -116
rect 11529 -116 11563 -92
rect 11529 -126 11563 -116
rect 11621 -116 11655 -92
rect 11621 -126 11655 -116
rect 11713 -116 11747 -92
rect 11713 -126 11747 -116
rect 11805 -116 11839 -92
rect 11805 -126 11839 -116
rect 11897 -116 11931 -92
rect 11897 -126 11931 -116
rect 11989 -116 12023 -92
rect 11989 -126 12023 -116
rect 12081 -116 12115 -92
rect 12081 -126 12115 -116
rect 12173 -116 12207 -92
rect 12173 -126 12207 -116
rect 12265 -116 12299 -92
rect 12265 -126 12299 -116
rect 12357 -116 12391 -92
rect 12357 -126 12391 -116
rect 12449 -116 12483 -92
rect 12449 -126 12483 -116
rect 12541 -116 12575 -92
rect 12541 -126 12575 -116
rect 12633 -116 12667 -92
rect 12633 -126 12667 -116
rect 12725 -116 12759 -92
rect 12725 -126 12759 -116
rect 12817 -116 12851 -92
rect 12817 -126 12851 -116
rect 12909 -116 12943 -92
rect 12909 -126 12943 -116
rect 13001 -116 13035 -92
rect 13001 -126 13035 -116
rect 13093 -116 13127 -92
rect 13093 -126 13127 -116
rect 13185 -116 13219 -92
rect 13185 -126 13219 -116
rect 13277 -116 13311 -92
rect 13277 -126 13311 -116
rect 13369 -116 13403 -92
rect 13369 -126 13403 -116
rect 13461 -116 13495 -92
rect 13461 -126 13495 -116
rect 13553 -116 13587 -92
rect 13553 -126 13587 -116
rect 13645 -116 13679 -92
rect 13645 -126 13679 -116
rect 13737 -116 13771 -92
rect 13737 -126 13771 -116
rect 13829 -116 13863 -92
rect 13829 -126 13863 -116
rect 13921 -116 13955 -92
rect 13921 -126 13955 -116
rect 14013 -116 14047 -92
rect 14013 -126 14047 -116
rect 14105 -116 14139 -92
rect 14105 -126 14139 -116
rect 14197 -116 14231 -92
rect 14197 -126 14231 -116
rect 14289 -116 14323 -92
rect 14289 -126 14323 -116
rect 14381 -116 14415 -92
rect 14381 -126 14415 -116
rect 14473 -116 14507 -92
rect 14473 -126 14507 -116
rect 14565 -116 14599 -92
rect 14565 -126 14599 -116
rect 14657 -116 14691 -92
rect 14657 -126 14691 -116
rect 14749 -116 14783 -92
rect 14749 -126 14783 -116
rect 14841 -116 14875 -92
rect 14841 -126 14875 -116
rect 14933 -116 14967 -92
rect 14933 -126 14967 -116
rect 15025 -116 15059 -92
rect 15025 -126 15059 -116
rect 15117 -116 15151 -92
rect 15117 -126 15151 -116
rect 15209 -116 15243 -92
rect 15209 -126 15243 -116
rect 15301 -116 15335 -92
rect 15301 -126 15335 -116
rect 15393 -116 15427 -92
rect 15393 -126 15427 -116
rect 15485 -116 15519 -92
rect 15485 -126 15519 -116
rect 15577 -116 15611 -92
rect 15577 -126 15611 -116
rect 15669 -116 15703 -92
rect 15669 -126 15703 -116
rect 15761 -116 15795 -92
rect 15761 -126 15795 -116
rect 15853 -116 15887 -92
rect 15853 -126 15887 -116
rect 15945 -116 15979 -92
rect 15945 -126 15979 -116
rect 16037 -116 16071 -92
rect 16037 -126 16071 -116
rect 16129 -116 16163 -92
rect 16129 -126 16163 -116
rect 16221 -116 16255 -92
rect 16221 -126 16255 -116
rect 16313 -116 16347 -92
rect 16313 -126 16347 -116
rect 16405 -116 16439 -92
rect 16405 -126 16439 -116
rect 16497 -116 16531 -92
rect 16497 -126 16531 -116
rect 16589 -116 16623 -92
rect 16589 -126 16623 -116
rect 16681 -116 16715 -92
rect 16681 -126 16715 -116
<< metal1 >>
rect -126 2980 15690 3002
rect -126 2978 1265 2980
rect -126 2976 255 2978
rect -126 2971 53 2976
rect 105 2971 255 2976
rect -126 2937 31 2971
rect 105 2937 123 2971
rect 157 2937 215 2971
rect 249 2937 255 2971
rect -126 2924 53 2937
rect 105 2926 255 2937
rect 307 2976 864 2978
rect 307 2971 466 2976
rect 518 2971 656 2976
rect 708 2971 864 2976
rect 916 2971 1066 2978
rect 1118 2971 1265 2978
rect 341 2937 399 2971
rect 433 2937 466 2971
rect 525 2937 583 2971
rect 617 2937 656 2971
rect 709 2937 767 2971
rect 801 2937 859 2971
rect 916 2937 951 2971
rect 985 2937 1043 2971
rect 1118 2937 1135 2971
rect 1169 2937 1227 2971
rect 1261 2937 1265 2971
rect 307 2926 466 2937
rect 105 2924 466 2926
rect 518 2924 656 2937
rect 708 2926 864 2937
rect 916 2926 1066 2937
rect 1118 2928 1265 2937
rect 1317 2979 2152 2980
rect 1317 2977 1661 2979
rect 1317 2971 1460 2977
rect 1512 2971 1661 2977
rect 1713 2977 2152 2979
rect 1713 2971 1878 2977
rect 1930 2971 2152 2977
rect 2204 2976 15690 2980
rect 2204 2973 2652 2976
rect 2204 2971 2429 2973
rect 2481 2971 2652 2973
rect 2704 2975 15690 2976
rect 2704 2971 2884 2975
rect 1317 2937 1319 2971
rect 1353 2937 1411 2971
rect 1445 2937 1460 2971
rect 1537 2937 1595 2971
rect 1629 2937 1661 2971
rect 1721 2937 1779 2971
rect 1813 2937 1871 2971
rect 1930 2937 1963 2971
rect 1997 2937 2055 2971
rect 2089 2937 2147 2971
rect 2204 2937 2239 2971
rect 2273 2937 2331 2971
rect 2365 2937 2423 2971
rect 2481 2937 2515 2971
rect 2549 2937 2607 2971
rect 2641 2937 2652 2971
rect 2733 2937 2791 2971
rect 2825 2937 2884 2971
rect 1317 2928 1460 2937
rect 1118 2926 1460 2928
rect 708 2925 1460 2926
rect 1512 2927 1661 2937
rect 1713 2927 1878 2937
rect 1512 2925 1878 2927
rect 1930 2928 2152 2937
rect 2204 2928 2429 2937
rect 1930 2925 2429 2928
rect 708 2924 2429 2925
rect -126 2921 2429 2924
rect 2481 2924 2652 2937
rect 2704 2924 2884 2937
rect 2481 2923 2884 2924
rect 2936 2974 5903 2975
rect 2936 2973 5028 2974
rect 2936 2972 4828 2973
rect 2936 2971 4520 2972
rect 4572 2971 4828 2972
rect 4880 2971 5028 2973
rect 5080 2973 5701 2974
rect 5080 2971 5247 2973
rect 5299 2972 5701 2973
rect 5299 2971 5493 2972
rect 5545 2971 5701 2972
rect 5753 2971 5903 2974
rect 5955 2974 15690 2975
rect 5955 2971 6096 2974
rect 6148 2973 15690 2974
rect 6148 2971 6468 2973
rect 6520 2971 7220 2973
rect 2936 2937 4415 2971
rect 4449 2937 4507 2971
rect 4572 2937 4599 2971
rect 4633 2937 4691 2971
rect 4725 2937 4783 2971
rect 4817 2937 4828 2971
rect 4909 2937 4967 2971
rect 5001 2937 5028 2971
rect 5093 2937 5151 2971
rect 5185 2937 5243 2971
rect 5299 2937 5335 2971
rect 5369 2937 5427 2971
rect 5461 2937 5493 2971
rect 5553 2937 5611 2971
rect 5645 2937 5701 2971
rect 5753 2937 5795 2971
rect 5829 2937 5887 2971
rect 5955 2937 5979 2971
rect 6013 2937 6071 2971
rect 6148 2937 6163 2971
rect 6197 2937 6255 2971
rect 6289 2937 6347 2971
rect 6381 2937 6439 2971
rect 6520 2937 6531 2971
rect 6565 2937 6623 2971
rect 2936 2923 4520 2937
rect 2481 2921 4520 2923
rect -126 2920 4520 2921
rect 4572 2921 4828 2937
rect 4880 2922 5028 2937
rect 5080 2922 5247 2937
rect 4880 2921 5247 2922
rect 5299 2921 5493 2937
rect 4572 2920 5493 2921
rect 5545 2922 5701 2937
rect 5753 2923 5903 2937
rect 5955 2923 6096 2937
rect 5753 2922 6096 2923
rect 6148 2922 6468 2937
rect 5545 2921 6468 2922
rect 6520 2921 6657 2937
rect 5545 2920 6657 2921
rect -126 2919 6657 2920
rect 6709 2937 6715 2971
rect 6749 2937 6807 2971
rect 6841 2937 6899 2971
rect 6933 2937 6947 2971
rect 7025 2937 7083 2971
rect 7117 2937 7175 2971
rect 7209 2937 7220 2971
rect 6709 2919 6947 2937
rect 6999 2921 7220 2937
rect 7272 2921 15690 2973
rect 6999 2919 15690 2921
rect -126 2906 15690 2919
rect -126 2722 -34 2756
rect -68 2681 -34 2722
rect 27 2681 85 2687
rect -68 2675 85 2681
rect -68 2647 39 2675
rect 26 2641 39 2647
rect 73 2641 85 2675
rect 26 2631 85 2641
rect 2860 2622 2866 2674
rect 2918 2622 2924 2674
rect 7164 2668 7216 2674
rect 7421 2668 7427 2674
rect 7164 2666 7427 2668
rect 4411 2658 4469 2664
rect 4411 2656 4423 2658
rect 4270 2624 4423 2656
rect 4457 2624 4469 2658
rect 4270 2560 4302 2624
rect 4411 2618 4469 2624
rect 7164 2632 7176 2666
rect 7210 2632 7427 2666
rect 7164 2626 7427 2632
rect 7164 2620 7216 2626
rect 7421 2622 7427 2626
rect 7479 2622 7485 2674
rect -126 2526 4302 2560
rect -126 2448 16861 2458
rect -126 2441 16876 2448
rect -126 2437 1390 2441
rect -126 2427 1171 2437
rect -126 2393 31 2427
rect 65 2393 123 2427
rect 157 2393 215 2427
rect 249 2393 307 2427
rect 341 2393 399 2427
rect 433 2393 491 2427
rect 525 2393 583 2427
rect 617 2393 675 2427
rect 709 2393 767 2427
rect 801 2393 859 2427
rect 893 2393 951 2427
rect 985 2393 1043 2427
rect 1077 2393 1135 2427
rect 1169 2393 1171 2427
rect -126 2385 1171 2393
rect 1223 2427 1390 2437
rect 1442 2427 1673 2441
rect 1725 2427 1882 2441
rect 1934 2440 16876 2441
rect 1934 2439 4477 2440
rect 1934 2427 2153 2439
rect 2205 2437 4477 2439
rect 2205 2427 4228 2437
rect 1223 2393 1227 2427
rect 1261 2393 1319 2427
rect 1353 2393 1390 2427
rect 1445 2393 1503 2427
rect 1537 2393 1595 2427
rect 1629 2393 1673 2427
rect 1725 2393 1779 2427
rect 1813 2393 1871 2427
rect 1934 2393 1963 2427
rect 1997 2393 2055 2427
rect 2089 2393 2147 2427
rect 2205 2393 2239 2427
rect 2273 2393 2331 2427
rect 2365 2393 2423 2427
rect 2457 2393 2515 2427
rect 2549 2393 2607 2427
rect 2641 2393 2699 2427
rect 2733 2393 2791 2427
rect 2825 2393 4228 2427
rect 1223 2389 1390 2393
rect 1442 2389 1673 2393
rect 1725 2389 1882 2393
rect 1934 2389 2153 2393
rect 1223 2387 2153 2389
rect 2205 2387 4228 2393
rect 1223 2385 4228 2387
rect 4280 2427 4477 2437
rect 4529 2439 16876 2440
rect 4529 2437 7226 2439
rect 4529 2432 7022 2437
rect 4529 2427 5075 2432
rect 5127 2427 5304 2432
rect 5356 2427 7022 2432
rect 7074 2427 7226 2437
rect 4280 2393 4415 2427
rect 4449 2393 4477 2427
rect 4541 2393 4599 2427
rect 4633 2393 4691 2427
rect 4725 2393 4783 2427
rect 4817 2426 4875 2427
rect 4817 2393 4821 2426
rect 4280 2388 4477 2393
rect 4529 2388 4821 2393
rect 4280 2385 4821 2388
rect -126 2374 4821 2385
rect 4873 2393 4875 2426
rect 4909 2393 4967 2427
rect 5001 2393 5059 2427
rect 5127 2393 5151 2427
rect 5185 2393 5243 2427
rect 5277 2393 5304 2427
rect 5369 2393 5427 2427
rect 5461 2393 5519 2427
rect 5553 2393 5611 2427
rect 5645 2393 5703 2427
rect 5737 2393 5795 2427
rect 5829 2393 5887 2427
rect 5921 2393 5979 2427
rect 6013 2393 6071 2427
rect 6105 2393 6163 2427
rect 6197 2393 6255 2427
rect 6289 2393 6347 2427
rect 6381 2393 6439 2427
rect 6473 2393 6531 2427
rect 6565 2393 6623 2427
rect 6657 2393 6715 2427
rect 6749 2393 6807 2427
rect 6841 2393 6899 2427
rect 6933 2393 6991 2427
rect 7074 2393 7083 2427
rect 7117 2393 7175 2427
rect 7209 2393 7226 2427
rect 4873 2380 5075 2393
rect 5127 2380 5304 2393
rect 5356 2385 7022 2393
rect 7074 2387 7226 2393
rect 7278 2437 16876 2439
rect 7278 2387 7549 2437
rect 7074 2385 7549 2387
rect 7601 2385 16876 2437
rect 5356 2380 16876 2385
rect 4873 2374 16876 2380
rect -126 2362 16876 2374
rect 1018 2294 1024 2303
rect 95 2260 1024 2294
rect 1018 2250 1024 2260
rect 1077 2294 1083 2303
rect 2860 2294 2866 2302
rect 1077 2260 2866 2294
rect 1077 2250 1083 2260
rect 2860 2250 2866 2260
rect 2918 2294 2924 2302
rect 3412 2294 3418 2309
rect 2918 2260 3418 2294
rect 2918 2250 2924 2260
rect 3412 2256 3418 2260
rect 3471 2294 3477 2309
rect 5803 2294 5809 2309
rect 3471 2260 5809 2294
rect 3471 2256 3477 2260
rect 3412 2255 3477 2256
rect 5803 2256 5809 2260
rect 5862 2294 5868 2309
rect 8194 2294 8200 2309
rect 5862 2260 8200 2294
rect 5862 2256 5868 2260
rect 7416 2259 7533 2260
rect 5803 2255 5868 2256
rect 8194 2256 8200 2260
rect 8253 2294 8259 2309
rect 10586 2294 10592 2309
rect 8253 2260 10592 2294
rect 8253 2256 8259 2260
rect 8194 2255 8259 2256
rect 10586 2256 10592 2260
rect 10645 2294 10651 2309
rect 12977 2294 12983 2309
rect 10645 2260 12983 2294
rect 10645 2256 10651 2260
rect 10586 2255 10651 2256
rect 12977 2256 12983 2260
rect 13036 2294 13042 2309
rect 15370 2294 15376 2309
rect 13036 2260 15376 2294
rect 13036 2256 13042 2260
rect 12977 2255 13042 2256
rect 15370 2256 15376 2260
rect 15429 2294 15435 2309
rect 15429 2260 16861 2294
rect 15429 2256 15435 2260
rect 15370 2255 15435 2256
rect 1018 2249 1083 2250
rect 95 2186 16861 2188
rect 95 2154 16876 2186
rect 7419 2153 7528 2154
rect 467 2082 474 2091
rect 95 2048 474 2082
rect 467 2039 474 2048
rect 526 2082 533 2091
rect 1729 2082 1736 2091
rect 526 2048 1736 2082
rect 526 2039 533 2048
rect 1729 2039 1736 2048
rect 1788 2082 1795 2091
rect 2860 2082 2867 2090
rect 1788 2048 2867 2082
rect 1788 2039 1795 2048
rect 2860 2038 2867 2048
rect 2919 2082 2926 2090
rect 4121 2082 4128 2091
rect 2919 2048 4128 2082
rect 2919 2038 2926 2048
rect 4121 2039 4128 2048
rect 4180 2082 4187 2091
rect 5252 2082 5259 2090
rect 4180 2048 5259 2082
rect 4180 2039 4187 2048
rect 5252 2038 5259 2048
rect 5311 2082 5318 2090
rect 6512 2082 6519 2092
rect 5311 2048 6519 2082
rect 5311 2038 5318 2048
rect 6512 2040 6519 2048
rect 6571 2082 6578 2092
rect 7421 2082 7427 2090
rect 6571 2048 7427 2082
rect 6571 2040 6578 2048
rect 7421 2038 7427 2048
rect 7479 2082 7485 2090
rect 7644 2082 7651 2091
rect 7479 2048 7651 2082
rect 7479 2038 7485 2048
rect 7644 2039 7651 2048
rect 7703 2082 7710 2091
rect 8905 2082 8912 2092
rect 7703 2048 8912 2082
rect 7703 2039 7710 2048
rect 8905 2040 8912 2048
rect 8964 2082 8971 2092
rect 10035 2082 10042 2090
rect 8964 2048 10042 2082
rect 8964 2040 8971 2048
rect 10035 2038 10042 2048
rect 10094 2082 10101 2090
rect 11298 2082 11305 2092
rect 10094 2048 11305 2082
rect 10094 2038 10101 2048
rect 11298 2040 11305 2048
rect 11357 2082 11364 2092
rect 12427 2082 12434 2089
rect 11357 2048 12434 2082
rect 11357 2040 11364 2048
rect 12427 2037 12434 2048
rect 12486 2082 12493 2089
rect 13687 2082 13694 2092
rect 12486 2048 13694 2082
rect 12486 2037 12493 2048
rect 13687 2040 13694 2048
rect 13746 2082 13753 2092
rect 14819 2082 14826 2090
rect 13746 2048 14826 2082
rect 13746 2040 13753 2048
rect 14819 2038 14826 2048
rect 14878 2082 14885 2090
rect 16082 2082 16089 2092
rect 14878 2048 16089 2082
rect 14878 2038 14885 2048
rect 16082 2040 16089 2048
rect 16141 2082 16148 2092
rect 16141 2048 16861 2082
rect 16141 2040 16148 2048
rect 95 1944 16876 1976
rect 95 1942 16861 1944
rect -126 1856 16861 1860
rect -144 1840 16861 1856
rect -144 1837 5962 1840
rect -144 1836 5596 1837
rect -144 1834 3028 1836
rect -144 1832 2703 1834
rect -144 1780 19 1832
rect 71 1830 2703 1832
rect 71 1829 259 1830
rect 311 1829 799 1830
rect 71 1795 121 1829
rect 155 1795 213 1829
rect 247 1795 259 1829
rect 339 1795 397 1829
rect 431 1795 489 1829
rect 523 1795 581 1829
rect 633 1795 673 1829
rect 707 1795 765 1829
rect 71 1780 259 1795
rect -144 1778 259 1780
rect 311 1778 581 1795
rect -144 1777 581 1778
rect 633 1778 799 1795
rect 851 1829 2703 1830
rect 2755 1829 3028 1834
rect 3080 1829 3296 1836
rect 851 1795 1463 1829
rect 1497 1795 1555 1829
rect 1589 1795 1647 1829
rect 1681 1795 1739 1829
rect 1773 1795 1831 1829
rect 1865 1795 1923 1829
rect 1957 1795 2015 1829
rect 2049 1795 2107 1829
rect 2141 1795 2199 1829
rect 2233 1795 2421 1829
rect 2455 1795 2513 1829
rect 2547 1795 2605 1829
rect 2639 1795 2697 1829
rect 2755 1795 2789 1829
rect 2823 1795 2881 1829
rect 2915 1795 2973 1829
rect 3007 1795 3028 1829
rect 3099 1795 3157 1829
rect 3191 1795 3296 1829
rect 851 1782 2703 1795
rect 2755 1784 3028 1795
rect 3080 1784 3296 1795
rect 3348 1784 3562 1836
rect 3614 1834 5596 1836
rect 3614 1784 3802 1834
rect 2755 1782 3802 1784
rect 3854 1829 5596 1834
rect 3854 1795 3855 1829
rect 3889 1795 3947 1829
rect 3981 1795 4039 1829
rect 4073 1795 4131 1829
rect 4165 1795 4223 1829
rect 4257 1795 4315 1829
rect 4349 1795 4407 1829
rect 4441 1795 4499 1829
rect 4533 1795 4591 1829
rect 4625 1795 4813 1829
rect 4847 1795 4905 1829
rect 4939 1795 4997 1829
rect 5031 1795 5089 1829
rect 5123 1795 5181 1829
rect 5215 1795 5273 1829
rect 5307 1795 5365 1829
rect 5399 1795 5457 1829
rect 5491 1795 5549 1829
rect 5583 1795 5596 1829
rect 3854 1785 5596 1795
rect 5648 1788 5962 1837
rect 6014 1788 6206 1840
rect 6258 1838 16861 1840
rect 6258 1833 9030 1838
rect 6258 1831 8572 1833
rect 6258 1829 6629 1831
rect 6681 1829 8572 1831
rect 6279 1795 6337 1829
rect 6371 1795 6429 1829
rect 6463 1795 6521 1829
rect 6555 1795 6613 1829
rect 6681 1795 6705 1829
rect 6739 1795 6797 1829
rect 6831 1795 6889 1829
rect 6923 1795 6981 1829
rect 7015 1795 7205 1829
rect 7239 1795 7297 1829
rect 7331 1795 7389 1829
rect 7423 1795 7481 1829
rect 7515 1795 7573 1829
rect 7607 1795 7665 1829
rect 7699 1795 7757 1829
rect 7791 1795 7849 1829
rect 7883 1795 7941 1829
rect 7975 1795 8572 1829
rect 6258 1788 6629 1795
rect 5648 1785 6629 1788
rect 3854 1782 6629 1785
rect 851 1779 6629 1782
rect 6681 1781 8572 1795
rect 8624 1830 9030 1833
rect 8624 1829 8824 1830
rect 8876 1829 9030 1830
rect 9082 1836 16861 1838
rect 9082 1834 11653 1836
rect 9082 1833 11443 1834
rect 9082 1832 9611 1833
rect 9082 1829 9313 1832
rect 9365 1829 9611 1832
rect 9663 1829 11443 1833
rect 11495 1829 11653 1834
rect 11705 1834 16861 1836
rect 11705 1829 12004 1834
rect 12056 1829 12284 1834
rect 12336 1833 15547 1834
rect 12336 1829 12601 1833
rect 12653 1831 15547 1833
rect 12653 1829 14391 1831
rect 14443 1829 14686 1831
rect 14738 1829 14973 1831
rect 8624 1795 8639 1829
rect 8673 1795 8731 1829
rect 8765 1795 8823 1829
rect 8876 1795 8915 1829
rect 8949 1795 9007 1829
rect 9082 1795 9099 1829
rect 9133 1795 9191 1829
rect 9225 1795 9283 1829
rect 9365 1795 9375 1829
rect 9409 1795 9597 1829
rect 9663 1795 9689 1829
rect 9723 1795 9781 1829
rect 9815 1795 9873 1829
rect 9907 1795 9965 1829
rect 9999 1795 10057 1829
rect 10091 1795 10149 1829
rect 10183 1795 10241 1829
rect 10275 1795 10333 1829
rect 10367 1795 11031 1829
rect 11065 1795 11123 1829
rect 11157 1795 11215 1829
rect 11249 1795 11307 1829
rect 11341 1795 11399 1829
rect 11433 1795 11443 1829
rect 11525 1795 11583 1829
rect 11617 1795 11653 1829
rect 11709 1795 11767 1829
rect 11801 1795 11989 1829
rect 12056 1795 12081 1829
rect 12115 1795 12173 1829
rect 12207 1795 12265 1829
rect 12336 1795 12357 1829
rect 12391 1795 12449 1829
rect 12483 1795 12541 1829
rect 12575 1795 12601 1829
rect 12667 1795 12725 1829
rect 12759 1795 13421 1829
rect 13455 1795 13513 1829
rect 13547 1795 13605 1829
rect 13639 1795 13697 1829
rect 13731 1795 13789 1829
rect 13823 1795 13881 1829
rect 13915 1795 13973 1829
rect 14007 1795 14065 1829
rect 14099 1795 14157 1829
rect 14191 1795 14381 1829
rect 14443 1795 14473 1829
rect 14507 1795 14565 1829
rect 14599 1795 14657 1829
rect 14738 1795 14749 1829
rect 14783 1795 14841 1829
rect 14875 1795 14933 1829
rect 14967 1795 14973 1829
rect 8624 1781 8824 1795
rect 6681 1779 8824 1781
rect 851 1778 8824 1779
rect 8876 1786 9030 1795
rect 9082 1786 9313 1795
rect 8876 1780 9313 1786
rect 9365 1781 9611 1795
rect 9663 1782 11443 1795
rect 11495 1784 11653 1795
rect 11705 1784 12004 1795
rect 11495 1782 12004 1784
rect 12056 1782 12284 1795
rect 12336 1782 12601 1795
rect 9663 1781 12601 1782
rect 12653 1781 14391 1795
rect 9365 1780 14391 1781
rect 8876 1779 14391 1780
rect 14443 1779 14686 1795
rect 14738 1779 14973 1795
rect 15025 1829 15263 1831
rect 15059 1795 15117 1829
rect 15151 1795 15263 1829
rect 15025 1779 15263 1795
rect 15315 1782 15547 1831
rect 15599 1829 16861 1834
rect 15599 1795 15815 1829
rect 15849 1795 15907 1829
rect 15941 1795 15999 1829
rect 16033 1795 16091 1829
rect 16125 1795 16183 1829
rect 16217 1795 16275 1829
rect 16309 1795 16367 1829
rect 16401 1795 16459 1829
rect 16493 1795 16551 1829
rect 16585 1795 16861 1829
rect 15599 1782 16861 1795
rect 15315 1779 16861 1782
rect 8876 1778 16861 1779
rect 633 1777 16861 1778
rect -144 1770 16861 1777
rect -126 1764 16861 1770
rect 468 1565 475 1617
rect 527 1565 534 1617
rect 641 1591 710 1608
rect 1551 1591 1557 1603
rect 641 1557 656 1591
rect 690 1557 1557 1591
rect 641 1542 710 1557
rect 1551 1550 1557 1557
rect 1609 1550 1616 1603
rect 1730 1565 1737 1617
rect 1789 1565 1796 1617
rect 2861 1564 2868 1616
rect 2920 1564 2927 1616
rect 3033 1590 3103 1611
rect 3943 1590 3949 1602
rect 1551 1549 1616 1550
rect 3033 1556 3048 1590
rect 3082 1556 3949 1590
rect 3033 1541 3103 1556
rect 3943 1549 3949 1556
rect 4001 1549 4008 1602
rect 4122 1565 4129 1617
rect 4181 1565 4188 1617
rect 5253 1564 5260 1616
rect 5312 1564 5319 1616
rect 5424 1602 5488 1605
rect 5424 1591 5489 1602
rect 3943 1548 4008 1549
rect 5424 1557 5439 1591
rect 5473 1590 5489 1591
rect 6333 1590 6339 1602
rect 5473 1559 6339 1590
rect 5473 1557 5489 1559
rect 5424 1548 5489 1557
rect 6333 1549 6339 1559
rect 6391 1549 6398 1602
rect 6513 1566 6520 1618
rect 6572 1566 6579 1618
rect 7645 1565 7652 1617
rect 7704 1565 7711 1617
rect 7817 1591 7884 1604
rect 8727 1591 8733 1603
rect 6333 1548 6398 1549
rect 7817 1557 7832 1591
rect 7866 1558 8733 1591
rect 7866 1557 7884 1558
rect 5424 1546 5488 1548
rect 7817 1543 7884 1557
rect 8727 1550 8733 1558
rect 8785 1550 8792 1603
rect 8906 1566 8913 1618
rect 8965 1566 8972 1618
rect 10036 1564 10043 1616
rect 10095 1564 10102 1616
rect 10208 1592 10270 1607
rect 8727 1549 8792 1550
rect 10208 1558 10223 1592
rect 10257 1591 10270 1592
rect 11119 1591 11125 1602
rect 10257 1559 11125 1591
rect 10257 1558 10270 1559
rect 10208 1544 10270 1558
rect 11119 1549 11125 1559
rect 11177 1549 11184 1602
rect 11299 1566 11306 1618
rect 11358 1566 11365 1618
rect 12428 1563 12435 1615
rect 12487 1563 12494 1615
rect 12600 1593 12658 1604
rect 13508 1593 13514 1602
rect 12600 1592 13514 1593
rect 11119 1548 11184 1549
rect 12600 1558 12615 1592
rect 12649 1559 13514 1592
rect 12649 1558 12658 1559
rect 12600 1546 12658 1558
rect 13508 1549 13514 1559
rect 13566 1549 13573 1602
rect 13688 1566 13695 1618
rect 13747 1566 13754 1618
rect 14820 1564 14827 1616
rect 14879 1564 14886 1616
rect 14996 1592 15048 1598
rect 15903 1592 15909 1603
rect 14996 1558 15008 1592
rect 15042 1558 15909 1592
rect 14996 1552 15048 1558
rect 15903 1550 15909 1558
rect 15961 1550 15968 1603
rect 16083 1566 16090 1618
rect 16142 1566 16149 1618
rect 15903 1549 15968 1550
rect 13508 1548 13573 1549
rect 17 1414 71 1420
rect 17 1362 18 1414
rect 70 1362 71 1414
rect 349 1400 356 1452
rect 408 1448 414 1452
rect 1950 1448 1957 1453
rect 408 1406 1957 1448
rect 408 1400 414 1406
rect 1950 1401 1957 1406
rect 2009 1401 2015 1453
rect 2409 1414 2463 1420
rect 2188 1362 2194 1414
rect 2246 1362 2254 1414
rect 2409 1362 2410 1414
rect 2462 1362 2463 1414
rect 2741 1400 2748 1452
rect 2800 1448 2806 1452
rect 4342 1448 4349 1453
rect 2800 1406 4349 1448
rect 2800 1400 2806 1406
rect 4342 1401 4349 1406
rect 4401 1401 4407 1453
rect 4801 1414 4855 1420
rect 4582 1362 4588 1414
rect 4640 1362 4648 1414
rect 4801 1362 4802 1414
rect 4854 1362 4855 1414
rect 5132 1401 5139 1453
rect 5191 1449 5197 1453
rect 6733 1449 6740 1454
rect 5191 1407 6740 1449
rect 5191 1401 5197 1407
rect 6733 1402 6740 1407
rect 6792 1402 6798 1454
rect 6972 1364 6978 1416
rect 7030 1364 7038 1416
rect 7193 1414 7247 1420
rect 17 1356 71 1362
rect 2409 1356 2463 1362
rect 4801 1356 4855 1362
rect 7193 1362 7194 1414
rect 7246 1362 7247 1414
rect 7525 1400 7532 1452
rect 7584 1448 7590 1452
rect 9126 1448 9133 1453
rect 7584 1406 9133 1448
rect 7584 1400 7590 1406
rect 9126 1401 9133 1406
rect 9185 1401 9191 1453
rect 9584 1415 9638 1421
rect 9364 1362 9370 1414
rect 9422 1362 9430 1414
rect 9584 1363 9585 1415
rect 9637 1363 9638 1415
rect 9917 1401 9924 1453
rect 9976 1449 9982 1453
rect 11518 1449 11525 1454
rect 9976 1407 11525 1449
rect 9976 1401 9982 1407
rect 11518 1402 11525 1407
rect 11577 1402 11583 1454
rect 11756 1364 11762 1416
rect 11814 1364 11822 1416
rect 11976 1414 12030 1420
rect 7193 1356 7247 1362
rect 9584 1357 9638 1363
rect 11976 1362 11977 1414
rect 12029 1362 12030 1414
rect 12309 1401 12316 1453
rect 12368 1449 12374 1453
rect 13910 1449 13917 1454
rect 12368 1407 13917 1449
rect 12368 1401 12374 1407
rect 13910 1402 13917 1407
rect 13969 1402 13975 1454
rect 14369 1415 14423 1421
rect 14148 1362 14154 1414
rect 14206 1362 14214 1414
rect 14369 1363 14370 1415
rect 14422 1363 14423 1415
rect 14704 1401 14711 1453
rect 14763 1449 14769 1453
rect 16305 1449 16312 1454
rect 14763 1407 16312 1449
rect 14763 1401 14769 1407
rect 16305 1402 16312 1407
rect 16364 1402 16370 1454
rect 16540 1364 16546 1416
rect 16598 1364 16606 1416
rect 11976 1356 12030 1362
rect 14369 1357 14423 1363
rect 16175 1316 16205 1362
rect -126 1314 16861 1316
rect -126 1301 16876 1314
rect -126 1299 10510 1301
rect -126 1297 7858 1299
rect -126 1294 7668 1297
rect -126 1285 1210 1294
rect -126 1251 29 1285
rect 63 1251 121 1285
rect 155 1251 213 1285
rect 247 1251 305 1285
rect 339 1251 397 1285
rect 431 1251 489 1285
rect 523 1251 581 1285
rect 615 1251 673 1285
rect 707 1251 765 1285
rect 799 1251 1210 1285
rect -126 1242 1210 1251
rect 1262 1242 1427 1294
rect 1479 1285 1646 1294
rect 1698 1290 5044 1294
rect 1698 1285 1859 1290
rect 1911 1285 2070 1290
rect 2122 1285 4194 1290
rect 4246 1289 5044 1290
rect 4246 1285 4472 1289
rect 4524 1285 5044 1289
rect 5096 1285 5283 1294
rect 5335 1292 7668 1294
rect 5335 1285 7441 1292
rect 7493 1285 7668 1292
rect 7720 1285 7858 1297
rect 7910 1296 10510 1299
rect 7910 1293 10284 1296
rect 7910 1290 10055 1293
rect 7910 1285 8074 1290
rect 1497 1251 1555 1285
rect 1589 1251 1646 1285
rect 1698 1251 1739 1285
rect 1773 1251 1831 1285
rect 1911 1251 1923 1285
rect 1957 1251 2015 1285
rect 2049 1251 2070 1285
rect 2141 1251 2199 1285
rect 2233 1251 2421 1285
rect 2455 1251 2513 1285
rect 2547 1251 2605 1285
rect 2639 1251 2697 1285
rect 2731 1251 2789 1285
rect 2823 1251 2881 1285
rect 2915 1251 2973 1285
rect 3007 1251 3065 1285
rect 3099 1251 3157 1285
rect 3191 1251 3855 1285
rect 3889 1251 3947 1285
rect 3981 1251 4039 1285
rect 4073 1251 4131 1285
rect 4165 1251 4194 1285
rect 4257 1251 4315 1285
rect 4349 1251 4407 1285
rect 4441 1251 4472 1285
rect 4533 1251 4591 1285
rect 4625 1251 4813 1285
rect 4847 1251 4905 1285
rect 4939 1251 4997 1285
rect 5031 1251 5044 1285
rect 5123 1251 5181 1285
rect 5215 1251 5273 1285
rect 5335 1251 5365 1285
rect 5399 1251 5457 1285
rect 5491 1251 5549 1285
rect 5583 1251 6245 1285
rect 6279 1251 6337 1285
rect 6371 1251 6429 1285
rect 6463 1251 6521 1285
rect 6555 1251 6613 1285
rect 6647 1251 6705 1285
rect 6739 1251 6797 1285
rect 6831 1251 6889 1285
rect 6923 1251 6981 1285
rect 7015 1251 7205 1285
rect 7239 1251 7297 1285
rect 7331 1251 7389 1285
rect 7423 1251 7441 1285
rect 7515 1251 7573 1285
rect 7607 1251 7665 1285
rect 7720 1251 7757 1285
rect 7791 1251 7849 1285
rect 7910 1251 7941 1285
rect 7975 1251 8074 1285
rect 1479 1242 1646 1251
rect 1698 1242 1859 1251
rect -126 1238 1859 1242
rect 1911 1238 2070 1251
rect 2122 1238 4194 1251
rect 4246 1238 4472 1251
rect -126 1237 4472 1238
rect 4524 1242 5044 1251
rect 5096 1242 5283 1251
rect 5335 1242 7441 1251
rect 4524 1240 7441 1242
rect 7493 1245 7668 1251
rect 7720 1247 7858 1251
rect 7910 1247 8074 1251
rect 7720 1245 8074 1247
rect 7493 1240 8074 1245
rect 4524 1238 8074 1240
rect 8126 1285 10055 1290
rect 10107 1285 10284 1293
rect 10336 1285 10510 1296
rect 8126 1251 8639 1285
rect 8673 1251 8731 1285
rect 8765 1251 8823 1285
rect 8857 1251 8915 1285
rect 8949 1251 9007 1285
rect 9041 1251 9099 1285
rect 9133 1251 9191 1285
rect 9225 1251 9283 1285
rect 9317 1251 9375 1285
rect 9409 1251 9597 1285
rect 9631 1251 9689 1285
rect 9723 1251 9781 1285
rect 9815 1251 9873 1285
rect 9907 1251 9965 1285
rect 9999 1251 10055 1285
rect 10107 1251 10149 1285
rect 10183 1251 10241 1285
rect 10275 1251 10284 1285
rect 10367 1251 10510 1285
rect 8126 1241 10055 1251
rect 10107 1244 10284 1251
rect 10336 1249 10510 1251
rect 10562 1299 16876 1301
rect 10562 1293 10974 1299
rect 10562 1249 10738 1293
rect 10336 1244 10738 1249
rect 10107 1241 10738 1244
rect 10790 1247 10974 1293
rect 11026 1298 16876 1299
rect 11026 1295 16022 1298
rect 11026 1290 13105 1295
rect 11026 1285 11166 1290
rect 11218 1285 12901 1290
rect 11026 1251 11031 1285
rect 11065 1251 11123 1285
rect 11157 1251 11166 1285
rect 11249 1251 11307 1285
rect 11341 1251 11399 1285
rect 11433 1251 11491 1285
rect 11525 1251 11583 1285
rect 11617 1251 11675 1285
rect 11709 1251 11767 1285
rect 11801 1251 11989 1285
rect 12023 1251 12081 1285
rect 12115 1251 12173 1285
rect 12207 1251 12265 1285
rect 12299 1251 12357 1285
rect 12391 1251 12449 1285
rect 12483 1251 12541 1285
rect 12575 1251 12633 1285
rect 12667 1251 12725 1285
rect 12759 1251 12901 1285
rect 11026 1247 11166 1251
rect 10790 1241 11166 1247
rect 8126 1238 11166 1241
rect 11218 1238 12901 1251
rect 12953 1243 13105 1290
rect 13157 1294 16022 1295
rect 13157 1290 15828 1294
rect 13157 1243 13296 1290
rect 12953 1238 13296 1243
rect 13348 1289 13788 1290
rect 13348 1285 13498 1289
rect 13550 1285 13788 1289
rect 13840 1289 15828 1290
rect 13840 1285 14073 1289
rect 14125 1285 15828 1289
rect 15880 1285 16022 1294
rect 16074 1297 16876 1298
rect 16074 1295 16434 1297
rect 16074 1285 16211 1295
rect 16263 1285 16434 1295
rect 16486 1285 16876 1297
rect 13348 1251 13421 1285
rect 13455 1251 13498 1285
rect 13550 1251 13605 1285
rect 13639 1251 13697 1285
rect 13731 1251 13788 1285
rect 13840 1251 13881 1285
rect 13915 1251 13973 1285
rect 14007 1251 14065 1285
rect 14125 1251 14157 1285
rect 14191 1251 14381 1285
rect 14415 1251 14473 1285
rect 14507 1251 14565 1285
rect 14599 1251 14657 1285
rect 14691 1251 14749 1285
rect 14783 1251 14841 1285
rect 14875 1251 14933 1285
rect 14967 1251 15025 1285
rect 15059 1251 15117 1285
rect 15151 1251 15815 1285
rect 15880 1251 15907 1285
rect 15941 1251 15999 1285
rect 16074 1251 16091 1285
rect 16125 1251 16183 1285
rect 16263 1251 16275 1285
rect 16309 1251 16367 1285
rect 16401 1251 16434 1285
rect 16493 1251 16551 1285
rect 16585 1251 16876 1285
rect 13348 1238 13498 1251
rect 4524 1237 13498 1238
rect 13550 1238 13788 1251
rect 13840 1238 14073 1251
rect 13550 1237 14073 1238
rect 14125 1242 15828 1251
rect 15880 1246 16022 1251
rect 16074 1246 16211 1251
rect 15880 1243 16211 1246
rect 16263 1245 16434 1251
rect 16486 1245 16876 1251
rect 16263 1243 16876 1245
rect 15880 1242 16876 1243
rect 14125 1237 16876 1242
rect -126 1228 16876 1237
rect -126 1220 16861 1228
rect 16237 1172 16303 1173
rect -126 1164 16782 1172
rect -144 1151 16782 1164
rect -144 1150 8753 1151
rect -144 1149 3262 1150
rect -144 1141 265 1149
rect 317 1146 3262 1149
rect 317 1145 2654 1146
rect 317 1141 467 1145
rect 519 1143 2654 1145
rect 519 1142 885 1143
rect 519 1141 656 1142
rect 708 1141 885 1142
rect 937 1141 2654 1143
rect 2706 1143 3262 1146
rect 2706 1141 2869 1143
rect 2921 1141 3262 1143
rect 3314 1149 8753 1150
rect 3314 1148 8563 1149
rect 3314 1141 3542 1148
rect 3594 1147 8563 1148
rect 3594 1146 6518 1147
rect 3594 1141 3761 1146
rect 3813 1145 6518 1146
rect 3813 1143 6327 1145
rect 3813 1141 5582 1143
rect 5634 1141 6327 1143
rect 6379 1141 6518 1145
rect 6570 1141 8563 1147
rect 8615 1141 8753 1149
rect 8805 1150 16782 1151
rect 8805 1149 14613 1150
rect 8805 1141 8947 1149
rect 8999 1145 14613 1149
rect 8999 1141 9258 1145
rect 9310 1144 14613 1145
rect 9310 1141 11441 1144
rect 11493 1141 11645 1144
rect 11697 1142 14613 1144
rect 11697 1141 12449 1142
rect 12501 1141 12653 1142
rect 12705 1141 14613 1142
rect 14665 1148 15542 1150
rect 14665 1141 14846 1148
rect 14898 1146 15262 1148
rect 14898 1141 15053 1146
rect 15105 1141 15262 1146
rect 15314 1141 15542 1148
rect 15594 1141 16782 1150
rect -144 1107 29 1141
rect 63 1107 121 1141
rect 155 1107 213 1141
rect 247 1107 265 1141
rect 339 1107 397 1141
rect 431 1107 467 1141
rect 523 1107 581 1141
rect 615 1107 656 1141
rect 708 1107 765 1141
rect 799 1107 857 1141
rect 937 1107 949 1141
rect 983 1107 1041 1141
rect 1075 1107 1133 1141
rect 1167 1107 1225 1141
rect 1259 1107 1317 1141
rect 1351 1107 1409 1141
rect 1443 1107 1501 1141
rect 1535 1107 1593 1141
rect 1627 1107 1685 1141
rect 1719 1107 1777 1141
rect 1811 1107 1869 1141
rect 1903 1107 1961 1141
rect 1995 1107 2053 1141
rect 2087 1107 2145 1141
rect 2179 1107 2237 1141
rect 2271 1107 2329 1141
rect 2363 1107 2421 1141
rect 2455 1107 2513 1141
rect 2547 1107 2605 1141
rect 2639 1107 2654 1141
rect 2731 1107 2789 1141
rect 2823 1107 2869 1141
rect 2921 1107 2973 1141
rect 3007 1107 3065 1141
rect 3099 1140 3157 1141
rect 3119 1107 3157 1140
rect 3191 1107 3249 1141
rect 3314 1107 3341 1141
rect 3375 1107 3433 1141
rect 3467 1107 3525 1141
rect 3594 1107 3617 1141
rect 3651 1107 3709 1141
rect 3743 1107 3761 1141
rect 3835 1107 3893 1141
rect 3927 1107 3985 1141
rect 4019 1107 4077 1141
rect 4111 1107 4169 1141
rect 4203 1107 4261 1141
rect 4295 1107 4353 1141
rect 4387 1107 4445 1141
rect 4479 1107 4537 1141
rect 4571 1107 4629 1141
rect 4663 1107 4721 1141
rect 4755 1107 4813 1141
rect 4847 1107 4905 1141
rect 4939 1107 4997 1141
rect 5031 1107 5089 1141
rect 5123 1107 5181 1141
rect 5215 1107 5273 1141
rect 5307 1107 5365 1141
rect 5399 1107 5457 1141
rect 5491 1107 5549 1141
rect 5634 1107 5641 1141
rect 5675 1107 5733 1141
rect 5767 1107 5825 1141
rect 5859 1107 5917 1141
rect 5951 1140 6009 1141
rect 5985 1107 6009 1140
rect 6043 1107 6101 1141
rect 6135 1138 6193 1141
rect 6174 1107 6193 1138
rect 6227 1107 6285 1141
rect 6319 1107 6327 1141
rect 6411 1107 6469 1141
rect 6503 1107 6518 1141
rect 6595 1107 6653 1141
rect 6687 1107 6745 1141
rect 6779 1107 6837 1141
rect 6871 1107 6929 1141
rect 6963 1107 7021 1141
rect 7055 1107 7113 1141
rect 7147 1107 7205 1141
rect 7239 1107 7297 1141
rect 7331 1107 7389 1141
rect 7423 1107 7481 1141
rect 7515 1107 7573 1141
rect 7607 1107 7665 1141
rect 7699 1107 7757 1141
rect 7791 1107 7849 1141
rect 7883 1107 7941 1141
rect 7975 1107 8033 1141
rect 8067 1107 8125 1141
rect 8159 1107 8217 1141
rect 8251 1107 8309 1141
rect 8343 1107 8401 1141
rect 8435 1107 8493 1141
rect 8527 1107 8563 1141
rect 8619 1107 8677 1141
rect 8711 1107 8753 1141
rect 8805 1107 8861 1141
rect 8895 1107 8947 1141
rect 8999 1107 9045 1141
rect 9079 1107 9137 1141
rect 9171 1107 9229 1141
rect 9310 1107 9321 1141
rect 9355 1107 9413 1141
rect 9447 1107 9505 1141
rect 9539 1107 9597 1141
rect 9631 1107 9689 1141
rect 9723 1107 9781 1141
rect 9815 1107 9873 1141
rect 9907 1107 9965 1141
rect 9999 1107 10057 1141
rect 10091 1107 10149 1141
rect 10183 1107 10241 1141
rect 10275 1107 10333 1141
rect 10367 1107 10425 1141
rect 10459 1107 10517 1141
rect 10551 1107 10609 1141
rect 10643 1107 10701 1141
rect 10735 1107 10793 1141
rect 10827 1107 10885 1141
rect 10919 1107 10977 1141
rect 11011 1107 11069 1141
rect 11103 1107 11161 1141
rect 11195 1107 11253 1141
rect 11287 1107 11345 1141
rect 11379 1107 11437 1141
rect 11493 1107 11529 1141
rect 11563 1107 11621 1141
rect 11697 1107 11713 1141
rect 11747 1107 11805 1141
rect 11839 1107 11897 1141
rect 11931 1107 11989 1141
rect 12023 1107 12081 1141
rect 12115 1107 12173 1141
rect 12207 1140 12265 1141
rect 12207 1107 12210 1140
rect -144 1097 265 1107
rect 317 1097 467 1107
rect -144 1093 467 1097
rect 519 1093 656 1107
rect -144 1090 656 1093
rect 708 1091 885 1107
rect 937 1094 2654 1107
rect 2706 1094 2869 1107
rect 937 1091 2869 1094
rect 2921 1091 3067 1107
rect 708 1090 3067 1091
rect -144 1088 3067 1090
rect 3119 1098 3262 1107
rect 3314 1098 3542 1107
rect 3119 1096 3542 1098
rect 3594 1096 3761 1107
rect 3119 1094 3761 1096
rect 3813 1094 5582 1107
rect 3119 1091 5582 1094
rect 5634 1091 5933 1107
rect 3119 1088 5933 1091
rect 5985 1088 6122 1107
rect -144 1086 6122 1088
rect 6174 1093 6327 1107
rect 6379 1095 6518 1107
rect 6570 1097 8563 1107
rect 8615 1099 8753 1107
rect 8805 1099 8947 1107
rect 8615 1097 8947 1099
rect 8999 1097 9258 1107
rect 6570 1095 9258 1097
rect 6379 1093 9258 1095
rect 9310 1093 11441 1107
rect 6174 1092 11441 1093
rect 11493 1092 11645 1107
rect 11697 1092 12210 1107
rect 6174 1088 12210 1092
rect 12262 1107 12265 1140
rect 12299 1107 12357 1141
rect 12391 1107 12449 1141
rect 12501 1107 12541 1141
rect 12575 1107 12633 1141
rect 12705 1107 12725 1141
rect 12759 1107 12817 1141
rect 12851 1107 12909 1141
rect 12943 1107 13001 1141
rect 13035 1107 13093 1141
rect 13127 1107 13185 1141
rect 13219 1107 13277 1141
rect 13311 1107 13369 1141
rect 13403 1107 13461 1141
rect 13495 1107 13553 1141
rect 13587 1107 13645 1141
rect 13679 1107 13737 1141
rect 13771 1107 13829 1141
rect 13863 1107 13921 1141
rect 13955 1107 14013 1141
rect 14047 1107 14105 1141
rect 14139 1107 14197 1141
rect 14231 1107 14289 1141
rect 14323 1107 14381 1141
rect 14415 1107 14473 1141
rect 14507 1107 14565 1141
rect 14599 1107 14613 1141
rect 14691 1107 14749 1141
rect 14783 1107 14841 1141
rect 14898 1107 14933 1141
rect 14967 1107 15025 1141
rect 15105 1107 15117 1141
rect 15151 1107 15209 1141
rect 15243 1107 15262 1141
rect 15335 1107 15393 1141
rect 15427 1107 15485 1141
rect 15519 1107 15542 1141
rect 15611 1107 15669 1141
rect 15703 1107 15761 1141
rect 15795 1107 15853 1141
rect 15887 1107 15945 1141
rect 15979 1107 16037 1141
rect 16071 1107 16129 1141
rect 16163 1107 16221 1141
rect 16255 1107 16313 1141
rect 16347 1107 16405 1141
rect 16439 1107 16497 1141
rect 16531 1107 16589 1141
rect 16623 1107 16681 1141
rect 16715 1107 16782 1141
rect 12262 1090 12449 1107
rect 12501 1090 12653 1107
rect 12705 1098 14613 1107
rect 14665 1098 14846 1107
rect 12705 1096 14846 1098
rect 14898 1096 15053 1107
rect 12705 1094 15053 1096
rect 15105 1096 15262 1107
rect 15314 1098 15542 1107
rect 15594 1098 16782 1107
rect 15314 1096 16782 1098
rect 15105 1094 16782 1096
rect 12705 1090 16782 1094
rect 12262 1088 16782 1090
rect 6174 1086 16782 1088
rect -144 1078 16782 1086
rect -126 1076 16782 1078
rect 2324 1042 2376 1048
rect 2324 984 2376 990
rect 4716 1042 4768 1048
rect 4716 984 4768 990
rect 7108 1042 7160 1048
rect 7108 984 7160 990
rect 9500 1042 9552 1048
rect 9500 984 9552 990
rect 11892 1042 11944 1048
rect 11892 984 11944 990
rect 14284 1042 14336 1048
rect 14284 984 14336 990
rect 16676 1042 16728 1048
rect 16676 984 16728 990
rect 201 971 259 977
rect 201 937 213 971
rect 247 968 259 971
rect 477 971 535 977
rect 477 968 489 971
rect 247 940 489 968
rect 247 937 259 940
rect 201 931 259 937
rect 477 937 489 940
rect 523 968 535 971
rect 1213 971 1271 977
rect 2593 971 2651 977
rect 1213 968 1225 971
rect 523 940 1225 968
rect 523 937 535 940
rect 477 931 535 937
rect 1213 937 1225 940
rect 1259 937 1271 971
rect 1213 931 1271 937
rect 2042 965 2094 971
rect 2593 937 2605 971
rect 2639 968 2651 971
rect 2869 971 2927 977
rect 2869 968 2881 971
rect 2639 940 2881 968
rect 2639 937 2651 940
rect 2593 931 2651 937
rect 2869 937 2881 940
rect 2915 968 2927 971
rect 3605 971 3663 977
rect 3605 968 3617 971
rect 2915 940 3617 968
rect 2915 937 2927 940
rect 2869 931 2927 937
rect 3605 937 3617 940
rect 3651 937 3663 971
rect 3605 931 3663 937
rect 4434 966 4486 972
rect 1121 903 1179 909
rect 17 869 71 875
rect 17 817 18 869
rect 70 817 71 869
rect 351 841 357 894
rect 409 841 416 894
rect 1121 869 1133 903
rect 1167 900 1179 903
rect 1759 903 1817 909
rect 2042 907 2094 913
rect 4985 971 5043 977
rect 4985 937 4997 971
rect 5031 968 5043 971
rect 5261 971 5319 977
rect 5261 968 5273 971
rect 5031 940 5273 968
rect 5031 937 5043 940
rect 4985 931 5043 937
rect 5261 937 5273 940
rect 5307 968 5319 971
rect 5997 971 6055 977
rect 5997 968 6009 971
rect 5307 940 6009 968
rect 5307 937 5319 940
rect 5261 931 5319 937
rect 5997 937 6009 940
rect 6043 937 6055 971
rect 5997 931 6055 937
rect 6825 966 6877 972
rect 1759 900 1771 903
rect 1167 872 1771 900
rect 1167 869 1179 872
rect 1121 863 1179 869
rect 1759 869 1771 872
rect 1805 869 1817 903
rect 3513 903 3571 909
rect 1759 863 1817 869
rect 2409 869 2463 875
rect 351 840 416 841
rect 1213 835 1271 841
rect 1213 832 1225 835
rect 17 811 71 817
rect 584 804 1225 832
rect 584 773 627 804
rect 1213 801 1225 804
rect 1259 801 1271 835
rect 2409 817 2410 869
rect 2462 817 2463 869
rect 2743 841 2749 894
rect 2801 841 2808 894
rect 3513 869 3525 903
rect 3559 900 3571 903
rect 4151 903 4209 909
rect 4434 908 4486 914
rect 7377 971 7435 977
rect 7377 937 7389 971
rect 7423 968 7435 971
rect 7653 971 7711 977
rect 7653 968 7665 971
rect 7423 940 7665 968
rect 7423 937 7435 940
rect 7377 931 7435 937
rect 7653 937 7665 940
rect 7699 968 7711 971
rect 8389 971 8447 977
rect 8389 968 8401 971
rect 7699 940 8401 968
rect 7699 937 7711 940
rect 7653 931 7711 937
rect 8389 937 8401 940
rect 8435 937 8447 971
rect 8389 931 8447 937
rect 9218 967 9270 973
rect 4151 900 4163 903
rect 3559 872 4163 900
rect 3559 869 3571 872
rect 3513 863 3571 869
rect 4151 869 4163 872
rect 4197 869 4209 903
rect 5905 903 5963 909
rect 4151 863 4209 869
rect 4801 869 4855 875
rect 2743 840 2808 841
rect 3605 835 3663 841
rect 3605 832 3617 835
rect 2409 811 2463 817
rect 1213 795 1271 801
rect 2976 804 3617 832
rect 110 767 168 773
rect 110 733 122 767
rect 156 764 168 767
rect 569 767 627 773
rect 569 764 581 767
rect 156 736 581 764
rect 156 733 168 736
rect 110 727 168 733
rect 569 733 581 736
rect 615 733 627 767
rect 569 727 627 733
rect 753 767 811 773
rect 753 733 765 767
rect 799 764 811 767
rect 1024 770 1078 776
rect 2976 773 3019 804
rect 3605 801 3617 804
rect 3651 801 3663 835
rect 4801 817 4802 869
rect 4854 817 4855 869
rect 5135 842 5141 895
rect 5193 842 5200 895
rect 5905 869 5917 903
rect 5951 900 5963 903
rect 6543 903 6601 909
rect 6825 908 6877 914
rect 9769 971 9827 977
rect 9769 937 9781 971
rect 9815 968 9827 971
rect 10045 971 10103 977
rect 10045 968 10057 971
rect 9815 940 10057 968
rect 9815 937 9827 940
rect 9769 931 9827 937
rect 10045 937 10057 940
rect 10091 968 10103 971
rect 10781 971 10839 977
rect 10781 968 10793 971
rect 10091 940 10793 968
rect 10091 937 10103 940
rect 10045 931 10103 937
rect 10781 937 10793 940
rect 10827 937 10839 971
rect 10781 931 10839 937
rect 11609 966 11661 972
rect 9218 909 9270 915
rect 12161 971 12219 977
rect 12161 937 12173 971
rect 12207 968 12219 971
rect 12437 971 12495 977
rect 12437 968 12449 971
rect 12207 940 12449 968
rect 12207 937 12219 940
rect 12161 931 12219 937
rect 12437 937 12449 940
rect 12483 968 12495 971
rect 13173 971 13231 977
rect 14553 971 14611 977
rect 13173 968 13185 971
rect 12483 940 13185 968
rect 12483 937 12495 940
rect 12437 931 12495 937
rect 13173 937 13185 940
rect 13219 937 13231 971
rect 13173 931 13231 937
rect 14002 965 14054 971
rect 6543 900 6555 903
rect 5951 872 6555 900
rect 5951 869 5963 872
rect 5905 863 5963 869
rect 6543 869 6555 872
rect 6589 869 6601 903
rect 8297 903 8355 909
rect 6543 863 6601 869
rect 7193 869 7247 875
rect 5135 841 5200 842
rect 5997 835 6055 841
rect 5997 832 6009 835
rect 4801 811 4855 817
rect 3605 795 3663 801
rect 5368 804 6009 832
rect 1024 764 1025 770
rect 799 736 1025 764
rect 799 733 811 736
rect 753 727 811 733
rect 1024 718 1025 736
rect 1077 764 1078 770
rect 1503 767 1561 773
rect 1503 764 1515 767
rect 1077 736 1515 764
rect 1077 718 1078 736
rect 1503 733 1515 736
rect 1549 733 1561 767
rect 1503 727 1561 733
rect 2502 767 2560 773
rect 2502 733 2514 767
rect 2548 764 2560 767
rect 2961 767 3019 773
rect 2961 764 2973 767
rect 2548 736 2973 764
rect 2548 733 2560 736
rect 2502 727 2560 733
rect 2961 733 2973 736
rect 3007 733 3019 767
rect 2961 727 3019 733
rect 3145 767 3203 773
rect 3145 733 3157 767
rect 3191 764 3203 767
rect 3417 770 3471 776
rect 5368 773 5411 804
rect 5997 801 6009 804
rect 6043 801 6055 835
rect 7193 817 7194 869
rect 7246 817 7247 869
rect 7527 842 7533 895
rect 7585 842 7592 895
rect 8297 869 8309 903
rect 8343 900 8355 903
rect 8935 903 8993 909
rect 8935 900 8947 903
rect 8343 872 8947 900
rect 8343 869 8355 872
rect 8297 863 8355 869
rect 8935 869 8947 872
rect 8981 869 8993 903
rect 10689 903 10747 909
rect 8935 863 8993 869
rect 9584 870 9638 876
rect 7527 841 7592 842
rect 8389 835 8447 841
rect 8389 832 8401 835
rect 7193 811 7247 817
rect 5997 795 6055 801
rect 7760 804 8401 832
rect 3417 764 3418 770
rect 3191 736 3418 764
rect 3191 733 3203 736
rect 3145 727 3203 733
rect 1024 712 1078 718
rect 3417 718 3418 736
rect 3470 764 3471 770
rect 3895 767 3953 773
rect 3895 764 3907 767
rect 3470 736 3907 764
rect 3470 718 3471 736
rect 3895 733 3907 736
rect 3941 733 3953 767
rect 3895 727 3953 733
rect 4894 767 4952 773
rect 4894 733 4906 767
rect 4940 764 4952 767
rect 5353 767 5411 773
rect 5353 764 5365 767
rect 4940 736 5365 764
rect 4940 733 4952 736
rect 4894 727 4952 733
rect 5353 733 5365 736
rect 5399 733 5411 767
rect 5353 727 5411 733
rect 5537 767 5595 773
rect 5537 733 5549 767
rect 5583 764 5595 767
rect 5809 770 5863 776
rect 7760 773 7803 804
rect 8389 801 8401 804
rect 8435 801 8447 835
rect 9584 818 9585 870
rect 9637 818 9638 870
rect 9919 841 9925 894
rect 9977 841 9984 894
rect 10689 869 10701 903
rect 10735 900 10747 903
rect 11327 903 11385 909
rect 11609 908 11661 914
rect 14553 937 14565 971
rect 14599 968 14611 971
rect 14829 971 14887 977
rect 14829 968 14841 971
rect 14599 940 14841 968
rect 14599 937 14611 940
rect 14553 931 14611 937
rect 14829 937 14841 940
rect 14875 968 14887 971
rect 15565 971 15623 977
rect 15565 968 15577 971
rect 14875 940 15577 968
rect 14875 937 14887 940
rect 14829 931 14887 937
rect 15565 937 15577 940
rect 15611 937 15623 971
rect 15565 931 15623 937
rect 16395 967 16447 973
rect 11327 900 11339 903
rect 10735 872 11339 900
rect 10735 869 10747 872
rect 10689 863 10747 869
rect 11327 869 11339 872
rect 11373 869 11385 903
rect 13081 903 13139 909
rect 11327 863 11385 869
rect 11976 869 12030 875
rect 9919 840 9984 841
rect 10781 835 10839 841
rect 10781 832 10793 835
rect 9584 812 9638 818
rect 8389 795 8447 801
rect 10152 804 10793 832
rect 5809 764 5810 770
rect 5583 736 5810 764
rect 5583 733 5595 736
rect 5537 727 5595 733
rect 3417 712 3471 718
rect 5809 718 5810 736
rect 5862 764 5863 770
rect 6287 767 6345 773
rect 6287 764 6299 767
rect 5862 736 6299 764
rect 5862 718 5863 736
rect 6287 733 6299 736
rect 6333 733 6345 767
rect 6287 727 6345 733
rect 7286 767 7344 773
rect 7286 733 7298 767
rect 7332 764 7344 767
rect 7745 767 7803 773
rect 7745 764 7757 767
rect 7332 736 7757 764
rect 7332 733 7344 736
rect 7286 727 7344 733
rect 7745 733 7757 736
rect 7791 733 7803 767
rect 7745 727 7803 733
rect 7929 767 7987 773
rect 7929 733 7941 767
rect 7975 764 7987 767
rect 8201 770 8255 776
rect 10152 773 10195 804
rect 10781 801 10793 804
rect 10827 801 10839 835
rect 11976 817 11977 869
rect 12029 817 12030 869
rect 12311 842 12317 895
rect 12369 842 12376 895
rect 13081 869 13093 903
rect 13127 900 13139 903
rect 13719 903 13777 909
rect 14002 907 14054 913
rect 16395 909 16447 915
rect 13719 900 13731 903
rect 13127 872 13731 900
rect 13127 869 13139 872
rect 13081 863 13139 869
rect 13719 869 13731 872
rect 13765 869 13777 903
rect 15473 903 15531 909
rect 13719 863 13777 869
rect 14369 870 14423 876
rect 12311 841 12376 842
rect 13173 835 13231 841
rect 13173 832 13185 835
rect 11976 811 12030 817
rect 10781 795 10839 801
rect 12544 804 13185 832
rect 8201 764 8202 770
rect 7975 736 8202 764
rect 7975 733 7987 736
rect 7929 727 7987 733
rect 5809 712 5863 718
rect 8201 718 8202 736
rect 8254 764 8255 770
rect 8679 767 8737 773
rect 8679 764 8691 767
rect 8254 736 8691 764
rect 8254 718 8255 736
rect 8679 733 8691 736
rect 8725 733 8737 767
rect 8679 727 8737 733
rect 9678 767 9736 773
rect 9678 733 9690 767
rect 9724 764 9736 767
rect 10137 767 10195 773
rect 10137 764 10149 767
rect 9724 736 10149 764
rect 9724 733 9736 736
rect 9678 727 9736 733
rect 10137 733 10149 736
rect 10183 733 10195 767
rect 10137 727 10195 733
rect 10321 767 10379 773
rect 10321 733 10333 767
rect 10367 764 10379 767
rect 10592 770 10646 776
rect 12544 773 12587 804
rect 13173 801 13185 804
rect 13219 801 13231 835
rect 14369 818 14370 870
rect 14422 818 14423 870
rect 14704 841 14710 894
rect 14762 841 14769 894
rect 15473 869 15485 903
rect 15519 900 15531 903
rect 16111 903 16169 909
rect 16111 900 16123 903
rect 15519 872 16123 900
rect 15519 869 15531 872
rect 15473 863 15531 869
rect 16111 869 16123 872
rect 16157 869 16169 903
rect 16111 863 16169 869
rect 14704 840 14769 841
rect 15565 835 15623 841
rect 15565 832 15577 835
rect 14369 812 14423 818
rect 13173 795 13231 801
rect 14936 804 15577 832
rect 10592 764 10593 770
rect 10367 736 10593 764
rect 10367 733 10379 736
rect 10321 727 10379 733
rect 8201 712 8255 718
rect 10592 718 10593 736
rect 10645 764 10646 770
rect 11071 767 11129 773
rect 11071 764 11083 767
rect 10645 736 11083 764
rect 10645 718 10646 736
rect 11071 733 11083 736
rect 11117 733 11129 767
rect 11071 727 11129 733
rect 12070 767 12128 773
rect 12070 733 12082 767
rect 12116 764 12128 767
rect 12529 767 12587 773
rect 12529 764 12541 767
rect 12116 736 12541 764
rect 12116 733 12128 736
rect 12070 727 12128 733
rect 12529 733 12541 736
rect 12575 733 12587 767
rect 12529 727 12587 733
rect 12713 767 12771 773
rect 12713 733 12725 767
rect 12759 764 12771 767
rect 12984 770 13038 776
rect 14936 773 14979 804
rect 15565 801 15577 804
rect 15611 801 15623 835
rect 15565 795 15623 801
rect 12984 764 12985 770
rect 12759 736 12985 764
rect 12759 733 12771 736
rect 12713 727 12771 733
rect 10592 710 10646 718
rect 12984 718 12985 736
rect 13037 764 13038 770
rect 13463 767 13521 773
rect 13463 764 13475 767
rect 13037 736 13475 764
rect 13037 718 13038 736
rect 13463 733 13475 736
rect 13509 733 13521 767
rect 13463 727 13521 733
rect 14462 767 14520 773
rect 14462 733 14474 767
rect 14508 764 14520 767
rect 14921 767 14979 773
rect 14921 764 14933 767
rect 14508 736 14933 764
rect 14508 733 14520 736
rect 14462 727 14520 733
rect 14921 733 14933 736
rect 14967 733 14979 767
rect 14921 727 14979 733
rect 15105 767 15163 773
rect 15105 733 15117 767
rect 15151 764 15163 767
rect 15376 770 15430 776
rect 15376 764 15377 770
rect 15151 736 15377 764
rect 15151 733 15163 736
rect 15105 727 15163 733
rect 12984 712 13038 718
rect 15376 718 15377 736
rect 15429 764 15430 770
rect 15855 767 15913 773
rect 15855 764 15867 767
rect 15429 736 15867 764
rect 15429 718 15430 736
rect 15855 733 15867 736
rect 15901 733 15913 767
rect 15855 727 15913 733
rect 15376 712 15430 718
rect 16816 628 16861 632
rect -126 612 16876 628
rect -126 600 1421 612
rect -126 597 1192 600
rect 1244 597 1421 600
rect 1473 611 16876 612
rect 1473 609 5038 611
rect 1473 606 4708 609
rect 1473 602 1832 606
rect 1473 597 1640 602
rect 1692 597 1832 602
rect 1884 604 4708 606
rect 1884 597 2326 604
rect 2378 603 4708 604
rect 2378 597 4118 603
rect 4170 601 4708 603
rect 4170 597 4511 601
rect 4563 597 4708 601
rect 4760 597 5038 609
rect 5090 597 5234 611
rect 5286 609 8069 611
rect 5286 608 7648 609
rect 5286 604 7442 608
rect 5286 597 7141 604
rect 7193 597 7442 604
rect 7494 597 7648 608
rect 7700 605 8069 609
rect 7700 597 7858 605
rect 7910 597 8069 605
rect -126 563 29 597
rect 63 563 121 597
rect 155 563 213 597
rect 247 563 305 597
rect 339 563 397 597
rect 431 563 489 597
rect 523 563 581 597
rect 615 563 673 597
rect 707 563 765 597
rect 799 563 857 597
rect 891 563 949 597
rect 983 563 1041 597
rect 1075 563 1133 597
rect 1167 563 1192 597
rect 1259 563 1317 597
rect 1351 563 1409 597
rect 1473 563 1501 597
rect 1535 563 1593 597
rect 1627 563 1640 597
rect 1719 563 1777 597
rect 1811 563 1832 597
rect 1903 563 1961 597
rect 1995 563 2053 597
rect 2087 563 2145 597
rect 2179 563 2237 597
rect 2271 563 2326 597
rect 2378 563 2421 597
rect 2455 563 2513 597
rect 2547 563 2605 597
rect 2639 563 2697 597
rect 2731 563 2789 597
rect 2823 563 2881 597
rect 2915 563 2973 597
rect 3007 563 3065 597
rect 3099 563 3157 597
rect 3191 563 3249 597
rect 3283 563 3341 597
rect 3375 563 3433 597
rect 3467 563 3525 597
rect 3559 563 3617 597
rect 3651 563 3709 597
rect 3743 563 3801 597
rect 3835 563 3893 597
rect 3927 563 3985 597
rect 4019 563 4077 597
rect 4111 563 4118 597
rect 4203 563 4261 597
rect 4295 563 4353 597
rect 4387 563 4445 597
rect 4479 563 4511 597
rect 4571 563 4629 597
rect 4663 563 4708 597
rect 4760 563 4813 597
rect 4847 563 4905 597
rect 4939 563 4997 597
rect 5031 563 5038 597
rect 5123 563 5181 597
rect 5215 563 5234 597
rect 5307 563 5365 597
rect 5399 563 5457 597
rect 5491 563 5549 597
rect 5583 563 5641 597
rect 5675 563 5733 597
rect 5767 563 5825 597
rect 5859 563 5917 597
rect 5951 563 6009 597
rect 6043 563 6101 597
rect 6135 563 6193 597
rect 6227 563 6285 597
rect 6319 563 6377 597
rect 6411 563 6469 597
rect 6503 563 6561 597
rect 6595 563 6653 597
rect 6687 563 6745 597
rect 6779 563 6837 597
rect 6871 563 6929 597
rect 6963 563 7021 597
rect 7055 563 7113 597
rect 7193 563 7205 597
rect 7239 563 7297 597
rect 7331 563 7389 597
rect 7423 563 7442 597
rect 7515 563 7573 597
rect 7607 563 7648 597
rect 7700 563 7757 597
rect 7791 563 7849 597
rect 7910 563 7941 597
rect 7975 563 8033 597
rect 8067 563 8069 597
rect -126 548 1192 563
rect 1244 560 1421 563
rect 1473 560 1640 563
rect 1244 550 1640 560
rect 1692 554 1832 563
rect 1884 554 2326 563
rect 1692 552 2326 554
rect 2378 552 4118 563
rect 1692 551 4118 552
rect 4170 551 4511 563
rect 1692 550 4511 551
rect 1244 549 4511 550
rect 4563 557 4708 563
rect 4760 559 5038 563
rect 5090 559 5234 563
rect 5286 559 7141 563
rect 4760 557 7141 559
rect 4563 552 7141 557
rect 7193 556 7442 563
rect 7494 557 7648 563
rect 7700 557 7858 563
rect 7494 556 7858 557
rect 7193 553 7858 556
rect 7910 559 8069 563
rect 8121 608 10968 611
rect 8121 607 10727 608
rect 8121 600 10206 607
rect 8121 597 9949 600
rect 10001 597 10206 600
rect 10258 603 10727 607
rect 10258 597 10456 603
rect 10508 597 10727 603
rect 10779 597 10968 608
rect 11020 610 16876 611
rect 11020 608 16216 610
rect 11020 607 16021 608
rect 11020 597 11193 607
rect 11245 606 16021 607
rect 11245 605 13101 606
rect 11245 597 12900 605
rect 12952 597 13101 605
rect 13153 602 13526 606
rect 13153 597 13319 602
rect 13371 597 13526 602
rect 13578 605 16021 606
rect 13578 597 13731 605
rect 13783 601 15830 605
rect 13783 597 14078 601
rect 14130 597 15830 601
rect 15882 597 16021 605
rect 16073 597 16216 608
rect 16268 605 16876 610
rect 16268 597 16663 605
rect 8121 563 8125 597
rect 8159 563 8217 597
rect 8251 563 8309 597
rect 8343 563 8401 597
rect 8435 563 8493 597
rect 8527 563 8585 597
rect 8619 563 8677 597
rect 8711 563 8769 597
rect 8803 563 8861 597
rect 8895 563 8953 597
rect 8987 563 9045 597
rect 9079 563 9137 597
rect 9171 563 9229 597
rect 9263 563 9321 597
rect 9355 563 9413 597
rect 9447 563 9505 597
rect 9539 563 9597 597
rect 9631 563 9689 597
rect 9723 563 9781 597
rect 9815 563 9873 597
rect 9907 563 9949 597
rect 10001 563 10057 597
rect 10091 563 10149 597
rect 10183 563 10206 597
rect 10275 563 10333 597
rect 10367 563 10425 597
rect 10508 563 10517 597
rect 10551 563 10609 597
rect 10643 563 10701 597
rect 10779 563 10793 597
rect 10827 563 10885 597
rect 10919 563 10968 597
rect 11020 563 11069 597
rect 11103 563 11161 597
rect 11245 563 11253 597
rect 11287 563 11345 597
rect 11379 563 11437 597
rect 11471 563 11529 597
rect 11563 563 11621 597
rect 11655 563 11713 597
rect 11747 563 11805 597
rect 11839 563 11897 597
rect 11931 563 11989 597
rect 12023 563 12081 597
rect 12115 563 12173 597
rect 12207 563 12265 597
rect 12299 563 12357 597
rect 12391 563 12449 597
rect 12483 563 12541 597
rect 12575 563 12633 597
rect 12667 563 12725 597
rect 12759 563 12817 597
rect 12851 563 12900 597
rect 12952 563 13001 597
rect 13035 563 13093 597
rect 13153 563 13185 597
rect 13219 563 13277 597
rect 13311 563 13319 597
rect 13403 563 13461 597
rect 13495 563 13526 597
rect 13587 563 13645 597
rect 13679 563 13731 597
rect 13783 563 13829 597
rect 13863 563 13921 597
rect 13955 563 14013 597
rect 14047 563 14078 597
rect 14139 563 14197 597
rect 14231 563 14289 597
rect 14323 563 14381 597
rect 14415 563 14473 597
rect 14507 563 14565 597
rect 14599 563 14657 597
rect 14691 563 14749 597
rect 14783 563 14841 597
rect 14875 563 14933 597
rect 14967 563 15025 597
rect 15059 563 15117 597
rect 15151 563 15209 597
rect 15243 563 15301 597
rect 15335 563 15393 597
rect 15427 563 15485 597
rect 15519 563 15577 597
rect 15611 563 15669 597
rect 15703 563 15761 597
rect 15795 563 15830 597
rect 15887 563 15945 597
rect 15979 563 16021 597
rect 16073 563 16129 597
rect 16163 563 16216 597
rect 16268 563 16313 597
rect 16347 563 16405 597
rect 16439 563 16497 597
rect 16531 563 16589 597
rect 16623 563 16663 597
rect 8121 559 9949 563
rect 7910 553 9949 559
rect 7193 552 9949 553
rect 4563 549 9949 552
rect 1244 548 9949 549
rect 10001 555 10206 563
rect 10258 555 10456 563
rect 10001 551 10456 555
rect 10508 556 10727 563
rect 10779 559 10968 563
rect 11020 559 11193 563
rect 10779 556 11193 559
rect 10508 555 11193 556
rect 11245 555 12900 563
rect 10508 553 12900 555
rect 12952 554 13101 563
rect 13153 554 13319 563
rect 12952 553 13319 554
rect 10508 551 13319 553
rect 10001 550 13319 551
rect 13371 554 13526 563
rect 13578 554 13731 563
rect 13371 553 13731 554
rect 13783 553 14078 563
rect 13371 550 14078 553
rect 10001 549 14078 550
rect 14130 553 15830 563
rect 15882 556 16021 563
rect 16073 558 16216 563
rect 16268 558 16663 563
rect 16073 556 16663 558
rect 15882 553 16663 556
rect 16715 553 16876 605
rect 14130 549 16876 553
rect 10001 548 16876 549
rect -126 542 16876 548
rect -126 536 16861 542
rect -126 532 16816 536
rect 1591 483 1657 487
rect 3983 483 4049 487
rect 6375 483 6441 487
rect 8767 483 8833 487
rect 11159 483 11225 487
rect 13551 483 13617 487
rect 15943 483 16009 485
rect 16816 483 16861 487
rect -126 476 16861 483
rect -144 464 16861 476
rect -144 461 15022 464
rect -144 459 3786 461
rect -144 456 495 459
rect -144 452 47 456
rect 99 452 495 456
rect 547 457 3786 459
rect 547 456 929 457
rect 547 452 713 456
rect -144 418 29 452
rect 99 418 121 452
rect 155 418 213 452
rect 247 418 280 452
rect 339 418 397 452
rect 431 418 489 452
rect 547 418 581 452
rect 615 418 673 452
rect 707 418 713 452
rect -144 404 47 418
rect 99 404 280 418
rect -144 400 280 404
rect 332 407 495 418
rect 547 407 713 418
rect 332 404 713 407
rect 765 452 929 456
rect 981 456 3786 457
rect 981 453 3050 456
rect 981 452 2650 453
rect 2702 452 2840 453
rect 2892 452 3050 453
rect 3102 453 3562 456
rect 3102 452 3267 453
rect 3319 452 3562 453
rect 799 418 857 452
rect 891 418 929 452
rect 983 418 1041 452
rect 1075 418 1133 452
rect 1167 418 1225 452
rect 1259 418 1317 452
rect 1351 418 1409 452
rect 1443 418 1501 452
rect 1535 418 1593 452
rect 1627 418 1685 452
rect 1719 418 1777 452
rect 1811 418 1869 452
rect 1903 418 1961 452
rect 1995 418 2053 452
rect 2087 418 2145 452
rect 2179 418 2237 452
rect 2271 418 2329 452
rect 2363 418 2421 452
rect 2455 418 2513 452
rect 2547 418 2605 452
rect 2639 418 2650 452
rect 2731 418 2789 452
rect 2823 418 2840 452
rect 2915 418 2973 452
rect 3007 418 3050 452
rect 3102 418 3157 452
rect 3191 418 3249 452
rect 3319 418 3341 452
rect 3375 418 3433 452
rect 3467 418 3525 452
rect 3559 418 3562 452
rect 765 405 929 418
rect 981 405 2650 418
rect 765 404 2650 405
rect 332 401 2650 404
rect 2702 401 2840 418
rect 2892 404 3050 418
rect 3102 404 3267 418
rect 2892 401 3267 404
rect 3319 404 3562 418
rect 3614 452 3786 456
rect 3838 456 6433 461
rect 3838 454 6216 456
rect 3838 452 5664 454
rect 5716 452 6216 454
rect 6268 452 6433 456
rect 6485 458 14390 461
rect 6485 452 6634 458
rect 6686 457 14390 458
rect 6686 452 9529 457
rect 9581 455 14390 457
rect 9581 453 12210 455
rect 9581 452 11430 453
rect 11482 452 11686 453
rect 11738 452 11921 453
rect 11973 452 12210 453
rect 3614 418 3617 452
rect 3651 418 3709 452
rect 3743 418 3786 452
rect 3838 418 3893 452
rect 3927 418 3985 452
rect 4019 418 4077 452
rect 4111 418 4169 452
rect 4203 418 4261 452
rect 4295 418 4353 452
rect 4387 418 4445 452
rect 4479 418 4537 452
rect 4571 418 4629 452
rect 4663 418 4721 452
rect 4755 418 4813 452
rect 4847 418 4905 452
rect 4939 418 4997 452
rect 5031 418 5089 452
rect 5123 418 5181 452
rect 5215 418 5273 452
rect 5307 418 5365 452
rect 5399 418 5457 452
rect 5491 418 5549 452
rect 5583 418 5641 452
rect 5716 418 5733 452
rect 5767 418 5825 452
rect 5859 418 5917 452
rect 5951 418 5964 452
rect 6043 418 6101 452
rect 6135 418 6193 452
rect 6268 418 6285 452
rect 6319 418 6377 452
rect 6411 418 6433 452
rect 6503 418 6561 452
rect 6595 418 6634 452
rect 6687 418 6745 452
rect 6779 418 6837 452
rect 6871 418 6929 452
rect 6963 418 7021 452
rect 7055 418 7113 452
rect 7147 418 7205 452
rect 7239 418 7297 452
rect 7331 418 7389 452
rect 7423 418 7481 452
rect 7515 418 7573 452
rect 7607 418 7665 452
rect 7699 418 7757 452
rect 7791 418 7849 452
rect 7883 418 7941 452
rect 7975 418 8033 452
rect 8067 418 8125 452
rect 8159 418 8217 452
rect 8251 418 8309 452
rect 8343 418 8401 452
rect 8435 418 8493 452
rect 8527 449 8585 452
rect 8571 418 8585 449
rect 8619 418 8677 452
rect 8711 449 8769 452
rect 3614 409 3786 418
rect 3838 409 5664 418
rect 3614 404 5664 409
rect 3319 402 5664 404
rect 5716 402 5964 418
rect 3319 401 5964 402
rect 332 400 5964 401
rect 6016 404 6216 418
rect 6268 409 6433 418
rect 6485 409 6634 418
rect 6268 406 6634 409
rect 6686 406 8519 418
rect 6268 404 8519 406
rect 6016 400 8519 404
rect -144 397 8519 400
rect 8571 397 8711 418
rect 8763 418 8769 449
rect 8803 418 8861 452
rect 8895 449 8953 452
rect 8895 418 8911 449
rect 8987 418 9045 452
rect 9079 418 9137 452
rect 9171 418 9229 452
rect 9263 418 9321 452
rect 9355 418 9413 452
rect 9447 418 9505 452
rect 9581 418 9597 452
rect 9631 418 9689 452
rect 9723 418 9781 452
rect 9815 418 9873 452
rect 9907 418 9965 452
rect 9999 418 10057 452
rect 10091 418 10149 452
rect 10183 418 10241 452
rect 10275 418 10333 452
rect 10367 418 10425 452
rect 10459 418 10517 452
rect 10551 418 10609 452
rect 10643 418 10701 452
rect 10735 418 10793 452
rect 10827 418 10885 452
rect 10919 418 10977 452
rect 11011 418 11069 452
rect 11103 418 11161 452
rect 11195 418 11253 452
rect 11287 418 11345 452
rect 11379 418 11430 452
rect 11482 418 11529 452
rect 11563 418 11621 452
rect 11655 418 11686 452
rect 11747 418 11805 452
rect 11839 418 11897 452
rect 11973 418 11989 452
rect 12023 418 12081 452
rect 12115 418 12173 452
rect 12207 418 12210 452
rect 8763 397 8911 418
rect 8963 405 9529 418
rect 9581 405 11430 418
rect 8963 401 11430 405
rect 11482 401 11686 418
rect 11738 401 11921 418
rect 11973 403 12210 418
rect 12262 453 12604 455
rect 12262 452 12400 453
rect 12452 452 12604 453
rect 12656 452 14390 455
rect 14442 457 15022 461
rect 14442 452 14632 457
rect 14684 456 15022 457
rect 14684 452 14832 456
rect 14884 452 15022 456
rect 15074 462 16861 464
rect 15074 452 15243 462
rect 12262 418 12265 452
rect 12299 418 12357 452
rect 12391 418 12400 452
rect 12483 418 12541 452
rect 12575 418 12604 452
rect 12667 418 12725 452
rect 12759 418 12817 452
rect 12851 418 12909 452
rect 12943 418 13001 452
rect 13035 418 13093 452
rect 13127 418 13185 452
rect 13219 418 13277 452
rect 13311 418 13369 452
rect 13403 418 13461 452
rect 13495 418 13553 452
rect 13587 418 13645 452
rect 13679 418 13737 452
rect 13771 418 13829 452
rect 13863 418 13921 452
rect 13955 418 14013 452
rect 14047 418 14105 452
rect 14139 418 14197 452
rect 14231 418 14289 452
rect 14323 418 14381 452
rect 14442 418 14473 452
rect 14507 418 14565 452
rect 14599 418 14632 452
rect 14691 418 14749 452
rect 14783 418 14832 452
rect 14884 418 14933 452
rect 14967 418 15022 452
rect 15074 418 15117 452
rect 15151 418 15209 452
rect 12262 403 12400 418
rect 11973 401 12400 403
rect 12452 403 12604 418
rect 12656 409 14390 418
rect 14442 409 14632 418
rect 12656 405 14632 409
rect 14684 405 14832 418
rect 12656 404 14832 405
rect 14884 412 15022 418
rect 15074 412 15243 418
rect 14884 410 15243 412
rect 15295 457 16861 462
rect 15295 452 15539 457
rect 15591 452 16861 457
rect 15295 418 15301 452
rect 15335 418 15393 452
rect 15427 418 15485 452
rect 15519 418 15539 452
rect 15611 418 15669 452
rect 15703 418 15761 452
rect 15795 418 15853 452
rect 15887 418 15945 452
rect 15979 418 16037 452
rect 16071 418 16129 452
rect 16163 418 16221 452
rect 16255 418 16313 452
rect 16347 418 16405 452
rect 16439 418 16497 452
rect 16531 418 16589 452
rect 16623 418 16681 452
rect 16715 418 16861 452
rect 15295 410 15539 418
rect 14884 405 15539 410
rect 15591 405 16861 418
rect 14884 404 16861 405
rect 12656 403 16861 404
rect 12452 401 16861 403
rect 8963 397 16861 401
rect -144 391 16861 397
rect -144 390 16816 391
rect -126 387 16816 390
rect 12384 386 12481 387
rect 17 350 69 356
rect 2409 350 2461 356
rect 1019 302 1025 314
rect 17 292 69 298
rect 297 286 349 292
rect 297 228 349 234
rect 508 271 1025 302
rect 508 154 537 271
rect 1019 262 1025 271
rect 1077 262 1083 314
rect 4802 350 4854 356
rect 3411 303 3417 315
rect 2409 292 2461 298
rect 1121 282 1179 288
rect 1121 248 1133 282
rect 1167 279 1179 282
rect 1857 282 1915 288
rect 1857 279 1869 282
rect 1167 251 1869 279
rect 1167 248 1179 251
rect 1121 242 1179 248
rect 1857 248 1869 251
rect 1903 279 1915 282
rect 2133 282 2191 288
rect 2133 279 2145 282
rect 1903 251 2145 279
rect 1903 248 1915 251
rect 1857 242 1915 248
rect 2133 248 2145 251
rect 2179 248 2191 282
rect 2133 242 2191 248
rect 2689 286 2741 292
rect 2689 228 2741 234
rect 2900 272 3417 303
rect 575 214 633 220
rect 575 180 587 214
rect 621 211 633 214
rect 1213 214 1271 220
rect 1213 211 1225 214
rect 621 183 1225 211
rect 621 180 633 183
rect 575 174 633 180
rect 1213 180 1225 183
rect 1259 180 1271 214
rect 1213 174 1271 180
rect 2298 163 2304 215
rect 2358 163 2364 215
rect 490 148 548 154
rect 490 114 502 148
rect 536 114 548 148
rect 490 108 548 114
rect 1121 146 1179 152
rect 1121 112 1133 146
rect 1167 143 1179 146
rect 1167 115 1808 143
rect 1167 112 1179 115
rect 508 107 537 108
rect 1121 106 1179 112
rect 1765 84 1808 115
rect 1953 107 1959 160
rect 2011 107 2018 160
rect 2900 156 2929 272
rect 3411 263 3417 272
rect 3469 263 3475 315
rect 7193 350 7245 356
rect 5803 302 5809 314
rect 4802 292 4854 298
rect 3513 282 3571 288
rect 3513 248 3525 282
rect 3559 279 3571 282
rect 4249 282 4307 288
rect 4249 279 4261 282
rect 3559 251 4261 279
rect 3559 248 3571 251
rect 3513 242 3571 248
rect 4249 248 4261 251
rect 4295 279 4307 282
rect 4525 282 4583 288
rect 4525 279 4537 282
rect 4295 251 4537 279
rect 4295 248 4307 251
rect 4249 242 4307 248
rect 4525 248 4537 251
rect 4571 248 4583 282
rect 4525 242 4583 248
rect 5080 286 5132 292
rect 5080 228 5132 234
rect 5292 271 5809 302
rect 2967 214 3025 220
rect 2967 180 2979 214
rect 3013 211 3025 214
rect 3605 214 3663 220
rect 3605 211 3617 214
rect 3013 183 3617 211
rect 3013 180 3025 183
rect 2967 174 3025 180
rect 3605 180 3617 183
rect 3651 180 3663 214
rect 3605 174 3663 180
rect 4692 163 4698 215
rect 4752 163 4758 215
rect 2879 150 2937 156
rect 2879 116 2891 150
rect 2925 116 2937 150
rect 2879 110 2937 116
rect 3513 146 3571 152
rect 3513 112 3525 146
rect 3559 143 3571 146
rect 3559 115 4200 143
rect 3559 112 3571 115
rect 2900 108 2929 110
rect 1953 106 2018 107
rect 3513 106 3571 112
rect 4157 84 4200 115
rect 4345 107 4351 160
rect 4403 107 4410 160
rect 5292 156 5321 271
rect 5803 262 5809 271
rect 5861 262 5867 314
rect 9585 349 9637 355
rect 8195 302 8201 314
rect 7193 292 7245 298
rect 5905 282 5963 288
rect 5905 248 5917 282
rect 5951 279 5963 282
rect 6641 282 6699 288
rect 6641 279 6653 282
rect 5951 251 6653 279
rect 5951 248 5963 251
rect 5905 242 5963 248
rect 6641 248 6653 251
rect 6687 279 6699 282
rect 6917 282 6975 288
rect 6917 279 6929 282
rect 6687 251 6929 279
rect 6687 248 6699 251
rect 6641 242 6699 248
rect 6917 248 6929 251
rect 6963 248 6975 282
rect 6917 242 6975 248
rect 7473 286 7525 292
rect 7473 228 7525 234
rect 7684 271 8201 302
rect 5359 214 5417 220
rect 5359 180 5371 214
rect 5405 211 5417 214
rect 5997 214 6055 220
rect 5997 211 6009 214
rect 5405 183 6009 211
rect 5405 180 5417 183
rect 5359 174 5417 180
rect 5997 180 6009 183
rect 6043 180 6055 214
rect 5997 174 6055 180
rect 7082 165 7088 217
rect 7142 165 7148 217
rect 6736 160 6801 161
rect 5272 150 5330 156
rect 5272 116 5284 150
rect 5318 116 5330 150
rect 5272 110 5330 116
rect 5905 146 5963 152
rect 5905 112 5917 146
rect 5951 143 5963 146
rect 5951 115 6592 143
rect 5951 112 5963 115
rect 5292 107 5321 110
rect 4345 106 4410 107
rect 5905 106 5963 112
rect 6549 84 6592 115
rect 6736 108 6742 160
rect 6794 108 6801 160
rect 7684 156 7713 271
rect 8195 262 8201 271
rect 8253 262 8259 314
rect 11978 351 12030 357
rect 10587 302 10593 314
rect 9585 291 9637 297
rect 8297 282 8355 288
rect 8297 248 8309 282
rect 8343 279 8355 282
rect 9033 282 9091 288
rect 9033 279 9045 282
rect 8343 251 9045 279
rect 8343 248 8355 251
rect 8297 242 8355 248
rect 9033 248 9045 251
rect 9079 279 9091 282
rect 9309 282 9367 288
rect 9309 279 9321 282
rect 9079 251 9321 279
rect 9079 248 9091 251
rect 9033 242 9091 248
rect 9309 248 9321 251
rect 9355 248 9367 282
rect 9309 242 9367 248
rect 9865 286 9917 292
rect 9865 228 9917 234
rect 10076 271 10593 302
rect 7751 214 7809 220
rect 7751 180 7763 214
rect 7797 211 7809 214
rect 8389 214 8447 220
rect 8389 211 8401 214
rect 7797 183 8401 211
rect 7797 180 7809 183
rect 7751 174 7809 180
rect 8389 180 8401 183
rect 8435 180 8447 214
rect 8389 174 8447 180
rect 9474 163 9480 215
rect 9534 163 9540 215
rect 7665 150 7723 156
rect 7665 116 7677 150
rect 7711 116 7723 150
rect 7665 110 7723 116
rect 8297 146 8355 152
rect 8297 112 8309 146
rect 8343 143 8355 146
rect 8343 115 8984 143
rect 8343 112 8355 115
rect 6736 107 6801 108
rect 7684 107 7713 110
rect 8297 106 8355 112
rect 8941 84 8984 115
rect 9129 107 9135 160
rect 9187 107 9194 160
rect 10076 156 10105 271
rect 10587 262 10593 271
rect 10645 262 10651 314
rect 14369 351 14421 357
rect 12979 303 12985 315
rect 11978 293 12030 299
rect 10689 282 10747 288
rect 10689 248 10701 282
rect 10735 279 10747 282
rect 11425 282 11483 288
rect 11425 279 11437 282
rect 10735 251 11437 279
rect 10735 248 10747 251
rect 10689 242 10747 248
rect 11425 248 11437 251
rect 11471 279 11483 282
rect 11701 282 11759 288
rect 11701 279 11713 282
rect 11471 251 11713 279
rect 11471 248 11483 251
rect 11425 242 11483 248
rect 11701 248 11713 251
rect 11747 248 11759 282
rect 11701 242 11759 248
rect 12256 287 12308 293
rect 12256 229 12308 235
rect 12468 272 12985 303
rect 10143 214 10201 220
rect 10143 180 10155 214
rect 10189 211 10201 214
rect 10781 214 10839 220
rect 10781 211 10793 214
rect 10189 183 10793 211
rect 10189 180 10201 183
rect 10143 174 10201 180
rect 10781 180 10793 183
rect 10827 180 10839 214
rect 10781 174 10839 180
rect 11866 165 11872 217
rect 11926 165 11932 217
rect 10056 150 10114 156
rect 10056 116 10068 150
rect 10102 116 10114 150
rect 10056 110 10114 116
rect 10689 146 10747 152
rect 10689 112 10701 146
rect 10735 143 10747 146
rect 10735 115 11376 143
rect 10735 112 10747 115
rect 10076 107 10105 110
rect 9129 106 9194 107
rect 10689 106 10747 112
rect 11333 84 11376 115
rect 11520 107 11526 160
rect 11578 107 11585 160
rect 12468 156 12497 272
rect 12979 263 12985 272
rect 13037 263 13043 315
rect 15371 303 15377 315
rect 14369 293 14421 299
rect 13081 282 13139 288
rect 13081 248 13093 282
rect 13127 279 13139 282
rect 13817 282 13875 288
rect 13817 279 13829 282
rect 13127 251 13829 279
rect 13127 248 13139 251
rect 13081 242 13139 248
rect 13817 248 13829 251
rect 13863 279 13875 282
rect 14093 282 14151 288
rect 14093 279 14105 282
rect 13863 251 14105 279
rect 13863 248 13875 251
rect 13817 242 13875 248
rect 14093 248 14105 251
rect 14139 248 14151 282
rect 14093 242 14151 248
rect 14649 286 14701 292
rect 14649 228 14701 234
rect 14860 272 15377 303
rect 12535 214 12593 220
rect 12535 180 12547 214
rect 12581 211 12593 214
rect 13173 214 13231 220
rect 13173 211 13185 214
rect 12581 183 13185 211
rect 12581 180 12593 183
rect 12535 174 12593 180
rect 13173 180 13185 183
rect 13219 180 13231 214
rect 13173 174 13231 180
rect 14258 163 14264 215
rect 14318 163 14324 215
rect 12449 150 12507 156
rect 12449 116 12461 150
rect 12495 116 12507 150
rect 12449 110 12507 116
rect 13081 146 13139 152
rect 13081 112 13093 146
rect 13127 143 13139 146
rect 13127 115 13768 143
rect 13127 112 13139 115
rect 12468 108 12497 110
rect 11520 106 11585 107
rect 13081 106 13139 112
rect 13725 84 13768 115
rect 13913 107 13919 160
rect 13971 107 13978 160
rect 14860 156 14889 272
rect 15371 263 15377 272
rect 15429 263 15435 315
rect 15473 282 15531 288
rect 15473 248 15485 282
rect 15519 279 15531 282
rect 16209 282 16267 288
rect 16209 279 16221 282
rect 15519 251 16221 279
rect 15519 248 15531 251
rect 15473 242 15531 248
rect 16209 248 16221 251
rect 16255 279 16267 282
rect 16485 282 16543 288
rect 16485 279 16497 282
rect 16255 251 16497 279
rect 16255 248 16267 251
rect 16209 242 16267 248
rect 16485 248 16497 251
rect 16531 248 16543 282
rect 16485 242 16543 248
rect 14927 214 14985 220
rect 14927 180 14939 214
rect 14973 211 14985 214
rect 15565 214 15623 220
rect 15565 211 15577 214
rect 14973 183 15577 211
rect 14973 180 14985 183
rect 14927 174 14985 180
rect 15565 180 15577 183
rect 15611 180 15623 214
rect 15565 174 15623 180
rect 16650 165 16656 217
rect 16710 165 16716 217
rect 14840 150 14898 156
rect 14840 116 14852 150
rect 14886 116 14898 150
rect 14840 110 14898 116
rect 15473 146 15531 152
rect 15473 112 15485 146
rect 15519 143 15531 146
rect 15519 115 16160 143
rect 15519 112 15531 115
rect 14860 108 14889 110
rect 13913 106 13978 107
rect 15473 106 15531 112
rect 16117 84 16160 115
rect 16306 107 16312 160
rect 16364 107 16371 160
rect 16306 106 16371 107
rect 831 78 889 84
rect 831 44 843 78
rect 877 75 889 78
rect 1581 78 1639 84
rect 1581 75 1593 78
rect 877 47 1593 75
rect 877 44 889 47
rect 831 38 889 44
rect 1581 44 1593 47
rect 1627 44 1639 78
rect 1581 38 1639 44
rect 1765 78 1823 84
rect 1765 44 1777 78
rect 1811 75 1823 78
rect 2224 78 2282 84
rect 2224 75 2236 78
rect 1811 47 2236 75
rect 1811 44 1823 47
rect 1765 38 1823 44
rect 2224 44 2236 47
rect 2270 44 2282 78
rect 2224 38 2282 44
rect 3223 78 3281 84
rect 3223 44 3235 78
rect 3269 75 3281 78
rect 3973 78 4031 84
rect 3973 75 3985 78
rect 3269 47 3985 75
rect 3269 44 3281 47
rect 3223 38 3281 44
rect 3973 44 3985 47
rect 4019 44 4031 78
rect 3973 38 4031 44
rect 4157 78 4215 84
rect 4157 44 4169 78
rect 4203 75 4215 78
rect 4616 78 4674 84
rect 4616 75 4628 78
rect 4203 47 4628 75
rect 4203 44 4215 47
rect 4157 38 4215 44
rect 4616 44 4628 47
rect 4662 44 4674 78
rect 4616 38 4674 44
rect 5615 78 5673 84
rect 5615 44 5627 78
rect 5661 75 5673 78
rect 6365 78 6423 84
rect 6365 75 6377 78
rect 5661 47 6377 75
rect 5661 44 5673 47
rect 5615 38 5673 44
rect 6365 44 6377 47
rect 6411 44 6423 78
rect 6365 38 6423 44
rect 6549 78 6607 84
rect 6549 44 6561 78
rect 6595 75 6607 78
rect 7008 78 7066 84
rect 7008 75 7020 78
rect 6595 47 7020 75
rect 6595 44 6607 47
rect 6549 38 6607 44
rect 7008 44 7020 47
rect 7054 44 7066 78
rect 7008 38 7066 44
rect 8007 78 8065 84
rect 8007 44 8019 78
rect 8053 75 8065 78
rect 8757 78 8815 84
rect 8757 75 8769 78
rect 8053 47 8769 75
rect 8053 44 8065 47
rect 8007 38 8065 44
rect 8757 44 8769 47
rect 8803 44 8815 78
rect 8757 38 8815 44
rect 8941 78 8999 84
rect 8941 44 8953 78
rect 8987 75 8999 78
rect 9400 78 9458 84
rect 9400 75 9412 78
rect 8987 47 9412 75
rect 8987 44 8999 47
rect 8941 38 8999 44
rect 9400 44 9412 47
rect 9446 44 9458 78
rect 9400 38 9458 44
rect 10399 78 10457 84
rect 10399 44 10411 78
rect 10445 75 10457 78
rect 11149 78 11207 84
rect 11149 75 11161 78
rect 10445 47 11161 75
rect 10445 44 10457 47
rect 10399 38 10457 44
rect 11149 44 11161 47
rect 11195 44 11207 78
rect 11149 38 11207 44
rect 11333 78 11391 84
rect 11333 44 11345 78
rect 11379 75 11391 78
rect 11792 78 11850 84
rect 11792 75 11804 78
rect 11379 47 11804 75
rect 11379 44 11391 47
rect 11333 38 11391 44
rect 11792 44 11804 47
rect 11838 44 11850 78
rect 11792 38 11850 44
rect 12791 78 12849 84
rect 12791 44 12803 78
rect 12837 75 12849 78
rect 13541 78 13599 84
rect 13541 75 13553 78
rect 12837 47 13553 75
rect 12837 44 12849 47
rect 12791 38 12849 44
rect 13541 44 13553 47
rect 13587 44 13599 78
rect 13541 38 13599 44
rect 13725 78 13783 84
rect 13725 44 13737 78
rect 13771 75 13783 78
rect 14184 78 14242 84
rect 14184 75 14196 78
rect 13771 47 14196 75
rect 13771 44 13783 47
rect 13725 38 13783 44
rect 14184 44 14196 47
rect 14230 44 14242 78
rect 14184 38 14242 44
rect 15183 78 15241 84
rect 15183 44 15195 78
rect 15229 75 15241 78
rect 15933 78 15991 84
rect 15933 75 15945 78
rect 15229 47 15945 75
rect 15229 44 15241 47
rect 15183 38 15241 44
rect 15933 44 15945 47
rect 15979 44 15991 78
rect 15933 38 15991 44
rect 16117 78 16175 84
rect 16117 44 16129 78
rect 16163 75 16175 78
rect 16576 78 16634 84
rect 16576 75 16588 78
rect 16163 47 16588 75
rect 16163 44 16175 47
rect 16117 38 16175 44
rect 16576 44 16588 47
rect 16622 44 16634 78
rect 16576 38 16634 44
rect 16816 -61 16861 -57
rect -126 -64 16861 -61
rect -126 -74 16876 -64
rect -126 -76 2163 -74
rect -126 -92 421 -76
rect 473 -79 2163 -76
rect 473 -92 620 -79
rect -126 -126 29 -92
rect 63 -126 121 -92
rect 155 -126 213 -92
rect 247 -126 305 -92
rect 339 -126 397 -92
rect 473 -126 489 -92
rect 523 -126 581 -92
rect 615 -126 620 -92
rect -126 -128 421 -126
rect 473 -128 620 -126
rect -126 -131 620 -128
rect 672 -92 831 -79
rect 883 -92 1037 -79
rect 1089 -81 1739 -79
rect 1089 -92 1265 -81
rect 672 -126 673 -92
rect 707 -126 765 -92
rect 799 -126 831 -92
rect 891 -126 949 -92
rect 983 -126 1037 -92
rect 1089 -126 1133 -92
rect 1167 -126 1225 -92
rect 1259 -126 1265 -92
rect 672 -131 831 -126
rect 883 -131 1037 -126
rect 1089 -131 1265 -126
rect -126 -133 1265 -131
rect 1317 -92 1509 -81
rect 1561 -92 1739 -81
rect 1791 -92 1945 -79
rect 1997 -92 2163 -79
rect 2215 -77 16876 -74
rect 2215 -80 2574 -77
rect 2215 -92 2366 -80
rect 1351 -126 1409 -92
rect 1443 -126 1501 -92
rect 1561 -126 1593 -92
rect 1627 -126 1685 -92
rect 1719 -126 1739 -92
rect 1811 -126 1869 -92
rect 1903 -126 1945 -92
rect 1997 -126 2053 -92
rect 2087 -126 2145 -92
rect 2215 -126 2237 -92
rect 2271 -126 2329 -92
rect 2363 -126 2366 -92
rect 1317 -133 1509 -126
rect 1561 -131 1739 -126
rect 1791 -131 1945 -126
rect 1997 -131 2366 -126
rect 1561 -132 2366 -131
rect 2418 -92 2574 -80
rect 2626 -80 3455 -77
rect 2626 -81 3045 -80
rect 2626 -92 2837 -81
rect 2889 -92 3045 -81
rect 3097 -83 3455 -80
rect 3097 -92 3255 -83
rect 3307 -92 3455 -83
rect 3507 -78 7335 -77
rect 3507 -79 4285 -78
rect 3507 -80 4069 -79
rect 3507 -92 3658 -80
rect 3710 -92 3868 -80
rect 3920 -92 4069 -80
rect 4121 -92 4285 -79
rect 4337 -80 5212 -78
rect 4337 -92 4566 -80
rect 4618 -84 5212 -80
rect 4618 -85 4991 -84
rect 4618 -92 4786 -85
rect 4838 -92 4991 -85
rect 5043 -92 5212 -84
rect 5264 -79 7335 -78
rect 5264 -84 6057 -79
rect 5264 -85 5626 -84
rect 5264 -92 5417 -85
rect 5469 -92 5626 -85
rect 5678 -92 5843 -84
rect 5895 -92 6057 -84
rect 6109 -80 7132 -79
rect 6109 -81 6933 -80
rect 6109 -92 6252 -81
rect 6304 -84 6649 -81
rect 6304 -92 6447 -84
rect 6499 -92 6649 -84
rect 6701 -92 6933 -81
rect 6985 -92 7132 -80
rect 7184 -92 7335 -79
rect 2418 -126 2421 -92
rect 2455 -126 2513 -92
rect 2547 -126 2574 -92
rect 2639 -126 2697 -92
rect 2731 -126 2789 -92
rect 2823 -126 2837 -92
rect 2915 -126 2973 -92
rect 3007 -126 3045 -92
rect 3099 -126 3157 -92
rect 3191 -126 3249 -92
rect 3307 -126 3341 -92
rect 3375 -126 3433 -92
rect 3507 -126 3525 -92
rect 3559 -126 3617 -92
rect 3651 -126 3658 -92
rect 3743 -126 3801 -92
rect 3835 -126 3868 -92
rect 3927 -126 3985 -92
rect 4019 -126 4069 -92
rect 4121 -126 4169 -92
rect 4203 -126 4261 -92
rect 4337 -126 4353 -92
rect 4387 -126 4445 -92
rect 4479 -126 4537 -92
rect 4618 -126 4629 -92
rect 4663 -126 4721 -92
rect 4755 -126 4786 -92
rect 4847 -126 4905 -92
rect 4939 -126 4991 -92
rect 5043 -126 5089 -92
rect 5123 -126 5181 -92
rect 5264 -126 5273 -92
rect 5307 -126 5365 -92
rect 5399 -126 5417 -92
rect 5491 -126 5549 -92
rect 5583 -126 5626 -92
rect 5678 -126 5733 -92
rect 5767 -126 5825 -92
rect 5895 -126 5917 -92
rect 5951 -126 6009 -92
rect 6043 -126 6057 -92
rect 6135 -126 6193 -92
rect 6227 -126 6252 -92
rect 6319 -126 6377 -92
rect 6411 -126 6447 -92
rect 6503 -126 6561 -92
rect 6595 -126 6649 -92
rect 6701 -126 6745 -92
rect 6779 -126 6837 -92
rect 6871 -126 6929 -92
rect 6985 -126 7021 -92
rect 7055 -126 7113 -92
rect 7184 -126 7205 -92
rect 7239 -126 7297 -92
rect 7331 -126 7335 -92
rect 2418 -129 2574 -126
rect 2626 -129 2837 -126
rect 2418 -132 2837 -129
rect 1561 -133 2837 -132
rect 2889 -132 3045 -126
rect 3097 -132 3255 -126
rect 2889 -133 3255 -132
rect -126 -135 3255 -133
rect 3307 -129 3455 -126
rect 3507 -129 3658 -126
rect 3307 -132 3658 -129
rect 3710 -132 3868 -126
rect 3920 -131 4069 -126
rect 4121 -130 4285 -126
rect 4337 -130 4566 -126
rect 4121 -131 4566 -130
rect 3920 -132 4566 -131
rect 4618 -132 4786 -126
rect 3307 -135 4786 -132
rect -126 -137 4786 -135
rect 4838 -136 4991 -126
rect 5043 -130 5212 -126
rect 5264 -130 5417 -126
rect 5043 -136 5417 -130
rect 4838 -137 5417 -136
rect 5469 -136 5626 -126
rect 5678 -136 5843 -126
rect 5895 -131 6057 -126
rect 6109 -131 6252 -126
rect 5895 -133 6252 -131
rect 6304 -133 6447 -126
rect 5895 -136 6447 -133
rect 6499 -133 6649 -126
rect 6701 -132 6933 -126
rect 6985 -131 7132 -126
rect 7184 -129 7335 -126
rect 7387 -78 10817 -77
rect 7387 -79 9034 -78
rect 7387 -80 7987 -79
rect 7387 -92 7600 -80
rect 7652 -81 7987 -80
rect 7652 -92 7798 -81
rect 7850 -92 7987 -81
rect 8039 -92 8199 -79
rect 8251 -92 8416 -79
rect 8468 -83 9034 -79
rect 8468 -92 8621 -83
rect 7387 -126 7389 -92
rect 7423 -126 7481 -92
rect 7515 -126 7573 -92
rect 7652 -126 7665 -92
rect 7699 -126 7757 -92
rect 7791 -126 7798 -92
rect 7883 -126 7941 -92
rect 7975 -126 7987 -92
rect 8067 -126 8125 -92
rect 8159 -126 8199 -92
rect 8251 -126 8309 -92
rect 8343 -126 8401 -92
rect 8468 -126 8493 -92
rect 8527 -126 8585 -92
rect 8619 -126 8621 -92
rect 7387 -129 7600 -126
rect 7184 -131 7600 -129
rect 6985 -132 7600 -131
rect 7652 -132 7798 -126
rect 6701 -133 7798 -132
rect 7850 -131 7987 -126
rect 8039 -131 8199 -126
rect 8251 -131 8416 -126
rect 8468 -131 8621 -126
rect 7850 -133 8621 -131
rect 6499 -135 8621 -133
rect 8673 -92 8826 -83
rect 8878 -92 9034 -83
rect 9086 -79 10817 -78
rect 9086 -92 9317 -79
rect 9369 -81 10195 -79
rect 9369 -92 9510 -81
rect 9562 -83 10195 -81
rect 9562 -92 9736 -83
rect 9788 -92 10001 -83
rect 8673 -126 8677 -92
rect 8711 -126 8769 -92
rect 8803 -126 8826 -92
rect 8895 -126 8953 -92
rect 8987 -126 9034 -92
rect 9086 -126 9137 -92
rect 9171 -126 9229 -92
rect 9263 -126 9317 -92
rect 9369 -126 9413 -92
rect 9447 -126 9505 -92
rect 9562 -126 9597 -92
rect 9631 -126 9689 -92
rect 9723 -126 9736 -92
rect 9815 -126 9873 -92
rect 9907 -126 9965 -92
rect 9999 -126 10001 -92
rect 8673 -135 8826 -126
rect 8878 -130 9034 -126
rect 9086 -130 9317 -126
rect 8878 -131 9317 -130
rect 9369 -131 9510 -126
rect 8878 -133 9510 -131
rect 9562 -133 9736 -126
rect 8878 -135 9736 -133
rect 9788 -135 10001 -126
rect 10053 -92 10195 -83
rect 10247 -80 10817 -79
rect 10247 -88 10597 -80
rect 10247 -92 10393 -88
rect 10445 -92 10597 -88
rect 10649 -92 10817 -80
rect 10869 -78 16876 -77
rect 10869 -81 11260 -78
rect 10869 -92 11032 -81
rect 11084 -92 11260 -81
rect 11312 -79 11895 -78
rect 11312 -81 11702 -79
rect 11312 -92 11464 -81
rect 11516 -92 11702 -81
rect 11754 -92 11895 -79
rect 11947 -80 16876 -78
rect 11947 -83 12348 -80
rect 11947 -92 12092 -83
rect 12144 -92 12348 -83
rect 12400 -81 16876 -80
rect 12400 -83 13460 -81
rect 12400 -84 13041 -83
rect 12400 -92 12587 -84
rect 12639 -88 13041 -84
rect 12639 -92 12820 -88
rect 12872 -92 13041 -88
rect 10053 -126 10057 -92
rect 10091 -126 10149 -92
rect 10183 -126 10195 -92
rect 10275 -126 10333 -92
rect 10367 -126 10393 -92
rect 10459 -126 10517 -92
rect 10551 -126 10597 -92
rect 10649 -126 10701 -92
rect 10735 -126 10793 -92
rect 10869 -126 10885 -92
rect 10919 -126 10977 -92
rect 11011 -126 11032 -92
rect 11103 -126 11161 -92
rect 11195 -126 11253 -92
rect 11312 -126 11345 -92
rect 11379 -126 11437 -92
rect 11516 -126 11529 -92
rect 11563 -126 11621 -92
rect 11655 -126 11702 -92
rect 11754 -126 11805 -92
rect 11839 -126 11895 -92
rect 11947 -126 11989 -92
rect 12023 -126 12081 -92
rect 12144 -126 12173 -92
rect 12207 -126 12265 -92
rect 12299 -126 12348 -92
rect 12400 -126 12449 -92
rect 12483 -126 12541 -92
rect 12575 -126 12587 -92
rect 12667 -126 12725 -92
rect 12759 -126 12817 -92
rect 12872 -126 12909 -92
rect 12943 -126 13001 -92
rect 13035 -126 13041 -92
rect 10053 -131 10195 -126
rect 10247 -131 10393 -126
rect 10053 -135 10393 -131
rect 6499 -136 10393 -135
rect 5469 -137 10393 -136
rect -126 -140 10393 -137
rect 10445 -132 10597 -126
rect 10649 -129 10817 -126
rect 10869 -129 11032 -126
rect 10649 -132 11032 -129
rect 10445 -133 11032 -132
rect 11084 -130 11260 -126
rect 11312 -130 11464 -126
rect 11084 -133 11464 -130
rect 11516 -131 11702 -126
rect 11754 -130 11895 -126
rect 11947 -130 12092 -126
rect 11754 -131 12092 -130
rect 11516 -133 12092 -131
rect 10445 -135 12092 -133
rect 12144 -132 12348 -126
rect 12400 -132 12587 -126
rect 12144 -135 12587 -132
rect 10445 -136 12587 -135
rect 12639 -136 12820 -126
rect 10445 -140 12820 -136
rect 12872 -135 13041 -126
rect 13093 -92 13232 -83
rect 13284 -92 13460 -83
rect 13512 -82 14511 -81
rect 13512 -83 14285 -82
rect 13512 -86 14096 -83
rect 13512 -92 13657 -86
rect 13709 -92 13869 -86
rect 13127 -126 13185 -92
rect 13219 -126 13232 -92
rect 13311 -126 13369 -92
rect 13403 -126 13460 -92
rect 13512 -126 13553 -92
rect 13587 -126 13645 -92
rect 13709 -126 13737 -92
rect 13771 -126 13829 -92
rect 13863 -126 13869 -92
rect 13093 -135 13232 -126
rect 13284 -133 13460 -126
rect 13512 -133 13657 -126
rect 13284 -135 13657 -133
rect 12872 -138 13657 -135
rect 13709 -138 13869 -126
rect 13921 -92 14096 -86
rect 14148 -92 14285 -83
rect 14337 -92 14511 -82
rect 13955 -126 14013 -92
rect 14047 -126 14096 -92
rect 14148 -126 14197 -92
rect 14231 -126 14285 -92
rect 14337 -126 14381 -92
rect 14415 -126 14473 -92
rect 14507 -126 14511 -92
rect 13921 -135 14096 -126
rect 14148 -134 14285 -126
rect 14337 -133 14511 -126
rect 14563 -92 14765 -81
rect 14817 -82 16497 -81
rect 14817 -84 15497 -82
rect 14817 -92 15009 -84
rect 15061 -85 15497 -84
rect 15061 -92 15239 -85
rect 15291 -92 15497 -85
rect 15549 -92 15707 -82
rect 14563 -126 14565 -92
rect 14599 -126 14657 -92
rect 14691 -126 14749 -92
rect 14817 -126 14841 -92
rect 14875 -126 14933 -92
rect 14967 -126 15009 -92
rect 15061 -126 15117 -92
rect 15151 -126 15209 -92
rect 15291 -126 15301 -92
rect 15335 -126 15393 -92
rect 15427 -126 15485 -92
rect 15549 -126 15577 -92
rect 15611 -126 15669 -92
rect 15703 -126 15707 -92
rect 14563 -133 14765 -126
rect 14817 -133 15009 -126
rect 14337 -134 15009 -133
rect 14148 -135 15009 -134
rect 13921 -136 15009 -135
rect 15061 -136 15239 -126
rect 13921 -137 15239 -136
rect 15291 -134 15497 -126
rect 15549 -134 15707 -126
rect 15759 -92 15932 -82
rect 15984 -85 16497 -82
rect 15984 -92 16151 -85
rect 16203 -92 16497 -85
rect 16549 -84 16876 -81
rect 16549 -92 16696 -84
rect 15759 -126 15761 -92
rect 15795 -126 15853 -92
rect 15887 -126 15932 -92
rect 15984 -126 16037 -92
rect 16071 -126 16129 -92
rect 16203 -126 16221 -92
rect 16255 -126 16313 -92
rect 16347 -126 16405 -92
rect 16439 -126 16497 -92
rect 16549 -126 16589 -92
rect 16623 -126 16681 -92
rect 15759 -134 15932 -126
rect 15984 -134 16151 -126
rect 15291 -137 16151 -134
rect 16203 -133 16497 -126
rect 16549 -133 16696 -126
rect 16203 -136 16696 -133
rect 16748 -136 16876 -84
rect 16203 -137 16876 -136
rect 13921 -138 16876 -137
rect 12872 -140 16876 -138
rect -126 -150 16876 -140
rect -126 -153 16861 -150
rect -126 -157 16816 -153
<< via1 >>
rect 53 2971 105 2976
rect 53 2937 65 2971
rect 65 2937 105 2971
rect 53 2924 105 2937
rect 255 2926 307 2978
rect 466 2971 518 2976
rect 656 2971 708 2976
rect 864 2971 916 2978
rect 1066 2971 1118 2978
rect 466 2937 491 2971
rect 491 2937 518 2971
rect 656 2937 675 2971
rect 675 2937 708 2971
rect 864 2937 893 2971
rect 893 2937 916 2971
rect 1066 2937 1077 2971
rect 1077 2937 1118 2971
rect 466 2924 518 2937
rect 656 2924 708 2937
rect 864 2926 916 2937
rect 1066 2926 1118 2937
rect 1265 2928 1317 2980
rect 1460 2971 1512 2977
rect 1661 2971 1713 2979
rect 1878 2971 1930 2977
rect 2152 2971 2204 2980
rect 2429 2971 2481 2973
rect 2652 2971 2704 2976
rect 1460 2937 1503 2971
rect 1503 2937 1512 2971
rect 1661 2937 1687 2971
rect 1687 2937 1713 2971
rect 1878 2937 1905 2971
rect 1905 2937 1930 2971
rect 2152 2937 2181 2971
rect 2181 2937 2204 2971
rect 2429 2937 2457 2971
rect 2457 2937 2481 2971
rect 2652 2937 2699 2971
rect 2699 2937 2704 2971
rect 1460 2925 1512 2937
rect 1661 2927 1713 2937
rect 1878 2925 1930 2937
rect 2152 2928 2204 2937
rect 2429 2921 2481 2937
rect 2652 2924 2704 2937
rect 2884 2923 2936 2975
rect 4520 2971 4572 2972
rect 4828 2971 4880 2973
rect 5028 2971 5080 2974
rect 5247 2971 5299 2973
rect 5493 2971 5545 2972
rect 5701 2971 5753 2974
rect 5903 2971 5955 2975
rect 6096 2971 6148 2974
rect 6468 2971 6520 2973
rect 4520 2937 4541 2971
rect 4541 2937 4572 2971
rect 4828 2937 4875 2971
rect 4875 2937 4880 2971
rect 5028 2937 5059 2971
rect 5059 2937 5080 2971
rect 5247 2937 5277 2971
rect 5277 2937 5299 2971
rect 5493 2937 5519 2971
rect 5519 2937 5545 2971
rect 5701 2937 5703 2971
rect 5703 2937 5737 2971
rect 5737 2937 5753 2971
rect 5903 2937 5921 2971
rect 5921 2937 5955 2971
rect 6096 2937 6105 2971
rect 6105 2937 6148 2971
rect 6468 2937 6473 2971
rect 6473 2937 6520 2971
rect 4520 2920 4572 2937
rect 4828 2921 4880 2937
rect 5028 2922 5080 2937
rect 5247 2921 5299 2937
rect 5493 2920 5545 2937
rect 5701 2922 5753 2937
rect 5903 2923 5955 2937
rect 6096 2922 6148 2937
rect 6468 2921 6520 2937
rect 6657 2919 6709 2971
rect 6947 2937 6991 2971
rect 6991 2937 6999 2971
rect 6947 2919 6999 2937
rect 7220 2921 7272 2973
rect 2866 2664 2918 2674
rect 2866 2630 2876 2664
rect 2876 2630 2910 2664
rect 2910 2630 2918 2664
rect 2866 2622 2918 2630
rect 7427 2622 7479 2674
rect 1171 2385 1223 2437
rect 1390 2427 1442 2441
rect 1673 2427 1725 2441
rect 1882 2427 1934 2441
rect 2153 2427 2205 2439
rect 1390 2393 1411 2427
rect 1411 2393 1442 2427
rect 1673 2393 1687 2427
rect 1687 2393 1721 2427
rect 1721 2393 1725 2427
rect 1882 2393 1905 2427
rect 1905 2393 1934 2427
rect 2153 2393 2181 2427
rect 2181 2393 2205 2427
rect 1390 2389 1442 2393
rect 1673 2389 1725 2393
rect 1882 2389 1934 2393
rect 2153 2387 2205 2393
rect 4228 2385 4280 2437
rect 4477 2427 4529 2440
rect 5075 2427 5127 2432
rect 5304 2427 5356 2432
rect 7022 2427 7074 2437
rect 4477 2393 4507 2427
rect 4507 2393 4529 2427
rect 4477 2388 4529 2393
rect 4821 2374 4873 2426
rect 5075 2393 5093 2427
rect 5093 2393 5127 2427
rect 5304 2393 5335 2427
rect 5335 2393 5356 2427
rect 7022 2393 7025 2427
rect 7025 2393 7074 2427
rect 5075 2380 5127 2393
rect 5304 2380 5356 2393
rect 7022 2385 7074 2393
rect 7226 2387 7278 2439
rect 7549 2385 7601 2437
rect 1024 2250 1077 2303
rect 2866 2250 2918 2302
rect 3418 2256 3471 2309
rect 5809 2256 5862 2309
rect 8200 2256 8253 2309
rect 10592 2256 10645 2309
rect 12983 2256 13036 2309
rect 15376 2256 15429 2309
rect 474 2039 526 2091
rect 1736 2039 1788 2091
rect 2867 2038 2919 2090
rect 4128 2039 4180 2091
rect 5259 2038 5311 2090
rect 6519 2040 6571 2092
rect 7427 2038 7479 2090
rect 7651 2039 7703 2091
rect 8912 2040 8964 2092
rect 10042 2038 10094 2090
rect 11305 2040 11357 2092
rect 12434 2037 12486 2089
rect 13694 2040 13746 2092
rect 14826 2038 14878 2090
rect 16089 2040 16141 2092
rect 19 1829 71 1832
rect 259 1829 311 1830
rect 19 1795 29 1829
rect 29 1795 63 1829
rect 63 1795 71 1829
rect 259 1795 305 1829
rect 305 1795 311 1829
rect 581 1795 615 1829
rect 615 1795 633 1829
rect 19 1780 71 1795
rect 259 1778 311 1795
rect 581 1777 633 1795
rect 799 1778 851 1830
rect 2703 1829 2755 1834
rect 3028 1829 3080 1836
rect 2703 1795 2731 1829
rect 2731 1795 2755 1829
rect 3028 1795 3065 1829
rect 3065 1795 3080 1829
rect 2703 1782 2755 1795
rect 3028 1784 3080 1795
rect 3296 1784 3348 1836
rect 3562 1784 3614 1836
rect 3802 1782 3854 1834
rect 5596 1785 5648 1837
rect 5962 1788 6014 1840
rect 6206 1829 6258 1840
rect 6629 1829 6681 1831
rect 6206 1795 6245 1829
rect 6245 1795 6258 1829
rect 6629 1795 6647 1829
rect 6647 1795 6681 1829
rect 6206 1788 6258 1795
rect 6629 1779 6681 1795
rect 8572 1781 8624 1833
rect 8824 1829 8876 1830
rect 9030 1829 9082 1838
rect 9313 1829 9365 1832
rect 9611 1829 9663 1833
rect 11443 1829 11495 1834
rect 11653 1829 11705 1836
rect 12004 1829 12056 1834
rect 12284 1829 12336 1834
rect 12601 1829 12653 1833
rect 14391 1829 14443 1831
rect 14686 1829 14738 1831
rect 8824 1795 8857 1829
rect 8857 1795 8876 1829
rect 9030 1795 9041 1829
rect 9041 1795 9082 1829
rect 9313 1795 9317 1829
rect 9317 1795 9365 1829
rect 9611 1795 9631 1829
rect 9631 1795 9663 1829
rect 11443 1795 11491 1829
rect 11491 1795 11495 1829
rect 11653 1795 11675 1829
rect 11675 1795 11705 1829
rect 12004 1795 12023 1829
rect 12023 1795 12056 1829
rect 12284 1795 12299 1829
rect 12299 1795 12336 1829
rect 12601 1795 12633 1829
rect 12633 1795 12653 1829
rect 14391 1795 14415 1829
rect 14415 1795 14443 1829
rect 14686 1795 14691 1829
rect 14691 1795 14738 1829
rect 8824 1778 8876 1795
rect 9030 1786 9082 1795
rect 9313 1780 9365 1795
rect 9611 1781 9663 1795
rect 11443 1782 11495 1795
rect 11653 1784 11705 1795
rect 12004 1782 12056 1795
rect 12284 1782 12336 1795
rect 12601 1781 12653 1795
rect 14391 1779 14443 1795
rect 14686 1779 14738 1795
rect 14973 1779 15025 1831
rect 15263 1779 15315 1831
rect 15547 1782 15599 1834
rect 475 1607 527 1617
rect 475 1573 484 1607
rect 484 1573 518 1607
rect 518 1573 527 1607
rect 475 1565 527 1573
rect 1557 1592 1609 1603
rect 1557 1558 1566 1592
rect 1566 1558 1600 1592
rect 1600 1558 1609 1592
rect 1557 1550 1609 1558
rect 1737 1607 1789 1617
rect 1737 1573 1746 1607
rect 1746 1573 1780 1607
rect 1780 1573 1789 1607
rect 1737 1565 1789 1573
rect 2868 1606 2920 1616
rect 2868 1572 2877 1606
rect 2877 1572 2911 1606
rect 2911 1572 2920 1606
rect 2868 1564 2920 1572
rect 3949 1591 4001 1602
rect 3949 1557 3958 1591
rect 3958 1557 3992 1591
rect 3992 1557 4001 1591
rect 3949 1549 4001 1557
rect 4129 1607 4181 1617
rect 4129 1573 4138 1607
rect 4138 1573 4172 1607
rect 4172 1573 4181 1607
rect 4129 1565 4181 1573
rect 5260 1606 5312 1616
rect 5260 1572 5269 1606
rect 5269 1572 5303 1606
rect 5303 1572 5312 1606
rect 5260 1564 5312 1572
rect 6339 1591 6391 1602
rect 6339 1557 6348 1591
rect 6348 1557 6382 1591
rect 6382 1557 6391 1591
rect 6339 1549 6391 1557
rect 6520 1608 6572 1618
rect 6520 1574 6529 1608
rect 6529 1574 6563 1608
rect 6563 1574 6572 1608
rect 6520 1566 6572 1574
rect 7652 1607 7704 1617
rect 7652 1573 7661 1607
rect 7661 1573 7695 1607
rect 7695 1573 7704 1607
rect 7652 1565 7704 1573
rect 8733 1592 8785 1603
rect 8733 1558 8742 1592
rect 8742 1558 8776 1592
rect 8776 1558 8785 1592
rect 8733 1550 8785 1558
rect 8913 1608 8965 1618
rect 8913 1574 8922 1608
rect 8922 1574 8956 1608
rect 8956 1574 8965 1608
rect 8913 1566 8965 1574
rect 10043 1606 10095 1616
rect 10043 1572 10052 1606
rect 10052 1572 10086 1606
rect 10086 1572 10095 1606
rect 10043 1564 10095 1572
rect 11125 1591 11177 1602
rect 11125 1557 11134 1591
rect 11134 1557 11168 1591
rect 11168 1557 11177 1591
rect 11125 1549 11177 1557
rect 11306 1608 11358 1618
rect 11306 1574 11315 1608
rect 11315 1574 11349 1608
rect 11349 1574 11358 1608
rect 11306 1566 11358 1574
rect 12435 1605 12487 1615
rect 12435 1571 12444 1605
rect 12444 1571 12478 1605
rect 12478 1571 12487 1605
rect 12435 1563 12487 1571
rect 13514 1591 13566 1602
rect 13514 1557 13523 1591
rect 13523 1557 13557 1591
rect 13557 1557 13566 1591
rect 13514 1549 13566 1557
rect 13695 1608 13747 1618
rect 13695 1574 13704 1608
rect 13704 1574 13738 1608
rect 13738 1574 13747 1608
rect 13695 1566 13747 1574
rect 14827 1606 14879 1616
rect 14827 1572 14836 1606
rect 14836 1572 14870 1606
rect 14870 1572 14879 1606
rect 14827 1564 14879 1572
rect 15909 1592 15961 1603
rect 15909 1558 15918 1592
rect 15918 1558 15952 1592
rect 15952 1558 15961 1592
rect 15909 1550 15961 1558
rect 16090 1608 16142 1618
rect 16090 1574 16099 1608
rect 16099 1574 16133 1608
rect 16133 1574 16142 1608
rect 16090 1566 16142 1574
rect 18 1406 70 1414
rect 18 1372 28 1406
rect 28 1372 62 1406
rect 62 1372 70 1406
rect 18 1362 70 1372
rect 356 1400 408 1452
rect 1957 1401 2009 1453
rect 2194 1404 2246 1414
rect 2194 1370 2204 1404
rect 2204 1370 2238 1404
rect 2238 1370 2246 1404
rect 2194 1362 2246 1370
rect 2410 1406 2462 1414
rect 2410 1372 2420 1406
rect 2420 1372 2454 1406
rect 2454 1372 2462 1406
rect 2410 1362 2462 1372
rect 2748 1400 2800 1452
rect 4349 1401 4401 1453
rect 4588 1404 4640 1414
rect 4588 1370 4598 1404
rect 4598 1370 4632 1404
rect 4632 1370 4640 1404
rect 4588 1362 4640 1370
rect 4802 1406 4854 1414
rect 4802 1372 4812 1406
rect 4812 1372 4846 1406
rect 4846 1372 4854 1406
rect 4802 1362 4854 1372
rect 5139 1401 5191 1453
rect 6740 1402 6792 1454
rect 6978 1406 7030 1416
rect 6978 1372 6988 1406
rect 6988 1372 7022 1406
rect 7022 1372 7030 1406
rect 6978 1364 7030 1372
rect 7194 1406 7246 1414
rect 7194 1372 7204 1406
rect 7204 1372 7238 1406
rect 7238 1372 7246 1406
rect 7194 1362 7246 1372
rect 7532 1400 7584 1452
rect 9133 1401 9185 1453
rect 9370 1404 9422 1414
rect 9370 1370 9380 1404
rect 9380 1370 9414 1404
rect 9414 1370 9422 1404
rect 9370 1362 9422 1370
rect 9585 1407 9637 1415
rect 9585 1373 9595 1407
rect 9595 1373 9629 1407
rect 9629 1373 9637 1407
rect 9585 1363 9637 1373
rect 9924 1401 9976 1453
rect 11525 1402 11577 1454
rect 11762 1406 11814 1416
rect 11762 1372 11772 1406
rect 11772 1372 11806 1406
rect 11806 1372 11814 1406
rect 11762 1364 11814 1372
rect 11977 1406 12029 1414
rect 11977 1372 11987 1406
rect 11987 1372 12021 1406
rect 12021 1372 12029 1406
rect 11977 1362 12029 1372
rect 12316 1401 12368 1453
rect 13917 1402 13969 1454
rect 14154 1404 14206 1414
rect 14154 1370 14164 1404
rect 14164 1370 14198 1404
rect 14198 1370 14206 1404
rect 14154 1362 14206 1370
rect 14370 1407 14422 1415
rect 14370 1373 14380 1407
rect 14380 1373 14414 1407
rect 14414 1373 14422 1407
rect 14370 1363 14422 1373
rect 14711 1401 14763 1453
rect 16312 1402 16364 1454
rect 16546 1406 16598 1416
rect 16546 1372 16556 1406
rect 16556 1372 16590 1406
rect 16590 1372 16598 1406
rect 16546 1364 16598 1372
rect 1210 1242 1262 1294
rect 1427 1285 1479 1294
rect 1646 1285 1698 1294
rect 1859 1285 1911 1290
rect 2070 1285 2122 1290
rect 4194 1285 4246 1290
rect 4472 1285 4524 1289
rect 5044 1285 5096 1294
rect 5283 1285 5335 1294
rect 7441 1285 7493 1292
rect 7668 1285 7720 1297
rect 7858 1285 7910 1299
rect 1427 1251 1463 1285
rect 1463 1251 1479 1285
rect 1646 1251 1647 1285
rect 1647 1251 1681 1285
rect 1681 1251 1698 1285
rect 1859 1251 1865 1285
rect 1865 1251 1911 1285
rect 2070 1251 2107 1285
rect 2107 1251 2122 1285
rect 4194 1251 4223 1285
rect 4223 1251 4246 1285
rect 4472 1251 4499 1285
rect 4499 1251 4524 1285
rect 5044 1251 5089 1285
rect 5089 1251 5096 1285
rect 5283 1251 5307 1285
rect 5307 1251 5335 1285
rect 7441 1251 7481 1285
rect 7481 1251 7493 1285
rect 7668 1251 7699 1285
rect 7699 1251 7720 1285
rect 7858 1251 7883 1285
rect 7883 1251 7910 1285
rect 1427 1242 1479 1251
rect 1646 1242 1698 1251
rect 1859 1238 1911 1251
rect 2070 1238 2122 1251
rect 4194 1238 4246 1251
rect 4472 1237 4524 1251
rect 5044 1242 5096 1251
rect 5283 1242 5335 1251
rect 7441 1240 7493 1251
rect 7668 1245 7720 1251
rect 7858 1247 7910 1251
rect 8074 1238 8126 1290
rect 10055 1285 10107 1293
rect 10284 1285 10336 1296
rect 10055 1251 10057 1285
rect 10057 1251 10091 1285
rect 10091 1251 10107 1285
rect 10284 1251 10333 1285
rect 10333 1251 10336 1285
rect 10055 1241 10107 1251
rect 10284 1244 10336 1251
rect 10510 1249 10562 1301
rect 10738 1241 10790 1293
rect 10974 1247 11026 1299
rect 11166 1285 11218 1290
rect 11166 1251 11215 1285
rect 11215 1251 11218 1285
rect 11166 1238 11218 1251
rect 12901 1238 12953 1290
rect 13105 1243 13157 1295
rect 13296 1238 13348 1290
rect 13498 1285 13550 1289
rect 13788 1285 13840 1290
rect 14073 1285 14125 1289
rect 15828 1285 15880 1294
rect 16022 1285 16074 1298
rect 16211 1285 16263 1295
rect 16434 1285 16486 1297
rect 13498 1251 13513 1285
rect 13513 1251 13547 1285
rect 13547 1251 13550 1285
rect 13788 1251 13789 1285
rect 13789 1251 13823 1285
rect 13823 1251 13840 1285
rect 14073 1251 14099 1285
rect 14099 1251 14125 1285
rect 15828 1251 15849 1285
rect 15849 1251 15880 1285
rect 16022 1251 16033 1285
rect 16033 1251 16074 1285
rect 16211 1251 16217 1285
rect 16217 1251 16263 1285
rect 16434 1251 16459 1285
rect 16459 1251 16486 1285
rect 13498 1237 13550 1251
rect 13788 1238 13840 1251
rect 14073 1237 14125 1251
rect 15828 1242 15880 1251
rect 16022 1246 16074 1251
rect 16211 1243 16263 1251
rect 16434 1245 16486 1251
rect 265 1141 317 1149
rect 467 1141 519 1145
rect 656 1141 708 1142
rect 885 1141 937 1143
rect 2654 1141 2706 1146
rect 2869 1141 2921 1143
rect 3262 1141 3314 1150
rect 3542 1141 3594 1148
rect 3761 1141 3813 1146
rect 5582 1141 5634 1143
rect 6327 1141 6379 1145
rect 6518 1141 6570 1147
rect 8563 1141 8615 1149
rect 8753 1141 8805 1151
rect 8947 1141 8999 1149
rect 9258 1141 9310 1145
rect 11441 1141 11493 1144
rect 11645 1141 11697 1144
rect 12449 1141 12501 1142
rect 12653 1141 12705 1142
rect 14613 1141 14665 1150
rect 14846 1141 14898 1148
rect 15053 1141 15105 1146
rect 15262 1141 15314 1148
rect 15542 1141 15594 1150
rect 265 1107 305 1141
rect 305 1107 317 1141
rect 467 1107 489 1141
rect 489 1107 519 1141
rect 656 1107 673 1141
rect 673 1107 707 1141
rect 707 1107 708 1141
rect 885 1107 891 1141
rect 891 1107 937 1141
rect 2654 1107 2697 1141
rect 2697 1107 2706 1141
rect 2869 1107 2881 1141
rect 2881 1107 2915 1141
rect 2915 1107 2921 1141
rect 3067 1107 3099 1140
rect 3099 1107 3119 1140
rect 3262 1107 3283 1141
rect 3283 1107 3314 1141
rect 3542 1107 3559 1141
rect 3559 1107 3594 1141
rect 3761 1107 3801 1141
rect 3801 1107 3813 1141
rect 5582 1107 5583 1141
rect 5583 1107 5634 1141
rect 5933 1107 5951 1140
rect 5951 1107 5985 1140
rect 6122 1107 6135 1138
rect 6135 1107 6174 1138
rect 6327 1107 6377 1141
rect 6377 1107 6379 1141
rect 6518 1107 6561 1141
rect 6561 1107 6570 1141
rect 8563 1107 8585 1141
rect 8585 1107 8615 1141
rect 8753 1107 8769 1141
rect 8769 1107 8803 1141
rect 8803 1107 8805 1141
rect 8947 1107 8953 1141
rect 8953 1107 8987 1141
rect 8987 1107 8999 1141
rect 9258 1107 9263 1141
rect 9263 1107 9310 1141
rect 11441 1107 11471 1141
rect 11471 1107 11493 1141
rect 11645 1107 11655 1141
rect 11655 1107 11697 1141
rect 265 1097 317 1107
rect 467 1093 519 1107
rect 656 1090 708 1107
rect 885 1091 937 1107
rect 2654 1094 2706 1107
rect 2869 1091 2921 1107
rect 3067 1088 3119 1107
rect 3262 1098 3314 1107
rect 3542 1096 3594 1107
rect 3761 1094 3813 1107
rect 5582 1091 5634 1107
rect 5933 1088 5985 1107
rect 6122 1086 6174 1107
rect 6327 1093 6379 1107
rect 6518 1095 6570 1107
rect 8563 1097 8615 1107
rect 8753 1099 8805 1107
rect 8947 1097 8999 1107
rect 9258 1093 9310 1107
rect 11441 1092 11493 1107
rect 11645 1092 11697 1107
rect 12210 1088 12262 1140
rect 12449 1107 12483 1141
rect 12483 1107 12501 1141
rect 12653 1107 12667 1141
rect 12667 1107 12705 1141
rect 14613 1107 14657 1141
rect 14657 1107 14665 1141
rect 14846 1107 14875 1141
rect 14875 1107 14898 1141
rect 15053 1107 15059 1141
rect 15059 1107 15105 1141
rect 15262 1107 15301 1141
rect 15301 1107 15314 1141
rect 15542 1107 15577 1141
rect 15577 1107 15594 1141
rect 12449 1090 12501 1107
rect 12653 1090 12705 1107
rect 14613 1098 14665 1107
rect 14846 1096 14898 1107
rect 15053 1094 15105 1107
rect 15262 1096 15314 1107
rect 15542 1098 15594 1107
rect 2324 1034 2376 1042
rect 2324 1000 2334 1034
rect 2334 1000 2368 1034
rect 2368 1000 2376 1034
rect 2324 990 2376 1000
rect 4716 1034 4768 1042
rect 4716 1000 4726 1034
rect 4726 1000 4760 1034
rect 4760 1000 4768 1034
rect 4716 990 4768 1000
rect 7108 1034 7160 1042
rect 7108 1000 7118 1034
rect 7118 1000 7152 1034
rect 7152 1000 7160 1034
rect 7108 990 7160 1000
rect 9500 1034 9552 1042
rect 9500 1000 9510 1034
rect 9510 1000 9544 1034
rect 9544 1000 9552 1034
rect 9500 990 9552 1000
rect 11892 1034 11944 1042
rect 11892 1000 11902 1034
rect 11902 1000 11936 1034
rect 11936 1000 11944 1034
rect 11892 990 11944 1000
rect 14284 1034 14336 1042
rect 14284 1000 14294 1034
rect 14294 1000 14328 1034
rect 14328 1000 14336 1034
rect 14284 990 14336 1000
rect 16676 1034 16728 1042
rect 16676 1000 16686 1034
rect 16686 1000 16720 1034
rect 16720 1000 16728 1034
rect 16676 990 16728 1000
rect 2042 955 2094 965
rect 2042 921 2051 955
rect 2051 921 2085 955
rect 2085 921 2094 955
rect 4434 956 4486 966
rect 2042 913 2094 921
rect 18 859 70 869
rect 18 825 26 859
rect 26 825 60 859
rect 60 825 70 859
rect 18 817 70 825
rect 357 883 409 894
rect 357 849 366 883
rect 366 849 400 883
rect 400 849 409 883
rect 357 841 409 849
rect 4434 922 4443 956
rect 4443 922 4477 956
rect 4477 922 4486 956
rect 6825 956 6877 966
rect 4434 914 4486 922
rect 2410 859 2462 869
rect 2410 825 2418 859
rect 2418 825 2452 859
rect 2452 825 2462 859
rect 2410 817 2462 825
rect 2749 883 2801 894
rect 2749 849 2758 883
rect 2758 849 2792 883
rect 2792 849 2801 883
rect 2749 841 2801 849
rect 6825 922 6834 956
rect 6834 922 6868 956
rect 6868 922 6877 956
rect 9218 957 9270 967
rect 6825 914 6877 922
rect 4802 859 4854 869
rect 4802 825 4810 859
rect 4810 825 4844 859
rect 4844 825 4854 859
rect 4802 817 4854 825
rect 5141 884 5193 895
rect 5141 850 5150 884
rect 5150 850 5184 884
rect 5184 850 5193 884
rect 5141 842 5193 850
rect 9218 923 9227 957
rect 9227 923 9261 957
rect 9261 923 9270 957
rect 11609 956 11661 966
rect 9218 915 9270 923
rect 11609 922 11618 956
rect 11618 922 11652 956
rect 11652 922 11661 956
rect 14002 955 14054 965
rect 11609 914 11661 922
rect 1025 718 1077 770
rect 7194 859 7246 869
rect 7194 825 7202 859
rect 7202 825 7236 859
rect 7236 825 7246 859
rect 7194 817 7246 825
rect 7533 884 7585 895
rect 7533 850 7542 884
rect 7542 850 7576 884
rect 7576 850 7585 884
rect 7533 842 7585 850
rect 3418 718 3470 770
rect 9585 860 9637 870
rect 9585 826 9593 860
rect 9593 826 9627 860
rect 9627 826 9637 860
rect 9585 818 9637 826
rect 9925 883 9977 894
rect 9925 849 9934 883
rect 9934 849 9968 883
rect 9968 849 9977 883
rect 9925 841 9977 849
rect 14002 921 14011 955
rect 14011 921 14045 955
rect 14045 921 14054 955
rect 16395 957 16447 967
rect 14002 913 14054 921
rect 5810 718 5862 770
rect 11977 859 12029 869
rect 11977 825 11985 859
rect 11985 825 12019 859
rect 12019 825 12029 859
rect 11977 817 12029 825
rect 12317 884 12369 895
rect 12317 850 12326 884
rect 12326 850 12360 884
rect 12360 850 12369 884
rect 12317 842 12369 850
rect 16395 923 16404 957
rect 16404 923 16438 957
rect 16438 923 16447 957
rect 16395 915 16447 923
rect 8202 718 8254 770
rect 14370 860 14422 870
rect 14370 826 14378 860
rect 14378 826 14412 860
rect 14412 826 14422 860
rect 14370 818 14422 826
rect 14710 883 14762 894
rect 14710 849 14719 883
rect 14719 849 14753 883
rect 14753 849 14762 883
rect 14710 841 14762 849
rect 10593 718 10645 770
rect 12985 718 13037 770
rect 15377 718 15429 770
rect 1192 597 1244 600
rect 1421 597 1473 612
rect 1640 597 1692 602
rect 1832 597 1884 606
rect 2326 597 2378 604
rect 4118 597 4170 603
rect 4511 597 4563 601
rect 4708 597 4760 609
rect 5038 597 5090 611
rect 5234 597 5286 611
rect 7141 597 7193 604
rect 7442 597 7494 608
rect 7648 597 7700 609
rect 7858 597 7910 605
rect 1192 563 1225 597
rect 1225 563 1244 597
rect 1421 563 1443 597
rect 1443 563 1473 597
rect 1640 563 1685 597
rect 1685 563 1692 597
rect 1832 563 1869 597
rect 1869 563 1884 597
rect 2326 563 2329 597
rect 2329 563 2363 597
rect 2363 563 2378 597
rect 4118 563 4169 597
rect 4169 563 4170 597
rect 4511 563 4537 597
rect 4537 563 4563 597
rect 4708 563 4721 597
rect 4721 563 4755 597
rect 4755 563 4760 597
rect 5038 563 5089 597
rect 5089 563 5090 597
rect 5234 563 5273 597
rect 5273 563 5286 597
rect 7141 563 7147 597
rect 7147 563 7193 597
rect 7442 563 7481 597
rect 7481 563 7494 597
rect 7648 563 7665 597
rect 7665 563 7699 597
rect 7699 563 7700 597
rect 7858 563 7883 597
rect 7883 563 7910 597
rect 1192 548 1244 563
rect 1421 560 1473 563
rect 1640 550 1692 563
rect 1832 554 1884 563
rect 2326 552 2378 563
rect 4118 551 4170 563
rect 4511 549 4563 563
rect 4708 557 4760 563
rect 5038 559 5090 563
rect 5234 559 5286 563
rect 7141 552 7193 563
rect 7442 556 7494 563
rect 7648 557 7700 563
rect 7858 553 7910 563
rect 8069 559 8121 611
rect 9949 597 10001 600
rect 10206 597 10258 607
rect 10456 597 10508 603
rect 10727 597 10779 608
rect 10968 597 11020 611
rect 11193 597 11245 607
rect 12900 597 12952 605
rect 13101 597 13153 606
rect 13319 597 13371 602
rect 13526 597 13578 606
rect 13731 597 13783 605
rect 14078 597 14130 601
rect 15830 597 15882 605
rect 16021 597 16073 608
rect 16216 597 16268 610
rect 16663 597 16715 605
rect 9949 563 9965 597
rect 9965 563 9999 597
rect 9999 563 10001 597
rect 10206 563 10241 597
rect 10241 563 10258 597
rect 10456 563 10459 597
rect 10459 563 10508 597
rect 10727 563 10735 597
rect 10735 563 10779 597
rect 10968 563 10977 597
rect 10977 563 11011 597
rect 11011 563 11020 597
rect 11193 563 11195 597
rect 11195 563 11245 597
rect 12900 563 12909 597
rect 12909 563 12943 597
rect 12943 563 12952 597
rect 13101 563 13127 597
rect 13127 563 13153 597
rect 13319 563 13369 597
rect 13369 563 13371 597
rect 13526 563 13553 597
rect 13553 563 13578 597
rect 13731 563 13737 597
rect 13737 563 13771 597
rect 13771 563 13783 597
rect 14078 563 14105 597
rect 14105 563 14130 597
rect 15830 563 15853 597
rect 15853 563 15882 597
rect 16021 563 16037 597
rect 16037 563 16071 597
rect 16071 563 16073 597
rect 16216 563 16221 597
rect 16221 563 16255 597
rect 16255 563 16268 597
rect 16663 563 16681 597
rect 16681 563 16715 597
rect 9949 548 10001 563
rect 10206 555 10258 563
rect 10456 551 10508 563
rect 10727 556 10779 563
rect 10968 559 11020 563
rect 11193 555 11245 563
rect 12900 553 12952 563
rect 13101 554 13153 563
rect 13319 550 13371 563
rect 13526 554 13578 563
rect 13731 553 13783 563
rect 14078 549 14130 563
rect 15830 553 15882 563
rect 16021 556 16073 563
rect 16216 558 16268 563
rect 16663 553 16715 563
rect 47 452 99 456
rect 495 452 547 459
rect 47 418 63 452
rect 63 418 99 452
rect 280 418 305 452
rect 305 418 332 452
rect 495 418 523 452
rect 523 418 547 452
rect 47 404 99 418
rect 280 400 332 418
rect 495 407 547 418
rect 713 404 765 456
rect 929 452 981 457
rect 2650 452 2702 453
rect 2840 452 2892 453
rect 3050 452 3102 456
rect 3267 452 3319 453
rect 929 418 949 452
rect 949 418 981 452
rect 2650 418 2697 452
rect 2697 418 2702 452
rect 2840 418 2881 452
rect 2881 418 2892 452
rect 3050 418 3065 452
rect 3065 418 3099 452
rect 3099 418 3102 452
rect 3267 418 3283 452
rect 3283 418 3319 452
rect 929 405 981 418
rect 2650 401 2702 418
rect 2840 401 2892 418
rect 3050 404 3102 418
rect 3267 401 3319 418
rect 3562 404 3614 456
rect 3786 452 3838 461
rect 5664 452 5716 454
rect 6216 452 6268 456
rect 6433 452 6485 461
rect 6634 452 6686 458
rect 9529 452 9581 457
rect 11430 452 11482 453
rect 11686 452 11738 453
rect 11921 452 11973 453
rect 3786 418 3801 452
rect 3801 418 3835 452
rect 3835 418 3838 452
rect 5664 418 5675 452
rect 5675 418 5716 452
rect 5964 418 6009 452
rect 6009 418 6016 452
rect 6216 418 6227 452
rect 6227 418 6268 452
rect 6433 418 6469 452
rect 6469 418 6485 452
rect 6634 418 6653 452
rect 6653 418 6686 452
rect 8519 418 8527 449
rect 8527 418 8571 449
rect 3786 409 3838 418
rect 5664 402 5716 418
rect 5964 400 6016 418
rect 6216 404 6268 418
rect 6433 409 6485 418
rect 6634 406 6686 418
rect 8519 397 8571 418
rect 8711 397 8763 449
rect 8911 418 8953 449
rect 8953 418 8963 449
rect 9529 418 9539 452
rect 9539 418 9581 452
rect 11430 418 11437 452
rect 11437 418 11471 452
rect 11471 418 11482 452
rect 11686 418 11713 452
rect 11713 418 11738 452
rect 11921 418 11931 452
rect 11931 418 11973 452
rect 8911 397 8963 418
rect 9529 405 9581 418
rect 11430 401 11482 418
rect 11686 401 11738 418
rect 11921 401 11973 418
rect 12210 403 12262 455
rect 12400 452 12452 453
rect 12604 452 12656 455
rect 14390 452 14442 461
rect 14632 452 14684 457
rect 14832 452 14884 456
rect 15022 452 15074 464
rect 12400 418 12449 452
rect 12449 418 12452 452
rect 12604 418 12633 452
rect 12633 418 12656 452
rect 14390 418 14415 452
rect 14415 418 14442 452
rect 14632 418 14657 452
rect 14657 418 14684 452
rect 14832 418 14841 452
rect 14841 418 14875 452
rect 14875 418 14884 452
rect 15022 418 15025 452
rect 15025 418 15059 452
rect 15059 418 15074 452
rect 12400 401 12452 418
rect 12604 403 12656 418
rect 14390 409 14442 418
rect 14632 405 14684 418
rect 14832 404 14884 418
rect 15022 412 15074 418
rect 15243 410 15295 462
rect 15539 452 15591 457
rect 15539 418 15577 452
rect 15577 418 15591 452
rect 15539 405 15591 418
rect 17 342 69 350
rect 17 308 26 342
rect 26 308 60 342
rect 60 308 69 342
rect 2409 342 2461 350
rect 17 298 69 308
rect 297 276 349 286
rect 297 242 306 276
rect 306 242 340 276
rect 340 242 349 276
rect 297 234 349 242
rect 1025 262 1077 314
rect 2409 308 2418 342
rect 2418 308 2452 342
rect 2452 308 2461 342
rect 4802 342 4854 350
rect 2409 298 2461 308
rect 2689 276 2741 286
rect 2689 242 2698 276
rect 2698 242 2732 276
rect 2732 242 2741 276
rect 2689 234 2741 242
rect 2304 205 2358 215
rect 2304 171 2314 205
rect 2314 171 2348 205
rect 2348 171 2358 205
rect 2304 163 2358 171
rect 1959 149 2011 160
rect 1959 115 1968 149
rect 1968 115 2002 149
rect 2002 115 2011 149
rect 1959 107 2011 115
rect 3417 263 3469 315
rect 4802 308 4811 342
rect 4811 308 4845 342
rect 4845 308 4854 342
rect 7193 342 7245 350
rect 4802 298 4854 308
rect 5080 276 5132 286
rect 5080 242 5089 276
rect 5089 242 5123 276
rect 5123 242 5132 276
rect 5080 234 5132 242
rect 4698 205 4752 215
rect 4698 171 4708 205
rect 4708 171 4742 205
rect 4742 171 4752 205
rect 4698 163 4752 171
rect 4351 149 4403 160
rect 4351 115 4360 149
rect 4360 115 4394 149
rect 4394 115 4403 149
rect 4351 107 4403 115
rect 5809 262 5861 314
rect 7193 308 7202 342
rect 7202 308 7236 342
rect 7236 308 7245 342
rect 9585 341 9637 349
rect 7193 298 7245 308
rect 7473 276 7525 286
rect 7473 242 7482 276
rect 7482 242 7516 276
rect 7516 242 7525 276
rect 7473 234 7525 242
rect 7088 207 7142 217
rect 7088 173 7098 207
rect 7098 173 7132 207
rect 7132 173 7142 207
rect 7088 165 7142 173
rect 6742 150 6794 160
rect 6742 116 6751 150
rect 6751 116 6785 150
rect 6785 116 6794 150
rect 6742 108 6794 116
rect 8201 262 8253 314
rect 9585 307 9594 341
rect 9594 307 9628 341
rect 9628 307 9637 341
rect 11978 343 12030 351
rect 9585 297 9637 307
rect 9865 276 9917 286
rect 9865 242 9874 276
rect 9874 242 9908 276
rect 9908 242 9917 276
rect 9865 234 9917 242
rect 9480 205 9534 215
rect 9480 171 9490 205
rect 9490 171 9524 205
rect 9524 171 9534 205
rect 9480 163 9534 171
rect 9135 149 9187 160
rect 9135 115 9144 149
rect 9144 115 9178 149
rect 9178 115 9187 149
rect 9135 107 9187 115
rect 10593 262 10645 314
rect 11978 309 11987 343
rect 11987 309 12021 343
rect 12021 309 12030 343
rect 14369 343 14421 351
rect 11978 299 12030 309
rect 12256 277 12308 287
rect 12256 243 12265 277
rect 12265 243 12299 277
rect 12299 243 12308 277
rect 12256 235 12308 243
rect 11872 207 11926 217
rect 11872 173 11882 207
rect 11882 173 11916 207
rect 11916 173 11926 207
rect 11872 165 11926 173
rect 11526 149 11578 160
rect 11526 115 11535 149
rect 11535 115 11569 149
rect 11569 115 11578 149
rect 11526 107 11578 115
rect 12985 263 13037 315
rect 14369 309 14378 343
rect 14378 309 14412 343
rect 14412 309 14421 343
rect 14369 299 14421 309
rect 14649 276 14701 286
rect 14649 242 14658 276
rect 14658 242 14692 276
rect 14692 242 14701 276
rect 14649 234 14701 242
rect 14264 205 14318 215
rect 14264 171 14274 205
rect 14274 171 14308 205
rect 14308 171 14318 205
rect 14264 163 14318 171
rect 13919 149 13971 160
rect 13919 115 13928 149
rect 13928 115 13962 149
rect 13962 115 13971 149
rect 13919 107 13971 115
rect 15377 263 15429 315
rect 16656 207 16710 217
rect 16656 173 16666 207
rect 16666 173 16700 207
rect 16700 173 16710 207
rect 16656 165 16710 173
rect 16312 149 16364 160
rect 16312 115 16321 149
rect 16321 115 16355 149
rect 16355 115 16364 149
rect 16312 107 16364 115
rect 421 -92 473 -76
rect 421 -126 431 -92
rect 431 -126 473 -92
rect 421 -128 473 -126
rect 620 -131 672 -79
rect 831 -92 883 -79
rect 1037 -92 1089 -79
rect 831 -126 857 -92
rect 857 -126 883 -92
rect 1037 -126 1041 -92
rect 1041 -126 1075 -92
rect 1075 -126 1089 -92
rect 831 -131 883 -126
rect 1037 -131 1089 -126
rect 1265 -133 1317 -81
rect 1509 -92 1561 -81
rect 1739 -92 1791 -79
rect 1945 -92 1997 -79
rect 2163 -92 2215 -74
rect 1509 -126 1535 -92
rect 1535 -126 1561 -92
rect 1739 -126 1777 -92
rect 1777 -126 1791 -92
rect 1945 -126 1961 -92
rect 1961 -126 1995 -92
rect 1995 -126 1997 -92
rect 2163 -126 2179 -92
rect 2179 -126 2215 -92
rect 1509 -133 1561 -126
rect 1739 -131 1791 -126
rect 1945 -131 1997 -126
rect 2366 -132 2418 -80
rect 2574 -92 2626 -77
rect 2837 -92 2889 -81
rect 3045 -92 3097 -80
rect 3255 -92 3307 -83
rect 3455 -92 3507 -77
rect 3658 -92 3710 -80
rect 3868 -92 3920 -80
rect 4069 -92 4121 -79
rect 4285 -92 4337 -78
rect 4566 -92 4618 -80
rect 4786 -92 4838 -85
rect 4991 -92 5043 -84
rect 5212 -92 5264 -78
rect 5417 -92 5469 -85
rect 5626 -92 5678 -84
rect 5843 -92 5895 -84
rect 6057 -92 6109 -79
rect 6252 -92 6304 -81
rect 6447 -92 6499 -84
rect 6649 -92 6701 -81
rect 6933 -92 6985 -80
rect 7132 -92 7184 -79
rect 2574 -126 2605 -92
rect 2605 -126 2626 -92
rect 2837 -126 2881 -92
rect 2881 -126 2889 -92
rect 3045 -126 3065 -92
rect 3065 -126 3097 -92
rect 3255 -126 3283 -92
rect 3283 -126 3307 -92
rect 3455 -126 3467 -92
rect 3467 -126 3507 -92
rect 3658 -126 3709 -92
rect 3709 -126 3710 -92
rect 3868 -126 3893 -92
rect 3893 -126 3920 -92
rect 4069 -126 4077 -92
rect 4077 -126 4111 -92
rect 4111 -126 4121 -92
rect 4285 -126 4295 -92
rect 4295 -126 4337 -92
rect 4566 -126 4571 -92
rect 4571 -126 4618 -92
rect 4786 -126 4813 -92
rect 4813 -126 4838 -92
rect 4991 -126 4997 -92
rect 4997 -126 5031 -92
rect 5031 -126 5043 -92
rect 5212 -126 5215 -92
rect 5215 -126 5264 -92
rect 5417 -126 5457 -92
rect 5457 -126 5469 -92
rect 5626 -126 5641 -92
rect 5641 -126 5675 -92
rect 5675 -126 5678 -92
rect 5843 -126 5859 -92
rect 5859 -126 5895 -92
rect 6057 -126 6101 -92
rect 6101 -126 6109 -92
rect 6252 -126 6285 -92
rect 6285 -126 6304 -92
rect 6447 -126 6469 -92
rect 6469 -126 6499 -92
rect 6649 -126 6653 -92
rect 6653 -126 6687 -92
rect 6687 -126 6701 -92
rect 6933 -126 6963 -92
rect 6963 -126 6985 -92
rect 7132 -126 7147 -92
rect 7147 -126 7184 -92
rect 2574 -129 2626 -126
rect 2837 -133 2889 -126
rect 3045 -132 3097 -126
rect 3255 -135 3307 -126
rect 3455 -129 3507 -126
rect 3658 -132 3710 -126
rect 3868 -132 3920 -126
rect 4069 -131 4121 -126
rect 4285 -130 4337 -126
rect 4566 -132 4618 -126
rect 4786 -137 4838 -126
rect 4991 -136 5043 -126
rect 5212 -130 5264 -126
rect 5417 -137 5469 -126
rect 5626 -136 5678 -126
rect 5843 -136 5895 -126
rect 6057 -131 6109 -126
rect 6252 -133 6304 -126
rect 6447 -136 6499 -126
rect 6649 -133 6701 -126
rect 6933 -132 6985 -126
rect 7132 -131 7184 -126
rect 7335 -129 7387 -77
rect 7600 -92 7652 -80
rect 7798 -92 7850 -81
rect 7987 -92 8039 -79
rect 8199 -92 8251 -79
rect 8416 -92 8468 -79
rect 7600 -126 7607 -92
rect 7607 -126 7652 -92
rect 7798 -126 7849 -92
rect 7849 -126 7850 -92
rect 7987 -126 8033 -92
rect 8033 -126 8039 -92
rect 8199 -126 8217 -92
rect 8217 -126 8251 -92
rect 8416 -126 8435 -92
rect 8435 -126 8468 -92
rect 7600 -132 7652 -126
rect 7798 -133 7850 -126
rect 7987 -131 8039 -126
rect 8199 -131 8251 -126
rect 8416 -131 8468 -126
rect 8621 -135 8673 -83
rect 8826 -92 8878 -83
rect 9034 -92 9086 -78
rect 9317 -92 9369 -79
rect 9510 -92 9562 -81
rect 9736 -92 9788 -83
rect 8826 -126 8861 -92
rect 8861 -126 8878 -92
rect 9034 -126 9045 -92
rect 9045 -126 9079 -92
rect 9079 -126 9086 -92
rect 9317 -126 9321 -92
rect 9321 -126 9355 -92
rect 9355 -126 9369 -92
rect 9510 -126 9539 -92
rect 9539 -126 9562 -92
rect 9736 -126 9781 -92
rect 9781 -126 9788 -92
rect 8826 -135 8878 -126
rect 9034 -130 9086 -126
rect 9317 -131 9369 -126
rect 9510 -133 9562 -126
rect 9736 -135 9788 -126
rect 10001 -135 10053 -83
rect 10195 -92 10247 -79
rect 10393 -92 10445 -88
rect 10597 -92 10649 -80
rect 10817 -92 10869 -77
rect 11032 -92 11084 -81
rect 11260 -92 11312 -78
rect 11464 -92 11516 -81
rect 11702 -92 11754 -79
rect 11895 -92 11947 -78
rect 12092 -92 12144 -83
rect 12348 -92 12400 -80
rect 12587 -92 12639 -84
rect 12820 -92 12872 -88
rect 10195 -126 10241 -92
rect 10241 -126 10247 -92
rect 10393 -126 10425 -92
rect 10425 -126 10445 -92
rect 10597 -126 10609 -92
rect 10609 -126 10643 -92
rect 10643 -126 10649 -92
rect 10817 -126 10827 -92
rect 10827 -126 10869 -92
rect 11032 -126 11069 -92
rect 11069 -126 11084 -92
rect 11260 -126 11287 -92
rect 11287 -126 11312 -92
rect 11464 -126 11471 -92
rect 11471 -126 11516 -92
rect 11702 -126 11713 -92
rect 11713 -126 11747 -92
rect 11747 -126 11754 -92
rect 11895 -126 11897 -92
rect 11897 -126 11931 -92
rect 11931 -126 11947 -92
rect 12092 -126 12115 -92
rect 12115 -126 12144 -92
rect 12348 -126 12357 -92
rect 12357 -126 12391 -92
rect 12391 -126 12400 -92
rect 12587 -126 12633 -92
rect 12633 -126 12639 -92
rect 12820 -126 12851 -92
rect 12851 -126 12872 -92
rect 10195 -131 10247 -126
rect 10393 -140 10445 -126
rect 10597 -132 10649 -126
rect 10817 -129 10869 -126
rect 11032 -133 11084 -126
rect 11260 -130 11312 -126
rect 11464 -133 11516 -126
rect 11702 -131 11754 -126
rect 11895 -130 11947 -126
rect 12092 -135 12144 -126
rect 12348 -132 12400 -126
rect 12587 -136 12639 -126
rect 12820 -140 12872 -126
rect 13041 -135 13093 -83
rect 13232 -92 13284 -83
rect 13460 -92 13512 -81
rect 13657 -92 13709 -86
rect 13232 -126 13277 -92
rect 13277 -126 13284 -92
rect 13460 -126 13461 -92
rect 13461 -126 13495 -92
rect 13495 -126 13512 -92
rect 13657 -126 13679 -92
rect 13679 -126 13709 -92
rect 13232 -135 13284 -126
rect 13460 -133 13512 -126
rect 13657 -138 13709 -126
rect 13869 -138 13921 -86
rect 14096 -92 14148 -83
rect 14285 -92 14337 -82
rect 14096 -126 14105 -92
rect 14105 -126 14139 -92
rect 14139 -126 14148 -92
rect 14285 -126 14289 -92
rect 14289 -126 14323 -92
rect 14323 -126 14337 -92
rect 14096 -135 14148 -126
rect 14285 -134 14337 -126
rect 14511 -133 14563 -81
rect 14765 -92 14817 -81
rect 15009 -92 15061 -84
rect 15239 -92 15291 -85
rect 15497 -92 15549 -82
rect 14765 -126 14783 -92
rect 14783 -126 14817 -92
rect 15009 -126 15025 -92
rect 15025 -126 15059 -92
rect 15059 -126 15061 -92
rect 15239 -126 15243 -92
rect 15243 -126 15291 -92
rect 15497 -126 15519 -92
rect 15519 -126 15549 -92
rect 14765 -133 14817 -126
rect 15009 -136 15061 -126
rect 15239 -137 15291 -126
rect 15497 -134 15549 -126
rect 15707 -134 15759 -82
rect 15932 -92 15984 -82
rect 16151 -92 16203 -85
rect 16497 -92 16549 -81
rect 16696 -92 16748 -84
rect 15932 -126 15945 -92
rect 15945 -126 15979 -92
rect 15979 -126 15984 -92
rect 16151 -126 16163 -92
rect 16163 -126 16203 -92
rect 16497 -126 16531 -92
rect 16531 -126 16549 -92
rect 16696 -126 16715 -92
rect 16715 -126 16748 -92
rect 15932 -134 15984 -126
rect 16151 -137 16203 -126
rect 16497 -133 16549 -126
rect 16696 -136 16748 -126
<< metal2 >>
rect 51 2978 107 2987
rect 51 2913 107 2922
rect 17 1834 73 1843
rect 17 1769 73 1778
rect 17 1414 71 1420
rect 17 1362 18 1414
rect 70 1362 71 1414
rect 17 1356 71 1362
rect 23 875 65 1356
rect 17 869 71 875
rect 17 817 18 869
rect 70 817 71 869
rect 17 811 71 817
rect 45 458 101 467
rect 45 393 101 402
rect 17 350 69 356
rect 141 346 183 3300
rect 253 2980 309 2989
rect 253 2915 309 2924
rect 464 2978 520 2987
rect 464 2913 520 2922
rect 654 2978 710 2987
rect 654 2913 710 2922
rect 862 2980 918 2989
rect 862 2915 918 2924
rect 1064 2980 1120 2989
rect 1064 2915 1120 2924
rect 1263 2982 1319 2991
rect 1263 2917 1319 2926
rect 1458 2979 1514 2988
rect 1458 2914 1514 2923
rect 1169 2439 1225 2448
rect 1169 2374 1225 2383
rect 1388 2443 1444 2452
rect 1388 2378 1444 2387
rect 1018 2250 1024 2303
rect 1077 2250 1083 2303
rect 1018 2249 1083 2250
rect 467 2039 474 2091
rect 526 2039 533 2091
rect 257 1832 313 1841
rect 257 1767 313 1776
rect 482 1617 519 2039
rect 579 1831 635 1840
rect 579 1766 635 1775
rect 797 1832 853 1841
rect 797 1767 853 1776
rect 468 1565 475 1617
rect 527 1565 534 1617
rect 349 1400 356 1452
rect 408 1400 414 1452
rect 263 1151 319 1160
rect 263 1086 319 1095
rect 362 894 404 1400
rect 465 1147 521 1156
rect 465 1082 521 1091
rect 654 1144 710 1153
rect 654 1079 710 1088
rect 883 1145 939 1154
rect 883 1080 939 1089
rect 351 841 357 894
rect 409 841 416 894
rect 351 840 416 841
rect 1030 776 1072 2249
rect 1562 1603 1604 3300
rect 1659 2981 1715 2990
rect 1659 2916 1715 2925
rect 1876 2979 1932 2988
rect 1876 2914 1932 2923
rect 1671 2443 1727 2452
rect 1671 2378 1727 2387
rect 1880 2443 1936 2452
rect 1880 2378 1936 2387
rect 1729 2039 1736 2091
rect 1788 2039 1795 2091
rect 1744 1617 1781 2039
rect 1551 1550 1557 1603
rect 1609 1550 1616 1603
rect 1730 1565 1737 1617
rect 1789 1565 1796 1617
rect 1551 1549 1616 1550
rect 1964 1453 2006 3300
rect 2150 2982 2206 2991
rect 2150 2917 2206 2926
rect 2151 2441 2207 2450
rect 2151 2376 2207 2385
rect 1950 1401 1957 1453
rect 2009 1401 2015 1453
rect 1208 1296 1264 1305
rect 1208 1231 1264 1240
rect 1425 1296 1481 1305
rect 1425 1231 1481 1240
rect 1644 1296 1700 1305
rect 1644 1231 1700 1240
rect 1857 1292 1913 1301
rect 1857 1227 1913 1236
rect 1024 770 1078 776
rect 1024 718 1025 770
rect 1077 718 1078 770
rect 1024 712 1078 718
rect 278 454 334 463
rect 278 389 334 398
rect 493 461 549 470
rect 493 396 549 405
rect 711 458 767 467
rect 711 393 767 402
rect 927 459 983 468
rect 927 394 983 403
rect 69 304 183 346
rect 1030 314 1072 712
rect 1419 614 1475 623
rect 1190 602 1246 611
rect 1419 549 1475 558
rect 1638 604 1694 613
rect 1190 537 1246 546
rect 1638 539 1694 548
rect 1830 608 1886 617
rect 1830 543 1886 552
rect 17 292 69 298
rect 297 286 349 292
rect 1019 262 1025 314
rect 1077 262 1083 314
rect 297 228 349 234
rect 301 -343 343 228
rect 1964 160 2006 1401
rect 2188 1362 2194 1414
rect 2246 1362 2254 1414
rect 2068 1292 2124 1301
rect 2068 1227 2124 1236
rect 2042 965 2094 971
rect 2042 907 2094 913
rect 1953 107 1959 160
rect 2011 107 2018 160
rect 1953 106 2018 107
rect 419 -74 475 -65
rect 419 -139 475 -130
rect 618 -77 674 -68
rect 618 -142 674 -133
rect 829 -77 885 -68
rect 829 -142 885 -133
rect 1035 -77 1091 -68
rect 1035 -142 1091 -133
rect 1263 -79 1319 -70
rect 1263 -144 1319 -135
rect 1507 -79 1563 -70
rect 1507 -144 1563 -135
rect 1737 -77 1793 -68
rect 1737 -142 1793 -133
rect 1943 -77 1999 -68
rect 1943 -142 1999 -133
rect 2046 -343 2088 907
rect 2200 215 2242 1362
rect 2330 1048 2372 3300
rect 2427 2975 2483 2984
rect 2427 2910 2483 2919
rect 2409 1414 2463 1420
rect 2409 1362 2410 1414
rect 2462 1362 2463 1414
rect 2409 1356 2463 1362
rect 2324 1042 2376 1048
rect 2324 984 2376 990
rect 2415 875 2457 1356
rect 2409 869 2463 875
rect 2409 817 2410 869
rect 2462 817 2463 869
rect 2409 811 2463 817
rect 2324 606 2380 615
rect 2324 541 2380 550
rect 2409 350 2461 356
rect 2533 346 2575 3300
rect 2650 2978 2706 2987
rect 2650 2913 2706 2922
rect 2882 2977 2938 2986
rect 2882 2912 2938 2921
rect 2860 2622 2866 2674
rect 2918 2622 2924 2674
rect 2866 2302 2918 2622
rect 2860 2250 2866 2302
rect 2918 2250 2924 2302
rect 3412 2256 3418 2309
rect 3471 2256 3477 2309
rect 3412 2255 3477 2256
rect 2860 2038 2867 2090
rect 2919 2038 2926 2090
rect 2701 1836 2757 1845
rect 2701 1771 2757 1780
rect 2875 1616 2912 2038
rect 3026 1838 3082 1847
rect 3026 1773 3082 1782
rect 3294 1838 3350 1847
rect 3294 1773 3350 1782
rect 2861 1564 2868 1616
rect 2920 1564 2927 1616
rect 2741 1400 2748 1452
rect 2800 1400 2806 1452
rect 2652 1148 2708 1157
rect 2652 1083 2708 1092
rect 2754 894 2796 1400
rect 2867 1145 2923 1154
rect 3260 1152 3316 1161
rect 2867 1080 2923 1089
rect 3065 1142 3121 1151
rect 3260 1087 3316 1096
rect 3065 1077 3121 1086
rect 2743 841 2749 894
rect 2801 841 2808 894
rect 2743 840 2808 841
rect 3424 776 3466 2255
rect 3560 1838 3616 1847
rect 3560 1773 3616 1782
rect 3800 1836 3856 1845
rect 3800 1771 3856 1780
rect 3954 1602 3996 3300
rect 4226 2439 4282 2448
rect 4226 2374 4282 2383
rect 4121 2039 4128 2091
rect 4180 2039 4187 2091
rect 4136 1617 4173 2039
rect 3943 1549 3949 1602
rect 4001 1549 4008 1602
rect 4122 1565 4129 1617
rect 4181 1565 4188 1617
rect 3943 1548 4008 1549
rect 4356 1453 4398 3300
rect 4518 2974 4574 2983
rect 4518 2909 4574 2918
rect 4475 2442 4531 2451
rect 4475 2377 4531 2386
rect 4342 1401 4349 1453
rect 4401 1401 4407 1453
rect 4192 1292 4248 1301
rect 4192 1227 4248 1236
rect 3540 1150 3596 1159
rect 3540 1085 3596 1094
rect 3759 1148 3815 1157
rect 3759 1083 3815 1092
rect 3417 770 3471 776
rect 3417 718 3418 770
rect 3470 718 3471 770
rect 3417 712 3471 718
rect 2648 455 2704 464
rect 2648 390 2704 399
rect 2838 455 2894 464
rect 2838 390 2894 399
rect 3048 458 3104 467
rect 3048 393 3104 402
rect 3265 455 3321 464
rect 3265 390 3321 399
rect 2461 304 2575 346
rect 3422 315 3464 712
rect 4116 605 4172 614
rect 4116 540 4172 549
rect 3560 458 3616 467
rect 3560 393 3616 402
rect 3784 463 3840 472
rect 3784 398 3840 407
rect 2409 292 2461 298
rect 2689 286 2741 292
rect 3411 263 3417 315
rect 3469 263 3475 315
rect 2689 228 2741 234
rect 2200 175 2304 215
rect 2298 163 2304 175
rect 2358 163 2364 215
rect 2161 -72 2217 -63
rect 2161 -137 2217 -128
rect 2364 -78 2420 -69
rect 2364 -143 2420 -134
rect 2572 -75 2628 -66
rect 2572 -140 2628 -131
rect 2693 -343 2735 228
rect 4356 160 4398 1401
rect 4582 1362 4588 1414
rect 4640 1362 4648 1414
rect 4470 1291 4526 1300
rect 4470 1226 4526 1235
rect 4434 966 4486 972
rect 4434 908 4486 914
rect 4345 107 4351 160
rect 4403 107 4410 160
rect 4345 106 4410 107
rect 2835 -79 2891 -70
rect 2835 -144 2891 -135
rect 3043 -78 3099 -69
rect 3043 -143 3099 -134
rect 3253 -81 3309 -72
rect 3253 -146 3309 -137
rect 3453 -75 3509 -66
rect 3453 -140 3509 -131
rect 3656 -78 3712 -69
rect 3656 -143 3712 -134
rect 3866 -78 3922 -69
rect 3866 -143 3922 -134
rect 4067 -77 4123 -68
rect 4067 -142 4123 -133
rect 4283 -76 4339 -67
rect 4283 -141 4339 -132
rect 4438 -343 4480 908
rect 4509 603 4565 612
rect 4509 538 4565 547
rect 4594 215 4636 1362
rect 4722 1048 4764 3300
rect 4826 2975 4882 2984
rect 4826 2910 4882 2919
rect 4819 2428 4875 2437
rect 4819 2363 4875 2372
rect 4801 1414 4855 1420
rect 4801 1362 4802 1414
rect 4854 1362 4855 1414
rect 4801 1356 4855 1362
rect 4716 1042 4768 1048
rect 4716 984 4768 990
rect 4807 875 4849 1356
rect 4801 869 4855 875
rect 4801 817 4802 869
rect 4854 817 4855 869
rect 4801 811 4855 817
rect 4706 611 4762 620
rect 4706 546 4762 555
rect 4802 350 4854 356
rect 4926 346 4968 3300
rect 5026 2976 5082 2985
rect 5026 2911 5082 2920
rect 5245 2975 5301 2984
rect 5245 2910 5301 2919
rect 5491 2974 5547 2983
rect 5491 2909 5547 2918
rect 5699 2976 5755 2985
rect 5699 2911 5755 2920
rect 5901 2977 5957 2986
rect 5901 2912 5957 2921
rect 6094 2976 6150 2985
rect 6094 2911 6150 2920
rect 5073 2434 5129 2443
rect 5073 2369 5129 2378
rect 5302 2434 5358 2443
rect 5302 2369 5358 2378
rect 5803 2256 5809 2309
rect 5862 2256 5868 2309
rect 5803 2255 5868 2256
rect 5252 2038 5259 2090
rect 5311 2038 5318 2090
rect 5267 1616 5304 2038
rect 5594 1839 5650 1848
rect 5594 1774 5650 1783
rect 5253 1564 5260 1616
rect 5312 1564 5319 1616
rect 5132 1401 5139 1453
rect 5191 1401 5197 1453
rect 5042 1296 5098 1305
rect 5042 1231 5098 1240
rect 5146 895 5188 1401
rect 5281 1296 5337 1305
rect 5281 1231 5337 1240
rect 5580 1145 5636 1154
rect 5580 1080 5636 1089
rect 5135 842 5141 895
rect 5193 842 5200 895
rect 5135 841 5200 842
rect 5815 776 5857 2255
rect 5960 1842 6016 1851
rect 5960 1777 6016 1786
rect 6204 1842 6260 1851
rect 6204 1777 6260 1786
rect 6344 1602 6386 3300
rect 6466 2975 6522 2984
rect 6466 2910 6522 2919
rect 6655 2973 6711 2982
rect 6655 2908 6711 2917
rect 6512 2040 6519 2092
rect 6571 2040 6578 2092
rect 6527 1853 6564 2040
rect 6521 1819 6564 1853
rect 6527 1618 6564 1819
rect 6627 1833 6683 1842
rect 6627 1768 6683 1777
rect 6333 1549 6339 1602
rect 6391 1549 6398 1602
rect 6513 1566 6520 1618
rect 6572 1566 6579 1618
rect 6333 1548 6398 1549
rect 6747 1454 6789 3300
rect 6945 2973 7001 2982
rect 6945 2908 7001 2917
rect 7020 2439 7076 2448
rect 7020 2374 7076 2383
rect 6733 1402 6740 1454
rect 6792 1402 6798 1454
rect 5931 1142 5987 1151
rect 5931 1077 5987 1086
rect 6120 1140 6176 1149
rect 6120 1075 6176 1084
rect 6325 1147 6381 1156
rect 6325 1082 6381 1091
rect 6516 1149 6572 1158
rect 6516 1084 6572 1093
rect 5809 770 5863 776
rect 5809 718 5810 770
rect 5862 718 5863 770
rect 5809 712 5863 718
rect 5036 613 5092 622
rect 5036 548 5092 557
rect 5232 613 5288 622
rect 5232 548 5288 557
rect 5662 456 5718 465
rect 5662 391 5718 400
rect 4854 304 4968 346
rect 5814 314 5856 712
rect 5962 454 6018 463
rect 5962 389 6018 398
rect 6214 458 6270 467
rect 6214 393 6270 402
rect 6431 463 6487 472
rect 6431 398 6487 407
rect 6632 460 6688 469
rect 6632 395 6688 404
rect 4802 292 4854 298
rect 5080 286 5132 292
rect 5803 262 5809 314
rect 5861 262 5867 314
rect 5080 228 5132 234
rect 4594 175 4698 215
rect 4692 163 4698 175
rect 4752 163 4758 215
rect 4564 -78 4620 -69
rect 4564 -143 4620 -134
rect 4784 -83 4840 -74
rect 4784 -148 4840 -139
rect 4989 -82 5045 -73
rect 4989 -147 5045 -138
rect 5084 -343 5126 228
rect 6747 161 6789 1402
rect 6972 1364 6978 1416
rect 7030 1364 7038 1416
rect 6825 966 6877 972
rect 6825 908 6877 914
rect 6736 160 6801 161
rect 6736 108 6742 160
rect 6794 108 6801 160
rect 6736 107 6801 108
rect 5210 -76 5266 -67
rect 5210 -141 5266 -132
rect 5415 -83 5471 -74
rect 5415 -148 5471 -139
rect 5624 -82 5680 -73
rect 5624 -147 5680 -138
rect 5841 -82 5897 -73
rect 5841 -147 5897 -138
rect 6055 -77 6111 -68
rect 6055 -142 6111 -133
rect 6250 -79 6306 -70
rect 6250 -144 6306 -135
rect 6445 -82 6501 -73
rect 6445 -147 6501 -138
rect 6647 -79 6703 -70
rect 6647 -144 6703 -135
rect 6829 -343 6871 908
rect 6984 217 7026 1364
rect 7114 1048 7156 3300
rect 7218 2975 7274 2984
rect 7218 2910 7274 2919
rect 7224 2441 7280 2450
rect 7224 2376 7280 2385
rect 7193 1414 7247 1420
rect 7193 1362 7194 1414
rect 7246 1362 7247 1414
rect 7193 1356 7247 1362
rect 7108 1042 7160 1048
rect 7108 984 7160 990
rect 7199 875 7241 1356
rect 7193 869 7247 875
rect 7193 817 7194 869
rect 7246 817 7247 869
rect 7193 811 7247 817
rect 7139 606 7195 615
rect 7139 541 7195 550
rect 7193 350 7245 356
rect 7317 346 7359 3300
rect 7421 2622 7427 2674
rect 7479 2622 7485 2674
rect 7427 2090 7479 2622
rect 7547 2439 7603 2448
rect 7547 2374 7603 2383
rect 8194 2256 8200 2309
rect 8253 2256 8259 2309
rect 8194 2255 8259 2256
rect 7421 2038 7427 2090
rect 7479 2038 7485 2090
rect 7644 2039 7651 2091
rect 7703 2039 7710 2091
rect 7659 1617 7696 2039
rect 7645 1565 7652 1617
rect 7704 1565 7711 1617
rect 7525 1400 7532 1452
rect 7584 1400 7590 1452
rect 7439 1294 7495 1303
rect 7439 1229 7495 1238
rect 7538 895 7580 1400
rect 7666 1299 7722 1308
rect 7666 1234 7722 1243
rect 7856 1301 7912 1310
rect 7856 1236 7912 1245
rect 8072 1292 8128 1301
rect 8072 1227 8128 1236
rect 7527 842 7533 895
rect 7585 842 7592 895
rect 7527 841 7592 842
rect 8206 776 8248 2255
rect 8570 1835 8626 1844
rect 8570 1770 8626 1779
rect 8738 1603 8780 3300
rect 8905 2040 8912 2092
rect 8964 2040 8971 2092
rect 8822 1832 8878 1841
rect 8822 1767 8878 1776
rect 8920 1618 8957 2040
rect 9028 1840 9084 1849
rect 9028 1775 9084 1784
rect 8727 1550 8733 1603
rect 8785 1550 8792 1603
rect 8906 1566 8913 1618
rect 8965 1566 8972 1618
rect 8727 1549 8792 1550
rect 9140 1453 9182 3300
rect 9311 1834 9367 1843
rect 9311 1769 9367 1778
rect 9126 1401 9133 1453
rect 9185 1401 9191 1453
rect 8561 1151 8617 1160
rect 8561 1086 8617 1095
rect 8751 1153 8807 1162
rect 8751 1088 8807 1097
rect 8945 1151 9001 1160
rect 8945 1086 9001 1095
rect 8201 770 8255 776
rect 8201 718 8202 770
rect 8254 718 8255 770
rect 8201 712 8255 718
rect 7440 610 7496 619
rect 7440 545 7496 554
rect 7646 611 7702 620
rect 7646 546 7702 555
rect 7856 607 7912 616
rect 7856 542 7912 551
rect 8067 613 8123 622
rect 8067 548 8123 557
rect 7245 304 7359 346
rect 8206 314 8248 712
rect 8517 451 8573 460
rect 8517 386 8573 395
rect 8709 451 8765 460
rect 8709 386 8765 395
rect 8909 451 8965 460
rect 8909 386 8965 395
rect 7193 292 7245 298
rect 7473 286 7525 292
rect 8195 262 8201 314
rect 8253 262 8259 314
rect 7473 228 7525 234
rect 6984 177 7088 217
rect 7082 165 7088 177
rect 7142 165 7148 217
rect 6931 -78 6987 -69
rect 6931 -143 6987 -134
rect 7130 -77 7186 -68
rect 7130 -142 7186 -133
rect 7333 -75 7389 -66
rect 7333 -140 7389 -131
rect 7477 -343 7519 228
rect 9140 160 9182 1401
rect 9364 1362 9370 1414
rect 9422 1362 9430 1414
rect 9256 1147 9312 1156
rect 9256 1082 9312 1091
rect 9218 967 9270 973
rect 9218 909 9270 915
rect 9129 107 9135 160
rect 9187 107 9194 160
rect 9129 106 9194 107
rect 7598 -78 7654 -69
rect 7598 -143 7654 -134
rect 7796 -79 7852 -70
rect 7796 -144 7852 -135
rect 7985 -77 8041 -68
rect 7985 -142 8041 -133
rect 8197 -77 8253 -68
rect 8197 -142 8253 -133
rect 8414 -77 8470 -68
rect 8414 -142 8470 -133
rect 8619 -81 8675 -72
rect 8619 -146 8675 -137
rect 8824 -81 8880 -72
rect 8824 -146 8880 -137
rect 9032 -76 9088 -67
rect 9032 -141 9088 -132
rect 9222 -343 9264 909
rect 9376 215 9418 1362
rect 9506 1048 9548 3300
rect 9609 1835 9665 1844
rect 9609 1770 9665 1779
rect 9584 1415 9638 1421
rect 9584 1363 9585 1415
rect 9637 1363 9638 1415
rect 9584 1357 9638 1363
rect 9500 1042 9552 1048
rect 9500 984 9552 990
rect 9590 876 9632 1357
rect 9584 870 9638 876
rect 9584 818 9585 870
rect 9637 818 9638 870
rect 9584 812 9638 818
rect 9527 459 9583 468
rect 9527 394 9583 403
rect 9585 349 9637 355
rect 9709 345 9751 3300
rect 10586 2256 10592 2309
rect 10645 2256 10651 2309
rect 10586 2255 10651 2256
rect 10035 2038 10042 2090
rect 10094 2038 10101 2090
rect 10050 1616 10087 2038
rect 10036 1564 10043 1616
rect 10095 1564 10102 1616
rect 9917 1401 9924 1453
rect 9976 1401 9982 1453
rect 9930 894 9972 1401
rect 10053 1295 10109 1304
rect 10053 1230 10109 1239
rect 10282 1298 10338 1307
rect 10282 1233 10338 1242
rect 10508 1303 10564 1312
rect 10508 1238 10564 1247
rect 9919 841 9925 894
rect 9977 841 9984 894
rect 9919 840 9984 841
rect 10598 776 10640 2255
rect 11130 1602 11172 3300
rect 11298 2040 11305 2092
rect 11357 2040 11364 2092
rect 11313 1618 11350 2040
rect 11441 1836 11497 1845
rect 11441 1771 11497 1780
rect 11119 1549 11125 1602
rect 11177 1549 11184 1602
rect 11299 1566 11306 1618
rect 11358 1566 11365 1618
rect 11119 1548 11184 1549
rect 11531 1454 11573 3300
rect 11651 1838 11707 1847
rect 11651 1773 11707 1782
rect 11518 1402 11525 1454
rect 11577 1402 11583 1454
rect 10736 1295 10792 1304
rect 10736 1230 10792 1239
rect 10972 1301 11028 1310
rect 10972 1236 11028 1245
rect 11164 1292 11220 1301
rect 11164 1227 11220 1236
rect 11439 1146 11495 1155
rect 11439 1081 11495 1090
rect 10592 770 10646 776
rect 10592 718 10593 770
rect 10645 718 10646 770
rect 10592 710 10646 718
rect 9947 602 10003 611
rect 9947 537 10003 546
rect 10204 609 10260 618
rect 10204 544 10260 553
rect 10454 605 10510 614
rect 10454 540 10510 549
rect 9637 303 9751 345
rect 10598 314 10640 710
rect 10725 610 10781 619
rect 10725 545 10781 554
rect 10966 613 11022 622
rect 10966 548 11022 557
rect 11191 609 11247 618
rect 11191 544 11247 553
rect 11428 455 11484 464
rect 11428 390 11484 399
rect 9585 291 9637 297
rect 9865 286 9917 292
rect 10587 262 10593 314
rect 10645 262 10651 314
rect 9865 228 9917 234
rect 9376 175 9480 215
rect 9474 163 9480 175
rect 9534 163 9540 215
rect 9315 -77 9371 -68
rect 9315 -142 9371 -133
rect 9508 -79 9564 -70
rect 9508 -144 9564 -135
rect 9734 -81 9790 -72
rect 9734 -146 9790 -137
rect 9869 -343 9911 228
rect 11531 160 11573 1402
rect 11756 1364 11762 1416
rect 11814 1364 11822 1416
rect 11643 1146 11699 1155
rect 11643 1081 11699 1090
rect 11609 966 11661 972
rect 11609 908 11661 914
rect 11520 107 11526 160
rect 11578 107 11585 160
rect 11520 106 11585 107
rect 9999 -81 10055 -72
rect 9999 -146 10055 -137
rect 10193 -77 10249 -68
rect 10193 -142 10249 -133
rect 10391 -86 10447 -77
rect 10391 -151 10447 -142
rect 10595 -78 10651 -69
rect 10595 -143 10651 -134
rect 10815 -75 10871 -66
rect 10815 -140 10871 -131
rect 11030 -79 11086 -70
rect 11030 -144 11086 -135
rect 11258 -76 11314 -67
rect 11258 -141 11314 -132
rect 11462 -79 11518 -70
rect 11462 -144 11518 -135
rect 11613 -343 11655 908
rect 11684 455 11740 464
rect 11684 390 11740 399
rect 11768 217 11810 1364
rect 11898 1048 11940 3300
rect 12002 1836 12058 1845
rect 12002 1771 12058 1780
rect 11976 1414 12030 1420
rect 11976 1362 11977 1414
rect 12029 1362 12030 1414
rect 11976 1356 12030 1362
rect 11892 1042 11944 1048
rect 11892 984 11944 990
rect 11982 875 12024 1356
rect 11976 869 12030 875
rect 11976 817 11977 869
rect 12029 817 12030 869
rect 11976 811 12030 817
rect 11919 455 11975 464
rect 11919 390 11975 399
rect 11978 351 12030 357
rect 12102 347 12144 3300
rect 12977 2256 12983 2309
rect 13036 2256 13042 2309
rect 12977 2255 13042 2256
rect 12427 2037 12434 2089
rect 12486 2037 12493 2089
rect 12282 1836 12338 1845
rect 12282 1771 12338 1780
rect 12442 1615 12479 2037
rect 12599 1835 12655 1844
rect 12599 1770 12655 1779
rect 12428 1563 12435 1615
rect 12487 1563 12494 1615
rect 12309 1401 12316 1453
rect 12368 1401 12374 1453
rect 12208 1142 12264 1151
rect 12208 1077 12264 1086
rect 12322 895 12364 1401
rect 12899 1292 12955 1301
rect 12899 1227 12955 1236
rect 12447 1144 12503 1153
rect 12447 1079 12503 1088
rect 12651 1144 12707 1153
rect 12651 1079 12707 1088
rect 12311 842 12317 895
rect 12369 842 12376 895
rect 12311 841 12376 842
rect 12989 776 13031 2255
rect 13519 1602 13561 3300
rect 13687 2040 13694 2092
rect 13746 2040 13753 2092
rect 13702 1618 13739 2040
rect 13508 1549 13514 1602
rect 13566 1549 13573 1602
rect 13688 1566 13695 1618
rect 13747 1566 13754 1618
rect 13508 1548 13573 1549
rect 13924 1454 13966 3300
rect 13910 1402 13917 1454
rect 13969 1402 13975 1454
rect 13103 1297 13159 1306
rect 13103 1232 13159 1241
rect 13294 1292 13350 1301
rect 13294 1227 13350 1236
rect 13496 1291 13552 1300
rect 13496 1226 13552 1235
rect 13786 1292 13842 1301
rect 13786 1227 13842 1236
rect 12984 770 13038 776
rect 12984 718 12985 770
rect 13037 718 13038 770
rect 12984 712 13038 718
rect 12898 607 12954 616
rect 12898 542 12954 551
rect 12208 457 12264 466
rect 12208 392 12264 401
rect 12398 455 12454 464
rect 12398 390 12454 399
rect 12602 457 12658 466
rect 12602 392 12658 401
rect 12030 305 12144 347
rect 12990 315 13032 712
rect 13099 608 13155 617
rect 13099 543 13155 552
rect 13317 604 13373 613
rect 13317 539 13373 548
rect 13524 608 13580 617
rect 13524 543 13580 552
rect 13729 607 13785 616
rect 13729 542 13785 551
rect 11978 293 12030 299
rect 12256 287 12308 293
rect 12979 263 12985 315
rect 13037 263 13043 315
rect 12256 229 12308 235
rect 11768 177 11872 217
rect 11866 165 11872 177
rect 11926 165 11932 217
rect 11700 -77 11756 -68
rect 11700 -142 11756 -133
rect 11893 -76 11949 -67
rect 11893 -141 11949 -132
rect 12090 -81 12146 -72
rect 12090 -146 12146 -137
rect 12260 -343 12302 229
rect 13924 160 13966 1402
rect 14148 1362 14154 1414
rect 14206 1362 14214 1414
rect 14071 1291 14127 1300
rect 14071 1226 14127 1235
rect 14002 965 14054 971
rect 14002 907 14054 913
rect 13913 107 13919 160
rect 13971 107 13978 160
rect 13913 106 13978 107
rect 12346 -78 12402 -69
rect 12346 -143 12402 -134
rect 12585 -82 12641 -73
rect 12585 -147 12641 -138
rect 12818 -86 12874 -77
rect 12818 -151 12874 -142
rect 13039 -81 13095 -72
rect 13039 -146 13095 -137
rect 13230 -81 13286 -72
rect 13230 -146 13286 -137
rect 13458 -79 13514 -70
rect 13458 -144 13514 -135
rect 13655 -84 13711 -75
rect 13655 -149 13711 -140
rect 13867 -84 13923 -75
rect 13867 -149 13923 -140
rect 14006 -343 14048 907
rect 14076 603 14132 612
rect 14076 538 14132 547
rect 14160 215 14202 1362
rect 14290 1048 14332 3300
rect 14389 1833 14445 1842
rect 14389 1768 14445 1777
rect 14369 1415 14423 1421
rect 14369 1363 14370 1415
rect 14422 1363 14423 1415
rect 14369 1357 14423 1363
rect 14284 1042 14336 1048
rect 14284 984 14336 990
rect 14375 876 14417 1357
rect 14369 870 14423 876
rect 14369 818 14370 870
rect 14422 818 14423 870
rect 14369 812 14423 818
rect 14388 463 14444 472
rect 14388 398 14444 407
rect 14369 351 14421 357
rect 14493 347 14535 3300
rect 15370 2256 15376 2309
rect 15429 2256 15435 2309
rect 15370 2255 15435 2256
rect 14819 2038 14826 2090
rect 14878 2038 14885 2090
rect 14684 1833 14740 1842
rect 14684 1768 14740 1777
rect 14834 1616 14871 2038
rect 14971 1833 15027 1842
rect 14971 1768 15027 1777
rect 15261 1833 15317 1842
rect 15261 1768 15317 1777
rect 14820 1564 14827 1616
rect 14879 1564 14886 1616
rect 14704 1401 14711 1453
rect 14763 1401 14769 1453
rect 14611 1152 14667 1161
rect 14611 1087 14667 1096
rect 14715 894 14757 1401
rect 14844 1150 14900 1159
rect 14844 1085 14900 1094
rect 15051 1148 15107 1157
rect 15051 1083 15107 1092
rect 15260 1150 15316 1159
rect 15260 1085 15316 1094
rect 14704 841 14710 894
rect 14762 841 14769 894
rect 14704 840 14769 841
rect 15382 776 15424 2255
rect 15545 1836 15601 1845
rect 15545 1771 15601 1780
rect 15914 1603 15956 3300
rect 16082 2040 16089 2092
rect 16141 2040 16148 2092
rect 16097 1618 16134 2040
rect 15903 1550 15909 1603
rect 15961 1550 15968 1603
rect 16083 1566 16090 1618
rect 16142 1566 16149 1618
rect 15903 1549 15968 1550
rect 16317 1454 16359 3300
rect 16305 1402 16312 1454
rect 16364 1402 16370 1454
rect 15826 1296 15882 1305
rect 15826 1231 15882 1240
rect 16020 1300 16076 1309
rect 16020 1235 16076 1244
rect 16209 1297 16265 1306
rect 16209 1232 16265 1241
rect 15540 1152 15596 1161
rect 15540 1087 15596 1096
rect 15376 770 15430 776
rect 15376 718 15377 770
rect 15429 718 15430 770
rect 15376 712 15430 718
rect 14630 459 14686 468
rect 14630 394 14686 403
rect 14830 458 14886 467
rect 14830 393 14886 402
rect 15020 466 15076 475
rect 15020 401 15076 410
rect 15241 464 15297 473
rect 15241 399 15297 408
rect 14421 305 14535 347
rect 15382 315 15424 712
rect 15828 607 15884 616
rect 15828 542 15884 551
rect 16019 610 16075 619
rect 16019 545 16075 554
rect 16214 612 16270 621
rect 16214 547 16270 556
rect 15537 459 15593 468
rect 15537 394 15593 403
rect 14369 293 14421 299
rect 14649 286 14701 292
rect 15371 263 15377 315
rect 15429 263 15435 315
rect 14649 228 14701 234
rect 14160 175 14264 215
rect 14258 163 14264 175
rect 14318 163 14324 215
rect 14094 -81 14150 -72
rect 14094 -146 14150 -137
rect 14283 -80 14339 -71
rect 14283 -145 14339 -136
rect 14509 -79 14565 -70
rect 14509 -144 14565 -135
rect 14653 -343 14695 228
rect 16317 160 16359 1402
rect 16540 1364 16546 1416
rect 16598 1364 16606 1416
rect 16432 1299 16488 1308
rect 16432 1234 16488 1243
rect 16395 967 16447 973
rect 16395 909 16447 915
rect 16306 107 16312 160
rect 16364 107 16371 160
rect 16306 106 16371 107
rect 14763 -79 14819 -70
rect 14763 -144 14819 -135
rect 15007 -82 15063 -73
rect 15007 -147 15063 -138
rect 15237 -83 15293 -74
rect 15237 -148 15293 -139
rect 15495 -80 15551 -71
rect 15495 -145 15551 -136
rect 15705 -80 15761 -71
rect 15705 -145 15761 -136
rect 15930 -80 15986 -71
rect 15930 -145 15986 -136
rect 16149 -83 16205 -74
rect 16149 -148 16205 -139
rect 16399 -343 16441 909
rect 16552 217 16594 1364
rect 16682 1048 16724 3300
rect 16676 1042 16728 1048
rect 16676 984 16728 990
rect 16661 607 16717 616
rect 16661 542 16717 551
rect 16552 177 16656 217
rect 16650 165 16656 177
rect 16710 165 16716 217
rect 16495 -79 16551 -70
rect 16495 -144 16551 -135
rect 16694 -82 16750 -73
rect 16694 -147 16750 -138
<< via2 >>
rect 51 2976 107 2978
rect 51 2924 53 2976
rect 53 2924 105 2976
rect 105 2924 107 2976
rect 51 2922 107 2924
rect 17 1832 73 1834
rect 17 1780 19 1832
rect 19 1780 71 1832
rect 71 1780 73 1832
rect 17 1778 73 1780
rect 45 456 101 458
rect 45 404 47 456
rect 47 404 99 456
rect 99 404 101 456
rect 45 402 101 404
rect 253 2978 309 2980
rect 253 2926 255 2978
rect 255 2926 307 2978
rect 307 2926 309 2978
rect 253 2924 309 2926
rect 464 2976 520 2978
rect 464 2924 466 2976
rect 466 2924 518 2976
rect 518 2924 520 2976
rect 464 2922 520 2924
rect 654 2976 710 2978
rect 654 2924 656 2976
rect 656 2924 708 2976
rect 708 2924 710 2976
rect 654 2922 710 2924
rect 862 2978 918 2980
rect 862 2926 864 2978
rect 864 2926 916 2978
rect 916 2926 918 2978
rect 862 2924 918 2926
rect 1064 2978 1120 2980
rect 1064 2926 1066 2978
rect 1066 2926 1118 2978
rect 1118 2926 1120 2978
rect 1064 2924 1120 2926
rect 1263 2980 1319 2982
rect 1263 2928 1265 2980
rect 1265 2928 1317 2980
rect 1317 2928 1319 2980
rect 1263 2926 1319 2928
rect 1458 2977 1514 2979
rect 1458 2925 1460 2977
rect 1460 2925 1512 2977
rect 1512 2925 1514 2977
rect 1458 2923 1514 2925
rect 1169 2437 1225 2439
rect 1169 2385 1171 2437
rect 1171 2385 1223 2437
rect 1223 2385 1225 2437
rect 1169 2383 1225 2385
rect 1388 2441 1444 2443
rect 1388 2389 1390 2441
rect 1390 2389 1442 2441
rect 1442 2389 1444 2441
rect 1388 2387 1444 2389
rect 257 1830 313 1832
rect 257 1778 259 1830
rect 259 1778 311 1830
rect 311 1778 313 1830
rect 257 1776 313 1778
rect 579 1829 635 1831
rect 579 1777 581 1829
rect 581 1777 633 1829
rect 633 1777 635 1829
rect 579 1775 635 1777
rect 797 1830 853 1832
rect 797 1778 799 1830
rect 799 1778 851 1830
rect 851 1778 853 1830
rect 797 1776 853 1778
rect 263 1149 319 1151
rect 263 1097 265 1149
rect 265 1097 317 1149
rect 317 1097 319 1149
rect 263 1095 319 1097
rect 465 1145 521 1147
rect 465 1093 467 1145
rect 467 1093 519 1145
rect 519 1093 521 1145
rect 465 1091 521 1093
rect 654 1142 710 1144
rect 654 1090 656 1142
rect 656 1090 708 1142
rect 708 1090 710 1142
rect 654 1088 710 1090
rect 883 1143 939 1145
rect 883 1091 885 1143
rect 885 1091 937 1143
rect 937 1091 939 1143
rect 883 1089 939 1091
rect 1659 2979 1715 2981
rect 1659 2927 1661 2979
rect 1661 2927 1713 2979
rect 1713 2927 1715 2979
rect 1659 2925 1715 2927
rect 1876 2977 1932 2979
rect 1876 2925 1878 2977
rect 1878 2925 1930 2977
rect 1930 2925 1932 2977
rect 1876 2923 1932 2925
rect 1671 2441 1727 2443
rect 1671 2389 1673 2441
rect 1673 2389 1725 2441
rect 1725 2389 1727 2441
rect 1671 2387 1727 2389
rect 1880 2441 1936 2443
rect 1880 2389 1882 2441
rect 1882 2389 1934 2441
rect 1934 2389 1936 2441
rect 1880 2387 1936 2389
rect 2150 2980 2206 2982
rect 2150 2928 2152 2980
rect 2152 2928 2204 2980
rect 2204 2928 2206 2980
rect 2150 2926 2206 2928
rect 2151 2439 2207 2441
rect 2151 2387 2153 2439
rect 2153 2387 2205 2439
rect 2205 2387 2207 2439
rect 2151 2385 2207 2387
rect 1208 1294 1264 1296
rect 1208 1242 1210 1294
rect 1210 1242 1262 1294
rect 1262 1242 1264 1294
rect 1208 1240 1264 1242
rect 1425 1294 1481 1296
rect 1425 1242 1427 1294
rect 1427 1242 1479 1294
rect 1479 1242 1481 1294
rect 1425 1240 1481 1242
rect 1644 1294 1700 1296
rect 1644 1242 1646 1294
rect 1646 1242 1698 1294
rect 1698 1242 1700 1294
rect 1644 1240 1700 1242
rect 1857 1290 1913 1292
rect 1857 1238 1859 1290
rect 1859 1238 1911 1290
rect 1911 1238 1913 1290
rect 1857 1236 1913 1238
rect 278 452 334 454
rect 278 400 280 452
rect 280 400 332 452
rect 332 400 334 452
rect 278 398 334 400
rect 493 459 549 461
rect 493 407 495 459
rect 495 407 547 459
rect 547 407 549 459
rect 493 405 549 407
rect 711 456 767 458
rect 711 404 713 456
rect 713 404 765 456
rect 765 404 767 456
rect 711 402 767 404
rect 927 457 983 459
rect 927 405 929 457
rect 929 405 981 457
rect 981 405 983 457
rect 927 403 983 405
rect 1419 612 1475 614
rect 1190 600 1246 602
rect 1190 548 1192 600
rect 1192 548 1244 600
rect 1244 548 1246 600
rect 1419 560 1421 612
rect 1421 560 1473 612
rect 1473 560 1475 612
rect 1419 558 1475 560
rect 1638 602 1694 604
rect 1638 550 1640 602
rect 1640 550 1692 602
rect 1692 550 1694 602
rect 1190 546 1246 548
rect 1638 548 1694 550
rect 1830 606 1886 608
rect 1830 554 1832 606
rect 1832 554 1884 606
rect 1884 554 1886 606
rect 1830 552 1886 554
rect 2068 1290 2124 1292
rect 2068 1238 2070 1290
rect 2070 1238 2122 1290
rect 2122 1238 2124 1290
rect 2068 1236 2124 1238
rect 419 -76 475 -74
rect 419 -128 421 -76
rect 421 -128 473 -76
rect 473 -128 475 -76
rect 419 -130 475 -128
rect 618 -79 674 -77
rect 618 -131 620 -79
rect 620 -131 672 -79
rect 672 -131 674 -79
rect 618 -133 674 -131
rect 829 -79 885 -77
rect 829 -131 831 -79
rect 831 -131 883 -79
rect 883 -131 885 -79
rect 829 -133 885 -131
rect 1035 -79 1091 -77
rect 1035 -131 1037 -79
rect 1037 -131 1089 -79
rect 1089 -131 1091 -79
rect 1035 -133 1091 -131
rect 1263 -81 1319 -79
rect 1263 -133 1265 -81
rect 1265 -133 1317 -81
rect 1317 -133 1319 -81
rect 1263 -135 1319 -133
rect 1507 -81 1563 -79
rect 1507 -133 1509 -81
rect 1509 -133 1561 -81
rect 1561 -133 1563 -81
rect 1507 -135 1563 -133
rect 1737 -79 1793 -77
rect 1737 -131 1739 -79
rect 1739 -131 1791 -79
rect 1791 -131 1793 -79
rect 1737 -133 1793 -131
rect 1943 -79 1999 -77
rect 1943 -131 1945 -79
rect 1945 -131 1997 -79
rect 1997 -131 1999 -79
rect 1943 -133 1999 -131
rect 2427 2973 2483 2975
rect 2427 2921 2429 2973
rect 2429 2921 2481 2973
rect 2481 2921 2483 2973
rect 2427 2919 2483 2921
rect 2324 604 2380 606
rect 2324 552 2326 604
rect 2326 552 2378 604
rect 2378 552 2380 604
rect 2324 550 2380 552
rect 2650 2976 2706 2978
rect 2650 2924 2652 2976
rect 2652 2924 2704 2976
rect 2704 2924 2706 2976
rect 2650 2922 2706 2924
rect 2882 2975 2938 2977
rect 2882 2923 2884 2975
rect 2884 2923 2936 2975
rect 2936 2923 2938 2975
rect 2882 2921 2938 2923
rect 2701 1834 2757 1836
rect 2701 1782 2703 1834
rect 2703 1782 2755 1834
rect 2755 1782 2757 1834
rect 2701 1780 2757 1782
rect 3026 1836 3082 1838
rect 3026 1784 3028 1836
rect 3028 1784 3080 1836
rect 3080 1784 3082 1836
rect 3026 1782 3082 1784
rect 3294 1836 3350 1838
rect 3294 1784 3296 1836
rect 3296 1784 3348 1836
rect 3348 1784 3350 1836
rect 3294 1782 3350 1784
rect 2652 1146 2708 1148
rect 2652 1094 2654 1146
rect 2654 1094 2706 1146
rect 2706 1094 2708 1146
rect 2652 1092 2708 1094
rect 2867 1143 2923 1145
rect 2867 1091 2869 1143
rect 2869 1091 2921 1143
rect 2921 1091 2923 1143
rect 2867 1089 2923 1091
rect 3065 1140 3121 1142
rect 3065 1088 3067 1140
rect 3067 1088 3119 1140
rect 3119 1088 3121 1140
rect 3065 1086 3121 1088
rect 3260 1150 3316 1152
rect 3260 1098 3262 1150
rect 3262 1098 3314 1150
rect 3314 1098 3316 1150
rect 3260 1096 3316 1098
rect 3560 1836 3616 1838
rect 3560 1784 3562 1836
rect 3562 1784 3614 1836
rect 3614 1784 3616 1836
rect 3560 1782 3616 1784
rect 3800 1834 3856 1836
rect 3800 1782 3802 1834
rect 3802 1782 3854 1834
rect 3854 1782 3856 1834
rect 3800 1780 3856 1782
rect 4226 2437 4282 2439
rect 4226 2385 4228 2437
rect 4228 2385 4280 2437
rect 4280 2385 4282 2437
rect 4226 2383 4282 2385
rect 4518 2972 4574 2974
rect 4518 2920 4520 2972
rect 4520 2920 4572 2972
rect 4572 2920 4574 2972
rect 4518 2918 4574 2920
rect 4475 2440 4531 2442
rect 4475 2388 4477 2440
rect 4477 2388 4529 2440
rect 4529 2388 4531 2440
rect 4475 2386 4531 2388
rect 4192 1290 4248 1292
rect 4192 1238 4194 1290
rect 4194 1238 4246 1290
rect 4246 1238 4248 1290
rect 4192 1236 4248 1238
rect 3540 1148 3596 1150
rect 3540 1096 3542 1148
rect 3542 1096 3594 1148
rect 3594 1096 3596 1148
rect 3540 1094 3596 1096
rect 3759 1146 3815 1148
rect 3759 1094 3761 1146
rect 3761 1094 3813 1146
rect 3813 1094 3815 1146
rect 3759 1092 3815 1094
rect 2648 453 2704 455
rect 2648 401 2650 453
rect 2650 401 2702 453
rect 2702 401 2704 453
rect 2648 399 2704 401
rect 2838 453 2894 455
rect 2838 401 2840 453
rect 2840 401 2892 453
rect 2892 401 2894 453
rect 2838 399 2894 401
rect 3048 456 3104 458
rect 3048 404 3050 456
rect 3050 404 3102 456
rect 3102 404 3104 456
rect 3048 402 3104 404
rect 3265 453 3321 455
rect 3265 401 3267 453
rect 3267 401 3319 453
rect 3319 401 3321 453
rect 3265 399 3321 401
rect 4116 603 4172 605
rect 4116 551 4118 603
rect 4118 551 4170 603
rect 4170 551 4172 603
rect 4116 549 4172 551
rect 3560 456 3616 458
rect 3560 404 3562 456
rect 3562 404 3614 456
rect 3614 404 3616 456
rect 3560 402 3616 404
rect 3784 461 3840 463
rect 3784 409 3786 461
rect 3786 409 3838 461
rect 3838 409 3840 461
rect 3784 407 3840 409
rect 2161 -74 2217 -72
rect 2161 -126 2163 -74
rect 2163 -126 2215 -74
rect 2215 -126 2217 -74
rect 2161 -128 2217 -126
rect 2364 -80 2420 -78
rect 2364 -132 2366 -80
rect 2366 -132 2418 -80
rect 2418 -132 2420 -80
rect 2364 -134 2420 -132
rect 2572 -77 2628 -75
rect 2572 -129 2574 -77
rect 2574 -129 2626 -77
rect 2626 -129 2628 -77
rect 2572 -131 2628 -129
rect 4470 1289 4526 1291
rect 4470 1237 4472 1289
rect 4472 1237 4524 1289
rect 4524 1237 4526 1289
rect 4470 1235 4526 1237
rect 2835 -81 2891 -79
rect 2835 -133 2837 -81
rect 2837 -133 2889 -81
rect 2889 -133 2891 -81
rect 2835 -135 2891 -133
rect 3043 -80 3099 -78
rect 3043 -132 3045 -80
rect 3045 -132 3097 -80
rect 3097 -132 3099 -80
rect 3043 -134 3099 -132
rect 3253 -83 3309 -81
rect 3253 -135 3255 -83
rect 3255 -135 3307 -83
rect 3307 -135 3309 -83
rect 3253 -137 3309 -135
rect 3453 -77 3509 -75
rect 3453 -129 3455 -77
rect 3455 -129 3507 -77
rect 3507 -129 3509 -77
rect 3453 -131 3509 -129
rect 3656 -80 3712 -78
rect 3656 -132 3658 -80
rect 3658 -132 3710 -80
rect 3710 -132 3712 -80
rect 3656 -134 3712 -132
rect 3866 -80 3922 -78
rect 3866 -132 3868 -80
rect 3868 -132 3920 -80
rect 3920 -132 3922 -80
rect 3866 -134 3922 -132
rect 4067 -79 4123 -77
rect 4067 -131 4069 -79
rect 4069 -131 4121 -79
rect 4121 -131 4123 -79
rect 4067 -133 4123 -131
rect 4283 -78 4339 -76
rect 4283 -130 4285 -78
rect 4285 -130 4337 -78
rect 4337 -130 4339 -78
rect 4283 -132 4339 -130
rect 4509 601 4565 603
rect 4509 549 4511 601
rect 4511 549 4563 601
rect 4563 549 4565 601
rect 4509 547 4565 549
rect 4826 2973 4882 2975
rect 4826 2921 4828 2973
rect 4828 2921 4880 2973
rect 4880 2921 4882 2973
rect 4826 2919 4882 2921
rect 4819 2426 4875 2428
rect 4819 2374 4821 2426
rect 4821 2374 4873 2426
rect 4873 2374 4875 2426
rect 4819 2372 4875 2374
rect 4706 609 4762 611
rect 4706 557 4708 609
rect 4708 557 4760 609
rect 4760 557 4762 609
rect 4706 555 4762 557
rect 5026 2974 5082 2976
rect 5026 2922 5028 2974
rect 5028 2922 5080 2974
rect 5080 2922 5082 2974
rect 5026 2920 5082 2922
rect 5245 2973 5301 2975
rect 5245 2921 5247 2973
rect 5247 2921 5299 2973
rect 5299 2921 5301 2973
rect 5245 2919 5301 2921
rect 5491 2972 5547 2974
rect 5491 2920 5493 2972
rect 5493 2920 5545 2972
rect 5545 2920 5547 2972
rect 5491 2918 5547 2920
rect 5699 2974 5755 2976
rect 5699 2922 5701 2974
rect 5701 2922 5753 2974
rect 5753 2922 5755 2974
rect 5699 2920 5755 2922
rect 5901 2975 5957 2977
rect 5901 2923 5903 2975
rect 5903 2923 5955 2975
rect 5955 2923 5957 2975
rect 5901 2921 5957 2923
rect 6094 2974 6150 2976
rect 6094 2922 6096 2974
rect 6096 2922 6148 2974
rect 6148 2922 6150 2974
rect 6094 2920 6150 2922
rect 5073 2432 5129 2434
rect 5073 2380 5075 2432
rect 5075 2380 5127 2432
rect 5127 2380 5129 2432
rect 5073 2378 5129 2380
rect 5302 2432 5358 2434
rect 5302 2380 5304 2432
rect 5304 2380 5356 2432
rect 5356 2380 5358 2432
rect 5302 2378 5358 2380
rect 5594 1837 5650 1839
rect 5594 1785 5596 1837
rect 5596 1785 5648 1837
rect 5648 1785 5650 1837
rect 5594 1783 5650 1785
rect 5042 1294 5098 1296
rect 5042 1242 5044 1294
rect 5044 1242 5096 1294
rect 5096 1242 5098 1294
rect 5042 1240 5098 1242
rect 5281 1294 5337 1296
rect 5281 1242 5283 1294
rect 5283 1242 5335 1294
rect 5335 1242 5337 1294
rect 5281 1240 5337 1242
rect 5580 1143 5636 1145
rect 5580 1091 5582 1143
rect 5582 1091 5634 1143
rect 5634 1091 5636 1143
rect 5580 1089 5636 1091
rect 5960 1840 6016 1842
rect 5960 1788 5962 1840
rect 5962 1788 6014 1840
rect 6014 1788 6016 1840
rect 5960 1786 6016 1788
rect 6204 1840 6260 1842
rect 6204 1788 6206 1840
rect 6206 1788 6258 1840
rect 6258 1788 6260 1840
rect 6204 1786 6260 1788
rect 6466 2973 6522 2975
rect 6466 2921 6468 2973
rect 6468 2921 6520 2973
rect 6520 2921 6522 2973
rect 6466 2919 6522 2921
rect 6655 2971 6711 2973
rect 6655 2919 6657 2971
rect 6657 2919 6709 2971
rect 6709 2919 6711 2971
rect 6655 2917 6711 2919
rect 6627 1831 6683 1833
rect 6627 1779 6629 1831
rect 6629 1779 6681 1831
rect 6681 1779 6683 1831
rect 6627 1777 6683 1779
rect 6945 2971 7001 2973
rect 6945 2919 6947 2971
rect 6947 2919 6999 2971
rect 6999 2919 7001 2971
rect 6945 2917 7001 2919
rect 7020 2437 7076 2439
rect 7020 2385 7022 2437
rect 7022 2385 7074 2437
rect 7074 2385 7076 2437
rect 7020 2383 7076 2385
rect 5931 1140 5987 1142
rect 5931 1088 5933 1140
rect 5933 1088 5985 1140
rect 5985 1088 5987 1140
rect 5931 1086 5987 1088
rect 6120 1138 6176 1140
rect 6120 1086 6122 1138
rect 6122 1086 6174 1138
rect 6174 1086 6176 1138
rect 6120 1084 6176 1086
rect 6325 1145 6381 1147
rect 6325 1093 6327 1145
rect 6327 1093 6379 1145
rect 6379 1093 6381 1145
rect 6325 1091 6381 1093
rect 6516 1147 6572 1149
rect 6516 1095 6518 1147
rect 6518 1095 6570 1147
rect 6570 1095 6572 1147
rect 6516 1093 6572 1095
rect 5036 611 5092 613
rect 5036 559 5038 611
rect 5038 559 5090 611
rect 5090 559 5092 611
rect 5036 557 5092 559
rect 5232 611 5288 613
rect 5232 559 5234 611
rect 5234 559 5286 611
rect 5286 559 5288 611
rect 5232 557 5288 559
rect 5662 454 5718 456
rect 5662 402 5664 454
rect 5664 402 5716 454
rect 5716 402 5718 454
rect 5662 400 5718 402
rect 5962 452 6018 454
rect 5962 400 5964 452
rect 5964 400 6016 452
rect 6016 400 6018 452
rect 5962 398 6018 400
rect 6214 456 6270 458
rect 6214 404 6216 456
rect 6216 404 6268 456
rect 6268 404 6270 456
rect 6214 402 6270 404
rect 6431 461 6487 463
rect 6431 409 6433 461
rect 6433 409 6485 461
rect 6485 409 6487 461
rect 6431 407 6487 409
rect 6632 458 6688 460
rect 6632 406 6634 458
rect 6634 406 6686 458
rect 6686 406 6688 458
rect 6632 404 6688 406
rect 4564 -80 4620 -78
rect 4564 -132 4566 -80
rect 4566 -132 4618 -80
rect 4618 -132 4620 -80
rect 4564 -134 4620 -132
rect 4784 -85 4840 -83
rect 4784 -137 4786 -85
rect 4786 -137 4838 -85
rect 4838 -137 4840 -85
rect 4784 -139 4840 -137
rect 4989 -84 5045 -82
rect 4989 -136 4991 -84
rect 4991 -136 5043 -84
rect 5043 -136 5045 -84
rect 4989 -138 5045 -136
rect 5210 -78 5266 -76
rect 5210 -130 5212 -78
rect 5212 -130 5264 -78
rect 5264 -130 5266 -78
rect 5210 -132 5266 -130
rect 5415 -85 5471 -83
rect 5415 -137 5417 -85
rect 5417 -137 5469 -85
rect 5469 -137 5471 -85
rect 5415 -139 5471 -137
rect 5624 -84 5680 -82
rect 5624 -136 5626 -84
rect 5626 -136 5678 -84
rect 5678 -136 5680 -84
rect 5624 -138 5680 -136
rect 5841 -84 5897 -82
rect 5841 -136 5843 -84
rect 5843 -136 5895 -84
rect 5895 -136 5897 -84
rect 5841 -138 5897 -136
rect 6055 -79 6111 -77
rect 6055 -131 6057 -79
rect 6057 -131 6109 -79
rect 6109 -131 6111 -79
rect 6055 -133 6111 -131
rect 6250 -81 6306 -79
rect 6250 -133 6252 -81
rect 6252 -133 6304 -81
rect 6304 -133 6306 -81
rect 6250 -135 6306 -133
rect 6445 -84 6501 -82
rect 6445 -136 6447 -84
rect 6447 -136 6499 -84
rect 6499 -136 6501 -84
rect 6445 -138 6501 -136
rect 6647 -81 6703 -79
rect 6647 -133 6649 -81
rect 6649 -133 6701 -81
rect 6701 -133 6703 -81
rect 6647 -135 6703 -133
rect 7218 2973 7274 2975
rect 7218 2921 7220 2973
rect 7220 2921 7272 2973
rect 7272 2921 7274 2973
rect 7218 2919 7274 2921
rect 7224 2439 7280 2441
rect 7224 2387 7226 2439
rect 7226 2387 7278 2439
rect 7278 2387 7280 2439
rect 7224 2385 7280 2387
rect 7139 604 7195 606
rect 7139 552 7141 604
rect 7141 552 7193 604
rect 7193 552 7195 604
rect 7139 550 7195 552
rect 7547 2437 7603 2439
rect 7547 2385 7549 2437
rect 7549 2385 7601 2437
rect 7601 2385 7603 2437
rect 7547 2383 7603 2385
rect 7439 1292 7495 1294
rect 7439 1240 7441 1292
rect 7441 1240 7493 1292
rect 7493 1240 7495 1292
rect 7439 1238 7495 1240
rect 7666 1297 7722 1299
rect 7666 1245 7668 1297
rect 7668 1245 7720 1297
rect 7720 1245 7722 1297
rect 7666 1243 7722 1245
rect 7856 1299 7912 1301
rect 7856 1247 7858 1299
rect 7858 1247 7910 1299
rect 7910 1247 7912 1299
rect 7856 1245 7912 1247
rect 8072 1290 8128 1292
rect 8072 1238 8074 1290
rect 8074 1238 8126 1290
rect 8126 1238 8128 1290
rect 8072 1236 8128 1238
rect 8570 1833 8626 1835
rect 8570 1781 8572 1833
rect 8572 1781 8624 1833
rect 8624 1781 8626 1833
rect 8570 1779 8626 1781
rect 8822 1830 8878 1832
rect 8822 1778 8824 1830
rect 8824 1778 8876 1830
rect 8876 1778 8878 1830
rect 8822 1776 8878 1778
rect 9028 1838 9084 1840
rect 9028 1786 9030 1838
rect 9030 1786 9082 1838
rect 9082 1786 9084 1838
rect 9028 1784 9084 1786
rect 9311 1832 9367 1834
rect 9311 1780 9313 1832
rect 9313 1780 9365 1832
rect 9365 1780 9367 1832
rect 9311 1778 9367 1780
rect 8561 1149 8617 1151
rect 8561 1097 8563 1149
rect 8563 1097 8615 1149
rect 8615 1097 8617 1149
rect 8561 1095 8617 1097
rect 8751 1151 8807 1153
rect 8751 1099 8753 1151
rect 8753 1099 8805 1151
rect 8805 1099 8807 1151
rect 8751 1097 8807 1099
rect 8945 1149 9001 1151
rect 8945 1097 8947 1149
rect 8947 1097 8999 1149
rect 8999 1097 9001 1149
rect 8945 1095 9001 1097
rect 7440 608 7496 610
rect 7440 556 7442 608
rect 7442 556 7494 608
rect 7494 556 7496 608
rect 7440 554 7496 556
rect 7646 609 7702 611
rect 7646 557 7648 609
rect 7648 557 7700 609
rect 7700 557 7702 609
rect 7646 555 7702 557
rect 7856 605 7912 607
rect 7856 553 7858 605
rect 7858 553 7910 605
rect 7910 553 7912 605
rect 7856 551 7912 553
rect 8067 611 8123 613
rect 8067 559 8069 611
rect 8069 559 8121 611
rect 8121 559 8123 611
rect 8067 557 8123 559
rect 8517 449 8573 451
rect 8517 397 8519 449
rect 8519 397 8571 449
rect 8571 397 8573 449
rect 8517 395 8573 397
rect 8709 449 8765 451
rect 8709 397 8711 449
rect 8711 397 8763 449
rect 8763 397 8765 449
rect 8709 395 8765 397
rect 8909 449 8965 451
rect 8909 397 8911 449
rect 8911 397 8963 449
rect 8963 397 8965 449
rect 8909 395 8965 397
rect 6931 -80 6987 -78
rect 6931 -132 6933 -80
rect 6933 -132 6985 -80
rect 6985 -132 6987 -80
rect 6931 -134 6987 -132
rect 7130 -79 7186 -77
rect 7130 -131 7132 -79
rect 7132 -131 7184 -79
rect 7184 -131 7186 -79
rect 7130 -133 7186 -131
rect 7333 -77 7389 -75
rect 7333 -129 7335 -77
rect 7335 -129 7387 -77
rect 7387 -129 7389 -77
rect 7333 -131 7389 -129
rect 9256 1145 9312 1147
rect 9256 1093 9258 1145
rect 9258 1093 9310 1145
rect 9310 1093 9312 1145
rect 9256 1091 9312 1093
rect 7598 -80 7654 -78
rect 7598 -132 7600 -80
rect 7600 -132 7652 -80
rect 7652 -132 7654 -80
rect 7598 -134 7654 -132
rect 7796 -81 7852 -79
rect 7796 -133 7798 -81
rect 7798 -133 7850 -81
rect 7850 -133 7852 -81
rect 7796 -135 7852 -133
rect 7985 -79 8041 -77
rect 7985 -131 7987 -79
rect 7987 -131 8039 -79
rect 8039 -131 8041 -79
rect 7985 -133 8041 -131
rect 8197 -79 8253 -77
rect 8197 -131 8199 -79
rect 8199 -131 8251 -79
rect 8251 -131 8253 -79
rect 8197 -133 8253 -131
rect 8414 -79 8470 -77
rect 8414 -131 8416 -79
rect 8416 -131 8468 -79
rect 8468 -131 8470 -79
rect 8414 -133 8470 -131
rect 8619 -83 8675 -81
rect 8619 -135 8621 -83
rect 8621 -135 8673 -83
rect 8673 -135 8675 -83
rect 8619 -137 8675 -135
rect 8824 -83 8880 -81
rect 8824 -135 8826 -83
rect 8826 -135 8878 -83
rect 8878 -135 8880 -83
rect 8824 -137 8880 -135
rect 9032 -78 9088 -76
rect 9032 -130 9034 -78
rect 9034 -130 9086 -78
rect 9086 -130 9088 -78
rect 9032 -132 9088 -130
rect 9609 1833 9665 1835
rect 9609 1781 9611 1833
rect 9611 1781 9663 1833
rect 9663 1781 9665 1833
rect 9609 1779 9665 1781
rect 9527 457 9583 459
rect 9527 405 9529 457
rect 9529 405 9581 457
rect 9581 405 9583 457
rect 9527 403 9583 405
rect 10053 1293 10109 1295
rect 10053 1241 10055 1293
rect 10055 1241 10107 1293
rect 10107 1241 10109 1293
rect 10053 1239 10109 1241
rect 10282 1296 10338 1298
rect 10282 1244 10284 1296
rect 10284 1244 10336 1296
rect 10336 1244 10338 1296
rect 10282 1242 10338 1244
rect 10508 1301 10564 1303
rect 10508 1249 10510 1301
rect 10510 1249 10562 1301
rect 10562 1249 10564 1301
rect 10508 1247 10564 1249
rect 11441 1834 11497 1836
rect 11441 1782 11443 1834
rect 11443 1782 11495 1834
rect 11495 1782 11497 1834
rect 11441 1780 11497 1782
rect 11651 1836 11707 1838
rect 11651 1784 11653 1836
rect 11653 1784 11705 1836
rect 11705 1784 11707 1836
rect 11651 1782 11707 1784
rect 10736 1293 10792 1295
rect 10736 1241 10738 1293
rect 10738 1241 10790 1293
rect 10790 1241 10792 1293
rect 10736 1239 10792 1241
rect 10972 1299 11028 1301
rect 10972 1247 10974 1299
rect 10974 1247 11026 1299
rect 11026 1247 11028 1299
rect 10972 1245 11028 1247
rect 11164 1290 11220 1292
rect 11164 1238 11166 1290
rect 11166 1238 11218 1290
rect 11218 1238 11220 1290
rect 11164 1236 11220 1238
rect 11439 1144 11495 1146
rect 11439 1092 11441 1144
rect 11441 1092 11493 1144
rect 11493 1092 11495 1144
rect 11439 1090 11495 1092
rect 9947 600 10003 602
rect 9947 548 9949 600
rect 9949 548 10001 600
rect 10001 548 10003 600
rect 9947 546 10003 548
rect 10204 607 10260 609
rect 10204 555 10206 607
rect 10206 555 10258 607
rect 10258 555 10260 607
rect 10204 553 10260 555
rect 10454 603 10510 605
rect 10454 551 10456 603
rect 10456 551 10508 603
rect 10508 551 10510 603
rect 10454 549 10510 551
rect 10725 608 10781 610
rect 10725 556 10727 608
rect 10727 556 10779 608
rect 10779 556 10781 608
rect 10725 554 10781 556
rect 10966 611 11022 613
rect 10966 559 10968 611
rect 10968 559 11020 611
rect 11020 559 11022 611
rect 10966 557 11022 559
rect 11191 607 11247 609
rect 11191 555 11193 607
rect 11193 555 11245 607
rect 11245 555 11247 607
rect 11191 553 11247 555
rect 11428 453 11484 455
rect 11428 401 11430 453
rect 11430 401 11482 453
rect 11482 401 11484 453
rect 11428 399 11484 401
rect 9315 -79 9371 -77
rect 9315 -131 9317 -79
rect 9317 -131 9369 -79
rect 9369 -131 9371 -79
rect 9315 -133 9371 -131
rect 9508 -81 9564 -79
rect 9508 -133 9510 -81
rect 9510 -133 9562 -81
rect 9562 -133 9564 -81
rect 9508 -135 9564 -133
rect 9734 -83 9790 -81
rect 9734 -135 9736 -83
rect 9736 -135 9788 -83
rect 9788 -135 9790 -83
rect 9734 -137 9790 -135
rect 11643 1144 11699 1146
rect 11643 1092 11645 1144
rect 11645 1092 11697 1144
rect 11697 1092 11699 1144
rect 11643 1090 11699 1092
rect 9999 -83 10055 -81
rect 9999 -135 10001 -83
rect 10001 -135 10053 -83
rect 10053 -135 10055 -83
rect 9999 -137 10055 -135
rect 10193 -79 10249 -77
rect 10193 -131 10195 -79
rect 10195 -131 10247 -79
rect 10247 -131 10249 -79
rect 10193 -133 10249 -131
rect 10391 -88 10447 -86
rect 10391 -140 10393 -88
rect 10393 -140 10445 -88
rect 10445 -140 10447 -88
rect 10391 -142 10447 -140
rect 10595 -80 10651 -78
rect 10595 -132 10597 -80
rect 10597 -132 10649 -80
rect 10649 -132 10651 -80
rect 10595 -134 10651 -132
rect 10815 -77 10871 -75
rect 10815 -129 10817 -77
rect 10817 -129 10869 -77
rect 10869 -129 10871 -77
rect 10815 -131 10871 -129
rect 11030 -81 11086 -79
rect 11030 -133 11032 -81
rect 11032 -133 11084 -81
rect 11084 -133 11086 -81
rect 11030 -135 11086 -133
rect 11258 -78 11314 -76
rect 11258 -130 11260 -78
rect 11260 -130 11312 -78
rect 11312 -130 11314 -78
rect 11258 -132 11314 -130
rect 11462 -81 11518 -79
rect 11462 -133 11464 -81
rect 11464 -133 11516 -81
rect 11516 -133 11518 -81
rect 11462 -135 11518 -133
rect 11684 453 11740 455
rect 11684 401 11686 453
rect 11686 401 11738 453
rect 11738 401 11740 453
rect 11684 399 11740 401
rect 12002 1834 12058 1836
rect 12002 1782 12004 1834
rect 12004 1782 12056 1834
rect 12056 1782 12058 1834
rect 12002 1780 12058 1782
rect 11919 453 11975 455
rect 11919 401 11921 453
rect 11921 401 11973 453
rect 11973 401 11975 453
rect 11919 399 11975 401
rect 12282 1834 12338 1836
rect 12282 1782 12284 1834
rect 12284 1782 12336 1834
rect 12336 1782 12338 1834
rect 12282 1780 12338 1782
rect 12599 1833 12655 1835
rect 12599 1781 12601 1833
rect 12601 1781 12653 1833
rect 12653 1781 12655 1833
rect 12599 1779 12655 1781
rect 12208 1140 12264 1142
rect 12208 1088 12210 1140
rect 12210 1088 12262 1140
rect 12262 1088 12264 1140
rect 12208 1086 12264 1088
rect 12899 1290 12955 1292
rect 12899 1238 12901 1290
rect 12901 1238 12953 1290
rect 12953 1238 12955 1290
rect 12899 1236 12955 1238
rect 12447 1142 12503 1144
rect 12447 1090 12449 1142
rect 12449 1090 12501 1142
rect 12501 1090 12503 1142
rect 12447 1088 12503 1090
rect 12651 1142 12707 1144
rect 12651 1090 12653 1142
rect 12653 1090 12705 1142
rect 12705 1090 12707 1142
rect 12651 1088 12707 1090
rect 13103 1295 13159 1297
rect 13103 1243 13105 1295
rect 13105 1243 13157 1295
rect 13157 1243 13159 1295
rect 13103 1241 13159 1243
rect 13294 1290 13350 1292
rect 13294 1238 13296 1290
rect 13296 1238 13348 1290
rect 13348 1238 13350 1290
rect 13294 1236 13350 1238
rect 13496 1289 13552 1291
rect 13496 1237 13498 1289
rect 13498 1237 13550 1289
rect 13550 1237 13552 1289
rect 13496 1235 13552 1237
rect 13786 1290 13842 1292
rect 13786 1238 13788 1290
rect 13788 1238 13840 1290
rect 13840 1238 13842 1290
rect 13786 1236 13842 1238
rect 12898 605 12954 607
rect 12898 553 12900 605
rect 12900 553 12952 605
rect 12952 553 12954 605
rect 12898 551 12954 553
rect 12208 455 12264 457
rect 12208 403 12210 455
rect 12210 403 12262 455
rect 12262 403 12264 455
rect 12208 401 12264 403
rect 12398 453 12454 455
rect 12398 401 12400 453
rect 12400 401 12452 453
rect 12452 401 12454 453
rect 12398 399 12454 401
rect 12602 455 12658 457
rect 12602 403 12604 455
rect 12604 403 12656 455
rect 12656 403 12658 455
rect 12602 401 12658 403
rect 13099 606 13155 608
rect 13099 554 13101 606
rect 13101 554 13153 606
rect 13153 554 13155 606
rect 13099 552 13155 554
rect 13317 602 13373 604
rect 13317 550 13319 602
rect 13319 550 13371 602
rect 13371 550 13373 602
rect 13317 548 13373 550
rect 13524 606 13580 608
rect 13524 554 13526 606
rect 13526 554 13578 606
rect 13578 554 13580 606
rect 13524 552 13580 554
rect 13729 605 13785 607
rect 13729 553 13731 605
rect 13731 553 13783 605
rect 13783 553 13785 605
rect 13729 551 13785 553
rect 11700 -79 11756 -77
rect 11700 -131 11702 -79
rect 11702 -131 11754 -79
rect 11754 -131 11756 -79
rect 11700 -133 11756 -131
rect 11893 -78 11949 -76
rect 11893 -130 11895 -78
rect 11895 -130 11947 -78
rect 11947 -130 11949 -78
rect 11893 -132 11949 -130
rect 12090 -83 12146 -81
rect 12090 -135 12092 -83
rect 12092 -135 12144 -83
rect 12144 -135 12146 -83
rect 12090 -137 12146 -135
rect 14071 1289 14127 1291
rect 14071 1237 14073 1289
rect 14073 1237 14125 1289
rect 14125 1237 14127 1289
rect 14071 1235 14127 1237
rect 12346 -80 12402 -78
rect 12346 -132 12348 -80
rect 12348 -132 12400 -80
rect 12400 -132 12402 -80
rect 12346 -134 12402 -132
rect 12585 -84 12641 -82
rect 12585 -136 12587 -84
rect 12587 -136 12639 -84
rect 12639 -136 12641 -84
rect 12585 -138 12641 -136
rect 12818 -88 12874 -86
rect 12818 -140 12820 -88
rect 12820 -140 12872 -88
rect 12872 -140 12874 -88
rect 12818 -142 12874 -140
rect 13039 -83 13095 -81
rect 13039 -135 13041 -83
rect 13041 -135 13093 -83
rect 13093 -135 13095 -83
rect 13039 -137 13095 -135
rect 13230 -83 13286 -81
rect 13230 -135 13232 -83
rect 13232 -135 13284 -83
rect 13284 -135 13286 -83
rect 13230 -137 13286 -135
rect 13458 -81 13514 -79
rect 13458 -133 13460 -81
rect 13460 -133 13512 -81
rect 13512 -133 13514 -81
rect 13458 -135 13514 -133
rect 13655 -86 13711 -84
rect 13655 -138 13657 -86
rect 13657 -138 13709 -86
rect 13709 -138 13711 -86
rect 13655 -140 13711 -138
rect 13867 -86 13923 -84
rect 13867 -138 13869 -86
rect 13869 -138 13921 -86
rect 13921 -138 13923 -86
rect 13867 -140 13923 -138
rect 14076 601 14132 603
rect 14076 549 14078 601
rect 14078 549 14130 601
rect 14130 549 14132 601
rect 14076 547 14132 549
rect 14389 1831 14445 1833
rect 14389 1779 14391 1831
rect 14391 1779 14443 1831
rect 14443 1779 14445 1831
rect 14389 1777 14445 1779
rect 14388 461 14444 463
rect 14388 409 14390 461
rect 14390 409 14442 461
rect 14442 409 14444 461
rect 14388 407 14444 409
rect 14684 1831 14740 1833
rect 14684 1779 14686 1831
rect 14686 1779 14738 1831
rect 14738 1779 14740 1831
rect 14684 1777 14740 1779
rect 14971 1831 15027 1833
rect 14971 1779 14973 1831
rect 14973 1779 15025 1831
rect 15025 1779 15027 1831
rect 14971 1777 15027 1779
rect 15261 1831 15317 1833
rect 15261 1779 15263 1831
rect 15263 1779 15315 1831
rect 15315 1779 15317 1831
rect 15261 1777 15317 1779
rect 14611 1150 14667 1152
rect 14611 1098 14613 1150
rect 14613 1098 14665 1150
rect 14665 1098 14667 1150
rect 14611 1096 14667 1098
rect 14844 1148 14900 1150
rect 14844 1096 14846 1148
rect 14846 1096 14898 1148
rect 14898 1096 14900 1148
rect 14844 1094 14900 1096
rect 15051 1146 15107 1148
rect 15051 1094 15053 1146
rect 15053 1094 15105 1146
rect 15105 1094 15107 1146
rect 15051 1092 15107 1094
rect 15260 1148 15316 1150
rect 15260 1096 15262 1148
rect 15262 1096 15314 1148
rect 15314 1096 15316 1148
rect 15260 1094 15316 1096
rect 15545 1834 15601 1836
rect 15545 1782 15547 1834
rect 15547 1782 15599 1834
rect 15599 1782 15601 1834
rect 15545 1780 15601 1782
rect 15826 1294 15882 1296
rect 15826 1242 15828 1294
rect 15828 1242 15880 1294
rect 15880 1242 15882 1294
rect 15826 1240 15882 1242
rect 16020 1298 16076 1300
rect 16020 1246 16022 1298
rect 16022 1246 16074 1298
rect 16074 1246 16076 1298
rect 16020 1244 16076 1246
rect 16209 1295 16265 1297
rect 16209 1243 16211 1295
rect 16211 1243 16263 1295
rect 16263 1243 16265 1295
rect 16209 1241 16265 1243
rect 15540 1150 15596 1152
rect 15540 1098 15542 1150
rect 15542 1098 15594 1150
rect 15594 1098 15596 1150
rect 15540 1096 15596 1098
rect 14630 457 14686 459
rect 14630 405 14632 457
rect 14632 405 14684 457
rect 14684 405 14686 457
rect 14630 403 14686 405
rect 14830 456 14886 458
rect 14830 404 14832 456
rect 14832 404 14884 456
rect 14884 404 14886 456
rect 14830 402 14886 404
rect 15020 464 15076 466
rect 15020 412 15022 464
rect 15022 412 15074 464
rect 15074 412 15076 464
rect 15020 410 15076 412
rect 15241 462 15297 464
rect 15241 410 15243 462
rect 15243 410 15295 462
rect 15295 410 15297 462
rect 15241 408 15297 410
rect 15828 605 15884 607
rect 15828 553 15830 605
rect 15830 553 15882 605
rect 15882 553 15884 605
rect 15828 551 15884 553
rect 16019 608 16075 610
rect 16019 556 16021 608
rect 16021 556 16073 608
rect 16073 556 16075 608
rect 16019 554 16075 556
rect 16214 610 16270 612
rect 16214 558 16216 610
rect 16216 558 16268 610
rect 16268 558 16270 610
rect 16214 556 16270 558
rect 15537 457 15593 459
rect 15537 405 15539 457
rect 15539 405 15591 457
rect 15591 405 15593 457
rect 15537 403 15593 405
rect 14094 -83 14150 -81
rect 14094 -135 14096 -83
rect 14096 -135 14148 -83
rect 14148 -135 14150 -83
rect 14094 -137 14150 -135
rect 14283 -82 14339 -80
rect 14283 -134 14285 -82
rect 14285 -134 14337 -82
rect 14337 -134 14339 -82
rect 14283 -136 14339 -134
rect 14509 -81 14565 -79
rect 14509 -133 14511 -81
rect 14511 -133 14563 -81
rect 14563 -133 14565 -81
rect 14509 -135 14565 -133
rect 16432 1297 16488 1299
rect 16432 1245 16434 1297
rect 16434 1245 16486 1297
rect 16486 1245 16488 1297
rect 16432 1243 16488 1245
rect 14763 -81 14819 -79
rect 14763 -133 14765 -81
rect 14765 -133 14817 -81
rect 14817 -133 14819 -81
rect 14763 -135 14819 -133
rect 15007 -84 15063 -82
rect 15007 -136 15009 -84
rect 15009 -136 15061 -84
rect 15061 -136 15063 -84
rect 15007 -138 15063 -136
rect 15237 -85 15293 -83
rect 15237 -137 15239 -85
rect 15239 -137 15291 -85
rect 15291 -137 15293 -85
rect 15237 -139 15293 -137
rect 15495 -82 15551 -80
rect 15495 -134 15497 -82
rect 15497 -134 15549 -82
rect 15549 -134 15551 -82
rect 15495 -136 15551 -134
rect 15705 -82 15761 -80
rect 15705 -134 15707 -82
rect 15707 -134 15759 -82
rect 15759 -134 15761 -82
rect 15705 -136 15761 -134
rect 15930 -82 15986 -80
rect 15930 -134 15932 -82
rect 15932 -134 15984 -82
rect 15984 -134 15986 -82
rect 15930 -136 15986 -134
rect 16149 -85 16205 -83
rect 16149 -137 16151 -85
rect 16151 -137 16203 -85
rect 16203 -137 16205 -85
rect 16149 -139 16205 -137
rect 16661 605 16717 607
rect 16661 553 16663 605
rect 16663 553 16715 605
rect 16715 553 16717 605
rect 16661 551 16717 553
rect 16495 -81 16551 -79
rect 16495 -133 16497 -81
rect 16497 -133 16549 -81
rect 16549 -133 16551 -81
rect 16495 -135 16551 -133
rect 16694 -84 16750 -82
rect 16694 -136 16696 -84
rect 16696 -136 16748 -84
rect 16748 -136 16750 -84
rect 16694 -138 16750 -136
<< metal3 >>
rect 16 2982 145 2993
rect 16 2918 47 2982
rect 111 2918 145 2982
rect 16 2907 145 2918
rect 218 2984 347 2995
rect 218 2920 249 2984
rect 313 2920 347 2984
rect 218 2909 347 2920
rect 429 2982 558 2993
rect 429 2918 460 2982
rect 524 2918 558 2982
rect 429 2907 558 2918
rect 619 2982 748 2993
rect 619 2918 650 2982
rect 714 2918 748 2982
rect 619 2907 748 2918
rect 827 2984 956 2995
rect 827 2920 858 2984
rect 922 2920 956 2984
rect 827 2909 956 2920
rect 1029 2984 1158 2995
rect 1029 2920 1060 2984
rect 1124 2920 1158 2984
rect 1029 2909 1158 2920
rect 1228 2986 1357 2997
rect 1228 2922 1259 2986
rect 1323 2922 1357 2986
rect 1228 2911 1357 2922
rect 1423 2983 1552 2994
rect 1423 2919 1454 2983
rect 1518 2919 1552 2983
rect 1423 2908 1552 2919
rect 1624 2985 1753 2996
rect 1624 2921 1655 2985
rect 1719 2921 1753 2985
rect 1624 2910 1753 2921
rect 1841 2983 1970 2994
rect 1841 2919 1872 2983
rect 1936 2919 1970 2983
rect 1841 2908 1970 2919
rect 2115 2986 2244 2997
rect 2115 2922 2146 2986
rect 2210 2922 2244 2986
rect 2115 2911 2244 2922
rect 2392 2979 2521 2990
rect 2392 2915 2423 2979
rect 2487 2915 2521 2979
rect 2392 2904 2521 2915
rect 2615 2982 2744 2993
rect 2615 2918 2646 2982
rect 2710 2918 2744 2982
rect 2615 2907 2744 2918
rect 2847 2981 2976 2992
rect 2847 2917 2878 2981
rect 2942 2917 2976 2981
rect 2847 2906 2976 2917
rect 4483 2978 4612 2989
rect 4483 2914 4514 2978
rect 4578 2914 4612 2978
rect 4483 2903 4612 2914
rect 4791 2979 4920 2990
rect 4791 2915 4822 2979
rect 4886 2915 4920 2979
rect 4791 2904 4920 2915
rect 4991 2980 5120 2991
rect 4991 2916 5022 2980
rect 5086 2916 5120 2980
rect 4991 2905 5120 2916
rect 5210 2979 5339 2990
rect 5210 2915 5241 2979
rect 5305 2915 5339 2979
rect 5210 2904 5339 2915
rect 5456 2978 5585 2989
rect 5456 2914 5487 2978
rect 5551 2914 5585 2978
rect 5456 2903 5585 2914
rect 5664 2980 5793 2991
rect 5664 2916 5695 2980
rect 5759 2916 5793 2980
rect 5664 2905 5793 2916
rect 5866 2981 5995 2992
rect 5866 2917 5897 2981
rect 5961 2917 5995 2981
rect 5866 2906 5995 2917
rect 6059 2980 6188 2991
rect 6059 2916 6090 2980
rect 6154 2916 6188 2980
rect 6059 2905 6188 2916
rect 6431 2979 6560 2990
rect 6431 2915 6462 2979
rect 6526 2915 6560 2979
rect 6431 2904 6560 2915
rect 6620 2977 6749 2988
rect 6620 2913 6651 2977
rect 6715 2913 6749 2977
rect 6620 2902 6749 2913
rect 6910 2977 7039 2988
rect 6910 2913 6941 2977
rect 7005 2913 7039 2977
rect 6910 2902 7039 2913
rect 7183 2979 7312 2990
rect 7183 2915 7214 2979
rect 7278 2915 7312 2979
rect 7183 2904 7312 2915
rect 1134 2443 1263 2454
rect 1134 2379 1165 2443
rect 1229 2379 1263 2443
rect 1134 2368 1263 2379
rect 1353 2447 1482 2458
rect 1353 2383 1384 2447
rect 1448 2383 1482 2447
rect 1353 2372 1482 2383
rect 1636 2447 1765 2458
rect 1636 2383 1667 2447
rect 1731 2383 1765 2447
rect 1636 2372 1765 2383
rect 1845 2447 1974 2458
rect 1845 2383 1876 2447
rect 1940 2383 1974 2447
rect 1845 2372 1974 2383
rect 2116 2445 2245 2456
rect 2116 2381 2147 2445
rect 2211 2381 2245 2445
rect 2116 2370 2245 2381
rect 4191 2443 4320 2454
rect 4191 2379 4222 2443
rect 4286 2379 4320 2443
rect 4191 2368 4320 2379
rect 4440 2446 4569 2457
rect 4440 2382 4471 2446
rect 4535 2382 4569 2446
rect 4440 2371 4569 2382
rect 4784 2432 4913 2443
rect 4784 2368 4815 2432
rect 4879 2368 4913 2432
rect 4784 2357 4913 2368
rect 5038 2438 5167 2449
rect 5038 2374 5069 2438
rect 5133 2374 5167 2438
rect 5038 2363 5167 2374
rect 5267 2438 5396 2449
rect 5267 2374 5298 2438
rect 5362 2374 5396 2438
rect 5267 2363 5396 2374
rect 6985 2443 7114 2454
rect 6985 2379 7016 2443
rect 7080 2379 7114 2443
rect 6985 2368 7114 2379
rect 7189 2445 7318 2456
rect 7189 2381 7220 2445
rect 7284 2381 7318 2445
rect 7189 2370 7318 2381
rect 7512 2443 7641 2454
rect 7512 2379 7543 2443
rect 7607 2379 7641 2443
rect 7512 2368 7641 2379
rect -18 1838 111 1849
rect -18 1774 13 1838
rect 77 1774 111 1838
rect -18 1763 111 1774
rect 222 1836 351 1847
rect 222 1772 253 1836
rect 317 1772 351 1836
rect 222 1761 351 1772
rect 544 1835 673 1846
rect 544 1771 575 1835
rect 639 1771 673 1835
rect 544 1760 673 1771
rect 762 1836 891 1847
rect 762 1772 793 1836
rect 857 1772 891 1836
rect 762 1761 891 1772
rect 2666 1840 2795 1851
rect 2666 1776 2697 1840
rect 2761 1776 2795 1840
rect 2666 1765 2795 1776
rect 2991 1842 3120 1853
rect 2991 1778 3022 1842
rect 3086 1778 3120 1842
rect 2991 1767 3120 1778
rect 3259 1842 3388 1853
rect 3259 1778 3290 1842
rect 3354 1778 3388 1842
rect 3259 1767 3388 1778
rect 3525 1842 3654 1853
rect 3525 1778 3556 1842
rect 3620 1778 3654 1842
rect 3525 1767 3654 1778
rect 3765 1840 3894 1851
rect 3765 1776 3796 1840
rect 3860 1776 3894 1840
rect 3765 1765 3894 1776
rect 5559 1843 5688 1854
rect 5559 1779 5590 1843
rect 5654 1779 5688 1843
rect 5559 1768 5688 1779
rect 5925 1846 6054 1857
rect 5925 1782 5956 1846
rect 6020 1782 6054 1846
rect 5925 1771 6054 1782
rect 6169 1846 6298 1857
rect 6169 1782 6200 1846
rect 6264 1782 6298 1846
rect 6169 1771 6298 1782
rect 6592 1837 6721 1848
rect 6592 1773 6623 1837
rect 6687 1773 6721 1837
rect 6592 1762 6721 1773
rect 8535 1839 8664 1850
rect 8535 1775 8566 1839
rect 8630 1775 8664 1839
rect 8535 1764 8664 1775
rect 8787 1836 8916 1847
rect 8787 1772 8818 1836
rect 8882 1772 8916 1836
rect 8787 1761 8916 1772
rect 8993 1844 9122 1855
rect 8993 1780 9024 1844
rect 9088 1780 9122 1844
rect 8993 1769 9122 1780
rect 9276 1838 9405 1849
rect 9276 1774 9307 1838
rect 9371 1774 9405 1838
rect 9276 1763 9405 1774
rect 9574 1839 9703 1850
rect 9574 1775 9605 1839
rect 9669 1775 9703 1839
rect 9574 1764 9703 1775
rect 11406 1840 11535 1851
rect 11406 1776 11437 1840
rect 11501 1776 11535 1840
rect 11406 1765 11535 1776
rect 11616 1842 11745 1853
rect 11616 1778 11647 1842
rect 11711 1778 11745 1842
rect 11616 1767 11745 1778
rect 11967 1840 12096 1851
rect 11967 1776 11998 1840
rect 12062 1776 12096 1840
rect 11967 1765 12096 1776
rect 12247 1840 12376 1851
rect 12247 1776 12278 1840
rect 12342 1776 12376 1840
rect 12247 1765 12376 1776
rect 12564 1839 12693 1850
rect 12564 1775 12595 1839
rect 12659 1775 12693 1839
rect 12564 1764 12693 1775
rect 14354 1837 14483 1848
rect 14354 1773 14385 1837
rect 14449 1773 14483 1837
rect 14354 1762 14483 1773
rect 14649 1837 14778 1848
rect 14649 1773 14680 1837
rect 14744 1773 14778 1837
rect 14649 1762 14778 1773
rect 14936 1837 15065 1848
rect 14936 1773 14967 1837
rect 15031 1773 15065 1837
rect 14936 1762 15065 1773
rect 15226 1837 15355 1848
rect 15226 1773 15257 1837
rect 15321 1773 15355 1837
rect 15226 1762 15355 1773
rect 15510 1840 15639 1851
rect 15510 1776 15541 1840
rect 15605 1776 15639 1840
rect 15510 1765 15639 1776
rect 1173 1300 1302 1311
rect 1173 1236 1204 1300
rect 1268 1236 1302 1300
rect 1173 1225 1302 1236
rect 1390 1300 1519 1311
rect 1390 1236 1421 1300
rect 1485 1236 1519 1300
rect 1390 1225 1519 1236
rect 1609 1300 1738 1311
rect 1609 1236 1640 1300
rect 1704 1236 1738 1300
rect 1609 1225 1738 1236
rect 1822 1296 1951 1307
rect 1822 1232 1853 1296
rect 1917 1232 1951 1296
rect 1822 1221 1951 1232
rect 2033 1296 2162 1307
rect 2033 1232 2064 1296
rect 2128 1232 2162 1296
rect 2033 1221 2162 1232
rect 4157 1296 4286 1307
rect 4157 1232 4188 1296
rect 4252 1232 4286 1296
rect 4157 1221 4286 1232
rect 4435 1295 4564 1306
rect 4435 1231 4466 1295
rect 4530 1231 4564 1295
rect 4435 1220 4564 1231
rect 5007 1300 5136 1311
rect 5007 1236 5038 1300
rect 5102 1236 5136 1300
rect 5007 1225 5136 1236
rect 5246 1300 5375 1311
rect 5246 1236 5277 1300
rect 5341 1236 5375 1300
rect 5246 1225 5375 1236
rect 7404 1298 7533 1309
rect 7404 1234 7435 1298
rect 7499 1234 7533 1298
rect 7404 1223 7533 1234
rect 7631 1303 7760 1314
rect 7631 1239 7662 1303
rect 7726 1239 7760 1303
rect 7631 1228 7760 1239
rect 7821 1305 7950 1316
rect 7821 1241 7852 1305
rect 7916 1241 7950 1305
rect 7821 1230 7950 1241
rect 8037 1296 8166 1307
rect 8037 1232 8068 1296
rect 8132 1232 8166 1296
rect 8037 1221 8166 1232
rect 10018 1299 10147 1310
rect 10018 1235 10049 1299
rect 10113 1235 10147 1299
rect 10018 1224 10147 1235
rect 10247 1302 10376 1313
rect 10247 1238 10278 1302
rect 10342 1238 10376 1302
rect 10247 1227 10376 1238
rect 10473 1307 10602 1318
rect 10473 1243 10504 1307
rect 10568 1243 10602 1307
rect 10473 1232 10602 1243
rect 10701 1299 10830 1310
rect 10701 1235 10732 1299
rect 10796 1235 10830 1299
rect 10701 1224 10830 1235
rect 10937 1305 11066 1316
rect 10937 1241 10968 1305
rect 11032 1241 11066 1305
rect 10937 1230 11066 1241
rect 11129 1296 11258 1307
rect 11129 1232 11160 1296
rect 11224 1232 11258 1296
rect 11129 1221 11258 1232
rect 12864 1296 12993 1307
rect 12864 1232 12895 1296
rect 12959 1232 12993 1296
rect 12864 1221 12993 1232
rect 13068 1301 13197 1312
rect 13068 1237 13099 1301
rect 13163 1237 13197 1301
rect 13068 1226 13197 1237
rect 13259 1296 13388 1307
rect 13259 1232 13290 1296
rect 13354 1232 13388 1296
rect 13259 1221 13388 1232
rect 13461 1295 13590 1306
rect 13461 1231 13492 1295
rect 13556 1231 13590 1295
rect 13461 1220 13590 1231
rect 13751 1296 13880 1307
rect 13751 1232 13782 1296
rect 13846 1232 13880 1296
rect 13751 1221 13880 1232
rect 14036 1295 14165 1306
rect 14036 1231 14067 1295
rect 14131 1231 14165 1295
rect 14036 1220 14165 1231
rect 15791 1300 15920 1311
rect 15791 1236 15822 1300
rect 15886 1236 15920 1300
rect 15791 1225 15920 1236
rect 15985 1304 16114 1315
rect 15985 1240 16016 1304
rect 16080 1240 16114 1304
rect 15985 1229 16114 1240
rect 16174 1301 16303 1312
rect 16174 1237 16205 1301
rect 16269 1237 16303 1301
rect 16174 1226 16303 1237
rect 16397 1303 16526 1314
rect 16397 1239 16428 1303
rect 16492 1239 16526 1303
rect 16397 1228 16526 1239
rect 228 1155 357 1166
rect 228 1091 259 1155
rect 323 1091 357 1155
rect 228 1080 357 1091
rect 430 1151 559 1162
rect 430 1087 461 1151
rect 525 1087 559 1151
rect 430 1076 559 1087
rect 619 1148 748 1159
rect 619 1084 650 1148
rect 714 1084 748 1148
rect 619 1073 748 1084
rect 848 1149 977 1160
rect 848 1085 879 1149
rect 943 1085 977 1149
rect 848 1074 977 1085
rect 2617 1152 2746 1163
rect 2617 1088 2648 1152
rect 2712 1088 2746 1152
rect 2617 1077 2746 1088
rect 2832 1149 2961 1160
rect 2832 1085 2863 1149
rect 2927 1085 2961 1149
rect 2832 1074 2961 1085
rect 3030 1146 3159 1157
rect 3030 1082 3061 1146
rect 3125 1082 3159 1146
rect 3030 1071 3159 1082
rect 3225 1156 3354 1167
rect 3225 1092 3256 1156
rect 3320 1092 3354 1156
rect 3225 1081 3354 1092
rect 3505 1154 3634 1165
rect 3505 1090 3536 1154
rect 3600 1090 3634 1154
rect 3505 1079 3634 1090
rect 3724 1152 3853 1163
rect 3724 1088 3755 1152
rect 3819 1088 3853 1152
rect 3724 1077 3853 1088
rect 5545 1149 5674 1160
rect 5545 1085 5576 1149
rect 5640 1085 5674 1149
rect 5545 1074 5674 1085
rect 5896 1146 6025 1157
rect 5896 1082 5927 1146
rect 5991 1082 6025 1146
rect 5896 1071 6025 1082
rect 6085 1144 6214 1155
rect 6085 1080 6116 1144
rect 6180 1080 6214 1144
rect 6085 1069 6214 1080
rect 6290 1151 6419 1162
rect 6290 1087 6321 1151
rect 6385 1087 6419 1151
rect 6290 1076 6419 1087
rect 6481 1153 6610 1164
rect 6481 1089 6512 1153
rect 6576 1089 6610 1153
rect 6481 1078 6610 1089
rect 8526 1155 8655 1166
rect 8526 1091 8557 1155
rect 8621 1091 8655 1155
rect 8526 1080 8655 1091
rect 8716 1157 8845 1168
rect 8716 1093 8747 1157
rect 8811 1093 8845 1157
rect 8716 1082 8845 1093
rect 8910 1155 9039 1166
rect 8910 1091 8941 1155
rect 9005 1091 9039 1155
rect 8910 1080 9039 1091
rect 9221 1151 9350 1162
rect 9221 1087 9252 1151
rect 9316 1087 9350 1151
rect 9221 1076 9350 1087
rect 11404 1150 11533 1161
rect 11404 1086 11435 1150
rect 11499 1086 11533 1150
rect 11404 1075 11533 1086
rect 11608 1150 11737 1161
rect 11608 1086 11639 1150
rect 11703 1086 11737 1150
rect 11608 1075 11737 1086
rect 12173 1146 12302 1157
rect 12173 1082 12204 1146
rect 12268 1082 12302 1146
rect 12173 1071 12302 1082
rect 12412 1148 12541 1159
rect 12412 1084 12443 1148
rect 12507 1084 12541 1148
rect 12412 1073 12541 1084
rect 12616 1148 12745 1159
rect 12616 1084 12647 1148
rect 12711 1084 12745 1148
rect 12616 1073 12745 1084
rect 14576 1156 14705 1167
rect 14576 1092 14607 1156
rect 14671 1092 14705 1156
rect 14576 1081 14705 1092
rect 14809 1154 14938 1165
rect 14809 1090 14840 1154
rect 14904 1090 14938 1154
rect 14809 1079 14938 1090
rect 15016 1152 15145 1163
rect 15016 1088 15047 1152
rect 15111 1088 15145 1152
rect 15016 1077 15145 1088
rect 15225 1154 15354 1165
rect 15225 1090 15256 1154
rect 15320 1090 15354 1154
rect 15225 1079 15354 1090
rect 15505 1156 15634 1167
rect 15505 1092 15536 1156
rect 15600 1092 15634 1156
rect 15505 1081 15634 1092
rect 1384 618 1513 629
rect 1155 606 1284 617
rect 1155 542 1186 606
rect 1250 542 1284 606
rect 1384 554 1415 618
rect 1479 554 1513 618
rect 1384 543 1513 554
rect 1603 608 1732 619
rect 1603 544 1634 608
rect 1698 544 1732 608
rect 1155 531 1284 542
rect 1603 533 1732 544
rect 1795 612 1924 623
rect 1795 548 1826 612
rect 1890 548 1924 612
rect 1795 537 1924 548
rect 2289 610 2418 621
rect 2289 546 2320 610
rect 2384 546 2418 610
rect 2289 535 2418 546
rect 4081 609 4210 620
rect 4081 545 4112 609
rect 4176 545 4210 609
rect 4081 534 4210 545
rect 4474 607 4603 618
rect 4474 543 4505 607
rect 4569 543 4603 607
rect 4474 532 4603 543
rect 4671 615 4800 626
rect 4671 551 4702 615
rect 4766 551 4800 615
rect 4671 540 4800 551
rect 5001 617 5130 628
rect 5001 553 5032 617
rect 5096 553 5130 617
rect 5001 542 5130 553
rect 5197 617 5326 628
rect 5197 553 5228 617
rect 5292 553 5326 617
rect 5197 542 5326 553
rect 7104 610 7233 621
rect 7104 546 7135 610
rect 7199 546 7233 610
rect 7104 535 7233 546
rect 7405 614 7534 625
rect 7405 550 7436 614
rect 7500 550 7534 614
rect 7405 539 7534 550
rect 7611 615 7740 626
rect 7611 551 7642 615
rect 7706 551 7740 615
rect 7611 540 7740 551
rect 7821 611 7950 622
rect 7821 547 7852 611
rect 7916 547 7950 611
rect 7821 536 7950 547
rect 8032 617 8161 628
rect 8032 553 8063 617
rect 8127 553 8161 617
rect 8032 542 8161 553
rect 9912 606 10041 617
rect 9912 542 9943 606
rect 10007 542 10041 606
rect 9912 531 10041 542
rect 10169 613 10298 624
rect 10169 549 10200 613
rect 10264 549 10298 613
rect 10169 538 10298 549
rect 10419 609 10548 620
rect 10419 545 10450 609
rect 10514 545 10548 609
rect 10419 534 10548 545
rect 10690 614 10819 625
rect 10690 550 10721 614
rect 10785 550 10819 614
rect 10690 539 10819 550
rect 10931 617 11060 628
rect 10931 553 10962 617
rect 11026 553 11060 617
rect 10931 542 11060 553
rect 11156 613 11285 624
rect 11156 549 11187 613
rect 11251 549 11285 613
rect 11156 538 11285 549
rect 12863 611 12992 622
rect 12863 547 12894 611
rect 12958 547 12992 611
rect 12863 536 12992 547
rect 13064 612 13193 623
rect 13064 548 13095 612
rect 13159 548 13193 612
rect 13064 537 13193 548
rect 13282 608 13411 619
rect 13282 544 13313 608
rect 13377 544 13411 608
rect 13282 533 13411 544
rect 13489 612 13618 623
rect 13489 548 13520 612
rect 13584 548 13618 612
rect 13489 537 13618 548
rect 13694 611 13823 622
rect 13694 547 13725 611
rect 13789 547 13823 611
rect 13694 536 13823 547
rect 14041 607 14170 618
rect 14041 543 14072 607
rect 14136 543 14170 607
rect 14041 532 14170 543
rect 15793 611 15922 622
rect 15793 547 15824 611
rect 15888 547 15922 611
rect 15793 536 15922 547
rect 15984 614 16113 625
rect 15984 550 16015 614
rect 16079 550 16113 614
rect 15984 539 16113 550
rect 16179 616 16308 627
rect 16179 552 16210 616
rect 16274 552 16308 616
rect 16179 541 16308 552
rect 16626 611 16755 622
rect 16626 547 16657 611
rect 16721 547 16755 611
rect 16626 536 16755 547
rect 10 462 139 473
rect 10 398 41 462
rect 105 398 139 462
rect 10 387 139 398
rect 243 458 372 469
rect 243 394 274 458
rect 338 394 372 458
rect 243 383 372 394
rect 458 465 587 476
rect 458 401 489 465
rect 553 401 587 465
rect 458 390 587 401
rect 676 462 805 473
rect 676 398 707 462
rect 771 398 805 462
rect 676 387 805 398
rect 892 463 1021 474
rect 892 399 923 463
rect 987 399 1021 463
rect 892 388 1021 399
rect 2613 459 2742 470
rect 2613 395 2644 459
rect 2708 395 2742 459
rect 2613 384 2742 395
rect 2803 459 2932 470
rect 2803 395 2834 459
rect 2898 395 2932 459
rect 2803 384 2932 395
rect 3013 462 3142 473
rect 3013 398 3044 462
rect 3108 398 3142 462
rect 3013 387 3142 398
rect 3230 459 3359 470
rect 3230 395 3261 459
rect 3325 395 3359 459
rect 3230 384 3359 395
rect 3525 462 3654 473
rect 3525 398 3556 462
rect 3620 398 3654 462
rect 3525 387 3654 398
rect 3749 467 3878 478
rect 3749 403 3780 467
rect 3844 403 3878 467
rect 3749 392 3878 403
rect 5627 460 5756 471
rect 5627 396 5658 460
rect 5722 396 5756 460
rect 5627 385 5756 396
rect 5927 458 6056 469
rect 5927 394 5958 458
rect 6022 394 6056 458
rect 5927 383 6056 394
rect 6179 462 6308 473
rect 6179 398 6210 462
rect 6274 398 6308 462
rect 6179 387 6308 398
rect 6396 467 6525 478
rect 6396 403 6427 467
rect 6491 403 6525 467
rect 6396 392 6525 403
rect 6597 464 6726 475
rect 6597 400 6628 464
rect 6692 400 6726 464
rect 6597 389 6726 400
rect 8482 455 8611 466
rect 8482 391 8513 455
rect 8577 391 8611 455
rect 8482 380 8611 391
rect 8674 455 8803 466
rect 8674 391 8705 455
rect 8769 391 8803 455
rect 8674 380 8803 391
rect 8874 455 9003 466
rect 8874 391 8905 455
rect 8969 391 9003 455
rect 8874 380 9003 391
rect 9492 463 9621 474
rect 9492 399 9523 463
rect 9587 399 9621 463
rect 9492 388 9621 399
rect 11393 459 11522 470
rect 11393 395 11424 459
rect 11488 395 11522 459
rect 11393 384 11522 395
rect 11649 459 11778 470
rect 11649 395 11680 459
rect 11744 395 11778 459
rect 11649 384 11778 395
rect 11884 459 12013 470
rect 11884 395 11915 459
rect 11979 395 12013 459
rect 11884 384 12013 395
rect 12173 461 12302 472
rect 12173 397 12204 461
rect 12268 397 12302 461
rect 12173 386 12302 397
rect 12363 459 12492 470
rect 12363 395 12394 459
rect 12458 395 12492 459
rect 12363 384 12492 395
rect 12567 461 12696 472
rect 12567 397 12598 461
rect 12662 397 12696 461
rect 12567 386 12696 397
rect 14353 467 14482 478
rect 14353 403 14384 467
rect 14448 403 14482 467
rect 14353 392 14482 403
rect 14595 463 14724 474
rect 14595 399 14626 463
rect 14690 399 14724 463
rect 14595 388 14724 399
rect 14795 462 14924 473
rect 14795 398 14826 462
rect 14890 398 14924 462
rect 14795 387 14924 398
rect 14985 470 15114 481
rect 14985 406 15016 470
rect 15080 406 15114 470
rect 14985 395 15114 406
rect 15206 468 15335 479
rect 15206 404 15237 468
rect 15301 404 15335 468
rect 15206 393 15335 404
rect 15502 463 15631 474
rect 15502 399 15533 463
rect 15597 399 15631 463
rect 15502 388 15631 399
rect 384 -70 513 -59
rect 384 -134 415 -70
rect 479 -134 513 -70
rect 384 -145 513 -134
rect 583 -73 712 -62
rect 583 -137 614 -73
rect 678 -137 712 -73
rect 583 -148 712 -137
rect 794 -73 923 -62
rect 794 -137 825 -73
rect 889 -137 923 -73
rect 794 -148 923 -137
rect 1000 -73 1129 -62
rect 1000 -137 1031 -73
rect 1095 -137 1129 -73
rect 1000 -148 1129 -137
rect 1228 -75 1357 -64
rect 1228 -139 1259 -75
rect 1323 -139 1357 -75
rect 1228 -150 1357 -139
rect 1472 -75 1601 -64
rect 1472 -139 1503 -75
rect 1567 -139 1601 -75
rect 1472 -150 1601 -139
rect 1702 -73 1831 -62
rect 1702 -137 1733 -73
rect 1797 -137 1831 -73
rect 1702 -148 1831 -137
rect 1908 -73 2037 -62
rect 1908 -137 1939 -73
rect 2003 -137 2037 -73
rect 1908 -148 2037 -137
rect 2126 -68 2255 -57
rect 2126 -132 2157 -68
rect 2221 -132 2255 -68
rect 2126 -143 2255 -132
rect 2329 -74 2458 -63
rect 2329 -138 2360 -74
rect 2424 -138 2458 -74
rect 2329 -149 2458 -138
rect 2537 -71 2666 -60
rect 2537 -135 2568 -71
rect 2632 -135 2666 -71
rect 2537 -146 2666 -135
rect 2800 -75 2929 -64
rect 2800 -139 2831 -75
rect 2895 -139 2929 -75
rect 2800 -150 2929 -139
rect 3008 -74 3137 -63
rect 3008 -138 3039 -74
rect 3103 -138 3137 -74
rect 3008 -149 3137 -138
rect 3218 -77 3347 -66
rect 3218 -141 3249 -77
rect 3313 -141 3347 -77
rect 3218 -152 3347 -141
rect 3418 -71 3547 -60
rect 3418 -135 3449 -71
rect 3513 -135 3547 -71
rect 3418 -146 3547 -135
rect 3621 -74 3750 -63
rect 3621 -138 3652 -74
rect 3716 -138 3750 -74
rect 3621 -149 3750 -138
rect 3831 -74 3960 -63
rect 3831 -138 3862 -74
rect 3926 -138 3960 -74
rect 3831 -149 3960 -138
rect 4032 -73 4161 -62
rect 4032 -137 4063 -73
rect 4127 -137 4161 -73
rect 4032 -148 4161 -137
rect 4248 -72 4377 -61
rect 4248 -136 4279 -72
rect 4343 -136 4377 -72
rect 4248 -147 4377 -136
rect 4529 -74 4658 -63
rect 4529 -138 4560 -74
rect 4624 -138 4658 -74
rect 4529 -149 4658 -138
rect 4749 -79 4878 -68
rect 4749 -143 4780 -79
rect 4844 -143 4878 -79
rect 4749 -154 4878 -143
rect 4954 -78 5083 -67
rect 4954 -142 4985 -78
rect 5049 -142 5083 -78
rect 4954 -153 5083 -142
rect 5175 -72 5304 -61
rect 5175 -136 5206 -72
rect 5270 -136 5304 -72
rect 5175 -147 5304 -136
rect 5380 -79 5509 -68
rect 5380 -143 5411 -79
rect 5475 -143 5509 -79
rect 5380 -154 5509 -143
rect 5589 -78 5718 -67
rect 5589 -142 5620 -78
rect 5684 -142 5718 -78
rect 5589 -153 5718 -142
rect 5806 -78 5935 -67
rect 5806 -142 5837 -78
rect 5901 -142 5935 -78
rect 5806 -153 5935 -142
rect 6020 -73 6149 -62
rect 6020 -137 6051 -73
rect 6115 -137 6149 -73
rect 6020 -148 6149 -137
rect 6215 -75 6344 -64
rect 6215 -139 6246 -75
rect 6310 -139 6344 -75
rect 6215 -150 6344 -139
rect 6410 -78 6539 -67
rect 6410 -142 6441 -78
rect 6505 -142 6539 -78
rect 6410 -153 6539 -142
rect 6612 -75 6741 -64
rect 6612 -139 6643 -75
rect 6707 -139 6741 -75
rect 6612 -150 6741 -139
rect 6896 -74 7025 -63
rect 6896 -138 6927 -74
rect 6991 -138 7025 -74
rect 6896 -149 7025 -138
rect 7095 -73 7224 -62
rect 7095 -137 7126 -73
rect 7190 -137 7224 -73
rect 7095 -148 7224 -137
rect 7298 -71 7427 -60
rect 7298 -135 7329 -71
rect 7393 -135 7427 -71
rect 7298 -146 7427 -135
rect 7563 -74 7692 -63
rect 7563 -138 7594 -74
rect 7658 -138 7692 -74
rect 7563 -149 7692 -138
rect 7761 -75 7890 -64
rect 7761 -139 7792 -75
rect 7856 -139 7890 -75
rect 7761 -150 7890 -139
rect 7950 -73 8079 -62
rect 7950 -137 7981 -73
rect 8045 -137 8079 -73
rect 7950 -148 8079 -137
rect 8162 -73 8291 -62
rect 8162 -137 8193 -73
rect 8257 -137 8291 -73
rect 8162 -148 8291 -137
rect 8379 -73 8508 -62
rect 8379 -137 8410 -73
rect 8474 -137 8508 -73
rect 8379 -148 8508 -137
rect 8584 -77 8713 -66
rect 8584 -141 8615 -77
rect 8679 -141 8713 -77
rect 8584 -152 8713 -141
rect 8789 -77 8918 -66
rect 8789 -141 8820 -77
rect 8884 -141 8918 -77
rect 8789 -152 8918 -141
rect 8997 -72 9126 -61
rect 8997 -136 9028 -72
rect 9092 -136 9126 -72
rect 8997 -147 9126 -136
rect 9280 -73 9409 -62
rect 9280 -137 9311 -73
rect 9375 -137 9409 -73
rect 9280 -148 9409 -137
rect 9473 -75 9602 -64
rect 9473 -139 9504 -75
rect 9568 -139 9602 -75
rect 9473 -150 9602 -139
rect 9699 -77 9828 -66
rect 9699 -141 9730 -77
rect 9794 -141 9828 -77
rect 9699 -152 9828 -141
rect 9964 -77 10093 -66
rect 9964 -141 9995 -77
rect 10059 -141 10093 -77
rect 9964 -152 10093 -141
rect 10158 -73 10287 -62
rect 10158 -137 10189 -73
rect 10253 -137 10287 -73
rect 10158 -148 10287 -137
rect 10356 -82 10485 -71
rect 10356 -146 10387 -82
rect 10451 -146 10485 -82
rect 10356 -157 10485 -146
rect 10560 -74 10689 -63
rect 10560 -138 10591 -74
rect 10655 -138 10689 -74
rect 10560 -149 10689 -138
rect 10780 -71 10909 -60
rect 10780 -135 10811 -71
rect 10875 -135 10909 -71
rect 10780 -146 10909 -135
rect 10995 -75 11124 -64
rect 10995 -139 11026 -75
rect 11090 -139 11124 -75
rect 10995 -150 11124 -139
rect 11223 -72 11352 -61
rect 11223 -136 11254 -72
rect 11318 -136 11352 -72
rect 11223 -147 11352 -136
rect 11427 -75 11556 -64
rect 11427 -139 11458 -75
rect 11522 -139 11556 -75
rect 11427 -150 11556 -139
rect 11665 -73 11794 -62
rect 11665 -137 11696 -73
rect 11760 -137 11794 -73
rect 11665 -148 11794 -137
rect 11858 -72 11987 -61
rect 11858 -136 11889 -72
rect 11953 -136 11987 -72
rect 11858 -147 11987 -136
rect 12055 -77 12184 -66
rect 12055 -141 12086 -77
rect 12150 -141 12184 -77
rect 12055 -152 12184 -141
rect 12311 -74 12440 -63
rect 12311 -138 12342 -74
rect 12406 -138 12440 -74
rect 12311 -149 12440 -138
rect 12550 -78 12679 -67
rect 12550 -142 12581 -78
rect 12645 -142 12679 -78
rect 12550 -153 12679 -142
rect 12783 -82 12912 -71
rect 12783 -146 12814 -82
rect 12878 -146 12912 -82
rect 12783 -157 12912 -146
rect 13004 -77 13133 -66
rect 13004 -141 13035 -77
rect 13099 -141 13133 -77
rect 13004 -152 13133 -141
rect 13195 -77 13324 -66
rect 13195 -141 13226 -77
rect 13290 -141 13324 -77
rect 13195 -152 13324 -141
rect 13423 -75 13552 -64
rect 13423 -139 13454 -75
rect 13518 -139 13552 -75
rect 13423 -150 13552 -139
rect 13620 -80 13749 -69
rect 13620 -144 13651 -80
rect 13715 -144 13749 -80
rect 13620 -155 13749 -144
rect 13832 -80 13961 -69
rect 13832 -144 13863 -80
rect 13927 -144 13961 -80
rect 13832 -155 13961 -144
rect 14059 -77 14188 -66
rect 14059 -141 14090 -77
rect 14154 -141 14188 -77
rect 14059 -152 14188 -141
rect 14248 -76 14377 -65
rect 14248 -140 14279 -76
rect 14343 -140 14377 -76
rect 14248 -151 14377 -140
rect 14474 -75 14603 -64
rect 14474 -139 14505 -75
rect 14569 -139 14603 -75
rect 14474 -150 14603 -139
rect 14728 -75 14857 -64
rect 14728 -139 14759 -75
rect 14823 -139 14857 -75
rect 14728 -150 14857 -139
rect 14972 -78 15101 -67
rect 14972 -142 15003 -78
rect 15067 -142 15101 -78
rect 14972 -153 15101 -142
rect 15202 -79 15331 -68
rect 15202 -143 15233 -79
rect 15297 -143 15331 -79
rect 15202 -154 15331 -143
rect 15460 -76 15589 -65
rect 15460 -140 15491 -76
rect 15555 -140 15589 -76
rect 15460 -151 15589 -140
rect 15670 -76 15799 -65
rect 15670 -140 15701 -76
rect 15765 -140 15799 -76
rect 15670 -151 15799 -140
rect 15895 -76 16024 -65
rect 15895 -140 15926 -76
rect 15990 -140 16024 -76
rect 15895 -151 16024 -140
rect 16114 -79 16243 -68
rect 16114 -143 16145 -79
rect 16209 -143 16243 -79
rect 16114 -154 16243 -143
rect 16460 -75 16589 -64
rect 16460 -139 16491 -75
rect 16555 -139 16589 -75
rect 16460 -150 16589 -139
rect 16659 -78 16788 -67
rect 16659 -142 16690 -78
rect 16754 -142 16788 -78
rect 16659 -153 16788 -142
<< via3 >>
rect 47 2978 111 2982
rect 47 2922 51 2978
rect 51 2922 107 2978
rect 107 2922 111 2978
rect 47 2918 111 2922
rect 249 2980 313 2984
rect 249 2924 253 2980
rect 253 2924 309 2980
rect 309 2924 313 2980
rect 249 2920 313 2924
rect 460 2978 524 2982
rect 460 2922 464 2978
rect 464 2922 520 2978
rect 520 2922 524 2978
rect 460 2918 524 2922
rect 650 2978 714 2982
rect 650 2922 654 2978
rect 654 2922 710 2978
rect 710 2922 714 2978
rect 650 2918 714 2922
rect 858 2980 922 2984
rect 858 2924 862 2980
rect 862 2924 918 2980
rect 918 2924 922 2980
rect 858 2920 922 2924
rect 1060 2980 1124 2984
rect 1060 2924 1064 2980
rect 1064 2924 1120 2980
rect 1120 2924 1124 2980
rect 1060 2920 1124 2924
rect 1259 2982 1323 2986
rect 1259 2926 1263 2982
rect 1263 2926 1319 2982
rect 1319 2926 1323 2982
rect 1259 2922 1323 2926
rect 1454 2979 1518 2983
rect 1454 2923 1458 2979
rect 1458 2923 1514 2979
rect 1514 2923 1518 2979
rect 1454 2919 1518 2923
rect 1655 2981 1719 2985
rect 1655 2925 1659 2981
rect 1659 2925 1715 2981
rect 1715 2925 1719 2981
rect 1655 2921 1719 2925
rect 1872 2979 1936 2983
rect 1872 2923 1876 2979
rect 1876 2923 1932 2979
rect 1932 2923 1936 2979
rect 1872 2919 1936 2923
rect 2146 2982 2210 2986
rect 2146 2926 2150 2982
rect 2150 2926 2206 2982
rect 2206 2926 2210 2982
rect 2146 2922 2210 2926
rect 2423 2975 2487 2979
rect 2423 2919 2427 2975
rect 2427 2919 2483 2975
rect 2483 2919 2487 2975
rect 2423 2915 2487 2919
rect 2646 2978 2710 2982
rect 2646 2922 2650 2978
rect 2650 2922 2706 2978
rect 2706 2922 2710 2978
rect 2646 2918 2710 2922
rect 2878 2977 2942 2981
rect 2878 2921 2882 2977
rect 2882 2921 2938 2977
rect 2938 2921 2942 2977
rect 2878 2917 2942 2921
rect 4514 2974 4578 2978
rect 4514 2918 4518 2974
rect 4518 2918 4574 2974
rect 4574 2918 4578 2974
rect 4514 2914 4578 2918
rect 4822 2975 4886 2979
rect 4822 2919 4826 2975
rect 4826 2919 4882 2975
rect 4882 2919 4886 2975
rect 4822 2915 4886 2919
rect 5022 2976 5086 2980
rect 5022 2920 5026 2976
rect 5026 2920 5082 2976
rect 5082 2920 5086 2976
rect 5022 2916 5086 2920
rect 5241 2975 5305 2979
rect 5241 2919 5245 2975
rect 5245 2919 5301 2975
rect 5301 2919 5305 2975
rect 5241 2915 5305 2919
rect 5487 2974 5551 2978
rect 5487 2918 5491 2974
rect 5491 2918 5547 2974
rect 5547 2918 5551 2974
rect 5487 2914 5551 2918
rect 5695 2976 5759 2980
rect 5695 2920 5699 2976
rect 5699 2920 5755 2976
rect 5755 2920 5759 2976
rect 5695 2916 5759 2920
rect 5897 2977 5961 2981
rect 5897 2921 5901 2977
rect 5901 2921 5957 2977
rect 5957 2921 5961 2977
rect 5897 2917 5961 2921
rect 6090 2976 6154 2980
rect 6090 2920 6094 2976
rect 6094 2920 6150 2976
rect 6150 2920 6154 2976
rect 6090 2916 6154 2920
rect 6462 2975 6526 2979
rect 6462 2919 6466 2975
rect 6466 2919 6522 2975
rect 6522 2919 6526 2975
rect 6462 2915 6526 2919
rect 6651 2973 6715 2977
rect 6651 2917 6655 2973
rect 6655 2917 6711 2973
rect 6711 2917 6715 2973
rect 6651 2913 6715 2917
rect 6941 2973 7005 2977
rect 6941 2917 6945 2973
rect 6945 2917 7001 2973
rect 7001 2917 7005 2973
rect 6941 2913 7005 2917
rect 7214 2975 7278 2979
rect 7214 2919 7218 2975
rect 7218 2919 7274 2975
rect 7274 2919 7278 2975
rect 7214 2915 7278 2919
rect 1165 2439 1229 2443
rect 1165 2383 1169 2439
rect 1169 2383 1225 2439
rect 1225 2383 1229 2439
rect 1165 2379 1229 2383
rect 1384 2443 1448 2447
rect 1384 2387 1388 2443
rect 1388 2387 1444 2443
rect 1444 2387 1448 2443
rect 1384 2383 1448 2387
rect 1667 2443 1731 2447
rect 1667 2387 1671 2443
rect 1671 2387 1727 2443
rect 1727 2387 1731 2443
rect 1667 2383 1731 2387
rect 1876 2443 1940 2447
rect 1876 2387 1880 2443
rect 1880 2387 1936 2443
rect 1936 2387 1940 2443
rect 1876 2383 1940 2387
rect 2147 2441 2211 2445
rect 2147 2385 2151 2441
rect 2151 2385 2207 2441
rect 2207 2385 2211 2441
rect 2147 2381 2211 2385
rect 4222 2439 4286 2443
rect 4222 2383 4226 2439
rect 4226 2383 4282 2439
rect 4282 2383 4286 2439
rect 4222 2379 4286 2383
rect 4471 2442 4535 2446
rect 4471 2386 4475 2442
rect 4475 2386 4531 2442
rect 4531 2386 4535 2442
rect 4471 2382 4535 2386
rect 4815 2428 4879 2432
rect 4815 2372 4819 2428
rect 4819 2372 4875 2428
rect 4875 2372 4879 2428
rect 4815 2368 4879 2372
rect 5069 2434 5133 2438
rect 5069 2378 5073 2434
rect 5073 2378 5129 2434
rect 5129 2378 5133 2434
rect 5069 2374 5133 2378
rect 5298 2434 5362 2438
rect 5298 2378 5302 2434
rect 5302 2378 5358 2434
rect 5358 2378 5362 2434
rect 5298 2374 5362 2378
rect 7016 2439 7080 2443
rect 7016 2383 7020 2439
rect 7020 2383 7076 2439
rect 7076 2383 7080 2439
rect 7016 2379 7080 2383
rect 7220 2441 7284 2445
rect 7220 2385 7224 2441
rect 7224 2385 7280 2441
rect 7280 2385 7284 2441
rect 7220 2381 7284 2385
rect 7543 2439 7607 2443
rect 7543 2383 7547 2439
rect 7547 2383 7603 2439
rect 7603 2383 7607 2439
rect 7543 2379 7607 2383
rect 13 1834 77 1838
rect 13 1778 17 1834
rect 17 1778 73 1834
rect 73 1778 77 1834
rect 13 1774 77 1778
rect 253 1832 317 1836
rect 253 1776 257 1832
rect 257 1776 313 1832
rect 313 1776 317 1832
rect 253 1772 317 1776
rect 575 1831 639 1835
rect 575 1775 579 1831
rect 579 1775 635 1831
rect 635 1775 639 1831
rect 575 1771 639 1775
rect 793 1832 857 1836
rect 793 1776 797 1832
rect 797 1776 853 1832
rect 853 1776 857 1832
rect 793 1772 857 1776
rect 2697 1836 2761 1840
rect 2697 1780 2701 1836
rect 2701 1780 2757 1836
rect 2757 1780 2761 1836
rect 2697 1776 2761 1780
rect 3022 1838 3086 1842
rect 3022 1782 3026 1838
rect 3026 1782 3082 1838
rect 3082 1782 3086 1838
rect 3022 1778 3086 1782
rect 3290 1838 3354 1842
rect 3290 1782 3294 1838
rect 3294 1782 3350 1838
rect 3350 1782 3354 1838
rect 3290 1778 3354 1782
rect 3556 1838 3620 1842
rect 3556 1782 3560 1838
rect 3560 1782 3616 1838
rect 3616 1782 3620 1838
rect 3556 1778 3620 1782
rect 3796 1836 3860 1840
rect 3796 1780 3800 1836
rect 3800 1780 3856 1836
rect 3856 1780 3860 1836
rect 3796 1776 3860 1780
rect 5590 1839 5654 1843
rect 5590 1783 5594 1839
rect 5594 1783 5650 1839
rect 5650 1783 5654 1839
rect 5590 1779 5654 1783
rect 5956 1842 6020 1846
rect 5956 1786 5960 1842
rect 5960 1786 6016 1842
rect 6016 1786 6020 1842
rect 5956 1782 6020 1786
rect 6200 1842 6264 1846
rect 6200 1786 6204 1842
rect 6204 1786 6260 1842
rect 6260 1786 6264 1842
rect 6200 1782 6264 1786
rect 6623 1833 6687 1837
rect 6623 1777 6627 1833
rect 6627 1777 6683 1833
rect 6683 1777 6687 1833
rect 6623 1773 6687 1777
rect 8566 1835 8630 1839
rect 8566 1779 8570 1835
rect 8570 1779 8626 1835
rect 8626 1779 8630 1835
rect 8566 1775 8630 1779
rect 8818 1832 8882 1836
rect 8818 1776 8822 1832
rect 8822 1776 8878 1832
rect 8878 1776 8882 1832
rect 8818 1772 8882 1776
rect 9024 1840 9088 1844
rect 9024 1784 9028 1840
rect 9028 1784 9084 1840
rect 9084 1784 9088 1840
rect 9024 1780 9088 1784
rect 9307 1834 9371 1838
rect 9307 1778 9311 1834
rect 9311 1778 9367 1834
rect 9367 1778 9371 1834
rect 9307 1774 9371 1778
rect 9605 1835 9669 1839
rect 9605 1779 9609 1835
rect 9609 1779 9665 1835
rect 9665 1779 9669 1835
rect 9605 1775 9669 1779
rect 11437 1836 11501 1840
rect 11437 1780 11441 1836
rect 11441 1780 11497 1836
rect 11497 1780 11501 1836
rect 11437 1776 11501 1780
rect 11647 1838 11711 1842
rect 11647 1782 11651 1838
rect 11651 1782 11707 1838
rect 11707 1782 11711 1838
rect 11647 1778 11711 1782
rect 11998 1836 12062 1840
rect 11998 1780 12002 1836
rect 12002 1780 12058 1836
rect 12058 1780 12062 1836
rect 11998 1776 12062 1780
rect 12278 1836 12342 1840
rect 12278 1780 12282 1836
rect 12282 1780 12338 1836
rect 12338 1780 12342 1836
rect 12278 1776 12342 1780
rect 12595 1835 12659 1839
rect 12595 1779 12599 1835
rect 12599 1779 12655 1835
rect 12655 1779 12659 1835
rect 12595 1775 12659 1779
rect 14385 1833 14449 1837
rect 14385 1777 14389 1833
rect 14389 1777 14445 1833
rect 14445 1777 14449 1833
rect 14385 1773 14449 1777
rect 14680 1833 14744 1837
rect 14680 1777 14684 1833
rect 14684 1777 14740 1833
rect 14740 1777 14744 1833
rect 14680 1773 14744 1777
rect 14967 1833 15031 1837
rect 14967 1777 14971 1833
rect 14971 1777 15027 1833
rect 15027 1777 15031 1833
rect 14967 1773 15031 1777
rect 15257 1833 15321 1837
rect 15257 1777 15261 1833
rect 15261 1777 15317 1833
rect 15317 1777 15321 1833
rect 15257 1773 15321 1777
rect 15541 1836 15605 1840
rect 15541 1780 15545 1836
rect 15545 1780 15601 1836
rect 15601 1780 15605 1836
rect 15541 1776 15605 1780
rect 1204 1296 1268 1300
rect 1204 1240 1208 1296
rect 1208 1240 1264 1296
rect 1264 1240 1268 1296
rect 1204 1236 1268 1240
rect 1421 1296 1485 1300
rect 1421 1240 1425 1296
rect 1425 1240 1481 1296
rect 1481 1240 1485 1296
rect 1421 1236 1485 1240
rect 1640 1296 1704 1300
rect 1640 1240 1644 1296
rect 1644 1240 1700 1296
rect 1700 1240 1704 1296
rect 1640 1236 1704 1240
rect 1853 1292 1917 1296
rect 1853 1236 1857 1292
rect 1857 1236 1913 1292
rect 1913 1236 1917 1292
rect 1853 1232 1917 1236
rect 2064 1292 2128 1296
rect 2064 1236 2068 1292
rect 2068 1236 2124 1292
rect 2124 1236 2128 1292
rect 2064 1232 2128 1236
rect 4188 1292 4252 1296
rect 4188 1236 4192 1292
rect 4192 1236 4248 1292
rect 4248 1236 4252 1292
rect 4188 1232 4252 1236
rect 4466 1291 4530 1295
rect 4466 1235 4470 1291
rect 4470 1235 4526 1291
rect 4526 1235 4530 1291
rect 4466 1231 4530 1235
rect 5038 1296 5102 1300
rect 5038 1240 5042 1296
rect 5042 1240 5098 1296
rect 5098 1240 5102 1296
rect 5038 1236 5102 1240
rect 5277 1296 5341 1300
rect 5277 1240 5281 1296
rect 5281 1240 5337 1296
rect 5337 1240 5341 1296
rect 5277 1236 5341 1240
rect 7435 1294 7499 1298
rect 7435 1238 7439 1294
rect 7439 1238 7495 1294
rect 7495 1238 7499 1294
rect 7435 1234 7499 1238
rect 7662 1299 7726 1303
rect 7662 1243 7666 1299
rect 7666 1243 7722 1299
rect 7722 1243 7726 1299
rect 7662 1239 7726 1243
rect 7852 1301 7916 1305
rect 7852 1245 7856 1301
rect 7856 1245 7912 1301
rect 7912 1245 7916 1301
rect 7852 1241 7916 1245
rect 8068 1292 8132 1296
rect 8068 1236 8072 1292
rect 8072 1236 8128 1292
rect 8128 1236 8132 1292
rect 8068 1232 8132 1236
rect 10049 1295 10113 1299
rect 10049 1239 10053 1295
rect 10053 1239 10109 1295
rect 10109 1239 10113 1295
rect 10049 1235 10113 1239
rect 10278 1298 10342 1302
rect 10278 1242 10282 1298
rect 10282 1242 10338 1298
rect 10338 1242 10342 1298
rect 10278 1238 10342 1242
rect 10504 1303 10568 1307
rect 10504 1247 10508 1303
rect 10508 1247 10564 1303
rect 10564 1247 10568 1303
rect 10504 1243 10568 1247
rect 10732 1295 10796 1299
rect 10732 1239 10736 1295
rect 10736 1239 10792 1295
rect 10792 1239 10796 1295
rect 10732 1235 10796 1239
rect 10968 1301 11032 1305
rect 10968 1245 10972 1301
rect 10972 1245 11028 1301
rect 11028 1245 11032 1301
rect 10968 1241 11032 1245
rect 11160 1292 11224 1296
rect 11160 1236 11164 1292
rect 11164 1236 11220 1292
rect 11220 1236 11224 1292
rect 11160 1232 11224 1236
rect 12895 1292 12959 1296
rect 12895 1236 12899 1292
rect 12899 1236 12955 1292
rect 12955 1236 12959 1292
rect 12895 1232 12959 1236
rect 13099 1297 13163 1301
rect 13099 1241 13103 1297
rect 13103 1241 13159 1297
rect 13159 1241 13163 1297
rect 13099 1237 13163 1241
rect 13290 1292 13354 1296
rect 13290 1236 13294 1292
rect 13294 1236 13350 1292
rect 13350 1236 13354 1292
rect 13290 1232 13354 1236
rect 13492 1291 13556 1295
rect 13492 1235 13496 1291
rect 13496 1235 13552 1291
rect 13552 1235 13556 1291
rect 13492 1231 13556 1235
rect 13782 1292 13846 1296
rect 13782 1236 13786 1292
rect 13786 1236 13842 1292
rect 13842 1236 13846 1292
rect 13782 1232 13846 1236
rect 14067 1291 14131 1295
rect 14067 1235 14071 1291
rect 14071 1235 14127 1291
rect 14127 1235 14131 1291
rect 14067 1231 14131 1235
rect 15822 1296 15886 1300
rect 15822 1240 15826 1296
rect 15826 1240 15882 1296
rect 15882 1240 15886 1296
rect 15822 1236 15886 1240
rect 16016 1300 16080 1304
rect 16016 1244 16020 1300
rect 16020 1244 16076 1300
rect 16076 1244 16080 1300
rect 16016 1240 16080 1244
rect 16205 1297 16269 1301
rect 16205 1241 16209 1297
rect 16209 1241 16265 1297
rect 16265 1241 16269 1297
rect 16205 1237 16269 1241
rect 16428 1299 16492 1303
rect 16428 1243 16432 1299
rect 16432 1243 16488 1299
rect 16488 1243 16492 1299
rect 16428 1239 16492 1243
rect 259 1151 323 1155
rect 259 1095 263 1151
rect 263 1095 319 1151
rect 319 1095 323 1151
rect 259 1091 323 1095
rect 461 1147 525 1151
rect 461 1091 465 1147
rect 465 1091 521 1147
rect 521 1091 525 1147
rect 461 1087 525 1091
rect 650 1144 714 1148
rect 650 1088 654 1144
rect 654 1088 710 1144
rect 710 1088 714 1144
rect 650 1084 714 1088
rect 879 1145 943 1149
rect 879 1089 883 1145
rect 883 1089 939 1145
rect 939 1089 943 1145
rect 879 1085 943 1089
rect 2648 1148 2712 1152
rect 2648 1092 2652 1148
rect 2652 1092 2708 1148
rect 2708 1092 2712 1148
rect 2648 1088 2712 1092
rect 2863 1145 2927 1149
rect 2863 1089 2867 1145
rect 2867 1089 2923 1145
rect 2923 1089 2927 1145
rect 2863 1085 2927 1089
rect 3061 1142 3125 1146
rect 3061 1086 3065 1142
rect 3065 1086 3121 1142
rect 3121 1086 3125 1142
rect 3061 1082 3125 1086
rect 3256 1152 3320 1156
rect 3256 1096 3260 1152
rect 3260 1096 3316 1152
rect 3316 1096 3320 1152
rect 3256 1092 3320 1096
rect 3536 1150 3600 1154
rect 3536 1094 3540 1150
rect 3540 1094 3596 1150
rect 3596 1094 3600 1150
rect 3536 1090 3600 1094
rect 3755 1148 3819 1152
rect 3755 1092 3759 1148
rect 3759 1092 3815 1148
rect 3815 1092 3819 1148
rect 3755 1088 3819 1092
rect 5576 1145 5640 1149
rect 5576 1089 5580 1145
rect 5580 1089 5636 1145
rect 5636 1089 5640 1145
rect 5576 1085 5640 1089
rect 5927 1142 5991 1146
rect 5927 1086 5931 1142
rect 5931 1086 5987 1142
rect 5987 1086 5991 1142
rect 5927 1082 5991 1086
rect 6116 1140 6180 1144
rect 6116 1084 6120 1140
rect 6120 1084 6176 1140
rect 6176 1084 6180 1140
rect 6116 1080 6180 1084
rect 6321 1147 6385 1151
rect 6321 1091 6325 1147
rect 6325 1091 6381 1147
rect 6381 1091 6385 1147
rect 6321 1087 6385 1091
rect 6512 1149 6576 1153
rect 6512 1093 6516 1149
rect 6516 1093 6572 1149
rect 6572 1093 6576 1149
rect 6512 1089 6576 1093
rect 8557 1151 8621 1155
rect 8557 1095 8561 1151
rect 8561 1095 8617 1151
rect 8617 1095 8621 1151
rect 8557 1091 8621 1095
rect 8747 1153 8811 1157
rect 8747 1097 8751 1153
rect 8751 1097 8807 1153
rect 8807 1097 8811 1153
rect 8747 1093 8811 1097
rect 8941 1151 9005 1155
rect 8941 1095 8945 1151
rect 8945 1095 9001 1151
rect 9001 1095 9005 1151
rect 8941 1091 9005 1095
rect 9252 1147 9316 1151
rect 9252 1091 9256 1147
rect 9256 1091 9312 1147
rect 9312 1091 9316 1147
rect 9252 1087 9316 1091
rect 11435 1146 11499 1150
rect 11435 1090 11439 1146
rect 11439 1090 11495 1146
rect 11495 1090 11499 1146
rect 11435 1086 11499 1090
rect 11639 1146 11703 1150
rect 11639 1090 11643 1146
rect 11643 1090 11699 1146
rect 11699 1090 11703 1146
rect 11639 1086 11703 1090
rect 12204 1142 12268 1146
rect 12204 1086 12208 1142
rect 12208 1086 12264 1142
rect 12264 1086 12268 1142
rect 12204 1082 12268 1086
rect 12443 1144 12507 1148
rect 12443 1088 12447 1144
rect 12447 1088 12503 1144
rect 12503 1088 12507 1144
rect 12443 1084 12507 1088
rect 12647 1144 12711 1148
rect 12647 1088 12651 1144
rect 12651 1088 12707 1144
rect 12707 1088 12711 1144
rect 12647 1084 12711 1088
rect 14607 1152 14671 1156
rect 14607 1096 14611 1152
rect 14611 1096 14667 1152
rect 14667 1096 14671 1152
rect 14607 1092 14671 1096
rect 14840 1150 14904 1154
rect 14840 1094 14844 1150
rect 14844 1094 14900 1150
rect 14900 1094 14904 1150
rect 14840 1090 14904 1094
rect 15047 1148 15111 1152
rect 15047 1092 15051 1148
rect 15051 1092 15107 1148
rect 15107 1092 15111 1148
rect 15047 1088 15111 1092
rect 15256 1150 15320 1154
rect 15256 1094 15260 1150
rect 15260 1094 15316 1150
rect 15316 1094 15320 1150
rect 15256 1090 15320 1094
rect 15536 1152 15600 1156
rect 15536 1096 15540 1152
rect 15540 1096 15596 1152
rect 15596 1096 15600 1152
rect 15536 1092 15600 1096
rect 1186 602 1250 606
rect 1186 546 1190 602
rect 1190 546 1246 602
rect 1246 546 1250 602
rect 1186 542 1250 546
rect 1415 614 1479 618
rect 1415 558 1419 614
rect 1419 558 1475 614
rect 1475 558 1479 614
rect 1415 554 1479 558
rect 1634 604 1698 608
rect 1634 548 1638 604
rect 1638 548 1694 604
rect 1694 548 1698 604
rect 1634 544 1698 548
rect 1826 608 1890 612
rect 1826 552 1830 608
rect 1830 552 1886 608
rect 1886 552 1890 608
rect 1826 548 1890 552
rect 2320 606 2384 610
rect 2320 550 2324 606
rect 2324 550 2380 606
rect 2380 550 2384 606
rect 2320 546 2384 550
rect 4112 605 4176 609
rect 4112 549 4116 605
rect 4116 549 4172 605
rect 4172 549 4176 605
rect 4112 545 4176 549
rect 4505 603 4569 607
rect 4505 547 4509 603
rect 4509 547 4565 603
rect 4565 547 4569 603
rect 4505 543 4569 547
rect 4702 611 4766 615
rect 4702 555 4706 611
rect 4706 555 4762 611
rect 4762 555 4766 611
rect 4702 551 4766 555
rect 5032 613 5096 617
rect 5032 557 5036 613
rect 5036 557 5092 613
rect 5092 557 5096 613
rect 5032 553 5096 557
rect 5228 613 5292 617
rect 5228 557 5232 613
rect 5232 557 5288 613
rect 5288 557 5292 613
rect 5228 553 5292 557
rect 7135 606 7199 610
rect 7135 550 7139 606
rect 7139 550 7195 606
rect 7195 550 7199 606
rect 7135 546 7199 550
rect 7436 610 7500 614
rect 7436 554 7440 610
rect 7440 554 7496 610
rect 7496 554 7500 610
rect 7436 550 7500 554
rect 7642 611 7706 615
rect 7642 555 7646 611
rect 7646 555 7702 611
rect 7702 555 7706 611
rect 7642 551 7706 555
rect 7852 607 7916 611
rect 7852 551 7856 607
rect 7856 551 7912 607
rect 7912 551 7916 607
rect 7852 547 7916 551
rect 8063 613 8127 617
rect 8063 557 8067 613
rect 8067 557 8123 613
rect 8123 557 8127 613
rect 8063 553 8127 557
rect 9943 602 10007 606
rect 9943 546 9947 602
rect 9947 546 10003 602
rect 10003 546 10007 602
rect 9943 542 10007 546
rect 10200 609 10264 613
rect 10200 553 10204 609
rect 10204 553 10260 609
rect 10260 553 10264 609
rect 10200 549 10264 553
rect 10450 605 10514 609
rect 10450 549 10454 605
rect 10454 549 10510 605
rect 10510 549 10514 605
rect 10450 545 10514 549
rect 10721 610 10785 614
rect 10721 554 10725 610
rect 10725 554 10781 610
rect 10781 554 10785 610
rect 10721 550 10785 554
rect 10962 613 11026 617
rect 10962 557 10966 613
rect 10966 557 11022 613
rect 11022 557 11026 613
rect 10962 553 11026 557
rect 11187 609 11251 613
rect 11187 553 11191 609
rect 11191 553 11247 609
rect 11247 553 11251 609
rect 11187 549 11251 553
rect 12894 607 12958 611
rect 12894 551 12898 607
rect 12898 551 12954 607
rect 12954 551 12958 607
rect 12894 547 12958 551
rect 13095 608 13159 612
rect 13095 552 13099 608
rect 13099 552 13155 608
rect 13155 552 13159 608
rect 13095 548 13159 552
rect 13313 604 13377 608
rect 13313 548 13317 604
rect 13317 548 13373 604
rect 13373 548 13377 604
rect 13313 544 13377 548
rect 13520 608 13584 612
rect 13520 552 13524 608
rect 13524 552 13580 608
rect 13580 552 13584 608
rect 13520 548 13584 552
rect 13725 607 13789 611
rect 13725 551 13729 607
rect 13729 551 13785 607
rect 13785 551 13789 607
rect 13725 547 13789 551
rect 14072 603 14136 607
rect 14072 547 14076 603
rect 14076 547 14132 603
rect 14132 547 14136 603
rect 14072 543 14136 547
rect 15824 607 15888 611
rect 15824 551 15828 607
rect 15828 551 15884 607
rect 15884 551 15888 607
rect 15824 547 15888 551
rect 16015 610 16079 614
rect 16015 554 16019 610
rect 16019 554 16075 610
rect 16075 554 16079 610
rect 16015 550 16079 554
rect 16210 612 16274 616
rect 16210 556 16214 612
rect 16214 556 16270 612
rect 16270 556 16274 612
rect 16210 552 16274 556
rect 16657 607 16721 611
rect 16657 551 16661 607
rect 16661 551 16717 607
rect 16717 551 16721 607
rect 16657 547 16721 551
rect 41 458 105 462
rect 41 402 45 458
rect 45 402 101 458
rect 101 402 105 458
rect 41 398 105 402
rect 274 454 338 458
rect 274 398 278 454
rect 278 398 334 454
rect 334 398 338 454
rect 274 394 338 398
rect 489 461 553 465
rect 489 405 493 461
rect 493 405 549 461
rect 549 405 553 461
rect 489 401 553 405
rect 707 458 771 462
rect 707 402 711 458
rect 711 402 767 458
rect 767 402 771 458
rect 707 398 771 402
rect 923 459 987 463
rect 923 403 927 459
rect 927 403 983 459
rect 983 403 987 459
rect 923 399 987 403
rect 2644 455 2708 459
rect 2644 399 2648 455
rect 2648 399 2704 455
rect 2704 399 2708 455
rect 2644 395 2708 399
rect 2834 455 2898 459
rect 2834 399 2838 455
rect 2838 399 2894 455
rect 2894 399 2898 455
rect 2834 395 2898 399
rect 3044 458 3108 462
rect 3044 402 3048 458
rect 3048 402 3104 458
rect 3104 402 3108 458
rect 3044 398 3108 402
rect 3261 455 3325 459
rect 3261 399 3265 455
rect 3265 399 3321 455
rect 3321 399 3325 455
rect 3261 395 3325 399
rect 3556 458 3620 462
rect 3556 402 3560 458
rect 3560 402 3616 458
rect 3616 402 3620 458
rect 3556 398 3620 402
rect 3780 463 3844 467
rect 3780 407 3784 463
rect 3784 407 3840 463
rect 3840 407 3844 463
rect 3780 403 3844 407
rect 5658 456 5722 460
rect 5658 400 5662 456
rect 5662 400 5718 456
rect 5718 400 5722 456
rect 5658 396 5722 400
rect 5958 454 6022 458
rect 5958 398 5962 454
rect 5962 398 6018 454
rect 6018 398 6022 454
rect 5958 394 6022 398
rect 6210 458 6274 462
rect 6210 402 6214 458
rect 6214 402 6270 458
rect 6270 402 6274 458
rect 6210 398 6274 402
rect 6427 463 6491 467
rect 6427 407 6431 463
rect 6431 407 6487 463
rect 6487 407 6491 463
rect 6427 403 6491 407
rect 6628 460 6692 464
rect 6628 404 6632 460
rect 6632 404 6688 460
rect 6688 404 6692 460
rect 6628 400 6692 404
rect 8513 451 8577 455
rect 8513 395 8517 451
rect 8517 395 8573 451
rect 8573 395 8577 451
rect 8513 391 8577 395
rect 8705 451 8769 455
rect 8705 395 8709 451
rect 8709 395 8765 451
rect 8765 395 8769 451
rect 8705 391 8769 395
rect 8905 451 8969 455
rect 8905 395 8909 451
rect 8909 395 8965 451
rect 8965 395 8969 451
rect 8905 391 8969 395
rect 9523 459 9587 463
rect 9523 403 9527 459
rect 9527 403 9583 459
rect 9583 403 9587 459
rect 9523 399 9587 403
rect 11424 455 11488 459
rect 11424 399 11428 455
rect 11428 399 11484 455
rect 11484 399 11488 455
rect 11424 395 11488 399
rect 11680 455 11744 459
rect 11680 399 11684 455
rect 11684 399 11740 455
rect 11740 399 11744 455
rect 11680 395 11744 399
rect 11915 455 11979 459
rect 11915 399 11919 455
rect 11919 399 11975 455
rect 11975 399 11979 455
rect 11915 395 11979 399
rect 12204 457 12268 461
rect 12204 401 12208 457
rect 12208 401 12264 457
rect 12264 401 12268 457
rect 12204 397 12268 401
rect 12394 455 12458 459
rect 12394 399 12398 455
rect 12398 399 12454 455
rect 12454 399 12458 455
rect 12394 395 12458 399
rect 12598 457 12662 461
rect 12598 401 12602 457
rect 12602 401 12658 457
rect 12658 401 12662 457
rect 12598 397 12662 401
rect 14384 463 14448 467
rect 14384 407 14388 463
rect 14388 407 14444 463
rect 14444 407 14448 463
rect 14384 403 14448 407
rect 14626 459 14690 463
rect 14626 403 14630 459
rect 14630 403 14686 459
rect 14686 403 14690 459
rect 14626 399 14690 403
rect 14826 458 14890 462
rect 14826 402 14830 458
rect 14830 402 14886 458
rect 14886 402 14890 458
rect 14826 398 14890 402
rect 15016 466 15080 470
rect 15016 410 15020 466
rect 15020 410 15076 466
rect 15076 410 15080 466
rect 15016 406 15080 410
rect 15237 464 15301 468
rect 15237 408 15241 464
rect 15241 408 15297 464
rect 15297 408 15301 464
rect 15237 404 15301 408
rect 15533 459 15597 463
rect 15533 403 15537 459
rect 15537 403 15593 459
rect 15593 403 15597 459
rect 15533 399 15597 403
rect 415 -74 479 -70
rect 415 -130 419 -74
rect 419 -130 475 -74
rect 475 -130 479 -74
rect 415 -134 479 -130
rect 614 -77 678 -73
rect 614 -133 618 -77
rect 618 -133 674 -77
rect 674 -133 678 -77
rect 614 -137 678 -133
rect 825 -77 889 -73
rect 825 -133 829 -77
rect 829 -133 885 -77
rect 885 -133 889 -77
rect 825 -137 889 -133
rect 1031 -77 1095 -73
rect 1031 -133 1035 -77
rect 1035 -133 1091 -77
rect 1091 -133 1095 -77
rect 1031 -137 1095 -133
rect 1259 -79 1323 -75
rect 1259 -135 1263 -79
rect 1263 -135 1319 -79
rect 1319 -135 1323 -79
rect 1259 -139 1323 -135
rect 1503 -79 1567 -75
rect 1503 -135 1507 -79
rect 1507 -135 1563 -79
rect 1563 -135 1567 -79
rect 1503 -139 1567 -135
rect 1733 -77 1797 -73
rect 1733 -133 1737 -77
rect 1737 -133 1793 -77
rect 1793 -133 1797 -77
rect 1733 -137 1797 -133
rect 1939 -77 2003 -73
rect 1939 -133 1943 -77
rect 1943 -133 1999 -77
rect 1999 -133 2003 -77
rect 1939 -137 2003 -133
rect 2157 -72 2221 -68
rect 2157 -128 2161 -72
rect 2161 -128 2217 -72
rect 2217 -128 2221 -72
rect 2157 -132 2221 -128
rect 2360 -78 2424 -74
rect 2360 -134 2364 -78
rect 2364 -134 2420 -78
rect 2420 -134 2424 -78
rect 2360 -138 2424 -134
rect 2568 -75 2632 -71
rect 2568 -131 2572 -75
rect 2572 -131 2628 -75
rect 2628 -131 2632 -75
rect 2568 -135 2632 -131
rect 2831 -79 2895 -75
rect 2831 -135 2835 -79
rect 2835 -135 2891 -79
rect 2891 -135 2895 -79
rect 2831 -139 2895 -135
rect 3039 -78 3103 -74
rect 3039 -134 3043 -78
rect 3043 -134 3099 -78
rect 3099 -134 3103 -78
rect 3039 -138 3103 -134
rect 3249 -81 3313 -77
rect 3249 -137 3253 -81
rect 3253 -137 3309 -81
rect 3309 -137 3313 -81
rect 3249 -141 3313 -137
rect 3449 -75 3513 -71
rect 3449 -131 3453 -75
rect 3453 -131 3509 -75
rect 3509 -131 3513 -75
rect 3449 -135 3513 -131
rect 3652 -78 3716 -74
rect 3652 -134 3656 -78
rect 3656 -134 3712 -78
rect 3712 -134 3716 -78
rect 3652 -138 3716 -134
rect 3862 -78 3926 -74
rect 3862 -134 3866 -78
rect 3866 -134 3922 -78
rect 3922 -134 3926 -78
rect 3862 -138 3926 -134
rect 4063 -77 4127 -73
rect 4063 -133 4067 -77
rect 4067 -133 4123 -77
rect 4123 -133 4127 -77
rect 4063 -137 4127 -133
rect 4279 -76 4343 -72
rect 4279 -132 4283 -76
rect 4283 -132 4339 -76
rect 4339 -132 4343 -76
rect 4279 -136 4343 -132
rect 4560 -78 4624 -74
rect 4560 -134 4564 -78
rect 4564 -134 4620 -78
rect 4620 -134 4624 -78
rect 4560 -138 4624 -134
rect 4780 -83 4844 -79
rect 4780 -139 4784 -83
rect 4784 -139 4840 -83
rect 4840 -139 4844 -83
rect 4780 -143 4844 -139
rect 4985 -82 5049 -78
rect 4985 -138 4989 -82
rect 4989 -138 5045 -82
rect 5045 -138 5049 -82
rect 4985 -142 5049 -138
rect 5206 -76 5270 -72
rect 5206 -132 5210 -76
rect 5210 -132 5266 -76
rect 5266 -132 5270 -76
rect 5206 -136 5270 -132
rect 5411 -83 5475 -79
rect 5411 -139 5415 -83
rect 5415 -139 5471 -83
rect 5471 -139 5475 -83
rect 5411 -143 5475 -139
rect 5620 -82 5684 -78
rect 5620 -138 5624 -82
rect 5624 -138 5680 -82
rect 5680 -138 5684 -82
rect 5620 -142 5684 -138
rect 5837 -82 5901 -78
rect 5837 -138 5841 -82
rect 5841 -138 5897 -82
rect 5897 -138 5901 -82
rect 5837 -142 5901 -138
rect 6051 -77 6115 -73
rect 6051 -133 6055 -77
rect 6055 -133 6111 -77
rect 6111 -133 6115 -77
rect 6051 -137 6115 -133
rect 6246 -79 6310 -75
rect 6246 -135 6250 -79
rect 6250 -135 6306 -79
rect 6306 -135 6310 -79
rect 6246 -139 6310 -135
rect 6441 -82 6505 -78
rect 6441 -138 6445 -82
rect 6445 -138 6501 -82
rect 6501 -138 6505 -82
rect 6441 -142 6505 -138
rect 6643 -79 6707 -75
rect 6643 -135 6647 -79
rect 6647 -135 6703 -79
rect 6703 -135 6707 -79
rect 6643 -139 6707 -135
rect 6927 -78 6991 -74
rect 6927 -134 6931 -78
rect 6931 -134 6987 -78
rect 6987 -134 6991 -78
rect 6927 -138 6991 -134
rect 7126 -77 7190 -73
rect 7126 -133 7130 -77
rect 7130 -133 7186 -77
rect 7186 -133 7190 -77
rect 7126 -137 7190 -133
rect 7329 -75 7393 -71
rect 7329 -131 7333 -75
rect 7333 -131 7389 -75
rect 7389 -131 7393 -75
rect 7329 -135 7393 -131
rect 7594 -78 7658 -74
rect 7594 -134 7598 -78
rect 7598 -134 7654 -78
rect 7654 -134 7658 -78
rect 7594 -138 7658 -134
rect 7792 -79 7856 -75
rect 7792 -135 7796 -79
rect 7796 -135 7852 -79
rect 7852 -135 7856 -79
rect 7792 -139 7856 -135
rect 7981 -77 8045 -73
rect 7981 -133 7985 -77
rect 7985 -133 8041 -77
rect 8041 -133 8045 -77
rect 7981 -137 8045 -133
rect 8193 -77 8257 -73
rect 8193 -133 8197 -77
rect 8197 -133 8253 -77
rect 8253 -133 8257 -77
rect 8193 -137 8257 -133
rect 8410 -77 8474 -73
rect 8410 -133 8414 -77
rect 8414 -133 8470 -77
rect 8470 -133 8474 -77
rect 8410 -137 8474 -133
rect 8615 -81 8679 -77
rect 8615 -137 8619 -81
rect 8619 -137 8675 -81
rect 8675 -137 8679 -81
rect 8615 -141 8679 -137
rect 8820 -81 8884 -77
rect 8820 -137 8824 -81
rect 8824 -137 8880 -81
rect 8880 -137 8884 -81
rect 8820 -141 8884 -137
rect 9028 -76 9092 -72
rect 9028 -132 9032 -76
rect 9032 -132 9088 -76
rect 9088 -132 9092 -76
rect 9028 -136 9092 -132
rect 9311 -77 9375 -73
rect 9311 -133 9315 -77
rect 9315 -133 9371 -77
rect 9371 -133 9375 -77
rect 9311 -137 9375 -133
rect 9504 -79 9568 -75
rect 9504 -135 9508 -79
rect 9508 -135 9564 -79
rect 9564 -135 9568 -79
rect 9504 -139 9568 -135
rect 9730 -81 9794 -77
rect 9730 -137 9734 -81
rect 9734 -137 9790 -81
rect 9790 -137 9794 -81
rect 9730 -141 9794 -137
rect 9995 -81 10059 -77
rect 9995 -137 9999 -81
rect 9999 -137 10055 -81
rect 10055 -137 10059 -81
rect 9995 -141 10059 -137
rect 10189 -77 10253 -73
rect 10189 -133 10193 -77
rect 10193 -133 10249 -77
rect 10249 -133 10253 -77
rect 10189 -137 10253 -133
rect 10387 -86 10451 -82
rect 10387 -142 10391 -86
rect 10391 -142 10447 -86
rect 10447 -142 10451 -86
rect 10387 -146 10451 -142
rect 10591 -78 10655 -74
rect 10591 -134 10595 -78
rect 10595 -134 10651 -78
rect 10651 -134 10655 -78
rect 10591 -138 10655 -134
rect 10811 -75 10875 -71
rect 10811 -131 10815 -75
rect 10815 -131 10871 -75
rect 10871 -131 10875 -75
rect 10811 -135 10875 -131
rect 11026 -79 11090 -75
rect 11026 -135 11030 -79
rect 11030 -135 11086 -79
rect 11086 -135 11090 -79
rect 11026 -139 11090 -135
rect 11254 -76 11318 -72
rect 11254 -132 11258 -76
rect 11258 -132 11314 -76
rect 11314 -132 11318 -76
rect 11254 -136 11318 -132
rect 11458 -79 11522 -75
rect 11458 -135 11462 -79
rect 11462 -135 11518 -79
rect 11518 -135 11522 -79
rect 11458 -139 11522 -135
rect 11696 -77 11760 -73
rect 11696 -133 11700 -77
rect 11700 -133 11756 -77
rect 11756 -133 11760 -77
rect 11696 -137 11760 -133
rect 11889 -76 11953 -72
rect 11889 -132 11893 -76
rect 11893 -132 11949 -76
rect 11949 -132 11953 -76
rect 11889 -136 11953 -132
rect 12086 -81 12150 -77
rect 12086 -137 12090 -81
rect 12090 -137 12146 -81
rect 12146 -137 12150 -81
rect 12086 -141 12150 -137
rect 12342 -78 12406 -74
rect 12342 -134 12346 -78
rect 12346 -134 12402 -78
rect 12402 -134 12406 -78
rect 12342 -138 12406 -134
rect 12581 -82 12645 -78
rect 12581 -138 12585 -82
rect 12585 -138 12641 -82
rect 12641 -138 12645 -82
rect 12581 -142 12645 -138
rect 12814 -86 12878 -82
rect 12814 -142 12818 -86
rect 12818 -142 12874 -86
rect 12874 -142 12878 -86
rect 12814 -146 12878 -142
rect 13035 -81 13099 -77
rect 13035 -137 13039 -81
rect 13039 -137 13095 -81
rect 13095 -137 13099 -81
rect 13035 -141 13099 -137
rect 13226 -81 13290 -77
rect 13226 -137 13230 -81
rect 13230 -137 13286 -81
rect 13286 -137 13290 -81
rect 13226 -141 13290 -137
rect 13454 -79 13518 -75
rect 13454 -135 13458 -79
rect 13458 -135 13514 -79
rect 13514 -135 13518 -79
rect 13454 -139 13518 -135
rect 13651 -84 13715 -80
rect 13651 -140 13655 -84
rect 13655 -140 13711 -84
rect 13711 -140 13715 -84
rect 13651 -144 13715 -140
rect 13863 -84 13927 -80
rect 13863 -140 13867 -84
rect 13867 -140 13923 -84
rect 13923 -140 13927 -84
rect 13863 -144 13927 -140
rect 14090 -81 14154 -77
rect 14090 -137 14094 -81
rect 14094 -137 14150 -81
rect 14150 -137 14154 -81
rect 14090 -141 14154 -137
rect 14279 -80 14343 -76
rect 14279 -136 14283 -80
rect 14283 -136 14339 -80
rect 14339 -136 14343 -80
rect 14279 -140 14343 -136
rect 14505 -79 14569 -75
rect 14505 -135 14509 -79
rect 14509 -135 14565 -79
rect 14565 -135 14569 -79
rect 14505 -139 14569 -135
rect 14759 -79 14823 -75
rect 14759 -135 14763 -79
rect 14763 -135 14819 -79
rect 14819 -135 14823 -79
rect 14759 -139 14823 -135
rect 15003 -82 15067 -78
rect 15003 -138 15007 -82
rect 15007 -138 15063 -82
rect 15063 -138 15067 -82
rect 15003 -142 15067 -138
rect 15233 -83 15297 -79
rect 15233 -139 15237 -83
rect 15237 -139 15293 -83
rect 15293 -139 15297 -83
rect 15233 -143 15297 -139
rect 15491 -80 15555 -76
rect 15491 -136 15495 -80
rect 15495 -136 15551 -80
rect 15551 -136 15555 -80
rect 15491 -140 15555 -136
rect 15701 -80 15765 -76
rect 15701 -136 15705 -80
rect 15705 -136 15761 -80
rect 15761 -136 15765 -80
rect 15701 -140 15765 -136
rect 15926 -80 15990 -76
rect 15926 -136 15930 -80
rect 15930 -136 15986 -80
rect 15986 -136 15990 -80
rect 15926 -140 15990 -136
rect 16145 -83 16209 -79
rect 16145 -139 16149 -83
rect 16149 -139 16205 -83
rect 16205 -139 16209 -83
rect 16145 -143 16209 -139
rect 16491 -79 16555 -75
rect 16491 -135 16495 -79
rect 16495 -135 16551 -79
rect 16551 -135 16555 -79
rect 16491 -139 16555 -135
rect 16690 -82 16754 -78
rect 16690 -138 16694 -82
rect 16694 -138 16750 -82
rect 16750 -138 16754 -82
rect 16690 -142 16754 -138
<< metal4 >>
rect -144 3018 7278 3041
rect -144 2986 15690 3018
rect -144 2984 1259 2986
rect -144 2982 249 2984
rect -144 2918 47 2982
rect 111 2920 249 2982
rect 313 2982 858 2984
rect 313 2920 460 2982
rect 111 2918 460 2920
rect 524 2918 650 2982
rect 714 2920 858 2982
rect 922 2920 1060 2984
rect 1124 2922 1259 2984
rect 1323 2985 2146 2986
rect 1323 2983 1655 2985
rect 1323 2922 1454 2983
rect 1124 2920 1454 2922
rect 714 2919 1454 2920
rect 1518 2921 1655 2983
rect 1719 2983 2146 2985
rect 1719 2921 1872 2983
rect 1518 2919 1872 2921
rect 1936 2922 2146 2983
rect 2210 2982 15690 2986
rect 2210 2979 2646 2982
rect 2210 2922 2423 2979
rect 1936 2919 2423 2922
rect 714 2918 2423 2919
rect -144 2915 2423 2918
rect 2487 2918 2646 2979
rect 2710 2981 15690 2982
rect 2710 2918 2878 2981
rect 2487 2917 2878 2918
rect 2942 2980 5897 2981
rect 2942 2979 5022 2980
rect 2942 2978 4822 2979
rect 2942 2917 4514 2978
rect 2487 2915 4514 2917
rect -144 2914 4514 2915
rect 4578 2915 4822 2978
rect 4886 2916 5022 2979
rect 5086 2979 5695 2980
rect 5086 2916 5241 2979
rect 4886 2915 5241 2916
rect 5305 2978 5695 2979
rect 5305 2915 5487 2978
rect 4578 2914 5487 2915
rect 5551 2916 5695 2978
rect 5759 2917 5897 2980
rect 5961 2980 15690 2981
rect 5961 2917 6090 2980
rect 5759 2916 6090 2917
rect 6154 2979 15690 2980
rect 6154 2916 6462 2979
rect 5551 2915 6462 2916
rect 6526 2977 7214 2979
rect 6526 2915 6651 2977
rect 5551 2914 6651 2915
rect -144 2913 6651 2914
rect 6715 2913 6941 2977
rect 7005 2915 7214 2977
rect 7278 2915 15690 2979
rect 7005 2913 15690 2915
rect -144 2721 15690 2913
rect -144 1838 1030 2721
rect -144 1774 13 1838
rect 77 1836 1030 1838
rect 77 1774 253 1836
rect -144 1772 253 1774
rect 317 1835 793 1836
rect 317 1772 575 1835
rect -144 1771 575 1772
rect 639 1772 793 1835
rect 857 1772 1030 1836
rect 639 1771 1030 1772
rect -144 1155 1030 1771
rect -144 1091 259 1155
rect 323 1151 1030 1155
rect 323 1091 461 1151
rect -144 1087 461 1091
rect 525 1149 1030 1151
rect 525 1148 879 1149
rect 525 1087 650 1148
rect -144 1084 650 1087
rect 714 1085 879 1148
rect 943 1085 1030 1149
rect 714 1084 1030 1085
rect -144 465 1030 1084
rect -144 462 489 465
rect -144 398 41 462
rect 105 458 489 462
rect 105 398 274 458
rect -144 394 274 398
rect 338 401 489 458
rect 553 463 1030 465
rect 553 462 923 463
rect 553 401 707 462
rect 338 398 707 401
rect 771 399 923 462
rect 987 399 1030 463
rect 771 398 1030 399
rect 338 394 1030 398
rect -144 195 1030 394
rect 1110 2447 2496 2640
rect 1110 2443 1384 2447
rect 1110 2379 1165 2443
rect 1229 2383 1384 2443
rect 1448 2383 1667 2447
rect 1731 2383 1876 2447
rect 1940 2445 2496 2447
rect 1940 2383 2147 2445
rect 1229 2381 2147 2383
rect 2211 2381 2496 2445
rect 1229 2379 2496 2381
rect 1110 1300 2496 2379
rect 1110 1236 1204 1300
rect 1268 1236 1421 1300
rect 1485 1236 1640 1300
rect 1704 1296 2496 1300
rect 1704 1236 1853 1296
rect 1110 1232 1853 1236
rect 1917 1232 2064 1296
rect 2128 1232 2496 1296
rect 1110 618 2496 1232
rect 1110 606 1415 618
rect 1110 542 1186 606
rect 1250 554 1415 606
rect 1479 612 2496 618
rect 1479 608 1826 612
rect 1479 554 1634 608
rect 1250 544 1634 554
rect 1698 548 1826 608
rect 1890 610 2496 612
rect 1890 548 2320 610
rect 1698 546 2320 548
rect 2384 546 2496 610
rect 1698 544 2496 546
rect 1250 542 2496 544
rect 1110 114 2496 542
rect 2576 1842 3962 2721
rect 2576 1840 3022 1842
rect 2576 1776 2697 1840
rect 2761 1778 3022 1840
rect 3086 1778 3290 1842
rect 3354 1778 3556 1842
rect 3620 1840 3962 1842
rect 3620 1778 3796 1840
rect 2761 1776 3796 1778
rect 3860 1776 3962 1840
rect 2576 1156 3962 1776
rect 2576 1152 3256 1156
rect 2576 1088 2648 1152
rect 2712 1149 3256 1152
rect 2712 1088 2863 1149
rect 2576 1085 2863 1088
rect 2927 1146 3256 1149
rect 2927 1085 3061 1146
rect 2576 1082 3061 1085
rect 3125 1092 3256 1146
rect 3320 1154 3962 1156
rect 3320 1092 3536 1154
rect 3125 1090 3536 1092
rect 3600 1152 3962 1154
rect 3600 1090 3755 1152
rect 3125 1088 3755 1090
rect 3819 1088 3962 1152
rect 3125 1082 3962 1088
rect 2576 467 3962 1082
rect 2576 462 3780 467
rect 2576 459 3044 462
rect 2576 395 2644 459
rect 2708 395 2834 459
rect 2898 398 3044 459
rect 3108 459 3556 462
rect 3108 398 3261 459
rect 2898 395 3261 398
rect 3325 398 3556 459
rect 3620 403 3780 462
rect 3844 403 3962 467
rect 3620 398 3962 403
rect 3325 395 3962 398
rect 2576 195 3962 395
rect 4042 2446 5428 2640
rect 4042 2443 4471 2446
rect 4042 2379 4222 2443
rect 4286 2382 4471 2443
rect 4535 2438 5428 2446
rect 4535 2432 5069 2438
rect 4535 2382 4815 2432
rect 4286 2379 4815 2382
rect 4042 2368 4815 2379
rect 4879 2374 5069 2432
rect 5133 2374 5298 2438
rect 5362 2374 5428 2438
rect 4879 2368 5428 2374
rect 4042 1300 5428 2368
rect 4042 1296 5038 1300
rect 4042 1232 4188 1296
rect 4252 1295 5038 1296
rect 4252 1232 4466 1295
rect 4042 1231 4466 1232
rect 4530 1236 5038 1295
rect 5102 1236 5277 1300
rect 5341 1236 5428 1300
rect 4530 1231 5428 1236
rect 4042 617 5428 1231
rect 4042 615 5032 617
rect 4042 609 4702 615
rect 4042 545 4112 609
rect 4176 607 4702 609
rect 4176 545 4505 607
rect 4042 543 4505 545
rect 4569 551 4702 607
rect 4766 553 5032 615
rect 5096 553 5228 617
rect 5292 553 5428 617
rect 4766 551 5428 553
rect 4569 543 5428 551
rect 4042 114 5428 543
rect 5508 1846 6894 2721
rect 5508 1843 5956 1846
rect 5508 1779 5590 1843
rect 5654 1782 5956 1843
rect 6020 1782 6200 1846
rect 6264 1837 6894 1846
rect 6264 1782 6623 1837
rect 5654 1779 6623 1782
rect 5508 1773 6623 1779
rect 6687 1773 6894 1837
rect 5508 1153 6894 1773
rect 5508 1151 6512 1153
rect 5508 1149 6321 1151
rect 5508 1085 5576 1149
rect 5640 1146 6321 1149
rect 5640 1085 5927 1146
rect 5508 1082 5927 1085
rect 5991 1144 6321 1146
rect 5991 1082 6116 1144
rect 5508 1080 6116 1082
rect 6180 1087 6321 1144
rect 6385 1089 6512 1151
rect 6576 1089 6894 1153
rect 6385 1087 6894 1089
rect 6180 1080 6894 1087
rect 5508 467 6894 1080
rect 5508 462 6427 467
rect 5508 460 6210 462
rect 5508 396 5658 460
rect 5722 458 6210 460
rect 5722 396 5958 458
rect 5508 394 5958 396
rect 6022 398 6210 458
rect 6274 403 6427 462
rect 6491 464 6894 467
rect 6491 403 6628 464
rect 6274 400 6628 403
rect 6692 400 6894 464
rect 6274 398 6894 400
rect 6022 394 6894 398
rect 5508 194 6894 394
rect 6974 2445 8360 2640
rect 6974 2443 7220 2445
rect 6974 2379 7016 2443
rect 7080 2381 7220 2443
rect 7284 2443 8360 2445
rect 7284 2381 7543 2443
rect 7080 2379 7543 2381
rect 7607 2379 8360 2443
rect 6974 1305 8360 2379
rect 6974 1303 7852 1305
rect 6974 1298 7662 1303
rect 6974 1234 7435 1298
rect 7499 1239 7662 1298
rect 7726 1241 7852 1303
rect 7916 1296 8360 1305
rect 7916 1241 8068 1296
rect 7726 1239 8068 1241
rect 7499 1234 8068 1239
rect 6974 1232 8068 1234
rect 8132 1232 8360 1296
rect 6974 617 8360 1232
rect 6974 615 8063 617
rect 6974 614 7642 615
rect 6974 610 7436 614
rect 6974 546 7135 610
rect 7199 550 7436 610
rect 7500 551 7642 614
rect 7706 611 8063 615
rect 7706 551 7852 611
rect 7500 550 7852 551
rect 7199 547 7852 550
rect 7916 553 8063 611
rect 8127 553 8360 617
rect 7916 547 8360 553
rect 7199 546 8360 547
rect 6974 114 8360 546
rect 8440 1844 9826 2721
rect 8440 1839 9024 1844
rect 8440 1775 8566 1839
rect 8630 1836 9024 1839
rect 8630 1775 8818 1836
rect 8440 1772 8818 1775
rect 8882 1780 9024 1836
rect 9088 1839 9826 1844
rect 9088 1838 9605 1839
rect 9088 1780 9307 1838
rect 8882 1774 9307 1780
rect 9371 1775 9605 1838
rect 9669 1775 9826 1839
rect 9371 1774 9826 1775
rect 8882 1772 9826 1774
rect 8440 1157 9826 1772
rect 8440 1155 8747 1157
rect 8440 1091 8557 1155
rect 8621 1093 8747 1155
rect 8811 1155 9826 1157
rect 8811 1093 8941 1155
rect 8621 1091 8941 1093
rect 9005 1151 9826 1155
rect 9005 1091 9252 1151
rect 8440 1087 9252 1091
rect 9316 1087 9826 1151
rect 8440 463 9826 1087
rect 8440 455 9523 463
rect 8440 391 8513 455
rect 8577 391 8705 455
rect 8769 391 8905 455
rect 8969 399 9523 455
rect 9587 399 9826 463
rect 8969 391 9826 399
rect 8440 195 9826 391
rect 9906 1307 11292 2641
rect 9906 1302 10504 1307
rect 9906 1299 10278 1302
rect 9906 1235 10049 1299
rect 10113 1238 10278 1299
rect 10342 1243 10504 1302
rect 10568 1305 11292 1307
rect 10568 1299 10968 1305
rect 10568 1243 10732 1299
rect 10342 1238 10732 1243
rect 10113 1235 10732 1238
rect 10796 1241 10968 1299
rect 11032 1296 11292 1305
rect 11032 1241 11160 1296
rect 10796 1235 11160 1241
rect 9906 1232 11160 1235
rect 11224 1232 11292 1296
rect 9906 617 11292 1232
rect 9906 614 10962 617
rect 9906 613 10721 614
rect 9906 606 10200 613
rect 9906 542 9943 606
rect 10007 549 10200 606
rect 10264 609 10721 613
rect 10264 549 10450 609
rect 10007 545 10450 549
rect 10514 550 10721 609
rect 10785 553 10962 614
rect 11026 613 11292 617
rect 11026 553 11187 613
rect 10785 550 11187 553
rect 10514 549 11187 550
rect 11251 549 11292 613
rect 10514 545 11292 549
rect 10007 542 11292 545
rect 9906 114 11292 542
rect 11372 1842 12758 2721
rect 11372 1840 11647 1842
rect 11372 1776 11437 1840
rect 11501 1778 11647 1840
rect 11711 1840 12758 1842
rect 11711 1778 11998 1840
rect 11501 1776 11998 1778
rect 12062 1776 12278 1840
rect 12342 1839 12758 1840
rect 12342 1776 12595 1839
rect 11372 1775 12595 1776
rect 12659 1775 12758 1839
rect 11372 1150 12758 1775
rect 11372 1086 11435 1150
rect 11499 1086 11639 1150
rect 11703 1148 12758 1150
rect 11703 1146 12443 1148
rect 11703 1086 12204 1146
rect 11372 1082 12204 1086
rect 12268 1084 12443 1146
rect 12507 1084 12647 1148
rect 12711 1084 12758 1148
rect 12268 1082 12758 1084
rect 11372 461 12758 1082
rect 11372 459 12204 461
rect 11372 395 11424 459
rect 11488 395 11680 459
rect 11744 395 11915 459
rect 11979 397 12204 459
rect 12268 459 12598 461
rect 12268 397 12394 459
rect 11979 395 12394 397
rect 12458 397 12598 459
rect 12662 397 12758 461
rect 12458 395 12758 397
rect 11372 195 12758 395
rect 12838 1301 14224 2640
rect 12838 1296 13099 1301
rect 12838 1232 12895 1296
rect 12959 1237 13099 1296
rect 13163 1296 14224 1301
rect 13163 1237 13290 1296
rect 12959 1232 13290 1237
rect 13354 1295 13782 1296
rect 13354 1232 13492 1295
rect 12838 1231 13492 1232
rect 13556 1232 13782 1295
rect 13846 1295 14224 1296
rect 13846 1232 14067 1295
rect 13556 1231 14067 1232
rect 14131 1231 14224 1295
rect 12838 612 14224 1231
rect 12838 611 13095 612
rect 12838 547 12894 611
rect 12958 548 13095 611
rect 13159 608 13520 612
rect 13159 548 13313 608
rect 12958 547 13313 548
rect 12838 544 13313 547
rect 13377 548 13520 608
rect 13584 611 14224 612
rect 13584 548 13725 611
rect 13377 547 13725 548
rect 13789 607 14224 611
rect 13789 547 14072 607
rect 13377 544 14072 547
rect 12838 543 14072 544
rect 14136 543 14224 607
rect 12838 114 14224 543
rect 14304 1840 15690 2721
rect 14304 1837 15541 1840
rect 14304 1773 14385 1837
rect 14449 1773 14680 1837
rect 14744 1773 14967 1837
rect 15031 1773 15257 1837
rect 15321 1776 15541 1837
rect 15605 1776 15690 1840
rect 15321 1773 15690 1776
rect 14304 1156 15690 1773
rect 14304 1092 14607 1156
rect 14671 1154 15536 1156
rect 14671 1092 14840 1154
rect 14304 1090 14840 1092
rect 14904 1152 15256 1154
rect 14904 1090 15047 1152
rect 14304 1088 15047 1090
rect 15111 1090 15256 1152
rect 15320 1092 15536 1154
rect 15600 1092 15690 1156
rect 15320 1090 15690 1092
rect 15111 1088 15690 1090
rect 14304 470 15690 1088
rect 14304 467 15016 470
rect 14304 403 14384 467
rect 14448 463 15016 467
rect 14448 403 14626 463
rect 14304 399 14626 403
rect 14690 462 15016 463
rect 14690 399 14826 462
rect 14304 398 14826 399
rect 14890 406 15016 462
rect 15080 468 15690 470
rect 15080 406 15237 468
rect 14890 404 15237 406
rect 15301 463 15690 468
rect 15301 404 15533 463
rect 14890 399 15533 404
rect 15597 399 15690 463
rect 14890 398 15690 399
rect 14304 195 15690 398
rect 15770 1304 16876 2640
rect 15770 1300 16016 1304
rect 15770 1236 15822 1300
rect 15886 1240 16016 1300
rect 16080 1303 16876 1304
rect 16080 1301 16428 1303
rect 16080 1240 16205 1301
rect 15886 1237 16205 1240
rect 16269 1239 16428 1301
rect 16492 1239 16876 1303
rect 16269 1237 16876 1239
rect 15886 1236 16876 1237
rect 15770 616 16876 1236
rect 15770 614 16210 616
rect 15770 611 16015 614
rect 15770 547 15824 611
rect 15888 550 16015 611
rect 16079 552 16210 614
rect 16274 611 16876 616
rect 16274 552 16657 611
rect 16079 550 16657 552
rect 15888 547 16657 550
rect 16721 547 16876 611
rect 15770 114 16876 547
rect 196 -68 16876 114
rect 196 -70 2157 -68
rect 196 -134 415 -70
rect 479 -73 2157 -70
rect 479 -134 614 -73
rect 196 -137 614 -134
rect 678 -137 825 -73
rect 889 -137 1031 -73
rect 1095 -75 1733 -73
rect 1095 -137 1259 -75
rect 196 -139 1259 -137
rect 1323 -139 1503 -75
rect 1567 -137 1733 -75
rect 1797 -137 1939 -73
rect 2003 -132 2157 -73
rect 2221 -71 16876 -68
rect 2221 -74 2568 -71
rect 2221 -132 2360 -74
rect 2003 -137 2360 -132
rect 1567 -138 2360 -137
rect 2424 -135 2568 -74
rect 2632 -74 3449 -71
rect 2632 -75 3039 -74
rect 2632 -135 2831 -75
rect 2424 -138 2831 -135
rect 1567 -139 2831 -138
rect 2895 -138 3039 -75
rect 3103 -77 3449 -74
rect 3103 -138 3249 -77
rect 2895 -139 3249 -138
rect 196 -141 3249 -139
rect 3313 -135 3449 -77
rect 3513 -72 7329 -71
rect 3513 -73 4279 -72
rect 3513 -74 4063 -73
rect 3513 -135 3652 -74
rect 3313 -138 3652 -135
rect 3716 -138 3862 -74
rect 3926 -137 4063 -74
rect 4127 -136 4279 -73
rect 4343 -74 5206 -72
rect 4343 -136 4560 -74
rect 4127 -137 4560 -136
rect 3926 -138 4560 -137
rect 4624 -78 5206 -74
rect 4624 -79 4985 -78
rect 4624 -138 4780 -79
rect 3313 -141 4780 -138
rect 196 -143 4780 -141
rect 4844 -142 4985 -79
rect 5049 -136 5206 -78
rect 5270 -73 7329 -72
rect 5270 -78 6051 -73
rect 5270 -79 5620 -78
rect 5270 -136 5411 -79
rect 5049 -142 5411 -136
rect 4844 -143 5411 -142
rect 5475 -142 5620 -79
rect 5684 -142 5837 -78
rect 5901 -137 6051 -78
rect 6115 -74 7126 -73
rect 6115 -75 6927 -74
rect 6115 -137 6246 -75
rect 5901 -139 6246 -137
rect 6310 -78 6643 -75
rect 6310 -139 6441 -78
rect 5901 -142 6441 -139
rect 6505 -139 6643 -78
rect 6707 -138 6927 -75
rect 6991 -137 7126 -74
rect 7190 -135 7329 -73
rect 7393 -72 10811 -71
rect 7393 -73 9028 -72
rect 7393 -74 7981 -73
rect 7393 -135 7594 -74
rect 7190 -137 7594 -135
rect 6991 -138 7594 -137
rect 7658 -75 7981 -74
rect 7658 -138 7792 -75
rect 6707 -139 7792 -138
rect 7856 -137 7981 -75
rect 8045 -137 8193 -73
rect 8257 -137 8410 -73
rect 8474 -77 9028 -73
rect 8474 -137 8615 -77
rect 7856 -139 8615 -137
rect 6505 -141 8615 -139
rect 8679 -141 8820 -77
rect 8884 -136 9028 -77
rect 9092 -73 10811 -72
rect 9092 -136 9311 -73
rect 8884 -137 9311 -136
rect 9375 -75 10189 -73
rect 9375 -137 9504 -75
rect 8884 -139 9504 -137
rect 9568 -77 10189 -75
rect 9568 -139 9730 -77
rect 8884 -141 9730 -139
rect 9794 -141 9995 -77
rect 10059 -137 10189 -77
rect 10253 -74 10811 -73
rect 10253 -82 10591 -74
rect 10253 -137 10387 -82
rect 10059 -141 10387 -137
rect 6505 -142 10387 -141
rect 5475 -143 10387 -142
rect 196 -146 10387 -143
rect 10451 -138 10591 -82
rect 10655 -135 10811 -74
rect 10875 -72 16876 -71
rect 10875 -75 11254 -72
rect 10875 -135 11026 -75
rect 10655 -138 11026 -135
rect 10451 -139 11026 -138
rect 11090 -136 11254 -75
rect 11318 -73 11889 -72
rect 11318 -75 11696 -73
rect 11318 -136 11458 -75
rect 11090 -139 11458 -136
rect 11522 -137 11696 -75
rect 11760 -136 11889 -73
rect 11953 -74 16876 -72
rect 11953 -77 12342 -74
rect 11953 -136 12086 -77
rect 11760 -137 12086 -136
rect 11522 -139 12086 -137
rect 10451 -141 12086 -139
rect 12150 -138 12342 -77
rect 12406 -75 16876 -74
rect 12406 -77 13454 -75
rect 12406 -78 13035 -77
rect 12406 -138 12581 -78
rect 12150 -141 12581 -138
rect 10451 -142 12581 -141
rect 12645 -82 13035 -78
rect 12645 -142 12814 -82
rect 10451 -146 12814 -142
rect 12878 -141 13035 -82
rect 13099 -141 13226 -77
rect 13290 -139 13454 -77
rect 13518 -76 14505 -75
rect 13518 -77 14279 -76
rect 13518 -80 14090 -77
rect 13518 -139 13651 -80
rect 13290 -141 13651 -139
rect 12878 -144 13651 -141
rect 13715 -144 13863 -80
rect 13927 -141 14090 -80
rect 14154 -140 14279 -77
rect 14343 -139 14505 -76
rect 14569 -139 14759 -75
rect 14823 -76 16491 -75
rect 14823 -78 15491 -76
rect 14823 -139 15003 -78
rect 14343 -140 15003 -139
rect 14154 -141 15003 -140
rect 13927 -142 15003 -141
rect 15067 -79 15491 -78
rect 15067 -142 15233 -79
rect 13927 -143 15233 -142
rect 15297 -140 15491 -79
rect 15555 -140 15701 -76
rect 15765 -140 15926 -76
rect 15990 -79 16491 -76
rect 15990 -140 16145 -79
rect 15297 -143 16145 -140
rect 16209 -139 16491 -79
rect 16555 -78 16876 -75
rect 16555 -139 16690 -78
rect 16209 -142 16690 -139
rect 16754 -142 16876 -78
rect 16209 -143 16876 -142
rect 13927 -144 16876 -143
rect 12878 -146 16876 -144
rect 196 -206 16876 -146
<< labels >>
flabel metal2 9709 344 9751 3300 0 FreeSans 320 0 0 0 VSS_SW[3]
port 6 nsew
flabel metal2 7317 345 7359 3300 0 FreeSans 320 0 0 0 VSS_SW[4]
port 7 nsew
flabel metal2 4926 345 4968 3300 0 FreeSans 320 0 0 0 VSS_SW[5]
port 8 nsew
flabel metal2 14290 1062 14332 3300 0 FreeSans 320 0 0 0 VDD_SW[2]
port 11 nsew
flabel metal2 11898 1062 11940 3300 0 FreeSans 320 0 0 0 VDD_SW[3]
port 12 nsew
flabel metal2 9506 1062 9548 3300 0 FreeSans 320 0 0 0 VDD_SW[4]
port 13 nsew
flabel metal2 7114 1062 7156 3300 0 FreeSans 320 0 0 0 VDD_SW[5]
port 14 nsew
flabel metal2 4722 1062 4764 3300 0 FreeSans 320 0 0 0 VDD_SW[6]
port 15 nsew
flabel metal2 13924 1454 13966 3300 0 FreeSans 320 0 0 0 D[2]
port 17 nsew
flabel metal2 11531 1454 11573 3300 0 FreeSans 320 0 0 0 D[3]
port 18 nsew
flabel metal2 9140 1453 9182 3300 0 FreeSans 320 0 0 0 D[4]
port 19 nsew
flabel metal2 6747 1454 6789 3300 0 FreeSans 320 0 0 0 D[5]
port 20 nsew
flabel metal2 4356 1453 4398 3300 0 FreeSans 320 0 0 0 D[6]
port 21 nsew
flabel metal2 13519 1602 13561 3300 0 FreeSans 320 0 0 0 check[1]
port 24 nsew
flabel metal2 11130 1602 11172 3300 0 FreeSans 320 0 0 0 check[2]
port 25 nsew
flabel metal2 8738 1603 8780 3300 0 FreeSans 320 0 0 0 check[3]
port 26 nsew
flabel metal2 6344 1602 6386 3300 0 FreeSans 320 0 0 0 check[4]
port 27 nsew
flabel metal2 3954 1602 3996 3300 0 FreeSans 320 0 0 0 check[5]
port 28 nsew
flabel metal2 16682 1062 16724 3300 0 FreeSans 320 0 0 0 VDD_SW[1]
port 49 nsew
flabel metal2 1562 1603 1604 3300 0 FreeSans 320 0 0 0 check[6]
port 29 nsew
flabel metal2 1964 1453 2006 3300 0 FreeSans 320 0 0 0 D[7]
port 22 nsew
flabel metal2 2330 1062 2372 3300 0 FreeSans 320 0 0 0 VDD_SW[7]
port 16 nsew
flabel metal2 2533 345 2575 3300 0 FreeSans 320 0 0 0 VSS_SW[6]
port 9 nsew
flabel metal2 141 345 183 3300 0 FreeSans 320 0 0 0 VSS_SW[7]
port 10 nsew
rlabel comment s 4386 2410 4386 2410 4 buf_1
rlabel comment s 5214 2410 5214 2410 4 buf_16
rlabel comment s 4662 2410 4662 2410 4 buf_4
rlabel comment s 276 1268 276 1268 4 buf_4
rlabel comment s 828 1268 828 1268 4 buf_16
rlabel comment s 0 1268 0 1268 4 buf_1
rlabel comment s 3128 1268 3128 1268 4 buf_4
rlabel comment s 3680 1268 3680 1268 4 buf_16
rlabel comment s 2852 1268 2852 1268 4 buf_1
rlabel comment s 6216 1268 6216 1268 4 buf_1
rlabel comment s 7044 1268 7044 1268 4 buf_16
rlabel comment s 6492 1268 6492 1268 4 buf_4
rlabel comment s 9068 1268 9068 1268 4 buf_1
rlabel comment s 9896 1268 9896 1268 4 buf_16
rlabel comment s 9344 1268 9344 1268 4 buf_4
rlabel comment s 11982 1268 11982 1268 4 buf_1
rlabel comment s 12810 1268 12810 1268 4 buf_16
rlabel comment s 12258 1268 12258 1268 4 buf_4
rlabel comment s 13730 1268 13730 1268 4 buf_1
rlabel comment s 14558 1268 14558 1268 4 buf_16
rlabel comment s 14006 1268 14006 1268 4 buf_4
flabel metal2 16399 -322 16441 915 0 FreeSans 320 0 0 0 VDD_SW_b[1]
port 30 nsew
flabel metal2 14006 -322 14048 913 0 FreeSans 320 0 0 0 VDD_SW_b[2]
port 31 nsew
flabel metal2 11613 -322 11655 914 0 FreeSans 320 0 0 0 VDD_SW_b[3]
port 32 nsew
flabel metal2 9222 -322 9264 915 0 FreeSans 320 0 0 0 VDD_SW_b[4]
port 33 nsew
flabel metal2 4438 -322 4480 914 0 FreeSans 320 0 0 0 VDD_SW_b[6]
port 35 nsew
flabel metal2 2046 -322 2088 913 0 FreeSans 320 0 0 0 VDD_SW_b[7]
port 36 nsew
rlabel comment s 276 580 276 580 4 buf_4
rlabel comment s 828 580 828 580 4 buf_16
rlabel comment s 0 580 0 580 4 buf_1
rlabel comment s 2852 580 2852 580 4 buf_1
rlabel comment s 3680 580 3680 580 4 buf_16
rlabel comment s 3128 580 3128 580 4 buf_4
rlabel comment s 5980 580 5980 580 4 buf_4
rlabel comment s 6532 580 6532 580 4 buf_16
rlabel comment s 5704 580 5704 580 4 buf_1
rlabel comment s 8556 580 8556 580 4 buf_1
rlabel comment s 9384 580 9384 580 4 buf_16
rlabel comment s 8832 580 8832 580 4 buf_4
rlabel comment s 11408 580 11408 580 4 buf_1
rlabel comment s 12236 580 12236 580 4 buf_16
rlabel comment s 11684 580 11684 580 4 buf_4
rlabel comment s 14260 580 14260 580 4 buf_1
rlabel comment s 15088 580 15088 580 4 buf_16
rlabel comment s 14536 580 14536 580 4 buf_4
flabel metal2 14653 -343 14695 234 0 FreeSans 320 0 0 0 VSS_SW_b[1]
port 37 nsew
flabel metal2 12260 -343 12302 235 0 FreeSans 320 0 0 0 VSS_SW_b[2]
port 38 nsew
flabel metal2 9869 -343 9911 234 0 FreeSans 320 0 0 0 VSS_SW_b[3]
port 39 nsew
flabel metal2 7477 -343 7519 234 0 FreeSans 320 0 0 0 VSS_SW_b[4]
port 40 nsew
flabel metal2 5084 -343 5126 234 0 FreeSans 320 0 0 0 VSS_SW_b[5]
port 41 nsew
flabel metal2 2693 -343 2735 234 0 FreeSans 320 0 0 0 VSS_SW_b[6]
port 42 nsew
flabel metal2 301 -343 343 234 0 FreeSans 320 0 0 0 VSS_SW_b[7]
port 44 nsew
flabel metal2 14493 346 14535 3300 0 FreeSans 320 0 0 0 VSS_SW[1]
port 4 nsew
flabel metal2 12102 346 12144 3300 0 FreeSans 320 0 0 0 VSS_SW[2]
port 5 nsew
flabel metal1 -126 2526 4302 2560 0 FreeSans 320 0 0 0 ready
port 51 nsew
flabel metal1 -126 2722 -34 2756 0 FreeSans 320 0 0 0 reset
port 52 nsew
flabel metal2 6829 -322 6871 914 0 FreeSans 320 0 0 0 VDD_SW_b[5]
port 34 nsew
flabel metal4 12406 -75 16876 114 0 FreeSans 1600 0 0 0 VSS
port 59 nsew
flabel metal2 15914 1603 15956 3300 0 FreeSans 320 0 0 0 check[0]
port 23 nsew
flabel metal2 16317 1454 16359 3300 0 FreeSans 320 0 0 0 D[1]
port 46 nsew
flabel metal4 7278 2721 15690 3018 0 FreeSans 1600 0 0 0 VDD
port 61 nsew
flabel locali 14841 112 14875 146 0 FreeSans 400 0 0 0 x35.RESET_B
flabel locali 16681 -126 16715 -92 7 FreeSans 400 0 0 0 x35.VGND
flabel locali 16681 112 16715 146 0 FreeSans 400 0 0 0 x35.CLK_N
flabel locali 16681 180 16715 214 0 FreeSans 400 0 0 0 x35.CLK_N
flabel locali 15945 44 15979 78 0 FreeSans 400 0 0 0 x35.SET_B
flabel locali 14381 -24 14415 10 0 FreeSans 400 0 0 0 x35.Q
flabel locali 14381 248 14415 282 0 FreeSans 400 0 0 0 x35.Q
flabel locali 14381 316 14415 350 0 FreeSans 400 0 0 0 x35.Q
flabel locali 16681 418 16715 452 7 FreeSans 400 0 0 0 x35.VPWR
flabel locali 16313 112 16347 146 0 FreeSans 200 0 0 0 x35.D
flabel locali 16313 180 16347 214 0 FreeSans 200 0 0 0 x35.D
flabel locali 14657 316 14691 350 0 FreeSans 400 0 0 0 x35.Q_N
flabel locali 14657 248 14691 282 0 FreeSans 400 0 0 0 x35.Q_N
flabel locali 14657 -24 14691 10 0 FreeSans 400 0 0 0 x35.Q_N
flabel metal1 16681 -126 16715 -92 0 FreeSans 200 0 0 0 x35.VGND
flabel metal1 16681 418 16715 452 0 FreeSans 200 0 0 0 x35.VPWR
flabel nwell 16681 418 16715 452 7 FreeSans 400 0 0 0 x35.VPB
flabel nwell 16698 435 16698 435 0 FreeSans 200 0 0 0 x35.VPB
flabel pwell 16681 -126 16715 -92 7 FreeSans 400 0 0 0 x35.VNB
flabel pwell 16698 -109 16698 -109 0 FreeSans 200 0 0 0 x35.VNB
rlabel comment 16744 -109 16744 -109 6 x35.dfbbn_1
rlabel locali 15179 38 15288 104 1 x35.SET_B
rlabel metal1 15183 75 15241 84 1 x35.SET_B
rlabel metal1 15183 38 15241 47 1 x35.SET_B
rlabel metal1 15933 75 15991 84 1 x35.SET_B
rlabel metal1 15183 47 15991 75 1 x35.SET_B
rlabel metal1 15933 38 15991 47 1 x35.SET_B
rlabel metal1 14352 -157 16744 -61 1 x35.VGND
rlabel metal1 14352 387 16744 483 1 x35.VPWR
flabel locali 16221 801 16255 835 0 FreeSans 400 0 0 0 x34.RESET_B
flabel locali 14381 563 14415 597 3 FreeSans 400 0 0 0 x34.VGND
flabel locali 14381 801 14415 835 0 FreeSans 400 0 0 0 x34.CLK_N
flabel locali 14381 869 14415 903 0 FreeSans 400 0 0 0 x34.CLK_N
flabel locali 15117 733 15151 767 0 FreeSans 400 0 0 0 x34.SET_B
flabel locali 16681 665 16715 699 0 FreeSans 400 0 0 0 x34.Q
flabel locali 16681 937 16715 971 0 FreeSans 400 0 0 0 x34.Q
flabel locali 16681 1005 16715 1039 0 FreeSans 400 0 0 0 x34.Q
flabel locali 14381 1107 14415 1141 3 FreeSans 400 0 0 0 x34.VPWR
flabel locali 14749 801 14783 835 0 FreeSans 200 0 0 0 x34.D
flabel locali 14749 869 14783 903 0 FreeSans 200 0 0 0 x34.D
flabel locali 16405 1005 16439 1039 0 FreeSans 400 0 0 0 x34.Q_N
flabel locali 16405 937 16439 971 0 FreeSans 400 0 0 0 x34.Q_N
flabel locali 16405 665 16439 699 0 FreeSans 400 0 0 0 x34.Q_N
flabel metal1 14381 563 14415 597 0 FreeSans 200 0 0 0 x34.VGND
flabel metal1 14381 1107 14415 1141 0 FreeSans 200 0 0 0 x34.VPWR
flabel nwell 14381 1107 14415 1141 3 FreeSans 400 0 0 0 x34.VPB
flabel nwell 14398 1124 14398 1124 0 FreeSans 200 0 0 0 x34.VPB
flabel pwell 14381 563 14415 597 3 FreeSans 400 0 0 0 x34.VNB
flabel pwell 14398 580 14398 580 0 FreeSans 200 0 0 0 x34.VNB
rlabel comment 14352 580 14352 580 4 x34.dfbbn_1
rlabel locali 15808 727 15917 793 1 x34.SET_B
rlabel metal1 15855 764 15913 773 1 x34.SET_B
rlabel metal1 15855 727 15913 736 1 x34.SET_B
rlabel metal1 15105 764 15163 773 1 x34.SET_B
rlabel metal1 15105 736 15913 764 1 x34.SET_B
rlabel metal1 15105 727 15163 736 1 x34.SET_B
rlabel metal1 14352 532 16744 628 1 x34.VGND
rlabel metal1 14352 1076 16744 1172 1 x34.VPWR
flabel locali 12449 112 12483 146 0 FreeSans 400 0 0 0 x32.RESET_B
flabel locali 14289 -126 14323 -92 7 FreeSans 400 0 0 0 x32.VGND
flabel locali 14289 112 14323 146 0 FreeSans 400 0 0 0 x32.CLK_N
flabel locali 14289 180 14323 214 0 FreeSans 400 0 0 0 x32.CLK_N
flabel locali 13553 44 13587 78 0 FreeSans 400 0 0 0 x32.SET_B
flabel locali 11989 -24 12023 10 0 FreeSans 400 0 0 0 x32.Q
flabel locali 11989 248 12023 282 0 FreeSans 400 0 0 0 x32.Q
flabel locali 11989 316 12023 350 0 FreeSans 400 0 0 0 x32.Q
flabel locali 14289 418 14323 452 7 FreeSans 400 0 0 0 x32.VPWR
flabel locali 13921 112 13955 146 0 FreeSans 200 0 0 0 x32.D
flabel locali 13921 180 13955 214 0 FreeSans 200 0 0 0 x32.D
flabel locali 12265 316 12299 350 0 FreeSans 400 0 0 0 x32.Q_N
flabel locali 12265 248 12299 282 0 FreeSans 400 0 0 0 x32.Q_N
flabel locali 12265 -24 12299 10 0 FreeSans 400 0 0 0 x32.Q_N
flabel metal1 14289 -126 14323 -92 0 FreeSans 200 0 0 0 x32.VGND
flabel metal1 14289 418 14323 452 0 FreeSans 200 0 0 0 x32.VPWR
flabel nwell 14289 418 14323 452 7 FreeSans 400 0 0 0 x32.VPB
flabel nwell 14306 435 14306 435 0 FreeSans 200 0 0 0 x32.VPB
flabel pwell 14289 -126 14323 -92 7 FreeSans 400 0 0 0 x32.VNB
flabel pwell 14306 -109 14306 -109 0 FreeSans 200 0 0 0 x32.VNB
rlabel comment 14352 -109 14352 -109 6 x32.dfbbn_1
rlabel locali 12787 38 12896 104 1 x32.SET_B
rlabel metal1 12791 75 12849 84 1 x32.SET_B
rlabel metal1 12791 38 12849 47 1 x32.SET_B
rlabel metal1 13541 75 13599 84 1 x32.SET_B
rlabel metal1 12791 47 13599 75 1 x32.SET_B
rlabel metal1 13541 38 13599 47 1 x32.SET_B
rlabel metal1 11960 -157 14352 -61 1 x32.VGND
rlabel metal1 11960 387 14352 483 1 x32.VPWR
flabel locali 13829 801 13863 835 0 FreeSans 400 0 0 0 x31.RESET_B
flabel locali 11989 563 12023 597 3 FreeSans 400 0 0 0 x31.VGND
flabel locali 11989 801 12023 835 0 FreeSans 400 0 0 0 x31.CLK_N
flabel locali 11989 869 12023 903 0 FreeSans 400 0 0 0 x31.CLK_N
flabel locali 12725 733 12759 767 0 FreeSans 400 0 0 0 x31.SET_B
flabel locali 14289 665 14323 699 0 FreeSans 400 0 0 0 x31.Q
flabel locali 14289 937 14323 971 0 FreeSans 400 0 0 0 x31.Q
flabel locali 14289 1005 14323 1039 0 FreeSans 400 0 0 0 x31.Q
flabel locali 11989 1107 12023 1141 3 FreeSans 400 0 0 0 x31.VPWR
flabel locali 12357 801 12391 835 0 FreeSans 200 0 0 0 x31.D
flabel locali 12357 869 12391 903 0 FreeSans 200 0 0 0 x31.D
flabel locali 14013 1005 14047 1039 0 FreeSans 400 0 0 0 x31.Q_N
flabel locali 14013 937 14047 971 0 FreeSans 400 0 0 0 x31.Q_N
flabel locali 14013 665 14047 699 0 FreeSans 400 0 0 0 x31.Q_N
flabel metal1 11989 563 12023 597 0 FreeSans 200 0 0 0 x31.VGND
flabel metal1 11989 1107 12023 1141 0 FreeSans 200 0 0 0 x31.VPWR
flabel nwell 11989 1107 12023 1141 3 FreeSans 400 0 0 0 x31.VPB
flabel nwell 12006 1124 12006 1124 0 FreeSans 200 0 0 0 x31.VPB
flabel pwell 11989 563 12023 597 3 FreeSans 400 0 0 0 x31.VNB
flabel pwell 12006 580 12006 580 0 FreeSans 200 0 0 0 x31.VNB
rlabel comment 11960 580 11960 580 4 x31.dfbbn_1
rlabel locali 13416 727 13525 793 1 x31.SET_B
rlabel metal1 13463 764 13521 773 1 x31.SET_B
rlabel metal1 13463 727 13521 736 1 x31.SET_B
rlabel metal1 12713 764 12771 773 1 x31.SET_B
rlabel metal1 12713 736 13521 764 1 x31.SET_B
rlabel metal1 12713 727 12771 736 1 x31.SET_B
rlabel metal1 11960 532 14352 628 1 x31.VGND
rlabel metal1 11960 1076 14352 1172 1 x31.VPWR
flabel locali 5612 2631 5646 2665 0 FreeSans 200 0 0 0 x30.A
flabel locali 5520 2631 5554 2665 0 FreeSans 200 0 0 0 x30.A
flabel locali 7175 2631 7209 2665 0 FreeSans 200 0 0 0 x30.X
flabel locali 7175 2699 7209 2733 0 FreeSans 200 0 0 0 x30.X
flabel pwell 5244 2393 5278 2427 0 FreeSans 200 0 0 0 x30.VNB
flabel nwell 5244 2937 5278 2971 0 FreeSans 200 0 0 0 x30.VPB
flabel metal1 5244 2393 5278 2427 0 FreeSans 200 0 0 0 x30.VGND
flabel metal1 5244 2937 5278 2971 0 FreeSans 200 0 0 0 x30.VPWR
rlabel comment 5214 2410 5214 2410 4 x30.buf_16
rlabel metal1 5214 2362 7238 2458 1 x30.VGND
rlabel metal1 5214 2906 7238 3002 1 x30.VPWR
flabel locali 10057 112 10091 146 0 FreeSans 400 0 0 0 x29.RESET_B
flabel locali 11897 -126 11931 -92 7 FreeSans 400 0 0 0 x29.VGND
flabel locali 11897 112 11931 146 0 FreeSans 400 0 0 0 x29.CLK_N
flabel locali 11897 180 11931 214 0 FreeSans 400 0 0 0 x29.CLK_N
flabel locali 11161 44 11195 78 0 FreeSans 400 0 0 0 x29.SET_B
flabel locali 9597 -24 9631 10 0 FreeSans 400 0 0 0 x29.Q
flabel locali 9597 248 9631 282 0 FreeSans 400 0 0 0 x29.Q
flabel locali 9597 316 9631 350 0 FreeSans 400 0 0 0 x29.Q
flabel locali 11897 418 11931 452 7 FreeSans 400 0 0 0 x29.VPWR
flabel locali 11529 112 11563 146 0 FreeSans 200 0 0 0 x29.D
flabel locali 11529 180 11563 214 0 FreeSans 200 0 0 0 x29.D
flabel locali 9873 316 9907 350 0 FreeSans 400 0 0 0 x29.Q_N
flabel locali 9873 248 9907 282 0 FreeSans 400 0 0 0 x29.Q_N
flabel locali 9873 -24 9907 10 0 FreeSans 400 0 0 0 x29.Q_N
flabel metal1 11897 -126 11931 -92 0 FreeSans 200 0 0 0 x29.VGND
flabel metal1 11897 418 11931 452 0 FreeSans 200 0 0 0 x29.VPWR
flabel nwell 11897 418 11931 452 7 FreeSans 400 0 0 0 x29.VPB
flabel nwell 11914 435 11914 435 0 FreeSans 200 0 0 0 x29.VPB
flabel pwell 11897 -126 11931 -92 7 FreeSans 400 0 0 0 x29.VNB
flabel pwell 11914 -109 11914 -109 0 FreeSans 200 0 0 0 x29.VNB
rlabel comment 11960 -109 11960 -109 6 x29.dfbbn_1
rlabel locali 10395 38 10504 104 1 x29.SET_B
rlabel metal1 10399 75 10457 84 1 x29.SET_B
rlabel metal1 10399 38 10457 47 1 x29.SET_B
rlabel metal1 11149 75 11207 84 1 x29.SET_B
rlabel metal1 10399 47 11207 75 1 x29.SET_B
rlabel metal1 11149 38 11207 47 1 x29.SET_B
rlabel metal1 9568 -157 11960 -61 1 x29.VGND
rlabel metal1 9568 387 11960 483 1 x29.VPWR
flabel locali 11437 801 11471 835 0 FreeSans 400 0 0 0 x28.RESET_B
flabel locali 9597 563 9631 597 3 FreeSans 400 0 0 0 x28.VGND
flabel locali 9597 801 9631 835 0 FreeSans 400 0 0 0 x28.CLK_N
flabel locali 9597 869 9631 903 0 FreeSans 400 0 0 0 x28.CLK_N
flabel locali 10333 733 10367 767 0 FreeSans 400 0 0 0 x28.SET_B
flabel locali 11897 665 11931 699 0 FreeSans 400 0 0 0 x28.Q
flabel locali 11897 937 11931 971 0 FreeSans 400 0 0 0 x28.Q
flabel locali 11897 1005 11931 1039 0 FreeSans 400 0 0 0 x28.Q
flabel locali 9597 1107 9631 1141 3 FreeSans 400 0 0 0 x28.VPWR
flabel locali 9965 801 9999 835 0 FreeSans 200 0 0 0 x28.D
flabel locali 9965 869 9999 903 0 FreeSans 200 0 0 0 x28.D
flabel locali 11621 1005 11655 1039 0 FreeSans 400 0 0 0 x28.Q_N
flabel locali 11621 937 11655 971 0 FreeSans 400 0 0 0 x28.Q_N
flabel locali 11621 665 11655 699 0 FreeSans 400 0 0 0 x28.Q_N
flabel metal1 9597 563 9631 597 0 FreeSans 200 0 0 0 x28.VGND
flabel metal1 9597 1107 9631 1141 0 FreeSans 200 0 0 0 x28.VPWR
flabel nwell 9597 1107 9631 1141 3 FreeSans 400 0 0 0 x28.VPB
flabel nwell 9614 1124 9614 1124 0 FreeSans 200 0 0 0 x28.VPB
flabel pwell 9597 563 9631 597 3 FreeSans 400 0 0 0 x28.VNB
flabel pwell 9614 580 9614 580 0 FreeSans 200 0 0 0 x28.VNB
rlabel comment 9568 580 9568 580 4 x28.dfbbn_1
rlabel locali 11024 727 11133 793 1 x28.SET_B
rlabel metal1 11071 764 11129 773 1 x28.SET_B
rlabel metal1 11071 727 11129 736 1 x28.SET_B
rlabel metal1 10321 764 10379 773 1 x28.SET_B
rlabel metal1 10321 736 11129 764 1 x28.SET_B
rlabel metal1 10321 727 10379 736 1 x28.SET_B
rlabel metal1 9568 532 11960 628 1 x28.VGND
rlabel metal1 9568 1076 11960 1172 1 x28.VPWR
flabel metal1 4692 2937 4726 2971 0 FreeSans 200 0 0 0 x27.VPWR
flabel metal1 4692 2393 4726 2427 0 FreeSans 200 0 0 0 x27.VGND
flabel locali 4968 2631 5002 2665 0 FreeSans 200 0 0 0 x27.X
flabel locali 4968 2699 5002 2733 0 FreeSans 200 0 0 0 x27.X
flabel locali 4968 2563 5002 2597 0 FreeSans 200 0 0 0 x27.X
flabel locali 4692 2937 4726 2971 0 FreeSans 200 0 0 0 x27.VPWR
flabel locali 4692 2393 4726 2427 0 FreeSans 200 0 0 0 x27.VGND
flabel locali 4692 2631 4726 2665 0 FreeSans 200 0 0 0 x27.A
flabel nwell 4692 2937 4726 2971 0 FreeSans 200 0 0 0 x27.VPB
flabel pwell 4692 2393 4726 2427 0 FreeSans 200 0 0 0 x27.VNB
rlabel comment 4662 2410 4662 2410 4 x27.buf_4
rlabel metal1 4662 2362 5214 2458 1 x27.VGND
rlabel metal1 4662 2906 5214 3002 1 x27.VPWR
flabel locali 7665 112 7699 146 0 FreeSans 400 0 0 0 x26.RESET_B
flabel locali 9505 -126 9539 -92 7 FreeSans 400 0 0 0 x26.VGND
flabel locali 9505 112 9539 146 0 FreeSans 400 0 0 0 x26.CLK_N
flabel locali 9505 180 9539 214 0 FreeSans 400 0 0 0 x26.CLK_N
flabel locali 8769 44 8803 78 0 FreeSans 400 0 0 0 x26.SET_B
flabel locali 7205 -24 7239 10 0 FreeSans 400 0 0 0 x26.Q
flabel locali 7205 248 7239 282 0 FreeSans 400 0 0 0 x26.Q
flabel locali 7205 316 7239 350 0 FreeSans 400 0 0 0 x26.Q
flabel locali 9505 418 9539 452 7 FreeSans 400 0 0 0 x26.VPWR
flabel locali 9137 112 9171 146 0 FreeSans 200 0 0 0 x26.D
flabel locali 9137 180 9171 214 0 FreeSans 200 0 0 0 x26.D
flabel locali 7481 316 7515 350 0 FreeSans 400 0 0 0 x26.Q_N
flabel locali 7481 248 7515 282 0 FreeSans 400 0 0 0 x26.Q_N
flabel locali 7481 -24 7515 10 0 FreeSans 400 0 0 0 x26.Q_N
flabel metal1 9505 -126 9539 -92 0 FreeSans 200 0 0 0 x26.VGND
flabel metal1 9505 418 9539 452 0 FreeSans 200 0 0 0 x26.VPWR
flabel nwell 9505 418 9539 452 7 FreeSans 400 0 0 0 x26.VPB
flabel nwell 9522 435 9522 435 0 FreeSans 200 0 0 0 x26.VPB
flabel pwell 9505 -126 9539 -92 7 FreeSans 400 0 0 0 x26.VNB
flabel pwell 9522 -109 9522 -109 0 FreeSans 200 0 0 0 x26.VNB
rlabel comment 9568 -109 9568 -109 6 x26.dfbbn_1
rlabel locali 8003 38 8112 104 1 x26.SET_B
rlabel metal1 8007 75 8065 84 1 x26.SET_B
rlabel metal1 8007 38 8065 47 1 x26.SET_B
rlabel metal1 8757 75 8815 84 1 x26.SET_B
rlabel metal1 8007 47 8815 75 1 x26.SET_B
rlabel metal1 8757 38 8815 47 1 x26.SET_B
rlabel metal1 7176 -157 9568 -61 1 x26.VGND
rlabel metal1 7176 387 9568 483 1 x26.VPWR
flabel locali 9045 801 9079 835 0 FreeSans 400 0 0 0 x25.RESET_B
flabel locali 7205 563 7239 597 3 FreeSans 400 0 0 0 x25.VGND
flabel locali 7205 801 7239 835 0 FreeSans 400 0 0 0 x25.CLK_N
flabel locali 7205 869 7239 903 0 FreeSans 400 0 0 0 x25.CLK_N
flabel locali 7941 733 7975 767 0 FreeSans 400 0 0 0 x25.SET_B
flabel locali 9505 665 9539 699 0 FreeSans 400 0 0 0 x25.Q
flabel locali 9505 937 9539 971 0 FreeSans 400 0 0 0 x25.Q
flabel locali 9505 1005 9539 1039 0 FreeSans 400 0 0 0 x25.Q
flabel locali 7205 1107 7239 1141 3 FreeSans 400 0 0 0 x25.VPWR
flabel locali 7573 801 7607 835 0 FreeSans 200 0 0 0 x25.D
flabel locali 7573 869 7607 903 0 FreeSans 200 0 0 0 x25.D
flabel locali 9229 1005 9263 1039 0 FreeSans 400 0 0 0 x25.Q_N
flabel locali 9229 937 9263 971 0 FreeSans 400 0 0 0 x25.Q_N
flabel locali 9229 665 9263 699 0 FreeSans 400 0 0 0 x25.Q_N
flabel metal1 7205 563 7239 597 0 FreeSans 200 0 0 0 x25.VGND
flabel metal1 7205 1107 7239 1141 0 FreeSans 200 0 0 0 x25.VPWR
flabel nwell 7205 1107 7239 1141 3 FreeSans 400 0 0 0 x25.VPB
flabel nwell 7222 1124 7222 1124 0 FreeSans 200 0 0 0 x25.VPB
flabel pwell 7205 563 7239 597 3 FreeSans 400 0 0 0 x25.VNB
flabel pwell 7222 580 7222 580 0 FreeSans 200 0 0 0 x25.VNB
rlabel comment 7176 580 7176 580 4 x25.dfbbn_1
rlabel locali 8632 727 8741 793 1 x25.SET_B
rlabel metal1 8679 764 8737 773 1 x25.SET_B
rlabel metal1 8679 727 8737 736 1 x25.SET_B
rlabel metal1 7929 764 7987 773 1 x25.SET_B
rlabel metal1 7929 736 8737 764 1 x25.SET_B
rlabel metal1 7929 727 7987 736 1 x25.SET_B
rlabel metal1 7176 532 9568 628 1 x25.VGND
rlabel metal1 7176 1076 9568 1172 1 x25.VPWR
flabel locali 5273 112 5307 146 0 FreeSans 400 0 0 0 x24.RESET_B
flabel locali 7113 -126 7147 -92 7 FreeSans 400 0 0 0 x24.VGND
flabel locali 7113 112 7147 146 0 FreeSans 400 0 0 0 x24.CLK_N
flabel locali 7113 180 7147 214 0 FreeSans 400 0 0 0 x24.CLK_N
flabel locali 6377 44 6411 78 0 FreeSans 400 0 0 0 x24.SET_B
flabel locali 4813 -24 4847 10 0 FreeSans 400 0 0 0 x24.Q
flabel locali 4813 248 4847 282 0 FreeSans 400 0 0 0 x24.Q
flabel locali 4813 316 4847 350 0 FreeSans 400 0 0 0 x24.Q
flabel locali 7113 418 7147 452 7 FreeSans 400 0 0 0 x24.VPWR
flabel locali 6745 112 6779 146 0 FreeSans 200 0 0 0 x24.D
flabel locali 6745 180 6779 214 0 FreeSans 200 0 0 0 x24.D
flabel locali 5089 316 5123 350 0 FreeSans 400 0 0 0 x24.Q_N
flabel locali 5089 248 5123 282 0 FreeSans 400 0 0 0 x24.Q_N
flabel locali 5089 -24 5123 10 0 FreeSans 400 0 0 0 x24.Q_N
flabel metal1 7113 -126 7147 -92 0 FreeSans 200 0 0 0 x24.VGND
flabel metal1 7113 418 7147 452 0 FreeSans 200 0 0 0 x24.VPWR
flabel nwell 7113 418 7147 452 7 FreeSans 400 0 0 0 x24.VPB
flabel nwell 7130 435 7130 435 0 FreeSans 200 0 0 0 x24.VPB
flabel pwell 7113 -126 7147 -92 7 FreeSans 400 0 0 0 x24.VNB
flabel pwell 7130 -109 7130 -109 0 FreeSans 200 0 0 0 x24.VNB
rlabel comment 7176 -109 7176 -109 6 x24.dfbbn_1
rlabel locali 5611 38 5720 104 1 x24.SET_B
rlabel metal1 5615 75 5673 84 1 x24.SET_B
rlabel metal1 5615 38 5673 47 1 x24.SET_B
rlabel metal1 6365 75 6423 84 1 x24.SET_B
rlabel metal1 5615 47 6423 75 1 x24.SET_B
rlabel metal1 6365 38 6423 47 1 x24.SET_B
rlabel metal1 4784 -157 7176 -61 1 x24.VGND
rlabel metal1 4784 387 7176 483 1 x24.VPWR
flabel locali 6653 801 6687 835 0 FreeSans 400 0 0 0 x23.RESET_B
flabel locali 4813 563 4847 597 3 FreeSans 400 0 0 0 x23.VGND
flabel locali 4813 801 4847 835 0 FreeSans 400 0 0 0 x23.CLK_N
flabel locali 4813 869 4847 903 0 FreeSans 400 0 0 0 x23.CLK_N
flabel locali 5549 733 5583 767 0 FreeSans 400 0 0 0 x23.SET_B
flabel locali 7113 665 7147 699 0 FreeSans 400 0 0 0 x23.Q
flabel locali 7113 937 7147 971 0 FreeSans 400 0 0 0 x23.Q
flabel locali 7113 1005 7147 1039 0 FreeSans 400 0 0 0 x23.Q
flabel locali 4813 1107 4847 1141 3 FreeSans 400 0 0 0 x23.VPWR
flabel locali 5181 801 5215 835 0 FreeSans 200 0 0 0 x23.D
flabel locali 5181 869 5215 903 0 FreeSans 200 0 0 0 x23.D
flabel locali 6837 1005 6871 1039 0 FreeSans 400 0 0 0 x23.Q_N
flabel locali 6837 937 6871 971 0 FreeSans 400 0 0 0 x23.Q_N
flabel locali 6837 665 6871 699 0 FreeSans 400 0 0 0 x23.Q_N
flabel metal1 4813 563 4847 597 0 FreeSans 200 0 0 0 x23.VGND
flabel metal1 4813 1107 4847 1141 0 FreeSans 200 0 0 0 x23.VPWR
flabel nwell 4813 1107 4847 1141 3 FreeSans 400 0 0 0 x23.VPB
flabel nwell 4830 1124 4830 1124 0 FreeSans 200 0 0 0 x23.VPB
flabel pwell 4813 563 4847 597 3 FreeSans 400 0 0 0 x23.VNB
flabel pwell 4830 580 4830 580 0 FreeSans 200 0 0 0 x23.VNB
rlabel comment 4784 580 4784 580 4 x23.dfbbn_1
rlabel locali 6240 727 6349 793 1 x23.SET_B
rlabel metal1 6287 764 6345 773 1 x23.SET_B
rlabel metal1 6287 727 6345 736 1 x23.SET_B
rlabel metal1 5537 764 5595 773 1 x23.SET_B
rlabel metal1 5537 736 6345 764 1 x23.SET_B
rlabel metal1 5537 727 5595 736 1 x23.SET_B
rlabel metal1 4784 532 7176 628 1 x23.VGND
rlabel metal1 4784 1076 7176 1172 1 x23.VPWR
flabel metal1 4417 2393 4451 2427 0 FreeSans 200 0 0 0 x22.VGND
flabel metal1 4415 2937 4449 2971 0 FreeSans 200 0 0 0 x22.VPWR
flabel locali 4415 2937 4449 2971 0 FreeSans 200 0 0 0 x22.VPWR
flabel locali 4417 2393 4451 2427 0 FreeSans 200 0 0 0 x22.VGND
flabel locali 4597 2495 4631 2529 0 FreeSans 200 0 0 0 x22.X
flabel locali 4597 2767 4631 2801 0 FreeSans 200 0 0 0 x22.X
flabel locali 4597 2835 4631 2869 0 FreeSans 200 0 0 0 x22.X
flabel locali 4415 2631 4449 2665 0 FreeSans 200 0 0 0 x22.A
flabel nwell 4415 2937 4449 2971 0 FreeSans 200 0 0 0 x22.VPB
flabel pwell 4417 2393 4451 2427 0 FreeSans 200 0 0 0 x22.VNB
rlabel comment 4386 2410 4386 2410 4 x22.buf_1
rlabel metal1 4386 2362 4662 2458 1 x22.VGND
rlabel metal1 4386 2906 4662 3002 1 x22.VPWR
flabel locali 2881 112 2915 146 0 FreeSans 400 0 0 0 x21.RESET_B
flabel locali 4721 -126 4755 -92 7 FreeSans 400 0 0 0 x21.VGND
flabel locali 4721 112 4755 146 0 FreeSans 400 0 0 0 x21.CLK_N
flabel locali 4721 180 4755 214 0 FreeSans 400 0 0 0 x21.CLK_N
flabel locali 3985 44 4019 78 0 FreeSans 400 0 0 0 x21.SET_B
flabel locali 2421 -24 2455 10 0 FreeSans 400 0 0 0 x21.Q
flabel locali 2421 248 2455 282 0 FreeSans 400 0 0 0 x21.Q
flabel locali 2421 316 2455 350 0 FreeSans 400 0 0 0 x21.Q
flabel locali 4721 418 4755 452 7 FreeSans 400 0 0 0 x21.VPWR
flabel locali 4353 112 4387 146 0 FreeSans 200 0 0 0 x21.D
flabel locali 4353 180 4387 214 0 FreeSans 200 0 0 0 x21.D
flabel locali 2697 316 2731 350 0 FreeSans 400 0 0 0 x21.Q_N
flabel locali 2697 248 2731 282 0 FreeSans 400 0 0 0 x21.Q_N
flabel locali 2697 -24 2731 10 0 FreeSans 400 0 0 0 x21.Q_N
flabel metal1 4721 -126 4755 -92 0 FreeSans 200 0 0 0 x21.VGND
flabel metal1 4721 418 4755 452 0 FreeSans 200 0 0 0 x21.VPWR
flabel nwell 4721 418 4755 452 7 FreeSans 400 0 0 0 x21.VPB
flabel nwell 4738 435 4738 435 0 FreeSans 200 0 0 0 x21.VPB
flabel pwell 4721 -126 4755 -92 7 FreeSans 400 0 0 0 x21.VNB
flabel pwell 4738 -109 4738 -109 0 FreeSans 200 0 0 0 x21.VNB
rlabel comment 4784 -109 4784 -109 6 x21.dfbbn_1
rlabel locali 3219 38 3328 104 1 x21.SET_B
rlabel metal1 3223 75 3281 84 1 x21.SET_B
rlabel metal1 3223 38 3281 47 1 x21.SET_B
rlabel metal1 3973 75 4031 84 1 x21.SET_B
rlabel metal1 3223 47 4031 75 1 x21.SET_B
rlabel metal1 3973 38 4031 47 1 x21.SET_B
rlabel metal1 2392 -157 4784 -61 1 x21.VGND
rlabel metal1 2392 387 4784 483 1 x21.VPWR
flabel metal1 16550 1251 16584 1285 0 FreeSans 200 0 0 0 x20.VGND
flabel metal1 16550 1795 16584 1829 0 FreeSans 200 0 0 0 x20.VPWR
flabel locali 15906 1557 15940 1591 0 FreeSans 250 0 0 0 x20.S
flabel locali 15998 1557 16032 1591 0 FreeSans 250 0 0 0 x20.S
flabel locali 16090 1421 16124 1455 0 FreeSans 250 0 0 0 x20.A1
flabel locali 16090 1489 16124 1523 0 FreeSans 250 0 0 0 x20.A1
flabel locali 16182 1489 16216 1523 0 FreeSans 250 0 0 0 x20.A0
flabel locali 16550 1353 16584 1387 0 FreeSans 250 0 0 0 x20.X
flabel locali 16550 1625 16584 1659 0 FreeSans 250 0 0 0 x20.X
flabel locali 16550 1693 16584 1727 0 FreeSans 250 0 0 0 x20.X
flabel nwell 16506 1795 16540 1829 0 FreeSans 250 0 0 0 x20.VPB
flabel pwell 16496 1251 16530 1285 0 FreeSans 250 0 0 0 x20.VNB
rlabel comment 16614 1268 16614 1268 6 x20.mux2_1
rlabel metal1 15786 1220 16614 1316 1 x20.VGND
rlabel metal1 15786 1764 16614 1860 1 x20.VPWR
flabel locali 4261 801 4295 835 0 FreeSans 400 0 0 0 x19.RESET_B
flabel locali 2421 563 2455 597 3 FreeSans 400 0 0 0 x19.VGND
flabel locali 2421 801 2455 835 0 FreeSans 400 0 0 0 x19.CLK_N
flabel locali 2421 869 2455 903 0 FreeSans 400 0 0 0 x19.CLK_N
flabel locali 3157 733 3191 767 0 FreeSans 400 0 0 0 x19.SET_B
flabel locali 4721 665 4755 699 0 FreeSans 400 0 0 0 x19.Q
flabel locali 4721 937 4755 971 0 FreeSans 400 0 0 0 x19.Q
flabel locali 4721 1005 4755 1039 0 FreeSans 400 0 0 0 x19.Q
flabel locali 2421 1107 2455 1141 3 FreeSans 400 0 0 0 x19.VPWR
flabel locali 2789 801 2823 835 0 FreeSans 200 0 0 0 x19.D
flabel locali 2789 869 2823 903 0 FreeSans 200 0 0 0 x19.D
flabel locali 4445 1005 4479 1039 0 FreeSans 400 0 0 0 x19.Q_N
flabel locali 4445 937 4479 971 0 FreeSans 400 0 0 0 x19.Q_N
flabel locali 4445 665 4479 699 0 FreeSans 400 0 0 0 x19.Q_N
flabel metal1 2421 563 2455 597 0 FreeSans 200 0 0 0 x19.VGND
flabel metal1 2421 1107 2455 1141 0 FreeSans 200 0 0 0 x19.VPWR
flabel nwell 2421 1107 2455 1141 3 FreeSans 400 0 0 0 x19.VPB
flabel nwell 2438 1124 2438 1124 0 FreeSans 200 0 0 0 x19.VPB
flabel pwell 2421 563 2455 597 3 FreeSans 400 0 0 0 x19.VNB
flabel pwell 2438 580 2438 580 0 FreeSans 200 0 0 0 x19.VNB
rlabel comment 2392 580 2392 580 4 x19.dfbbn_1
rlabel locali 3848 727 3957 793 1 x19.SET_B
rlabel metal1 3895 764 3953 773 1 x19.SET_B
rlabel metal1 3895 727 3953 736 1 x19.SET_B
rlabel metal1 3145 764 3203 773 1 x19.SET_B
rlabel metal1 3145 736 3953 764 1 x19.SET_B
rlabel metal1 3145 727 3203 736 1 x19.SET_B
rlabel metal1 2392 532 4784 628 1 x19.VGND
rlabel metal1 2392 1076 4784 1172 1 x19.VPWR
flabel metal1 14382 1251 14416 1285 0 FreeSans 200 0 0 0 x18.VGND
flabel metal1 14382 1795 14416 1829 0 FreeSans 200 0 0 0 x18.VPWR
flabel locali 15026 1557 15060 1591 0 FreeSans 250 0 0 0 x18.S
flabel locali 14934 1557 14968 1591 0 FreeSans 250 0 0 0 x18.S
flabel locali 14842 1421 14876 1455 0 FreeSans 250 0 0 0 x18.A1
flabel locali 14842 1489 14876 1523 0 FreeSans 250 0 0 0 x18.A1
flabel locali 14750 1489 14784 1523 0 FreeSans 250 0 0 0 x18.A0
flabel locali 14382 1353 14416 1387 0 FreeSans 250 0 0 0 x18.X
flabel locali 14382 1625 14416 1659 0 FreeSans 250 0 0 0 x18.X
flabel locali 14382 1693 14416 1727 0 FreeSans 250 0 0 0 x18.X
flabel nwell 14426 1795 14460 1829 0 FreeSans 250 0 0 0 x18.VPB
flabel pwell 14436 1251 14470 1285 0 FreeSans 250 0 0 0 x18.VNB
rlabel comment 14352 1268 14352 1268 4 x18.mux2_1
rlabel metal1 14352 1220 15180 1316 1 x18.VGND
rlabel metal1 14352 1764 15180 1860 1 x18.VPWR
flabel metal1 14156 1251 14190 1285 0 FreeSans 200 0 0 0 x17.VGND
flabel metal1 14156 1795 14190 1829 0 FreeSans 200 0 0 0 x17.VPWR
flabel locali 13512 1557 13546 1591 0 FreeSans 250 0 0 0 x17.S
flabel locali 13604 1557 13638 1591 0 FreeSans 250 0 0 0 x17.S
flabel locali 13696 1421 13730 1455 0 FreeSans 250 0 0 0 x17.A1
flabel locali 13696 1489 13730 1523 0 FreeSans 250 0 0 0 x17.A1
flabel locali 13788 1489 13822 1523 0 FreeSans 250 0 0 0 x17.A0
flabel locali 14156 1353 14190 1387 0 FreeSans 250 0 0 0 x17.X
flabel locali 14156 1625 14190 1659 0 FreeSans 250 0 0 0 x17.X
flabel locali 14156 1693 14190 1727 0 FreeSans 250 0 0 0 x17.X
flabel nwell 14112 1795 14146 1829 0 FreeSans 250 0 0 0 x17.VPB
flabel pwell 14102 1251 14136 1285 0 FreeSans 250 0 0 0 x17.VNB
rlabel comment 14220 1268 14220 1268 6 x17.mux2_1
rlabel metal1 13392 1220 14220 1316 1 x17.VGND
rlabel metal1 13392 1764 14220 1860 1 x17.VPWR
flabel metal1 11990 1251 12024 1285 0 FreeSans 200 0 0 0 x16.VGND
flabel metal1 11990 1795 12024 1829 0 FreeSans 200 0 0 0 x16.VPWR
flabel locali 12634 1557 12668 1591 0 FreeSans 250 0 0 0 x16.S
flabel locali 12542 1557 12576 1591 0 FreeSans 250 0 0 0 x16.S
flabel locali 12450 1421 12484 1455 0 FreeSans 250 0 0 0 x16.A1
flabel locali 12450 1489 12484 1523 0 FreeSans 250 0 0 0 x16.A1
flabel locali 12358 1489 12392 1523 0 FreeSans 250 0 0 0 x16.A0
flabel locali 11990 1353 12024 1387 0 FreeSans 250 0 0 0 x16.X
flabel locali 11990 1625 12024 1659 0 FreeSans 250 0 0 0 x16.X
flabel locali 11990 1693 12024 1727 0 FreeSans 250 0 0 0 x16.X
flabel nwell 12034 1795 12068 1829 0 FreeSans 250 0 0 0 x16.VPB
flabel pwell 12044 1251 12078 1285 0 FreeSans 250 0 0 0 x16.VNB
rlabel comment 11960 1268 11960 1268 4 x16.mux2_1
rlabel metal1 11960 1220 12788 1316 1 x16.VGND
rlabel metal1 11960 1764 12788 1860 1 x16.VPWR
flabel metal1 11766 1251 11800 1285 0 FreeSans 200 0 0 0 x15.VGND
flabel metal1 11766 1795 11800 1829 0 FreeSans 200 0 0 0 x15.VPWR
flabel locali 11122 1557 11156 1591 0 FreeSans 250 0 0 0 x15.S
flabel locali 11214 1557 11248 1591 0 FreeSans 250 0 0 0 x15.S
flabel locali 11306 1421 11340 1455 0 FreeSans 250 0 0 0 x15.A1
flabel locali 11306 1489 11340 1523 0 FreeSans 250 0 0 0 x15.A1
flabel locali 11398 1489 11432 1523 0 FreeSans 250 0 0 0 x15.A0
flabel locali 11766 1353 11800 1387 0 FreeSans 250 0 0 0 x15.X
flabel locali 11766 1625 11800 1659 0 FreeSans 250 0 0 0 x15.X
flabel locali 11766 1693 11800 1727 0 FreeSans 250 0 0 0 x15.X
flabel nwell 11722 1795 11756 1829 0 FreeSans 250 0 0 0 x15.VPB
flabel pwell 11712 1251 11746 1285 0 FreeSans 250 0 0 0 x15.VNB
rlabel comment 11830 1268 11830 1268 6 x15.mux2_1
rlabel metal1 11002 1220 11830 1316 1 x15.VGND
rlabel metal1 11002 1764 11830 1860 1 x15.VPWR
flabel metal1 9598 1251 9632 1285 0 FreeSans 200 0 0 0 x14.VGND
flabel metal1 9598 1795 9632 1829 0 FreeSans 200 0 0 0 x14.VPWR
flabel locali 10242 1557 10276 1591 0 FreeSans 250 0 0 0 x14.S
flabel locali 10150 1557 10184 1591 0 FreeSans 250 0 0 0 x14.S
flabel locali 10058 1421 10092 1455 0 FreeSans 250 0 0 0 x14.A1
flabel locali 10058 1489 10092 1523 0 FreeSans 250 0 0 0 x14.A1
flabel locali 9966 1489 10000 1523 0 FreeSans 250 0 0 0 x14.A0
flabel locali 9598 1353 9632 1387 0 FreeSans 250 0 0 0 x14.X
flabel locali 9598 1625 9632 1659 0 FreeSans 250 0 0 0 x14.X
flabel locali 9598 1693 9632 1727 0 FreeSans 250 0 0 0 x14.X
flabel nwell 9642 1795 9676 1829 0 FreeSans 250 0 0 0 x14.VPB
flabel pwell 9652 1251 9686 1285 0 FreeSans 250 0 0 0 x14.VNB
rlabel comment 9568 1268 9568 1268 4 x14.mux2_1
rlabel metal1 9568 1220 10396 1316 1 x14.VGND
rlabel metal1 9568 1764 10396 1860 1 x14.VPWR
flabel metal1 9374 1251 9408 1285 0 FreeSans 200 0 0 0 x13.VGND
flabel metal1 9374 1795 9408 1829 0 FreeSans 200 0 0 0 x13.VPWR
flabel locali 8730 1557 8764 1591 0 FreeSans 250 0 0 0 x13.S
flabel locali 8822 1557 8856 1591 0 FreeSans 250 0 0 0 x13.S
flabel locali 8914 1421 8948 1455 0 FreeSans 250 0 0 0 x13.A1
flabel locali 8914 1489 8948 1523 0 FreeSans 250 0 0 0 x13.A1
flabel locali 9006 1489 9040 1523 0 FreeSans 250 0 0 0 x13.A0
flabel locali 9374 1353 9408 1387 0 FreeSans 250 0 0 0 x13.X
flabel locali 9374 1625 9408 1659 0 FreeSans 250 0 0 0 x13.X
flabel locali 9374 1693 9408 1727 0 FreeSans 250 0 0 0 x13.X
flabel nwell 9330 1795 9364 1829 0 FreeSans 250 0 0 0 x13.VPB
flabel pwell 9320 1251 9354 1285 0 FreeSans 250 0 0 0 x13.VNB
rlabel comment 9438 1268 9438 1268 6 x13.mux2_1
rlabel metal1 8610 1220 9438 1316 1 x13.VGND
rlabel metal1 8610 1764 9438 1860 1 x13.VPWR
flabel metal1 7206 1251 7240 1285 0 FreeSans 200 0 0 0 x12.VGND
flabel metal1 7206 1795 7240 1829 0 FreeSans 200 0 0 0 x12.VPWR
flabel locali 7850 1557 7884 1591 0 FreeSans 250 0 0 0 x12.S
flabel locali 7758 1557 7792 1591 0 FreeSans 250 0 0 0 x12.S
flabel locali 7666 1421 7700 1455 0 FreeSans 250 0 0 0 x12.A1
flabel locali 7666 1489 7700 1523 0 FreeSans 250 0 0 0 x12.A1
flabel locali 7574 1489 7608 1523 0 FreeSans 250 0 0 0 x12.A0
flabel locali 7206 1353 7240 1387 0 FreeSans 250 0 0 0 x12.X
flabel locali 7206 1625 7240 1659 0 FreeSans 250 0 0 0 x12.X
flabel locali 7206 1693 7240 1727 0 FreeSans 250 0 0 0 x12.X
flabel nwell 7250 1795 7284 1829 0 FreeSans 250 0 0 0 x12.VPB
flabel pwell 7260 1251 7294 1285 0 FreeSans 250 0 0 0 x12.VNB
rlabel comment 7176 1268 7176 1268 4 x12.mux2_1
rlabel metal1 7176 1220 8004 1316 1 x12.VGND
rlabel metal1 7176 1764 8004 1860 1 x12.VPWR
flabel metal1 6980 1251 7014 1285 0 FreeSans 200 0 0 0 x11.VGND
flabel metal1 6980 1795 7014 1829 0 FreeSans 200 0 0 0 x11.VPWR
flabel locali 6336 1557 6370 1591 0 FreeSans 250 0 0 0 x11.S
flabel locali 6428 1557 6462 1591 0 FreeSans 250 0 0 0 x11.S
flabel locali 6520 1421 6554 1455 0 FreeSans 250 0 0 0 x11.A1
flabel locali 6520 1489 6554 1523 0 FreeSans 250 0 0 0 x11.A1
flabel locali 6612 1489 6646 1523 0 FreeSans 250 0 0 0 x11.A0
flabel locali 6980 1353 7014 1387 0 FreeSans 250 0 0 0 x11.X
flabel locali 6980 1625 7014 1659 0 FreeSans 250 0 0 0 x11.X
flabel locali 6980 1693 7014 1727 0 FreeSans 250 0 0 0 x11.X
flabel nwell 6936 1795 6970 1829 0 FreeSans 250 0 0 0 x11.VPB
flabel pwell 6926 1251 6960 1285 0 FreeSans 250 0 0 0 x11.VNB
rlabel comment 7044 1268 7044 1268 6 x11.mux2_1
rlabel metal1 6216 1220 7044 1316 1 x11.VGND
rlabel metal1 6216 1764 7044 1860 1 x11.VPWR
flabel metal1 4814 1251 4848 1285 0 FreeSans 200 0 0 0 x10.VGND
flabel metal1 4814 1795 4848 1829 0 FreeSans 200 0 0 0 x10.VPWR
flabel locali 5458 1557 5492 1591 0 FreeSans 250 0 0 0 x10.S
flabel locali 5366 1557 5400 1591 0 FreeSans 250 0 0 0 x10.S
flabel locali 5274 1421 5308 1455 0 FreeSans 250 0 0 0 x10.A1
flabel locali 5274 1489 5308 1523 0 FreeSans 250 0 0 0 x10.A1
flabel locali 5182 1489 5216 1523 0 FreeSans 250 0 0 0 x10.A0
flabel locali 4814 1353 4848 1387 0 FreeSans 250 0 0 0 x10.X
flabel locali 4814 1625 4848 1659 0 FreeSans 250 0 0 0 x10.X
flabel locali 4814 1693 4848 1727 0 FreeSans 250 0 0 0 x10.X
flabel nwell 4858 1795 4892 1829 0 FreeSans 250 0 0 0 x10.VPB
flabel pwell 4868 1251 4902 1285 0 FreeSans 250 0 0 0 x10.VNB
rlabel comment 4784 1268 4784 1268 4 x10.mux2_1
rlabel metal1 4784 1220 5612 1316 1 x10.VGND
rlabel metal1 4784 1764 5612 1860 1 x10.VPWR
flabel metal1 4590 1251 4624 1285 0 FreeSans 200 0 0 0 x9.VGND
flabel metal1 4590 1795 4624 1829 0 FreeSans 200 0 0 0 x9.VPWR
flabel locali 3946 1557 3980 1591 0 FreeSans 250 0 0 0 x9.S
flabel locali 4038 1557 4072 1591 0 FreeSans 250 0 0 0 x9.S
flabel locali 4130 1421 4164 1455 0 FreeSans 250 0 0 0 x9.A1
flabel locali 4130 1489 4164 1523 0 FreeSans 250 0 0 0 x9.A1
flabel locali 4222 1489 4256 1523 0 FreeSans 250 0 0 0 x9.A0
flabel locali 4590 1353 4624 1387 0 FreeSans 250 0 0 0 x9.X
flabel locali 4590 1625 4624 1659 0 FreeSans 250 0 0 0 x9.X
flabel locali 4590 1693 4624 1727 0 FreeSans 250 0 0 0 x9.X
flabel nwell 4546 1795 4580 1829 0 FreeSans 250 0 0 0 x9.VPB
flabel pwell 4536 1251 4570 1285 0 FreeSans 250 0 0 0 x9.VNB
rlabel comment 4654 1268 4654 1268 6 x9.mux2_1
rlabel metal1 3826 1220 4654 1316 1 x9.VGND
rlabel metal1 3826 1764 4654 1860 1 x9.VPWR
flabel metal1 2422 1251 2456 1285 0 FreeSans 200 0 0 0 x8.VGND
flabel metal1 2422 1795 2456 1829 0 FreeSans 200 0 0 0 x8.VPWR
flabel locali 3066 1557 3100 1591 0 FreeSans 250 0 0 0 x8.S
flabel locali 2974 1557 3008 1591 0 FreeSans 250 0 0 0 x8.S
flabel locali 2882 1421 2916 1455 0 FreeSans 250 0 0 0 x8.A1
flabel locali 2882 1489 2916 1523 0 FreeSans 250 0 0 0 x8.A1
flabel locali 2790 1489 2824 1523 0 FreeSans 250 0 0 0 x8.A0
flabel locali 2422 1353 2456 1387 0 FreeSans 250 0 0 0 x8.X
flabel locali 2422 1625 2456 1659 0 FreeSans 250 0 0 0 x8.X
flabel locali 2422 1693 2456 1727 0 FreeSans 250 0 0 0 x8.X
flabel nwell 2466 1795 2500 1829 0 FreeSans 250 0 0 0 x8.VPB
flabel pwell 2476 1251 2510 1285 0 FreeSans 250 0 0 0 x8.VNB
rlabel comment 2392 1268 2392 1268 4 x8.mux2_1
rlabel metal1 2392 1220 3220 1316 1 x8.VGND
rlabel metal1 2392 1764 3220 1860 1 x8.VPWR
flabel metal1 2198 1251 2232 1285 0 FreeSans 200 0 0 0 x7.VGND
flabel metal1 2198 1795 2232 1829 0 FreeSans 200 0 0 0 x7.VPWR
flabel locali 1554 1557 1588 1591 0 FreeSans 250 0 0 0 x7.S
flabel locali 1646 1557 1680 1591 0 FreeSans 250 0 0 0 x7.S
flabel locali 1738 1421 1772 1455 0 FreeSans 250 0 0 0 x7.A1
flabel locali 1738 1489 1772 1523 0 FreeSans 250 0 0 0 x7.A1
flabel locali 1830 1489 1864 1523 0 FreeSans 250 0 0 0 x7.A0
flabel locali 2198 1353 2232 1387 0 FreeSans 250 0 0 0 x7.X
flabel locali 2198 1625 2232 1659 0 FreeSans 250 0 0 0 x7.X
flabel locali 2198 1693 2232 1727 0 FreeSans 250 0 0 0 x7.X
flabel nwell 2154 1795 2188 1829 0 FreeSans 250 0 0 0 x7.VPB
flabel pwell 2144 1251 2178 1285 0 FreeSans 250 0 0 0 x7.VNB
rlabel comment 2262 1268 2262 1268 6 x7.mux2_1
rlabel metal1 1434 1220 2262 1316 1 x7.VGND
rlabel metal1 1434 1764 2262 1860 1 x7.VPWR
flabel metal1 30 1251 64 1285 0 FreeSans 200 0 0 0 x6.VGND
flabel metal1 30 1795 64 1829 0 FreeSans 200 0 0 0 x6.VPWR
flabel locali 674 1557 708 1591 0 FreeSans 250 0 0 0 x6.S
flabel locali 582 1557 616 1591 0 FreeSans 250 0 0 0 x6.S
flabel locali 490 1421 524 1455 0 FreeSans 250 0 0 0 x6.A1
flabel locali 490 1489 524 1523 0 FreeSans 250 0 0 0 x6.A1
flabel locali 398 1489 432 1523 0 FreeSans 250 0 0 0 x6.A0
flabel locali 30 1353 64 1387 0 FreeSans 250 0 0 0 x6.X
flabel locali 30 1625 64 1659 0 FreeSans 250 0 0 0 x6.X
flabel locali 30 1693 64 1727 0 FreeSans 250 0 0 0 x6.X
flabel nwell 74 1795 108 1829 0 FreeSans 250 0 0 0 x6.VPB
flabel pwell 84 1251 118 1285 0 FreeSans 250 0 0 0 x6.VNB
rlabel comment 0 1268 0 1268 4 x6.mux2_1
rlabel metal1 0 1220 828 1316 1 x6.VGND
rlabel metal1 0 1764 828 1860 1 x6.VPWR
flabel locali 489 112 523 146 0 FreeSans 400 0 0 0 x5.RESET_B
flabel locali 2329 -126 2363 -92 7 FreeSans 400 0 0 0 x5.VGND
flabel locali 2329 112 2363 146 0 FreeSans 400 0 0 0 x5.CLK_N
flabel locali 2329 180 2363 214 0 FreeSans 400 0 0 0 x5.CLK_N
flabel locali 1593 44 1627 78 0 FreeSans 400 0 0 0 x5.SET_B
flabel locali 29 -24 63 10 0 FreeSans 400 0 0 0 x5.Q
flabel locali 29 248 63 282 0 FreeSans 400 0 0 0 x5.Q
flabel locali 29 316 63 350 0 FreeSans 400 0 0 0 x5.Q
flabel locali 2329 418 2363 452 7 FreeSans 400 0 0 0 x5.VPWR
flabel locali 1961 112 1995 146 0 FreeSans 200 0 0 0 x5.D
flabel locali 1961 180 1995 214 0 FreeSans 200 0 0 0 x5.D
flabel locali 305 316 339 350 0 FreeSans 400 0 0 0 x5.Q_N
flabel locali 305 248 339 282 0 FreeSans 400 0 0 0 x5.Q_N
flabel locali 305 -24 339 10 0 FreeSans 400 0 0 0 x5.Q_N
flabel metal1 2329 -126 2363 -92 0 FreeSans 200 0 0 0 x5.VGND
flabel metal1 2329 418 2363 452 0 FreeSans 200 0 0 0 x5.VPWR
flabel nwell 2329 418 2363 452 7 FreeSans 400 0 0 0 x5.VPB
flabel nwell 2346 435 2346 435 0 FreeSans 200 0 0 0 x5.VPB
flabel pwell 2329 -126 2363 -92 7 FreeSans 400 0 0 0 x5.VNB
flabel pwell 2346 -109 2346 -109 0 FreeSans 200 0 0 0 x5.VNB
rlabel comment 2392 -109 2392 -109 6 x5.dfbbn_1
rlabel locali 827 38 936 104 1 x5.SET_B
rlabel metal1 831 75 889 84 1 x5.SET_B
rlabel metal1 831 38 889 47 1 x5.SET_B
rlabel metal1 1581 75 1639 84 1 x5.SET_B
rlabel metal1 831 47 1639 75 1 x5.SET_B
rlabel metal1 1581 38 1639 47 1 x5.SET_B
rlabel metal1 0 -157 2392 -61 1 x5.VGND
rlabel metal1 0 387 2392 483 1 x5.VPWR
flabel metal1 308 2937 342 2971 0 FreeSans 200 0 0 0 x3.VPWR
flabel metal1 308 2393 342 2427 0 FreeSans 200 0 0 0 x3.VGND
flabel locali 584 2631 618 2665 0 FreeSans 200 0 0 0 x3.X
flabel locali 584 2699 618 2733 0 FreeSans 200 0 0 0 x3.X
flabel locali 584 2563 618 2597 0 FreeSans 200 0 0 0 x3.X
flabel locali 308 2937 342 2971 0 FreeSans 200 0 0 0 x3.VPWR
flabel locali 308 2393 342 2427 0 FreeSans 200 0 0 0 x3.VGND
flabel locali 308 2631 342 2665 0 FreeSans 200 0 0 0 x3.A
flabel nwell 308 2937 342 2971 0 FreeSans 200 0 0 0 x3.VPB
flabel pwell 308 2393 342 2427 0 FreeSans 200 0 0 0 x3.VNB
rlabel comment 278 2410 278 2410 4 x3.buf_4
rlabel metal1 278 2362 830 2458 1 x3.VGND
rlabel metal1 278 2906 830 3002 1 x3.VPWR
flabel locali 1228 2631 1262 2665 0 FreeSans 200 0 0 0 x2.A
flabel locali 1136 2631 1170 2665 0 FreeSans 200 0 0 0 x2.A
flabel locali 2791 2631 2825 2665 0 FreeSans 200 0 0 0 x2.X
flabel locali 2791 2699 2825 2733 0 FreeSans 200 0 0 0 x2.X
flabel pwell 860 2393 894 2427 0 FreeSans 200 0 0 0 x2.VNB
flabel nwell 860 2937 894 2971 0 FreeSans 200 0 0 0 x2.VPB
flabel metal1 860 2393 894 2427 0 FreeSans 200 0 0 0 x2.VGND
flabel metal1 860 2937 894 2971 0 FreeSans 200 0 0 0 x2.VPWR
rlabel comment 830 2410 830 2410 4 x2.buf_16
rlabel metal1 830 2362 2854 2458 1 x2.VGND
rlabel metal1 830 2906 2854 3002 1 x2.VPWR
flabel metal1 33 2393 67 2427 0 FreeSans 200 0 0 0 x1.VGND
flabel metal1 31 2937 65 2971 0 FreeSans 200 0 0 0 x1.VPWR
flabel locali 31 2937 65 2971 0 FreeSans 200 0 0 0 x1.VPWR
flabel locali 33 2393 67 2427 0 FreeSans 200 0 0 0 x1.VGND
flabel locali 213 2495 247 2529 0 FreeSans 200 0 0 0 x1.X
flabel locali 213 2767 247 2801 0 FreeSans 200 0 0 0 x1.X
flabel locali 213 2835 247 2869 0 FreeSans 200 0 0 0 x1.X
flabel locali 31 2631 65 2665 0 FreeSans 200 0 0 0 x1.A
flabel nwell 31 2937 65 2971 0 FreeSans 200 0 0 0 x1.VPB
flabel pwell 33 2393 67 2427 0 FreeSans 200 0 0 0 x1.VNB
rlabel comment 2 2410 2 2410 4 x1.buf_1
rlabel metal1 2 2362 278 2458 1 x1.VGND
rlabel metal1 2 2906 278 3002 1 x1.VPWR
flabel locali 1869 801 1903 835 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfbbn_1_0.RESET_B
flabel locali 29 563 63 597 3 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfbbn_1_0.VGND
flabel locali 29 801 63 835 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfbbn_1_0.CLK_N
flabel locali 29 869 63 903 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfbbn_1_0.CLK_N
flabel locali 765 733 799 767 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfbbn_1_0.SET_B
flabel locali 2329 665 2363 699 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfbbn_1_0.Q
flabel locali 2329 937 2363 971 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfbbn_1_0.Q
flabel locali 2329 1005 2363 1039 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfbbn_1_0.Q
flabel locali 29 1107 63 1141 3 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfbbn_1_0.VPWR
flabel locali 397 801 431 835 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfbbn_1_0.D
flabel locali 397 869 431 903 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfbbn_1_0.D
flabel locali 2053 1005 2087 1039 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfbbn_1_0.Q_N
flabel locali 2053 937 2087 971 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfbbn_1_0.Q_N
flabel locali 2053 665 2087 699 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfbbn_1_0.Q_N
flabel metal1 29 563 63 597 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfbbn_1_0.VGND
flabel metal1 29 1107 63 1141 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfbbn_1_0.VPWR
flabel nwell 29 1107 63 1141 3 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfbbn_1_0.VPB
flabel nwell 46 1124 46 1124 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfbbn_1_0.VPB
flabel pwell 29 563 63 597 3 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfbbn_1_0.VNB
flabel pwell 46 580 46 580 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfbbn_1_0.VNB
rlabel comment 0 580 0 580 4 sky130_fd_sc_hd__dfbbn_1_0.dfbbn_1
rlabel locali 1456 727 1565 793 1 sky130_fd_sc_hd__dfbbn_1_0.SET_B
rlabel metal1 1503 764 1561 773 1 sky130_fd_sc_hd__dfbbn_1_0.SET_B
rlabel metal1 1503 727 1561 736 1 sky130_fd_sc_hd__dfbbn_1_0.SET_B
rlabel metal1 753 764 811 773 1 sky130_fd_sc_hd__dfbbn_1_0.SET_B
rlabel metal1 753 736 1561 764 1 sky130_fd_sc_hd__dfbbn_1_0.SET_B
rlabel metal1 753 727 811 736 1 sky130_fd_sc_hd__dfbbn_1_0.SET_B
rlabel metal1 0 532 2392 628 1 sky130_fd_sc_hd__dfbbn_1_0.VGND
rlabel metal1 0 1076 2392 1172 1 sky130_fd_sc_hd__dfbbn_1_0.VPWR
<< end >>
