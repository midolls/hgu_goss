magic
tech sky130A
magscale 1 2
timestamp 1698857008
<< checkpaint >>
rect -1260 -660 28280 4586
rect -1260 -10460 1460 -660
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 0 -6400 200 -6200
rect 0 -6800 200 -6600
rect 0 -7200 200 -7000
rect 0 -7600 200 -7400
rect 0 -8000 200 -7800
rect 0 -8400 200 -8200
rect 0 -8800 200 -8600
rect 0 -9200 200 -9000
use hgu_delay_no_code  x1
timestamp 1698844916
transform 1 0 -2483 0 1 333
box 9238 267 15993 2993
use hgu_delay_no_code  x2
timestamp 1698844916
transform 1 0 4272 0 1 333
box 9238 267 15993 2993
use hgu_delay_no_code  x3
timestamp 1698844916
transform 1 0 11027 0 1 333
box 9238 267 15993 2993
use hgu_delay_no_code  x4
timestamp 1698844916
transform 1 0 -9238 0 1 333
box 9238 267 15993 2993
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 IN
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 OUT
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE1\[0\]}
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE1\[1\]}
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE1\[2\]}
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 {}
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE1\[3\]}
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE2\[0\]}
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE2\[1\]}
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE2\[2\]}
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE2\[3\]}
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE3\[0\]}
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 {}
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE3\[1\]}
port 15 nsew
flabel metal1 0 -6400 200 -6200 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE3\[2\]}
port 16 nsew
flabel metal1 0 -6800 200 -6600 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE3\[3\]}
port 17 nsew
flabel metal1 0 -7200 200 -7000 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE0\[0\]}
port 18 nsew
flabel metal1 0 -7600 200 -7400 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE0\[1\]}
port 19 nsew
flabel metal1 0 -8000 200 -7800 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE0\[2\]}
port 20 nsew
flabel metal1 0 -8400 200 -8200 0 FreeSans 256 0 0 0 {}
port 21 nsew
flabel metal1 0 -8800 200 -8600 0 FreeSans 256 0 0 0 {CAP_CTRL_CODE0\[3\]}
port 22 nsew
flabel metal1 0 -9200 200 -9000 0 FreeSans 256 0 0 0 sample_delay_offset
port 23 nsew
<< end >>
