* NGSPICE file created from hgu_cdac_half_flat.ext - technology: sky130A

.subckt hgu_cdac_half_flat tu tub
X0 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X1 inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF a_3540_5180# hgu_cdac_8bit_array_2.drv<7:0> inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X2 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X4 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X5 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X6 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X7 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X8 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X9 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X10 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X11 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X12 hgu_inverter_1.VSS a_5521_5720# hgu_cdac_8bit_array_3.drv<15:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X13 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X14 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X15 hgu_inverter_1.VSS a_8105_5185# hgu_cdac_8bit_array_2.drv<15:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X16 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X17 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X18 hgu_cdac_8bit_array_3.drv<7:0> a_2970_5870# inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X19 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X20 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X21 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X22 hgu_cdac_8bit_array_2.drv<1:0> a_657_5185# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X23 hgu_inverter_1.VSS a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X24 hgu_inverter_1.VSS a_5521_5720# hgu_cdac_8bit_array_3.drv<15:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X25 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X26 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X27 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X28 hgu_cdac_8bit_array_2.drv<7:0> a_3540_5180# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X29 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X30 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_8105_5185# hgu_cdac_8bit_array_2.drv<15:0> inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X31 hgu_cdac_8bit_array_3.drv<7:0> a_2970_5870# inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X32 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X33 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X34 hgu_cdac_8bit_array_3.drv<15:0> a_5521_5720# inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X35 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X36 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_5521_5720# hgu_cdac_8bit_array_3.drv<15:0> inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X37 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X38 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X39 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X40 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X41 hgu_cdac_8bit_array_2.drv<7:0> a_3540_5180# inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X42 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X43 hgu_inverter_1.VSS a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X44 hgu_cdac_8bit_array_2.drv<1:0> a_657_5185# inv_2_test_0/x2.VREF inv_2_test_0/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X45 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X46 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X47 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X48 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X49 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X50 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X51 inv_4_test_2/inv_2_test_1/x2.VREF a_1437_5881# hgu_cdac_8bit_array_3.drv<3:0> inv_4_test_2/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X52 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X53 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X54 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X55 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X56 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X57 hgu_inverter_1.VSS a_5521_5720# hgu_cdac_8bit_array_3.drv<15:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X58 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X59 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X60 hgu_cdac_8bit_array_2.drv<3:0> a_1921_5185# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X61 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X62 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X63 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X64 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X65 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_5521_5720# hgu_cdac_8bit_array_3.drv<15:0> inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X66 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X67 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X68 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X69 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X70 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X71 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X72 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X73 hgu_cdac_8bit_array_3.drv<15:0> a_5521_5720# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X74 hgu_cdac_8bit_array_2.drv<3:0> a_1921_5185# inv_4_test_1/inv_2_test_1/x2.VREF inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X75 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X76 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X77 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_5521_5720# hgu_cdac_8bit_array_3.drv<15:0> inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X78 hgu_cdac_8bit_array_2.drv<15:0> a_8105_5185# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X79 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X80 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X81 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X82 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X83 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X84 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X85 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X86 hgu_cdac_8bit_array_2.drv<15:0> a_8105_5185# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X87 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X88 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X89 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X90 hgu_cdac_8bit_array_2.drv<15:0> a_8105_5185# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X91 hgu_cdac_8bit_array_2.drv<15:0> a_8105_5185# inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X92 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X93 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X94 inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF a_3540_5180# hgu_cdac_8bit_array_2.drv<7:0> inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X95 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X96 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X97 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X98 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X99 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X100 hgu_inverter_1.VSS a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X101 hgu_cdac_8bit_array_2.drv<15:0> a_8105_5185# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X102 hgu_cdac_8bit_array_2.drv<15:0> a_8105_5185# inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X103 hgu_cdac_8bit_array_2.drv<15:0> a_8105_5185# inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X104 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X105 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X106 hgu_inverter_1.VSS a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X107 hgu_inverter_1.VSS a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X108 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X109 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X110 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X111 hgu_cdac_8bit_array_3.drv<15:0> a_5521_5720# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X112 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X113 hgu_inverter_1.VSS a_1437_5881# hgu_cdac_8bit_array_3.drv<3:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X114 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X115 hgu_cdac_8bit_array_2.drv<7:0> a_3540_5180# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X116 hgu_cdac_8bit_array_2.drv<15:0> a_8105_5185# inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X117 hgu_cdac_8bit_array_3.drv<3:0> a_1437_5881# inv_4_test_2/inv_2_test_1/x2.VREF inv_4_test_2/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X118 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X119 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X120 hgu_inverter_1.VSS a_1921_5185# hgu_cdac_8bit_array_2.drv<3:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X121 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X122 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X123 hgu_cdac_8bit_array_3.drv<15:0> a_5521_5720# inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X124 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X125 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X126 hgu_inverter_1.VSS a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X127 hgu_inverter_1.VSS a_5521_5720# hgu_cdac_8bit_array_3.drv<15:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X128 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X129 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X130 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X131 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X132 hgu_cdac_8bit_array_3.drv<15:0> a_5521_5720# inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X133 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X134 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X135 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X136 inv_4_test_1/inv_2_test_1/x2.VREF a_1921_5185# hgu_cdac_8bit_array_2.drv<3:0> inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X137 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X138 hgu_inverter_1.VSS a_2970_5870# hgu_cdac_8bit_array_3.drv<7:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X139 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X140 hgu_inverter_1.VSS a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X141 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X142 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X143 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X144 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X145 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X146 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X147 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X148 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X149 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X150 hgu_cdac_8bit_array_2.drv<7:0> a_3540_5180# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X151 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X152 hgu_cdac_8bit_array_2.drv<3:0> a_1921_5185# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X153 hgu_inverter_1.VSS a_2970_5870# hgu_cdac_8bit_array_3.drv<7:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X154 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X155 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X156 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X157 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X158 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X159 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X160 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X161 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X162 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X163 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X164 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X165 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X166 hgu_inverter_1.VSS a_8105_5185# hgu_cdac_8bit_array_2.drv<15:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X167 hgu_cdac_8bit_array_2.drv<3:0> a_1921_5185# inv_4_test_1/inv_2_test_1/x2.VREF inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X168 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X169 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X170 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X171 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X172 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X173 hgu_inverter_1.VSS a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X174 hgu_cdac_8bit_array_3.drv<1:0> a_528_5873# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X175 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X176 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X177 hgu_inverter_1.VSS a_3540_5180# hgu_cdac_8bit_array_2.drv<7:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X178 hgu_inverter_1.VSS a_8105_5185# hgu_cdac_8bit_array_2.drv<15:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X179 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X180 hgu_cdac_8bit_array_3.drv<7:0> a_2970_5870# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X181 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_5521_5720# hgu_cdac_8bit_array_3.drv<15:0> inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X182 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X183 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X184 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X185 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_8105_5185# hgu_cdac_8bit_array_2.drv<15:0> inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X186 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X187 hgu_inverter_1.VSS a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X188 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X189 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X190 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X191 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X192 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X193 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X194 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X195 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_5521_5720# hgu_cdac_8bit_array_3.drv<15:0> inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X196 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X197 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_8105_5185# hgu_cdac_8bit_array_2.drv<15:0> inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X198 hgu_inverter_1.VSS a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X199 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X200 hgu_cdac_8bit_array_2.drv<7:0> a_3540_5180# inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X201 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X202 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X203 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X204 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X205 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X206 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X207 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X208 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X209 inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_2970_5870# hgu_cdac_8bit_array_3.drv<7:0> inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X210 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X211 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X212 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X213 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X214 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X215 hgu_inverter_1.VSS a_657_5185# hgu_cdac_8bit_array_2.drv<1:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X216 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X217 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X218 hgu_cdac_8bit_array_3.drv<15:0> a_5521_5720# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X219 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X220 hgu_inverter_1.VSS a_3540_5180# hgu_cdac_8bit_array_2.drv<7:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X221 inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_2970_5870# hgu_cdac_8bit_array_3.drv<7:0> inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X222 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X223 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_5521_5720# hgu_cdac_8bit_array_3.drv<15:0> inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X224 hgu_inverter_1.VSS a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X225 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X226 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X227 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X228 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X229 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X230 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X231 inv_2_test_0/x2.VREF a_657_5185# hgu_cdac_8bit_array_2.drv<1:0> inv_2_test_0/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X232 hgu_cdac_8bit_array_3.drv<15:0> a_5521_5720# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X233 hgu_inverter_1.VSS a_8105_5185# hgu_cdac_8bit_array_2.drv<15:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X234 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X235 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X236 hgu_cdac_8bit_array_3.drv<15:0> a_5521_5720# inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X237 hgu_cdac_8bit_array_2.drv<15:0> a_8105_5185# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X238 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X239 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X240 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X241 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X242 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X243 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X244 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X245 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_8105_5185# hgu_cdac_8bit_array_2.drv<15:0> inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X246 hgu_cdac_8bit_array_3.drv<1:0> a_528_5873# inv_2_test_1/x2.VREF inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X247 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X248 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X249 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X250 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X251 hgu_cdac_8bit_array_3.drv<7:0> a_2970_5870# inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X252 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X253 hgu_cdac_8bit_array_2.drv<15:0> a_8105_5185# inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X254 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X255 hgu_inverter_1.VSS a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X256 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X257 hgu_inverter_1.VSS a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X258 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X259 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X260 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X261 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X262 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X263 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X264 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X265 hgu_inverter_1.VSS a_8105_5185# hgu_cdac_8bit_array_2.drv<15:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X266 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X267 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X268 hgu_inverter_1.VSS a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X269 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X270 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X271 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X272 hgu_inverter_1.VSS a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X273 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X274 hgu_inverter_1.VSS a_8105_5185# hgu_cdac_8bit_array_2.drv<15:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X275 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X276 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X277 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X278 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_8105_5185# hgu_cdac_8bit_array_2.drv<15:0> inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X279 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X280 hgu_cdac_8bit_array_3.drv<15:0> a_5521_5720# inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X281 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X282 hgu_cdac_8bit_array_2.drv<7:0> a_3540_5180# inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X283 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X284 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X285 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X286 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X287 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X288 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X289 hgu_inverter_1.VSS a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X290 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X291 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_5521_5720# hgu_cdac_8bit_array_3.drv<15:0> inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X292 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X293 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_8105_5185# hgu_cdac_8bit_array_2.drv<15:0> inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X294 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X295 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X296 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X297 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X298 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X299 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X300 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X301 hgu_inverter_1.VSS a_5521_5720# hgu_cdac_8bit_array_3.drv<15:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X302 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X303 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X304 hgu_inverter_1.VSS a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X305 hgu_cdac_8bit_array_3.drv<3:0> a_1437_5881# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X306 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X307 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X308 inv_4_test_2/inv_2_test_1/x2.VREF a_1437_5881# hgu_cdac_8bit_array_3.drv<3:0> inv_4_test_2/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X309 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X310 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X311 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X312 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X313 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X314 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X315 hgu_cdac_8bit_array_3.drv<15:0> a_5521_5720# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X316 hgu_cdac_8bit_array_2.drv<7:0> a_3540_5180# inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X317 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X318 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X319 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X320 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X321 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X322 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X323 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X324 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X325 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X326 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X327 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X328 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X329 hgu_inverter_1.VSS a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X330 hgu_inverter_1.VSS a_3540_5180# hgu_cdac_8bit_array_2.drv<7:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X331 hgu_cdac_8bit_array_3.drv<7:0> a_2970_5870# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X332 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X333 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X334 hgu_inverter_1.VSS a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X335 hgu_inverter_1.VSS a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X336 inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF a_3540_5180# hgu_cdac_8bit_array_2.drv<7:0> inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X337 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X338 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X339 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X340 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X341 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X342 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X343 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X344 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X345 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X346 hgu_cdac_8bit_array_2.drv<15:0> a_8105_5185# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X347 hgu_inverter_1.VSS a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X348 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X349 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X350 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X351 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X352 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X353 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X354 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X355 hgu_inverter_1.VSS a_528_5873# hgu_cdac_8bit_array_3.drv<1:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X356 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X357 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X358 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X359 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X360 hgu_inverter_1.VSS a_1437_5881# hgu_cdac_8bit_array_3.drv<3:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X361 hgu_inverter_1.VSS a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X362 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X363 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X364 hgu_cdac_8bit_array_2.drv<15:0> a_8105_5185# inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X365 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X366 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X367 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X368 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X369 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X370 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X371 hgu_cdac_8bit_array_3.drv<15:0> a_5521_5720# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X372 hgu_inverter_1.VSS a_5521_5720# hgu_cdac_8bit_array_3.drv<15:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X373 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X374 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X375 hgu_inverter_1.VSS a_1921_5185# hgu_cdac_8bit_array_2.drv<3:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X376 hgu_cdac_8bit_array_2.drv<7:0> a_3540_5180# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X377 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X378 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X379 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X380 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X381 hgu_cdac_8bit_array_3.drv<15:0> a_5521_5720# inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X382 hgu_inverter_1.VSS a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X383 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X384 inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF a_3540_5180# hgu_cdac_8bit_array_2.drv<7:0> inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X385 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X386 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X387 hgu_inverter_1.VSS a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X388 hgu_inverter_1.VSS a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X389 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X390 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X391 inv_4_test_1/inv_2_test_1/x2.VREF a_1921_5185# hgu_cdac_8bit_array_2.drv<3:0> inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X392 hgu_cdac_8bit_array_3.drv<0> a_n249_5874# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.35
X393 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X394 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X395 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X396 hgu_cdac_8bit_array_3.drv<15:0> a_5521_5720# inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X397 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X398 hgu_cdac_8bit_array_2.drv<0> a_n271_5184# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.35
X399 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X400 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X401 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X402 hgu_inverter_1.VSS a_2970_5870# hgu_cdac_8bit_array_3.drv<7:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X403 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X404 hgu_inverter_1.VSS a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X405 hgu_inverter_1.VSS a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X406 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X407 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X408 hgu_inverter_1.VSS a_5521_5720# hgu_cdac_8bit_array_3.drv<15:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X409 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X410 hgu_cdac_8bit_array_3.drv<7:0> a_2970_5870# inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X411 hgu_inverter_1.VSS a_2970_5870# hgu_cdac_8bit_array_3.drv<7:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X412 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X413 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X414 hgu_inverter_1.VSS a_8105_5185# hgu_cdac_8bit_array_2.drv<15:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X415 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X416 hgu_cdac_8bit_array_2.drv<0> a_n271_5184# hgu_inverter_0.VREF hgu_inverter_0.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.35
X417 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X418 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X419 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X420 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X421 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X422 hgu_inverter_1.VSS a_5521_5720# hgu_cdac_8bit_array_3.drv<15:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X423 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X424 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X425 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X426 hgu_inverter_1.VSS a_8105_5185# hgu_cdac_8bit_array_2.drv<15:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X427 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X428 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X429 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X430 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X431 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_8105_5185# hgu_cdac_8bit_array_2.drv<15:0> inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X432 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X433 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X434 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X435 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X436 inv_2_test_1/x2.VREF a_528_5873# hgu_cdac_8bit_array_3.drv<1:0> inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X437 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X438 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X439 hgu_cdac_8bit_array_3.drv<0> a_n249_5874# hgu_inverter_1.VREF hgu_inverter_1.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.35
X440 hgu_inverter_1.VSS a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X441 hgu_cdac_8bit_array_3.drv<3:0> a_1437_5881# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X442 hgu_inverter_1.VSS a_3540_5180# hgu_cdac_8bit_array_2.drv<7:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X443 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X444 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_8105_5185# hgu_cdac_8bit_array_2.drv<15:0> inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X445 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X446 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X447 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X448 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X449 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X450 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X451 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X452 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X453 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X454 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X455 hgu_inverter_1.VSS a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X456 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X457 hgu_cdac_8bit_array_2.drv<15:0> a_8105_5185# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X458 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X459 hgu_cdac_8bit_array_3.drv<7:0> a_2970_5870# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X460 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X461 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X462 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X463 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X464 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X465 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X466 hgu_cdac_8bit_array_3.drv<15:0> a_5521_5720# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X467 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X468 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X469 hgu_cdac_8bit_array_2.drv<15:0> a_8105_5185# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X470 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X471 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X472 hgu_cdac_8bit_array_2.drv<15:0> a_8105_5185# inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X473 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X474 inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_2970_5870# hgu_cdac_8bit_array_3.drv<7:0> inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X475 hgu_cdac_8bit_array_3.drv<7:0> a_2970_5870# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X476 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_5521_5720# hgu_cdac_8bit_array_3.drv<15:0> inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X477 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X478 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X479 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X480 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X481 hgu_cdac_8bit_array_3.drv<15:0> a_5521_5720# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X482 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X483 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X484 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X485 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X486 hgu_cdac_8bit_array_3.drv<31:0> a_10713_5389# inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X487 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X488 inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_2970_5870# hgu_cdac_8bit_array_3.drv<7:0> inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X489 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X490 hgu_cdac_8bit_array_3.drv<15:0> a_5521_5720# inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X491 hgu_cdac_8bit_array_2.drv<15:0> a_8105_5185# inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X492 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X493 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X494 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X495 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X496 hgu_inverter_1.VSS a_20359_5189# hgu_cdac_8bit_array_2.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X497 hgu_inverter_1.VSS a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X498 hgu_cdac_8bit_array_2.drv<31:0> a_15263_5235# hgu_inverter_1.VSS hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X499 hgu_cdac_8bit_array_3.drv<63:0> a_29809_5455# inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X500 hgu_inverter_1.VSS a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X501 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X502 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X503 hgu_cdac_8bit_array_3.drv<3:0> a_1437_5881# inv_4_test_2/inv_2_test_1/x2.VREF inv_4_test_2/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X504 hgu_inverter_1.VSS a_15263_5235# hgu_cdac_8bit_array_2.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X505 hgu_cdac_8bit_array_2.drv<63:0> a_20359_5189# inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X506 hgu_inverter_1.VSS a_10713_5389# hgu_cdac_8bit_array_3.drv<31:0> hgu_inverter_1.VSS sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X507 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF a_29809_5455# hgu_cdac_8bit_array_3.drv<63:0> inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
.ends

