* NGSPICE file created from hgu_sarlogic_flat.ext - technology: sky130A

.subckt hgu_sarlogic_flat ready ext_clk sample_clk sample_clk_b sar_clk sel_bit[0]
+ sel_bit[1] sar_result[1] sar_result[2] sar_result[3] sar_result[6] sar_result[0]
+ sample_delay_cap_ctrl_code[2] sample_delay_cap_ctrl_code[1] sample_delay_cap_ctrl_code[0]
+ sample_delay_cap_ctrl_code[6] sample_delay_cap_ctrl_code[5] sample_delay_cap_ctrl_code[4]
+ sample_delay_cap_ctrl_code[3] sample_delay_cap_ctrl_code[11] sample_delay_cap_ctrl_code[15]
+ async_setb_delay_cap_ctrl_code[2] async_setb_delay_cap_ctrl_code[1] async_setb_delay_cap_ctrl_code[0]
+ async_resetb_delay_cap_ctrl_code[0] async_resetb_delay_cap_ctrl_code[1] async_resetb_delay_cap_ctrl_code[2]
+ async_setb_delay_cap_ctrl_code[3] async_delay_offset retimer_eob_delay_offset retimer_delay_code[2]
+ retimer_delay_code[1] vss_sw[7] vss_sw[6] vss_sw[5] vss_sw[4] vss_sw[3] vss_sw[2]
+ vss_sw[1] vdd_sw[7] vdd_sw[6] vdd_sw[5] vdd_sw[4] vdd_sw[3] vdd_sw[2] vdd_sw[1]
+ vss_sw_b[7] vss_sw_b[6] vss_sw_b[5] vss_sw_b[4] vdd_sw_b[1] vdd_sw_b[2] vdd_sw_b[3]
+ vdd_sw_b[4] vdd_sw_b[6] vdd_sw_b[7] sample_delay_cap_ctrl_code[9] sample_delay_cap_ctrl_code[14]
+ sample_delay_cap_ctrl_code[13] sample_delay_cap_ctrl_code[12] sample_delay_cap_ctrl_code[10]
+ comp_result retimer_delay_code[0] retimer_delay_code[3] vdd_sw_b[5] sar_result[4]
+ sar_result[5] sar_result[7] async_resetb_delay_cap_ctrl_code[3] vss_sw_b[1] vss_sw_b[2]
+ vss_sw_b[3] sample_delay_cap_ctrl_code[8] sample_delay_cap_ctrl_code[7] sample_delay_offset
+ VDD VSS
X0 a_9687_n656# a_9222_n964# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1 VSS a_13898_892# x4.x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_22178_5989# a_21713_5681# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X3 x4.x2.X a_9514_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_28443_2504# a_28162_2510# a_28350_2504# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X5 VDD VDD a_11141_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X6 a_15829_n1475# a_15925_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X7 a_21957_5989# a_21539_6073# a_21713_5681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X8 a_9990_n670# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X9 a_13898_892# x4.x30.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 VSS a_27006_1838# a_26941_1864# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X11 VDD a_21950_n670# a_21875_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X12 VSS a_27006_3758# a_26941_4162# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X13 a_15944_n938# a_15778_n938# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_16455_4992# a_17010_4992# a_16968_5300# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X15 x3.x5.X a_11801_6580# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_19700_3246# x4.D[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VDD a_12261_8772# a_11883_8462# VDD sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X18 vdd_sw_b[1] a_24342_n670# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X19 a_10549_8788# a_10817_8528# a_10763_8554# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X20 a_26737_2826# a_26225_2478# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X21 VDD retimer_eob_delay_offset x5.x2.x6.SW VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X22 a_15433_4145# x3.x77.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 x2.x2.x3.IN x2.x2.x2.x9.output_stack a_19961_8655# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X24 a_30402_5732# x5.x2.x9.output_stack x5.x3.A VSS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X25 a_14860_n1443# a_14387_n1353# a_15104_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X26 x3.x4.X a_11974_5018# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_28350_3144# x4.D[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X28 a_15433_4145# a_14830_4119# a_15317_4119# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X29 x1.x4.x9.output_stack async_resetb_delay_cap_ctrl_code[2] x1.x4.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X30 a_15334_3554# a_14375_3272# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X31 a_11075_11958# a_10909_11958# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X32 a_23484_n572# a_23120_n938# a_23400_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X33 a_26051_2230# a_25770_1864# a_25958_1864# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X34 vdd_sw_b[6] a_12382_n670# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X35 VDD a_16928_4119# a_16838_4511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X36 a_14250_n656# a_13832_n572# a_14006_n964# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X37 a_9938_n938# a_8768_n938# a_9831_n572# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X38 a_16398_n964# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X39 a_22290_n250# a_22036_77# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X40 VSS a_9514_892# x4.x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X41 a_10004_8554# a_9804_8920# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X42 a_21752_5300# a_21552_5018# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X43 a_26051_9043# x2.x2.x2.IN a_25979_9181# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X44 a_21538_4511# a_21257_4145# a_21445_4145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X45 x3.x4.X a_11974_5018# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X46 a_19053_4145# x3.x7.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X47 a_21512_n1261# a_20709_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X48 VDD a_23003_n98# x4.x18.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X49 a_14917_4992# x3.x5.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X50 a_8956_n938# x4.x5.D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X51 VDD a_10957_7987# x1.x3.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X52 VSS VDD a_20041_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X53 a_11524_n572# a_11160_n938# a_11440_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X54 a_26365_2870# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X55 VSS x3.D[0] a_18699_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X56 VDD x5.x3.X a_27996_3790# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X57 a_13577_n250# x4.x11.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X58 a_18752_4992# a_18847_4992# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X59 a_23818_n656# a_23400_n572# a_23574_n964# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X60 VSS a_15317_4119# a_16024_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X61 x1.x10.Y x1.x10.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X62 a_19159_3272# x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X63 x5.x1[4].Q_N a_27006_2478# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X64 a_24664_5133# x5.eob a_24592_5133# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X65 a_27240_2146# a_26832_1864# a_27006_1838# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X66 a_18934_n938# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X67 a_9552_n1261# a_8749_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X68 a_22036_n1443# a_21563_n1353# a_22280_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X69 a_26386_12029# x2.x2.x1.x9.output_stack x2.x2.x2.IN VSS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X70 a_3051_11231# ready a_2979_11231# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X71 a_19636_5384# a_18847_4992# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X72 VSS a_13898_892# x4.x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X73 a_10332_77# VSS a_10332_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X74 a_18336_n938# a_18170_n938# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X75 a_19321_5681# a_19147_6073# a_19461_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X76 a_19838_5384# a_19701_4992# a_19402_4992# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X77 a_27122_3144# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X78 VDD a_27006_3758# a_27713_3800# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X79 a_21852_4145# x3.x39.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X80 VDD a_18317_n1653# vss_sw_b[3] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X81 a_27122_3144# a_26519_3118# a_27006_3118# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X82 a_23120_n938# a_22954_n938# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X83 x3.x4.X a_11974_5018# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X84 a_23145_77# x4.x20.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X85 a_15335_n250# x4.x9.A1 a_15114_77# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X86 a_22224_4145# a_21712_4119# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X87 a_12942_3554# a_11983_3272# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X88 a_19255_5707# a_18866_5707# a_19147_6073# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X89 x4.x9.A1 a_13898_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X90 a_2979_9193# sar_clk a_2891_9055# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X91 a_21768_n1653# a_22036_n1443# a_21982_n1345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X92 VSS VDD a_11263_8932# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X93 a_21713_5681# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X94 VSS x4.x30.A a_13898_892# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X95 a_9514_892# x4.x3.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X96 a_23366_n250# VSS a_23003_n98# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X97 a_22231_3272# a_22091_3546# a_21793_3246# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X98 a_12545_11952# a_12137_12330# a_12311_11926# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X99 a_16661_4145# x3.x7.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X100 a_15042_77# a_14860_77# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X101 x1.x4.x4[3].floating async_resetb_delay_cap_ctrl_code[2] x1.x4.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X102 a_23308_n938# x4.D[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X103 x3.x4.A a_11360_5018# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X104 a_10272_7835# x5.eob VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X105 a_26469_2504# a_26051_2504# a_26225_2478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X106 a_26051_9319# x2.x2.x2.IN a_25979_9457# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X107 a_18025_5384# a_17513_4992# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X108 a_28551_2882# a_28162_2510# a_28443_2504# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X109 VDD VDD a_26519_1838# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X110 VDD x5.x3.X a_25604_3790# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X111 a_14081_4145# a_13915_4145# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X112 a_16873_3272# a_17009_3246# a_16454_3246# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X113 VSS x4.x15.S a_20121_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X114 a_9080_n276# x4.x7.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X115 VDD a_11883_7842# sample_clk_b VDD sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X116 a_11406_n250# VSS a_11043_n98# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X117 a_26225_3758# a_26051_3784# a_26365_4150# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X118 x4.x3.A a_8604_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X119 a_11099_7835# sample_clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X120 VDD a_16360_4992# x4.x20.S VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X121 a_24070_n1627# a_23955_n1353# a_23647_n1459# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X122 a_16767_3272# x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X123 x2.x2.x2.x6.SW sample_delay_offset VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X124 a_22493_4119# a_22319_4145# a_22609_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X125 VSS a_19320_4119# a_19254_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X126 sample_clk a_11883_8462# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X127 VDD a_8653_n1475# vss_sw[7] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X128 VDD a_28911_1838# a_29632_2146# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X129 a_17441_5707# a_16929_5681# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X130 a_19302_n938# a_18790_n964# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X131 a_12330_n938# a_11160_n938# a_12223_n572# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X132 a_28757_3144# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X133 a_10280_8554# a_9491_8544# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X134 a_20709_n1653# a_21022_n1627# a_21128_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X135 x4.x17.X a_22290_77# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X136 a_15121_4992# a_15389_5202# a_15335_5300# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X137 a_10482_8554# a_10345_8772# a_10046_8528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X138 a_15944_n938# a_15778_n938# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X139 VDD a_14774_n670# a_15495_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X140 VSS a_27006_2478# a_27713_2520# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X141 a_15053_3638# a_14916_3246# a_14617_3246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X142 a_24664_5409# x5.eob a_24592_5409# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X143 x3.x4.X a_11974_5018# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X144 a_29129_3144# a_28617_3118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X145 VSS x4.D[4] a_17697_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X146 a_12223_11952# a_11075_11958# a_12137_12330# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X147 a_11974_5018# x3.x4.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X148 a_10521_n1627# a_9604_n1653# a_10076_n1443# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X149 a_19317_7792# x2.x2.x3.IN a_19229_7654# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X150 x3.x75.Q a_16024_4145# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X151 x1.x2.x9.output_stack ready a_2979_11507# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X152 VSS a_19558_n670# a_20279_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X153 VDD a_17710_5681# a_17622_6073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X154 VSS a_9491_8544# x1.x27.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X155 a_16863_5707# a_16474_5707# a_16755_6073# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X156 a_18724_n938# a_18170_n938# a_18616_n572# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X157 a_29224_2882# a_28162_2510# a_29129_2826# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X158 a_13252_8858# x2.x7.A VDD VSS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X159 VDD a_16929_5681# a_16839_6073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X160 a_29310_2504# a_28162_2510# a_29224_2882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X161 x3.x30.Q_N a_17710_5681# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X162 a_17010_4992# a_17308_5292# a_17244_5384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X163 a_21898_n938# a_20728_n938# a_21791_n572# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X164 VSS a_14006_n964# a_13940_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X165 sar_result[3] a_30105_3144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X166 a_21539_6073# a_21258_5707# a_21446_5707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X167 x5.x1[7].Q_N a_29398_1838# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X168 a_8749_n1653# a_9062_n1627# a_9168_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X169 a_13832_n572# a_13386_n938# a_13740_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X170 a_20974_n250# VSS a_20611_n98# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X171 a_24612_77# a_24430_77# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X172 a_17535_4145# a_16473_4145# a_17440_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X173 VSS a_18648_n276# a_18582_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X174 VSS a_22296_3246# a_22231_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X175 x2.x7.A x2.x2.x3.x9.output_stack a_13252_8655# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X176 x4.x9.A1 a_13898_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X177 x4.x20.X a_24684_77# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X178 x3.x75.Q_N a_15317_4119# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X179 a_20601_13233# x2.x2.x1.IN a_20513_13095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X180 a_2979_9469# sar_clk a_2891_9331# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X181 a_20916_n938# x4.D[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X182 a_9110_77# x4.x9.A1 a_8651_n98# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X183 a_17710_5681# a_17536_5707# a_17826_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X184 VDD a_26519_3118# a_27240_3426# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X185 VDD a_11530_11926# a_11440_11952# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X186 a_14481_3272# a_14617_3246# a_14062_3246# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X187 VSS a_24342_n670# a_24290_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X188 a_24374_n1345# a_23414_n1627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X189 a_28551_3144# a_28162_3144# a_28443_3510# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X190 a_13846_n1627# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X191 VSS x3.x4.X a_19614_4119# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X192 a_19342_9043# x2.x2.x3.IN a_19270_9181# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X193 x2.x2.x2.x5[7].floating x2.x2.x2.x10.Y x2.x2.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X194 VDD x2.x3.Y a_12261_8772# VDD sky130_fd_pr__pfet_01v8 ad=0.406 pd=3.38 as=0.406 ps=3.38 w=1.4 l=0.15
X195 a_3004_7942# sar_clk a_2916_7804# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X196 VDD a_27006_1838# a_27713_1864# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X197 a_23400_n572# a_23120_n938# a_23308_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X198 a_10130_7987# x1.x3.X a_10272_8162# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X199 a_8789_11554# x1.x9.A VDD VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X200 a_19270_9871# x2.x2.x3.IN a_19182_9733# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X201 a_22405_4511# a_21257_4145# a_22319_4145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X202 VSS x4.D[1] a_24873_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X203 a_16910_n938# a_16398_n964# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X204 VSS a_12382_n670# a_12330_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X205 x3.x7.X a_11392_4144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X206 a_14081_4145# a_13915_4145# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X207 x5.x2.x9.output_stack x5.x2.x10.Y x5.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X208 a_9366_n938# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X209 a_29398_3118# a_29224_3144# a_29514_3144# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X210 a_19230_4511# a_18699_4145# a_19146_4511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X211 a_15317_4119# x3.x77.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X212 x3.x66.Q_N a_22493_4119# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X213 VDD a_11360_5018# x3.x4.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X214 a_12661_3638# a_12524_3246# a_12225_3246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X215 VDD x1.x9.Y a_9491_8544# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X216 a_11687_n1459# a_11996_n1653# a_11931_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X217 x4.x2.X a_9514_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X218 a_29398_3758# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X219 a_20172_3456# a_19699_3546# a_20416_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X220 a_26026_7516# x2.x2.x2.IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X221 a_19677_12029# x2.x2.x1.IN VDD VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X222 VDD VDD a_19376_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X223 a_25979_9595# x2.x2.x2.IN a_25891_9457# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X224 VSS x4.x17.S a_22036_77# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X225 a_28162_2510# a_27996_2510# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X226 VDD x3.x75.Q a_16307_4145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X227 a_13898_892# x4.x30.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X228 VDD VDD a_21239_4992# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X229 vdd_sw[3] a_20279_n938# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X230 a_13892_12957# x2.x3.A a_13804_12819# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X231 VDD a_10130_7987# sar_clk VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X232 a_10272_8162# x5.eob VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X233 a_20040_3272# a_20172_3456# a_19904_3246# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X234 a_21040_n276# x4.x17.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X235 a_14618_4992# a_14916_5292# a_14852_5384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X236 VSS a_11614_n964# a_11548_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X237 a_13867_11844# x2.x3.A a_13779_11844# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X238 a_29224_3144# a_28162_3144# a_29129_3144# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X239 a_22027_3638# a_21238_3246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X240 a_21904_n1627# a_22036_n1443# a_21768_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X241 a_11099_8162# sample_clk VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X242 a_11645_n1345# a_11454_n1627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X243 a_14615_n572# a_13386_n938# a_14518_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X244 a_17436_77# a_17254_77# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X245 VDD a_11974_5018# x3.x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X246 VDD a_8880_892# x4.x3.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X247 a_9491_8544# a_9804_8920# a_9910_8876# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X248 a_18821_n1345# a_18630_n1627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X249 VDD x2.x2.x1.IN a_20513_13371# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X250 VSS a_21950_n670# a_21898_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X251 a_13432_6946# a_13316_6554# a_13346_6580# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.16 as=0.0567 ps=0.69 w=0.42 l=0.15
X252 x5.x2.x5[7].floating x5.x2.x10.Y x5.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X253 VSS a_20709_n1653# vss_sw_b[2] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X254 x5.x3.X a_30706_5822# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X255 VDD VDD a_19084_n964# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X256 a_20172_3456# a_19700_3246# a_20416_3638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X257 a_22093_4992# x3.x5.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X258 a_21008_n572# a_20728_n938# a_20916_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X259 VDD a_15318_5681# a_16025_5707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X260 a_19342_9319# x2.x2.x3.IN a_19270_9457# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X261 a_19266_5018# a_19402_4992# a_18847_4992# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X262 a_22809_5018# a_22297_4992# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X263 a_17091_n572# a_15778_n938# a_17007_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X264 VSS a_13968_4992# x3.x48.Q VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X265 a_28617_1838# a_28443_2230# a_28757_1864# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X266 a_11670_3246# a_11983_3272# a_12089_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X267 VDD x4.x15.S a_20114_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X268 VDD a_12200_n1653# a_12133_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X269 VDD a_14062_3246# x3.x54.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X270 x3.x4.X a_11974_5018# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X271 a_22511_5300# a_21552_5018# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X272 VSS x3.x20.Q_N a_12089_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X273 x3.x69.Q_N a_20101_4119# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X274 a_15143_4145# a_13915_4145# a_15001_4427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X275 VSS x4.x11.S a_14860_77# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X276 VDD x3.x20.Q_N a_11670_3246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X277 VDD x4.x20.S a_14339_6946# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X278 a_18866_5707# a_18700_5707# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X279 VDD a_15317_4119# a_15229_4511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X280 a_28350_1864# x4.x5.D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X281 VSS x1.x10.A a_8789_8529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X282 x2.x2.x3.x6.SW sample_delay_offset VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X283 VSS a_8749_n1653# vss_sw_b[7] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X284 a_10546_77# VSS a_10332_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X285 x4.x27.A a_12988_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X286 a_16429_n1345# a_16238_n1627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X287 a_8793_77# x4.x7.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X288 a_28350_3784# x4.D[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X289 VDD VSS a_13915_4145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X290 a_25770_2510# a_25604_2510# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X291 a_16360_4992# a_16455_4992# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X292 VDD a_21768_n1653# a_21701_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X293 a_13836_6580# sel_bit[0] a_14134_6580# VSS sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0671 ps=0.75 w=0.36 l=0.15
X294 VSS a_11045_n1475# vss_sw[6] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X295 VDD VDD a_13533_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X296 a_18221_n1475# a_18317_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X297 x3.x4.A a_11360_5018# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X298 a_29224_1864# a_27996_1864# a_29082_2146# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X299 a_21551_3272# x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X300 x2.x2.x1.x9.output_stack x2.x2.x1.x10.Y x2.x2.x1.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X301 VDD a_29398_1838# a_29310_2230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X302 a_25958_1864# x4.D[6] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X303 a_19558_n670# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X304 x3.x27.Q_N a_15318_5681# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X305 a_22481_n1627# a_21563_n1353# a_22036_n1443# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X306 VDD x4.x17.S a_22036_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X307 VDD x3.x36.Q_N a_21238_3246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X308 VDD a_18847_4992# x3.x42.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X309 VSS x3.x75.Q a_16307_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X310 VSS a_19905_4992# a_19840_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X311 a_8651_n98# x4.x9.A1 a_8793_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X312 VDD x5.x3.X a_27996_2510# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X313 a_22207_n656# a_21791_n572# a_21950_n670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X314 VDD VDD a_23101_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X315 VSS a_20613_n1475# vss_sw[2] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X316 a_14617_3246# a_14915_3546# a_14851_3638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X317 a_18866_5707# a_18700_5707# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X318 x5.x2.x9.output_stack retimer_delay_code[2] x5.x2.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X319 a_14592_n1653# a_14860_n1443# a_14806_n1345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X320 vdd_sw_b[4] a_17166_n670# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X321 VDD a_9514_892# x4.x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X322 VDD sar_clk a_12988_892# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X323 VSS x3.x36.Q_N a_21657_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X324 a_26918_3510# a_25770_3144# a_26832_3144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X325 a_13346_6580# a_13316_6554# a_13251_6580# VSS sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.066 ps=0.745 w=0.36 l=0.15
X326 a_26737_1864# a_26225_1838# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X327 a_19785_4427# a_19320_4119# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X328 a_13836_6580# a_13316_6554# a_14111_6878# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.164 ps=1.33 w=0.42 l=0.15
X329 a_10076_n1443# a_9604_n1653# a_10320_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X330 a_12468_n1443# a_11995_n1353# a_12712_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X331 a_3004_12482# ready a_2916_12344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X332 VDD a_28617_1838# a_28527_2230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X333 a_13939_11706# x2.x3.A a_13867_11844# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X334 a_19701_4992# x3.x5.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X335 a_24684_n250# a_24430_77# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X336 a_13042_5707# x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X337 VDD a_12926_5681# a_13633_5707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X338 a_22406_6073# a_21258_5707# a_22320_5707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X339 x3.x4.X a_11974_5018# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X340 VSS x4.x18.X a_22954_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X341 a_17496_n1627# a_16984_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X342 x5.x1[2].Q_N a_27006_3118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X343 VDD x3.x4.X a_17222_4119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X344 x2.x2.x2.x9.output_stack sample_delay_cap_ctrl_code[9] x2.x2.x2.x3[1].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X345 VDD a_21143_3246# x4.D[3] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X346 a_19786_5989# a_19321_5681# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X347 a_13042_5707# a_12439_5681# a_12926_5681# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X348 a_11454_n1627# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X349 a_15318_5681# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X350 a_19231_6073# a_18700_5707# a_19147_6073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X351 a_21326_n938# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X352 a_16929_5681# a_16755_6073# a_17069_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X353 sar_result[1] a_30105_3800# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X354 VDD x3.x5.A a_11801_6580# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X355 a_12852_6554# a_13721_6554# a_13346_6580# VSS sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X356 VDD x2.x1.x4.Y a_11824_12152# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X357 a_3051_9745# sar_clk a_2979_9745# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X358 x2.x2.x3.x5[7].floating x2.x2.x3.x10.Y x2.x2.x3.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X359 VSS a_11883_7842# sample_clk_b VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X360 a_18317_n1653# a_18863_n1459# a_18821_n1345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X361 a_12724_n250# a_12470_77# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X362 a_19317_8068# x2.x2.x3.IN a_19229_7930# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X363 a_26832_4162# a_25604_3790# a_26690_3784# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X364 VSS x2.x2.x2.IN a_26386_12370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X365 VSS x4.x8.X a_10994_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X366 x4.x9.A1 a_13898_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X367 a_22093_4992# x3.x5.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X368 VDD a_14300_n964# a_15031_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X369 a_12200_n1653# a_12468_n1443# a_12414_n1345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X370 a_18790_n964# a_18616_n572# a_18934_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X371 a_17308_3246# x4.D[4] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X372 a_22290_77# x4.x9.A1 a_22218_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X373 a_15252_4145# a_13915_4145# a_15143_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X374 VSS x3.x5.X a_16308_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X375 a_19270_9043# x2.x2.x3.IN x2.x2.x3.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X376 a_10559_7809# x5.eob VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X377 a_14269_4145# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X378 a_8789_8870# x1.x4.x9.output_stack x1.x10.A VSS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X379 x5.x2.x9.output_stack retimer_eob_delay_offset x5.x2.x7.floating VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X380 a_22230_5384# a_22093_4992# a_21794_4992# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X381 VDD a_9514_892# x4.x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X382 a_19399_n572# a_18336_n938# a_19255_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X383 x4.x7.X a_10332_77# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X384 a_26159_2882# a_25770_2510# a_26051_2504# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X385 a_10817_8528# a_10344_8676# a_11061_8920# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X386 VDD a_16455_4992# x3.x45.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X387 VDD a_26225_3118# a_26135_3510# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X388 VSS VSS a_13915_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X389 VDD a_11974_5018# x3.x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X390 a_14860_n1443# a_14388_n1653# a_15104_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X391 VDD x5.x3.X a_25604_2510# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X392 a_2979_10541# ready a_2891_10541# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X393 a_14502_n1627# a_14387_n1353# a_14079_n1459# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X394 VSS VDD a_17649_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X395 x1.x4.x9.output_stack async_delay_offset x1.x4.x7.floating VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X396 a_26051_9871# x2.x2.x2.IN a_25979_9871# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X397 a_15633_5384# a_15121_4992# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X398 x2.x2.x1.x2.floating sample_delay_cap_ctrl_code[4] x2.x2.x1.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X399 x1.x4.x9.output_stack sar_clk a_2916_8080# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X400 a_14575_3554# a_14375_3272# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X401 a_24428_n1443# a_23956_n1653# a_24672_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X402 a_23003_n98# x4.x9.A1 a_23145_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X403 a_15049_5707# a_14537_5681# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X404 a_19900_77# VSS a_19900_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X405 VDD x3.x5.X a_16308_5707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X406 VDD a_28911_3984# a_28861_3784# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X407 a_13867_11016# x2.x3.A a_13779_11016# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X408 VSS x4.x16.X a_20562_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X409 VDD x3.x4.X a_14830_4119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X410 VDD a_23868_n964# a_24599_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X411 x1.x4.x10.Y async_resetb_delay_cap_ctrl_code[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X412 a_3004_12758# ready a_2916_12620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X413 x2.x2.x1.x4[3].floating sample_delay_cap_ctrl_code[6] x2.x2.x1.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X414 a_15144_5707# a_13916_5707# a_15002_5989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X415 a_14537_5681# a_14363_6073# a_14677_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X416 x2.x2.x1.x9.output_stack x2.x2.x1.x10.Y x2.x2.x1.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X417 VSS a_12852_6554# x5.eob VSS sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X418 x4.x9.S a_18417_5707# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X419 x2.x3.A a_13018_11968# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X420 VDD a_15318_5681# a_15230_6073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X421 VDD a_23574_n964# a_23484_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X422 a_18226_3272# a_17307_3546# a_17780_3456# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X423 a_20101_4119# a_19927_4145# a_20217_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X424 a_11043_n98# x4.x9.A1 a_11185_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X425 a_26832_1864# a_25770_1864# a_26737_1864# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X426 a_18846_3246# a_19401_3246# a_19359_3554# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X427 a_19701_4992# x3.x5.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X428 VDD a_11908_n964# a_12639_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X429 VDD a_17222_4119# a_17172_4427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X430 a_14270_5707# x3.x27.D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X431 VDD a_11883_8462# sample_clk VDD sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X432 x3.x7.A a_11116_4144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X433 VSS a_22494_5681# a_23201_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X434 VSS a_18219_n98# x4.x14.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X435 sar_result[7] a_30105_1864# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X436 a_21257_4145# a_21091_4145# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X437 VDD a_17223_5681# a_17173_5989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X438 a_11670_12318# a_11824_12152# a_11530_11926# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X439 a_11974_5018# x3.x4.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X440 a_26225_3118# a_26051_3510# a_26365_3144# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X441 a_17007_n572# a_15944_n938# a_16863_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X442 a_21678_n1627# a_21563_n1353# a_21255_n1459# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X443 a_16332_n938# a_15778_n938# a_16224_n572# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X444 a_19270_9319# x2.x2.x3.IN a_19182_9181# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X445 a_14806_n1345# a_13846_n1627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X446 VDD x4.x20.S a_24430_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X447 VSS a_29398_2478# a_29333_2882# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X448 a_17166_n670# a_17007_n572# a_17306_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X449 a_25958_2504# x4.D[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X450 a_26159_3144# a_25770_3144# a_26051_3510# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X451 VSS a_13898_892# x4.x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X452 x3.x77.Y x5.eob VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X453 a_18630_n1627# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X454 x1.x2.x10.Y async_setb_delay_cap_ctrl_code[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X455 a_2979_9883# sar_clk a_2891_9883# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X456 a_14362_4511# a_13915_4145# a_14269_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X457 VDD a_8880_892# x4.x3.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X458 x4.x2.X a_9514_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X459 x4.D[2] a_23200_4145# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X460 a_11530_11926# x2.x1.x3.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X461 VSS a_21040_n276# a_20974_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X462 VSS a_14536_4119# a_14470_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X463 a_2979_10817# ready a_2891_10817# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X464 VSS x4.x13.S a_17729_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X465 a_12657_5707# a_12145_5681# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X466 a_14518_n938# a_14006_n964# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X467 a_22481_n1627# a_21564_n1653# a_22036_n1443# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X468 x5.x2.x10.Y retimer_delay_code[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X469 VDD x4.x18.X a_22954_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X470 VSS x4.x17.S a_22511_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X471 a_12752_5707# a_11524_5707# a_12610_5989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X472 x2.x2.x3.x3[1].floating sample_delay_cap_ctrl_code[13] x2.x2.x3.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X473 a_29398_2478# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X474 VSS a_28617_2478# a_28551_2882# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X475 a_16471_n1459# a_16780_n1653# a_16715_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X476 a_10559_7809# x5.eob VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X477 VDD a_12926_5681# a_12838_6073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X478 a_9366_n938# a_9516_n964# a_9222_n964# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X479 VSS async_delay_offset x1.x2.x6.SW VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X480 VDD x3.x4.X a_17223_5681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X481 VDD a_9990_n670# a_9915_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X482 VSS a_9990_n670# a_9938_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X483 x2.x1.x4.Y VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X484 a_15144_5707# a_14082_5707# a_15049_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X485 a_20416_3638# a_19904_3246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X486 VDD x4.x20.S a_15835_5018# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X487 VSS x5.x3.X a_27996_1864# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X488 VDD a_14830_4119# a_14780_4427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X489 a_16238_n1627# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X490 VDD x4.x8.X a_10994_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X491 x2.x2.x3.x9.output_stack sample_delay_cap_ctrl_code[13] x2.x2.x3.x3[1].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X492 VDD a_12261_7986# a_11883_7842# VDD sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X493 x3.x20.Q_N a_12926_5681# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X494 VSS a_8880_892# x4.x3.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X495 VDD a_19084_n964# a_19034_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X496 VSS x5.x3.X a_27996_3790# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X497 a_19961_8655# x2.x2.x3.IN VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X498 VSS a_20102_5681# a_20809_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X499 a_12336_n1627# a_12468_n1443# a_12200_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X500 VSS a_15827_n98# x4.x12.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X501 a_23010_3272# a_22092_3246# a_22564_3456# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X502 a_26026_7792# x2.x2.x2.IN a_25938_7930# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X503 a_19888_n1261# a_19376_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X504 a_27122_2870# a_26519_2704# a_27006_2478# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X505 VSS x2.x3.A a_13867_11016# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X506 VDD a_14831_5681# a_14781_5989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X507 a_22027_3272# a_21238_3246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X508 a_19053_4145# x3.x7.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X509 a_20089_n1627# a_19172_n1653# a_19644_n1443# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X510 VDD a_8651_n98# x4.x6.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X511 a_24684_77# x4.x9.A1 a_24612_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X512 VSS VDD a_14300_n964# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X513 a_8653_n1475# a_8749_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X514 a_13940_n938# a_13386_n938# a_13832_n572# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X515 sar_result[2] a_27713_3144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X516 a_27006_1838# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X517 a_22232_5018# a_22092_5292# a_21794_4992# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X518 a_14079_n1459# a_14388_n1653# a_14323_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X519 VDD a_9080_n276# a_9110_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X520 VDD x3.x7.X a_23010_3272# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X521 VDD a_11392_4144# x3.x7.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X522 a_21257_4145# a_21091_4145# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X523 x2.x2.x4.x9.output_stack sample_delay_cap_ctrl_code[1] x2.x2.x4.x3[1].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X524 a_14774_n670# a_14615_n572# a_14914_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X525 VSS x4.x20.S a_24430_77# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X526 x4.x9.A1 a_13898_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X527 x2.x2.x1.x4[3].floating sample_delay_cap_ctrl_code[6] x2.x2.x1.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X528 x3.x4.X a_11974_5018# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X529 x3.x3.A a_11084_5018# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X530 VDD x5.x3.X a_27996_1864# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X531 a_19399_n572# a_18170_n938# a_19302_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X532 a_17306_n938# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X533 x4.D[1] a_20808_4145# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X534 x2.x2.x2.x7.floating sample_delay_offset x2.x2.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X535 a_24617_6936# x5.eob a_24529_7074# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X536 a_13836_6580# sel_bit[1] a_12852_6554# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X537 a_23647_n1459# a_23956_n1653# a_23891_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X538 VSS a_13898_892# x4.x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X539 x1.x2.x9.output_stack x1.x2.x10.Y x1.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X540 VDD x4.x3.X a_9514_892# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X541 a_14446_4511# a_13915_4145# a_14362_4511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X542 a_20119_5300# a_19160_5018# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X543 VDD a_16984_n1653# a_16917_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X544 VDD x4.x16.X a_20562_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X545 VDD VDD a_28911_3984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X546 VDD x2.x2.x2.x9.output_stack a_19961_8655# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X547 a_16768_5018# x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X548 a_14037_n1345# a_13846_n1627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X549 a_15114_77# x4.x9.A1 a_15042_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X550 VDD x2.x2.x3.IN a_19961_8858# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X551 a_30402_5732# x5.x2.x9.output_stack VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X552 VDD a_19558_n670# a_19483_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X553 x2.x2.x2.x9.output_stack x2.x2.x2.x10.Y x2.x2.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X554 x2.x2.x4.x2.floating sample_delay_cap_ctrl_code[0] x2.x2.x4.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X555 a_20013_4511# a_18865_4145# a_19927_4145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X556 a_21853_5707# a_22007_5681# a_21713_5681# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X557 a_19342_9871# x2.x2.x3.IN a_19270_9871# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X558 VDD x3.x4.X a_14831_5681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X559 VDD x3.x27.Q_N a_15120_3246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X560 x2.x2.x4.x9.output_stack x2.x2.x4.x10.Y x2.x2.x4.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X561 VSS a_10559_7809# a_10493_7835# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X562 a_12752_5707# a_11690_5707# a_12657_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X563 VSS VDD a_23868_n964# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X564 a_28527_2230# a_27996_1864# a_28443_2230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X565 VSS x5.x3.X a_25604_1864# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X566 VSS a_23101_n1653# vss_sw_b[1] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X567 a_11043_n98# VSS a_11185_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X568 a_29129_2826# a_28617_2478# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X569 a_26225_3758# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X570 VDD a_9514_892# x4.x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X571 a_26051_9043# x2.x2.x2.IN a_25979_9043# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X572 VDD async_delay_offset x1.x4.x6.SW VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X573 VDD a_16692_n964# a_16642_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X574 VSS x5.x3.X a_25604_3790# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X575 a_12913_n1627# a_11995_n1353# a_12468_n1443# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X576 a_12427_12318# a_11824_12152# a_12311_11926# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X577 a_29333_4162# a_27996_3790# a_29224_4162# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X578 a_16661_4145# x3.x7.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X579 VDD a_10345_8772# a_10344_8676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X580 a_17648_3272# a_17780_3456# a_17512_3246# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X581 VSS VDD a_11908_n964# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X582 a_27240_3784# a_26832_4162# a_27006_3758# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X583 x4.x9.A1 a_13898_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X584 x5.x2.x9.output_stack retimer_delay_code[1] x5.x2.x3[1].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X585 a_24267_n572# a_22954_n938# a_24183_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X586 vdd_sw_b[5] a_14774_n670# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X587 a_19677_12370# x2.x2.x4.x9.output_stack VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X588 VSS a_22297_4992# a_22232_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X589 VDD x3.x7.X a_20618_3272# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X590 VDD a_27006_1838# a_26918_2230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X591 VDD a_21238_3246# x3.x63.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X592 VDD a_11974_5018# x3.x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X593 VDD a_29398_2478# a_30105_2520# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X594 a_14592_n1653# a_13846_n1627# a_14728_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X595 VDD x5.x3.X a_25604_1864# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X596 a_14914_n938# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X597 a_17252_n1443# a_16779_n1353# a_17496_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X598 VDD a_24160_n1653# a_24093_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X599 a_21950_n670# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X600 VDD a_12311_11926# a_13018_11968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X601 VDD a_19320_4119# a_19230_4511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X602 a_26386_12029# x2.x2.x1.x9.output_stack VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X603 a_14482_5018# a_14618_4992# a_14063_4992# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X604 a_12307_n572# a_10994_n938# a_12223_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X605 a_16238_n1627# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X606 a_12938_77# VSS a_12724_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X607 VDD VDD a_16692_n964# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X608 sar_result[5] a_30105_2520# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X609 VDD x3.x3.A a_11360_5018# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X610 VSS a_18846_3246# x3.x60.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X611 a_26386_12370# x2.x2.x2.IN VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X612 a_26832_2882# a_25604_2510# a_26690_2504# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X613 a_21326_n938# a_21476_n964# a_21182_n964# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X614 VSS a_23005_n1475# vss_sw[1] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X615 a_23904_n1261# a_23101_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X616 a_16984_n1653# a_17252_n1443# a_17198_n1345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X617 x3.x7.A a_11116_4144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X618 a_29398_2478# a_29224_2882# a_29514_2870# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X619 a_2979_9055# sar_clk a_2891_9055# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X620 x1.x4.x9.output_stack x1.x4.x6.SW x1.x4.x6.floating VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X621 a_12200_n1653# a_11454_n1627# a_12336_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X622 a_21128_n1627# a_21255_n1459# a_20709_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X623 a_13892_13233# x2.x3.A a_13804_13371# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X624 a_20173_5202# a_19700_5292# a_20417_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X625 a_26051_3784# a_25770_3790# a_25958_3784# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X626 vdd_sw_b[1] a_24342_n670# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X627 VSS a_14916_3246# a_14915_3546# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X628 a_26941_4162# a_25604_3790# a_26832_4162# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X629 VSS a_10957_7987# x1.x3.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X630 a_10332_n250# a_10078_77# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X631 a_19054_5707# x4.x9.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X632 a_26051_2230# a_25604_1864# a_25958_1864# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X633 x5.x1[5].Q_N a_29398_2478# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X634 a_11061_8920# a_10549_8788# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X635 a_26051_9319# x2.x2.x2.IN a_25979_9319# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X636 a_16968_5300# a_16768_5018# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X637 a_20041_5018# a_20173_5202# a_19905_4992# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X638 VSS a_26225_1838# a_26159_1864# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X639 VDD a_28911_3984# a_29632_3784# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X640 a_21768_n1653# a_21022_n1627# a_21904_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X641 a_29514_2870# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X642 x5.eob a_12852_6554# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X643 VSS a_26225_3758# a_26159_4162# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X644 a_21875_n572# a_20562_n938# a_21791_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X645 vdd_sw_b[6] a_12382_n670# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X646 x1.x2.x9.output_stack x1.x2.x10.Y x1.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X647 a_24428_n1443# a_23955_n1353# a_24672_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X648 x3.x5.X a_11801_6580# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X649 a_9014_n250# VSS a_8651_n98# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X650 a_9168_n1627# a_9295_n1459# a_8749_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X651 a_28443_3784# a_27996_3790# a_28350_3784# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X652 VDD sample_delay_cap_ctrl_code[11] x2.x2.x2.x10.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X653 x3.x5.A a_11525_6580# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X654 a_19815_n656# a_19399_n572# a_19558_n670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X655 a_22090_n938# a_21476_n964# a_21950_n670# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X656 a_28617_3118# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X657 a_19320_4119# a_19146_4511# a_19460_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X658 a_19828_77# a_19646_77# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X659 VSS a_19171_n1353# a_19172_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X660 VDD a_28911_2704# a_28861_2504# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X661 x2.x2.x2.x9.output_stack x2.x2.x2.x10.Y x2.x2.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X662 VDD a_21476_n964# a_22207_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X663 x2.x2.x4.x9.output_stack x2.x2.x4.x10.Y x2.x2.x4.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X664 x2.x2.x1.x9.output_stack x2.x2.x1.x6.SW x2.x2.x1.x6.floating VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X665 x2.x2.x1.x10.Y sample_delay_cap_ctrl_code[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X666 a_25979_9181# x2.x2.x2.IN a_25891_9181# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X667 a_10589_8162# VSS a_10130_7987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X668 a_14447_6073# a_13916_5707# a_14363_6073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X669 a_19254_4145# a_18865_4145# a_19146_4511# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X670 x4.x9.X a_12724_77# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X671 a_13160_5989# a_12752_5707# a_12926_5681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X672 a_24160_n1653# a_24428_n1443# a_24374_n1345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X673 a_28757_4150# a_28911_3984# a_28617_3758# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X674 a_19461_5707# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X675 a_11045_n1475# a_11141_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X676 a_29082_3426# a_28617_3118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X677 VSS a_16454_3246# x3.x57.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X678 a_10130_n938# a_9516_n964# a_9990_n670# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X679 a_19317_7516# x2.x2.x3.IN a_19229_7654# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X680 a_20014_6073# a_18866_5707# a_19928_5707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X681 a_13898_892# x4.x30.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X682 a_28861_3426# a_28443_3510# a_28617_3118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X683 a_16454_3246# a_17009_3246# a_16967_3554# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X684 VDD a_18751_3246# x4.D[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X685 a_17508_77# x4.x9.A1 a_17436_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X686 a_19255_n656# a_18790_n964# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X687 a_13867_11430# x2.x3.A a_13779_11292# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X688 VDD a_9516_n964# a_10247_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X689 a_15827_n98# VSS a_15969_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X690 a_12145_5681# x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X691 a_8789_11895# x1.x2.x9.output_stack VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X692 sar_result[0] a_27713_3800# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X693 VSS sel_bit[1] a_13721_6554# VSS sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.113 ps=1.38 w=0.42 l=0.15
X694 a_14006_n964# a_13832_n572# a_14150_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X695 a_22727_4427# a_22319_4145# a_22493_4119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X696 VDD a_17309_4992# a_17308_5292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X697 a_12524_3246# x4.D[6] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X698 sample_clk a_11883_8462# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X699 VSS x3.x5.X a_11524_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X700 a_11263_8932# a_10344_8676# a_10817_8528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X701 VDD x2.x2.x3.x9.output_stack a_13252_8655# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X702 VSS a_12524_3246# a_12523_3546# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X703 VDD x2.x7.A a_13252_8858# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X704 a_26026_8068# x2.x2.x2.IN x2.x2.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X705 a_20611_n98# VSS a_20753_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X706 x2.x2.x3.x9.output_stack x2.x2.x3.x10.Y x2.x2.x3.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X707 a_16662_5707# x4.x7.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X708 a_22728_5989# a_22320_5707# a_22494_5681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X709 a_11502_77# x4.x9.A1 a_11043_n98# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X710 VDD x3.x7.A a_11392_4144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X711 a_23011_5018# a_22092_5292# a_22565_5202# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X712 a_24592_4995# x5.eob a_24504_4995# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X713 a_17447_3272# a_17307_3546# a_17009_3246# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X714 a_19590_n1345# a_18630_n1627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X715 a_13967_3246# a_14062_3246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X716 a_22429_5707# a_21092_5707# a_22320_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X717 VSS VDD a_28911_1838# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X718 VDD x3.x4.X a_22006_4119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X719 VDD a_17513_4992# a_17446_5384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X720 a_17440_4145# a_16928_4119# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X721 a_17781_5202# a_17309_4992# a_18025_5384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X722 a_23101_n1653# a_23414_n1627# a_23520_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X723 a_16224_n572# a_15778_n938# a_16132_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X724 VSS VDD a_28911_3984# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X725 a_19342_9043# x2.x2.x3.IN a_19270_9043# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X726 VSS a_11530_11926# a_11464_12330# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X727 a_3004_7666# sar_clk a_2916_7804# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X728 VDD x3.x4.A a_11974_5018# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X729 VDD a_15317_4119# a_16024_4145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X730 VDD x4.x3.X a_9514_892# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X731 a_12913_n1627# a_11996_n1653# a_12468_n1443# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X732 a_28443_3510# a_28162_3144# a_28350_3144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X733 a_19270_9733# x2.x2.x3.IN a_19182_9733# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X734 x2.x2.x3.x5[7].floating x2.x2.x3.x10.Y x2.x2.x3.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X735 VDD a_19321_5681# a_19231_6073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X736 VDD x3.x5.X a_11524_5707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X737 x3.x4.X a_11974_5018# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X738 a_21239_4992# a_21552_5018# a_21658_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X739 VDD a_14830_4119# a_15551_4427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X740 a_24290_n938# a_23120_n938# a_24183_n572# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X741 VSS a_27006_2478# a_26941_2882# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X742 x2.x2.x1.x9.output_stack sample_delay_cap_ctrl_code[6] x2.x2.x1.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X743 a_21446_5707# x4.x11.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X744 VSS VDD a_21658_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X745 a_16862_4145# a_16473_4145# a_16754_4511# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X746 VDD x2.x7.A x2.x7.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X747 x2.x2.x3.x4[3].floating sample_delay_cap_ctrl_code[14] x2.x2.x3.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X748 VDD a_14831_5681# a_15552_5989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X749 x3.x72.Q_N a_17709_4119# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X750 a_26690_3426# a_26225_3118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X751 x4.x30.A a_13264_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X752 a_14062_3246# a_14617_3246# a_14575_3554# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X753 a_25979_9457# x2.x2.x2.IN a_25891_9457# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X754 VDD a_13435_n98# x4.x10.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X755 x4.x2.X a_9514_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X756 a_17198_n1345# a_16238_n1627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X757 VDD a_9514_892# x4.x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X758 x5.eob a_12852_6554# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X759 a_16863_n656# a_16398_n964# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X760 x2.x2.x4.x9.output_stack x2.x3.A a_13804_12819# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X761 a_9491_8544# a_10046_8528# a_10004_8554# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X762 a_19160_5018# x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X763 a_20416_3272# a_19904_3246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X764 VSS a_11575_3246# x4.x5.D VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X765 VSS a_14774_n670# a_15495_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X766 a_11614_n964# a_11440_n572# a_11758_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X767 VSS a_13435_n98# x4.x10.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X768 a_17709_4119# a_17535_4145# a_17825_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X769 x1.x2.x9.output_stack x1.x2.x10.Y x1.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X770 VDD a_22092_3246# a_22091_3546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X771 a_20618_3272# a_19700_3246# a_20172_3456# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X772 a_13867_11706# x2.x3.A a_13779_11568# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X773 VSS x5.x3.A a_30706_5822# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X774 VDD x4.x17.S a_22504_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X775 a_11472_n276# x4.x9.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X776 VDD VDD a_18847_4992# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X777 a_13442_3272# a_12523_3546# a_12996_3456# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X778 a_2979_10021# sar_clk a_2891_9883# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X779 a_8789_8529# x1.x4.x9.output_stack x1.x10.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X780 VDD x4.x27.A a_13264_892# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X781 a_29632_3426# a_29224_3144# a_29398_3118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X782 a_11548_n938# a_10994_n938# a_11440_n572# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X783 x4.x3.X a_8880_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X784 sar_result[6] a_27713_1864# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X785 a_18865_4145# a_18699_4145# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X786 VDD a_11974_5018# x3.x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X787 a_13967_3246# a_14062_3246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X788 VDD VDD a_22297_4992# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X789 a_11575_3246# a_11670_3246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X790 vdd_sw[4] a_17887_n938# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X791 a_13939_11430# x2.x3.A a_13867_11430# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X792 VDD a_11801_6580# x3.x5.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X793 VSS a_12145_5681# a_12079_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X794 a_18863_n1459# a_19172_n1653# a_19107_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X795 VDD a_22296_3246# a_22229_3638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X796 VSS a_17309_4992# a_17308_5292# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X797 VSS x3.x7.X a_23010_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X798 a_30402_6073# x5.x2.x9.output_stack x5.x3.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X799 a_3051_10679# ready a_2979_10679# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X800 VSS x3.x4.X a_17223_5681# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X801 a_15389_5202# a_14917_4992# a_15633_5384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X802 VSS a_29398_3118# a_30105_3144# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X803 a_27006_3758# a_26832_4162# a_27122_4150# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X804 a_9132_n572# a_8768_n938# a_9048_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X805 VDD a_26519_1838# a_26469_2146# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X806 VSS VDD a_9944_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X807 a_19635_3638# a_18846_3246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X808 a_3051_9193# sar_clk a_2979_9331# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X809 a_19342_9319# x2.x2.x3.IN a_19270_9319# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X810 VDD a_12852_6554# x5.eob VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X811 VSS a_17512_3246# a_17447_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X812 a_19837_3638# a_19700_3246# a_19401_3246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X813 x2.x2.x1.x9.output_stack x2.x2.x1.x10.Y x2.x2.x1.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X814 VSS a_22494_5681# a_22429_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X815 a_12382_n670# a_12223_n572# a_12522_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X816 VDD a_19171_n1353# a_19172_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X817 a_18616_n572# a_18336_n938# a_18524_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X818 x5.x1[0].Q_N a_27006_3758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X819 VDD a_9514_892# x4.x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X820 a_17007_n572# a_15778_n938# a_16910_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X821 a_27122_1864# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X822 VSS x2.x2.x2.x9.output_stack a_19961_8858# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X823 VDD sample_delay_cap_ctrl_code[15] x2.x2.x3.x10.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X824 a_30402_5732# x5.x3.A VDD VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X825 a_27122_4150# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X826 x2.x2.x2.x9.output_stack sample_delay_cap_ctrl_code[10] x2.x2.x2.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X827 VSS a_10130_7987# sar_clk VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X828 a_27122_1864# a_26519_1838# a_27006_1838# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X829 a_24296_n1627# a_24428_n1443# a_24160_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X830 x2.x2.x4.x10.Y sample_delay_cap_ctrl_code[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X831 a_20576_11292# x2.x2.x1.IN a_20488_11292# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X832 a_16768_5018# x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X833 VSS x4.x7.S a_10078_77# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X834 a_26225_2478# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X835 a_15388_3456# a_14915_3546# a_15632_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X836 x1.x4.x9.output_stack x1.x4.x10.Y x1.x4.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X837 a_21539_6073# a_21092_5707# a_21446_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X838 a_9466_n656# a_9048_n572# a_9222_n964# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X839 a_12852_6554# sel_bit[1] a_13346_6580# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0729 pd=0.81 as=0.14 ps=1.6 w=0.54 l=0.15
X840 a_17722_77# VSS a_17508_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X841 VDD a_19700_3246# a_19699_3546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X842 a_17697_n1627# a_16779_n1353# a_17252_n1443# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X843 VSS a_21713_5681# a_21647_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X844 VSS a_23574_n964# a_23508_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X845 x4.x3.A a_8604_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X846 a_14134_6580# x3.x48.Q VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0819 ps=0.81 w=0.42 l=0.15
X847 a_14269_4145# VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X848 VDD a_11974_5018# x3.x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X849 a_18024_3638# a_17512_3246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X850 VDD VDD a_12439_5681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X851 VDD x3.x20.Q_N a_12728_3246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X852 VSS a_16360_4992# x4.x20.S VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X853 VSS a_15829_n1475# vss_sw[4] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X854 a_27240_2504# a_26832_2882# a_27006_2478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X855 x2.x2.x1.x9.output_stack sample_delay_cap_ctrl_code[6] x2.x2.x1.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X856 a_26135_2230# a_25604_1864# a_26051_2230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X857 a_11575_3246# a_11670_3246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X858 a_8789_11895# x1.x9.A VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X859 VDD a_14300_n964# a_14250_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X860 a_19904_3246# a_20172_3456# a_20118_3554# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X861 vdd_sw[5] a_15495_n938# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X862 x3.x5.A a_11525_6580# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X863 VSS x3.x7.X a_20618_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X864 a_10957_7987# x1.x3.A0 a_11099_8162# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X865 x5.x3.X a_30706_5822# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X866 VDD a_14592_n1653# a_14525_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X867 a_26225_2478# a_26051_2504# a_26365_2870# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X868 x1.x4.x5[7].floating x1.x4.x10.Y x1.x4.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X869 VSS x3.x4.X a_14831_5681# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X870 VDD x5.x3.A a_30706_5822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X871 x1.x2.x9.output_stack ready a_2916_12344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X872 a_13939_11706# x2.x3.A a_13867_11706# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X873 a_24617_6660# x5.eob a_24529_6522# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X874 a_19840_5018# a_19700_5292# a_19402_4992# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X875 a_18846_3246# a_19159_3272# a_19265_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X876 a_11974_5018# x3.x4.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X877 a_18865_4145# a_18699_4145# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X878 VDD x3.x4.X a_22007_5681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X879 a_15305_n1627# a_14387_n1353# a_14860_n1443# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X880 a_19120_n1261# a_18317_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X881 VSS x3.x33.Q_N a_19265_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X882 a_13898_892# x4.x30.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X883 a_28757_1864# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X884 a_2979_11231# ready a_2891_11093# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X885 VSS x4.x20.S a_14340_6580# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.066 ps=0.745 w=0.42 l=0.15
X886 a_28757_4150# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X887 a_28350_1864# x4.x5.D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X888 a_13251_6580# x4.x15.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.107 ps=1 w=0.42 l=0.15
X889 x3.x30.Q_N a_17710_5681# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X890 VSS a_13437_n1475# vss_sw[5] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X891 VDD VDD a_15925_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X892 VSS x3.x27.Q_N a_15256_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X893 a_3051_9469# sar_clk a_2979_9607# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X894 a_29129_1864# a_28617_1838# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X895 sar_result[3] a_30105_3144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X896 VDD a_20709_n1653# vss_sw_b[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X897 a_16256_n276# x4.x13.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X898 VSS VDD a_26519_3118# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X899 a_17727_5300# a_16768_5018# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X900 a_11560_n1627# a_11687_n1459# a_11141_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X901 VSS x4.x6.X a_8602_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X902 a_24873_n1627# a_23955_n1353# a_24428_n1443# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X903 a_17009_3246# a_17307_3546# a_17243_3638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X904 x3.x75.Q_N a_15317_4119# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X905 VDD a_9396_8528# x1.x3.A0 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X906 a_16984_n1653# a_16238_n1627# a_17120_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X907 a_26051_2504# a_25770_2510# a_25958_2504# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X908 a_19461_5707# a_19615_5681# a_19321_5681# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X909 VSS a_10345_8772# a_10344_8676# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X910 a_29310_3510# a_28162_3144# a_29224_3144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X911 a_20576_11568# x2.x2.x1.IN a_20488_11568# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X912 a_8749_n1653# a_9295_n1459# a_9253_n1345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X913 x2.x2.x2.x4[3].floating sample_delay_cap_ctrl_code[10] x2.x2.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X914 a_29224_4162# a_27996_3790# a_29082_3784# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X915 x1.x2.x9.output_stack x1.x2.x6.SW x1.x2.x6.floating VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X916 a_13552_n938# a_13386_n938# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X917 VDD a_28911_2704# a_29632_2504# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X918 a_16767_3272# x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X919 VDD a_29398_3758# a_29310_3784# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X920 a_25958_3784# x3.D[0] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X921 vdd_sw_b[2] a_21950_n670# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X922 VDD a_8749_n1653# vss_sw_b[7] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X923 a_12311_11926# a_12137_12330# a_12427_12318# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X924 a_12468_n1443# a_11996_n1653# a_12712_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X925 a_23011_5018# a_22093_4992# a_22565_5202# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X926 a_22028_5018# a_21239_4992# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X927 a_19888_n1627# a_19376_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X928 VDD a_11908_n964# a_11858_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X929 a_10320_n1261# a_9808_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X930 VDD x4.x3.X a_9514_892# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X931 a_20648_11154# x2.x2.x1.IN a_20576_11292# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X932 a_13898_892# x4.x30.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X933 VDD a_11045_n1475# vss_sw[6] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X934 a_13846_n1627# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X935 x4.x9.A1 a_13898_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X936 a_28551_1864# a_28162_1864# a_28443_2230# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X937 a_26051_9595# x2.x2.x2.IN a_25979_9733# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X938 VSS a_9603_n1353# a_9604_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X939 a_16928_4119# a_16754_4511# a_17068_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X940 VSS a_11360_5018# x3.x4.A VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X941 a_21701_n1261# a_21564_n1653# a_21255_n1459# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X942 x2.x2.x1.x9.output_stack sample_delay_offset x2.x2.x1.x7.floating VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X943 a_21092_n572# a_20728_n938# a_21008_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X944 a_16454_3246# a_16767_3272# a_16873_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X945 vdd_sw_b[7] a_9990_n670# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X946 VDD a_14536_4119# a_14446_4511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X947 a_14006_n964# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X948 VDD a_27006_2478# a_27713_2520# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X949 VDD a_28617_3758# a_28527_3784# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X950 x2.x2.x2.x9.output_stack sample_delay_cap_ctrl_code[10] x2.x2.x2.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X951 VDD a_20613_n1475# vss_sw[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X952 a_18524_n938# x4.D[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X953 a_23145_n250# x4.x20.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X954 a_26365_4150# a_26519_3984# a_26225_3758# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X955 a_24617_6936# x5.eob a_24529_6798# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X956 a_17069_5707# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X957 a_29398_1838# a_29224_1864# a_29514_1864# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X958 a_22609_4145# x3.x39.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X959 a_26469_3426# a_26051_3510# a_26225_3118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X960 x4.x9.X a_12724_77# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X961 VDD a_16359_3246# x4.D[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X962 VSS a_9080_n276# a_9014_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X963 VDD a_11392_4144# x3.x7.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X964 a_2979_11507# ready a_2891_11369# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X965 a_10484_8932# a_10344_8676# a_10046_8528# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X966 a_24160_n1653# a_23414_n1627# a_24296_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X967 sar_result[4] a_27713_2520# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X968 x5.x2.x4[3].floating retimer_delay_code[2] x5.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X969 a_9741_n1261# a_9604_n1653# a_9295_n1459# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X970 VDD x2.x7.Y x2.x3.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X971 VDD a_14917_4992# a_14916_5292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X972 a_16360_4992# a_16455_4992# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X973 a_11185_n250# x4.x9.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X974 a_21426_n656# a_21008_n572# a_21182_n964# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X975 a_17252_n1443# a_16780_n1653# a_17496_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X976 VSS a_11974_5018# x3.x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X977 a_9048_n572# a_8768_n938# a_8956_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X978 VDD x3.x4.A a_11974_5018# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X979 a_29224_1864# a_28162_1864# a_29129_1864# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X980 a_16894_n1627# a_16779_n1353# a_16471_n1459# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X981 VSS sample_delay_offset x2.x2.x4.x6.SW VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X982 a_22296_3246# a_21551_3272# a_22432_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X983 VSS x2.x2.x3.x9.output_stack a_13252_8858# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X984 a_16542_n938# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X985 x2.x2.x3.x9.output_stack sample_delay_cap_ctrl_code[14] x2.x2.x3.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X986 a_17244_5384# a_16455_4992# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X987 x1.x4.x9.output_stack async_resetb_delay_cap_ctrl_code[2] x1.x4.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X988 a_12758_8861# x2.x3.A x2.x3.Y VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X989 x4.x9.A1 a_13898_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X990 a_20335_4427# a_19927_4145# a_20101_4119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X991 VDD a_15121_4992# a_15054_5384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X992 a_17446_5384# a_17309_4992# a_17010_4992# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X993 a_15048_4145# a_14536_4119# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X994 a_2979_9745# sar_clk a_2891_9607# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X995 VSS x2.x3.Y a_12261_8772# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X996 a_20336_5989# a_19928_5707# a_20102_5681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X997 a_17649_5018# a_17781_5202# a_17513_4992# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X998 VSS a_11883_8462# sample_clk VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X999 VDD a_11801_6580# x3.x5.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1000 a_14536_4119# a_14362_4511# a_14676_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X1001 a_28757_3144# a_28911_3118# a_28617_3118# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1002 x3.D[0] a_18416_4145# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X1003 a_20648_11430# x2.x2.x1.IN a_20576_11568# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1004 a_20037_5707# a_18700_5707# a_19928_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X1005 a_22610_5707# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X1006 a_23005_n1475# a_23101_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1007 a_11614_n964# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X1008 a_15114_77# VSS a_15114_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1009 a_21239_4992# a_21794_4992# a_21752_5300# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X1010 a_18219_n98# VSS a_18361_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X1011 a_22610_5707# a_22007_5681# a_22494_5681# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1012 a_19698_n938# a_19084_n964# a_19558_n670# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1013 a_17729_n250# x4.x9.A1 a_17508_77# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X1014 VDD a_11883_7842# sample_clk_b VDD sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X1015 a_20753_n250# x4.x17.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X1016 a_14677_5707# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X1017 a_9062_n1627# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1018 a_18219_n98# x4.x9.A1 a_18361_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1019 VSS a_11670_3246# x3.x51.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1020 VDD a_13264_892# x4.x30.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1021 VSS a_22493_4119# a_23200_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1022 VDD a_19084_n964# a_19815_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X1023 VDD a_13967_3246# x4.D[6] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1024 a_11386_7809# sample_clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X1025 a_13894_77# x4.x9.A1 a_13435_n98# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X1026 a_28350_2504# x4.D[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1027 VDD a_11974_5018# x3.x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1028 VSS a_18847_4992# x3.x42.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1029 VDD x4.x6.X a_8602_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1030 a_21143_3246# a_21238_3246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1031 VDD a_12439_5681# a_13160_5989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X1032 VDD a_24342_n670# a_25063_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1033 VSS x4.x27.A a_13264_892# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1034 a_14375_3272# x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1035 a_15305_n1627# a_14388_n1653# a_14860_n1443# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X1036 a_25979_9871# x2.x2.x2.IN a_25891_9733# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1037 x2.x2.x2.x9.output_stack sample_delay_cap_ctrl_code[8] x2.x2.x2.x2.floating VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.43 as=0.122 ps=1.42 w=0.42 l=0.15
X1038 a_11878_5707# x5.eob VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X1039 VDD a_12311_11926# a_12223_11952# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X1040 VSS a_13533_n1653# vss_sw_b[5] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1041 VDD a_26519_1838# a_27240_2146# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X1042 VSS a_17710_5681# a_18417_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1043 a_26365_3144# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X1044 a_8789_11554# x1.x2.x9.output_stack x1.x9.A VSS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X1045 VDD a_11360_5018# x3.x4.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1046 VDD x4.x17.S a_18227_5018# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X1047 a_14852_5384# a_14063_4992# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X1048 VDD a_11472_n276# a_11502_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1049 a_13552_n938# a_13386_n938# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1050 VDD a_12382_n670# a_13103_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1051 VDD a_22006_4119# a_22727_4427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X1052 x1.x10.Y x1.x10.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1053 a_9396_8528# a_9491_8544# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1054 VSS a_14917_4992# a_14916_5292# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1055 a_26051_9871# x2.x2.x2.IN a_25979_10009# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1056 VDD VDD a_16455_4992# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X1057 a_24873_n1627# a_23956_n1653# a_24428_n1443# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X1058 a_19677_12029# x2.x2.x4.x9.output_stack x2.x2.x1.IN VSS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X1059 a_21255_n1459# a_21563_n1353# a_21512_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X1060 x2.x2.x3.x4[3].floating sample_delay_cap_ctrl_code[14] x2.x2.x3.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X1061 a_14471_5707# a_14082_5707# a_14363_6073# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X1062 VDD a_14537_5681# a_14447_6073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X1063 a_24664_4857# x5.eob a_24592_4995# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1064 a_19635_3272# a_18846_3246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X1065 x3.x3.A a_11084_5018# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1066 VDD a_9603_n1353# a_9604_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1067 a_9990_n670# a_9831_n572# a_10130_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X1068 x5.x1[6].Q_N a_27006_1838# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1069 a_11440_n572# a_10994_n938# a_11348_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X1070 VDD a_20611_n98# x4.x16.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X1071 a_15143_4145# a_14081_4145# a_15048_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X1072 VSS a_11141_n1653# vss_sw_b[6] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1073 VSS a_16256_n276# a_16190_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1074 a_22229_3638# a_22092_3246# a_21793_3246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X1075 VDD a_11974_5018# x3.x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1076 a_14728_n1627# a_14860_n1443# a_14592_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X1077 VSS a_20101_4119# a_20808_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1078 VDD a_30706_5822# x5.x3.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1079 VSS x4.x7.S a_10553_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X1080 a_15318_5681# a_15144_5707# a_15434_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X1081 a_19342_9595# x2.x2.x3.IN a_19270_9733# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1082 x4.x27.A a_12988_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1083 a_14376_5018# x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X1084 x1.x2.x2.floating async_setb_delay_cap_ctrl_code[0] x1.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X1085 a_9295_n1459# a_9603_n1353# a_9552_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X1086 VDD x4.D[3] a_20089_n1627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1087 VSS a_20102_5681# a_20037_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X1088 a_12089_3272# a_12225_3246# a_11670_3246# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X1089 VSS x1.x9.Y a_9910_8876# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X1090 VSS a_16455_4992# x3.x45.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1091 a_21143_3246# a_21238_3246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1092 x5.x2.x9.output_stack x5.x2.x6.SW x5.x2.x6.floating VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1093 VSS a_11974_5018# x3.x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1094 a_22297_4992# a_22565_5202# a_22511_5300# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X1095 VDD a_21950_n670# a_22671_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1096 x2.x2.x2.x9.output_stack x2.x2.x2.x10.Y x2.x2.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X1097 a_11995_n1353# x4.x9.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1098 a_11983_3272# x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1099 a_21008_n572# a_20562_n938# a_20916_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X1100 VSS x4.x30.A a_13898_892# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1101 x1.x2.x4[3].floating async_setb_delay_cap_ctrl_code[2] x1.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X1102 a_8789_8870# x1.x4.x9.output_stack VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1103 a_18024_3272# a_17512_3246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X1104 a_11263_11952# x2.x1.x2.D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X1105 x4.x9.A1 a_13898_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1106 a_12996_3456# a_12523_3546# a_13240_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X1107 a_27006_3118# a_26832_3144# a_27122_3144# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X1108 a_12137_12330# a_10909_11958# a_11995_11952# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X1109 a_19160_5018# x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1110 VDD a_9990_n670# a_10711_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1111 a_11774_11952# a_11356_11952# a_11530_11926# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X1112 x2.x2.x2.x6.SW sample_delay_offset VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1113 VDD VDD a_14063_4992# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X1114 VSS VDD a_21904_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X1115 a_27006_3758# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X1116 a_10260_77# a_10078_77# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1117 a_15632_3638# a_15120_3246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X1118 VDD a_19376_n1653# a_19309_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X1119 a_17448_5018# a_17308_5292# a_17010_4992# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X1120 a_28162_3144# a_27996_3144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1121 x4.x9.S a_18417_5707# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1122 a_8653_n1475# a_8749_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1123 VDD a_19904_3246# a_19837_3638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X1124 VSS a_12728_3246# a_12663_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X1125 a_11944_n1261# a_11141_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X1126 a_9915_n572# a_8602_n938# a_9831_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X1127 VSS a_9514_892# x4.x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1128 a_21852_4145# a_22006_4119# a_21712_4119# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1129 a_11386_7809# sample_clk VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1130 VSS a_27006_3118# a_27713_3144# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1131 VSS VDD a_12439_5681# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1132 VDD a_9491_8544# x1.x27.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X1133 VSS a_13864_n276# a_13798_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1134 VSS x1.x9.Y a_10685_8876# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X1135 VDD sample_delay_offset x2.x2.x1.x6.SW VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1136 a_12223_n572# a_10994_n938# a_12126_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X1137 x1.x4.x9.output_stack x1.x4.x10.Y x1.x4.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X1138 VSS a_18221_n1475# vss_sw[3] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1139 a_19320_4119# x3.x42.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X1140 x2.x2.x2.x5[7].floating x2.x2.x2.x10.Y x2.x2.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X1141 a_14339_6946# sel_bit[0] a_13836_6580# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0974 pd=0.97 as=0.0567 ps=0.69 w=0.42 l=0.15
X1142 VDD a_9514_892# x4.x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1143 a_10046_8528# a_10344_8676# a_10280_8554# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X1144 VSS x4.x15.S a_19646_77# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X1145 a_16344_n1627# a_16471_n1459# a_15925_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X1146 a_19401_3246# a_19700_3246# a_19635_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X1147 a_19171_n1353# x4.x15.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1148 VDD x3.x4.A a_11974_5018# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1149 a_13832_n572# a_13552_n938# a_13740_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X1150 a_22493_4119# x3.x39.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X1151 a_13892_13233# x2.x3.A a_13804_13095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1152 VSS x3.x20.Q_N a_12864_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X1153 vdd_sw[2] a_22671_n938# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1154 x3.x5.X a_11801_6580# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1155 a_28527_3784# a_27996_3790# a_28443_3784# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X1156 x5.x2.x9.output_stack x5.x2.x10.Y x5.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X1157 a_20114_77# VSS a_19900_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X1158 a_19564_4427# a_19146_4511# a_19320_4119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X1159 a_29224_2882# a_27996_2510# a_29082_2504# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X1160 x3.x77.Y x5.eob VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1161 x4.x9.A1 a_13898_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1162 a_15335_5300# a_14376_5018# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X1163 VSS a_24160_n1653# a_24070_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X1164 x1.x2.x10.Y async_setb_delay_cap_ctrl_code[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1165 a_8789_8870# x1.x10.A VDD VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1166 a_16874_5018# a_17010_4992# a_16455_4992# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X1167 a_20417_5018# a_19905_4992# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X1168 a_26225_1838# a_26051_2230# a_26365_1864# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X1169 VDD a_29398_2478# a_29310_2504# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X1170 a_25958_2504# x4.D[4] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X1171 a_22218_77# a_22036_77# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1172 a_19565_5989# a_19147_6073# a_19321_5681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X1173 VSS sar_clk a_12988_892# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1174 a_19644_n1443# a_19171_n1353# a_19888_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X1175 a_20619_5018# a_19701_4992# a_20173_5202# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1176 vdd_sw[7] a_10711_n938# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1177 x5.x1[3].Q_N a_29398_3118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X1178 a_20576_11982# x2.x2.x1.IN a_20488_11844# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1179 a_16728_n1261# a_15925_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X1180 a_26918_2230# a_25770_1864# a_26832_1864# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X1181 VDD a_23101_n1653# vss_sw_b[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X1182 a_16474_5707# a_16308_5707# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1183 a_18630_n1627# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X1184 VDD a_9222_n964# a_9132_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X1185 a_26159_1864# a_25770_1864# a_26051_2230# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X1186 a_17308_3246# x4.D[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1187 a_13952_n1627# a_14079_n1459# a_13533_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X1188 VDD sample_clk_b a_8604_892# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1189 VSS x3.x36.Q_N a_22432_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X1190 x5.x2.x5[7].floating x5.x2.x10.Y x5.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X1191 VDD a_27006_3758# a_26918_3784# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X1192 a_3051_10955# ready a_2979_11093# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1193 a_25770_3144# a_25604_3144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1194 a_17512_3246# a_17780_3456# a_17726_3554# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X1195 a_13968_4992# a_14063_4992# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1196 VDD x3.x7.X a_15834_3272# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X1197 a_11995_11952# a_11530_11926# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1198 a_24592_5685# x5.eob a_24504_5547# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1199 VSS x4.x13.S a_23011_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1200 a_25979_9043# x2.x2.x2.IN x2.x2.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1201 VDD a_13264_892# x4.x30.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1202 VDD a_28617_2478# a_28527_2504# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X1203 a_19376_n1653# a_19644_n1443# a_19590_n1345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X1204 x1.x4.x3[1].floating async_resetb_delay_cap_ctrl_code[1] x1.x4.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X1205 a_17166_n670# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X1206 x3.x20.Q_N a_12926_5681# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1207 a_23520_n1627# a_23647_n1459# a_23101_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X1208 VSS a_11386_7809# a_11320_7835# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1209 a_19317_7516# x2.x2.x3.IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1210 a_19360_5300# a_19160_5018# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X1211 VSS a_17513_4992# a_17448_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X1212 a_28162_3144# a_27996_3144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1213 a_19146_4511# a_18865_4145# a_19053_4145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X1214 a_29398_3118# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X1215 a_16474_5707# a_16308_5707# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1216 VDD a_22494_5681# a_23201_5707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1217 a_12225_3246# a_12523_3546# a_12459_3638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X1218 a_16132_n938# x4.D[4] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1219 sar_result[2] a_27713_3144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1220 x2.x2.x1.x3[1].floating sample_delay_cap_ctrl_code[5] x2.x2.x1.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X1221 x2.x2.x1.x5[7].floating x2.x2.x1.x10.Y x2.x2.x1.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X1222 VSS a_11995_n1353# a_11996_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1223 VSS x5.x3.X a_27996_2510# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1224 a_24093_n1261# a_23956_n1653# a_23647_n1459# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X1225 a_17393_4427# a_16928_4119# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1226 VSS a_11392_4144# x3.x7.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1227 a_11141_n1653# a_11454_n1627# a_11560_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1228 VDD a_26225_1838# a_26135_2230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X1229 a_11995_n1353# x4.x9.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1230 a_22280_n1261# a_21768_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X1231 VDD x2.x3.A a_13804_13371# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1232 a_17394_5989# a_16929_5681# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1233 a_15389_5202# a_14916_5292# a_15633_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X1234 a_24592_4857# x5.eob a_24504_4719# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1235 VDD a_23005_n1475# vss_sw[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1236 a_12926_5681# x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X1237 VSS a_21563_n1353# a_21564_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1238 VDD VDD a_9808_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X1239 a_21022_n1627# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1240 x2.x2.x3.x9.output_stack x2.x2.x3.x10.Y x2.x2.x3.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X1241 a_26365_3144# a_26519_3118# a_26225_3118# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1242 x4.x11.X a_15114_77# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X1243 a_13437_n1475# a_13533_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1244 a_19460_4145# x3.x42.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X1245 a_13346_6580# sel_bit[0] a_13247_6902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.105 ps=0.995 w=0.42 l=0.15
X1246 a_20218_5707# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X1247 VDD a_11974_5018# x3.x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1248 VSS x4.x15.S a_20619_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1249 x4.x13.X a_17508_77# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X1250 a_14916_3246# x4.D[5] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1251 a_17306_n938# a_16692_n964# a_17166_n670# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1252 a_3051_11231# ready a_2979_11369# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1253 a_19286_n1627# a_19171_n1353# a_18863_n1459# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X1254 a_18700_n572# a_18336_n938# a_18616_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X1255 a_14774_n670# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X1256 x4.x9.A1 a_13898_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1257 x2.x2.x3.x6.SW sample_delay_offset VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1258 a_12639_n656# a_12223_n572# a_12382_n670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X1259 a_10685_8876# a_10817_8528# a_10549_8788# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X1260 a_18847_4992# a_19160_5018# a_19266_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1261 a_19321_5681# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X1262 VSS VDD a_21128_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X1263 x2.x2.x1.x9.output_stack x2.x2.x1.IN a_20576_11982# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1264 a_25979_9319# x2.x2.x2.IN a_25891_9181# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1265 VDD a_14063_4992# x3.x48.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X1266 a_15925_n1653# a_16238_n1627# a_16344_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1267 VSS x4.x3.X a_9514_892# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1268 a_25770_3144# a_25604_3144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1269 a_16754_4511# a_16473_4145# a_16661_4145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X1270 VSS a_12261_8772# a_11883_8462# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1271 a_9734_n938# a_9222_n964# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X1272 VDD a_20102_5681# a_20809_5707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1273 a_10280_8920# a_9491_8544# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X1274 a_13740_n938# x4.D[5] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1275 a_22494_5681# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X1276 VSS VDD a_15257_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X1277 a_13252_8655# x2.x7.A VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X1278 a_19171_n1353# x4.x15.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1279 a_11045_n1475# a_11141_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1280 a_12838_6073# a_11690_5707# a_12752_5707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X1281 a_20601_12957# x2.x2.x1.IN a_20513_13095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1282 VSS x5.x3.X a_25604_2510# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1283 a_22428_4145# a_21091_4145# a_22319_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X1284 a_20121_n250# x4.x9.A1 a_19900_77# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X1285 a_29333_2882# a_27996_2510# a_29224_2882# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X1286 a_15001_4427# a_14536_4119# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1287 a_8789_8529# x1.x4.x9.output_stack VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1288 a_12183_3554# a_11983_3272# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X1289 VSS a_11974_5018# x3.x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1290 a_11758_n938# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X1291 a_17508_77# VSS a_17508_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1292 VDD a_26519_3984# a_26469_3784# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X1293 x2.x2.x3.x5[7].floating x2.x2.x3.x10.Y x2.x2.x3.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X1294 x4.x11.X a_15114_77# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X1295 x2.x2.x3.x7.floating sample_delay_offset x2.x2.x3.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1296 x1.x4.x5[7].floating x1.x4.x10.Y x1.x4.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X1297 a_15002_5989# a_14537_5681# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1298 VSS VDD a_9168_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X1299 x2.x2.x2.x3[1].floating sample_delay_cap_ctrl_code[9] x2.x2.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X1300 VDD a_11883_8462# sample_clk VDD sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X1301 a_12145_5681# a_11971_6073# a_12285_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X1302 x1.x9.Y x1.x9.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1303 a_20613_n1475# a_20709_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1304 a_22290_77# VSS a_22290_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1305 x4.x2.X a_9514_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1306 VSS retimer_eob_delay_offset x5.x2.x6.SW VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1307 x4.x7.S a_16025_5707# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X1308 VDD a_21182_n964# a_21092_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X1309 a_21445_4145# x3.x7.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1310 a_11416_8162# VSS a_10957_7987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X1311 a_12079_5707# a_11690_5707# a_11971_6073# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X1312 VSS x3.x3.A a_11360_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1313 a_17943_4427# a_17535_4145# a_17709_4119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X1314 a_29514_4150# a_28911_3984# a_29398_3758# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1315 a_22809_5384# a_22297_4992# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X1316 a_10320_n1627# a_9808_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X1317 a_17944_5989# a_17536_5707# a_17710_5681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X1318 VSS x2.x2.x1.IN a_19677_12370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X1319 VDD a_9514_892# x4.x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1320 VSS VDD a_14728_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X1321 a_26832_4162# a_25770_3790# a_26737_4106# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X1322 VSS a_15925_n1653# vss_sw_b[4] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1323 x2.x2.x1.x5[7].floating x2.x2.x1.x10.Y x2.x2.x1.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X1324 VDD a_21144_4992# x4.x15.S VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1325 x2.x2.x3.IN x2.x2.x2.x9.output_stack a_19961_8858# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X1326 a_16455_4992# a_16768_5018# a_16874_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1327 a_14615_n572# a_13552_n938# a_14471_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X1328 a_17645_5707# a_16308_5707# a_17536_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X1329 a_19506_n938# a_18336_n938# a_19399_n572# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X1330 VDD ready a_2916_12896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1331 a_19147_6073# a_18866_5707# a_19054_5707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X1332 VDD x4.x5.D a_10521_n1627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1333 a_21751_3554# a_21551_3272# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X1334 a_18582_n250# VSS a_18219_n98# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X1335 a_20576_11154# x2.x2.x1.IN a_20488_11016# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1336 a_24086_n938# a_23574_n964# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X1337 sar_result[1] a_30105_3800# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1338 a_26832_3144# a_25604_3144# a_26690_3426# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X1339 VDD x5.x3.A a_30402_5732# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X1340 a_18524_n938# x4.D[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1341 a_12945_n250# x4.x9.A1 a_12724_77# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X1342 x5.x1[1].Q_N a_29398_3758# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X1343 a_21713_5681# a_21539_6073# a_21853_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X1344 a_23574_n964# a_23400_n572# a_23718_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X1345 VDD a_13864_n276# a_13894_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1346 VDD x4.x17.S a_13432_6946# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.138 ps=1.16 w=0.64 l=0.15
X1347 a_14323_n1627# a_13533_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X1348 a_26941_2882# a_25604_2510# a_26832_2882# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X1349 a_19147_6073# a_18700_5707# a_19054_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1350 VDD a_11995_n1353# a_11996_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1351 VDD a_18219_n98# x4.x14.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X1352 VSS x3.x4.X a_17222_4119# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1353 a_12126_n938# a_11614_n964# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X1354 a_18751_3246# a_18846_3246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1355 VDD a_17308_3246# a_17307_3546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1356 a_21647_5707# a_21258_5707# a_21539_6073# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X1357 a_23508_n938# a_22954_n938# a_23400_n572# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X1358 a_29333_3144# a_27996_3144# a_29224_3144# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X1359 VSS VDD a_12336_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X1360 x3.x36.Q_N a_22494_5681# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X1361 VSS a_17709_4119# a_17644_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X1362 a_21794_4992# a_22092_5292# a_22028_5384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X1363 x4.x2.X a_9514_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1364 x1.x4.x9.output_stack x1.x4.x10.Y x1.x4.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X1365 a_13898_892# x4.x30.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1366 VSS a_26225_2478# a_26159_2882# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X1367 a_17120_n1627# a_17252_n1443# a_16984_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X1368 a_23891_n1627# a_23101_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X1369 a_27006_2478# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X1370 x3.x27.D a_13633_5707# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X1371 a_22297_4992# a_21552_5018# a_22433_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1372 VDD a_21563_n1353# a_21564_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1373 a_9080_n276# x4.x7.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1374 VSS a_22493_4119# a_22428_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X1375 a_15632_3272# a_15120_3246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X1376 a_28443_2504# a_27996_2510# a_28350_2504# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1377 x5.x2.x9.output_stack x5.eob a_24529_6522# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1378 VDD VDD a_17513_4992# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X1379 a_15834_3272# a_14916_3246# a_15388_3456# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1380 VDD a_17512_3246# a_17445_3638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X1381 x2.x2.x4.x4[3].floating sample_delay_cap_ctrl_code[2] x2.x2.x4.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X1382 a_10130_7987# VSS a_10272_7835# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1383 a_17780_3456# a_17307_3546# a_18024_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X1384 VDD VDD a_28911_2704# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X1385 x2.x2.x4.x9.output_stack x2.x2.x4.x10.Y x2.x2.x4.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X1386 VDD x4.x7.S a_10078_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X1387 VDD a_12439_5681# a_12389_5989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X1388 a_24342_n670# a_24183_n572# a_24482_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X1389 vdd_sw[4] a_17887_n938# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X1390 x1.x4.x5[7].floating x1.x4.x10.Y x1.x4.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X1391 x4.x9.A1 a_13898_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1392 a_28757_2870# a_28911_2704# a_28617_2478# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1393 a_21538_4511# a_21091_4145# a_21445_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1394 VDD VDD a_11263_8932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X1395 VDD VDD a_28911_3118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X1396 a_9603_n1353# x4.x7.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1397 a_16755_6073# a_16474_5707# a_16662_5707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X1398 VSS a_21712_4119# a_21646_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X1399 VSS x4.x20.S a_24905_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X1400 a_17009_3246# a_17308_3246# a_17243_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X1401 a_21694_n938# a_21182_n964# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X1402 a_23955_n1353# x4.x20.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1403 a_21499_n1627# a_20709_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X1404 a_14340_6580# a_13316_6554# a_13836_6580# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.072 ps=0.76 w=0.36 l=0.15
X1405 VSS x3.x7.A a_11392_4144# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1406 a_20101_4119# x3.x42.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X1407 a_21793_3246# a_22092_3246# a_22027_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X1408 a_28527_2504# a_27996_2510# a_28443_2504# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X1409 VSS a_14592_n1653# a_14502_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X1410 VSS a_17710_5681# a_17645_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X1411 VSS a_19558_n670# a_19506_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X1412 VDD x2.x2.x2.IN a_26386_12029# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X1413 a_23010_3272# a_22091_3546# a_22564_3456# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1414 a_16755_6073# a_16308_5707# a_16662_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1415 a_14336_n1261# a_13533_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X1416 a_2979_9331# sar_clk a_2891_9331# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1417 a_12652_77# a_12470_77# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1418 VSS x3.x4.X a_14830_4119# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1419 a_18751_3246# a_18846_3246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1420 a_9910_8876# a_10046_8528# a_9491_8544# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X1421 VSS x3.x4.A a_11974_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1422 VSS a_16929_5681# a_16863_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X1423 a_26941_3144# a_25604_3144# a_26832_3144# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X1424 VSS a_29398_3118# a_29333_3144# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X1425 a_25958_3144# x4.D[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1426 a_17780_3456# a_17308_3246# a_18024_3638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X1427 x3.x33.Q_N a_20102_5681# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X1428 VDD VDD a_26519_3984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X1429 x2.x1.x3.Y VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1430 a_14376_5018# x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1431 VDD a_17166_n670# a_17091_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X1432 x5.x1[7].Q_N a_29398_1838# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X1433 a_20648_11154# x2.x2.x1.IN a_20576_11154# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1434 a_26135_3784# a_25604_3790# a_26051_3784# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X1435 a_17621_4511# a_16473_4145# a_17535_4145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X1436 a_9539_n1627# a_8749_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X1437 a_26386_12370# x2.x2.x1.x9.output_stack x2.x2.x2.IN VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X1438 VSS VDD a_28911_2704# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1439 x2.x2.x1.x5[7].floating x2.x2.x1.x10.Y x2.x2.x1.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X1440 a_13456_6580# sel_bit[0] a_13346_6580# VSS sky130_fd_pr__nfet_01v8 ad=0.0786 pd=0.805 as=0.072 ps=0.76 w=0.36 l=0.15
X1441 a_11185_77# x4.x9.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X1442 x4.x9.A1 a_13898_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1443 VDD a_27006_2478# a_26918_2504# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X1444 VDD a_29398_3118# a_30105_3144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1445 a_15120_3246# a_15388_3456# a_15334_3554# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X1446 VDD VDD a_18317_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X1447 x3.x72.Q_N a_17709_4119# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1448 VSS VDD a_21476_n964# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1449 a_10332_77# x4.x9.A1 a_10260_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1450 VSS x3.x7.X a_15834_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1451 VDD a_15829_n1475# vss_sw[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1452 a_9514_892# x4.x3.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1453 VDD a_10549_8788# a_10482_8554# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X1454 x4.x3.X a_8880_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1455 a_28443_3510# a_27996_3144# a_28350_3144# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1456 VSS a_28617_3118# a_28551_3144# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X1457 vdd_sw[5] a_15495_n938# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X1458 a_19376_n1653# a_18630_n1627# a_19512_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1459 a_15256_3272# a_15388_3456# a_15120_3246# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X1460 a_19636_5018# a_18847_4992# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X1461 a_24482_n938# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X1462 a_19159_3272# x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X1463 VDD x3.x7.X a_13442_3272# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X1464 a_19460_4145# a_19614_4119# a_19320_4119# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1465 VSS VDD a_9516_n964# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1466 a_28350_3784# x4.D[1] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X1467 VSS a_10549_8788# a_10484_8932# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X1468 a_14617_3246# a_14916_3246# a_14851_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X1469 VSS a_21768_n1653# a_21678_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X1470 a_21070_77# x4.x9.A1 a_20611_n98# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X1471 VDD a_18648_n276# a_18678_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1472 a_14525_n1261# a_14388_n1653# a_14079_n1459# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X1473 VDD x3.x33.Q_N a_18846_3246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X1474 x1.x2.x4[3].floating async_setb_delay_cap_ctrl_code[2] x1.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X1475 a_19317_7792# x2.x2.x3.IN a_19229_7930# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1476 VSS a_11974_5018# x3.x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1477 VDD comp_result a_11116_4144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1478 a_8793_n250# x4.x7.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X1479 x1.x2.x9.output_stack x1.x2.x10.Y x1.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X1480 a_12522_n938# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X1481 VSS a_9514_892# x4.x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1482 x5.x2.x2.floating retimer_delay_code[0] x5.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X1483 a_12712_n1261# a_12200_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X1484 VDD a_28911_3118# a_28861_3426# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X1485 VDD a_13437_n1475# vss_sw[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1486 x2.x7.A x2.x2.x3.x9.output_stack a_13252_8858# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X1487 VSS x4.D[3] a_20089_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1488 VDD x3.x36.Q_N a_22296_3246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X1489 a_28162_3790# a_27996_3790# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1490 a_21144_4992# a_21239_4992# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1491 x2.x2.x4.x4[3].floating sample_delay_cap_ctrl_code[2] x2.x2.x4.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X1492 VDD VDD a_14300_n964# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X1493 x2.x2.x4.x9.output_stack x2.x2.x4.x10.Y x2.x2.x4.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X1494 a_15388_3456# a_14916_3246# a_15632_3638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X1495 a_17309_4992# x3.x5.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1496 VDD a_14774_n670# a_14699_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X1497 x2.x1.x2.D a_12311_11926# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1498 VDD a_23868_n964# a_23818_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X1499 a_2979_9607# sar_clk a_2891_9607# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1500 VSS a_9808_n1653# a_9718_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X1501 a_18025_5018# a_17513_4992# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X1502 a_28617_1838# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X1503 a_12524_3246# x4.D[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1504 a_19034_n656# a_18616_n572# a_18790_n964# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X1505 VSS a_29398_1838# a_30105_1864# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1506 a_17068_4145# x3.x45.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X1507 x3.x7.X a_11392_4144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1508 a_12728_3246# a_12996_3456# a_12942_3554# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X1509 a_27006_2478# a_26832_2882# a_27122_2870# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X1510 VSS a_29398_3758# a_30105_3800# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1511 x2.x2.x2.x6.floating x2.x2.x2.x6.SW x2.x2.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1512 vdd_sw_b[2] a_21950_n670# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X1513 a_29082_2146# a_28617_1838# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1514 a_11974_5018# x3.x4.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1515 a_13533_n1653# a_13846_n1627# a_13952_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1516 a_16308_n572# a_15944_n938# a_16224_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X1517 a_28861_2146# a_28443_2230# a_28617_1838# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X1518 x5.x1[4].Q_N a_27006_2478# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1519 a_19644_n1443# a_19172_n1653# a_19888_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X1520 a_10022_n1345# a_9062_n1627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X1521 a_15114_n250# a_14860_77# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X1522 a_14576_5300# a_14376_5018# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X1523 x4.x20.X a_24684_77# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X1524 VDD a_26519_3984# a_27240_3784# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X1525 x5.x2.x9.output_stack x5.eob a_24592_5685# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1526 VSS a_23955_n1353# a_23956_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1527 a_27122_2870# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X1528 VSS a_11974_5018# x3.x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1529 a_9603_n1353# x4.x7.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1530 vdd_sw_b[7] a_9990_n670# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X1531 a_11348_n938# x4.D[6] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1532 VSS a_13898_892# x4.x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1533 a_19927_4145# a_18699_4145# a_19785_4427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X1534 a_23414_n1627# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1535 VDD VDD a_23868_n964# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X1536 a_23955_n1353# x4.x20.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1537 a_12382_n670# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X1538 a_26051_3784# a_25604_3790# a_25958_3784# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1539 a_25979_9733# x2.x2.x2.IN a_25891_9733# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1540 a_17423_n656# a_17007_n572# a_17166_n670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X1541 a_26225_3118# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X1542 a_11263_8932# a_10345_8772# a_10817_8528# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1543 a_18847_4992# a_19402_4992# a_19360_5300# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X1544 a_19402_4992# a_19701_4992# a_19636_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X1545 VDD a_26519_2704# a_26469_2504# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X1546 a_8789_11554# x1.x2.x9.output_stack VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1547 a_8789_8529# x1.x10.A VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1548 VDD a_12852_6554# x5.eob VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X1549 VSS a_9514_892# x4.x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1550 a_25770_3790# a_25604_3790# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1551 a_12055_6073# a_11524_5707# a_11971_6073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X1552 VSS x4.x3.A a_8880_892# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1553 VSS a_12311_11926# a_12246_12330# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X1554 VDD VDD a_21768_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X1555 VDD VDD a_11908_n964# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X1556 a_11758_n938# a_11908_n964# a_11614_n964# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1557 a_19900_n250# a_19646_77# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X1558 a_22092_3246# x4.D[2] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1559 VSS a_14062_3246# x3.x54.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1560 VSS x3.x5.X a_21092_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1561 VSS x4.x14.X a_18170_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1562 a_20036_4145# a_18699_4145# a_19927_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X1563 a_17622_6073# a_16474_5707# a_17536_5707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X1564 x4.x7.X a_10332_77# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X1565 VSS a_22092_3246# a_22091_3546# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1566 a_2979_10679# ready a_2891_10541# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1567 a_30402_6073# x5.x3.A VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1568 a_28443_2230# a_28162_1864# a_28350_1864# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X1569 a_19677_12029# x2.x2.x4.x9.output_stack VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1570 x2.x3.Y VDD a_12261_7986# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1571 a_22609_4145# a_22006_4119# a_22493_4119# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1572 VSS sample_clk_b a_11084_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1573 a_16642_n656# a_16224_n572# a_16398_n964# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X1574 a_14676_4145# x3.x77.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X1575 a_22510_3554# a_21551_3272# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X1576 a_24664_4857# x5.eob a_24592_4857# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1577 VDD a_21239_4992# x3.x39.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X1578 x3.x4.X a_11974_5018# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1579 a_20753_77# x4.x17.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X1580 a_19677_12370# x2.x2.x1.IN VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1581 a_3051_10955# ready a_2979_10955# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1582 a_17512_3246# a_16767_3272# a_17648_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1583 a_23574_n964# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X1584 VSS a_9222_n964# a_9156_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X1585 a_17309_4992# x3.x5.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1586 a_26690_2146# a_26225_1838# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1587 VDD a_11824_12152# a_11774_11952# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X1588 x4.x13.X a_17508_77# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X1589 a_11440_11952# a_10909_11958# a_11356_11952# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X1590 a_15835_5018# a_14916_5292# a_15389_5202# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1591 VSS VDD a_22433_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X1592 a_13916_n572# a_13552_n938# a_13832_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X1593 a_14270_5707# x3.x27.D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X1594 a_28757_2870# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X1595 a_21213_n1345# a_21022_n1627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X1596 a_17826_5707# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X1597 sar_result[7] a_30105_1864# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1598 VDD x4.D[5] a_15305_n1627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1599 a_17697_n1627# a_16780_n1653# a_17252_n1443# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X1600 a_15055_3272# a_14915_3546# a_14617_3246# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X1601 a_20619_5018# a_19700_5292# a_20173_5202# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1602 a_17826_5707# a_17223_5681# a_17710_5681# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1603 a_23005_n1475# a_23101_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1604 VDD x3.x5.X a_21092_5707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1605 a_15969_n250# x4.x13.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X1606 VSS VDD a_26519_1838# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1607 VDD x3.x4.X a_19614_4119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X1608 a_26026_7792# x2.x2.x2.IN a_25938_7654# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1609 VSS a_17709_4119# a_18416_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1610 VSS VDD a_26519_3984# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1611 x5.x1[5].Q_N a_29398_2478# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X1612 a_29632_2146# a_29224_1864# a_29398_1838# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X1613 x4.x13.S a_23201_5707# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X1614 sample_clk_b a_11883_7842# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1615 a_26051_3510# a_25770_3144# a_25958_3144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X1616 VSS a_13898_892# x4.x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1617 a_23647_n1459# a_23955_n1353# a_23904_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X1618 VDD a_9514_892# x4.x2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1619 a_9253_n1345# a_9062_n1627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X1620 a_16132_n938# x4.D[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1621 a_29514_3144# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X1622 VSS VDD a_17120_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X1623 VSS a_21143_3246# x4.D[3] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1624 a_14470_4145# a_14081_4145# a_14362_4511# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X1625 VSS a_24342_n670# a_25063_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1626 a_29514_3144# a_28911_3118# a_29398_3118# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1627 VSS a_23003_n98# x4.x18.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X1628 a_11263_11952# x2.x1.x2.D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1629 a_13836_6580# a_13721_6554# a_12852_6554# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.6 as=0.0729 ps=0.81 w=0.54 l=0.15
X1630 a_24592_5271# x5.eob a_24504_5271# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1631 a_19700_3246# x4.D[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1632 VSS x4.x12.X a_15778_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1633 VSS x3.x5.A a_11801_6580# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1634 VSS x4.x9.S a_12945_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X1635 a_11670_3246# a_12225_3246# a_12183_3554# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X1636 VSS a_19700_3246# a_19699_3546# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1637 a_22280_n1627# a_21768_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X1638 x2.x2.x4.x9.output_stack x2.x2.x4.x6.SW x2.x2.x4.x6.floating VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1639 a_10046_8528# a_10345_8772# a_10280_8920# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X1640 a_10763_8554# a_9804_8920# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X1641 a_14471_n656# a_14006_n964# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1642 a_22511_n250# x4.x9.A1 a_22290_77# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X1643 a_23003_n98# VSS a_23145_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X1644 a_22504_77# VSS a_22290_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X1645 x2.x2.x3.x9.output_stack x2.x2.x3.x10.Y x2.x2.x3.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X1646 VDD a_13533_n1653# vss_sw_b[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X1647 VSS a_11392_4144# x3.x7.X VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1648 VDD a_10559_7809# a_10589_8162# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1649 VSS a_12382_n670# a_13103_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1650 VSS a_11043_n98# x4.x8.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X1651 a_15317_4119# a_15143_4145# a_15433_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X1652 VDD a_18790_n964# a_18700_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X1653 a_21950_n670# a_21791_n572# a_22090_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X1654 VDD x4.x9.S a_12938_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X1655 VDD x4.D[2] a_22481_n1627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1656 a_23400_n572# a_22954_n938# a_23308_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X1657 VSS a_20101_4119# a_20036_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X1658 VSS a_30706_5822# x5.x3.X VSS sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X1659 a_26365_2870# a_26519_2704# a_26225_2478# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1660 a_3004_12482# ready a_2916_12620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1661 a_27240_3426# a_26832_3144# a_27006_3118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X1662 VDD a_11386_7809# a_11416_8162# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1663 a_9831_n572# a_8602_n938# a_9734_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X1664 VDD VDD a_28911_1838# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X1665 VSS x2.x2.x3.IN a_19961_8655# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1666 VDD a_22493_4119# a_23200_4145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1667 a_16473_4145# a_16307_4145# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1668 a_14387_n1353# x4.x11.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1669 VDD x4.x30.A a_13898_892# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1670 VSS x3.x4.A a_11974_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1671 a_13798_n250# VSS a_13435_n98# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X1672 a_12663_3272# a_12523_3546# a_12225_3246# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X1673 VDD VDD a_19905_4992# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X1674 VSS a_12200_n1653# a_12110_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X1675 a_28617_3758# a_28443_3784# a_28757_4150# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X1676 VDD a_11043_n98# x4.x8.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X1677 VSS comp_result a_11116_4144# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1678 a_8789_11895# x1.x2.x9.output_stack x1.x9.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X1679 VDD a_18752_4992# x4.x17.S VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1680 VDD a_23955_n1353# a_23956_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1681 x2.x2.x3.x6.floating x2.x2.x3.x6.SW x2.x2.x3.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1682 a_19317_8068# x2.x2.x3.IN x2.x2.x3.x9.output_stack VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1683 a_26386_12029# x2.x2.x2.IN VDD VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1684 VDD a_22007_5681# a_22728_5989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X1685 x4.x11.S a_20809_5707# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X1686 VDD a_11141_n1653# vss_sw_b[6] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X1687 VSS a_15318_5681# a_15253_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X1688 a_19833_5707# a_19321_5681# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X1689 sar_result[0] a_27713_3800# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1690 VSS VDD a_24296_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X1691 VSS a_17166_n670# a_17114_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X1692 a_17243_3638# a_16454_3246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X1693 a_20601_12957# x2.x2.x1.IN a_20513_12819# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1694 VSS a_15120_3246# a_15055_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X1695 a_8768_n938# a_8602_n938# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1696 VDD a_17166_n670# a_17887_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1697 a_17445_3638# a_17308_3246# a_17009_3246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X1698 a_20709_n1653# a_21255_n1459# a_21213_n1345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X1699 a_19928_5707# a_18700_5707# a_19786_5989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X1700 a_13740_n938# x4.D[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1701 a_16224_n572# a_15944_n938# a_16132_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X1702 x3.D[0] a_18416_4145# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1703 VSS a_21950_n670# a_22671_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1704 a_20576_11844# x2.x2.x1.IN a_20488_11844# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1705 VSS a_20611_n98# x4.x16.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X1706 a_26135_2504# a_25604_2510# a_26051_2504# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X1707 a_15229_4511# a_14081_4145# a_15143_4145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X1708 VDD x4.x9.S a_12470_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X1709 a_22565_5202# a_22093_4992# a_22809_5384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X1710 a_13316_6554# sel_bit[0] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1711 VDD x4.x14.X a_18170_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1712 a_13864_n276# x4.x11.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1713 VDD sar_clk a_11525_6580# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1714 x2.x2.x4.x9.output_stack sample_delay_cap_ctrl_code[2] x2.x2.x4.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X1715 a_19402_4992# a_19700_5292# a_19636_5384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X1716 VSS VDD a_19084_n964# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1717 a_24592_5547# x5.eob a_24504_5547# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1718 a_28757_1864# a_28911_1838# a_28617_1838# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1719 VSS a_27006_3118# a_26941_3144# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X1720 VSS a_9990_n670# a_10711_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1721 a_9222_n964# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X1722 vdd_sw[1] a_25063_n938# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1723 a_18736_n1627# a_18863_n1459# a_18317_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X1724 a_11356_11952# a_11075_11958# a_11263_11952# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X1725 VSS a_21182_n964# a_21116_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X1726 a_21563_n1353# x4.x17.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1727 a_10493_7835# x1.x3.X a_10130_7987# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X1728 x4.x9.A1 a_13898_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1729 a_9062_n1627# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X1730 VDD a_13898_892# x4.x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1731 VSS a_11974_5018# x3.x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1732 a_26737_4106# a_26225_3758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X1733 a_24183_n572# a_22954_n938# a_24086_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X1734 VDD a_28911_3118# a_29632_3426# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X1735 a_12133_n1261# a_11996_n1653# a_11687_n1459# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X1736 VSS x4.x3.X a_9514_892# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1737 a_28350_2504# x4.D[5] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X1738 VSS x3.x7.X a_13442_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1739 VDD a_20101_4119# a_20808_4145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1740 VSS x3.x4.X a_22006_4119# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1741 vdd_sw[6] a_13103_n938# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1742 VSS a_11360_5018# x3.x4.A VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1743 a_29310_2230# a_28162_1864# a_29224_1864# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X1744 a_21657_3272# a_21793_3246# a_21238_3246# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X1745 a_12864_3272# a_12996_3456# a_12728_3246# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X1746 VSS x4.x5.D a_10521_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1747 VSS a_12926_5681# a_12861_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X1748 x5.x2.x5[7].floating x5.x2.x10.Y x5.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X1749 a_19928_5707# a_18866_5707# a_19833_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X1750 VSS a_14774_n670# a_14722_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X1751 VDD x3.x7.X a_18226_3272# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X1752 a_14851_3638# a_14062_3246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X1753 VDD a_18221_n1475# vss_sw[3] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1754 a_16473_4145# a_16307_4145# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1755 VDD x3.x4.X a_19615_5681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X1756 VDD a_18846_3246# x3.x60.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X1757 a_28162_2510# a_27996_2510# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1758 VSS x3.x30.Q_N a_16873_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X1759 a_17709_4119# x3.x45.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X1760 a_24592_4719# x5.eob a_24504_4719# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1761 a_13577_77# x4.x11.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X1762 VSS a_16779_n1353# a_16780_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1763 a_26365_1864# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X1764 VDD x3.x30.Q_N a_16454_3246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X1765 a_26365_4150# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X1766 x5.x2.x10.Y retimer_delay_code[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1767 x4.x2.X a_9514_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1768 a_22564_3456# a_22091_3546# a_22808_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X1769 a_12042_12274# a_11530_11926# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X1770 a_10130_n938# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X1771 x3.x4.X a_11974_5018# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1772 VDD x1.x9.A a_8789_11554# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X1773 vdd_sw[2] a_22671_n938# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X1774 a_13864_n276# x4.x11.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X1775 a_21445_4145# x3.x7.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X1776 a_26918_3784# a_25770_3790# a_26832_4162# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X1777 VDD x4.x12.X a_15778_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1778 a_22432_3272# a_22564_3456# a_22296_3246# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X1779 VSS a_11974_5018# x3.x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1780 a_17069_5707# a_17223_5681# a_16929_5681# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1781 a_18934_n938# a_19084_n964# a_18790_n964# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1782 a_24898_77# VSS a_24684_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X1783 a_15633_5018# a_15121_4992# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X1784 a_15104_n1261# a_14592_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X1785 a_9048_n572# a_8602_n938# a_8956_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X1786 a_26469_2146# a_26051_2230# a_26225_1838# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X1787 VSS a_12311_11926# a_13018_11968# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1788 a_23462_77# x4.x9.A1 a_23003_n98# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X1789 VDD a_27006_3118# a_27713_3144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1790 vdd_sw[7] a_10711_n938# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X1791 a_13867_11292# x2.x3.A a_13779_11292# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1792 x5.eob a_12852_6554# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X1793 VSS x3.x4.X a_22007_5681# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1794 a_15835_5018# a_14917_4992# a_15389_5202# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1795 x4.x2.X a_9514_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1796 VSS a_14387_n1353# a_14388_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1797 a_11160_n938# a_10994_n938# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1798 a_20648_11706# x2.x2.x1.IN a_20576_11844# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1799 x1.x2.x9.output_stack async_setb_delay_cap_ctrl_code[2] x1.x2.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X1800 x3.x5.X a_11801_6580# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1801 a_21791_n572# a_20562_n938# a_21694_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X1802 a_14375_3272# x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X1803 a_17781_5202# a_17308_5292# a_18025_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X1804 VDD a_26519_2704# a_27240_2504# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X1805 vdd_sw_b[3] a_19558_n670# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1806 x4.x9.A1 a_13898_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1807 a_14387_n1353# x4.x11.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1808 a_24672_n1261# a_24160_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X1809 VSS sample_clk_b a_8604_892# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1810 a_26026_8068# x2.x2.x2.IN a_25938_7930# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1811 VDD VDD a_21476_n964# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X1812 x5.x2.x9.output_stack retimer_delay_code[2] x5.x2.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X1813 VDD a_21040_n276# a_21070_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1814 VDD ext_clk a_10909_11958# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1815 x2.x2.x4.x9.output_stack sample_delay_cap_ctrl_code[2] x2.x2.x4.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X1816 a_19961_8858# x2.x2.x3.IN VDD VSS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
X1817 x2.x2.x1.x10.Y sample_delay_cap_ctrl_code[7] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1818 VDD a_17710_5681# a_18417_5707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1819 VDD a_11824_12152# a_12545_11952# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X1820 a_19483_n572# a_18170_n938# a_19399_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X1821 a_17010_4992# a_17309_4992# a_17244_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X1822 a_14062_3246# a_14375_3272# a_14481_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1823 VSS x2.x7.A a_13252_8655# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1824 a_15328_77# VSS a_15114_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X1825 x3.x4.X a_11974_5018# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1826 VDD VDD a_12200_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X1827 a_14079_n1459# a_14387_n1353# a_14336_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X1828 a_23432_n276# x4.x20.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X1829 VDD a_16454_3246# x3.x57.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X1830 a_25770_2510# a_25604_2510# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1831 VSS x3.x27.Q_N a_14481_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X1832 a_20728_n938# a_20562_n938# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1833 VDD a_26225_3758# a_26135_3784# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X1834 a_17535_4145# a_16307_4145# a_17393_4427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X1835 a_21794_4992# a_22093_4992# a_22028_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X1836 VSS VDD a_13952_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X1837 a_15829_n1475# a_15925_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1838 VDD VDD a_9516_n964# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X1839 VDD x4.x13.S a_17254_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X1840 VDD x3.x27.Q_N a_14062_3246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X1841 a_28551_4162# a_28162_3790# a_28443_3784# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X1842 a_8768_n938# a_8602_n938# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1843 a_17508_n250# a_17254_77# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X1844 a_27006_1838# a_26832_1864# a_27122_1864# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X1845 VDD a_17709_4119# a_17621_4511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X1846 a_3004_7666# sar_clk a_2916_7528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1847 a_15031_n656# a_14615_n572# a_14774_n670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X1848 a_20217_4145# x3.x42.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X1849 a_22319_4145# a_21091_4145# a_22177_4427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X1850 a_25979_10009# x2.x2.x2.IN VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1851 a_19270_9595# x2.x2.x3.IN a_19182_9457# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1852 x4.x2.X a_9514_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1853 a_18752_4992# a_18847_4992# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1854 a_20217_4145# a_19614_4119# a_20101_4119# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1855 a_11472_n276# x4.x9.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X1856 VDD a_22493_4119# a_22405_4511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X1857 a_20118_3554# a_19159_3272# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X1858 x3.x4.A a_11360_5018# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1859 VSS VDD a_23520_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X1860 VDD x4.x7.S a_10546_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X1861 a_8651_n98# VSS a_8793_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X1862 a_13968_4992# a_14063_4992# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1863 a_23432_n276# x4.x20.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1864 a_18317_n1653# a_18630_n1627# a_18736_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1865 a_15120_3246# a_14375_3272# a_15256_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1866 a_21182_n964# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X1867 a_15230_6073# a_14082_5707# a_15144_5707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X1868 a_14677_5707# a_14831_5681# a_14537_5681# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1869 a_16542_n938# a_16692_n964# a_16398_n964# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1870 VSS a_27006_1838# a_27713_1864# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1871 VSS x3.x4.A a_11974_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1872 a_11687_n1459# a_11995_n1353# a_11944_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X1873 a_19904_3246# a_19159_3272# a_20040_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1874 VSS a_27006_3758# a_27713_3800# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1875 a_21563_n1353# x4.x17.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1876 a_14150_n938# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X1877 a_24599_n656# a_24183_n572# a_24342_n670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X1878 a_13437_n1475# a_13533_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1879 a_12724_77# x4.x9.A1 a_12652_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1880 VSS a_11883_8462# sample_clk VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1881 VDD x5.eob a_24529_7074# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1882 x4.x15.X a_19900_77# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X1883 a_11983_3272# x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X1884 a_20576_11016# x2.x2.x1.IN a_20488_11016# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1885 x1.x4.x10.Y async_resetb_delay_cap_ctrl_code[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1886 VDD a_21712_4119# a_21622_4511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X1887 a_15054_5384# a_14917_4992# a_14618_4992# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X1888 a_18863_n1459# a_19171_n1353# a_19120_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X1889 a_13867_11568# x2.x3.A a_13779_11568# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1890 a_29224_4162# a_28162_3790# a_29129_4106# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X1891 a_19359_3554# a_19159_3272# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X1892 a_15257_5018# a_15389_5202# a_15121_4992# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X1893 a_15434_5707# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X1894 VSS a_21238_3246# x3.x63.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1895 x3.x4.X a_11974_5018# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1896 x4.x3.X a_8880_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1897 x1.x2.x9.output_stack async_delay_offset x1.x2.x7.floating VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1898 VSS x4.x20.S a_15835_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1899 a_11931_n1627# a_11141_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X1900 a_18361_77# x4.x15.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X1901 x5.x1[3].Q_N a_29398_3118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1902 a_14063_4992# a_14618_4992# a_14576_5300# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X1903 a_14618_4992# a_14917_4992# a_14852_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X1904 x3.x75.Q a_16024_4145# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X1905 a_15434_5707# a_14831_5681# a_15318_5681# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1906 a_24039_n656# a_23574_n964# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1907 a_17710_5681# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X1908 a_23718_n938# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X1909 a_13939_11154# x2.x3.A a_13867_11292# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1910 a_29224_3144# a_27996_3144# a_29082_3426# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X1911 a_20218_5707# a_19615_5681# a_20102_5681# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1912 x5.x2.x4[3].floating retimer_delay_code[2] x5.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X1913 VDD a_22093_4992# a_22092_5292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1914 a_15827_n98# x4.x9.A1 a_15969_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1915 VDD a_29398_3118# a_29310_3510# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X1916 a_25958_3144# x4.D[2] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X1917 a_12285_5707# x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X1918 VDD a_16779_n1353# a_16780_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1919 x2.x2.x4.x9.output_stack sample_delay_offset x2.x2.x4.x7.floating VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1920 a_12712_n1627# a_12200_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X1921 VSS x4.x10.X a_13386_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1922 VDD a_16692_n964# a_17423_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X1923 x1.x2.x3[1].floating async_setb_delay_cap_ctrl_code[1] x1.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X1924 VSS sar_clk a_11525_6580# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1925 VDD a_11575_3246# x4.x5.D VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1926 a_19054_5707# x4.x9.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1927 a_21446_5707# x4.x11.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X1928 a_12079_n656# a_11614_n964# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1929 VSS x2.x1.x4.Y a_11824_12152# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1930 VSS VDD a_19266_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X1931 a_3051_9193# sar_clk a_2979_9193# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1932 VSS a_18317_n1653# vss_sw_b[3] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1933 a_11858_n656# a_11440_n572# a_11614_n964# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X1934 x1.x2.x9.output_stack async_setb_delay_cap_ctrl_code[2] x1.x2.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X1935 a_9514_892# x4.x3.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1936 VSS a_11883_7842# sample_clk_b VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1937 VDD a_13898_892# x4.x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1938 a_17644_4145# a_16307_4145# a_17535_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X1939 VSS x3.x5.X a_18700_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1940 VDD x4.D[6] a_12913_n1627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1941 VDD a_16398_n964# a_16308_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X1942 VSS a_13264_892# x4.x30.A VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1943 x2.x2.x3.x9.output_stack sample_delay_cap_ctrl_code[14] x2.x2.x3.x4[3].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X1944 a_20613_n1475# a_20709_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1945 VDD a_22297_4992# a_22230_5384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X1946 a_12728_3246# a_11983_3272# a_12864_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1947 x2.x2.x4.x3[1].floating sample_delay_cap_ctrl_code[1] x2.x2.x4.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X1948 VDD a_28617_3118# a_28527_3510# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X1949 a_19270_10009# x2.x2.x3.IN VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X1950 VSS a_15318_5681# a_16025_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1951 a_18226_3272# a_17308_3246# a_17780_3456# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1952 a_21712_4119# a_21538_4511# a_21852_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X1953 a_16715_n1627# a_15925_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X1954 a_28162_1864# a_27996_1864# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1955 VDD a_14387_n1353# a_14388_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1956 a_11160_n938# a_10994_n938# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1957 VDD a_19614_4119# a_20335_4427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X1958 x2.x2.x1.x5[7].floating x2.x2.x1.x10.Y x2.x2.x1.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X1959 VDD a_9808_n1653# a_9741_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X1960 VSS a_9514_892# x4.x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1961 a_19146_4511# a_18699_4145# a_19053_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1962 a_28162_3790# a_27996_3790# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1963 x3.x7.X a_11392_4144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1964 a_11061_8554# a_10549_8788# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X1965 VSS a_8880_892# x4.x3.X VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1966 a_21646_4145# a_21257_4145# a_21538_4511# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X1967 a_24905_n250# x4.x9.A1 a_24684_77# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X1968 a_16967_3554# a_16767_3272# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X1969 VDD a_19615_5681# a_20336_5989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X1970 sar_result[6] a_27713_1864# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1971 a_21853_5707# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X1972 VSS a_9514_892# x4.x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1973 x3.x66.Q_N a_22493_4119# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X1974 VDD x3.x5.X a_18700_5707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1975 VDD a_15925_n1653# vss_sw_b[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X1976 a_19512_n1627# a_19644_n1443# a_19376_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X1977 VDD a_12145_5681# a_12055_6073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X1978 x2.x3.Y x2.x3.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1979 a_11141_n1653# a_11687_n1459# a_11645_n1345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X1980 a_17243_3272# a_16454_3246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X1981 x4.x2.X a_9514_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1982 a_21647_n656# a_21182_n964# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X1983 a_22225_5707# a_21713_5681# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X1984 a_17536_5707# a_16308_5707# a_17394_5989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X1985 a_11348_n938# x4.D[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1986 a_22028_5384# a_21239_4992# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X1987 VSS a_8653_n1475# vss_sw[7] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1988 x4.x2.X a_9514_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1989 VSS x2.x2.x1.IN a_20576_11016# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X1990 VDD a_19701_4992# a_19700_5292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1991 a_20728_n938# a_20562_n938# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1992 a_13435_n98# x4.x9.A1 a_13577_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1993 a_16286_77# x4.x9.A1 a_15827_n98# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X1994 VDD a_13898_892# x4.x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1995 x2.x2.x4.x10.Y sample_delay_cap_ctrl_code[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1996 a_22320_5707# a_21092_5707# a_22178_5989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X1997 VSS a_11974_5018# x3.x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1998 a_16779_n1353# x4.x13.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1999 a_28162_1864# a_27996_1864# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2000 a_21551_3272# x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2001 a_13939_11430# x2.x3.A a_13867_11568# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2002 a_12926_5681# a_12752_5707# a_13042_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X2003 VDD a_19614_4119# a_19564_4427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X2004 a_16662_5707# x4.x7.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2005 a_21022_n1627# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X2006 VDD a_22494_5681# a_22406_6073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X2007 VDD a_13898_892# x4.x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2008 VSS a_18751_3246# x4.D[4] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2009 a_2979_11093# ready a_2891_11093# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2010 a_26365_1864# a_26519_1838# a_26225_1838# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2011 VSS a_13898_892# x4.x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2012 VDD a_19615_5681# a_19565_5989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X2013 VSS a_14063_4992# x3.x48.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2014 a_19905_4992# a_20173_5202# a_20119_5300# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X2015 VDD a_19558_n670# a_20279_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2016 a_3051_9469# sar_clk a_2979_9469# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2017 a_24664_5133# x5.eob a_24592_5271# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2018 VSS a_22093_4992# a_22092_5292# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2019 a_28617_3118# a_28443_3510# a_28757_3144# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X2020 a_20173_5202# a_19701_4992# a_20417_5384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X2021 a_22319_4145# a_21257_4145# a_22224_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X2022 VSS a_12926_5681# a_13633_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2023 VSS x4.x11.S a_15335_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X2024 VSS x4.x17.S a_13456_6580# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0786 ps=0.805 w=0.42 l=0.15
X2025 VSS a_16984_n1653# a_16894_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X2026 VSS a_19321_5681# a_19255_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X2027 a_22494_5681# a_22320_5707# a_22610_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X2028 a_19558_n670# a_19399_n572# a_19698_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X2029 x2.x3.A a_13018_11968# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2030 VDD a_21713_5681# a_21623_6073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X2031 a_17513_4992# a_16768_5018# a_17649_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2032 a_25770_1864# a_25604_1864# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2033 a_28350_3144# x4.D[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2034 x4.x15.X a_19900_77# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X2035 x4.x30.A a_13264_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2036 a_16754_4511# a_16307_4145# a_16661_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2037 VDD a_13968_4992# x3.x48.Q VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2038 a_25770_3790# a_25604_3790# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2039 a_13240_3638# a_12728_3246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X2040 x1.x2.x5[7].floating x1.x2.x10.Y x1.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X2041 VSS a_16928_4119# a_16862_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X2042 x3.x4.X a_11974_5018# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2043 VSS a_23432_n276# a_23366_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2044 x2.x2.x3.x9.output_stack sample_delay_cap_ctrl_code[12] x2.x2.x3.x2.floating VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.43 as=0.122 ps=1.42 w=0.42 l=0.15
X2045 x3.x69.Q_N a_20101_4119# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X2046 x1.x9.Y x1.x9.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2047 a_15056_5018# a_14916_5292# a_14618_4992# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X2048 a_10345_8772# sample_clk VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2049 VSS x4.D[5] a_15305_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2050 x4.x7.S a_16025_5707# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2051 a_12459_3638# a_11670_3246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X2052 VSS x3.x7.X a_18226_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2053 x2.x2.x1.x9.output_stack x2.x2.x1.x10.Y x2.x2.x1.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X2054 VSS a_9514_892# x4.x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2055 a_14851_3272# a_14062_3246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X2056 a_19342_9871# x2.x2.x3.IN a_19270_10009# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2057 VDD a_13898_892# x4.x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2058 a_11075_11958# a_10909_11958# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2059 a_21552_5018# x3.x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X2060 a_16256_n276# x4.x13.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2061 VSS async_delay_offset x1.x4.x6.SW VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2062 VSS a_11472_n276# a_11406_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2063 a_29082_3784# a_28617_3758# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X2064 a_26051_9595# x2.x2.x2.IN a_25979_9595# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2065 x3.x4.A a_11360_5018# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2066 a_28861_3784# a_28443_3784# a_28617_3758# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X2067 a_10957_7987# VSS a_11099_7835# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2068 a_16928_4119# x3.x45.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X2069 VSS ready a_2979_10541# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2070 a_17536_5707# a_16474_5707# a_17441_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X2071 a_25770_1864# a_25604_1864# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2072 a_22808_3638# a_22296_3246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X2073 VSS x4.x13.S a_17254_77# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X2074 a_26918_2504# a_25770_2510# a_26832_2882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X2075 x2.x2.x2.x9.output_stack x2.x2.x2.x10.Y x2.x2.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X2076 VDD x4.x10.X a_13386_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2077 x3.x27.Q_N a_15318_5681# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X2078 VSS a_21144_4992# x4.x15.S VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2079 x5.eob a_12852_6554# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.218 ps=1.97 w=0.65 l=0.15
X2080 a_26737_3144# a_26225_3118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X2081 a_22320_5707# a_21258_5707# a_22225_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X2082 a_29514_2870# a_28911_2704# a_29398_2478# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2083 a_26386_12370# x2.x2.x1.x9.output_stack VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2084 a_11440_n572# a_11160_n938# a_11348_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X2085 a_24617_6660# x5.eob a_24529_6798# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2086 vdd_sw[3] a_20279_n938# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2087 VSS a_19701_4992# a_19700_5292# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2088 a_17172_4427# a_16754_4511# a_16928_4119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X2089 a_2979_11369# ready a_2891_11369# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2090 VSS x3.x4.X a_19615_5681# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2091 a_16917_n1261# a_16780_n1653# a_16471_n1459# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X2092 VSS VDD a_16692_n964# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2093 a_11454_n1627# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2094 a_26832_2882# a_25770_2510# a_26737_2826# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X2095 a_29398_1838# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X2096 x1.x4.x9.output_stack async_resetb_delay_cap_ctrl_code[1] x1.x4.x3[1].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X2097 VDD x4.D[1] a_21091_4145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2098 a_17173_5989# a_16755_6073# a_16929_5681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X2099 a_24664_5409# x5.eob a_24592_5547# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2100 VSS a_18790_n964# a_18724_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X2101 x2.x2.x2.x5[7].floating x2.x2.x2.x10.Y x2.x2.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X2102 x3.x4.X a_11974_5018# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2103 sar_result[5] a_30105_2520# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2104 x5.x1[2].Q_N a_27006_3118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X2105 VSS x4.D[2] a_22481_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2106 a_14082_5707# a_13916_5707# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2107 a_19698_n938# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X2108 VSS a_11801_6580# x3.x5.X VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2109 a_8956_n938# x4.x5.D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2110 a_15969_77# x4.x13.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X2111 a_14916_3246# x4.D[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2112 x3.x36.Q_N a_22494_5681# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2113 VSS x3.x33.Q_N a_20040_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X2114 x3.x27.D a_13633_5707# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2115 VSS a_13898_892# x4.x9.A1 VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2116 a_21040_n276# x4.x17.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X2117 a_16838_4511# a_16307_4145# a_16754_4511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X2118 x2.x2.x4.x5[7].floating x2.x2.x4.x10.Y x2.x2.x4.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X2119 a_9718_n1627# a_9603_n1353# a_9295_n1459# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X2120 VDD VDD a_16984_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X2121 VDD a_26225_2478# a_26135_2504# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X2122 a_21793_3246# a_22091_3546# a_22027_3638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X2123 VSS a_12852_6554# x5.eob VSS sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X2124 a_26159_4162# a_25770_3790# a_26051_3784# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X2125 a_29333_1864# a_27996_1864# a_29224_1864# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X2126 a_20601_13233# x2.x2.x1.IN a_20513_13371# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2127 a_21622_4511# a_21091_4145# a_21538_4511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X2128 a_26690_3784# a_26225_3758# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X2129 a_11464_12330# a_11075_11958# a_11356_11952# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X2130 VDD x3.x30.Q_N a_17512_3246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X2131 a_14536_4119# x3.x77.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X2132 VDD x4.x30.A a_13898_892# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2133 VSS a_15121_4992# a_15056_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X2134 x5.x2.x9.output_stack x5.x2.x10.Y x5.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X2135 a_27006_3118# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X2136 a_14082_5707# a_13916_5707# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2137 VSS x5.eob a_24592_4719# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2138 a_16779_n1353# x4.x13.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2139 a_28617_3758# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X2140 a_30402_6073# x5.x2.x9.output_stack VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2141 VSS x5.x3.A a_30402_6073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X2142 a_9396_8528# a_9491_8544# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2143 VDD sample_delay_offset x2.x2.x4.x6.SW VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2144 a_3051_10679# ready a_2979_10817# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2145 VDD sample_clk_b a_11084_5018# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2146 a_12285_5707# a_12439_5681# a_12145_5681# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2147 a_9222_n964# a_9048_n572# a_9366_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X2148 x4.x2.X a_9514_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2149 VDD x5.x3.X a_27996_3144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2150 VSS sample_delay_cap_ctrl_code[11] x2.x2.x2.x10.Y VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2151 x4.x3.X a_8880_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2152 a_29632_3784# a_29224_4162# a_29398_3758# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X2153 a_14780_4427# a_14362_4511# a_14536_4119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X2154 VDD a_20101_4119# a_20013_4511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X2155 VDD a_23432_n276# a_23462_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2156 a_9156_n938# a_8602_n938# a_9048_n572# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X2157 a_18221_n1475# a_18317_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X2158 a_21238_3246# a_21551_3272# a_21657_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2159 a_14781_5989# a_14363_6073# a_14537_5681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X2160 x5.x2.x5[7].floating x5.x2.x10.Y x5.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X2161 a_26832_3144# a_25770_3144# a_26737_3144# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X2162 a_26026_7516# x2.x2.x2.IN a_25938_7654# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2163 a_14150_n938# a_14300_n964# a_14006_n964# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2164 a_23308_n938# x4.D[1] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2165 a_11690_5707# a_11524_5707# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2166 a_18227_5018# a_17308_5292# a_17781_5202# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2167 x4.x2.X a_9514_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2168 VDD VDD a_24160_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X2169 a_24342_n670# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X2170 x3.x33.Q_N a_20102_5681# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2171 vdd_sw_b[4] a_17166_n670# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2172 VDD x4.x15.S a_19646_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X2173 VDD x4.x11.S a_15328_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X2174 x2.x1.x3.Y VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2175 a_9831_n572# a_8768_n938# a_9687_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X2176 a_14699_n572# a_13386_n938# a_14615_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X2177 a_20576_11430# x2.x2.x1.IN a_20488_11292# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2178 a_28527_3510# a_27996_3144# a_28443_3510# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X2179 VSS x4.D[1] a_21091_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2180 VDD a_13898_892# x4.x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2181 VDD a_11670_3246# x3.x51.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X2182 a_13867_11982# x2.x3.A a_13779_11844# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2183 a_13247_6902# x4.x15.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=0.995 as=0.154 ps=1.34 w=0.64 l=0.15
X2184 a_21658_5018# a_21794_4992# a_21239_4992# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X2185 a_14914_n938# a_14300_n964# a_14774_n670# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2186 x5.x2.x3[1].floating retimer_delay_code[1] x5.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X2187 a_21144_4992# a_21239_4992# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X2188 a_26941_1864# a_25604_1864# a_26832_1864# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X2189 a_24592_5133# x5.eob a_24504_4995# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2190 VSS a_29398_1838# a_29333_1864# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X2191 a_25958_1864# x4.D[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2192 a_10247_n656# a_9831_n572# a_9990_n670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X2193 a_16929_5681# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X2194 a_23718_n938# a_23868_n964# a_23574_n964# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2195 VSS x4.x30.A a_13898_892# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2196 VSS a_29398_3758# a_29333_4162# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X2197 a_25958_3784# x3.D[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2198 a_11974_5018# x3.x4.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2199 VSS VDD a_16874_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X2200 a_9514_892# x4.x3.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2201 a_14362_4511# a_14081_4145# a_14269_4145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X2202 a_20089_n1627# a_19171_n1353# a_19644_n1443# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X2203 a_18361_n250# x4.x15.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X2204 a_11690_5707# a_11524_5707# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2205 a_23605_n1345# a_23414_n1627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X2206 a_28443_3784# a_28162_3790# a_28350_3784# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X2207 a_22565_5202# a_22092_5292# a_22809_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X2208 a_17825_4145# x3.x45.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X2209 VDD x4.D[4] a_17697_n1627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2210 a_13435_n98# VSS a_13577_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X2211 VDD a_27006_3118# a_26918_3510# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X2212 VSS a_17308_3246# a_17307_3546# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2213 a_20102_5681# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X2214 VDD a_29398_3758# a_30105_3800# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2215 x1.x2.x5[7].floating x1.x2.x10.Y x1.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X2216 VSS a_8651_n98# x4.x6.X VSS sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X2217 VDD VDD a_20709_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X2218 a_17825_4145# a_17222_4119# a_17709_4119# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2219 a_28443_2230# a_27996_1864# a_28350_1864# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2220 VDD x5.x3.X a_25604_3144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2221 a_17726_3554# a_16767_3272# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X2222 x2.x2.x2.x5[7].floating x2.x2.x2.x10.Y x2.x2.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X2223 a_19342_9595# x2.x2.x3.IN a_19270_9595# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2224 a_22433_5018# a_22565_5202# a_22297_4992# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X2225 VSS a_28617_1838# a_28551_1864# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X2226 VSS x4.x3.X a_9514_892# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2227 x4.x2.X a_9514_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2228 x4.x30.A a_13264_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2229 VSS a_28617_3758# a_28551_4162# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X2230 a_12610_5989# a_12145_5681# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X2231 VDD x4.x11.S a_14860_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X2232 a_26832_1864# a_25604_1864# a_26690_2146# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X2233 x2.x2.x3.x9.output_stack x2.x2.x3.x10.Y x2.x2.x3.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X2234 a_18790_n964# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X2235 x4.D[2] a_23200_4145# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X2236 a_10076_n1443# a_9603_n1353# a_10320_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X2237 VDD a_14006_n964# a_13916_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X2238 x2.x2.x4.x5[7].floating x2.x2.x4.x10.Y x2.x2.x4.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X2239 x4.x2.X a_9514_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2240 a_15104_n1627# a_14592_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X2241 a_12427_12318# x2.x1.x3.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X2242 VSS x2.x7.A x2.x7.Y VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2243 a_24482_n938# a_23868_n964# a_24342_n670# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2244 a_20916_n938# x4.D[2] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2245 VDD x4.x20.S a_24898_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X2246 VSS x5.x3.X a_27996_3144# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2247 VSS VDD a_19512_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X2248 VDD a_13898_892# x4.x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2249 a_15551_4427# a_15143_4145# a_15317_4119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X2250 a_12246_12330# a_10909_11958# a_12137_12330# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X2251 a_24183_n572# a_23120_n938# a_24039_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X2252 VDD VDD a_8749_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X2253 x4.x30.A a_13264_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2254 a_27122_4150# a_26519_3984# a_27006_3758# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2255 a_20417_5384# a_19905_4992# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X2256 a_15925_n1653# a_16471_n1459# a_16429_n1345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X2257 x2.x2.x1.x9.output_stack x2.x2.x1.IN a_20513_12819# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2258 a_16839_6073# a_16308_5707# a_16755_6073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X2259 VDD async_delay_offset x1.x2.x6.SW VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2260 x4.x17.X a_22290_77# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X2261 a_15552_5989# a_15144_5707# a_15318_5681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X2262 a_24672_n1627# a_24160_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X2263 a_9808_n1653# a_10076_n1443# a_10022_n1345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X2264 x3.x7.X a_11392_4144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2265 x2.x1.x4.Y VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2266 x2.x2.x3.x5[7].floating x2.x2.x3.x10.Y x2.x2.x3.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X2267 x5.x2.x9.output_stack x5.x2.x10.Y x5.x2.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X2268 a_12522_n938# a_11908_n964# a_12382_n670# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2269 a_21623_6073# a_21092_5707# a_21539_6073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X2270 a_20576_11706# x2.x2.x1.IN a_20488_11568# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2271 a_14063_4992# a_14376_5018# a_14482_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2272 a_12223_n572# a_11160_n938# a_12079_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X2273 a_15253_5707# a_13916_5707# a_15144_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X2274 a_17114_n938# a_15944_n938# a_17007_n572# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X2275 a_14537_5681# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X2276 a_19107_n1627# a_18317_n1653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X2277 a_11974_5018# x3.x4.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2278 VDD x4.D[1] a_24873_n1627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2279 a_3004_7942# sar_clk a_2916_8080# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2280 VSS VDD a_14482_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X2281 a_16190_n250# VSS a_15827_n98# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X2282 VSS a_16359_3246# x4.D[5] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2283 a_14111_6878# x3.x48.Q VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.164 pd=1.33 as=0.0864 ps=0.91 w=0.64 l=0.15
X2284 a_24684_77# VSS a_24684_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2285 a_24592_5409# x5.eob a_24504_5271# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2286 a_16398_n964# a_16224_n572# a_16542_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X2287 VDD x4.x13.S a_23011_5018# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X2288 VSS x3.x5.X a_13916_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2289 a_20648_11430# x2.x2.x1.IN a_20576_11430# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2290 a_10553_n250# x4.x9.A1 a_10332_77# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X2291 VSS a_29398_2478# a_30105_2520# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2292 x5.x1[0].Q_N a_27006_3758# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X2293 a_21182_n964# a_21008_n572# a_21326_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X2294 x2.x2.x4.x9.output_stack x2.x3.A a_13867_11982# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2295 a_9804_8920# x1.x10.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X2296 a_12110_n1627# a_11995_n1353# a_11687_n1459# VSS sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X2297 a_13533_n1653# a_14079_n1459# a_14037_n1345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X2298 VDD a_20102_5681# a_20014_6073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X2299 a_19839_3272# a_19699_3546# a_19401_3246# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X2300 x3.x4.X a_11974_5018# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2301 a_12724_77# VSS a_12724_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2302 x4.x9.A1 a_13898_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2303 a_16359_3246# a_16454_3246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X2304 VDD a_14916_3246# a_14915_3546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2305 VSS ext_clk a_10909_11958# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2306 x2.x2.x1.x9.output_stack sample_delay_cap_ctrl_code[5] x2.x2.x1.x3[1].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X2307 a_21116_n938# a_20562_n938# a_21008_n572# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X2308 VDD x4.x3.A a_8880_892# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2309 VDD a_19905_4992# a_19838_5384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X2310 VDD a_22006_4119# a_21956_4427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X2311 x4.D[1] a_20808_4145# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X2312 a_15121_4992# a_14376_5018# a_15257_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2313 VDD a_11614_n964# a_11524_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X2314 a_19832_4145# a_19320_4119# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X2315 VSS a_15317_4119# a_15252_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X2316 a_22036_n1443# a_21564_n1653# a_22280_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X2317 a_18616_n572# a_18170_n938# a_18524_n938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X2318 x4.x9.A1 a_13898_892# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2319 a_13892_12957# x2.x3.A a_13804_13095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2320 a_3051_9745# sar_clk a_2979_9883# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2321 a_10549_8788# a_9804_8920# a_10685_8876# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2322 VDD a_9516_n964# a_9466_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X2323 VDD a_22007_5681# a_21957_5989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X2324 a_23101_n1653# a_23647_n1459# a_23605_n1345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X2325 VDD a_17709_4119# a_18416_4145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2326 a_19905_4992# a_19160_5018# a_20041_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2327 a_23414_n1627# x4.x2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X2328 VSS x5.x3.X a_25604_3144# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2329 a_13240_3272# a_12728_3246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X2330 sample_clk_b a_11883_7842# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X2331 a_29129_4106# a_28617_3758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X2332 VSS sample_delay_cap_ctrl_code[15] x2.x2.x3.x10.Y VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2333 a_20611_n98# x4.x9.A1 a_20753_n250# VSS sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2334 VDD VDD a_15121_4992# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X2335 a_26051_2504# a_25604_2510# a_25958_2504# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2336 VDD x3.x5.X a_13916_5707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2337 VDD a_17222_4119# a_17943_4427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X2338 a_21791_n572# a_20728_n938# a_21647_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X2339 a_18678_77# x4.x9.A1 a_18219_n98# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X2340 VDD a_15120_3246# a_15053_3638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X2341 a_13442_3272# a_12524_3246# a_12996_3456# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2342 a_12459_3272# a_11670_3246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X2343 VSS a_11801_6580# x3.x5.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2344 a_20102_5681# a_19928_5707# a_20218_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X2345 VDD VDD a_26519_2704# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X2346 a_19270_9181# x2.x2.x3.IN a_19182_9181# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2347 VDD a_17223_5681# a_17944_5989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X2348 a_9808_n1653# a_9062_n1627# a_9944_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2349 a_12311_11926# x2.x1.x3.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X2350 a_13316_6554# sel_bit[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2351 VSS a_21239_4992# x3.x39.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2352 a_29082_2504# a_28617_2478# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X2353 x1.x2.x5[7].floating x1.x2.x10.Y x1.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X2354 x3.x4.X a_11974_5018# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2355 a_26469_3784# a_26051_3784# a_26225_3758# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X2356 a_28861_2504# a_28443_2504# a_28617_2478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X2357 VSS a_19376_n1653# a_19286_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X2358 VDD a_29398_1838# a_30105_1864# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2359 VDD VDD a_26519_3118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X2360 a_12137_12330# a_11075_11958# a_12042_12274# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X2361 a_12861_5707# a_11524_5707# a_12752_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X2362 VSS a_9514_892# x4.x2.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2363 a_14722_n938# a_13552_n938# a_14615_n572# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X2364 a_11878_5707# x5.eob VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2365 a_14363_6073# a_14082_5707# a_14270_5707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X2366 a_19900_77# x4.x9.A1 a_19828_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2367 VDD a_16256_n276# a_16286_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2368 a_22808_3272# a_22296_3246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X2369 a_21238_3246# a_21793_3246# a_21751_3554# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X2370 a_19265_3272# a_19401_3246# a_18846_3246# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X2371 VSS a_13967_3246# x4.D[6] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2372 VSS a_17166_n670# a_17887_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2373 VSS a_12261_7986# a_11883_7842# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2374 VDD x4.x15.S a_20619_5018# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X2375 VDD x4.x30.A a_13898_892# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2376 x2.x2.x4.x5[7].floating x2.x2.x4.x10.Y x2.x2.x4.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X2377 a_15834_3272# a_14915_3546# a_15388_3456# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2378 a_12414_n1345# a_11454_n1627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X2379 x1.x4.x9.output_stack x1.x4.x10.Y x1.x4.x5[7].floating VDD sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X2380 a_13867_11154# x2.x3.A a_13779_11016# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2381 a_20618_3272# a_19699_3546# a_20172_3456# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2382 a_14363_6073# a_13916_5707# a_14270_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2383 a_20648_11706# x2.x2.x1.IN a_20576_11706# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2384 a_16359_3246# a_16454_3246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2385 a_17513_4992# a_17781_5202# a_17727_5300# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X2386 VDD a_12524_3246# a_12523_3546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2387 a_3004_12758# ready a_2916_12896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2388 x4.x13.S a_23201_5707# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2389 VSS a_14537_5681# a_14471_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X2390 VSS x4.D[6] a_12913_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2391 VSS a_16398_n964# a_16332_n938# VSS sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X2392 a_10817_8528# a_10345_8772# a_11061_8554# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X2393 x1.x2.x9.output_stack async_setb_delay_cap_ctrl_code[1] x1.x2.x3[1].floating VSS sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X2394 a_21982_n1345# a_21022_n1627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X2395 a_19927_4145# a_18865_4145# a_19832_4145# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X2396 x5.x1[6].Q_N a_27006_1838# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X2397 VDD x1.x10.A a_8789_8870# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X2398 x1.x4.x2.floating async_resetb_delay_cap_ctrl_code[0] x1.x4.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X2399 a_10345_8772# sample_clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2400 a_18648_n276# x4.x15.S VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2401 a_29398_3758# a_29224_4162# a_29514_4150# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X2402 VDD a_28911_1838# a_28861_2146# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X2403 VSS VDD a_26519_2704# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2404 vdd_sw[1] a_25063_n938# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X2405 a_18227_5018# a_17309_4992# a_17781_5202# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2406 a_29310_3784# a_28162_3790# a_29224_4162# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X2407 VSS a_19904_3246# a_19839_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X2408 x1.x4.x5[7].floating x1.x4.x10.Y x1.x4.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X2409 a_11670_12318# x2.x1.x3.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X2410 VDD a_12728_3246# a_12661_3638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X2411 VSS a_9396_8528# x1.x3.A0 VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2412 a_26051_3510# a_25604_3144# a_25958_3144# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2413 x5.x1[1].Q_N a_29398_3758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2414 VSS VDD a_11560_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X2415 a_29514_1864# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X2416 a_19309_n1261# a_19172_n1653# a_18863_n1459# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X2417 a_9514_892# x4.x3.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2418 VSS a_26225_3118# a_26159_3144# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X2419 VDD sar_clk a_2916_7528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2420 vdd_sw[6] a_13103_n938# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X2421 a_26690_2504# a_26225_2478# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X2422 a_29514_4150# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X2423 a_29514_1864# a_28911_1838# a_29398_1838# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2424 x2.x1.x2.D a_12311_11926# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X2425 a_9804_8920# x1.x10.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2426 a_9944_n1627# a_10076_n1443# a_9808_n1653# VSS sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X2427 a_17244_5018# a_16455_4992# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X2428 a_22090_n938# x4.x2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X2429 a_19270_9457# x2.x2.x3.IN a_19182_9457# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2430 a_17496_n1261# a_16984_n1653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X2431 a_17068_4145# a_17222_4119# a_16928_4119# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2432 a_11971_6073# a_11690_5707# a_11878_5707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X2433 VSS VDD a_18736_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X2434 VSS x4.x9.S a_12470_77# VSS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X2435 a_28617_2478# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X2436 a_12225_3246# a_12524_3246# a_12459_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X2437 a_11320_7835# x1.x3.A0 a_10957_7987# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X2438 a_9514_892# x4.x3.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2439 VSS a_13264_892# x4.x30.A VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2440 x2.x3.Y VSS a_12261_7986# VDD sky130_fd_pr__pfet_01v8 ad=0.551 pd=4.38 as=0.551 ps=4.38 w=1.9 l=0.15
X2441 x4.x2.X a_9514_892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2442 a_2979_10955# ready a_2891_10817# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X2443 VDD x1.x9.Y a_10549_8788# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X2444 a_21552_5018# x3.x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2445 VDD a_24342_n670# a_24267_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X2446 VDD x4.x13.S a_17722_77# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X2447 a_21258_5707# a_21092_5707# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2448 a_18336_n938# a_18170_n938# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2449 VDD a_15827_n98# x4.x12.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X2450 a_29632_2504# a_29224_2882# a_29398_2478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X2451 VDD a_26519_3118# a_26469_3426# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X2452 VSS a_18752_4992# x4.x17.S VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2453 a_22092_3246# x4.D[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2454 a_11971_6073# a_11524_5707# a_11878_5707# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2455 VDD x3.x33.Q_N a_19904_3246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X2456 a_11530_11926# a_11356_11952# a_11670_12318# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X2457 a_12389_5989# a_11971_6073# a_12145_5681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X2458 a_23120_n938# a_22954_n938# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2459 a_22296_3246# a_22564_3456# a_22510_3554# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X2460 x2.x2.x2.x4[3].floating sample_delay_cap_ctrl_code[10] x2.x2.x2.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X2461 x4.x11.S a_20809_5707# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2462 a_12996_3456# a_12524_3246# a_13240_3638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X2463 a_14917_4992# x3.x5.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2464 VDD a_13898_892# x4.x9.A1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2465 a_28617_2478# a_28443_2504# a_28757_2870# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X2466 VDD VDD a_14592_n1653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X2467 a_16471_n1459# a_16779_n1353# a_16728_n1261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X2468 VDD a_12382_n670# a_12307_n572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X2469 VDD a_21476_n964# a_21426_n656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X2470 a_21255_n1459# a_21564_n1653# a_21499_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X2471 a_26225_1838# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X2472 VDD x2.x2.x1.IN a_19677_12029# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X2473 VSS VDD a_16344_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X2474 VDD x3.D[0] a_18699_4145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2475 x1.x2.x5[7].floating x1.x2.x10.Y x1.x2.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X2476 vdd_sw_b[5] a_14774_n670# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2477 VDD sel_bit[1] a_13721_6554# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2478 a_21712_4119# x3.x39.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X2479 sar_result[4] a_27713_2520# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2480 VSS x1.x9.A a_8789_11895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X2481 a_13939_11154# x2.x3.A a_13867_11154# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2482 VSS x2.x7.Y a_12758_8861# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2483 a_21258_5707# a_21092_5707# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2484 VSS sar_clk a_2979_10021# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2485 vdd_sw_b[3] a_19558_n670# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X2486 a_19677_12370# x2.x2.x4.x9.output_stack x2.x2.x1.IN VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X2487 VSS x3.x30.Q_N a_17648_3272# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X2488 x2.x2.x4.x5[7].floating x2.x2.x4.x10.Y x2.x2.x4.x9.output_stack VDD sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X2489 a_22564_3456# a_22092_3246# a_22808_3638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X2490 a_18648_n276# x4.x15.S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X2491 VSS VDD a_28911_3118# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2492 a_22177_4427# a_21712_4119# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X2493 VSS x4.x17.S a_18227_5018# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2494 a_10521_n1627# a_9603_n1353# a_10076_n1443# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X2495 a_14852_5018# a_14063_4992# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X2496 a_9295_n1459# a_9604_n1653# a_9539_n1627# VSS sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X2497 a_19401_3246# a_19699_3546# a_19635_3638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X2498 VSS sample_delay_offset x2.x2.x1.x6.SW VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2499 a_21956_4427# a_21538_4511# a_21712_4119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X2500 a_14676_4145# a_14830_4119# a_14536_4119# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2501 a_11356_11952# a_10909_11958# a_11263_11952# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2502 x1.x4.x9.output_stack sar_clk a_2979_9055# VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X2503 x1.x4.x4[3].floating async_resetb_delay_cap_ctrl_code[2] x1.x4.x9.output_stack VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X2504 a_26135_3510# a_25604_3144# a_26051_3510# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

