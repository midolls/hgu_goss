magic
tech sky130A
magscale 1 2
timestamp 1699094131
<< pwell >>
rect 312 2604 338 2636
rect 306 1080 332 1112
<< psubdiff >>
rect 300 2029 348 2143
<< metal3 >>
rect -14 3050 658 3052
rect -14 2986 90 3050
rect 154 2986 170 3050
rect 234 2986 250 3050
rect 314 2986 330 3050
rect 394 2986 410 3050
rect 474 2986 490 3050
rect 554 2986 658 3050
rect -14 2984 658 2986
rect -14 2830 52 2920
rect -14 2766 -13 2830
rect 51 2766 52 2830
rect -14 2750 52 2766
rect -14 2686 -13 2750
rect 51 2686 52 2750
rect -14 2670 52 2686
rect -14 2606 -13 2670
rect 51 2606 52 2670
rect -14 2590 52 2606
rect -14 2526 -13 2590
rect 51 2526 52 2590
rect -14 2510 52 2526
rect -14 2446 -13 2510
rect 51 2446 52 2510
rect -14 2430 52 2446
rect -14 2366 -13 2430
rect 51 2366 52 2430
rect -14 2350 52 2366
rect -14 2286 -13 2350
rect 51 2286 52 2350
rect -14 2270 52 2286
rect -14 2206 -13 2270
rect 51 2206 52 2270
rect -14 2190 52 2206
rect -14 2126 -13 2190
rect 51 2126 52 2190
rect -14 2110 52 2126
rect -14 2046 -13 2110
rect 51 2046 52 2110
rect -14 1892 52 2046
rect 112 1954 172 2984
rect 232 1892 292 2924
rect 352 1954 412 2984
rect 472 1892 532 2924
rect 592 2830 658 2920
rect 592 2766 593 2830
rect 657 2766 658 2830
rect 592 2750 658 2766
rect 592 2686 593 2750
rect 657 2686 658 2750
rect 592 2670 658 2686
rect 592 2606 593 2670
rect 657 2606 658 2670
rect 592 2590 658 2606
rect 592 2526 593 2590
rect 657 2526 658 2590
rect 592 2510 658 2526
rect 592 2446 593 2510
rect 657 2446 658 2510
rect 592 2430 658 2446
rect 592 2366 593 2430
rect 657 2366 658 2430
rect 592 2350 658 2366
rect 592 2286 593 2350
rect 657 2286 658 2350
rect 592 2270 658 2286
rect 592 2206 593 2270
rect 657 2206 658 2270
rect 592 2190 658 2206
rect 592 2126 593 2190
rect 657 2126 658 2190
rect 592 2110 658 2126
rect 592 2046 593 2110
rect 657 2046 658 2110
rect 592 1892 658 2046
rect -14 1890 658 1892
rect -14 1826 90 1890
rect 154 1826 170 1890
rect 234 1826 250 1890
rect 314 1826 330 1890
rect 394 1826 410 1890
rect 474 1826 490 1890
rect 554 1826 658 1890
rect -14 1824 658 1826
rect -14 1670 52 1824
rect -14 1606 -13 1670
rect 51 1606 52 1670
rect -14 1590 52 1606
rect -14 1526 -13 1590
rect 51 1526 52 1590
rect -14 1510 52 1526
rect -14 1446 -13 1510
rect 51 1446 52 1510
rect -14 1430 52 1446
rect -14 1366 -13 1430
rect 51 1366 52 1430
rect -14 1350 52 1366
rect -14 1286 -13 1350
rect 51 1286 52 1350
rect -14 1270 52 1286
rect -14 1206 -13 1270
rect 51 1206 52 1270
rect -14 1190 52 1206
rect -14 1126 -13 1190
rect 51 1126 52 1190
rect -14 1110 52 1126
rect -14 1046 -13 1110
rect 51 1046 52 1110
rect -14 1030 52 1046
rect -14 966 -13 1030
rect 51 966 52 1030
rect -14 950 52 966
rect -14 886 -13 950
rect 51 886 52 950
rect -14 796 52 886
rect 112 792 172 1824
rect 232 732 292 1762
rect 352 792 412 1824
rect 472 732 532 1762
rect 592 1670 658 1824
rect 592 1606 593 1670
rect 657 1606 658 1670
rect 592 1590 658 1606
rect 592 1526 593 1590
rect 657 1526 658 1590
rect 592 1510 658 1526
rect 592 1446 593 1510
rect 657 1446 658 1510
rect 592 1430 658 1446
rect 592 1366 593 1430
rect 657 1366 658 1430
rect 592 1350 658 1366
rect 592 1286 593 1350
rect 657 1286 658 1350
rect 592 1270 658 1286
rect 592 1206 593 1270
rect 657 1206 658 1270
rect 592 1190 658 1206
rect 592 1126 593 1190
rect 657 1126 658 1190
rect 592 1110 658 1126
rect 592 1046 593 1110
rect 657 1046 658 1110
rect 592 1030 658 1046
rect 592 966 593 1030
rect 657 966 658 1030
rect 592 950 658 966
rect 592 886 593 950
rect 657 886 658 950
rect 592 796 658 886
rect -14 730 658 732
rect -14 666 90 730
rect 154 666 170 730
rect 234 666 250 730
rect 314 666 330 730
rect 394 666 410 730
rect 474 666 490 730
rect 554 666 658 730
rect -14 664 658 666
<< via3 >>
rect 90 2986 154 3050
rect 170 2986 234 3050
rect 250 2986 314 3050
rect 330 2986 394 3050
rect 410 2986 474 3050
rect 490 2986 554 3050
rect -13 2766 51 2830
rect -13 2686 51 2750
rect -13 2606 51 2670
rect -13 2526 51 2590
rect -13 2446 51 2510
rect -13 2366 51 2430
rect -13 2286 51 2350
rect -13 2206 51 2270
rect -13 2126 51 2190
rect -13 2046 51 2110
rect 593 2766 657 2830
rect 593 2686 657 2750
rect 593 2606 657 2670
rect 593 2526 657 2590
rect 593 2446 657 2510
rect 593 2366 657 2430
rect 593 2286 657 2350
rect 593 2206 657 2270
rect 593 2126 657 2190
rect 593 2046 657 2110
rect 90 1826 154 1890
rect 170 1826 234 1890
rect 250 1826 314 1890
rect 330 1826 394 1890
rect 410 1826 474 1890
rect 490 1826 554 1890
rect -13 1606 51 1670
rect -13 1526 51 1590
rect -13 1446 51 1510
rect -13 1366 51 1430
rect -13 1286 51 1350
rect -13 1206 51 1270
rect -13 1126 51 1190
rect -13 1046 51 1110
rect -13 966 51 1030
rect -13 886 51 950
rect 593 1606 657 1670
rect 593 1526 657 1590
rect 593 1446 657 1510
rect 593 1366 657 1430
rect 593 1286 657 1350
rect 593 1206 657 1270
rect 593 1126 657 1190
rect 593 1046 657 1110
rect 593 966 657 1030
rect 593 886 657 950
rect 90 666 154 730
rect 170 666 234 730
rect 250 666 314 730
rect 330 666 394 730
rect 410 666 474 730
rect 490 666 554 730
<< metal4 >>
rect -14 3050 658 3052
rect -14 2986 90 3050
rect 154 2986 170 3050
rect 234 2986 250 3050
rect 314 2986 330 3050
rect 394 2986 410 3050
rect 474 2986 490 3050
rect 554 2986 658 3050
rect -14 2984 658 2986
rect -14 2830 52 2920
rect -14 2766 -13 2830
rect 51 2766 52 2830
rect -14 2750 52 2766
rect -14 2686 -13 2750
rect 51 2686 52 2750
rect -14 2670 52 2686
rect -14 2606 -13 2670
rect 51 2606 52 2670
rect -14 2590 52 2606
rect -14 2526 -13 2590
rect 51 2526 52 2590
rect -14 2510 52 2526
rect -14 2446 -13 2510
rect 51 2446 52 2510
rect -14 2430 52 2446
rect -14 2366 -13 2430
rect 51 2366 52 2430
rect -14 2350 52 2366
rect -14 2286 -13 2350
rect 51 2286 52 2350
rect -14 2270 52 2286
rect -14 2206 -13 2270
rect 51 2206 52 2270
rect -14 2190 52 2206
rect -14 2126 -13 2190
rect 51 2126 52 2190
rect -14 2110 52 2126
rect -14 2046 -13 2110
rect 51 2046 52 2110
rect -14 1892 52 2046
rect 112 1892 172 2924
rect 232 1954 292 2984
rect 352 1892 412 2924
rect 472 1954 532 2984
rect 592 2830 658 2920
rect 592 2766 593 2830
rect 657 2766 658 2830
rect 592 2750 658 2766
rect 592 2686 593 2750
rect 657 2686 658 2750
rect 592 2670 658 2686
rect 592 2606 593 2670
rect 657 2606 658 2670
rect 592 2590 658 2606
rect 592 2526 593 2590
rect 657 2526 658 2590
rect 592 2510 658 2526
rect 592 2446 593 2510
rect 657 2446 658 2510
rect 592 2430 658 2446
rect 592 2366 593 2430
rect 657 2366 658 2430
rect 592 2350 658 2366
rect 592 2286 593 2350
rect 657 2286 658 2350
rect 592 2270 658 2286
rect 592 2206 593 2270
rect 657 2206 658 2270
rect 592 2190 658 2206
rect 592 2126 593 2190
rect 657 2126 658 2190
rect 592 2110 658 2126
rect 592 2046 593 2110
rect 657 2046 658 2110
rect 592 1892 658 2046
rect -14 1890 658 1892
rect -14 1826 90 1890
rect 154 1826 170 1890
rect 234 1826 250 1890
rect 314 1826 330 1890
rect 394 1826 410 1890
rect 474 1826 490 1890
rect 554 1826 658 1890
rect -14 1824 658 1826
rect -14 1670 52 1824
rect -14 1606 -13 1670
rect 51 1606 52 1670
rect -14 1590 52 1606
rect -14 1526 -13 1590
rect 51 1526 52 1590
rect -14 1510 52 1526
rect -14 1446 -13 1510
rect 51 1446 52 1510
rect -14 1430 52 1446
rect -14 1366 -13 1430
rect 51 1366 52 1430
rect -14 1350 52 1366
rect -14 1286 -13 1350
rect 51 1286 52 1350
rect -14 1270 52 1286
rect -14 1206 -13 1270
rect 51 1206 52 1270
rect -14 1190 52 1206
rect -14 1126 -13 1190
rect 51 1126 52 1190
rect -14 1110 52 1126
rect -14 1046 -13 1110
rect 51 1046 52 1110
rect -14 1030 52 1046
rect -14 966 -13 1030
rect 51 966 52 1030
rect -14 950 52 966
rect -14 886 -13 950
rect 51 886 52 950
rect -14 796 52 886
rect 112 732 172 1762
rect 232 792 292 1824
rect 352 732 412 1762
rect 472 792 532 1824
rect 592 1670 658 1824
rect 592 1606 593 1670
rect 657 1606 658 1670
rect 592 1590 658 1606
rect 592 1526 593 1590
rect 657 1526 658 1590
rect 592 1510 658 1526
rect 592 1446 593 1510
rect 657 1446 658 1510
rect 592 1430 658 1446
rect 592 1366 593 1430
rect 657 1366 658 1430
rect 592 1350 658 1366
rect 592 1286 593 1350
rect 657 1286 658 1350
rect 592 1270 658 1286
rect 592 1206 593 1270
rect 657 1206 658 1270
rect 592 1190 658 1206
rect 592 1126 593 1190
rect 657 1126 658 1190
rect 592 1110 658 1126
rect 592 1046 593 1110
rect 657 1046 658 1110
rect 592 1030 658 1046
rect 592 966 593 1030
rect 657 966 658 1030
rect 592 950 658 966
rect 592 886 593 950
rect 657 886 658 950
rect 592 796 658 886
rect -14 730 658 732
rect -14 666 90 730
rect 154 666 170 730
rect 234 666 250 730
rect 314 666 330 730
rect 394 666 410 730
rect 474 666 490 730
rect 554 666 658 730
rect -14 664 658 666
<< labels >>
flabel psubdiff 300 2029 348 2143 0 FreeSans 160 0 0 0 SUB
port 1 nsew
flabel metal4 364 2058 400 2148 0 FreeSans 320 0 0 0 CBOT
port 4 nsew
flabel metal4 244 2488 280 2590 0 FreeSans 320 0 0 0 CTOP
port 6 nsew
flabel metal4 362 928 402 1006 0 FreeSans 320 0 0 0 CTOP
port 8 nsew
flabel pwell 312 2604 338 2636 0 FreeSans 160 0 0 0 x2.SUB
flabel metal4 370 2270 396 2302 0 FreeSans 320 0 0 0 x2.CBOT
flabel metal4 252 2860 278 2892 0 FreeSans 320 0 0 0 x2.CTOP
flabel pwell 306 1080 332 1112 0 FreeSans 160 0 0 0 x1.SUB
flabel metal4 248 1414 274 1446 0 FreeSans 320 0 0 0 x1.CBOT
flabel metal4 366 824 392 856 0 FreeSans 320 0 0 0 x1.CTOP
<< end >>
