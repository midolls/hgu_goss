magic
tech sky130A
magscale 1 2
timestamp 1698674545
<< nwell >>
rect -38 861 314 1182
<< pwell >>
rect 42 621 228 803
rect 42 617 63 621
rect 29 583 63 617
<< scnmos >>
rect 120 647 150 777
<< scpmoshvt >>
rect 120 897 150 1097
<< ndiff >>
rect 68 765 120 777
rect 68 731 76 765
rect 110 731 120 765
rect 68 697 120 731
rect 68 663 76 697
rect 110 663 120 697
rect 68 647 120 663
rect 150 765 202 777
rect 150 731 160 765
rect 194 731 202 765
rect 150 697 202 731
rect 150 663 160 697
rect 194 663 202 697
rect 150 647 202 663
<< pdiff >>
rect 68 1085 120 1097
rect 68 1051 76 1085
rect 110 1051 120 1085
rect 68 1017 120 1051
rect 68 983 76 1017
rect 110 983 120 1017
rect 68 949 120 983
rect 68 915 76 949
rect 110 915 120 949
rect 68 897 120 915
rect 150 1085 202 1097
rect 150 1051 160 1085
rect 194 1051 202 1085
rect 150 1017 202 1051
rect 150 983 160 1017
rect 194 983 202 1017
rect 150 949 202 983
rect 150 915 160 949
rect 194 915 202 949
rect 150 897 202 915
<< ndiffc >>
rect 76 731 110 765
rect 76 663 110 697
rect 160 731 194 765
rect 160 663 194 697
<< pdiffc >>
rect 76 1051 110 1085
rect 76 983 110 1017
rect 76 915 110 949
rect 160 1051 194 1085
rect 160 983 194 1017
rect 160 915 194 949
<< poly >>
rect 120 1097 150 1123
rect 120 865 150 897
rect 64 849 150 865
rect 64 815 80 849
rect 114 815 150 849
rect 64 799 150 815
rect 120 777 150 799
rect 120 621 150 647
<< polycont >>
rect 80 815 114 849
<< locali >>
rect 0 1127 29 1161
rect 63 1127 121 1161
rect 155 1127 213 1161
rect 247 1127 276 1161
rect 68 1085 110 1127
rect 68 1051 76 1085
rect 68 1017 110 1051
rect 68 983 76 1017
rect 68 949 110 983
rect 68 915 76 949
rect 68 899 110 915
rect 144 1085 210 1093
rect 144 1051 160 1085
rect 194 1051 210 1085
rect 144 1017 210 1051
rect 144 983 160 1017
rect 194 983 210 1017
rect 144 949 210 983
rect 144 915 160 949
rect 194 915 210 949
rect 144 897 210 915
rect 64 849 130 863
rect 64 815 80 849
rect 114 815 130 849
rect 64 765 110 781
rect 164 777 210 897
rect 64 731 76 765
rect 64 697 110 731
rect 64 663 76 697
rect 64 617 110 663
rect 144 765 210 777
rect 144 731 160 765
rect 194 731 210 765
rect 144 697 210 731
rect 144 663 160 697
rect 194 663 210 697
rect 144 651 210 663
rect 0 583 29 617
rect 63 583 121 617
rect 155 583 213 617
rect 247 583 276 617
<< viali >>
rect 29 1127 63 1161
rect 121 1127 155 1161
rect 213 1127 247 1161
rect 29 583 63 617
rect 121 583 155 617
rect 213 583 247 617
<< metal1 >>
rect 0 1161 276 1192
rect 0 1127 29 1161
rect 63 1127 121 1161
rect 155 1127 213 1161
rect 247 1127 276 1161
rect 0 1096 276 1127
rect 0 617 276 648
rect 0 583 29 617
rect 63 583 121 617
rect 155 583 213 617
rect 247 583 276 617
rect 0 552 276 583
<< labels >>
flabel locali 164 889 198 923 0 FreeSans 340 0 0 0 x11.Y
flabel locali 164 821 198 855 0 FreeSans 340 0 0 0 x11.Y
flabel locali 72 821 106 855 0 FreeSans 340 0 0 0 x11.A
flabel metal1 29 583 63 617 0 FreeSans 200 0 0 0 x11.VGND
flabel metal1 29 1127 63 1161 0 FreeSans 200 0 0 0 x11.VPWR
rlabel comment 0 600 0 600 4 x11.inv_1
rlabel metal1 0 552 276 648 1 x11.VGND
rlabel metal1 0 1096 276 1192 1 x11.VPWR
flabel pwell 29 583 63 617 0 FreeSans 200 0 0 0 x11.VNB
flabel nwell 29 1127 63 1161 0 FreeSans 200 0 0 0 x11.VPB
<< end >>
