magic
tech sky130A
magscale 1 2
timestamp 1700302578
<< nwell >>
rect 19900 13675 20720 13706
rect 13765 13674 26680 13675
rect 2877 12603 9083 13200
rect 13239 13077 26680 13674
rect 13236 12710 26680 13077
rect 2828 12602 9083 12603
rect 2348 12345 9083 12602
rect 2348 12235 9375 12345
rect 13765 12381 19971 12710
rect 20474 12381 26680 12710
rect 14410 12315 14628 12381
rect 15142 12318 15486 12381
rect 16354 12318 16698 12381
rect 17566 12318 17910 12381
rect 18778 12318 19122 12381
rect 19552 12333 19963 12381
rect 19552 12332 19771 12333
rect 21119 12315 21337 12381
rect 21851 12318 22195 12381
rect 23063 12318 23407 12381
rect 24275 12318 24619 12381
rect 25487 12318 25831 12381
rect 26261 12333 26672 12381
rect 26261 12332 26480 12333
rect 2877 11906 9375 12235
rect 3522 11840 3740 11906
rect 4254 11843 4598 11906
rect 5466 11843 5810 11906
rect 6678 11843 7022 11906
rect 7890 11843 8234 11906
rect 8664 11858 9375 11906
rect 8664 11857 8883 11858
rect 10844 11783 13312 12189
rect 10844 11524 12932 11783
rect 3522 8740 3740 8806
rect 4254 8740 4598 8803
rect 5466 8740 5810 8803
rect 6678 8740 7022 8803
rect 7890 8740 8234 8803
rect 8604 8790 11744 8794
rect 8604 8777 11747 8790
rect 8604 8740 13627 8777
rect 2877 8728 13627 8740
rect 14057 8728 14401 8791
rect 15269 8728 15613 8791
rect 16481 8728 16825 8791
rect 17693 8728 18037 8791
rect 18551 8728 18769 8794
rect 20117 8776 20336 8777
rect 19925 8728 20336 8776
rect 20766 8728 21110 8791
rect 21978 8728 22322 8791
rect 23190 8728 23534 8791
rect 24402 8728 24746 8791
rect 25260 8728 25478 8794
rect 2877 8411 19414 8728
rect 2348 8399 19414 8411
rect 19917 8399 26123 8728
rect 2348 8255 26652 8399
rect 2348 8051 12403 8255
rect 2348 8044 9139 8051
rect 10016 8049 12403 8051
rect 11513 8048 12403 8049
rect 11785 8047 12403 8048
rect 2828 8043 9139 8044
rect 2877 8024 9139 8043
rect 13208 8032 26652 8255
rect 13208 8031 26172 8032
rect 2877 7663 9138 8024
rect 13208 8000 26123 8031
rect 2877 7446 9083 7663
rect 12653 7546 26123 8000
rect 13208 7434 26123 7546
rect 19400 7430 20204 7434
rect 19433 7427 20204 7430
rect 24490 7378 26123 7434
rect 11454 6796 14647 7156
rect 11455 6794 14639 6796
rect 24490 6781 31087 7378
rect 24441 6780 31087 6781
rect 23961 6413 31087 6780
rect 11447 5920 23503 6281
rect 24490 6351 31087 6413
rect 24490 6084 31085 6351
rect 25135 6018 25353 6084
rect 25867 6021 26211 6084
rect 27079 6021 27423 6084
rect 28291 6021 28635 6084
rect 29503 6021 29847 6084
rect 30277 6036 31085 6084
rect 30277 6035 30496 6036
rect 11007 5227 23503 5592
rect 11052 4679 11955 4728
rect 11051 4358 11955 4679
rect 13593 4363 23497 4727
rect 13593 4359 23494 4363
rect 11459 3807 23494 3846
rect 11458 3486 23494 3807
rect 25539 3358 30399 4020
rect 25539 2078 30399 2740
rect 8539 1106 11467 1466
rect 12923 1106 15851 1466
rect 8533 -39 25245 325
rect 8537 -724 25357 -364
rect 8537 -1413 25357 -1052
<< pwell >>
rect 13316 12470 13502 12652
rect 13506 12470 13692 12652
rect 13316 12466 13337 12470
rect 10912 12428 10946 12466
rect 13303 12432 13337 12466
rect 13671 12466 13692 12470
rect 13671 12432 13705 12466
rect 10883 12292 13273 12428
rect 20025 12470 20211 12652
rect 20215 12470 20401 12652
rect 20025 12466 20046 12470
rect 20012 12432 20046 12466
rect 20380 12466 20401 12470
rect 20380 12432 20414 12466
rect 11664 12248 12118 12292
rect 12439 12248 13273 12292
rect 12806 12246 13273 12248
rect 2428 11995 2614 12177
rect 2618 11995 2804 12177
rect 2428 11991 2449 11995
rect 2415 11957 2449 11991
rect 2783 11991 2804 11995
rect 2783 11957 2817 11991
rect 9103 11618 9289 11800
rect 9103 11614 9124 11618
rect 9090 11580 9124 11614
rect 10924 11286 11110 11468
rect 11200 11286 11386 11468
rect 10924 11282 10945 11286
rect 11200 11282 11221 11286
rect 10911 11248 10945 11282
rect 11187 11248 11221 11282
rect 9090 9034 9124 9068
rect 9103 9030 9124 9034
rect 11645 9030 11679 9068
rect 9103 8848 9289 9030
rect 9318 8894 11708 9030
rect 12863 9017 12897 9055
rect 13138 9021 13172 9055
rect 13138 9017 13159 9021
rect 9318 8850 10152 8894
rect 10473 8850 10927 8894
rect 9318 8848 9785 8850
rect 12650 8835 12920 9017
rect 12973 8835 13159 9017
rect 2415 8655 2449 8689
rect 2428 8651 2449 8655
rect 2783 8655 2817 8689
rect 2783 8651 2804 8655
rect 2428 8469 2614 8651
rect 2618 8469 2804 8651
rect 19474 8643 19508 8677
rect 19487 8639 19508 8643
rect 19842 8643 19876 8677
rect 19842 8639 19863 8643
rect 19487 8457 19673 8639
rect 19677 8457 19863 8639
rect 26183 8643 26217 8677
rect 26196 8639 26217 8643
rect 26551 8643 26585 8677
rect 26551 8639 26572 8643
rect 26196 8457 26382 8639
rect 26386 8457 26572 8639
rect 10055 7945 10241 7991
rect 10882 7945 11068 7991
rect 10055 7809 10835 7945
rect 10882 7809 11662 7945
rect 10138 7771 10172 7809
rect 10965 7771 10999 7809
rect 11456 6482 14630 6755
rect 24041 6173 24227 6355
rect 24231 6173 24417 6355
rect 24041 6169 24062 6173
rect 24028 6135 24062 6169
rect 24396 6169 24417 6173
rect 24396 6135 24430 6169
rect 30777 5932 31046 5978
rect 11493 5612 23457 5884
rect 30680 5796 31046 5932
rect 30708 5758 30742 5796
rect 11060 5148 23457 5188
rect 11058 4992 23457 5148
rect 11060 4922 23457 4992
rect 11090 4118 11364 4274
rect 11366 4118 11888 4300
rect 11120 4080 11154 4118
rect 11395 4080 11429 4118
rect 13673 4115 23456 4310
rect 25607 4260 25641 4298
rect 27999 4260 28033 4298
rect 25578 4124 27968 4260
rect 27970 4124 30360 4260
rect 13660 4081 23456 4115
rect 13673 4050 23456 4081
rect 26359 4080 26813 4124
rect 27134 4080 27968 4124
rect 28751 4080 29205 4124
rect 29526 4080 30360 4124
rect 27501 4078 27968 4080
rect 29893 4078 30360 4080
rect 11497 3177 23456 3461
rect 27501 3298 27968 3300
rect 29893 3298 30360 3300
rect 26359 3254 26813 3298
rect 27134 3254 27968 3298
rect 28751 3254 29205 3298
rect 29526 3254 30360 3298
rect 25578 3118 27968 3254
rect 27970 3118 30360 3254
rect 25607 3080 25641 3118
rect 27999 3080 28033 3118
rect 25607 2980 25641 3018
rect 27999 2980 28033 3018
rect 25578 2844 27968 2980
rect 27970 2844 30360 2980
rect 26359 2800 26813 2844
rect 27134 2800 27968 2844
rect 28751 2800 29205 2844
rect 29526 2800 30360 2844
rect 27501 2798 27968 2800
rect 29893 2798 30360 2800
rect 27501 2018 27968 2020
rect 29893 2018 30360 2020
rect 26359 1974 26813 2018
rect 27134 1974 27968 2018
rect 28751 1974 29205 2018
rect 29526 1974 30360 2018
rect 25578 1838 27968 1974
rect 27970 1838 30360 1974
rect 25607 1800 25641 1838
rect 27999 1800 28033 1838
rect 8578 866 8852 1022
rect 8854 866 9376 1048
rect 9406 866 11356 1048
rect 12962 866 13236 1022
rect 13238 866 13760 1048
rect 13790 866 15740 1048
rect 8608 828 8642 866
rect 8883 828 8917 866
rect 9435 828 9469 866
rect 12992 828 13026 866
rect 13267 828 13301 866
rect 13819 828 13853 866
rect 8576 -140 8762 -94
rect 10650 -140 10836 -94
rect 8576 -276 9356 -140
rect 10056 -276 10836 -140
rect 10968 -140 11154 -94
rect 13042 -140 13228 -94
rect 10968 -276 11748 -140
rect 12448 -276 13228 -140
rect 13360 -140 13546 -94
rect 15432 -140 15618 -94
rect 13360 -276 14140 -140
rect 14838 -276 15618 -140
rect 15752 -140 15938 -94
rect 17826 -140 18012 -94
rect 15752 -276 16532 -140
rect 17232 -276 18012 -140
rect 18144 -140 18330 -94
rect 20218 -140 20404 -94
rect 18144 -276 18924 -140
rect 19624 -276 20404 -140
rect 20536 -140 20722 -94
rect 22608 -140 22794 -94
rect 20536 -276 21316 -140
rect 22014 -276 22794 -140
rect 22928 -140 23114 -94
rect 25002 -140 25188 -94
rect 22928 -276 23708 -140
rect 24408 -276 25188 -140
rect 8659 -314 8693 -276
rect 10719 -314 10753 -276
rect 11051 -314 11085 -276
rect 13111 -314 13145 -276
rect 13443 -314 13477 -276
rect 15501 -314 15535 -276
rect 15835 -314 15869 -276
rect 17895 -314 17929 -276
rect 18227 -314 18261 -276
rect 20287 -314 20321 -276
rect 20619 -314 20653 -276
rect 22677 -314 22711 -276
rect 23011 -314 23045 -276
rect 25071 -314 25105 -276
rect 10499 -784 10966 -782
rect 12891 -784 13358 -782
rect 15283 -784 15750 -782
rect 17675 -784 18142 -782
rect 20067 -784 20534 -782
rect 22459 -784 22926 -782
rect 24851 -784 25318 -782
rect 9355 -828 9810 -784
rect 10132 -828 10966 -784
rect 11747 -828 12202 -784
rect 12524 -828 13358 -784
rect 14139 -828 14594 -784
rect 14916 -828 15750 -784
rect 16531 -828 16986 -784
rect 17308 -828 18142 -784
rect 18923 -828 19378 -784
rect 19700 -828 20534 -784
rect 21315 -828 21770 -784
rect 22092 -828 22926 -784
rect 23707 -828 24162 -784
rect 24484 -828 25318 -784
rect 8576 -964 10966 -828
rect 10968 -964 13358 -828
rect 13360 -964 15750 -828
rect 15752 -964 18142 -828
rect 18144 -964 20534 -828
rect 20536 -964 22926 -828
rect 22928 -964 25318 -828
rect 8604 -1002 8638 -964
rect 10996 -1002 11030 -964
rect 13388 -1002 13422 -964
rect 15780 -1002 15814 -964
rect 18172 -1002 18206 -964
rect 20564 -1002 20598 -964
rect 22956 -1002 22990 -964
rect 8576 -1473 9043 -1471
rect 10968 -1473 11435 -1471
rect 13360 -1473 13827 -1471
rect 15752 -1473 16219 -1471
rect 18144 -1473 18611 -1471
rect 20536 -1473 21003 -1471
rect 22928 -1473 23395 -1471
rect 8576 -1517 9410 -1473
rect 9732 -1517 10187 -1473
rect 10968 -1517 11802 -1473
rect 12124 -1517 12579 -1473
rect 13360 -1517 14194 -1473
rect 14516 -1517 14971 -1473
rect 15752 -1517 16586 -1473
rect 16908 -1517 17363 -1473
rect 18144 -1517 18978 -1473
rect 19300 -1517 19755 -1473
rect 20536 -1517 21370 -1473
rect 21692 -1517 22147 -1473
rect 22928 -1517 23762 -1473
rect 24084 -1517 24539 -1473
rect 8576 -1653 10966 -1517
rect 10968 -1653 13358 -1517
rect 13360 -1653 15750 -1517
rect 15752 -1653 18142 -1517
rect 18144 -1653 20534 -1517
rect 20536 -1653 22926 -1517
rect 22928 -1653 25318 -1517
rect 10904 -1691 10938 -1653
rect 13296 -1691 13330 -1653
rect 15688 -1691 15722 -1653
rect 18080 -1691 18114 -1653
rect 20472 -1691 20506 -1653
rect 22864 -1691 22898 -1653
rect 25256 -1691 25290 -1653
<< nmos >>
rect 14857 12166 14887 12250
rect 15589 12166 15619 12250
rect 15711 12166 15741 12250
rect 16801 12166 16831 12250
rect 16923 12166 16953 12250
rect 18139 12166 18169 12250
rect 18261 12166 18291 12250
rect 18995 12166 19025 12250
rect 19647 12167 19677 12251
rect 19739 12167 19769 12251
rect 19835 12167 19865 12251
rect 21566 12166 21596 12250
rect 22298 12166 22328 12250
rect 22420 12166 22450 12250
rect 23510 12166 23540 12250
rect 23632 12166 23662 12250
rect 24848 12166 24878 12250
rect 24970 12166 25000 12250
rect 25704 12166 25734 12250
rect 26356 12167 26386 12251
rect 26448 12167 26478 12251
rect 26544 12167 26574 12251
rect 13837 11982 13867 12066
rect 13909 11982 13939 12066
rect 19647 12029 19677 12113
rect 20546 11982 20576 12066
rect 20618 11982 20648 12066
rect 26356 12029 26386 12113
rect 13837 11844 13867 11928
rect 13909 11844 13939 11928
rect 20546 11844 20576 11928
rect 20618 11844 20648 11928
rect 3969 11691 3999 11775
rect 4701 11691 4731 11775
rect 4823 11691 4853 11775
rect 5913 11691 5943 11775
rect 6035 11691 6065 11775
rect 7251 11691 7281 11775
rect 7373 11691 7403 11775
rect 8107 11691 8137 11775
rect 8759 11692 8789 11776
rect 8851 11692 8881 11776
rect 8947 11692 8977 11776
rect 2949 11507 2979 11591
rect 3021 11507 3051 11591
rect 8759 11554 8789 11638
rect 13837 11706 13867 11790
rect 13909 11706 13939 11790
rect 20546 11706 20576 11790
rect 20618 11706 20648 11790
rect 13837 11568 13867 11652
rect 13909 11568 13939 11652
rect 20546 11568 20576 11652
rect 20618 11568 20648 11652
rect 2949 11369 2979 11453
rect 3021 11369 3051 11453
rect 2949 11231 2979 11315
rect 3021 11231 3051 11315
rect 13837 11430 13867 11514
rect 13909 11430 13939 11514
rect 20546 11430 20576 11514
rect 20618 11430 20648 11514
rect 13837 11292 13867 11376
rect 13909 11292 13939 11376
rect 20546 11292 20576 11376
rect 20618 11292 20648 11376
rect 2949 11093 2979 11177
rect 3021 11093 3051 11177
rect 13837 11154 13867 11238
rect 13909 11154 13939 11238
rect 20546 11154 20576 11238
rect 20618 11154 20648 11238
rect 2949 10955 2979 11039
rect 3021 10955 3051 11039
rect 13837 11016 13867 11100
rect 13909 11016 13939 11100
rect 20546 11016 20576 11100
rect 20618 11016 20648 11100
rect 2949 10817 2979 10901
rect 3021 10817 3051 10901
rect 2949 10679 2979 10763
rect 3021 10679 3051 10763
rect 2949 10541 2979 10625
rect 3021 10541 3051 10625
rect 2949 10021 2979 10105
rect 3021 10021 3051 10105
rect 19240 10009 19270 10093
rect 19312 10009 19342 10093
rect 25949 10009 25979 10093
rect 26021 10009 26051 10093
rect 2949 9883 2979 9967
rect 3021 9883 3051 9967
rect 19240 9871 19270 9955
rect 19312 9871 19342 9955
rect 2949 9745 2979 9829
rect 3021 9745 3051 9829
rect 25949 9871 25979 9955
rect 26021 9871 26051 9955
rect 19240 9733 19270 9817
rect 19312 9733 19342 9817
rect 25949 9733 25979 9817
rect 26021 9733 26051 9817
rect 2949 9607 2979 9691
rect 3021 9607 3051 9691
rect 19240 9595 19270 9679
rect 19312 9595 19342 9679
rect 25949 9595 25979 9679
rect 26021 9595 26051 9679
rect 2949 9469 2979 9553
rect 3021 9469 3051 9553
rect 19240 9457 19270 9541
rect 19312 9457 19342 9541
rect 25949 9457 25979 9541
rect 26021 9457 26051 9541
rect 2949 9331 2979 9415
rect 3021 9331 3051 9415
rect 19240 9319 19270 9403
rect 19312 9319 19342 9403
rect 25949 9319 25979 9403
rect 26021 9319 26051 9403
rect 2949 9193 2979 9277
rect 3021 9193 3051 9277
rect 19240 9181 19270 9265
rect 19312 9181 19342 9265
rect 25949 9181 25979 9265
rect 26021 9181 26051 9265
rect 2949 9055 2979 9139
rect 3021 9055 3051 9139
rect 8759 9008 8789 9092
rect 3969 8871 3999 8955
rect 4701 8871 4731 8955
rect 4823 8871 4853 8955
rect 5913 8871 5943 8955
rect 6035 8871 6065 8955
rect 7251 8871 7281 8955
rect 7373 8871 7403 8955
rect 8107 8871 8137 8955
rect 8759 8870 8789 8954
rect 8851 8870 8881 8954
rect 8947 8870 8977 8954
rect 13502 8996 13532 9080
rect 19240 9043 19270 9127
rect 19312 9043 19342 9127
rect 11883 8872 11913 8956
rect 11979 8872 12009 8956
rect 12075 8872 12105 8956
rect 12279 8860 12309 8944
rect 12480 8859 12510 8943
rect 20211 8996 20241 9080
rect 25949 9043 25979 9127
rect 26021 9043 26051 9127
rect 13314 8858 13344 8942
rect 13410 8858 13440 8942
rect 13502 8858 13532 8942
rect 14154 8859 14184 8943
rect 14888 8859 14918 8943
rect 15010 8859 15040 8943
rect 16226 8859 16256 8943
rect 16348 8859 16378 8943
rect 17438 8859 17468 8943
rect 17560 8859 17590 8943
rect 18292 8859 18322 8943
rect 20023 8858 20053 8942
rect 20119 8858 20149 8942
rect 20211 8858 20241 8942
rect 20863 8859 20893 8943
rect 21597 8859 21627 8943
rect 21719 8859 21749 8943
rect 22935 8859 22965 8943
rect 23057 8859 23087 8943
rect 24147 8859 24177 8943
rect 24269 8859 24299 8943
rect 25001 8859 25031 8943
rect 12748 8068 12778 8152
rect 11883 7868 11913 7952
rect 11979 7868 12009 7952
rect 12075 7868 12105 7952
rect 12279 7880 12309 7964
rect 25582 5869 25612 5953
rect 26314 5869 26344 5953
rect 26436 5869 26466 5953
rect 27526 5869 27556 5953
rect 27648 5869 27678 5953
rect 28864 5869 28894 5953
rect 28986 5869 29016 5953
rect 29720 5869 29750 5953
rect 30372 5870 30402 5954
rect 30464 5870 30494 5954
rect 30560 5870 30590 5954
rect 24562 5685 24592 5769
rect 24634 5685 24664 5769
rect 30372 5732 30402 5816
rect 24562 5547 24592 5631
rect 24634 5547 24664 5631
rect 24562 5409 24592 5493
rect 24634 5409 24664 5493
rect 24562 5271 24592 5355
rect 24634 5271 24664 5355
rect 24562 5133 24592 5217
rect 24634 5133 24664 5217
rect 24562 4995 24592 5079
rect 24634 4995 24664 5079
rect 24562 4857 24592 4941
rect 24634 4857 24664 4941
rect 24562 4719 24592 4803
rect 24634 4719 24664 4803
<< scnmos >>
rect 13394 12496 13424 12626
rect 13584 12496 13614 12626
rect 20103 12496 20133 12626
rect 20293 12496 20323 12626
rect 10961 12318 10991 12402
rect 11045 12318 11075 12402
rect 11233 12318 11263 12402
rect 11328 12330 11358 12402
rect 11434 12330 11464 12402
rect 11530 12318 11560 12402
rect 11640 12318 11670 12402
rect 2506 12021 2536 12151
rect 2696 12021 2726 12151
rect 11740 12274 11770 12402
rect 11824 12274 11854 12402
rect 12012 12274 12042 12402
rect 12107 12330 12137 12402
rect 12216 12330 12246 12402
rect 12311 12318 12341 12402
rect 12397 12318 12427 12402
rect 12515 12274 12545 12402
rect 12599 12274 12629 12402
rect 12787 12318 12817 12402
rect 12882 12272 12912 12402
rect 13070 12318 13100 12402
rect 13165 12272 13195 12402
rect 9181 11644 9211 11774
rect 11002 11312 11032 11442
rect 11278 11312 11308 11442
rect 9181 8874 9211 9004
rect 9396 8874 9426 9004
rect 9491 8920 9521 9004
rect 9679 8874 9709 9004
rect 9774 8920 9804 9004
rect 9962 8876 9992 9004
rect 10046 8876 10076 9004
rect 10164 8920 10194 9004
rect 10250 8920 10280 9004
rect 10345 8932 10375 9004
rect 10454 8932 10484 9004
rect 2506 8495 2536 8625
rect 2696 8495 2726 8625
rect 10549 8876 10579 9004
rect 10737 8876 10767 9004
rect 10821 8876 10851 9004
rect 10921 8920 10951 9004
rect 11031 8920 11061 9004
rect 11127 8932 11157 9004
rect 11233 8932 11263 9004
rect 11328 8920 11358 9004
rect 11516 8920 11546 9004
rect 11600 8920 11630 9004
rect 12728 8861 12758 8991
rect 12812 8861 12842 8991
rect 13051 8861 13081 8991
rect 19565 8483 19595 8613
rect 19755 8483 19785 8613
rect 26274 8483 26304 8613
rect 26464 8483 26494 8613
rect 10133 7835 10163 7965
rect 10242 7835 10272 7919
rect 10338 7835 10368 7919
rect 10463 7835 10493 7919
rect 10559 7835 10589 7919
rect 10727 7835 10757 7919
rect 10960 7835 10990 7965
rect 11069 7835 11099 7919
rect 11165 7835 11195 7919
rect 11290 7835 11320 7919
rect 11386 7835 11416 7919
rect 11554 7835 11584 7919
rect 11577 6580 11607 6684
rect 11665 6580 11695 6684
rect 11853 6580 11883 6710
rect 11937 6580 11967 6710
rect 12021 6580 12051 6710
rect 12105 6580 12135 6710
rect 12189 6580 12219 6710
rect 12852 6580 12882 6710
rect 12936 6580 12966 6710
rect 13036 6580 13066 6710
rect 13120 6580 13150 6710
rect 13221 6580 13251 6664
rect 13316 6580 13346 6652
rect 13426 6580 13456 6652
rect 13533 6580 13563 6664
rect 13721 6580 13751 6664
rect 13806 6580 13836 6664
rect 13996 6580 14026 6664
rect 14104 6580 14134 6664
rect 14200 6580 14230 6652
rect 14310 6580 14340 6652
rect 14405 6580 14435 6664
rect 14489 6580 14519 6664
rect 24119 6199 24149 6329
rect 24309 6199 24339 6329
rect 11576 5707 11606 5791
rect 11660 5707 11690 5791
rect 11848 5707 11878 5791
rect 11943 5707 11973 5779
rect 12049 5707 12079 5779
rect 12145 5707 12175 5791
rect 12255 5707 12285 5791
rect 12355 5707 12385 5835
rect 12439 5707 12469 5835
rect 12627 5707 12657 5835
rect 12722 5707 12752 5779
rect 12831 5707 12861 5779
rect 12926 5707 12956 5791
rect 13012 5707 13042 5791
rect 13130 5707 13160 5835
rect 13214 5707 13244 5835
rect 13402 5707 13432 5791
rect 13497 5707 13527 5837
rect 13685 5707 13715 5791
rect 13780 5707 13810 5837
rect 13968 5707 13998 5791
rect 14052 5707 14082 5791
rect 14240 5707 14270 5791
rect 14335 5707 14365 5779
rect 14441 5707 14471 5779
rect 14537 5707 14567 5791
rect 14647 5707 14677 5791
rect 14747 5707 14777 5835
rect 14831 5707 14861 5835
rect 15019 5707 15049 5835
rect 15114 5707 15144 5779
rect 15223 5707 15253 5779
rect 15318 5707 15348 5791
rect 15404 5707 15434 5791
rect 15522 5707 15552 5835
rect 15606 5707 15636 5835
rect 15794 5707 15824 5791
rect 15889 5707 15919 5837
rect 16077 5707 16107 5791
rect 16172 5707 16202 5837
rect 16360 5707 16390 5791
rect 16444 5707 16474 5791
rect 16632 5707 16662 5791
rect 16727 5707 16757 5779
rect 16833 5707 16863 5779
rect 16929 5707 16959 5791
rect 17039 5707 17069 5791
rect 17139 5707 17169 5835
rect 17223 5707 17253 5835
rect 17411 5707 17441 5835
rect 17506 5707 17536 5779
rect 17615 5707 17645 5779
rect 17710 5707 17740 5791
rect 17796 5707 17826 5791
rect 17914 5707 17944 5835
rect 17998 5707 18028 5835
rect 18186 5707 18216 5791
rect 18281 5707 18311 5837
rect 18469 5707 18499 5791
rect 18564 5707 18594 5837
rect 18752 5707 18782 5791
rect 18836 5707 18866 5791
rect 19024 5707 19054 5791
rect 19119 5707 19149 5779
rect 19225 5707 19255 5779
rect 19321 5707 19351 5791
rect 19431 5707 19461 5791
rect 19531 5707 19561 5835
rect 19615 5707 19645 5835
rect 19803 5707 19833 5835
rect 19898 5707 19928 5779
rect 20007 5707 20037 5779
rect 20102 5707 20132 5791
rect 20188 5707 20218 5791
rect 20306 5707 20336 5835
rect 20390 5707 20420 5835
rect 20578 5707 20608 5791
rect 20673 5707 20703 5837
rect 20861 5707 20891 5791
rect 20956 5707 20986 5837
rect 21144 5707 21174 5791
rect 21228 5707 21258 5791
rect 21416 5707 21446 5791
rect 21511 5707 21541 5779
rect 21617 5707 21647 5779
rect 21713 5707 21743 5791
rect 21823 5707 21853 5791
rect 21923 5707 21953 5835
rect 22007 5707 22037 5835
rect 22195 5707 22225 5835
rect 22290 5707 22320 5779
rect 22399 5707 22429 5779
rect 22494 5707 22524 5791
rect 22580 5707 22610 5791
rect 22698 5707 22728 5835
rect 22782 5707 22812 5835
rect 22970 5707 23000 5791
rect 23065 5707 23095 5837
rect 23253 5707 23283 5791
rect 23348 5707 23378 5837
rect 30758 5822 30788 5906
rect 30853 5822 30883 5952
rect 30937 5822 30967 5952
rect 11136 5018 11166 5122
rect 11224 5018 11254 5122
rect 11412 5018 11442 5148
rect 11496 5018 11526 5148
rect 11580 5018 11610 5148
rect 11664 5018 11694 5148
rect 11748 5018 11778 5148
rect 11944 5018 11974 5148
rect 12028 5018 12058 5148
rect 12112 5018 12142 5148
rect 12196 5018 12226 5148
rect 12280 5018 12310 5148
rect 12364 5018 12394 5148
rect 12448 5018 12478 5148
rect 12532 5018 12562 5148
rect 12616 5018 12646 5148
rect 12700 5018 12730 5148
rect 12784 5018 12814 5148
rect 12868 5018 12898 5148
rect 12952 5018 12982 5148
rect 13036 5018 13066 5148
rect 13120 5018 13150 5148
rect 13204 5018 13234 5148
rect 13288 5018 13318 5148
rect 13372 5018 13402 5148
rect 13456 5018 13486 5148
rect 13540 5018 13570 5148
rect 13624 5018 13654 5148
rect 13708 5018 13738 5148
rect 13968 5018 13998 5148
rect 14063 5018 14093 5102
rect 14251 5018 14281 5148
rect 14346 5018 14376 5102
rect 14534 5018 14564 5146
rect 14618 5018 14648 5146
rect 14736 5018 14766 5102
rect 14822 5018 14852 5102
rect 14917 5018 14947 5090
rect 15026 5018 15056 5090
rect 15121 5018 15151 5146
rect 15309 5018 15339 5146
rect 15393 5018 15423 5146
rect 15493 5018 15523 5102
rect 15603 5018 15633 5102
rect 15699 5018 15729 5090
rect 15805 5018 15835 5090
rect 15900 5018 15930 5102
rect 16088 5018 16118 5102
rect 16172 5018 16202 5102
rect 16360 5018 16390 5148
rect 16455 5018 16485 5102
rect 16643 5018 16673 5148
rect 16738 5018 16768 5102
rect 16926 5018 16956 5146
rect 17010 5018 17040 5146
rect 17128 5018 17158 5102
rect 17214 5018 17244 5102
rect 17309 5018 17339 5090
rect 17418 5018 17448 5090
rect 17513 5018 17543 5146
rect 17701 5018 17731 5146
rect 17785 5018 17815 5146
rect 17885 5018 17915 5102
rect 17995 5018 18025 5102
rect 18091 5018 18121 5090
rect 18197 5018 18227 5090
rect 18292 5018 18322 5102
rect 18480 5018 18510 5102
rect 18564 5018 18594 5102
rect 18752 5018 18782 5148
rect 18847 5018 18877 5102
rect 19035 5018 19065 5148
rect 19130 5018 19160 5102
rect 19318 5018 19348 5146
rect 19402 5018 19432 5146
rect 19520 5018 19550 5102
rect 19606 5018 19636 5102
rect 19701 5018 19731 5090
rect 19810 5018 19840 5090
rect 19905 5018 19935 5146
rect 20093 5018 20123 5146
rect 20177 5018 20207 5146
rect 20277 5018 20307 5102
rect 20387 5018 20417 5102
rect 20483 5018 20513 5090
rect 20589 5018 20619 5090
rect 20684 5018 20714 5102
rect 20872 5018 20902 5102
rect 20956 5018 20986 5102
rect 21144 5018 21174 5148
rect 21239 5018 21269 5102
rect 21427 5018 21457 5148
rect 21522 5018 21552 5102
rect 21710 5018 21740 5146
rect 21794 5018 21824 5146
rect 21912 5018 21942 5102
rect 21998 5018 22028 5102
rect 22093 5018 22123 5090
rect 22202 5018 22232 5090
rect 22297 5018 22327 5146
rect 22485 5018 22515 5146
rect 22569 5018 22599 5146
rect 22669 5018 22699 5102
rect 22779 5018 22809 5102
rect 22875 5018 22905 5090
rect 22981 5018 23011 5090
rect 23076 5018 23106 5102
rect 23264 5018 23294 5102
rect 23348 5018 23378 5102
rect 11168 4144 11198 4248
rect 11256 4144 11286 4248
rect 11444 4144 11474 4274
rect 11528 4144 11558 4274
rect 11612 4144 11642 4274
rect 11696 4144 11726 4274
rect 11780 4144 11810 4274
rect 13751 4145 13781 4275
rect 13967 4145 13997 4229
rect 14051 4145 14081 4229
rect 14239 4145 14269 4229
rect 14334 4145 14364 4217
rect 14440 4145 14470 4217
rect 14536 4145 14566 4229
rect 14646 4145 14676 4229
rect 14746 4145 14776 4273
rect 14830 4145 14860 4273
rect 15018 4145 15048 4273
rect 15113 4145 15143 4217
rect 15222 4145 15252 4217
rect 15317 4145 15347 4229
rect 15403 4145 15433 4229
rect 15521 4145 15551 4273
rect 15605 4145 15635 4273
rect 15793 4145 15823 4229
rect 15888 4145 15918 4275
rect 16076 4145 16106 4229
rect 16171 4145 16201 4275
rect 16359 4145 16389 4229
rect 16443 4145 16473 4229
rect 16631 4145 16661 4229
rect 16726 4145 16756 4217
rect 16832 4145 16862 4217
rect 16928 4145 16958 4229
rect 17038 4145 17068 4229
rect 17138 4145 17168 4273
rect 17222 4145 17252 4273
rect 17410 4145 17440 4273
rect 17505 4145 17535 4217
rect 17614 4145 17644 4217
rect 17709 4145 17739 4229
rect 17795 4145 17825 4229
rect 17913 4145 17943 4273
rect 17997 4145 18027 4273
rect 18185 4145 18215 4229
rect 18280 4145 18310 4275
rect 18468 4145 18498 4229
rect 18563 4145 18593 4275
rect 18751 4145 18781 4229
rect 18835 4145 18865 4229
rect 19023 4145 19053 4229
rect 19118 4145 19148 4217
rect 19224 4145 19254 4217
rect 19320 4145 19350 4229
rect 19430 4145 19460 4229
rect 19530 4145 19560 4273
rect 19614 4145 19644 4273
rect 19802 4145 19832 4273
rect 19897 4145 19927 4217
rect 20006 4145 20036 4217
rect 20101 4145 20131 4229
rect 20187 4145 20217 4229
rect 20305 4145 20335 4273
rect 20389 4145 20419 4273
rect 20577 4145 20607 4229
rect 20672 4145 20702 4275
rect 20860 4145 20890 4229
rect 20955 4145 20985 4275
rect 21143 4145 21173 4229
rect 21227 4145 21257 4229
rect 21415 4145 21445 4229
rect 21510 4145 21540 4217
rect 21616 4145 21646 4217
rect 21712 4145 21742 4229
rect 21822 4145 21852 4229
rect 21922 4145 21952 4273
rect 22006 4145 22036 4273
rect 22194 4145 22224 4273
rect 22289 4145 22319 4217
rect 22398 4145 22428 4217
rect 22493 4145 22523 4229
rect 22579 4145 22609 4229
rect 22697 4145 22727 4273
rect 22781 4145 22811 4273
rect 22969 4145 22999 4229
rect 23064 4145 23094 4275
rect 23252 4145 23282 4229
rect 23347 4145 23377 4275
rect 25656 4150 25686 4234
rect 25740 4150 25770 4234
rect 25928 4150 25958 4234
rect 26023 4162 26053 4234
rect 26129 4162 26159 4234
rect 26225 4150 26255 4234
rect 26335 4150 26365 4234
rect 26435 4106 26465 4234
rect 26519 4106 26549 4234
rect 26707 4106 26737 4234
rect 26802 4162 26832 4234
rect 26911 4162 26941 4234
rect 27006 4150 27036 4234
rect 27092 4150 27122 4234
rect 27210 4106 27240 4234
rect 27294 4106 27324 4234
rect 27482 4150 27512 4234
rect 27577 4104 27607 4234
rect 27765 4150 27795 4234
rect 27860 4104 27890 4234
rect 28048 4150 28078 4234
rect 28132 4150 28162 4234
rect 28320 4150 28350 4234
rect 28415 4162 28445 4234
rect 28521 4162 28551 4234
rect 28617 4150 28647 4234
rect 28727 4150 28757 4234
rect 28827 4106 28857 4234
rect 28911 4106 28941 4234
rect 29099 4106 29129 4234
rect 29194 4162 29224 4234
rect 29303 4162 29333 4234
rect 29398 4150 29428 4234
rect 29484 4150 29514 4234
rect 29602 4106 29632 4234
rect 29686 4106 29716 4234
rect 29874 4150 29904 4234
rect 29969 4104 29999 4234
rect 30157 4150 30187 4234
rect 30252 4104 30282 4234
rect 11575 3272 11605 3402
rect 11670 3272 11700 3356
rect 11858 3272 11888 3402
rect 11953 3272 11983 3356
rect 12141 3272 12171 3400
rect 12225 3272 12255 3400
rect 12343 3272 12373 3356
rect 12429 3272 12459 3356
rect 12524 3272 12554 3344
rect 12633 3272 12663 3344
rect 12728 3272 12758 3400
rect 12916 3272 12946 3400
rect 13000 3272 13030 3400
rect 13100 3272 13130 3356
rect 13210 3272 13240 3356
rect 13306 3272 13336 3344
rect 13412 3272 13442 3344
rect 13507 3272 13537 3356
rect 13695 3272 13725 3356
rect 13779 3272 13809 3356
rect 13967 3272 13997 3402
rect 14062 3272 14092 3356
rect 14250 3272 14280 3402
rect 14345 3272 14375 3356
rect 14533 3272 14563 3400
rect 14617 3272 14647 3400
rect 14735 3272 14765 3356
rect 14821 3272 14851 3356
rect 14916 3272 14946 3344
rect 15025 3272 15055 3344
rect 15120 3272 15150 3400
rect 15308 3272 15338 3400
rect 15392 3272 15422 3400
rect 15492 3272 15522 3356
rect 15602 3272 15632 3356
rect 15698 3272 15728 3344
rect 15804 3272 15834 3344
rect 15899 3272 15929 3356
rect 16087 3272 16117 3356
rect 16171 3272 16201 3356
rect 16359 3272 16389 3402
rect 16454 3272 16484 3356
rect 16642 3272 16672 3402
rect 16737 3272 16767 3356
rect 16925 3272 16955 3400
rect 17009 3272 17039 3400
rect 17127 3272 17157 3356
rect 17213 3272 17243 3356
rect 17308 3272 17338 3344
rect 17417 3272 17447 3344
rect 17512 3272 17542 3400
rect 17700 3272 17730 3400
rect 17784 3272 17814 3400
rect 17884 3272 17914 3356
rect 17994 3272 18024 3356
rect 18090 3272 18120 3344
rect 18196 3272 18226 3344
rect 18291 3272 18321 3356
rect 18479 3272 18509 3356
rect 18563 3272 18593 3356
rect 18751 3272 18781 3402
rect 18846 3272 18876 3356
rect 19034 3272 19064 3402
rect 19129 3272 19159 3356
rect 19317 3272 19347 3400
rect 19401 3272 19431 3400
rect 19519 3272 19549 3356
rect 19605 3272 19635 3356
rect 19700 3272 19730 3344
rect 19809 3272 19839 3344
rect 19904 3272 19934 3400
rect 20092 3272 20122 3400
rect 20176 3272 20206 3400
rect 20276 3272 20306 3356
rect 20386 3272 20416 3356
rect 20482 3272 20512 3344
rect 20588 3272 20618 3344
rect 20683 3272 20713 3356
rect 20871 3272 20901 3356
rect 20955 3272 20985 3356
rect 21143 3272 21173 3402
rect 21238 3272 21268 3356
rect 21426 3272 21456 3402
rect 21521 3272 21551 3356
rect 21709 3272 21739 3400
rect 21793 3272 21823 3400
rect 21911 3272 21941 3356
rect 21997 3272 22027 3356
rect 22092 3272 22122 3344
rect 22201 3272 22231 3344
rect 22296 3272 22326 3400
rect 22484 3272 22514 3400
rect 22568 3272 22598 3400
rect 22668 3272 22698 3356
rect 22778 3272 22808 3356
rect 22874 3272 22904 3344
rect 22980 3272 23010 3344
rect 23075 3272 23105 3356
rect 23263 3272 23293 3356
rect 23347 3272 23377 3356
rect 25656 3144 25686 3228
rect 25740 3144 25770 3228
rect 25928 3144 25958 3228
rect 26023 3144 26053 3216
rect 26129 3144 26159 3216
rect 26225 3144 26255 3228
rect 26335 3144 26365 3228
rect 26435 3144 26465 3272
rect 26519 3144 26549 3272
rect 26707 3144 26737 3272
rect 26802 3144 26832 3216
rect 26911 3144 26941 3216
rect 27006 3144 27036 3228
rect 27092 3144 27122 3228
rect 27210 3144 27240 3272
rect 27294 3144 27324 3272
rect 27482 3144 27512 3228
rect 27577 3144 27607 3274
rect 27765 3144 27795 3228
rect 27860 3144 27890 3274
rect 28048 3144 28078 3228
rect 28132 3144 28162 3228
rect 28320 3144 28350 3228
rect 28415 3144 28445 3216
rect 28521 3144 28551 3216
rect 28617 3144 28647 3228
rect 28727 3144 28757 3228
rect 28827 3144 28857 3272
rect 28911 3144 28941 3272
rect 29099 3144 29129 3272
rect 29194 3144 29224 3216
rect 29303 3144 29333 3216
rect 29398 3144 29428 3228
rect 29484 3144 29514 3228
rect 29602 3144 29632 3272
rect 29686 3144 29716 3272
rect 29874 3144 29904 3228
rect 29969 3144 29999 3274
rect 30157 3144 30187 3228
rect 30252 3144 30282 3274
rect 25656 2870 25686 2954
rect 25740 2870 25770 2954
rect 25928 2870 25958 2954
rect 26023 2882 26053 2954
rect 26129 2882 26159 2954
rect 26225 2870 26255 2954
rect 26335 2870 26365 2954
rect 26435 2826 26465 2954
rect 26519 2826 26549 2954
rect 26707 2826 26737 2954
rect 26802 2882 26832 2954
rect 26911 2882 26941 2954
rect 27006 2870 27036 2954
rect 27092 2870 27122 2954
rect 27210 2826 27240 2954
rect 27294 2826 27324 2954
rect 27482 2870 27512 2954
rect 27577 2824 27607 2954
rect 27765 2870 27795 2954
rect 27860 2824 27890 2954
rect 28048 2870 28078 2954
rect 28132 2870 28162 2954
rect 28320 2870 28350 2954
rect 28415 2882 28445 2954
rect 28521 2882 28551 2954
rect 28617 2870 28647 2954
rect 28727 2870 28757 2954
rect 28827 2826 28857 2954
rect 28911 2826 28941 2954
rect 29099 2826 29129 2954
rect 29194 2882 29224 2954
rect 29303 2882 29333 2954
rect 29398 2870 29428 2954
rect 29484 2870 29514 2954
rect 29602 2826 29632 2954
rect 29686 2826 29716 2954
rect 29874 2870 29904 2954
rect 29969 2824 29999 2954
rect 30157 2870 30187 2954
rect 30252 2824 30282 2954
rect 25656 1864 25686 1948
rect 25740 1864 25770 1948
rect 25928 1864 25958 1948
rect 26023 1864 26053 1936
rect 26129 1864 26159 1936
rect 26225 1864 26255 1948
rect 26335 1864 26365 1948
rect 26435 1864 26465 1992
rect 26519 1864 26549 1992
rect 26707 1864 26737 1992
rect 26802 1864 26832 1936
rect 26911 1864 26941 1936
rect 27006 1864 27036 1948
rect 27092 1864 27122 1948
rect 27210 1864 27240 1992
rect 27294 1864 27324 1992
rect 27482 1864 27512 1948
rect 27577 1864 27607 1994
rect 27765 1864 27795 1948
rect 27860 1864 27890 1994
rect 28048 1864 28078 1948
rect 28132 1864 28162 1948
rect 28320 1864 28350 1948
rect 28415 1864 28445 1936
rect 28521 1864 28551 1936
rect 28617 1864 28647 1948
rect 28727 1864 28757 1948
rect 28827 1864 28857 1992
rect 28911 1864 28941 1992
rect 29099 1864 29129 1992
rect 29194 1864 29224 1936
rect 29303 1864 29333 1936
rect 29398 1864 29428 1948
rect 29484 1864 29514 1948
rect 29602 1864 29632 1992
rect 29686 1864 29716 1992
rect 29874 1864 29904 1948
rect 29969 1864 29999 1994
rect 30157 1864 30187 1948
rect 30252 1864 30282 1994
rect 8656 892 8686 996
rect 8744 892 8774 996
rect 8932 892 8962 1022
rect 9016 892 9046 1022
rect 9100 892 9130 1022
rect 9184 892 9214 1022
rect 9268 892 9298 1022
rect 9484 892 9514 1022
rect 9568 892 9598 1022
rect 9652 892 9682 1022
rect 9736 892 9766 1022
rect 9820 892 9850 1022
rect 9904 892 9934 1022
rect 9988 892 10018 1022
rect 10072 892 10102 1022
rect 10156 892 10186 1022
rect 10240 892 10270 1022
rect 10324 892 10354 1022
rect 10408 892 10438 1022
rect 10492 892 10522 1022
rect 10576 892 10606 1022
rect 10660 892 10690 1022
rect 10744 892 10774 1022
rect 10828 892 10858 1022
rect 10912 892 10942 1022
rect 10996 892 11026 1022
rect 11080 892 11110 1022
rect 11164 892 11194 1022
rect 11248 892 11278 1022
rect 13040 892 13070 996
rect 13128 892 13158 996
rect 13316 892 13346 1022
rect 13400 892 13430 1022
rect 13484 892 13514 1022
rect 13568 892 13598 1022
rect 13652 892 13682 1022
rect 13868 892 13898 1022
rect 13952 892 13982 1022
rect 14036 892 14066 1022
rect 14120 892 14150 1022
rect 14204 892 14234 1022
rect 14288 892 14318 1022
rect 14372 892 14402 1022
rect 14456 892 14486 1022
rect 14540 892 14570 1022
rect 14624 892 14654 1022
rect 14708 892 14738 1022
rect 14792 892 14822 1022
rect 14876 892 14906 1022
rect 14960 892 14990 1022
rect 15044 892 15074 1022
rect 15128 892 15158 1022
rect 15212 892 15242 1022
rect 15296 892 15326 1022
rect 15380 892 15410 1022
rect 15464 892 15494 1022
rect 15548 892 15578 1022
rect 15632 892 15662 1022
rect 8654 -250 8684 -120
rect 8763 -250 8793 -166
rect 8859 -250 8889 -166
rect 8984 -250 9014 -166
rect 9080 -250 9110 -166
rect 9248 -250 9278 -166
rect 10134 -250 10164 -166
rect 10302 -250 10332 -166
rect 10398 -250 10428 -166
rect 10523 -250 10553 -166
rect 10619 -250 10649 -166
rect 10728 -250 10758 -120
rect 11046 -250 11076 -120
rect 11155 -250 11185 -166
rect 11251 -250 11281 -166
rect 11376 -250 11406 -166
rect 11472 -250 11502 -166
rect 11640 -250 11670 -166
rect 12526 -250 12556 -166
rect 12694 -250 12724 -166
rect 12790 -250 12820 -166
rect 12915 -250 12945 -166
rect 13011 -250 13041 -166
rect 13120 -250 13150 -120
rect 13438 -250 13468 -120
rect 13547 -250 13577 -166
rect 13643 -250 13673 -166
rect 13768 -250 13798 -166
rect 13864 -250 13894 -166
rect 14032 -250 14062 -166
rect 14916 -250 14946 -166
rect 15084 -250 15114 -166
rect 15180 -250 15210 -166
rect 15305 -250 15335 -166
rect 15401 -250 15431 -166
rect 15510 -250 15540 -120
rect 15830 -250 15860 -120
rect 15939 -250 15969 -166
rect 16035 -250 16065 -166
rect 16160 -250 16190 -166
rect 16256 -250 16286 -166
rect 16424 -250 16454 -166
rect 17310 -250 17340 -166
rect 17478 -250 17508 -166
rect 17574 -250 17604 -166
rect 17699 -250 17729 -166
rect 17795 -250 17825 -166
rect 17904 -250 17934 -120
rect 18222 -250 18252 -120
rect 18331 -250 18361 -166
rect 18427 -250 18457 -166
rect 18552 -250 18582 -166
rect 18648 -250 18678 -166
rect 18816 -250 18846 -166
rect 19702 -250 19732 -166
rect 19870 -250 19900 -166
rect 19966 -250 19996 -166
rect 20091 -250 20121 -166
rect 20187 -250 20217 -166
rect 20296 -250 20326 -120
rect 20614 -250 20644 -120
rect 20723 -250 20753 -166
rect 20819 -250 20849 -166
rect 20944 -250 20974 -166
rect 21040 -250 21070 -166
rect 21208 -250 21238 -166
rect 22092 -250 22122 -166
rect 22260 -250 22290 -166
rect 22356 -250 22386 -166
rect 22481 -250 22511 -166
rect 22577 -250 22607 -166
rect 22686 -250 22716 -120
rect 23006 -250 23036 -120
rect 23115 -250 23145 -166
rect 23211 -250 23241 -166
rect 23336 -250 23366 -166
rect 23432 -250 23462 -166
rect 23600 -250 23630 -166
rect 24486 -250 24516 -166
rect 24654 -250 24684 -166
rect 24750 -250 24780 -166
rect 24875 -250 24905 -166
rect 24971 -250 25001 -166
rect 25080 -250 25110 -120
rect 8654 -938 8684 -854
rect 8738 -938 8768 -854
rect 8926 -938 8956 -854
rect 9021 -938 9051 -866
rect 9126 -938 9156 -866
rect 9222 -938 9252 -854
rect 9336 -938 9366 -854
rect 9432 -938 9462 -810
rect 9516 -938 9546 -810
rect 9704 -938 9734 -810
rect 9824 -938 9854 -866
rect 9908 -938 9938 -866
rect 10003 -938 10033 -854
rect 10100 -938 10130 -854
rect 10208 -938 10238 -810
rect 10292 -938 10322 -810
rect 10480 -938 10510 -854
rect 10575 -938 10605 -808
rect 10763 -938 10793 -854
rect 10858 -938 10888 -808
rect 11046 -938 11076 -854
rect 11130 -938 11160 -854
rect 11318 -938 11348 -854
rect 11413 -938 11443 -866
rect 11518 -938 11548 -866
rect 11614 -938 11644 -854
rect 11728 -938 11758 -854
rect 11824 -938 11854 -810
rect 11908 -938 11938 -810
rect 12096 -938 12126 -810
rect 12216 -938 12246 -866
rect 12300 -938 12330 -866
rect 12395 -938 12425 -854
rect 12492 -938 12522 -854
rect 12600 -938 12630 -810
rect 12684 -938 12714 -810
rect 12872 -938 12902 -854
rect 12967 -938 12997 -808
rect 13155 -938 13185 -854
rect 13250 -938 13280 -808
rect 13438 -938 13468 -854
rect 13522 -938 13552 -854
rect 13710 -938 13740 -854
rect 13805 -938 13835 -866
rect 13910 -938 13940 -866
rect 14006 -938 14036 -854
rect 14120 -938 14150 -854
rect 14216 -938 14246 -810
rect 14300 -938 14330 -810
rect 14488 -938 14518 -810
rect 14608 -938 14638 -866
rect 14692 -938 14722 -866
rect 14787 -938 14817 -854
rect 14884 -938 14914 -854
rect 14992 -938 15022 -810
rect 15076 -938 15106 -810
rect 15264 -938 15294 -854
rect 15359 -938 15389 -808
rect 15547 -938 15577 -854
rect 15642 -938 15672 -808
rect 15830 -938 15860 -854
rect 15914 -938 15944 -854
rect 16102 -938 16132 -854
rect 16197 -938 16227 -866
rect 16302 -938 16332 -866
rect 16398 -938 16428 -854
rect 16512 -938 16542 -854
rect 16608 -938 16638 -810
rect 16692 -938 16722 -810
rect 16880 -938 16910 -810
rect 17000 -938 17030 -866
rect 17084 -938 17114 -866
rect 17179 -938 17209 -854
rect 17276 -938 17306 -854
rect 17384 -938 17414 -810
rect 17468 -938 17498 -810
rect 17656 -938 17686 -854
rect 17751 -938 17781 -808
rect 17939 -938 17969 -854
rect 18034 -938 18064 -808
rect 18222 -938 18252 -854
rect 18306 -938 18336 -854
rect 18494 -938 18524 -854
rect 18589 -938 18619 -866
rect 18694 -938 18724 -866
rect 18790 -938 18820 -854
rect 18904 -938 18934 -854
rect 19000 -938 19030 -810
rect 19084 -938 19114 -810
rect 19272 -938 19302 -810
rect 19392 -938 19422 -866
rect 19476 -938 19506 -866
rect 19571 -938 19601 -854
rect 19668 -938 19698 -854
rect 19776 -938 19806 -810
rect 19860 -938 19890 -810
rect 20048 -938 20078 -854
rect 20143 -938 20173 -808
rect 20331 -938 20361 -854
rect 20426 -938 20456 -808
rect 20614 -938 20644 -854
rect 20698 -938 20728 -854
rect 20886 -938 20916 -854
rect 20981 -938 21011 -866
rect 21086 -938 21116 -866
rect 21182 -938 21212 -854
rect 21296 -938 21326 -854
rect 21392 -938 21422 -810
rect 21476 -938 21506 -810
rect 21664 -938 21694 -810
rect 21784 -938 21814 -866
rect 21868 -938 21898 -866
rect 21963 -938 21993 -854
rect 22060 -938 22090 -854
rect 22168 -938 22198 -810
rect 22252 -938 22282 -810
rect 22440 -938 22470 -854
rect 22535 -938 22565 -808
rect 22723 -938 22753 -854
rect 22818 -938 22848 -808
rect 23006 -938 23036 -854
rect 23090 -938 23120 -854
rect 23278 -938 23308 -854
rect 23373 -938 23403 -866
rect 23478 -938 23508 -866
rect 23574 -938 23604 -854
rect 23688 -938 23718 -854
rect 23784 -938 23814 -810
rect 23868 -938 23898 -810
rect 24056 -938 24086 -810
rect 24176 -938 24206 -866
rect 24260 -938 24290 -866
rect 24355 -938 24385 -854
rect 24452 -938 24482 -854
rect 24560 -938 24590 -810
rect 24644 -938 24674 -810
rect 24832 -938 24862 -854
rect 24927 -938 24957 -808
rect 25115 -938 25145 -854
rect 25210 -938 25240 -808
rect 8654 -1627 8684 -1497
rect 8749 -1627 8779 -1543
rect 8937 -1627 8967 -1497
rect 9032 -1627 9062 -1543
rect 9220 -1627 9250 -1499
rect 9304 -1627 9334 -1499
rect 9412 -1627 9442 -1543
rect 9509 -1627 9539 -1543
rect 9604 -1627 9634 -1555
rect 9688 -1627 9718 -1555
rect 9808 -1627 9838 -1499
rect 9996 -1627 10026 -1499
rect 10080 -1627 10110 -1499
rect 10176 -1627 10206 -1543
rect 10290 -1627 10320 -1543
rect 10386 -1627 10416 -1555
rect 10491 -1627 10521 -1555
rect 10586 -1627 10616 -1543
rect 10774 -1627 10804 -1543
rect 10858 -1627 10888 -1543
rect 11046 -1627 11076 -1497
rect 11141 -1627 11171 -1543
rect 11329 -1627 11359 -1497
rect 11424 -1627 11454 -1543
rect 11612 -1627 11642 -1499
rect 11696 -1627 11726 -1499
rect 11804 -1627 11834 -1543
rect 11901 -1627 11931 -1543
rect 11996 -1627 12026 -1555
rect 12080 -1627 12110 -1555
rect 12200 -1627 12230 -1499
rect 12388 -1627 12418 -1499
rect 12472 -1627 12502 -1499
rect 12568 -1627 12598 -1543
rect 12682 -1627 12712 -1543
rect 12778 -1627 12808 -1555
rect 12883 -1627 12913 -1555
rect 12978 -1627 13008 -1543
rect 13166 -1627 13196 -1543
rect 13250 -1627 13280 -1543
rect 13438 -1627 13468 -1497
rect 13533 -1627 13563 -1543
rect 13721 -1627 13751 -1497
rect 13816 -1627 13846 -1543
rect 14004 -1627 14034 -1499
rect 14088 -1627 14118 -1499
rect 14196 -1627 14226 -1543
rect 14293 -1627 14323 -1543
rect 14388 -1627 14418 -1555
rect 14472 -1627 14502 -1555
rect 14592 -1627 14622 -1499
rect 14780 -1627 14810 -1499
rect 14864 -1627 14894 -1499
rect 14960 -1627 14990 -1543
rect 15074 -1627 15104 -1543
rect 15170 -1627 15200 -1555
rect 15275 -1627 15305 -1555
rect 15370 -1627 15400 -1543
rect 15558 -1627 15588 -1543
rect 15642 -1627 15672 -1543
rect 15830 -1627 15860 -1497
rect 15925 -1627 15955 -1543
rect 16113 -1627 16143 -1497
rect 16208 -1627 16238 -1543
rect 16396 -1627 16426 -1499
rect 16480 -1627 16510 -1499
rect 16588 -1627 16618 -1543
rect 16685 -1627 16715 -1543
rect 16780 -1627 16810 -1555
rect 16864 -1627 16894 -1555
rect 16984 -1627 17014 -1499
rect 17172 -1627 17202 -1499
rect 17256 -1627 17286 -1499
rect 17352 -1627 17382 -1543
rect 17466 -1627 17496 -1543
rect 17562 -1627 17592 -1555
rect 17667 -1627 17697 -1555
rect 17762 -1627 17792 -1543
rect 17950 -1627 17980 -1543
rect 18034 -1627 18064 -1543
rect 18222 -1627 18252 -1497
rect 18317 -1627 18347 -1543
rect 18505 -1627 18535 -1497
rect 18600 -1627 18630 -1543
rect 18788 -1627 18818 -1499
rect 18872 -1627 18902 -1499
rect 18980 -1627 19010 -1543
rect 19077 -1627 19107 -1543
rect 19172 -1627 19202 -1555
rect 19256 -1627 19286 -1555
rect 19376 -1627 19406 -1499
rect 19564 -1627 19594 -1499
rect 19648 -1627 19678 -1499
rect 19744 -1627 19774 -1543
rect 19858 -1627 19888 -1543
rect 19954 -1627 19984 -1555
rect 20059 -1627 20089 -1555
rect 20154 -1627 20184 -1543
rect 20342 -1627 20372 -1543
rect 20426 -1627 20456 -1543
rect 20614 -1627 20644 -1497
rect 20709 -1627 20739 -1543
rect 20897 -1627 20927 -1497
rect 20992 -1627 21022 -1543
rect 21180 -1627 21210 -1499
rect 21264 -1627 21294 -1499
rect 21372 -1627 21402 -1543
rect 21469 -1627 21499 -1543
rect 21564 -1627 21594 -1555
rect 21648 -1627 21678 -1555
rect 21768 -1627 21798 -1499
rect 21956 -1627 21986 -1499
rect 22040 -1627 22070 -1499
rect 22136 -1627 22166 -1543
rect 22250 -1627 22280 -1543
rect 22346 -1627 22376 -1555
rect 22451 -1627 22481 -1555
rect 22546 -1627 22576 -1543
rect 22734 -1627 22764 -1543
rect 22818 -1627 22848 -1543
rect 23006 -1627 23036 -1497
rect 23101 -1627 23131 -1543
rect 23289 -1627 23319 -1497
rect 23384 -1627 23414 -1543
rect 23572 -1627 23602 -1499
rect 23656 -1627 23686 -1499
rect 23764 -1627 23794 -1543
rect 23861 -1627 23891 -1543
rect 23956 -1627 23986 -1555
rect 24040 -1627 24070 -1555
rect 24160 -1627 24190 -1499
rect 24348 -1627 24378 -1499
rect 24432 -1627 24462 -1499
rect 24528 -1627 24558 -1543
rect 24642 -1627 24672 -1543
rect 24738 -1627 24768 -1555
rect 24843 -1627 24873 -1555
rect 24938 -1627 24968 -1543
rect 25126 -1627 25156 -1543
rect 25210 -1627 25240 -1543
<< pmos >>
rect 3616 11889 3646 11973
rect 4348 11892 4378 11976
rect 4474 11892 4504 11976
rect 5560 11892 5590 11976
rect 5686 11892 5716 11976
rect 6772 11892 6802 11976
rect 6898 11892 6928 11976
rect 7984 11892 8014 11976
rect 8110 11892 8140 11976
rect 14504 12364 14534 12448
rect 15236 12367 15266 12451
rect 15362 12367 15392 12451
rect 16448 12367 16478 12451
rect 16574 12367 16604 12451
rect 17660 12367 17690 12451
rect 17786 12367 17816 12451
rect 18872 12367 18902 12451
rect 18998 12367 19028 12451
rect 21213 12364 21243 12448
rect 21945 12367 21975 12451
rect 22071 12367 22101 12451
rect 23157 12367 23187 12451
rect 23283 12367 23313 12451
rect 24369 12367 24399 12451
rect 24495 12367 24525 12451
rect 25581 12367 25611 12451
rect 25707 12367 25737 12451
rect 3616 8673 3646 8757
rect 4348 8670 4378 8754
rect 4474 8670 4504 8754
rect 5560 8670 5590 8754
rect 5686 8670 5716 8754
rect 6772 8670 6802 8754
rect 6898 8670 6928 8754
rect 7984 8670 8014 8754
rect 8110 8670 8140 8754
rect 11883 8488 11913 8740
rect 11979 8488 12009 8740
rect 12075 8488 12105 8740
rect 12279 8489 12309 8741
rect 12480 8460 12510 8740
rect 14151 8658 14181 8742
rect 14277 8658 14307 8742
rect 15363 8658 15393 8742
rect 15489 8658 15519 8742
rect 16575 8658 16605 8742
rect 16701 8658 16731 8742
rect 17787 8658 17817 8742
rect 17913 8658 17943 8742
rect 18645 8661 18675 8745
rect 20860 8658 20890 8742
rect 20986 8658 21016 8742
rect 22072 8658 22102 8742
rect 22198 8658 22228 8742
rect 23284 8658 23314 8742
rect 23410 8658 23440 8742
rect 24496 8658 24526 8742
rect 24622 8658 24652 8742
rect 25354 8661 25384 8745
rect 11883 8084 11913 8336
rect 11979 8084 12009 8336
rect 12075 8084 12105 8336
rect 12279 8083 12309 8335
rect 12748 7584 12778 7964
rect 25229 6067 25259 6151
rect 25961 6070 25991 6154
rect 26087 6070 26117 6154
rect 27173 6070 27203 6154
rect 27299 6070 27329 6154
rect 28385 6070 28415 6154
rect 28511 6070 28541 6154
rect 29597 6070 29627 6154
rect 29723 6070 29753 6154
<< scpmoshvt >>
rect 13394 12746 13424 12946
rect 13584 12746 13614 12946
rect 20103 12746 20133 12946
rect 20293 12746 20323 12946
rect 2506 12271 2536 12471
rect 2696 12271 2726 12471
rect 9181 11894 9211 12094
rect 10961 11958 10991 12086
rect 11045 11958 11075 12086
rect 11233 11952 11263 12036
rect 11326 11952 11356 12036
rect 11410 11952 11440 12036
rect 11530 11952 11560 12036
rect 11636 11952 11666 12036
rect 11744 11952 11774 12120
rect 11828 11952 11858 12120
rect 11965 11952 11995 12120
rect 12109 11952 12139 12036
rect 12193 11952 12223 12036
rect 12311 11952 12341 12036
rect 12419 11952 12449 12036
rect 12515 11952 12545 12120
rect 12587 11952 12617 12120
rect 12785 12020 12815 12148
rect 12882 11952 12912 12152
rect 13070 11968 13100 12096
rect 13165 11952 13195 12152
rect 11002 11562 11032 11762
rect 11278 11562 11308 11762
rect 9181 8554 9211 8754
rect 9396 8554 9426 8754
rect 9491 8570 9521 8698
rect 9679 8554 9709 8754
rect 9776 8622 9806 8750
rect 9974 8554 10004 8722
rect 10046 8554 10076 8722
rect 10142 8554 10172 8638
rect 10250 8554 10280 8638
rect 10368 8554 10398 8638
rect 10452 8554 10482 8638
rect 10596 8554 10626 8722
rect 10733 8554 10763 8722
rect 10817 8554 10847 8722
rect 10925 8554 10955 8638
rect 11031 8554 11061 8638
rect 11151 8554 11181 8638
rect 11235 8554 11265 8638
rect 11328 8554 11358 8638
rect 11516 8560 11546 8688
rect 11600 8560 11630 8688
rect 12728 8541 12758 8741
rect 12812 8541 12842 8741
rect 13051 8541 13081 8741
rect 2506 8175 2536 8375
rect 2696 8175 2726 8375
rect 10133 8085 10163 8285
rect 10242 8162 10272 8246
rect 10345 8162 10375 8246
rect 10559 8162 10589 8246
rect 10631 8162 10661 8246
rect 10727 8162 10757 8246
rect 10960 8085 10990 8285
rect 11069 8162 11099 8246
rect 11172 8162 11202 8246
rect 11386 8162 11416 8246
rect 11458 8162 11488 8246
rect 11554 8162 11584 8246
rect 19565 8163 19595 8363
rect 19755 8163 19785 8363
rect 26274 8163 26304 8363
rect 26464 8163 26494 8363
rect 11577 6872 11607 7030
rect 11665 6872 11695 7030
rect 11853 6830 11883 7030
rect 11937 6830 11967 7030
rect 12021 6830 12051 7030
rect 12105 6830 12135 7030
rect 12189 6830 12219 7030
rect 12852 6830 12882 7030
rect 12936 6830 12966 7030
rect 13036 6830 13066 7030
rect 13120 6830 13150 7030
rect 13217 6902 13247 7030
rect 13318 6946 13348 7030
rect 13402 6946 13432 7030
rect 13537 6902 13567 7030
rect 13725 6849 13755 6957
rect 13809 6849 13839 6957
rect 13997 6878 14027 7006
rect 14081 6878 14111 7006
rect 14225 6946 14255 7030
rect 14309 6946 14339 7030
rect 14405 6902 14435 7030
rect 14489 6902 14519 7030
rect 24119 6449 24149 6649
rect 24309 6449 24339 6649
rect 11576 6023 11606 6151
rect 11660 6023 11690 6151
rect 11848 6073 11878 6157
rect 11941 6073 11971 6157
rect 12025 6073 12055 6157
rect 12145 6073 12175 6157
rect 12251 6073 12281 6157
rect 12359 5989 12389 6157
rect 12443 5989 12473 6157
rect 12580 5989 12610 6157
rect 12724 6073 12754 6157
rect 12808 6073 12838 6157
rect 12926 6073 12956 6157
rect 13034 6073 13064 6157
rect 13130 5989 13160 6157
rect 13202 5989 13232 6157
rect 13400 5961 13430 6089
rect 13497 5957 13527 6157
rect 13685 6013 13715 6141
rect 13780 5957 13810 6157
rect 13968 6023 13998 6151
rect 14052 6023 14082 6151
rect 14240 6073 14270 6157
rect 14333 6073 14363 6157
rect 14417 6073 14447 6157
rect 14537 6073 14567 6157
rect 14643 6073 14673 6157
rect 14751 5989 14781 6157
rect 14835 5989 14865 6157
rect 14972 5989 15002 6157
rect 15116 6073 15146 6157
rect 15200 6073 15230 6157
rect 15318 6073 15348 6157
rect 15426 6073 15456 6157
rect 15522 5989 15552 6157
rect 15594 5989 15624 6157
rect 15792 5961 15822 6089
rect 15889 5957 15919 6157
rect 16077 6013 16107 6141
rect 16172 5957 16202 6157
rect 16360 6023 16390 6151
rect 16444 6023 16474 6151
rect 16632 6073 16662 6157
rect 16725 6073 16755 6157
rect 16809 6073 16839 6157
rect 16929 6073 16959 6157
rect 17035 6073 17065 6157
rect 17143 5989 17173 6157
rect 17227 5989 17257 6157
rect 17364 5989 17394 6157
rect 17508 6073 17538 6157
rect 17592 6073 17622 6157
rect 17710 6073 17740 6157
rect 17818 6073 17848 6157
rect 17914 5989 17944 6157
rect 17986 5989 18016 6157
rect 18184 5961 18214 6089
rect 18281 5957 18311 6157
rect 18469 6013 18499 6141
rect 18564 5957 18594 6157
rect 18752 6023 18782 6151
rect 18836 6023 18866 6151
rect 19024 6073 19054 6157
rect 19117 6073 19147 6157
rect 19201 6073 19231 6157
rect 19321 6073 19351 6157
rect 19427 6073 19457 6157
rect 19535 5989 19565 6157
rect 19619 5989 19649 6157
rect 19756 5989 19786 6157
rect 19900 6073 19930 6157
rect 19984 6073 20014 6157
rect 20102 6073 20132 6157
rect 20210 6073 20240 6157
rect 20306 5989 20336 6157
rect 20378 5989 20408 6157
rect 20576 5961 20606 6089
rect 20673 5957 20703 6157
rect 20861 6013 20891 6141
rect 20956 5957 20986 6157
rect 21144 6023 21174 6151
rect 21228 6023 21258 6151
rect 21416 6073 21446 6157
rect 21509 6073 21539 6157
rect 21593 6073 21623 6157
rect 21713 6073 21743 6157
rect 21819 6073 21849 6157
rect 21927 5989 21957 6157
rect 22011 5989 22041 6157
rect 22148 5989 22178 6157
rect 22292 6073 22322 6157
rect 22376 6073 22406 6157
rect 22494 6073 22524 6157
rect 22602 6073 22632 6157
rect 22698 5989 22728 6157
rect 22770 5989 22800 6157
rect 22968 5961 22998 6089
rect 23065 5957 23095 6157
rect 23253 6013 23283 6141
rect 23348 5957 23378 6157
rect 30758 6136 30788 6264
rect 30853 6072 30883 6272
rect 30937 6072 30967 6272
rect 11136 5310 11166 5468
rect 11224 5310 11254 5468
rect 11412 5268 11442 5468
rect 11496 5268 11526 5468
rect 11580 5268 11610 5468
rect 11664 5268 11694 5468
rect 11748 5268 11778 5468
rect 11944 5268 11974 5468
rect 12028 5268 12058 5468
rect 12112 5268 12142 5468
rect 12196 5268 12226 5468
rect 12280 5268 12310 5468
rect 12364 5268 12394 5468
rect 12448 5268 12478 5468
rect 12532 5268 12562 5468
rect 12616 5268 12646 5468
rect 12700 5268 12730 5468
rect 12784 5268 12814 5468
rect 12868 5268 12898 5468
rect 12952 5268 12982 5468
rect 13036 5268 13066 5468
rect 13120 5268 13150 5468
rect 13204 5268 13234 5468
rect 13288 5268 13318 5468
rect 13372 5268 13402 5468
rect 13456 5268 13486 5468
rect 13540 5268 13570 5468
rect 13624 5268 13654 5468
rect 13708 5268 13738 5468
rect 13968 5268 13998 5468
rect 14063 5324 14093 5452
rect 14251 5268 14281 5468
rect 14348 5272 14378 5400
rect 14546 5300 14576 5468
rect 14618 5300 14648 5468
rect 14714 5384 14744 5468
rect 14822 5384 14852 5468
rect 14940 5384 14970 5468
rect 15024 5384 15054 5468
rect 15168 5300 15198 5468
rect 15305 5300 15335 5468
rect 15389 5300 15419 5468
rect 15497 5384 15527 5468
rect 15603 5384 15633 5468
rect 15723 5384 15753 5468
rect 15807 5384 15837 5468
rect 15900 5384 15930 5468
rect 16088 5334 16118 5462
rect 16172 5334 16202 5462
rect 16360 5268 16390 5468
rect 16455 5324 16485 5452
rect 16643 5268 16673 5468
rect 16740 5272 16770 5400
rect 16938 5300 16968 5468
rect 17010 5300 17040 5468
rect 17106 5384 17136 5468
rect 17214 5384 17244 5468
rect 17332 5384 17362 5468
rect 17416 5384 17446 5468
rect 17560 5300 17590 5468
rect 17697 5300 17727 5468
rect 17781 5300 17811 5468
rect 17889 5384 17919 5468
rect 17995 5384 18025 5468
rect 18115 5384 18145 5468
rect 18199 5384 18229 5468
rect 18292 5384 18322 5468
rect 18480 5334 18510 5462
rect 18564 5334 18594 5462
rect 18752 5268 18782 5468
rect 18847 5324 18877 5452
rect 19035 5268 19065 5468
rect 19132 5272 19162 5400
rect 19330 5300 19360 5468
rect 19402 5300 19432 5468
rect 19498 5384 19528 5468
rect 19606 5384 19636 5468
rect 19724 5384 19754 5468
rect 19808 5384 19838 5468
rect 19952 5300 19982 5468
rect 20089 5300 20119 5468
rect 20173 5300 20203 5468
rect 20281 5384 20311 5468
rect 20387 5384 20417 5468
rect 20507 5384 20537 5468
rect 20591 5384 20621 5468
rect 20684 5384 20714 5468
rect 20872 5334 20902 5462
rect 20956 5334 20986 5462
rect 21144 5268 21174 5468
rect 21239 5324 21269 5452
rect 21427 5268 21457 5468
rect 21524 5272 21554 5400
rect 21722 5300 21752 5468
rect 21794 5300 21824 5468
rect 21890 5384 21920 5468
rect 21998 5384 22028 5468
rect 22116 5384 22146 5468
rect 22200 5384 22230 5468
rect 22344 5300 22374 5468
rect 22481 5300 22511 5468
rect 22565 5300 22595 5468
rect 22673 5384 22703 5468
rect 22779 5384 22809 5468
rect 22899 5384 22929 5468
rect 22983 5384 23013 5468
rect 23076 5384 23106 5468
rect 23264 5334 23294 5462
rect 23348 5334 23378 5462
rect 11168 4436 11198 4594
rect 11256 4436 11286 4594
rect 11444 4394 11474 4594
rect 11528 4394 11558 4594
rect 11612 4394 11642 4594
rect 11696 4394 11726 4594
rect 11780 4394 11810 4594
rect 13751 4395 13781 4595
rect 13967 4461 13997 4589
rect 14051 4461 14081 4589
rect 14239 4511 14269 4595
rect 14332 4511 14362 4595
rect 14416 4511 14446 4595
rect 14536 4511 14566 4595
rect 14642 4511 14672 4595
rect 14750 4427 14780 4595
rect 14834 4427 14864 4595
rect 14971 4427 15001 4595
rect 15115 4511 15145 4595
rect 15199 4511 15229 4595
rect 15317 4511 15347 4595
rect 15425 4511 15455 4595
rect 15521 4427 15551 4595
rect 15593 4427 15623 4595
rect 15791 4399 15821 4527
rect 15888 4395 15918 4595
rect 16076 4451 16106 4579
rect 16171 4395 16201 4595
rect 16359 4461 16389 4589
rect 16443 4461 16473 4589
rect 16631 4511 16661 4595
rect 16724 4511 16754 4595
rect 16808 4511 16838 4595
rect 16928 4511 16958 4595
rect 17034 4511 17064 4595
rect 17142 4427 17172 4595
rect 17226 4427 17256 4595
rect 17363 4427 17393 4595
rect 17507 4511 17537 4595
rect 17591 4511 17621 4595
rect 17709 4511 17739 4595
rect 17817 4511 17847 4595
rect 17913 4427 17943 4595
rect 17985 4427 18015 4595
rect 18183 4399 18213 4527
rect 18280 4395 18310 4595
rect 18468 4451 18498 4579
rect 18563 4395 18593 4595
rect 18751 4461 18781 4589
rect 18835 4461 18865 4589
rect 19023 4511 19053 4595
rect 19116 4511 19146 4595
rect 19200 4511 19230 4595
rect 19320 4511 19350 4595
rect 19426 4511 19456 4595
rect 19534 4427 19564 4595
rect 19618 4427 19648 4595
rect 19755 4427 19785 4595
rect 19899 4511 19929 4595
rect 19983 4511 20013 4595
rect 20101 4511 20131 4595
rect 20209 4511 20239 4595
rect 20305 4427 20335 4595
rect 20377 4427 20407 4595
rect 20575 4399 20605 4527
rect 20672 4395 20702 4595
rect 20860 4451 20890 4579
rect 20955 4395 20985 4595
rect 21143 4461 21173 4589
rect 21227 4461 21257 4589
rect 21415 4511 21445 4595
rect 21508 4511 21538 4595
rect 21592 4511 21622 4595
rect 21712 4511 21742 4595
rect 21818 4511 21848 4595
rect 21926 4427 21956 4595
rect 22010 4427 22040 4595
rect 22147 4427 22177 4595
rect 22291 4511 22321 4595
rect 22375 4511 22405 4595
rect 22493 4511 22523 4595
rect 22601 4511 22631 4595
rect 22697 4427 22727 4595
rect 22769 4427 22799 4595
rect 22967 4399 22997 4527
rect 23064 4395 23094 4595
rect 23252 4451 23282 4579
rect 23347 4395 23377 4595
rect 25656 3790 25686 3918
rect 25740 3790 25770 3918
rect 25928 3784 25958 3868
rect 26021 3784 26051 3868
rect 26105 3784 26135 3868
rect 26225 3784 26255 3868
rect 26331 3784 26361 3868
rect 26439 3784 26469 3952
rect 26523 3784 26553 3952
rect 26660 3784 26690 3952
rect 26804 3784 26834 3868
rect 26888 3784 26918 3868
rect 27006 3784 27036 3868
rect 27114 3784 27144 3868
rect 27210 3784 27240 3952
rect 27282 3784 27312 3952
rect 27480 3852 27510 3980
rect 27577 3784 27607 3984
rect 27765 3800 27795 3928
rect 27860 3784 27890 3984
rect 28048 3790 28078 3918
rect 28132 3790 28162 3918
rect 28320 3784 28350 3868
rect 28413 3784 28443 3868
rect 28497 3784 28527 3868
rect 28617 3784 28647 3868
rect 28723 3784 28753 3868
rect 28831 3784 28861 3952
rect 28915 3784 28945 3952
rect 29052 3784 29082 3952
rect 29196 3784 29226 3868
rect 29280 3784 29310 3868
rect 29398 3784 29428 3868
rect 29506 3784 29536 3868
rect 29602 3784 29632 3952
rect 29674 3784 29704 3952
rect 29872 3852 29902 3980
rect 29969 3784 29999 3984
rect 30157 3800 30187 3928
rect 30252 3784 30282 3984
rect 11575 3522 11605 3722
rect 11670 3578 11700 3706
rect 11858 3522 11888 3722
rect 11955 3526 11985 3654
rect 12153 3554 12183 3722
rect 12225 3554 12255 3722
rect 12321 3638 12351 3722
rect 12429 3638 12459 3722
rect 12547 3638 12577 3722
rect 12631 3638 12661 3722
rect 12775 3554 12805 3722
rect 12912 3554 12942 3722
rect 12996 3554 13026 3722
rect 13104 3638 13134 3722
rect 13210 3638 13240 3722
rect 13330 3638 13360 3722
rect 13414 3638 13444 3722
rect 13507 3638 13537 3722
rect 13695 3588 13725 3716
rect 13779 3588 13809 3716
rect 13967 3522 13997 3722
rect 14062 3578 14092 3706
rect 14250 3522 14280 3722
rect 14347 3526 14377 3654
rect 14545 3554 14575 3722
rect 14617 3554 14647 3722
rect 14713 3638 14743 3722
rect 14821 3638 14851 3722
rect 14939 3638 14969 3722
rect 15023 3638 15053 3722
rect 15167 3554 15197 3722
rect 15304 3554 15334 3722
rect 15388 3554 15418 3722
rect 15496 3638 15526 3722
rect 15602 3638 15632 3722
rect 15722 3638 15752 3722
rect 15806 3638 15836 3722
rect 15899 3638 15929 3722
rect 16087 3588 16117 3716
rect 16171 3588 16201 3716
rect 16359 3522 16389 3722
rect 16454 3578 16484 3706
rect 16642 3522 16672 3722
rect 16739 3526 16769 3654
rect 16937 3554 16967 3722
rect 17009 3554 17039 3722
rect 17105 3638 17135 3722
rect 17213 3638 17243 3722
rect 17331 3638 17361 3722
rect 17415 3638 17445 3722
rect 17559 3554 17589 3722
rect 17696 3554 17726 3722
rect 17780 3554 17810 3722
rect 17888 3638 17918 3722
rect 17994 3638 18024 3722
rect 18114 3638 18144 3722
rect 18198 3638 18228 3722
rect 18291 3638 18321 3722
rect 18479 3588 18509 3716
rect 18563 3588 18593 3716
rect 18751 3522 18781 3722
rect 18846 3578 18876 3706
rect 19034 3522 19064 3722
rect 19131 3526 19161 3654
rect 19329 3554 19359 3722
rect 19401 3554 19431 3722
rect 19497 3638 19527 3722
rect 19605 3638 19635 3722
rect 19723 3638 19753 3722
rect 19807 3638 19837 3722
rect 19951 3554 19981 3722
rect 20088 3554 20118 3722
rect 20172 3554 20202 3722
rect 20280 3638 20310 3722
rect 20386 3638 20416 3722
rect 20506 3638 20536 3722
rect 20590 3638 20620 3722
rect 20683 3638 20713 3722
rect 20871 3588 20901 3716
rect 20955 3588 20985 3716
rect 21143 3522 21173 3722
rect 21238 3578 21268 3706
rect 21426 3522 21456 3722
rect 21523 3526 21553 3654
rect 21721 3554 21751 3722
rect 21793 3554 21823 3722
rect 21889 3638 21919 3722
rect 21997 3638 22027 3722
rect 22115 3638 22145 3722
rect 22199 3638 22229 3722
rect 22343 3554 22373 3722
rect 22480 3554 22510 3722
rect 22564 3554 22594 3722
rect 22672 3638 22702 3722
rect 22778 3638 22808 3722
rect 22898 3638 22928 3722
rect 22982 3638 23012 3722
rect 23075 3638 23105 3722
rect 23263 3588 23293 3716
rect 23347 3588 23377 3716
rect 25656 3460 25686 3588
rect 25740 3460 25770 3588
rect 25928 3510 25958 3594
rect 26021 3510 26051 3594
rect 26105 3510 26135 3594
rect 26225 3510 26255 3594
rect 26331 3510 26361 3594
rect 26439 3426 26469 3594
rect 26523 3426 26553 3594
rect 26660 3426 26690 3594
rect 26804 3510 26834 3594
rect 26888 3510 26918 3594
rect 27006 3510 27036 3594
rect 27114 3510 27144 3594
rect 27210 3426 27240 3594
rect 27282 3426 27312 3594
rect 27480 3398 27510 3526
rect 27577 3394 27607 3594
rect 27765 3450 27795 3578
rect 27860 3394 27890 3594
rect 28048 3460 28078 3588
rect 28132 3460 28162 3588
rect 28320 3510 28350 3594
rect 28413 3510 28443 3594
rect 28497 3510 28527 3594
rect 28617 3510 28647 3594
rect 28723 3510 28753 3594
rect 28831 3426 28861 3594
rect 28915 3426 28945 3594
rect 29052 3426 29082 3594
rect 29196 3510 29226 3594
rect 29280 3510 29310 3594
rect 29398 3510 29428 3594
rect 29506 3510 29536 3594
rect 29602 3426 29632 3594
rect 29674 3426 29704 3594
rect 29872 3398 29902 3526
rect 29969 3394 29999 3594
rect 30157 3450 30187 3578
rect 30252 3394 30282 3594
rect 25656 2510 25686 2638
rect 25740 2510 25770 2638
rect 25928 2504 25958 2588
rect 26021 2504 26051 2588
rect 26105 2504 26135 2588
rect 26225 2504 26255 2588
rect 26331 2504 26361 2588
rect 26439 2504 26469 2672
rect 26523 2504 26553 2672
rect 26660 2504 26690 2672
rect 26804 2504 26834 2588
rect 26888 2504 26918 2588
rect 27006 2504 27036 2588
rect 27114 2504 27144 2588
rect 27210 2504 27240 2672
rect 27282 2504 27312 2672
rect 27480 2572 27510 2700
rect 27577 2504 27607 2704
rect 27765 2520 27795 2648
rect 27860 2504 27890 2704
rect 28048 2510 28078 2638
rect 28132 2510 28162 2638
rect 28320 2504 28350 2588
rect 28413 2504 28443 2588
rect 28497 2504 28527 2588
rect 28617 2504 28647 2588
rect 28723 2504 28753 2588
rect 28831 2504 28861 2672
rect 28915 2504 28945 2672
rect 29052 2504 29082 2672
rect 29196 2504 29226 2588
rect 29280 2504 29310 2588
rect 29398 2504 29428 2588
rect 29506 2504 29536 2588
rect 29602 2504 29632 2672
rect 29674 2504 29704 2672
rect 29872 2572 29902 2700
rect 29969 2504 29999 2704
rect 30157 2520 30187 2648
rect 30252 2504 30282 2704
rect 25656 2180 25686 2308
rect 25740 2180 25770 2308
rect 25928 2230 25958 2314
rect 26021 2230 26051 2314
rect 26105 2230 26135 2314
rect 26225 2230 26255 2314
rect 26331 2230 26361 2314
rect 26439 2146 26469 2314
rect 26523 2146 26553 2314
rect 26660 2146 26690 2314
rect 26804 2230 26834 2314
rect 26888 2230 26918 2314
rect 27006 2230 27036 2314
rect 27114 2230 27144 2314
rect 27210 2146 27240 2314
rect 27282 2146 27312 2314
rect 27480 2118 27510 2246
rect 27577 2114 27607 2314
rect 27765 2170 27795 2298
rect 27860 2114 27890 2314
rect 28048 2180 28078 2308
rect 28132 2180 28162 2308
rect 28320 2230 28350 2314
rect 28413 2230 28443 2314
rect 28497 2230 28527 2314
rect 28617 2230 28647 2314
rect 28723 2230 28753 2314
rect 28831 2146 28861 2314
rect 28915 2146 28945 2314
rect 29052 2146 29082 2314
rect 29196 2230 29226 2314
rect 29280 2230 29310 2314
rect 29398 2230 29428 2314
rect 29506 2230 29536 2314
rect 29602 2146 29632 2314
rect 29674 2146 29704 2314
rect 29872 2118 29902 2246
rect 29969 2114 29999 2314
rect 30157 2170 30187 2298
rect 30252 2114 30282 2314
rect 8656 1184 8686 1342
rect 8744 1184 8774 1342
rect 8932 1142 8962 1342
rect 9016 1142 9046 1342
rect 9100 1142 9130 1342
rect 9184 1142 9214 1342
rect 9268 1142 9298 1342
rect 9484 1142 9514 1342
rect 9568 1142 9598 1342
rect 9652 1142 9682 1342
rect 9736 1142 9766 1342
rect 9820 1142 9850 1342
rect 9904 1142 9934 1342
rect 9988 1142 10018 1342
rect 10072 1142 10102 1342
rect 10156 1142 10186 1342
rect 10240 1142 10270 1342
rect 10324 1142 10354 1342
rect 10408 1142 10438 1342
rect 10492 1142 10522 1342
rect 10576 1142 10606 1342
rect 10660 1142 10690 1342
rect 10744 1142 10774 1342
rect 10828 1142 10858 1342
rect 10912 1142 10942 1342
rect 10996 1142 11026 1342
rect 11080 1142 11110 1342
rect 11164 1142 11194 1342
rect 11248 1142 11278 1342
rect 13040 1184 13070 1342
rect 13128 1184 13158 1342
rect 13316 1142 13346 1342
rect 13400 1142 13430 1342
rect 13484 1142 13514 1342
rect 13568 1142 13598 1342
rect 13652 1142 13682 1342
rect 13868 1142 13898 1342
rect 13952 1142 13982 1342
rect 14036 1142 14066 1342
rect 14120 1142 14150 1342
rect 14204 1142 14234 1342
rect 14288 1142 14318 1342
rect 14372 1142 14402 1342
rect 14456 1142 14486 1342
rect 14540 1142 14570 1342
rect 14624 1142 14654 1342
rect 14708 1142 14738 1342
rect 14792 1142 14822 1342
rect 14876 1142 14906 1342
rect 14960 1142 14990 1342
rect 15044 1142 15074 1342
rect 15128 1142 15158 1342
rect 15212 1142 15242 1342
rect 15296 1142 15326 1342
rect 15380 1142 15410 1342
rect 15464 1142 15494 1342
rect 15548 1142 15578 1342
rect 15632 1142 15662 1342
rect 8654 0 8684 200
rect 8763 77 8793 161
rect 8866 77 8896 161
rect 9080 77 9110 161
rect 9152 77 9182 161
rect 9248 77 9278 161
rect 10134 77 10164 161
rect 10230 77 10260 161
rect 10302 77 10332 161
rect 10516 77 10546 161
rect 10619 77 10649 161
rect 10728 0 10758 200
rect 11046 0 11076 200
rect 11155 77 11185 161
rect 11258 77 11288 161
rect 11472 77 11502 161
rect 11544 77 11574 161
rect 11640 77 11670 161
rect 12526 77 12556 161
rect 12622 77 12652 161
rect 12694 77 12724 161
rect 12908 77 12938 161
rect 13011 77 13041 161
rect 13120 0 13150 200
rect 13438 0 13468 200
rect 13547 77 13577 161
rect 13650 77 13680 161
rect 13864 77 13894 161
rect 13936 77 13966 161
rect 14032 77 14062 161
rect 14916 77 14946 161
rect 15012 77 15042 161
rect 15084 77 15114 161
rect 15298 77 15328 161
rect 15401 77 15431 161
rect 15510 0 15540 200
rect 15830 0 15860 200
rect 15939 77 15969 161
rect 16042 77 16072 161
rect 16256 77 16286 161
rect 16328 77 16358 161
rect 16424 77 16454 161
rect 17310 77 17340 161
rect 17406 77 17436 161
rect 17478 77 17508 161
rect 17692 77 17722 161
rect 17795 77 17825 161
rect 17904 0 17934 200
rect 18222 0 18252 200
rect 18331 77 18361 161
rect 18434 77 18464 161
rect 18648 77 18678 161
rect 18720 77 18750 161
rect 18816 77 18846 161
rect 19702 77 19732 161
rect 19798 77 19828 161
rect 19870 77 19900 161
rect 20084 77 20114 161
rect 20187 77 20217 161
rect 20296 0 20326 200
rect 20614 0 20644 200
rect 20723 77 20753 161
rect 20826 77 20856 161
rect 21040 77 21070 161
rect 21112 77 21142 161
rect 21208 77 21238 161
rect 22092 77 22122 161
rect 22188 77 22218 161
rect 22260 77 22290 161
rect 22474 77 22504 161
rect 22577 77 22607 161
rect 22686 0 22716 200
rect 23006 0 23036 200
rect 23115 77 23145 161
rect 23218 77 23248 161
rect 23432 77 23462 161
rect 23504 77 23534 161
rect 23600 77 23630 161
rect 24486 77 24516 161
rect 24582 77 24612 161
rect 24654 77 24684 161
rect 24868 77 24898 161
rect 24971 77 25001 161
rect 25080 0 25110 200
rect 8654 -622 8684 -494
rect 8738 -622 8768 -494
rect 8926 -572 8956 -488
rect 9018 -572 9048 -488
rect 9102 -572 9132 -488
rect 9222 -572 9252 -488
rect 9328 -572 9358 -488
rect 9436 -656 9466 -488
rect 9520 -656 9550 -488
rect 9657 -656 9687 -488
rect 9801 -572 9831 -488
rect 9885 -572 9915 -488
rect 9990 -572 10020 -488
rect 10111 -572 10141 -488
rect 10217 -656 10247 -488
rect 10289 -656 10319 -488
rect 10478 -684 10508 -556
rect 10575 -688 10605 -488
rect 10763 -632 10793 -504
rect 10858 -688 10888 -488
rect 11046 -622 11076 -494
rect 11130 -622 11160 -494
rect 11318 -572 11348 -488
rect 11410 -572 11440 -488
rect 11494 -572 11524 -488
rect 11614 -572 11644 -488
rect 11720 -572 11750 -488
rect 11828 -656 11858 -488
rect 11912 -656 11942 -488
rect 12049 -656 12079 -488
rect 12193 -572 12223 -488
rect 12277 -572 12307 -488
rect 12382 -572 12412 -488
rect 12503 -572 12533 -488
rect 12609 -656 12639 -488
rect 12681 -656 12711 -488
rect 12870 -684 12900 -556
rect 12967 -688 12997 -488
rect 13155 -632 13185 -504
rect 13250 -688 13280 -488
rect 13438 -622 13468 -494
rect 13522 -622 13552 -494
rect 13710 -572 13740 -488
rect 13802 -572 13832 -488
rect 13886 -572 13916 -488
rect 14006 -572 14036 -488
rect 14112 -572 14142 -488
rect 14220 -656 14250 -488
rect 14304 -656 14334 -488
rect 14441 -656 14471 -488
rect 14585 -572 14615 -488
rect 14669 -572 14699 -488
rect 14774 -572 14804 -488
rect 14895 -572 14925 -488
rect 15001 -656 15031 -488
rect 15073 -656 15103 -488
rect 15262 -684 15292 -556
rect 15359 -688 15389 -488
rect 15547 -632 15577 -504
rect 15642 -688 15672 -488
rect 15830 -622 15860 -494
rect 15914 -622 15944 -494
rect 16102 -572 16132 -488
rect 16194 -572 16224 -488
rect 16278 -572 16308 -488
rect 16398 -572 16428 -488
rect 16504 -572 16534 -488
rect 16612 -656 16642 -488
rect 16696 -656 16726 -488
rect 16833 -656 16863 -488
rect 16977 -572 17007 -488
rect 17061 -572 17091 -488
rect 17166 -572 17196 -488
rect 17287 -572 17317 -488
rect 17393 -656 17423 -488
rect 17465 -656 17495 -488
rect 17654 -684 17684 -556
rect 17751 -688 17781 -488
rect 17939 -632 17969 -504
rect 18034 -688 18064 -488
rect 18222 -622 18252 -494
rect 18306 -622 18336 -494
rect 18494 -572 18524 -488
rect 18586 -572 18616 -488
rect 18670 -572 18700 -488
rect 18790 -572 18820 -488
rect 18896 -572 18926 -488
rect 19004 -656 19034 -488
rect 19088 -656 19118 -488
rect 19225 -656 19255 -488
rect 19369 -572 19399 -488
rect 19453 -572 19483 -488
rect 19558 -572 19588 -488
rect 19679 -572 19709 -488
rect 19785 -656 19815 -488
rect 19857 -656 19887 -488
rect 20046 -684 20076 -556
rect 20143 -688 20173 -488
rect 20331 -632 20361 -504
rect 20426 -688 20456 -488
rect 20614 -622 20644 -494
rect 20698 -622 20728 -494
rect 20886 -572 20916 -488
rect 20978 -572 21008 -488
rect 21062 -572 21092 -488
rect 21182 -572 21212 -488
rect 21288 -572 21318 -488
rect 21396 -656 21426 -488
rect 21480 -656 21510 -488
rect 21617 -656 21647 -488
rect 21761 -572 21791 -488
rect 21845 -572 21875 -488
rect 21950 -572 21980 -488
rect 22071 -572 22101 -488
rect 22177 -656 22207 -488
rect 22249 -656 22279 -488
rect 22438 -684 22468 -556
rect 22535 -688 22565 -488
rect 22723 -632 22753 -504
rect 22818 -688 22848 -488
rect 23006 -622 23036 -494
rect 23090 -622 23120 -494
rect 23278 -572 23308 -488
rect 23370 -572 23400 -488
rect 23454 -572 23484 -488
rect 23574 -572 23604 -488
rect 23680 -572 23710 -488
rect 23788 -656 23818 -488
rect 23872 -656 23902 -488
rect 24009 -656 24039 -488
rect 24153 -572 24183 -488
rect 24237 -572 24267 -488
rect 24342 -572 24372 -488
rect 24463 -572 24493 -488
rect 24569 -656 24599 -488
rect 24641 -656 24671 -488
rect 24830 -684 24860 -556
rect 24927 -688 24957 -488
rect 25115 -632 25145 -504
rect 25210 -688 25240 -488
rect 8654 -1377 8684 -1177
rect 8749 -1321 8779 -1193
rect 8937 -1377 8967 -1177
rect 9034 -1373 9064 -1245
rect 9223 -1345 9253 -1177
rect 9295 -1345 9325 -1177
rect 9401 -1261 9431 -1177
rect 9522 -1261 9552 -1177
rect 9627 -1261 9657 -1177
rect 9711 -1261 9741 -1177
rect 9855 -1345 9885 -1177
rect 9992 -1345 10022 -1177
rect 10076 -1345 10106 -1177
rect 10184 -1261 10214 -1177
rect 10290 -1261 10320 -1177
rect 10410 -1261 10440 -1177
rect 10494 -1261 10524 -1177
rect 10586 -1261 10616 -1177
rect 10774 -1311 10804 -1183
rect 10858 -1311 10888 -1183
rect 11046 -1377 11076 -1177
rect 11141 -1321 11171 -1193
rect 11329 -1377 11359 -1177
rect 11426 -1373 11456 -1245
rect 11615 -1345 11645 -1177
rect 11687 -1345 11717 -1177
rect 11793 -1261 11823 -1177
rect 11914 -1261 11944 -1177
rect 12019 -1261 12049 -1177
rect 12103 -1261 12133 -1177
rect 12247 -1345 12277 -1177
rect 12384 -1345 12414 -1177
rect 12468 -1345 12498 -1177
rect 12576 -1261 12606 -1177
rect 12682 -1261 12712 -1177
rect 12802 -1261 12832 -1177
rect 12886 -1261 12916 -1177
rect 12978 -1261 13008 -1177
rect 13166 -1311 13196 -1183
rect 13250 -1311 13280 -1183
rect 13438 -1377 13468 -1177
rect 13533 -1321 13563 -1193
rect 13721 -1377 13751 -1177
rect 13818 -1373 13848 -1245
rect 14007 -1345 14037 -1177
rect 14079 -1345 14109 -1177
rect 14185 -1261 14215 -1177
rect 14306 -1261 14336 -1177
rect 14411 -1261 14441 -1177
rect 14495 -1261 14525 -1177
rect 14639 -1345 14669 -1177
rect 14776 -1345 14806 -1177
rect 14860 -1345 14890 -1177
rect 14968 -1261 14998 -1177
rect 15074 -1261 15104 -1177
rect 15194 -1261 15224 -1177
rect 15278 -1261 15308 -1177
rect 15370 -1261 15400 -1177
rect 15558 -1311 15588 -1183
rect 15642 -1311 15672 -1183
rect 15830 -1377 15860 -1177
rect 15925 -1321 15955 -1193
rect 16113 -1377 16143 -1177
rect 16210 -1373 16240 -1245
rect 16399 -1345 16429 -1177
rect 16471 -1345 16501 -1177
rect 16577 -1261 16607 -1177
rect 16698 -1261 16728 -1177
rect 16803 -1261 16833 -1177
rect 16887 -1261 16917 -1177
rect 17031 -1345 17061 -1177
rect 17168 -1345 17198 -1177
rect 17252 -1345 17282 -1177
rect 17360 -1261 17390 -1177
rect 17466 -1261 17496 -1177
rect 17586 -1261 17616 -1177
rect 17670 -1261 17700 -1177
rect 17762 -1261 17792 -1177
rect 17950 -1311 17980 -1183
rect 18034 -1311 18064 -1183
rect 18222 -1377 18252 -1177
rect 18317 -1321 18347 -1193
rect 18505 -1377 18535 -1177
rect 18602 -1373 18632 -1245
rect 18791 -1345 18821 -1177
rect 18863 -1345 18893 -1177
rect 18969 -1261 18999 -1177
rect 19090 -1261 19120 -1177
rect 19195 -1261 19225 -1177
rect 19279 -1261 19309 -1177
rect 19423 -1345 19453 -1177
rect 19560 -1345 19590 -1177
rect 19644 -1345 19674 -1177
rect 19752 -1261 19782 -1177
rect 19858 -1261 19888 -1177
rect 19978 -1261 20008 -1177
rect 20062 -1261 20092 -1177
rect 20154 -1261 20184 -1177
rect 20342 -1311 20372 -1183
rect 20426 -1311 20456 -1183
rect 20614 -1377 20644 -1177
rect 20709 -1321 20739 -1193
rect 20897 -1377 20927 -1177
rect 20994 -1373 21024 -1245
rect 21183 -1345 21213 -1177
rect 21255 -1345 21285 -1177
rect 21361 -1261 21391 -1177
rect 21482 -1261 21512 -1177
rect 21587 -1261 21617 -1177
rect 21671 -1261 21701 -1177
rect 21815 -1345 21845 -1177
rect 21952 -1345 21982 -1177
rect 22036 -1345 22066 -1177
rect 22144 -1261 22174 -1177
rect 22250 -1261 22280 -1177
rect 22370 -1261 22400 -1177
rect 22454 -1261 22484 -1177
rect 22546 -1261 22576 -1177
rect 22734 -1311 22764 -1183
rect 22818 -1311 22848 -1183
rect 23006 -1377 23036 -1177
rect 23101 -1321 23131 -1193
rect 23289 -1377 23319 -1177
rect 23386 -1373 23416 -1245
rect 23575 -1345 23605 -1177
rect 23647 -1345 23677 -1177
rect 23753 -1261 23783 -1177
rect 23874 -1261 23904 -1177
rect 23979 -1261 24009 -1177
rect 24063 -1261 24093 -1177
rect 24207 -1345 24237 -1177
rect 24344 -1345 24374 -1177
rect 24428 -1345 24458 -1177
rect 24536 -1261 24566 -1177
rect 24642 -1261 24672 -1177
rect 24762 -1261 24792 -1177
rect 24846 -1261 24876 -1177
rect 24938 -1261 24968 -1177
rect 25126 -1311 25156 -1183
rect 25210 -1311 25240 -1183
<< pmoshvt >>
rect 13862 13509 13892 13593
rect 20571 13509 20601 13593
rect 13862 13371 13892 13455
rect 20571 13371 20601 13455
rect 13862 13233 13892 13317
rect 20571 13233 20601 13317
rect 2974 13034 3004 13118
rect 13862 13095 13892 13179
rect 20571 13095 20601 13179
rect 2974 12896 3004 12980
rect 13862 12957 13892 13041
rect 2974 12758 3004 12842
rect 20571 12957 20601 13041
rect 13862 12819 13892 12903
rect 2974 12620 3004 12704
rect 20571 12819 20601 12903
rect 2974 12482 3004 12566
rect 19647 12508 19677 12592
rect 2974 12344 3004 12428
rect 26356 12508 26386 12592
rect 8759 12033 8789 12117
rect 8759 11895 8789 11979
rect 8851 11895 8881 11979
rect 8947 11895 8977 11979
rect 19647 12370 19677 12454
rect 19739 12370 19769 12454
rect 19835 12370 19865 12454
rect 26356 12370 26386 12454
rect 26448 12370 26478 12454
rect 26544 12370 26574 12454
rect 8759 8667 8789 8751
rect 8851 8667 8881 8751
rect 8947 8667 8977 8751
rect 8759 8529 8789 8613
rect 13314 8655 13344 8739
rect 13410 8655 13440 8739
rect 13502 8655 13532 8739
rect 20023 8655 20053 8739
rect 20119 8655 20149 8739
rect 20211 8655 20241 8739
rect 13502 8517 13532 8601
rect 20211 8517 20241 8601
rect 2974 8218 3004 8302
rect 2974 8080 3004 8164
rect 2974 7942 3004 8026
rect 2974 7804 3004 7888
rect 19287 8206 19317 8290
rect 25996 8206 26026 8290
rect 19287 8068 19317 8152
rect 25996 8068 26026 8152
rect 2974 7666 3004 7750
rect 2974 7528 3004 7612
rect 19287 7930 19317 8014
rect 25996 7930 26026 8014
rect 19287 7792 19317 7876
rect 25996 7792 26026 7876
rect 19287 7654 19317 7738
rect 25996 7654 26026 7738
rect 19287 7516 19317 7600
rect 25996 7516 26026 7600
rect 24587 7212 24617 7296
rect 24587 7074 24617 7158
rect 24587 6936 24617 7020
rect 24587 6798 24617 6882
rect 24587 6660 24617 6744
rect 24587 6522 24617 6606
rect 30372 6211 30402 6295
rect 30372 6073 30402 6157
rect 30464 6073 30494 6157
rect 30560 6073 30590 6157
<< ndiff >>
rect 13342 12614 13394 12626
rect 13342 12580 13350 12614
rect 13384 12580 13394 12614
rect 13342 12546 13394 12580
rect 13342 12512 13350 12546
rect 13384 12512 13394 12546
rect 13342 12496 13394 12512
rect 13424 12614 13476 12626
rect 13424 12580 13434 12614
rect 13468 12580 13476 12614
rect 13424 12546 13476 12580
rect 13424 12512 13434 12546
rect 13468 12512 13476 12546
rect 13424 12496 13476 12512
rect 13532 12614 13584 12626
rect 13532 12580 13540 12614
rect 13574 12580 13584 12614
rect 13532 12546 13584 12580
rect 13532 12512 13540 12546
rect 13574 12512 13584 12546
rect 13532 12496 13584 12512
rect 13614 12614 13666 12626
rect 13614 12580 13624 12614
rect 13658 12580 13666 12614
rect 20051 12614 20103 12626
rect 13614 12546 13666 12580
rect 13614 12512 13624 12546
rect 13658 12512 13666 12546
rect 13614 12496 13666 12512
rect 20051 12580 20059 12614
rect 20093 12580 20103 12614
rect 20051 12546 20103 12580
rect 20051 12512 20059 12546
rect 20093 12512 20103 12546
rect 20051 12496 20103 12512
rect 20133 12614 20185 12626
rect 20133 12580 20143 12614
rect 20177 12580 20185 12614
rect 20133 12546 20185 12580
rect 20133 12512 20143 12546
rect 20177 12512 20185 12546
rect 20133 12496 20185 12512
rect 20241 12614 20293 12626
rect 20241 12580 20249 12614
rect 20283 12580 20293 12614
rect 20241 12546 20293 12580
rect 20241 12512 20249 12546
rect 20283 12512 20293 12546
rect 20241 12496 20293 12512
rect 20323 12614 20375 12626
rect 20323 12580 20333 12614
rect 20367 12580 20375 12614
rect 20323 12546 20375 12580
rect 20323 12512 20333 12546
rect 20367 12512 20375 12546
rect 20323 12496 20375 12512
rect 10909 12364 10961 12402
rect 10909 12330 10917 12364
rect 10951 12330 10961 12364
rect 10909 12318 10961 12330
rect 10991 12390 11045 12402
rect 10991 12356 11001 12390
rect 11035 12356 11045 12390
rect 10991 12318 11045 12356
rect 11075 12364 11127 12402
rect 11075 12330 11085 12364
rect 11119 12330 11127 12364
rect 11075 12318 11127 12330
rect 11181 12390 11233 12402
rect 11181 12356 11189 12390
rect 11223 12356 11233 12390
rect 11181 12318 11233 12356
rect 11263 12372 11328 12402
rect 11263 12338 11273 12372
rect 11307 12338 11328 12372
rect 11263 12330 11328 12338
rect 11358 12390 11434 12402
rect 11358 12356 11379 12390
rect 11413 12356 11434 12390
rect 11358 12330 11434 12356
rect 11464 12330 11530 12402
rect 11263 12318 11313 12330
rect 11479 12318 11530 12330
rect 11560 12394 11640 12402
rect 11560 12360 11596 12394
rect 11630 12360 11640 12394
rect 11560 12318 11640 12360
rect 11670 12374 11740 12402
rect 11670 12340 11680 12374
rect 11714 12340 11740 12374
rect 11670 12318 11740 12340
rect 2454 12139 2506 12151
rect 2454 12105 2462 12139
rect 2496 12105 2506 12139
rect 2454 12071 2506 12105
rect 2454 12037 2462 12071
rect 2496 12037 2506 12071
rect 2454 12021 2506 12037
rect 2536 12139 2588 12151
rect 2536 12105 2546 12139
rect 2580 12105 2588 12139
rect 2536 12071 2588 12105
rect 2536 12037 2546 12071
rect 2580 12037 2588 12071
rect 2536 12021 2588 12037
rect 2644 12139 2696 12151
rect 2644 12105 2652 12139
rect 2686 12105 2696 12139
rect 2644 12071 2696 12105
rect 2644 12037 2652 12071
rect 2686 12037 2696 12071
rect 2644 12021 2696 12037
rect 2726 12139 2778 12151
rect 2726 12105 2736 12139
rect 2770 12105 2778 12139
rect 2726 12071 2778 12105
rect 2726 12037 2736 12071
rect 2770 12037 2778 12071
rect 2726 12021 2778 12037
rect 11690 12274 11740 12318
rect 11770 12330 11824 12402
rect 11770 12296 11780 12330
rect 11814 12296 11824 12330
rect 11770 12274 11824 12296
rect 11854 12356 11906 12402
rect 11854 12322 11864 12356
rect 11898 12322 11906 12356
rect 11854 12274 11906 12322
rect 11960 12390 12012 12402
rect 11960 12356 11968 12390
rect 12002 12356 12012 12390
rect 11960 12274 12012 12356
rect 12042 12330 12107 12402
rect 12137 12390 12216 12402
rect 12137 12356 12162 12390
rect 12196 12356 12216 12390
rect 12137 12330 12216 12356
rect 12246 12330 12311 12402
rect 12042 12274 12092 12330
rect 12261 12318 12311 12330
rect 12341 12394 12397 12402
rect 12341 12360 12353 12394
rect 12387 12360 12397 12394
rect 12341 12318 12397 12360
rect 12427 12374 12515 12402
rect 12427 12340 12455 12374
rect 12489 12340 12515 12374
rect 12427 12318 12515 12340
rect 12465 12274 12515 12318
rect 12545 12330 12599 12402
rect 12545 12296 12555 12330
rect 12589 12296 12599 12330
rect 12545 12274 12599 12296
rect 12629 12382 12681 12402
rect 12629 12348 12639 12382
rect 12673 12348 12681 12382
rect 12629 12274 12681 12348
rect 12735 12380 12787 12402
rect 12735 12346 12743 12380
rect 12777 12346 12787 12380
rect 12735 12318 12787 12346
rect 12817 12390 12882 12402
rect 12817 12356 12838 12390
rect 12872 12356 12882 12390
rect 12817 12318 12882 12356
rect 12832 12272 12882 12318
rect 12912 12356 12964 12402
rect 12912 12322 12922 12356
rect 12956 12322 12964 12356
rect 12912 12272 12964 12322
rect 13018 12364 13070 12402
rect 13018 12330 13026 12364
rect 13060 12330 13070 12364
rect 13018 12318 13070 12330
rect 13100 12390 13165 12402
rect 13100 12356 13121 12390
rect 13155 12356 13165 12390
rect 13100 12318 13165 12356
rect 13115 12272 13165 12318
rect 13195 12354 13247 12402
rect 13195 12320 13205 12354
rect 13239 12320 13247 12354
rect 13195 12272 13247 12320
rect 14799 12238 14857 12250
rect 14799 12178 14811 12238
rect 14845 12178 14857 12238
rect 14799 12166 14857 12178
rect 14887 12238 14945 12250
rect 14887 12178 14901 12238
rect 14935 12178 14945 12238
rect 14887 12166 14945 12178
rect 15531 12238 15589 12250
rect 15531 12178 15543 12238
rect 15577 12178 15589 12238
rect 15531 12166 15589 12178
rect 15619 12238 15711 12250
rect 15619 12178 15650 12238
rect 15684 12178 15711 12238
rect 15619 12166 15711 12178
rect 15741 12238 15799 12250
rect 15741 12178 15753 12238
rect 15787 12178 15799 12238
rect 15741 12166 15799 12178
rect 16743 12238 16801 12250
rect 16743 12178 16755 12238
rect 16789 12178 16801 12238
rect 16743 12166 16801 12178
rect 16831 12238 16923 12250
rect 16831 12178 16861 12238
rect 16895 12178 16923 12238
rect 16831 12166 16923 12178
rect 16953 12238 17011 12250
rect 16953 12178 16965 12238
rect 16999 12178 17011 12238
rect 16953 12166 17011 12178
rect 18081 12238 18139 12250
rect 18081 12178 18093 12238
rect 18127 12178 18139 12238
rect 18081 12166 18139 12178
rect 18169 12238 18261 12250
rect 18169 12178 18201 12238
rect 18235 12178 18261 12238
rect 18169 12166 18261 12178
rect 18291 12238 18349 12250
rect 18291 12178 18303 12238
rect 18337 12178 18349 12238
rect 18291 12166 18349 12178
rect 18936 12238 18995 12250
rect 18936 12178 18948 12238
rect 18982 12178 18995 12238
rect 18936 12166 18995 12178
rect 19025 12238 19083 12250
rect 19025 12178 19037 12238
rect 19071 12178 19083 12238
rect 19025 12166 19083 12178
rect 19589 12239 19647 12251
rect 19589 12179 19601 12239
rect 19635 12179 19647 12239
rect 19589 12167 19647 12179
rect 19677 12239 19739 12251
rect 19677 12179 19689 12239
rect 19723 12179 19739 12239
rect 19677 12167 19739 12179
rect 19769 12239 19835 12251
rect 19769 12179 19785 12239
rect 19819 12179 19835 12239
rect 19769 12167 19835 12179
rect 19865 12239 19927 12251
rect 19865 12179 19881 12239
rect 19915 12179 19927 12239
rect 19865 12167 19927 12179
rect 21508 12238 21566 12250
rect 21508 12178 21520 12238
rect 21554 12178 21566 12238
rect 21508 12166 21566 12178
rect 21596 12238 21654 12250
rect 21596 12178 21610 12238
rect 21644 12178 21654 12238
rect 21596 12166 21654 12178
rect 22240 12238 22298 12250
rect 22240 12178 22252 12238
rect 22286 12178 22298 12238
rect 22240 12166 22298 12178
rect 22328 12238 22420 12250
rect 22328 12178 22359 12238
rect 22393 12178 22420 12238
rect 22328 12166 22420 12178
rect 22450 12238 22508 12250
rect 22450 12178 22462 12238
rect 22496 12178 22508 12238
rect 22450 12166 22508 12178
rect 23452 12238 23510 12250
rect 23452 12178 23464 12238
rect 23498 12178 23510 12238
rect 23452 12166 23510 12178
rect 23540 12238 23632 12250
rect 23540 12178 23570 12238
rect 23604 12178 23632 12238
rect 23540 12166 23632 12178
rect 23662 12238 23720 12250
rect 23662 12178 23674 12238
rect 23708 12178 23720 12238
rect 23662 12166 23720 12178
rect 24790 12238 24848 12250
rect 24790 12178 24802 12238
rect 24836 12178 24848 12238
rect 24790 12166 24848 12178
rect 24878 12238 24970 12250
rect 24878 12178 24910 12238
rect 24944 12178 24970 12238
rect 24878 12166 24970 12178
rect 25000 12238 25058 12250
rect 25000 12178 25012 12238
rect 25046 12178 25058 12238
rect 25000 12166 25058 12178
rect 25645 12238 25704 12250
rect 25645 12178 25657 12238
rect 25691 12178 25704 12238
rect 25645 12166 25704 12178
rect 25734 12238 25792 12250
rect 25734 12178 25746 12238
rect 25780 12178 25792 12238
rect 25734 12166 25792 12178
rect 26298 12239 26356 12251
rect 26298 12179 26310 12239
rect 26344 12179 26356 12239
rect 26298 12167 26356 12179
rect 26386 12239 26448 12251
rect 26386 12179 26398 12239
rect 26432 12179 26448 12239
rect 26386 12167 26448 12179
rect 26478 12239 26544 12251
rect 26478 12179 26494 12239
rect 26528 12179 26544 12239
rect 26478 12167 26544 12179
rect 26574 12239 26636 12251
rect 26574 12179 26590 12239
rect 26624 12179 26636 12239
rect 26574 12167 26636 12179
rect 19589 12101 19647 12113
rect 13779 12054 13837 12066
rect 13779 11994 13791 12054
rect 13825 11994 13837 12054
rect 13779 11982 13837 11994
rect 13867 11982 13909 12066
rect 13939 12054 13997 12066
rect 13939 11994 13951 12054
rect 13985 11994 13997 12054
rect 19589 12041 19601 12101
rect 19635 12041 19647 12101
rect 19589 12029 19647 12041
rect 19677 12101 19735 12113
rect 19677 12041 19689 12101
rect 19723 12041 19735 12101
rect 26298 12101 26356 12113
rect 19677 12029 19735 12041
rect 20488 12054 20546 12066
rect 13939 11982 13997 11994
rect 20488 11994 20500 12054
rect 20534 11994 20546 12054
rect 20488 11982 20546 11994
rect 20576 11982 20618 12066
rect 20648 12054 20706 12066
rect 20648 11994 20660 12054
rect 20694 11994 20706 12054
rect 26298 12041 26310 12101
rect 26344 12041 26356 12101
rect 26298 12029 26356 12041
rect 26386 12101 26444 12113
rect 26386 12041 26398 12101
rect 26432 12041 26444 12101
rect 26386 12029 26444 12041
rect 20648 11982 20706 11994
rect 13779 11916 13837 11928
rect 13779 11856 13791 11916
rect 13825 11856 13837 11916
rect 13779 11844 13837 11856
rect 13867 11844 13909 11928
rect 13939 11916 13997 11928
rect 13939 11856 13951 11916
rect 13985 11856 13997 11916
rect 13939 11844 13997 11856
rect 20488 11916 20546 11928
rect 20488 11856 20500 11916
rect 20534 11856 20546 11916
rect 20488 11844 20546 11856
rect 20576 11844 20618 11928
rect 20648 11916 20706 11928
rect 20648 11856 20660 11916
rect 20694 11856 20706 11916
rect 20648 11844 20706 11856
rect 3911 11763 3969 11775
rect 3911 11703 3923 11763
rect 3957 11703 3969 11763
rect 3911 11691 3969 11703
rect 3999 11763 4057 11775
rect 3999 11703 4013 11763
rect 4047 11703 4057 11763
rect 3999 11691 4057 11703
rect 4643 11763 4701 11775
rect 4643 11703 4655 11763
rect 4689 11703 4701 11763
rect 4643 11691 4701 11703
rect 4731 11763 4823 11775
rect 4731 11703 4762 11763
rect 4796 11703 4823 11763
rect 4731 11691 4823 11703
rect 4853 11763 4911 11775
rect 4853 11703 4865 11763
rect 4899 11703 4911 11763
rect 4853 11691 4911 11703
rect 5855 11763 5913 11775
rect 5855 11703 5867 11763
rect 5901 11703 5913 11763
rect 5855 11691 5913 11703
rect 5943 11763 6035 11775
rect 5943 11703 5973 11763
rect 6007 11703 6035 11763
rect 5943 11691 6035 11703
rect 6065 11763 6123 11775
rect 6065 11703 6077 11763
rect 6111 11703 6123 11763
rect 6065 11691 6123 11703
rect 7193 11763 7251 11775
rect 7193 11703 7205 11763
rect 7239 11703 7251 11763
rect 7193 11691 7251 11703
rect 7281 11763 7373 11775
rect 7281 11703 7313 11763
rect 7347 11703 7373 11763
rect 7281 11691 7373 11703
rect 7403 11763 7461 11775
rect 7403 11703 7415 11763
rect 7449 11703 7461 11763
rect 7403 11691 7461 11703
rect 8048 11763 8107 11775
rect 8048 11703 8060 11763
rect 8094 11703 8107 11763
rect 8048 11691 8107 11703
rect 8137 11763 8195 11775
rect 8137 11703 8149 11763
rect 8183 11703 8195 11763
rect 8137 11691 8195 11703
rect 8701 11764 8759 11776
rect 8701 11704 8713 11764
rect 8747 11704 8759 11764
rect 8701 11692 8759 11704
rect 8789 11764 8851 11776
rect 8789 11704 8801 11764
rect 8835 11704 8851 11764
rect 8789 11692 8851 11704
rect 8881 11764 8947 11776
rect 8881 11704 8897 11764
rect 8931 11704 8947 11764
rect 8881 11692 8947 11704
rect 8977 11764 9039 11776
rect 8977 11704 8993 11764
rect 9027 11704 9039 11764
rect 8977 11692 9039 11704
rect 9129 11762 9181 11774
rect 9129 11728 9137 11762
rect 9171 11728 9181 11762
rect 9129 11694 9181 11728
rect 9129 11660 9137 11694
rect 9171 11660 9181 11694
rect 9129 11644 9181 11660
rect 9211 11762 9263 11774
rect 13779 11778 13837 11790
rect 9211 11728 9221 11762
rect 9255 11728 9263 11762
rect 9211 11694 9263 11728
rect 9211 11660 9221 11694
rect 9255 11660 9263 11694
rect 9211 11644 9263 11660
rect 8701 11626 8759 11638
rect 2891 11579 2949 11591
rect 2891 11519 2903 11579
rect 2937 11519 2949 11579
rect 2891 11507 2949 11519
rect 2979 11507 3021 11591
rect 3051 11579 3109 11591
rect 3051 11519 3063 11579
rect 3097 11519 3109 11579
rect 8701 11566 8713 11626
rect 8747 11566 8759 11626
rect 8701 11554 8759 11566
rect 8789 11626 8847 11638
rect 8789 11566 8801 11626
rect 8835 11566 8847 11626
rect 8789 11554 8847 11566
rect 13779 11718 13791 11778
rect 13825 11718 13837 11778
rect 13779 11706 13837 11718
rect 13867 11706 13909 11790
rect 13939 11778 13997 11790
rect 13939 11718 13951 11778
rect 13985 11718 13997 11778
rect 13939 11706 13997 11718
rect 20488 11778 20546 11790
rect 20488 11718 20500 11778
rect 20534 11718 20546 11778
rect 20488 11706 20546 11718
rect 20576 11706 20618 11790
rect 20648 11778 20706 11790
rect 20648 11718 20660 11778
rect 20694 11718 20706 11778
rect 20648 11706 20706 11718
rect 13779 11640 13837 11652
rect 3051 11507 3109 11519
rect 13779 11580 13791 11640
rect 13825 11580 13837 11640
rect 13779 11568 13837 11580
rect 13867 11568 13909 11652
rect 13939 11640 13997 11652
rect 13939 11580 13951 11640
rect 13985 11580 13997 11640
rect 13939 11568 13997 11580
rect 20488 11640 20546 11652
rect 20488 11580 20500 11640
rect 20534 11580 20546 11640
rect 20488 11568 20546 11580
rect 20576 11568 20618 11652
rect 20648 11640 20706 11652
rect 20648 11580 20660 11640
rect 20694 11580 20706 11640
rect 20648 11568 20706 11580
rect 2891 11441 2949 11453
rect 2891 11381 2903 11441
rect 2937 11381 2949 11441
rect 2891 11369 2949 11381
rect 2979 11369 3021 11453
rect 3051 11441 3109 11453
rect 13779 11502 13837 11514
rect 13779 11442 13791 11502
rect 13825 11442 13837 11502
rect 3051 11381 3063 11441
rect 3097 11381 3109 11441
rect 3051 11369 3109 11381
rect 10950 11430 11002 11442
rect 10950 11396 10958 11430
rect 10992 11396 11002 11430
rect 10950 11362 11002 11396
rect 10950 11328 10958 11362
rect 10992 11328 11002 11362
rect 2891 11303 2949 11315
rect 2891 11243 2903 11303
rect 2937 11243 2949 11303
rect 2891 11231 2949 11243
rect 2979 11231 3021 11315
rect 3051 11303 3109 11315
rect 10950 11312 11002 11328
rect 11032 11430 11084 11442
rect 11032 11396 11042 11430
rect 11076 11396 11084 11430
rect 11032 11362 11084 11396
rect 11032 11328 11042 11362
rect 11076 11328 11084 11362
rect 11032 11312 11084 11328
rect 11226 11430 11278 11442
rect 11226 11396 11234 11430
rect 11268 11396 11278 11430
rect 11226 11362 11278 11396
rect 11226 11328 11234 11362
rect 11268 11328 11278 11362
rect 11226 11312 11278 11328
rect 11308 11430 11360 11442
rect 13779 11430 13837 11442
rect 13867 11430 13909 11514
rect 13939 11502 13997 11514
rect 13939 11442 13951 11502
rect 13985 11442 13997 11502
rect 13939 11430 13997 11442
rect 20488 11502 20546 11514
rect 20488 11442 20500 11502
rect 20534 11442 20546 11502
rect 20488 11430 20546 11442
rect 20576 11430 20618 11514
rect 20648 11502 20706 11514
rect 20648 11442 20660 11502
rect 20694 11442 20706 11502
rect 20648 11430 20706 11442
rect 11308 11396 11318 11430
rect 11352 11396 11360 11430
rect 11308 11362 11360 11396
rect 11308 11328 11318 11362
rect 11352 11328 11360 11362
rect 11308 11312 11360 11328
rect 13779 11364 13837 11376
rect 3051 11243 3063 11303
rect 3097 11243 3109 11303
rect 13779 11304 13791 11364
rect 13825 11304 13837 11364
rect 13779 11292 13837 11304
rect 13867 11292 13909 11376
rect 13939 11364 13997 11376
rect 13939 11304 13951 11364
rect 13985 11304 13997 11364
rect 13939 11292 13997 11304
rect 20488 11364 20546 11376
rect 20488 11304 20500 11364
rect 20534 11304 20546 11364
rect 20488 11292 20546 11304
rect 20576 11292 20618 11376
rect 20648 11364 20706 11376
rect 20648 11304 20660 11364
rect 20694 11304 20706 11364
rect 20648 11292 20706 11304
rect 3051 11231 3109 11243
rect 13779 11226 13837 11238
rect 2891 11165 2949 11177
rect 2891 11105 2903 11165
rect 2937 11105 2949 11165
rect 2891 11093 2949 11105
rect 2979 11093 3021 11177
rect 3051 11165 3109 11177
rect 3051 11105 3063 11165
rect 3097 11105 3109 11165
rect 13779 11166 13791 11226
rect 13825 11166 13837 11226
rect 13779 11154 13837 11166
rect 13867 11154 13909 11238
rect 13939 11226 13997 11238
rect 13939 11166 13951 11226
rect 13985 11166 13997 11226
rect 13939 11154 13997 11166
rect 3051 11093 3109 11105
rect 20488 11226 20546 11238
rect 20488 11166 20500 11226
rect 20534 11166 20546 11226
rect 20488 11154 20546 11166
rect 20576 11154 20618 11238
rect 20648 11226 20706 11238
rect 20648 11166 20660 11226
rect 20694 11166 20706 11226
rect 20648 11154 20706 11166
rect 13779 11088 13837 11100
rect 2891 11027 2949 11039
rect 2891 10967 2903 11027
rect 2937 10967 2949 11027
rect 2891 10955 2949 10967
rect 2979 10955 3021 11039
rect 3051 11027 3109 11039
rect 3051 10967 3063 11027
rect 3097 10967 3109 11027
rect 13779 11028 13791 11088
rect 13825 11028 13837 11088
rect 13779 11016 13837 11028
rect 13867 11016 13909 11100
rect 13939 11088 13997 11100
rect 13939 11028 13951 11088
rect 13985 11028 13997 11088
rect 20488 11088 20546 11100
rect 13939 11016 13997 11028
rect 20488 11028 20500 11088
rect 20534 11028 20546 11088
rect 20488 11016 20546 11028
rect 20576 11016 20618 11100
rect 20648 11088 20706 11100
rect 20648 11028 20660 11088
rect 20694 11028 20706 11088
rect 20648 11016 20706 11028
rect 3051 10955 3109 10967
rect 2891 10889 2949 10901
rect 2891 10829 2903 10889
rect 2937 10829 2949 10889
rect 2891 10817 2949 10829
rect 2979 10817 3021 10901
rect 3051 10889 3109 10901
rect 3051 10829 3063 10889
rect 3097 10829 3109 10889
rect 3051 10817 3109 10829
rect 2891 10751 2949 10763
rect 2891 10691 2903 10751
rect 2937 10691 2949 10751
rect 2891 10679 2949 10691
rect 2979 10679 3021 10763
rect 3051 10751 3109 10763
rect 3051 10691 3063 10751
rect 3097 10691 3109 10751
rect 3051 10679 3109 10691
rect 2891 10613 2949 10625
rect 2891 10553 2903 10613
rect 2937 10553 2949 10613
rect 2891 10541 2949 10553
rect 2979 10541 3021 10625
rect 3051 10613 3109 10625
rect 3051 10553 3063 10613
rect 3097 10553 3109 10613
rect 3051 10541 3109 10553
rect 2891 10093 2949 10105
rect 2891 10033 2903 10093
rect 2937 10033 2949 10093
rect 2891 10021 2949 10033
rect 2979 10021 3021 10105
rect 3051 10093 3109 10105
rect 3051 10033 3063 10093
rect 3097 10033 3109 10093
rect 19182 10081 19240 10093
rect 3051 10021 3109 10033
rect 19182 10021 19194 10081
rect 19228 10021 19240 10081
rect 19182 10009 19240 10021
rect 19270 10009 19312 10093
rect 19342 10081 19400 10093
rect 19342 10021 19354 10081
rect 19388 10021 19400 10081
rect 25891 10081 25949 10093
rect 19342 10009 19400 10021
rect 25891 10021 25903 10081
rect 25937 10021 25949 10081
rect 25891 10009 25949 10021
rect 25979 10009 26021 10093
rect 26051 10081 26109 10093
rect 26051 10021 26063 10081
rect 26097 10021 26109 10081
rect 26051 10009 26109 10021
rect 2891 9955 2949 9967
rect 2891 9895 2903 9955
rect 2937 9895 2949 9955
rect 2891 9883 2949 9895
rect 2979 9883 3021 9967
rect 3051 9955 3109 9967
rect 3051 9895 3063 9955
rect 3097 9895 3109 9955
rect 3051 9883 3109 9895
rect 19182 9943 19240 9955
rect 19182 9883 19194 9943
rect 19228 9883 19240 9943
rect 19182 9871 19240 9883
rect 19270 9871 19312 9955
rect 19342 9943 19400 9955
rect 19342 9883 19354 9943
rect 19388 9883 19400 9943
rect 19342 9871 19400 9883
rect 2891 9817 2949 9829
rect 2891 9757 2903 9817
rect 2937 9757 2949 9817
rect 2891 9745 2949 9757
rect 2979 9745 3021 9829
rect 3051 9817 3109 9829
rect 25891 9943 25949 9955
rect 25891 9883 25903 9943
rect 25937 9883 25949 9943
rect 25891 9871 25949 9883
rect 25979 9871 26021 9955
rect 26051 9943 26109 9955
rect 26051 9883 26063 9943
rect 26097 9883 26109 9943
rect 26051 9871 26109 9883
rect 3051 9757 3063 9817
rect 3097 9757 3109 9817
rect 3051 9745 3109 9757
rect 19182 9805 19240 9817
rect 19182 9745 19194 9805
rect 19228 9745 19240 9805
rect 19182 9733 19240 9745
rect 19270 9733 19312 9817
rect 19342 9805 19400 9817
rect 19342 9745 19354 9805
rect 19388 9745 19400 9805
rect 19342 9733 19400 9745
rect 25891 9805 25949 9817
rect 25891 9745 25903 9805
rect 25937 9745 25949 9805
rect 25891 9733 25949 9745
rect 25979 9733 26021 9817
rect 26051 9805 26109 9817
rect 26051 9745 26063 9805
rect 26097 9745 26109 9805
rect 26051 9733 26109 9745
rect 2891 9679 2949 9691
rect 2891 9619 2903 9679
rect 2937 9619 2949 9679
rect 2891 9607 2949 9619
rect 2979 9607 3021 9691
rect 3051 9679 3109 9691
rect 3051 9619 3063 9679
rect 3097 9619 3109 9679
rect 3051 9607 3109 9619
rect 19182 9667 19240 9679
rect 19182 9607 19194 9667
rect 19228 9607 19240 9667
rect 19182 9595 19240 9607
rect 19270 9595 19312 9679
rect 19342 9667 19400 9679
rect 19342 9607 19354 9667
rect 19388 9607 19400 9667
rect 19342 9595 19400 9607
rect 25891 9667 25949 9679
rect 25891 9607 25903 9667
rect 25937 9607 25949 9667
rect 25891 9595 25949 9607
rect 25979 9595 26021 9679
rect 26051 9667 26109 9679
rect 26051 9607 26063 9667
rect 26097 9607 26109 9667
rect 26051 9595 26109 9607
rect 2891 9541 2949 9553
rect 2891 9481 2903 9541
rect 2937 9481 2949 9541
rect 2891 9469 2949 9481
rect 2979 9469 3021 9553
rect 3051 9541 3109 9553
rect 3051 9481 3063 9541
rect 3097 9481 3109 9541
rect 3051 9469 3109 9481
rect 19182 9529 19240 9541
rect 19182 9469 19194 9529
rect 19228 9469 19240 9529
rect 19182 9457 19240 9469
rect 19270 9457 19312 9541
rect 19342 9529 19400 9541
rect 19342 9469 19354 9529
rect 19388 9469 19400 9529
rect 19342 9457 19400 9469
rect 25891 9529 25949 9541
rect 25891 9469 25903 9529
rect 25937 9469 25949 9529
rect 25891 9457 25949 9469
rect 25979 9457 26021 9541
rect 26051 9529 26109 9541
rect 26051 9469 26063 9529
rect 26097 9469 26109 9529
rect 26051 9457 26109 9469
rect 2891 9403 2949 9415
rect 2891 9343 2903 9403
rect 2937 9343 2949 9403
rect 2891 9331 2949 9343
rect 2979 9331 3021 9415
rect 3051 9403 3109 9415
rect 3051 9343 3063 9403
rect 3097 9343 3109 9403
rect 3051 9331 3109 9343
rect 19182 9391 19240 9403
rect 19182 9331 19194 9391
rect 19228 9331 19240 9391
rect 19182 9319 19240 9331
rect 19270 9319 19312 9403
rect 19342 9391 19400 9403
rect 19342 9331 19354 9391
rect 19388 9331 19400 9391
rect 19342 9319 19400 9331
rect 25891 9391 25949 9403
rect 25891 9331 25903 9391
rect 25937 9331 25949 9391
rect 25891 9319 25949 9331
rect 25979 9319 26021 9403
rect 26051 9391 26109 9403
rect 26051 9331 26063 9391
rect 26097 9331 26109 9391
rect 26051 9319 26109 9331
rect 2891 9265 2949 9277
rect 2891 9205 2903 9265
rect 2937 9205 2949 9265
rect 2891 9193 2949 9205
rect 2979 9193 3021 9277
rect 3051 9265 3109 9277
rect 3051 9205 3063 9265
rect 3097 9205 3109 9265
rect 3051 9193 3109 9205
rect 19182 9253 19240 9265
rect 19182 9193 19194 9253
rect 19228 9193 19240 9253
rect 19182 9181 19240 9193
rect 19270 9181 19312 9265
rect 19342 9253 19400 9265
rect 19342 9193 19354 9253
rect 19388 9193 19400 9253
rect 19342 9181 19400 9193
rect 25891 9253 25949 9265
rect 25891 9193 25903 9253
rect 25937 9193 25949 9253
rect 25891 9181 25949 9193
rect 25979 9181 26021 9265
rect 26051 9253 26109 9265
rect 26051 9193 26063 9253
rect 26097 9193 26109 9253
rect 26051 9181 26109 9193
rect 2891 9127 2949 9139
rect 2891 9067 2903 9127
rect 2937 9067 2949 9127
rect 2891 9055 2949 9067
rect 2979 9055 3021 9139
rect 3051 9127 3109 9139
rect 3051 9067 3063 9127
rect 3097 9067 3109 9127
rect 19182 9115 19240 9127
rect 3051 9055 3109 9067
rect 8701 9080 8759 9092
rect 8701 9020 8713 9080
rect 8747 9020 8759 9080
rect 8701 9008 8759 9020
rect 8789 9080 8847 9092
rect 8789 9020 8801 9080
rect 8835 9020 8847 9080
rect 13444 9068 13502 9080
rect 8789 9008 8847 9020
rect 3911 8943 3969 8955
rect 3911 8883 3923 8943
rect 3957 8883 3969 8943
rect 3911 8871 3969 8883
rect 3999 8943 4057 8955
rect 3999 8883 4013 8943
rect 4047 8883 4057 8943
rect 3999 8871 4057 8883
rect 4643 8943 4701 8955
rect 4643 8883 4655 8943
rect 4689 8883 4701 8943
rect 4643 8871 4701 8883
rect 4731 8943 4823 8955
rect 4731 8883 4762 8943
rect 4796 8883 4823 8943
rect 4731 8871 4823 8883
rect 4853 8943 4911 8955
rect 4853 8883 4865 8943
rect 4899 8883 4911 8943
rect 4853 8871 4911 8883
rect 5855 8943 5913 8955
rect 5855 8883 5867 8943
rect 5901 8883 5913 8943
rect 5855 8871 5913 8883
rect 5943 8943 6035 8955
rect 5943 8883 5973 8943
rect 6007 8883 6035 8943
rect 5943 8871 6035 8883
rect 6065 8943 6123 8955
rect 6065 8883 6077 8943
rect 6111 8883 6123 8943
rect 6065 8871 6123 8883
rect 7193 8943 7251 8955
rect 7193 8883 7205 8943
rect 7239 8883 7251 8943
rect 7193 8871 7251 8883
rect 7281 8943 7373 8955
rect 7281 8883 7313 8943
rect 7347 8883 7373 8943
rect 7281 8871 7373 8883
rect 7403 8943 7461 8955
rect 7403 8883 7415 8943
rect 7449 8883 7461 8943
rect 7403 8871 7461 8883
rect 8048 8943 8107 8955
rect 8048 8883 8060 8943
rect 8094 8883 8107 8943
rect 8048 8871 8107 8883
rect 8137 8943 8195 8955
rect 9129 8988 9181 9004
rect 9129 8954 9137 8988
rect 9171 8954 9181 8988
rect 8137 8883 8149 8943
rect 8183 8883 8195 8943
rect 8137 8871 8195 8883
rect 8701 8942 8759 8954
rect 8701 8882 8713 8942
rect 8747 8882 8759 8942
rect 8701 8870 8759 8882
rect 8789 8942 8851 8954
rect 8789 8882 8801 8942
rect 8835 8882 8851 8942
rect 8789 8870 8851 8882
rect 8881 8942 8947 8954
rect 8881 8882 8897 8942
rect 8931 8882 8947 8942
rect 8881 8870 8947 8882
rect 8977 8942 9039 8954
rect 8977 8882 8993 8942
rect 9027 8882 9039 8942
rect 8977 8870 9039 8882
rect 9129 8920 9181 8954
rect 9129 8886 9137 8920
rect 9171 8886 9181 8920
rect 9129 8874 9181 8886
rect 9211 8988 9263 9004
rect 9211 8954 9221 8988
rect 9255 8954 9263 8988
rect 9211 8920 9263 8954
rect 9211 8886 9221 8920
rect 9255 8886 9263 8920
rect 9211 8874 9263 8886
rect 9344 8956 9396 9004
rect 9344 8922 9352 8956
rect 9386 8922 9396 8956
rect 9344 8874 9396 8922
rect 9426 8992 9491 9004
rect 9426 8958 9436 8992
rect 9470 8958 9491 8992
rect 9426 8920 9491 8958
rect 9521 8966 9573 9004
rect 9521 8932 9531 8966
rect 9565 8932 9573 8966
rect 9521 8920 9573 8932
rect 9627 8958 9679 9004
rect 9627 8924 9635 8958
rect 9669 8924 9679 8958
rect 9426 8874 9476 8920
rect 9627 8874 9679 8924
rect 9709 8992 9774 9004
rect 9709 8958 9719 8992
rect 9753 8958 9774 8992
rect 9709 8920 9774 8958
rect 9804 8982 9856 9004
rect 9804 8948 9814 8982
rect 9848 8948 9856 8982
rect 9804 8920 9856 8948
rect 9910 8984 9962 9004
rect 9910 8950 9918 8984
rect 9952 8950 9962 8984
rect 9709 8874 9759 8920
rect 9910 8876 9962 8950
rect 9992 8932 10046 9004
rect 9992 8898 10002 8932
rect 10036 8898 10046 8932
rect 9992 8876 10046 8898
rect 10076 8976 10164 9004
rect 10076 8942 10102 8976
rect 10136 8942 10164 8976
rect 10076 8920 10164 8942
rect 10194 8996 10250 9004
rect 10194 8962 10204 8996
rect 10238 8962 10250 8996
rect 10194 8920 10250 8962
rect 10280 8932 10345 9004
rect 10375 8992 10454 9004
rect 10375 8958 10395 8992
rect 10429 8958 10454 8992
rect 10375 8932 10454 8958
rect 10484 8932 10549 9004
rect 10280 8920 10330 8932
rect 10076 8876 10126 8920
rect 2454 8609 2506 8625
rect 2454 8575 2462 8609
rect 2496 8575 2506 8609
rect 2454 8541 2506 8575
rect 2454 8507 2462 8541
rect 2496 8507 2506 8541
rect 2454 8495 2506 8507
rect 2536 8609 2588 8625
rect 2536 8575 2546 8609
rect 2580 8575 2588 8609
rect 2536 8541 2588 8575
rect 2536 8507 2546 8541
rect 2580 8507 2588 8541
rect 2536 8495 2588 8507
rect 2644 8609 2696 8625
rect 2644 8575 2652 8609
rect 2686 8575 2696 8609
rect 2644 8541 2696 8575
rect 2644 8507 2652 8541
rect 2686 8507 2696 8541
rect 2644 8495 2696 8507
rect 2726 8609 2778 8625
rect 2726 8575 2736 8609
rect 2770 8575 2778 8609
rect 2726 8541 2778 8575
rect 2726 8507 2736 8541
rect 2770 8507 2778 8541
rect 2726 8495 2778 8507
rect 10499 8876 10549 8932
rect 10579 8992 10631 9004
rect 10579 8958 10589 8992
rect 10623 8958 10631 8992
rect 10579 8876 10631 8958
rect 10685 8958 10737 9004
rect 10685 8924 10693 8958
rect 10727 8924 10737 8958
rect 10685 8876 10737 8924
rect 10767 8932 10821 9004
rect 10767 8898 10777 8932
rect 10811 8898 10821 8932
rect 10767 8876 10821 8898
rect 10851 8976 10921 9004
rect 10851 8942 10877 8976
rect 10911 8942 10921 8976
rect 10851 8920 10921 8942
rect 10951 8996 11031 9004
rect 10951 8962 10961 8996
rect 10995 8962 11031 8996
rect 10951 8920 11031 8962
rect 11061 8932 11127 9004
rect 11157 8992 11233 9004
rect 11157 8958 11178 8992
rect 11212 8958 11233 8992
rect 11157 8932 11233 8958
rect 11263 8974 11328 9004
rect 11263 8940 11284 8974
rect 11318 8940 11328 8974
rect 11263 8932 11328 8940
rect 11061 8920 11112 8932
rect 10851 8876 10901 8920
rect 11278 8920 11328 8932
rect 11358 8992 11410 9004
rect 11358 8958 11368 8992
rect 11402 8958 11410 8992
rect 11358 8920 11410 8958
rect 11464 8966 11516 9004
rect 11464 8932 11472 8966
rect 11506 8932 11516 8966
rect 11464 8920 11516 8932
rect 11546 8992 11600 9004
rect 11546 8958 11556 8992
rect 11590 8958 11600 8992
rect 11546 8920 11600 8958
rect 11630 8966 11682 9004
rect 13444 9008 13456 9068
rect 13490 9008 13502 9068
rect 13444 8996 13502 9008
rect 13532 9068 13590 9080
rect 13532 9008 13544 9068
rect 13578 9008 13590 9068
rect 19182 9055 19194 9115
rect 19228 9055 19240 9115
rect 19182 9043 19240 9055
rect 19270 9043 19312 9127
rect 19342 9115 19400 9127
rect 19342 9055 19354 9115
rect 19388 9055 19400 9115
rect 25891 9115 25949 9127
rect 19342 9043 19400 9055
rect 20153 9068 20211 9080
rect 13532 8996 13590 9008
rect 11630 8932 11640 8966
rect 11674 8932 11682 8966
rect 12676 8979 12728 8991
rect 11630 8920 11682 8932
rect 11821 8944 11883 8956
rect 11821 8884 11833 8944
rect 11867 8884 11883 8944
rect 11821 8872 11883 8884
rect 11913 8944 11979 8956
rect 11913 8884 11929 8944
rect 11963 8884 11979 8944
rect 11913 8872 11979 8884
rect 12009 8944 12075 8956
rect 12009 8884 12025 8944
rect 12059 8884 12075 8944
rect 12009 8872 12075 8884
rect 12105 8944 12167 8956
rect 12105 8884 12121 8944
rect 12155 8884 12167 8944
rect 12105 8872 12167 8884
rect 12221 8932 12279 8944
rect 12221 8872 12233 8932
rect 12267 8872 12279 8932
rect 12221 8860 12279 8872
rect 12309 8932 12367 8944
rect 12676 8945 12684 8979
rect 12718 8945 12728 8979
rect 12309 8872 12321 8932
rect 12355 8872 12367 8932
rect 12309 8860 12367 8872
rect 12422 8931 12480 8943
rect 12422 8871 12434 8931
rect 12468 8871 12480 8931
rect 12422 8859 12480 8871
rect 12510 8931 12568 8943
rect 12510 8871 12522 8931
rect 12556 8871 12568 8931
rect 12510 8859 12568 8871
rect 12676 8911 12728 8945
rect 12676 8877 12684 8911
rect 12718 8877 12728 8911
rect 12676 8861 12728 8877
rect 12758 8861 12812 8991
rect 12842 8979 12894 8991
rect 12842 8945 12852 8979
rect 12886 8945 12894 8979
rect 12842 8911 12894 8945
rect 12842 8877 12852 8911
rect 12886 8877 12894 8911
rect 12842 8861 12894 8877
rect 12999 8975 13051 8991
rect 12999 8941 13007 8975
rect 13041 8941 13051 8975
rect 12999 8907 13051 8941
rect 12999 8873 13007 8907
rect 13041 8873 13051 8907
rect 12999 8861 13051 8873
rect 13081 8975 13133 8991
rect 13081 8941 13091 8975
rect 13125 8941 13133 8975
rect 20153 9008 20165 9068
rect 20199 9008 20211 9068
rect 20153 8996 20211 9008
rect 20241 9068 20299 9080
rect 20241 9008 20253 9068
rect 20287 9008 20299 9068
rect 25891 9055 25903 9115
rect 25937 9055 25949 9115
rect 25891 9043 25949 9055
rect 25979 9043 26021 9127
rect 26051 9115 26109 9127
rect 26051 9055 26063 9115
rect 26097 9055 26109 9115
rect 26051 9043 26109 9055
rect 20241 8996 20299 9008
rect 13081 8907 13133 8941
rect 13081 8873 13091 8907
rect 13125 8873 13133 8907
rect 13081 8861 13133 8873
rect 13252 8930 13314 8942
rect 13252 8870 13264 8930
rect 13298 8870 13314 8930
rect 13252 8858 13314 8870
rect 13344 8930 13410 8942
rect 13344 8870 13360 8930
rect 13394 8870 13410 8930
rect 13344 8858 13410 8870
rect 13440 8930 13502 8942
rect 13440 8870 13456 8930
rect 13490 8870 13502 8930
rect 13440 8858 13502 8870
rect 13532 8930 13590 8942
rect 13532 8870 13544 8930
rect 13578 8870 13590 8930
rect 13532 8858 13590 8870
rect 14096 8931 14154 8943
rect 14096 8871 14108 8931
rect 14142 8871 14154 8931
rect 14096 8859 14154 8871
rect 14184 8931 14243 8943
rect 14184 8871 14197 8931
rect 14231 8871 14243 8931
rect 14184 8859 14243 8871
rect 14830 8931 14888 8943
rect 14830 8871 14842 8931
rect 14876 8871 14888 8931
rect 14830 8859 14888 8871
rect 14918 8931 15010 8943
rect 14918 8871 14944 8931
rect 14978 8871 15010 8931
rect 14918 8859 15010 8871
rect 15040 8931 15098 8943
rect 15040 8871 15052 8931
rect 15086 8871 15098 8931
rect 15040 8859 15098 8871
rect 16168 8931 16226 8943
rect 16168 8871 16180 8931
rect 16214 8871 16226 8931
rect 16168 8859 16226 8871
rect 16256 8931 16348 8943
rect 16256 8871 16284 8931
rect 16318 8871 16348 8931
rect 16256 8859 16348 8871
rect 16378 8931 16436 8943
rect 16378 8871 16390 8931
rect 16424 8871 16436 8931
rect 16378 8859 16436 8871
rect 17380 8931 17438 8943
rect 17380 8871 17392 8931
rect 17426 8871 17438 8931
rect 17380 8859 17438 8871
rect 17468 8931 17560 8943
rect 17468 8871 17495 8931
rect 17529 8871 17560 8931
rect 17468 8859 17560 8871
rect 17590 8931 17648 8943
rect 17590 8871 17602 8931
rect 17636 8871 17648 8931
rect 17590 8859 17648 8871
rect 18234 8931 18292 8943
rect 18234 8871 18244 8931
rect 18278 8871 18292 8931
rect 18234 8859 18292 8871
rect 18322 8931 18380 8943
rect 18322 8871 18334 8931
rect 18368 8871 18380 8931
rect 18322 8859 18380 8871
rect 19961 8930 20023 8942
rect 19961 8870 19973 8930
rect 20007 8870 20023 8930
rect 19961 8858 20023 8870
rect 20053 8930 20119 8942
rect 20053 8870 20069 8930
rect 20103 8870 20119 8930
rect 20053 8858 20119 8870
rect 20149 8930 20211 8942
rect 20149 8870 20165 8930
rect 20199 8870 20211 8930
rect 20149 8858 20211 8870
rect 20241 8930 20299 8942
rect 20241 8870 20253 8930
rect 20287 8870 20299 8930
rect 20241 8858 20299 8870
rect 20805 8931 20863 8943
rect 20805 8871 20817 8931
rect 20851 8871 20863 8931
rect 20805 8859 20863 8871
rect 20893 8931 20952 8943
rect 20893 8871 20906 8931
rect 20940 8871 20952 8931
rect 20893 8859 20952 8871
rect 21539 8931 21597 8943
rect 21539 8871 21551 8931
rect 21585 8871 21597 8931
rect 21539 8859 21597 8871
rect 21627 8931 21719 8943
rect 21627 8871 21653 8931
rect 21687 8871 21719 8931
rect 21627 8859 21719 8871
rect 21749 8931 21807 8943
rect 21749 8871 21761 8931
rect 21795 8871 21807 8931
rect 21749 8859 21807 8871
rect 22877 8931 22935 8943
rect 22877 8871 22889 8931
rect 22923 8871 22935 8931
rect 22877 8859 22935 8871
rect 22965 8931 23057 8943
rect 22965 8871 22993 8931
rect 23027 8871 23057 8931
rect 22965 8859 23057 8871
rect 23087 8931 23145 8943
rect 23087 8871 23099 8931
rect 23133 8871 23145 8931
rect 23087 8859 23145 8871
rect 24089 8931 24147 8943
rect 24089 8871 24101 8931
rect 24135 8871 24147 8931
rect 24089 8859 24147 8871
rect 24177 8931 24269 8943
rect 24177 8871 24204 8931
rect 24238 8871 24269 8931
rect 24177 8859 24269 8871
rect 24299 8931 24357 8943
rect 24299 8871 24311 8931
rect 24345 8871 24357 8931
rect 24299 8859 24357 8871
rect 24943 8931 25001 8943
rect 24943 8871 24953 8931
rect 24987 8871 25001 8931
rect 24943 8859 25001 8871
rect 25031 8931 25089 8943
rect 25031 8871 25043 8931
rect 25077 8871 25089 8931
rect 25031 8859 25089 8871
rect 19513 8597 19565 8613
rect 19513 8563 19521 8597
rect 19555 8563 19565 8597
rect 19513 8529 19565 8563
rect 19513 8495 19521 8529
rect 19555 8495 19565 8529
rect 19513 8483 19565 8495
rect 19595 8597 19647 8613
rect 19595 8563 19605 8597
rect 19639 8563 19647 8597
rect 19595 8529 19647 8563
rect 19595 8495 19605 8529
rect 19639 8495 19647 8529
rect 19595 8483 19647 8495
rect 19703 8597 19755 8613
rect 19703 8563 19711 8597
rect 19745 8563 19755 8597
rect 19703 8529 19755 8563
rect 19703 8495 19711 8529
rect 19745 8495 19755 8529
rect 19703 8483 19755 8495
rect 19785 8597 19837 8613
rect 19785 8563 19795 8597
rect 19829 8563 19837 8597
rect 19785 8529 19837 8563
rect 19785 8495 19795 8529
rect 19829 8495 19837 8529
rect 26222 8597 26274 8613
rect 26222 8563 26230 8597
rect 26264 8563 26274 8597
rect 26222 8529 26274 8563
rect 19785 8483 19837 8495
rect 26222 8495 26230 8529
rect 26264 8495 26274 8529
rect 26222 8483 26274 8495
rect 26304 8597 26356 8613
rect 26304 8563 26314 8597
rect 26348 8563 26356 8597
rect 26304 8529 26356 8563
rect 26304 8495 26314 8529
rect 26348 8495 26356 8529
rect 26304 8483 26356 8495
rect 26412 8597 26464 8613
rect 26412 8563 26420 8597
rect 26454 8563 26464 8597
rect 26412 8529 26464 8563
rect 26412 8495 26420 8529
rect 26454 8495 26464 8529
rect 26412 8483 26464 8495
rect 26494 8597 26546 8613
rect 26494 8563 26504 8597
rect 26538 8563 26546 8597
rect 26494 8529 26546 8563
rect 26494 8495 26504 8529
rect 26538 8495 26546 8529
rect 26494 8483 26546 8495
rect 10081 7900 10133 7965
rect 10081 7866 10089 7900
rect 10123 7866 10133 7900
rect 10081 7835 10133 7866
rect 10163 7919 10215 7965
rect 10163 7881 10242 7919
rect 10163 7847 10173 7881
rect 10207 7847 10242 7881
rect 10163 7835 10242 7847
rect 10272 7835 10338 7919
rect 10368 7896 10463 7919
rect 10368 7862 10380 7896
rect 10414 7862 10463 7896
rect 10368 7835 10463 7862
rect 10493 7835 10559 7919
rect 10589 7896 10727 7919
rect 10589 7862 10615 7896
rect 10649 7862 10683 7896
rect 10717 7862 10727 7896
rect 10589 7835 10727 7862
rect 10757 7896 10809 7919
rect 10757 7862 10767 7896
rect 10801 7862 10809 7896
rect 10757 7835 10809 7862
rect 10908 7900 10960 7965
rect 10908 7866 10916 7900
rect 10950 7866 10960 7900
rect 10908 7835 10960 7866
rect 10990 7919 11042 7965
rect 12690 8140 12748 8152
rect 12690 8080 12702 8140
rect 12736 8080 12748 8140
rect 12690 8068 12748 8080
rect 12778 8140 12836 8152
rect 12778 8080 12790 8140
rect 12824 8080 12836 8140
rect 12778 8068 12836 8080
rect 12221 7952 12279 7964
rect 11821 7940 11883 7952
rect 10990 7881 11069 7919
rect 10990 7847 11000 7881
rect 11034 7847 11069 7881
rect 10990 7835 11069 7847
rect 11099 7835 11165 7919
rect 11195 7896 11290 7919
rect 11195 7862 11207 7896
rect 11241 7862 11290 7896
rect 11195 7835 11290 7862
rect 11320 7835 11386 7919
rect 11416 7896 11554 7919
rect 11416 7862 11442 7896
rect 11476 7862 11510 7896
rect 11544 7862 11554 7896
rect 11416 7835 11554 7862
rect 11584 7896 11636 7919
rect 11584 7862 11594 7896
rect 11628 7862 11636 7896
rect 11821 7880 11833 7940
rect 11867 7880 11883 7940
rect 11821 7868 11883 7880
rect 11913 7940 11979 7952
rect 11913 7880 11929 7940
rect 11963 7880 11979 7940
rect 11913 7868 11979 7880
rect 12009 7940 12075 7952
rect 12009 7880 12025 7940
rect 12059 7880 12075 7940
rect 12009 7868 12075 7880
rect 12105 7940 12167 7952
rect 12105 7880 12121 7940
rect 12155 7880 12167 7940
rect 12221 7892 12233 7952
rect 12267 7892 12279 7952
rect 12221 7880 12279 7892
rect 12309 7952 12367 7964
rect 12309 7892 12321 7952
rect 12355 7892 12367 7952
rect 12309 7880 12367 7892
rect 12105 7868 12167 7880
rect 11584 7835 11636 7862
rect 11525 6639 11577 6684
rect 11525 6605 11533 6639
rect 11567 6605 11577 6639
rect 11525 6580 11577 6605
rect 11607 6626 11665 6684
rect 11607 6592 11619 6626
rect 11653 6592 11665 6626
rect 11607 6580 11665 6592
rect 11695 6656 11747 6684
rect 11695 6622 11705 6656
rect 11739 6622 11747 6656
rect 11695 6580 11747 6622
rect 11801 6662 11853 6710
rect 11801 6628 11809 6662
rect 11843 6628 11853 6662
rect 11801 6580 11853 6628
rect 11883 6630 11937 6710
rect 11883 6596 11893 6630
rect 11927 6596 11937 6630
rect 11883 6580 11937 6596
rect 11967 6662 12021 6710
rect 11967 6628 11977 6662
rect 12011 6628 12021 6662
rect 11967 6580 12021 6628
rect 12051 6630 12105 6710
rect 12051 6596 12061 6630
rect 12095 6596 12105 6630
rect 12051 6580 12105 6596
rect 12135 6662 12189 6710
rect 12135 6628 12145 6662
rect 12179 6628 12189 6662
rect 12135 6580 12189 6628
rect 12219 6694 12271 6710
rect 12219 6660 12229 6694
rect 12263 6660 12271 6694
rect 12219 6626 12271 6660
rect 12219 6592 12229 6626
rect 12263 6592 12271 6626
rect 12219 6580 12271 6592
rect 12785 6694 12852 6710
rect 12785 6660 12793 6694
rect 12827 6660 12852 6694
rect 12785 6626 12852 6660
rect 12785 6592 12793 6626
rect 12827 6592 12852 6626
rect 12785 6580 12852 6592
rect 12882 6662 12936 6710
rect 12882 6628 12892 6662
rect 12926 6628 12936 6662
rect 12882 6580 12936 6628
rect 12966 6694 13036 6710
rect 12966 6660 12976 6694
rect 13010 6660 13036 6694
rect 12966 6626 13036 6660
rect 12966 6592 12976 6626
rect 13010 6592 13036 6626
rect 12966 6580 13036 6592
rect 13066 6662 13120 6710
rect 13066 6628 13076 6662
rect 13110 6628 13120 6662
rect 13066 6580 13120 6628
rect 13150 6664 13206 6710
rect 13150 6652 13221 6664
rect 13150 6618 13160 6652
rect 13194 6618 13221 6652
rect 13150 6580 13221 6618
rect 13251 6652 13301 6664
rect 13471 6652 13533 6664
rect 13251 6580 13316 6652
rect 13346 6626 13426 6652
rect 13346 6592 13369 6626
rect 13403 6592 13426 6626
rect 13346 6580 13426 6592
rect 13456 6580 13533 6652
rect 13563 6626 13615 6664
rect 13563 6592 13573 6626
rect 13607 6592 13615 6626
rect 13563 6580 13615 6592
rect 13669 6634 13721 6664
rect 13669 6600 13677 6634
rect 13711 6600 13721 6634
rect 13669 6580 13721 6600
rect 13751 6652 13806 6664
rect 13751 6618 13761 6652
rect 13795 6618 13806 6652
rect 13751 6580 13806 6618
rect 13836 6652 13888 6664
rect 13836 6618 13846 6652
rect 13880 6618 13888 6652
rect 13836 6580 13888 6618
rect 13942 6626 13996 6664
rect 13942 6592 13950 6626
rect 13984 6592 13996 6626
rect 13942 6580 13996 6592
rect 14026 6626 14104 6664
rect 14026 6592 14049 6626
rect 14083 6592 14104 6626
rect 14026 6580 14104 6592
rect 14134 6652 14185 6664
rect 14355 6652 14405 6664
rect 14134 6580 14200 6652
rect 14230 6640 14310 6652
rect 14230 6606 14253 6640
rect 14287 6606 14310 6640
rect 14230 6580 14310 6606
rect 14340 6580 14405 6652
rect 14435 6626 14489 6664
rect 14435 6592 14445 6626
rect 14479 6592 14489 6626
rect 14435 6580 14489 6592
rect 14519 6652 14571 6664
rect 14519 6618 14529 6652
rect 14563 6618 14571 6652
rect 14519 6580 14571 6618
rect 24067 6317 24119 6329
rect 24067 6283 24075 6317
rect 24109 6283 24119 6317
rect 24067 6249 24119 6283
rect 24067 6215 24075 6249
rect 24109 6215 24119 6249
rect 24067 6199 24119 6215
rect 24149 6317 24201 6329
rect 24149 6283 24159 6317
rect 24193 6283 24201 6317
rect 24149 6249 24201 6283
rect 24149 6215 24159 6249
rect 24193 6215 24201 6249
rect 24149 6199 24201 6215
rect 24257 6317 24309 6329
rect 24257 6283 24265 6317
rect 24299 6283 24309 6317
rect 24257 6249 24309 6283
rect 24257 6215 24265 6249
rect 24299 6215 24309 6249
rect 24257 6199 24309 6215
rect 24339 6317 24391 6329
rect 24339 6283 24349 6317
rect 24383 6283 24391 6317
rect 24339 6249 24391 6283
rect 24339 6215 24349 6249
rect 24383 6215 24391 6249
rect 24339 6199 24391 6215
rect 11524 5779 11576 5791
rect 11524 5745 11532 5779
rect 11566 5745 11576 5779
rect 11524 5707 11576 5745
rect 11606 5753 11660 5791
rect 11606 5719 11616 5753
rect 11650 5719 11660 5753
rect 11606 5707 11660 5719
rect 11690 5779 11742 5791
rect 11690 5745 11700 5779
rect 11734 5745 11742 5779
rect 11690 5707 11742 5745
rect 11796 5753 11848 5791
rect 11796 5719 11804 5753
rect 11838 5719 11848 5753
rect 11796 5707 11848 5719
rect 11878 5779 11928 5791
rect 12305 5791 12355 5835
rect 12094 5779 12145 5791
rect 11878 5771 11943 5779
rect 11878 5737 11888 5771
rect 11922 5737 11943 5771
rect 11878 5707 11943 5737
rect 11973 5753 12049 5779
rect 11973 5719 11994 5753
rect 12028 5719 12049 5753
rect 11973 5707 12049 5719
rect 12079 5707 12145 5779
rect 12175 5749 12255 5791
rect 12175 5715 12211 5749
rect 12245 5715 12255 5749
rect 12175 5707 12255 5715
rect 12285 5769 12355 5791
rect 12285 5735 12295 5769
rect 12329 5735 12355 5769
rect 12285 5707 12355 5735
rect 12385 5813 12439 5835
rect 12385 5779 12395 5813
rect 12429 5779 12439 5813
rect 12385 5707 12439 5779
rect 12469 5787 12521 5835
rect 12469 5753 12479 5787
rect 12513 5753 12521 5787
rect 12469 5707 12521 5753
rect 12575 5753 12627 5835
rect 12575 5719 12583 5753
rect 12617 5719 12627 5753
rect 12575 5707 12627 5719
rect 12657 5779 12707 5835
rect 13080 5791 13130 5835
rect 12876 5779 12926 5791
rect 12657 5707 12722 5779
rect 12752 5753 12831 5779
rect 12752 5719 12777 5753
rect 12811 5719 12831 5753
rect 12752 5707 12831 5719
rect 12861 5707 12926 5779
rect 12956 5749 13012 5791
rect 12956 5715 12968 5749
rect 13002 5715 13012 5749
rect 12956 5707 13012 5715
rect 13042 5769 13130 5791
rect 13042 5735 13070 5769
rect 13104 5735 13130 5769
rect 13042 5707 13130 5735
rect 13160 5813 13214 5835
rect 13160 5779 13170 5813
rect 13204 5779 13214 5813
rect 13160 5707 13214 5779
rect 13244 5761 13296 5835
rect 13447 5791 13497 5837
rect 13244 5727 13254 5761
rect 13288 5727 13296 5761
rect 13244 5707 13296 5727
rect 13350 5763 13402 5791
rect 13350 5729 13358 5763
rect 13392 5729 13402 5763
rect 13350 5707 13402 5729
rect 13432 5753 13497 5791
rect 13432 5719 13453 5753
rect 13487 5719 13497 5753
rect 13432 5707 13497 5719
rect 13527 5787 13579 5837
rect 13730 5791 13780 5837
rect 13527 5753 13537 5787
rect 13571 5753 13579 5787
rect 13527 5707 13579 5753
rect 13633 5779 13685 5791
rect 13633 5745 13641 5779
rect 13675 5745 13685 5779
rect 13633 5707 13685 5745
rect 13715 5753 13780 5791
rect 13715 5719 13736 5753
rect 13770 5719 13780 5753
rect 13715 5707 13780 5719
rect 13810 5789 13862 5837
rect 13810 5755 13820 5789
rect 13854 5755 13862 5789
rect 13810 5707 13862 5755
rect 13916 5779 13968 5791
rect 13916 5745 13924 5779
rect 13958 5745 13968 5779
rect 13916 5707 13968 5745
rect 13998 5753 14052 5791
rect 13998 5719 14008 5753
rect 14042 5719 14052 5753
rect 13998 5707 14052 5719
rect 14082 5779 14134 5791
rect 14082 5745 14092 5779
rect 14126 5745 14134 5779
rect 14082 5707 14134 5745
rect 14188 5753 14240 5791
rect 14188 5719 14196 5753
rect 14230 5719 14240 5753
rect 14188 5707 14240 5719
rect 14270 5779 14320 5791
rect 14697 5791 14747 5835
rect 14486 5779 14537 5791
rect 14270 5771 14335 5779
rect 14270 5737 14280 5771
rect 14314 5737 14335 5771
rect 14270 5707 14335 5737
rect 14365 5753 14441 5779
rect 14365 5719 14386 5753
rect 14420 5719 14441 5753
rect 14365 5707 14441 5719
rect 14471 5707 14537 5779
rect 14567 5749 14647 5791
rect 14567 5715 14603 5749
rect 14637 5715 14647 5749
rect 14567 5707 14647 5715
rect 14677 5769 14747 5791
rect 14677 5735 14687 5769
rect 14721 5735 14747 5769
rect 14677 5707 14747 5735
rect 14777 5813 14831 5835
rect 14777 5779 14787 5813
rect 14821 5779 14831 5813
rect 14777 5707 14831 5779
rect 14861 5787 14913 5835
rect 14861 5753 14871 5787
rect 14905 5753 14913 5787
rect 14861 5707 14913 5753
rect 14967 5753 15019 5835
rect 14967 5719 14975 5753
rect 15009 5719 15019 5753
rect 14967 5707 15019 5719
rect 15049 5779 15099 5835
rect 15472 5791 15522 5835
rect 15268 5779 15318 5791
rect 15049 5707 15114 5779
rect 15144 5753 15223 5779
rect 15144 5719 15169 5753
rect 15203 5719 15223 5753
rect 15144 5707 15223 5719
rect 15253 5707 15318 5779
rect 15348 5749 15404 5791
rect 15348 5715 15360 5749
rect 15394 5715 15404 5749
rect 15348 5707 15404 5715
rect 15434 5769 15522 5791
rect 15434 5735 15462 5769
rect 15496 5735 15522 5769
rect 15434 5707 15522 5735
rect 15552 5813 15606 5835
rect 15552 5779 15562 5813
rect 15596 5779 15606 5813
rect 15552 5707 15606 5779
rect 15636 5761 15688 5835
rect 15839 5791 15889 5837
rect 15636 5727 15646 5761
rect 15680 5727 15688 5761
rect 15636 5707 15688 5727
rect 15742 5763 15794 5791
rect 15742 5729 15750 5763
rect 15784 5729 15794 5763
rect 15742 5707 15794 5729
rect 15824 5753 15889 5791
rect 15824 5719 15845 5753
rect 15879 5719 15889 5753
rect 15824 5707 15889 5719
rect 15919 5787 15971 5837
rect 16122 5791 16172 5837
rect 15919 5753 15929 5787
rect 15963 5753 15971 5787
rect 15919 5707 15971 5753
rect 16025 5779 16077 5791
rect 16025 5745 16033 5779
rect 16067 5745 16077 5779
rect 16025 5707 16077 5745
rect 16107 5753 16172 5791
rect 16107 5719 16128 5753
rect 16162 5719 16172 5753
rect 16107 5707 16172 5719
rect 16202 5789 16254 5837
rect 16202 5755 16212 5789
rect 16246 5755 16254 5789
rect 16202 5707 16254 5755
rect 16308 5779 16360 5791
rect 16308 5745 16316 5779
rect 16350 5745 16360 5779
rect 16308 5707 16360 5745
rect 16390 5753 16444 5791
rect 16390 5719 16400 5753
rect 16434 5719 16444 5753
rect 16390 5707 16444 5719
rect 16474 5779 16526 5791
rect 16474 5745 16484 5779
rect 16518 5745 16526 5779
rect 16474 5707 16526 5745
rect 16580 5753 16632 5791
rect 16580 5719 16588 5753
rect 16622 5719 16632 5753
rect 16580 5707 16632 5719
rect 16662 5779 16712 5791
rect 17089 5791 17139 5835
rect 16878 5779 16929 5791
rect 16662 5771 16727 5779
rect 16662 5737 16672 5771
rect 16706 5737 16727 5771
rect 16662 5707 16727 5737
rect 16757 5753 16833 5779
rect 16757 5719 16778 5753
rect 16812 5719 16833 5753
rect 16757 5707 16833 5719
rect 16863 5707 16929 5779
rect 16959 5749 17039 5791
rect 16959 5715 16995 5749
rect 17029 5715 17039 5749
rect 16959 5707 17039 5715
rect 17069 5769 17139 5791
rect 17069 5735 17079 5769
rect 17113 5735 17139 5769
rect 17069 5707 17139 5735
rect 17169 5813 17223 5835
rect 17169 5779 17179 5813
rect 17213 5779 17223 5813
rect 17169 5707 17223 5779
rect 17253 5787 17305 5835
rect 17253 5753 17263 5787
rect 17297 5753 17305 5787
rect 17253 5707 17305 5753
rect 17359 5753 17411 5835
rect 17359 5719 17367 5753
rect 17401 5719 17411 5753
rect 17359 5707 17411 5719
rect 17441 5779 17491 5835
rect 17864 5791 17914 5835
rect 17660 5779 17710 5791
rect 17441 5707 17506 5779
rect 17536 5753 17615 5779
rect 17536 5719 17561 5753
rect 17595 5719 17615 5753
rect 17536 5707 17615 5719
rect 17645 5707 17710 5779
rect 17740 5749 17796 5791
rect 17740 5715 17752 5749
rect 17786 5715 17796 5749
rect 17740 5707 17796 5715
rect 17826 5769 17914 5791
rect 17826 5735 17854 5769
rect 17888 5735 17914 5769
rect 17826 5707 17914 5735
rect 17944 5813 17998 5835
rect 17944 5779 17954 5813
rect 17988 5779 17998 5813
rect 17944 5707 17998 5779
rect 18028 5761 18080 5835
rect 18231 5791 18281 5837
rect 18028 5727 18038 5761
rect 18072 5727 18080 5761
rect 18028 5707 18080 5727
rect 18134 5763 18186 5791
rect 18134 5729 18142 5763
rect 18176 5729 18186 5763
rect 18134 5707 18186 5729
rect 18216 5753 18281 5791
rect 18216 5719 18237 5753
rect 18271 5719 18281 5753
rect 18216 5707 18281 5719
rect 18311 5787 18363 5837
rect 18514 5791 18564 5837
rect 18311 5753 18321 5787
rect 18355 5753 18363 5787
rect 18311 5707 18363 5753
rect 18417 5779 18469 5791
rect 18417 5745 18425 5779
rect 18459 5745 18469 5779
rect 18417 5707 18469 5745
rect 18499 5753 18564 5791
rect 18499 5719 18520 5753
rect 18554 5719 18564 5753
rect 18499 5707 18564 5719
rect 18594 5789 18646 5837
rect 18594 5755 18604 5789
rect 18638 5755 18646 5789
rect 18594 5707 18646 5755
rect 18700 5779 18752 5791
rect 18700 5745 18708 5779
rect 18742 5745 18752 5779
rect 18700 5707 18752 5745
rect 18782 5753 18836 5791
rect 18782 5719 18792 5753
rect 18826 5719 18836 5753
rect 18782 5707 18836 5719
rect 18866 5779 18918 5791
rect 18866 5745 18876 5779
rect 18910 5745 18918 5779
rect 18866 5707 18918 5745
rect 18972 5753 19024 5791
rect 18972 5719 18980 5753
rect 19014 5719 19024 5753
rect 18972 5707 19024 5719
rect 19054 5779 19104 5791
rect 19481 5791 19531 5835
rect 19270 5779 19321 5791
rect 19054 5771 19119 5779
rect 19054 5737 19064 5771
rect 19098 5737 19119 5771
rect 19054 5707 19119 5737
rect 19149 5753 19225 5779
rect 19149 5719 19170 5753
rect 19204 5719 19225 5753
rect 19149 5707 19225 5719
rect 19255 5707 19321 5779
rect 19351 5749 19431 5791
rect 19351 5715 19387 5749
rect 19421 5715 19431 5749
rect 19351 5707 19431 5715
rect 19461 5769 19531 5791
rect 19461 5735 19471 5769
rect 19505 5735 19531 5769
rect 19461 5707 19531 5735
rect 19561 5813 19615 5835
rect 19561 5779 19571 5813
rect 19605 5779 19615 5813
rect 19561 5707 19615 5779
rect 19645 5787 19697 5835
rect 19645 5753 19655 5787
rect 19689 5753 19697 5787
rect 19645 5707 19697 5753
rect 19751 5753 19803 5835
rect 19751 5719 19759 5753
rect 19793 5719 19803 5753
rect 19751 5707 19803 5719
rect 19833 5779 19883 5835
rect 20256 5791 20306 5835
rect 20052 5779 20102 5791
rect 19833 5707 19898 5779
rect 19928 5753 20007 5779
rect 19928 5719 19953 5753
rect 19987 5719 20007 5753
rect 19928 5707 20007 5719
rect 20037 5707 20102 5779
rect 20132 5749 20188 5791
rect 20132 5715 20144 5749
rect 20178 5715 20188 5749
rect 20132 5707 20188 5715
rect 20218 5769 20306 5791
rect 20218 5735 20246 5769
rect 20280 5735 20306 5769
rect 20218 5707 20306 5735
rect 20336 5813 20390 5835
rect 20336 5779 20346 5813
rect 20380 5779 20390 5813
rect 20336 5707 20390 5779
rect 20420 5761 20472 5835
rect 20623 5791 20673 5837
rect 20420 5727 20430 5761
rect 20464 5727 20472 5761
rect 20420 5707 20472 5727
rect 20526 5763 20578 5791
rect 20526 5729 20534 5763
rect 20568 5729 20578 5763
rect 20526 5707 20578 5729
rect 20608 5753 20673 5791
rect 20608 5719 20629 5753
rect 20663 5719 20673 5753
rect 20608 5707 20673 5719
rect 20703 5787 20755 5837
rect 20906 5791 20956 5837
rect 20703 5753 20713 5787
rect 20747 5753 20755 5787
rect 20703 5707 20755 5753
rect 20809 5779 20861 5791
rect 20809 5745 20817 5779
rect 20851 5745 20861 5779
rect 20809 5707 20861 5745
rect 20891 5753 20956 5791
rect 20891 5719 20912 5753
rect 20946 5719 20956 5753
rect 20891 5707 20956 5719
rect 20986 5789 21038 5837
rect 20986 5755 20996 5789
rect 21030 5755 21038 5789
rect 20986 5707 21038 5755
rect 21092 5779 21144 5791
rect 21092 5745 21100 5779
rect 21134 5745 21144 5779
rect 21092 5707 21144 5745
rect 21174 5753 21228 5791
rect 21174 5719 21184 5753
rect 21218 5719 21228 5753
rect 21174 5707 21228 5719
rect 21258 5779 21310 5791
rect 21258 5745 21268 5779
rect 21302 5745 21310 5779
rect 21258 5707 21310 5745
rect 21364 5753 21416 5791
rect 21364 5719 21372 5753
rect 21406 5719 21416 5753
rect 21364 5707 21416 5719
rect 21446 5779 21496 5791
rect 21873 5791 21923 5835
rect 21662 5779 21713 5791
rect 21446 5771 21511 5779
rect 21446 5737 21456 5771
rect 21490 5737 21511 5771
rect 21446 5707 21511 5737
rect 21541 5753 21617 5779
rect 21541 5719 21562 5753
rect 21596 5719 21617 5753
rect 21541 5707 21617 5719
rect 21647 5707 21713 5779
rect 21743 5749 21823 5791
rect 21743 5715 21779 5749
rect 21813 5715 21823 5749
rect 21743 5707 21823 5715
rect 21853 5769 21923 5791
rect 21853 5735 21863 5769
rect 21897 5735 21923 5769
rect 21853 5707 21923 5735
rect 21953 5813 22007 5835
rect 21953 5779 21963 5813
rect 21997 5779 22007 5813
rect 21953 5707 22007 5779
rect 22037 5787 22089 5835
rect 22037 5753 22047 5787
rect 22081 5753 22089 5787
rect 22037 5707 22089 5753
rect 22143 5753 22195 5835
rect 22143 5719 22151 5753
rect 22185 5719 22195 5753
rect 22143 5707 22195 5719
rect 22225 5779 22275 5835
rect 22648 5791 22698 5835
rect 22444 5779 22494 5791
rect 22225 5707 22290 5779
rect 22320 5753 22399 5779
rect 22320 5719 22345 5753
rect 22379 5719 22399 5753
rect 22320 5707 22399 5719
rect 22429 5707 22494 5779
rect 22524 5749 22580 5791
rect 22524 5715 22536 5749
rect 22570 5715 22580 5749
rect 22524 5707 22580 5715
rect 22610 5769 22698 5791
rect 22610 5735 22638 5769
rect 22672 5735 22698 5769
rect 22610 5707 22698 5735
rect 22728 5813 22782 5835
rect 22728 5779 22738 5813
rect 22772 5779 22782 5813
rect 22728 5707 22782 5779
rect 22812 5761 22864 5835
rect 23015 5791 23065 5837
rect 22812 5727 22822 5761
rect 22856 5727 22864 5761
rect 22812 5707 22864 5727
rect 22918 5763 22970 5791
rect 22918 5729 22926 5763
rect 22960 5729 22970 5763
rect 22918 5707 22970 5729
rect 23000 5753 23065 5791
rect 23000 5719 23021 5753
rect 23055 5719 23065 5753
rect 23000 5707 23065 5719
rect 23095 5787 23147 5837
rect 25524 5941 25582 5953
rect 25524 5881 25536 5941
rect 25570 5881 25582 5941
rect 25524 5869 25582 5881
rect 25612 5941 25670 5953
rect 25612 5881 25626 5941
rect 25660 5881 25670 5941
rect 25612 5869 25670 5881
rect 26256 5941 26314 5953
rect 26256 5881 26268 5941
rect 26302 5881 26314 5941
rect 26256 5869 26314 5881
rect 26344 5941 26436 5953
rect 26344 5881 26375 5941
rect 26409 5881 26436 5941
rect 26344 5869 26436 5881
rect 26466 5941 26524 5953
rect 26466 5881 26478 5941
rect 26512 5881 26524 5941
rect 26466 5869 26524 5881
rect 27468 5941 27526 5953
rect 27468 5881 27480 5941
rect 27514 5881 27526 5941
rect 27468 5869 27526 5881
rect 27556 5941 27648 5953
rect 27556 5881 27586 5941
rect 27620 5881 27648 5941
rect 27556 5869 27648 5881
rect 27678 5941 27736 5953
rect 27678 5881 27690 5941
rect 27724 5881 27736 5941
rect 27678 5869 27736 5881
rect 28806 5941 28864 5953
rect 28806 5881 28818 5941
rect 28852 5881 28864 5941
rect 28806 5869 28864 5881
rect 28894 5941 28986 5953
rect 28894 5881 28926 5941
rect 28960 5881 28986 5941
rect 28894 5869 28986 5881
rect 29016 5941 29074 5953
rect 29016 5881 29028 5941
rect 29062 5881 29074 5941
rect 29016 5869 29074 5881
rect 29661 5941 29720 5953
rect 29661 5881 29673 5941
rect 29707 5881 29720 5941
rect 29661 5869 29720 5881
rect 29750 5941 29808 5953
rect 29750 5881 29762 5941
rect 29796 5881 29808 5941
rect 29750 5869 29808 5881
rect 30314 5942 30372 5954
rect 30314 5882 30326 5942
rect 30360 5882 30372 5942
rect 30314 5870 30372 5882
rect 30402 5942 30464 5954
rect 30402 5882 30414 5942
rect 30448 5882 30464 5942
rect 30402 5870 30464 5882
rect 30494 5942 30560 5954
rect 30494 5882 30510 5942
rect 30544 5882 30560 5942
rect 30494 5870 30560 5882
rect 30590 5942 30652 5954
rect 30590 5882 30606 5942
rect 30640 5882 30652 5942
rect 30803 5906 30853 5952
rect 30590 5870 30652 5882
rect 30706 5881 30758 5906
rect 23298 5791 23348 5837
rect 23095 5753 23105 5787
rect 23139 5753 23147 5787
rect 23095 5707 23147 5753
rect 23201 5779 23253 5791
rect 23201 5745 23209 5779
rect 23243 5745 23253 5779
rect 23201 5707 23253 5745
rect 23283 5753 23348 5791
rect 23283 5719 23304 5753
rect 23338 5719 23348 5753
rect 23283 5707 23348 5719
rect 23378 5789 23430 5837
rect 23378 5755 23388 5789
rect 23422 5755 23430 5789
rect 30706 5847 30714 5881
rect 30748 5847 30758 5881
rect 30706 5822 30758 5847
rect 30788 5868 30853 5906
rect 30788 5834 30807 5868
rect 30841 5834 30853 5868
rect 30788 5822 30853 5834
rect 30883 5898 30937 5952
rect 30883 5864 30893 5898
rect 30927 5864 30937 5898
rect 30883 5822 30937 5864
rect 30967 5940 31020 5952
rect 30967 5906 30977 5940
rect 31011 5906 31020 5940
rect 30967 5872 31020 5906
rect 30967 5838 30977 5872
rect 31011 5838 31020 5872
rect 30967 5822 31020 5838
rect 30314 5804 30372 5816
rect 23378 5707 23430 5755
rect 24504 5757 24562 5769
rect 24504 5697 24516 5757
rect 24550 5697 24562 5757
rect 24504 5685 24562 5697
rect 24592 5685 24634 5769
rect 24664 5757 24722 5769
rect 24664 5697 24676 5757
rect 24710 5697 24722 5757
rect 30314 5744 30326 5804
rect 30360 5744 30372 5804
rect 30314 5732 30372 5744
rect 30402 5804 30460 5816
rect 30402 5744 30414 5804
rect 30448 5744 30460 5804
rect 30402 5732 30460 5744
rect 24664 5685 24722 5697
rect 24504 5619 24562 5631
rect 24504 5559 24516 5619
rect 24550 5559 24562 5619
rect 24504 5547 24562 5559
rect 24592 5547 24634 5631
rect 24664 5619 24722 5631
rect 24664 5559 24676 5619
rect 24710 5559 24722 5619
rect 24664 5547 24722 5559
rect 11084 5077 11136 5122
rect 11084 5043 11092 5077
rect 11126 5043 11136 5077
rect 11084 5018 11136 5043
rect 11166 5064 11224 5122
rect 11166 5030 11178 5064
rect 11212 5030 11224 5064
rect 11166 5018 11224 5030
rect 11254 5094 11306 5122
rect 11254 5060 11264 5094
rect 11298 5060 11306 5094
rect 11254 5018 11306 5060
rect 11360 5100 11412 5148
rect 11360 5066 11368 5100
rect 11402 5066 11412 5100
rect 11360 5018 11412 5066
rect 11442 5068 11496 5148
rect 11442 5034 11452 5068
rect 11486 5034 11496 5068
rect 11442 5018 11496 5034
rect 11526 5100 11580 5148
rect 11526 5066 11536 5100
rect 11570 5066 11580 5100
rect 11526 5018 11580 5066
rect 11610 5068 11664 5148
rect 11610 5034 11620 5068
rect 11654 5034 11664 5068
rect 11610 5018 11664 5034
rect 11694 5100 11748 5148
rect 11694 5066 11704 5100
rect 11738 5066 11748 5100
rect 11694 5018 11748 5066
rect 11778 5132 11830 5148
rect 11778 5098 11788 5132
rect 11822 5098 11830 5132
rect 11778 5064 11830 5098
rect 11778 5030 11788 5064
rect 11822 5030 11830 5064
rect 11778 5018 11830 5030
rect 11892 5136 11944 5148
rect 11892 5102 11900 5136
rect 11934 5102 11944 5136
rect 11892 5068 11944 5102
rect 11892 5034 11900 5068
rect 11934 5034 11944 5068
rect 11892 5018 11944 5034
rect 11974 5136 12028 5148
rect 11974 5102 11984 5136
rect 12018 5102 12028 5136
rect 11974 5068 12028 5102
rect 11974 5034 11984 5068
rect 12018 5034 12028 5068
rect 11974 5018 12028 5034
rect 12058 5068 12112 5148
rect 12058 5034 12068 5068
rect 12102 5034 12112 5068
rect 12058 5018 12112 5034
rect 12142 5136 12196 5148
rect 12142 5102 12152 5136
rect 12186 5102 12196 5136
rect 12142 5068 12196 5102
rect 12142 5034 12152 5068
rect 12186 5034 12196 5068
rect 12142 5018 12196 5034
rect 12226 5068 12280 5148
rect 12226 5034 12236 5068
rect 12270 5034 12280 5068
rect 12226 5018 12280 5034
rect 12310 5136 12364 5148
rect 12310 5102 12320 5136
rect 12354 5102 12364 5136
rect 12310 5068 12364 5102
rect 12310 5034 12320 5068
rect 12354 5034 12364 5068
rect 12310 5018 12364 5034
rect 12394 5068 12448 5148
rect 12394 5034 12404 5068
rect 12438 5034 12448 5068
rect 12394 5018 12448 5034
rect 12478 5136 12532 5148
rect 12478 5102 12488 5136
rect 12522 5102 12532 5136
rect 12478 5068 12532 5102
rect 12478 5034 12488 5068
rect 12522 5034 12532 5068
rect 12478 5018 12532 5034
rect 12562 5068 12616 5148
rect 12562 5034 12572 5068
rect 12606 5034 12616 5068
rect 12562 5018 12616 5034
rect 12646 5136 12700 5148
rect 12646 5102 12656 5136
rect 12690 5102 12700 5136
rect 12646 5068 12700 5102
rect 12646 5034 12656 5068
rect 12690 5034 12700 5068
rect 12646 5018 12700 5034
rect 12730 5068 12784 5148
rect 12730 5034 12740 5068
rect 12774 5034 12784 5068
rect 12730 5018 12784 5034
rect 12814 5136 12868 5148
rect 12814 5102 12824 5136
rect 12858 5102 12868 5136
rect 12814 5068 12868 5102
rect 12814 5034 12824 5068
rect 12858 5034 12868 5068
rect 12814 5018 12868 5034
rect 12898 5068 12952 5148
rect 12898 5034 12908 5068
rect 12942 5034 12952 5068
rect 12898 5018 12952 5034
rect 12982 5136 13036 5148
rect 12982 5102 12992 5136
rect 13026 5102 13036 5136
rect 12982 5068 13036 5102
rect 12982 5034 12992 5068
rect 13026 5034 13036 5068
rect 12982 5018 13036 5034
rect 13066 5068 13120 5148
rect 13066 5034 13076 5068
rect 13110 5034 13120 5068
rect 13066 5018 13120 5034
rect 13150 5136 13204 5148
rect 13150 5102 13160 5136
rect 13194 5102 13204 5136
rect 13150 5068 13204 5102
rect 13150 5034 13160 5068
rect 13194 5034 13204 5068
rect 13150 5018 13204 5034
rect 13234 5068 13288 5148
rect 13234 5034 13244 5068
rect 13278 5034 13288 5068
rect 13234 5018 13288 5034
rect 13318 5136 13372 5148
rect 13318 5102 13328 5136
rect 13362 5102 13372 5136
rect 13318 5068 13372 5102
rect 13318 5034 13328 5068
rect 13362 5034 13372 5068
rect 13318 5018 13372 5034
rect 13402 5068 13456 5148
rect 13402 5034 13412 5068
rect 13446 5034 13456 5068
rect 13402 5018 13456 5034
rect 13486 5136 13540 5148
rect 13486 5102 13496 5136
rect 13530 5102 13540 5136
rect 13486 5068 13540 5102
rect 13486 5034 13496 5068
rect 13530 5034 13540 5068
rect 13486 5018 13540 5034
rect 13570 5068 13624 5148
rect 13570 5034 13580 5068
rect 13614 5034 13624 5068
rect 13570 5018 13624 5034
rect 13654 5136 13708 5148
rect 13654 5102 13664 5136
rect 13698 5102 13708 5136
rect 13654 5068 13708 5102
rect 13654 5034 13664 5068
rect 13698 5034 13708 5068
rect 13654 5018 13708 5034
rect 13738 5068 13790 5148
rect 13738 5034 13748 5068
rect 13782 5034 13790 5068
rect 13738 5018 13790 5034
rect 13916 5100 13968 5148
rect 13916 5066 13924 5100
rect 13958 5066 13968 5100
rect 13916 5018 13968 5066
rect 13998 5102 14048 5148
rect 13998 5064 14063 5102
rect 13998 5030 14008 5064
rect 14042 5030 14063 5064
rect 13998 5018 14063 5030
rect 14093 5090 14145 5102
rect 14093 5056 14103 5090
rect 14137 5056 14145 5090
rect 14093 5018 14145 5056
rect 14199 5098 14251 5148
rect 14199 5064 14207 5098
rect 14241 5064 14251 5098
rect 14199 5018 14251 5064
rect 14281 5102 14331 5148
rect 14281 5064 14346 5102
rect 14281 5030 14291 5064
rect 14325 5030 14346 5064
rect 14281 5018 14346 5030
rect 14376 5074 14428 5102
rect 14376 5040 14386 5074
rect 14420 5040 14428 5074
rect 14376 5018 14428 5040
rect 14482 5072 14534 5146
rect 14482 5038 14490 5072
rect 14524 5038 14534 5072
rect 14482 5018 14534 5038
rect 14564 5124 14618 5146
rect 14564 5090 14574 5124
rect 14608 5090 14618 5124
rect 14564 5018 14618 5090
rect 14648 5102 14698 5146
rect 14648 5080 14736 5102
rect 14648 5046 14674 5080
rect 14708 5046 14736 5080
rect 14648 5018 14736 5046
rect 14766 5060 14822 5102
rect 14766 5026 14776 5060
rect 14810 5026 14822 5060
rect 14766 5018 14822 5026
rect 14852 5090 14902 5102
rect 15071 5090 15121 5146
rect 14852 5018 14917 5090
rect 14947 5064 15026 5090
rect 14947 5030 14967 5064
rect 15001 5030 15026 5064
rect 14947 5018 15026 5030
rect 15056 5018 15121 5090
rect 15151 5064 15203 5146
rect 15151 5030 15161 5064
rect 15195 5030 15203 5064
rect 15151 5018 15203 5030
rect 15257 5098 15309 5146
rect 15257 5064 15265 5098
rect 15299 5064 15309 5098
rect 15257 5018 15309 5064
rect 15339 5124 15393 5146
rect 15339 5090 15349 5124
rect 15383 5090 15393 5124
rect 15339 5018 15393 5090
rect 15423 5102 15473 5146
rect 15423 5080 15493 5102
rect 15423 5046 15449 5080
rect 15483 5046 15493 5080
rect 15423 5018 15493 5046
rect 15523 5060 15603 5102
rect 15523 5026 15533 5060
rect 15567 5026 15603 5060
rect 15523 5018 15603 5026
rect 15633 5090 15684 5102
rect 15850 5090 15900 5102
rect 15633 5018 15699 5090
rect 15729 5064 15805 5090
rect 15729 5030 15750 5064
rect 15784 5030 15805 5064
rect 15729 5018 15805 5030
rect 15835 5082 15900 5090
rect 15835 5048 15856 5082
rect 15890 5048 15900 5082
rect 15835 5018 15900 5048
rect 15930 5064 15982 5102
rect 15930 5030 15940 5064
rect 15974 5030 15982 5064
rect 15930 5018 15982 5030
rect 16036 5090 16088 5102
rect 16036 5056 16044 5090
rect 16078 5056 16088 5090
rect 16036 5018 16088 5056
rect 16118 5064 16172 5102
rect 16118 5030 16128 5064
rect 16162 5030 16172 5064
rect 16118 5018 16172 5030
rect 16202 5090 16254 5102
rect 16202 5056 16212 5090
rect 16246 5056 16254 5090
rect 16202 5018 16254 5056
rect 16308 5100 16360 5148
rect 16308 5066 16316 5100
rect 16350 5066 16360 5100
rect 16308 5018 16360 5066
rect 16390 5102 16440 5148
rect 16390 5064 16455 5102
rect 16390 5030 16400 5064
rect 16434 5030 16455 5064
rect 16390 5018 16455 5030
rect 16485 5090 16537 5102
rect 16485 5056 16495 5090
rect 16529 5056 16537 5090
rect 16485 5018 16537 5056
rect 16591 5098 16643 5148
rect 16591 5064 16599 5098
rect 16633 5064 16643 5098
rect 16591 5018 16643 5064
rect 16673 5102 16723 5148
rect 16673 5064 16738 5102
rect 16673 5030 16683 5064
rect 16717 5030 16738 5064
rect 16673 5018 16738 5030
rect 16768 5074 16820 5102
rect 16768 5040 16778 5074
rect 16812 5040 16820 5074
rect 16768 5018 16820 5040
rect 16874 5072 16926 5146
rect 16874 5038 16882 5072
rect 16916 5038 16926 5072
rect 16874 5018 16926 5038
rect 16956 5124 17010 5146
rect 16956 5090 16966 5124
rect 17000 5090 17010 5124
rect 16956 5018 17010 5090
rect 17040 5102 17090 5146
rect 17040 5080 17128 5102
rect 17040 5046 17066 5080
rect 17100 5046 17128 5080
rect 17040 5018 17128 5046
rect 17158 5060 17214 5102
rect 17158 5026 17168 5060
rect 17202 5026 17214 5060
rect 17158 5018 17214 5026
rect 17244 5090 17294 5102
rect 17463 5090 17513 5146
rect 17244 5018 17309 5090
rect 17339 5064 17418 5090
rect 17339 5030 17359 5064
rect 17393 5030 17418 5064
rect 17339 5018 17418 5030
rect 17448 5018 17513 5090
rect 17543 5064 17595 5146
rect 17543 5030 17553 5064
rect 17587 5030 17595 5064
rect 17543 5018 17595 5030
rect 17649 5098 17701 5146
rect 17649 5064 17657 5098
rect 17691 5064 17701 5098
rect 17649 5018 17701 5064
rect 17731 5124 17785 5146
rect 17731 5090 17741 5124
rect 17775 5090 17785 5124
rect 17731 5018 17785 5090
rect 17815 5102 17865 5146
rect 17815 5080 17885 5102
rect 17815 5046 17841 5080
rect 17875 5046 17885 5080
rect 17815 5018 17885 5046
rect 17915 5060 17995 5102
rect 17915 5026 17925 5060
rect 17959 5026 17995 5060
rect 17915 5018 17995 5026
rect 18025 5090 18076 5102
rect 18242 5090 18292 5102
rect 18025 5018 18091 5090
rect 18121 5064 18197 5090
rect 18121 5030 18142 5064
rect 18176 5030 18197 5064
rect 18121 5018 18197 5030
rect 18227 5082 18292 5090
rect 18227 5048 18248 5082
rect 18282 5048 18292 5082
rect 18227 5018 18292 5048
rect 18322 5064 18374 5102
rect 18322 5030 18332 5064
rect 18366 5030 18374 5064
rect 18322 5018 18374 5030
rect 18428 5090 18480 5102
rect 18428 5056 18436 5090
rect 18470 5056 18480 5090
rect 18428 5018 18480 5056
rect 18510 5064 18564 5102
rect 18510 5030 18520 5064
rect 18554 5030 18564 5064
rect 18510 5018 18564 5030
rect 18594 5090 18646 5102
rect 18594 5056 18604 5090
rect 18638 5056 18646 5090
rect 18594 5018 18646 5056
rect 18700 5100 18752 5148
rect 18700 5066 18708 5100
rect 18742 5066 18752 5100
rect 18700 5018 18752 5066
rect 18782 5102 18832 5148
rect 18782 5064 18847 5102
rect 18782 5030 18792 5064
rect 18826 5030 18847 5064
rect 18782 5018 18847 5030
rect 18877 5090 18929 5102
rect 18877 5056 18887 5090
rect 18921 5056 18929 5090
rect 18877 5018 18929 5056
rect 18983 5098 19035 5148
rect 18983 5064 18991 5098
rect 19025 5064 19035 5098
rect 18983 5018 19035 5064
rect 19065 5102 19115 5148
rect 19065 5064 19130 5102
rect 19065 5030 19075 5064
rect 19109 5030 19130 5064
rect 19065 5018 19130 5030
rect 19160 5074 19212 5102
rect 19160 5040 19170 5074
rect 19204 5040 19212 5074
rect 19160 5018 19212 5040
rect 19266 5072 19318 5146
rect 19266 5038 19274 5072
rect 19308 5038 19318 5072
rect 19266 5018 19318 5038
rect 19348 5124 19402 5146
rect 19348 5090 19358 5124
rect 19392 5090 19402 5124
rect 19348 5018 19402 5090
rect 19432 5102 19482 5146
rect 19432 5080 19520 5102
rect 19432 5046 19458 5080
rect 19492 5046 19520 5080
rect 19432 5018 19520 5046
rect 19550 5060 19606 5102
rect 19550 5026 19560 5060
rect 19594 5026 19606 5060
rect 19550 5018 19606 5026
rect 19636 5090 19686 5102
rect 19855 5090 19905 5146
rect 19636 5018 19701 5090
rect 19731 5064 19810 5090
rect 19731 5030 19751 5064
rect 19785 5030 19810 5064
rect 19731 5018 19810 5030
rect 19840 5018 19905 5090
rect 19935 5064 19987 5146
rect 19935 5030 19945 5064
rect 19979 5030 19987 5064
rect 19935 5018 19987 5030
rect 20041 5098 20093 5146
rect 20041 5064 20049 5098
rect 20083 5064 20093 5098
rect 20041 5018 20093 5064
rect 20123 5124 20177 5146
rect 20123 5090 20133 5124
rect 20167 5090 20177 5124
rect 20123 5018 20177 5090
rect 20207 5102 20257 5146
rect 20207 5080 20277 5102
rect 20207 5046 20233 5080
rect 20267 5046 20277 5080
rect 20207 5018 20277 5046
rect 20307 5060 20387 5102
rect 20307 5026 20317 5060
rect 20351 5026 20387 5060
rect 20307 5018 20387 5026
rect 20417 5090 20468 5102
rect 20634 5090 20684 5102
rect 20417 5018 20483 5090
rect 20513 5064 20589 5090
rect 20513 5030 20534 5064
rect 20568 5030 20589 5064
rect 20513 5018 20589 5030
rect 20619 5082 20684 5090
rect 20619 5048 20640 5082
rect 20674 5048 20684 5082
rect 20619 5018 20684 5048
rect 20714 5064 20766 5102
rect 20714 5030 20724 5064
rect 20758 5030 20766 5064
rect 20714 5018 20766 5030
rect 20820 5090 20872 5102
rect 20820 5056 20828 5090
rect 20862 5056 20872 5090
rect 20820 5018 20872 5056
rect 20902 5064 20956 5102
rect 20902 5030 20912 5064
rect 20946 5030 20956 5064
rect 20902 5018 20956 5030
rect 20986 5090 21038 5102
rect 20986 5056 20996 5090
rect 21030 5056 21038 5090
rect 20986 5018 21038 5056
rect 21092 5100 21144 5148
rect 21092 5066 21100 5100
rect 21134 5066 21144 5100
rect 21092 5018 21144 5066
rect 21174 5102 21224 5148
rect 21174 5064 21239 5102
rect 21174 5030 21184 5064
rect 21218 5030 21239 5064
rect 21174 5018 21239 5030
rect 21269 5090 21321 5102
rect 21269 5056 21279 5090
rect 21313 5056 21321 5090
rect 21269 5018 21321 5056
rect 21375 5098 21427 5148
rect 21375 5064 21383 5098
rect 21417 5064 21427 5098
rect 21375 5018 21427 5064
rect 21457 5102 21507 5148
rect 21457 5064 21522 5102
rect 21457 5030 21467 5064
rect 21501 5030 21522 5064
rect 21457 5018 21522 5030
rect 21552 5074 21604 5102
rect 21552 5040 21562 5074
rect 21596 5040 21604 5074
rect 21552 5018 21604 5040
rect 21658 5072 21710 5146
rect 21658 5038 21666 5072
rect 21700 5038 21710 5072
rect 21658 5018 21710 5038
rect 21740 5124 21794 5146
rect 21740 5090 21750 5124
rect 21784 5090 21794 5124
rect 21740 5018 21794 5090
rect 21824 5102 21874 5146
rect 24504 5481 24562 5493
rect 21824 5080 21912 5102
rect 21824 5046 21850 5080
rect 21884 5046 21912 5080
rect 21824 5018 21912 5046
rect 21942 5060 21998 5102
rect 21942 5026 21952 5060
rect 21986 5026 21998 5060
rect 21942 5018 21998 5026
rect 22028 5090 22078 5102
rect 22247 5090 22297 5146
rect 22028 5018 22093 5090
rect 22123 5064 22202 5090
rect 22123 5030 22143 5064
rect 22177 5030 22202 5064
rect 22123 5018 22202 5030
rect 22232 5018 22297 5090
rect 22327 5064 22379 5146
rect 22327 5030 22337 5064
rect 22371 5030 22379 5064
rect 22327 5018 22379 5030
rect 22433 5098 22485 5146
rect 22433 5064 22441 5098
rect 22475 5064 22485 5098
rect 22433 5018 22485 5064
rect 22515 5124 22569 5146
rect 22515 5090 22525 5124
rect 22559 5090 22569 5124
rect 22515 5018 22569 5090
rect 22599 5102 22649 5146
rect 24504 5421 24516 5481
rect 24550 5421 24562 5481
rect 24504 5409 24562 5421
rect 24592 5409 24634 5493
rect 24664 5481 24722 5493
rect 24664 5421 24676 5481
rect 24710 5421 24722 5481
rect 24664 5409 24722 5421
rect 24504 5343 24562 5355
rect 24504 5283 24516 5343
rect 24550 5283 24562 5343
rect 24504 5271 24562 5283
rect 24592 5271 24634 5355
rect 24664 5343 24722 5355
rect 24664 5283 24676 5343
rect 24710 5283 24722 5343
rect 24664 5271 24722 5283
rect 22599 5080 22669 5102
rect 22599 5046 22625 5080
rect 22659 5046 22669 5080
rect 22599 5018 22669 5046
rect 22699 5060 22779 5102
rect 22699 5026 22709 5060
rect 22743 5026 22779 5060
rect 22699 5018 22779 5026
rect 22809 5090 22860 5102
rect 24504 5205 24562 5217
rect 24504 5145 24516 5205
rect 24550 5145 24562 5205
rect 24504 5133 24562 5145
rect 24592 5133 24634 5217
rect 24664 5205 24722 5217
rect 24664 5145 24676 5205
rect 24710 5145 24722 5205
rect 24664 5133 24722 5145
rect 23026 5090 23076 5102
rect 22809 5018 22875 5090
rect 22905 5064 22981 5090
rect 22905 5030 22926 5064
rect 22960 5030 22981 5064
rect 22905 5018 22981 5030
rect 23011 5082 23076 5090
rect 23011 5048 23032 5082
rect 23066 5048 23076 5082
rect 23011 5018 23076 5048
rect 23106 5064 23158 5102
rect 23106 5030 23116 5064
rect 23150 5030 23158 5064
rect 23106 5018 23158 5030
rect 23212 5090 23264 5102
rect 23212 5056 23220 5090
rect 23254 5056 23264 5090
rect 23212 5018 23264 5056
rect 23294 5064 23348 5102
rect 23294 5030 23304 5064
rect 23338 5030 23348 5064
rect 23294 5018 23348 5030
rect 23378 5090 23430 5102
rect 23378 5056 23388 5090
rect 23422 5056 23430 5090
rect 23378 5018 23430 5056
rect 24504 5067 24562 5079
rect 24504 5007 24516 5067
rect 24550 5007 24562 5067
rect 24504 4995 24562 5007
rect 24592 4995 24634 5079
rect 24664 5067 24722 5079
rect 24664 5007 24676 5067
rect 24710 5007 24722 5067
rect 24664 4995 24722 5007
rect 24504 4929 24562 4941
rect 24504 4869 24516 4929
rect 24550 4869 24562 4929
rect 24504 4857 24562 4869
rect 24592 4857 24634 4941
rect 24664 4929 24722 4941
rect 24664 4869 24676 4929
rect 24710 4869 24722 4929
rect 24664 4857 24722 4869
rect 24504 4791 24562 4803
rect 24504 4731 24516 4791
rect 24550 4731 24562 4791
rect 24504 4719 24562 4731
rect 24592 4719 24634 4803
rect 24664 4791 24722 4803
rect 24664 4731 24676 4791
rect 24710 4731 24722 4791
rect 24664 4719 24722 4731
rect 11116 4203 11168 4248
rect 11116 4169 11124 4203
rect 11158 4169 11168 4203
rect 11116 4144 11168 4169
rect 11198 4190 11256 4248
rect 11198 4156 11210 4190
rect 11244 4156 11256 4190
rect 11198 4144 11256 4156
rect 11286 4220 11338 4248
rect 11286 4186 11296 4220
rect 11330 4186 11338 4220
rect 11286 4144 11338 4186
rect 11392 4226 11444 4274
rect 11392 4192 11400 4226
rect 11434 4192 11444 4226
rect 11392 4144 11444 4192
rect 11474 4194 11528 4274
rect 11474 4160 11484 4194
rect 11518 4160 11528 4194
rect 11474 4144 11528 4160
rect 11558 4226 11612 4274
rect 11558 4192 11568 4226
rect 11602 4192 11612 4226
rect 11558 4144 11612 4192
rect 11642 4194 11696 4274
rect 11642 4160 11652 4194
rect 11686 4160 11696 4194
rect 11642 4144 11696 4160
rect 11726 4226 11780 4274
rect 11726 4192 11736 4226
rect 11770 4192 11780 4226
rect 11726 4144 11780 4192
rect 11810 4258 11862 4274
rect 11810 4224 11820 4258
rect 11854 4224 11862 4258
rect 11810 4190 11862 4224
rect 11810 4156 11820 4190
rect 11854 4156 11862 4190
rect 11810 4144 11862 4156
rect 13699 4263 13751 4275
rect 13699 4229 13707 4263
rect 13741 4229 13751 4263
rect 13699 4195 13751 4229
rect 13699 4161 13707 4195
rect 13741 4161 13751 4195
rect 13699 4145 13751 4161
rect 13781 4263 13833 4275
rect 13781 4229 13791 4263
rect 13825 4229 13833 4263
rect 13781 4195 13833 4229
rect 13781 4161 13791 4195
rect 13825 4161 13833 4195
rect 13781 4145 13833 4161
rect 13915 4217 13967 4229
rect 13915 4183 13923 4217
rect 13957 4183 13967 4217
rect 13915 4145 13967 4183
rect 13997 4191 14051 4229
rect 13997 4157 14007 4191
rect 14041 4157 14051 4191
rect 13997 4145 14051 4157
rect 14081 4217 14133 4229
rect 14081 4183 14091 4217
rect 14125 4183 14133 4217
rect 14081 4145 14133 4183
rect 14187 4191 14239 4229
rect 14187 4157 14195 4191
rect 14229 4157 14239 4191
rect 14187 4145 14239 4157
rect 14269 4217 14319 4229
rect 14696 4229 14746 4273
rect 14485 4217 14536 4229
rect 14269 4209 14334 4217
rect 14269 4175 14279 4209
rect 14313 4175 14334 4209
rect 14269 4145 14334 4175
rect 14364 4191 14440 4217
rect 14364 4157 14385 4191
rect 14419 4157 14440 4191
rect 14364 4145 14440 4157
rect 14470 4145 14536 4217
rect 14566 4187 14646 4229
rect 14566 4153 14602 4187
rect 14636 4153 14646 4187
rect 14566 4145 14646 4153
rect 14676 4207 14746 4229
rect 14676 4173 14686 4207
rect 14720 4173 14746 4207
rect 14676 4145 14746 4173
rect 14776 4251 14830 4273
rect 14776 4217 14786 4251
rect 14820 4217 14830 4251
rect 14776 4145 14830 4217
rect 14860 4225 14912 4273
rect 14860 4191 14870 4225
rect 14904 4191 14912 4225
rect 14860 4145 14912 4191
rect 14966 4191 15018 4273
rect 14966 4157 14974 4191
rect 15008 4157 15018 4191
rect 14966 4145 15018 4157
rect 15048 4217 15098 4273
rect 15471 4229 15521 4273
rect 15267 4217 15317 4229
rect 15048 4145 15113 4217
rect 15143 4191 15222 4217
rect 15143 4157 15168 4191
rect 15202 4157 15222 4191
rect 15143 4145 15222 4157
rect 15252 4145 15317 4217
rect 15347 4187 15403 4229
rect 15347 4153 15359 4187
rect 15393 4153 15403 4187
rect 15347 4145 15403 4153
rect 15433 4207 15521 4229
rect 15433 4173 15461 4207
rect 15495 4173 15521 4207
rect 15433 4145 15521 4173
rect 15551 4251 15605 4273
rect 15551 4217 15561 4251
rect 15595 4217 15605 4251
rect 15551 4145 15605 4217
rect 15635 4199 15687 4273
rect 15838 4229 15888 4275
rect 15635 4165 15645 4199
rect 15679 4165 15687 4199
rect 15635 4145 15687 4165
rect 15741 4201 15793 4229
rect 15741 4167 15749 4201
rect 15783 4167 15793 4201
rect 15741 4145 15793 4167
rect 15823 4191 15888 4229
rect 15823 4157 15844 4191
rect 15878 4157 15888 4191
rect 15823 4145 15888 4157
rect 15918 4225 15970 4275
rect 16121 4229 16171 4275
rect 15918 4191 15928 4225
rect 15962 4191 15970 4225
rect 15918 4145 15970 4191
rect 16024 4217 16076 4229
rect 16024 4183 16032 4217
rect 16066 4183 16076 4217
rect 16024 4145 16076 4183
rect 16106 4191 16171 4229
rect 16106 4157 16127 4191
rect 16161 4157 16171 4191
rect 16106 4145 16171 4157
rect 16201 4227 16253 4275
rect 16201 4193 16211 4227
rect 16245 4193 16253 4227
rect 16201 4145 16253 4193
rect 16307 4217 16359 4229
rect 16307 4183 16315 4217
rect 16349 4183 16359 4217
rect 16307 4145 16359 4183
rect 16389 4191 16443 4229
rect 16389 4157 16399 4191
rect 16433 4157 16443 4191
rect 16389 4145 16443 4157
rect 16473 4217 16525 4229
rect 16473 4183 16483 4217
rect 16517 4183 16525 4217
rect 16473 4145 16525 4183
rect 16579 4191 16631 4229
rect 16579 4157 16587 4191
rect 16621 4157 16631 4191
rect 16579 4145 16631 4157
rect 16661 4217 16711 4229
rect 17088 4229 17138 4273
rect 16877 4217 16928 4229
rect 16661 4209 16726 4217
rect 16661 4175 16671 4209
rect 16705 4175 16726 4209
rect 16661 4145 16726 4175
rect 16756 4191 16832 4217
rect 16756 4157 16777 4191
rect 16811 4157 16832 4191
rect 16756 4145 16832 4157
rect 16862 4145 16928 4217
rect 16958 4187 17038 4229
rect 16958 4153 16994 4187
rect 17028 4153 17038 4187
rect 16958 4145 17038 4153
rect 17068 4207 17138 4229
rect 17068 4173 17078 4207
rect 17112 4173 17138 4207
rect 17068 4145 17138 4173
rect 17168 4251 17222 4273
rect 17168 4217 17178 4251
rect 17212 4217 17222 4251
rect 17168 4145 17222 4217
rect 17252 4225 17304 4273
rect 17252 4191 17262 4225
rect 17296 4191 17304 4225
rect 17252 4145 17304 4191
rect 17358 4191 17410 4273
rect 17358 4157 17366 4191
rect 17400 4157 17410 4191
rect 17358 4145 17410 4157
rect 17440 4217 17490 4273
rect 17863 4229 17913 4273
rect 17659 4217 17709 4229
rect 17440 4145 17505 4217
rect 17535 4191 17614 4217
rect 17535 4157 17560 4191
rect 17594 4157 17614 4191
rect 17535 4145 17614 4157
rect 17644 4145 17709 4217
rect 17739 4187 17795 4229
rect 17739 4153 17751 4187
rect 17785 4153 17795 4187
rect 17739 4145 17795 4153
rect 17825 4207 17913 4229
rect 17825 4173 17853 4207
rect 17887 4173 17913 4207
rect 17825 4145 17913 4173
rect 17943 4251 17997 4273
rect 17943 4217 17953 4251
rect 17987 4217 17997 4251
rect 17943 4145 17997 4217
rect 18027 4199 18079 4273
rect 18230 4229 18280 4275
rect 18027 4165 18037 4199
rect 18071 4165 18079 4199
rect 18027 4145 18079 4165
rect 18133 4201 18185 4229
rect 18133 4167 18141 4201
rect 18175 4167 18185 4201
rect 18133 4145 18185 4167
rect 18215 4191 18280 4229
rect 18215 4157 18236 4191
rect 18270 4157 18280 4191
rect 18215 4145 18280 4157
rect 18310 4225 18362 4275
rect 18513 4229 18563 4275
rect 18310 4191 18320 4225
rect 18354 4191 18362 4225
rect 18310 4145 18362 4191
rect 18416 4217 18468 4229
rect 18416 4183 18424 4217
rect 18458 4183 18468 4217
rect 18416 4145 18468 4183
rect 18498 4191 18563 4229
rect 18498 4157 18519 4191
rect 18553 4157 18563 4191
rect 18498 4145 18563 4157
rect 18593 4227 18645 4275
rect 18593 4193 18603 4227
rect 18637 4193 18645 4227
rect 18593 4145 18645 4193
rect 18699 4217 18751 4229
rect 18699 4183 18707 4217
rect 18741 4183 18751 4217
rect 18699 4145 18751 4183
rect 18781 4191 18835 4229
rect 18781 4157 18791 4191
rect 18825 4157 18835 4191
rect 18781 4145 18835 4157
rect 18865 4217 18917 4229
rect 18865 4183 18875 4217
rect 18909 4183 18917 4217
rect 18865 4145 18917 4183
rect 18971 4191 19023 4229
rect 18971 4157 18979 4191
rect 19013 4157 19023 4191
rect 18971 4145 19023 4157
rect 19053 4217 19103 4229
rect 19480 4229 19530 4273
rect 19269 4217 19320 4229
rect 19053 4209 19118 4217
rect 19053 4175 19063 4209
rect 19097 4175 19118 4209
rect 19053 4145 19118 4175
rect 19148 4191 19224 4217
rect 19148 4157 19169 4191
rect 19203 4157 19224 4191
rect 19148 4145 19224 4157
rect 19254 4145 19320 4217
rect 19350 4187 19430 4229
rect 19350 4153 19386 4187
rect 19420 4153 19430 4187
rect 19350 4145 19430 4153
rect 19460 4207 19530 4229
rect 19460 4173 19470 4207
rect 19504 4173 19530 4207
rect 19460 4145 19530 4173
rect 19560 4251 19614 4273
rect 19560 4217 19570 4251
rect 19604 4217 19614 4251
rect 19560 4145 19614 4217
rect 19644 4225 19696 4273
rect 19644 4191 19654 4225
rect 19688 4191 19696 4225
rect 19644 4145 19696 4191
rect 19750 4191 19802 4273
rect 19750 4157 19758 4191
rect 19792 4157 19802 4191
rect 19750 4145 19802 4157
rect 19832 4217 19882 4273
rect 20255 4229 20305 4273
rect 20051 4217 20101 4229
rect 19832 4145 19897 4217
rect 19927 4191 20006 4217
rect 19927 4157 19952 4191
rect 19986 4157 20006 4191
rect 19927 4145 20006 4157
rect 20036 4145 20101 4217
rect 20131 4187 20187 4229
rect 20131 4153 20143 4187
rect 20177 4153 20187 4187
rect 20131 4145 20187 4153
rect 20217 4207 20305 4229
rect 20217 4173 20245 4207
rect 20279 4173 20305 4207
rect 20217 4145 20305 4173
rect 20335 4251 20389 4273
rect 20335 4217 20345 4251
rect 20379 4217 20389 4251
rect 20335 4145 20389 4217
rect 20419 4199 20471 4273
rect 20622 4229 20672 4275
rect 20419 4165 20429 4199
rect 20463 4165 20471 4199
rect 20419 4145 20471 4165
rect 20525 4201 20577 4229
rect 20525 4167 20533 4201
rect 20567 4167 20577 4201
rect 20525 4145 20577 4167
rect 20607 4191 20672 4229
rect 20607 4157 20628 4191
rect 20662 4157 20672 4191
rect 20607 4145 20672 4157
rect 20702 4225 20754 4275
rect 20905 4229 20955 4275
rect 20702 4191 20712 4225
rect 20746 4191 20754 4225
rect 20702 4145 20754 4191
rect 20808 4217 20860 4229
rect 20808 4183 20816 4217
rect 20850 4183 20860 4217
rect 20808 4145 20860 4183
rect 20890 4191 20955 4229
rect 20890 4157 20911 4191
rect 20945 4157 20955 4191
rect 20890 4145 20955 4157
rect 20985 4227 21037 4275
rect 20985 4193 20995 4227
rect 21029 4193 21037 4227
rect 20985 4145 21037 4193
rect 21091 4217 21143 4229
rect 21091 4183 21099 4217
rect 21133 4183 21143 4217
rect 21091 4145 21143 4183
rect 21173 4191 21227 4229
rect 21173 4157 21183 4191
rect 21217 4157 21227 4191
rect 21173 4145 21227 4157
rect 21257 4217 21309 4229
rect 21257 4183 21267 4217
rect 21301 4183 21309 4217
rect 21257 4145 21309 4183
rect 21363 4191 21415 4229
rect 21363 4157 21371 4191
rect 21405 4157 21415 4191
rect 21363 4145 21415 4157
rect 21445 4217 21495 4229
rect 21872 4229 21922 4273
rect 21661 4217 21712 4229
rect 21445 4209 21510 4217
rect 21445 4175 21455 4209
rect 21489 4175 21510 4209
rect 21445 4145 21510 4175
rect 21540 4191 21616 4217
rect 21540 4157 21561 4191
rect 21595 4157 21616 4191
rect 21540 4145 21616 4157
rect 21646 4145 21712 4217
rect 21742 4187 21822 4229
rect 21742 4153 21778 4187
rect 21812 4153 21822 4187
rect 21742 4145 21822 4153
rect 21852 4207 21922 4229
rect 21852 4173 21862 4207
rect 21896 4173 21922 4207
rect 21852 4145 21922 4173
rect 21952 4251 22006 4273
rect 21952 4217 21962 4251
rect 21996 4217 22006 4251
rect 21952 4145 22006 4217
rect 22036 4225 22088 4273
rect 22036 4191 22046 4225
rect 22080 4191 22088 4225
rect 22036 4145 22088 4191
rect 22142 4191 22194 4273
rect 22142 4157 22150 4191
rect 22184 4157 22194 4191
rect 22142 4145 22194 4157
rect 22224 4217 22274 4273
rect 22647 4229 22697 4273
rect 22443 4217 22493 4229
rect 22224 4145 22289 4217
rect 22319 4191 22398 4217
rect 22319 4157 22344 4191
rect 22378 4157 22398 4191
rect 22319 4145 22398 4157
rect 22428 4145 22493 4217
rect 22523 4187 22579 4229
rect 22523 4153 22535 4187
rect 22569 4153 22579 4187
rect 22523 4145 22579 4153
rect 22609 4207 22697 4229
rect 22609 4173 22637 4207
rect 22671 4173 22697 4207
rect 22609 4145 22697 4173
rect 22727 4251 22781 4273
rect 22727 4217 22737 4251
rect 22771 4217 22781 4251
rect 22727 4145 22781 4217
rect 22811 4199 22863 4273
rect 23014 4229 23064 4275
rect 22811 4165 22821 4199
rect 22855 4165 22863 4199
rect 22811 4145 22863 4165
rect 22917 4201 22969 4229
rect 22917 4167 22925 4201
rect 22959 4167 22969 4201
rect 22917 4145 22969 4167
rect 22999 4191 23064 4229
rect 22999 4157 23020 4191
rect 23054 4157 23064 4191
rect 22999 4145 23064 4157
rect 23094 4225 23146 4275
rect 23297 4229 23347 4275
rect 23094 4191 23104 4225
rect 23138 4191 23146 4225
rect 23094 4145 23146 4191
rect 23200 4217 23252 4229
rect 23200 4183 23208 4217
rect 23242 4183 23252 4217
rect 23200 4145 23252 4183
rect 23282 4191 23347 4229
rect 23282 4157 23303 4191
rect 23337 4157 23347 4191
rect 23282 4145 23347 4157
rect 23377 4227 23429 4275
rect 23377 4193 23387 4227
rect 23421 4193 23429 4227
rect 23377 4145 23429 4193
rect 25604 4196 25656 4234
rect 25604 4162 25612 4196
rect 25646 4162 25656 4196
rect 25604 4150 25656 4162
rect 25686 4222 25740 4234
rect 25686 4188 25696 4222
rect 25730 4188 25740 4222
rect 25686 4150 25740 4188
rect 25770 4196 25822 4234
rect 25770 4162 25780 4196
rect 25814 4162 25822 4196
rect 25770 4150 25822 4162
rect 25876 4222 25928 4234
rect 25876 4188 25884 4222
rect 25918 4188 25928 4222
rect 25876 4150 25928 4188
rect 25958 4204 26023 4234
rect 25958 4170 25968 4204
rect 26002 4170 26023 4204
rect 25958 4162 26023 4170
rect 26053 4222 26129 4234
rect 26053 4188 26074 4222
rect 26108 4188 26129 4222
rect 26053 4162 26129 4188
rect 26159 4162 26225 4234
rect 25958 4150 26008 4162
rect 26174 4150 26225 4162
rect 26255 4226 26335 4234
rect 26255 4192 26291 4226
rect 26325 4192 26335 4226
rect 26255 4150 26335 4192
rect 26365 4206 26435 4234
rect 26365 4172 26375 4206
rect 26409 4172 26435 4206
rect 26365 4150 26435 4172
rect 26385 4106 26435 4150
rect 26465 4162 26519 4234
rect 26465 4128 26475 4162
rect 26509 4128 26519 4162
rect 26465 4106 26519 4128
rect 26549 4188 26601 4234
rect 26549 4154 26559 4188
rect 26593 4154 26601 4188
rect 26549 4106 26601 4154
rect 26655 4222 26707 4234
rect 26655 4188 26663 4222
rect 26697 4188 26707 4222
rect 26655 4106 26707 4188
rect 26737 4162 26802 4234
rect 26832 4222 26911 4234
rect 26832 4188 26857 4222
rect 26891 4188 26911 4222
rect 26832 4162 26911 4188
rect 26941 4162 27006 4234
rect 26737 4106 26787 4162
rect 26956 4150 27006 4162
rect 27036 4226 27092 4234
rect 27036 4192 27048 4226
rect 27082 4192 27092 4226
rect 27036 4150 27092 4192
rect 27122 4206 27210 4234
rect 27122 4172 27150 4206
rect 27184 4172 27210 4206
rect 27122 4150 27210 4172
rect 27160 4106 27210 4150
rect 27240 4162 27294 4234
rect 27240 4128 27250 4162
rect 27284 4128 27294 4162
rect 27240 4106 27294 4128
rect 27324 4214 27376 4234
rect 27324 4180 27334 4214
rect 27368 4180 27376 4214
rect 27324 4106 27376 4180
rect 27430 4212 27482 4234
rect 27430 4178 27438 4212
rect 27472 4178 27482 4212
rect 27430 4150 27482 4178
rect 27512 4222 27577 4234
rect 27512 4188 27533 4222
rect 27567 4188 27577 4222
rect 27512 4150 27577 4188
rect 27527 4104 27577 4150
rect 27607 4188 27659 4234
rect 27607 4154 27617 4188
rect 27651 4154 27659 4188
rect 27607 4104 27659 4154
rect 27713 4196 27765 4234
rect 27713 4162 27721 4196
rect 27755 4162 27765 4196
rect 27713 4150 27765 4162
rect 27795 4222 27860 4234
rect 27795 4188 27816 4222
rect 27850 4188 27860 4222
rect 27795 4150 27860 4188
rect 27810 4104 27860 4150
rect 27890 4186 27942 4234
rect 27890 4152 27900 4186
rect 27934 4152 27942 4186
rect 27890 4104 27942 4152
rect 27996 4196 28048 4234
rect 27996 4162 28004 4196
rect 28038 4162 28048 4196
rect 27996 4150 28048 4162
rect 28078 4222 28132 4234
rect 28078 4188 28088 4222
rect 28122 4188 28132 4222
rect 28078 4150 28132 4188
rect 28162 4196 28214 4234
rect 28162 4162 28172 4196
rect 28206 4162 28214 4196
rect 28162 4150 28214 4162
rect 28268 4222 28320 4234
rect 28268 4188 28276 4222
rect 28310 4188 28320 4222
rect 28268 4150 28320 4188
rect 28350 4204 28415 4234
rect 28350 4170 28360 4204
rect 28394 4170 28415 4204
rect 28350 4162 28415 4170
rect 28445 4222 28521 4234
rect 28445 4188 28466 4222
rect 28500 4188 28521 4222
rect 28445 4162 28521 4188
rect 28551 4162 28617 4234
rect 28350 4150 28400 4162
rect 28566 4150 28617 4162
rect 28647 4226 28727 4234
rect 28647 4192 28683 4226
rect 28717 4192 28727 4226
rect 28647 4150 28727 4192
rect 28757 4206 28827 4234
rect 28757 4172 28767 4206
rect 28801 4172 28827 4206
rect 28757 4150 28827 4172
rect 28777 4106 28827 4150
rect 28857 4162 28911 4234
rect 28857 4128 28867 4162
rect 28901 4128 28911 4162
rect 28857 4106 28911 4128
rect 28941 4188 28993 4234
rect 28941 4154 28951 4188
rect 28985 4154 28993 4188
rect 28941 4106 28993 4154
rect 29047 4222 29099 4234
rect 29047 4188 29055 4222
rect 29089 4188 29099 4222
rect 29047 4106 29099 4188
rect 29129 4162 29194 4234
rect 29224 4222 29303 4234
rect 29224 4188 29249 4222
rect 29283 4188 29303 4222
rect 29224 4162 29303 4188
rect 29333 4162 29398 4234
rect 29129 4106 29179 4162
rect 29348 4150 29398 4162
rect 29428 4226 29484 4234
rect 29428 4192 29440 4226
rect 29474 4192 29484 4226
rect 29428 4150 29484 4192
rect 29514 4206 29602 4234
rect 29514 4172 29542 4206
rect 29576 4172 29602 4206
rect 29514 4150 29602 4172
rect 29552 4106 29602 4150
rect 29632 4162 29686 4234
rect 29632 4128 29642 4162
rect 29676 4128 29686 4162
rect 29632 4106 29686 4128
rect 29716 4214 29768 4234
rect 29716 4180 29726 4214
rect 29760 4180 29768 4214
rect 29716 4106 29768 4180
rect 29822 4212 29874 4234
rect 29822 4178 29830 4212
rect 29864 4178 29874 4212
rect 29822 4150 29874 4178
rect 29904 4222 29969 4234
rect 29904 4188 29925 4222
rect 29959 4188 29969 4222
rect 29904 4150 29969 4188
rect 29919 4104 29969 4150
rect 29999 4188 30051 4234
rect 29999 4154 30009 4188
rect 30043 4154 30051 4188
rect 29999 4104 30051 4154
rect 30105 4196 30157 4234
rect 30105 4162 30113 4196
rect 30147 4162 30157 4196
rect 30105 4150 30157 4162
rect 30187 4222 30252 4234
rect 30187 4188 30208 4222
rect 30242 4188 30252 4222
rect 30187 4150 30252 4188
rect 30202 4104 30252 4150
rect 30282 4186 30334 4234
rect 30282 4152 30292 4186
rect 30326 4152 30334 4186
rect 30282 4104 30334 4152
rect 11523 3354 11575 3402
rect 11523 3320 11531 3354
rect 11565 3320 11575 3354
rect 11523 3272 11575 3320
rect 11605 3356 11655 3402
rect 11605 3318 11670 3356
rect 11605 3284 11615 3318
rect 11649 3284 11670 3318
rect 11605 3272 11670 3284
rect 11700 3344 11752 3356
rect 11700 3310 11710 3344
rect 11744 3310 11752 3344
rect 11700 3272 11752 3310
rect 11806 3352 11858 3402
rect 11806 3318 11814 3352
rect 11848 3318 11858 3352
rect 11806 3272 11858 3318
rect 11888 3356 11938 3402
rect 11888 3318 11953 3356
rect 11888 3284 11898 3318
rect 11932 3284 11953 3318
rect 11888 3272 11953 3284
rect 11983 3328 12035 3356
rect 11983 3294 11993 3328
rect 12027 3294 12035 3328
rect 11983 3272 12035 3294
rect 12089 3326 12141 3400
rect 12089 3292 12097 3326
rect 12131 3292 12141 3326
rect 12089 3272 12141 3292
rect 12171 3378 12225 3400
rect 12171 3344 12181 3378
rect 12215 3344 12225 3378
rect 12171 3272 12225 3344
rect 12255 3356 12305 3400
rect 12255 3334 12343 3356
rect 12255 3300 12281 3334
rect 12315 3300 12343 3334
rect 12255 3272 12343 3300
rect 12373 3314 12429 3356
rect 12373 3280 12383 3314
rect 12417 3280 12429 3314
rect 12373 3272 12429 3280
rect 12459 3344 12509 3356
rect 12678 3344 12728 3400
rect 12459 3272 12524 3344
rect 12554 3318 12633 3344
rect 12554 3284 12574 3318
rect 12608 3284 12633 3318
rect 12554 3272 12633 3284
rect 12663 3272 12728 3344
rect 12758 3318 12810 3400
rect 12758 3284 12768 3318
rect 12802 3284 12810 3318
rect 12758 3272 12810 3284
rect 12864 3352 12916 3400
rect 12864 3318 12872 3352
rect 12906 3318 12916 3352
rect 12864 3272 12916 3318
rect 12946 3378 13000 3400
rect 12946 3344 12956 3378
rect 12990 3344 13000 3378
rect 12946 3272 13000 3344
rect 13030 3356 13080 3400
rect 13030 3334 13100 3356
rect 13030 3300 13056 3334
rect 13090 3300 13100 3334
rect 13030 3272 13100 3300
rect 13130 3314 13210 3356
rect 13130 3280 13140 3314
rect 13174 3280 13210 3314
rect 13130 3272 13210 3280
rect 13240 3344 13291 3356
rect 13457 3344 13507 3356
rect 13240 3272 13306 3344
rect 13336 3318 13412 3344
rect 13336 3284 13357 3318
rect 13391 3284 13412 3318
rect 13336 3272 13412 3284
rect 13442 3336 13507 3344
rect 13442 3302 13463 3336
rect 13497 3302 13507 3336
rect 13442 3272 13507 3302
rect 13537 3318 13589 3356
rect 13537 3284 13547 3318
rect 13581 3284 13589 3318
rect 13537 3272 13589 3284
rect 13643 3344 13695 3356
rect 13643 3310 13651 3344
rect 13685 3310 13695 3344
rect 13643 3272 13695 3310
rect 13725 3318 13779 3356
rect 13725 3284 13735 3318
rect 13769 3284 13779 3318
rect 13725 3272 13779 3284
rect 13809 3344 13861 3356
rect 13809 3310 13819 3344
rect 13853 3310 13861 3344
rect 13809 3272 13861 3310
rect 13915 3354 13967 3402
rect 13915 3320 13923 3354
rect 13957 3320 13967 3354
rect 13915 3272 13967 3320
rect 13997 3356 14047 3402
rect 13997 3318 14062 3356
rect 13997 3284 14007 3318
rect 14041 3284 14062 3318
rect 13997 3272 14062 3284
rect 14092 3344 14144 3356
rect 14092 3310 14102 3344
rect 14136 3310 14144 3344
rect 14092 3272 14144 3310
rect 14198 3352 14250 3402
rect 14198 3318 14206 3352
rect 14240 3318 14250 3352
rect 14198 3272 14250 3318
rect 14280 3356 14330 3402
rect 14280 3318 14345 3356
rect 14280 3284 14290 3318
rect 14324 3284 14345 3318
rect 14280 3272 14345 3284
rect 14375 3328 14427 3356
rect 14375 3294 14385 3328
rect 14419 3294 14427 3328
rect 14375 3272 14427 3294
rect 14481 3326 14533 3400
rect 14481 3292 14489 3326
rect 14523 3292 14533 3326
rect 14481 3272 14533 3292
rect 14563 3378 14617 3400
rect 14563 3344 14573 3378
rect 14607 3344 14617 3378
rect 14563 3272 14617 3344
rect 14647 3356 14697 3400
rect 14647 3334 14735 3356
rect 14647 3300 14673 3334
rect 14707 3300 14735 3334
rect 14647 3272 14735 3300
rect 14765 3314 14821 3356
rect 14765 3280 14775 3314
rect 14809 3280 14821 3314
rect 14765 3272 14821 3280
rect 14851 3344 14901 3356
rect 15070 3344 15120 3400
rect 14851 3272 14916 3344
rect 14946 3318 15025 3344
rect 14946 3284 14966 3318
rect 15000 3284 15025 3318
rect 14946 3272 15025 3284
rect 15055 3272 15120 3344
rect 15150 3318 15202 3400
rect 15150 3284 15160 3318
rect 15194 3284 15202 3318
rect 15150 3272 15202 3284
rect 15256 3352 15308 3400
rect 15256 3318 15264 3352
rect 15298 3318 15308 3352
rect 15256 3272 15308 3318
rect 15338 3378 15392 3400
rect 15338 3344 15348 3378
rect 15382 3344 15392 3378
rect 15338 3272 15392 3344
rect 15422 3356 15472 3400
rect 15422 3334 15492 3356
rect 15422 3300 15448 3334
rect 15482 3300 15492 3334
rect 15422 3272 15492 3300
rect 15522 3314 15602 3356
rect 15522 3280 15532 3314
rect 15566 3280 15602 3314
rect 15522 3272 15602 3280
rect 15632 3344 15683 3356
rect 15849 3344 15899 3356
rect 15632 3272 15698 3344
rect 15728 3318 15804 3344
rect 15728 3284 15749 3318
rect 15783 3284 15804 3318
rect 15728 3272 15804 3284
rect 15834 3336 15899 3344
rect 15834 3302 15855 3336
rect 15889 3302 15899 3336
rect 15834 3272 15899 3302
rect 15929 3318 15981 3356
rect 15929 3284 15939 3318
rect 15973 3284 15981 3318
rect 15929 3272 15981 3284
rect 16035 3344 16087 3356
rect 16035 3310 16043 3344
rect 16077 3310 16087 3344
rect 16035 3272 16087 3310
rect 16117 3318 16171 3356
rect 16117 3284 16127 3318
rect 16161 3284 16171 3318
rect 16117 3272 16171 3284
rect 16201 3344 16253 3356
rect 16201 3310 16211 3344
rect 16245 3310 16253 3344
rect 16201 3272 16253 3310
rect 16307 3354 16359 3402
rect 16307 3320 16315 3354
rect 16349 3320 16359 3354
rect 16307 3272 16359 3320
rect 16389 3356 16439 3402
rect 16389 3318 16454 3356
rect 16389 3284 16399 3318
rect 16433 3284 16454 3318
rect 16389 3272 16454 3284
rect 16484 3344 16536 3356
rect 16484 3310 16494 3344
rect 16528 3310 16536 3344
rect 16484 3272 16536 3310
rect 16590 3352 16642 3402
rect 16590 3318 16598 3352
rect 16632 3318 16642 3352
rect 16590 3272 16642 3318
rect 16672 3356 16722 3402
rect 16672 3318 16737 3356
rect 16672 3284 16682 3318
rect 16716 3284 16737 3318
rect 16672 3272 16737 3284
rect 16767 3328 16819 3356
rect 16767 3294 16777 3328
rect 16811 3294 16819 3328
rect 16767 3272 16819 3294
rect 16873 3326 16925 3400
rect 16873 3292 16881 3326
rect 16915 3292 16925 3326
rect 16873 3272 16925 3292
rect 16955 3378 17009 3400
rect 16955 3344 16965 3378
rect 16999 3344 17009 3378
rect 16955 3272 17009 3344
rect 17039 3356 17089 3400
rect 17039 3334 17127 3356
rect 17039 3300 17065 3334
rect 17099 3300 17127 3334
rect 17039 3272 17127 3300
rect 17157 3314 17213 3356
rect 17157 3280 17167 3314
rect 17201 3280 17213 3314
rect 17157 3272 17213 3280
rect 17243 3344 17293 3356
rect 17462 3344 17512 3400
rect 17243 3272 17308 3344
rect 17338 3318 17417 3344
rect 17338 3284 17358 3318
rect 17392 3284 17417 3318
rect 17338 3272 17417 3284
rect 17447 3272 17512 3344
rect 17542 3318 17594 3400
rect 17542 3284 17552 3318
rect 17586 3284 17594 3318
rect 17542 3272 17594 3284
rect 17648 3352 17700 3400
rect 17648 3318 17656 3352
rect 17690 3318 17700 3352
rect 17648 3272 17700 3318
rect 17730 3378 17784 3400
rect 17730 3344 17740 3378
rect 17774 3344 17784 3378
rect 17730 3272 17784 3344
rect 17814 3356 17864 3400
rect 17814 3334 17884 3356
rect 17814 3300 17840 3334
rect 17874 3300 17884 3334
rect 17814 3272 17884 3300
rect 17914 3314 17994 3356
rect 17914 3280 17924 3314
rect 17958 3280 17994 3314
rect 17914 3272 17994 3280
rect 18024 3344 18075 3356
rect 18241 3344 18291 3356
rect 18024 3272 18090 3344
rect 18120 3318 18196 3344
rect 18120 3284 18141 3318
rect 18175 3284 18196 3318
rect 18120 3272 18196 3284
rect 18226 3336 18291 3344
rect 18226 3302 18247 3336
rect 18281 3302 18291 3336
rect 18226 3272 18291 3302
rect 18321 3318 18373 3356
rect 18321 3284 18331 3318
rect 18365 3284 18373 3318
rect 18321 3272 18373 3284
rect 18427 3344 18479 3356
rect 18427 3310 18435 3344
rect 18469 3310 18479 3344
rect 18427 3272 18479 3310
rect 18509 3318 18563 3356
rect 18509 3284 18519 3318
rect 18553 3284 18563 3318
rect 18509 3272 18563 3284
rect 18593 3344 18645 3356
rect 18593 3310 18603 3344
rect 18637 3310 18645 3344
rect 18593 3272 18645 3310
rect 18699 3354 18751 3402
rect 18699 3320 18707 3354
rect 18741 3320 18751 3354
rect 18699 3272 18751 3320
rect 18781 3356 18831 3402
rect 18781 3318 18846 3356
rect 18781 3284 18791 3318
rect 18825 3284 18846 3318
rect 18781 3272 18846 3284
rect 18876 3344 18928 3356
rect 18876 3310 18886 3344
rect 18920 3310 18928 3344
rect 18876 3272 18928 3310
rect 18982 3352 19034 3402
rect 18982 3318 18990 3352
rect 19024 3318 19034 3352
rect 18982 3272 19034 3318
rect 19064 3356 19114 3402
rect 19064 3318 19129 3356
rect 19064 3284 19074 3318
rect 19108 3284 19129 3318
rect 19064 3272 19129 3284
rect 19159 3328 19211 3356
rect 19159 3294 19169 3328
rect 19203 3294 19211 3328
rect 19159 3272 19211 3294
rect 19265 3326 19317 3400
rect 19265 3292 19273 3326
rect 19307 3292 19317 3326
rect 19265 3272 19317 3292
rect 19347 3378 19401 3400
rect 19347 3344 19357 3378
rect 19391 3344 19401 3378
rect 19347 3272 19401 3344
rect 19431 3356 19481 3400
rect 19431 3334 19519 3356
rect 19431 3300 19457 3334
rect 19491 3300 19519 3334
rect 19431 3272 19519 3300
rect 19549 3314 19605 3356
rect 19549 3280 19559 3314
rect 19593 3280 19605 3314
rect 19549 3272 19605 3280
rect 19635 3344 19685 3356
rect 19854 3344 19904 3400
rect 19635 3272 19700 3344
rect 19730 3318 19809 3344
rect 19730 3284 19750 3318
rect 19784 3284 19809 3318
rect 19730 3272 19809 3284
rect 19839 3272 19904 3344
rect 19934 3318 19986 3400
rect 19934 3284 19944 3318
rect 19978 3284 19986 3318
rect 19934 3272 19986 3284
rect 20040 3352 20092 3400
rect 20040 3318 20048 3352
rect 20082 3318 20092 3352
rect 20040 3272 20092 3318
rect 20122 3378 20176 3400
rect 20122 3344 20132 3378
rect 20166 3344 20176 3378
rect 20122 3272 20176 3344
rect 20206 3356 20256 3400
rect 20206 3334 20276 3356
rect 20206 3300 20232 3334
rect 20266 3300 20276 3334
rect 20206 3272 20276 3300
rect 20306 3314 20386 3356
rect 20306 3280 20316 3314
rect 20350 3280 20386 3314
rect 20306 3272 20386 3280
rect 20416 3344 20467 3356
rect 20633 3344 20683 3356
rect 20416 3272 20482 3344
rect 20512 3318 20588 3344
rect 20512 3284 20533 3318
rect 20567 3284 20588 3318
rect 20512 3272 20588 3284
rect 20618 3336 20683 3344
rect 20618 3302 20639 3336
rect 20673 3302 20683 3336
rect 20618 3272 20683 3302
rect 20713 3318 20765 3356
rect 20713 3284 20723 3318
rect 20757 3284 20765 3318
rect 20713 3272 20765 3284
rect 20819 3344 20871 3356
rect 20819 3310 20827 3344
rect 20861 3310 20871 3344
rect 20819 3272 20871 3310
rect 20901 3318 20955 3356
rect 20901 3284 20911 3318
rect 20945 3284 20955 3318
rect 20901 3272 20955 3284
rect 20985 3344 21037 3356
rect 20985 3310 20995 3344
rect 21029 3310 21037 3344
rect 20985 3272 21037 3310
rect 21091 3354 21143 3402
rect 21091 3320 21099 3354
rect 21133 3320 21143 3354
rect 21091 3272 21143 3320
rect 21173 3356 21223 3402
rect 21173 3318 21238 3356
rect 21173 3284 21183 3318
rect 21217 3284 21238 3318
rect 21173 3272 21238 3284
rect 21268 3344 21320 3356
rect 21268 3310 21278 3344
rect 21312 3310 21320 3344
rect 21268 3272 21320 3310
rect 21374 3352 21426 3402
rect 21374 3318 21382 3352
rect 21416 3318 21426 3352
rect 21374 3272 21426 3318
rect 21456 3356 21506 3402
rect 21456 3318 21521 3356
rect 21456 3284 21466 3318
rect 21500 3284 21521 3318
rect 21456 3272 21521 3284
rect 21551 3328 21603 3356
rect 21551 3294 21561 3328
rect 21595 3294 21603 3328
rect 21551 3272 21603 3294
rect 21657 3326 21709 3400
rect 21657 3292 21665 3326
rect 21699 3292 21709 3326
rect 21657 3272 21709 3292
rect 21739 3378 21793 3400
rect 21739 3344 21749 3378
rect 21783 3344 21793 3378
rect 21739 3272 21793 3344
rect 21823 3356 21873 3400
rect 21823 3334 21911 3356
rect 21823 3300 21849 3334
rect 21883 3300 21911 3334
rect 21823 3272 21911 3300
rect 21941 3314 21997 3356
rect 21941 3280 21951 3314
rect 21985 3280 21997 3314
rect 21941 3272 21997 3280
rect 22027 3344 22077 3356
rect 22246 3344 22296 3400
rect 22027 3272 22092 3344
rect 22122 3318 22201 3344
rect 22122 3284 22142 3318
rect 22176 3284 22201 3318
rect 22122 3272 22201 3284
rect 22231 3272 22296 3344
rect 22326 3318 22378 3400
rect 22326 3284 22336 3318
rect 22370 3284 22378 3318
rect 22326 3272 22378 3284
rect 22432 3352 22484 3400
rect 22432 3318 22440 3352
rect 22474 3318 22484 3352
rect 22432 3272 22484 3318
rect 22514 3378 22568 3400
rect 22514 3344 22524 3378
rect 22558 3344 22568 3378
rect 22514 3272 22568 3344
rect 22598 3356 22648 3400
rect 22598 3334 22668 3356
rect 22598 3300 22624 3334
rect 22658 3300 22668 3334
rect 22598 3272 22668 3300
rect 22698 3314 22778 3356
rect 22698 3280 22708 3314
rect 22742 3280 22778 3314
rect 22698 3272 22778 3280
rect 22808 3344 22859 3356
rect 23025 3344 23075 3356
rect 22808 3272 22874 3344
rect 22904 3318 22980 3344
rect 22904 3284 22925 3318
rect 22959 3284 22980 3318
rect 22904 3272 22980 3284
rect 23010 3336 23075 3344
rect 23010 3302 23031 3336
rect 23065 3302 23075 3336
rect 23010 3272 23075 3302
rect 23105 3318 23157 3356
rect 23105 3284 23115 3318
rect 23149 3284 23157 3318
rect 23105 3272 23157 3284
rect 23211 3344 23263 3356
rect 23211 3310 23219 3344
rect 23253 3310 23263 3344
rect 23211 3272 23263 3310
rect 23293 3318 23347 3356
rect 23293 3284 23303 3318
rect 23337 3284 23347 3318
rect 23293 3272 23347 3284
rect 23377 3344 23429 3356
rect 23377 3310 23387 3344
rect 23421 3310 23429 3344
rect 23377 3272 23429 3310
rect 25604 3216 25656 3228
rect 25604 3182 25612 3216
rect 25646 3182 25656 3216
rect 25604 3144 25656 3182
rect 25686 3190 25740 3228
rect 25686 3156 25696 3190
rect 25730 3156 25740 3190
rect 25686 3144 25740 3156
rect 25770 3216 25822 3228
rect 25770 3182 25780 3216
rect 25814 3182 25822 3216
rect 25770 3144 25822 3182
rect 25876 3190 25928 3228
rect 25876 3156 25884 3190
rect 25918 3156 25928 3190
rect 25876 3144 25928 3156
rect 25958 3216 26008 3228
rect 26385 3228 26435 3272
rect 26174 3216 26225 3228
rect 25958 3208 26023 3216
rect 25958 3174 25968 3208
rect 26002 3174 26023 3208
rect 25958 3144 26023 3174
rect 26053 3190 26129 3216
rect 26053 3156 26074 3190
rect 26108 3156 26129 3190
rect 26053 3144 26129 3156
rect 26159 3144 26225 3216
rect 26255 3186 26335 3228
rect 26255 3152 26291 3186
rect 26325 3152 26335 3186
rect 26255 3144 26335 3152
rect 26365 3206 26435 3228
rect 26365 3172 26375 3206
rect 26409 3172 26435 3206
rect 26365 3144 26435 3172
rect 26465 3250 26519 3272
rect 26465 3216 26475 3250
rect 26509 3216 26519 3250
rect 26465 3144 26519 3216
rect 26549 3224 26601 3272
rect 26549 3190 26559 3224
rect 26593 3190 26601 3224
rect 26549 3144 26601 3190
rect 26655 3190 26707 3272
rect 26655 3156 26663 3190
rect 26697 3156 26707 3190
rect 26655 3144 26707 3156
rect 26737 3216 26787 3272
rect 27160 3228 27210 3272
rect 26956 3216 27006 3228
rect 26737 3144 26802 3216
rect 26832 3190 26911 3216
rect 26832 3156 26857 3190
rect 26891 3156 26911 3190
rect 26832 3144 26911 3156
rect 26941 3144 27006 3216
rect 27036 3186 27092 3228
rect 27036 3152 27048 3186
rect 27082 3152 27092 3186
rect 27036 3144 27092 3152
rect 27122 3206 27210 3228
rect 27122 3172 27150 3206
rect 27184 3172 27210 3206
rect 27122 3144 27210 3172
rect 27240 3250 27294 3272
rect 27240 3216 27250 3250
rect 27284 3216 27294 3250
rect 27240 3144 27294 3216
rect 27324 3198 27376 3272
rect 27527 3228 27577 3274
rect 27324 3164 27334 3198
rect 27368 3164 27376 3198
rect 27324 3144 27376 3164
rect 27430 3200 27482 3228
rect 27430 3166 27438 3200
rect 27472 3166 27482 3200
rect 27430 3144 27482 3166
rect 27512 3190 27577 3228
rect 27512 3156 27533 3190
rect 27567 3156 27577 3190
rect 27512 3144 27577 3156
rect 27607 3224 27659 3274
rect 27810 3228 27860 3274
rect 27607 3190 27617 3224
rect 27651 3190 27659 3224
rect 27607 3144 27659 3190
rect 27713 3216 27765 3228
rect 27713 3182 27721 3216
rect 27755 3182 27765 3216
rect 27713 3144 27765 3182
rect 27795 3190 27860 3228
rect 27795 3156 27816 3190
rect 27850 3156 27860 3190
rect 27795 3144 27860 3156
rect 27890 3226 27942 3274
rect 27890 3192 27900 3226
rect 27934 3192 27942 3226
rect 27890 3144 27942 3192
rect 27996 3216 28048 3228
rect 27996 3182 28004 3216
rect 28038 3182 28048 3216
rect 27996 3144 28048 3182
rect 28078 3190 28132 3228
rect 28078 3156 28088 3190
rect 28122 3156 28132 3190
rect 28078 3144 28132 3156
rect 28162 3216 28214 3228
rect 28162 3182 28172 3216
rect 28206 3182 28214 3216
rect 28162 3144 28214 3182
rect 28268 3190 28320 3228
rect 28268 3156 28276 3190
rect 28310 3156 28320 3190
rect 28268 3144 28320 3156
rect 28350 3216 28400 3228
rect 28777 3228 28827 3272
rect 28566 3216 28617 3228
rect 28350 3208 28415 3216
rect 28350 3174 28360 3208
rect 28394 3174 28415 3208
rect 28350 3144 28415 3174
rect 28445 3190 28521 3216
rect 28445 3156 28466 3190
rect 28500 3156 28521 3190
rect 28445 3144 28521 3156
rect 28551 3144 28617 3216
rect 28647 3186 28727 3228
rect 28647 3152 28683 3186
rect 28717 3152 28727 3186
rect 28647 3144 28727 3152
rect 28757 3206 28827 3228
rect 28757 3172 28767 3206
rect 28801 3172 28827 3206
rect 28757 3144 28827 3172
rect 28857 3250 28911 3272
rect 28857 3216 28867 3250
rect 28901 3216 28911 3250
rect 28857 3144 28911 3216
rect 28941 3224 28993 3272
rect 28941 3190 28951 3224
rect 28985 3190 28993 3224
rect 28941 3144 28993 3190
rect 29047 3190 29099 3272
rect 29047 3156 29055 3190
rect 29089 3156 29099 3190
rect 29047 3144 29099 3156
rect 29129 3216 29179 3272
rect 29552 3228 29602 3272
rect 29348 3216 29398 3228
rect 29129 3144 29194 3216
rect 29224 3190 29303 3216
rect 29224 3156 29249 3190
rect 29283 3156 29303 3190
rect 29224 3144 29303 3156
rect 29333 3144 29398 3216
rect 29428 3186 29484 3228
rect 29428 3152 29440 3186
rect 29474 3152 29484 3186
rect 29428 3144 29484 3152
rect 29514 3206 29602 3228
rect 29514 3172 29542 3206
rect 29576 3172 29602 3206
rect 29514 3144 29602 3172
rect 29632 3250 29686 3272
rect 29632 3216 29642 3250
rect 29676 3216 29686 3250
rect 29632 3144 29686 3216
rect 29716 3198 29768 3272
rect 29919 3228 29969 3274
rect 29716 3164 29726 3198
rect 29760 3164 29768 3198
rect 29716 3144 29768 3164
rect 29822 3200 29874 3228
rect 29822 3166 29830 3200
rect 29864 3166 29874 3200
rect 29822 3144 29874 3166
rect 29904 3190 29969 3228
rect 29904 3156 29925 3190
rect 29959 3156 29969 3190
rect 29904 3144 29969 3156
rect 29999 3224 30051 3274
rect 30202 3228 30252 3274
rect 29999 3190 30009 3224
rect 30043 3190 30051 3224
rect 29999 3144 30051 3190
rect 30105 3216 30157 3228
rect 30105 3182 30113 3216
rect 30147 3182 30157 3216
rect 30105 3144 30157 3182
rect 30187 3190 30252 3228
rect 30187 3156 30208 3190
rect 30242 3156 30252 3190
rect 30187 3144 30252 3156
rect 30282 3226 30334 3274
rect 30282 3192 30292 3226
rect 30326 3192 30334 3226
rect 30282 3144 30334 3192
rect 25604 2916 25656 2954
rect 25604 2882 25612 2916
rect 25646 2882 25656 2916
rect 25604 2870 25656 2882
rect 25686 2942 25740 2954
rect 25686 2908 25696 2942
rect 25730 2908 25740 2942
rect 25686 2870 25740 2908
rect 25770 2916 25822 2954
rect 25770 2882 25780 2916
rect 25814 2882 25822 2916
rect 25770 2870 25822 2882
rect 25876 2942 25928 2954
rect 25876 2908 25884 2942
rect 25918 2908 25928 2942
rect 25876 2870 25928 2908
rect 25958 2924 26023 2954
rect 25958 2890 25968 2924
rect 26002 2890 26023 2924
rect 25958 2882 26023 2890
rect 26053 2942 26129 2954
rect 26053 2908 26074 2942
rect 26108 2908 26129 2942
rect 26053 2882 26129 2908
rect 26159 2882 26225 2954
rect 25958 2870 26008 2882
rect 26174 2870 26225 2882
rect 26255 2946 26335 2954
rect 26255 2912 26291 2946
rect 26325 2912 26335 2946
rect 26255 2870 26335 2912
rect 26365 2926 26435 2954
rect 26365 2892 26375 2926
rect 26409 2892 26435 2926
rect 26365 2870 26435 2892
rect 26385 2826 26435 2870
rect 26465 2882 26519 2954
rect 26465 2848 26475 2882
rect 26509 2848 26519 2882
rect 26465 2826 26519 2848
rect 26549 2908 26601 2954
rect 26549 2874 26559 2908
rect 26593 2874 26601 2908
rect 26549 2826 26601 2874
rect 26655 2942 26707 2954
rect 26655 2908 26663 2942
rect 26697 2908 26707 2942
rect 26655 2826 26707 2908
rect 26737 2882 26802 2954
rect 26832 2942 26911 2954
rect 26832 2908 26857 2942
rect 26891 2908 26911 2942
rect 26832 2882 26911 2908
rect 26941 2882 27006 2954
rect 26737 2826 26787 2882
rect 26956 2870 27006 2882
rect 27036 2946 27092 2954
rect 27036 2912 27048 2946
rect 27082 2912 27092 2946
rect 27036 2870 27092 2912
rect 27122 2926 27210 2954
rect 27122 2892 27150 2926
rect 27184 2892 27210 2926
rect 27122 2870 27210 2892
rect 27160 2826 27210 2870
rect 27240 2882 27294 2954
rect 27240 2848 27250 2882
rect 27284 2848 27294 2882
rect 27240 2826 27294 2848
rect 27324 2934 27376 2954
rect 27324 2900 27334 2934
rect 27368 2900 27376 2934
rect 27324 2826 27376 2900
rect 27430 2932 27482 2954
rect 27430 2898 27438 2932
rect 27472 2898 27482 2932
rect 27430 2870 27482 2898
rect 27512 2942 27577 2954
rect 27512 2908 27533 2942
rect 27567 2908 27577 2942
rect 27512 2870 27577 2908
rect 27527 2824 27577 2870
rect 27607 2908 27659 2954
rect 27607 2874 27617 2908
rect 27651 2874 27659 2908
rect 27607 2824 27659 2874
rect 27713 2916 27765 2954
rect 27713 2882 27721 2916
rect 27755 2882 27765 2916
rect 27713 2870 27765 2882
rect 27795 2942 27860 2954
rect 27795 2908 27816 2942
rect 27850 2908 27860 2942
rect 27795 2870 27860 2908
rect 27810 2824 27860 2870
rect 27890 2906 27942 2954
rect 27890 2872 27900 2906
rect 27934 2872 27942 2906
rect 27890 2824 27942 2872
rect 27996 2916 28048 2954
rect 27996 2882 28004 2916
rect 28038 2882 28048 2916
rect 27996 2870 28048 2882
rect 28078 2942 28132 2954
rect 28078 2908 28088 2942
rect 28122 2908 28132 2942
rect 28078 2870 28132 2908
rect 28162 2916 28214 2954
rect 28162 2882 28172 2916
rect 28206 2882 28214 2916
rect 28162 2870 28214 2882
rect 28268 2942 28320 2954
rect 28268 2908 28276 2942
rect 28310 2908 28320 2942
rect 28268 2870 28320 2908
rect 28350 2924 28415 2954
rect 28350 2890 28360 2924
rect 28394 2890 28415 2924
rect 28350 2882 28415 2890
rect 28445 2942 28521 2954
rect 28445 2908 28466 2942
rect 28500 2908 28521 2942
rect 28445 2882 28521 2908
rect 28551 2882 28617 2954
rect 28350 2870 28400 2882
rect 28566 2870 28617 2882
rect 28647 2946 28727 2954
rect 28647 2912 28683 2946
rect 28717 2912 28727 2946
rect 28647 2870 28727 2912
rect 28757 2926 28827 2954
rect 28757 2892 28767 2926
rect 28801 2892 28827 2926
rect 28757 2870 28827 2892
rect 28777 2826 28827 2870
rect 28857 2882 28911 2954
rect 28857 2848 28867 2882
rect 28901 2848 28911 2882
rect 28857 2826 28911 2848
rect 28941 2908 28993 2954
rect 28941 2874 28951 2908
rect 28985 2874 28993 2908
rect 28941 2826 28993 2874
rect 29047 2942 29099 2954
rect 29047 2908 29055 2942
rect 29089 2908 29099 2942
rect 29047 2826 29099 2908
rect 29129 2882 29194 2954
rect 29224 2942 29303 2954
rect 29224 2908 29249 2942
rect 29283 2908 29303 2942
rect 29224 2882 29303 2908
rect 29333 2882 29398 2954
rect 29129 2826 29179 2882
rect 29348 2870 29398 2882
rect 29428 2946 29484 2954
rect 29428 2912 29440 2946
rect 29474 2912 29484 2946
rect 29428 2870 29484 2912
rect 29514 2926 29602 2954
rect 29514 2892 29542 2926
rect 29576 2892 29602 2926
rect 29514 2870 29602 2892
rect 29552 2826 29602 2870
rect 29632 2882 29686 2954
rect 29632 2848 29642 2882
rect 29676 2848 29686 2882
rect 29632 2826 29686 2848
rect 29716 2934 29768 2954
rect 29716 2900 29726 2934
rect 29760 2900 29768 2934
rect 29716 2826 29768 2900
rect 29822 2932 29874 2954
rect 29822 2898 29830 2932
rect 29864 2898 29874 2932
rect 29822 2870 29874 2898
rect 29904 2942 29969 2954
rect 29904 2908 29925 2942
rect 29959 2908 29969 2942
rect 29904 2870 29969 2908
rect 29919 2824 29969 2870
rect 29999 2908 30051 2954
rect 29999 2874 30009 2908
rect 30043 2874 30051 2908
rect 29999 2824 30051 2874
rect 30105 2916 30157 2954
rect 30105 2882 30113 2916
rect 30147 2882 30157 2916
rect 30105 2870 30157 2882
rect 30187 2942 30252 2954
rect 30187 2908 30208 2942
rect 30242 2908 30252 2942
rect 30187 2870 30252 2908
rect 30202 2824 30252 2870
rect 30282 2906 30334 2954
rect 30282 2872 30292 2906
rect 30326 2872 30334 2906
rect 30282 2824 30334 2872
rect 25604 1936 25656 1948
rect 25604 1902 25612 1936
rect 25646 1902 25656 1936
rect 25604 1864 25656 1902
rect 25686 1910 25740 1948
rect 25686 1876 25696 1910
rect 25730 1876 25740 1910
rect 25686 1864 25740 1876
rect 25770 1936 25822 1948
rect 25770 1902 25780 1936
rect 25814 1902 25822 1936
rect 25770 1864 25822 1902
rect 25876 1910 25928 1948
rect 25876 1876 25884 1910
rect 25918 1876 25928 1910
rect 25876 1864 25928 1876
rect 25958 1936 26008 1948
rect 26385 1948 26435 1992
rect 26174 1936 26225 1948
rect 25958 1928 26023 1936
rect 25958 1894 25968 1928
rect 26002 1894 26023 1928
rect 25958 1864 26023 1894
rect 26053 1910 26129 1936
rect 26053 1876 26074 1910
rect 26108 1876 26129 1910
rect 26053 1864 26129 1876
rect 26159 1864 26225 1936
rect 26255 1906 26335 1948
rect 26255 1872 26291 1906
rect 26325 1872 26335 1906
rect 26255 1864 26335 1872
rect 26365 1926 26435 1948
rect 26365 1892 26375 1926
rect 26409 1892 26435 1926
rect 26365 1864 26435 1892
rect 26465 1970 26519 1992
rect 26465 1936 26475 1970
rect 26509 1936 26519 1970
rect 26465 1864 26519 1936
rect 26549 1944 26601 1992
rect 26549 1910 26559 1944
rect 26593 1910 26601 1944
rect 26549 1864 26601 1910
rect 26655 1910 26707 1992
rect 26655 1876 26663 1910
rect 26697 1876 26707 1910
rect 26655 1864 26707 1876
rect 26737 1936 26787 1992
rect 27160 1948 27210 1992
rect 26956 1936 27006 1948
rect 26737 1864 26802 1936
rect 26832 1910 26911 1936
rect 26832 1876 26857 1910
rect 26891 1876 26911 1910
rect 26832 1864 26911 1876
rect 26941 1864 27006 1936
rect 27036 1906 27092 1948
rect 27036 1872 27048 1906
rect 27082 1872 27092 1906
rect 27036 1864 27092 1872
rect 27122 1926 27210 1948
rect 27122 1892 27150 1926
rect 27184 1892 27210 1926
rect 27122 1864 27210 1892
rect 27240 1970 27294 1992
rect 27240 1936 27250 1970
rect 27284 1936 27294 1970
rect 27240 1864 27294 1936
rect 27324 1918 27376 1992
rect 27527 1948 27577 1994
rect 27324 1884 27334 1918
rect 27368 1884 27376 1918
rect 27324 1864 27376 1884
rect 27430 1920 27482 1948
rect 27430 1886 27438 1920
rect 27472 1886 27482 1920
rect 27430 1864 27482 1886
rect 27512 1910 27577 1948
rect 27512 1876 27533 1910
rect 27567 1876 27577 1910
rect 27512 1864 27577 1876
rect 27607 1944 27659 1994
rect 27810 1948 27860 1994
rect 27607 1910 27617 1944
rect 27651 1910 27659 1944
rect 27607 1864 27659 1910
rect 27713 1936 27765 1948
rect 27713 1902 27721 1936
rect 27755 1902 27765 1936
rect 27713 1864 27765 1902
rect 27795 1910 27860 1948
rect 27795 1876 27816 1910
rect 27850 1876 27860 1910
rect 27795 1864 27860 1876
rect 27890 1946 27942 1994
rect 27890 1912 27900 1946
rect 27934 1912 27942 1946
rect 27890 1864 27942 1912
rect 27996 1936 28048 1948
rect 27996 1902 28004 1936
rect 28038 1902 28048 1936
rect 27996 1864 28048 1902
rect 28078 1910 28132 1948
rect 28078 1876 28088 1910
rect 28122 1876 28132 1910
rect 28078 1864 28132 1876
rect 28162 1936 28214 1948
rect 28162 1902 28172 1936
rect 28206 1902 28214 1936
rect 28162 1864 28214 1902
rect 28268 1910 28320 1948
rect 28268 1876 28276 1910
rect 28310 1876 28320 1910
rect 28268 1864 28320 1876
rect 28350 1936 28400 1948
rect 28777 1948 28827 1992
rect 28566 1936 28617 1948
rect 28350 1928 28415 1936
rect 28350 1894 28360 1928
rect 28394 1894 28415 1928
rect 28350 1864 28415 1894
rect 28445 1910 28521 1936
rect 28445 1876 28466 1910
rect 28500 1876 28521 1910
rect 28445 1864 28521 1876
rect 28551 1864 28617 1936
rect 28647 1906 28727 1948
rect 28647 1872 28683 1906
rect 28717 1872 28727 1906
rect 28647 1864 28727 1872
rect 28757 1926 28827 1948
rect 28757 1892 28767 1926
rect 28801 1892 28827 1926
rect 28757 1864 28827 1892
rect 28857 1970 28911 1992
rect 28857 1936 28867 1970
rect 28901 1936 28911 1970
rect 28857 1864 28911 1936
rect 28941 1944 28993 1992
rect 28941 1910 28951 1944
rect 28985 1910 28993 1944
rect 28941 1864 28993 1910
rect 29047 1910 29099 1992
rect 29047 1876 29055 1910
rect 29089 1876 29099 1910
rect 29047 1864 29099 1876
rect 29129 1936 29179 1992
rect 29552 1948 29602 1992
rect 29348 1936 29398 1948
rect 29129 1864 29194 1936
rect 29224 1910 29303 1936
rect 29224 1876 29249 1910
rect 29283 1876 29303 1910
rect 29224 1864 29303 1876
rect 29333 1864 29398 1936
rect 29428 1906 29484 1948
rect 29428 1872 29440 1906
rect 29474 1872 29484 1906
rect 29428 1864 29484 1872
rect 29514 1926 29602 1948
rect 29514 1892 29542 1926
rect 29576 1892 29602 1926
rect 29514 1864 29602 1892
rect 29632 1970 29686 1992
rect 29632 1936 29642 1970
rect 29676 1936 29686 1970
rect 29632 1864 29686 1936
rect 29716 1918 29768 1992
rect 29919 1948 29969 1994
rect 29716 1884 29726 1918
rect 29760 1884 29768 1918
rect 29716 1864 29768 1884
rect 29822 1920 29874 1948
rect 29822 1886 29830 1920
rect 29864 1886 29874 1920
rect 29822 1864 29874 1886
rect 29904 1910 29969 1948
rect 29904 1876 29925 1910
rect 29959 1876 29969 1910
rect 29904 1864 29969 1876
rect 29999 1944 30051 1994
rect 30202 1948 30252 1994
rect 29999 1910 30009 1944
rect 30043 1910 30051 1944
rect 29999 1864 30051 1910
rect 30105 1936 30157 1948
rect 30105 1902 30113 1936
rect 30147 1902 30157 1936
rect 30105 1864 30157 1902
rect 30187 1910 30252 1948
rect 30187 1876 30208 1910
rect 30242 1876 30252 1910
rect 30187 1864 30252 1876
rect 30282 1946 30334 1994
rect 30282 1912 30292 1946
rect 30326 1912 30334 1946
rect 30282 1864 30334 1912
rect 8604 951 8656 996
rect 8604 917 8612 951
rect 8646 917 8656 951
rect 8604 892 8656 917
rect 8686 938 8744 996
rect 8686 904 8698 938
rect 8732 904 8744 938
rect 8686 892 8744 904
rect 8774 968 8826 996
rect 8774 934 8784 968
rect 8818 934 8826 968
rect 8774 892 8826 934
rect 8880 974 8932 1022
rect 8880 940 8888 974
rect 8922 940 8932 974
rect 8880 892 8932 940
rect 8962 942 9016 1022
rect 8962 908 8972 942
rect 9006 908 9016 942
rect 8962 892 9016 908
rect 9046 974 9100 1022
rect 9046 940 9056 974
rect 9090 940 9100 974
rect 9046 892 9100 940
rect 9130 942 9184 1022
rect 9130 908 9140 942
rect 9174 908 9184 942
rect 9130 892 9184 908
rect 9214 974 9268 1022
rect 9214 940 9224 974
rect 9258 940 9268 974
rect 9214 892 9268 940
rect 9298 1006 9350 1022
rect 9298 972 9308 1006
rect 9342 972 9350 1006
rect 9298 938 9350 972
rect 9298 904 9308 938
rect 9342 904 9350 938
rect 9298 892 9350 904
rect 9432 1010 9484 1022
rect 9432 976 9440 1010
rect 9474 976 9484 1010
rect 9432 942 9484 976
rect 9432 908 9440 942
rect 9474 908 9484 942
rect 9432 892 9484 908
rect 9514 1010 9568 1022
rect 9514 976 9524 1010
rect 9558 976 9568 1010
rect 9514 942 9568 976
rect 9514 908 9524 942
rect 9558 908 9568 942
rect 9514 892 9568 908
rect 9598 942 9652 1022
rect 9598 908 9608 942
rect 9642 908 9652 942
rect 9598 892 9652 908
rect 9682 1010 9736 1022
rect 9682 976 9692 1010
rect 9726 976 9736 1010
rect 9682 942 9736 976
rect 9682 908 9692 942
rect 9726 908 9736 942
rect 9682 892 9736 908
rect 9766 942 9820 1022
rect 9766 908 9776 942
rect 9810 908 9820 942
rect 9766 892 9820 908
rect 9850 1010 9904 1022
rect 9850 976 9860 1010
rect 9894 976 9904 1010
rect 9850 942 9904 976
rect 9850 908 9860 942
rect 9894 908 9904 942
rect 9850 892 9904 908
rect 9934 942 9988 1022
rect 9934 908 9944 942
rect 9978 908 9988 942
rect 9934 892 9988 908
rect 10018 1010 10072 1022
rect 10018 976 10028 1010
rect 10062 976 10072 1010
rect 10018 942 10072 976
rect 10018 908 10028 942
rect 10062 908 10072 942
rect 10018 892 10072 908
rect 10102 942 10156 1022
rect 10102 908 10112 942
rect 10146 908 10156 942
rect 10102 892 10156 908
rect 10186 1010 10240 1022
rect 10186 976 10196 1010
rect 10230 976 10240 1010
rect 10186 942 10240 976
rect 10186 908 10196 942
rect 10230 908 10240 942
rect 10186 892 10240 908
rect 10270 942 10324 1022
rect 10270 908 10280 942
rect 10314 908 10324 942
rect 10270 892 10324 908
rect 10354 1010 10408 1022
rect 10354 976 10364 1010
rect 10398 976 10408 1010
rect 10354 942 10408 976
rect 10354 908 10364 942
rect 10398 908 10408 942
rect 10354 892 10408 908
rect 10438 942 10492 1022
rect 10438 908 10448 942
rect 10482 908 10492 942
rect 10438 892 10492 908
rect 10522 1010 10576 1022
rect 10522 976 10532 1010
rect 10566 976 10576 1010
rect 10522 942 10576 976
rect 10522 908 10532 942
rect 10566 908 10576 942
rect 10522 892 10576 908
rect 10606 942 10660 1022
rect 10606 908 10616 942
rect 10650 908 10660 942
rect 10606 892 10660 908
rect 10690 1010 10744 1022
rect 10690 976 10700 1010
rect 10734 976 10744 1010
rect 10690 942 10744 976
rect 10690 908 10700 942
rect 10734 908 10744 942
rect 10690 892 10744 908
rect 10774 942 10828 1022
rect 10774 908 10784 942
rect 10818 908 10828 942
rect 10774 892 10828 908
rect 10858 1010 10912 1022
rect 10858 976 10868 1010
rect 10902 976 10912 1010
rect 10858 942 10912 976
rect 10858 908 10868 942
rect 10902 908 10912 942
rect 10858 892 10912 908
rect 10942 942 10996 1022
rect 10942 908 10952 942
rect 10986 908 10996 942
rect 10942 892 10996 908
rect 11026 1010 11080 1022
rect 11026 976 11036 1010
rect 11070 976 11080 1010
rect 11026 942 11080 976
rect 11026 908 11036 942
rect 11070 908 11080 942
rect 11026 892 11080 908
rect 11110 942 11164 1022
rect 11110 908 11120 942
rect 11154 908 11164 942
rect 11110 892 11164 908
rect 11194 1010 11248 1022
rect 11194 976 11204 1010
rect 11238 976 11248 1010
rect 11194 942 11248 976
rect 11194 908 11204 942
rect 11238 908 11248 942
rect 11194 892 11248 908
rect 11278 942 11330 1022
rect 11278 908 11288 942
rect 11322 908 11330 942
rect 11278 892 11330 908
rect 12988 951 13040 996
rect 12988 917 12996 951
rect 13030 917 13040 951
rect 12988 892 13040 917
rect 13070 938 13128 996
rect 13070 904 13082 938
rect 13116 904 13128 938
rect 13070 892 13128 904
rect 13158 968 13210 996
rect 13158 934 13168 968
rect 13202 934 13210 968
rect 13158 892 13210 934
rect 13264 974 13316 1022
rect 13264 940 13272 974
rect 13306 940 13316 974
rect 13264 892 13316 940
rect 13346 942 13400 1022
rect 13346 908 13356 942
rect 13390 908 13400 942
rect 13346 892 13400 908
rect 13430 974 13484 1022
rect 13430 940 13440 974
rect 13474 940 13484 974
rect 13430 892 13484 940
rect 13514 942 13568 1022
rect 13514 908 13524 942
rect 13558 908 13568 942
rect 13514 892 13568 908
rect 13598 974 13652 1022
rect 13598 940 13608 974
rect 13642 940 13652 974
rect 13598 892 13652 940
rect 13682 1006 13734 1022
rect 13682 972 13692 1006
rect 13726 972 13734 1006
rect 13682 938 13734 972
rect 13682 904 13692 938
rect 13726 904 13734 938
rect 13682 892 13734 904
rect 13816 1010 13868 1022
rect 13816 976 13824 1010
rect 13858 976 13868 1010
rect 13816 942 13868 976
rect 13816 908 13824 942
rect 13858 908 13868 942
rect 13816 892 13868 908
rect 13898 1010 13952 1022
rect 13898 976 13908 1010
rect 13942 976 13952 1010
rect 13898 942 13952 976
rect 13898 908 13908 942
rect 13942 908 13952 942
rect 13898 892 13952 908
rect 13982 942 14036 1022
rect 13982 908 13992 942
rect 14026 908 14036 942
rect 13982 892 14036 908
rect 14066 1010 14120 1022
rect 14066 976 14076 1010
rect 14110 976 14120 1010
rect 14066 942 14120 976
rect 14066 908 14076 942
rect 14110 908 14120 942
rect 14066 892 14120 908
rect 14150 942 14204 1022
rect 14150 908 14160 942
rect 14194 908 14204 942
rect 14150 892 14204 908
rect 14234 1010 14288 1022
rect 14234 976 14244 1010
rect 14278 976 14288 1010
rect 14234 942 14288 976
rect 14234 908 14244 942
rect 14278 908 14288 942
rect 14234 892 14288 908
rect 14318 942 14372 1022
rect 14318 908 14328 942
rect 14362 908 14372 942
rect 14318 892 14372 908
rect 14402 1010 14456 1022
rect 14402 976 14412 1010
rect 14446 976 14456 1010
rect 14402 942 14456 976
rect 14402 908 14412 942
rect 14446 908 14456 942
rect 14402 892 14456 908
rect 14486 942 14540 1022
rect 14486 908 14496 942
rect 14530 908 14540 942
rect 14486 892 14540 908
rect 14570 1010 14624 1022
rect 14570 976 14580 1010
rect 14614 976 14624 1010
rect 14570 942 14624 976
rect 14570 908 14580 942
rect 14614 908 14624 942
rect 14570 892 14624 908
rect 14654 942 14708 1022
rect 14654 908 14664 942
rect 14698 908 14708 942
rect 14654 892 14708 908
rect 14738 1010 14792 1022
rect 14738 976 14748 1010
rect 14782 976 14792 1010
rect 14738 942 14792 976
rect 14738 908 14748 942
rect 14782 908 14792 942
rect 14738 892 14792 908
rect 14822 942 14876 1022
rect 14822 908 14832 942
rect 14866 908 14876 942
rect 14822 892 14876 908
rect 14906 1010 14960 1022
rect 14906 976 14916 1010
rect 14950 976 14960 1010
rect 14906 942 14960 976
rect 14906 908 14916 942
rect 14950 908 14960 942
rect 14906 892 14960 908
rect 14990 942 15044 1022
rect 14990 908 15000 942
rect 15034 908 15044 942
rect 14990 892 15044 908
rect 15074 1010 15128 1022
rect 15074 976 15084 1010
rect 15118 976 15128 1010
rect 15074 942 15128 976
rect 15074 908 15084 942
rect 15118 908 15128 942
rect 15074 892 15128 908
rect 15158 942 15212 1022
rect 15158 908 15168 942
rect 15202 908 15212 942
rect 15158 892 15212 908
rect 15242 1010 15296 1022
rect 15242 976 15252 1010
rect 15286 976 15296 1010
rect 15242 942 15296 976
rect 15242 908 15252 942
rect 15286 908 15296 942
rect 15242 892 15296 908
rect 15326 942 15380 1022
rect 15326 908 15336 942
rect 15370 908 15380 942
rect 15326 892 15380 908
rect 15410 1010 15464 1022
rect 15410 976 15420 1010
rect 15454 976 15464 1010
rect 15410 942 15464 976
rect 15410 908 15420 942
rect 15454 908 15464 942
rect 15410 892 15464 908
rect 15494 942 15548 1022
rect 15494 908 15504 942
rect 15538 908 15548 942
rect 15494 892 15548 908
rect 15578 1010 15632 1022
rect 15578 976 15588 1010
rect 15622 976 15632 1010
rect 15578 942 15632 976
rect 15578 908 15588 942
rect 15622 908 15632 942
rect 15578 892 15632 908
rect 15662 942 15714 1022
rect 15662 908 15672 942
rect 15706 908 15714 942
rect 15662 892 15714 908
rect 8602 -185 8654 -120
rect 8602 -219 8610 -185
rect 8644 -219 8654 -185
rect 8602 -250 8654 -219
rect 8684 -166 8736 -120
rect 10676 -166 10728 -120
rect 8684 -204 8763 -166
rect 8684 -238 8694 -204
rect 8728 -238 8763 -204
rect 8684 -250 8763 -238
rect 8793 -250 8859 -166
rect 8889 -189 8984 -166
rect 8889 -223 8901 -189
rect 8935 -223 8984 -189
rect 8889 -250 8984 -223
rect 9014 -250 9080 -166
rect 9110 -189 9248 -166
rect 9110 -223 9136 -189
rect 9170 -223 9204 -189
rect 9238 -223 9248 -189
rect 9110 -250 9248 -223
rect 9278 -189 9330 -166
rect 9278 -223 9288 -189
rect 9322 -223 9330 -189
rect 9278 -250 9330 -223
rect 10082 -189 10134 -166
rect 10082 -223 10090 -189
rect 10124 -223 10134 -189
rect 10082 -250 10134 -223
rect 10164 -189 10302 -166
rect 10164 -223 10174 -189
rect 10208 -223 10242 -189
rect 10276 -223 10302 -189
rect 10164 -250 10302 -223
rect 10332 -250 10398 -166
rect 10428 -189 10523 -166
rect 10428 -223 10477 -189
rect 10511 -223 10523 -189
rect 10428 -250 10523 -223
rect 10553 -250 10619 -166
rect 10649 -204 10728 -166
rect 10649 -238 10684 -204
rect 10718 -238 10728 -204
rect 10649 -250 10728 -238
rect 10758 -185 10810 -120
rect 10758 -219 10768 -185
rect 10802 -219 10810 -185
rect 10758 -250 10810 -219
rect 10994 -185 11046 -120
rect 10994 -219 11002 -185
rect 11036 -219 11046 -185
rect 10994 -250 11046 -219
rect 11076 -166 11128 -120
rect 13068 -166 13120 -120
rect 11076 -204 11155 -166
rect 11076 -238 11086 -204
rect 11120 -238 11155 -204
rect 11076 -250 11155 -238
rect 11185 -250 11251 -166
rect 11281 -189 11376 -166
rect 11281 -223 11293 -189
rect 11327 -223 11376 -189
rect 11281 -250 11376 -223
rect 11406 -250 11472 -166
rect 11502 -189 11640 -166
rect 11502 -223 11528 -189
rect 11562 -223 11596 -189
rect 11630 -223 11640 -189
rect 11502 -250 11640 -223
rect 11670 -189 11722 -166
rect 11670 -223 11680 -189
rect 11714 -223 11722 -189
rect 11670 -250 11722 -223
rect 12474 -189 12526 -166
rect 12474 -223 12482 -189
rect 12516 -223 12526 -189
rect 12474 -250 12526 -223
rect 12556 -189 12694 -166
rect 12556 -223 12566 -189
rect 12600 -223 12634 -189
rect 12668 -223 12694 -189
rect 12556 -250 12694 -223
rect 12724 -250 12790 -166
rect 12820 -189 12915 -166
rect 12820 -223 12869 -189
rect 12903 -223 12915 -189
rect 12820 -250 12915 -223
rect 12945 -250 13011 -166
rect 13041 -204 13120 -166
rect 13041 -238 13076 -204
rect 13110 -238 13120 -204
rect 13041 -250 13120 -238
rect 13150 -185 13202 -120
rect 13150 -219 13160 -185
rect 13194 -219 13202 -185
rect 13150 -250 13202 -219
rect 13386 -185 13438 -120
rect 13386 -219 13394 -185
rect 13428 -219 13438 -185
rect 13386 -250 13438 -219
rect 13468 -166 13520 -120
rect 15458 -166 15510 -120
rect 13468 -204 13547 -166
rect 13468 -238 13478 -204
rect 13512 -238 13547 -204
rect 13468 -250 13547 -238
rect 13577 -250 13643 -166
rect 13673 -189 13768 -166
rect 13673 -223 13685 -189
rect 13719 -223 13768 -189
rect 13673 -250 13768 -223
rect 13798 -250 13864 -166
rect 13894 -189 14032 -166
rect 13894 -223 13920 -189
rect 13954 -223 13988 -189
rect 14022 -223 14032 -189
rect 13894 -250 14032 -223
rect 14062 -189 14114 -166
rect 14062 -223 14072 -189
rect 14106 -223 14114 -189
rect 14062 -250 14114 -223
rect 14864 -189 14916 -166
rect 14864 -223 14872 -189
rect 14906 -223 14916 -189
rect 14864 -250 14916 -223
rect 14946 -189 15084 -166
rect 14946 -223 14956 -189
rect 14990 -223 15024 -189
rect 15058 -223 15084 -189
rect 14946 -250 15084 -223
rect 15114 -250 15180 -166
rect 15210 -189 15305 -166
rect 15210 -223 15259 -189
rect 15293 -223 15305 -189
rect 15210 -250 15305 -223
rect 15335 -250 15401 -166
rect 15431 -204 15510 -166
rect 15431 -238 15466 -204
rect 15500 -238 15510 -204
rect 15431 -250 15510 -238
rect 15540 -185 15592 -120
rect 15540 -219 15550 -185
rect 15584 -219 15592 -185
rect 15540 -250 15592 -219
rect 15778 -185 15830 -120
rect 15778 -219 15786 -185
rect 15820 -219 15830 -185
rect 15778 -250 15830 -219
rect 15860 -166 15912 -120
rect 17852 -166 17904 -120
rect 15860 -204 15939 -166
rect 15860 -238 15870 -204
rect 15904 -238 15939 -204
rect 15860 -250 15939 -238
rect 15969 -250 16035 -166
rect 16065 -189 16160 -166
rect 16065 -223 16077 -189
rect 16111 -223 16160 -189
rect 16065 -250 16160 -223
rect 16190 -250 16256 -166
rect 16286 -189 16424 -166
rect 16286 -223 16312 -189
rect 16346 -223 16380 -189
rect 16414 -223 16424 -189
rect 16286 -250 16424 -223
rect 16454 -189 16506 -166
rect 16454 -223 16464 -189
rect 16498 -223 16506 -189
rect 16454 -250 16506 -223
rect 17258 -189 17310 -166
rect 17258 -223 17266 -189
rect 17300 -223 17310 -189
rect 17258 -250 17310 -223
rect 17340 -189 17478 -166
rect 17340 -223 17350 -189
rect 17384 -223 17418 -189
rect 17452 -223 17478 -189
rect 17340 -250 17478 -223
rect 17508 -250 17574 -166
rect 17604 -189 17699 -166
rect 17604 -223 17653 -189
rect 17687 -223 17699 -189
rect 17604 -250 17699 -223
rect 17729 -250 17795 -166
rect 17825 -204 17904 -166
rect 17825 -238 17860 -204
rect 17894 -238 17904 -204
rect 17825 -250 17904 -238
rect 17934 -185 17986 -120
rect 17934 -219 17944 -185
rect 17978 -219 17986 -185
rect 17934 -250 17986 -219
rect 18170 -185 18222 -120
rect 18170 -219 18178 -185
rect 18212 -219 18222 -185
rect 18170 -250 18222 -219
rect 18252 -166 18304 -120
rect 20244 -166 20296 -120
rect 18252 -204 18331 -166
rect 18252 -238 18262 -204
rect 18296 -238 18331 -204
rect 18252 -250 18331 -238
rect 18361 -250 18427 -166
rect 18457 -189 18552 -166
rect 18457 -223 18469 -189
rect 18503 -223 18552 -189
rect 18457 -250 18552 -223
rect 18582 -250 18648 -166
rect 18678 -189 18816 -166
rect 18678 -223 18704 -189
rect 18738 -223 18772 -189
rect 18806 -223 18816 -189
rect 18678 -250 18816 -223
rect 18846 -189 18898 -166
rect 18846 -223 18856 -189
rect 18890 -223 18898 -189
rect 18846 -250 18898 -223
rect 19650 -189 19702 -166
rect 19650 -223 19658 -189
rect 19692 -223 19702 -189
rect 19650 -250 19702 -223
rect 19732 -189 19870 -166
rect 19732 -223 19742 -189
rect 19776 -223 19810 -189
rect 19844 -223 19870 -189
rect 19732 -250 19870 -223
rect 19900 -250 19966 -166
rect 19996 -189 20091 -166
rect 19996 -223 20045 -189
rect 20079 -223 20091 -189
rect 19996 -250 20091 -223
rect 20121 -250 20187 -166
rect 20217 -204 20296 -166
rect 20217 -238 20252 -204
rect 20286 -238 20296 -204
rect 20217 -250 20296 -238
rect 20326 -185 20378 -120
rect 20326 -219 20336 -185
rect 20370 -219 20378 -185
rect 20326 -250 20378 -219
rect 20562 -185 20614 -120
rect 20562 -219 20570 -185
rect 20604 -219 20614 -185
rect 20562 -250 20614 -219
rect 20644 -166 20696 -120
rect 22634 -166 22686 -120
rect 20644 -204 20723 -166
rect 20644 -238 20654 -204
rect 20688 -238 20723 -204
rect 20644 -250 20723 -238
rect 20753 -250 20819 -166
rect 20849 -189 20944 -166
rect 20849 -223 20861 -189
rect 20895 -223 20944 -189
rect 20849 -250 20944 -223
rect 20974 -250 21040 -166
rect 21070 -189 21208 -166
rect 21070 -223 21096 -189
rect 21130 -223 21164 -189
rect 21198 -223 21208 -189
rect 21070 -250 21208 -223
rect 21238 -189 21290 -166
rect 21238 -223 21248 -189
rect 21282 -223 21290 -189
rect 21238 -250 21290 -223
rect 22040 -189 22092 -166
rect 22040 -223 22048 -189
rect 22082 -223 22092 -189
rect 22040 -250 22092 -223
rect 22122 -189 22260 -166
rect 22122 -223 22132 -189
rect 22166 -223 22200 -189
rect 22234 -223 22260 -189
rect 22122 -250 22260 -223
rect 22290 -250 22356 -166
rect 22386 -189 22481 -166
rect 22386 -223 22435 -189
rect 22469 -223 22481 -189
rect 22386 -250 22481 -223
rect 22511 -250 22577 -166
rect 22607 -204 22686 -166
rect 22607 -238 22642 -204
rect 22676 -238 22686 -204
rect 22607 -250 22686 -238
rect 22716 -185 22768 -120
rect 22716 -219 22726 -185
rect 22760 -219 22768 -185
rect 22716 -250 22768 -219
rect 22954 -185 23006 -120
rect 22954 -219 22962 -185
rect 22996 -219 23006 -185
rect 22954 -250 23006 -219
rect 23036 -166 23088 -120
rect 25028 -166 25080 -120
rect 23036 -204 23115 -166
rect 23036 -238 23046 -204
rect 23080 -238 23115 -204
rect 23036 -250 23115 -238
rect 23145 -250 23211 -166
rect 23241 -189 23336 -166
rect 23241 -223 23253 -189
rect 23287 -223 23336 -189
rect 23241 -250 23336 -223
rect 23366 -250 23432 -166
rect 23462 -189 23600 -166
rect 23462 -223 23488 -189
rect 23522 -223 23556 -189
rect 23590 -223 23600 -189
rect 23462 -250 23600 -223
rect 23630 -189 23682 -166
rect 23630 -223 23640 -189
rect 23674 -223 23682 -189
rect 23630 -250 23682 -223
rect 24434 -189 24486 -166
rect 24434 -223 24442 -189
rect 24476 -223 24486 -189
rect 24434 -250 24486 -223
rect 24516 -189 24654 -166
rect 24516 -223 24526 -189
rect 24560 -223 24594 -189
rect 24628 -223 24654 -189
rect 24516 -250 24654 -223
rect 24684 -250 24750 -166
rect 24780 -189 24875 -166
rect 24780 -223 24829 -189
rect 24863 -223 24875 -189
rect 24780 -250 24875 -223
rect 24905 -250 24971 -166
rect 25001 -204 25080 -166
rect 25001 -238 25036 -204
rect 25070 -238 25080 -204
rect 25001 -250 25080 -238
rect 25110 -185 25162 -120
rect 25110 -219 25120 -185
rect 25154 -219 25162 -185
rect 25110 -250 25162 -219
rect 8602 -866 8654 -854
rect 8602 -900 8610 -866
rect 8644 -900 8654 -866
rect 8602 -938 8654 -900
rect 8684 -892 8738 -854
rect 8684 -926 8694 -892
rect 8728 -926 8738 -892
rect 8684 -938 8738 -926
rect 8768 -866 8820 -854
rect 8768 -900 8778 -866
rect 8812 -900 8820 -866
rect 8768 -938 8820 -900
rect 8874 -892 8926 -854
rect 8874 -926 8882 -892
rect 8916 -926 8926 -892
rect 8874 -938 8926 -926
rect 8956 -866 9006 -854
rect 9381 -854 9432 -810
rect 9171 -866 9222 -854
rect 8956 -874 9021 -866
rect 8956 -908 8966 -874
rect 9000 -908 9021 -874
rect 8956 -938 9021 -908
rect 9051 -892 9126 -866
rect 9051 -926 9071 -892
rect 9105 -926 9126 -892
rect 9051 -938 9126 -926
rect 9156 -938 9222 -866
rect 9252 -896 9336 -854
rect 9252 -930 9292 -896
rect 9326 -930 9336 -896
rect 9252 -938 9336 -930
rect 9366 -890 9432 -854
rect 9366 -924 9376 -890
rect 9410 -924 9432 -890
rect 9366 -938 9432 -924
rect 9462 -832 9516 -810
rect 9462 -866 9472 -832
rect 9506 -866 9516 -832
rect 9462 -938 9516 -866
rect 9546 -858 9598 -810
rect 9546 -892 9556 -858
rect 9590 -892 9598 -858
rect 9546 -938 9598 -892
rect 9652 -892 9704 -810
rect 9652 -926 9660 -892
rect 9694 -926 9704 -892
rect 9652 -938 9704 -926
rect 9734 -866 9784 -810
rect 10158 -854 10208 -810
rect 9953 -866 10003 -854
rect 9734 -938 9824 -866
rect 9854 -892 9908 -866
rect 9854 -926 9864 -892
rect 9898 -926 9908 -892
rect 9854 -938 9908 -926
rect 9938 -938 10003 -866
rect 10033 -896 10100 -854
rect 10033 -930 10056 -896
rect 10090 -930 10100 -896
rect 10033 -938 10100 -930
rect 10130 -876 10208 -854
rect 10130 -910 10140 -876
rect 10174 -910 10208 -876
rect 10130 -938 10208 -910
rect 10238 -818 10292 -810
rect 10238 -852 10248 -818
rect 10282 -852 10292 -818
rect 10238 -938 10292 -852
rect 10322 -884 10374 -810
rect 10525 -854 10575 -808
rect 10322 -918 10332 -884
rect 10366 -918 10374 -884
rect 10322 -938 10374 -918
rect 10428 -882 10480 -854
rect 10428 -916 10436 -882
rect 10470 -916 10480 -882
rect 10428 -938 10480 -916
rect 10510 -892 10575 -854
rect 10510 -926 10531 -892
rect 10565 -926 10575 -892
rect 10510 -938 10575 -926
rect 10605 -858 10657 -808
rect 10808 -854 10858 -808
rect 10605 -892 10615 -858
rect 10649 -892 10657 -858
rect 10605 -938 10657 -892
rect 10711 -866 10763 -854
rect 10711 -900 10719 -866
rect 10753 -900 10763 -866
rect 10711 -938 10763 -900
rect 10793 -892 10858 -854
rect 10793 -926 10814 -892
rect 10848 -926 10858 -892
rect 10793 -938 10858 -926
rect 10888 -856 10940 -808
rect 10888 -890 10898 -856
rect 10932 -890 10940 -856
rect 10888 -938 10940 -890
rect 10994 -866 11046 -854
rect 10994 -900 11002 -866
rect 11036 -900 11046 -866
rect 10994 -938 11046 -900
rect 11076 -892 11130 -854
rect 11076 -926 11086 -892
rect 11120 -926 11130 -892
rect 11076 -938 11130 -926
rect 11160 -866 11212 -854
rect 11160 -900 11170 -866
rect 11204 -900 11212 -866
rect 11160 -938 11212 -900
rect 11266 -892 11318 -854
rect 11266 -926 11274 -892
rect 11308 -926 11318 -892
rect 11266 -938 11318 -926
rect 11348 -866 11398 -854
rect 11773 -854 11824 -810
rect 11563 -866 11614 -854
rect 11348 -874 11413 -866
rect 11348 -908 11358 -874
rect 11392 -908 11413 -874
rect 11348 -938 11413 -908
rect 11443 -892 11518 -866
rect 11443 -926 11463 -892
rect 11497 -926 11518 -892
rect 11443 -938 11518 -926
rect 11548 -938 11614 -866
rect 11644 -896 11728 -854
rect 11644 -930 11684 -896
rect 11718 -930 11728 -896
rect 11644 -938 11728 -930
rect 11758 -890 11824 -854
rect 11758 -924 11768 -890
rect 11802 -924 11824 -890
rect 11758 -938 11824 -924
rect 11854 -832 11908 -810
rect 11854 -866 11864 -832
rect 11898 -866 11908 -832
rect 11854 -938 11908 -866
rect 11938 -858 11990 -810
rect 11938 -892 11948 -858
rect 11982 -892 11990 -858
rect 11938 -938 11990 -892
rect 12044 -892 12096 -810
rect 12044 -926 12052 -892
rect 12086 -926 12096 -892
rect 12044 -938 12096 -926
rect 12126 -866 12176 -810
rect 12550 -854 12600 -810
rect 12345 -866 12395 -854
rect 12126 -938 12216 -866
rect 12246 -892 12300 -866
rect 12246 -926 12256 -892
rect 12290 -926 12300 -892
rect 12246 -938 12300 -926
rect 12330 -938 12395 -866
rect 12425 -896 12492 -854
rect 12425 -930 12448 -896
rect 12482 -930 12492 -896
rect 12425 -938 12492 -930
rect 12522 -876 12600 -854
rect 12522 -910 12532 -876
rect 12566 -910 12600 -876
rect 12522 -938 12600 -910
rect 12630 -818 12684 -810
rect 12630 -852 12640 -818
rect 12674 -852 12684 -818
rect 12630 -938 12684 -852
rect 12714 -884 12766 -810
rect 12917 -854 12967 -808
rect 12714 -918 12724 -884
rect 12758 -918 12766 -884
rect 12714 -938 12766 -918
rect 12820 -882 12872 -854
rect 12820 -916 12828 -882
rect 12862 -916 12872 -882
rect 12820 -938 12872 -916
rect 12902 -892 12967 -854
rect 12902 -926 12923 -892
rect 12957 -926 12967 -892
rect 12902 -938 12967 -926
rect 12997 -858 13049 -808
rect 13200 -854 13250 -808
rect 12997 -892 13007 -858
rect 13041 -892 13049 -858
rect 12997 -938 13049 -892
rect 13103 -866 13155 -854
rect 13103 -900 13111 -866
rect 13145 -900 13155 -866
rect 13103 -938 13155 -900
rect 13185 -892 13250 -854
rect 13185 -926 13206 -892
rect 13240 -926 13250 -892
rect 13185 -938 13250 -926
rect 13280 -856 13332 -808
rect 13280 -890 13290 -856
rect 13324 -890 13332 -856
rect 13280 -938 13332 -890
rect 13386 -866 13438 -854
rect 13386 -900 13394 -866
rect 13428 -900 13438 -866
rect 13386 -938 13438 -900
rect 13468 -892 13522 -854
rect 13468 -926 13478 -892
rect 13512 -926 13522 -892
rect 13468 -938 13522 -926
rect 13552 -866 13604 -854
rect 13552 -900 13562 -866
rect 13596 -900 13604 -866
rect 13552 -938 13604 -900
rect 13658 -892 13710 -854
rect 13658 -926 13666 -892
rect 13700 -926 13710 -892
rect 13658 -938 13710 -926
rect 13740 -866 13790 -854
rect 14165 -854 14216 -810
rect 13955 -866 14006 -854
rect 13740 -874 13805 -866
rect 13740 -908 13750 -874
rect 13784 -908 13805 -874
rect 13740 -938 13805 -908
rect 13835 -892 13910 -866
rect 13835 -926 13855 -892
rect 13889 -926 13910 -892
rect 13835 -938 13910 -926
rect 13940 -938 14006 -866
rect 14036 -896 14120 -854
rect 14036 -930 14076 -896
rect 14110 -930 14120 -896
rect 14036 -938 14120 -930
rect 14150 -890 14216 -854
rect 14150 -924 14160 -890
rect 14194 -924 14216 -890
rect 14150 -938 14216 -924
rect 14246 -832 14300 -810
rect 14246 -866 14256 -832
rect 14290 -866 14300 -832
rect 14246 -938 14300 -866
rect 14330 -858 14382 -810
rect 14330 -892 14340 -858
rect 14374 -892 14382 -858
rect 14330 -938 14382 -892
rect 14436 -892 14488 -810
rect 14436 -926 14444 -892
rect 14478 -926 14488 -892
rect 14436 -938 14488 -926
rect 14518 -866 14568 -810
rect 14942 -854 14992 -810
rect 14737 -866 14787 -854
rect 14518 -938 14608 -866
rect 14638 -892 14692 -866
rect 14638 -926 14648 -892
rect 14682 -926 14692 -892
rect 14638 -938 14692 -926
rect 14722 -938 14787 -866
rect 14817 -896 14884 -854
rect 14817 -930 14840 -896
rect 14874 -930 14884 -896
rect 14817 -938 14884 -930
rect 14914 -876 14992 -854
rect 14914 -910 14924 -876
rect 14958 -910 14992 -876
rect 14914 -938 14992 -910
rect 15022 -818 15076 -810
rect 15022 -852 15032 -818
rect 15066 -852 15076 -818
rect 15022 -938 15076 -852
rect 15106 -884 15158 -810
rect 15309 -854 15359 -808
rect 15106 -918 15116 -884
rect 15150 -918 15158 -884
rect 15106 -938 15158 -918
rect 15212 -882 15264 -854
rect 15212 -916 15220 -882
rect 15254 -916 15264 -882
rect 15212 -938 15264 -916
rect 15294 -892 15359 -854
rect 15294 -926 15315 -892
rect 15349 -926 15359 -892
rect 15294 -938 15359 -926
rect 15389 -858 15441 -808
rect 15592 -854 15642 -808
rect 15389 -892 15399 -858
rect 15433 -892 15441 -858
rect 15389 -938 15441 -892
rect 15495 -866 15547 -854
rect 15495 -900 15503 -866
rect 15537 -900 15547 -866
rect 15495 -938 15547 -900
rect 15577 -892 15642 -854
rect 15577 -926 15598 -892
rect 15632 -926 15642 -892
rect 15577 -938 15642 -926
rect 15672 -856 15724 -808
rect 15672 -890 15682 -856
rect 15716 -890 15724 -856
rect 15672 -938 15724 -890
rect 15778 -866 15830 -854
rect 15778 -900 15786 -866
rect 15820 -900 15830 -866
rect 15778 -938 15830 -900
rect 15860 -892 15914 -854
rect 15860 -926 15870 -892
rect 15904 -926 15914 -892
rect 15860 -938 15914 -926
rect 15944 -866 15996 -854
rect 15944 -900 15954 -866
rect 15988 -900 15996 -866
rect 15944 -938 15996 -900
rect 16050 -892 16102 -854
rect 16050 -926 16058 -892
rect 16092 -926 16102 -892
rect 16050 -938 16102 -926
rect 16132 -866 16182 -854
rect 16557 -854 16608 -810
rect 16347 -866 16398 -854
rect 16132 -874 16197 -866
rect 16132 -908 16142 -874
rect 16176 -908 16197 -874
rect 16132 -938 16197 -908
rect 16227 -892 16302 -866
rect 16227 -926 16247 -892
rect 16281 -926 16302 -892
rect 16227 -938 16302 -926
rect 16332 -938 16398 -866
rect 16428 -896 16512 -854
rect 16428 -930 16468 -896
rect 16502 -930 16512 -896
rect 16428 -938 16512 -930
rect 16542 -890 16608 -854
rect 16542 -924 16552 -890
rect 16586 -924 16608 -890
rect 16542 -938 16608 -924
rect 16638 -832 16692 -810
rect 16638 -866 16648 -832
rect 16682 -866 16692 -832
rect 16638 -938 16692 -866
rect 16722 -858 16774 -810
rect 16722 -892 16732 -858
rect 16766 -892 16774 -858
rect 16722 -938 16774 -892
rect 16828 -892 16880 -810
rect 16828 -926 16836 -892
rect 16870 -926 16880 -892
rect 16828 -938 16880 -926
rect 16910 -866 16960 -810
rect 17334 -854 17384 -810
rect 17129 -866 17179 -854
rect 16910 -938 17000 -866
rect 17030 -892 17084 -866
rect 17030 -926 17040 -892
rect 17074 -926 17084 -892
rect 17030 -938 17084 -926
rect 17114 -938 17179 -866
rect 17209 -896 17276 -854
rect 17209 -930 17232 -896
rect 17266 -930 17276 -896
rect 17209 -938 17276 -930
rect 17306 -876 17384 -854
rect 17306 -910 17316 -876
rect 17350 -910 17384 -876
rect 17306 -938 17384 -910
rect 17414 -818 17468 -810
rect 17414 -852 17424 -818
rect 17458 -852 17468 -818
rect 17414 -938 17468 -852
rect 17498 -884 17550 -810
rect 17701 -854 17751 -808
rect 17498 -918 17508 -884
rect 17542 -918 17550 -884
rect 17498 -938 17550 -918
rect 17604 -882 17656 -854
rect 17604 -916 17612 -882
rect 17646 -916 17656 -882
rect 17604 -938 17656 -916
rect 17686 -892 17751 -854
rect 17686 -926 17707 -892
rect 17741 -926 17751 -892
rect 17686 -938 17751 -926
rect 17781 -858 17833 -808
rect 17984 -854 18034 -808
rect 17781 -892 17791 -858
rect 17825 -892 17833 -858
rect 17781 -938 17833 -892
rect 17887 -866 17939 -854
rect 17887 -900 17895 -866
rect 17929 -900 17939 -866
rect 17887 -938 17939 -900
rect 17969 -892 18034 -854
rect 17969 -926 17990 -892
rect 18024 -926 18034 -892
rect 17969 -938 18034 -926
rect 18064 -856 18116 -808
rect 18064 -890 18074 -856
rect 18108 -890 18116 -856
rect 18064 -938 18116 -890
rect 18170 -866 18222 -854
rect 18170 -900 18178 -866
rect 18212 -900 18222 -866
rect 18170 -938 18222 -900
rect 18252 -892 18306 -854
rect 18252 -926 18262 -892
rect 18296 -926 18306 -892
rect 18252 -938 18306 -926
rect 18336 -866 18388 -854
rect 18336 -900 18346 -866
rect 18380 -900 18388 -866
rect 18336 -938 18388 -900
rect 18442 -892 18494 -854
rect 18442 -926 18450 -892
rect 18484 -926 18494 -892
rect 18442 -938 18494 -926
rect 18524 -866 18574 -854
rect 18949 -854 19000 -810
rect 18739 -866 18790 -854
rect 18524 -874 18589 -866
rect 18524 -908 18534 -874
rect 18568 -908 18589 -874
rect 18524 -938 18589 -908
rect 18619 -892 18694 -866
rect 18619 -926 18639 -892
rect 18673 -926 18694 -892
rect 18619 -938 18694 -926
rect 18724 -938 18790 -866
rect 18820 -896 18904 -854
rect 18820 -930 18860 -896
rect 18894 -930 18904 -896
rect 18820 -938 18904 -930
rect 18934 -890 19000 -854
rect 18934 -924 18944 -890
rect 18978 -924 19000 -890
rect 18934 -938 19000 -924
rect 19030 -832 19084 -810
rect 19030 -866 19040 -832
rect 19074 -866 19084 -832
rect 19030 -938 19084 -866
rect 19114 -858 19166 -810
rect 19114 -892 19124 -858
rect 19158 -892 19166 -858
rect 19114 -938 19166 -892
rect 19220 -892 19272 -810
rect 19220 -926 19228 -892
rect 19262 -926 19272 -892
rect 19220 -938 19272 -926
rect 19302 -866 19352 -810
rect 19726 -854 19776 -810
rect 19521 -866 19571 -854
rect 19302 -938 19392 -866
rect 19422 -892 19476 -866
rect 19422 -926 19432 -892
rect 19466 -926 19476 -892
rect 19422 -938 19476 -926
rect 19506 -938 19571 -866
rect 19601 -896 19668 -854
rect 19601 -930 19624 -896
rect 19658 -930 19668 -896
rect 19601 -938 19668 -930
rect 19698 -876 19776 -854
rect 19698 -910 19708 -876
rect 19742 -910 19776 -876
rect 19698 -938 19776 -910
rect 19806 -818 19860 -810
rect 19806 -852 19816 -818
rect 19850 -852 19860 -818
rect 19806 -938 19860 -852
rect 19890 -884 19942 -810
rect 20093 -854 20143 -808
rect 19890 -918 19900 -884
rect 19934 -918 19942 -884
rect 19890 -938 19942 -918
rect 19996 -882 20048 -854
rect 19996 -916 20004 -882
rect 20038 -916 20048 -882
rect 19996 -938 20048 -916
rect 20078 -892 20143 -854
rect 20078 -926 20099 -892
rect 20133 -926 20143 -892
rect 20078 -938 20143 -926
rect 20173 -858 20225 -808
rect 20376 -854 20426 -808
rect 20173 -892 20183 -858
rect 20217 -892 20225 -858
rect 20173 -938 20225 -892
rect 20279 -866 20331 -854
rect 20279 -900 20287 -866
rect 20321 -900 20331 -866
rect 20279 -938 20331 -900
rect 20361 -892 20426 -854
rect 20361 -926 20382 -892
rect 20416 -926 20426 -892
rect 20361 -938 20426 -926
rect 20456 -856 20508 -808
rect 20456 -890 20466 -856
rect 20500 -890 20508 -856
rect 20456 -938 20508 -890
rect 20562 -866 20614 -854
rect 20562 -900 20570 -866
rect 20604 -900 20614 -866
rect 20562 -938 20614 -900
rect 20644 -892 20698 -854
rect 20644 -926 20654 -892
rect 20688 -926 20698 -892
rect 20644 -938 20698 -926
rect 20728 -866 20780 -854
rect 20728 -900 20738 -866
rect 20772 -900 20780 -866
rect 20728 -938 20780 -900
rect 20834 -892 20886 -854
rect 20834 -926 20842 -892
rect 20876 -926 20886 -892
rect 20834 -938 20886 -926
rect 20916 -866 20966 -854
rect 21341 -854 21392 -810
rect 21131 -866 21182 -854
rect 20916 -874 20981 -866
rect 20916 -908 20926 -874
rect 20960 -908 20981 -874
rect 20916 -938 20981 -908
rect 21011 -892 21086 -866
rect 21011 -926 21031 -892
rect 21065 -926 21086 -892
rect 21011 -938 21086 -926
rect 21116 -938 21182 -866
rect 21212 -896 21296 -854
rect 21212 -930 21252 -896
rect 21286 -930 21296 -896
rect 21212 -938 21296 -930
rect 21326 -890 21392 -854
rect 21326 -924 21336 -890
rect 21370 -924 21392 -890
rect 21326 -938 21392 -924
rect 21422 -832 21476 -810
rect 21422 -866 21432 -832
rect 21466 -866 21476 -832
rect 21422 -938 21476 -866
rect 21506 -858 21558 -810
rect 21506 -892 21516 -858
rect 21550 -892 21558 -858
rect 21506 -938 21558 -892
rect 21612 -892 21664 -810
rect 21612 -926 21620 -892
rect 21654 -926 21664 -892
rect 21612 -938 21664 -926
rect 21694 -866 21744 -810
rect 22118 -854 22168 -810
rect 21913 -866 21963 -854
rect 21694 -938 21784 -866
rect 21814 -892 21868 -866
rect 21814 -926 21824 -892
rect 21858 -926 21868 -892
rect 21814 -938 21868 -926
rect 21898 -938 21963 -866
rect 21993 -896 22060 -854
rect 21993 -930 22016 -896
rect 22050 -930 22060 -896
rect 21993 -938 22060 -930
rect 22090 -876 22168 -854
rect 22090 -910 22100 -876
rect 22134 -910 22168 -876
rect 22090 -938 22168 -910
rect 22198 -818 22252 -810
rect 22198 -852 22208 -818
rect 22242 -852 22252 -818
rect 22198 -938 22252 -852
rect 22282 -884 22334 -810
rect 22485 -854 22535 -808
rect 22282 -918 22292 -884
rect 22326 -918 22334 -884
rect 22282 -938 22334 -918
rect 22388 -882 22440 -854
rect 22388 -916 22396 -882
rect 22430 -916 22440 -882
rect 22388 -938 22440 -916
rect 22470 -892 22535 -854
rect 22470 -926 22491 -892
rect 22525 -926 22535 -892
rect 22470 -938 22535 -926
rect 22565 -858 22617 -808
rect 22768 -854 22818 -808
rect 22565 -892 22575 -858
rect 22609 -892 22617 -858
rect 22565 -938 22617 -892
rect 22671 -866 22723 -854
rect 22671 -900 22679 -866
rect 22713 -900 22723 -866
rect 22671 -938 22723 -900
rect 22753 -892 22818 -854
rect 22753 -926 22774 -892
rect 22808 -926 22818 -892
rect 22753 -938 22818 -926
rect 22848 -856 22900 -808
rect 22848 -890 22858 -856
rect 22892 -890 22900 -856
rect 22848 -938 22900 -890
rect 22954 -866 23006 -854
rect 22954 -900 22962 -866
rect 22996 -900 23006 -866
rect 22954 -938 23006 -900
rect 23036 -892 23090 -854
rect 23036 -926 23046 -892
rect 23080 -926 23090 -892
rect 23036 -938 23090 -926
rect 23120 -866 23172 -854
rect 23120 -900 23130 -866
rect 23164 -900 23172 -866
rect 23120 -938 23172 -900
rect 23226 -892 23278 -854
rect 23226 -926 23234 -892
rect 23268 -926 23278 -892
rect 23226 -938 23278 -926
rect 23308 -866 23358 -854
rect 23733 -854 23784 -810
rect 23523 -866 23574 -854
rect 23308 -874 23373 -866
rect 23308 -908 23318 -874
rect 23352 -908 23373 -874
rect 23308 -938 23373 -908
rect 23403 -892 23478 -866
rect 23403 -926 23423 -892
rect 23457 -926 23478 -892
rect 23403 -938 23478 -926
rect 23508 -938 23574 -866
rect 23604 -896 23688 -854
rect 23604 -930 23644 -896
rect 23678 -930 23688 -896
rect 23604 -938 23688 -930
rect 23718 -890 23784 -854
rect 23718 -924 23728 -890
rect 23762 -924 23784 -890
rect 23718 -938 23784 -924
rect 23814 -832 23868 -810
rect 23814 -866 23824 -832
rect 23858 -866 23868 -832
rect 23814 -938 23868 -866
rect 23898 -858 23950 -810
rect 23898 -892 23908 -858
rect 23942 -892 23950 -858
rect 23898 -938 23950 -892
rect 24004 -892 24056 -810
rect 24004 -926 24012 -892
rect 24046 -926 24056 -892
rect 24004 -938 24056 -926
rect 24086 -866 24136 -810
rect 24510 -854 24560 -810
rect 24305 -866 24355 -854
rect 24086 -938 24176 -866
rect 24206 -892 24260 -866
rect 24206 -926 24216 -892
rect 24250 -926 24260 -892
rect 24206 -938 24260 -926
rect 24290 -938 24355 -866
rect 24385 -896 24452 -854
rect 24385 -930 24408 -896
rect 24442 -930 24452 -896
rect 24385 -938 24452 -930
rect 24482 -876 24560 -854
rect 24482 -910 24492 -876
rect 24526 -910 24560 -876
rect 24482 -938 24560 -910
rect 24590 -818 24644 -810
rect 24590 -852 24600 -818
rect 24634 -852 24644 -818
rect 24590 -938 24644 -852
rect 24674 -884 24726 -810
rect 24877 -854 24927 -808
rect 24674 -918 24684 -884
rect 24718 -918 24726 -884
rect 24674 -938 24726 -918
rect 24780 -882 24832 -854
rect 24780 -916 24788 -882
rect 24822 -916 24832 -882
rect 24780 -938 24832 -916
rect 24862 -892 24927 -854
rect 24862 -926 24883 -892
rect 24917 -926 24927 -892
rect 24862 -938 24927 -926
rect 24957 -858 25009 -808
rect 25160 -854 25210 -808
rect 24957 -892 24967 -858
rect 25001 -892 25009 -858
rect 24957 -938 25009 -892
rect 25063 -866 25115 -854
rect 25063 -900 25071 -866
rect 25105 -900 25115 -866
rect 25063 -938 25115 -900
rect 25145 -892 25210 -854
rect 25145 -926 25166 -892
rect 25200 -926 25210 -892
rect 25145 -938 25210 -926
rect 25240 -856 25292 -808
rect 25240 -890 25250 -856
rect 25284 -890 25292 -856
rect 25240 -938 25292 -890
rect 8602 -1545 8654 -1497
rect 8602 -1579 8610 -1545
rect 8644 -1579 8654 -1545
rect 8602 -1627 8654 -1579
rect 8684 -1543 8734 -1497
rect 8684 -1581 8749 -1543
rect 8684 -1615 8694 -1581
rect 8728 -1615 8749 -1581
rect 8684 -1627 8749 -1615
rect 8779 -1555 8831 -1543
rect 8779 -1589 8789 -1555
rect 8823 -1589 8831 -1555
rect 8779 -1627 8831 -1589
rect 8885 -1547 8937 -1497
rect 8885 -1581 8893 -1547
rect 8927 -1581 8937 -1547
rect 8885 -1627 8937 -1581
rect 8967 -1543 9017 -1497
rect 8967 -1581 9032 -1543
rect 8967 -1615 8977 -1581
rect 9011 -1615 9032 -1581
rect 8967 -1627 9032 -1615
rect 9062 -1571 9114 -1543
rect 9062 -1605 9072 -1571
rect 9106 -1605 9114 -1571
rect 9062 -1627 9114 -1605
rect 9168 -1573 9220 -1499
rect 9168 -1607 9176 -1573
rect 9210 -1607 9220 -1573
rect 9168 -1627 9220 -1607
rect 9250 -1507 9304 -1499
rect 9250 -1541 9260 -1507
rect 9294 -1541 9304 -1507
rect 9250 -1627 9304 -1541
rect 9334 -1543 9384 -1499
rect 9334 -1565 9412 -1543
rect 9334 -1599 9368 -1565
rect 9402 -1599 9412 -1565
rect 9334 -1627 9412 -1599
rect 9442 -1585 9509 -1543
rect 9442 -1619 9452 -1585
rect 9486 -1619 9509 -1585
rect 9442 -1627 9509 -1619
rect 9539 -1555 9589 -1543
rect 9758 -1555 9808 -1499
rect 9539 -1627 9604 -1555
rect 9634 -1581 9688 -1555
rect 9634 -1615 9644 -1581
rect 9678 -1615 9688 -1581
rect 9634 -1627 9688 -1615
rect 9718 -1627 9808 -1555
rect 9838 -1581 9890 -1499
rect 9838 -1615 9848 -1581
rect 9882 -1615 9890 -1581
rect 9838 -1627 9890 -1615
rect 9944 -1547 9996 -1499
rect 9944 -1581 9952 -1547
rect 9986 -1581 9996 -1547
rect 9944 -1627 9996 -1581
rect 10026 -1521 10080 -1499
rect 10026 -1555 10036 -1521
rect 10070 -1555 10080 -1521
rect 10026 -1627 10080 -1555
rect 10110 -1543 10161 -1499
rect 10110 -1579 10176 -1543
rect 10110 -1613 10132 -1579
rect 10166 -1613 10176 -1579
rect 10110 -1627 10176 -1613
rect 10206 -1585 10290 -1543
rect 10206 -1619 10216 -1585
rect 10250 -1619 10290 -1585
rect 10206 -1627 10290 -1619
rect 10320 -1555 10371 -1543
rect 10536 -1555 10586 -1543
rect 10320 -1627 10386 -1555
rect 10416 -1581 10491 -1555
rect 10416 -1615 10437 -1581
rect 10471 -1615 10491 -1581
rect 10416 -1627 10491 -1615
rect 10521 -1563 10586 -1555
rect 10521 -1597 10542 -1563
rect 10576 -1597 10586 -1563
rect 10521 -1627 10586 -1597
rect 10616 -1581 10668 -1543
rect 10616 -1615 10626 -1581
rect 10660 -1615 10668 -1581
rect 10616 -1627 10668 -1615
rect 10722 -1555 10774 -1543
rect 10722 -1589 10730 -1555
rect 10764 -1589 10774 -1555
rect 10722 -1627 10774 -1589
rect 10804 -1581 10858 -1543
rect 10804 -1615 10814 -1581
rect 10848 -1615 10858 -1581
rect 10804 -1627 10858 -1615
rect 10888 -1555 10940 -1543
rect 10888 -1589 10898 -1555
rect 10932 -1589 10940 -1555
rect 10888 -1627 10940 -1589
rect 10994 -1545 11046 -1497
rect 10994 -1579 11002 -1545
rect 11036 -1579 11046 -1545
rect 10994 -1627 11046 -1579
rect 11076 -1543 11126 -1497
rect 11076 -1581 11141 -1543
rect 11076 -1615 11086 -1581
rect 11120 -1615 11141 -1581
rect 11076 -1627 11141 -1615
rect 11171 -1555 11223 -1543
rect 11171 -1589 11181 -1555
rect 11215 -1589 11223 -1555
rect 11171 -1627 11223 -1589
rect 11277 -1547 11329 -1497
rect 11277 -1581 11285 -1547
rect 11319 -1581 11329 -1547
rect 11277 -1627 11329 -1581
rect 11359 -1543 11409 -1497
rect 11359 -1581 11424 -1543
rect 11359 -1615 11369 -1581
rect 11403 -1615 11424 -1581
rect 11359 -1627 11424 -1615
rect 11454 -1571 11506 -1543
rect 11454 -1605 11464 -1571
rect 11498 -1605 11506 -1571
rect 11454 -1627 11506 -1605
rect 11560 -1573 11612 -1499
rect 11560 -1607 11568 -1573
rect 11602 -1607 11612 -1573
rect 11560 -1627 11612 -1607
rect 11642 -1507 11696 -1499
rect 11642 -1541 11652 -1507
rect 11686 -1541 11696 -1507
rect 11642 -1627 11696 -1541
rect 11726 -1543 11776 -1499
rect 11726 -1565 11804 -1543
rect 11726 -1599 11760 -1565
rect 11794 -1599 11804 -1565
rect 11726 -1627 11804 -1599
rect 11834 -1585 11901 -1543
rect 11834 -1619 11844 -1585
rect 11878 -1619 11901 -1585
rect 11834 -1627 11901 -1619
rect 11931 -1555 11981 -1543
rect 12150 -1555 12200 -1499
rect 11931 -1627 11996 -1555
rect 12026 -1581 12080 -1555
rect 12026 -1615 12036 -1581
rect 12070 -1615 12080 -1581
rect 12026 -1627 12080 -1615
rect 12110 -1627 12200 -1555
rect 12230 -1581 12282 -1499
rect 12230 -1615 12240 -1581
rect 12274 -1615 12282 -1581
rect 12230 -1627 12282 -1615
rect 12336 -1547 12388 -1499
rect 12336 -1581 12344 -1547
rect 12378 -1581 12388 -1547
rect 12336 -1627 12388 -1581
rect 12418 -1521 12472 -1499
rect 12418 -1555 12428 -1521
rect 12462 -1555 12472 -1521
rect 12418 -1627 12472 -1555
rect 12502 -1543 12553 -1499
rect 12502 -1579 12568 -1543
rect 12502 -1613 12524 -1579
rect 12558 -1613 12568 -1579
rect 12502 -1627 12568 -1613
rect 12598 -1585 12682 -1543
rect 12598 -1619 12608 -1585
rect 12642 -1619 12682 -1585
rect 12598 -1627 12682 -1619
rect 12712 -1555 12763 -1543
rect 12928 -1555 12978 -1543
rect 12712 -1627 12778 -1555
rect 12808 -1581 12883 -1555
rect 12808 -1615 12829 -1581
rect 12863 -1615 12883 -1581
rect 12808 -1627 12883 -1615
rect 12913 -1563 12978 -1555
rect 12913 -1597 12934 -1563
rect 12968 -1597 12978 -1563
rect 12913 -1627 12978 -1597
rect 13008 -1581 13060 -1543
rect 13008 -1615 13018 -1581
rect 13052 -1615 13060 -1581
rect 13008 -1627 13060 -1615
rect 13114 -1555 13166 -1543
rect 13114 -1589 13122 -1555
rect 13156 -1589 13166 -1555
rect 13114 -1627 13166 -1589
rect 13196 -1581 13250 -1543
rect 13196 -1615 13206 -1581
rect 13240 -1615 13250 -1581
rect 13196 -1627 13250 -1615
rect 13280 -1555 13332 -1543
rect 13280 -1589 13290 -1555
rect 13324 -1589 13332 -1555
rect 13280 -1627 13332 -1589
rect 13386 -1545 13438 -1497
rect 13386 -1579 13394 -1545
rect 13428 -1579 13438 -1545
rect 13386 -1627 13438 -1579
rect 13468 -1543 13518 -1497
rect 13468 -1581 13533 -1543
rect 13468 -1615 13478 -1581
rect 13512 -1615 13533 -1581
rect 13468 -1627 13533 -1615
rect 13563 -1555 13615 -1543
rect 13563 -1589 13573 -1555
rect 13607 -1589 13615 -1555
rect 13563 -1627 13615 -1589
rect 13669 -1547 13721 -1497
rect 13669 -1581 13677 -1547
rect 13711 -1581 13721 -1547
rect 13669 -1627 13721 -1581
rect 13751 -1543 13801 -1497
rect 13751 -1581 13816 -1543
rect 13751 -1615 13761 -1581
rect 13795 -1615 13816 -1581
rect 13751 -1627 13816 -1615
rect 13846 -1571 13898 -1543
rect 13846 -1605 13856 -1571
rect 13890 -1605 13898 -1571
rect 13846 -1627 13898 -1605
rect 13952 -1573 14004 -1499
rect 13952 -1607 13960 -1573
rect 13994 -1607 14004 -1573
rect 13952 -1627 14004 -1607
rect 14034 -1507 14088 -1499
rect 14034 -1541 14044 -1507
rect 14078 -1541 14088 -1507
rect 14034 -1627 14088 -1541
rect 14118 -1543 14168 -1499
rect 14118 -1565 14196 -1543
rect 14118 -1599 14152 -1565
rect 14186 -1599 14196 -1565
rect 14118 -1627 14196 -1599
rect 14226 -1585 14293 -1543
rect 14226 -1619 14236 -1585
rect 14270 -1619 14293 -1585
rect 14226 -1627 14293 -1619
rect 14323 -1555 14373 -1543
rect 14542 -1555 14592 -1499
rect 14323 -1627 14388 -1555
rect 14418 -1581 14472 -1555
rect 14418 -1615 14428 -1581
rect 14462 -1615 14472 -1581
rect 14418 -1627 14472 -1615
rect 14502 -1627 14592 -1555
rect 14622 -1581 14674 -1499
rect 14622 -1615 14632 -1581
rect 14666 -1615 14674 -1581
rect 14622 -1627 14674 -1615
rect 14728 -1547 14780 -1499
rect 14728 -1581 14736 -1547
rect 14770 -1581 14780 -1547
rect 14728 -1627 14780 -1581
rect 14810 -1521 14864 -1499
rect 14810 -1555 14820 -1521
rect 14854 -1555 14864 -1521
rect 14810 -1627 14864 -1555
rect 14894 -1543 14945 -1499
rect 14894 -1579 14960 -1543
rect 14894 -1613 14916 -1579
rect 14950 -1613 14960 -1579
rect 14894 -1627 14960 -1613
rect 14990 -1585 15074 -1543
rect 14990 -1619 15000 -1585
rect 15034 -1619 15074 -1585
rect 14990 -1627 15074 -1619
rect 15104 -1555 15155 -1543
rect 15320 -1555 15370 -1543
rect 15104 -1627 15170 -1555
rect 15200 -1581 15275 -1555
rect 15200 -1615 15221 -1581
rect 15255 -1615 15275 -1581
rect 15200 -1627 15275 -1615
rect 15305 -1563 15370 -1555
rect 15305 -1597 15326 -1563
rect 15360 -1597 15370 -1563
rect 15305 -1627 15370 -1597
rect 15400 -1581 15452 -1543
rect 15400 -1615 15410 -1581
rect 15444 -1615 15452 -1581
rect 15400 -1627 15452 -1615
rect 15506 -1555 15558 -1543
rect 15506 -1589 15514 -1555
rect 15548 -1589 15558 -1555
rect 15506 -1627 15558 -1589
rect 15588 -1581 15642 -1543
rect 15588 -1615 15598 -1581
rect 15632 -1615 15642 -1581
rect 15588 -1627 15642 -1615
rect 15672 -1555 15724 -1543
rect 15672 -1589 15682 -1555
rect 15716 -1589 15724 -1555
rect 15672 -1627 15724 -1589
rect 15778 -1545 15830 -1497
rect 15778 -1579 15786 -1545
rect 15820 -1579 15830 -1545
rect 15778 -1627 15830 -1579
rect 15860 -1543 15910 -1497
rect 15860 -1581 15925 -1543
rect 15860 -1615 15870 -1581
rect 15904 -1615 15925 -1581
rect 15860 -1627 15925 -1615
rect 15955 -1555 16007 -1543
rect 15955 -1589 15965 -1555
rect 15999 -1589 16007 -1555
rect 15955 -1627 16007 -1589
rect 16061 -1547 16113 -1497
rect 16061 -1581 16069 -1547
rect 16103 -1581 16113 -1547
rect 16061 -1627 16113 -1581
rect 16143 -1543 16193 -1497
rect 16143 -1581 16208 -1543
rect 16143 -1615 16153 -1581
rect 16187 -1615 16208 -1581
rect 16143 -1627 16208 -1615
rect 16238 -1571 16290 -1543
rect 16238 -1605 16248 -1571
rect 16282 -1605 16290 -1571
rect 16238 -1627 16290 -1605
rect 16344 -1573 16396 -1499
rect 16344 -1607 16352 -1573
rect 16386 -1607 16396 -1573
rect 16344 -1627 16396 -1607
rect 16426 -1507 16480 -1499
rect 16426 -1541 16436 -1507
rect 16470 -1541 16480 -1507
rect 16426 -1627 16480 -1541
rect 16510 -1543 16560 -1499
rect 16510 -1565 16588 -1543
rect 16510 -1599 16544 -1565
rect 16578 -1599 16588 -1565
rect 16510 -1627 16588 -1599
rect 16618 -1585 16685 -1543
rect 16618 -1619 16628 -1585
rect 16662 -1619 16685 -1585
rect 16618 -1627 16685 -1619
rect 16715 -1555 16765 -1543
rect 16934 -1555 16984 -1499
rect 16715 -1627 16780 -1555
rect 16810 -1581 16864 -1555
rect 16810 -1615 16820 -1581
rect 16854 -1615 16864 -1581
rect 16810 -1627 16864 -1615
rect 16894 -1627 16984 -1555
rect 17014 -1581 17066 -1499
rect 17014 -1615 17024 -1581
rect 17058 -1615 17066 -1581
rect 17014 -1627 17066 -1615
rect 17120 -1547 17172 -1499
rect 17120 -1581 17128 -1547
rect 17162 -1581 17172 -1547
rect 17120 -1627 17172 -1581
rect 17202 -1521 17256 -1499
rect 17202 -1555 17212 -1521
rect 17246 -1555 17256 -1521
rect 17202 -1627 17256 -1555
rect 17286 -1543 17337 -1499
rect 17286 -1579 17352 -1543
rect 17286 -1613 17308 -1579
rect 17342 -1613 17352 -1579
rect 17286 -1627 17352 -1613
rect 17382 -1585 17466 -1543
rect 17382 -1619 17392 -1585
rect 17426 -1619 17466 -1585
rect 17382 -1627 17466 -1619
rect 17496 -1555 17547 -1543
rect 17712 -1555 17762 -1543
rect 17496 -1627 17562 -1555
rect 17592 -1581 17667 -1555
rect 17592 -1615 17613 -1581
rect 17647 -1615 17667 -1581
rect 17592 -1627 17667 -1615
rect 17697 -1563 17762 -1555
rect 17697 -1597 17718 -1563
rect 17752 -1597 17762 -1563
rect 17697 -1627 17762 -1597
rect 17792 -1581 17844 -1543
rect 17792 -1615 17802 -1581
rect 17836 -1615 17844 -1581
rect 17792 -1627 17844 -1615
rect 17898 -1555 17950 -1543
rect 17898 -1589 17906 -1555
rect 17940 -1589 17950 -1555
rect 17898 -1627 17950 -1589
rect 17980 -1581 18034 -1543
rect 17980 -1615 17990 -1581
rect 18024 -1615 18034 -1581
rect 17980 -1627 18034 -1615
rect 18064 -1555 18116 -1543
rect 18064 -1589 18074 -1555
rect 18108 -1589 18116 -1555
rect 18064 -1627 18116 -1589
rect 18170 -1545 18222 -1497
rect 18170 -1579 18178 -1545
rect 18212 -1579 18222 -1545
rect 18170 -1627 18222 -1579
rect 18252 -1543 18302 -1497
rect 18252 -1581 18317 -1543
rect 18252 -1615 18262 -1581
rect 18296 -1615 18317 -1581
rect 18252 -1627 18317 -1615
rect 18347 -1555 18399 -1543
rect 18347 -1589 18357 -1555
rect 18391 -1589 18399 -1555
rect 18347 -1627 18399 -1589
rect 18453 -1547 18505 -1497
rect 18453 -1581 18461 -1547
rect 18495 -1581 18505 -1547
rect 18453 -1627 18505 -1581
rect 18535 -1543 18585 -1497
rect 18535 -1581 18600 -1543
rect 18535 -1615 18545 -1581
rect 18579 -1615 18600 -1581
rect 18535 -1627 18600 -1615
rect 18630 -1571 18682 -1543
rect 18630 -1605 18640 -1571
rect 18674 -1605 18682 -1571
rect 18630 -1627 18682 -1605
rect 18736 -1573 18788 -1499
rect 18736 -1607 18744 -1573
rect 18778 -1607 18788 -1573
rect 18736 -1627 18788 -1607
rect 18818 -1507 18872 -1499
rect 18818 -1541 18828 -1507
rect 18862 -1541 18872 -1507
rect 18818 -1627 18872 -1541
rect 18902 -1543 18952 -1499
rect 18902 -1565 18980 -1543
rect 18902 -1599 18936 -1565
rect 18970 -1599 18980 -1565
rect 18902 -1627 18980 -1599
rect 19010 -1585 19077 -1543
rect 19010 -1619 19020 -1585
rect 19054 -1619 19077 -1585
rect 19010 -1627 19077 -1619
rect 19107 -1555 19157 -1543
rect 19326 -1555 19376 -1499
rect 19107 -1627 19172 -1555
rect 19202 -1581 19256 -1555
rect 19202 -1615 19212 -1581
rect 19246 -1615 19256 -1581
rect 19202 -1627 19256 -1615
rect 19286 -1627 19376 -1555
rect 19406 -1581 19458 -1499
rect 19406 -1615 19416 -1581
rect 19450 -1615 19458 -1581
rect 19406 -1627 19458 -1615
rect 19512 -1547 19564 -1499
rect 19512 -1581 19520 -1547
rect 19554 -1581 19564 -1547
rect 19512 -1627 19564 -1581
rect 19594 -1521 19648 -1499
rect 19594 -1555 19604 -1521
rect 19638 -1555 19648 -1521
rect 19594 -1627 19648 -1555
rect 19678 -1543 19729 -1499
rect 19678 -1579 19744 -1543
rect 19678 -1613 19700 -1579
rect 19734 -1613 19744 -1579
rect 19678 -1627 19744 -1613
rect 19774 -1585 19858 -1543
rect 19774 -1619 19784 -1585
rect 19818 -1619 19858 -1585
rect 19774 -1627 19858 -1619
rect 19888 -1555 19939 -1543
rect 20104 -1555 20154 -1543
rect 19888 -1627 19954 -1555
rect 19984 -1581 20059 -1555
rect 19984 -1615 20005 -1581
rect 20039 -1615 20059 -1581
rect 19984 -1627 20059 -1615
rect 20089 -1563 20154 -1555
rect 20089 -1597 20110 -1563
rect 20144 -1597 20154 -1563
rect 20089 -1627 20154 -1597
rect 20184 -1581 20236 -1543
rect 20184 -1615 20194 -1581
rect 20228 -1615 20236 -1581
rect 20184 -1627 20236 -1615
rect 20290 -1555 20342 -1543
rect 20290 -1589 20298 -1555
rect 20332 -1589 20342 -1555
rect 20290 -1627 20342 -1589
rect 20372 -1581 20426 -1543
rect 20372 -1615 20382 -1581
rect 20416 -1615 20426 -1581
rect 20372 -1627 20426 -1615
rect 20456 -1555 20508 -1543
rect 20456 -1589 20466 -1555
rect 20500 -1589 20508 -1555
rect 20456 -1627 20508 -1589
rect 20562 -1545 20614 -1497
rect 20562 -1579 20570 -1545
rect 20604 -1579 20614 -1545
rect 20562 -1627 20614 -1579
rect 20644 -1543 20694 -1497
rect 20644 -1581 20709 -1543
rect 20644 -1615 20654 -1581
rect 20688 -1615 20709 -1581
rect 20644 -1627 20709 -1615
rect 20739 -1555 20791 -1543
rect 20739 -1589 20749 -1555
rect 20783 -1589 20791 -1555
rect 20739 -1627 20791 -1589
rect 20845 -1547 20897 -1497
rect 20845 -1581 20853 -1547
rect 20887 -1581 20897 -1547
rect 20845 -1627 20897 -1581
rect 20927 -1543 20977 -1497
rect 20927 -1581 20992 -1543
rect 20927 -1615 20937 -1581
rect 20971 -1615 20992 -1581
rect 20927 -1627 20992 -1615
rect 21022 -1571 21074 -1543
rect 21022 -1605 21032 -1571
rect 21066 -1605 21074 -1571
rect 21022 -1627 21074 -1605
rect 21128 -1573 21180 -1499
rect 21128 -1607 21136 -1573
rect 21170 -1607 21180 -1573
rect 21128 -1627 21180 -1607
rect 21210 -1507 21264 -1499
rect 21210 -1541 21220 -1507
rect 21254 -1541 21264 -1507
rect 21210 -1627 21264 -1541
rect 21294 -1543 21344 -1499
rect 21294 -1565 21372 -1543
rect 21294 -1599 21328 -1565
rect 21362 -1599 21372 -1565
rect 21294 -1627 21372 -1599
rect 21402 -1585 21469 -1543
rect 21402 -1619 21412 -1585
rect 21446 -1619 21469 -1585
rect 21402 -1627 21469 -1619
rect 21499 -1555 21549 -1543
rect 21718 -1555 21768 -1499
rect 21499 -1627 21564 -1555
rect 21594 -1581 21648 -1555
rect 21594 -1615 21604 -1581
rect 21638 -1615 21648 -1581
rect 21594 -1627 21648 -1615
rect 21678 -1627 21768 -1555
rect 21798 -1581 21850 -1499
rect 21798 -1615 21808 -1581
rect 21842 -1615 21850 -1581
rect 21798 -1627 21850 -1615
rect 21904 -1547 21956 -1499
rect 21904 -1581 21912 -1547
rect 21946 -1581 21956 -1547
rect 21904 -1627 21956 -1581
rect 21986 -1521 22040 -1499
rect 21986 -1555 21996 -1521
rect 22030 -1555 22040 -1521
rect 21986 -1627 22040 -1555
rect 22070 -1543 22121 -1499
rect 22070 -1579 22136 -1543
rect 22070 -1613 22092 -1579
rect 22126 -1613 22136 -1579
rect 22070 -1627 22136 -1613
rect 22166 -1585 22250 -1543
rect 22166 -1619 22176 -1585
rect 22210 -1619 22250 -1585
rect 22166 -1627 22250 -1619
rect 22280 -1555 22331 -1543
rect 22496 -1555 22546 -1543
rect 22280 -1627 22346 -1555
rect 22376 -1581 22451 -1555
rect 22376 -1615 22397 -1581
rect 22431 -1615 22451 -1581
rect 22376 -1627 22451 -1615
rect 22481 -1563 22546 -1555
rect 22481 -1597 22502 -1563
rect 22536 -1597 22546 -1563
rect 22481 -1627 22546 -1597
rect 22576 -1581 22628 -1543
rect 22576 -1615 22586 -1581
rect 22620 -1615 22628 -1581
rect 22576 -1627 22628 -1615
rect 22682 -1555 22734 -1543
rect 22682 -1589 22690 -1555
rect 22724 -1589 22734 -1555
rect 22682 -1627 22734 -1589
rect 22764 -1581 22818 -1543
rect 22764 -1615 22774 -1581
rect 22808 -1615 22818 -1581
rect 22764 -1627 22818 -1615
rect 22848 -1555 22900 -1543
rect 22848 -1589 22858 -1555
rect 22892 -1589 22900 -1555
rect 22848 -1627 22900 -1589
rect 22954 -1545 23006 -1497
rect 22954 -1579 22962 -1545
rect 22996 -1579 23006 -1545
rect 22954 -1627 23006 -1579
rect 23036 -1543 23086 -1497
rect 23036 -1581 23101 -1543
rect 23036 -1615 23046 -1581
rect 23080 -1615 23101 -1581
rect 23036 -1627 23101 -1615
rect 23131 -1555 23183 -1543
rect 23131 -1589 23141 -1555
rect 23175 -1589 23183 -1555
rect 23131 -1627 23183 -1589
rect 23237 -1547 23289 -1497
rect 23237 -1581 23245 -1547
rect 23279 -1581 23289 -1547
rect 23237 -1627 23289 -1581
rect 23319 -1543 23369 -1497
rect 23319 -1581 23384 -1543
rect 23319 -1615 23329 -1581
rect 23363 -1615 23384 -1581
rect 23319 -1627 23384 -1615
rect 23414 -1571 23466 -1543
rect 23414 -1605 23424 -1571
rect 23458 -1605 23466 -1571
rect 23414 -1627 23466 -1605
rect 23520 -1573 23572 -1499
rect 23520 -1607 23528 -1573
rect 23562 -1607 23572 -1573
rect 23520 -1627 23572 -1607
rect 23602 -1507 23656 -1499
rect 23602 -1541 23612 -1507
rect 23646 -1541 23656 -1507
rect 23602 -1627 23656 -1541
rect 23686 -1543 23736 -1499
rect 23686 -1565 23764 -1543
rect 23686 -1599 23720 -1565
rect 23754 -1599 23764 -1565
rect 23686 -1627 23764 -1599
rect 23794 -1585 23861 -1543
rect 23794 -1619 23804 -1585
rect 23838 -1619 23861 -1585
rect 23794 -1627 23861 -1619
rect 23891 -1555 23941 -1543
rect 24110 -1555 24160 -1499
rect 23891 -1627 23956 -1555
rect 23986 -1581 24040 -1555
rect 23986 -1615 23996 -1581
rect 24030 -1615 24040 -1581
rect 23986 -1627 24040 -1615
rect 24070 -1627 24160 -1555
rect 24190 -1581 24242 -1499
rect 24190 -1615 24200 -1581
rect 24234 -1615 24242 -1581
rect 24190 -1627 24242 -1615
rect 24296 -1547 24348 -1499
rect 24296 -1581 24304 -1547
rect 24338 -1581 24348 -1547
rect 24296 -1627 24348 -1581
rect 24378 -1521 24432 -1499
rect 24378 -1555 24388 -1521
rect 24422 -1555 24432 -1521
rect 24378 -1627 24432 -1555
rect 24462 -1543 24513 -1499
rect 24462 -1579 24528 -1543
rect 24462 -1613 24484 -1579
rect 24518 -1613 24528 -1579
rect 24462 -1627 24528 -1613
rect 24558 -1585 24642 -1543
rect 24558 -1619 24568 -1585
rect 24602 -1619 24642 -1585
rect 24558 -1627 24642 -1619
rect 24672 -1555 24723 -1543
rect 24888 -1555 24938 -1543
rect 24672 -1627 24738 -1555
rect 24768 -1581 24843 -1555
rect 24768 -1615 24789 -1581
rect 24823 -1615 24843 -1581
rect 24768 -1627 24843 -1615
rect 24873 -1563 24938 -1555
rect 24873 -1597 24894 -1563
rect 24928 -1597 24938 -1563
rect 24873 -1627 24938 -1597
rect 24968 -1581 25020 -1543
rect 24968 -1615 24978 -1581
rect 25012 -1615 25020 -1581
rect 24968 -1627 25020 -1615
rect 25074 -1555 25126 -1543
rect 25074 -1589 25082 -1555
rect 25116 -1589 25126 -1555
rect 25074 -1627 25126 -1589
rect 25156 -1581 25210 -1543
rect 25156 -1615 25166 -1581
rect 25200 -1615 25210 -1581
rect 25156 -1627 25210 -1615
rect 25240 -1555 25292 -1543
rect 25240 -1589 25250 -1555
rect 25284 -1589 25292 -1555
rect 25240 -1627 25292 -1589
<< pdiff >>
rect 13804 13581 13862 13593
rect 13804 13521 13816 13581
rect 13850 13521 13862 13581
rect 13804 13509 13862 13521
rect 13892 13581 13950 13593
rect 13892 13521 13904 13581
rect 13938 13521 13950 13581
rect 13892 13509 13950 13521
rect 20513 13581 20571 13593
rect 20513 13521 20525 13581
rect 20559 13521 20571 13581
rect 20513 13509 20571 13521
rect 20601 13581 20659 13593
rect 20601 13521 20613 13581
rect 20647 13521 20659 13581
rect 20601 13509 20659 13521
rect 13804 13443 13862 13455
rect 13804 13383 13816 13443
rect 13850 13383 13862 13443
rect 13804 13371 13862 13383
rect 13892 13443 13950 13455
rect 13892 13383 13904 13443
rect 13938 13383 13950 13443
rect 13892 13371 13950 13383
rect 20513 13443 20571 13455
rect 20513 13383 20525 13443
rect 20559 13383 20571 13443
rect 20513 13371 20571 13383
rect 20601 13443 20659 13455
rect 20601 13383 20613 13443
rect 20647 13383 20659 13443
rect 20601 13371 20659 13383
rect 13804 13305 13862 13317
rect 13804 13245 13816 13305
rect 13850 13245 13862 13305
rect 13804 13233 13862 13245
rect 13892 13305 13950 13317
rect 13892 13245 13904 13305
rect 13938 13245 13950 13305
rect 20513 13305 20571 13317
rect 13892 13233 13950 13245
rect 20513 13245 20525 13305
rect 20559 13245 20571 13305
rect 20513 13233 20571 13245
rect 20601 13305 20659 13317
rect 20601 13245 20613 13305
rect 20647 13245 20659 13305
rect 20601 13233 20659 13245
rect 13804 13167 13862 13179
rect 2916 13106 2974 13118
rect 2916 13046 2928 13106
rect 2962 13046 2974 13106
rect 2916 13034 2974 13046
rect 3004 13106 3062 13118
rect 3004 13046 3016 13106
rect 3050 13046 3062 13106
rect 13804 13107 13816 13167
rect 13850 13107 13862 13167
rect 13804 13095 13862 13107
rect 13892 13167 13950 13179
rect 13892 13107 13904 13167
rect 13938 13107 13950 13167
rect 20513 13167 20571 13179
rect 13892 13095 13950 13107
rect 3004 13034 3062 13046
rect 20513 13107 20525 13167
rect 20559 13107 20571 13167
rect 20513 13095 20571 13107
rect 20601 13167 20659 13179
rect 20601 13107 20613 13167
rect 20647 13107 20659 13167
rect 20601 13095 20659 13107
rect 13804 13029 13862 13041
rect 2916 12968 2974 12980
rect 2916 12908 2928 12968
rect 2962 12908 2974 12968
rect 2916 12896 2974 12908
rect 3004 12968 3062 12980
rect 3004 12908 3016 12968
rect 3050 12908 3062 12968
rect 3004 12896 3062 12908
rect 13804 12969 13816 13029
rect 13850 12969 13862 13029
rect 13804 12957 13862 12969
rect 13892 13029 13950 13041
rect 13892 12969 13904 13029
rect 13938 12969 13950 13029
rect 20513 13029 20571 13041
rect 13892 12957 13950 12969
rect 13342 12934 13394 12946
rect 13342 12900 13350 12934
rect 13384 12900 13394 12934
rect 13342 12866 13394 12900
rect 2916 12830 2974 12842
rect 2916 12770 2928 12830
rect 2962 12770 2974 12830
rect 2916 12758 2974 12770
rect 3004 12830 3062 12842
rect 3004 12770 3016 12830
rect 3050 12770 3062 12830
rect 13342 12832 13350 12866
rect 13384 12832 13394 12866
rect 3004 12758 3062 12770
rect 13342 12798 13394 12832
rect 13342 12764 13350 12798
rect 13384 12764 13394 12798
rect 13342 12746 13394 12764
rect 13424 12934 13476 12946
rect 13424 12900 13434 12934
rect 13468 12900 13476 12934
rect 13424 12866 13476 12900
rect 13424 12832 13434 12866
rect 13468 12832 13476 12866
rect 13424 12798 13476 12832
rect 13424 12764 13434 12798
rect 13468 12764 13476 12798
rect 13424 12746 13476 12764
rect 13532 12934 13584 12946
rect 13532 12900 13540 12934
rect 13574 12900 13584 12934
rect 13532 12866 13584 12900
rect 13532 12832 13540 12866
rect 13574 12832 13584 12866
rect 13532 12798 13584 12832
rect 13532 12764 13540 12798
rect 13574 12764 13584 12798
rect 13532 12746 13584 12764
rect 13614 12934 13666 12946
rect 13614 12900 13624 12934
rect 13658 12900 13666 12934
rect 20513 12969 20525 13029
rect 20559 12969 20571 13029
rect 20513 12957 20571 12969
rect 20601 13029 20659 13041
rect 20601 12969 20613 13029
rect 20647 12969 20659 13029
rect 20601 12957 20659 12969
rect 13614 12866 13666 12900
rect 13614 12832 13624 12866
rect 13658 12832 13666 12866
rect 13614 12798 13666 12832
rect 13804 12891 13862 12903
rect 13804 12831 13816 12891
rect 13850 12831 13862 12891
rect 13804 12819 13862 12831
rect 13892 12891 13950 12903
rect 13892 12831 13904 12891
rect 13938 12831 13950 12891
rect 20051 12934 20103 12946
rect 20051 12900 20059 12934
rect 20093 12900 20103 12934
rect 13892 12819 13950 12831
rect 20051 12866 20103 12900
rect 20051 12832 20059 12866
rect 20093 12832 20103 12866
rect 13614 12764 13624 12798
rect 13658 12764 13666 12798
rect 20051 12798 20103 12832
rect 13614 12746 13666 12764
rect 2916 12692 2974 12704
rect 2916 12632 2928 12692
rect 2962 12632 2974 12692
rect 2916 12620 2974 12632
rect 3004 12692 3062 12704
rect 3004 12632 3016 12692
rect 3050 12632 3062 12692
rect 3004 12620 3062 12632
rect 20051 12764 20059 12798
rect 20093 12764 20103 12798
rect 20051 12746 20103 12764
rect 20133 12934 20185 12946
rect 20133 12900 20143 12934
rect 20177 12900 20185 12934
rect 20133 12866 20185 12900
rect 20133 12832 20143 12866
rect 20177 12832 20185 12866
rect 20133 12798 20185 12832
rect 20133 12764 20143 12798
rect 20177 12764 20185 12798
rect 20133 12746 20185 12764
rect 20241 12934 20293 12946
rect 20241 12900 20249 12934
rect 20283 12900 20293 12934
rect 20241 12866 20293 12900
rect 20241 12832 20249 12866
rect 20283 12832 20293 12866
rect 20241 12798 20293 12832
rect 20241 12764 20249 12798
rect 20283 12764 20293 12798
rect 20241 12746 20293 12764
rect 20323 12934 20375 12946
rect 20323 12900 20333 12934
rect 20367 12900 20375 12934
rect 20323 12866 20375 12900
rect 20323 12832 20333 12866
rect 20367 12832 20375 12866
rect 20323 12798 20375 12832
rect 20513 12891 20571 12903
rect 20513 12831 20525 12891
rect 20559 12831 20571 12891
rect 20513 12819 20571 12831
rect 20601 12891 20659 12903
rect 20601 12831 20613 12891
rect 20647 12831 20659 12891
rect 20601 12819 20659 12831
rect 20323 12764 20333 12798
rect 20367 12764 20375 12798
rect 20323 12746 20375 12764
rect 2916 12554 2974 12566
rect 2916 12494 2928 12554
rect 2962 12494 2974 12554
rect 2916 12482 2974 12494
rect 3004 12554 3062 12566
rect 3004 12494 3016 12554
rect 3050 12494 3062 12554
rect 3004 12482 3062 12494
rect 2454 12459 2506 12471
rect 2454 12425 2462 12459
rect 2496 12425 2506 12459
rect 2454 12391 2506 12425
rect 2454 12357 2462 12391
rect 2496 12357 2506 12391
rect 2454 12323 2506 12357
rect 2454 12289 2462 12323
rect 2496 12289 2506 12323
rect 2454 12271 2506 12289
rect 2536 12459 2588 12471
rect 2536 12425 2546 12459
rect 2580 12425 2588 12459
rect 2536 12391 2588 12425
rect 2536 12357 2546 12391
rect 2580 12357 2588 12391
rect 2536 12323 2588 12357
rect 2536 12289 2546 12323
rect 2580 12289 2588 12323
rect 2536 12271 2588 12289
rect 2644 12459 2696 12471
rect 2644 12425 2652 12459
rect 2686 12425 2696 12459
rect 2644 12391 2696 12425
rect 2644 12357 2652 12391
rect 2686 12357 2696 12391
rect 2644 12323 2696 12357
rect 2644 12289 2652 12323
rect 2686 12289 2696 12323
rect 2644 12271 2696 12289
rect 2726 12459 2778 12471
rect 2726 12425 2736 12459
rect 2770 12425 2778 12459
rect 19589 12580 19647 12592
rect 19589 12520 19601 12580
rect 19635 12520 19647 12580
rect 19589 12508 19647 12520
rect 19677 12580 19735 12592
rect 19677 12520 19689 12580
rect 19723 12520 19735 12580
rect 19677 12508 19735 12520
rect 2726 12391 2778 12425
rect 2726 12357 2736 12391
rect 2770 12357 2778 12391
rect 2726 12323 2778 12357
rect 2916 12416 2974 12428
rect 2916 12356 2928 12416
rect 2962 12356 2974 12416
rect 2916 12344 2974 12356
rect 3004 12416 3062 12428
rect 3004 12356 3016 12416
rect 3050 12356 3062 12416
rect 26298 12580 26356 12592
rect 26298 12520 26310 12580
rect 26344 12520 26356 12580
rect 26298 12508 26356 12520
rect 26386 12580 26444 12592
rect 26386 12520 26398 12580
rect 26432 12520 26444 12580
rect 26386 12508 26444 12520
rect 3004 12344 3062 12356
rect 2726 12289 2736 12323
rect 2770 12289 2778 12323
rect 2726 12271 2778 12289
rect 8701 12105 8759 12117
rect 8701 12045 8713 12105
rect 8747 12045 8759 12105
rect 8701 12033 8759 12045
rect 8789 12105 8847 12117
rect 8789 12045 8801 12105
rect 8835 12045 8847 12105
rect 8789 12033 8847 12045
rect 9129 12082 9181 12094
rect 9129 12048 9137 12082
rect 9171 12048 9181 12082
rect 9129 12014 9181 12048
rect 9129 11980 9137 12014
rect 9171 11980 9181 12014
rect 3558 11961 3616 11973
rect 3558 11901 3570 11961
rect 3604 11901 3616 11961
rect 3558 11889 3616 11901
rect 3646 11964 3704 11973
rect 3646 11904 3658 11964
rect 3692 11904 3704 11964
rect 3646 11889 3704 11904
rect 4290 11964 4348 11976
rect 4290 11904 4302 11964
rect 4336 11904 4348 11964
rect 4290 11892 4348 11904
rect 4378 11964 4474 11976
rect 4378 11904 4407 11964
rect 4441 11904 4474 11964
rect 4378 11892 4474 11904
rect 4504 11964 4562 11976
rect 4504 11904 4516 11964
rect 4550 11904 4562 11964
rect 4504 11892 4562 11904
rect 5502 11964 5560 11976
rect 5502 11904 5514 11964
rect 5548 11904 5560 11964
rect 5502 11892 5560 11904
rect 5590 11964 5686 11976
rect 5590 11904 5618 11964
rect 5652 11904 5686 11964
rect 5590 11892 5686 11904
rect 5716 11964 5774 11976
rect 5716 11904 5728 11964
rect 5762 11904 5774 11964
rect 5716 11892 5774 11904
rect 6714 11964 6772 11976
rect 6714 11904 6726 11964
rect 6760 11904 6772 11964
rect 6714 11892 6772 11904
rect 6802 11964 6898 11976
rect 6802 11904 6831 11964
rect 6865 11904 6898 11964
rect 6802 11892 6898 11904
rect 6928 11964 6986 11976
rect 6928 11904 6940 11964
rect 6974 11904 6986 11964
rect 6928 11892 6986 11904
rect 7926 11964 7984 11976
rect 7926 11904 7938 11964
rect 7972 11904 7984 11964
rect 7926 11892 7984 11904
rect 8014 11964 8110 11976
rect 8014 11904 8045 11964
rect 8079 11904 8110 11964
rect 8014 11892 8110 11904
rect 8140 11964 8198 11976
rect 8140 11904 8152 11964
rect 8186 11904 8198 11964
rect 8140 11892 8198 11904
rect 8701 11967 8759 11979
rect 8701 11907 8713 11967
rect 8747 11907 8759 11967
rect 8701 11895 8759 11907
rect 8789 11967 8851 11979
rect 8789 11907 8801 11967
rect 8835 11907 8851 11967
rect 8789 11895 8851 11907
rect 8881 11967 8947 11979
rect 8881 11907 8897 11967
rect 8931 11907 8947 11967
rect 8881 11895 8947 11907
rect 8977 11967 9039 11979
rect 8977 11907 8993 11967
rect 9027 11907 9039 11967
rect 8977 11895 9039 11907
rect 9129 11946 9181 11980
rect 9129 11912 9137 11946
rect 9171 11912 9181 11946
rect 9129 11894 9181 11912
rect 9211 12082 9263 12094
rect 9211 12048 9221 12082
rect 9255 12048 9263 12082
rect 9211 12014 9263 12048
rect 9211 11980 9221 12014
rect 9255 11980 9263 12014
rect 9211 11946 9263 11980
rect 10909 12074 10961 12086
rect 10909 12040 10917 12074
rect 10951 12040 10961 12074
rect 10909 12006 10961 12040
rect 10909 11972 10917 12006
rect 10951 11972 10961 12006
rect 10909 11958 10961 11972
rect 10991 12022 11045 12086
rect 10991 11988 11001 12022
rect 11035 11988 11045 12022
rect 10991 11958 11045 11988
rect 11075 12074 11127 12086
rect 11075 12040 11085 12074
rect 11119 12040 11127 12074
rect 11075 12006 11127 12040
rect 11682 12092 11744 12120
rect 11682 12058 11700 12092
rect 11734 12058 11744 12092
rect 11682 12036 11744 12058
rect 11075 11972 11085 12006
rect 11119 11972 11127 12006
rect 11075 11958 11127 11972
rect 11181 12022 11233 12036
rect 11181 11988 11189 12022
rect 11223 11988 11233 12022
rect 9211 11912 9221 11946
rect 9255 11912 9263 11946
rect 11181 11952 11233 11988
rect 11263 12006 11326 12036
rect 11263 11972 11273 12006
rect 11307 11972 11326 12006
rect 11263 11952 11326 11972
rect 11356 11999 11410 12036
rect 11356 11965 11366 11999
rect 11400 11965 11410 11999
rect 11356 11952 11410 11965
rect 11440 11952 11530 12036
rect 11560 12008 11636 12036
rect 11560 11974 11580 12008
rect 11614 11974 11636 12008
rect 11560 11952 11636 11974
rect 11666 12024 11744 12036
rect 11666 11990 11700 12024
rect 11734 11990 11744 12024
rect 11666 11952 11744 11990
rect 11774 11952 11828 12120
rect 11858 12066 11965 12120
rect 11858 12032 11874 12066
rect 11908 12032 11965 12066
rect 11858 11998 11965 12032
rect 11858 11964 11874 11998
rect 11908 11964 11965 11998
rect 11858 11952 11965 11964
rect 11995 12036 12047 12120
rect 14446 12436 14504 12448
rect 14446 12376 14458 12436
rect 14492 12376 14504 12436
rect 14446 12364 14504 12376
rect 14534 12439 14592 12448
rect 14534 12379 14546 12439
rect 14580 12379 14592 12439
rect 14534 12364 14592 12379
rect 15178 12439 15236 12451
rect 15178 12379 15190 12439
rect 15224 12379 15236 12439
rect 15178 12367 15236 12379
rect 15266 12439 15362 12451
rect 15266 12379 15295 12439
rect 15329 12379 15362 12439
rect 15266 12367 15362 12379
rect 15392 12439 15450 12451
rect 15392 12379 15404 12439
rect 15438 12379 15450 12439
rect 15392 12367 15450 12379
rect 16390 12439 16448 12451
rect 16390 12379 16402 12439
rect 16436 12379 16448 12439
rect 16390 12367 16448 12379
rect 16478 12439 16574 12451
rect 16478 12379 16506 12439
rect 16540 12379 16574 12439
rect 16478 12367 16574 12379
rect 16604 12439 16662 12451
rect 16604 12379 16616 12439
rect 16650 12379 16662 12439
rect 16604 12367 16662 12379
rect 17602 12439 17660 12451
rect 17602 12379 17614 12439
rect 17648 12379 17660 12439
rect 17602 12367 17660 12379
rect 17690 12439 17786 12451
rect 17690 12379 17719 12439
rect 17753 12379 17786 12439
rect 17690 12367 17786 12379
rect 17816 12439 17874 12451
rect 17816 12379 17828 12439
rect 17862 12379 17874 12439
rect 17816 12367 17874 12379
rect 18814 12439 18872 12451
rect 18814 12379 18826 12439
rect 18860 12379 18872 12439
rect 18814 12367 18872 12379
rect 18902 12439 18998 12451
rect 18902 12379 18933 12439
rect 18967 12379 18998 12439
rect 18902 12367 18998 12379
rect 19028 12439 19086 12451
rect 19028 12379 19040 12439
rect 19074 12379 19086 12439
rect 19028 12367 19086 12379
rect 19589 12442 19647 12454
rect 19589 12382 19601 12442
rect 19635 12382 19647 12442
rect 19589 12370 19647 12382
rect 19677 12442 19739 12454
rect 19677 12382 19689 12442
rect 19723 12382 19739 12442
rect 19677 12370 19739 12382
rect 19769 12442 19835 12454
rect 19769 12382 19785 12442
rect 19819 12382 19835 12442
rect 19769 12370 19835 12382
rect 19865 12442 19927 12454
rect 19865 12382 19881 12442
rect 19915 12382 19927 12442
rect 21155 12436 21213 12448
rect 19865 12370 19927 12382
rect 21155 12376 21167 12436
rect 21201 12376 21213 12436
rect 21155 12364 21213 12376
rect 21243 12439 21301 12448
rect 21243 12379 21255 12439
rect 21289 12379 21301 12439
rect 21243 12364 21301 12379
rect 21887 12439 21945 12451
rect 21887 12379 21899 12439
rect 21933 12379 21945 12439
rect 21887 12367 21945 12379
rect 21975 12439 22071 12451
rect 21975 12379 22004 12439
rect 22038 12379 22071 12439
rect 21975 12367 22071 12379
rect 22101 12439 22159 12451
rect 22101 12379 22113 12439
rect 22147 12379 22159 12439
rect 22101 12367 22159 12379
rect 23099 12439 23157 12451
rect 23099 12379 23111 12439
rect 23145 12379 23157 12439
rect 23099 12367 23157 12379
rect 23187 12439 23283 12451
rect 23187 12379 23215 12439
rect 23249 12379 23283 12439
rect 23187 12367 23283 12379
rect 23313 12439 23371 12451
rect 23313 12379 23325 12439
rect 23359 12379 23371 12439
rect 23313 12367 23371 12379
rect 24311 12439 24369 12451
rect 24311 12379 24323 12439
rect 24357 12379 24369 12439
rect 24311 12367 24369 12379
rect 24399 12439 24495 12451
rect 24399 12379 24428 12439
rect 24462 12379 24495 12439
rect 24399 12367 24495 12379
rect 24525 12439 24583 12451
rect 24525 12379 24537 12439
rect 24571 12379 24583 12439
rect 24525 12367 24583 12379
rect 25523 12439 25581 12451
rect 25523 12379 25535 12439
rect 25569 12379 25581 12439
rect 25523 12367 25581 12379
rect 25611 12439 25707 12451
rect 25611 12379 25642 12439
rect 25676 12379 25707 12439
rect 25611 12367 25707 12379
rect 25737 12439 25795 12451
rect 25737 12379 25749 12439
rect 25783 12379 25795 12439
rect 25737 12367 25795 12379
rect 26298 12442 26356 12454
rect 26298 12382 26310 12442
rect 26344 12382 26356 12442
rect 26298 12370 26356 12382
rect 26386 12442 26448 12454
rect 26386 12382 26398 12442
rect 26432 12382 26448 12442
rect 26386 12370 26448 12382
rect 26478 12442 26544 12454
rect 26478 12382 26494 12442
rect 26528 12382 26544 12442
rect 26478 12370 26544 12382
rect 26574 12442 26636 12454
rect 26574 12382 26590 12442
rect 26624 12382 26636 12442
rect 26574 12370 26636 12382
rect 12832 12148 12882 12152
rect 12733 12134 12785 12148
rect 12464 12036 12515 12120
rect 11995 11952 12109 12036
rect 12139 11999 12193 12036
rect 12139 11965 12149 11999
rect 12183 11965 12193 11999
rect 12139 11952 12193 11965
rect 12223 11952 12311 12036
rect 12341 11998 12419 12036
rect 12341 11964 12363 11998
rect 12397 11964 12419 11998
rect 12341 11952 12419 11964
rect 12449 12024 12515 12036
rect 12449 11990 12471 12024
rect 12505 11990 12515 12024
rect 12449 11952 12515 11990
rect 12545 11952 12587 12120
rect 12617 11998 12669 12120
rect 12733 12100 12741 12134
rect 12775 12100 12785 12134
rect 12733 12020 12785 12100
rect 12815 12020 12882 12148
rect 12617 11964 12627 11998
rect 12661 11964 12669 11998
rect 12830 11998 12882 12020
rect 12617 11952 12669 11964
rect 12830 11964 12838 11998
rect 12872 11964 12882 11998
rect 12830 11952 12882 11964
rect 12912 12103 12964 12152
rect 12912 12069 12922 12103
rect 12956 12069 12964 12103
rect 13115 12096 13165 12152
rect 12912 12035 12964 12069
rect 12912 12001 12922 12035
rect 12956 12001 12964 12035
rect 12912 11952 12964 12001
rect 13018 12084 13070 12096
rect 13018 12050 13026 12084
rect 13060 12050 13070 12084
rect 13018 12016 13070 12050
rect 13018 11982 13026 12016
rect 13060 11982 13070 12016
rect 13018 11968 13070 11982
rect 13100 12078 13165 12096
rect 13100 12044 13121 12078
rect 13155 12044 13165 12078
rect 13100 12010 13165 12044
rect 13100 11976 13121 12010
rect 13155 11976 13165 12010
rect 13100 11968 13165 11976
rect 13115 11952 13165 11968
rect 13195 12102 13247 12152
rect 13195 12068 13205 12102
rect 13239 12068 13247 12102
rect 13195 12034 13247 12068
rect 13195 12000 13205 12034
rect 13239 12000 13247 12034
rect 13195 11952 13247 12000
rect 9211 11894 9263 11912
rect 10950 11750 11002 11762
rect 10950 11716 10958 11750
rect 10992 11716 11002 11750
rect 10950 11682 11002 11716
rect 10950 11648 10958 11682
rect 10992 11648 11002 11682
rect 10950 11614 11002 11648
rect 10950 11580 10958 11614
rect 10992 11580 11002 11614
rect 10950 11562 11002 11580
rect 11032 11750 11084 11762
rect 11032 11716 11042 11750
rect 11076 11716 11084 11750
rect 11032 11682 11084 11716
rect 11032 11648 11042 11682
rect 11076 11648 11084 11682
rect 11032 11614 11084 11648
rect 11032 11580 11042 11614
rect 11076 11580 11084 11614
rect 11032 11562 11084 11580
rect 11226 11750 11278 11762
rect 11226 11716 11234 11750
rect 11268 11716 11278 11750
rect 11226 11682 11278 11716
rect 11226 11648 11234 11682
rect 11268 11648 11278 11682
rect 11226 11614 11278 11648
rect 11226 11580 11234 11614
rect 11268 11580 11278 11614
rect 11226 11562 11278 11580
rect 11308 11750 11360 11762
rect 11308 11716 11318 11750
rect 11352 11716 11360 11750
rect 11308 11682 11360 11716
rect 11308 11648 11318 11682
rect 11352 11648 11360 11682
rect 11308 11614 11360 11648
rect 11308 11580 11318 11614
rect 11352 11580 11360 11614
rect 11308 11562 11360 11580
rect 3558 8745 3616 8757
rect 3558 8685 3570 8745
rect 3604 8685 3616 8745
rect 3558 8673 3616 8685
rect 3646 8742 3704 8757
rect 3646 8682 3658 8742
rect 3692 8682 3704 8742
rect 3646 8673 3704 8682
rect 4290 8742 4348 8754
rect 4290 8682 4302 8742
rect 4336 8682 4348 8742
rect 4290 8670 4348 8682
rect 4378 8742 4474 8754
rect 4378 8682 4407 8742
rect 4441 8682 4474 8742
rect 4378 8670 4474 8682
rect 4504 8742 4562 8754
rect 4504 8682 4516 8742
rect 4550 8682 4562 8742
rect 4504 8670 4562 8682
rect 5502 8742 5560 8754
rect 5502 8682 5514 8742
rect 5548 8682 5560 8742
rect 5502 8670 5560 8682
rect 5590 8742 5686 8754
rect 5590 8682 5618 8742
rect 5652 8682 5686 8742
rect 5590 8670 5686 8682
rect 5716 8742 5774 8754
rect 5716 8682 5728 8742
rect 5762 8682 5774 8742
rect 5716 8670 5774 8682
rect 6714 8742 6772 8754
rect 6714 8682 6726 8742
rect 6760 8682 6772 8742
rect 6714 8670 6772 8682
rect 6802 8742 6898 8754
rect 6802 8682 6831 8742
rect 6865 8682 6898 8742
rect 6802 8670 6898 8682
rect 6928 8742 6986 8754
rect 6928 8682 6940 8742
rect 6974 8682 6986 8742
rect 6928 8670 6986 8682
rect 7926 8742 7984 8754
rect 7926 8682 7938 8742
rect 7972 8682 7984 8742
rect 7926 8670 7984 8682
rect 8014 8742 8110 8754
rect 8014 8682 8045 8742
rect 8079 8682 8110 8742
rect 8014 8670 8110 8682
rect 8140 8742 8198 8754
rect 8140 8682 8152 8742
rect 8186 8682 8198 8742
rect 8140 8670 8198 8682
rect 8701 8739 8759 8751
rect 8701 8679 8713 8739
rect 8747 8679 8759 8739
rect 8701 8667 8759 8679
rect 8789 8739 8851 8751
rect 8789 8679 8801 8739
rect 8835 8679 8851 8739
rect 8789 8667 8851 8679
rect 8881 8739 8947 8751
rect 8881 8679 8897 8739
rect 8931 8679 8947 8739
rect 8881 8667 8947 8679
rect 8977 8739 9039 8751
rect 8977 8679 8993 8739
rect 9027 8679 9039 8739
rect 8977 8667 9039 8679
rect 9129 8736 9181 8754
rect 9129 8702 9137 8736
rect 9171 8702 9181 8736
rect 9129 8668 9181 8702
rect 9129 8634 9137 8668
rect 9171 8634 9181 8668
rect 8701 8601 8759 8613
rect 8701 8541 8713 8601
rect 8747 8541 8759 8601
rect 8701 8529 8759 8541
rect 8789 8601 8847 8613
rect 8789 8541 8801 8601
rect 8835 8541 8847 8601
rect 9129 8600 9181 8634
rect 9129 8566 9137 8600
rect 9171 8566 9181 8600
rect 9129 8554 9181 8566
rect 9211 8736 9263 8754
rect 9211 8702 9221 8736
rect 9255 8702 9263 8736
rect 9211 8668 9263 8702
rect 9211 8634 9221 8668
rect 9255 8634 9263 8668
rect 9211 8600 9263 8634
rect 9211 8566 9221 8600
rect 9255 8566 9263 8600
rect 9211 8554 9263 8566
rect 9344 8704 9396 8754
rect 9344 8670 9352 8704
rect 9386 8670 9396 8704
rect 9344 8636 9396 8670
rect 9344 8602 9352 8636
rect 9386 8602 9396 8636
rect 9344 8554 9396 8602
rect 9426 8698 9476 8754
rect 9627 8705 9679 8754
rect 9426 8680 9491 8698
rect 9426 8646 9436 8680
rect 9470 8646 9491 8680
rect 9426 8612 9491 8646
rect 9426 8578 9436 8612
rect 9470 8578 9491 8612
rect 9426 8570 9491 8578
rect 9521 8686 9573 8698
rect 9521 8652 9531 8686
rect 9565 8652 9573 8686
rect 9521 8618 9573 8652
rect 9521 8584 9531 8618
rect 9565 8584 9573 8618
rect 9521 8570 9573 8584
rect 9627 8671 9635 8705
rect 9669 8671 9679 8705
rect 9627 8637 9679 8671
rect 9627 8603 9635 8637
rect 9669 8603 9679 8637
rect 9426 8554 9476 8570
rect 8789 8529 8847 8541
rect 9627 8554 9679 8603
rect 9709 8750 9759 8754
rect 9709 8622 9776 8750
rect 9806 8736 9858 8750
rect 9806 8702 9816 8736
rect 9850 8702 9858 8736
rect 9806 8622 9858 8702
rect 9709 8600 9761 8622
rect 9709 8566 9719 8600
rect 9753 8566 9761 8600
rect 9922 8600 9974 8722
rect 9709 8554 9761 8566
rect 9922 8566 9930 8600
rect 9964 8566 9974 8600
rect 9922 8554 9974 8566
rect 10004 8554 10046 8722
rect 10076 8638 10127 8722
rect 10544 8638 10596 8722
rect 10076 8626 10142 8638
rect 10076 8592 10086 8626
rect 10120 8592 10142 8626
rect 10076 8554 10142 8592
rect 10172 8600 10250 8638
rect 10172 8566 10194 8600
rect 10228 8566 10250 8600
rect 10172 8554 10250 8566
rect 10280 8554 10368 8638
rect 10398 8601 10452 8638
rect 10398 8567 10408 8601
rect 10442 8567 10452 8601
rect 10398 8554 10452 8567
rect 10482 8554 10596 8638
rect 10626 8668 10733 8722
rect 10626 8634 10683 8668
rect 10717 8634 10733 8668
rect 10626 8600 10733 8634
rect 10626 8566 10683 8600
rect 10717 8566 10733 8600
rect 10626 8554 10733 8566
rect 10763 8554 10817 8722
rect 10847 8694 10909 8722
rect 10847 8660 10857 8694
rect 10891 8660 10909 8694
rect 10847 8638 10909 8660
rect 11821 8728 11883 8740
rect 11464 8676 11516 8688
rect 11464 8642 11472 8676
rect 11506 8642 11516 8676
rect 10847 8626 10925 8638
rect 10847 8592 10857 8626
rect 10891 8592 10925 8626
rect 10847 8554 10925 8592
rect 10955 8610 11031 8638
rect 10955 8576 10977 8610
rect 11011 8576 11031 8610
rect 10955 8554 11031 8576
rect 11061 8554 11151 8638
rect 11181 8601 11235 8638
rect 11181 8567 11191 8601
rect 11225 8567 11235 8601
rect 11181 8554 11235 8567
rect 11265 8608 11328 8638
rect 11265 8574 11284 8608
rect 11318 8574 11328 8608
rect 11265 8554 11328 8574
rect 11358 8624 11410 8638
rect 11358 8590 11368 8624
rect 11402 8590 11410 8624
rect 11358 8554 11410 8590
rect 11464 8608 11516 8642
rect 11464 8574 11472 8608
rect 11506 8574 11516 8608
rect 11464 8560 11516 8574
rect 11546 8624 11600 8688
rect 11546 8590 11556 8624
rect 11590 8590 11600 8624
rect 11546 8560 11600 8590
rect 11630 8676 11682 8688
rect 11630 8642 11640 8676
rect 11674 8642 11682 8676
rect 11630 8608 11682 8642
rect 11630 8574 11640 8608
rect 11674 8574 11682 8608
rect 11630 8560 11682 8574
rect 11821 8500 11833 8728
rect 11867 8500 11883 8728
rect 11821 8488 11883 8500
rect 11913 8728 11979 8740
rect 11913 8500 11929 8728
rect 11963 8500 11979 8728
rect 11913 8488 11979 8500
rect 12009 8728 12075 8740
rect 12009 8500 12025 8728
rect 12059 8500 12075 8728
rect 12009 8488 12075 8500
rect 12105 8728 12167 8740
rect 12105 8500 12121 8728
rect 12155 8500 12167 8728
rect 12105 8488 12167 8500
rect 12221 8729 12279 8741
rect 12221 8501 12233 8729
rect 12267 8501 12279 8729
rect 12221 8489 12279 8501
rect 12309 8729 12367 8741
rect 12309 8501 12321 8729
rect 12355 8501 12367 8729
rect 12309 8489 12367 8501
rect 12422 8728 12480 8740
rect 12422 8472 12434 8728
rect 12468 8472 12480 8728
rect 12422 8460 12480 8472
rect 12510 8728 12568 8740
rect 12510 8472 12522 8728
rect 12556 8472 12568 8728
rect 12676 8723 12728 8741
rect 12676 8689 12684 8723
rect 12718 8689 12728 8723
rect 12676 8655 12728 8689
rect 12676 8621 12684 8655
rect 12718 8621 12728 8655
rect 12676 8587 12728 8621
rect 12676 8553 12684 8587
rect 12718 8553 12728 8587
rect 12676 8541 12728 8553
rect 12758 8723 12812 8741
rect 12758 8689 12768 8723
rect 12802 8689 12812 8723
rect 12758 8655 12812 8689
rect 12758 8621 12768 8655
rect 12802 8621 12812 8655
rect 12758 8587 12812 8621
rect 12758 8553 12768 8587
rect 12802 8553 12812 8587
rect 12758 8541 12812 8553
rect 12842 8723 12894 8741
rect 12842 8689 12852 8723
rect 12886 8689 12894 8723
rect 12842 8655 12894 8689
rect 12842 8621 12852 8655
rect 12886 8621 12894 8655
rect 12842 8587 12894 8621
rect 12842 8553 12852 8587
rect 12886 8553 12894 8587
rect 12842 8541 12894 8553
rect 12999 8723 13051 8741
rect 12999 8689 13007 8723
rect 13041 8689 13051 8723
rect 12999 8655 13051 8689
rect 12999 8621 13007 8655
rect 13041 8621 13051 8655
rect 12999 8587 13051 8621
rect 12999 8553 13007 8587
rect 13041 8553 13051 8587
rect 12999 8541 13051 8553
rect 13081 8723 13133 8741
rect 13081 8689 13091 8723
rect 13125 8689 13133 8723
rect 13081 8655 13133 8689
rect 13252 8727 13314 8739
rect 13252 8667 13264 8727
rect 13298 8667 13314 8727
rect 13252 8655 13314 8667
rect 13344 8727 13410 8739
rect 13344 8667 13360 8727
rect 13394 8667 13410 8727
rect 13344 8655 13410 8667
rect 13440 8727 13502 8739
rect 13440 8667 13456 8727
rect 13490 8667 13502 8727
rect 13440 8655 13502 8667
rect 13532 8727 13590 8739
rect 13532 8667 13544 8727
rect 13578 8667 13590 8727
rect 13532 8655 13590 8667
rect 14093 8730 14151 8742
rect 14093 8670 14105 8730
rect 14139 8670 14151 8730
rect 14093 8658 14151 8670
rect 14181 8730 14277 8742
rect 14181 8670 14212 8730
rect 14246 8670 14277 8730
rect 14181 8658 14277 8670
rect 14307 8730 14365 8742
rect 14307 8670 14319 8730
rect 14353 8670 14365 8730
rect 14307 8658 14365 8670
rect 15305 8730 15363 8742
rect 15305 8670 15317 8730
rect 15351 8670 15363 8730
rect 15305 8658 15363 8670
rect 15393 8730 15489 8742
rect 15393 8670 15426 8730
rect 15460 8670 15489 8730
rect 15393 8658 15489 8670
rect 15519 8730 15577 8742
rect 15519 8670 15531 8730
rect 15565 8670 15577 8730
rect 15519 8658 15577 8670
rect 16517 8730 16575 8742
rect 16517 8670 16529 8730
rect 16563 8670 16575 8730
rect 16517 8658 16575 8670
rect 16605 8730 16701 8742
rect 16605 8670 16639 8730
rect 16673 8670 16701 8730
rect 16605 8658 16701 8670
rect 16731 8730 16789 8742
rect 16731 8670 16743 8730
rect 16777 8670 16789 8730
rect 16731 8658 16789 8670
rect 17729 8730 17787 8742
rect 17729 8670 17741 8730
rect 17775 8670 17787 8730
rect 17729 8658 17787 8670
rect 17817 8730 17913 8742
rect 17817 8670 17850 8730
rect 17884 8670 17913 8730
rect 17817 8658 17913 8670
rect 17943 8730 18001 8742
rect 17943 8670 17955 8730
rect 17989 8670 18001 8730
rect 17943 8658 18001 8670
rect 18587 8730 18645 8745
rect 18587 8670 18599 8730
rect 18633 8670 18645 8730
rect 18587 8661 18645 8670
rect 18675 8733 18733 8745
rect 18675 8673 18687 8733
rect 18721 8673 18733 8733
rect 19961 8727 20023 8739
rect 18675 8661 18733 8673
rect 19961 8667 19973 8727
rect 20007 8667 20023 8727
rect 13081 8621 13091 8655
rect 13125 8621 13133 8655
rect 13081 8587 13133 8621
rect 19961 8655 20023 8667
rect 20053 8727 20119 8739
rect 20053 8667 20069 8727
rect 20103 8667 20119 8727
rect 20053 8655 20119 8667
rect 20149 8727 20211 8739
rect 20149 8667 20165 8727
rect 20199 8667 20211 8727
rect 20149 8655 20211 8667
rect 20241 8727 20299 8739
rect 20241 8667 20253 8727
rect 20287 8667 20299 8727
rect 20241 8655 20299 8667
rect 20802 8730 20860 8742
rect 20802 8670 20814 8730
rect 20848 8670 20860 8730
rect 20802 8658 20860 8670
rect 20890 8730 20986 8742
rect 20890 8670 20921 8730
rect 20955 8670 20986 8730
rect 20890 8658 20986 8670
rect 21016 8730 21074 8742
rect 21016 8670 21028 8730
rect 21062 8670 21074 8730
rect 21016 8658 21074 8670
rect 22014 8730 22072 8742
rect 22014 8670 22026 8730
rect 22060 8670 22072 8730
rect 22014 8658 22072 8670
rect 22102 8730 22198 8742
rect 22102 8670 22135 8730
rect 22169 8670 22198 8730
rect 22102 8658 22198 8670
rect 22228 8730 22286 8742
rect 22228 8670 22240 8730
rect 22274 8670 22286 8730
rect 22228 8658 22286 8670
rect 23226 8730 23284 8742
rect 23226 8670 23238 8730
rect 23272 8670 23284 8730
rect 23226 8658 23284 8670
rect 23314 8730 23410 8742
rect 23314 8670 23348 8730
rect 23382 8670 23410 8730
rect 23314 8658 23410 8670
rect 23440 8730 23498 8742
rect 23440 8670 23452 8730
rect 23486 8670 23498 8730
rect 23440 8658 23498 8670
rect 24438 8730 24496 8742
rect 24438 8670 24450 8730
rect 24484 8670 24496 8730
rect 24438 8658 24496 8670
rect 24526 8730 24622 8742
rect 24526 8670 24559 8730
rect 24593 8670 24622 8730
rect 24526 8658 24622 8670
rect 24652 8730 24710 8742
rect 24652 8670 24664 8730
rect 24698 8670 24710 8730
rect 24652 8658 24710 8670
rect 25296 8730 25354 8745
rect 25296 8670 25308 8730
rect 25342 8670 25354 8730
rect 25296 8661 25354 8670
rect 25384 8733 25442 8745
rect 25384 8673 25396 8733
rect 25430 8673 25442 8733
rect 25384 8661 25442 8673
rect 13081 8553 13091 8587
rect 13125 8553 13133 8587
rect 13081 8541 13133 8553
rect 13444 8589 13502 8601
rect 13444 8529 13456 8589
rect 13490 8529 13502 8589
rect 13444 8517 13502 8529
rect 13532 8589 13590 8601
rect 13532 8529 13544 8589
rect 13578 8529 13590 8589
rect 13532 8517 13590 8529
rect 20153 8589 20211 8601
rect 20153 8529 20165 8589
rect 20199 8529 20211 8589
rect 20153 8517 20211 8529
rect 20241 8589 20299 8601
rect 20241 8529 20253 8589
rect 20287 8529 20299 8589
rect 20241 8517 20299 8529
rect 12510 8460 12568 8472
rect 2454 8357 2506 8375
rect 2454 8323 2462 8357
rect 2496 8323 2506 8357
rect 2454 8289 2506 8323
rect 2454 8255 2462 8289
rect 2496 8255 2506 8289
rect 2454 8221 2506 8255
rect 2454 8187 2462 8221
rect 2496 8187 2506 8221
rect 2454 8175 2506 8187
rect 2536 8357 2588 8375
rect 2536 8323 2546 8357
rect 2580 8323 2588 8357
rect 2536 8289 2588 8323
rect 2536 8255 2546 8289
rect 2580 8255 2588 8289
rect 2536 8221 2588 8255
rect 2536 8187 2546 8221
rect 2580 8187 2588 8221
rect 2536 8175 2588 8187
rect 2644 8357 2696 8375
rect 2644 8323 2652 8357
rect 2686 8323 2696 8357
rect 2644 8289 2696 8323
rect 2644 8255 2652 8289
rect 2686 8255 2696 8289
rect 2644 8221 2696 8255
rect 2644 8187 2652 8221
rect 2686 8187 2696 8221
rect 2644 8175 2696 8187
rect 2726 8357 2778 8375
rect 2726 8323 2736 8357
rect 2770 8323 2778 8357
rect 2726 8289 2778 8323
rect 11821 8324 11883 8336
rect 2726 8255 2736 8289
rect 2770 8255 2778 8289
rect 2726 8221 2778 8255
rect 2726 8187 2736 8221
rect 2770 8187 2778 8221
rect 2916 8290 2974 8302
rect 2916 8230 2928 8290
rect 2962 8230 2974 8290
rect 2916 8218 2974 8230
rect 3004 8290 3062 8302
rect 3004 8230 3016 8290
rect 3050 8230 3062 8290
rect 10081 8273 10133 8285
rect 3004 8218 3062 8230
rect 2726 8175 2778 8187
rect 2916 8152 2974 8164
rect 2916 8092 2928 8152
rect 2962 8092 2974 8152
rect 2916 8080 2974 8092
rect 3004 8152 3062 8164
rect 10081 8239 10089 8273
rect 10123 8239 10133 8273
rect 10081 8205 10133 8239
rect 10081 8171 10089 8205
rect 10123 8171 10133 8205
rect 3004 8092 3016 8152
rect 3050 8092 3062 8152
rect 3004 8080 3062 8092
rect 10081 8137 10133 8171
rect 10081 8103 10089 8137
rect 10123 8103 10133 8137
rect 10081 8085 10133 8103
rect 10163 8273 10215 8285
rect 10163 8239 10173 8273
rect 10207 8246 10215 8273
rect 10908 8273 10960 8285
rect 10207 8239 10242 8246
rect 10163 8205 10242 8239
rect 10163 8171 10173 8205
rect 10207 8171 10242 8205
rect 10163 8162 10242 8171
rect 10272 8162 10345 8246
rect 10375 8213 10559 8246
rect 10375 8179 10409 8213
rect 10443 8179 10484 8213
rect 10518 8179 10559 8213
rect 10375 8162 10559 8179
rect 10589 8162 10631 8246
rect 10661 8213 10727 8246
rect 10661 8179 10681 8213
rect 10715 8179 10727 8213
rect 10661 8162 10727 8179
rect 10757 8213 10813 8246
rect 10757 8179 10767 8213
rect 10801 8179 10813 8213
rect 10757 8162 10813 8179
rect 10908 8239 10916 8273
rect 10950 8239 10960 8273
rect 10908 8205 10960 8239
rect 10908 8171 10916 8205
rect 10950 8171 10960 8205
rect 10163 8137 10215 8162
rect 10163 8103 10173 8137
rect 10207 8103 10215 8137
rect 10163 8085 10215 8103
rect 2916 8014 2974 8026
rect 2916 7954 2928 8014
rect 2962 7954 2974 8014
rect 2916 7942 2974 7954
rect 3004 8014 3062 8026
rect 3004 7954 3016 8014
rect 3050 7954 3062 8014
rect 3004 7942 3062 7954
rect 2916 7876 2974 7888
rect 2916 7816 2928 7876
rect 2962 7816 2974 7876
rect 2916 7804 2974 7816
rect 3004 7876 3062 7888
rect 3004 7816 3016 7876
rect 3050 7816 3062 7876
rect 10908 8137 10960 8171
rect 10908 8103 10916 8137
rect 10950 8103 10960 8137
rect 10908 8085 10960 8103
rect 10990 8273 11042 8285
rect 10990 8239 11000 8273
rect 11034 8246 11042 8273
rect 11034 8239 11069 8246
rect 10990 8205 11069 8239
rect 10990 8171 11000 8205
rect 11034 8171 11069 8205
rect 10990 8162 11069 8171
rect 11099 8162 11172 8246
rect 11202 8213 11386 8246
rect 11202 8179 11236 8213
rect 11270 8179 11311 8213
rect 11345 8179 11386 8213
rect 11202 8162 11386 8179
rect 11416 8162 11458 8246
rect 11488 8213 11554 8246
rect 11488 8179 11508 8213
rect 11542 8179 11554 8213
rect 11488 8162 11554 8179
rect 11584 8213 11640 8246
rect 11584 8179 11594 8213
rect 11628 8179 11640 8213
rect 11584 8162 11640 8179
rect 10990 8137 11042 8162
rect 10990 8103 11000 8137
rect 11034 8103 11042 8137
rect 10990 8085 11042 8103
rect 11821 8096 11833 8324
rect 11867 8096 11883 8324
rect 11821 8084 11883 8096
rect 11913 8324 11979 8336
rect 11913 8096 11929 8324
rect 11963 8096 11979 8324
rect 11913 8084 11979 8096
rect 12009 8324 12075 8336
rect 12009 8096 12025 8324
rect 12059 8096 12075 8324
rect 12009 8084 12075 8096
rect 12105 8324 12167 8336
rect 12105 8096 12121 8324
rect 12155 8096 12167 8324
rect 12105 8084 12167 8096
rect 12221 8323 12279 8335
rect 12221 8095 12233 8323
rect 12267 8095 12279 8323
rect 12221 8083 12279 8095
rect 12309 8323 12367 8335
rect 12309 8095 12321 8323
rect 12355 8095 12367 8323
rect 19513 8345 19565 8363
rect 19513 8311 19521 8345
rect 19555 8311 19565 8345
rect 19229 8278 19287 8290
rect 19229 8218 19241 8278
rect 19275 8218 19287 8278
rect 19229 8206 19287 8218
rect 19317 8278 19375 8290
rect 19317 8218 19329 8278
rect 19363 8218 19375 8278
rect 19317 8206 19375 8218
rect 19513 8277 19565 8311
rect 19513 8243 19521 8277
rect 19555 8243 19565 8277
rect 19513 8209 19565 8243
rect 12309 8083 12367 8095
rect 19513 8175 19521 8209
rect 19555 8175 19565 8209
rect 19513 8163 19565 8175
rect 19595 8345 19647 8363
rect 19595 8311 19605 8345
rect 19639 8311 19647 8345
rect 19595 8277 19647 8311
rect 19595 8243 19605 8277
rect 19639 8243 19647 8277
rect 19595 8209 19647 8243
rect 19595 8175 19605 8209
rect 19639 8175 19647 8209
rect 19595 8163 19647 8175
rect 19703 8345 19755 8363
rect 19703 8311 19711 8345
rect 19745 8311 19755 8345
rect 19703 8277 19755 8311
rect 19703 8243 19711 8277
rect 19745 8243 19755 8277
rect 19703 8209 19755 8243
rect 19703 8175 19711 8209
rect 19745 8175 19755 8209
rect 19703 8163 19755 8175
rect 19785 8345 19837 8363
rect 19785 8311 19795 8345
rect 19829 8311 19837 8345
rect 26222 8345 26274 8363
rect 19785 8277 19837 8311
rect 26222 8311 26230 8345
rect 26264 8311 26274 8345
rect 19785 8243 19795 8277
rect 19829 8243 19837 8277
rect 19785 8209 19837 8243
rect 25938 8278 25996 8290
rect 19785 8175 19795 8209
rect 19829 8175 19837 8209
rect 19785 8163 19837 8175
rect 25938 8218 25950 8278
rect 25984 8218 25996 8278
rect 25938 8206 25996 8218
rect 26026 8278 26084 8290
rect 26026 8218 26038 8278
rect 26072 8218 26084 8278
rect 26026 8206 26084 8218
rect 26222 8277 26274 8311
rect 26222 8243 26230 8277
rect 26264 8243 26274 8277
rect 26222 8209 26274 8243
rect 19229 8140 19287 8152
rect 19229 8080 19241 8140
rect 19275 8080 19287 8140
rect 19229 8068 19287 8080
rect 19317 8140 19375 8152
rect 19317 8080 19329 8140
rect 19363 8080 19375 8140
rect 26222 8175 26230 8209
rect 26264 8175 26274 8209
rect 26222 8163 26274 8175
rect 26304 8345 26356 8363
rect 26304 8311 26314 8345
rect 26348 8311 26356 8345
rect 26304 8277 26356 8311
rect 26304 8243 26314 8277
rect 26348 8243 26356 8277
rect 26304 8209 26356 8243
rect 26304 8175 26314 8209
rect 26348 8175 26356 8209
rect 26304 8163 26356 8175
rect 26412 8345 26464 8363
rect 26412 8311 26420 8345
rect 26454 8311 26464 8345
rect 26412 8277 26464 8311
rect 26412 8243 26420 8277
rect 26454 8243 26464 8277
rect 26412 8209 26464 8243
rect 26412 8175 26420 8209
rect 26454 8175 26464 8209
rect 26412 8163 26464 8175
rect 26494 8345 26546 8363
rect 26494 8311 26504 8345
rect 26538 8311 26546 8345
rect 26494 8277 26546 8311
rect 26494 8243 26504 8277
rect 26538 8243 26546 8277
rect 26494 8209 26546 8243
rect 26494 8175 26504 8209
rect 26538 8175 26546 8209
rect 26494 8163 26546 8175
rect 25938 8140 25996 8152
rect 19317 8068 19375 8080
rect 25938 8080 25950 8140
rect 25984 8080 25996 8140
rect 25938 8068 25996 8080
rect 26026 8140 26084 8152
rect 26026 8080 26038 8140
rect 26072 8080 26084 8140
rect 26026 8068 26084 8080
rect 19229 8002 19287 8014
rect 12690 7952 12748 7964
rect 3004 7804 3062 7816
rect 2916 7738 2974 7750
rect 2916 7678 2928 7738
rect 2962 7678 2974 7738
rect 2916 7666 2974 7678
rect 3004 7738 3062 7750
rect 3004 7678 3016 7738
rect 3050 7678 3062 7738
rect 3004 7666 3062 7678
rect 2916 7600 2974 7612
rect 2916 7540 2928 7600
rect 2962 7540 2974 7600
rect 2916 7528 2974 7540
rect 3004 7600 3062 7612
rect 3004 7540 3016 7600
rect 3050 7540 3062 7600
rect 12690 7596 12702 7952
rect 12736 7596 12748 7952
rect 12690 7584 12748 7596
rect 12778 7952 12836 7964
rect 12778 7596 12790 7952
rect 12824 7596 12836 7952
rect 19229 7942 19241 8002
rect 19275 7942 19287 8002
rect 19229 7930 19287 7942
rect 19317 8002 19375 8014
rect 19317 7942 19329 8002
rect 19363 7942 19375 8002
rect 19317 7930 19375 7942
rect 25938 8002 25996 8014
rect 25938 7942 25950 8002
rect 25984 7942 25996 8002
rect 25938 7930 25996 7942
rect 26026 8002 26084 8014
rect 26026 7942 26038 8002
rect 26072 7942 26084 8002
rect 26026 7930 26084 7942
rect 19229 7864 19287 7876
rect 19229 7804 19241 7864
rect 19275 7804 19287 7864
rect 19229 7792 19287 7804
rect 19317 7864 19375 7876
rect 19317 7804 19329 7864
rect 19363 7804 19375 7864
rect 25938 7864 25996 7876
rect 19317 7792 19375 7804
rect 25938 7804 25950 7864
rect 25984 7804 25996 7864
rect 25938 7792 25996 7804
rect 26026 7864 26084 7876
rect 26026 7804 26038 7864
rect 26072 7804 26084 7864
rect 26026 7792 26084 7804
rect 19229 7726 19287 7738
rect 19229 7666 19241 7726
rect 19275 7666 19287 7726
rect 19229 7654 19287 7666
rect 19317 7726 19375 7738
rect 19317 7666 19329 7726
rect 19363 7666 19375 7726
rect 19317 7654 19375 7666
rect 25938 7726 25996 7738
rect 25938 7666 25950 7726
rect 25984 7666 25996 7726
rect 25938 7654 25996 7666
rect 26026 7726 26084 7738
rect 26026 7666 26038 7726
rect 26072 7666 26084 7726
rect 26026 7654 26084 7666
rect 12778 7584 12836 7596
rect 3004 7528 3062 7540
rect 19229 7588 19287 7600
rect 19229 7528 19241 7588
rect 19275 7528 19287 7588
rect 19229 7516 19287 7528
rect 19317 7588 19375 7600
rect 19317 7528 19329 7588
rect 19363 7528 19375 7588
rect 25938 7588 25996 7600
rect 19317 7516 19375 7528
rect 25938 7528 25950 7588
rect 25984 7528 25996 7588
rect 25938 7516 25996 7528
rect 26026 7588 26084 7600
rect 26026 7528 26038 7588
rect 26072 7528 26084 7588
rect 26026 7516 26084 7528
rect 24529 7284 24587 7296
rect 24529 7224 24541 7284
rect 24575 7224 24587 7284
rect 24529 7212 24587 7224
rect 24617 7284 24675 7296
rect 24617 7224 24629 7284
rect 24663 7224 24675 7284
rect 24617 7212 24675 7224
rect 24529 7146 24587 7158
rect 24529 7086 24541 7146
rect 24575 7086 24587 7146
rect 24529 7074 24587 7086
rect 24617 7146 24675 7158
rect 24617 7086 24629 7146
rect 24663 7086 24675 7146
rect 24617 7074 24675 7086
rect 11525 7010 11577 7030
rect 11525 6976 11533 7010
rect 11567 6976 11577 7010
rect 11525 6942 11577 6976
rect 11525 6908 11533 6942
rect 11567 6908 11577 6942
rect 11525 6872 11577 6908
rect 11607 7010 11665 7030
rect 11607 6976 11619 7010
rect 11653 6976 11665 7010
rect 11607 6942 11665 6976
rect 11607 6908 11619 6942
rect 11653 6908 11665 6942
rect 11607 6872 11665 6908
rect 11695 7010 11747 7030
rect 11695 6976 11705 7010
rect 11739 6976 11747 7010
rect 11695 6929 11747 6976
rect 11695 6895 11705 6929
rect 11739 6895 11747 6929
rect 11695 6872 11747 6895
rect 11801 7012 11853 7030
rect 11801 6978 11809 7012
rect 11843 6978 11853 7012
rect 11801 6944 11853 6978
rect 11801 6910 11809 6944
rect 11843 6910 11853 6944
rect 11801 6876 11853 6910
rect 11801 6842 11809 6876
rect 11843 6842 11853 6876
rect 11801 6830 11853 6842
rect 11883 7018 11937 7030
rect 11883 6984 11893 7018
rect 11927 6984 11937 7018
rect 11883 6950 11937 6984
rect 11883 6916 11893 6950
rect 11927 6916 11937 6950
rect 11883 6830 11937 6916
rect 11967 6996 12021 7030
rect 11967 6962 11977 6996
rect 12011 6962 12021 6996
rect 11967 6901 12021 6962
rect 11967 6867 11977 6901
rect 12011 6867 12021 6901
rect 11967 6830 12021 6867
rect 12051 7018 12105 7030
rect 12051 6984 12061 7018
rect 12095 6984 12105 7018
rect 12051 6950 12105 6984
rect 12051 6916 12061 6950
rect 12095 6916 12105 6950
rect 12051 6830 12105 6916
rect 12135 6996 12189 7030
rect 12135 6962 12145 6996
rect 12179 6962 12189 6996
rect 12135 6901 12189 6962
rect 12135 6867 12145 6901
rect 12179 6867 12189 6901
rect 12135 6830 12189 6867
rect 12219 7018 12271 7030
rect 12219 6984 12229 7018
rect 12263 6984 12271 7018
rect 12219 6950 12271 6984
rect 12219 6916 12229 6950
rect 12263 6916 12271 6950
rect 12219 6882 12271 6916
rect 12219 6848 12229 6882
rect 12263 6848 12271 6882
rect 12219 6830 12271 6848
rect 12785 7018 12852 7030
rect 12785 6984 12793 7018
rect 12827 6984 12852 7018
rect 12785 6950 12852 6984
rect 12785 6916 12793 6950
rect 12827 6916 12852 6950
rect 12785 6882 12852 6916
rect 12785 6848 12793 6882
rect 12827 6848 12852 6882
rect 12785 6830 12852 6848
rect 12882 7008 12936 7030
rect 12882 6974 12892 7008
rect 12926 6974 12936 7008
rect 12882 6882 12936 6974
rect 12882 6848 12892 6882
rect 12926 6848 12936 6882
rect 12882 6830 12936 6848
rect 12966 7018 13036 7030
rect 12966 6984 12976 7018
rect 13010 6984 13036 7018
rect 12966 6950 13036 6984
rect 12966 6916 12976 6950
rect 13010 6916 13036 6950
rect 12966 6882 13036 6916
rect 12966 6848 12976 6882
rect 13010 6848 13036 6882
rect 12966 6830 13036 6848
rect 13066 7008 13120 7030
rect 13066 6974 13076 7008
rect 13110 6974 13120 7008
rect 13066 6934 13120 6974
rect 13066 6900 13076 6934
rect 13110 6900 13120 6934
rect 13066 6830 13120 6900
rect 13150 7018 13217 7030
rect 13150 6984 13160 7018
rect 13194 6984 13217 7018
rect 13150 6950 13217 6984
rect 13150 6916 13160 6950
rect 13194 6916 13217 6950
rect 13150 6902 13217 6916
rect 13247 6946 13318 7030
rect 13348 6998 13402 7030
rect 13348 6964 13358 6998
rect 13392 6964 13402 6998
rect 13348 6946 13402 6964
rect 13432 6946 13537 7030
rect 13247 6902 13303 6946
rect 13150 6830 13202 6902
rect 13487 6902 13537 6946
rect 13567 6984 13619 7030
rect 13567 6950 13577 6984
rect 13611 6950 13619 6984
rect 14126 7006 14225 7030
rect 13567 6902 13619 6950
rect 13673 6896 13725 6957
rect 13673 6862 13681 6896
rect 13715 6862 13725 6896
rect 13673 6849 13725 6862
rect 13755 6895 13809 6957
rect 13755 6861 13765 6895
rect 13799 6861 13809 6895
rect 13755 6849 13809 6861
rect 13839 6945 13891 6957
rect 13839 6911 13849 6945
rect 13883 6911 13891 6945
rect 13839 6849 13891 6911
rect 13945 6924 13997 7006
rect 13945 6890 13953 6924
rect 13987 6890 13997 6924
rect 13945 6878 13997 6890
rect 14027 6994 14081 7006
rect 14027 6960 14037 6994
rect 14071 6960 14081 6994
rect 14027 6878 14081 6960
rect 14111 6946 14225 7006
rect 14255 6992 14309 7030
rect 14255 6958 14265 6992
rect 14299 6958 14309 6992
rect 14255 6946 14309 6958
rect 14339 6946 14405 7030
rect 14111 6878 14169 6946
rect 14354 6902 14405 6946
rect 14435 7018 14489 7030
rect 14435 6984 14445 7018
rect 14479 6984 14489 7018
rect 14435 6902 14489 6984
rect 14519 6992 14571 7030
rect 14519 6958 14529 6992
rect 14563 6958 14571 6992
rect 14519 6902 14571 6958
rect 24529 7008 24587 7020
rect 24529 6948 24541 7008
rect 24575 6948 24587 7008
rect 24529 6936 24587 6948
rect 24617 7008 24675 7020
rect 24617 6948 24629 7008
rect 24663 6948 24675 7008
rect 24617 6936 24675 6948
rect 24529 6870 24587 6882
rect 24529 6810 24541 6870
rect 24575 6810 24587 6870
rect 24529 6798 24587 6810
rect 24617 6870 24675 6882
rect 24617 6810 24629 6870
rect 24663 6810 24675 6870
rect 24617 6798 24675 6810
rect 24529 6732 24587 6744
rect 24529 6672 24541 6732
rect 24575 6672 24587 6732
rect 24529 6660 24587 6672
rect 24617 6732 24675 6744
rect 24617 6672 24629 6732
rect 24663 6672 24675 6732
rect 24617 6660 24675 6672
rect 24067 6637 24119 6649
rect 24067 6603 24075 6637
rect 24109 6603 24119 6637
rect 24067 6569 24119 6603
rect 24067 6535 24075 6569
rect 24109 6535 24119 6569
rect 24067 6501 24119 6535
rect 24067 6467 24075 6501
rect 24109 6467 24119 6501
rect 24067 6449 24119 6467
rect 24149 6637 24201 6649
rect 24149 6603 24159 6637
rect 24193 6603 24201 6637
rect 24149 6569 24201 6603
rect 24149 6535 24159 6569
rect 24193 6535 24201 6569
rect 24149 6501 24201 6535
rect 24149 6467 24159 6501
rect 24193 6467 24201 6501
rect 24149 6449 24201 6467
rect 24257 6637 24309 6649
rect 24257 6603 24265 6637
rect 24299 6603 24309 6637
rect 24257 6569 24309 6603
rect 24257 6535 24265 6569
rect 24299 6535 24309 6569
rect 24257 6501 24309 6535
rect 24257 6467 24265 6501
rect 24299 6467 24309 6501
rect 24257 6449 24309 6467
rect 24339 6637 24391 6649
rect 24339 6603 24349 6637
rect 24383 6603 24391 6637
rect 24339 6569 24391 6603
rect 24339 6535 24349 6569
rect 24383 6535 24391 6569
rect 24339 6501 24391 6535
rect 24529 6594 24587 6606
rect 24529 6534 24541 6594
rect 24575 6534 24587 6594
rect 24529 6522 24587 6534
rect 24617 6594 24675 6606
rect 24617 6534 24629 6594
rect 24663 6534 24675 6594
rect 24617 6522 24675 6534
rect 24339 6467 24349 6501
rect 24383 6467 24391 6501
rect 24339 6449 24391 6467
rect 30314 6283 30372 6295
rect 11524 6137 11576 6151
rect 11524 6103 11532 6137
rect 11566 6103 11576 6137
rect 11524 6069 11576 6103
rect 11524 6035 11532 6069
rect 11566 6035 11576 6069
rect 11524 6023 11576 6035
rect 11606 6121 11660 6151
rect 11606 6087 11616 6121
rect 11650 6087 11660 6121
rect 11606 6023 11660 6087
rect 11690 6137 11742 6151
rect 11690 6103 11700 6137
rect 11734 6103 11742 6137
rect 11690 6069 11742 6103
rect 11796 6121 11848 6157
rect 11796 6087 11804 6121
rect 11838 6087 11848 6121
rect 11796 6073 11848 6087
rect 11878 6137 11941 6157
rect 11878 6103 11888 6137
rect 11922 6103 11941 6137
rect 11878 6073 11941 6103
rect 11971 6144 12025 6157
rect 11971 6110 11981 6144
rect 12015 6110 12025 6144
rect 11971 6073 12025 6110
rect 12055 6073 12145 6157
rect 12175 6135 12251 6157
rect 12175 6101 12195 6135
rect 12229 6101 12251 6135
rect 12175 6073 12251 6101
rect 12281 6119 12359 6157
rect 12281 6085 12315 6119
rect 12349 6085 12359 6119
rect 12281 6073 12359 6085
rect 11690 6035 11700 6069
rect 11734 6035 11742 6069
rect 11690 6023 11742 6035
rect 12297 6051 12359 6073
rect 12297 6017 12315 6051
rect 12349 6017 12359 6051
rect 12297 5989 12359 6017
rect 12389 5989 12443 6157
rect 12473 6145 12580 6157
rect 12473 6111 12489 6145
rect 12523 6111 12580 6145
rect 12473 6077 12580 6111
rect 12473 6043 12489 6077
rect 12523 6043 12580 6077
rect 12473 5989 12580 6043
rect 12610 6073 12724 6157
rect 12754 6144 12808 6157
rect 12754 6110 12764 6144
rect 12798 6110 12808 6144
rect 12754 6073 12808 6110
rect 12838 6073 12926 6157
rect 12956 6145 13034 6157
rect 12956 6111 12978 6145
rect 13012 6111 13034 6145
rect 12956 6073 13034 6111
rect 13064 6119 13130 6157
rect 13064 6085 13086 6119
rect 13120 6085 13130 6119
rect 13064 6073 13130 6085
rect 12610 5989 12662 6073
rect 13079 5989 13130 6073
rect 13160 5989 13202 6157
rect 13232 6145 13284 6157
rect 13232 6111 13242 6145
rect 13276 6111 13284 6145
rect 13232 5989 13284 6111
rect 13445 6145 13497 6157
rect 13445 6111 13453 6145
rect 13487 6111 13497 6145
rect 13445 6089 13497 6111
rect 13348 6009 13400 6089
rect 13348 5975 13356 6009
rect 13390 5975 13400 6009
rect 13348 5961 13400 5975
rect 13430 5961 13497 6089
rect 13447 5957 13497 5961
rect 13527 6108 13579 6157
rect 13730 6141 13780 6157
rect 13527 6074 13537 6108
rect 13571 6074 13579 6108
rect 13527 6040 13579 6074
rect 13527 6006 13537 6040
rect 13571 6006 13579 6040
rect 13633 6127 13685 6141
rect 13633 6093 13641 6127
rect 13675 6093 13685 6127
rect 13633 6059 13685 6093
rect 13633 6025 13641 6059
rect 13675 6025 13685 6059
rect 13633 6013 13685 6025
rect 13715 6133 13780 6141
rect 13715 6099 13736 6133
rect 13770 6099 13780 6133
rect 13715 6065 13780 6099
rect 13715 6031 13736 6065
rect 13770 6031 13780 6065
rect 13715 6013 13780 6031
rect 13527 5957 13579 6006
rect 13730 5957 13780 6013
rect 13810 6109 13862 6157
rect 13810 6075 13820 6109
rect 13854 6075 13862 6109
rect 13810 6041 13862 6075
rect 13810 6007 13820 6041
rect 13854 6007 13862 6041
rect 13916 6137 13968 6151
rect 13916 6103 13924 6137
rect 13958 6103 13968 6137
rect 13916 6069 13968 6103
rect 13916 6035 13924 6069
rect 13958 6035 13968 6069
rect 13916 6023 13968 6035
rect 13998 6121 14052 6151
rect 13998 6087 14008 6121
rect 14042 6087 14052 6121
rect 13998 6023 14052 6087
rect 14082 6137 14134 6151
rect 14082 6103 14092 6137
rect 14126 6103 14134 6137
rect 14082 6069 14134 6103
rect 14188 6121 14240 6157
rect 14188 6087 14196 6121
rect 14230 6087 14240 6121
rect 14188 6073 14240 6087
rect 14270 6137 14333 6157
rect 14270 6103 14280 6137
rect 14314 6103 14333 6137
rect 14270 6073 14333 6103
rect 14363 6144 14417 6157
rect 14363 6110 14373 6144
rect 14407 6110 14417 6144
rect 14363 6073 14417 6110
rect 14447 6073 14537 6157
rect 14567 6135 14643 6157
rect 14567 6101 14587 6135
rect 14621 6101 14643 6135
rect 14567 6073 14643 6101
rect 14673 6119 14751 6157
rect 14673 6085 14707 6119
rect 14741 6085 14751 6119
rect 14673 6073 14751 6085
rect 14082 6035 14092 6069
rect 14126 6035 14134 6069
rect 14082 6023 14134 6035
rect 13810 5957 13862 6007
rect 14689 6051 14751 6073
rect 14689 6017 14707 6051
rect 14741 6017 14751 6051
rect 14689 5989 14751 6017
rect 14781 5989 14835 6157
rect 14865 6145 14972 6157
rect 14865 6111 14881 6145
rect 14915 6111 14972 6145
rect 14865 6077 14972 6111
rect 14865 6043 14881 6077
rect 14915 6043 14972 6077
rect 14865 5989 14972 6043
rect 15002 6073 15116 6157
rect 15146 6144 15200 6157
rect 15146 6110 15156 6144
rect 15190 6110 15200 6144
rect 15146 6073 15200 6110
rect 15230 6073 15318 6157
rect 15348 6145 15426 6157
rect 15348 6111 15370 6145
rect 15404 6111 15426 6145
rect 15348 6073 15426 6111
rect 15456 6119 15522 6157
rect 15456 6085 15478 6119
rect 15512 6085 15522 6119
rect 15456 6073 15522 6085
rect 15002 5989 15054 6073
rect 15471 5989 15522 6073
rect 15552 5989 15594 6157
rect 15624 6145 15676 6157
rect 15624 6111 15634 6145
rect 15668 6111 15676 6145
rect 15837 6145 15889 6157
rect 15624 5989 15676 6111
rect 15837 6111 15845 6145
rect 15879 6111 15889 6145
rect 15837 6089 15889 6111
rect 15740 6009 15792 6089
rect 15740 5975 15748 6009
rect 15782 5975 15792 6009
rect 15740 5961 15792 5975
rect 15822 5961 15889 6089
rect 15839 5957 15889 5961
rect 15919 6108 15971 6157
rect 16122 6141 16172 6157
rect 15919 6074 15929 6108
rect 15963 6074 15971 6108
rect 15919 6040 15971 6074
rect 15919 6006 15929 6040
rect 15963 6006 15971 6040
rect 16025 6127 16077 6141
rect 16025 6093 16033 6127
rect 16067 6093 16077 6127
rect 16025 6059 16077 6093
rect 16025 6025 16033 6059
rect 16067 6025 16077 6059
rect 16025 6013 16077 6025
rect 16107 6133 16172 6141
rect 16107 6099 16128 6133
rect 16162 6099 16172 6133
rect 16107 6065 16172 6099
rect 16107 6031 16128 6065
rect 16162 6031 16172 6065
rect 16107 6013 16172 6031
rect 15919 5957 15971 6006
rect 16122 5957 16172 6013
rect 16202 6109 16254 6157
rect 16202 6075 16212 6109
rect 16246 6075 16254 6109
rect 16202 6041 16254 6075
rect 16202 6007 16212 6041
rect 16246 6007 16254 6041
rect 16308 6137 16360 6151
rect 16308 6103 16316 6137
rect 16350 6103 16360 6137
rect 16308 6069 16360 6103
rect 16308 6035 16316 6069
rect 16350 6035 16360 6069
rect 16308 6023 16360 6035
rect 16390 6121 16444 6151
rect 16390 6087 16400 6121
rect 16434 6087 16444 6121
rect 16390 6023 16444 6087
rect 16474 6137 16526 6151
rect 16474 6103 16484 6137
rect 16518 6103 16526 6137
rect 16474 6069 16526 6103
rect 16580 6121 16632 6157
rect 16580 6087 16588 6121
rect 16622 6087 16632 6121
rect 16580 6073 16632 6087
rect 16662 6137 16725 6157
rect 16662 6103 16672 6137
rect 16706 6103 16725 6137
rect 16662 6073 16725 6103
rect 16755 6144 16809 6157
rect 16755 6110 16765 6144
rect 16799 6110 16809 6144
rect 16755 6073 16809 6110
rect 16839 6073 16929 6157
rect 16959 6135 17035 6157
rect 16959 6101 16979 6135
rect 17013 6101 17035 6135
rect 16959 6073 17035 6101
rect 17065 6119 17143 6157
rect 17065 6085 17099 6119
rect 17133 6085 17143 6119
rect 17065 6073 17143 6085
rect 16474 6035 16484 6069
rect 16518 6035 16526 6069
rect 16474 6023 16526 6035
rect 16202 5957 16254 6007
rect 17081 6051 17143 6073
rect 17081 6017 17099 6051
rect 17133 6017 17143 6051
rect 17081 5989 17143 6017
rect 17173 5989 17227 6157
rect 17257 6145 17364 6157
rect 17257 6111 17273 6145
rect 17307 6111 17364 6145
rect 17257 6077 17364 6111
rect 17257 6043 17273 6077
rect 17307 6043 17364 6077
rect 17257 5989 17364 6043
rect 17394 6073 17508 6157
rect 17538 6144 17592 6157
rect 17538 6110 17548 6144
rect 17582 6110 17592 6144
rect 17538 6073 17592 6110
rect 17622 6073 17710 6157
rect 17740 6145 17818 6157
rect 17740 6111 17762 6145
rect 17796 6111 17818 6145
rect 17740 6073 17818 6111
rect 17848 6119 17914 6157
rect 17848 6085 17870 6119
rect 17904 6085 17914 6119
rect 17848 6073 17914 6085
rect 17394 5989 17446 6073
rect 17863 5989 17914 6073
rect 17944 5989 17986 6157
rect 18016 6145 18068 6157
rect 18016 6111 18026 6145
rect 18060 6111 18068 6145
rect 18229 6145 18281 6157
rect 18016 5989 18068 6111
rect 18229 6111 18237 6145
rect 18271 6111 18281 6145
rect 18229 6089 18281 6111
rect 18132 6009 18184 6089
rect 18132 5975 18140 6009
rect 18174 5975 18184 6009
rect 18132 5961 18184 5975
rect 18214 5961 18281 6089
rect 18231 5957 18281 5961
rect 18311 6108 18363 6157
rect 18514 6141 18564 6157
rect 18311 6074 18321 6108
rect 18355 6074 18363 6108
rect 18311 6040 18363 6074
rect 18311 6006 18321 6040
rect 18355 6006 18363 6040
rect 18417 6127 18469 6141
rect 18417 6093 18425 6127
rect 18459 6093 18469 6127
rect 18417 6059 18469 6093
rect 18417 6025 18425 6059
rect 18459 6025 18469 6059
rect 18417 6013 18469 6025
rect 18499 6133 18564 6141
rect 18499 6099 18520 6133
rect 18554 6099 18564 6133
rect 18499 6065 18564 6099
rect 18499 6031 18520 6065
rect 18554 6031 18564 6065
rect 18499 6013 18564 6031
rect 18311 5957 18363 6006
rect 18514 5957 18564 6013
rect 18594 6109 18646 6157
rect 18594 6075 18604 6109
rect 18638 6075 18646 6109
rect 18594 6041 18646 6075
rect 18594 6007 18604 6041
rect 18638 6007 18646 6041
rect 18700 6137 18752 6151
rect 18700 6103 18708 6137
rect 18742 6103 18752 6137
rect 18700 6069 18752 6103
rect 18700 6035 18708 6069
rect 18742 6035 18752 6069
rect 18700 6023 18752 6035
rect 18782 6121 18836 6151
rect 18782 6087 18792 6121
rect 18826 6087 18836 6121
rect 18782 6023 18836 6087
rect 18866 6137 18918 6151
rect 18866 6103 18876 6137
rect 18910 6103 18918 6137
rect 18866 6069 18918 6103
rect 18972 6121 19024 6157
rect 18972 6087 18980 6121
rect 19014 6087 19024 6121
rect 18972 6073 19024 6087
rect 19054 6137 19117 6157
rect 19054 6103 19064 6137
rect 19098 6103 19117 6137
rect 19054 6073 19117 6103
rect 19147 6144 19201 6157
rect 19147 6110 19157 6144
rect 19191 6110 19201 6144
rect 19147 6073 19201 6110
rect 19231 6073 19321 6157
rect 19351 6135 19427 6157
rect 19351 6101 19371 6135
rect 19405 6101 19427 6135
rect 19351 6073 19427 6101
rect 19457 6119 19535 6157
rect 19457 6085 19491 6119
rect 19525 6085 19535 6119
rect 19457 6073 19535 6085
rect 18866 6035 18876 6069
rect 18910 6035 18918 6069
rect 18866 6023 18918 6035
rect 18594 5957 18646 6007
rect 19473 6051 19535 6073
rect 19473 6017 19491 6051
rect 19525 6017 19535 6051
rect 19473 5989 19535 6017
rect 19565 5989 19619 6157
rect 19649 6145 19756 6157
rect 19649 6111 19665 6145
rect 19699 6111 19756 6145
rect 19649 6077 19756 6111
rect 19649 6043 19665 6077
rect 19699 6043 19756 6077
rect 19649 5989 19756 6043
rect 19786 6073 19900 6157
rect 19930 6144 19984 6157
rect 19930 6110 19940 6144
rect 19974 6110 19984 6144
rect 19930 6073 19984 6110
rect 20014 6073 20102 6157
rect 20132 6145 20210 6157
rect 20132 6111 20154 6145
rect 20188 6111 20210 6145
rect 20132 6073 20210 6111
rect 20240 6119 20306 6157
rect 20240 6085 20262 6119
rect 20296 6085 20306 6119
rect 20240 6073 20306 6085
rect 19786 5989 19838 6073
rect 20255 5989 20306 6073
rect 20336 5989 20378 6157
rect 20408 6145 20460 6157
rect 20408 6111 20418 6145
rect 20452 6111 20460 6145
rect 20621 6145 20673 6157
rect 20408 5989 20460 6111
rect 20621 6111 20629 6145
rect 20663 6111 20673 6145
rect 20621 6089 20673 6111
rect 20524 6009 20576 6089
rect 20524 5975 20532 6009
rect 20566 5975 20576 6009
rect 20524 5961 20576 5975
rect 20606 5961 20673 6089
rect 20623 5957 20673 5961
rect 20703 6108 20755 6157
rect 20906 6141 20956 6157
rect 20703 6074 20713 6108
rect 20747 6074 20755 6108
rect 20703 6040 20755 6074
rect 20703 6006 20713 6040
rect 20747 6006 20755 6040
rect 20809 6127 20861 6141
rect 20809 6093 20817 6127
rect 20851 6093 20861 6127
rect 20809 6059 20861 6093
rect 20809 6025 20817 6059
rect 20851 6025 20861 6059
rect 20809 6013 20861 6025
rect 20891 6133 20956 6141
rect 20891 6099 20912 6133
rect 20946 6099 20956 6133
rect 20891 6065 20956 6099
rect 20891 6031 20912 6065
rect 20946 6031 20956 6065
rect 20891 6013 20956 6031
rect 20703 5957 20755 6006
rect 20906 5957 20956 6013
rect 20986 6109 21038 6157
rect 20986 6075 20996 6109
rect 21030 6075 21038 6109
rect 20986 6041 21038 6075
rect 20986 6007 20996 6041
rect 21030 6007 21038 6041
rect 21092 6137 21144 6151
rect 21092 6103 21100 6137
rect 21134 6103 21144 6137
rect 21092 6069 21144 6103
rect 21092 6035 21100 6069
rect 21134 6035 21144 6069
rect 21092 6023 21144 6035
rect 21174 6121 21228 6151
rect 21174 6087 21184 6121
rect 21218 6087 21228 6121
rect 21174 6023 21228 6087
rect 21258 6137 21310 6151
rect 21258 6103 21268 6137
rect 21302 6103 21310 6137
rect 21258 6069 21310 6103
rect 21364 6121 21416 6157
rect 21364 6087 21372 6121
rect 21406 6087 21416 6121
rect 21364 6073 21416 6087
rect 21446 6137 21509 6157
rect 21446 6103 21456 6137
rect 21490 6103 21509 6137
rect 21446 6073 21509 6103
rect 21539 6144 21593 6157
rect 21539 6110 21549 6144
rect 21583 6110 21593 6144
rect 21539 6073 21593 6110
rect 21623 6073 21713 6157
rect 21743 6135 21819 6157
rect 21743 6101 21763 6135
rect 21797 6101 21819 6135
rect 21743 6073 21819 6101
rect 21849 6119 21927 6157
rect 21849 6085 21883 6119
rect 21917 6085 21927 6119
rect 21849 6073 21927 6085
rect 21258 6035 21268 6069
rect 21302 6035 21310 6069
rect 21258 6023 21310 6035
rect 20986 5957 21038 6007
rect 21865 6051 21927 6073
rect 21865 6017 21883 6051
rect 21917 6017 21927 6051
rect 21865 5989 21927 6017
rect 21957 5989 22011 6157
rect 22041 6145 22148 6157
rect 22041 6111 22057 6145
rect 22091 6111 22148 6145
rect 22041 6077 22148 6111
rect 22041 6043 22057 6077
rect 22091 6043 22148 6077
rect 22041 5989 22148 6043
rect 22178 6073 22292 6157
rect 22322 6144 22376 6157
rect 22322 6110 22332 6144
rect 22366 6110 22376 6144
rect 22322 6073 22376 6110
rect 22406 6073 22494 6157
rect 22524 6145 22602 6157
rect 22524 6111 22546 6145
rect 22580 6111 22602 6145
rect 22524 6073 22602 6111
rect 22632 6119 22698 6157
rect 22632 6085 22654 6119
rect 22688 6085 22698 6119
rect 22632 6073 22698 6085
rect 22178 5989 22230 6073
rect 22647 5989 22698 6073
rect 22728 5989 22770 6157
rect 22800 6145 22852 6157
rect 22800 6111 22810 6145
rect 22844 6111 22852 6145
rect 23013 6145 23065 6157
rect 22800 5989 22852 6111
rect 23013 6111 23021 6145
rect 23055 6111 23065 6145
rect 23013 6089 23065 6111
rect 22916 6009 22968 6089
rect 22916 5975 22924 6009
rect 22958 5975 22968 6009
rect 22916 5961 22968 5975
rect 22998 5961 23065 6089
rect 23015 5957 23065 5961
rect 23095 6108 23147 6157
rect 30314 6223 30326 6283
rect 30360 6223 30372 6283
rect 30314 6211 30372 6223
rect 30402 6283 30460 6295
rect 30402 6223 30414 6283
rect 30448 6223 30460 6283
rect 30803 6264 30853 6272
rect 30402 6211 30460 6223
rect 30706 6252 30758 6264
rect 30706 6218 30714 6252
rect 30748 6218 30758 6252
rect 23298 6141 23348 6157
rect 23095 6074 23105 6108
rect 23139 6074 23147 6108
rect 23095 6040 23147 6074
rect 23095 6006 23105 6040
rect 23139 6006 23147 6040
rect 23201 6127 23253 6141
rect 23201 6093 23209 6127
rect 23243 6093 23253 6127
rect 23201 6059 23253 6093
rect 23201 6025 23209 6059
rect 23243 6025 23253 6059
rect 23201 6013 23253 6025
rect 23283 6133 23348 6141
rect 23283 6099 23304 6133
rect 23338 6099 23348 6133
rect 23283 6065 23348 6099
rect 23283 6031 23304 6065
rect 23338 6031 23348 6065
rect 23283 6013 23348 6031
rect 23095 5957 23147 6006
rect 23298 5957 23348 6013
rect 23378 6109 23430 6157
rect 30706 6184 30758 6218
rect 23378 6075 23388 6109
rect 23422 6075 23430 6109
rect 25171 6139 25229 6151
rect 23378 6041 23430 6075
rect 25171 6079 25183 6139
rect 25217 6079 25229 6139
rect 25171 6067 25229 6079
rect 25259 6142 25317 6151
rect 25259 6082 25271 6142
rect 25305 6082 25317 6142
rect 25259 6067 25317 6082
rect 25903 6142 25961 6154
rect 25903 6082 25915 6142
rect 25949 6082 25961 6142
rect 25903 6070 25961 6082
rect 25991 6142 26087 6154
rect 25991 6082 26020 6142
rect 26054 6082 26087 6142
rect 25991 6070 26087 6082
rect 26117 6142 26175 6154
rect 26117 6082 26129 6142
rect 26163 6082 26175 6142
rect 26117 6070 26175 6082
rect 27115 6142 27173 6154
rect 27115 6082 27127 6142
rect 27161 6082 27173 6142
rect 27115 6070 27173 6082
rect 27203 6142 27299 6154
rect 27203 6082 27231 6142
rect 27265 6082 27299 6142
rect 27203 6070 27299 6082
rect 27329 6142 27387 6154
rect 27329 6082 27341 6142
rect 27375 6082 27387 6142
rect 27329 6070 27387 6082
rect 28327 6142 28385 6154
rect 28327 6082 28339 6142
rect 28373 6082 28385 6142
rect 28327 6070 28385 6082
rect 28415 6142 28511 6154
rect 28415 6082 28444 6142
rect 28478 6082 28511 6142
rect 28415 6070 28511 6082
rect 28541 6142 28599 6154
rect 28541 6082 28553 6142
rect 28587 6082 28599 6142
rect 28541 6070 28599 6082
rect 29539 6142 29597 6154
rect 29539 6082 29551 6142
rect 29585 6082 29597 6142
rect 29539 6070 29597 6082
rect 29627 6142 29723 6154
rect 29627 6082 29658 6142
rect 29692 6082 29723 6142
rect 29627 6070 29723 6082
rect 29753 6142 29811 6154
rect 29753 6082 29765 6142
rect 29799 6082 29811 6142
rect 29753 6070 29811 6082
rect 30314 6145 30372 6157
rect 30314 6085 30326 6145
rect 30360 6085 30372 6145
rect 30314 6073 30372 6085
rect 30402 6145 30464 6157
rect 30402 6085 30414 6145
rect 30448 6085 30464 6145
rect 30402 6073 30464 6085
rect 30494 6145 30560 6157
rect 30494 6085 30510 6145
rect 30544 6085 30560 6145
rect 30494 6073 30560 6085
rect 30590 6145 30652 6157
rect 30590 6085 30606 6145
rect 30640 6085 30652 6145
rect 30706 6150 30714 6184
rect 30748 6150 30758 6184
rect 30706 6136 30758 6150
rect 30788 6252 30853 6264
rect 30788 6218 30807 6252
rect 30841 6218 30853 6252
rect 30788 6184 30853 6218
rect 30788 6150 30807 6184
rect 30841 6150 30853 6184
rect 30788 6136 30853 6150
rect 30590 6073 30652 6085
rect 23378 6007 23388 6041
rect 23422 6007 23430 6041
rect 23378 5957 23430 6007
rect 30803 6072 30853 6136
rect 30883 6236 30937 6272
rect 30883 6202 30893 6236
rect 30927 6202 30937 6236
rect 30883 6155 30937 6202
rect 30883 6121 30893 6155
rect 30927 6121 30937 6155
rect 30883 6072 30937 6121
rect 30967 6260 31020 6272
rect 30967 6226 30977 6260
rect 31011 6226 31020 6260
rect 30967 6192 31020 6226
rect 30967 6158 30977 6192
rect 31011 6158 31020 6192
rect 30967 6124 31020 6158
rect 30967 6090 30977 6124
rect 31011 6090 31020 6124
rect 30967 6072 31020 6090
rect 11084 5448 11136 5468
rect 11084 5414 11092 5448
rect 11126 5414 11136 5448
rect 11084 5380 11136 5414
rect 11084 5346 11092 5380
rect 11126 5346 11136 5380
rect 11084 5310 11136 5346
rect 11166 5448 11224 5468
rect 11166 5414 11178 5448
rect 11212 5414 11224 5448
rect 11166 5380 11224 5414
rect 11166 5346 11178 5380
rect 11212 5346 11224 5380
rect 11166 5310 11224 5346
rect 11254 5448 11306 5468
rect 11254 5414 11264 5448
rect 11298 5414 11306 5448
rect 11254 5367 11306 5414
rect 11254 5333 11264 5367
rect 11298 5333 11306 5367
rect 11254 5310 11306 5333
rect 11360 5450 11412 5468
rect 11360 5416 11368 5450
rect 11402 5416 11412 5450
rect 11360 5382 11412 5416
rect 11360 5348 11368 5382
rect 11402 5348 11412 5382
rect 11360 5314 11412 5348
rect 11360 5280 11368 5314
rect 11402 5280 11412 5314
rect 11360 5268 11412 5280
rect 11442 5456 11496 5468
rect 11442 5422 11452 5456
rect 11486 5422 11496 5456
rect 11442 5388 11496 5422
rect 11442 5354 11452 5388
rect 11486 5354 11496 5388
rect 11442 5268 11496 5354
rect 11526 5434 11580 5468
rect 11526 5400 11536 5434
rect 11570 5400 11580 5434
rect 11526 5339 11580 5400
rect 11526 5305 11536 5339
rect 11570 5305 11580 5339
rect 11526 5268 11580 5305
rect 11610 5456 11664 5468
rect 11610 5422 11620 5456
rect 11654 5422 11664 5456
rect 11610 5388 11664 5422
rect 11610 5354 11620 5388
rect 11654 5354 11664 5388
rect 11610 5268 11664 5354
rect 11694 5434 11748 5468
rect 11694 5400 11704 5434
rect 11738 5400 11748 5434
rect 11694 5339 11748 5400
rect 11694 5305 11704 5339
rect 11738 5305 11748 5339
rect 11694 5268 11748 5305
rect 11778 5456 11830 5468
rect 11778 5422 11788 5456
rect 11822 5422 11830 5456
rect 11778 5388 11830 5422
rect 11778 5354 11788 5388
rect 11822 5354 11830 5388
rect 11778 5320 11830 5354
rect 11778 5286 11788 5320
rect 11822 5286 11830 5320
rect 11778 5268 11830 5286
rect 11892 5456 11944 5468
rect 11892 5422 11900 5456
rect 11934 5422 11944 5456
rect 11892 5388 11944 5422
rect 11892 5354 11900 5388
rect 11934 5354 11944 5388
rect 11892 5320 11944 5354
rect 11892 5286 11900 5320
rect 11934 5286 11944 5320
rect 11892 5268 11944 5286
rect 11974 5450 12028 5468
rect 11974 5416 11984 5450
rect 12018 5416 12028 5450
rect 11974 5382 12028 5416
rect 11974 5348 11984 5382
rect 12018 5348 12028 5382
rect 11974 5314 12028 5348
rect 11974 5280 11984 5314
rect 12018 5280 12028 5314
rect 11974 5268 12028 5280
rect 12058 5456 12112 5468
rect 12058 5422 12068 5456
rect 12102 5422 12112 5456
rect 12058 5388 12112 5422
rect 12058 5354 12068 5388
rect 12102 5354 12112 5388
rect 12058 5268 12112 5354
rect 12142 5450 12196 5468
rect 12142 5416 12152 5450
rect 12186 5416 12196 5450
rect 12142 5382 12196 5416
rect 12142 5348 12152 5382
rect 12186 5348 12196 5382
rect 12142 5314 12196 5348
rect 12142 5280 12152 5314
rect 12186 5280 12196 5314
rect 12142 5268 12196 5280
rect 12226 5456 12280 5468
rect 12226 5422 12236 5456
rect 12270 5422 12280 5456
rect 12226 5388 12280 5422
rect 12226 5354 12236 5388
rect 12270 5354 12280 5388
rect 12226 5268 12280 5354
rect 12310 5450 12364 5468
rect 12310 5416 12320 5450
rect 12354 5416 12364 5450
rect 12310 5382 12364 5416
rect 12310 5348 12320 5382
rect 12354 5348 12364 5382
rect 12310 5314 12364 5348
rect 12310 5280 12320 5314
rect 12354 5280 12364 5314
rect 12310 5268 12364 5280
rect 12394 5456 12448 5468
rect 12394 5422 12404 5456
rect 12438 5422 12448 5456
rect 12394 5388 12448 5422
rect 12394 5354 12404 5388
rect 12438 5354 12448 5388
rect 12394 5268 12448 5354
rect 12478 5450 12532 5468
rect 12478 5416 12488 5450
rect 12522 5416 12532 5450
rect 12478 5382 12532 5416
rect 12478 5348 12488 5382
rect 12522 5348 12532 5382
rect 12478 5314 12532 5348
rect 12478 5280 12488 5314
rect 12522 5280 12532 5314
rect 12478 5268 12532 5280
rect 12562 5456 12616 5468
rect 12562 5422 12572 5456
rect 12606 5422 12616 5456
rect 12562 5388 12616 5422
rect 12562 5354 12572 5388
rect 12606 5354 12616 5388
rect 12562 5268 12616 5354
rect 12646 5450 12700 5468
rect 12646 5416 12656 5450
rect 12690 5416 12700 5450
rect 12646 5382 12700 5416
rect 12646 5348 12656 5382
rect 12690 5348 12700 5382
rect 12646 5314 12700 5348
rect 12646 5280 12656 5314
rect 12690 5280 12700 5314
rect 12646 5268 12700 5280
rect 12730 5456 12784 5468
rect 12730 5422 12740 5456
rect 12774 5422 12784 5456
rect 12730 5388 12784 5422
rect 12730 5354 12740 5388
rect 12774 5354 12784 5388
rect 12730 5268 12784 5354
rect 12814 5450 12868 5468
rect 12814 5416 12824 5450
rect 12858 5416 12868 5450
rect 12814 5382 12868 5416
rect 12814 5348 12824 5382
rect 12858 5348 12868 5382
rect 12814 5314 12868 5348
rect 12814 5280 12824 5314
rect 12858 5280 12868 5314
rect 12814 5268 12868 5280
rect 12898 5456 12952 5468
rect 12898 5422 12908 5456
rect 12942 5422 12952 5456
rect 12898 5388 12952 5422
rect 12898 5354 12908 5388
rect 12942 5354 12952 5388
rect 12898 5268 12952 5354
rect 12982 5450 13036 5468
rect 12982 5416 12992 5450
rect 13026 5416 13036 5450
rect 12982 5382 13036 5416
rect 12982 5348 12992 5382
rect 13026 5348 13036 5382
rect 12982 5314 13036 5348
rect 12982 5280 12992 5314
rect 13026 5280 13036 5314
rect 12982 5268 13036 5280
rect 13066 5456 13120 5468
rect 13066 5422 13076 5456
rect 13110 5422 13120 5456
rect 13066 5388 13120 5422
rect 13066 5354 13076 5388
rect 13110 5354 13120 5388
rect 13066 5268 13120 5354
rect 13150 5450 13204 5468
rect 13150 5416 13160 5450
rect 13194 5416 13204 5450
rect 13150 5382 13204 5416
rect 13150 5348 13160 5382
rect 13194 5348 13204 5382
rect 13150 5314 13204 5348
rect 13150 5280 13160 5314
rect 13194 5280 13204 5314
rect 13150 5268 13204 5280
rect 13234 5456 13288 5468
rect 13234 5422 13244 5456
rect 13278 5422 13288 5456
rect 13234 5388 13288 5422
rect 13234 5354 13244 5388
rect 13278 5354 13288 5388
rect 13234 5268 13288 5354
rect 13318 5450 13372 5468
rect 13318 5416 13328 5450
rect 13362 5416 13372 5450
rect 13318 5382 13372 5416
rect 13318 5348 13328 5382
rect 13362 5348 13372 5382
rect 13318 5314 13372 5348
rect 13318 5280 13328 5314
rect 13362 5280 13372 5314
rect 13318 5268 13372 5280
rect 13402 5456 13456 5468
rect 13402 5422 13412 5456
rect 13446 5422 13456 5456
rect 13402 5388 13456 5422
rect 13402 5354 13412 5388
rect 13446 5354 13456 5388
rect 13402 5268 13456 5354
rect 13486 5450 13540 5468
rect 13486 5416 13496 5450
rect 13530 5416 13540 5450
rect 13486 5382 13540 5416
rect 13486 5348 13496 5382
rect 13530 5348 13540 5382
rect 13486 5314 13540 5348
rect 13486 5280 13496 5314
rect 13530 5280 13540 5314
rect 13486 5268 13540 5280
rect 13570 5456 13624 5468
rect 13570 5422 13580 5456
rect 13614 5422 13624 5456
rect 13570 5388 13624 5422
rect 13570 5354 13580 5388
rect 13614 5354 13624 5388
rect 13570 5268 13624 5354
rect 13654 5450 13708 5468
rect 13654 5416 13664 5450
rect 13698 5416 13708 5450
rect 13654 5382 13708 5416
rect 13654 5348 13664 5382
rect 13698 5348 13708 5382
rect 13654 5314 13708 5348
rect 13654 5280 13664 5314
rect 13698 5280 13708 5314
rect 13654 5268 13708 5280
rect 13738 5456 13790 5468
rect 13738 5422 13748 5456
rect 13782 5422 13790 5456
rect 13738 5388 13790 5422
rect 13738 5354 13748 5388
rect 13782 5354 13790 5388
rect 13738 5268 13790 5354
rect 13916 5420 13968 5468
rect 13916 5386 13924 5420
rect 13958 5386 13968 5420
rect 13916 5352 13968 5386
rect 13916 5318 13924 5352
rect 13958 5318 13968 5352
rect 13916 5268 13968 5318
rect 13998 5452 14048 5468
rect 13998 5444 14063 5452
rect 13998 5410 14008 5444
rect 14042 5410 14063 5444
rect 13998 5376 14063 5410
rect 13998 5342 14008 5376
rect 14042 5342 14063 5376
rect 13998 5324 14063 5342
rect 14093 5438 14145 5452
rect 14093 5404 14103 5438
rect 14137 5404 14145 5438
rect 14093 5370 14145 5404
rect 14093 5336 14103 5370
rect 14137 5336 14145 5370
rect 14093 5324 14145 5336
rect 14199 5419 14251 5468
rect 14199 5385 14207 5419
rect 14241 5385 14251 5419
rect 14199 5351 14251 5385
rect 13998 5268 14048 5324
rect 14199 5317 14207 5351
rect 14241 5317 14251 5351
rect 14199 5268 14251 5317
rect 14281 5456 14333 5468
rect 14281 5422 14291 5456
rect 14325 5422 14333 5456
rect 14494 5456 14546 5468
rect 14281 5400 14333 5422
rect 14494 5422 14502 5456
rect 14536 5422 14546 5456
rect 14281 5272 14348 5400
rect 14378 5320 14430 5400
rect 14378 5286 14388 5320
rect 14422 5286 14430 5320
rect 14494 5300 14546 5422
rect 14576 5300 14618 5468
rect 14648 5430 14714 5468
rect 14648 5396 14658 5430
rect 14692 5396 14714 5430
rect 14648 5384 14714 5396
rect 14744 5456 14822 5468
rect 14744 5422 14766 5456
rect 14800 5422 14822 5456
rect 14744 5384 14822 5422
rect 14852 5384 14940 5468
rect 14970 5455 15024 5468
rect 14970 5421 14980 5455
rect 15014 5421 15024 5455
rect 14970 5384 15024 5421
rect 15054 5384 15168 5468
rect 14648 5300 14699 5384
rect 14378 5272 14430 5286
rect 14281 5268 14331 5272
rect 15116 5300 15168 5384
rect 15198 5456 15305 5468
rect 15198 5422 15255 5456
rect 15289 5422 15305 5456
rect 15198 5388 15305 5422
rect 15198 5354 15255 5388
rect 15289 5354 15305 5388
rect 15198 5300 15305 5354
rect 15335 5300 15389 5468
rect 15419 5430 15497 5468
rect 15419 5396 15429 5430
rect 15463 5396 15497 5430
rect 15419 5384 15497 5396
rect 15527 5446 15603 5468
rect 15527 5412 15549 5446
rect 15583 5412 15603 5446
rect 15527 5384 15603 5412
rect 15633 5384 15723 5468
rect 15753 5455 15807 5468
rect 15753 5421 15763 5455
rect 15797 5421 15807 5455
rect 15753 5384 15807 5421
rect 15837 5448 15900 5468
rect 15837 5414 15856 5448
rect 15890 5414 15900 5448
rect 15837 5384 15900 5414
rect 15930 5432 15982 5468
rect 15930 5398 15940 5432
rect 15974 5398 15982 5432
rect 15930 5384 15982 5398
rect 16036 5448 16088 5462
rect 16036 5414 16044 5448
rect 16078 5414 16088 5448
rect 15419 5362 15481 5384
rect 15419 5328 15429 5362
rect 15463 5328 15481 5362
rect 15419 5300 15481 5328
rect 16036 5380 16088 5414
rect 16036 5346 16044 5380
rect 16078 5346 16088 5380
rect 16036 5334 16088 5346
rect 16118 5432 16172 5462
rect 16118 5398 16128 5432
rect 16162 5398 16172 5432
rect 16118 5334 16172 5398
rect 16202 5448 16254 5462
rect 16202 5414 16212 5448
rect 16246 5414 16254 5448
rect 16202 5380 16254 5414
rect 16202 5346 16212 5380
rect 16246 5346 16254 5380
rect 16202 5334 16254 5346
rect 16308 5420 16360 5468
rect 16308 5386 16316 5420
rect 16350 5386 16360 5420
rect 16308 5352 16360 5386
rect 16308 5318 16316 5352
rect 16350 5318 16360 5352
rect 16308 5268 16360 5318
rect 16390 5452 16440 5468
rect 16390 5444 16455 5452
rect 16390 5410 16400 5444
rect 16434 5410 16455 5444
rect 16390 5376 16455 5410
rect 16390 5342 16400 5376
rect 16434 5342 16455 5376
rect 16390 5324 16455 5342
rect 16485 5438 16537 5452
rect 16485 5404 16495 5438
rect 16529 5404 16537 5438
rect 16485 5370 16537 5404
rect 16485 5336 16495 5370
rect 16529 5336 16537 5370
rect 16485 5324 16537 5336
rect 16591 5419 16643 5468
rect 16591 5385 16599 5419
rect 16633 5385 16643 5419
rect 16591 5351 16643 5385
rect 16390 5268 16440 5324
rect 16591 5317 16599 5351
rect 16633 5317 16643 5351
rect 16591 5268 16643 5317
rect 16673 5456 16725 5468
rect 16673 5422 16683 5456
rect 16717 5422 16725 5456
rect 16886 5456 16938 5468
rect 16673 5400 16725 5422
rect 16886 5422 16894 5456
rect 16928 5422 16938 5456
rect 16673 5272 16740 5400
rect 16770 5320 16822 5400
rect 16770 5286 16780 5320
rect 16814 5286 16822 5320
rect 16886 5300 16938 5422
rect 16968 5300 17010 5468
rect 17040 5430 17106 5468
rect 17040 5396 17050 5430
rect 17084 5396 17106 5430
rect 17040 5384 17106 5396
rect 17136 5456 17214 5468
rect 17136 5422 17158 5456
rect 17192 5422 17214 5456
rect 17136 5384 17214 5422
rect 17244 5384 17332 5468
rect 17362 5455 17416 5468
rect 17362 5421 17372 5455
rect 17406 5421 17416 5455
rect 17362 5384 17416 5421
rect 17446 5384 17560 5468
rect 17040 5300 17091 5384
rect 16770 5272 16822 5286
rect 16673 5268 16723 5272
rect 17508 5300 17560 5384
rect 17590 5456 17697 5468
rect 17590 5422 17647 5456
rect 17681 5422 17697 5456
rect 17590 5388 17697 5422
rect 17590 5354 17647 5388
rect 17681 5354 17697 5388
rect 17590 5300 17697 5354
rect 17727 5300 17781 5468
rect 17811 5430 17889 5468
rect 17811 5396 17821 5430
rect 17855 5396 17889 5430
rect 17811 5384 17889 5396
rect 17919 5446 17995 5468
rect 17919 5412 17941 5446
rect 17975 5412 17995 5446
rect 17919 5384 17995 5412
rect 18025 5384 18115 5468
rect 18145 5455 18199 5468
rect 18145 5421 18155 5455
rect 18189 5421 18199 5455
rect 18145 5384 18199 5421
rect 18229 5448 18292 5468
rect 18229 5414 18248 5448
rect 18282 5414 18292 5448
rect 18229 5384 18292 5414
rect 18322 5432 18374 5468
rect 18322 5398 18332 5432
rect 18366 5398 18374 5432
rect 18322 5384 18374 5398
rect 18428 5448 18480 5462
rect 18428 5414 18436 5448
rect 18470 5414 18480 5448
rect 17811 5362 17873 5384
rect 17811 5328 17821 5362
rect 17855 5328 17873 5362
rect 17811 5300 17873 5328
rect 18428 5380 18480 5414
rect 18428 5346 18436 5380
rect 18470 5346 18480 5380
rect 18428 5334 18480 5346
rect 18510 5432 18564 5462
rect 18510 5398 18520 5432
rect 18554 5398 18564 5432
rect 18510 5334 18564 5398
rect 18594 5448 18646 5462
rect 18594 5414 18604 5448
rect 18638 5414 18646 5448
rect 18594 5380 18646 5414
rect 18594 5346 18604 5380
rect 18638 5346 18646 5380
rect 18594 5334 18646 5346
rect 18700 5420 18752 5468
rect 18700 5386 18708 5420
rect 18742 5386 18752 5420
rect 18700 5352 18752 5386
rect 18700 5318 18708 5352
rect 18742 5318 18752 5352
rect 18700 5268 18752 5318
rect 18782 5452 18832 5468
rect 18782 5444 18847 5452
rect 18782 5410 18792 5444
rect 18826 5410 18847 5444
rect 18782 5376 18847 5410
rect 18782 5342 18792 5376
rect 18826 5342 18847 5376
rect 18782 5324 18847 5342
rect 18877 5438 18929 5452
rect 18877 5404 18887 5438
rect 18921 5404 18929 5438
rect 18877 5370 18929 5404
rect 18877 5336 18887 5370
rect 18921 5336 18929 5370
rect 18877 5324 18929 5336
rect 18983 5419 19035 5468
rect 18983 5385 18991 5419
rect 19025 5385 19035 5419
rect 18983 5351 19035 5385
rect 18782 5268 18832 5324
rect 18983 5317 18991 5351
rect 19025 5317 19035 5351
rect 18983 5268 19035 5317
rect 19065 5456 19117 5468
rect 19065 5422 19075 5456
rect 19109 5422 19117 5456
rect 19278 5456 19330 5468
rect 19065 5400 19117 5422
rect 19278 5422 19286 5456
rect 19320 5422 19330 5456
rect 19065 5272 19132 5400
rect 19162 5320 19214 5400
rect 19162 5286 19172 5320
rect 19206 5286 19214 5320
rect 19278 5300 19330 5422
rect 19360 5300 19402 5468
rect 19432 5430 19498 5468
rect 19432 5396 19442 5430
rect 19476 5396 19498 5430
rect 19432 5384 19498 5396
rect 19528 5456 19606 5468
rect 19528 5422 19550 5456
rect 19584 5422 19606 5456
rect 19528 5384 19606 5422
rect 19636 5384 19724 5468
rect 19754 5455 19808 5468
rect 19754 5421 19764 5455
rect 19798 5421 19808 5455
rect 19754 5384 19808 5421
rect 19838 5384 19952 5468
rect 19432 5300 19483 5384
rect 19162 5272 19214 5286
rect 19065 5268 19115 5272
rect 19900 5300 19952 5384
rect 19982 5456 20089 5468
rect 19982 5422 20039 5456
rect 20073 5422 20089 5456
rect 19982 5388 20089 5422
rect 19982 5354 20039 5388
rect 20073 5354 20089 5388
rect 19982 5300 20089 5354
rect 20119 5300 20173 5468
rect 20203 5430 20281 5468
rect 20203 5396 20213 5430
rect 20247 5396 20281 5430
rect 20203 5384 20281 5396
rect 20311 5446 20387 5468
rect 20311 5412 20333 5446
rect 20367 5412 20387 5446
rect 20311 5384 20387 5412
rect 20417 5384 20507 5468
rect 20537 5455 20591 5468
rect 20537 5421 20547 5455
rect 20581 5421 20591 5455
rect 20537 5384 20591 5421
rect 20621 5448 20684 5468
rect 20621 5414 20640 5448
rect 20674 5414 20684 5448
rect 20621 5384 20684 5414
rect 20714 5432 20766 5468
rect 20714 5398 20724 5432
rect 20758 5398 20766 5432
rect 20714 5384 20766 5398
rect 20820 5448 20872 5462
rect 20820 5414 20828 5448
rect 20862 5414 20872 5448
rect 20203 5362 20265 5384
rect 20203 5328 20213 5362
rect 20247 5328 20265 5362
rect 20203 5300 20265 5328
rect 20820 5380 20872 5414
rect 20820 5346 20828 5380
rect 20862 5346 20872 5380
rect 20820 5334 20872 5346
rect 20902 5432 20956 5462
rect 20902 5398 20912 5432
rect 20946 5398 20956 5432
rect 20902 5334 20956 5398
rect 20986 5448 21038 5462
rect 20986 5414 20996 5448
rect 21030 5414 21038 5448
rect 20986 5380 21038 5414
rect 20986 5346 20996 5380
rect 21030 5346 21038 5380
rect 20986 5334 21038 5346
rect 21092 5420 21144 5468
rect 21092 5386 21100 5420
rect 21134 5386 21144 5420
rect 21092 5352 21144 5386
rect 21092 5318 21100 5352
rect 21134 5318 21144 5352
rect 21092 5268 21144 5318
rect 21174 5452 21224 5468
rect 21174 5444 21239 5452
rect 21174 5410 21184 5444
rect 21218 5410 21239 5444
rect 21174 5376 21239 5410
rect 21174 5342 21184 5376
rect 21218 5342 21239 5376
rect 21174 5324 21239 5342
rect 21269 5438 21321 5452
rect 21269 5404 21279 5438
rect 21313 5404 21321 5438
rect 21269 5370 21321 5404
rect 21269 5336 21279 5370
rect 21313 5336 21321 5370
rect 21269 5324 21321 5336
rect 21375 5419 21427 5468
rect 21375 5385 21383 5419
rect 21417 5385 21427 5419
rect 21375 5351 21427 5385
rect 21174 5268 21224 5324
rect 21375 5317 21383 5351
rect 21417 5317 21427 5351
rect 21375 5268 21427 5317
rect 21457 5456 21509 5468
rect 21457 5422 21467 5456
rect 21501 5422 21509 5456
rect 21670 5456 21722 5468
rect 21457 5400 21509 5422
rect 21670 5422 21678 5456
rect 21712 5422 21722 5456
rect 21457 5272 21524 5400
rect 21554 5320 21606 5400
rect 21554 5286 21564 5320
rect 21598 5286 21606 5320
rect 21670 5300 21722 5422
rect 21752 5300 21794 5468
rect 21824 5430 21890 5468
rect 21824 5396 21834 5430
rect 21868 5396 21890 5430
rect 21824 5384 21890 5396
rect 21920 5456 21998 5468
rect 21920 5422 21942 5456
rect 21976 5422 21998 5456
rect 21920 5384 21998 5422
rect 22028 5384 22116 5468
rect 22146 5455 22200 5468
rect 22146 5421 22156 5455
rect 22190 5421 22200 5455
rect 22146 5384 22200 5421
rect 22230 5384 22344 5468
rect 21824 5300 21875 5384
rect 21554 5272 21606 5286
rect 21457 5268 21507 5272
rect 22292 5300 22344 5384
rect 22374 5456 22481 5468
rect 22374 5422 22431 5456
rect 22465 5422 22481 5456
rect 22374 5388 22481 5422
rect 22374 5354 22431 5388
rect 22465 5354 22481 5388
rect 22374 5300 22481 5354
rect 22511 5300 22565 5468
rect 22595 5430 22673 5468
rect 22595 5396 22605 5430
rect 22639 5396 22673 5430
rect 22595 5384 22673 5396
rect 22703 5446 22779 5468
rect 22703 5412 22725 5446
rect 22759 5412 22779 5446
rect 22703 5384 22779 5412
rect 22809 5384 22899 5468
rect 22929 5455 22983 5468
rect 22929 5421 22939 5455
rect 22973 5421 22983 5455
rect 22929 5384 22983 5421
rect 23013 5448 23076 5468
rect 23013 5414 23032 5448
rect 23066 5414 23076 5448
rect 23013 5384 23076 5414
rect 23106 5432 23158 5468
rect 23106 5398 23116 5432
rect 23150 5398 23158 5432
rect 23106 5384 23158 5398
rect 23212 5448 23264 5462
rect 23212 5414 23220 5448
rect 23254 5414 23264 5448
rect 22595 5362 22657 5384
rect 22595 5328 22605 5362
rect 22639 5328 22657 5362
rect 22595 5300 22657 5328
rect 23212 5380 23264 5414
rect 23212 5346 23220 5380
rect 23254 5346 23264 5380
rect 23212 5334 23264 5346
rect 23294 5432 23348 5462
rect 23294 5398 23304 5432
rect 23338 5398 23348 5432
rect 23294 5334 23348 5398
rect 23378 5448 23430 5462
rect 23378 5414 23388 5448
rect 23422 5414 23430 5448
rect 23378 5380 23430 5414
rect 23378 5346 23388 5380
rect 23422 5346 23430 5380
rect 23378 5334 23430 5346
rect 11116 4574 11168 4594
rect 11116 4540 11124 4574
rect 11158 4540 11168 4574
rect 11116 4506 11168 4540
rect 11116 4472 11124 4506
rect 11158 4472 11168 4506
rect 11116 4436 11168 4472
rect 11198 4574 11256 4594
rect 11198 4540 11210 4574
rect 11244 4540 11256 4574
rect 11198 4506 11256 4540
rect 11198 4472 11210 4506
rect 11244 4472 11256 4506
rect 11198 4436 11256 4472
rect 11286 4574 11338 4594
rect 11286 4540 11296 4574
rect 11330 4540 11338 4574
rect 11286 4493 11338 4540
rect 11286 4459 11296 4493
rect 11330 4459 11338 4493
rect 11286 4436 11338 4459
rect 11392 4576 11444 4594
rect 11392 4542 11400 4576
rect 11434 4542 11444 4576
rect 11392 4508 11444 4542
rect 11392 4474 11400 4508
rect 11434 4474 11444 4508
rect 11392 4440 11444 4474
rect 11392 4406 11400 4440
rect 11434 4406 11444 4440
rect 11392 4394 11444 4406
rect 11474 4582 11528 4594
rect 11474 4548 11484 4582
rect 11518 4548 11528 4582
rect 11474 4514 11528 4548
rect 11474 4480 11484 4514
rect 11518 4480 11528 4514
rect 11474 4394 11528 4480
rect 11558 4560 11612 4594
rect 11558 4526 11568 4560
rect 11602 4526 11612 4560
rect 11558 4465 11612 4526
rect 11558 4431 11568 4465
rect 11602 4431 11612 4465
rect 11558 4394 11612 4431
rect 11642 4582 11696 4594
rect 11642 4548 11652 4582
rect 11686 4548 11696 4582
rect 11642 4514 11696 4548
rect 11642 4480 11652 4514
rect 11686 4480 11696 4514
rect 11642 4394 11696 4480
rect 11726 4560 11780 4594
rect 11726 4526 11736 4560
rect 11770 4526 11780 4560
rect 11726 4465 11780 4526
rect 11726 4431 11736 4465
rect 11770 4431 11780 4465
rect 11726 4394 11780 4431
rect 11810 4582 11862 4594
rect 11810 4548 11820 4582
rect 11854 4548 11862 4582
rect 11810 4514 11862 4548
rect 11810 4480 11820 4514
rect 11854 4480 11862 4514
rect 11810 4446 11862 4480
rect 11810 4412 11820 4446
rect 11854 4412 11862 4446
rect 11810 4394 11862 4412
rect 13699 4583 13751 4595
rect 13699 4549 13707 4583
rect 13741 4549 13751 4583
rect 13699 4515 13751 4549
rect 13699 4481 13707 4515
rect 13741 4481 13751 4515
rect 13699 4447 13751 4481
rect 13699 4413 13707 4447
rect 13741 4413 13751 4447
rect 13699 4395 13751 4413
rect 13781 4583 13833 4595
rect 13781 4549 13791 4583
rect 13825 4549 13833 4583
rect 13781 4515 13833 4549
rect 13781 4481 13791 4515
rect 13825 4481 13833 4515
rect 13781 4447 13833 4481
rect 13915 4575 13967 4589
rect 13915 4541 13923 4575
rect 13957 4541 13967 4575
rect 13915 4507 13967 4541
rect 13915 4473 13923 4507
rect 13957 4473 13967 4507
rect 13915 4461 13967 4473
rect 13997 4559 14051 4589
rect 13997 4525 14007 4559
rect 14041 4525 14051 4559
rect 13997 4461 14051 4525
rect 14081 4575 14133 4589
rect 14081 4541 14091 4575
rect 14125 4541 14133 4575
rect 14081 4507 14133 4541
rect 14187 4559 14239 4595
rect 14187 4525 14195 4559
rect 14229 4525 14239 4559
rect 14187 4511 14239 4525
rect 14269 4575 14332 4595
rect 14269 4541 14279 4575
rect 14313 4541 14332 4575
rect 14269 4511 14332 4541
rect 14362 4582 14416 4595
rect 14362 4548 14372 4582
rect 14406 4548 14416 4582
rect 14362 4511 14416 4548
rect 14446 4511 14536 4595
rect 14566 4573 14642 4595
rect 14566 4539 14586 4573
rect 14620 4539 14642 4573
rect 14566 4511 14642 4539
rect 14672 4557 14750 4595
rect 14672 4523 14706 4557
rect 14740 4523 14750 4557
rect 14672 4511 14750 4523
rect 14081 4473 14091 4507
rect 14125 4473 14133 4507
rect 14081 4461 14133 4473
rect 13781 4413 13791 4447
rect 13825 4413 13833 4447
rect 13781 4395 13833 4413
rect 14688 4489 14750 4511
rect 14688 4455 14706 4489
rect 14740 4455 14750 4489
rect 14688 4427 14750 4455
rect 14780 4427 14834 4595
rect 14864 4583 14971 4595
rect 14864 4549 14880 4583
rect 14914 4549 14971 4583
rect 14864 4515 14971 4549
rect 14864 4481 14880 4515
rect 14914 4481 14971 4515
rect 14864 4427 14971 4481
rect 15001 4511 15115 4595
rect 15145 4582 15199 4595
rect 15145 4548 15155 4582
rect 15189 4548 15199 4582
rect 15145 4511 15199 4548
rect 15229 4511 15317 4595
rect 15347 4583 15425 4595
rect 15347 4549 15369 4583
rect 15403 4549 15425 4583
rect 15347 4511 15425 4549
rect 15455 4557 15521 4595
rect 15455 4523 15477 4557
rect 15511 4523 15521 4557
rect 15455 4511 15521 4523
rect 15001 4427 15053 4511
rect 15470 4427 15521 4511
rect 15551 4427 15593 4595
rect 15623 4583 15675 4595
rect 15623 4549 15633 4583
rect 15667 4549 15675 4583
rect 15836 4583 15888 4595
rect 15623 4427 15675 4549
rect 15836 4549 15844 4583
rect 15878 4549 15888 4583
rect 15836 4527 15888 4549
rect 15739 4447 15791 4527
rect 15739 4413 15747 4447
rect 15781 4413 15791 4447
rect 15739 4399 15791 4413
rect 15821 4399 15888 4527
rect 15838 4395 15888 4399
rect 15918 4546 15970 4595
rect 16121 4579 16171 4595
rect 15918 4512 15928 4546
rect 15962 4512 15970 4546
rect 15918 4478 15970 4512
rect 15918 4444 15928 4478
rect 15962 4444 15970 4478
rect 16024 4565 16076 4579
rect 16024 4531 16032 4565
rect 16066 4531 16076 4565
rect 16024 4497 16076 4531
rect 16024 4463 16032 4497
rect 16066 4463 16076 4497
rect 16024 4451 16076 4463
rect 16106 4571 16171 4579
rect 16106 4537 16127 4571
rect 16161 4537 16171 4571
rect 16106 4503 16171 4537
rect 16106 4469 16127 4503
rect 16161 4469 16171 4503
rect 16106 4451 16171 4469
rect 15918 4395 15970 4444
rect 16121 4395 16171 4451
rect 16201 4547 16253 4595
rect 16201 4513 16211 4547
rect 16245 4513 16253 4547
rect 16201 4479 16253 4513
rect 16201 4445 16211 4479
rect 16245 4445 16253 4479
rect 16307 4575 16359 4589
rect 16307 4541 16315 4575
rect 16349 4541 16359 4575
rect 16307 4507 16359 4541
rect 16307 4473 16315 4507
rect 16349 4473 16359 4507
rect 16307 4461 16359 4473
rect 16389 4559 16443 4589
rect 16389 4525 16399 4559
rect 16433 4525 16443 4559
rect 16389 4461 16443 4525
rect 16473 4575 16525 4589
rect 16473 4541 16483 4575
rect 16517 4541 16525 4575
rect 16473 4507 16525 4541
rect 16579 4559 16631 4595
rect 16579 4525 16587 4559
rect 16621 4525 16631 4559
rect 16579 4511 16631 4525
rect 16661 4575 16724 4595
rect 16661 4541 16671 4575
rect 16705 4541 16724 4575
rect 16661 4511 16724 4541
rect 16754 4582 16808 4595
rect 16754 4548 16764 4582
rect 16798 4548 16808 4582
rect 16754 4511 16808 4548
rect 16838 4511 16928 4595
rect 16958 4573 17034 4595
rect 16958 4539 16978 4573
rect 17012 4539 17034 4573
rect 16958 4511 17034 4539
rect 17064 4557 17142 4595
rect 17064 4523 17098 4557
rect 17132 4523 17142 4557
rect 17064 4511 17142 4523
rect 16473 4473 16483 4507
rect 16517 4473 16525 4507
rect 16473 4461 16525 4473
rect 16201 4395 16253 4445
rect 17080 4489 17142 4511
rect 17080 4455 17098 4489
rect 17132 4455 17142 4489
rect 17080 4427 17142 4455
rect 17172 4427 17226 4595
rect 17256 4583 17363 4595
rect 17256 4549 17272 4583
rect 17306 4549 17363 4583
rect 17256 4515 17363 4549
rect 17256 4481 17272 4515
rect 17306 4481 17363 4515
rect 17256 4427 17363 4481
rect 17393 4511 17507 4595
rect 17537 4582 17591 4595
rect 17537 4548 17547 4582
rect 17581 4548 17591 4582
rect 17537 4511 17591 4548
rect 17621 4511 17709 4595
rect 17739 4583 17817 4595
rect 17739 4549 17761 4583
rect 17795 4549 17817 4583
rect 17739 4511 17817 4549
rect 17847 4557 17913 4595
rect 17847 4523 17869 4557
rect 17903 4523 17913 4557
rect 17847 4511 17913 4523
rect 17393 4427 17445 4511
rect 17862 4427 17913 4511
rect 17943 4427 17985 4595
rect 18015 4583 18067 4595
rect 18015 4549 18025 4583
rect 18059 4549 18067 4583
rect 18228 4583 18280 4595
rect 18015 4427 18067 4549
rect 18228 4549 18236 4583
rect 18270 4549 18280 4583
rect 18228 4527 18280 4549
rect 18131 4447 18183 4527
rect 18131 4413 18139 4447
rect 18173 4413 18183 4447
rect 18131 4399 18183 4413
rect 18213 4399 18280 4527
rect 18230 4395 18280 4399
rect 18310 4546 18362 4595
rect 18513 4579 18563 4595
rect 18310 4512 18320 4546
rect 18354 4512 18362 4546
rect 18310 4478 18362 4512
rect 18310 4444 18320 4478
rect 18354 4444 18362 4478
rect 18416 4565 18468 4579
rect 18416 4531 18424 4565
rect 18458 4531 18468 4565
rect 18416 4497 18468 4531
rect 18416 4463 18424 4497
rect 18458 4463 18468 4497
rect 18416 4451 18468 4463
rect 18498 4571 18563 4579
rect 18498 4537 18519 4571
rect 18553 4537 18563 4571
rect 18498 4503 18563 4537
rect 18498 4469 18519 4503
rect 18553 4469 18563 4503
rect 18498 4451 18563 4469
rect 18310 4395 18362 4444
rect 18513 4395 18563 4451
rect 18593 4547 18645 4595
rect 18593 4513 18603 4547
rect 18637 4513 18645 4547
rect 18593 4479 18645 4513
rect 18593 4445 18603 4479
rect 18637 4445 18645 4479
rect 18699 4575 18751 4589
rect 18699 4541 18707 4575
rect 18741 4541 18751 4575
rect 18699 4507 18751 4541
rect 18699 4473 18707 4507
rect 18741 4473 18751 4507
rect 18699 4461 18751 4473
rect 18781 4559 18835 4589
rect 18781 4525 18791 4559
rect 18825 4525 18835 4559
rect 18781 4461 18835 4525
rect 18865 4575 18917 4589
rect 18865 4541 18875 4575
rect 18909 4541 18917 4575
rect 18865 4507 18917 4541
rect 18971 4559 19023 4595
rect 18971 4525 18979 4559
rect 19013 4525 19023 4559
rect 18971 4511 19023 4525
rect 19053 4575 19116 4595
rect 19053 4541 19063 4575
rect 19097 4541 19116 4575
rect 19053 4511 19116 4541
rect 19146 4582 19200 4595
rect 19146 4548 19156 4582
rect 19190 4548 19200 4582
rect 19146 4511 19200 4548
rect 19230 4511 19320 4595
rect 19350 4573 19426 4595
rect 19350 4539 19370 4573
rect 19404 4539 19426 4573
rect 19350 4511 19426 4539
rect 19456 4557 19534 4595
rect 19456 4523 19490 4557
rect 19524 4523 19534 4557
rect 19456 4511 19534 4523
rect 18865 4473 18875 4507
rect 18909 4473 18917 4507
rect 18865 4461 18917 4473
rect 18593 4395 18645 4445
rect 19472 4489 19534 4511
rect 19472 4455 19490 4489
rect 19524 4455 19534 4489
rect 19472 4427 19534 4455
rect 19564 4427 19618 4595
rect 19648 4583 19755 4595
rect 19648 4549 19664 4583
rect 19698 4549 19755 4583
rect 19648 4515 19755 4549
rect 19648 4481 19664 4515
rect 19698 4481 19755 4515
rect 19648 4427 19755 4481
rect 19785 4511 19899 4595
rect 19929 4582 19983 4595
rect 19929 4548 19939 4582
rect 19973 4548 19983 4582
rect 19929 4511 19983 4548
rect 20013 4511 20101 4595
rect 20131 4583 20209 4595
rect 20131 4549 20153 4583
rect 20187 4549 20209 4583
rect 20131 4511 20209 4549
rect 20239 4557 20305 4595
rect 20239 4523 20261 4557
rect 20295 4523 20305 4557
rect 20239 4511 20305 4523
rect 19785 4427 19837 4511
rect 20254 4427 20305 4511
rect 20335 4427 20377 4595
rect 20407 4583 20459 4595
rect 20407 4549 20417 4583
rect 20451 4549 20459 4583
rect 20620 4583 20672 4595
rect 20407 4427 20459 4549
rect 20620 4549 20628 4583
rect 20662 4549 20672 4583
rect 20620 4527 20672 4549
rect 20523 4447 20575 4527
rect 20523 4413 20531 4447
rect 20565 4413 20575 4447
rect 20523 4399 20575 4413
rect 20605 4399 20672 4527
rect 20622 4395 20672 4399
rect 20702 4546 20754 4595
rect 20905 4579 20955 4595
rect 20702 4512 20712 4546
rect 20746 4512 20754 4546
rect 20702 4478 20754 4512
rect 20702 4444 20712 4478
rect 20746 4444 20754 4478
rect 20808 4565 20860 4579
rect 20808 4531 20816 4565
rect 20850 4531 20860 4565
rect 20808 4497 20860 4531
rect 20808 4463 20816 4497
rect 20850 4463 20860 4497
rect 20808 4451 20860 4463
rect 20890 4571 20955 4579
rect 20890 4537 20911 4571
rect 20945 4537 20955 4571
rect 20890 4503 20955 4537
rect 20890 4469 20911 4503
rect 20945 4469 20955 4503
rect 20890 4451 20955 4469
rect 20702 4395 20754 4444
rect 20905 4395 20955 4451
rect 20985 4547 21037 4595
rect 20985 4513 20995 4547
rect 21029 4513 21037 4547
rect 20985 4479 21037 4513
rect 20985 4445 20995 4479
rect 21029 4445 21037 4479
rect 21091 4575 21143 4589
rect 21091 4541 21099 4575
rect 21133 4541 21143 4575
rect 21091 4507 21143 4541
rect 21091 4473 21099 4507
rect 21133 4473 21143 4507
rect 21091 4461 21143 4473
rect 21173 4559 21227 4589
rect 21173 4525 21183 4559
rect 21217 4525 21227 4559
rect 21173 4461 21227 4525
rect 21257 4575 21309 4589
rect 21257 4541 21267 4575
rect 21301 4541 21309 4575
rect 21257 4507 21309 4541
rect 21363 4559 21415 4595
rect 21363 4525 21371 4559
rect 21405 4525 21415 4559
rect 21363 4511 21415 4525
rect 21445 4575 21508 4595
rect 21445 4541 21455 4575
rect 21489 4541 21508 4575
rect 21445 4511 21508 4541
rect 21538 4582 21592 4595
rect 21538 4548 21548 4582
rect 21582 4548 21592 4582
rect 21538 4511 21592 4548
rect 21622 4511 21712 4595
rect 21742 4573 21818 4595
rect 21742 4539 21762 4573
rect 21796 4539 21818 4573
rect 21742 4511 21818 4539
rect 21848 4557 21926 4595
rect 21848 4523 21882 4557
rect 21916 4523 21926 4557
rect 21848 4511 21926 4523
rect 21257 4473 21267 4507
rect 21301 4473 21309 4507
rect 21257 4461 21309 4473
rect 20985 4395 21037 4445
rect 21864 4489 21926 4511
rect 21864 4455 21882 4489
rect 21916 4455 21926 4489
rect 21864 4427 21926 4455
rect 21956 4427 22010 4595
rect 22040 4583 22147 4595
rect 22040 4549 22056 4583
rect 22090 4549 22147 4583
rect 22040 4515 22147 4549
rect 22040 4481 22056 4515
rect 22090 4481 22147 4515
rect 22040 4427 22147 4481
rect 22177 4511 22291 4595
rect 22321 4582 22375 4595
rect 22321 4548 22331 4582
rect 22365 4548 22375 4582
rect 22321 4511 22375 4548
rect 22405 4511 22493 4595
rect 22523 4583 22601 4595
rect 22523 4549 22545 4583
rect 22579 4549 22601 4583
rect 22523 4511 22601 4549
rect 22631 4557 22697 4595
rect 22631 4523 22653 4557
rect 22687 4523 22697 4557
rect 22631 4511 22697 4523
rect 22177 4427 22229 4511
rect 22646 4427 22697 4511
rect 22727 4427 22769 4595
rect 22799 4583 22851 4595
rect 22799 4549 22809 4583
rect 22843 4549 22851 4583
rect 23012 4583 23064 4595
rect 22799 4427 22851 4549
rect 23012 4549 23020 4583
rect 23054 4549 23064 4583
rect 23012 4527 23064 4549
rect 22915 4447 22967 4527
rect 22915 4413 22923 4447
rect 22957 4413 22967 4447
rect 22915 4399 22967 4413
rect 22997 4399 23064 4527
rect 23014 4395 23064 4399
rect 23094 4546 23146 4595
rect 23297 4579 23347 4595
rect 23094 4512 23104 4546
rect 23138 4512 23146 4546
rect 23094 4478 23146 4512
rect 23094 4444 23104 4478
rect 23138 4444 23146 4478
rect 23200 4565 23252 4579
rect 23200 4531 23208 4565
rect 23242 4531 23252 4565
rect 23200 4497 23252 4531
rect 23200 4463 23208 4497
rect 23242 4463 23252 4497
rect 23200 4451 23252 4463
rect 23282 4571 23347 4579
rect 23282 4537 23303 4571
rect 23337 4537 23347 4571
rect 23282 4503 23347 4537
rect 23282 4469 23303 4503
rect 23337 4469 23347 4503
rect 23282 4451 23347 4469
rect 23094 4395 23146 4444
rect 23297 4395 23347 4451
rect 23377 4547 23429 4595
rect 23377 4513 23387 4547
rect 23421 4513 23429 4547
rect 23377 4479 23429 4513
rect 23377 4445 23387 4479
rect 23421 4445 23429 4479
rect 23377 4395 23429 4445
rect 25604 3906 25656 3918
rect 25604 3872 25612 3906
rect 25646 3872 25656 3906
rect 25604 3838 25656 3872
rect 25604 3804 25612 3838
rect 25646 3804 25656 3838
rect 25604 3790 25656 3804
rect 25686 3854 25740 3918
rect 25686 3820 25696 3854
rect 25730 3820 25740 3854
rect 25686 3790 25740 3820
rect 25770 3906 25822 3918
rect 25770 3872 25780 3906
rect 25814 3872 25822 3906
rect 25770 3838 25822 3872
rect 26377 3924 26439 3952
rect 26377 3890 26395 3924
rect 26429 3890 26439 3924
rect 26377 3868 26439 3890
rect 25770 3804 25780 3838
rect 25814 3804 25822 3838
rect 25770 3790 25822 3804
rect 25876 3854 25928 3868
rect 25876 3820 25884 3854
rect 25918 3820 25928 3854
rect 25876 3784 25928 3820
rect 25958 3838 26021 3868
rect 25958 3804 25968 3838
rect 26002 3804 26021 3838
rect 25958 3784 26021 3804
rect 26051 3831 26105 3868
rect 26051 3797 26061 3831
rect 26095 3797 26105 3831
rect 26051 3784 26105 3797
rect 26135 3784 26225 3868
rect 26255 3840 26331 3868
rect 26255 3806 26275 3840
rect 26309 3806 26331 3840
rect 26255 3784 26331 3806
rect 26361 3856 26439 3868
rect 26361 3822 26395 3856
rect 26429 3822 26439 3856
rect 26361 3784 26439 3822
rect 26469 3784 26523 3952
rect 26553 3898 26660 3952
rect 26553 3864 26569 3898
rect 26603 3864 26660 3898
rect 26553 3830 26660 3864
rect 26553 3796 26569 3830
rect 26603 3796 26660 3830
rect 26553 3784 26660 3796
rect 26690 3868 26742 3952
rect 27527 3980 27577 3984
rect 27428 3966 27480 3980
rect 27159 3868 27210 3952
rect 26690 3784 26804 3868
rect 26834 3831 26888 3868
rect 26834 3797 26844 3831
rect 26878 3797 26888 3831
rect 26834 3784 26888 3797
rect 26918 3784 27006 3868
rect 27036 3830 27114 3868
rect 27036 3796 27058 3830
rect 27092 3796 27114 3830
rect 27036 3784 27114 3796
rect 27144 3856 27210 3868
rect 27144 3822 27166 3856
rect 27200 3822 27210 3856
rect 27144 3784 27210 3822
rect 27240 3784 27282 3952
rect 27312 3830 27364 3952
rect 27428 3932 27436 3966
rect 27470 3932 27480 3966
rect 27428 3852 27480 3932
rect 27510 3852 27577 3980
rect 27312 3796 27322 3830
rect 27356 3796 27364 3830
rect 27525 3830 27577 3852
rect 27312 3784 27364 3796
rect 27525 3796 27533 3830
rect 27567 3796 27577 3830
rect 27525 3784 27577 3796
rect 27607 3935 27659 3984
rect 27607 3901 27617 3935
rect 27651 3901 27659 3935
rect 27810 3928 27860 3984
rect 27607 3867 27659 3901
rect 27607 3833 27617 3867
rect 27651 3833 27659 3867
rect 27607 3784 27659 3833
rect 27713 3916 27765 3928
rect 27713 3882 27721 3916
rect 27755 3882 27765 3916
rect 27713 3848 27765 3882
rect 27713 3814 27721 3848
rect 27755 3814 27765 3848
rect 27713 3800 27765 3814
rect 27795 3910 27860 3928
rect 27795 3876 27816 3910
rect 27850 3876 27860 3910
rect 27795 3842 27860 3876
rect 27795 3808 27816 3842
rect 27850 3808 27860 3842
rect 27795 3800 27860 3808
rect 27810 3784 27860 3800
rect 27890 3934 27942 3984
rect 27890 3900 27900 3934
rect 27934 3900 27942 3934
rect 27890 3866 27942 3900
rect 27890 3832 27900 3866
rect 27934 3832 27942 3866
rect 27890 3784 27942 3832
rect 27996 3906 28048 3918
rect 27996 3872 28004 3906
rect 28038 3872 28048 3906
rect 27996 3838 28048 3872
rect 27996 3804 28004 3838
rect 28038 3804 28048 3838
rect 27996 3790 28048 3804
rect 28078 3854 28132 3918
rect 28078 3820 28088 3854
rect 28122 3820 28132 3854
rect 28078 3790 28132 3820
rect 28162 3906 28214 3918
rect 28162 3872 28172 3906
rect 28206 3872 28214 3906
rect 28162 3838 28214 3872
rect 28769 3924 28831 3952
rect 28769 3890 28787 3924
rect 28821 3890 28831 3924
rect 28769 3868 28831 3890
rect 28162 3804 28172 3838
rect 28206 3804 28214 3838
rect 28162 3790 28214 3804
rect 28268 3854 28320 3868
rect 28268 3820 28276 3854
rect 28310 3820 28320 3854
rect 28268 3784 28320 3820
rect 28350 3838 28413 3868
rect 28350 3804 28360 3838
rect 28394 3804 28413 3838
rect 28350 3784 28413 3804
rect 28443 3831 28497 3868
rect 28443 3797 28453 3831
rect 28487 3797 28497 3831
rect 28443 3784 28497 3797
rect 28527 3784 28617 3868
rect 28647 3840 28723 3868
rect 28647 3806 28667 3840
rect 28701 3806 28723 3840
rect 28647 3784 28723 3806
rect 28753 3856 28831 3868
rect 28753 3822 28787 3856
rect 28821 3822 28831 3856
rect 28753 3784 28831 3822
rect 28861 3784 28915 3952
rect 28945 3898 29052 3952
rect 28945 3864 28961 3898
rect 28995 3864 29052 3898
rect 28945 3830 29052 3864
rect 28945 3796 28961 3830
rect 28995 3796 29052 3830
rect 28945 3784 29052 3796
rect 29082 3868 29134 3952
rect 29919 3980 29969 3984
rect 29820 3966 29872 3980
rect 29551 3868 29602 3952
rect 29082 3784 29196 3868
rect 29226 3831 29280 3868
rect 29226 3797 29236 3831
rect 29270 3797 29280 3831
rect 29226 3784 29280 3797
rect 29310 3784 29398 3868
rect 29428 3830 29506 3868
rect 29428 3796 29450 3830
rect 29484 3796 29506 3830
rect 29428 3784 29506 3796
rect 29536 3856 29602 3868
rect 29536 3822 29558 3856
rect 29592 3822 29602 3856
rect 29536 3784 29602 3822
rect 29632 3784 29674 3952
rect 29704 3830 29756 3952
rect 29820 3932 29828 3966
rect 29862 3932 29872 3966
rect 29820 3852 29872 3932
rect 29902 3852 29969 3980
rect 29704 3796 29714 3830
rect 29748 3796 29756 3830
rect 29917 3830 29969 3852
rect 29704 3784 29756 3796
rect 29917 3796 29925 3830
rect 29959 3796 29969 3830
rect 29917 3784 29969 3796
rect 29999 3935 30051 3984
rect 29999 3901 30009 3935
rect 30043 3901 30051 3935
rect 30202 3928 30252 3984
rect 29999 3867 30051 3901
rect 29999 3833 30009 3867
rect 30043 3833 30051 3867
rect 29999 3784 30051 3833
rect 30105 3916 30157 3928
rect 30105 3882 30113 3916
rect 30147 3882 30157 3916
rect 30105 3848 30157 3882
rect 30105 3814 30113 3848
rect 30147 3814 30157 3848
rect 30105 3800 30157 3814
rect 30187 3910 30252 3928
rect 30187 3876 30208 3910
rect 30242 3876 30252 3910
rect 30187 3842 30252 3876
rect 30187 3808 30208 3842
rect 30242 3808 30252 3842
rect 30187 3800 30252 3808
rect 30202 3784 30252 3800
rect 30282 3934 30334 3984
rect 30282 3900 30292 3934
rect 30326 3900 30334 3934
rect 30282 3866 30334 3900
rect 30282 3832 30292 3866
rect 30326 3832 30334 3866
rect 30282 3784 30334 3832
rect 11523 3674 11575 3722
rect 11523 3640 11531 3674
rect 11565 3640 11575 3674
rect 11523 3606 11575 3640
rect 11523 3572 11531 3606
rect 11565 3572 11575 3606
rect 11523 3522 11575 3572
rect 11605 3706 11655 3722
rect 11605 3698 11670 3706
rect 11605 3664 11615 3698
rect 11649 3664 11670 3698
rect 11605 3630 11670 3664
rect 11605 3596 11615 3630
rect 11649 3596 11670 3630
rect 11605 3578 11670 3596
rect 11700 3692 11752 3706
rect 11700 3658 11710 3692
rect 11744 3658 11752 3692
rect 11700 3624 11752 3658
rect 11700 3590 11710 3624
rect 11744 3590 11752 3624
rect 11700 3578 11752 3590
rect 11806 3673 11858 3722
rect 11806 3639 11814 3673
rect 11848 3639 11858 3673
rect 11806 3605 11858 3639
rect 11605 3522 11655 3578
rect 11806 3571 11814 3605
rect 11848 3571 11858 3605
rect 11806 3522 11858 3571
rect 11888 3710 11940 3722
rect 11888 3676 11898 3710
rect 11932 3676 11940 3710
rect 12101 3710 12153 3722
rect 11888 3654 11940 3676
rect 12101 3676 12109 3710
rect 12143 3676 12153 3710
rect 11888 3526 11955 3654
rect 11985 3574 12037 3654
rect 11985 3540 11995 3574
rect 12029 3540 12037 3574
rect 12101 3554 12153 3676
rect 12183 3554 12225 3722
rect 12255 3684 12321 3722
rect 12255 3650 12265 3684
rect 12299 3650 12321 3684
rect 12255 3638 12321 3650
rect 12351 3710 12429 3722
rect 12351 3676 12373 3710
rect 12407 3676 12429 3710
rect 12351 3638 12429 3676
rect 12459 3638 12547 3722
rect 12577 3709 12631 3722
rect 12577 3675 12587 3709
rect 12621 3675 12631 3709
rect 12577 3638 12631 3675
rect 12661 3638 12775 3722
rect 12255 3554 12306 3638
rect 11985 3526 12037 3540
rect 11888 3522 11938 3526
rect 12723 3554 12775 3638
rect 12805 3710 12912 3722
rect 12805 3676 12862 3710
rect 12896 3676 12912 3710
rect 12805 3642 12912 3676
rect 12805 3608 12862 3642
rect 12896 3608 12912 3642
rect 12805 3554 12912 3608
rect 12942 3554 12996 3722
rect 13026 3684 13104 3722
rect 13026 3650 13036 3684
rect 13070 3650 13104 3684
rect 13026 3638 13104 3650
rect 13134 3700 13210 3722
rect 13134 3666 13156 3700
rect 13190 3666 13210 3700
rect 13134 3638 13210 3666
rect 13240 3638 13330 3722
rect 13360 3709 13414 3722
rect 13360 3675 13370 3709
rect 13404 3675 13414 3709
rect 13360 3638 13414 3675
rect 13444 3702 13507 3722
rect 13444 3668 13463 3702
rect 13497 3668 13507 3702
rect 13444 3638 13507 3668
rect 13537 3686 13589 3722
rect 13537 3652 13547 3686
rect 13581 3652 13589 3686
rect 13537 3638 13589 3652
rect 13643 3702 13695 3716
rect 13643 3668 13651 3702
rect 13685 3668 13695 3702
rect 13026 3616 13088 3638
rect 13026 3582 13036 3616
rect 13070 3582 13088 3616
rect 13026 3554 13088 3582
rect 13643 3634 13695 3668
rect 13643 3600 13651 3634
rect 13685 3600 13695 3634
rect 13643 3588 13695 3600
rect 13725 3686 13779 3716
rect 13725 3652 13735 3686
rect 13769 3652 13779 3686
rect 13725 3588 13779 3652
rect 13809 3702 13861 3716
rect 13809 3668 13819 3702
rect 13853 3668 13861 3702
rect 13809 3634 13861 3668
rect 13809 3600 13819 3634
rect 13853 3600 13861 3634
rect 13809 3588 13861 3600
rect 13915 3674 13967 3722
rect 13915 3640 13923 3674
rect 13957 3640 13967 3674
rect 13915 3606 13967 3640
rect 13915 3572 13923 3606
rect 13957 3572 13967 3606
rect 13915 3522 13967 3572
rect 13997 3706 14047 3722
rect 13997 3698 14062 3706
rect 13997 3664 14007 3698
rect 14041 3664 14062 3698
rect 13997 3630 14062 3664
rect 13997 3596 14007 3630
rect 14041 3596 14062 3630
rect 13997 3578 14062 3596
rect 14092 3692 14144 3706
rect 14092 3658 14102 3692
rect 14136 3658 14144 3692
rect 14092 3624 14144 3658
rect 14092 3590 14102 3624
rect 14136 3590 14144 3624
rect 14092 3578 14144 3590
rect 14198 3673 14250 3722
rect 14198 3639 14206 3673
rect 14240 3639 14250 3673
rect 14198 3605 14250 3639
rect 13997 3522 14047 3578
rect 14198 3571 14206 3605
rect 14240 3571 14250 3605
rect 14198 3522 14250 3571
rect 14280 3710 14332 3722
rect 14280 3676 14290 3710
rect 14324 3676 14332 3710
rect 14493 3710 14545 3722
rect 14280 3654 14332 3676
rect 14493 3676 14501 3710
rect 14535 3676 14545 3710
rect 14280 3526 14347 3654
rect 14377 3574 14429 3654
rect 14377 3540 14387 3574
rect 14421 3540 14429 3574
rect 14493 3554 14545 3676
rect 14575 3554 14617 3722
rect 14647 3684 14713 3722
rect 14647 3650 14657 3684
rect 14691 3650 14713 3684
rect 14647 3638 14713 3650
rect 14743 3710 14821 3722
rect 14743 3676 14765 3710
rect 14799 3676 14821 3710
rect 14743 3638 14821 3676
rect 14851 3638 14939 3722
rect 14969 3709 15023 3722
rect 14969 3675 14979 3709
rect 15013 3675 15023 3709
rect 14969 3638 15023 3675
rect 15053 3638 15167 3722
rect 14647 3554 14698 3638
rect 14377 3526 14429 3540
rect 14280 3522 14330 3526
rect 15115 3554 15167 3638
rect 15197 3710 15304 3722
rect 15197 3676 15254 3710
rect 15288 3676 15304 3710
rect 15197 3642 15304 3676
rect 15197 3608 15254 3642
rect 15288 3608 15304 3642
rect 15197 3554 15304 3608
rect 15334 3554 15388 3722
rect 15418 3684 15496 3722
rect 15418 3650 15428 3684
rect 15462 3650 15496 3684
rect 15418 3638 15496 3650
rect 15526 3700 15602 3722
rect 15526 3666 15548 3700
rect 15582 3666 15602 3700
rect 15526 3638 15602 3666
rect 15632 3638 15722 3722
rect 15752 3709 15806 3722
rect 15752 3675 15762 3709
rect 15796 3675 15806 3709
rect 15752 3638 15806 3675
rect 15836 3702 15899 3722
rect 15836 3668 15855 3702
rect 15889 3668 15899 3702
rect 15836 3638 15899 3668
rect 15929 3686 15981 3722
rect 15929 3652 15939 3686
rect 15973 3652 15981 3686
rect 15929 3638 15981 3652
rect 16035 3702 16087 3716
rect 16035 3668 16043 3702
rect 16077 3668 16087 3702
rect 15418 3616 15480 3638
rect 15418 3582 15428 3616
rect 15462 3582 15480 3616
rect 15418 3554 15480 3582
rect 16035 3634 16087 3668
rect 16035 3600 16043 3634
rect 16077 3600 16087 3634
rect 16035 3588 16087 3600
rect 16117 3686 16171 3716
rect 16117 3652 16127 3686
rect 16161 3652 16171 3686
rect 16117 3588 16171 3652
rect 16201 3702 16253 3716
rect 16201 3668 16211 3702
rect 16245 3668 16253 3702
rect 16201 3634 16253 3668
rect 16201 3600 16211 3634
rect 16245 3600 16253 3634
rect 16201 3588 16253 3600
rect 16307 3674 16359 3722
rect 16307 3640 16315 3674
rect 16349 3640 16359 3674
rect 16307 3606 16359 3640
rect 16307 3572 16315 3606
rect 16349 3572 16359 3606
rect 16307 3522 16359 3572
rect 16389 3706 16439 3722
rect 16389 3698 16454 3706
rect 16389 3664 16399 3698
rect 16433 3664 16454 3698
rect 16389 3630 16454 3664
rect 16389 3596 16399 3630
rect 16433 3596 16454 3630
rect 16389 3578 16454 3596
rect 16484 3692 16536 3706
rect 16484 3658 16494 3692
rect 16528 3658 16536 3692
rect 16484 3624 16536 3658
rect 16484 3590 16494 3624
rect 16528 3590 16536 3624
rect 16484 3578 16536 3590
rect 16590 3673 16642 3722
rect 16590 3639 16598 3673
rect 16632 3639 16642 3673
rect 16590 3605 16642 3639
rect 16389 3522 16439 3578
rect 16590 3571 16598 3605
rect 16632 3571 16642 3605
rect 16590 3522 16642 3571
rect 16672 3710 16724 3722
rect 16672 3676 16682 3710
rect 16716 3676 16724 3710
rect 16885 3710 16937 3722
rect 16672 3654 16724 3676
rect 16885 3676 16893 3710
rect 16927 3676 16937 3710
rect 16672 3526 16739 3654
rect 16769 3574 16821 3654
rect 16769 3540 16779 3574
rect 16813 3540 16821 3574
rect 16885 3554 16937 3676
rect 16967 3554 17009 3722
rect 17039 3684 17105 3722
rect 17039 3650 17049 3684
rect 17083 3650 17105 3684
rect 17039 3638 17105 3650
rect 17135 3710 17213 3722
rect 17135 3676 17157 3710
rect 17191 3676 17213 3710
rect 17135 3638 17213 3676
rect 17243 3638 17331 3722
rect 17361 3709 17415 3722
rect 17361 3675 17371 3709
rect 17405 3675 17415 3709
rect 17361 3638 17415 3675
rect 17445 3638 17559 3722
rect 17039 3554 17090 3638
rect 16769 3526 16821 3540
rect 16672 3522 16722 3526
rect 17507 3554 17559 3638
rect 17589 3710 17696 3722
rect 17589 3676 17646 3710
rect 17680 3676 17696 3710
rect 17589 3642 17696 3676
rect 17589 3608 17646 3642
rect 17680 3608 17696 3642
rect 17589 3554 17696 3608
rect 17726 3554 17780 3722
rect 17810 3684 17888 3722
rect 17810 3650 17820 3684
rect 17854 3650 17888 3684
rect 17810 3638 17888 3650
rect 17918 3700 17994 3722
rect 17918 3666 17940 3700
rect 17974 3666 17994 3700
rect 17918 3638 17994 3666
rect 18024 3638 18114 3722
rect 18144 3709 18198 3722
rect 18144 3675 18154 3709
rect 18188 3675 18198 3709
rect 18144 3638 18198 3675
rect 18228 3702 18291 3722
rect 18228 3668 18247 3702
rect 18281 3668 18291 3702
rect 18228 3638 18291 3668
rect 18321 3686 18373 3722
rect 18321 3652 18331 3686
rect 18365 3652 18373 3686
rect 18321 3638 18373 3652
rect 18427 3702 18479 3716
rect 18427 3668 18435 3702
rect 18469 3668 18479 3702
rect 17810 3616 17872 3638
rect 17810 3582 17820 3616
rect 17854 3582 17872 3616
rect 17810 3554 17872 3582
rect 18427 3634 18479 3668
rect 18427 3600 18435 3634
rect 18469 3600 18479 3634
rect 18427 3588 18479 3600
rect 18509 3686 18563 3716
rect 18509 3652 18519 3686
rect 18553 3652 18563 3686
rect 18509 3588 18563 3652
rect 18593 3702 18645 3716
rect 18593 3668 18603 3702
rect 18637 3668 18645 3702
rect 18593 3634 18645 3668
rect 18593 3600 18603 3634
rect 18637 3600 18645 3634
rect 18593 3588 18645 3600
rect 18699 3674 18751 3722
rect 18699 3640 18707 3674
rect 18741 3640 18751 3674
rect 18699 3606 18751 3640
rect 18699 3572 18707 3606
rect 18741 3572 18751 3606
rect 18699 3522 18751 3572
rect 18781 3706 18831 3722
rect 18781 3698 18846 3706
rect 18781 3664 18791 3698
rect 18825 3664 18846 3698
rect 18781 3630 18846 3664
rect 18781 3596 18791 3630
rect 18825 3596 18846 3630
rect 18781 3578 18846 3596
rect 18876 3692 18928 3706
rect 18876 3658 18886 3692
rect 18920 3658 18928 3692
rect 18876 3624 18928 3658
rect 18876 3590 18886 3624
rect 18920 3590 18928 3624
rect 18876 3578 18928 3590
rect 18982 3673 19034 3722
rect 18982 3639 18990 3673
rect 19024 3639 19034 3673
rect 18982 3605 19034 3639
rect 18781 3522 18831 3578
rect 18982 3571 18990 3605
rect 19024 3571 19034 3605
rect 18982 3522 19034 3571
rect 19064 3710 19116 3722
rect 19064 3676 19074 3710
rect 19108 3676 19116 3710
rect 19277 3710 19329 3722
rect 19064 3654 19116 3676
rect 19277 3676 19285 3710
rect 19319 3676 19329 3710
rect 19064 3526 19131 3654
rect 19161 3574 19213 3654
rect 19161 3540 19171 3574
rect 19205 3540 19213 3574
rect 19277 3554 19329 3676
rect 19359 3554 19401 3722
rect 19431 3684 19497 3722
rect 19431 3650 19441 3684
rect 19475 3650 19497 3684
rect 19431 3638 19497 3650
rect 19527 3710 19605 3722
rect 19527 3676 19549 3710
rect 19583 3676 19605 3710
rect 19527 3638 19605 3676
rect 19635 3638 19723 3722
rect 19753 3709 19807 3722
rect 19753 3675 19763 3709
rect 19797 3675 19807 3709
rect 19753 3638 19807 3675
rect 19837 3638 19951 3722
rect 19431 3554 19482 3638
rect 19161 3526 19213 3540
rect 19064 3522 19114 3526
rect 19899 3554 19951 3638
rect 19981 3710 20088 3722
rect 19981 3676 20038 3710
rect 20072 3676 20088 3710
rect 19981 3642 20088 3676
rect 19981 3608 20038 3642
rect 20072 3608 20088 3642
rect 19981 3554 20088 3608
rect 20118 3554 20172 3722
rect 20202 3684 20280 3722
rect 20202 3650 20212 3684
rect 20246 3650 20280 3684
rect 20202 3638 20280 3650
rect 20310 3700 20386 3722
rect 20310 3666 20332 3700
rect 20366 3666 20386 3700
rect 20310 3638 20386 3666
rect 20416 3638 20506 3722
rect 20536 3709 20590 3722
rect 20536 3675 20546 3709
rect 20580 3675 20590 3709
rect 20536 3638 20590 3675
rect 20620 3702 20683 3722
rect 20620 3668 20639 3702
rect 20673 3668 20683 3702
rect 20620 3638 20683 3668
rect 20713 3686 20765 3722
rect 20713 3652 20723 3686
rect 20757 3652 20765 3686
rect 20713 3638 20765 3652
rect 20819 3702 20871 3716
rect 20819 3668 20827 3702
rect 20861 3668 20871 3702
rect 20202 3616 20264 3638
rect 20202 3582 20212 3616
rect 20246 3582 20264 3616
rect 20202 3554 20264 3582
rect 20819 3634 20871 3668
rect 20819 3600 20827 3634
rect 20861 3600 20871 3634
rect 20819 3588 20871 3600
rect 20901 3686 20955 3716
rect 20901 3652 20911 3686
rect 20945 3652 20955 3686
rect 20901 3588 20955 3652
rect 20985 3702 21037 3716
rect 20985 3668 20995 3702
rect 21029 3668 21037 3702
rect 20985 3634 21037 3668
rect 20985 3600 20995 3634
rect 21029 3600 21037 3634
rect 20985 3588 21037 3600
rect 21091 3674 21143 3722
rect 21091 3640 21099 3674
rect 21133 3640 21143 3674
rect 21091 3606 21143 3640
rect 21091 3572 21099 3606
rect 21133 3572 21143 3606
rect 21091 3522 21143 3572
rect 21173 3706 21223 3722
rect 21173 3698 21238 3706
rect 21173 3664 21183 3698
rect 21217 3664 21238 3698
rect 21173 3630 21238 3664
rect 21173 3596 21183 3630
rect 21217 3596 21238 3630
rect 21173 3578 21238 3596
rect 21268 3692 21320 3706
rect 21268 3658 21278 3692
rect 21312 3658 21320 3692
rect 21268 3624 21320 3658
rect 21268 3590 21278 3624
rect 21312 3590 21320 3624
rect 21268 3578 21320 3590
rect 21374 3673 21426 3722
rect 21374 3639 21382 3673
rect 21416 3639 21426 3673
rect 21374 3605 21426 3639
rect 21173 3522 21223 3578
rect 21374 3571 21382 3605
rect 21416 3571 21426 3605
rect 21374 3522 21426 3571
rect 21456 3710 21508 3722
rect 21456 3676 21466 3710
rect 21500 3676 21508 3710
rect 21669 3710 21721 3722
rect 21456 3654 21508 3676
rect 21669 3676 21677 3710
rect 21711 3676 21721 3710
rect 21456 3526 21523 3654
rect 21553 3574 21605 3654
rect 21553 3540 21563 3574
rect 21597 3540 21605 3574
rect 21669 3554 21721 3676
rect 21751 3554 21793 3722
rect 21823 3684 21889 3722
rect 21823 3650 21833 3684
rect 21867 3650 21889 3684
rect 21823 3638 21889 3650
rect 21919 3710 21997 3722
rect 21919 3676 21941 3710
rect 21975 3676 21997 3710
rect 21919 3638 21997 3676
rect 22027 3638 22115 3722
rect 22145 3709 22199 3722
rect 22145 3675 22155 3709
rect 22189 3675 22199 3709
rect 22145 3638 22199 3675
rect 22229 3638 22343 3722
rect 21823 3554 21874 3638
rect 21553 3526 21605 3540
rect 21456 3522 21506 3526
rect 22291 3554 22343 3638
rect 22373 3710 22480 3722
rect 22373 3676 22430 3710
rect 22464 3676 22480 3710
rect 22373 3642 22480 3676
rect 22373 3608 22430 3642
rect 22464 3608 22480 3642
rect 22373 3554 22480 3608
rect 22510 3554 22564 3722
rect 22594 3684 22672 3722
rect 22594 3650 22604 3684
rect 22638 3650 22672 3684
rect 22594 3638 22672 3650
rect 22702 3700 22778 3722
rect 22702 3666 22724 3700
rect 22758 3666 22778 3700
rect 22702 3638 22778 3666
rect 22808 3638 22898 3722
rect 22928 3709 22982 3722
rect 22928 3675 22938 3709
rect 22972 3675 22982 3709
rect 22928 3638 22982 3675
rect 23012 3702 23075 3722
rect 23012 3668 23031 3702
rect 23065 3668 23075 3702
rect 23012 3638 23075 3668
rect 23105 3686 23157 3722
rect 23105 3652 23115 3686
rect 23149 3652 23157 3686
rect 23105 3638 23157 3652
rect 23211 3702 23263 3716
rect 23211 3668 23219 3702
rect 23253 3668 23263 3702
rect 22594 3616 22656 3638
rect 22594 3582 22604 3616
rect 22638 3582 22656 3616
rect 22594 3554 22656 3582
rect 23211 3634 23263 3668
rect 23211 3600 23219 3634
rect 23253 3600 23263 3634
rect 23211 3588 23263 3600
rect 23293 3686 23347 3716
rect 23293 3652 23303 3686
rect 23337 3652 23347 3686
rect 23293 3588 23347 3652
rect 23377 3702 23429 3716
rect 23377 3668 23387 3702
rect 23421 3668 23429 3702
rect 23377 3634 23429 3668
rect 23377 3600 23387 3634
rect 23421 3600 23429 3634
rect 23377 3588 23429 3600
rect 25604 3574 25656 3588
rect 25604 3540 25612 3574
rect 25646 3540 25656 3574
rect 25604 3506 25656 3540
rect 25604 3472 25612 3506
rect 25646 3472 25656 3506
rect 25604 3460 25656 3472
rect 25686 3558 25740 3588
rect 25686 3524 25696 3558
rect 25730 3524 25740 3558
rect 25686 3460 25740 3524
rect 25770 3574 25822 3588
rect 25770 3540 25780 3574
rect 25814 3540 25822 3574
rect 25770 3506 25822 3540
rect 25876 3558 25928 3594
rect 25876 3524 25884 3558
rect 25918 3524 25928 3558
rect 25876 3510 25928 3524
rect 25958 3574 26021 3594
rect 25958 3540 25968 3574
rect 26002 3540 26021 3574
rect 25958 3510 26021 3540
rect 26051 3581 26105 3594
rect 26051 3547 26061 3581
rect 26095 3547 26105 3581
rect 26051 3510 26105 3547
rect 26135 3510 26225 3594
rect 26255 3572 26331 3594
rect 26255 3538 26275 3572
rect 26309 3538 26331 3572
rect 26255 3510 26331 3538
rect 26361 3556 26439 3594
rect 26361 3522 26395 3556
rect 26429 3522 26439 3556
rect 26361 3510 26439 3522
rect 25770 3472 25780 3506
rect 25814 3472 25822 3506
rect 25770 3460 25822 3472
rect 26377 3488 26439 3510
rect 26377 3454 26395 3488
rect 26429 3454 26439 3488
rect 26377 3426 26439 3454
rect 26469 3426 26523 3594
rect 26553 3582 26660 3594
rect 26553 3548 26569 3582
rect 26603 3548 26660 3582
rect 26553 3514 26660 3548
rect 26553 3480 26569 3514
rect 26603 3480 26660 3514
rect 26553 3426 26660 3480
rect 26690 3510 26804 3594
rect 26834 3581 26888 3594
rect 26834 3547 26844 3581
rect 26878 3547 26888 3581
rect 26834 3510 26888 3547
rect 26918 3510 27006 3594
rect 27036 3582 27114 3594
rect 27036 3548 27058 3582
rect 27092 3548 27114 3582
rect 27036 3510 27114 3548
rect 27144 3556 27210 3594
rect 27144 3522 27166 3556
rect 27200 3522 27210 3556
rect 27144 3510 27210 3522
rect 26690 3426 26742 3510
rect 27159 3426 27210 3510
rect 27240 3426 27282 3594
rect 27312 3582 27364 3594
rect 27312 3548 27322 3582
rect 27356 3548 27364 3582
rect 27525 3582 27577 3594
rect 27312 3426 27364 3548
rect 27525 3548 27533 3582
rect 27567 3548 27577 3582
rect 27525 3526 27577 3548
rect 27428 3446 27480 3526
rect 27428 3412 27436 3446
rect 27470 3412 27480 3446
rect 27428 3398 27480 3412
rect 27510 3398 27577 3526
rect 27527 3394 27577 3398
rect 27607 3545 27659 3594
rect 27810 3578 27860 3594
rect 27607 3511 27617 3545
rect 27651 3511 27659 3545
rect 27607 3477 27659 3511
rect 27607 3443 27617 3477
rect 27651 3443 27659 3477
rect 27713 3564 27765 3578
rect 27713 3530 27721 3564
rect 27755 3530 27765 3564
rect 27713 3496 27765 3530
rect 27713 3462 27721 3496
rect 27755 3462 27765 3496
rect 27713 3450 27765 3462
rect 27795 3570 27860 3578
rect 27795 3536 27816 3570
rect 27850 3536 27860 3570
rect 27795 3502 27860 3536
rect 27795 3468 27816 3502
rect 27850 3468 27860 3502
rect 27795 3450 27860 3468
rect 27607 3394 27659 3443
rect 27810 3394 27860 3450
rect 27890 3546 27942 3594
rect 27890 3512 27900 3546
rect 27934 3512 27942 3546
rect 27890 3478 27942 3512
rect 27890 3444 27900 3478
rect 27934 3444 27942 3478
rect 27996 3574 28048 3588
rect 27996 3540 28004 3574
rect 28038 3540 28048 3574
rect 27996 3506 28048 3540
rect 27996 3472 28004 3506
rect 28038 3472 28048 3506
rect 27996 3460 28048 3472
rect 28078 3558 28132 3588
rect 28078 3524 28088 3558
rect 28122 3524 28132 3558
rect 28078 3460 28132 3524
rect 28162 3574 28214 3588
rect 28162 3540 28172 3574
rect 28206 3540 28214 3574
rect 28162 3506 28214 3540
rect 28268 3558 28320 3594
rect 28268 3524 28276 3558
rect 28310 3524 28320 3558
rect 28268 3510 28320 3524
rect 28350 3574 28413 3594
rect 28350 3540 28360 3574
rect 28394 3540 28413 3574
rect 28350 3510 28413 3540
rect 28443 3581 28497 3594
rect 28443 3547 28453 3581
rect 28487 3547 28497 3581
rect 28443 3510 28497 3547
rect 28527 3510 28617 3594
rect 28647 3572 28723 3594
rect 28647 3538 28667 3572
rect 28701 3538 28723 3572
rect 28647 3510 28723 3538
rect 28753 3556 28831 3594
rect 28753 3522 28787 3556
rect 28821 3522 28831 3556
rect 28753 3510 28831 3522
rect 28162 3472 28172 3506
rect 28206 3472 28214 3506
rect 28162 3460 28214 3472
rect 27890 3394 27942 3444
rect 28769 3488 28831 3510
rect 28769 3454 28787 3488
rect 28821 3454 28831 3488
rect 28769 3426 28831 3454
rect 28861 3426 28915 3594
rect 28945 3582 29052 3594
rect 28945 3548 28961 3582
rect 28995 3548 29052 3582
rect 28945 3514 29052 3548
rect 28945 3480 28961 3514
rect 28995 3480 29052 3514
rect 28945 3426 29052 3480
rect 29082 3510 29196 3594
rect 29226 3581 29280 3594
rect 29226 3547 29236 3581
rect 29270 3547 29280 3581
rect 29226 3510 29280 3547
rect 29310 3510 29398 3594
rect 29428 3582 29506 3594
rect 29428 3548 29450 3582
rect 29484 3548 29506 3582
rect 29428 3510 29506 3548
rect 29536 3556 29602 3594
rect 29536 3522 29558 3556
rect 29592 3522 29602 3556
rect 29536 3510 29602 3522
rect 29082 3426 29134 3510
rect 29551 3426 29602 3510
rect 29632 3426 29674 3594
rect 29704 3582 29756 3594
rect 29704 3548 29714 3582
rect 29748 3548 29756 3582
rect 29917 3582 29969 3594
rect 29704 3426 29756 3548
rect 29917 3548 29925 3582
rect 29959 3548 29969 3582
rect 29917 3526 29969 3548
rect 29820 3446 29872 3526
rect 29820 3412 29828 3446
rect 29862 3412 29872 3446
rect 29820 3398 29872 3412
rect 29902 3398 29969 3526
rect 29919 3394 29969 3398
rect 29999 3545 30051 3594
rect 30202 3578 30252 3594
rect 29999 3511 30009 3545
rect 30043 3511 30051 3545
rect 29999 3477 30051 3511
rect 29999 3443 30009 3477
rect 30043 3443 30051 3477
rect 30105 3564 30157 3578
rect 30105 3530 30113 3564
rect 30147 3530 30157 3564
rect 30105 3496 30157 3530
rect 30105 3462 30113 3496
rect 30147 3462 30157 3496
rect 30105 3450 30157 3462
rect 30187 3570 30252 3578
rect 30187 3536 30208 3570
rect 30242 3536 30252 3570
rect 30187 3502 30252 3536
rect 30187 3468 30208 3502
rect 30242 3468 30252 3502
rect 30187 3450 30252 3468
rect 29999 3394 30051 3443
rect 30202 3394 30252 3450
rect 30282 3546 30334 3594
rect 30282 3512 30292 3546
rect 30326 3512 30334 3546
rect 30282 3478 30334 3512
rect 30282 3444 30292 3478
rect 30326 3444 30334 3478
rect 30282 3394 30334 3444
rect 25604 2626 25656 2638
rect 25604 2592 25612 2626
rect 25646 2592 25656 2626
rect 25604 2558 25656 2592
rect 25604 2524 25612 2558
rect 25646 2524 25656 2558
rect 25604 2510 25656 2524
rect 25686 2574 25740 2638
rect 25686 2540 25696 2574
rect 25730 2540 25740 2574
rect 25686 2510 25740 2540
rect 25770 2626 25822 2638
rect 25770 2592 25780 2626
rect 25814 2592 25822 2626
rect 25770 2558 25822 2592
rect 26377 2644 26439 2672
rect 26377 2610 26395 2644
rect 26429 2610 26439 2644
rect 26377 2588 26439 2610
rect 25770 2524 25780 2558
rect 25814 2524 25822 2558
rect 25770 2510 25822 2524
rect 25876 2574 25928 2588
rect 25876 2540 25884 2574
rect 25918 2540 25928 2574
rect 25876 2504 25928 2540
rect 25958 2558 26021 2588
rect 25958 2524 25968 2558
rect 26002 2524 26021 2558
rect 25958 2504 26021 2524
rect 26051 2551 26105 2588
rect 26051 2517 26061 2551
rect 26095 2517 26105 2551
rect 26051 2504 26105 2517
rect 26135 2504 26225 2588
rect 26255 2560 26331 2588
rect 26255 2526 26275 2560
rect 26309 2526 26331 2560
rect 26255 2504 26331 2526
rect 26361 2576 26439 2588
rect 26361 2542 26395 2576
rect 26429 2542 26439 2576
rect 26361 2504 26439 2542
rect 26469 2504 26523 2672
rect 26553 2618 26660 2672
rect 26553 2584 26569 2618
rect 26603 2584 26660 2618
rect 26553 2550 26660 2584
rect 26553 2516 26569 2550
rect 26603 2516 26660 2550
rect 26553 2504 26660 2516
rect 26690 2588 26742 2672
rect 27527 2700 27577 2704
rect 27428 2686 27480 2700
rect 27159 2588 27210 2672
rect 26690 2504 26804 2588
rect 26834 2551 26888 2588
rect 26834 2517 26844 2551
rect 26878 2517 26888 2551
rect 26834 2504 26888 2517
rect 26918 2504 27006 2588
rect 27036 2550 27114 2588
rect 27036 2516 27058 2550
rect 27092 2516 27114 2550
rect 27036 2504 27114 2516
rect 27144 2576 27210 2588
rect 27144 2542 27166 2576
rect 27200 2542 27210 2576
rect 27144 2504 27210 2542
rect 27240 2504 27282 2672
rect 27312 2550 27364 2672
rect 27428 2652 27436 2686
rect 27470 2652 27480 2686
rect 27428 2572 27480 2652
rect 27510 2572 27577 2700
rect 27312 2516 27322 2550
rect 27356 2516 27364 2550
rect 27525 2550 27577 2572
rect 27312 2504 27364 2516
rect 27525 2516 27533 2550
rect 27567 2516 27577 2550
rect 27525 2504 27577 2516
rect 27607 2655 27659 2704
rect 27607 2621 27617 2655
rect 27651 2621 27659 2655
rect 27810 2648 27860 2704
rect 27607 2587 27659 2621
rect 27607 2553 27617 2587
rect 27651 2553 27659 2587
rect 27607 2504 27659 2553
rect 27713 2636 27765 2648
rect 27713 2602 27721 2636
rect 27755 2602 27765 2636
rect 27713 2568 27765 2602
rect 27713 2534 27721 2568
rect 27755 2534 27765 2568
rect 27713 2520 27765 2534
rect 27795 2630 27860 2648
rect 27795 2596 27816 2630
rect 27850 2596 27860 2630
rect 27795 2562 27860 2596
rect 27795 2528 27816 2562
rect 27850 2528 27860 2562
rect 27795 2520 27860 2528
rect 27810 2504 27860 2520
rect 27890 2654 27942 2704
rect 27890 2620 27900 2654
rect 27934 2620 27942 2654
rect 27890 2586 27942 2620
rect 27890 2552 27900 2586
rect 27934 2552 27942 2586
rect 27890 2504 27942 2552
rect 27996 2626 28048 2638
rect 27996 2592 28004 2626
rect 28038 2592 28048 2626
rect 27996 2558 28048 2592
rect 27996 2524 28004 2558
rect 28038 2524 28048 2558
rect 27996 2510 28048 2524
rect 28078 2574 28132 2638
rect 28078 2540 28088 2574
rect 28122 2540 28132 2574
rect 28078 2510 28132 2540
rect 28162 2626 28214 2638
rect 28162 2592 28172 2626
rect 28206 2592 28214 2626
rect 28162 2558 28214 2592
rect 28769 2644 28831 2672
rect 28769 2610 28787 2644
rect 28821 2610 28831 2644
rect 28769 2588 28831 2610
rect 28162 2524 28172 2558
rect 28206 2524 28214 2558
rect 28162 2510 28214 2524
rect 28268 2574 28320 2588
rect 28268 2540 28276 2574
rect 28310 2540 28320 2574
rect 28268 2504 28320 2540
rect 28350 2558 28413 2588
rect 28350 2524 28360 2558
rect 28394 2524 28413 2558
rect 28350 2504 28413 2524
rect 28443 2551 28497 2588
rect 28443 2517 28453 2551
rect 28487 2517 28497 2551
rect 28443 2504 28497 2517
rect 28527 2504 28617 2588
rect 28647 2560 28723 2588
rect 28647 2526 28667 2560
rect 28701 2526 28723 2560
rect 28647 2504 28723 2526
rect 28753 2576 28831 2588
rect 28753 2542 28787 2576
rect 28821 2542 28831 2576
rect 28753 2504 28831 2542
rect 28861 2504 28915 2672
rect 28945 2618 29052 2672
rect 28945 2584 28961 2618
rect 28995 2584 29052 2618
rect 28945 2550 29052 2584
rect 28945 2516 28961 2550
rect 28995 2516 29052 2550
rect 28945 2504 29052 2516
rect 29082 2588 29134 2672
rect 29919 2700 29969 2704
rect 29820 2686 29872 2700
rect 29551 2588 29602 2672
rect 29082 2504 29196 2588
rect 29226 2551 29280 2588
rect 29226 2517 29236 2551
rect 29270 2517 29280 2551
rect 29226 2504 29280 2517
rect 29310 2504 29398 2588
rect 29428 2550 29506 2588
rect 29428 2516 29450 2550
rect 29484 2516 29506 2550
rect 29428 2504 29506 2516
rect 29536 2576 29602 2588
rect 29536 2542 29558 2576
rect 29592 2542 29602 2576
rect 29536 2504 29602 2542
rect 29632 2504 29674 2672
rect 29704 2550 29756 2672
rect 29820 2652 29828 2686
rect 29862 2652 29872 2686
rect 29820 2572 29872 2652
rect 29902 2572 29969 2700
rect 29704 2516 29714 2550
rect 29748 2516 29756 2550
rect 29917 2550 29969 2572
rect 29704 2504 29756 2516
rect 29917 2516 29925 2550
rect 29959 2516 29969 2550
rect 29917 2504 29969 2516
rect 29999 2655 30051 2704
rect 29999 2621 30009 2655
rect 30043 2621 30051 2655
rect 30202 2648 30252 2704
rect 29999 2587 30051 2621
rect 29999 2553 30009 2587
rect 30043 2553 30051 2587
rect 29999 2504 30051 2553
rect 30105 2636 30157 2648
rect 30105 2602 30113 2636
rect 30147 2602 30157 2636
rect 30105 2568 30157 2602
rect 30105 2534 30113 2568
rect 30147 2534 30157 2568
rect 30105 2520 30157 2534
rect 30187 2630 30252 2648
rect 30187 2596 30208 2630
rect 30242 2596 30252 2630
rect 30187 2562 30252 2596
rect 30187 2528 30208 2562
rect 30242 2528 30252 2562
rect 30187 2520 30252 2528
rect 30202 2504 30252 2520
rect 30282 2654 30334 2704
rect 30282 2620 30292 2654
rect 30326 2620 30334 2654
rect 30282 2586 30334 2620
rect 30282 2552 30292 2586
rect 30326 2552 30334 2586
rect 30282 2504 30334 2552
rect 25604 2294 25656 2308
rect 25604 2260 25612 2294
rect 25646 2260 25656 2294
rect 25604 2226 25656 2260
rect 25604 2192 25612 2226
rect 25646 2192 25656 2226
rect 25604 2180 25656 2192
rect 25686 2278 25740 2308
rect 25686 2244 25696 2278
rect 25730 2244 25740 2278
rect 25686 2180 25740 2244
rect 25770 2294 25822 2308
rect 25770 2260 25780 2294
rect 25814 2260 25822 2294
rect 25770 2226 25822 2260
rect 25876 2278 25928 2314
rect 25876 2244 25884 2278
rect 25918 2244 25928 2278
rect 25876 2230 25928 2244
rect 25958 2294 26021 2314
rect 25958 2260 25968 2294
rect 26002 2260 26021 2294
rect 25958 2230 26021 2260
rect 26051 2301 26105 2314
rect 26051 2267 26061 2301
rect 26095 2267 26105 2301
rect 26051 2230 26105 2267
rect 26135 2230 26225 2314
rect 26255 2292 26331 2314
rect 26255 2258 26275 2292
rect 26309 2258 26331 2292
rect 26255 2230 26331 2258
rect 26361 2276 26439 2314
rect 26361 2242 26395 2276
rect 26429 2242 26439 2276
rect 26361 2230 26439 2242
rect 25770 2192 25780 2226
rect 25814 2192 25822 2226
rect 25770 2180 25822 2192
rect 26377 2208 26439 2230
rect 26377 2174 26395 2208
rect 26429 2174 26439 2208
rect 26377 2146 26439 2174
rect 26469 2146 26523 2314
rect 26553 2302 26660 2314
rect 26553 2268 26569 2302
rect 26603 2268 26660 2302
rect 26553 2234 26660 2268
rect 26553 2200 26569 2234
rect 26603 2200 26660 2234
rect 26553 2146 26660 2200
rect 26690 2230 26804 2314
rect 26834 2301 26888 2314
rect 26834 2267 26844 2301
rect 26878 2267 26888 2301
rect 26834 2230 26888 2267
rect 26918 2230 27006 2314
rect 27036 2302 27114 2314
rect 27036 2268 27058 2302
rect 27092 2268 27114 2302
rect 27036 2230 27114 2268
rect 27144 2276 27210 2314
rect 27144 2242 27166 2276
rect 27200 2242 27210 2276
rect 27144 2230 27210 2242
rect 26690 2146 26742 2230
rect 27159 2146 27210 2230
rect 27240 2146 27282 2314
rect 27312 2302 27364 2314
rect 27312 2268 27322 2302
rect 27356 2268 27364 2302
rect 27525 2302 27577 2314
rect 27312 2146 27364 2268
rect 27525 2268 27533 2302
rect 27567 2268 27577 2302
rect 27525 2246 27577 2268
rect 27428 2166 27480 2246
rect 27428 2132 27436 2166
rect 27470 2132 27480 2166
rect 27428 2118 27480 2132
rect 27510 2118 27577 2246
rect 27527 2114 27577 2118
rect 27607 2265 27659 2314
rect 27810 2298 27860 2314
rect 27607 2231 27617 2265
rect 27651 2231 27659 2265
rect 27607 2197 27659 2231
rect 27607 2163 27617 2197
rect 27651 2163 27659 2197
rect 27713 2284 27765 2298
rect 27713 2250 27721 2284
rect 27755 2250 27765 2284
rect 27713 2216 27765 2250
rect 27713 2182 27721 2216
rect 27755 2182 27765 2216
rect 27713 2170 27765 2182
rect 27795 2290 27860 2298
rect 27795 2256 27816 2290
rect 27850 2256 27860 2290
rect 27795 2222 27860 2256
rect 27795 2188 27816 2222
rect 27850 2188 27860 2222
rect 27795 2170 27860 2188
rect 27607 2114 27659 2163
rect 27810 2114 27860 2170
rect 27890 2266 27942 2314
rect 27890 2232 27900 2266
rect 27934 2232 27942 2266
rect 27890 2198 27942 2232
rect 27890 2164 27900 2198
rect 27934 2164 27942 2198
rect 27996 2294 28048 2308
rect 27996 2260 28004 2294
rect 28038 2260 28048 2294
rect 27996 2226 28048 2260
rect 27996 2192 28004 2226
rect 28038 2192 28048 2226
rect 27996 2180 28048 2192
rect 28078 2278 28132 2308
rect 28078 2244 28088 2278
rect 28122 2244 28132 2278
rect 28078 2180 28132 2244
rect 28162 2294 28214 2308
rect 28162 2260 28172 2294
rect 28206 2260 28214 2294
rect 28162 2226 28214 2260
rect 28268 2278 28320 2314
rect 28268 2244 28276 2278
rect 28310 2244 28320 2278
rect 28268 2230 28320 2244
rect 28350 2294 28413 2314
rect 28350 2260 28360 2294
rect 28394 2260 28413 2294
rect 28350 2230 28413 2260
rect 28443 2301 28497 2314
rect 28443 2267 28453 2301
rect 28487 2267 28497 2301
rect 28443 2230 28497 2267
rect 28527 2230 28617 2314
rect 28647 2292 28723 2314
rect 28647 2258 28667 2292
rect 28701 2258 28723 2292
rect 28647 2230 28723 2258
rect 28753 2276 28831 2314
rect 28753 2242 28787 2276
rect 28821 2242 28831 2276
rect 28753 2230 28831 2242
rect 28162 2192 28172 2226
rect 28206 2192 28214 2226
rect 28162 2180 28214 2192
rect 27890 2114 27942 2164
rect 28769 2208 28831 2230
rect 28769 2174 28787 2208
rect 28821 2174 28831 2208
rect 28769 2146 28831 2174
rect 28861 2146 28915 2314
rect 28945 2302 29052 2314
rect 28945 2268 28961 2302
rect 28995 2268 29052 2302
rect 28945 2234 29052 2268
rect 28945 2200 28961 2234
rect 28995 2200 29052 2234
rect 28945 2146 29052 2200
rect 29082 2230 29196 2314
rect 29226 2301 29280 2314
rect 29226 2267 29236 2301
rect 29270 2267 29280 2301
rect 29226 2230 29280 2267
rect 29310 2230 29398 2314
rect 29428 2302 29506 2314
rect 29428 2268 29450 2302
rect 29484 2268 29506 2302
rect 29428 2230 29506 2268
rect 29536 2276 29602 2314
rect 29536 2242 29558 2276
rect 29592 2242 29602 2276
rect 29536 2230 29602 2242
rect 29082 2146 29134 2230
rect 29551 2146 29602 2230
rect 29632 2146 29674 2314
rect 29704 2302 29756 2314
rect 29704 2268 29714 2302
rect 29748 2268 29756 2302
rect 29917 2302 29969 2314
rect 29704 2146 29756 2268
rect 29917 2268 29925 2302
rect 29959 2268 29969 2302
rect 29917 2246 29969 2268
rect 29820 2166 29872 2246
rect 29820 2132 29828 2166
rect 29862 2132 29872 2166
rect 29820 2118 29872 2132
rect 29902 2118 29969 2246
rect 29919 2114 29969 2118
rect 29999 2265 30051 2314
rect 30202 2298 30252 2314
rect 29999 2231 30009 2265
rect 30043 2231 30051 2265
rect 29999 2197 30051 2231
rect 29999 2163 30009 2197
rect 30043 2163 30051 2197
rect 30105 2284 30157 2298
rect 30105 2250 30113 2284
rect 30147 2250 30157 2284
rect 30105 2216 30157 2250
rect 30105 2182 30113 2216
rect 30147 2182 30157 2216
rect 30105 2170 30157 2182
rect 30187 2290 30252 2298
rect 30187 2256 30208 2290
rect 30242 2256 30252 2290
rect 30187 2222 30252 2256
rect 30187 2188 30208 2222
rect 30242 2188 30252 2222
rect 30187 2170 30252 2188
rect 29999 2114 30051 2163
rect 30202 2114 30252 2170
rect 30282 2266 30334 2314
rect 30282 2232 30292 2266
rect 30326 2232 30334 2266
rect 30282 2198 30334 2232
rect 30282 2164 30292 2198
rect 30326 2164 30334 2198
rect 30282 2114 30334 2164
rect 8604 1322 8656 1342
rect 8604 1288 8612 1322
rect 8646 1288 8656 1322
rect 8604 1254 8656 1288
rect 8604 1220 8612 1254
rect 8646 1220 8656 1254
rect 8604 1184 8656 1220
rect 8686 1322 8744 1342
rect 8686 1288 8698 1322
rect 8732 1288 8744 1322
rect 8686 1254 8744 1288
rect 8686 1220 8698 1254
rect 8732 1220 8744 1254
rect 8686 1184 8744 1220
rect 8774 1322 8826 1342
rect 8774 1288 8784 1322
rect 8818 1288 8826 1322
rect 8774 1241 8826 1288
rect 8774 1207 8784 1241
rect 8818 1207 8826 1241
rect 8774 1184 8826 1207
rect 8880 1324 8932 1342
rect 8880 1290 8888 1324
rect 8922 1290 8932 1324
rect 8880 1256 8932 1290
rect 8880 1222 8888 1256
rect 8922 1222 8932 1256
rect 8880 1188 8932 1222
rect 8880 1154 8888 1188
rect 8922 1154 8932 1188
rect 8880 1142 8932 1154
rect 8962 1330 9016 1342
rect 8962 1296 8972 1330
rect 9006 1296 9016 1330
rect 8962 1262 9016 1296
rect 8962 1228 8972 1262
rect 9006 1228 9016 1262
rect 8962 1142 9016 1228
rect 9046 1308 9100 1342
rect 9046 1274 9056 1308
rect 9090 1274 9100 1308
rect 9046 1213 9100 1274
rect 9046 1179 9056 1213
rect 9090 1179 9100 1213
rect 9046 1142 9100 1179
rect 9130 1330 9184 1342
rect 9130 1296 9140 1330
rect 9174 1296 9184 1330
rect 9130 1262 9184 1296
rect 9130 1228 9140 1262
rect 9174 1228 9184 1262
rect 9130 1142 9184 1228
rect 9214 1308 9268 1342
rect 9214 1274 9224 1308
rect 9258 1274 9268 1308
rect 9214 1213 9268 1274
rect 9214 1179 9224 1213
rect 9258 1179 9268 1213
rect 9214 1142 9268 1179
rect 9298 1330 9350 1342
rect 9298 1296 9308 1330
rect 9342 1296 9350 1330
rect 9298 1262 9350 1296
rect 9298 1228 9308 1262
rect 9342 1228 9350 1262
rect 9298 1194 9350 1228
rect 9298 1160 9308 1194
rect 9342 1160 9350 1194
rect 9298 1142 9350 1160
rect 9432 1330 9484 1342
rect 9432 1296 9440 1330
rect 9474 1296 9484 1330
rect 9432 1262 9484 1296
rect 9432 1228 9440 1262
rect 9474 1228 9484 1262
rect 9432 1194 9484 1228
rect 9432 1160 9440 1194
rect 9474 1160 9484 1194
rect 9432 1142 9484 1160
rect 9514 1324 9568 1342
rect 9514 1290 9524 1324
rect 9558 1290 9568 1324
rect 9514 1256 9568 1290
rect 9514 1222 9524 1256
rect 9558 1222 9568 1256
rect 9514 1188 9568 1222
rect 9514 1154 9524 1188
rect 9558 1154 9568 1188
rect 9514 1142 9568 1154
rect 9598 1330 9652 1342
rect 9598 1296 9608 1330
rect 9642 1296 9652 1330
rect 9598 1262 9652 1296
rect 9598 1228 9608 1262
rect 9642 1228 9652 1262
rect 9598 1142 9652 1228
rect 9682 1324 9736 1342
rect 9682 1290 9692 1324
rect 9726 1290 9736 1324
rect 9682 1256 9736 1290
rect 9682 1222 9692 1256
rect 9726 1222 9736 1256
rect 9682 1188 9736 1222
rect 9682 1154 9692 1188
rect 9726 1154 9736 1188
rect 9682 1142 9736 1154
rect 9766 1330 9820 1342
rect 9766 1296 9776 1330
rect 9810 1296 9820 1330
rect 9766 1262 9820 1296
rect 9766 1228 9776 1262
rect 9810 1228 9820 1262
rect 9766 1142 9820 1228
rect 9850 1324 9904 1342
rect 9850 1290 9860 1324
rect 9894 1290 9904 1324
rect 9850 1256 9904 1290
rect 9850 1222 9860 1256
rect 9894 1222 9904 1256
rect 9850 1188 9904 1222
rect 9850 1154 9860 1188
rect 9894 1154 9904 1188
rect 9850 1142 9904 1154
rect 9934 1330 9988 1342
rect 9934 1296 9944 1330
rect 9978 1296 9988 1330
rect 9934 1262 9988 1296
rect 9934 1228 9944 1262
rect 9978 1228 9988 1262
rect 9934 1142 9988 1228
rect 10018 1324 10072 1342
rect 10018 1290 10028 1324
rect 10062 1290 10072 1324
rect 10018 1256 10072 1290
rect 10018 1222 10028 1256
rect 10062 1222 10072 1256
rect 10018 1188 10072 1222
rect 10018 1154 10028 1188
rect 10062 1154 10072 1188
rect 10018 1142 10072 1154
rect 10102 1330 10156 1342
rect 10102 1296 10112 1330
rect 10146 1296 10156 1330
rect 10102 1262 10156 1296
rect 10102 1228 10112 1262
rect 10146 1228 10156 1262
rect 10102 1142 10156 1228
rect 10186 1324 10240 1342
rect 10186 1290 10196 1324
rect 10230 1290 10240 1324
rect 10186 1256 10240 1290
rect 10186 1222 10196 1256
rect 10230 1222 10240 1256
rect 10186 1188 10240 1222
rect 10186 1154 10196 1188
rect 10230 1154 10240 1188
rect 10186 1142 10240 1154
rect 10270 1330 10324 1342
rect 10270 1296 10280 1330
rect 10314 1296 10324 1330
rect 10270 1262 10324 1296
rect 10270 1228 10280 1262
rect 10314 1228 10324 1262
rect 10270 1142 10324 1228
rect 10354 1324 10408 1342
rect 10354 1290 10364 1324
rect 10398 1290 10408 1324
rect 10354 1256 10408 1290
rect 10354 1222 10364 1256
rect 10398 1222 10408 1256
rect 10354 1188 10408 1222
rect 10354 1154 10364 1188
rect 10398 1154 10408 1188
rect 10354 1142 10408 1154
rect 10438 1330 10492 1342
rect 10438 1296 10448 1330
rect 10482 1296 10492 1330
rect 10438 1262 10492 1296
rect 10438 1228 10448 1262
rect 10482 1228 10492 1262
rect 10438 1142 10492 1228
rect 10522 1324 10576 1342
rect 10522 1290 10532 1324
rect 10566 1290 10576 1324
rect 10522 1256 10576 1290
rect 10522 1222 10532 1256
rect 10566 1222 10576 1256
rect 10522 1188 10576 1222
rect 10522 1154 10532 1188
rect 10566 1154 10576 1188
rect 10522 1142 10576 1154
rect 10606 1330 10660 1342
rect 10606 1296 10616 1330
rect 10650 1296 10660 1330
rect 10606 1262 10660 1296
rect 10606 1228 10616 1262
rect 10650 1228 10660 1262
rect 10606 1142 10660 1228
rect 10690 1324 10744 1342
rect 10690 1290 10700 1324
rect 10734 1290 10744 1324
rect 10690 1256 10744 1290
rect 10690 1222 10700 1256
rect 10734 1222 10744 1256
rect 10690 1188 10744 1222
rect 10690 1154 10700 1188
rect 10734 1154 10744 1188
rect 10690 1142 10744 1154
rect 10774 1330 10828 1342
rect 10774 1296 10784 1330
rect 10818 1296 10828 1330
rect 10774 1262 10828 1296
rect 10774 1228 10784 1262
rect 10818 1228 10828 1262
rect 10774 1142 10828 1228
rect 10858 1324 10912 1342
rect 10858 1290 10868 1324
rect 10902 1290 10912 1324
rect 10858 1256 10912 1290
rect 10858 1222 10868 1256
rect 10902 1222 10912 1256
rect 10858 1188 10912 1222
rect 10858 1154 10868 1188
rect 10902 1154 10912 1188
rect 10858 1142 10912 1154
rect 10942 1330 10996 1342
rect 10942 1296 10952 1330
rect 10986 1296 10996 1330
rect 10942 1262 10996 1296
rect 10942 1228 10952 1262
rect 10986 1228 10996 1262
rect 10942 1142 10996 1228
rect 11026 1324 11080 1342
rect 11026 1290 11036 1324
rect 11070 1290 11080 1324
rect 11026 1256 11080 1290
rect 11026 1222 11036 1256
rect 11070 1222 11080 1256
rect 11026 1188 11080 1222
rect 11026 1154 11036 1188
rect 11070 1154 11080 1188
rect 11026 1142 11080 1154
rect 11110 1330 11164 1342
rect 11110 1296 11120 1330
rect 11154 1296 11164 1330
rect 11110 1262 11164 1296
rect 11110 1228 11120 1262
rect 11154 1228 11164 1262
rect 11110 1142 11164 1228
rect 11194 1324 11248 1342
rect 11194 1290 11204 1324
rect 11238 1290 11248 1324
rect 11194 1256 11248 1290
rect 11194 1222 11204 1256
rect 11238 1222 11248 1256
rect 11194 1188 11248 1222
rect 11194 1154 11204 1188
rect 11238 1154 11248 1188
rect 11194 1142 11248 1154
rect 11278 1330 11330 1342
rect 11278 1296 11288 1330
rect 11322 1296 11330 1330
rect 11278 1262 11330 1296
rect 11278 1228 11288 1262
rect 11322 1228 11330 1262
rect 11278 1142 11330 1228
rect 12988 1322 13040 1342
rect 12988 1288 12996 1322
rect 13030 1288 13040 1322
rect 12988 1254 13040 1288
rect 12988 1220 12996 1254
rect 13030 1220 13040 1254
rect 12988 1184 13040 1220
rect 13070 1322 13128 1342
rect 13070 1288 13082 1322
rect 13116 1288 13128 1322
rect 13070 1254 13128 1288
rect 13070 1220 13082 1254
rect 13116 1220 13128 1254
rect 13070 1184 13128 1220
rect 13158 1322 13210 1342
rect 13158 1288 13168 1322
rect 13202 1288 13210 1322
rect 13158 1241 13210 1288
rect 13158 1207 13168 1241
rect 13202 1207 13210 1241
rect 13158 1184 13210 1207
rect 13264 1324 13316 1342
rect 13264 1290 13272 1324
rect 13306 1290 13316 1324
rect 13264 1256 13316 1290
rect 13264 1222 13272 1256
rect 13306 1222 13316 1256
rect 13264 1188 13316 1222
rect 13264 1154 13272 1188
rect 13306 1154 13316 1188
rect 13264 1142 13316 1154
rect 13346 1330 13400 1342
rect 13346 1296 13356 1330
rect 13390 1296 13400 1330
rect 13346 1262 13400 1296
rect 13346 1228 13356 1262
rect 13390 1228 13400 1262
rect 13346 1142 13400 1228
rect 13430 1308 13484 1342
rect 13430 1274 13440 1308
rect 13474 1274 13484 1308
rect 13430 1213 13484 1274
rect 13430 1179 13440 1213
rect 13474 1179 13484 1213
rect 13430 1142 13484 1179
rect 13514 1330 13568 1342
rect 13514 1296 13524 1330
rect 13558 1296 13568 1330
rect 13514 1262 13568 1296
rect 13514 1228 13524 1262
rect 13558 1228 13568 1262
rect 13514 1142 13568 1228
rect 13598 1308 13652 1342
rect 13598 1274 13608 1308
rect 13642 1274 13652 1308
rect 13598 1213 13652 1274
rect 13598 1179 13608 1213
rect 13642 1179 13652 1213
rect 13598 1142 13652 1179
rect 13682 1330 13734 1342
rect 13682 1296 13692 1330
rect 13726 1296 13734 1330
rect 13682 1262 13734 1296
rect 13682 1228 13692 1262
rect 13726 1228 13734 1262
rect 13682 1194 13734 1228
rect 13682 1160 13692 1194
rect 13726 1160 13734 1194
rect 13682 1142 13734 1160
rect 13816 1330 13868 1342
rect 13816 1296 13824 1330
rect 13858 1296 13868 1330
rect 13816 1262 13868 1296
rect 13816 1228 13824 1262
rect 13858 1228 13868 1262
rect 13816 1194 13868 1228
rect 13816 1160 13824 1194
rect 13858 1160 13868 1194
rect 13816 1142 13868 1160
rect 13898 1324 13952 1342
rect 13898 1290 13908 1324
rect 13942 1290 13952 1324
rect 13898 1256 13952 1290
rect 13898 1222 13908 1256
rect 13942 1222 13952 1256
rect 13898 1188 13952 1222
rect 13898 1154 13908 1188
rect 13942 1154 13952 1188
rect 13898 1142 13952 1154
rect 13982 1330 14036 1342
rect 13982 1296 13992 1330
rect 14026 1296 14036 1330
rect 13982 1262 14036 1296
rect 13982 1228 13992 1262
rect 14026 1228 14036 1262
rect 13982 1142 14036 1228
rect 14066 1324 14120 1342
rect 14066 1290 14076 1324
rect 14110 1290 14120 1324
rect 14066 1256 14120 1290
rect 14066 1222 14076 1256
rect 14110 1222 14120 1256
rect 14066 1188 14120 1222
rect 14066 1154 14076 1188
rect 14110 1154 14120 1188
rect 14066 1142 14120 1154
rect 14150 1330 14204 1342
rect 14150 1296 14160 1330
rect 14194 1296 14204 1330
rect 14150 1262 14204 1296
rect 14150 1228 14160 1262
rect 14194 1228 14204 1262
rect 14150 1142 14204 1228
rect 14234 1324 14288 1342
rect 14234 1290 14244 1324
rect 14278 1290 14288 1324
rect 14234 1256 14288 1290
rect 14234 1222 14244 1256
rect 14278 1222 14288 1256
rect 14234 1188 14288 1222
rect 14234 1154 14244 1188
rect 14278 1154 14288 1188
rect 14234 1142 14288 1154
rect 14318 1330 14372 1342
rect 14318 1296 14328 1330
rect 14362 1296 14372 1330
rect 14318 1262 14372 1296
rect 14318 1228 14328 1262
rect 14362 1228 14372 1262
rect 14318 1142 14372 1228
rect 14402 1324 14456 1342
rect 14402 1290 14412 1324
rect 14446 1290 14456 1324
rect 14402 1256 14456 1290
rect 14402 1222 14412 1256
rect 14446 1222 14456 1256
rect 14402 1188 14456 1222
rect 14402 1154 14412 1188
rect 14446 1154 14456 1188
rect 14402 1142 14456 1154
rect 14486 1330 14540 1342
rect 14486 1296 14496 1330
rect 14530 1296 14540 1330
rect 14486 1262 14540 1296
rect 14486 1228 14496 1262
rect 14530 1228 14540 1262
rect 14486 1142 14540 1228
rect 14570 1324 14624 1342
rect 14570 1290 14580 1324
rect 14614 1290 14624 1324
rect 14570 1256 14624 1290
rect 14570 1222 14580 1256
rect 14614 1222 14624 1256
rect 14570 1188 14624 1222
rect 14570 1154 14580 1188
rect 14614 1154 14624 1188
rect 14570 1142 14624 1154
rect 14654 1330 14708 1342
rect 14654 1296 14664 1330
rect 14698 1296 14708 1330
rect 14654 1262 14708 1296
rect 14654 1228 14664 1262
rect 14698 1228 14708 1262
rect 14654 1142 14708 1228
rect 14738 1324 14792 1342
rect 14738 1290 14748 1324
rect 14782 1290 14792 1324
rect 14738 1256 14792 1290
rect 14738 1222 14748 1256
rect 14782 1222 14792 1256
rect 14738 1188 14792 1222
rect 14738 1154 14748 1188
rect 14782 1154 14792 1188
rect 14738 1142 14792 1154
rect 14822 1330 14876 1342
rect 14822 1296 14832 1330
rect 14866 1296 14876 1330
rect 14822 1262 14876 1296
rect 14822 1228 14832 1262
rect 14866 1228 14876 1262
rect 14822 1142 14876 1228
rect 14906 1324 14960 1342
rect 14906 1290 14916 1324
rect 14950 1290 14960 1324
rect 14906 1256 14960 1290
rect 14906 1222 14916 1256
rect 14950 1222 14960 1256
rect 14906 1188 14960 1222
rect 14906 1154 14916 1188
rect 14950 1154 14960 1188
rect 14906 1142 14960 1154
rect 14990 1330 15044 1342
rect 14990 1296 15000 1330
rect 15034 1296 15044 1330
rect 14990 1262 15044 1296
rect 14990 1228 15000 1262
rect 15034 1228 15044 1262
rect 14990 1142 15044 1228
rect 15074 1324 15128 1342
rect 15074 1290 15084 1324
rect 15118 1290 15128 1324
rect 15074 1256 15128 1290
rect 15074 1222 15084 1256
rect 15118 1222 15128 1256
rect 15074 1188 15128 1222
rect 15074 1154 15084 1188
rect 15118 1154 15128 1188
rect 15074 1142 15128 1154
rect 15158 1330 15212 1342
rect 15158 1296 15168 1330
rect 15202 1296 15212 1330
rect 15158 1262 15212 1296
rect 15158 1228 15168 1262
rect 15202 1228 15212 1262
rect 15158 1142 15212 1228
rect 15242 1324 15296 1342
rect 15242 1290 15252 1324
rect 15286 1290 15296 1324
rect 15242 1256 15296 1290
rect 15242 1222 15252 1256
rect 15286 1222 15296 1256
rect 15242 1188 15296 1222
rect 15242 1154 15252 1188
rect 15286 1154 15296 1188
rect 15242 1142 15296 1154
rect 15326 1330 15380 1342
rect 15326 1296 15336 1330
rect 15370 1296 15380 1330
rect 15326 1262 15380 1296
rect 15326 1228 15336 1262
rect 15370 1228 15380 1262
rect 15326 1142 15380 1228
rect 15410 1324 15464 1342
rect 15410 1290 15420 1324
rect 15454 1290 15464 1324
rect 15410 1256 15464 1290
rect 15410 1222 15420 1256
rect 15454 1222 15464 1256
rect 15410 1188 15464 1222
rect 15410 1154 15420 1188
rect 15454 1154 15464 1188
rect 15410 1142 15464 1154
rect 15494 1330 15548 1342
rect 15494 1296 15504 1330
rect 15538 1296 15548 1330
rect 15494 1262 15548 1296
rect 15494 1228 15504 1262
rect 15538 1228 15548 1262
rect 15494 1142 15548 1228
rect 15578 1324 15632 1342
rect 15578 1290 15588 1324
rect 15622 1290 15632 1324
rect 15578 1256 15632 1290
rect 15578 1222 15588 1256
rect 15622 1222 15632 1256
rect 15578 1188 15632 1222
rect 15578 1154 15588 1188
rect 15622 1154 15632 1188
rect 15578 1142 15632 1154
rect 15662 1330 15714 1342
rect 15662 1296 15672 1330
rect 15706 1296 15714 1330
rect 15662 1262 15714 1296
rect 15662 1228 15672 1262
rect 15706 1228 15714 1262
rect 15662 1142 15714 1228
rect 8602 188 8654 200
rect 8602 154 8610 188
rect 8644 154 8654 188
rect 8602 120 8654 154
rect 8602 86 8610 120
rect 8644 86 8654 120
rect 8602 52 8654 86
rect 8602 18 8610 52
rect 8644 18 8654 52
rect 8602 0 8654 18
rect 8684 188 8736 200
rect 8684 154 8694 188
rect 8728 161 8736 188
rect 10676 188 10728 200
rect 10676 161 10684 188
rect 8728 154 8763 161
rect 8684 120 8763 154
rect 8684 86 8694 120
rect 8728 86 8763 120
rect 8684 77 8763 86
rect 8793 77 8866 161
rect 8896 128 9080 161
rect 8896 94 8930 128
rect 8964 94 9005 128
rect 9039 94 9080 128
rect 8896 77 9080 94
rect 9110 77 9152 161
rect 9182 128 9248 161
rect 9182 94 9202 128
rect 9236 94 9248 128
rect 9182 77 9248 94
rect 9278 128 9334 161
rect 9278 94 9288 128
rect 9322 94 9334 128
rect 9278 77 9334 94
rect 10078 128 10134 161
rect 10078 94 10090 128
rect 10124 94 10134 128
rect 10078 77 10134 94
rect 10164 128 10230 161
rect 10164 94 10176 128
rect 10210 94 10230 128
rect 10164 77 10230 94
rect 10260 77 10302 161
rect 10332 128 10516 161
rect 10332 94 10373 128
rect 10407 94 10448 128
rect 10482 94 10516 128
rect 10332 77 10516 94
rect 10546 77 10619 161
rect 10649 154 10684 161
rect 10718 154 10728 188
rect 10649 120 10728 154
rect 10649 86 10684 120
rect 10718 86 10728 120
rect 10649 77 10728 86
rect 8684 52 8736 77
rect 8684 18 8694 52
rect 8728 18 8736 52
rect 8684 0 8736 18
rect 10676 52 10728 77
rect 10676 18 10684 52
rect 10718 18 10728 52
rect 10676 0 10728 18
rect 10758 188 10810 200
rect 10758 154 10768 188
rect 10802 154 10810 188
rect 10758 120 10810 154
rect 10758 86 10768 120
rect 10802 86 10810 120
rect 10758 52 10810 86
rect 10758 18 10768 52
rect 10802 18 10810 52
rect 10758 0 10810 18
rect 10994 188 11046 200
rect 10994 154 11002 188
rect 11036 154 11046 188
rect 10994 120 11046 154
rect 10994 86 11002 120
rect 11036 86 11046 120
rect 10994 52 11046 86
rect 10994 18 11002 52
rect 11036 18 11046 52
rect 10994 0 11046 18
rect 11076 188 11128 200
rect 11076 154 11086 188
rect 11120 161 11128 188
rect 13068 188 13120 200
rect 13068 161 13076 188
rect 11120 154 11155 161
rect 11076 120 11155 154
rect 11076 86 11086 120
rect 11120 86 11155 120
rect 11076 77 11155 86
rect 11185 77 11258 161
rect 11288 128 11472 161
rect 11288 94 11322 128
rect 11356 94 11397 128
rect 11431 94 11472 128
rect 11288 77 11472 94
rect 11502 77 11544 161
rect 11574 128 11640 161
rect 11574 94 11594 128
rect 11628 94 11640 128
rect 11574 77 11640 94
rect 11670 128 11726 161
rect 11670 94 11680 128
rect 11714 94 11726 128
rect 11670 77 11726 94
rect 12470 128 12526 161
rect 12470 94 12482 128
rect 12516 94 12526 128
rect 12470 77 12526 94
rect 12556 128 12622 161
rect 12556 94 12568 128
rect 12602 94 12622 128
rect 12556 77 12622 94
rect 12652 77 12694 161
rect 12724 128 12908 161
rect 12724 94 12765 128
rect 12799 94 12840 128
rect 12874 94 12908 128
rect 12724 77 12908 94
rect 12938 77 13011 161
rect 13041 154 13076 161
rect 13110 154 13120 188
rect 13041 120 13120 154
rect 13041 86 13076 120
rect 13110 86 13120 120
rect 13041 77 13120 86
rect 11076 52 11128 77
rect 11076 18 11086 52
rect 11120 18 11128 52
rect 11076 0 11128 18
rect 13068 52 13120 77
rect 13068 18 13076 52
rect 13110 18 13120 52
rect 13068 0 13120 18
rect 13150 188 13202 200
rect 13150 154 13160 188
rect 13194 154 13202 188
rect 13150 120 13202 154
rect 13150 86 13160 120
rect 13194 86 13202 120
rect 13150 52 13202 86
rect 13150 18 13160 52
rect 13194 18 13202 52
rect 13150 0 13202 18
rect 13386 188 13438 200
rect 13386 154 13394 188
rect 13428 154 13438 188
rect 13386 120 13438 154
rect 13386 86 13394 120
rect 13428 86 13438 120
rect 13386 52 13438 86
rect 13386 18 13394 52
rect 13428 18 13438 52
rect 13386 0 13438 18
rect 13468 188 13520 200
rect 13468 154 13478 188
rect 13512 161 13520 188
rect 15458 188 15510 200
rect 15458 161 15466 188
rect 13512 154 13547 161
rect 13468 120 13547 154
rect 13468 86 13478 120
rect 13512 86 13547 120
rect 13468 77 13547 86
rect 13577 77 13650 161
rect 13680 128 13864 161
rect 13680 94 13714 128
rect 13748 94 13789 128
rect 13823 94 13864 128
rect 13680 77 13864 94
rect 13894 77 13936 161
rect 13966 128 14032 161
rect 13966 94 13986 128
rect 14020 94 14032 128
rect 13966 77 14032 94
rect 14062 128 14118 161
rect 14062 94 14072 128
rect 14106 94 14118 128
rect 14062 77 14118 94
rect 14860 128 14916 161
rect 14860 94 14872 128
rect 14906 94 14916 128
rect 14860 77 14916 94
rect 14946 128 15012 161
rect 14946 94 14958 128
rect 14992 94 15012 128
rect 14946 77 15012 94
rect 15042 77 15084 161
rect 15114 128 15298 161
rect 15114 94 15155 128
rect 15189 94 15230 128
rect 15264 94 15298 128
rect 15114 77 15298 94
rect 15328 77 15401 161
rect 15431 154 15466 161
rect 15500 154 15510 188
rect 15431 120 15510 154
rect 15431 86 15466 120
rect 15500 86 15510 120
rect 15431 77 15510 86
rect 13468 52 13520 77
rect 13468 18 13478 52
rect 13512 18 13520 52
rect 13468 0 13520 18
rect 15458 52 15510 77
rect 15458 18 15466 52
rect 15500 18 15510 52
rect 15458 0 15510 18
rect 15540 188 15592 200
rect 15540 154 15550 188
rect 15584 154 15592 188
rect 15540 120 15592 154
rect 15540 86 15550 120
rect 15584 86 15592 120
rect 15540 52 15592 86
rect 15540 18 15550 52
rect 15584 18 15592 52
rect 15540 0 15592 18
rect 15778 188 15830 200
rect 15778 154 15786 188
rect 15820 154 15830 188
rect 15778 120 15830 154
rect 15778 86 15786 120
rect 15820 86 15830 120
rect 15778 52 15830 86
rect 15778 18 15786 52
rect 15820 18 15830 52
rect 15778 0 15830 18
rect 15860 188 15912 200
rect 15860 154 15870 188
rect 15904 161 15912 188
rect 17852 188 17904 200
rect 17852 161 17860 188
rect 15904 154 15939 161
rect 15860 120 15939 154
rect 15860 86 15870 120
rect 15904 86 15939 120
rect 15860 77 15939 86
rect 15969 77 16042 161
rect 16072 128 16256 161
rect 16072 94 16106 128
rect 16140 94 16181 128
rect 16215 94 16256 128
rect 16072 77 16256 94
rect 16286 77 16328 161
rect 16358 128 16424 161
rect 16358 94 16378 128
rect 16412 94 16424 128
rect 16358 77 16424 94
rect 16454 128 16510 161
rect 16454 94 16464 128
rect 16498 94 16510 128
rect 16454 77 16510 94
rect 17254 128 17310 161
rect 17254 94 17266 128
rect 17300 94 17310 128
rect 17254 77 17310 94
rect 17340 128 17406 161
rect 17340 94 17352 128
rect 17386 94 17406 128
rect 17340 77 17406 94
rect 17436 77 17478 161
rect 17508 128 17692 161
rect 17508 94 17549 128
rect 17583 94 17624 128
rect 17658 94 17692 128
rect 17508 77 17692 94
rect 17722 77 17795 161
rect 17825 154 17860 161
rect 17894 154 17904 188
rect 17825 120 17904 154
rect 17825 86 17860 120
rect 17894 86 17904 120
rect 17825 77 17904 86
rect 15860 52 15912 77
rect 15860 18 15870 52
rect 15904 18 15912 52
rect 15860 0 15912 18
rect 17852 52 17904 77
rect 17852 18 17860 52
rect 17894 18 17904 52
rect 17852 0 17904 18
rect 17934 188 17986 200
rect 17934 154 17944 188
rect 17978 154 17986 188
rect 17934 120 17986 154
rect 17934 86 17944 120
rect 17978 86 17986 120
rect 17934 52 17986 86
rect 17934 18 17944 52
rect 17978 18 17986 52
rect 17934 0 17986 18
rect 18170 188 18222 200
rect 18170 154 18178 188
rect 18212 154 18222 188
rect 18170 120 18222 154
rect 18170 86 18178 120
rect 18212 86 18222 120
rect 18170 52 18222 86
rect 18170 18 18178 52
rect 18212 18 18222 52
rect 18170 0 18222 18
rect 18252 188 18304 200
rect 18252 154 18262 188
rect 18296 161 18304 188
rect 20244 188 20296 200
rect 20244 161 20252 188
rect 18296 154 18331 161
rect 18252 120 18331 154
rect 18252 86 18262 120
rect 18296 86 18331 120
rect 18252 77 18331 86
rect 18361 77 18434 161
rect 18464 128 18648 161
rect 18464 94 18498 128
rect 18532 94 18573 128
rect 18607 94 18648 128
rect 18464 77 18648 94
rect 18678 77 18720 161
rect 18750 128 18816 161
rect 18750 94 18770 128
rect 18804 94 18816 128
rect 18750 77 18816 94
rect 18846 128 18902 161
rect 18846 94 18856 128
rect 18890 94 18902 128
rect 18846 77 18902 94
rect 19646 128 19702 161
rect 19646 94 19658 128
rect 19692 94 19702 128
rect 19646 77 19702 94
rect 19732 128 19798 161
rect 19732 94 19744 128
rect 19778 94 19798 128
rect 19732 77 19798 94
rect 19828 77 19870 161
rect 19900 128 20084 161
rect 19900 94 19941 128
rect 19975 94 20016 128
rect 20050 94 20084 128
rect 19900 77 20084 94
rect 20114 77 20187 161
rect 20217 154 20252 161
rect 20286 154 20296 188
rect 20217 120 20296 154
rect 20217 86 20252 120
rect 20286 86 20296 120
rect 20217 77 20296 86
rect 18252 52 18304 77
rect 18252 18 18262 52
rect 18296 18 18304 52
rect 18252 0 18304 18
rect 20244 52 20296 77
rect 20244 18 20252 52
rect 20286 18 20296 52
rect 20244 0 20296 18
rect 20326 188 20378 200
rect 20326 154 20336 188
rect 20370 154 20378 188
rect 20326 120 20378 154
rect 20326 86 20336 120
rect 20370 86 20378 120
rect 20326 52 20378 86
rect 20326 18 20336 52
rect 20370 18 20378 52
rect 20326 0 20378 18
rect 20562 188 20614 200
rect 20562 154 20570 188
rect 20604 154 20614 188
rect 20562 120 20614 154
rect 20562 86 20570 120
rect 20604 86 20614 120
rect 20562 52 20614 86
rect 20562 18 20570 52
rect 20604 18 20614 52
rect 20562 0 20614 18
rect 20644 188 20696 200
rect 20644 154 20654 188
rect 20688 161 20696 188
rect 22634 188 22686 200
rect 22634 161 22642 188
rect 20688 154 20723 161
rect 20644 120 20723 154
rect 20644 86 20654 120
rect 20688 86 20723 120
rect 20644 77 20723 86
rect 20753 77 20826 161
rect 20856 128 21040 161
rect 20856 94 20890 128
rect 20924 94 20965 128
rect 20999 94 21040 128
rect 20856 77 21040 94
rect 21070 77 21112 161
rect 21142 128 21208 161
rect 21142 94 21162 128
rect 21196 94 21208 128
rect 21142 77 21208 94
rect 21238 128 21294 161
rect 21238 94 21248 128
rect 21282 94 21294 128
rect 21238 77 21294 94
rect 22036 128 22092 161
rect 22036 94 22048 128
rect 22082 94 22092 128
rect 22036 77 22092 94
rect 22122 128 22188 161
rect 22122 94 22134 128
rect 22168 94 22188 128
rect 22122 77 22188 94
rect 22218 77 22260 161
rect 22290 128 22474 161
rect 22290 94 22331 128
rect 22365 94 22406 128
rect 22440 94 22474 128
rect 22290 77 22474 94
rect 22504 77 22577 161
rect 22607 154 22642 161
rect 22676 154 22686 188
rect 22607 120 22686 154
rect 22607 86 22642 120
rect 22676 86 22686 120
rect 22607 77 22686 86
rect 20644 52 20696 77
rect 20644 18 20654 52
rect 20688 18 20696 52
rect 20644 0 20696 18
rect 22634 52 22686 77
rect 22634 18 22642 52
rect 22676 18 22686 52
rect 22634 0 22686 18
rect 22716 188 22768 200
rect 22716 154 22726 188
rect 22760 154 22768 188
rect 22716 120 22768 154
rect 22716 86 22726 120
rect 22760 86 22768 120
rect 22716 52 22768 86
rect 22716 18 22726 52
rect 22760 18 22768 52
rect 22716 0 22768 18
rect 22954 188 23006 200
rect 22954 154 22962 188
rect 22996 154 23006 188
rect 22954 120 23006 154
rect 22954 86 22962 120
rect 22996 86 23006 120
rect 22954 52 23006 86
rect 22954 18 22962 52
rect 22996 18 23006 52
rect 22954 0 23006 18
rect 23036 188 23088 200
rect 23036 154 23046 188
rect 23080 161 23088 188
rect 25028 188 25080 200
rect 25028 161 25036 188
rect 23080 154 23115 161
rect 23036 120 23115 154
rect 23036 86 23046 120
rect 23080 86 23115 120
rect 23036 77 23115 86
rect 23145 77 23218 161
rect 23248 128 23432 161
rect 23248 94 23282 128
rect 23316 94 23357 128
rect 23391 94 23432 128
rect 23248 77 23432 94
rect 23462 77 23504 161
rect 23534 128 23600 161
rect 23534 94 23554 128
rect 23588 94 23600 128
rect 23534 77 23600 94
rect 23630 128 23686 161
rect 23630 94 23640 128
rect 23674 94 23686 128
rect 23630 77 23686 94
rect 24430 128 24486 161
rect 24430 94 24442 128
rect 24476 94 24486 128
rect 24430 77 24486 94
rect 24516 128 24582 161
rect 24516 94 24528 128
rect 24562 94 24582 128
rect 24516 77 24582 94
rect 24612 77 24654 161
rect 24684 128 24868 161
rect 24684 94 24725 128
rect 24759 94 24800 128
rect 24834 94 24868 128
rect 24684 77 24868 94
rect 24898 77 24971 161
rect 25001 154 25036 161
rect 25070 154 25080 188
rect 25001 120 25080 154
rect 25001 86 25036 120
rect 25070 86 25080 120
rect 25001 77 25080 86
rect 23036 52 23088 77
rect 23036 18 23046 52
rect 23080 18 23088 52
rect 23036 0 23088 18
rect 25028 52 25080 77
rect 25028 18 25036 52
rect 25070 18 25080 52
rect 25028 0 25080 18
rect 25110 188 25162 200
rect 25110 154 25120 188
rect 25154 154 25162 188
rect 25110 120 25162 154
rect 25110 86 25120 120
rect 25154 86 25162 120
rect 25110 52 25162 86
rect 25110 18 25120 52
rect 25154 18 25162 52
rect 25110 0 25162 18
rect 8602 -508 8654 -494
rect 8602 -542 8610 -508
rect 8644 -542 8654 -508
rect 8602 -576 8654 -542
rect 8602 -610 8610 -576
rect 8644 -610 8654 -576
rect 8602 -622 8654 -610
rect 8684 -524 8738 -494
rect 8684 -558 8694 -524
rect 8728 -558 8738 -524
rect 8684 -622 8738 -558
rect 8768 -508 8820 -494
rect 8768 -542 8778 -508
rect 8812 -542 8820 -508
rect 8768 -576 8820 -542
rect 8874 -524 8926 -488
rect 8874 -558 8882 -524
rect 8916 -558 8926 -524
rect 8874 -572 8926 -558
rect 8956 -508 9018 -488
rect 8956 -542 8966 -508
rect 9000 -542 9018 -508
rect 8956 -572 9018 -542
rect 9048 -501 9102 -488
rect 9048 -535 9058 -501
rect 9092 -535 9102 -501
rect 9048 -572 9102 -535
rect 9132 -572 9222 -488
rect 9252 -510 9328 -488
rect 9252 -544 9272 -510
rect 9306 -544 9328 -510
rect 9252 -572 9328 -544
rect 9358 -526 9436 -488
rect 9358 -560 9392 -526
rect 9426 -560 9436 -526
rect 9358 -572 9436 -560
rect 8768 -610 8778 -576
rect 8812 -610 8820 -576
rect 8768 -622 8820 -610
rect 9374 -594 9436 -572
rect 9374 -628 9392 -594
rect 9426 -628 9436 -594
rect 9374 -656 9436 -628
rect 9466 -656 9520 -488
rect 9550 -500 9657 -488
rect 9550 -534 9566 -500
rect 9600 -534 9657 -500
rect 9550 -568 9657 -534
rect 9550 -602 9566 -568
rect 9600 -602 9657 -568
rect 9550 -656 9657 -602
rect 9687 -572 9801 -488
rect 9831 -501 9885 -488
rect 9831 -535 9841 -501
rect 9875 -535 9885 -501
rect 9831 -572 9885 -535
rect 9915 -572 9990 -488
rect 10020 -500 10111 -488
rect 10020 -534 10055 -500
rect 10089 -534 10111 -500
rect 10020 -572 10111 -534
rect 10141 -526 10217 -488
rect 10141 -560 10163 -526
rect 10197 -560 10217 -526
rect 10141 -572 10217 -560
rect 9687 -656 9739 -572
rect 10167 -656 10217 -572
rect 10247 -656 10289 -488
rect 10319 -500 10371 -488
rect 10319 -534 10329 -500
rect 10363 -534 10371 -500
rect 10319 -656 10371 -534
rect 10523 -500 10575 -488
rect 10523 -534 10531 -500
rect 10565 -534 10575 -500
rect 10523 -556 10575 -534
rect 10425 -636 10478 -556
rect 10425 -670 10433 -636
rect 10467 -670 10478 -636
rect 10425 -684 10478 -670
rect 10508 -684 10575 -556
rect 10525 -688 10575 -684
rect 10605 -537 10657 -488
rect 10808 -504 10858 -488
rect 10605 -571 10615 -537
rect 10649 -571 10657 -537
rect 10605 -605 10657 -571
rect 10605 -639 10615 -605
rect 10649 -639 10657 -605
rect 10711 -518 10763 -504
rect 10711 -552 10719 -518
rect 10753 -552 10763 -518
rect 10711 -586 10763 -552
rect 10711 -620 10719 -586
rect 10753 -620 10763 -586
rect 10711 -632 10763 -620
rect 10793 -512 10858 -504
rect 10793 -546 10814 -512
rect 10848 -546 10858 -512
rect 10793 -580 10858 -546
rect 10793 -614 10814 -580
rect 10848 -614 10858 -580
rect 10793 -632 10858 -614
rect 10605 -688 10657 -639
rect 10808 -688 10858 -632
rect 10888 -536 10940 -488
rect 10888 -570 10898 -536
rect 10932 -570 10940 -536
rect 10888 -604 10940 -570
rect 10888 -638 10898 -604
rect 10932 -638 10940 -604
rect 10994 -508 11046 -494
rect 10994 -542 11002 -508
rect 11036 -542 11046 -508
rect 10994 -576 11046 -542
rect 10994 -610 11002 -576
rect 11036 -610 11046 -576
rect 10994 -622 11046 -610
rect 11076 -524 11130 -494
rect 11076 -558 11086 -524
rect 11120 -558 11130 -524
rect 11076 -622 11130 -558
rect 11160 -508 11212 -494
rect 11160 -542 11170 -508
rect 11204 -542 11212 -508
rect 11160 -576 11212 -542
rect 11266 -524 11318 -488
rect 11266 -558 11274 -524
rect 11308 -558 11318 -524
rect 11266 -572 11318 -558
rect 11348 -508 11410 -488
rect 11348 -542 11358 -508
rect 11392 -542 11410 -508
rect 11348 -572 11410 -542
rect 11440 -501 11494 -488
rect 11440 -535 11450 -501
rect 11484 -535 11494 -501
rect 11440 -572 11494 -535
rect 11524 -572 11614 -488
rect 11644 -510 11720 -488
rect 11644 -544 11664 -510
rect 11698 -544 11720 -510
rect 11644 -572 11720 -544
rect 11750 -526 11828 -488
rect 11750 -560 11784 -526
rect 11818 -560 11828 -526
rect 11750 -572 11828 -560
rect 11160 -610 11170 -576
rect 11204 -610 11212 -576
rect 11160 -622 11212 -610
rect 10888 -688 10940 -638
rect 11766 -594 11828 -572
rect 11766 -628 11784 -594
rect 11818 -628 11828 -594
rect 11766 -656 11828 -628
rect 11858 -656 11912 -488
rect 11942 -500 12049 -488
rect 11942 -534 11958 -500
rect 11992 -534 12049 -500
rect 11942 -568 12049 -534
rect 11942 -602 11958 -568
rect 11992 -602 12049 -568
rect 11942 -656 12049 -602
rect 12079 -572 12193 -488
rect 12223 -501 12277 -488
rect 12223 -535 12233 -501
rect 12267 -535 12277 -501
rect 12223 -572 12277 -535
rect 12307 -572 12382 -488
rect 12412 -500 12503 -488
rect 12412 -534 12447 -500
rect 12481 -534 12503 -500
rect 12412 -572 12503 -534
rect 12533 -526 12609 -488
rect 12533 -560 12555 -526
rect 12589 -560 12609 -526
rect 12533 -572 12609 -560
rect 12079 -656 12131 -572
rect 12559 -656 12609 -572
rect 12639 -656 12681 -488
rect 12711 -500 12763 -488
rect 12711 -534 12721 -500
rect 12755 -534 12763 -500
rect 12711 -656 12763 -534
rect 12915 -500 12967 -488
rect 12915 -534 12923 -500
rect 12957 -534 12967 -500
rect 12915 -556 12967 -534
rect 12817 -636 12870 -556
rect 12817 -670 12825 -636
rect 12859 -670 12870 -636
rect 12817 -684 12870 -670
rect 12900 -684 12967 -556
rect 12917 -688 12967 -684
rect 12997 -537 13049 -488
rect 13200 -504 13250 -488
rect 12997 -571 13007 -537
rect 13041 -571 13049 -537
rect 12997 -605 13049 -571
rect 12997 -639 13007 -605
rect 13041 -639 13049 -605
rect 13103 -518 13155 -504
rect 13103 -552 13111 -518
rect 13145 -552 13155 -518
rect 13103 -586 13155 -552
rect 13103 -620 13111 -586
rect 13145 -620 13155 -586
rect 13103 -632 13155 -620
rect 13185 -512 13250 -504
rect 13185 -546 13206 -512
rect 13240 -546 13250 -512
rect 13185 -580 13250 -546
rect 13185 -614 13206 -580
rect 13240 -614 13250 -580
rect 13185 -632 13250 -614
rect 12997 -688 13049 -639
rect 13200 -688 13250 -632
rect 13280 -536 13332 -488
rect 13280 -570 13290 -536
rect 13324 -570 13332 -536
rect 13280 -604 13332 -570
rect 13280 -638 13290 -604
rect 13324 -638 13332 -604
rect 13386 -508 13438 -494
rect 13386 -542 13394 -508
rect 13428 -542 13438 -508
rect 13386 -576 13438 -542
rect 13386 -610 13394 -576
rect 13428 -610 13438 -576
rect 13386 -622 13438 -610
rect 13468 -524 13522 -494
rect 13468 -558 13478 -524
rect 13512 -558 13522 -524
rect 13468 -622 13522 -558
rect 13552 -508 13604 -494
rect 13552 -542 13562 -508
rect 13596 -542 13604 -508
rect 13552 -576 13604 -542
rect 13658 -524 13710 -488
rect 13658 -558 13666 -524
rect 13700 -558 13710 -524
rect 13658 -572 13710 -558
rect 13740 -508 13802 -488
rect 13740 -542 13750 -508
rect 13784 -542 13802 -508
rect 13740 -572 13802 -542
rect 13832 -501 13886 -488
rect 13832 -535 13842 -501
rect 13876 -535 13886 -501
rect 13832 -572 13886 -535
rect 13916 -572 14006 -488
rect 14036 -510 14112 -488
rect 14036 -544 14056 -510
rect 14090 -544 14112 -510
rect 14036 -572 14112 -544
rect 14142 -526 14220 -488
rect 14142 -560 14176 -526
rect 14210 -560 14220 -526
rect 14142 -572 14220 -560
rect 13552 -610 13562 -576
rect 13596 -610 13604 -576
rect 13552 -622 13604 -610
rect 13280 -688 13332 -638
rect 14158 -594 14220 -572
rect 14158 -628 14176 -594
rect 14210 -628 14220 -594
rect 14158 -656 14220 -628
rect 14250 -656 14304 -488
rect 14334 -500 14441 -488
rect 14334 -534 14350 -500
rect 14384 -534 14441 -500
rect 14334 -568 14441 -534
rect 14334 -602 14350 -568
rect 14384 -602 14441 -568
rect 14334 -656 14441 -602
rect 14471 -572 14585 -488
rect 14615 -501 14669 -488
rect 14615 -535 14625 -501
rect 14659 -535 14669 -501
rect 14615 -572 14669 -535
rect 14699 -572 14774 -488
rect 14804 -500 14895 -488
rect 14804 -534 14839 -500
rect 14873 -534 14895 -500
rect 14804 -572 14895 -534
rect 14925 -526 15001 -488
rect 14925 -560 14947 -526
rect 14981 -560 15001 -526
rect 14925 -572 15001 -560
rect 14471 -656 14523 -572
rect 14951 -656 15001 -572
rect 15031 -656 15073 -488
rect 15103 -500 15155 -488
rect 15103 -534 15113 -500
rect 15147 -534 15155 -500
rect 15103 -656 15155 -534
rect 15307 -500 15359 -488
rect 15307 -534 15315 -500
rect 15349 -534 15359 -500
rect 15307 -556 15359 -534
rect 15209 -636 15262 -556
rect 15209 -670 15217 -636
rect 15251 -670 15262 -636
rect 15209 -684 15262 -670
rect 15292 -684 15359 -556
rect 15309 -688 15359 -684
rect 15389 -537 15441 -488
rect 15592 -504 15642 -488
rect 15389 -571 15399 -537
rect 15433 -571 15441 -537
rect 15389 -605 15441 -571
rect 15389 -639 15399 -605
rect 15433 -639 15441 -605
rect 15495 -518 15547 -504
rect 15495 -552 15503 -518
rect 15537 -552 15547 -518
rect 15495 -586 15547 -552
rect 15495 -620 15503 -586
rect 15537 -620 15547 -586
rect 15495 -632 15547 -620
rect 15577 -512 15642 -504
rect 15577 -546 15598 -512
rect 15632 -546 15642 -512
rect 15577 -580 15642 -546
rect 15577 -614 15598 -580
rect 15632 -614 15642 -580
rect 15577 -632 15642 -614
rect 15389 -688 15441 -639
rect 15592 -688 15642 -632
rect 15672 -536 15724 -488
rect 15672 -570 15682 -536
rect 15716 -570 15724 -536
rect 15672 -604 15724 -570
rect 15672 -638 15682 -604
rect 15716 -638 15724 -604
rect 15778 -508 15830 -494
rect 15778 -542 15786 -508
rect 15820 -542 15830 -508
rect 15778 -576 15830 -542
rect 15778 -610 15786 -576
rect 15820 -610 15830 -576
rect 15778 -622 15830 -610
rect 15860 -524 15914 -494
rect 15860 -558 15870 -524
rect 15904 -558 15914 -524
rect 15860 -622 15914 -558
rect 15944 -508 15996 -494
rect 15944 -542 15954 -508
rect 15988 -542 15996 -508
rect 15944 -576 15996 -542
rect 16050 -524 16102 -488
rect 16050 -558 16058 -524
rect 16092 -558 16102 -524
rect 16050 -572 16102 -558
rect 16132 -508 16194 -488
rect 16132 -542 16142 -508
rect 16176 -542 16194 -508
rect 16132 -572 16194 -542
rect 16224 -501 16278 -488
rect 16224 -535 16234 -501
rect 16268 -535 16278 -501
rect 16224 -572 16278 -535
rect 16308 -572 16398 -488
rect 16428 -510 16504 -488
rect 16428 -544 16448 -510
rect 16482 -544 16504 -510
rect 16428 -572 16504 -544
rect 16534 -526 16612 -488
rect 16534 -560 16568 -526
rect 16602 -560 16612 -526
rect 16534 -572 16612 -560
rect 15944 -610 15954 -576
rect 15988 -610 15996 -576
rect 15944 -622 15996 -610
rect 15672 -688 15724 -638
rect 16550 -594 16612 -572
rect 16550 -628 16568 -594
rect 16602 -628 16612 -594
rect 16550 -656 16612 -628
rect 16642 -656 16696 -488
rect 16726 -500 16833 -488
rect 16726 -534 16742 -500
rect 16776 -534 16833 -500
rect 16726 -568 16833 -534
rect 16726 -602 16742 -568
rect 16776 -602 16833 -568
rect 16726 -656 16833 -602
rect 16863 -572 16977 -488
rect 17007 -501 17061 -488
rect 17007 -535 17017 -501
rect 17051 -535 17061 -501
rect 17007 -572 17061 -535
rect 17091 -572 17166 -488
rect 17196 -500 17287 -488
rect 17196 -534 17231 -500
rect 17265 -534 17287 -500
rect 17196 -572 17287 -534
rect 17317 -526 17393 -488
rect 17317 -560 17339 -526
rect 17373 -560 17393 -526
rect 17317 -572 17393 -560
rect 16863 -656 16915 -572
rect 17343 -656 17393 -572
rect 17423 -656 17465 -488
rect 17495 -500 17547 -488
rect 17495 -534 17505 -500
rect 17539 -534 17547 -500
rect 17495 -656 17547 -534
rect 17699 -500 17751 -488
rect 17699 -534 17707 -500
rect 17741 -534 17751 -500
rect 17699 -556 17751 -534
rect 17601 -636 17654 -556
rect 17601 -670 17609 -636
rect 17643 -670 17654 -636
rect 17601 -684 17654 -670
rect 17684 -684 17751 -556
rect 17701 -688 17751 -684
rect 17781 -537 17833 -488
rect 17984 -504 18034 -488
rect 17781 -571 17791 -537
rect 17825 -571 17833 -537
rect 17781 -605 17833 -571
rect 17781 -639 17791 -605
rect 17825 -639 17833 -605
rect 17887 -518 17939 -504
rect 17887 -552 17895 -518
rect 17929 -552 17939 -518
rect 17887 -586 17939 -552
rect 17887 -620 17895 -586
rect 17929 -620 17939 -586
rect 17887 -632 17939 -620
rect 17969 -512 18034 -504
rect 17969 -546 17990 -512
rect 18024 -546 18034 -512
rect 17969 -580 18034 -546
rect 17969 -614 17990 -580
rect 18024 -614 18034 -580
rect 17969 -632 18034 -614
rect 17781 -688 17833 -639
rect 17984 -688 18034 -632
rect 18064 -536 18116 -488
rect 18064 -570 18074 -536
rect 18108 -570 18116 -536
rect 18064 -604 18116 -570
rect 18064 -638 18074 -604
rect 18108 -638 18116 -604
rect 18170 -508 18222 -494
rect 18170 -542 18178 -508
rect 18212 -542 18222 -508
rect 18170 -576 18222 -542
rect 18170 -610 18178 -576
rect 18212 -610 18222 -576
rect 18170 -622 18222 -610
rect 18252 -524 18306 -494
rect 18252 -558 18262 -524
rect 18296 -558 18306 -524
rect 18252 -622 18306 -558
rect 18336 -508 18388 -494
rect 18336 -542 18346 -508
rect 18380 -542 18388 -508
rect 18336 -576 18388 -542
rect 18442 -524 18494 -488
rect 18442 -558 18450 -524
rect 18484 -558 18494 -524
rect 18442 -572 18494 -558
rect 18524 -508 18586 -488
rect 18524 -542 18534 -508
rect 18568 -542 18586 -508
rect 18524 -572 18586 -542
rect 18616 -501 18670 -488
rect 18616 -535 18626 -501
rect 18660 -535 18670 -501
rect 18616 -572 18670 -535
rect 18700 -572 18790 -488
rect 18820 -510 18896 -488
rect 18820 -544 18840 -510
rect 18874 -544 18896 -510
rect 18820 -572 18896 -544
rect 18926 -526 19004 -488
rect 18926 -560 18960 -526
rect 18994 -560 19004 -526
rect 18926 -572 19004 -560
rect 18336 -610 18346 -576
rect 18380 -610 18388 -576
rect 18336 -622 18388 -610
rect 18064 -688 18116 -638
rect 18942 -594 19004 -572
rect 18942 -628 18960 -594
rect 18994 -628 19004 -594
rect 18942 -656 19004 -628
rect 19034 -656 19088 -488
rect 19118 -500 19225 -488
rect 19118 -534 19134 -500
rect 19168 -534 19225 -500
rect 19118 -568 19225 -534
rect 19118 -602 19134 -568
rect 19168 -602 19225 -568
rect 19118 -656 19225 -602
rect 19255 -572 19369 -488
rect 19399 -501 19453 -488
rect 19399 -535 19409 -501
rect 19443 -535 19453 -501
rect 19399 -572 19453 -535
rect 19483 -572 19558 -488
rect 19588 -500 19679 -488
rect 19588 -534 19623 -500
rect 19657 -534 19679 -500
rect 19588 -572 19679 -534
rect 19709 -526 19785 -488
rect 19709 -560 19731 -526
rect 19765 -560 19785 -526
rect 19709 -572 19785 -560
rect 19255 -656 19307 -572
rect 19735 -656 19785 -572
rect 19815 -656 19857 -488
rect 19887 -500 19939 -488
rect 19887 -534 19897 -500
rect 19931 -534 19939 -500
rect 19887 -656 19939 -534
rect 20091 -500 20143 -488
rect 20091 -534 20099 -500
rect 20133 -534 20143 -500
rect 20091 -556 20143 -534
rect 19993 -636 20046 -556
rect 19993 -670 20001 -636
rect 20035 -670 20046 -636
rect 19993 -684 20046 -670
rect 20076 -684 20143 -556
rect 20093 -688 20143 -684
rect 20173 -537 20225 -488
rect 20376 -504 20426 -488
rect 20173 -571 20183 -537
rect 20217 -571 20225 -537
rect 20173 -605 20225 -571
rect 20173 -639 20183 -605
rect 20217 -639 20225 -605
rect 20279 -518 20331 -504
rect 20279 -552 20287 -518
rect 20321 -552 20331 -518
rect 20279 -586 20331 -552
rect 20279 -620 20287 -586
rect 20321 -620 20331 -586
rect 20279 -632 20331 -620
rect 20361 -512 20426 -504
rect 20361 -546 20382 -512
rect 20416 -546 20426 -512
rect 20361 -580 20426 -546
rect 20361 -614 20382 -580
rect 20416 -614 20426 -580
rect 20361 -632 20426 -614
rect 20173 -688 20225 -639
rect 20376 -688 20426 -632
rect 20456 -536 20508 -488
rect 20456 -570 20466 -536
rect 20500 -570 20508 -536
rect 20456 -604 20508 -570
rect 20456 -638 20466 -604
rect 20500 -638 20508 -604
rect 20562 -508 20614 -494
rect 20562 -542 20570 -508
rect 20604 -542 20614 -508
rect 20562 -576 20614 -542
rect 20562 -610 20570 -576
rect 20604 -610 20614 -576
rect 20562 -622 20614 -610
rect 20644 -524 20698 -494
rect 20644 -558 20654 -524
rect 20688 -558 20698 -524
rect 20644 -622 20698 -558
rect 20728 -508 20780 -494
rect 20728 -542 20738 -508
rect 20772 -542 20780 -508
rect 20728 -576 20780 -542
rect 20834 -524 20886 -488
rect 20834 -558 20842 -524
rect 20876 -558 20886 -524
rect 20834 -572 20886 -558
rect 20916 -508 20978 -488
rect 20916 -542 20926 -508
rect 20960 -542 20978 -508
rect 20916 -572 20978 -542
rect 21008 -501 21062 -488
rect 21008 -535 21018 -501
rect 21052 -535 21062 -501
rect 21008 -572 21062 -535
rect 21092 -572 21182 -488
rect 21212 -510 21288 -488
rect 21212 -544 21232 -510
rect 21266 -544 21288 -510
rect 21212 -572 21288 -544
rect 21318 -526 21396 -488
rect 21318 -560 21352 -526
rect 21386 -560 21396 -526
rect 21318 -572 21396 -560
rect 20728 -610 20738 -576
rect 20772 -610 20780 -576
rect 20728 -622 20780 -610
rect 20456 -688 20508 -638
rect 21334 -594 21396 -572
rect 21334 -628 21352 -594
rect 21386 -628 21396 -594
rect 21334 -656 21396 -628
rect 21426 -656 21480 -488
rect 21510 -500 21617 -488
rect 21510 -534 21526 -500
rect 21560 -534 21617 -500
rect 21510 -568 21617 -534
rect 21510 -602 21526 -568
rect 21560 -602 21617 -568
rect 21510 -656 21617 -602
rect 21647 -572 21761 -488
rect 21791 -501 21845 -488
rect 21791 -535 21801 -501
rect 21835 -535 21845 -501
rect 21791 -572 21845 -535
rect 21875 -572 21950 -488
rect 21980 -500 22071 -488
rect 21980 -534 22015 -500
rect 22049 -534 22071 -500
rect 21980 -572 22071 -534
rect 22101 -526 22177 -488
rect 22101 -560 22123 -526
rect 22157 -560 22177 -526
rect 22101 -572 22177 -560
rect 21647 -656 21699 -572
rect 22127 -656 22177 -572
rect 22207 -656 22249 -488
rect 22279 -500 22331 -488
rect 22279 -534 22289 -500
rect 22323 -534 22331 -500
rect 22279 -656 22331 -534
rect 22483 -500 22535 -488
rect 22483 -534 22491 -500
rect 22525 -534 22535 -500
rect 22483 -556 22535 -534
rect 22385 -636 22438 -556
rect 22385 -670 22393 -636
rect 22427 -670 22438 -636
rect 22385 -684 22438 -670
rect 22468 -684 22535 -556
rect 22485 -688 22535 -684
rect 22565 -537 22617 -488
rect 22768 -504 22818 -488
rect 22565 -571 22575 -537
rect 22609 -571 22617 -537
rect 22565 -605 22617 -571
rect 22565 -639 22575 -605
rect 22609 -639 22617 -605
rect 22671 -518 22723 -504
rect 22671 -552 22679 -518
rect 22713 -552 22723 -518
rect 22671 -586 22723 -552
rect 22671 -620 22679 -586
rect 22713 -620 22723 -586
rect 22671 -632 22723 -620
rect 22753 -512 22818 -504
rect 22753 -546 22774 -512
rect 22808 -546 22818 -512
rect 22753 -580 22818 -546
rect 22753 -614 22774 -580
rect 22808 -614 22818 -580
rect 22753 -632 22818 -614
rect 22565 -688 22617 -639
rect 22768 -688 22818 -632
rect 22848 -536 22900 -488
rect 22848 -570 22858 -536
rect 22892 -570 22900 -536
rect 22848 -604 22900 -570
rect 22848 -638 22858 -604
rect 22892 -638 22900 -604
rect 22954 -508 23006 -494
rect 22954 -542 22962 -508
rect 22996 -542 23006 -508
rect 22954 -576 23006 -542
rect 22954 -610 22962 -576
rect 22996 -610 23006 -576
rect 22954 -622 23006 -610
rect 23036 -524 23090 -494
rect 23036 -558 23046 -524
rect 23080 -558 23090 -524
rect 23036 -622 23090 -558
rect 23120 -508 23172 -494
rect 23120 -542 23130 -508
rect 23164 -542 23172 -508
rect 23120 -576 23172 -542
rect 23226 -524 23278 -488
rect 23226 -558 23234 -524
rect 23268 -558 23278 -524
rect 23226 -572 23278 -558
rect 23308 -508 23370 -488
rect 23308 -542 23318 -508
rect 23352 -542 23370 -508
rect 23308 -572 23370 -542
rect 23400 -501 23454 -488
rect 23400 -535 23410 -501
rect 23444 -535 23454 -501
rect 23400 -572 23454 -535
rect 23484 -572 23574 -488
rect 23604 -510 23680 -488
rect 23604 -544 23624 -510
rect 23658 -544 23680 -510
rect 23604 -572 23680 -544
rect 23710 -526 23788 -488
rect 23710 -560 23744 -526
rect 23778 -560 23788 -526
rect 23710 -572 23788 -560
rect 23120 -610 23130 -576
rect 23164 -610 23172 -576
rect 23120 -622 23172 -610
rect 22848 -688 22900 -638
rect 23726 -594 23788 -572
rect 23726 -628 23744 -594
rect 23778 -628 23788 -594
rect 23726 -656 23788 -628
rect 23818 -656 23872 -488
rect 23902 -500 24009 -488
rect 23902 -534 23918 -500
rect 23952 -534 24009 -500
rect 23902 -568 24009 -534
rect 23902 -602 23918 -568
rect 23952 -602 24009 -568
rect 23902 -656 24009 -602
rect 24039 -572 24153 -488
rect 24183 -501 24237 -488
rect 24183 -535 24193 -501
rect 24227 -535 24237 -501
rect 24183 -572 24237 -535
rect 24267 -572 24342 -488
rect 24372 -500 24463 -488
rect 24372 -534 24407 -500
rect 24441 -534 24463 -500
rect 24372 -572 24463 -534
rect 24493 -526 24569 -488
rect 24493 -560 24515 -526
rect 24549 -560 24569 -526
rect 24493 -572 24569 -560
rect 24039 -656 24091 -572
rect 24519 -656 24569 -572
rect 24599 -656 24641 -488
rect 24671 -500 24723 -488
rect 24671 -534 24681 -500
rect 24715 -534 24723 -500
rect 24671 -656 24723 -534
rect 24875 -500 24927 -488
rect 24875 -534 24883 -500
rect 24917 -534 24927 -500
rect 24875 -556 24927 -534
rect 24777 -636 24830 -556
rect 24777 -670 24785 -636
rect 24819 -670 24830 -636
rect 24777 -684 24830 -670
rect 24860 -684 24927 -556
rect 24877 -688 24927 -684
rect 24957 -537 25009 -488
rect 25160 -504 25210 -488
rect 24957 -571 24967 -537
rect 25001 -571 25009 -537
rect 24957 -605 25009 -571
rect 24957 -639 24967 -605
rect 25001 -639 25009 -605
rect 25063 -518 25115 -504
rect 25063 -552 25071 -518
rect 25105 -552 25115 -518
rect 25063 -586 25115 -552
rect 25063 -620 25071 -586
rect 25105 -620 25115 -586
rect 25063 -632 25115 -620
rect 25145 -512 25210 -504
rect 25145 -546 25166 -512
rect 25200 -546 25210 -512
rect 25145 -580 25210 -546
rect 25145 -614 25166 -580
rect 25200 -614 25210 -580
rect 25145 -632 25210 -614
rect 24957 -688 25009 -639
rect 25160 -688 25210 -632
rect 25240 -536 25292 -488
rect 25240 -570 25250 -536
rect 25284 -570 25292 -536
rect 25240 -604 25292 -570
rect 25240 -638 25250 -604
rect 25284 -638 25292 -604
rect 25240 -688 25292 -638
rect 8602 -1225 8654 -1177
rect 8602 -1259 8610 -1225
rect 8644 -1259 8654 -1225
rect 8602 -1293 8654 -1259
rect 8602 -1327 8610 -1293
rect 8644 -1327 8654 -1293
rect 8602 -1377 8654 -1327
rect 8684 -1193 8734 -1177
rect 8684 -1201 8749 -1193
rect 8684 -1235 8694 -1201
rect 8728 -1235 8749 -1201
rect 8684 -1269 8749 -1235
rect 8684 -1303 8694 -1269
rect 8728 -1303 8749 -1269
rect 8684 -1321 8749 -1303
rect 8779 -1207 8831 -1193
rect 8779 -1241 8789 -1207
rect 8823 -1241 8831 -1207
rect 8779 -1275 8831 -1241
rect 8779 -1309 8789 -1275
rect 8823 -1309 8831 -1275
rect 8779 -1321 8831 -1309
rect 8885 -1226 8937 -1177
rect 8885 -1260 8893 -1226
rect 8927 -1260 8937 -1226
rect 8885 -1294 8937 -1260
rect 8684 -1377 8734 -1321
rect 8885 -1328 8893 -1294
rect 8927 -1328 8937 -1294
rect 8885 -1377 8937 -1328
rect 8967 -1189 9019 -1177
rect 8967 -1223 8977 -1189
rect 9011 -1223 9019 -1189
rect 9171 -1189 9223 -1177
rect 8967 -1245 9019 -1223
rect 9171 -1223 9179 -1189
rect 9213 -1223 9223 -1189
rect 8967 -1373 9034 -1245
rect 9064 -1325 9117 -1245
rect 9064 -1359 9075 -1325
rect 9109 -1359 9117 -1325
rect 9171 -1345 9223 -1223
rect 9253 -1345 9295 -1177
rect 9325 -1215 9401 -1177
rect 9325 -1249 9345 -1215
rect 9379 -1249 9401 -1215
rect 9325 -1261 9401 -1249
rect 9431 -1189 9522 -1177
rect 9431 -1223 9453 -1189
rect 9487 -1223 9522 -1189
rect 9431 -1261 9522 -1223
rect 9552 -1261 9627 -1177
rect 9657 -1190 9711 -1177
rect 9657 -1224 9667 -1190
rect 9701 -1224 9711 -1190
rect 9657 -1261 9711 -1224
rect 9741 -1261 9855 -1177
rect 9325 -1345 9375 -1261
rect 9064 -1373 9117 -1359
rect 8967 -1377 9017 -1373
rect 9803 -1345 9855 -1261
rect 9885 -1189 9992 -1177
rect 9885 -1223 9942 -1189
rect 9976 -1223 9992 -1189
rect 9885 -1257 9992 -1223
rect 9885 -1291 9942 -1257
rect 9976 -1291 9992 -1257
rect 9885 -1345 9992 -1291
rect 10022 -1345 10076 -1177
rect 10106 -1215 10184 -1177
rect 10106 -1249 10116 -1215
rect 10150 -1249 10184 -1215
rect 10106 -1261 10184 -1249
rect 10214 -1199 10290 -1177
rect 10214 -1233 10236 -1199
rect 10270 -1233 10290 -1199
rect 10214 -1261 10290 -1233
rect 10320 -1261 10410 -1177
rect 10440 -1190 10494 -1177
rect 10440 -1224 10450 -1190
rect 10484 -1224 10494 -1190
rect 10440 -1261 10494 -1224
rect 10524 -1197 10586 -1177
rect 10524 -1231 10542 -1197
rect 10576 -1231 10586 -1197
rect 10524 -1261 10586 -1231
rect 10616 -1213 10668 -1177
rect 10616 -1247 10626 -1213
rect 10660 -1247 10668 -1213
rect 10616 -1261 10668 -1247
rect 10722 -1197 10774 -1183
rect 10722 -1231 10730 -1197
rect 10764 -1231 10774 -1197
rect 10106 -1283 10168 -1261
rect 10106 -1317 10116 -1283
rect 10150 -1317 10168 -1283
rect 10106 -1345 10168 -1317
rect 10722 -1265 10774 -1231
rect 10722 -1299 10730 -1265
rect 10764 -1299 10774 -1265
rect 10722 -1311 10774 -1299
rect 10804 -1213 10858 -1183
rect 10804 -1247 10814 -1213
rect 10848 -1247 10858 -1213
rect 10804 -1311 10858 -1247
rect 10888 -1197 10940 -1183
rect 10888 -1231 10898 -1197
rect 10932 -1231 10940 -1197
rect 10888 -1265 10940 -1231
rect 10888 -1299 10898 -1265
rect 10932 -1299 10940 -1265
rect 10888 -1311 10940 -1299
rect 10994 -1225 11046 -1177
rect 10994 -1259 11002 -1225
rect 11036 -1259 11046 -1225
rect 10994 -1293 11046 -1259
rect 10994 -1327 11002 -1293
rect 11036 -1327 11046 -1293
rect 10994 -1377 11046 -1327
rect 11076 -1193 11126 -1177
rect 11076 -1201 11141 -1193
rect 11076 -1235 11086 -1201
rect 11120 -1235 11141 -1201
rect 11076 -1269 11141 -1235
rect 11076 -1303 11086 -1269
rect 11120 -1303 11141 -1269
rect 11076 -1321 11141 -1303
rect 11171 -1207 11223 -1193
rect 11171 -1241 11181 -1207
rect 11215 -1241 11223 -1207
rect 11171 -1275 11223 -1241
rect 11171 -1309 11181 -1275
rect 11215 -1309 11223 -1275
rect 11171 -1321 11223 -1309
rect 11277 -1226 11329 -1177
rect 11277 -1260 11285 -1226
rect 11319 -1260 11329 -1226
rect 11277 -1294 11329 -1260
rect 11076 -1377 11126 -1321
rect 11277 -1328 11285 -1294
rect 11319 -1328 11329 -1294
rect 11277 -1377 11329 -1328
rect 11359 -1189 11411 -1177
rect 11359 -1223 11369 -1189
rect 11403 -1223 11411 -1189
rect 11563 -1189 11615 -1177
rect 11359 -1245 11411 -1223
rect 11563 -1223 11571 -1189
rect 11605 -1223 11615 -1189
rect 11359 -1373 11426 -1245
rect 11456 -1325 11509 -1245
rect 11456 -1359 11467 -1325
rect 11501 -1359 11509 -1325
rect 11563 -1345 11615 -1223
rect 11645 -1345 11687 -1177
rect 11717 -1215 11793 -1177
rect 11717 -1249 11737 -1215
rect 11771 -1249 11793 -1215
rect 11717 -1261 11793 -1249
rect 11823 -1189 11914 -1177
rect 11823 -1223 11845 -1189
rect 11879 -1223 11914 -1189
rect 11823 -1261 11914 -1223
rect 11944 -1261 12019 -1177
rect 12049 -1190 12103 -1177
rect 12049 -1224 12059 -1190
rect 12093 -1224 12103 -1190
rect 12049 -1261 12103 -1224
rect 12133 -1261 12247 -1177
rect 11717 -1345 11767 -1261
rect 11456 -1373 11509 -1359
rect 11359 -1377 11409 -1373
rect 12195 -1345 12247 -1261
rect 12277 -1189 12384 -1177
rect 12277 -1223 12334 -1189
rect 12368 -1223 12384 -1189
rect 12277 -1257 12384 -1223
rect 12277 -1291 12334 -1257
rect 12368 -1291 12384 -1257
rect 12277 -1345 12384 -1291
rect 12414 -1345 12468 -1177
rect 12498 -1215 12576 -1177
rect 12498 -1249 12508 -1215
rect 12542 -1249 12576 -1215
rect 12498 -1261 12576 -1249
rect 12606 -1199 12682 -1177
rect 12606 -1233 12628 -1199
rect 12662 -1233 12682 -1199
rect 12606 -1261 12682 -1233
rect 12712 -1261 12802 -1177
rect 12832 -1190 12886 -1177
rect 12832 -1224 12842 -1190
rect 12876 -1224 12886 -1190
rect 12832 -1261 12886 -1224
rect 12916 -1197 12978 -1177
rect 12916 -1231 12934 -1197
rect 12968 -1231 12978 -1197
rect 12916 -1261 12978 -1231
rect 13008 -1213 13060 -1177
rect 13008 -1247 13018 -1213
rect 13052 -1247 13060 -1213
rect 13008 -1261 13060 -1247
rect 13114 -1197 13166 -1183
rect 13114 -1231 13122 -1197
rect 13156 -1231 13166 -1197
rect 12498 -1283 12560 -1261
rect 12498 -1317 12508 -1283
rect 12542 -1317 12560 -1283
rect 12498 -1345 12560 -1317
rect 13114 -1265 13166 -1231
rect 13114 -1299 13122 -1265
rect 13156 -1299 13166 -1265
rect 13114 -1311 13166 -1299
rect 13196 -1213 13250 -1183
rect 13196 -1247 13206 -1213
rect 13240 -1247 13250 -1213
rect 13196 -1311 13250 -1247
rect 13280 -1197 13332 -1183
rect 13280 -1231 13290 -1197
rect 13324 -1231 13332 -1197
rect 13280 -1265 13332 -1231
rect 13280 -1299 13290 -1265
rect 13324 -1299 13332 -1265
rect 13280 -1311 13332 -1299
rect 13386 -1225 13438 -1177
rect 13386 -1259 13394 -1225
rect 13428 -1259 13438 -1225
rect 13386 -1293 13438 -1259
rect 13386 -1327 13394 -1293
rect 13428 -1327 13438 -1293
rect 13386 -1377 13438 -1327
rect 13468 -1193 13518 -1177
rect 13468 -1201 13533 -1193
rect 13468 -1235 13478 -1201
rect 13512 -1235 13533 -1201
rect 13468 -1269 13533 -1235
rect 13468 -1303 13478 -1269
rect 13512 -1303 13533 -1269
rect 13468 -1321 13533 -1303
rect 13563 -1207 13615 -1193
rect 13563 -1241 13573 -1207
rect 13607 -1241 13615 -1207
rect 13563 -1275 13615 -1241
rect 13563 -1309 13573 -1275
rect 13607 -1309 13615 -1275
rect 13563 -1321 13615 -1309
rect 13669 -1226 13721 -1177
rect 13669 -1260 13677 -1226
rect 13711 -1260 13721 -1226
rect 13669 -1294 13721 -1260
rect 13468 -1377 13518 -1321
rect 13669 -1328 13677 -1294
rect 13711 -1328 13721 -1294
rect 13669 -1377 13721 -1328
rect 13751 -1189 13803 -1177
rect 13751 -1223 13761 -1189
rect 13795 -1223 13803 -1189
rect 13955 -1189 14007 -1177
rect 13751 -1245 13803 -1223
rect 13955 -1223 13963 -1189
rect 13997 -1223 14007 -1189
rect 13751 -1373 13818 -1245
rect 13848 -1325 13901 -1245
rect 13848 -1359 13859 -1325
rect 13893 -1359 13901 -1325
rect 13955 -1345 14007 -1223
rect 14037 -1345 14079 -1177
rect 14109 -1215 14185 -1177
rect 14109 -1249 14129 -1215
rect 14163 -1249 14185 -1215
rect 14109 -1261 14185 -1249
rect 14215 -1189 14306 -1177
rect 14215 -1223 14237 -1189
rect 14271 -1223 14306 -1189
rect 14215 -1261 14306 -1223
rect 14336 -1261 14411 -1177
rect 14441 -1190 14495 -1177
rect 14441 -1224 14451 -1190
rect 14485 -1224 14495 -1190
rect 14441 -1261 14495 -1224
rect 14525 -1261 14639 -1177
rect 14109 -1345 14159 -1261
rect 13848 -1373 13901 -1359
rect 13751 -1377 13801 -1373
rect 14587 -1345 14639 -1261
rect 14669 -1189 14776 -1177
rect 14669 -1223 14726 -1189
rect 14760 -1223 14776 -1189
rect 14669 -1257 14776 -1223
rect 14669 -1291 14726 -1257
rect 14760 -1291 14776 -1257
rect 14669 -1345 14776 -1291
rect 14806 -1345 14860 -1177
rect 14890 -1215 14968 -1177
rect 14890 -1249 14900 -1215
rect 14934 -1249 14968 -1215
rect 14890 -1261 14968 -1249
rect 14998 -1199 15074 -1177
rect 14998 -1233 15020 -1199
rect 15054 -1233 15074 -1199
rect 14998 -1261 15074 -1233
rect 15104 -1261 15194 -1177
rect 15224 -1190 15278 -1177
rect 15224 -1224 15234 -1190
rect 15268 -1224 15278 -1190
rect 15224 -1261 15278 -1224
rect 15308 -1197 15370 -1177
rect 15308 -1231 15326 -1197
rect 15360 -1231 15370 -1197
rect 15308 -1261 15370 -1231
rect 15400 -1213 15452 -1177
rect 15400 -1247 15410 -1213
rect 15444 -1247 15452 -1213
rect 15400 -1261 15452 -1247
rect 15506 -1197 15558 -1183
rect 15506 -1231 15514 -1197
rect 15548 -1231 15558 -1197
rect 14890 -1283 14952 -1261
rect 14890 -1317 14900 -1283
rect 14934 -1317 14952 -1283
rect 14890 -1345 14952 -1317
rect 15506 -1265 15558 -1231
rect 15506 -1299 15514 -1265
rect 15548 -1299 15558 -1265
rect 15506 -1311 15558 -1299
rect 15588 -1213 15642 -1183
rect 15588 -1247 15598 -1213
rect 15632 -1247 15642 -1213
rect 15588 -1311 15642 -1247
rect 15672 -1197 15724 -1183
rect 15672 -1231 15682 -1197
rect 15716 -1231 15724 -1197
rect 15672 -1265 15724 -1231
rect 15672 -1299 15682 -1265
rect 15716 -1299 15724 -1265
rect 15672 -1311 15724 -1299
rect 15778 -1225 15830 -1177
rect 15778 -1259 15786 -1225
rect 15820 -1259 15830 -1225
rect 15778 -1293 15830 -1259
rect 15778 -1327 15786 -1293
rect 15820 -1327 15830 -1293
rect 15778 -1377 15830 -1327
rect 15860 -1193 15910 -1177
rect 15860 -1201 15925 -1193
rect 15860 -1235 15870 -1201
rect 15904 -1235 15925 -1201
rect 15860 -1269 15925 -1235
rect 15860 -1303 15870 -1269
rect 15904 -1303 15925 -1269
rect 15860 -1321 15925 -1303
rect 15955 -1207 16007 -1193
rect 15955 -1241 15965 -1207
rect 15999 -1241 16007 -1207
rect 15955 -1275 16007 -1241
rect 15955 -1309 15965 -1275
rect 15999 -1309 16007 -1275
rect 15955 -1321 16007 -1309
rect 16061 -1226 16113 -1177
rect 16061 -1260 16069 -1226
rect 16103 -1260 16113 -1226
rect 16061 -1294 16113 -1260
rect 15860 -1377 15910 -1321
rect 16061 -1328 16069 -1294
rect 16103 -1328 16113 -1294
rect 16061 -1377 16113 -1328
rect 16143 -1189 16195 -1177
rect 16143 -1223 16153 -1189
rect 16187 -1223 16195 -1189
rect 16347 -1189 16399 -1177
rect 16143 -1245 16195 -1223
rect 16347 -1223 16355 -1189
rect 16389 -1223 16399 -1189
rect 16143 -1373 16210 -1245
rect 16240 -1325 16293 -1245
rect 16240 -1359 16251 -1325
rect 16285 -1359 16293 -1325
rect 16347 -1345 16399 -1223
rect 16429 -1345 16471 -1177
rect 16501 -1215 16577 -1177
rect 16501 -1249 16521 -1215
rect 16555 -1249 16577 -1215
rect 16501 -1261 16577 -1249
rect 16607 -1189 16698 -1177
rect 16607 -1223 16629 -1189
rect 16663 -1223 16698 -1189
rect 16607 -1261 16698 -1223
rect 16728 -1261 16803 -1177
rect 16833 -1190 16887 -1177
rect 16833 -1224 16843 -1190
rect 16877 -1224 16887 -1190
rect 16833 -1261 16887 -1224
rect 16917 -1261 17031 -1177
rect 16501 -1345 16551 -1261
rect 16240 -1373 16293 -1359
rect 16143 -1377 16193 -1373
rect 16979 -1345 17031 -1261
rect 17061 -1189 17168 -1177
rect 17061 -1223 17118 -1189
rect 17152 -1223 17168 -1189
rect 17061 -1257 17168 -1223
rect 17061 -1291 17118 -1257
rect 17152 -1291 17168 -1257
rect 17061 -1345 17168 -1291
rect 17198 -1345 17252 -1177
rect 17282 -1215 17360 -1177
rect 17282 -1249 17292 -1215
rect 17326 -1249 17360 -1215
rect 17282 -1261 17360 -1249
rect 17390 -1199 17466 -1177
rect 17390 -1233 17412 -1199
rect 17446 -1233 17466 -1199
rect 17390 -1261 17466 -1233
rect 17496 -1261 17586 -1177
rect 17616 -1190 17670 -1177
rect 17616 -1224 17626 -1190
rect 17660 -1224 17670 -1190
rect 17616 -1261 17670 -1224
rect 17700 -1197 17762 -1177
rect 17700 -1231 17718 -1197
rect 17752 -1231 17762 -1197
rect 17700 -1261 17762 -1231
rect 17792 -1213 17844 -1177
rect 17792 -1247 17802 -1213
rect 17836 -1247 17844 -1213
rect 17792 -1261 17844 -1247
rect 17898 -1197 17950 -1183
rect 17898 -1231 17906 -1197
rect 17940 -1231 17950 -1197
rect 17282 -1283 17344 -1261
rect 17282 -1317 17292 -1283
rect 17326 -1317 17344 -1283
rect 17282 -1345 17344 -1317
rect 17898 -1265 17950 -1231
rect 17898 -1299 17906 -1265
rect 17940 -1299 17950 -1265
rect 17898 -1311 17950 -1299
rect 17980 -1213 18034 -1183
rect 17980 -1247 17990 -1213
rect 18024 -1247 18034 -1213
rect 17980 -1311 18034 -1247
rect 18064 -1197 18116 -1183
rect 18064 -1231 18074 -1197
rect 18108 -1231 18116 -1197
rect 18064 -1265 18116 -1231
rect 18064 -1299 18074 -1265
rect 18108 -1299 18116 -1265
rect 18064 -1311 18116 -1299
rect 18170 -1225 18222 -1177
rect 18170 -1259 18178 -1225
rect 18212 -1259 18222 -1225
rect 18170 -1293 18222 -1259
rect 18170 -1327 18178 -1293
rect 18212 -1327 18222 -1293
rect 18170 -1377 18222 -1327
rect 18252 -1193 18302 -1177
rect 18252 -1201 18317 -1193
rect 18252 -1235 18262 -1201
rect 18296 -1235 18317 -1201
rect 18252 -1269 18317 -1235
rect 18252 -1303 18262 -1269
rect 18296 -1303 18317 -1269
rect 18252 -1321 18317 -1303
rect 18347 -1207 18399 -1193
rect 18347 -1241 18357 -1207
rect 18391 -1241 18399 -1207
rect 18347 -1275 18399 -1241
rect 18347 -1309 18357 -1275
rect 18391 -1309 18399 -1275
rect 18347 -1321 18399 -1309
rect 18453 -1226 18505 -1177
rect 18453 -1260 18461 -1226
rect 18495 -1260 18505 -1226
rect 18453 -1294 18505 -1260
rect 18252 -1377 18302 -1321
rect 18453 -1328 18461 -1294
rect 18495 -1328 18505 -1294
rect 18453 -1377 18505 -1328
rect 18535 -1189 18587 -1177
rect 18535 -1223 18545 -1189
rect 18579 -1223 18587 -1189
rect 18739 -1189 18791 -1177
rect 18535 -1245 18587 -1223
rect 18739 -1223 18747 -1189
rect 18781 -1223 18791 -1189
rect 18535 -1373 18602 -1245
rect 18632 -1325 18685 -1245
rect 18632 -1359 18643 -1325
rect 18677 -1359 18685 -1325
rect 18739 -1345 18791 -1223
rect 18821 -1345 18863 -1177
rect 18893 -1215 18969 -1177
rect 18893 -1249 18913 -1215
rect 18947 -1249 18969 -1215
rect 18893 -1261 18969 -1249
rect 18999 -1189 19090 -1177
rect 18999 -1223 19021 -1189
rect 19055 -1223 19090 -1189
rect 18999 -1261 19090 -1223
rect 19120 -1261 19195 -1177
rect 19225 -1190 19279 -1177
rect 19225 -1224 19235 -1190
rect 19269 -1224 19279 -1190
rect 19225 -1261 19279 -1224
rect 19309 -1261 19423 -1177
rect 18893 -1345 18943 -1261
rect 18632 -1373 18685 -1359
rect 18535 -1377 18585 -1373
rect 19371 -1345 19423 -1261
rect 19453 -1189 19560 -1177
rect 19453 -1223 19510 -1189
rect 19544 -1223 19560 -1189
rect 19453 -1257 19560 -1223
rect 19453 -1291 19510 -1257
rect 19544 -1291 19560 -1257
rect 19453 -1345 19560 -1291
rect 19590 -1345 19644 -1177
rect 19674 -1215 19752 -1177
rect 19674 -1249 19684 -1215
rect 19718 -1249 19752 -1215
rect 19674 -1261 19752 -1249
rect 19782 -1199 19858 -1177
rect 19782 -1233 19804 -1199
rect 19838 -1233 19858 -1199
rect 19782 -1261 19858 -1233
rect 19888 -1261 19978 -1177
rect 20008 -1190 20062 -1177
rect 20008 -1224 20018 -1190
rect 20052 -1224 20062 -1190
rect 20008 -1261 20062 -1224
rect 20092 -1197 20154 -1177
rect 20092 -1231 20110 -1197
rect 20144 -1231 20154 -1197
rect 20092 -1261 20154 -1231
rect 20184 -1213 20236 -1177
rect 20184 -1247 20194 -1213
rect 20228 -1247 20236 -1213
rect 20184 -1261 20236 -1247
rect 20290 -1197 20342 -1183
rect 20290 -1231 20298 -1197
rect 20332 -1231 20342 -1197
rect 19674 -1283 19736 -1261
rect 19674 -1317 19684 -1283
rect 19718 -1317 19736 -1283
rect 19674 -1345 19736 -1317
rect 20290 -1265 20342 -1231
rect 20290 -1299 20298 -1265
rect 20332 -1299 20342 -1265
rect 20290 -1311 20342 -1299
rect 20372 -1213 20426 -1183
rect 20372 -1247 20382 -1213
rect 20416 -1247 20426 -1213
rect 20372 -1311 20426 -1247
rect 20456 -1197 20508 -1183
rect 20456 -1231 20466 -1197
rect 20500 -1231 20508 -1197
rect 20456 -1265 20508 -1231
rect 20456 -1299 20466 -1265
rect 20500 -1299 20508 -1265
rect 20456 -1311 20508 -1299
rect 20562 -1225 20614 -1177
rect 20562 -1259 20570 -1225
rect 20604 -1259 20614 -1225
rect 20562 -1293 20614 -1259
rect 20562 -1327 20570 -1293
rect 20604 -1327 20614 -1293
rect 20562 -1377 20614 -1327
rect 20644 -1193 20694 -1177
rect 20644 -1201 20709 -1193
rect 20644 -1235 20654 -1201
rect 20688 -1235 20709 -1201
rect 20644 -1269 20709 -1235
rect 20644 -1303 20654 -1269
rect 20688 -1303 20709 -1269
rect 20644 -1321 20709 -1303
rect 20739 -1207 20791 -1193
rect 20739 -1241 20749 -1207
rect 20783 -1241 20791 -1207
rect 20739 -1275 20791 -1241
rect 20739 -1309 20749 -1275
rect 20783 -1309 20791 -1275
rect 20739 -1321 20791 -1309
rect 20845 -1226 20897 -1177
rect 20845 -1260 20853 -1226
rect 20887 -1260 20897 -1226
rect 20845 -1294 20897 -1260
rect 20644 -1377 20694 -1321
rect 20845 -1328 20853 -1294
rect 20887 -1328 20897 -1294
rect 20845 -1377 20897 -1328
rect 20927 -1189 20979 -1177
rect 20927 -1223 20937 -1189
rect 20971 -1223 20979 -1189
rect 21131 -1189 21183 -1177
rect 20927 -1245 20979 -1223
rect 21131 -1223 21139 -1189
rect 21173 -1223 21183 -1189
rect 20927 -1373 20994 -1245
rect 21024 -1325 21077 -1245
rect 21024 -1359 21035 -1325
rect 21069 -1359 21077 -1325
rect 21131 -1345 21183 -1223
rect 21213 -1345 21255 -1177
rect 21285 -1215 21361 -1177
rect 21285 -1249 21305 -1215
rect 21339 -1249 21361 -1215
rect 21285 -1261 21361 -1249
rect 21391 -1189 21482 -1177
rect 21391 -1223 21413 -1189
rect 21447 -1223 21482 -1189
rect 21391 -1261 21482 -1223
rect 21512 -1261 21587 -1177
rect 21617 -1190 21671 -1177
rect 21617 -1224 21627 -1190
rect 21661 -1224 21671 -1190
rect 21617 -1261 21671 -1224
rect 21701 -1261 21815 -1177
rect 21285 -1345 21335 -1261
rect 21024 -1373 21077 -1359
rect 20927 -1377 20977 -1373
rect 21763 -1345 21815 -1261
rect 21845 -1189 21952 -1177
rect 21845 -1223 21902 -1189
rect 21936 -1223 21952 -1189
rect 21845 -1257 21952 -1223
rect 21845 -1291 21902 -1257
rect 21936 -1291 21952 -1257
rect 21845 -1345 21952 -1291
rect 21982 -1345 22036 -1177
rect 22066 -1215 22144 -1177
rect 22066 -1249 22076 -1215
rect 22110 -1249 22144 -1215
rect 22066 -1261 22144 -1249
rect 22174 -1199 22250 -1177
rect 22174 -1233 22196 -1199
rect 22230 -1233 22250 -1199
rect 22174 -1261 22250 -1233
rect 22280 -1261 22370 -1177
rect 22400 -1190 22454 -1177
rect 22400 -1224 22410 -1190
rect 22444 -1224 22454 -1190
rect 22400 -1261 22454 -1224
rect 22484 -1197 22546 -1177
rect 22484 -1231 22502 -1197
rect 22536 -1231 22546 -1197
rect 22484 -1261 22546 -1231
rect 22576 -1213 22628 -1177
rect 22576 -1247 22586 -1213
rect 22620 -1247 22628 -1213
rect 22576 -1261 22628 -1247
rect 22682 -1197 22734 -1183
rect 22682 -1231 22690 -1197
rect 22724 -1231 22734 -1197
rect 22066 -1283 22128 -1261
rect 22066 -1317 22076 -1283
rect 22110 -1317 22128 -1283
rect 22066 -1345 22128 -1317
rect 22682 -1265 22734 -1231
rect 22682 -1299 22690 -1265
rect 22724 -1299 22734 -1265
rect 22682 -1311 22734 -1299
rect 22764 -1213 22818 -1183
rect 22764 -1247 22774 -1213
rect 22808 -1247 22818 -1213
rect 22764 -1311 22818 -1247
rect 22848 -1197 22900 -1183
rect 22848 -1231 22858 -1197
rect 22892 -1231 22900 -1197
rect 22848 -1265 22900 -1231
rect 22848 -1299 22858 -1265
rect 22892 -1299 22900 -1265
rect 22848 -1311 22900 -1299
rect 22954 -1225 23006 -1177
rect 22954 -1259 22962 -1225
rect 22996 -1259 23006 -1225
rect 22954 -1293 23006 -1259
rect 22954 -1327 22962 -1293
rect 22996 -1327 23006 -1293
rect 22954 -1377 23006 -1327
rect 23036 -1193 23086 -1177
rect 23036 -1201 23101 -1193
rect 23036 -1235 23046 -1201
rect 23080 -1235 23101 -1201
rect 23036 -1269 23101 -1235
rect 23036 -1303 23046 -1269
rect 23080 -1303 23101 -1269
rect 23036 -1321 23101 -1303
rect 23131 -1207 23183 -1193
rect 23131 -1241 23141 -1207
rect 23175 -1241 23183 -1207
rect 23131 -1275 23183 -1241
rect 23131 -1309 23141 -1275
rect 23175 -1309 23183 -1275
rect 23131 -1321 23183 -1309
rect 23237 -1226 23289 -1177
rect 23237 -1260 23245 -1226
rect 23279 -1260 23289 -1226
rect 23237 -1294 23289 -1260
rect 23036 -1377 23086 -1321
rect 23237 -1328 23245 -1294
rect 23279 -1328 23289 -1294
rect 23237 -1377 23289 -1328
rect 23319 -1189 23371 -1177
rect 23319 -1223 23329 -1189
rect 23363 -1223 23371 -1189
rect 23523 -1189 23575 -1177
rect 23319 -1245 23371 -1223
rect 23523 -1223 23531 -1189
rect 23565 -1223 23575 -1189
rect 23319 -1373 23386 -1245
rect 23416 -1325 23469 -1245
rect 23416 -1359 23427 -1325
rect 23461 -1359 23469 -1325
rect 23523 -1345 23575 -1223
rect 23605 -1345 23647 -1177
rect 23677 -1215 23753 -1177
rect 23677 -1249 23697 -1215
rect 23731 -1249 23753 -1215
rect 23677 -1261 23753 -1249
rect 23783 -1189 23874 -1177
rect 23783 -1223 23805 -1189
rect 23839 -1223 23874 -1189
rect 23783 -1261 23874 -1223
rect 23904 -1261 23979 -1177
rect 24009 -1190 24063 -1177
rect 24009 -1224 24019 -1190
rect 24053 -1224 24063 -1190
rect 24009 -1261 24063 -1224
rect 24093 -1261 24207 -1177
rect 23677 -1345 23727 -1261
rect 23416 -1373 23469 -1359
rect 23319 -1377 23369 -1373
rect 24155 -1345 24207 -1261
rect 24237 -1189 24344 -1177
rect 24237 -1223 24294 -1189
rect 24328 -1223 24344 -1189
rect 24237 -1257 24344 -1223
rect 24237 -1291 24294 -1257
rect 24328 -1291 24344 -1257
rect 24237 -1345 24344 -1291
rect 24374 -1345 24428 -1177
rect 24458 -1215 24536 -1177
rect 24458 -1249 24468 -1215
rect 24502 -1249 24536 -1215
rect 24458 -1261 24536 -1249
rect 24566 -1199 24642 -1177
rect 24566 -1233 24588 -1199
rect 24622 -1233 24642 -1199
rect 24566 -1261 24642 -1233
rect 24672 -1261 24762 -1177
rect 24792 -1190 24846 -1177
rect 24792 -1224 24802 -1190
rect 24836 -1224 24846 -1190
rect 24792 -1261 24846 -1224
rect 24876 -1197 24938 -1177
rect 24876 -1231 24894 -1197
rect 24928 -1231 24938 -1197
rect 24876 -1261 24938 -1231
rect 24968 -1213 25020 -1177
rect 24968 -1247 24978 -1213
rect 25012 -1247 25020 -1213
rect 24968 -1261 25020 -1247
rect 25074 -1197 25126 -1183
rect 25074 -1231 25082 -1197
rect 25116 -1231 25126 -1197
rect 24458 -1283 24520 -1261
rect 24458 -1317 24468 -1283
rect 24502 -1317 24520 -1283
rect 24458 -1345 24520 -1317
rect 25074 -1265 25126 -1231
rect 25074 -1299 25082 -1265
rect 25116 -1299 25126 -1265
rect 25074 -1311 25126 -1299
rect 25156 -1213 25210 -1183
rect 25156 -1247 25166 -1213
rect 25200 -1247 25210 -1213
rect 25156 -1311 25210 -1247
rect 25240 -1197 25292 -1183
rect 25240 -1231 25250 -1197
rect 25284 -1231 25292 -1197
rect 25240 -1265 25292 -1231
rect 25240 -1299 25250 -1265
rect 25284 -1299 25292 -1265
rect 25240 -1311 25292 -1299
<< ndiffc >>
rect 13350 12580 13384 12614
rect 13350 12512 13384 12546
rect 13434 12580 13468 12614
rect 13434 12512 13468 12546
rect 13540 12580 13574 12614
rect 13540 12512 13574 12546
rect 13624 12580 13658 12614
rect 13624 12512 13658 12546
rect 20059 12580 20093 12614
rect 20059 12512 20093 12546
rect 20143 12580 20177 12614
rect 20143 12512 20177 12546
rect 20249 12580 20283 12614
rect 20249 12512 20283 12546
rect 20333 12580 20367 12614
rect 20333 12512 20367 12546
rect 10917 12330 10951 12364
rect 11001 12356 11035 12390
rect 11085 12330 11119 12364
rect 11189 12356 11223 12390
rect 11273 12338 11307 12372
rect 11379 12356 11413 12390
rect 11596 12360 11630 12394
rect 11680 12340 11714 12374
rect 2462 12105 2496 12139
rect 2462 12037 2496 12071
rect 2546 12105 2580 12139
rect 2546 12037 2580 12071
rect 2652 12105 2686 12139
rect 2652 12037 2686 12071
rect 2736 12105 2770 12139
rect 2736 12037 2770 12071
rect 11780 12296 11814 12330
rect 11864 12322 11898 12356
rect 11968 12356 12002 12390
rect 12162 12356 12196 12390
rect 12353 12360 12387 12394
rect 12455 12340 12489 12374
rect 12555 12296 12589 12330
rect 12639 12348 12673 12382
rect 12743 12346 12777 12380
rect 12838 12356 12872 12390
rect 12922 12322 12956 12356
rect 13026 12330 13060 12364
rect 13121 12356 13155 12390
rect 13205 12320 13239 12354
rect 14811 12178 14845 12238
rect 14901 12178 14935 12238
rect 15543 12178 15577 12238
rect 15650 12178 15684 12238
rect 15753 12178 15787 12238
rect 16755 12178 16789 12238
rect 16861 12178 16895 12238
rect 16965 12178 16999 12238
rect 18093 12178 18127 12238
rect 18201 12178 18235 12238
rect 18303 12178 18337 12238
rect 18948 12178 18982 12238
rect 19037 12178 19071 12238
rect 19601 12179 19635 12239
rect 19689 12179 19723 12239
rect 19785 12179 19819 12239
rect 19881 12179 19915 12239
rect 21520 12178 21554 12238
rect 21610 12178 21644 12238
rect 22252 12178 22286 12238
rect 22359 12178 22393 12238
rect 22462 12178 22496 12238
rect 23464 12178 23498 12238
rect 23570 12178 23604 12238
rect 23674 12178 23708 12238
rect 24802 12178 24836 12238
rect 24910 12178 24944 12238
rect 25012 12178 25046 12238
rect 25657 12178 25691 12238
rect 25746 12178 25780 12238
rect 26310 12179 26344 12239
rect 26398 12179 26432 12239
rect 26494 12179 26528 12239
rect 26590 12179 26624 12239
rect 13791 11994 13825 12054
rect 13951 11994 13985 12054
rect 19601 12041 19635 12101
rect 19689 12041 19723 12101
rect 20500 11994 20534 12054
rect 20660 11994 20694 12054
rect 26310 12041 26344 12101
rect 26398 12041 26432 12101
rect 13791 11856 13825 11916
rect 13951 11856 13985 11916
rect 20500 11856 20534 11916
rect 20660 11856 20694 11916
rect 3923 11703 3957 11763
rect 4013 11703 4047 11763
rect 4655 11703 4689 11763
rect 4762 11703 4796 11763
rect 4865 11703 4899 11763
rect 5867 11703 5901 11763
rect 5973 11703 6007 11763
rect 6077 11703 6111 11763
rect 7205 11703 7239 11763
rect 7313 11703 7347 11763
rect 7415 11703 7449 11763
rect 8060 11703 8094 11763
rect 8149 11703 8183 11763
rect 8713 11704 8747 11764
rect 8801 11704 8835 11764
rect 8897 11704 8931 11764
rect 8993 11704 9027 11764
rect 9137 11728 9171 11762
rect 9137 11660 9171 11694
rect 9221 11728 9255 11762
rect 9221 11660 9255 11694
rect 2903 11519 2937 11579
rect 3063 11519 3097 11579
rect 8713 11566 8747 11626
rect 8801 11566 8835 11626
rect 13791 11718 13825 11778
rect 13951 11718 13985 11778
rect 20500 11718 20534 11778
rect 20660 11718 20694 11778
rect 13791 11580 13825 11640
rect 13951 11580 13985 11640
rect 20500 11580 20534 11640
rect 20660 11580 20694 11640
rect 2903 11381 2937 11441
rect 13791 11442 13825 11502
rect 3063 11381 3097 11441
rect 10958 11396 10992 11430
rect 10958 11328 10992 11362
rect 2903 11243 2937 11303
rect 11042 11396 11076 11430
rect 11042 11328 11076 11362
rect 11234 11396 11268 11430
rect 11234 11328 11268 11362
rect 13951 11442 13985 11502
rect 20500 11442 20534 11502
rect 20660 11442 20694 11502
rect 11318 11396 11352 11430
rect 11318 11328 11352 11362
rect 3063 11243 3097 11303
rect 13791 11304 13825 11364
rect 13951 11304 13985 11364
rect 20500 11304 20534 11364
rect 20660 11304 20694 11364
rect 2903 11105 2937 11165
rect 3063 11105 3097 11165
rect 13791 11166 13825 11226
rect 13951 11166 13985 11226
rect 20500 11166 20534 11226
rect 20660 11166 20694 11226
rect 2903 10967 2937 11027
rect 3063 10967 3097 11027
rect 13791 11028 13825 11088
rect 13951 11028 13985 11088
rect 20500 11028 20534 11088
rect 20660 11028 20694 11088
rect 2903 10829 2937 10889
rect 3063 10829 3097 10889
rect 2903 10691 2937 10751
rect 3063 10691 3097 10751
rect 2903 10553 2937 10613
rect 3063 10553 3097 10613
rect 2903 10033 2937 10093
rect 3063 10033 3097 10093
rect 19194 10021 19228 10081
rect 19354 10021 19388 10081
rect 25903 10021 25937 10081
rect 26063 10021 26097 10081
rect 2903 9895 2937 9955
rect 3063 9895 3097 9955
rect 19194 9883 19228 9943
rect 19354 9883 19388 9943
rect 2903 9757 2937 9817
rect 25903 9883 25937 9943
rect 26063 9883 26097 9943
rect 3063 9757 3097 9817
rect 19194 9745 19228 9805
rect 19354 9745 19388 9805
rect 25903 9745 25937 9805
rect 26063 9745 26097 9805
rect 2903 9619 2937 9679
rect 3063 9619 3097 9679
rect 19194 9607 19228 9667
rect 19354 9607 19388 9667
rect 25903 9607 25937 9667
rect 26063 9607 26097 9667
rect 2903 9481 2937 9541
rect 3063 9481 3097 9541
rect 19194 9469 19228 9529
rect 19354 9469 19388 9529
rect 25903 9469 25937 9529
rect 26063 9469 26097 9529
rect 2903 9343 2937 9403
rect 3063 9343 3097 9403
rect 19194 9331 19228 9391
rect 19354 9331 19388 9391
rect 25903 9331 25937 9391
rect 26063 9331 26097 9391
rect 2903 9205 2937 9265
rect 3063 9205 3097 9265
rect 19194 9193 19228 9253
rect 19354 9193 19388 9253
rect 25903 9193 25937 9253
rect 26063 9193 26097 9253
rect 2903 9067 2937 9127
rect 3063 9067 3097 9127
rect 8713 9020 8747 9080
rect 8801 9020 8835 9080
rect 3923 8883 3957 8943
rect 4013 8883 4047 8943
rect 4655 8883 4689 8943
rect 4762 8883 4796 8943
rect 4865 8883 4899 8943
rect 5867 8883 5901 8943
rect 5973 8883 6007 8943
rect 6077 8883 6111 8943
rect 7205 8883 7239 8943
rect 7313 8883 7347 8943
rect 7415 8883 7449 8943
rect 8060 8883 8094 8943
rect 9137 8954 9171 8988
rect 8149 8883 8183 8943
rect 8713 8882 8747 8942
rect 8801 8882 8835 8942
rect 8897 8882 8931 8942
rect 8993 8882 9027 8942
rect 9137 8886 9171 8920
rect 9221 8954 9255 8988
rect 9221 8886 9255 8920
rect 9352 8922 9386 8956
rect 9436 8958 9470 8992
rect 9531 8932 9565 8966
rect 9635 8924 9669 8958
rect 9719 8958 9753 8992
rect 9814 8948 9848 8982
rect 9918 8950 9952 8984
rect 10002 8898 10036 8932
rect 10102 8942 10136 8976
rect 10204 8962 10238 8996
rect 10395 8958 10429 8992
rect 2462 8575 2496 8609
rect 2462 8507 2496 8541
rect 2546 8575 2580 8609
rect 2546 8507 2580 8541
rect 2652 8575 2686 8609
rect 2652 8507 2686 8541
rect 2736 8575 2770 8609
rect 2736 8507 2770 8541
rect 10589 8958 10623 8992
rect 10693 8924 10727 8958
rect 10777 8898 10811 8932
rect 10877 8942 10911 8976
rect 10961 8962 10995 8996
rect 11178 8958 11212 8992
rect 11284 8940 11318 8974
rect 11368 8958 11402 8992
rect 11472 8932 11506 8966
rect 11556 8958 11590 8992
rect 13456 9008 13490 9068
rect 13544 9008 13578 9068
rect 19194 9055 19228 9115
rect 19354 9055 19388 9115
rect 11640 8932 11674 8966
rect 11833 8884 11867 8944
rect 11929 8884 11963 8944
rect 12025 8884 12059 8944
rect 12121 8884 12155 8944
rect 12233 8872 12267 8932
rect 12684 8945 12718 8979
rect 12321 8872 12355 8932
rect 12434 8871 12468 8931
rect 12522 8871 12556 8931
rect 12684 8877 12718 8911
rect 12852 8945 12886 8979
rect 12852 8877 12886 8911
rect 13007 8941 13041 8975
rect 13007 8873 13041 8907
rect 13091 8941 13125 8975
rect 20165 9008 20199 9068
rect 20253 9008 20287 9068
rect 25903 9055 25937 9115
rect 26063 9055 26097 9115
rect 13091 8873 13125 8907
rect 13264 8870 13298 8930
rect 13360 8870 13394 8930
rect 13456 8870 13490 8930
rect 13544 8870 13578 8930
rect 14108 8871 14142 8931
rect 14197 8871 14231 8931
rect 14842 8871 14876 8931
rect 14944 8871 14978 8931
rect 15052 8871 15086 8931
rect 16180 8871 16214 8931
rect 16284 8871 16318 8931
rect 16390 8871 16424 8931
rect 17392 8871 17426 8931
rect 17495 8871 17529 8931
rect 17602 8871 17636 8931
rect 18244 8871 18278 8931
rect 18334 8871 18368 8931
rect 19973 8870 20007 8930
rect 20069 8870 20103 8930
rect 20165 8870 20199 8930
rect 20253 8870 20287 8930
rect 20817 8871 20851 8931
rect 20906 8871 20940 8931
rect 21551 8871 21585 8931
rect 21653 8871 21687 8931
rect 21761 8871 21795 8931
rect 22889 8871 22923 8931
rect 22993 8871 23027 8931
rect 23099 8871 23133 8931
rect 24101 8871 24135 8931
rect 24204 8871 24238 8931
rect 24311 8871 24345 8931
rect 24953 8871 24987 8931
rect 25043 8871 25077 8931
rect 19521 8563 19555 8597
rect 19521 8495 19555 8529
rect 19605 8563 19639 8597
rect 19605 8495 19639 8529
rect 19711 8563 19745 8597
rect 19711 8495 19745 8529
rect 19795 8563 19829 8597
rect 19795 8495 19829 8529
rect 26230 8563 26264 8597
rect 26230 8495 26264 8529
rect 26314 8563 26348 8597
rect 26314 8495 26348 8529
rect 26420 8563 26454 8597
rect 26420 8495 26454 8529
rect 26504 8563 26538 8597
rect 26504 8495 26538 8529
rect 10089 7866 10123 7900
rect 10173 7847 10207 7881
rect 10380 7862 10414 7896
rect 10615 7862 10649 7896
rect 10683 7862 10717 7896
rect 10767 7862 10801 7896
rect 10916 7866 10950 7900
rect 12702 8080 12736 8140
rect 12790 8080 12824 8140
rect 11000 7847 11034 7881
rect 11207 7862 11241 7896
rect 11442 7862 11476 7896
rect 11510 7862 11544 7896
rect 11594 7862 11628 7896
rect 11833 7880 11867 7940
rect 11929 7880 11963 7940
rect 12025 7880 12059 7940
rect 12121 7880 12155 7940
rect 12233 7892 12267 7952
rect 12321 7892 12355 7952
rect 11533 6605 11567 6639
rect 11619 6592 11653 6626
rect 11705 6622 11739 6656
rect 11809 6628 11843 6662
rect 11893 6596 11927 6630
rect 11977 6628 12011 6662
rect 12061 6596 12095 6630
rect 12145 6628 12179 6662
rect 12229 6660 12263 6694
rect 12229 6592 12263 6626
rect 12793 6660 12827 6694
rect 12793 6592 12827 6626
rect 12892 6628 12926 6662
rect 12976 6660 13010 6694
rect 12976 6592 13010 6626
rect 13076 6628 13110 6662
rect 13160 6618 13194 6652
rect 13369 6592 13403 6626
rect 13573 6592 13607 6626
rect 13677 6600 13711 6634
rect 13761 6618 13795 6652
rect 13846 6618 13880 6652
rect 13950 6592 13984 6626
rect 14049 6592 14083 6626
rect 14253 6606 14287 6640
rect 14445 6592 14479 6626
rect 14529 6618 14563 6652
rect 24075 6283 24109 6317
rect 24075 6215 24109 6249
rect 24159 6283 24193 6317
rect 24159 6215 24193 6249
rect 24265 6283 24299 6317
rect 24265 6215 24299 6249
rect 24349 6283 24383 6317
rect 24349 6215 24383 6249
rect 11532 5745 11566 5779
rect 11616 5719 11650 5753
rect 11700 5745 11734 5779
rect 11804 5719 11838 5753
rect 11888 5737 11922 5771
rect 11994 5719 12028 5753
rect 12211 5715 12245 5749
rect 12295 5735 12329 5769
rect 12395 5779 12429 5813
rect 12479 5753 12513 5787
rect 12583 5719 12617 5753
rect 12777 5719 12811 5753
rect 12968 5715 13002 5749
rect 13070 5735 13104 5769
rect 13170 5779 13204 5813
rect 13254 5727 13288 5761
rect 13358 5729 13392 5763
rect 13453 5719 13487 5753
rect 13537 5753 13571 5787
rect 13641 5745 13675 5779
rect 13736 5719 13770 5753
rect 13820 5755 13854 5789
rect 13924 5745 13958 5779
rect 14008 5719 14042 5753
rect 14092 5745 14126 5779
rect 14196 5719 14230 5753
rect 14280 5737 14314 5771
rect 14386 5719 14420 5753
rect 14603 5715 14637 5749
rect 14687 5735 14721 5769
rect 14787 5779 14821 5813
rect 14871 5753 14905 5787
rect 14975 5719 15009 5753
rect 15169 5719 15203 5753
rect 15360 5715 15394 5749
rect 15462 5735 15496 5769
rect 15562 5779 15596 5813
rect 15646 5727 15680 5761
rect 15750 5729 15784 5763
rect 15845 5719 15879 5753
rect 15929 5753 15963 5787
rect 16033 5745 16067 5779
rect 16128 5719 16162 5753
rect 16212 5755 16246 5789
rect 16316 5745 16350 5779
rect 16400 5719 16434 5753
rect 16484 5745 16518 5779
rect 16588 5719 16622 5753
rect 16672 5737 16706 5771
rect 16778 5719 16812 5753
rect 16995 5715 17029 5749
rect 17079 5735 17113 5769
rect 17179 5779 17213 5813
rect 17263 5753 17297 5787
rect 17367 5719 17401 5753
rect 17561 5719 17595 5753
rect 17752 5715 17786 5749
rect 17854 5735 17888 5769
rect 17954 5779 17988 5813
rect 18038 5727 18072 5761
rect 18142 5729 18176 5763
rect 18237 5719 18271 5753
rect 18321 5753 18355 5787
rect 18425 5745 18459 5779
rect 18520 5719 18554 5753
rect 18604 5755 18638 5789
rect 18708 5745 18742 5779
rect 18792 5719 18826 5753
rect 18876 5745 18910 5779
rect 18980 5719 19014 5753
rect 19064 5737 19098 5771
rect 19170 5719 19204 5753
rect 19387 5715 19421 5749
rect 19471 5735 19505 5769
rect 19571 5779 19605 5813
rect 19655 5753 19689 5787
rect 19759 5719 19793 5753
rect 19953 5719 19987 5753
rect 20144 5715 20178 5749
rect 20246 5735 20280 5769
rect 20346 5779 20380 5813
rect 20430 5727 20464 5761
rect 20534 5729 20568 5763
rect 20629 5719 20663 5753
rect 20713 5753 20747 5787
rect 20817 5745 20851 5779
rect 20912 5719 20946 5753
rect 20996 5755 21030 5789
rect 21100 5745 21134 5779
rect 21184 5719 21218 5753
rect 21268 5745 21302 5779
rect 21372 5719 21406 5753
rect 21456 5737 21490 5771
rect 21562 5719 21596 5753
rect 21779 5715 21813 5749
rect 21863 5735 21897 5769
rect 21963 5779 21997 5813
rect 22047 5753 22081 5787
rect 22151 5719 22185 5753
rect 22345 5719 22379 5753
rect 22536 5715 22570 5749
rect 22638 5735 22672 5769
rect 22738 5779 22772 5813
rect 22822 5727 22856 5761
rect 22926 5729 22960 5763
rect 23021 5719 23055 5753
rect 25536 5881 25570 5941
rect 25626 5881 25660 5941
rect 26268 5881 26302 5941
rect 26375 5881 26409 5941
rect 26478 5881 26512 5941
rect 27480 5881 27514 5941
rect 27586 5881 27620 5941
rect 27690 5881 27724 5941
rect 28818 5881 28852 5941
rect 28926 5881 28960 5941
rect 29028 5881 29062 5941
rect 29673 5881 29707 5941
rect 29762 5881 29796 5941
rect 30326 5882 30360 5942
rect 30414 5882 30448 5942
rect 30510 5882 30544 5942
rect 30606 5882 30640 5942
rect 23105 5753 23139 5787
rect 23209 5745 23243 5779
rect 23304 5719 23338 5753
rect 23388 5755 23422 5789
rect 30714 5847 30748 5881
rect 30807 5834 30841 5868
rect 30893 5864 30927 5898
rect 30977 5906 31011 5940
rect 30977 5838 31011 5872
rect 24516 5697 24550 5757
rect 24676 5697 24710 5757
rect 30326 5744 30360 5804
rect 30414 5744 30448 5804
rect 24516 5559 24550 5619
rect 24676 5559 24710 5619
rect 11092 5043 11126 5077
rect 11178 5030 11212 5064
rect 11264 5060 11298 5094
rect 11368 5066 11402 5100
rect 11452 5034 11486 5068
rect 11536 5066 11570 5100
rect 11620 5034 11654 5068
rect 11704 5066 11738 5100
rect 11788 5098 11822 5132
rect 11788 5030 11822 5064
rect 11900 5102 11934 5136
rect 11900 5034 11934 5068
rect 11984 5102 12018 5136
rect 11984 5034 12018 5068
rect 12068 5034 12102 5068
rect 12152 5102 12186 5136
rect 12152 5034 12186 5068
rect 12236 5034 12270 5068
rect 12320 5102 12354 5136
rect 12320 5034 12354 5068
rect 12404 5034 12438 5068
rect 12488 5102 12522 5136
rect 12488 5034 12522 5068
rect 12572 5034 12606 5068
rect 12656 5102 12690 5136
rect 12656 5034 12690 5068
rect 12740 5034 12774 5068
rect 12824 5102 12858 5136
rect 12824 5034 12858 5068
rect 12908 5034 12942 5068
rect 12992 5102 13026 5136
rect 12992 5034 13026 5068
rect 13076 5034 13110 5068
rect 13160 5102 13194 5136
rect 13160 5034 13194 5068
rect 13244 5034 13278 5068
rect 13328 5102 13362 5136
rect 13328 5034 13362 5068
rect 13412 5034 13446 5068
rect 13496 5102 13530 5136
rect 13496 5034 13530 5068
rect 13580 5034 13614 5068
rect 13664 5102 13698 5136
rect 13664 5034 13698 5068
rect 13748 5034 13782 5068
rect 13924 5066 13958 5100
rect 14008 5030 14042 5064
rect 14103 5056 14137 5090
rect 14207 5064 14241 5098
rect 14291 5030 14325 5064
rect 14386 5040 14420 5074
rect 14490 5038 14524 5072
rect 14574 5090 14608 5124
rect 14674 5046 14708 5080
rect 14776 5026 14810 5060
rect 14967 5030 15001 5064
rect 15161 5030 15195 5064
rect 15265 5064 15299 5098
rect 15349 5090 15383 5124
rect 15449 5046 15483 5080
rect 15533 5026 15567 5060
rect 15750 5030 15784 5064
rect 15856 5048 15890 5082
rect 15940 5030 15974 5064
rect 16044 5056 16078 5090
rect 16128 5030 16162 5064
rect 16212 5056 16246 5090
rect 16316 5066 16350 5100
rect 16400 5030 16434 5064
rect 16495 5056 16529 5090
rect 16599 5064 16633 5098
rect 16683 5030 16717 5064
rect 16778 5040 16812 5074
rect 16882 5038 16916 5072
rect 16966 5090 17000 5124
rect 17066 5046 17100 5080
rect 17168 5026 17202 5060
rect 17359 5030 17393 5064
rect 17553 5030 17587 5064
rect 17657 5064 17691 5098
rect 17741 5090 17775 5124
rect 17841 5046 17875 5080
rect 17925 5026 17959 5060
rect 18142 5030 18176 5064
rect 18248 5048 18282 5082
rect 18332 5030 18366 5064
rect 18436 5056 18470 5090
rect 18520 5030 18554 5064
rect 18604 5056 18638 5090
rect 18708 5066 18742 5100
rect 18792 5030 18826 5064
rect 18887 5056 18921 5090
rect 18991 5064 19025 5098
rect 19075 5030 19109 5064
rect 19170 5040 19204 5074
rect 19274 5038 19308 5072
rect 19358 5090 19392 5124
rect 19458 5046 19492 5080
rect 19560 5026 19594 5060
rect 19751 5030 19785 5064
rect 19945 5030 19979 5064
rect 20049 5064 20083 5098
rect 20133 5090 20167 5124
rect 20233 5046 20267 5080
rect 20317 5026 20351 5060
rect 20534 5030 20568 5064
rect 20640 5048 20674 5082
rect 20724 5030 20758 5064
rect 20828 5056 20862 5090
rect 20912 5030 20946 5064
rect 20996 5056 21030 5090
rect 21100 5066 21134 5100
rect 21184 5030 21218 5064
rect 21279 5056 21313 5090
rect 21383 5064 21417 5098
rect 21467 5030 21501 5064
rect 21562 5040 21596 5074
rect 21666 5038 21700 5072
rect 21750 5090 21784 5124
rect 21850 5046 21884 5080
rect 21952 5026 21986 5060
rect 22143 5030 22177 5064
rect 22337 5030 22371 5064
rect 22441 5064 22475 5098
rect 22525 5090 22559 5124
rect 24516 5421 24550 5481
rect 24676 5421 24710 5481
rect 24516 5283 24550 5343
rect 24676 5283 24710 5343
rect 22625 5046 22659 5080
rect 22709 5026 22743 5060
rect 24516 5145 24550 5205
rect 24676 5145 24710 5205
rect 22926 5030 22960 5064
rect 23032 5048 23066 5082
rect 23116 5030 23150 5064
rect 23220 5056 23254 5090
rect 23304 5030 23338 5064
rect 23388 5056 23422 5090
rect 24516 5007 24550 5067
rect 24676 5007 24710 5067
rect 24516 4869 24550 4929
rect 24676 4869 24710 4929
rect 24516 4731 24550 4791
rect 24676 4731 24710 4791
rect 11124 4169 11158 4203
rect 11210 4156 11244 4190
rect 11296 4186 11330 4220
rect 11400 4192 11434 4226
rect 11484 4160 11518 4194
rect 11568 4192 11602 4226
rect 11652 4160 11686 4194
rect 11736 4192 11770 4226
rect 11820 4224 11854 4258
rect 11820 4156 11854 4190
rect 13707 4229 13741 4263
rect 13707 4161 13741 4195
rect 13791 4229 13825 4263
rect 13791 4161 13825 4195
rect 13923 4183 13957 4217
rect 14007 4157 14041 4191
rect 14091 4183 14125 4217
rect 14195 4157 14229 4191
rect 14279 4175 14313 4209
rect 14385 4157 14419 4191
rect 14602 4153 14636 4187
rect 14686 4173 14720 4207
rect 14786 4217 14820 4251
rect 14870 4191 14904 4225
rect 14974 4157 15008 4191
rect 15168 4157 15202 4191
rect 15359 4153 15393 4187
rect 15461 4173 15495 4207
rect 15561 4217 15595 4251
rect 15645 4165 15679 4199
rect 15749 4167 15783 4201
rect 15844 4157 15878 4191
rect 15928 4191 15962 4225
rect 16032 4183 16066 4217
rect 16127 4157 16161 4191
rect 16211 4193 16245 4227
rect 16315 4183 16349 4217
rect 16399 4157 16433 4191
rect 16483 4183 16517 4217
rect 16587 4157 16621 4191
rect 16671 4175 16705 4209
rect 16777 4157 16811 4191
rect 16994 4153 17028 4187
rect 17078 4173 17112 4207
rect 17178 4217 17212 4251
rect 17262 4191 17296 4225
rect 17366 4157 17400 4191
rect 17560 4157 17594 4191
rect 17751 4153 17785 4187
rect 17853 4173 17887 4207
rect 17953 4217 17987 4251
rect 18037 4165 18071 4199
rect 18141 4167 18175 4201
rect 18236 4157 18270 4191
rect 18320 4191 18354 4225
rect 18424 4183 18458 4217
rect 18519 4157 18553 4191
rect 18603 4193 18637 4227
rect 18707 4183 18741 4217
rect 18791 4157 18825 4191
rect 18875 4183 18909 4217
rect 18979 4157 19013 4191
rect 19063 4175 19097 4209
rect 19169 4157 19203 4191
rect 19386 4153 19420 4187
rect 19470 4173 19504 4207
rect 19570 4217 19604 4251
rect 19654 4191 19688 4225
rect 19758 4157 19792 4191
rect 19952 4157 19986 4191
rect 20143 4153 20177 4187
rect 20245 4173 20279 4207
rect 20345 4217 20379 4251
rect 20429 4165 20463 4199
rect 20533 4167 20567 4201
rect 20628 4157 20662 4191
rect 20712 4191 20746 4225
rect 20816 4183 20850 4217
rect 20911 4157 20945 4191
rect 20995 4193 21029 4227
rect 21099 4183 21133 4217
rect 21183 4157 21217 4191
rect 21267 4183 21301 4217
rect 21371 4157 21405 4191
rect 21455 4175 21489 4209
rect 21561 4157 21595 4191
rect 21778 4153 21812 4187
rect 21862 4173 21896 4207
rect 21962 4217 21996 4251
rect 22046 4191 22080 4225
rect 22150 4157 22184 4191
rect 22344 4157 22378 4191
rect 22535 4153 22569 4187
rect 22637 4173 22671 4207
rect 22737 4217 22771 4251
rect 22821 4165 22855 4199
rect 22925 4167 22959 4201
rect 23020 4157 23054 4191
rect 23104 4191 23138 4225
rect 23208 4183 23242 4217
rect 23303 4157 23337 4191
rect 23387 4193 23421 4227
rect 25612 4162 25646 4196
rect 25696 4188 25730 4222
rect 25780 4162 25814 4196
rect 25884 4188 25918 4222
rect 25968 4170 26002 4204
rect 26074 4188 26108 4222
rect 26291 4192 26325 4226
rect 26375 4172 26409 4206
rect 26475 4128 26509 4162
rect 26559 4154 26593 4188
rect 26663 4188 26697 4222
rect 26857 4188 26891 4222
rect 27048 4192 27082 4226
rect 27150 4172 27184 4206
rect 27250 4128 27284 4162
rect 27334 4180 27368 4214
rect 27438 4178 27472 4212
rect 27533 4188 27567 4222
rect 27617 4154 27651 4188
rect 27721 4162 27755 4196
rect 27816 4188 27850 4222
rect 27900 4152 27934 4186
rect 28004 4162 28038 4196
rect 28088 4188 28122 4222
rect 28172 4162 28206 4196
rect 28276 4188 28310 4222
rect 28360 4170 28394 4204
rect 28466 4188 28500 4222
rect 28683 4192 28717 4226
rect 28767 4172 28801 4206
rect 28867 4128 28901 4162
rect 28951 4154 28985 4188
rect 29055 4188 29089 4222
rect 29249 4188 29283 4222
rect 29440 4192 29474 4226
rect 29542 4172 29576 4206
rect 29642 4128 29676 4162
rect 29726 4180 29760 4214
rect 29830 4178 29864 4212
rect 29925 4188 29959 4222
rect 30009 4154 30043 4188
rect 30113 4162 30147 4196
rect 30208 4188 30242 4222
rect 30292 4152 30326 4186
rect 11531 3320 11565 3354
rect 11615 3284 11649 3318
rect 11710 3310 11744 3344
rect 11814 3318 11848 3352
rect 11898 3284 11932 3318
rect 11993 3294 12027 3328
rect 12097 3292 12131 3326
rect 12181 3344 12215 3378
rect 12281 3300 12315 3334
rect 12383 3280 12417 3314
rect 12574 3284 12608 3318
rect 12768 3284 12802 3318
rect 12872 3318 12906 3352
rect 12956 3344 12990 3378
rect 13056 3300 13090 3334
rect 13140 3280 13174 3314
rect 13357 3284 13391 3318
rect 13463 3302 13497 3336
rect 13547 3284 13581 3318
rect 13651 3310 13685 3344
rect 13735 3284 13769 3318
rect 13819 3310 13853 3344
rect 13923 3320 13957 3354
rect 14007 3284 14041 3318
rect 14102 3310 14136 3344
rect 14206 3318 14240 3352
rect 14290 3284 14324 3318
rect 14385 3294 14419 3328
rect 14489 3292 14523 3326
rect 14573 3344 14607 3378
rect 14673 3300 14707 3334
rect 14775 3280 14809 3314
rect 14966 3284 15000 3318
rect 15160 3284 15194 3318
rect 15264 3318 15298 3352
rect 15348 3344 15382 3378
rect 15448 3300 15482 3334
rect 15532 3280 15566 3314
rect 15749 3284 15783 3318
rect 15855 3302 15889 3336
rect 15939 3284 15973 3318
rect 16043 3310 16077 3344
rect 16127 3284 16161 3318
rect 16211 3310 16245 3344
rect 16315 3320 16349 3354
rect 16399 3284 16433 3318
rect 16494 3310 16528 3344
rect 16598 3318 16632 3352
rect 16682 3284 16716 3318
rect 16777 3294 16811 3328
rect 16881 3292 16915 3326
rect 16965 3344 16999 3378
rect 17065 3300 17099 3334
rect 17167 3280 17201 3314
rect 17358 3284 17392 3318
rect 17552 3284 17586 3318
rect 17656 3318 17690 3352
rect 17740 3344 17774 3378
rect 17840 3300 17874 3334
rect 17924 3280 17958 3314
rect 18141 3284 18175 3318
rect 18247 3302 18281 3336
rect 18331 3284 18365 3318
rect 18435 3310 18469 3344
rect 18519 3284 18553 3318
rect 18603 3310 18637 3344
rect 18707 3320 18741 3354
rect 18791 3284 18825 3318
rect 18886 3310 18920 3344
rect 18990 3318 19024 3352
rect 19074 3284 19108 3318
rect 19169 3294 19203 3328
rect 19273 3292 19307 3326
rect 19357 3344 19391 3378
rect 19457 3300 19491 3334
rect 19559 3280 19593 3314
rect 19750 3284 19784 3318
rect 19944 3284 19978 3318
rect 20048 3318 20082 3352
rect 20132 3344 20166 3378
rect 20232 3300 20266 3334
rect 20316 3280 20350 3314
rect 20533 3284 20567 3318
rect 20639 3302 20673 3336
rect 20723 3284 20757 3318
rect 20827 3310 20861 3344
rect 20911 3284 20945 3318
rect 20995 3310 21029 3344
rect 21099 3320 21133 3354
rect 21183 3284 21217 3318
rect 21278 3310 21312 3344
rect 21382 3318 21416 3352
rect 21466 3284 21500 3318
rect 21561 3294 21595 3328
rect 21665 3292 21699 3326
rect 21749 3344 21783 3378
rect 21849 3300 21883 3334
rect 21951 3280 21985 3314
rect 22142 3284 22176 3318
rect 22336 3284 22370 3318
rect 22440 3318 22474 3352
rect 22524 3344 22558 3378
rect 22624 3300 22658 3334
rect 22708 3280 22742 3314
rect 22925 3284 22959 3318
rect 23031 3302 23065 3336
rect 23115 3284 23149 3318
rect 23219 3310 23253 3344
rect 23303 3284 23337 3318
rect 23387 3310 23421 3344
rect 25612 3182 25646 3216
rect 25696 3156 25730 3190
rect 25780 3182 25814 3216
rect 25884 3156 25918 3190
rect 25968 3174 26002 3208
rect 26074 3156 26108 3190
rect 26291 3152 26325 3186
rect 26375 3172 26409 3206
rect 26475 3216 26509 3250
rect 26559 3190 26593 3224
rect 26663 3156 26697 3190
rect 26857 3156 26891 3190
rect 27048 3152 27082 3186
rect 27150 3172 27184 3206
rect 27250 3216 27284 3250
rect 27334 3164 27368 3198
rect 27438 3166 27472 3200
rect 27533 3156 27567 3190
rect 27617 3190 27651 3224
rect 27721 3182 27755 3216
rect 27816 3156 27850 3190
rect 27900 3192 27934 3226
rect 28004 3182 28038 3216
rect 28088 3156 28122 3190
rect 28172 3182 28206 3216
rect 28276 3156 28310 3190
rect 28360 3174 28394 3208
rect 28466 3156 28500 3190
rect 28683 3152 28717 3186
rect 28767 3172 28801 3206
rect 28867 3216 28901 3250
rect 28951 3190 28985 3224
rect 29055 3156 29089 3190
rect 29249 3156 29283 3190
rect 29440 3152 29474 3186
rect 29542 3172 29576 3206
rect 29642 3216 29676 3250
rect 29726 3164 29760 3198
rect 29830 3166 29864 3200
rect 29925 3156 29959 3190
rect 30009 3190 30043 3224
rect 30113 3182 30147 3216
rect 30208 3156 30242 3190
rect 30292 3192 30326 3226
rect 25612 2882 25646 2916
rect 25696 2908 25730 2942
rect 25780 2882 25814 2916
rect 25884 2908 25918 2942
rect 25968 2890 26002 2924
rect 26074 2908 26108 2942
rect 26291 2912 26325 2946
rect 26375 2892 26409 2926
rect 26475 2848 26509 2882
rect 26559 2874 26593 2908
rect 26663 2908 26697 2942
rect 26857 2908 26891 2942
rect 27048 2912 27082 2946
rect 27150 2892 27184 2926
rect 27250 2848 27284 2882
rect 27334 2900 27368 2934
rect 27438 2898 27472 2932
rect 27533 2908 27567 2942
rect 27617 2874 27651 2908
rect 27721 2882 27755 2916
rect 27816 2908 27850 2942
rect 27900 2872 27934 2906
rect 28004 2882 28038 2916
rect 28088 2908 28122 2942
rect 28172 2882 28206 2916
rect 28276 2908 28310 2942
rect 28360 2890 28394 2924
rect 28466 2908 28500 2942
rect 28683 2912 28717 2946
rect 28767 2892 28801 2926
rect 28867 2848 28901 2882
rect 28951 2874 28985 2908
rect 29055 2908 29089 2942
rect 29249 2908 29283 2942
rect 29440 2912 29474 2946
rect 29542 2892 29576 2926
rect 29642 2848 29676 2882
rect 29726 2900 29760 2934
rect 29830 2898 29864 2932
rect 29925 2908 29959 2942
rect 30009 2874 30043 2908
rect 30113 2882 30147 2916
rect 30208 2908 30242 2942
rect 30292 2872 30326 2906
rect 25612 1902 25646 1936
rect 25696 1876 25730 1910
rect 25780 1902 25814 1936
rect 25884 1876 25918 1910
rect 25968 1894 26002 1928
rect 26074 1876 26108 1910
rect 26291 1872 26325 1906
rect 26375 1892 26409 1926
rect 26475 1936 26509 1970
rect 26559 1910 26593 1944
rect 26663 1876 26697 1910
rect 26857 1876 26891 1910
rect 27048 1872 27082 1906
rect 27150 1892 27184 1926
rect 27250 1936 27284 1970
rect 27334 1884 27368 1918
rect 27438 1886 27472 1920
rect 27533 1876 27567 1910
rect 27617 1910 27651 1944
rect 27721 1902 27755 1936
rect 27816 1876 27850 1910
rect 27900 1912 27934 1946
rect 28004 1902 28038 1936
rect 28088 1876 28122 1910
rect 28172 1902 28206 1936
rect 28276 1876 28310 1910
rect 28360 1894 28394 1928
rect 28466 1876 28500 1910
rect 28683 1872 28717 1906
rect 28767 1892 28801 1926
rect 28867 1936 28901 1970
rect 28951 1910 28985 1944
rect 29055 1876 29089 1910
rect 29249 1876 29283 1910
rect 29440 1872 29474 1906
rect 29542 1892 29576 1926
rect 29642 1936 29676 1970
rect 29726 1884 29760 1918
rect 29830 1886 29864 1920
rect 29925 1876 29959 1910
rect 30009 1910 30043 1944
rect 30113 1902 30147 1936
rect 30208 1876 30242 1910
rect 30292 1912 30326 1946
rect 8612 917 8646 951
rect 8698 904 8732 938
rect 8784 934 8818 968
rect 8888 940 8922 974
rect 8972 908 9006 942
rect 9056 940 9090 974
rect 9140 908 9174 942
rect 9224 940 9258 974
rect 9308 972 9342 1006
rect 9308 904 9342 938
rect 9440 976 9474 1010
rect 9440 908 9474 942
rect 9524 976 9558 1010
rect 9524 908 9558 942
rect 9608 908 9642 942
rect 9692 976 9726 1010
rect 9692 908 9726 942
rect 9776 908 9810 942
rect 9860 976 9894 1010
rect 9860 908 9894 942
rect 9944 908 9978 942
rect 10028 976 10062 1010
rect 10028 908 10062 942
rect 10112 908 10146 942
rect 10196 976 10230 1010
rect 10196 908 10230 942
rect 10280 908 10314 942
rect 10364 976 10398 1010
rect 10364 908 10398 942
rect 10448 908 10482 942
rect 10532 976 10566 1010
rect 10532 908 10566 942
rect 10616 908 10650 942
rect 10700 976 10734 1010
rect 10700 908 10734 942
rect 10784 908 10818 942
rect 10868 976 10902 1010
rect 10868 908 10902 942
rect 10952 908 10986 942
rect 11036 976 11070 1010
rect 11036 908 11070 942
rect 11120 908 11154 942
rect 11204 976 11238 1010
rect 11204 908 11238 942
rect 11288 908 11322 942
rect 12996 917 13030 951
rect 13082 904 13116 938
rect 13168 934 13202 968
rect 13272 940 13306 974
rect 13356 908 13390 942
rect 13440 940 13474 974
rect 13524 908 13558 942
rect 13608 940 13642 974
rect 13692 972 13726 1006
rect 13692 904 13726 938
rect 13824 976 13858 1010
rect 13824 908 13858 942
rect 13908 976 13942 1010
rect 13908 908 13942 942
rect 13992 908 14026 942
rect 14076 976 14110 1010
rect 14076 908 14110 942
rect 14160 908 14194 942
rect 14244 976 14278 1010
rect 14244 908 14278 942
rect 14328 908 14362 942
rect 14412 976 14446 1010
rect 14412 908 14446 942
rect 14496 908 14530 942
rect 14580 976 14614 1010
rect 14580 908 14614 942
rect 14664 908 14698 942
rect 14748 976 14782 1010
rect 14748 908 14782 942
rect 14832 908 14866 942
rect 14916 976 14950 1010
rect 14916 908 14950 942
rect 15000 908 15034 942
rect 15084 976 15118 1010
rect 15084 908 15118 942
rect 15168 908 15202 942
rect 15252 976 15286 1010
rect 15252 908 15286 942
rect 15336 908 15370 942
rect 15420 976 15454 1010
rect 15420 908 15454 942
rect 15504 908 15538 942
rect 15588 976 15622 1010
rect 15588 908 15622 942
rect 15672 908 15706 942
rect 8610 -219 8644 -185
rect 8694 -238 8728 -204
rect 8901 -223 8935 -189
rect 9136 -223 9170 -189
rect 9204 -223 9238 -189
rect 9288 -223 9322 -189
rect 10090 -223 10124 -189
rect 10174 -223 10208 -189
rect 10242 -223 10276 -189
rect 10477 -223 10511 -189
rect 10684 -238 10718 -204
rect 10768 -219 10802 -185
rect 11002 -219 11036 -185
rect 11086 -238 11120 -204
rect 11293 -223 11327 -189
rect 11528 -223 11562 -189
rect 11596 -223 11630 -189
rect 11680 -223 11714 -189
rect 12482 -223 12516 -189
rect 12566 -223 12600 -189
rect 12634 -223 12668 -189
rect 12869 -223 12903 -189
rect 13076 -238 13110 -204
rect 13160 -219 13194 -185
rect 13394 -219 13428 -185
rect 13478 -238 13512 -204
rect 13685 -223 13719 -189
rect 13920 -223 13954 -189
rect 13988 -223 14022 -189
rect 14072 -223 14106 -189
rect 14872 -223 14906 -189
rect 14956 -223 14990 -189
rect 15024 -223 15058 -189
rect 15259 -223 15293 -189
rect 15466 -238 15500 -204
rect 15550 -219 15584 -185
rect 15786 -219 15820 -185
rect 15870 -238 15904 -204
rect 16077 -223 16111 -189
rect 16312 -223 16346 -189
rect 16380 -223 16414 -189
rect 16464 -223 16498 -189
rect 17266 -223 17300 -189
rect 17350 -223 17384 -189
rect 17418 -223 17452 -189
rect 17653 -223 17687 -189
rect 17860 -238 17894 -204
rect 17944 -219 17978 -185
rect 18178 -219 18212 -185
rect 18262 -238 18296 -204
rect 18469 -223 18503 -189
rect 18704 -223 18738 -189
rect 18772 -223 18806 -189
rect 18856 -223 18890 -189
rect 19658 -223 19692 -189
rect 19742 -223 19776 -189
rect 19810 -223 19844 -189
rect 20045 -223 20079 -189
rect 20252 -238 20286 -204
rect 20336 -219 20370 -185
rect 20570 -219 20604 -185
rect 20654 -238 20688 -204
rect 20861 -223 20895 -189
rect 21096 -223 21130 -189
rect 21164 -223 21198 -189
rect 21248 -223 21282 -189
rect 22048 -223 22082 -189
rect 22132 -223 22166 -189
rect 22200 -223 22234 -189
rect 22435 -223 22469 -189
rect 22642 -238 22676 -204
rect 22726 -219 22760 -185
rect 22962 -219 22996 -185
rect 23046 -238 23080 -204
rect 23253 -223 23287 -189
rect 23488 -223 23522 -189
rect 23556 -223 23590 -189
rect 23640 -223 23674 -189
rect 24442 -223 24476 -189
rect 24526 -223 24560 -189
rect 24594 -223 24628 -189
rect 24829 -223 24863 -189
rect 25036 -238 25070 -204
rect 25120 -219 25154 -185
rect 8610 -900 8644 -866
rect 8694 -926 8728 -892
rect 8778 -900 8812 -866
rect 8882 -926 8916 -892
rect 8966 -908 9000 -874
rect 9071 -926 9105 -892
rect 9292 -930 9326 -896
rect 9376 -924 9410 -890
rect 9472 -866 9506 -832
rect 9556 -892 9590 -858
rect 9660 -926 9694 -892
rect 9864 -926 9898 -892
rect 10056 -930 10090 -896
rect 10140 -910 10174 -876
rect 10248 -852 10282 -818
rect 10332 -918 10366 -884
rect 10436 -916 10470 -882
rect 10531 -926 10565 -892
rect 10615 -892 10649 -858
rect 10719 -900 10753 -866
rect 10814 -926 10848 -892
rect 10898 -890 10932 -856
rect 11002 -900 11036 -866
rect 11086 -926 11120 -892
rect 11170 -900 11204 -866
rect 11274 -926 11308 -892
rect 11358 -908 11392 -874
rect 11463 -926 11497 -892
rect 11684 -930 11718 -896
rect 11768 -924 11802 -890
rect 11864 -866 11898 -832
rect 11948 -892 11982 -858
rect 12052 -926 12086 -892
rect 12256 -926 12290 -892
rect 12448 -930 12482 -896
rect 12532 -910 12566 -876
rect 12640 -852 12674 -818
rect 12724 -918 12758 -884
rect 12828 -916 12862 -882
rect 12923 -926 12957 -892
rect 13007 -892 13041 -858
rect 13111 -900 13145 -866
rect 13206 -926 13240 -892
rect 13290 -890 13324 -856
rect 13394 -900 13428 -866
rect 13478 -926 13512 -892
rect 13562 -900 13596 -866
rect 13666 -926 13700 -892
rect 13750 -908 13784 -874
rect 13855 -926 13889 -892
rect 14076 -930 14110 -896
rect 14160 -924 14194 -890
rect 14256 -866 14290 -832
rect 14340 -892 14374 -858
rect 14444 -926 14478 -892
rect 14648 -926 14682 -892
rect 14840 -930 14874 -896
rect 14924 -910 14958 -876
rect 15032 -852 15066 -818
rect 15116 -918 15150 -884
rect 15220 -916 15254 -882
rect 15315 -926 15349 -892
rect 15399 -892 15433 -858
rect 15503 -900 15537 -866
rect 15598 -926 15632 -892
rect 15682 -890 15716 -856
rect 15786 -900 15820 -866
rect 15870 -926 15904 -892
rect 15954 -900 15988 -866
rect 16058 -926 16092 -892
rect 16142 -908 16176 -874
rect 16247 -926 16281 -892
rect 16468 -930 16502 -896
rect 16552 -924 16586 -890
rect 16648 -866 16682 -832
rect 16732 -892 16766 -858
rect 16836 -926 16870 -892
rect 17040 -926 17074 -892
rect 17232 -930 17266 -896
rect 17316 -910 17350 -876
rect 17424 -852 17458 -818
rect 17508 -918 17542 -884
rect 17612 -916 17646 -882
rect 17707 -926 17741 -892
rect 17791 -892 17825 -858
rect 17895 -900 17929 -866
rect 17990 -926 18024 -892
rect 18074 -890 18108 -856
rect 18178 -900 18212 -866
rect 18262 -926 18296 -892
rect 18346 -900 18380 -866
rect 18450 -926 18484 -892
rect 18534 -908 18568 -874
rect 18639 -926 18673 -892
rect 18860 -930 18894 -896
rect 18944 -924 18978 -890
rect 19040 -866 19074 -832
rect 19124 -892 19158 -858
rect 19228 -926 19262 -892
rect 19432 -926 19466 -892
rect 19624 -930 19658 -896
rect 19708 -910 19742 -876
rect 19816 -852 19850 -818
rect 19900 -918 19934 -884
rect 20004 -916 20038 -882
rect 20099 -926 20133 -892
rect 20183 -892 20217 -858
rect 20287 -900 20321 -866
rect 20382 -926 20416 -892
rect 20466 -890 20500 -856
rect 20570 -900 20604 -866
rect 20654 -926 20688 -892
rect 20738 -900 20772 -866
rect 20842 -926 20876 -892
rect 20926 -908 20960 -874
rect 21031 -926 21065 -892
rect 21252 -930 21286 -896
rect 21336 -924 21370 -890
rect 21432 -866 21466 -832
rect 21516 -892 21550 -858
rect 21620 -926 21654 -892
rect 21824 -926 21858 -892
rect 22016 -930 22050 -896
rect 22100 -910 22134 -876
rect 22208 -852 22242 -818
rect 22292 -918 22326 -884
rect 22396 -916 22430 -882
rect 22491 -926 22525 -892
rect 22575 -892 22609 -858
rect 22679 -900 22713 -866
rect 22774 -926 22808 -892
rect 22858 -890 22892 -856
rect 22962 -900 22996 -866
rect 23046 -926 23080 -892
rect 23130 -900 23164 -866
rect 23234 -926 23268 -892
rect 23318 -908 23352 -874
rect 23423 -926 23457 -892
rect 23644 -930 23678 -896
rect 23728 -924 23762 -890
rect 23824 -866 23858 -832
rect 23908 -892 23942 -858
rect 24012 -926 24046 -892
rect 24216 -926 24250 -892
rect 24408 -930 24442 -896
rect 24492 -910 24526 -876
rect 24600 -852 24634 -818
rect 24684 -918 24718 -884
rect 24788 -916 24822 -882
rect 24883 -926 24917 -892
rect 24967 -892 25001 -858
rect 25071 -900 25105 -866
rect 25166 -926 25200 -892
rect 25250 -890 25284 -856
rect 8610 -1579 8644 -1545
rect 8694 -1615 8728 -1581
rect 8789 -1589 8823 -1555
rect 8893 -1581 8927 -1547
rect 8977 -1615 9011 -1581
rect 9072 -1605 9106 -1571
rect 9176 -1607 9210 -1573
rect 9260 -1541 9294 -1507
rect 9368 -1599 9402 -1565
rect 9452 -1619 9486 -1585
rect 9644 -1615 9678 -1581
rect 9848 -1615 9882 -1581
rect 9952 -1581 9986 -1547
rect 10036 -1555 10070 -1521
rect 10132 -1613 10166 -1579
rect 10216 -1619 10250 -1585
rect 10437 -1615 10471 -1581
rect 10542 -1597 10576 -1563
rect 10626 -1615 10660 -1581
rect 10730 -1589 10764 -1555
rect 10814 -1615 10848 -1581
rect 10898 -1589 10932 -1555
rect 11002 -1579 11036 -1545
rect 11086 -1615 11120 -1581
rect 11181 -1589 11215 -1555
rect 11285 -1581 11319 -1547
rect 11369 -1615 11403 -1581
rect 11464 -1605 11498 -1571
rect 11568 -1607 11602 -1573
rect 11652 -1541 11686 -1507
rect 11760 -1599 11794 -1565
rect 11844 -1619 11878 -1585
rect 12036 -1615 12070 -1581
rect 12240 -1615 12274 -1581
rect 12344 -1581 12378 -1547
rect 12428 -1555 12462 -1521
rect 12524 -1613 12558 -1579
rect 12608 -1619 12642 -1585
rect 12829 -1615 12863 -1581
rect 12934 -1597 12968 -1563
rect 13018 -1615 13052 -1581
rect 13122 -1589 13156 -1555
rect 13206 -1615 13240 -1581
rect 13290 -1589 13324 -1555
rect 13394 -1579 13428 -1545
rect 13478 -1615 13512 -1581
rect 13573 -1589 13607 -1555
rect 13677 -1581 13711 -1547
rect 13761 -1615 13795 -1581
rect 13856 -1605 13890 -1571
rect 13960 -1607 13994 -1573
rect 14044 -1541 14078 -1507
rect 14152 -1599 14186 -1565
rect 14236 -1619 14270 -1585
rect 14428 -1615 14462 -1581
rect 14632 -1615 14666 -1581
rect 14736 -1581 14770 -1547
rect 14820 -1555 14854 -1521
rect 14916 -1613 14950 -1579
rect 15000 -1619 15034 -1585
rect 15221 -1615 15255 -1581
rect 15326 -1597 15360 -1563
rect 15410 -1615 15444 -1581
rect 15514 -1589 15548 -1555
rect 15598 -1615 15632 -1581
rect 15682 -1589 15716 -1555
rect 15786 -1579 15820 -1545
rect 15870 -1615 15904 -1581
rect 15965 -1589 15999 -1555
rect 16069 -1581 16103 -1547
rect 16153 -1615 16187 -1581
rect 16248 -1605 16282 -1571
rect 16352 -1607 16386 -1573
rect 16436 -1541 16470 -1507
rect 16544 -1599 16578 -1565
rect 16628 -1619 16662 -1585
rect 16820 -1615 16854 -1581
rect 17024 -1615 17058 -1581
rect 17128 -1581 17162 -1547
rect 17212 -1555 17246 -1521
rect 17308 -1613 17342 -1579
rect 17392 -1619 17426 -1585
rect 17613 -1615 17647 -1581
rect 17718 -1597 17752 -1563
rect 17802 -1615 17836 -1581
rect 17906 -1589 17940 -1555
rect 17990 -1615 18024 -1581
rect 18074 -1589 18108 -1555
rect 18178 -1579 18212 -1545
rect 18262 -1615 18296 -1581
rect 18357 -1589 18391 -1555
rect 18461 -1581 18495 -1547
rect 18545 -1615 18579 -1581
rect 18640 -1605 18674 -1571
rect 18744 -1607 18778 -1573
rect 18828 -1541 18862 -1507
rect 18936 -1599 18970 -1565
rect 19020 -1619 19054 -1585
rect 19212 -1615 19246 -1581
rect 19416 -1615 19450 -1581
rect 19520 -1581 19554 -1547
rect 19604 -1555 19638 -1521
rect 19700 -1613 19734 -1579
rect 19784 -1619 19818 -1585
rect 20005 -1615 20039 -1581
rect 20110 -1597 20144 -1563
rect 20194 -1615 20228 -1581
rect 20298 -1589 20332 -1555
rect 20382 -1615 20416 -1581
rect 20466 -1589 20500 -1555
rect 20570 -1579 20604 -1545
rect 20654 -1615 20688 -1581
rect 20749 -1589 20783 -1555
rect 20853 -1581 20887 -1547
rect 20937 -1615 20971 -1581
rect 21032 -1605 21066 -1571
rect 21136 -1607 21170 -1573
rect 21220 -1541 21254 -1507
rect 21328 -1599 21362 -1565
rect 21412 -1619 21446 -1585
rect 21604 -1615 21638 -1581
rect 21808 -1615 21842 -1581
rect 21912 -1581 21946 -1547
rect 21996 -1555 22030 -1521
rect 22092 -1613 22126 -1579
rect 22176 -1619 22210 -1585
rect 22397 -1615 22431 -1581
rect 22502 -1597 22536 -1563
rect 22586 -1615 22620 -1581
rect 22690 -1589 22724 -1555
rect 22774 -1615 22808 -1581
rect 22858 -1589 22892 -1555
rect 22962 -1579 22996 -1545
rect 23046 -1615 23080 -1581
rect 23141 -1589 23175 -1555
rect 23245 -1581 23279 -1547
rect 23329 -1615 23363 -1581
rect 23424 -1605 23458 -1571
rect 23528 -1607 23562 -1573
rect 23612 -1541 23646 -1507
rect 23720 -1599 23754 -1565
rect 23804 -1619 23838 -1585
rect 23996 -1615 24030 -1581
rect 24200 -1615 24234 -1581
rect 24304 -1581 24338 -1547
rect 24388 -1555 24422 -1521
rect 24484 -1613 24518 -1579
rect 24568 -1619 24602 -1585
rect 24789 -1615 24823 -1581
rect 24894 -1597 24928 -1563
rect 24978 -1615 25012 -1581
rect 25082 -1589 25116 -1555
rect 25166 -1615 25200 -1581
rect 25250 -1589 25284 -1555
<< pdiffc >>
rect 13816 13521 13850 13581
rect 13904 13521 13938 13581
rect 20525 13521 20559 13581
rect 20613 13521 20647 13581
rect 13816 13383 13850 13443
rect 13904 13383 13938 13443
rect 20525 13383 20559 13443
rect 20613 13383 20647 13443
rect 13816 13245 13850 13305
rect 13904 13245 13938 13305
rect 20525 13245 20559 13305
rect 20613 13245 20647 13305
rect 2928 13046 2962 13106
rect 3016 13046 3050 13106
rect 13816 13107 13850 13167
rect 13904 13107 13938 13167
rect 20525 13107 20559 13167
rect 20613 13107 20647 13167
rect 2928 12908 2962 12968
rect 3016 12908 3050 12968
rect 13816 12969 13850 13029
rect 13904 12969 13938 13029
rect 13350 12900 13384 12934
rect 2928 12770 2962 12830
rect 3016 12770 3050 12830
rect 13350 12832 13384 12866
rect 13350 12764 13384 12798
rect 13434 12900 13468 12934
rect 13434 12832 13468 12866
rect 13434 12764 13468 12798
rect 13540 12900 13574 12934
rect 13540 12832 13574 12866
rect 13540 12764 13574 12798
rect 13624 12900 13658 12934
rect 20525 12969 20559 13029
rect 20613 12969 20647 13029
rect 13624 12832 13658 12866
rect 13816 12831 13850 12891
rect 13904 12831 13938 12891
rect 20059 12900 20093 12934
rect 20059 12832 20093 12866
rect 13624 12764 13658 12798
rect 2928 12632 2962 12692
rect 3016 12632 3050 12692
rect 20059 12764 20093 12798
rect 20143 12900 20177 12934
rect 20143 12832 20177 12866
rect 20143 12764 20177 12798
rect 20249 12900 20283 12934
rect 20249 12832 20283 12866
rect 20249 12764 20283 12798
rect 20333 12900 20367 12934
rect 20333 12832 20367 12866
rect 20525 12831 20559 12891
rect 20613 12831 20647 12891
rect 20333 12764 20367 12798
rect 2928 12494 2962 12554
rect 3016 12494 3050 12554
rect 2462 12425 2496 12459
rect 2462 12357 2496 12391
rect 2462 12289 2496 12323
rect 2546 12425 2580 12459
rect 2546 12357 2580 12391
rect 2546 12289 2580 12323
rect 2652 12425 2686 12459
rect 2652 12357 2686 12391
rect 2652 12289 2686 12323
rect 2736 12425 2770 12459
rect 19601 12520 19635 12580
rect 19689 12520 19723 12580
rect 2736 12357 2770 12391
rect 2928 12356 2962 12416
rect 3016 12356 3050 12416
rect 26310 12520 26344 12580
rect 26398 12520 26432 12580
rect 2736 12289 2770 12323
rect 8713 12045 8747 12105
rect 8801 12045 8835 12105
rect 9137 12048 9171 12082
rect 9137 11980 9171 12014
rect 3570 11901 3604 11961
rect 3658 11904 3692 11964
rect 4302 11904 4336 11964
rect 4407 11904 4441 11964
rect 4516 11904 4550 11964
rect 5514 11904 5548 11964
rect 5618 11904 5652 11964
rect 5728 11904 5762 11964
rect 6726 11904 6760 11964
rect 6831 11904 6865 11964
rect 6940 11904 6974 11964
rect 7938 11904 7972 11964
rect 8045 11904 8079 11964
rect 8152 11904 8186 11964
rect 8713 11907 8747 11967
rect 8801 11907 8835 11967
rect 8897 11907 8931 11967
rect 8993 11907 9027 11967
rect 9137 11912 9171 11946
rect 9221 12048 9255 12082
rect 9221 11980 9255 12014
rect 10917 12040 10951 12074
rect 10917 11972 10951 12006
rect 11001 11988 11035 12022
rect 11085 12040 11119 12074
rect 11700 12058 11734 12092
rect 11085 11972 11119 12006
rect 11189 11988 11223 12022
rect 9221 11912 9255 11946
rect 11273 11972 11307 12006
rect 11366 11965 11400 11999
rect 11580 11974 11614 12008
rect 11700 11990 11734 12024
rect 11874 12032 11908 12066
rect 11874 11964 11908 11998
rect 14458 12376 14492 12436
rect 14546 12379 14580 12439
rect 15190 12379 15224 12439
rect 15295 12379 15329 12439
rect 15404 12379 15438 12439
rect 16402 12379 16436 12439
rect 16506 12379 16540 12439
rect 16616 12379 16650 12439
rect 17614 12379 17648 12439
rect 17719 12379 17753 12439
rect 17828 12379 17862 12439
rect 18826 12379 18860 12439
rect 18933 12379 18967 12439
rect 19040 12379 19074 12439
rect 19601 12382 19635 12442
rect 19689 12382 19723 12442
rect 19785 12382 19819 12442
rect 19881 12382 19915 12442
rect 21167 12376 21201 12436
rect 21255 12379 21289 12439
rect 21899 12379 21933 12439
rect 22004 12379 22038 12439
rect 22113 12379 22147 12439
rect 23111 12379 23145 12439
rect 23215 12379 23249 12439
rect 23325 12379 23359 12439
rect 24323 12379 24357 12439
rect 24428 12379 24462 12439
rect 24537 12379 24571 12439
rect 25535 12379 25569 12439
rect 25642 12379 25676 12439
rect 25749 12379 25783 12439
rect 26310 12382 26344 12442
rect 26398 12382 26432 12442
rect 26494 12382 26528 12442
rect 26590 12382 26624 12442
rect 12149 11965 12183 11999
rect 12363 11964 12397 11998
rect 12471 11990 12505 12024
rect 12741 12100 12775 12134
rect 12627 11964 12661 11998
rect 12838 11964 12872 11998
rect 12922 12069 12956 12103
rect 12922 12001 12956 12035
rect 13026 12050 13060 12084
rect 13026 11982 13060 12016
rect 13121 12044 13155 12078
rect 13121 11976 13155 12010
rect 13205 12068 13239 12102
rect 13205 12000 13239 12034
rect 10958 11716 10992 11750
rect 10958 11648 10992 11682
rect 10958 11580 10992 11614
rect 11042 11716 11076 11750
rect 11042 11648 11076 11682
rect 11042 11580 11076 11614
rect 11234 11716 11268 11750
rect 11234 11648 11268 11682
rect 11234 11580 11268 11614
rect 11318 11716 11352 11750
rect 11318 11648 11352 11682
rect 11318 11580 11352 11614
rect 3570 8685 3604 8745
rect 3658 8682 3692 8742
rect 4302 8682 4336 8742
rect 4407 8682 4441 8742
rect 4516 8682 4550 8742
rect 5514 8682 5548 8742
rect 5618 8682 5652 8742
rect 5728 8682 5762 8742
rect 6726 8682 6760 8742
rect 6831 8682 6865 8742
rect 6940 8682 6974 8742
rect 7938 8682 7972 8742
rect 8045 8682 8079 8742
rect 8152 8682 8186 8742
rect 8713 8679 8747 8739
rect 8801 8679 8835 8739
rect 8897 8679 8931 8739
rect 8993 8679 9027 8739
rect 9137 8702 9171 8736
rect 9137 8634 9171 8668
rect 8713 8541 8747 8601
rect 8801 8541 8835 8601
rect 9137 8566 9171 8600
rect 9221 8702 9255 8736
rect 9221 8634 9255 8668
rect 9221 8566 9255 8600
rect 9352 8670 9386 8704
rect 9352 8602 9386 8636
rect 9436 8646 9470 8680
rect 9436 8578 9470 8612
rect 9531 8652 9565 8686
rect 9531 8584 9565 8618
rect 9635 8671 9669 8705
rect 9635 8603 9669 8637
rect 9816 8702 9850 8736
rect 9719 8566 9753 8600
rect 9930 8566 9964 8600
rect 10086 8592 10120 8626
rect 10194 8566 10228 8600
rect 10408 8567 10442 8601
rect 10683 8634 10717 8668
rect 10683 8566 10717 8600
rect 10857 8660 10891 8694
rect 11472 8642 11506 8676
rect 10857 8592 10891 8626
rect 10977 8576 11011 8610
rect 11191 8567 11225 8601
rect 11284 8574 11318 8608
rect 11368 8590 11402 8624
rect 11472 8574 11506 8608
rect 11556 8590 11590 8624
rect 11640 8642 11674 8676
rect 11640 8574 11674 8608
rect 11833 8500 11867 8728
rect 11929 8500 11963 8728
rect 12025 8500 12059 8728
rect 12121 8500 12155 8728
rect 12233 8501 12267 8729
rect 12321 8501 12355 8729
rect 12434 8472 12468 8728
rect 12522 8472 12556 8728
rect 12684 8689 12718 8723
rect 12684 8621 12718 8655
rect 12684 8553 12718 8587
rect 12768 8689 12802 8723
rect 12768 8621 12802 8655
rect 12768 8553 12802 8587
rect 12852 8689 12886 8723
rect 12852 8621 12886 8655
rect 12852 8553 12886 8587
rect 13007 8689 13041 8723
rect 13007 8621 13041 8655
rect 13007 8553 13041 8587
rect 13091 8689 13125 8723
rect 13264 8667 13298 8727
rect 13360 8667 13394 8727
rect 13456 8667 13490 8727
rect 13544 8667 13578 8727
rect 14105 8670 14139 8730
rect 14212 8670 14246 8730
rect 14319 8670 14353 8730
rect 15317 8670 15351 8730
rect 15426 8670 15460 8730
rect 15531 8670 15565 8730
rect 16529 8670 16563 8730
rect 16639 8670 16673 8730
rect 16743 8670 16777 8730
rect 17741 8670 17775 8730
rect 17850 8670 17884 8730
rect 17955 8670 17989 8730
rect 18599 8670 18633 8730
rect 18687 8673 18721 8733
rect 19973 8667 20007 8727
rect 13091 8621 13125 8655
rect 20069 8667 20103 8727
rect 20165 8667 20199 8727
rect 20253 8667 20287 8727
rect 20814 8670 20848 8730
rect 20921 8670 20955 8730
rect 21028 8670 21062 8730
rect 22026 8670 22060 8730
rect 22135 8670 22169 8730
rect 22240 8670 22274 8730
rect 23238 8670 23272 8730
rect 23348 8670 23382 8730
rect 23452 8670 23486 8730
rect 24450 8670 24484 8730
rect 24559 8670 24593 8730
rect 24664 8670 24698 8730
rect 25308 8670 25342 8730
rect 25396 8673 25430 8733
rect 13091 8553 13125 8587
rect 13456 8529 13490 8589
rect 13544 8529 13578 8589
rect 20165 8529 20199 8589
rect 20253 8529 20287 8589
rect 2462 8323 2496 8357
rect 2462 8255 2496 8289
rect 2462 8187 2496 8221
rect 2546 8323 2580 8357
rect 2546 8255 2580 8289
rect 2546 8187 2580 8221
rect 2652 8323 2686 8357
rect 2652 8255 2686 8289
rect 2652 8187 2686 8221
rect 2736 8323 2770 8357
rect 2736 8255 2770 8289
rect 2736 8187 2770 8221
rect 2928 8230 2962 8290
rect 3016 8230 3050 8290
rect 2928 8092 2962 8152
rect 10089 8239 10123 8273
rect 10089 8171 10123 8205
rect 3016 8092 3050 8152
rect 10089 8103 10123 8137
rect 10173 8239 10207 8273
rect 10173 8171 10207 8205
rect 10409 8179 10443 8213
rect 10484 8179 10518 8213
rect 10681 8179 10715 8213
rect 10767 8179 10801 8213
rect 10916 8239 10950 8273
rect 10916 8171 10950 8205
rect 10173 8103 10207 8137
rect 2928 7954 2962 8014
rect 3016 7954 3050 8014
rect 2928 7816 2962 7876
rect 3016 7816 3050 7876
rect 10916 8103 10950 8137
rect 11000 8239 11034 8273
rect 11000 8171 11034 8205
rect 11236 8179 11270 8213
rect 11311 8179 11345 8213
rect 11508 8179 11542 8213
rect 11594 8179 11628 8213
rect 11000 8103 11034 8137
rect 11833 8096 11867 8324
rect 11929 8096 11963 8324
rect 12025 8096 12059 8324
rect 12121 8096 12155 8324
rect 12233 8095 12267 8323
rect 12321 8095 12355 8323
rect 19521 8311 19555 8345
rect 19241 8218 19275 8278
rect 19329 8218 19363 8278
rect 19521 8243 19555 8277
rect 19521 8175 19555 8209
rect 19605 8311 19639 8345
rect 19605 8243 19639 8277
rect 19605 8175 19639 8209
rect 19711 8311 19745 8345
rect 19711 8243 19745 8277
rect 19711 8175 19745 8209
rect 19795 8311 19829 8345
rect 26230 8311 26264 8345
rect 19795 8243 19829 8277
rect 19795 8175 19829 8209
rect 25950 8218 25984 8278
rect 26038 8218 26072 8278
rect 26230 8243 26264 8277
rect 19241 8080 19275 8140
rect 19329 8080 19363 8140
rect 26230 8175 26264 8209
rect 26314 8311 26348 8345
rect 26314 8243 26348 8277
rect 26314 8175 26348 8209
rect 26420 8311 26454 8345
rect 26420 8243 26454 8277
rect 26420 8175 26454 8209
rect 26504 8311 26538 8345
rect 26504 8243 26538 8277
rect 26504 8175 26538 8209
rect 25950 8080 25984 8140
rect 26038 8080 26072 8140
rect 2928 7678 2962 7738
rect 3016 7678 3050 7738
rect 2928 7540 2962 7600
rect 3016 7540 3050 7600
rect 12702 7596 12736 7952
rect 12790 7596 12824 7952
rect 19241 7942 19275 8002
rect 19329 7942 19363 8002
rect 25950 7942 25984 8002
rect 26038 7942 26072 8002
rect 19241 7804 19275 7864
rect 19329 7804 19363 7864
rect 25950 7804 25984 7864
rect 26038 7804 26072 7864
rect 19241 7666 19275 7726
rect 19329 7666 19363 7726
rect 25950 7666 25984 7726
rect 26038 7666 26072 7726
rect 19241 7528 19275 7588
rect 19329 7528 19363 7588
rect 25950 7528 25984 7588
rect 26038 7528 26072 7588
rect 24541 7224 24575 7284
rect 24629 7224 24663 7284
rect 24541 7086 24575 7146
rect 24629 7086 24663 7146
rect 11533 6976 11567 7010
rect 11533 6908 11567 6942
rect 11619 6976 11653 7010
rect 11619 6908 11653 6942
rect 11705 6976 11739 7010
rect 11705 6895 11739 6929
rect 11809 6978 11843 7012
rect 11809 6910 11843 6944
rect 11809 6842 11843 6876
rect 11893 6984 11927 7018
rect 11893 6916 11927 6950
rect 11977 6962 12011 6996
rect 11977 6867 12011 6901
rect 12061 6984 12095 7018
rect 12061 6916 12095 6950
rect 12145 6962 12179 6996
rect 12145 6867 12179 6901
rect 12229 6984 12263 7018
rect 12229 6916 12263 6950
rect 12229 6848 12263 6882
rect 12793 6984 12827 7018
rect 12793 6916 12827 6950
rect 12793 6848 12827 6882
rect 12892 6974 12926 7008
rect 12892 6848 12926 6882
rect 12976 6984 13010 7018
rect 12976 6916 13010 6950
rect 12976 6848 13010 6882
rect 13076 6974 13110 7008
rect 13076 6900 13110 6934
rect 13160 6984 13194 7018
rect 13160 6916 13194 6950
rect 13358 6964 13392 6998
rect 13577 6950 13611 6984
rect 13681 6862 13715 6896
rect 13765 6861 13799 6895
rect 13849 6911 13883 6945
rect 13953 6890 13987 6924
rect 14037 6960 14071 6994
rect 14265 6958 14299 6992
rect 14445 6984 14479 7018
rect 14529 6958 14563 6992
rect 24541 6948 24575 7008
rect 24629 6948 24663 7008
rect 24541 6810 24575 6870
rect 24629 6810 24663 6870
rect 24541 6672 24575 6732
rect 24629 6672 24663 6732
rect 24075 6603 24109 6637
rect 24075 6535 24109 6569
rect 24075 6467 24109 6501
rect 24159 6603 24193 6637
rect 24159 6535 24193 6569
rect 24159 6467 24193 6501
rect 24265 6603 24299 6637
rect 24265 6535 24299 6569
rect 24265 6467 24299 6501
rect 24349 6603 24383 6637
rect 24349 6535 24383 6569
rect 24541 6534 24575 6594
rect 24629 6534 24663 6594
rect 24349 6467 24383 6501
rect 11532 6103 11566 6137
rect 11532 6035 11566 6069
rect 11616 6087 11650 6121
rect 11700 6103 11734 6137
rect 11804 6087 11838 6121
rect 11888 6103 11922 6137
rect 11981 6110 12015 6144
rect 12195 6101 12229 6135
rect 12315 6085 12349 6119
rect 11700 6035 11734 6069
rect 12315 6017 12349 6051
rect 12489 6111 12523 6145
rect 12489 6043 12523 6077
rect 12764 6110 12798 6144
rect 12978 6111 13012 6145
rect 13086 6085 13120 6119
rect 13242 6111 13276 6145
rect 13453 6111 13487 6145
rect 13356 5975 13390 6009
rect 13537 6074 13571 6108
rect 13537 6006 13571 6040
rect 13641 6093 13675 6127
rect 13641 6025 13675 6059
rect 13736 6099 13770 6133
rect 13736 6031 13770 6065
rect 13820 6075 13854 6109
rect 13820 6007 13854 6041
rect 13924 6103 13958 6137
rect 13924 6035 13958 6069
rect 14008 6087 14042 6121
rect 14092 6103 14126 6137
rect 14196 6087 14230 6121
rect 14280 6103 14314 6137
rect 14373 6110 14407 6144
rect 14587 6101 14621 6135
rect 14707 6085 14741 6119
rect 14092 6035 14126 6069
rect 14707 6017 14741 6051
rect 14881 6111 14915 6145
rect 14881 6043 14915 6077
rect 15156 6110 15190 6144
rect 15370 6111 15404 6145
rect 15478 6085 15512 6119
rect 15634 6111 15668 6145
rect 15845 6111 15879 6145
rect 15748 5975 15782 6009
rect 15929 6074 15963 6108
rect 15929 6006 15963 6040
rect 16033 6093 16067 6127
rect 16033 6025 16067 6059
rect 16128 6099 16162 6133
rect 16128 6031 16162 6065
rect 16212 6075 16246 6109
rect 16212 6007 16246 6041
rect 16316 6103 16350 6137
rect 16316 6035 16350 6069
rect 16400 6087 16434 6121
rect 16484 6103 16518 6137
rect 16588 6087 16622 6121
rect 16672 6103 16706 6137
rect 16765 6110 16799 6144
rect 16979 6101 17013 6135
rect 17099 6085 17133 6119
rect 16484 6035 16518 6069
rect 17099 6017 17133 6051
rect 17273 6111 17307 6145
rect 17273 6043 17307 6077
rect 17548 6110 17582 6144
rect 17762 6111 17796 6145
rect 17870 6085 17904 6119
rect 18026 6111 18060 6145
rect 18237 6111 18271 6145
rect 18140 5975 18174 6009
rect 18321 6074 18355 6108
rect 18321 6006 18355 6040
rect 18425 6093 18459 6127
rect 18425 6025 18459 6059
rect 18520 6099 18554 6133
rect 18520 6031 18554 6065
rect 18604 6075 18638 6109
rect 18604 6007 18638 6041
rect 18708 6103 18742 6137
rect 18708 6035 18742 6069
rect 18792 6087 18826 6121
rect 18876 6103 18910 6137
rect 18980 6087 19014 6121
rect 19064 6103 19098 6137
rect 19157 6110 19191 6144
rect 19371 6101 19405 6135
rect 19491 6085 19525 6119
rect 18876 6035 18910 6069
rect 19491 6017 19525 6051
rect 19665 6111 19699 6145
rect 19665 6043 19699 6077
rect 19940 6110 19974 6144
rect 20154 6111 20188 6145
rect 20262 6085 20296 6119
rect 20418 6111 20452 6145
rect 20629 6111 20663 6145
rect 20532 5975 20566 6009
rect 20713 6074 20747 6108
rect 20713 6006 20747 6040
rect 20817 6093 20851 6127
rect 20817 6025 20851 6059
rect 20912 6099 20946 6133
rect 20912 6031 20946 6065
rect 20996 6075 21030 6109
rect 20996 6007 21030 6041
rect 21100 6103 21134 6137
rect 21100 6035 21134 6069
rect 21184 6087 21218 6121
rect 21268 6103 21302 6137
rect 21372 6087 21406 6121
rect 21456 6103 21490 6137
rect 21549 6110 21583 6144
rect 21763 6101 21797 6135
rect 21883 6085 21917 6119
rect 21268 6035 21302 6069
rect 21883 6017 21917 6051
rect 22057 6111 22091 6145
rect 22057 6043 22091 6077
rect 22332 6110 22366 6144
rect 22546 6111 22580 6145
rect 22654 6085 22688 6119
rect 22810 6111 22844 6145
rect 23021 6111 23055 6145
rect 22924 5975 22958 6009
rect 30326 6223 30360 6283
rect 30414 6223 30448 6283
rect 30714 6218 30748 6252
rect 23105 6074 23139 6108
rect 23105 6006 23139 6040
rect 23209 6093 23243 6127
rect 23209 6025 23243 6059
rect 23304 6099 23338 6133
rect 23304 6031 23338 6065
rect 23388 6075 23422 6109
rect 25183 6079 25217 6139
rect 25271 6082 25305 6142
rect 25915 6082 25949 6142
rect 26020 6082 26054 6142
rect 26129 6082 26163 6142
rect 27127 6082 27161 6142
rect 27231 6082 27265 6142
rect 27341 6082 27375 6142
rect 28339 6082 28373 6142
rect 28444 6082 28478 6142
rect 28553 6082 28587 6142
rect 29551 6082 29585 6142
rect 29658 6082 29692 6142
rect 29765 6082 29799 6142
rect 30326 6085 30360 6145
rect 30414 6085 30448 6145
rect 30510 6085 30544 6145
rect 30606 6085 30640 6145
rect 30714 6150 30748 6184
rect 30807 6218 30841 6252
rect 30807 6150 30841 6184
rect 23388 6007 23422 6041
rect 30893 6202 30927 6236
rect 30893 6121 30927 6155
rect 30977 6226 31011 6260
rect 30977 6158 31011 6192
rect 30977 6090 31011 6124
rect 11092 5414 11126 5448
rect 11092 5346 11126 5380
rect 11178 5414 11212 5448
rect 11178 5346 11212 5380
rect 11264 5414 11298 5448
rect 11264 5333 11298 5367
rect 11368 5416 11402 5450
rect 11368 5348 11402 5382
rect 11368 5280 11402 5314
rect 11452 5422 11486 5456
rect 11452 5354 11486 5388
rect 11536 5400 11570 5434
rect 11536 5305 11570 5339
rect 11620 5422 11654 5456
rect 11620 5354 11654 5388
rect 11704 5400 11738 5434
rect 11704 5305 11738 5339
rect 11788 5422 11822 5456
rect 11788 5354 11822 5388
rect 11788 5286 11822 5320
rect 11900 5422 11934 5456
rect 11900 5354 11934 5388
rect 11900 5286 11934 5320
rect 11984 5416 12018 5450
rect 11984 5348 12018 5382
rect 11984 5280 12018 5314
rect 12068 5422 12102 5456
rect 12068 5354 12102 5388
rect 12152 5416 12186 5450
rect 12152 5348 12186 5382
rect 12152 5280 12186 5314
rect 12236 5422 12270 5456
rect 12236 5354 12270 5388
rect 12320 5416 12354 5450
rect 12320 5348 12354 5382
rect 12320 5280 12354 5314
rect 12404 5422 12438 5456
rect 12404 5354 12438 5388
rect 12488 5416 12522 5450
rect 12488 5348 12522 5382
rect 12488 5280 12522 5314
rect 12572 5422 12606 5456
rect 12572 5354 12606 5388
rect 12656 5416 12690 5450
rect 12656 5348 12690 5382
rect 12656 5280 12690 5314
rect 12740 5422 12774 5456
rect 12740 5354 12774 5388
rect 12824 5416 12858 5450
rect 12824 5348 12858 5382
rect 12824 5280 12858 5314
rect 12908 5422 12942 5456
rect 12908 5354 12942 5388
rect 12992 5416 13026 5450
rect 12992 5348 13026 5382
rect 12992 5280 13026 5314
rect 13076 5422 13110 5456
rect 13076 5354 13110 5388
rect 13160 5416 13194 5450
rect 13160 5348 13194 5382
rect 13160 5280 13194 5314
rect 13244 5422 13278 5456
rect 13244 5354 13278 5388
rect 13328 5416 13362 5450
rect 13328 5348 13362 5382
rect 13328 5280 13362 5314
rect 13412 5422 13446 5456
rect 13412 5354 13446 5388
rect 13496 5416 13530 5450
rect 13496 5348 13530 5382
rect 13496 5280 13530 5314
rect 13580 5422 13614 5456
rect 13580 5354 13614 5388
rect 13664 5416 13698 5450
rect 13664 5348 13698 5382
rect 13664 5280 13698 5314
rect 13748 5422 13782 5456
rect 13748 5354 13782 5388
rect 13924 5386 13958 5420
rect 13924 5318 13958 5352
rect 14008 5410 14042 5444
rect 14008 5342 14042 5376
rect 14103 5404 14137 5438
rect 14103 5336 14137 5370
rect 14207 5385 14241 5419
rect 14207 5317 14241 5351
rect 14291 5422 14325 5456
rect 14502 5422 14536 5456
rect 14388 5286 14422 5320
rect 14658 5396 14692 5430
rect 14766 5422 14800 5456
rect 14980 5421 15014 5455
rect 15255 5422 15289 5456
rect 15255 5354 15289 5388
rect 15429 5396 15463 5430
rect 15549 5412 15583 5446
rect 15763 5421 15797 5455
rect 15856 5414 15890 5448
rect 15940 5398 15974 5432
rect 16044 5414 16078 5448
rect 15429 5328 15463 5362
rect 16044 5346 16078 5380
rect 16128 5398 16162 5432
rect 16212 5414 16246 5448
rect 16212 5346 16246 5380
rect 16316 5386 16350 5420
rect 16316 5318 16350 5352
rect 16400 5410 16434 5444
rect 16400 5342 16434 5376
rect 16495 5404 16529 5438
rect 16495 5336 16529 5370
rect 16599 5385 16633 5419
rect 16599 5317 16633 5351
rect 16683 5422 16717 5456
rect 16894 5422 16928 5456
rect 16780 5286 16814 5320
rect 17050 5396 17084 5430
rect 17158 5422 17192 5456
rect 17372 5421 17406 5455
rect 17647 5422 17681 5456
rect 17647 5354 17681 5388
rect 17821 5396 17855 5430
rect 17941 5412 17975 5446
rect 18155 5421 18189 5455
rect 18248 5414 18282 5448
rect 18332 5398 18366 5432
rect 18436 5414 18470 5448
rect 17821 5328 17855 5362
rect 18436 5346 18470 5380
rect 18520 5398 18554 5432
rect 18604 5414 18638 5448
rect 18604 5346 18638 5380
rect 18708 5386 18742 5420
rect 18708 5318 18742 5352
rect 18792 5410 18826 5444
rect 18792 5342 18826 5376
rect 18887 5404 18921 5438
rect 18887 5336 18921 5370
rect 18991 5385 19025 5419
rect 18991 5317 19025 5351
rect 19075 5422 19109 5456
rect 19286 5422 19320 5456
rect 19172 5286 19206 5320
rect 19442 5396 19476 5430
rect 19550 5422 19584 5456
rect 19764 5421 19798 5455
rect 20039 5422 20073 5456
rect 20039 5354 20073 5388
rect 20213 5396 20247 5430
rect 20333 5412 20367 5446
rect 20547 5421 20581 5455
rect 20640 5414 20674 5448
rect 20724 5398 20758 5432
rect 20828 5414 20862 5448
rect 20213 5328 20247 5362
rect 20828 5346 20862 5380
rect 20912 5398 20946 5432
rect 20996 5414 21030 5448
rect 20996 5346 21030 5380
rect 21100 5386 21134 5420
rect 21100 5318 21134 5352
rect 21184 5410 21218 5444
rect 21184 5342 21218 5376
rect 21279 5404 21313 5438
rect 21279 5336 21313 5370
rect 21383 5385 21417 5419
rect 21383 5317 21417 5351
rect 21467 5422 21501 5456
rect 21678 5422 21712 5456
rect 21564 5286 21598 5320
rect 21834 5396 21868 5430
rect 21942 5422 21976 5456
rect 22156 5421 22190 5455
rect 22431 5422 22465 5456
rect 22431 5354 22465 5388
rect 22605 5396 22639 5430
rect 22725 5412 22759 5446
rect 22939 5421 22973 5455
rect 23032 5414 23066 5448
rect 23116 5398 23150 5432
rect 23220 5414 23254 5448
rect 22605 5328 22639 5362
rect 23220 5346 23254 5380
rect 23304 5398 23338 5432
rect 23388 5414 23422 5448
rect 23388 5346 23422 5380
rect 11124 4540 11158 4574
rect 11124 4472 11158 4506
rect 11210 4540 11244 4574
rect 11210 4472 11244 4506
rect 11296 4540 11330 4574
rect 11296 4459 11330 4493
rect 11400 4542 11434 4576
rect 11400 4474 11434 4508
rect 11400 4406 11434 4440
rect 11484 4548 11518 4582
rect 11484 4480 11518 4514
rect 11568 4526 11602 4560
rect 11568 4431 11602 4465
rect 11652 4548 11686 4582
rect 11652 4480 11686 4514
rect 11736 4526 11770 4560
rect 11736 4431 11770 4465
rect 11820 4548 11854 4582
rect 11820 4480 11854 4514
rect 11820 4412 11854 4446
rect 13707 4549 13741 4583
rect 13707 4481 13741 4515
rect 13707 4413 13741 4447
rect 13791 4549 13825 4583
rect 13791 4481 13825 4515
rect 13923 4541 13957 4575
rect 13923 4473 13957 4507
rect 14007 4525 14041 4559
rect 14091 4541 14125 4575
rect 14195 4525 14229 4559
rect 14279 4541 14313 4575
rect 14372 4548 14406 4582
rect 14586 4539 14620 4573
rect 14706 4523 14740 4557
rect 14091 4473 14125 4507
rect 13791 4413 13825 4447
rect 14706 4455 14740 4489
rect 14880 4549 14914 4583
rect 14880 4481 14914 4515
rect 15155 4548 15189 4582
rect 15369 4549 15403 4583
rect 15477 4523 15511 4557
rect 15633 4549 15667 4583
rect 15844 4549 15878 4583
rect 15747 4413 15781 4447
rect 15928 4512 15962 4546
rect 15928 4444 15962 4478
rect 16032 4531 16066 4565
rect 16032 4463 16066 4497
rect 16127 4537 16161 4571
rect 16127 4469 16161 4503
rect 16211 4513 16245 4547
rect 16211 4445 16245 4479
rect 16315 4541 16349 4575
rect 16315 4473 16349 4507
rect 16399 4525 16433 4559
rect 16483 4541 16517 4575
rect 16587 4525 16621 4559
rect 16671 4541 16705 4575
rect 16764 4548 16798 4582
rect 16978 4539 17012 4573
rect 17098 4523 17132 4557
rect 16483 4473 16517 4507
rect 17098 4455 17132 4489
rect 17272 4549 17306 4583
rect 17272 4481 17306 4515
rect 17547 4548 17581 4582
rect 17761 4549 17795 4583
rect 17869 4523 17903 4557
rect 18025 4549 18059 4583
rect 18236 4549 18270 4583
rect 18139 4413 18173 4447
rect 18320 4512 18354 4546
rect 18320 4444 18354 4478
rect 18424 4531 18458 4565
rect 18424 4463 18458 4497
rect 18519 4537 18553 4571
rect 18519 4469 18553 4503
rect 18603 4513 18637 4547
rect 18603 4445 18637 4479
rect 18707 4541 18741 4575
rect 18707 4473 18741 4507
rect 18791 4525 18825 4559
rect 18875 4541 18909 4575
rect 18979 4525 19013 4559
rect 19063 4541 19097 4575
rect 19156 4548 19190 4582
rect 19370 4539 19404 4573
rect 19490 4523 19524 4557
rect 18875 4473 18909 4507
rect 19490 4455 19524 4489
rect 19664 4549 19698 4583
rect 19664 4481 19698 4515
rect 19939 4548 19973 4582
rect 20153 4549 20187 4583
rect 20261 4523 20295 4557
rect 20417 4549 20451 4583
rect 20628 4549 20662 4583
rect 20531 4413 20565 4447
rect 20712 4512 20746 4546
rect 20712 4444 20746 4478
rect 20816 4531 20850 4565
rect 20816 4463 20850 4497
rect 20911 4537 20945 4571
rect 20911 4469 20945 4503
rect 20995 4513 21029 4547
rect 20995 4445 21029 4479
rect 21099 4541 21133 4575
rect 21099 4473 21133 4507
rect 21183 4525 21217 4559
rect 21267 4541 21301 4575
rect 21371 4525 21405 4559
rect 21455 4541 21489 4575
rect 21548 4548 21582 4582
rect 21762 4539 21796 4573
rect 21882 4523 21916 4557
rect 21267 4473 21301 4507
rect 21882 4455 21916 4489
rect 22056 4549 22090 4583
rect 22056 4481 22090 4515
rect 22331 4548 22365 4582
rect 22545 4549 22579 4583
rect 22653 4523 22687 4557
rect 22809 4549 22843 4583
rect 23020 4549 23054 4583
rect 22923 4413 22957 4447
rect 23104 4512 23138 4546
rect 23104 4444 23138 4478
rect 23208 4531 23242 4565
rect 23208 4463 23242 4497
rect 23303 4537 23337 4571
rect 23303 4469 23337 4503
rect 23387 4513 23421 4547
rect 23387 4445 23421 4479
rect 25612 3872 25646 3906
rect 25612 3804 25646 3838
rect 25696 3820 25730 3854
rect 25780 3872 25814 3906
rect 26395 3890 26429 3924
rect 25780 3804 25814 3838
rect 25884 3820 25918 3854
rect 25968 3804 26002 3838
rect 26061 3797 26095 3831
rect 26275 3806 26309 3840
rect 26395 3822 26429 3856
rect 26569 3864 26603 3898
rect 26569 3796 26603 3830
rect 26844 3797 26878 3831
rect 27058 3796 27092 3830
rect 27166 3822 27200 3856
rect 27436 3932 27470 3966
rect 27322 3796 27356 3830
rect 27533 3796 27567 3830
rect 27617 3901 27651 3935
rect 27617 3833 27651 3867
rect 27721 3882 27755 3916
rect 27721 3814 27755 3848
rect 27816 3876 27850 3910
rect 27816 3808 27850 3842
rect 27900 3900 27934 3934
rect 27900 3832 27934 3866
rect 28004 3872 28038 3906
rect 28004 3804 28038 3838
rect 28088 3820 28122 3854
rect 28172 3872 28206 3906
rect 28787 3890 28821 3924
rect 28172 3804 28206 3838
rect 28276 3820 28310 3854
rect 28360 3804 28394 3838
rect 28453 3797 28487 3831
rect 28667 3806 28701 3840
rect 28787 3822 28821 3856
rect 28961 3864 28995 3898
rect 28961 3796 28995 3830
rect 29236 3797 29270 3831
rect 29450 3796 29484 3830
rect 29558 3822 29592 3856
rect 29828 3932 29862 3966
rect 29714 3796 29748 3830
rect 29925 3796 29959 3830
rect 30009 3901 30043 3935
rect 30009 3833 30043 3867
rect 30113 3882 30147 3916
rect 30113 3814 30147 3848
rect 30208 3876 30242 3910
rect 30208 3808 30242 3842
rect 30292 3900 30326 3934
rect 30292 3832 30326 3866
rect 11531 3640 11565 3674
rect 11531 3572 11565 3606
rect 11615 3664 11649 3698
rect 11615 3596 11649 3630
rect 11710 3658 11744 3692
rect 11710 3590 11744 3624
rect 11814 3639 11848 3673
rect 11814 3571 11848 3605
rect 11898 3676 11932 3710
rect 12109 3676 12143 3710
rect 11995 3540 12029 3574
rect 12265 3650 12299 3684
rect 12373 3676 12407 3710
rect 12587 3675 12621 3709
rect 12862 3676 12896 3710
rect 12862 3608 12896 3642
rect 13036 3650 13070 3684
rect 13156 3666 13190 3700
rect 13370 3675 13404 3709
rect 13463 3668 13497 3702
rect 13547 3652 13581 3686
rect 13651 3668 13685 3702
rect 13036 3582 13070 3616
rect 13651 3600 13685 3634
rect 13735 3652 13769 3686
rect 13819 3668 13853 3702
rect 13819 3600 13853 3634
rect 13923 3640 13957 3674
rect 13923 3572 13957 3606
rect 14007 3664 14041 3698
rect 14007 3596 14041 3630
rect 14102 3658 14136 3692
rect 14102 3590 14136 3624
rect 14206 3639 14240 3673
rect 14206 3571 14240 3605
rect 14290 3676 14324 3710
rect 14501 3676 14535 3710
rect 14387 3540 14421 3574
rect 14657 3650 14691 3684
rect 14765 3676 14799 3710
rect 14979 3675 15013 3709
rect 15254 3676 15288 3710
rect 15254 3608 15288 3642
rect 15428 3650 15462 3684
rect 15548 3666 15582 3700
rect 15762 3675 15796 3709
rect 15855 3668 15889 3702
rect 15939 3652 15973 3686
rect 16043 3668 16077 3702
rect 15428 3582 15462 3616
rect 16043 3600 16077 3634
rect 16127 3652 16161 3686
rect 16211 3668 16245 3702
rect 16211 3600 16245 3634
rect 16315 3640 16349 3674
rect 16315 3572 16349 3606
rect 16399 3664 16433 3698
rect 16399 3596 16433 3630
rect 16494 3658 16528 3692
rect 16494 3590 16528 3624
rect 16598 3639 16632 3673
rect 16598 3571 16632 3605
rect 16682 3676 16716 3710
rect 16893 3676 16927 3710
rect 16779 3540 16813 3574
rect 17049 3650 17083 3684
rect 17157 3676 17191 3710
rect 17371 3675 17405 3709
rect 17646 3676 17680 3710
rect 17646 3608 17680 3642
rect 17820 3650 17854 3684
rect 17940 3666 17974 3700
rect 18154 3675 18188 3709
rect 18247 3668 18281 3702
rect 18331 3652 18365 3686
rect 18435 3668 18469 3702
rect 17820 3582 17854 3616
rect 18435 3600 18469 3634
rect 18519 3652 18553 3686
rect 18603 3668 18637 3702
rect 18603 3600 18637 3634
rect 18707 3640 18741 3674
rect 18707 3572 18741 3606
rect 18791 3664 18825 3698
rect 18791 3596 18825 3630
rect 18886 3658 18920 3692
rect 18886 3590 18920 3624
rect 18990 3639 19024 3673
rect 18990 3571 19024 3605
rect 19074 3676 19108 3710
rect 19285 3676 19319 3710
rect 19171 3540 19205 3574
rect 19441 3650 19475 3684
rect 19549 3676 19583 3710
rect 19763 3675 19797 3709
rect 20038 3676 20072 3710
rect 20038 3608 20072 3642
rect 20212 3650 20246 3684
rect 20332 3666 20366 3700
rect 20546 3675 20580 3709
rect 20639 3668 20673 3702
rect 20723 3652 20757 3686
rect 20827 3668 20861 3702
rect 20212 3582 20246 3616
rect 20827 3600 20861 3634
rect 20911 3652 20945 3686
rect 20995 3668 21029 3702
rect 20995 3600 21029 3634
rect 21099 3640 21133 3674
rect 21099 3572 21133 3606
rect 21183 3664 21217 3698
rect 21183 3596 21217 3630
rect 21278 3658 21312 3692
rect 21278 3590 21312 3624
rect 21382 3639 21416 3673
rect 21382 3571 21416 3605
rect 21466 3676 21500 3710
rect 21677 3676 21711 3710
rect 21563 3540 21597 3574
rect 21833 3650 21867 3684
rect 21941 3676 21975 3710
rect 22155 3675 22189 3709
rect 22430 3676 22464 3710
rect 22430 3608 22464 3642
rect 22604 3650 22638 3684
rect 22724 3666 22758 3700
rect 22938 3675 22972 3709
rect 23031 3668 23065 3702
rect 23115 3652 23149 3686
rect 23219 3668 23253 3702
rect 22604 3582 22638 3616
rect 23219 3600 23253 3634
rect 23303 3652 23337 3686
rect 23387 3668 23421 3702
rect 23387 3600 23421 3634
rect 25612 3540 25646 3574
rect 25612 3472 25646 3506
rect 25696 3524 25730 3558
rect 25780 3540 25814 3574
rect 25884 3524 25918 3558
rect 25968 3540 26002 3574
rect 26061 3547 26095 3581
rect 26275 3538 26309 3572
rect 26395 3522 26429 3556
rect 25780 3472 25814 3506
rect 26395 3454 26429 3488
rect 26569 3548 26603 3582
rect 26569 3480 26603 3514
rect 26844 3547 26878 3581
rect 27058 3548 27092 3582
rect 27166 3522 27200 3556
rect 27322 3548 27356 3582
rect 27533 3548 27567 3582
rect 27436 3412 27470 3446
rect 27617 3511 27651 3545
rect 27617 3443 27651 3477
rect 27721 3530 27755 3564
rect 27721 3462 27755 3496
rect 27816 3536 27850 3570
rect 27816 3468 27850 3502
rect 27900 3512 27934 3546
rect 27900 3444 27934 3478
rect 28004 3540 28038 3574
rect 28004 3472 28038 3506
rect 28088 3524 28122 3558
rect 28172 3540 28206 3574
rect 28276 3524 28310 3558
rect 28360 3540 28394 3574
rect 28453 3547 28487 3581
rect 28667 3538 28701 3572
rect 28787 3522 28821 3556
rect 28172 3472 28206 3506
rect 28787 3454 28821 3488
rect 28961 3548 28995 3582
rect 28961 3480 28995 3514
rect 29236 3547 29270 3581
rect 29450 3548 29484 3582
rect 29558 3522 29592 3556
rect 29714 3548 29748 3582
rect 29925 3548 29959 3582
rect 29828 3412 29862 3446
rect 30009 3511 30043 3545
rect 30009 3443 30043 3477
rect 30113 3530 30147 3564
rect 30113 3462 30147 3496
rect 30208 3536 30242 3570
rect 30208 3468 30242 3502
rect 30292 3512 30326 3546
rect 30292 3444 30326 3478
rect 25612 2592 25646 2626
rect 25612 2524 25646 2558
rect 25696 2540 25730 2574
rect 25780 2592 25814 2626
rect 26395 2610 26429 2644
rect 25780 2524 25814 2558
rect 25884 2540 25918 2574
rect 25968 2524 26002 2558
rect 26061 2517 26095 2551
rect 26275 2526 26309 2560
rect 26395 2542 26429 2576
rect 26569 2584 26603 2618
rect 26569 2516 26603 2550
rect 26844 2517 26878 2551
rect 27058 2516 27092 2550
rect 27166 2542 27200 2576
rect 27436 2652 27470 2686
rect 27322 2516 27356 2550
rect 27533 2516 27567 2550
rect 27617 2621 27651 2655
rect 27617 2553 27651 2587
rect 27721 2602 27755 2636
rect 27721 2534 27755 2568
rect 27816 2596 27850 2630
rect 27816 2528 27850 2562
rect 27900 2620 27934 2654
rect 27900 2552 27934 2586
rect 28004 2592 28038 2626
rect 28004 2524 28038 2558
rect 28088 2540 28122 2574
rect 28172 2592 28206 2626
rect 28787 2610 28821 2644
rect 28172 2524 28206 2558
rect 28276 2540 28310 2574
rect 28360 2524 28394 2558
rect 28453 2517 28487 2551
rect 28667 2526 28701 2560
rect 28787 2542 28821 2576
rect 28961 2584 28995 2618
rect 28961 2516 28995 2550
rect 29236 2517 29270 2551
rect 29450 2516 29484 2550
rect 29558 2542 29592 2576
rect 29828 2652 29862 2686
rect 29714 2516 29748 2550
rect 29925 2516 29959 2550
rect 30009 2621 30043 2655
rect 30009 2553 30043 2587
rect 30113 2602 30147 2636
rect 30113 2534 30147 2568
rect 30208 2596 30242 2630
rect 30208 2528 30242 2562
rect 30292 2620 30326 2654
rect 30292 2552 30326 2586
rect 25612 2260 25646 2294
rect 25612 2192 25646 2226
rect 25696 2244 25730 2278
rect 25780 2260 25814 2294
rect 25884 2244 25918 2278
rect 25968 2260 26002 2294
rect 26061 2267 26095 2301
rect 26275 2258 26309 2292
rect 26395 2242 26429 2276
rect 25780 2192 25814 2226
rect 26395 2174 26429 2208
rect 26569 2268 26603 2302
rect 26569 2200 26603 2234
rect 26844 2267 26878 2301
rect 27058 2268 27092 2302
rect 27166 2242 27200 2276
rect 27322 2268 27356 2302
rect 27533 2268 27567 2302
rect 27436 2132 27470 2166
rect 27617 2231 27651 2265
rect 27617 2163 27651 2197
rect 27721 2250 27755 2284
rect 27721 2182 27755 2216
rect 27816 2256 27850 2290
rect 27816 2188 27850 2222
rect 27900 2232 27934 2266
rect 27900 2164 27934 2198
rect 28004 2260 28038 2294
rect 28004 2192 28038 2226
rect 28088 2244 28122 2278
rect 28172 2260 28206 2294
rect 28276 2244 28310 2278
rect 28360 2260 28394 2294
rect 28453 2267 28487 2301
rect 28667 2258 28701 2292
rect 28787 2242 28821 2276
rect 28172 2192 28206 2226
rect 28787 2174 28821 2208
rect 28961 2268 28995 2302
rect 28961 2200 28995 2234
rect 29236 2267 29270 2301
rect 29450 2268 29484 2302
rect 29558 2242 29592 2276
rect 29714 2268 29748 2302
rect 29925 2268 29959 2302
rect 29828 2132 29862 2166
rect 30009 2231 30043 2265
rect 30009 2163 30043 2197
rect 30113 2250 30147 2284
rect 30113 2182 30147 2216
rect 30208 2256 30242 2290
rect 30208 2188 30242 2222
rect 30292 2232 30326 2266
rect 30292 2164 30326 2198
rect 8612 1288 8646 1322
rect 8612 1220 8646 1254
rect 8698 1288 8732 1322
rect 8698 1220 8732 1254
rect 8784 1288 8818 1322
rect 8784 1207 8818 1241
rect 8888 1290 8922 1324
rect 8888 1222 8922 1256
rect 8888 1154 8922 1188
rect 8972 1296 9006 1330
rect 8972 1228 9006 1262
rect 9056 1274 9090 1308
rect 9056 1179 9090 1213
rect 9140 1296 9174 1330
rect 9140 1228 9174 1262
rect 9224 1274 9258 1308
rect 9224 1179 9258 1213
rect 9308 1296 9342 1330
rect 9308 1228 9342 1262
rect 9308 1160 9342 1194
rect 9440 1296 9474 1330
rect 9440 1228 9474 1262
rect 9440 1160 9474 1194
rect 9524 1290 9558 1324
rect 9524 1222 9558 1256
rect 9524 1154 9558 1188
rect 9608 1296 9642 1330
rect 9608 1228 9642 1262
rect 9692 1290 9726 1324
rect 9692 1222 9726 1256
rect 9692 1154 9726 1188
rect 9776 1296 9810 1330
rect 9776 1228 9810 1262
rect 9860 1290 9894 1324
rect 9860 1222 9894 1256
rect 9860 1154 9894 1188
rect 9944 1296 9978 1330
rect 9944 1228 9978 1262
rect 10028 1290 10062 1324
rect 10028 1222 10062 1256
rect 10028 1154 10062 1188
rect 10112 1296 10146 1330
rect 10112 1228 10146 1262
rect 10196 1290 10230 1324
rect 10196 1222 10230 1256
rect 10196 1154 10230 1188
rect 10280 1296 10314 1330
rect 10280 1228 10314 1262
rect 10364 1290 10398 1324
rect 10364 1222 10398 1256
rect 10364 1154 10398 1188
rect 10448 1296 10482 1330
rect 10448 1228 10482 1262
rect 10532 1290 10566 1324
rect 10532 1222 10566 1256
rect 10532 1154 10566 1188
rect 10616 1296 10650 1330
rect 10616 1228 10650 1262
rect 10700 1290 10734 1324
rect 10700 1222 10734 1256
rect 10700 1154 10734 1188
rect 10784 1296 10818 1330
rect 10784 1228 10818 1262
rect 10868 1290 10902 1324
rect 10868 1222 10902 1256
rect 10868 1154 10902 1188
rect 10952 1296 10986 1330
rect 10952 1228 10986 1262
rect 11036 1290 11070 1324
rect 11036 1222 11070 1256
rect 11036 1154 11070 1188
rect 11120 1296 11154 1330
rect 11120 1228 11154 1262
rect 11204 1290 11238 1324
rect 11204 1222 11238 1256
rect 11204 1154 11238 1188
rect 11288 1296 11322 1330
rect 11288 1228 11322 1262
rect 12996 1288 13030 1322
rect 12996 1220 13030 1254
rect 13082 1288 13116 1322
rect 13082 1220 13116 1254
rect 13168 1288 13202 1322
rect 13168 1207 13202 1241
rect 13272 1290 13306 1324
rect 13272 1222 13306 1256
rect 13272 1154 13306 1188
rect 13356 1296 13390 1330
rect 13356 1228 13390 1262
rect 13440 1274 13474 1308
rect 13440 1179 13474 1213
rect 13524 1296 13558 1330
rect 13524 1228 13558 1262
rect 13608 1274 13642 1308
rect 13608 1179 13642 1213
rect 13692 1296 13726 1330
rect 13692 1228 13726 1262
rect 13692 1160 13726 1194
rect 13824 1296 13858 1330
rect 13824 1228 13858 1262
rect 13824 1160 13858 1194
rect 13908 1290 13942 1324
rect 13908 1222 13942 1256
rect 13908 1154 13942 1188
rect 13992 1296 14026 1330
rect 13992 1228 14026 1262
rect 14076 1290 14110 1324
rect 14076 1222 14110 1256
rect 14076 1154 14110 1188
rect 14160 1296 14194 1330
rect 14160 1228 14194 1262
rect 14244 1290 14278 1324
rect 14244 1222 14278 1256
rect 14244 1154 14278 1188
rect 14328 1296 14362 1330
rect 14328 1228 14362 1262
rect 14412 1290 14446 1324
rect 14412 1222 14446 1256
rect 14412 1154 14446 1188
rect 14496 1296 14530 1330
rect 14496 1228 14530 1262
rect 14580 1290 14614 1324
rect 14580 1222 14614 1256
rect 14580 1154 14614 1188
rect 14664 1296 14698 1330
rect 14664 1228 14698 1262
rect 14748 1290 14782 1324
rect 14748 1222 14782 1256
rect 14748 1154 14782 1188
rect 14832 1296 14866 1330
rect 14832 1228 14866 1262
rect 14916 1290 14950 1324
rect 14916 1222 14950 1256
rect 14916 1154 14950 1188
rect 15000 1296 15034 1330
rect 15000 1228 15034 1262
rect 15084 1290 15118 1324
rect 15084 1222 15118 1256
rect 15084 1154 15118 1188
rect 15168 1296 15202 1330
rect 15168 1228 15202 1262
rect 15252 1290 15286 1324
rect 15252 1222 15286 1256
rect 15252 1154 15286 1188
rect 15336 1296 15370 1330
rect 15336 1228 15370 1262
rect 15420 1290 15454 1324
rect 15420 1222 15454 1256
rect 15420 1154 15454 1188
rect 15504 1296 15538 1330
rect 15504 1228 15538 1262
rect 15588 1290 15622 1324
rect 15588 1222 15622 1256
rect 15588 1154 15622 1188
rect 15672 1296 15706 1330
rect 15672 1228 15706 1262
rect 8610 154 8644 188
rect 8610 86 8644 120
rect 8610 18 8644 52
rect 8694 154 8728 188
rect 8694 86 8728 120
rect 8930 94 8964 128
rect 9005 94 9039 128
rect 9202 94 9236 128
rect 9288 94 9322 128
rect 10090 94 10124 128
rect 10176 94 10210 128
rect 10373 94 10407 128
rect 10448 94 10482 128
rect 10684 154 10718 188
rect 10684 86 10718 120
rect 8694 18 8728 52
rect 10684 18 10718 52
rect 10768 154 10802 188
rect 10768 86 10802 120
rect 10768 18 10802 52
rect 11002 154 11036 188
rect 11002 86 11036 120
rect 11002 18 11036 52
rect 11086 154 11120 188
rect 11086 86 11120 120
rect 11322 94 11356 128
rect 11397 94 11431 128
rect 11594 94 11628 128
rect 11680 94 11714 128
rect 12482 94 12516 128
rect 12568 94 12602 128
rect 12765 94 12799 128
rect 12840 94 12874 128
rect 13076 154 13110 188
rect 13076 86 13110 120
rect 11086 18 11120 52
rect 13076 18 13110 52
rect 13160 154 13194 188
rect 13160 86 13194 120
rect 13160 18 13194 52
rect 13394 154 13428 188
rect 13394 86 13428 120
rect 13394 18 13428 52
rect 13478 154 13512 188
rect 13478 86 13512 120
rect 13714 94 13748 128
rect 13789 94 13823 128
rect 13986 94 14020 128
rect 14072 94 14106 128
rect 14872 94 14906 128
rect 14958 94 14992 128
rect 15155 94 15189 128
rect 15230 94 15264 128
rect 15466 154 15500 188
rect 15466 86 15500 120
rect 13478 18 13512 52
rect 15466 18 15500 52
rect 15550 154 15584 188
rect 15550 86 15584 120
rect 15550 18 15584 52
rect 15786 154 15820 188
rect 15786 86 15820 120
rect 15786 18 15820 52
rect 15870 154 15904 188
rect 15870 86 15904 120
rect 16106 94 16140 128
rect 16181 94 16215 128
rect 16378 94 16412 128
rect 16464 94 16498 128
rect 17266 94 17300 128
rect 17352 94 17386 128
rect 17549 94 17583 128
rect 17624 94 17658 128
rect 17860 154 17894 188
rect 17860 86 17894 120
rect 15870 18 15904 52
rect 17860 18 17894 52
rect 17944 154 17978 188
rect 17944 86 17978 120
rect 17944 18 17978 52
rect 18178 154 18212 188
rect 18178 86 18212 120
rect 18178 18 18212 52
rect 18262 154 18296 188
rect 18262 86 18296 120
rect 18498 94 18532 128
rect 18573 94 18607 128
rect 18770 94 18804 128
rect 18856 94 18890 128
rect 19658 94 19692 128
rect 19744 94 19778 128
rect 19941 94 19975 128
rect 20016 94 20050 128
rect 20252 154 20286 188
rect 20252 86 20286 120
rect 18262 18 18296 52
rect 20252 18 20286 52
rect 20336 154 20370 188
rect 20336 86 20370 120
rect 20336 18 20370 52
rect 20570 154 20604 188
rect 20570 86 20604 120
rect 20570 18 20604 52
rect 20654 154 20688 188
rect 20654 86 20688 120
rect 20890 94 20924 128
rect 20965 94 20999 128
rect 21162 94 21196 128
rect 21248 94 21282 128
rect 22048 94 22082 128
rect 22134 94 22168 128
rect 22331 94 22365 128
rect 22406 94 22440 128
rect 22642 154 22676 188
rect 22642 86 22676 120
rect 20654 18 20688 52
rect 22642 18 22676 52
rect 22726 154 22760 188
rect 22726 86 22760 120
rect 22726 18 22760 52
rect 22962 154 22996 188
rect 22962 86 22996 120
rect 22962 18 22996 52
rect 23046 154 23080 188
rect 23046 86 23080 120
rect 23282 94 23316 128
rect 23357 94 23391 128
rect 23554 94 23588 128
rect 23640 94 23674 128
rect 24442 94 24476 128
rect 24528 94 24562 128
rect 24725 94 24759 128
rect 24800 94 24834 128
rect 25036 154 25070 188
rect 25036 86 25070 120
rect 23046 18 23080 52
rect 25036 18 25070 52
rect 25120 154 25154 188
rect 25120 86 25154 120
rect 25120 18 25154 52
rect 8610 -542 8644 -508
rect 8610 -610 8644 -576
rect 8694 -558 8728 -524
rect 8778 -542 8812 -508
rect 8882 -558 8916 -524
rect 8966 -542 9000 -508
rect 9058 -535 9092 -501
rect 9272 -544 9306 -510
rect 9392 -560 9426 -526
rect 8778 -610 8812 -576
rect 9392 -628 9426 -594
rect 9566 -534 9600 -500
rect 9566 -602 9600 -568
rect 9841 -535 9875 -501
rect 10055 -534 10089 -500
rect 10163 -560 10197 -526
rect 10329 -534 10363 -500
rect 10531 -534 10565 -500
rect 10433 -670 10467 -636
rect 10615 -571 10649 -537
rect 10615 -639 10649 -605
rect 10719 -552 10753 -518
rect 10719 -620 10753 -586
rect 10814 -546 10848 -512
rect 10814 -614 10848 -580
rect 10898 -570 10932 -536
rect 10898 -638 10932 -604
rect 11002 -542 11036 -508
rect 11002 -610 11036 -576
rect 11086 -558 11120 -524
rect 11170 -542 11204 -508
rect 11274 -558 11308 -524
rect 11358 -542 11392 -508
rect 11450 -535 11484 -501
rect 11664 -544 11698 -510
rect 11784 -560 11818 -526
rect 11170 -610 11204 -576
rect 11784 -628 11818 -594
rect 11958 -534 11992 -500
rect 11958 -602 11992 -568
rect 12233 -535 12267 -501
rect 12447 -534 12481 -500
rect 12555 -560 12589 -526
rect 12721 -534 12755 -500
rect 12923 -534 12957 -500
rect 12825 -670 12859 -636
rect 13007 -571 13041 -537
rect 13007 -639 13041 -605
rect 13111 -552 13145 -518
rect 13111 -620 13145 -586
rect 13206 -546 13240 -512
rect 13206 -614 13240 -580
rect 13290 -570 13324 -536
rect 13290 -638 13324 -604
rect 13394 -542 13428 -508
rect 13394 -610 13428 -576
rect 13478 -558 13512 -524
rect 13562 -542 13596 -508
rect 13666 -558 13700 -524
rect 13750 -542 13784 -508
rect 13842 -535 13876 -501
rect 14056 -544 14090 -510
rect 14176 -560 14210 -526
rect 13562 -610 13596 -576
rect 14176 -628 14210 -594
rect 14350 -534 14384 -500
rect 14350 -602 14384 -568
rect 14625 -535 14659 -501
rect 14839 -534 14873 -500
rect 14947 -560 14981 -526
rect 15113 -534 15147 -500
rect 15315 -534 15349 -500
rect 15217 -670 15251 -636
rect 15399 -571 15433 -537
rect 15399 -639 15433 -605
rect 15503 -552 15537 -518
rect 15503 -620 15537 -586
rect 15598 -546 15632 -512
rect 15598 -614 15632 -580
rect 15682 -570 15716 -536
rect 15682 -638 15716 -604
rect 15786 -542 15820 -508
rect 15786 -610 15820 -576
rect 15870 -558 15904 -524
rect 15954 -542 15988 -508
rect 16058 -558 16092 -524
rect 16142 -542 16176 -508
rect 16234 -535 16268 -501
rect 16448 -544 16482 -510
rect 16568 -560 16602 -526
rect 15954 -610 15988 -576
rect 16568 -628 16602 -594
rect 16742 -534 16776 -500
rect 16742 -602 16776 -568
rect 17017 -535 17051 -501
rect 17231 -534 17265 -500
rect 17339 -560 17373 -526
rect 17505 -534 17539 -500
rect 17707 -534 17741 -500
rect 17609 -670 17643 -636
rect 17791 -571 17825 -537
rect 17791 -639 17825 -605
rect 17895 -552 17929 -518
rect 17895 -620 17929 -586
rect 17990 -546 18024 -512
rect 17990 -614 18024 -580
rect 18074 -570 18108 -536
rect 18074 -638 18108 -604
rect 18178 -542 18212 -508
rect 18178 -610 18212 -576
rect 18262 -558 18296 -524
rect 18346 -542 18380 -508
rect 18450 -558 18484 -524
rect 18534 -542 18568 -508
rect 18626 -535 18660 -501
rect 18840 -544 18874 -510
rect 18960 -560 18994 -526
rect 18346 -610 18380 -576
rect 18960 -628 18994 -594
rect 19134 -534 19168 -500
rect 19134 -602 19168 -568
rect 19409 -535 19443 -501
rect 19623 -534 19657 -500
rect 19731 -560 19765 -526
rect 19897 -534 19931 -500
rect 20099 -534 20133 -500
rect 20001 -670 20035 -636
rect 20183 -571 20217 -537
rect 20183 -639 20217 -605
rect 20287 -552 20321 -518
rect 20287 -620 20321 -586
rect 20382 -546 20416 -512
rect 20382 -614 20416 -580
rect 20466 -570 20500 -536
rect 20466 -638 20500 -604
rect 20570 -542 20604 -508
rect 20570 -610 20604 -576
rect 20654 -558 20688 -524
rect 20738 -542 20772 -508
rect 20842 -558 20876 -524
rect 20926 -542 20960 -508
rect 21018 -535 21052 -501
rect 21232 -544 21266 -510
rect 21352 -560 21386 -526
rect 20738 -610 20772 -576
rect 21352 -628 21386 -594
rect 21526 -534 21560 -500
rect 21526 -602 21560 -568
rect 21801 -535 21835 -501
rect 22015 -534 22049 -500
rect 22123 -560 22157 -526
rect 22289 -534 22323 -500
rect 22491 -534 22525 -500
rect 22393 -670 22427 -636
rect 22575 -571 22609 -537
rect 22575 -639 22609 -605
rect 22679 -552 22713 -518
rect 22679 -620 22713 -586
rect 22774 -546 22808 -512
rect 22774 -614 22808 -580
rect 22858 -570 22892 -536
rect 22858 -638 22892 -604
rect 22962 -542 22996 -508
rect 22962 -610 22996 -576
rect 23046 -558 23080 -524
rect 23130 -542 23164 -508
rect 23234 -558 23268 -524
rect 23318 -542 23352 -508
rect 23410 -535 23444 -501
rect 23624 -544 23658 -510
rect 23744 -560 23778 -526
rect 23130 -610 23164 -576
rect 23744 -628 23778 -594
rect 23918 -534 23952 -500
rect 23918 -602 23952 -568
rect 24193 -535 24227 -501
rect 24407 -534 24441 -500
rect 24515 -560 24549 -526
rect 24681 -534 24715 -500
rect 24883 -534 24917 -500
rect 24785 -670 24819 -636
rect 24967 -571 25001 -537
rect 24967 -639 25001 -605
rect 25071 -552 25105 -518
rect 25071 -620 25105 -586
rect 25166 -546 25200 -512
rect 25166 -614 25200 -580
rect 25250 -570 25284 -536
rect 25250 -638 25284 -604
rect 8610 -1259 8644 -1225
rect 8610 -1327 8644 -1293
rect 8694 -1235 8728 -1201
rect 8694 -1303 8728 -1269
rect 8789 -1241 8823 -1207
rect 8789 -1309 8823 -1275
rect 8893 -1260 8927 -1226
rect 8893 -1328 8927 -1294
rect 8977 -1223 9011 -1189
rect 9179 -1223 9213 -1189
rect 9075 -1359 9109 -1325
rect 9345 -1249 9379 -1215
rect 9453 -1223 9487 -1189
rect 9667 -1224 9701 -1190
rect 9942 -1223 9976 -1189
rect 9942 -1291 9976 -1257
rect 10116 -1249 10150 -1215
rect 10236 -1233 10270 -1199
rect 10450 -1224 10484 -1190
rect 10542 -1231 10576 -1197
rect 10626 -1247 10660 -1213
rect 10730 -1231 10764 -1197
rect 10116 -1317 10150 -1283
rect 10730 -1299 10764 -1265
rect 10814 -1247 10848 -1213
rect 10898 -1231 10932 -1197
rect 10898 -1299 10932 -1265
rect 11002 -1259 11036 -1225
rect 11002 -1327 11036 -1293
rect 11086 -1235 11120 -1201
rect 11086 -1303 11120 -1269
rect 11181 -1241 11215 -1207
rect 11181 -1309 11215 -1275
rect 11285 -1260 11319 -1226
rect 11285 -1328 11319 -1294
rect 11369 -1223 11403 -1189
rect 11571 -1223 11605 -1189
rect 11467 -1359 11501 -1325
rect 11737 -1249 11771 -1215
rect 11845 -1223 11879 -1189
rect 12059 -1224 12093 -1190
rect 12334 -1223 12368 -1189
rect 12334 -1291 12368 -1257
rect 12508 -1249 12542 -1215
rect 12628 -1233 12662 -1199
rect 12842 -1224 12876 -1190
rect 12934 -1231 12968 -1197
rect 13018 -1247 13052 -1213
rect 13122 -1231 13156 -1197
rect 12508 -1317 12542 -1283
rect 13122 -1299 13156 -1265
rect 13206 -1247 13240 -1213
rect 13290 -1231 13324 -1197
rect 13290 -1299 13324 -1265
rect 13394 -1259 13428 -1225
rect 13394 -1327 13428 -1293
rect 13478 -1235 13512 -1201
rect 13478 -1303 13512 -1269
rect 13573 -1241 13607 -1207
rect 13573 -1309 13607 -1275
rect 13677 -1260 13711 -1226
rect 13677 -1328 13711 -1294
rect 13761 -1223 13795 -1189
rect 13963 -1223 13997 -1189
rect 13859 -1359 13893 -1325
rect 14129 -1249 14163 -1215
rect 14237 -1223 14271 -1189
rect 14451 -1224 14485 -1190
rect 14726 -1223 14760 -1189
rect 14726 -1291 14760 -1257
rect 14900 -1249 14934 -1215
rect 15020 -1233 15054 -1199
rect 15234 -1224 15268 -1190
rect 15326 -1231 15360 -1197
rect 15410 -1247 15444 -1213
rect 15514 -1231 15548 -1197
rect 14900 -1317 14934 -1283
rect 15514 -1299 15548 -1265
rect 15598 -1247 15632 -1213
rect 15682 -1231 15716 -1197
rect 15682 -1299 15716 -1265
rect 15786 -1259 15820 -1225
rect 15786 -1327 15820 -1293
rect 15870 -1235 15904 -1201
rect 15870 -1303 15904 -1269
rect 15965 -1241 15999 -1207
rect 15965 -1309 15999 -1275
rect 16069 -1260 16103 -1226
rect 16069 -1328 16103 -1294
rect 16153 -1223 16187 -1189
rect 16355 -1223 16389 -1189
rect 16251 -1359 16285 -1325
rect 16521 -1249 16555 -1215
rect 16629 -1223 16663 -1189
rect 16843 -1224 16877 -1190
rect 17118 -1223 17152 -1189
rect 17118 -1291 17152 -1257
rect 17292 -1249 17326 -1215
rect 17412 -1233 17446 -1199
rect 17626 -1224 17660 -1190
rect 17718 -1231 17752 -1197
rect 17802 -1247 17836 -1213
rect 17906 -1231 17940 -1197
rect 17292 -1317 17326 -1283
rect 17906 -1299 17940 -1265
rect 17990 -1247 18024 -1213
rect 18074 -1231 18108 -1197
rect 18074 -1299 18108 -1265
rect 18178 -1259 18212 -1225
rect 18178 -1327 18212 -1293
rect 18262 -1235 18296 -1201
rect 18262 -1303 18296 -1269
rect 18357 -1241 18391 -1207
rect 18357 -1309 18391 -1275
rect 18461 -1260 18495 -1226
rect 18461 -1328 18495 -1294
rect 18545 -1223 18579 -1189
rect 18747 -1223 18781 -1189
rect 18643 -1359 18677 -1325
rect 18913 -1249 18947 -1215
rect 19021 -1223 19055 -1189
rect 19235 -1224 19269 -1190
rect 19510 -1223 19544 -1189
rect 19510 -1291 19544 -1257
rect 19684 -1249 19718 -1215
rect 19804 -1233 19838 -1199
rect 20018 -1224 20052 -1190
rect 20110 -1231 20144 -1197
rect 20194 -1247 20228 -1213
rect 20298 -1231 20332 -1197
rect 19684 -1317 19718 -1283
rect 20298 -1299 20332 -1265
rect 20382 -1247 20416 -1213
rect 20466 -1231 20500 -1197
rect 20466 -1299 20500 -1265
rect 20570 -1259 20604 -1225
rect 20570 -1327 20604 -1293
rect 20654 -1235 20688 -1201
rect 20654 -1303 20688 -1269
rect 20749 -1241 20783 -1207
rect 20749 -1309 20783 -1275
rect 20853 -1260 20887 -1226
rect 20853 -1328 20887 -1294
rect 20937 -1223 20971 -1189
rect 21139 -1223 21173 -1189
rect 21035 -1359 21069 -1325
rect 21305 -1249 21339 -1215
rect 21413 -1223 21447 -1189
rect 21627 -1224 21661 -1190
rect 21902 -1223 21936 -1189
rect 21902 -1291 21936 -1257
rect 22076 -1249 22110 -1215
rect 22196 -1233 22230 -1199
rect 22410 -1224 22444 -1190
rect 22502 -1231 22536 -1197
rect 22586 -1247 22620 -1213
rect 22690 -1231 22724 -1197
rect 22076 -1317 22110 -1283
rect 22690 -1299 22724 -1265
rect 22774 -1247 22808 -1213
rect 22858 -1231 22892 -1197
rect 22858 -1299 22892 -1265
rect 22962 -1259 22996 -1225
rect 22962 -1327 22996 -1293
rect 23046 -1235 23080 -1201
rect 23046 -1303 23080 -1269
rect 23141 -1241 23175 -1207
rect 23141 -1309 23175 -1275
rect 23245 -1260 23279 -1226
rect 23245 -1328 23279 -1294
rect 23329 -1223 23363 -1189
rect 23531 -1223 23565 -1189
rect 23427 -1359 23461 -1325
rect 23697 -1249 23731 -1215
rect 23805 -1223 23839 -1189
rect 24019 -1224 24053 -1190
rect 24294 -1223 24328 -1189
rect 24294 -1291 24328 -1257
rect 24468 -1249 24502 -1215
rect 24588 -1233 24622 -1199
rect 24802 -1224 24836 -1190
rect 24894 -1231 24928 -1197
rect 24978 -1247 25012 -1213
rect 25082 -1231 25116 -1197
rect 24468 -1317 24502 -1283
rect 25082 -1299 25116 -1265
rect 25166 -1247 25200 -1213
rect 25250 -1231 25284 -1197
rect 25250 -1299 25284 -1265
<< psubdiff >>
rect 10882 12466 10911 12500
rect 10945 12466 11003 12500
rect 11037 12466 11095 12500
rect 11129 12466 11187 12500
rect 11221 12466 11279 12500
rect 11313 12466 11371 12500
rect 11405 12466 11463 12500
rect 11497 12466 11555 12500
rect 11589 12466 11647 12500
rect 11681 12466 11739 12500
rect 11773 12466 11831 12500
rect 11865 12466 11923 12500
rect 11957 12466 12015 12500
rect 12049 12466 12107 12500
rect 12141 12466 12199 12500
rect 12233 12466 12291 12500
rect 12325 12466 12383 12500
rect 12417 12466 12475 12500
rect 12509 12466 12567 12500
rect 12601 12466 12659 12500
rect 12693 12466 12751 12500
rect 12785 12466 12843 12500
rect 12877 12466 12935 12500
rect 12969 12466 13027 12500
rect 13061 12466 13119 12500
rect 13153 12466 13211 12500
rect 13245 12466 13274 12500
rect 13344 12403 13368 12437
rect 13402 12403 13486 12437
rect 13520 12403 13630 12437
rect 13664 12403 13706 12437
rect 2456 11928 2480 11962
rect 2514 11928 2598 11962
rect 2632 11928 2742 11962
rect 2776 11928 2818 11962
rect 2456 11926 2818 11928
rect 13344 12401 13706 12403
rect 20053 12403 20077 12437
rect 20111 12403 20195 12437
rect 20229 12403 20339 12437
rect 20373 12403 20415 12437
rect 20053 12401 20415 12403
rect 9061 11572 9336 11581
rect 9061 11538 9091 11572
rect 9125 11538 9183 11572
rect 9217 11570 9336 11572
rect 9217 11538 9277 11570
rect 9061 11536 9277 11538
rect 9311 11536 9336 11570
rect 13288 11596 13406 11616
rect 9061 11531 9336 11536
rect 13288 11539 13315 11596
rect 13381 11539 13406 11596
rect 13288 11517 13406 11539
rect 10882 11214 10911 11248
rect 10945 11214 11003 11248
rect 11037 11214 11095 11248
rect 11129 11214 11187 11248
rect 11221 11214 11279 11248
rect 11313 11214 11371 11248
rect 11405 11214 11434 11248
rect 14068 11212 14172 11247
rect 14068 11178 14099 11212
rect 14133 11178 14172 11212
rect 14068 11149 14172 11178
rect 20777 11212 20881 11247
rect 20777 11178 20808 11212
rect 20842 11178 20881 11212
rect 20777 11149 20881 11178
rect 14466 11041 14798 11057
rect 14466 11007 14492 11041
rect 14526 11007 14572 11041
rect 14606 11007 14652 11041
rect 14686 11007 14732 11041
rect 14766 11007 14798 11041
rect 14466 10989 14798 11007
rect 15198 11041 15530 11057
rect 15198 11007 15224 11041
rect 15258 11007 15304 11041
rect 15338 11007 15384 11041
rect 15418 11007 15464 11041
rect 15498 11007 15530 11041
rect 15198 10989 15530 11007
rect 15800 11041 16132 11057
rect 15800 11007 15832 11041
rect 15866 11007 15912 11041
rect 15946 11007 15992 11041
rect 16026 11007 16072 11041
rect 16106 11007 16132 11041
rect 15800 10989 16132 11007
rect 16410 11041 16742 11057
rect 16410 11007 16436 11041
rect 16470 11007 16516 11041
rect 16550 11007 16596 11041
rect 16630 11007 16676 11041
rect 16710 11007 16742 11041
rect 16410 10989 16742 11007
rect 17012 11041 17344 11057
rect 17012 11007 17044 11041
rect 17078 11007 17124 11041
rect 17158 11007 17204 11041
rect 17238 11007 17284 11041
rect 17318 11007 17344 11041
rect 17012 10989 17344 11007
rect 17748 11041 18080 11057
rect 17748 11007 17774 11041
rect 17808 11007 17854 11041
rect 17888 11007 17934 11041
rect 17968 11007 18014 11041
rect 18048 11007 18080 11041
rect 17748 10989 18080 11007
rect 18350 11041 18682 11057
rect 18350 11007 18382 11041
rect 18416 11007 18462 11041
rect 18496 11007 18542 11041
rect 18576 11007 18622 11041
rect 18656 11007 18682 11041
rect 18350 10989 18682 11007
rect 19084 11041 19416 11057
rect 19084 11007 19116 11041
rect 19150 11007 19196 11041
rect 19230 11007 19276 11041
rect 19310 11007 19356 11041
rect 19390 11007 19416 11041
rect 21175 11041 21507 11057
rect 19084 10989 19416 11007
rect 21175 11007 21201 11041
rect 21235 11007 21281 11041
rect 21315 11007 21361 11041
rect 21395 11007 21441 11041
rect 21475 11007 21507 11041
rect 21175 10989 21507 11007
rect 21907 11041 22239 11057
rect 21907 11007 21933 11041
rect 21967 11007 22013 11041
rect 22047 11007 22093 11041
rect 22127 11007 22173 11041
rect 22207 11007 22239 11041
rect 21907 10989 22239 11007
rect 22509 11041 22841 11057
rect 22509 11007 22541 11041
rect 22575 11007 22621 11041
rect 22655 11007 22701 11041
rect 22735 11007 22781 11041
rect 22815 11007 22841 11041
rect 22509 10989 22841 11007
rect 23119 11041 23451 11057
rect 23119 11007 23145 11041
rect 23179 11007 23225 11041
rect 23259 11007 23305 11041
rect 23339 11007 23385 11041
rect 23419 11007 23451 11041
rect 23119 10989 23451 11007
rect 23721 11041 24053 11057
rect 23721 11007 23753 11041
rect 23787 11007 23833 11041
rect 23867 11007 23913 11041
rect 23947 11007 23993 11041
rect 24027 11007 24053 11041
rect 23721 10989 24053 11007
rect 24457 11041 24789 11057
rect 24457 11007 24483 11041
rect 24517 11007 24563 11041
rect 24597 11007 24643 11041
rect 24677 11007 24723 11041
rect 24757 11007 24789 11041
rect 24457 10989 24789 11007
rect 25059 11041 25391 11057
rect 25059 11007 25091 11041
rect 25125 11007 25171 11041
rect 25205 11007 25251 11041
rect 25285 11007 25331 11041
rect 25365 11007 25391 11041
rect 25059 10989 25391 11007
rect 25793 11041 26125 11057
rect 25793 11007 25825 11041
rect 25859 11007 25905 11041
rect 25939 11007 25985 11041
rect 26019 11007 26065 11041
rect 26099 11007 26125 11041
rect 25793 10989 26125 11007
rect 3180 10737 3284 10772
rect 3180 10703 3211 10737
rect 3245 10703 3284 10737
rect 3180 10674 3284 10703
rect 3578 10566 3910 10582
rect 3578 10532 3604 10566
rect 3638 10532 3684 10566
rect 3718 10532 3764 10566
rect 3798 10532 3844 10566
rect 3878 10532 3910 10566
rect 3578 10514 3910 10532
rect 4310 10566 4642 10582
rect 4310 10532 4336 10566
rect 4370 10532 4416 10566
rect 4450 10532 4496 10566
rect 4530 10532 4576 10566
rect 4610 10532 4642 10566
rect 4310 10514 4642 10532
rect 4912 10566 5244 10582
rect 4912 10532 4944 10566
rect 4978 10532 5024 10566
rect 5058 10532 5104 10566
rect 5138 10532 5184 10566
rect 5218 10532 5244 10566
rect 4912 10514 5244 10532
rect 5522 10566 5854 10582
rect 5522 10532 5548 10566
rect 5582 10532 5628 10566
rect 5662 10532 5708 10566
rect 5742 10532 5788 10566
rect 5822 10532 5854 10566
rect 5522 10514 5854 10532
rect 6124 10566 6456 10582
rect 6124 10532 6156 10566
rect 6190 10532 6236 10566
rect 6270 10532 6316 10566
rect 6350 10532 6396 10566
rect 6430 10532 6456 10566
rect 6124 10514 6456 10532
rect 6860 10566 7192 10582
rect 6860 10532 6886 10566
rect 6920 10532 6966 10566
rect 7000 10532 7046 10566
rect 7080 10532 7126 10566
rect 7160 10532 7192 10566
rect 6860 10514 7192 10532
rect 7462 10566 7794 10582
rect 7462 10532 7494 10566
rect 7528 10532 7574 10566
rect 7608 10532 7654 10566
rect 7688 10532 7734 10566
rect 7768 10532 7794 10566
rect 7462 10514 7794 10532
rect 8196 10566 8528 10582
rect 8196 10532 8228 10566
rect 8262 10532 8308 10566
rect 8342 10532 8388 10566
rect 8422 10532 8468 10566
rect 8502 10532 8528 10566
rect 8196 10514 8528 10532
rect 3578 10114 3910 10132
rect 3578 10080 3604 10114
rect 3638 10080 3684 10114
rect 3718 10080 3764 10114
rect 3798 10080 3844 10114
rect 3878 10080 3910 10114
rect 3578 10064 3910 10080
rect 4310 10114 4642 10132
rect 4310 10080 4336 10114
rect 4370 10080 4416 10114
rect 4450 10080 4496 10114
rect 4530 10080 4576 10114
rect 4610 10080 4642 10114
rect 4310 10064 4642 10080
rect 4912 10114 5244 10132
rect 4912 10080 4944 10114
rect 4978 10080 5024 10114
rect 5058 10080 5104 10114
rect 5138 10080 5184 10114
rect 5218 10080 5244 10114
rect 4912 10064 5244 10080
rect 5522 10114 5854 10132
rect 5522 10080 5548 10114
rect 5582 10080 5628 10114
rect 5662 10080 5708 10114
rect 5742 10080 5788 10114
rect 5822 10080 5854 10114
rect 5522 10064 5854 10080
rect 6124 10114 6456 10132
rect 6124 10080 6156 10114
rect 6190 10080 6236 10114
rect 6270 10080 6316 10114
rect 6350 10080 6396 10114
rect 6430 10080 6456 10114
rect 6124 10064 6456 10080
rect 6860 10114 7192 10132
rect 6860 10080 6886 10114
rect 6920 10080 6966 10114
rect 7000 10080 7046 10114
rect 7080 10080 7126 10114
rect 7160 10080 7192 10114
rect 6860 10064 7192 10080
rect 7462 10114 7794 10132
rect 7462 10080 7494 10114
rect 7528 10080 7574 10114
rect 7608 10080 7654 10114
rect 7688 10080 7734 10114
rect 7768 10080 7794 10114
rect 7462 10064 7794 10080
rect 8196 10114 8528 10132
rect 8196 10080 8228 10114
rect 8262 10080 8308 10114
rect 8342 10080 8388 10114
rect 8422 10080 8468 10114
rect 8502 10080 8528 10114
rect 8196 10064 8528 10080
rect 13763 10102 14095 10120
rect 13763 10068 13789 10102
rect 13823 10068 13869 10102
rect 13903 10068 13949 10102
rect 13983 10068 14029 10102
rect 14063 10068 14095 10102
rect 13763 10052 14095 10068
rect 14497 10102 14829 10120
rect 14497 10068 14523 10102
rect 14557 10068 14603 10102
rect 14637 10068 14683 10102
rect 14717 10068 14763 10102
rect 14797 10068 14829 10102
rect 14497 10052 14829 10068
rect 15099 10102 15431 10120
rect 15099 10068 15131 10102
rect 15165 10068 15211 10102
rect 15245 10068 15291 10102
rect 15325 10068 15371 10102
rect 15405 10068 15431 10102
rect 15099 10052 15431 10068
rect 15835 10102 16167 10120
rect 15835 10068 15861 10102
rect 15895 10068 15941 10102
rect 15975 10068 16021 10102
rect 16055 10068 16101 10102
rect 16135 10068 16167 10102
rect 15835 10052 16167 10068
rect 16437 10102 16769 10120
rect 16437 10068 16469 10102
rect 16503 10068 16549 10102
rect 16583 10068 16629 10102
rect 16663 10068 16709 10102
rect 16743 10068 16769 10102
rect 16437 10052 16769 10068
rect 17047 10102 17379 10120
rect 17047 10068 17073 10102
rect 17107 10068 17153 10102
rect 17187 10068 17233 10102
rect 17267 10068 17313 10102
rect 17347 10068 17379 10102
rect 17047 10052 17379 10068
rect 17649 10102 17981 10120
rect 17649 10068 17681 10102
rect 17715 10068 17761 10102
rect 17795 10068 17841 10102
rect 17875 10068 17921 10102
rect 17955 10068 17981 10102
rect 17649 10052 17981 10068
rect 18381 10102 18713 10120
rect 18381 10068 18413 10102
rect 18447 10068 18493 10102
rect 18527 10068 18573 10102
rect 18607 10068 18653 10102
rect 18687 10068 18713 10102
rect 20472 10102 20804 10120
rect 18381 10052 18713 10068
rect 20472 10068 20498 10102
rect 20532 10068 20578 10102
rect 20612 10068 20658 10102
rect 20692 10068 20738 10102
rect 20772 10068 20804 10102
rect 20472 10052 20804 10068
rect 21206 10102 21538 10120
rect 21206 10068 21232 10102
rect 21266 10068 21312 10102
rect 21346 10068 21392 10102
rect 21426 10068 21472 10102
rect 21506 10068 21538 10102
rect 21206 10052 21538 10068
rect 21808 10102 22140 10120
rect 21808 10068 21840 10102
rect 21874 10068 21920 10102
rect 21954 10068 22000 10102
rect 22034 10068 22080 10102
rect 22114 10068 22140 10102
rect 21808 10052 22140 10068
rect 22544 10102 22876 10120
rect 22544 10068 22570 10102
rect 22604 10068 22650 10102
rect 22684 10068 22730 10102
rect 22764 10068 22810 10102
rect 22844 10068 22876 10102
rect 22544 10052 22876 10068
rect 23146 10102 23478 10120
rect 23146 10068 23178 10102
rect 23212 10068 23258 10102
rect 23292 10068 23338 10102
rect 23372 10068 23418 10102
rect 23452 10068 23478 10102
rect 23146 10052 23478 10068
rect 23756 10102 24088 10120
rect 23756 10068 23782 10102
rect 23816 10068 23862 10102
rect 23896 10068 23942 10102
rect 23976 10068 24022 10102
rect 24056 10068 24088 10102
rect 23756 10052 24088 10068
rect 24358 10102 24690 10120
rect 24358 10068 24390 10102
rect 24424 10068 24470 10102
rect 24504 10068 24550 10102
rect 24584 10068 24630 10102
rect 24664 10068 24690 10102
rect 24358 10052 24690 10068
rect 25090 10102 25422 10120
rect 25090 10068 25122 10102
rect 25156 10068 25202 10102
rect 25236 10068 25282 10102
rect 25316 10068 25362 10102
rect 25396 10068 25422 10102
rect 25090 10052 25422 10068
rect 3180 9943 3284 9972
rect 3180 9909 3211 9943
rect 3245 9909 3284 9943
rect 3180 9874 3284 9909
rect 19007 9931 19111 9960
rect 19007 9897 19046 9931
rect 19080 9897 19111 9931
rect 19007 9862 19111 9897
rect 25716 9931 25820 9960
rect 25716 9897 25755 9931
rect 25789 9897 25820 9931
rect 25716 9862 25820 9897
rect 9061 9103 11710 9106
rect 9061 9102 9898 9103
rect 9061 9068 9090 9102
rect 9124 9068 9182 9102
rect 9216 9068 9274 9102
rect 9308 9068 9346 9102
rect 9380 9101 9530 9102
rect 9380 9068 9438 9101
rect 9061 9067 9438 9068
rect 9472 9068 9530 9101
rect 9564 9068 9714 9102
rect 9748 9068 9806 9102
rect 9840 9069 9898 9102
rect 9932 9102 11710 9103
rect 9932 9069 9990 9102
rect 9840 9068 9990 9069
rect 10024 9101 10174 9102
rect 10024 9068 10082 9101
rect 9472 9067 10082 9068
rect 10116 9068 10174 9101
rect 10208 9068 10266 9102
rect 10300 9068 10358 9102
rect 10392 9068 10450 9102
rect 10484 9068 10542 9102
rect 10576 9068 10634 9102
rect 10668 9068 10726 9102
rect 10760 9068 10818 9102
rect 10852 9101 11002 9102
rect 10852 9068 10910 9101
rect 10116 9067 10910 9068
rect 10944 9068 11002 9101
rect 11036 9068 11094 9102
rect 11128 9068 11278 9102
rect 11312 9068 11370 9102
rect 11404 9068 11462 9102
rect 11496 9068 11554 9102
rect 11588 9101 11710 9102
rect 11588 9068 11646 9101
rect 10944 9067 11646 9068
rect 11680 9067 11710 9101
rect 2456 8718 2818 8720
rect 2456 8684 2480 8718
rect 2514 8684 2598 8718
rect 2632 8684 2742 8718
rect 2776 8684 2818 8718
rect 19473 8706 19835 8708
rect 19473 8672 19515 8706
rect 19549 8672 19659 8706
rect 19693 8672 19777 8706
rect 19811 8672 19835 8706
rect 26182 8706 26544 8708
rect 26182 8672 26224 8706
rect 26258 8672 26368 8706
rect 26402 8672 26486 8706
rect 26520 8672 26544 8706
rect 10054 7771 10534 7773
rect 10054 7737 10083 7771
rect 10117 7737 10175 7771
rect 10209 7737 10267 7771
rect 10301 7737 10359 7771
rect 10393 7737 10451 7771
rect 10485 7737 10534 7771
rect 10054 7734 10534 7737
rect 10668 7737 10727 7771
rect 10761 7770 10910 7771
rect 10761 7737 10819 7770
rect 10668 7736 10819 7737
rect 10853 7737 10910 7770
rect 10944 7737 11002 7771
rect 11036 7737 11095 7771
rect 11129 7737 11186 7771
rect 11220 7737 11278 7771
rect 11312 7737 11336 7771
rect 10853 7736 11336 7737
rect 10668 7732 11336 7736
rect 11494 7736 11554 7770
rect 11588 7736 11646 7770
rect 11680 7736 11707 7770
rect 11494 7732 11707 7736
rect 11498 6492 11527 6526
rect 11561 6492 11619 6526
rect 11653 6492 11711 6526
rect 11745 6492 11803 6526
rect 11837 6492 11895 6526
rect 11929 6492 11987 6526
rect 12021 6492 12079 6526
rect 12113 6492 12171 6526
rect 12205 6492 12263 6526
rect 12297 6492 12355 6526
rect 12389 6492 12447 6526
rect 12481 6492 12539 6526
rect 12573 6492 12631 6526
rect 12665 6492 12723 6526
rect 12757 6492 12815 6526
rect 12849 6492 12907 6526
rect 12941 6492 12999 6526
rect 13033 6492 13091 6526
rect 13125 6492 13183 6526
rect 13217 6492 13275 6526
rect 13309 6492 13367 6526
rect 13401 6492 13459 6526
rect 13493 6492 13551 6526
rect 13585 6492 13643 6526
rect 13677 6492 13735 6526
rect 13769 6492 13827 6526
rect 13861 6492 13919 6526
rect 13953 6492 14011 6526
rect 14045 6492 14103 6526
rect 14137 6492 14195 6526
rect 14229 6492 14287 6526
rect 14321 6492 14379 6526
rect 14413 6492 14471 6526
rect 14505 6492 14598 6526
rect 24069 6106 24093 6140
rect 24127 6106 24211 6140
rect 24245 6106 24355 6140
rect 24389 6106 24431 6140
rect 24069 6104 24431 6106
rect 30680 5757 30800 5758
rect 30680 5723 30708 5757
rect 30742 5724 30800 5757
rect 30834 5724 30892 5758
rect 30926 5724 30985 5758
rect 31019 5724 31049 5758
rect 30742 5723 31049 5724
rect 30680 5722 31049 5723
rect 11497 5619 11526 5653
rect 11560 5619 11618 5653
rect 11652 5619 11710 5653
rect 11744 5619 11802 5653
rect 11836 5619 11894 5653
rect 11928 5619 11986 5653
rect 12020 5619 12078 5653
rect 12112 5619 12170 5653
rect 12204 5619 12262 5653
rect 12296 5619 12354 5653
rect 12388 5619 12446 5653
rect 12480 5619 12538 5653
rect 12572 5619 12630 5653
rect 12664 5619 12722 5653
rect 12756 5619 12814 5653
rect 12848 5619 12906 5653
rect 12940 5619 12998 5653
rect 13032 5619 13090 5653
rect 13124 5619 13182 5653
rect 13216 5619 13274 5653
rect 13308 5619 13366 5653
rect 13400 5619 13458 5653
rect 13492 5619 13550 5653
rect 13584 5619 13642 5653
rect 13676 5619 13734 5653
rect 13768 5619 13826 5653
rect 13860 5619 13918 5653
rect 13952 5619 14010 5653
rect 14044 5619 14102 5653
rect 14136 5619 14194 5653
rect 14228 5619 14286 5653
rect 14320 5619 14378 5653
rect 14412 5619 14470 5653
rect 14504 5619 14562 5653
rect 14596 5619 14654 5653
rect 14688 5619 14746 5653
rect 14780 5619 14838 5653
rect 14872 5619 14930 5653
rect 14964 5619 15022 5653
rect 15056 5619 15114 5653
rect 15148 5619 15206 5653
rect 15240 5619 15298 5653
rect 15332 5619 15390 5653
rect 15424 5619 15482 5653
rect 15516 5619 15574 5653
rect 15608 5619 15666 5653
rect 15700 5619 15758 5653
rect 15792 5619 15850 5653
rect 15884 5619 15942 5653
rect 15976 5619 16034 5653
rect 16068 5619 16126 5653
rect 16160 5619 16218 5653
rect 16252 5619 16310 5653
rect 16344 5619 16402 5653
rect 16436 5619 16494 5653
rect 16528 5619 16586 5653
rect 16620 5619 16678 5653
rect 16712 5619 16770 5653
rect 16804 5619 16862 5653
rect 16896 5619 16954 5653
rect 16988 5619 17046 5653
rect 17080 5619 17138 5653
rect 17172 5619 17230 5653
rect 17264 5619 17322 5653
rect 17356 5619 17414 5653
rect 17448 5619 17506 5653
rect 17540 5619 17598 5653
rect 17632 5619 17690 5653
rect 17724 5619 17782 5653
rect 17816 5619 17874 5653
rect 17908 5619 17966 5653
rect 18000 5619 18058 5653
rect 18092 5619 18150 5653
rect 18184 5619 18242 5653
rect 18276 5619 18334 5653
rect 18368 5619 18426 5653
rect 18460 5619 18518 5653
rect 18552 5619 18610 5653
rect 18644 5619 18702 5653
rect 18736 5619 18794 5653
rect 18828 5619 18886 5653
rect 18920 5619 18978 5653
rect 19012 5619 19070 5653
rect 19104 5619 19162 5653
rect 19196 5619 19254 5653
rect 19288 5619 19346 5653
rect 19380 5619 19438 5653
rect 19472 5619 19530 5653
rect 19564 5619 19622 5653
rect 19656 5619 19714 5653
rect 19748 5619 19806 5653
rect 19840 5619 19898 5653
rect 19932 5619 19990 5653
rect 20024 5619 20082 5653
rect 20116 5619 20174 5653
rect 20208 5619 20266 5653
rect 20300 5619 20358 5653
rect 20392 5619 20450 5653
rect 20484 5619 20542 5653
rect 20576 5619 20634 5653
rect 20668 5619 20726 5653
rect 20760 5619 20818 5653
rect 20852 5619 20910 5653
rect 20944 5619 21002 5653
rect 21036 5619 21094 5653
rect 21128 5619 21186 5653
rect 21220 5619 21278 5653
rect 21312 5619 21370 5653
rect 21404 5619 21462 5653
rect 21496 5619 21554 5653
rect 21588 5619 21646 5653
rect 21680 5619 21738 5653
rect 21772 5619 21830 5653
rect 21864 5619 21922 5653
rect 21956 5619 22014 5653
rect 22048 5619 22106 5653
rect 22140 5619 22198 5653
rect 22232 5619 22290 5653
rect 22324 5619 22382 5653
rect 22416 5619 22474 5653
rect 22508 5619 22566 5653
rect 22600 5619 22658 5653
rect 22692 5619 22750 5653
rect 22784 5619 22842 5653
rect 22876 5619 22934 5653
rect 22968 5619 23026 5653
rect 23060 5619 23118 5653
rect 23152 5619 23210 5653
rect 23244 5619 23302 5653
rect 23336 5619 23394 5653
rect 23428 5619 23457 5653
rect 11057 4930 11086 4964
rect 11120 4930 11178 4964
rect 11212 4930 11270 4964
rect 11304 4930 11362 4964
rect 11396 4930 11454 4964
rect 11488 4930 11546 4964
rect 11580 4930 11638 4964
rect 11672 4930 11730 4964
rect 11764 4930 11822 4964
rect 11856 4930 11914 4964
rect 11948 4930 12006 4964
rect 12040 4930 12098 4964
rect 12132 4930 12190 4964
rect 12224 4930 12282 4964
rect 12316 4930 12374 4964
rect 12408 4930 12466 4964
rect 12500 4930 12558 4964
rect 12592 4930 12650 4964
rect 12684 4930 12742 4964
rect 12776 4930 12834 4964
rect 12868 4930 12926 4964
rect 12960 4930 13018 4964
rect 13052 4930 13110 4964
rect 13144 4930 13202 4964
rect 13236 4930 13294 4964
rect 13328 4930 13386 4964
rect 13420 4930 13478 4964
rect 13512 4930 13570 4964
rect 13604 4930 13662 4964
rect 13696 4930 13754 4964
rect 13788 4930 13846 4964
rect 13880 4930 13938 4964
rect 13972 4930 14030 4964
rect 14064 4930 14122 4964
rect 14156 4930 14214 4964
rect 14248 4930 14306 4964
rect 14340 4930 14398 4964
rect 14432 4930 14490 4964
rect 14524 4930 14582 4964
rect 14616 4930 14674 4964
rect 14708 4930 14766 4964
rect 14800 4930 14858 4964
rect 14892 4930 14950 4964
rect 14984 4930 15042 4964
rect 15076 4930 15134 4964
rect 15168 4930 15226 4964
rect 15260 4930 15318 4964
rect 15352 4930 15410 4964
rect 15444 4930 15502 4964
rect 15536 4930 15594 4964
rect 15628 4930 15686 4964
rect 15720 4930 15778 4964
rect 15812 4930 15870 4964
rect 15904 4930 15962 4964
rect 15996 4930 16054 4964
rect 16088 4930 16146 4964
rect 16180 4930 16238 4964
rect 16272 4930 16330 4964
rect 16364 4930 16422 4964
rect 16456 4930 16514 4964
rect 16548 4930 16606 4964
rect 16640 4930 16698 4964
rect 16732 4930 16790 4964
rect 16824 4930 16882 4964
rect 16916 4930 16974 4964
rect 17008 4930 17066 4964
rect 17100 4930 17158 4964
rect 17192 4930 17250 4964
rect 17284 4930 17342 4964
rect 17376 4930 17434 4964
rect 17468 4930 17526 4964
rect 17560 4930 17618 4964
rect 17652 4930 17710 4964
rect 17744 4930 17802 4964
rect 17836 4930 17894 4964
rect 17928 4930 17986 4964
rect 18020 4930 18078 4964
rect 18112 4930 18170 4964
rect 18204 4930 18262 4964
rect 18296 4930 18354 4964
rect 18388 4930 18446 4964
rect 18480 4930 18538 4964
rect 18572 4930 18630 4964
rect 18664 4930 18722 4964
rect 18756 4930 18814 4964
rect 18848 4930 18906 4964
rect 18940 4930 18998 4964
rect 19032 4930 19090 4964
rect 19124 4930 19182 4964
rect 19216 4930 19274 4964
rect 19308 4930 19366 4964
rect 19400 4930 19458 4964
rect 19492 4930 19550 4964
rect 19584 4930 19642 4964
rect 19676 4930 19734 4964
rect 19768 4930 19826 4964
rect 19860 4930 19898 4964
rect 19932 4930 19990 4964
rect 20024 4930 20082 4964
rect 20116 4930 20174 4964
rect 20208 4930 20266 4964
rect 20300 4930 20358 4964
rect 20392 4930 20450 4964
rect 20484 4930 20542 4964
rect 20576 4930 20634 4964
rect 20668 4930 20726 4964
rect 20760 4930 20818 4964
rect 20852 4930 20910 4964
rect 20944 4930 21002 4964
rect 21036 4930 21094 4964
rect 21128 4930 21186 4964
rect 21220 4930 21278 4964
rect 21312 4930 21370 4964
rect 21404 4930 21462 4964
rect 21496 4930 21554 4964
rect 21588 4930 21646 4964
rect 21680 4930 21738 4964
rect 21772 4930 21830 4964
rect 21864 4930 21922 4964
rect 21956 4930 22014 4964
rect 22048 4930 22106 4964
rect 22140 4930 22198 4964
rect 22232 4930 22290 4964
rect 22324 4930 22382 4964
rect 22416 4930 22474 4964
rect 22508 4930 22566 4964
rect 22600 4930 22658 4964
rect 22692 4930 22750 4964
rect 22784 4930 22842 4964
rect 22876 4930 22934 4964
rect 22968 4930 23026 4964
rect 23060 4930 23118 4964
rect 23152 4930 23210 4964
rect 23244 4930 23302 4964
rect 23336 4930 23394 4964
rect 23428 4930 23457 4964
rect 24793 4915 24897 4950
rect 24793 4881 24824 4915
rect 24858 4881 24897 4915
rect 24793 4852 24897 4881
rect 25191 4744 25523 4760
rect 25191 4710 25217 4744
rect 25251 4710 25297 4744
rect 25331 4710 25377 4744
rect 25411 4710 25457 4744
rect 25491 4710 25523 4744
rect 25191 4692 25523 4710
rect 25923 4744 26255 4760
rect 25923 4710 25949 4744
rect 25983 4710 26029 4744
rect 26063 4710 26109 4744
rect 26143 4710 26189 4744
rect 26223 4710 26255 4744
rect 25923 4692 26255 4710
rect 26525 4744 26857 4760
rect 26525 4710 26557 4744
rect 26591 4710 26637 4744
rect 26671 4710 26717 4744
rect 26751 4710 26797 4744
rect 26831 4710 26857 4744
rect 26525 4692 26857 4710
rect 27135 4744 27467 4760
rect 27135 4710 27161 4744
rect 27195 4710 27241 4744
rect 27275 4710 27321 4744
rect 27355 4710 27401 4744
rect 27435 4710 27467 4744
rect 27135 4692 27467 4710
rect 27737 4744 28069 4760
rect 27737 4710 27769 4744
rect 27803 4710 27849 4744
rect 27883 4710 27929 4744
rect 27963 4710 28009 4744
rect 28043 4710 28069 4744
rect 27737 4692 28069 4710
rect 28473 4744 28805 4760
rect 28473 4710 28499 4744
rect 28533 4710 28579 4744
rect 28613 4710 28659 4744
rect 28693 4710 28739 4744
rect 28773 4710 28805 4744
rect 28473 4692 28805 4710
rect 29075 4744 29407 4760
rect 29075 4710 29107 4744
rect 29141 4710 29187 4744
rect 29221 4710 29267 4744
rect 29301 4710 29347 4744
rect 29381 4710 29407 4744
rect 29075 4692 29407 4710
rect 29809 4744 30141 4760
rect 29809 4710 29841 4744
rect 29875 4710 29921 4744
rect 29955 4710 30001 4744
rect 30035 4710 30081 4744
rect 30115 4710 30141 4744
rect 29809 4692 30141 4710
rect 25577 4298 25606 4332
rect 25640 4298 25698 4332
rect 25732 4298 25790 4332
rect 25824 4298 25882 4332
rect 25916 4298 25974 4332
rect 26008 4298 26066 4332
rect 26100 4298 26158 4332
rect 26192 4298 26250 4332
rect 26284 4298 26342 4332
rect 26376 4298 26433 4332
rect 26467 4298 26526 4332
rect 26560 4298 26618 4332
rect 26652 4298 26710 4332
rect 26744 4298 26802 4332
rect 26836 4298 26894 4332
rect 26928 4298 26986 4332
rect 27020 4298 27078 4332
rect 27112 4298 27170 4332
rect 27204 4298 27262 4332
rect 27296 4298 27354 4332
rect 27388 4298 27446 4332
rect 27480 4298 27538 4332
rect 27572 4298 27630 4332
rect 27664 4298 27722 4332
rect 27756 4298 27814 4332
rect 27848 4298 27906 4332
rect 27940 4298 27998 4332
rect 28032 4298 28090 4332
rect 28124 4298 28182 4332
rect 28216 4298 28274 4332
rect 28308 4298 28366 4332
rect 28400 4298 28458 4332
rect 28492 4298 28550 4332
rect 28584 4298 28642 4332
rect 28676 4298 28734 4332
rect 28768 4298 28826 4332
rect 28860 4298 28918 4332
rect 28952 4298 29010 4332
rect 29044 4298 29102 4332
rect 29136 4298 29194 4332
rect 29228 4298 29286 4332
rect 29320 4298 29378 4332
rect 29412 4298 29470 4332
rect 29504 4298 29562 4332
rect 29596 4298 29654 4332
rect 29688 4298 29746 4332
rect 29780 4298 29838 4332
rect 29872 4298 29930 4332
rect 29964 4298 30022 4332
rect 30056 4298 30114 4332
rect 30148 4298 30206 4332
rect 30240 4298 30298 4332
rect 30332 4298 30361 4332
rect 11089 4045 11117 4079
rect 11151 4045 11210 4079
rect 11244 4045 11302 4079
rect 11336 4045 11394 4079
rect 11428 4045 11486 4079
rect 11520 4045 11578 4079
rect 11612 4045 11670 4079
rect 11704 4045 11762 4079
rect 11796 4045 11854 4079
rect 11888 4045 11917 4079
rect 13630 4057 13660 4091
rect 13694 4057 13752 4091
rect 13786 4057 13844 4091
rect 13878 4057 13936 4091
rect 13970 4057 14028 4091
rect 14062 4057 14120 4091
rect 14154 4057 14212 4091
rect 14246 4057 14304 4091
rect 14338 4057 14396 4091
rect 14430 4057 14488 4091
rect 14522 4057 14580 4091
rect 14614 4057 14672 4091
rect 14706 4057 14764 4091
rect 14798 4057 14856 4091
rect 14890 4057 14948 4091
rect 14982 4057 15040 4091
rect 15074 4057 15132 4091
rect 15166 4057 15224 4091
rect 15258 4057 15316 4091
rect 15350 4057 15408 4091
rect 15442 4057 15500 4091
rect 15534 4057 15592 4091
rect 15626 4057 15684 4091
rect 15718 4057 15776 4091
rect 15810 4057 15868 4091
rect 15902 4057 15960 4091
rect 15994 4057 16052 4091
rect 16086 4057 16144 4091
rect 16178 4057 16236 4091
rect 16270 4057 16328 4091
rect 16362 4057 16420 4091
rect 16454 4057 16512 4091
rect 16546 4057 16604 4091
rect 16638 4057 16696 4091
rect 16730 4057 16788 4091
rect 16822 4057 16880 4091
rect 16914 4057 16972 4091
rect 17006 4057 17064 4091
rect 17098 4057 17156 4091
rect 17190 4057 17248 4091
rect 17282 4057 17340 4091
rect 17374 4057 17432 4091
rect 17466 4057 17524 4091
rect 17558 4057 17616 4091
rect 17650 4057 17708 4091
rect 17742 4057 17800 4091
rect 17834 4057 17892 4091
rect 17926 4057 17984 4091
rect 18018 4057 18076 4091
rect 18110 4057 18168 4091
rect 18202 4057 18260 4091
rect 18294 4057 18352 4091
rect 18386 4057 18444 4091
rect 18478 4057 18536 4091
rect 18570 4057 18628 4091
rect 18662 4057 18720 4091
rect 18754 4057 18812 4091
rect 18846 4057 18904 4091
rect 18938 4057 18996 4091
rect 19030 4057 19088 4091
rect 19122 4057 19180 4091
rect 19214 4057 19272 4091
rect 19306 4057 19364 4091
rect 19398 4057 19456 4091
rect 19490 4057 19548 4091
rect 19582 4057 19640 4091
rect 19674 4057 19732 4091
rect 19766 4057 19824 4091
rect 19858 4057 19916 4091
rect 19950 4057 20008 4091
rect 20042 4057 20100 4091
rect 20134 4057 20192 4091
rect 20226 4057 20284 4091
rect 20318 4057 20357 4091
rect 20410 4057 20449 4091
rect 20502 4057 20541 4091
rect 20594 4057 20633 4091
rect 20686 4057 20725 4091
rect 20778 4057 20817 4091
rect 20870 4057 20909 4091
rect 20962 4057 21001 4091
rect 21054 4057 21093 4091
rect 21146 4057 21185 4091
rect 21238 4057 21277 4091
rect 21330 4057 21369 4091
rect 21422 4057 21461 4091
rect 21514 4057 21553 4091
rect 21606 4057 21645 4091
rect 21698 4057 21737 4091
rect 21790 4057 21829 4091
rect 21882 4057 21921 4091
rect 21974 4057 22013 4091
rect 22066 4057 22105 4091
rect 22158 4057 22197 4091
rect 22250 4057 22289 4091
rect 22342 4057 22381 4091
rect 22434 4057 22473 4091
rect 22507 4057 22565 4091
rect 22599 4057 22657 4091
rect 22691 4057 22749 4091
rect 22783 4057 22841 4091
rect 22875 4057 22933 4091
rect 22967 4057 23025 4091
rect 23059 4057 23117 4091
rect 23151 4057 23209 4091
rect 23243 4057 23301 4091
rect 23335 4057 23393 4091
rect 23427 4057 23455 4091
rect 11496 3184 11525 3218
rect 11559 3184 11617 3218
rect 11651 3184 11709 3218
rect 11743 3184 11801 3218
rect 11835 3184 11893 3218
rect 11927 3184 11985 3218
rect 12019 3184 12077 3218
rect 12111 3184 12169 3218
rect 12203 3184 12261 3218
rect 12295 3184 12353 3218
rect 12387 3184 12445 3218
rect 12479 3184 12537 3218
rect 12571 3184 12629 3218
rect 12663 3184 12721 3218
rect 12755 3184 12813 3218
rect 12847 3184 12905 3218
rect 12939 3184 12997 3218
rect 13031 3184 13089 3218
rect 13123 3184 13181 3218
rect 13215 3184 13273 3218
rect 13307 3184 13365 3218
rect 13399 3184 13457 3218
rect 13491 3184 13549 3218
rect 13583 3184 13641 3218
rect 13675 3184 13733 3218
rect 13767 3184 13825 3218
rect 13859 3184 13917 3218
rect 13951 3184 14009 3218
rect 14043 3184 14101 3218
rect 14135 3184 14193 3218
rect 14227 3184 14285 3218
rect 14319 3184 14377 3218
rect 14411 3184 14469 3218
rect 14503 3184 14561 3218
rect 14595 3184 14653 3218
rect 14687 3184 14745 3218
rect 14779 3184 14837 3218
rect 14871 3184 14929 3218
rect 14963 3184 15021 3218
rect 15055 3184 15113 3218
rect 15147 3184 15205 3218
rect 15239 3184 15297 3218
rect 15331 3184 15389 3218
rect 15423 3184 15481 3218
rect 15515 3184 15573 3218
rect 15607 3184 15665 3218
rect 15699 3184 15757 3218
rect 15791 3184 15849 3218
rect 15883 3184 15941 3218
rect 15975 3184 16033 3218
rect 16067 3184 16125 3218
rect 16159 3184 16217 3218
rect 16251 3184 16309 3218
rect 16343 3184 16401 3218
rect 16435 3184 16493 3218
rect 16527 3184 16585 3218
rect 16619 3184 16677 3218
rect 16711 3184 16769 3218
rect 16803 3184 16861 3218
rect 16895 3184 16953 3218
rect 16987 3184 17045 3218
rect 17079 3184 17137 3218
rect 17171 3184 17229 3218
rect 17263 3184 17321 3218
rect 17355 3184 17413 3218
rect 17447 3184 17505 3218
rect 17539 3184 17597 3218
rect 17631 3184 17689 3218
rect 17723 3184 17781 3218
rect 17815 3184 17873 3218
rect 17907 3184 17965 3218
rect 17999 3184 18057 3218
rect 18091 3184 18149 3218
rect 18183 3184 18241 3218
rect 18275 3184 18333 3218
rect 18367 3184 18425 3218
rect 18459 3184 18517 3218
rect 18551 3184 18609 3218
rect 18643 3184 18701 3218
rect 18735 3184 18793 3218
rect 18827 3184 18885 3218
rect 18919 3184 18977 3218
rect 19011 3184 19069 3218
rect 19103 3184 19161 3218
rect 19195 3184 19253 3218
rect 19287 3184 19345 3218
rect 19379 3184 19437 3218
rect 19471 3184 19529 3218
rect 19563 3184 19621 3218
rect 19655 3184 19713 3218
rect 19747 3184 19805 3218
rect 19839 3184 19897 3218
rect 19931 3184 19989 3218
rect 20023 3184 20081 3218
rect 20115 3184 20173 3218
rect 20207 3184 20265 3218
rect 20299 3184 20357 3218
rect 20391 3184 20449 3218
rect 20483 3184 20541 3218
rect 20575 3184 20633 3218
rect 20667 3184 20725 3218
rect 20759 3184 20817 3218
rect 20851 3184 20909 3218
rect 20943 3184 21001 3218
rect 21035 3184 21093 3218
rect 21127 3184 21185 3218
rect 21219 3184 21277 3218
rect 21311 3184 21369 3218
rect 21403 3184 21461 3218
rect 21495 3184 21553 3218
rect 21587 3184 21645 3218
rect 21679 3184 21737 3218
rect 21771 3184 21829 3218
rect 21863 3184 21921 3218
rect 21955 3184 22013 3218
rect 22047 3184 22105 3218
rect 22139 3184 22197 3218
rect 22231 3184 22289 3218
rect 22323 3184 22381 3218
rect 22415 3184 22473 3218
rect 22507 3184 22565 3218
rect 22599 3184 22657 3218
rect 22691 3184 22749 3218
rect 22783 3184 22841 3218
rect 22875 3184 22933 3218
rect 22967 3184 23025 3218
rect 23059 3184 23117 3218
rect 23151 3184 23209 3218
rect 23243 3184 23301 3218
rect 23335 3184 23393 3218
rect 23427 3184 23456 3218
rect 25577 3033 25606 3067
rect 25640 3033 25698 3067
rect 25732 3033 25790 3067
rect 25824 3033 25882 3067
rect 25916 3033 25974 3067
rect 26008 3033 26066 3067
rect 26100 3033 26158 3067
rect 26192 3033 26250 3067
rect 26284 3033 26342 3067
rect 26376 3033 26434 3067
rect 26468 3033 26526 3067
rect 26560 3033 26618 3067
rect 26652 3033 26710 3067
rect 26744 3033 26802 3067
rect 26836 3033 26894 3067
rect 26928 3033 26986 3067
rect 27020 3033 27078 3067
rect 27112 3033 27171 3067
rect 27205 3033 27262 3067
rect 27296 3033 27354 3067
rect 27388 3033 27446 3067
rect 27480 3033 27539 3067
rect 27573 3033 27630 3067
rect 27664 3033 27722 3067
rect 27756 3033 27814 3067
rect 27848 3033 27906 3067
rect 27940 3033 27998 3067
rect 28032 3033 28090 3067
rect 28124 3033 28182 3067
rect 28216 3033 28274 3067
rect 28308 3033 28366 3067
rect 28400 3033 28458 3067
rect 28492 3033 28550 3067
rect 28584 3033 28642 3067
rect 28676 3033 28733 3067
rect 28767 3033 28825 3067
rect 28859 3033 28918 3067
rect 28952 3033 29010 3067
rect 29044 3033 29102 3067
rect 29136 3033 29193 3067
rect 29227 3033 29286 3067
rect 29320 3033 29377 3067
rect 29411 3033 29470 3067
rect 29504 3033 29562 3067
rect 29596 3033 29654 3067
rect 29688 3033 29746 3067
rect 29780 3033 29838 3067
rect 29872 3033 29930 3067
rect 29964 3033 30022 3067
rect 30056 3033 30114 3067
rect 30148 3033 30206 3067
rect 30240 3033 30298 3067
rect 30332 3033 30361 3067
rect 25577 1766 25606 1800
rect 25640 1766 25698 1800
rect 25732 1766 25790 1800
rect 25824 1766 25882 1800
rect 25916 1766 25974 1800
rect 26008 1766 26066 1800
rect 26100 1766 26158 1800
rect 26192 1766 26250 1800
rect 26284 1766 26342 1800
rect 26376 1766 26434 1800
rect 26468 1766 26526 1800
rect 26560 1766 26618 1800
rect 26652 1766 26710 1800
rect 26744 1766 26802 1800
rect 26836 1766 26894 1800
rect 26928 1766 26986 1800
rect 27020 1766 27078 1800
rect 27112 1766 27170 1800
rect 27204 1766 27262 1800
rect 27296 1766 27354 1800
rect 27388 1766 27446 1800
rect 27480 1766 27538 1800
rect 27572 1766 27630 1800
rect 27664 1766 27722 1800
rect 27756 1766 27814 1800
rect 27848 1766 27906 1800
rect 27940 1766 27998 1800
rect 28032 1766 28090 1800
rect 28124 1766 28182 1800
rect 28216 1766 28274 1800
rect 28308 1766 28366 1800
rect 28400 1766 28458 1800
rect 28492 1766 28550 1800
rect 28584 1766 28642 1800
rect 28676 1766 28734 1800
rect 28768 1766 28826 1800
rect 28860 1766 28918 1800
rect 28952 1766 29010 1800
rect 29044 1766 29102 1800
rect 29136 1766 29194 1800
rect 29228 1766 29286 1800
rect 29320 1766 29378 1800
rect 29412 1766 29470 1800
rect 29504 1766 29562 1800
rect 29596 1766 29654 1800
rect 29688 1766 29746 1800
rect 29780 1766 29838 1800
rect 29872 1766 29930 1800
rect 29964 1766 30022 1800
rect 30056 1766 30114 1800
rect 30148 1766 30206 1800
rect 30240 1766 30298 1800
rect 30332 1766 30361 1800
rect 8577 804 8606 838
rect 8640 804 8698 838
rect 8732 804 8790 838
rect 8824 804 8882 838
rect 8916 804 8974 838
rect 9008 804 9066 838
rect 9100 804 9158 838
rect 9192 804 9250 838
rect 9284 804 9342 838
rect 9376 804 9434 838
rect 9468 804 9526 838
rect 9560 804 9618 838
rect 9652 804 9710 838
rect 9744 804 9802 838
rect 9836 804 9894 838
rect 9928 804 9986 838
rect 10020 804 10078 838
rect 10112 804 10170 838
rect 10204 804 10262 838
rect 10296 804 10354 838
rect 10388 804 10446 838
rect 10480 804 10538 838
rect 10572 804 10630 838
rect 10664 804 10722 838
rect 10756 804 10814 838
rect 10848 804 10906 838
rect 10940 804 10998 838
rect 11032 804 11090 838
rect 11124 804 11182 838
rect 11216 804 11274 838
rect 11308 804 11366 838
rect 11400 804 11429 838
rect 12961 804 12990 838
rect 13024 804 13082 838
rect 13116 804 13174 838
rect 13208 804 13266 838
rect 13300 804 13358 838
rect 13392 804 13450 838
rect 13484 804 13542 838
rect 13576 804 13634 838
rect 13668 804 13726 838
rect 13760 804 13818 838
rect 13852 804 13910 838
rect 13944 804 14002 838
rect 14036 804 14094 838
rect 14128 804 14186 838
rect 14220 804 14278 838
rect 14312 804 14370 838
rect 14404 804 14462 838
rect 14496 804 14554 838
rect 14588 804 14646 838
rect 14680 804 14738 838
rect 14772 804 14830 838
rect 14864 804 14922 838
rect 14956 804 15014 838
rect 15048 804 15106 838
rect 15140 804 15198 838
rect 15232 804 15290 838
rect 15324 804 15382 838
rect 15416 804 15474 838
rect 15508 804 15566 838
rect 15600 804 15658 838
rect 15692 804 15750 838
rect 15784 804 15813 838
rect 8575 -338 8604 -304
rect 8638 -338 8696 -304
rect 8730 -338 8788 -304
rect 8822 -338 8880 -304
rect 8914 -338 8972 -304
rect 9006 -338 9064 -304
rect 9098 -338 9156 -304
rect 9190 -338 9248 -304
rect 9282 -338 9340 -304
rect 9374 -338 9432 -304
rect 9466 -338 9524 -304
rect 9558 -338 9616 -304
rect 9650 -338 9708 -304
rect 9742 -338 9800 -304
rect 9834 -338 9892 -304
rect 9926 -338 9984 -304
rect 10018 -338 10076 -304
rect 10110 -338 10168 -304
rect 10202 -338 10260 -304
rect 10294 -338 10352 -304
rect 10386 -338 10444 -304
rect 10478 -338 10536 -304
rect 10570 -338 10628 -304
rect 10662 -338 10720 -304
rect 10754 -338 10812 -304
rect 10846 -338 10904 -304
rect 10938 -338 10996 -304
rect 11030 -338 11088 -304
rect 11122 -338 11180 -304
rect 11214 -338 11272 -304
rect 11306 -338 11364 -304
rect 11398 -338 11456 -304
rect 11490 -338 11548 -304
rect 11582 -338 11640 -304
rect 11674 -338 11732 -304
rect 11766 -338 11824 -304
rect 11858 -338 11916 -304
rect 11950 -338 12008 -304
rect 12042 -338 12100 -304
rect 12134 -338 12192 -304
rect 12226 -338 12284 -304
rect 12318 -338 12376 -304
rect 12410 -338 12468 -304
rect 12502 -338 12560 -304
rect 12594 -338 12652 -304
rect 12686 -338 12744 -304
rect 12778 -338 12836 -304
rect 12870 -338 12928 -304
rect 12962 -338 13020 -304
rect 13054 -338 13112 -304
rect 13146 -338 13204 -304
rect 13238 -338 13296 -304
rect 13330 -338 13388 -304
rect 13422 -338 13480 -304
rect 13514 -338 13572 -304
rect 13606 -338 13664 -304
rect 13698 -338 13756 -304
rect 13790 -338 13848 -304
rect 13882 -338 13940 -304
rect 13974 -338 14032 -304
rect 14066 -338 14124 -304
rect 14158 -338 14216 -304
rect 14250 -334 14820 -304
rect 14250 -338 14279 -334
rect 14791 -338 14820 -334
rect 14854 -338 14912 -304
rect 14946 -338 15004 -304
rect 15038 -338 15096 -304
rect 15130 -338 15188 -304
rect 15222 -338 15280 -304
rect 15314 -338 15372 -304
rect 15406 -338 15464 -304
rect 15498 -338 15556 -304
rect 15590 -338 15648 -304
rect 15682 -338 15740 -304
rect 15774 -338 15832 -304
rect 15866 -338 15924 -304
rect 15958 -338 16016 -304
rect 16050 -338 16108 -304
rect 16142 -338 16200 -304
rect 16234 -338 16292 -304
rect 16326 -338 16384 -304
rect 16418 -338 16476 -304
rect 16510 -338 16568 -304
rect 16602 -338 16660 -304
rect 16694 -338 16752 -304
rect 16786 -338 16844 -304
rect 16878 -338 16936 -304
rect 16970 -338 17028 -304
rect 17062 -338 17120 -304
rect 17154 -338 17212 -304
rect 17246 -338 17304 -304
rect 17338 -338 17396 -304
rect 17430 -338 17488 -304
rect 17522 -338 17580 -304
rect 17614 -338 17672 -304
rect 17706 -338 17764 -304
rect 17798 -338 17856 -304
rect 17890 -338 17948 -304
rect 17982 -338 18040 -304
rect 18074 -338 18132 -304
rect 18166 -338 18224 -304
rect 18258 -338 18316 -304
rect 18350 -338 18408 -304
rect 18442 -338 18500 -304
rect 18534 -338 18592 -304
rect 18626 -338 18684 -304
rect 18718 -338 18776 -304
rect 18810 -338 18868 -304
rect 18902 -338 18960 -304
rect 18994 -338 19052 -304
rect 19086 -338 19144 -304
rect 19178 -338 19236 -304
rect 19270 -338 19328 -304
rect 19362 -338 19420 -304
rect 19454 -338 19512 -304
rect 19546 -338 19604 -304
rect 19638 -338 19696 -304
rect 19730 -338 19788 -304
rect 19822 -338 19880 -304
rect 19914 -338 19972 -304
rect 20006 -338 20064 -304
rect 20098 -338 20156 -304
rect 20190 -338 20248 -304
rect 20282 -338 20340 -304
rect 20374 -338 20432 -304
rect 20466 -334 20586 -304
rect 20466 -338 20495 -334
rect 20557 -338 20586 -334
rect 20620 -338 20678 -304
rect 20712 -338 20770 -304
rect 20804 -338 20862 -304
rect 20896 -338 20954 -304
rect 20988 -338 21046 -304
rect 21080 -338 21138 -304
rect 21172 -338 21230 -304
rect 21264 -338 21322 -304
rect 21356 -338 21414 -304
rect 21448 -338 21506 -304
rect 21540 -338 21598 -304
rect 21632 -338 21690 -304
rect 21724 -338 21782 -304
rect 21816 -338 21874 -304
rect 21908 -338 21966 -304
rect 22000 -338 22058 -304
rect 22092 -338 22150 -304
rect 22184 -338 22242 -304
rect 22276 -338 22334 -304
rect 22368 -338 22426 -304
rect 22460 -338 22518 -304
rect 22552 -338 22610 -304
rect 22644 -338 22702 -304
rect 22736 -338 22794 -304
rect 22828 -338 22886 -304
rect 22920 -338 22978 -304
rect 23012 -338 23070 -304
rect 23104 -338 23162 -304
rect 23196 -338 23254 -304
rect 23288 -338 23346 -304
rect 23380 -338 23438 -304
rect 23472 -338 23530 -304
rect 23564 -338 23622 -304
rect 23656 -338 23714 -304
rect 23748 -338 23806 -304
rect 23840 -338 23898 -304
rect 23932 -338 23990 -304
rect 24024 -338 24082 -304
rect 24116 -338 24174 -304
rect 24208 -338 24266 -304
rect 24300 -338 24358 -304
rect 24392 -338 24450 -304
rect 24484 -338 24542 -304
rect 24576 -338 24634 -304
rect 24668 -338 24726 -304
rect 24760 -338 24818 -304
rect 24852 -338 24910 -304
rect 24944 -338 25002 -304
rect 25036 -338 25094 -304
rect 25128 -334 25189 -304
rect 25128 -338 25157 -334
rect 8574 -1022 8604 -992
rect 8575 -1026 8604 -1022
rect 8638 -1026 8696 -992
rect 8730 -1026 8788 -992
rect 8822 -1026 8880 -992
rect 8914 -1026 8972 -992
rect 9006 -1026 9064 -992
rect 9098 -1026 9156 -992
rect 9190 -1026 9248 -992
rect 9282 -1026 9340 -992
rect 9374 -1026 9432 -992
rect 9466 -1026 9524 -992
rect 9558 -1026 9616 -992
rect 9650 -1026 9708 -992
rect 9742 -1026 9800 -992
rect 9834 -1026 9892 -992
rect 9926 -1026 9984 -992
rect 10018 -1026 10076 -992
rect 10110 -1026 10168 -992
rect 10202 -1026 10260 -992
rect 10294 -1026 10352 -992
rect 10386 -1026 10444 -992
rect 10478 -1026 10536 -992
rect 10570 -1026 10628 -992
rect 10662 -1026 10720 -992
rect 10754 -1026 10812 -992
rect 10846 -1026 10904 -992
rect 10938 -1026 10996 -992
rect 11030 -1026 11088 -992
rect 11122 -1026 11180 -992
rect 11214 -1026 11272 -992
rect 11306 -1026 11364 -992
rect 11398 -1026 11456 -992
rect 11490 -1026 11548 -992
rect 11582 -1026 11640 -992
rect 11674 -1026 11732 -992
rect 11766 -1026 11824 -992
rect 11858 -1026 11916 -992
rect 11950 -1026 12008 -992
rect 12042 -1026 12100 -992
rect 12134 -1026 12192 -992
rect 12226 -1026 12284 -992
rect 12318 -1026 12376 -992
rect 12410 -1026 12468 -992
rect 12502 -1026 12560 -992
rect 12594 -1026 12652 -992
rect 12686 -1026 12744 -992
rect 12778 -1026 12836 -992
rect 12870 -1026 12928 -992
rect 12962 -1026 13020 -992
rect 13054 -1026 13112 -992
rect 13146 -1026 13204 -992
rect 13238 -1026 13296 -992
rect 13330 -1026 13388 -992
rect 13422 -1026 13480 -992
rect 13514 -1026 13572 -992
rect 13606 -1026 13664 -992
rect 13698 -1026 13756 -992
rect 13790 -1026 13848 -992
rect 13882 -1026 13940 -992
rect 13974 -1026 14032 -992
rect 14066 -1026 14124 -992
rect 14158 -1026 14216 -992
rect 14250 -1026 14308 -992
rect 14342 -1026 14400 -992
rect 14434 -1026 14492 -992
rect 14526 -1026 14584 -992
rect 14618 -1026 14676 -992
rect 14710 -1026 14768 -992
rect 14802 -1026 14860 -992
rect 14894 -1026 14952 -992
rect 14986 -1026 15044 -992
rect 15078 -1026 15136 -992
rect 15170 -1026 15228 -992
rect 15262 -1026 15320 -992
rect 15354 -1026 15412 -992
rect 15446 -1026 15504 -992
rect 15538 -1026 15596 -992
rect 15630 -1026 15688 -992
rect 15722 -1026 15780 -992
rect 15814 -1026 15872 -992
rect 15906 -1026 15964 -992
rect 15998 -1026 16056 -992
rect 16090 -1026 16148 -992
rect 16182 -1026 16240 -992
rect 16274 -1026 16332 -992
rect 16366 -1026 16424 -992
rect 16458 -1026 16516 -992
rect 16550 -1026 16608 -992
rect 16642 -1026 16700 -992
rect 16734 -1026 16792 -992
rect 16826 -1026 16884 -992
rect 16918 -1026 16976 -992
rect 17010 -1026 17068 -992
rect 17102 -1026 17160 -992
rect 17194 -1026 17252 -992
rect 17286 -1026 17344 -992
rect 17378 -1026 17436 -992
rect 17470 -1026 17528 -992
rect 17562 -1026 17620 -992
rect 17654 -1026 17712 -992
rect 17746 -1026 17804 -992
rect 17838 -1026 17896 -992
rect 17930 -1026 17988 -992
rect 18022 -1026 18080 -992
rect 18114 -1026 18172 -992
rect 18206 -1026 18264 -992
rect 18298 -1026 18356 -992
rect 18390 -1026 18448 -992
rect 18482 -1026 18540 -992
rect 18574 -1026 18632 -992
rect 18666 -1026 18724 -992
rect 18758 -1026 18816 -992
rect 18850 -1026 18908 -992
rect 18942 -1026 19000 -992
rect 19034 -1026 19092 -992
rect 19126 -1026 19184 -992
rect 19218 -1026 19276 -992
rect 19310 -1026 19368 -992
rect 19402 -1026 19460 -992
rect 19494 -1026 19552 -992
rect 19586 -1026 19644 -992
rect 19678 -1026 19736 -992
rect 19770 -1026 19828 -992
rect 19862 -1026 19920 -992
rect 19954 -1026 20012 -992
rect 20046 -1026 20104 -992
rect 20138 -1026 20196 -992
rect 20230 -1026 20288 -992
rect 20322 -1026 20380 -992
rect 20414 -1026 20472 -992
rect 20506 -1026 20564 -992
rect 20598 -1026 20656 -992
rect 20690 -1026 20748 -992
rect 20782 -1026 20840 -992
rect 20874 -1026 20932 -992
rect 20966 -1026 21024 -992
rect 21058 -1026 21116 -992
rect 21150 -1026 21208 -992
rect 21242 -1026 21300 -992
rect 21334 -1026 21392 -992
rect 21426 -1026 21484 -992
rect 21518 -1026 21576 -992
rect 21610 -1026 21668 -992
rect 21702 -1026 21760 -992
rect 21794 -1026 21852 -992
rect 21886 -1026 21944 -992
rect 21978 -1026 22036 -992
rect 22070 -1026 22128 -992
rect 22162 -1026 22220 -992
rect 22254 -1026 22312 -992
rect 22346 -1026 22404 -992
rect 22438 -1026 22496 -992
rect 22530 -1026 22588 -992
rect 22622 -1026 22680 -992
rect 22714 -1026 22772 -992
rect 22806 -1026 22864 -992
rect 22898 -1026 22956 -992
rect 22990 -1026 23048 -992
rect 23082 -1026 23140 -992
rect 23174 -1026 23232 -992
rect 23266 -1026 23324 -992
rect 23358 -1026 23416 -992
rect 23450 -1026 23508 -992
rect 23542 -1026 23600 -992
rect 23634 -1026 23692 -992
rect 23726 -1026 23784 -992
rect 23818 -1026 23876 -992
rect 23910 -1026 23968 -992
rect 24002 -1026 24060 -992
rect 24094 -1026 24152 -992
rect 24186 -1026 24244 -992
rect 24278 -1026 24336 -992
rect 24370 -1026 24428 -992
rect 24462 -1026 24520 -992
rect 24554 -1026 24612 -992
rect 24646 -1026 24704 -992
rect 24738 -1026 24796 -992
rect 24830 -1026 24888 -992
rect 24922 -1026 24980 -992
rect 25014 -1026 25072 -992
rect 25106 -1026 25164 -992
rect 25198 -1026 25256 -992
rect 25290 -1026 25319 -992
rect 8575 -1715 8604 -1681
rect 8638 -1715 8696 -1681
rect 8730 -1715 8788 -1681
rect 8822 -1715 8880 -1681
rect 8914 -1715 8972 -1681
rect 9006 -1715 9064 -1681
rect 9098 -1715 9156 -1681
rect 9190 -1715 9248 -1681
rect 9282 -1715 9340 -1681
rect 9374 -1715 9432 -1681
rect 9466 -1715 9524 -1681
rect 9558 -1715 9616 -1681
rect 9650 -1715 9708 -1681
rect 9742 -1715 9800 -1681
rect 9834 -1715 9892 -1681
rect 9926 -1715 9984 -1681
rect 10018 -1715 10076 -1681
rect 10110 -1715 10168 -1681
rect 10202 -1715 10260 -1681
rect 10294 -1715 10352 -1681
rect 10386 -1715 10444 -1681
rect 10478 -1715 10536 -1681
rect 10570 -1715 10628 -1681
rect 10662 -1715 10720 -1681
rect 10754 -1715 10812 -1681
rect 10846 -1715 10904 -1681
rect 10938 -1715 10996 -1681
rect 11030 -1715 11088 -1681
rect 11122 -1715 11180 -1681
rect 11214 -1715 11272 -1681
rect 11306 -1715 11364 -1681
rect 11398 -1715 11456 -1681
rect 11490 -1715 11548 -1681
rect 11582 -1715 11640 -1681
rect 11674 -1715 11732 -1681
rect 11766 -1715 11824 -1681
rect 11858 -1715 11916 -1681
rect 11950 -1715 12008 -1681
rect 12042 -1715 12100 -1681
rect 12134 -1715 12192 -1681
rect 12226 -1715 12284 -1681
rect 12318 -1715 12376 -1681
rect 12410 -1715 12468 -1681
rect 12502 -1715 12560 -1681
rect 12594 -1715 12652 -1681
rect 12686 -1715 12744 -1681
rect 12778 -1715 12836 -1681
rect 12870 -1715 12928 -1681
rect 12962 -1715 13020 -1681
rect 13054 -1715 13112 -1681
rect 13146 -1715 13204 -1681
rect 13238 -1715 13296 -1681
rect 13330 -1715 13388 -1681
rect 13422 -1715 13480 -1681
rect 13514 -1715 13572 -1681
rect 13606 -1715 13664 -1681
rect 13698 -1715 13756 -1681
rect 13790 -1715 13848 -1681
rect 13882 -1715 13940 -1681
rect 13974 -1715 14032 -1681
rect 14066 -1715 14124 -1681
rect 14158 -1715 14216 -1681
rect 14250 -1715 14308 -1681
rect 14342 -1715 14400 -1681
rect 14434 -1715 14492 -1681
rect 14526 -1715 14584 -1681
rect 14618 -1715 14676 -1681
rect 14710 -1715 14768 -1681
rect 14802 -1715 14860 -1681
rect 14894 -1715 14952 -1681
rect 14986 -1715 15044 -1681
rect 15078 -1715 15136 -1681
rect 15170 -1715 15228 -1681
rect 15262 -1715 15320 -1681
rect 15354 -1715 15412 -1681
rect 15446 -1715 15504 -1681
rect 15538 -1715 15596 -1681
rect 15630 -1715 15688 -1681
rect 15722 -1715 15780 -1681
rect 15814 -1715 15872 -1681
rect 15906 -1715 15964 -1681
rect 15998 -1715 16056 -1681
rect 16090 -1715 16148 -1681
rect 16182 -1715 16240 -1681
rect 16274 -1715 16332 -1681
rect 16366 -1715 16424 -1681
rect 16458 -1715 16516 -1681
rect 16550 -1715 16608 -1681
rect 16642 -1715 16700 -1681
rect 16734 -1715 16792 -1681
rect 16826 -1715 16884 -1681
rect 16918 -1715 16976 -1681
rect 17010 -1715 17068 -1681
rect 17102 -1715 17160 -1681
rect 17194 -1715 17252 -1681
rect 17286 -1715 17344 -1681
rect 17378 -1715 17436 -1681
rect 17470 -1715 17528 -1681
rect 17562 -1715 17620 -1681
rect 17654 -1715 17712 -1681
rect 17746 -1715 17804 -1681
rect 17838 -1715 17896 -1681
rect 17930 -1715 17988 -1681
rect 18022 -1715 18080 -1681
rect 18114 -1715 18172 -1681
rect 18206 -1715 18264 -1681
rect 18298 -1715 18356 -1681
rect 18390 -1715 18448 -1681
rect 18482 -1715 18540 -1681
rect 18574 -1715 18632 -1681
rect 18666 -1715 18724 -1681
rect 18758 -1715 18816 -1681
rect 18850 -1715 18908 -1681
rect 18942 -1715 19000 -1681
rect 19034 -1715 19092 -1681
rect 19126 -1715 19184 -1681
rect 19218 -1715 19276 -1681
rect 19310 -1715 19368 -1681
rect 19402 -1715 19460 -1681
rect 19494 -1715 19552 -1681
rect 19586 -1715 19644 -1681
rect 19678 -1715 19736 -1681
rect 19770 -1715 19828 -1681
rect 19862 -1715 19920 -1681
rect 19954 -1715 20012 -1681
rect 20046 -1715 20104 -1681
rect 20138 -1715 20196 -1681
rect 20230 -1715 20288 -1681
rect 20322 -1715 20380 -1681
rect 20414 -1715 20472 -1681
rect 20506 -1715 20564 -1681
rect 20598 -1715 20656 -1681
rect 20690 -1715 20748 -1681
rect 20782 -1715 20840 -1681
rect 20874 -1715 20932 -1681
rect 20966 -1715 21024 -1681
rect 21058 -1715 21116 -1681
rect 21150 -1715 21208 -1681
rect 21242 -1715 21300 -1681
rect 21334 -1715 21392 -1681
rect 21426 -1715 21484 -1681
rect 21518 -1715 21576 -1681
rect 21610 -1715 21668 -1681
rect 21702 -1715 21760 -1681
rect 21794 -1715 21852 -1681
rect 21886 -1715 21944 -1681
rect 21978 -1715 22036 -1681
rect 22070 -1715 22128 -1681
rect 22162 -1715 22220 -1681
rect 22254 -1715 22312 -1681
rect 22346 -1715 22404 -1681
rect 22438 -1715 22496 -1681
rect 22530 -1715 22588 -1681
rect 22622 -1715 22680 -1681
rect 22714 -1715 22772 -1681
rect 22806 -1715 22864 -1681
rect 22898 -1715 22956 -1681
rect 22990 -1715 23048 -1681
rect 23082 -1715 23140 -1681
rect 23174 -1715 23232 -1681
rect 23266 -1715 23324 -1681
rect 23358 -1715 23416 -1681
rect 23450 -1715 23508 -1681
rect 23542 -1715 23600 -1681
rect 23634 -1715 23692 -1681
rect 23726 -1715 23784 -1681
rect 23818 -1715 23876 -1681
rect 23910 -1715 23968 -1681
rect 24002 -1715 24060 -1681
rect 24094 -1715 24152 -1681
rect 24186 -1715 24244 -1681
rect 24278 -1715 24336 -1681
rect 24370 -1715 24428 -1681
rect 24462 -1715 24520 -1681
rect 24554 -1715 24612 -1681
rect 24646 -1715 24704 -1681
rect 24738 -1715 24796 -1681
rect 24830 -1715 24888 -1681
rect 24922 -1715 24980 -1681
rect 25014 -1715 25072 -1681
rect 25106 -1715 25164 -1681
rect 25198 -1715 25256 -1681
rect 25290 -1715 25319 -1681
<< nsubdiff >>
rect 14014 13605 14552 13625
rect 14014 13571 14062 13605
rect 14096 13571 14142 13605
rect 14176 13571 14222 13605
rect 14256 13571 14302 13605
rect 14336 13571 14382 13605
rect 14416 13571 14462 13605
rect 14496 13571 14552 13605
rect 14014 13557 14552 13571
rect 14746 13608 15284 13628
rect 14746 13574 14794 13608
rect 14828 13574 14874 13608
rect 14908 13574 14954 13608
rect 14988 13574 15034 13608
rect 15068 13574 15114 13608
rect 15148 13574 15194 13608
rect 15228 13574 15284 13608
rect 14746 13560 15284 13574
rect 15344 13608 15882 13628
rect 15344 13574 15400 13608
rect 15434 13574 15480 13608
rect 15514 13574 15560 13608
rect 15594 13574 15640 13608
rect 15674 13574 15720 13608
rect 15754 13574 15800 13608
rect 15834 13574 15882 13608
rect 15344 13560 15882 13574
rect 15958 13608 16496 13628
rect 15958 13574 16006 13608
rect 16040 13574 16086 13608
rect 16120 13574 16166 13608
rect 16200 13574 16246 13608
rect 16280 13574 16326 13608
rect 16360 13574 16406 13608
rect 16440 13574 16496 13608
rect 15958 13560 16496 13574
rect 16556 13608 17094 13628
rect 16556 13574 16612 13608
rect 16646 13574 16692 13608
rect 16726 13574 16772 13608
rect 16806 13574 16852 13608
rect 16886 13574 16932 13608
rect 16966 13574 17012 13608
rect 17046 13574 17094 13608
rect 16556 13560 17094 13574
rect 17170 13608 17708 13628
rect 17170 13574 17218 13608
rect 17252 13574 17298 13608
rect 17332 13574 17378 13608
rect 17412 13574 17458 13608
rect 17492 13574 17538 13608
rect 17572 13574 17618 13608
rect 17652 13574 17708 13608
rect 17170 13560 17708 13574
rect 17768 13608 18306 13628
rect 17768 13574 17824 13608
rect 17858 13574 17904 13608
rect 17938 13574 17984 13608
rect 18018 13574 18064 13608
rect 18098 13574 18144 13608
rect 18178 13574 18224 13608
rect 18258 13574 18306 13608
rect 17768 13560 18306 13574
rect 18382 13608 18920 13628
rect 18382 13574 18430 13608
rect 18464 13574 18510 13608
rect 18544 13574 18590 13608
rect 18624 13574 18670 13608
rect 18704 13574 18750 13608
rect 18784 13574 18830 13608
rect 18864 13574 18920 13608
rect 18382 13560 18920 13574
rect 18980 13608 19518 13628
rect 18980 13574 19036 13608
rect 19070 13574 19116 13608
rect 19150 13574 19196 13608
rect 19230 13574 19276 13608
rect 19310 13574 19356 13608
rect 19390 13574 19436 13608
rect 19470 13574 19518 13608
rect 20723 13605 21261 13625
rect 18980 13560 19518 13574
rect 19750 13557 19836 13583
rect 19750 13523 19776 13557
rect 19810 13523 19836 13557
rect 19750 13497 19836 13523
rect 20227 13560 20313 13586
rect 20227 13526 20253 13560
rect 20287 13526 20313 13560
rect 20227 13500 20313 13526
rect 20723 13571 20771 13605
rect 20805 13571 20851 13605
rect 20885 13571 20931 13605
rect 20965 13571 21011 13605
rect 21045 13571 21091 13605
rect 21125 13571 21171 13605
rect 21205 13571 21261 13605
rect 20723 13557 21261 13571
rect 21455 13608 21993 13628
rect 21455 13574 21503 13608
rect 21537 13574 21583 13608
rect 21617 13574 21663 13608
rect 21697 13574 21743 13608
rect 21777 13574 21823 13608
rect 21857 13574 21903 13608
rect 21937 13574 21993 13608
rect 21455 13560 21993 13574
rect 22053 13608 22591 13628
rect 22053 13574 22109 13608
rect 22143 13574 22189 13608
rect 22223 13574 22269 13608
rect 22303 13574 22349 13608
rect 22383 13574 22429 13608
rect 22463 13574 22509 13608
rect 22543 13574 22591 13608
rect 22053 13560 22591 13574
rect 22667 13608 23205 13628
rect 22667 13574 22715 13608
rect 22749 13574 22795 13608
rect 22829 13574 22875 13608
rect 22909 13574 22955 13608
rect 22989 13574 23035 13608
rect 23069 13574 23115 13608
rect 23149 13574 23205 13608
rect 22667 13560 23205 13574
rect 23265 13608 23803 13628
rect 23265 13574 23321 13608
rect 23355 13574 23401 13608
rect 23435 13574 23481 13608
rect 23515 13574 23561 13608
rect 23595 13574 23641 13608
rect 23675 13574 23721 13608
rect 23755 13574 23803 13608
rect 23265 13560 23803 13574
rect 23879 13608 24417 13628
rect 23879 13574 23927 13608
rect 23961 13574 24007 13608
rect 24041 13574 24087 13608
rect 24121 13574 24167 13608
rect 24201 13574 24247 13608
rect 24281 13574 24327 13608
rect 24361 13574 24417 13608
rect 23879 13560 24417 13574
rect 24477 13608 25015 13628
rect 24477 13574 24533 13608
rect 24567 13574 24613 13608
rect 24647 13574 24693 13608
rect 24727 13574 24773 13608
rect 24807 13574 24853 13608
rect 24887 13574 24933 13608
rect 24967 13574 25015 13608
rect 24477 13560 25015 13574
rect 25091 13608 25629 13628
rect 25091 13574 25139 13608
rect 25173 13574 25219 13608
rect 25253 13574 25299 13608
rect 25333 13574 25379 13608
rect 25413 13574 25459 13608
rect 25493 13574 25539 13608
rect 25573 13574 25629 13608
rect 25091 13560 25629 13574
rect 25689 13608 26227 13628
rect 25689 13574 25745 13608
rect 25779 13574 25825 13608
rect 25859 13574 25905 13608
rect 25939 13574 25985 13608
rect 26019 13574 26065 13608
rect 26099 13574 26145 13608
rect 26179 13574 26227 13608
rect 25689 13560 26227 13574
rect 26459 13557 26545 13583
rect 26459 13523 26485 13557
rect 26519 13523 26545 13557
rect 26459 13497 26545 13523
rect 14004 13427 14087 13452
rect 14004 13392 14029 13427
rect 14063 13392 14087 13427
rect 14004 13368 14087 13392
rect 19755 13413 19841 13439
rect 19755 13379 19781 13413
rect 19815 13379 19841 13413
rect 19755 13353 19841 13379
rect 20216 13388 20302 13414
rect 20216 13354 20242 13388
rect 20276 13354 20302 13388
rect 20713 13427 20796 13452
rect 20713 13392 20738 13427
rect 20772 13392 20796 13427
rect 20216 13328 20302 13354
rect 20713 13368 20796 13392
rect 26464 13413 26550 13439
rect 26464 13379 26490 13413
rect 26524 13379 26550 13413
rect 26464 13353 26550 13379
rect 19756 13261 19842 13287
rect 19756 13227 19782 13261
rect 19816 13227 19842 13261
rect 26465 13261 26551 13287
rect 19756 13201 19842 13227
rect 20216 13196 20302 13222
rect 3126 13130 3664 13150
rect 3126 13096 3174 13130
rect 3208 13096 3254 13130
rect 3288 13096 3334 13130
rect 3368 13096 3414 13130
rect 3448 13096 3494 13130
rect 3528 13096 3574 13130
rect 3608 13096 3664 13130
rect 3126 13082 3664 13096
rect 3858 13133 4396 13153
rect 3858 13099 3906 13133
rect 3940 13099 3986 13133
rect 4020 13099 4066 13133
rect 4100 13099 4146 13133
rect 4180 13099 4226 13133
rect 4260 13099 4306 13133
rect 4340 13099 4396 13133
rect 3858 13085 4396 13099
rect 4456 13133 4994 13153
rect 4456 13099 4512 13133
rect 4546 13099 4592 13133
rect 4626 13099 4672 13133
rect 4706 13099 4752 13133
rect 4786 13099 4832 13133
rect 4866 13099 4912 13133
rect 4946 13099 4994 13133
rect 4456 13085 4994 13099
rect 5070 13133 5608 13153
rect 5070 13099 5118 13133
rect 5152 13099 5198 13133
rect 5232 13099 5278 13133
rect 5312 13099 5358 13133
rect 5392 13099 5438 13133
rect 5472 13099 5518 13133
rect 5552 13099 5608 13133
rect 5070 13085 5608 13099
rect 5668 13133 6206 13153
rect 5668 13099 5724 13133
rect 5758 13099 5804 13133
rect 5838 13099 5884 13133
rect 5918 13099 5964 13133
rect 5998 13099 6044 13133
rect 6078 13099 6124 13133
rect 6158 13099 6206 13133
rect 5668 13085 6206 13099
rect 6282 13133 6820 13153
rect 6282 13099 6330 13133
rect 6364 13099 6410 13133
rect 6444 13099 6490 13133
rect 6524 13099 6570 13133
rect 6604 13099 6650 13133
rect 6684 13099 6730 13133
rect 6764 13099 6820 13133
rect 6282 13085 6820 13099
rect 6880 13133 7418 13153
rect 6880 13099 6936 13133
rect 6970 13099 7016 13133
rect 7050 13099 7096 13133
rect 7130 13099 7176 13133
rect 7210 13099 7256 13133
rect 7290 13099 7336 13133
rect 7370 13099 7418 13133
rect 6880 13085 7418 13099
rect 7494 13133 8032 13153
rect 7494 13099 7542 13133
rect 7576 13099 7622 13133
rect 7656 13099 7702 13133
rect 7736 13099 7782 13133
rect 7816 13099 7862 13133
rect 7896 13099 7942 13133
rect 7976 13099 8032 13133
rect 7494 13085 8032 13099
rect 8092 13133 8630 13153
rect 8092 13099 8148 13133
rect 8182 13099 8228 13133
rect 8262 13099 8308 13133
rect 8342 13099 8388 13133
rect 8422 13099 8468 13133
rect 8502 13099 8548 13133
rect 8582 13099 8630 13133
rect 8092 13085 8630 13099
rect 8862 13082 8948 13108
rect 20216 13162 20242 13196
rect 20276 13162 20302 13196
rect 26465 13227 26491 13261
rect 26525 13227 26551 13261
rect 26465 13201 26551 13227
rect 20216 13136 20302 13162
rect 8862 13048 8888 13082
rect 8922 13048 8948 13082
rect 8862 13022 8948 13048
rect 19756 13091 19842 13117
rect 19756 13057 19782 13091
rect 19816 13057 19842 13091
rect 13318 13039 13734 13041
rect 13318 13005 13348 13039
rect 13382 13005 13478 13039
rect 13512 13005 13624 13039
rect 13658 13005 13734 13039
rect 13318 13001 13734 13005
rect 3116 12952 3199 12977
rect 3116 12917 3141 12952
rect 3175 12917 3199 12952
rect 3116 12893 3199 12917
rect 8867 12938 8953 12964
rect 19756 13031 19842 13057
rect 26465 13091 26551 13117
rect 26465 13057 26491 13091
rect 26525 13057 26551 13091
rect 20027 13039 20443 13041
rect 20027 13005 20057 13039
rect 20091 13005 20187 13039
rect 20221 13005 20333 13039
rect 20367 13005 20443 13039
rect 20027 13001 20443 13005
rect 8867 12904 8893 12938
rect 8927 12904 8953 12938
rect 8867 12878 8953 12904
rect 8868 12786 8954 12812
rect 8868 12752 8894 12786
rect 8928 12752 8954 12786
rect 8868 12726 8954 12752
rect 19755 12934 19841 12960
rect 26465 13031 26551 13057
rect 19755 12900 19781 12934
rect 19815 12900 19841 12934
rect 19755 12874 19841 12900
rect 8868 12616 8954 12642
rect 26464 12934 26550 12960
rect 26464 12900 26490 12934
rect 26524 12900 26550 12934
rect 26464 12874 26550 12900
rect 8868 12582 8894 12616
rect 8928 12582 8954 12616
rect 2430 12564 2846 12566
rect 2430 12530 2460 12564
rect 2494 12530 2590 12564
rect 2624 12530 2736 12564
rect 2770 12530 2846 12564
rect 2430 12526 2846 12530
rect 8868 12556 8954 12582
rect 8867 12459 8953 12485
rect 8867 12425 8893 12459
rect 8927 12425 8953 12459
rect 8867 12399 8953 12425
rect 9061 12194 9338 12217
rect 9061 12193 9182 12194
rect 9061 12159 9090 12193
rect 9124 12160 9182 12193
rect 9216 12160 9274 12194
rect 9308 12160 9338 12194
rect 9124 12159 9338 12160
rect 9061 12153 9338 12159
rect 10885 11888 13274 11889
rect 10885 11876 11463 11888
rect 10885 11875 11372 11876
rect 10885 11874 11186 11875
rect 10885 11840 10911 11874
rect 10945 11873 11096 11874
rect 10945 11840 11004 11873
rect 10885 11839 11004 11840
rect 11038 11840 11096 11873
rect 11130 11841 11186 11874
rect 11220 11841 11281 11875
rect 11315 11842 11372 11875
rect 11406 11854 11463 11876
rect 11497 11854 11555 11888
rect 11589 11854 11647 11888
rect 11681 11854 11739 11888
rect 11773 11854 11831 11888
rect 11865 11854 11923 11888
rect 11957 11854 12015 11888
rect 12049 11854 12107 11888
rect 12141 11854 12199 11888
rect 12233 11854 12291 11888
rect 12325 11854 12383 11888
rect 12417 11854 12475 11888
rect 12509 11854 12567 11888
rect 12601 11854 12659 11888
rect 12693 11854 12751 11888
rect 12785 11854 12843 11888
rect 12877 11854 12935 11888
rect 12969 11854 13027 11888
rect 13061 11854 13119 11888
rect 13153 11854 13211 11888
rect 13245 11854 13274 11888
rect 11406 11842 13274 11854
rect 11315 11841 13274 11842
rect 11130 11840 13274 11841
rect 11038 11839 13274 11840
rect 10885 11829 13274 11839
rect 9061 8455 11295 8457
rect 9061 8454 9709 8455
rect 9061 8450 9288 8454
rect 9061 8416 9152 8450
rect 9186 8420 9288 8450
rect 9322 8453 9624 8454
rect 9322 8420 9406 8453
rect 9186 8419 9406 8420
rect 9440 8419 9549 8453
rect 9583 8420 9624 8453
rect 9658 8421 9709 8454
rect 9743 8450 9997 8455
rect 9743 8448 9900 8450
rect 9743 8421 9811 8448
rect 9658 8420 9811 8421
rect 9583 8419 9811 8420
rect 9186 8416 9811 8419
rect 9061 8414 9811 8416
rect 9845 8416 9900 8448
rect 9934 8421 9997 8450
rect 10031 8452 11295 8455
rect 10031 8444 10175 8452
rect 10031 8421 10083 8444
rect 9934 8416 10083 8421
rect 9845 8414 10083 8416
rect 9061 8410 10083 8414
rect 10117 8418 10175 8444
rect 10209 8451 11295 8452
rect 10209 8418 10267 8451
rect 10117 8417 10267 8418
rect 10301 8449 11295 8451
rect 10301 8446 10919 8449
rect 10301 8443 10822 8446
rect 10301 8442 10637 8443
rect 10301 8440 10544 8442
rect 10301 8438 10456 8440
rect 10301 8417 10355 8438
rect 10117 8410 10355 8417
rect 9061 8404 10355 8410
rect 10389 8406 10456 8438
rect 10490 8408 10544 8440
rect 10578 8409 10637 8442
rect 10671 8442 10822 8443
rect 10671 8409 10733 8442
rect 10578 8408 10733 8409
rect 10767 8412 10822 8442
rect 10856 8415 10919 8446
rect 10953 8447 11295 8449
rect 10953 8445 11093 8447
rect 10953 8415 11003 8445
rect 10856 8412 11003 8415
rect 10767 8411 11003 8412
rect 11037 8413 11093 8445
rect 11127 8443 11295 8447
rect 11127 8413 11191 8443
rect 11037 8411 11191 8413
rect 10767 8409 11191 8411
rect 11225 8434 11295 8443
rect 11405 8448 11708 8457
rect 11405 8434 11462 8448
rect 11225 8414 11462 8434
rect 11496 8414 11560 8448
rect 11594 8446 11708 8448
rect 11594 8414 11643 8446
rect 11225 8412 11643 8414
rect 11677 8412 11708 8446
rect 11225 8409 11708 8412
rect 10767 8408 11708 8409
rect 10490 8406 11708 8408
rect 10389 8404 11708 8406
rect 9061 8387 11708 8404
rect 12426 8371 12589 8393
rect 8867 8221 8953 8247
rect 8867 8187 8893 8221
rect 8927 8187 8953 8221
rect 2430 8116 2846 8120
rect 2430 8082 2460 8116
rect 2494 8082 2590 8116
rect 2624 8082 2736 8116
rect 2770 8082 2846 8116
rect 2430 8080 2846 8082
rect 8867 8161 8953 8187
rect 8868 8064 8954 8090
rect 8868 8030 8894 8064
rect 8928 8030 8954 8064
rect 8868 8004 8954 8030
rect 8868 7894 8954 7920
rect 8868 7860 8894 7894
rect 8928 7860 8954 7894
rect 8868 7834 8954 7860
rect 12426 8337 12452 8371
rect 12486 8370 12589 8371
rect 12486 8337 12531 8370
rect 12426 8336 12531 8337
rect 12565 8336 12589 8370
rect 12426 8309 12589 8336
rect 13338 8209 13424 8235
rect 13338 8175 13364 8209
rect 13398 8175 13424 8209
rect 13338 8149 13424 8175
rect 20047 8209 20133 8235
rect 20047 8175 20073 8209
rect 20107 8175 20133 8209
rect 13337 8052 13423 8078
rect 20047 8149 20133 8175
rect 19445 8104 19861 8108
rect 19445 8070 19521 8104
rect 19555 8070 19667 8104
rect 19701 8070 19797 8104
rect 19831 8070 19861 8104
rect 19445 8068 19861 8070
rect 13337 8018 13363 8052
rect 13397 8018 13423 8052
rect 13337 7992 13423 8018
rect 20046 8052 20132 8078
rect 26154 8104 26570 8108
rect 26154 8070 26230 8104
rect 26264 8070 26376 8104
rect 26410 8070 26506 8104
rect 26540 8070 26570 8104
rect 26154 8068 26570 8070
rect 20046 8018 20072 8052
rect 20106 8018 20132 8052
rect 3116 7729 3199 7753
rect 3116 7694 3141 7729
rect 3175 7694 3199 7729
rect 3116 7669 3199 7694
rect 8867 7742 8953 7768
rect 8867 7708 8893 7742
rect 8927 7708 8953 7742
rect 8867 7682 8953 7708
rect 8862 7598 8948 7624
rect 8862 7564 8888 7598
rect 8922 7564 8948 7598
rect 12921 7918 13007 7944
rect 19624 7980 19710 8006
rect 20046 7992 20132 8018
rect 19624 7946 19650 7980
rect 19684 7946 19710 7980
rect 12921 7884 12947 7918
rect 12981 7884 13007 7918
rect 12921 7858 13007 7884
rect 13337 7882 13423 7908
rect 13337 7848 13363 7882
rect 13397 7848 13423 7882
rect 19624 7920 19710 7946
rect 20046 7882 20132 7908
rect 13337 7822 13423 7848
rect 20046 7848 20072 7882
rect 20106 7848 20132 7882
rect 20046 7822 20132 7848
rect 13338 7730 13424 7756
rect 12913 7698 12999 7724
rect 12913 7664 12939 7698
rect 12973 7664 12999 7698
rect 13338 7696 13364 7730
rect 13398 7696 13424 7730
rect 13338 7670 13424 7696
rect 19092 7717 19175 7741
rect 19624 7784 19710 7810
rect 19624 7750 19650 7784
rect 19684 7750 19710 7784
rect 19092 7682 19116 7717
rect 19150 7682 19175 7717
rect 12913 7638 12999 7664
rect 19092 7657 19175 7682
rect 19624 7724 19710 7750
rect 20047 7730 20133 7756
rect 20047 7696 20073 7730
rect 20107 7696 20133 7730
rect 20047 7670 20133 7696
rect 25801 7717 25884 7741
rect 25801 7682 25825 7717
rect 25859 7682 25884 7717
rect 25801 7657 25884 7682
rect 13343 7586 13429 7612
rect 19624 7609 19710 7635
rect 3126 7550 3664 7564
rect 3126 7516 3174 7550
rect 3208 7516 3254 7550
rect 3288 7516 3334 7550
rect 3368 7516 3414 7550
rect 3448 7516 3494 7550
rect 3528 7516 3574 7550
rect 3608 7516 3664 7550
rect 3126 7496 3664 7516
rect 3858 7547 4396 7561
rect 3858 7513 3906 7547
rect 3940 7513 3986 7547
rect 4020 7513 4066 7547
rect 4100 7513 4146 7547
rect 4180 7513 4226 7547
rect 4260 7513 4306 7547
rect 4340 7513 4396 7547
rect 3858 7493 4396 7513
rect 4456 7547 4994 7561
rect 4456 7513 4512 7547
rect 4546 7513 4592 7547
rect 4626 7513 4672 7547
rect 4706 7513 4752 7547
rect 4786 7513 4832 7547
rect 4866 7513 4912 7547
rect 4946 7513 4994 7547
rect 4456 7493 4994 7513
rect 5070 7547 5608 7561
rect 5070 7513 5118 7547
rect 5152 7513 5198 7547
rect 5232 7513 5278 7547
rect 5312 7513 5358 7547
rect 5392 7513 5438 7547
rect 5472 7513 5518 7547
rect 5552 7513 5608 7547
rect 5070 7493 5608 7513
rect 5668 7547 6206 7561
rect 5668 7513 5724 7547
rect 5758 7513 5804 7547
rect 5838 7513 5884 7547
rect 5918 7513 5964 7547
rect 5998 7513 6044 7547
rect 6078 7513 6124 7547
rect 6158 7513 6206 7547
rect 5668 7493 6206 7513
rect 6282 7547 6820 7561
rect 6282 7513 6330 7547
rect 6364 7513 6410 7547
rect 6444 7513 6490 7547
rect 6524 7513 6570 7547
rect 6604 7513 6650 7547
rect 6684 7513 6730 7547
rect 6764 7513 6820 7547
rect 6282 7493 6820 7513
rect 6880 7547 7418 7561
rect 6880 7513 6936 7547
rect 6970 7513 7016 7547
rect 7050 7513 7096 7547
rect 7130 7513 7176 7547
rect 7210 7513 7256 7547
rect 7290 7513 7336 7547
rect 7370 7513 7418 7547
rect 6880 7493 7418 7513
rect 7494 7547 8032 7561
rect 7494 7513 7542 7547
rect 7576 7513 7622 7547
rect 7656 7513 7702 7547
rect 7736 7513 7782 7547
rect 7816 7513 7862 7547
rect 7896 7513 7942 7547
rect 7976 7513 8032 7547
rect 7494 7493 8032 7513
rect 8092 7547 8630 7561
rect 8092 7513 8148 7547
rect 8182 7513 8228 7547
rect 8262 7513 8308 7547
rect 8342 7513 8388 7547
rect 8422 7513 8468 7547
rect 8502 7513 8548 7547
rect 8582 7513 8630 7547
rect 8862 7538 8948 7564
rect 8092 7493 8630 7513
rect 13343 7552 13369 7586
rect 13403 7552 13429 7586
rect 13343 7526 13429 7552
rect 13661 7535 14199 7549
rect 13661 7501 13709 7535
rect 13743 7501 13789 7535
rect 13823 7501 13869 7535
rect 13903 7501 13949 7535
rect 13983 7501 14029 7535
rect 14063 7501 14109 7535
rect 14143 7501 14199 7535
rect 13661 7481 14199 7501
rect 14259 7535 14797 7549
rect 14259 7501 14315 7535
rect 14349 7501 14395 7535
rect 14429 7501 14475 7535
rect 14509 7501 14555 7535
rect 14589 7501 14635 7535
rect 14669 7501 14715 7535
rect 14749 7501 14797 7535
rect 14259 7481 14797 7501
rect 14873 7535 15411 7549
rect 14873 7501 14921 7535
rect 14955 7501 15001 7535
rect 15035 7501 15081 7535
rect 15115 7501 15161 7535
rect 15195 7501 15241 7535
rect 15275 7501 15321 7535
rect 15355 7501 15411 7535
rect 14873 7481 15411 7501
rect 15471 7535 16009 7549
rect 15471 7501 15527 7535
rect 15561 7501 15607 7535
rect 15641 7501 15687 7535
rect 15721 7501 15767 7535
rect 15801 7501 15847 7535
rect 15881 7501 15927 7535
rect 15961 7501 16009 7535
rect 15471 7481 16009 7501
rect 16085 7535 16623 7549
rect 16085 7501 16133 7535
rect 16167 7501 16213 7535
rect 16247 7501 16293 7535
rect 16327 7501 16373 7535
rect 16407 7501 16453 7535
rect 16487 7501 16533 7535
rect 16567 7501 16623 7535
rect 16085 7481 16623 7501
rect 16683 7535 17221 7549
rect 16683 7501 16739 7535
rect 16773 7501 16819 7535
rect 16853 7501 16899 7535
rect 16933 7501 16979 7535
rect 17013 7501 17059 7535
rect 17093 7501 17139 7535
rect 17173 7501 17221 7535
rect 16683 7481 17221 7501
rect 17297 7535 17835 7549
rect 17297 7501 17345 7535
rect 17379 7501 17425 7535
rect 17459 7501 17505 7535
rect 17539 7501 17585 7535
rect 17619 7501 17665 7535
rect 17699 7501 17745 7535
rect 17779 7501 17835 7535
rect 17297 7481 17835 7501
rect 17895 7535 18433 7549
rect 17895 7501 17951 7535
rect 17985 7501 18031 7535
rect 18065 7501 18111 7535
rect 18145 7501 18191 7535
rect 18225 7501 18271 7535
rect 18305 7501 18351 7535
rect 18385 7501 18433 7535
rect 17895 7481 18433 7501
rect 18627 7538 19165 7552
rect 18627 7504 18683 7538
rect 18717 7504 18763 7538
rect 18797 7504 18843 7538
rect 18877 7504 18923 7538
rect 18957 7504 19003 7538
rect 19037 7504 19083 7538
rect 19117 7504 19165 7538
rect 19624 7575 19650 7609
rect 19684 7575 19710 7609
rect 19624 7549 19710 7575
rect 20052 7586 20138 7612
rect 20052 7552 20078 7586
rect 20112 7552 20138 7586
rect 20052 7526 20138 7552
rect 20370 7535 20908 7549
rect 18627 7484 19165 7504
rect 20370 7501 20418 7535
rect 20452 7501 20498 7535
rect 20532 7501 20578 7535
rect 20612 7501 20658 7535
rect 20692 7501 20738 7535
rect 20772 7501 20818 7535
rect 20852 7501 20908 7535
rect 20370 7481 20908 7501
rect 20968 7535 21506 7549
rect 20968 7501 21024 7535
rect 21058 7501 21104 7535
rect 21138 7501 21184 7535
rect 21218 7501 21264 7535
rect 21298 7501 21344 7535
rect 21378 7501 21424 7535
rect 21458 7501 21506 7535
rect 20968 7481 21506 7501
rect 21582 7535 22120 7549
rect 21582 7501 21630 7535
rect 21664 7501 21710 7535
rect 21744 7501 21790 7535
rect 21824 7501 21870 7535
rect 21904 7501 21950 7535
rect 21984 7501 22030 7535
rect 22064 7501 22120 7535
rect 21582 7481 22120 7501
rect 22180 7535 22718 7549
rect 22180 7501 22236 7535
rect 22270 7501 22316 7535
rect 22350 7501 22396 7535
rect 22430 7501 22476 7535
rect 22510 7501 22556 7535
rect 22590 7501 22636 7535
rect 22670 7501 22718 7535
rect 22180 7481 22718 7501
rect 22794 7535 23332 7549
rect 22794 7501 22842 7535
rect 22876 7501 22922 7535
rect 22956 7501 23002 7535
rect 23036 7501 23082 7535
rect 23116 7501 23162 7535
rect 23196 7501 23242 7535
rect 23276 7501 23332 7535
rect 22794 7481 23332 7501
rect 23392 7535 23930 7549
rect 23392 7501 23448 7535
rect 23482 7501 23528 7535
rect 23562 7501 23608 7535
rect 23642 7501 23688 7535
rect 23722 7501 23768 7535
rect 23802 7501 23848 7535
rect 23882 7501 23930 7535
rect 23392 7481 23930 7501
rect 24006 7535 24544 7549
rect 24006 7501 24054 7535
rect 24088 7501 24134 7535
rect 24168 7501 24214 7535
rect 24248 7501 24294 7535
rect 24328 7501 24374 7535
rect 24408 7501 24454 7535
rect 24488 7501 24544 7535
rect 24006 7481 24544 7501
rect 24604 7535 25142 7549
rect 24604 7501 24660 7535
rect 24694 7501 24740 7535
rect 24774 7501 24820 7535
rect 24854 7501 24900 7535
rect 24934 7501 24980 7535
rect 25014 7501 25060 7535
rect 25094 7501 25142 7535
rect 24604 7481 25142 7501
rect 25336 7538 25874 7552
rect 25336 7504 25392 7538
rect 25426 7504 25472 7538
rect 25506 7504 25552 7538
rect 25586 7504 25632 7538
rect 25666 7504 25712 7538
rect 25746 7504 25792 7538
rect 25826 7504 25874 7538
rect 25336 7484 25874 7504
rect 24739 7308 25277 7328
rect 24739 7274 24787 7308
rect 24821 7274 24867 7308
rect 24901 7274 24947 7308
rect 24981 7274 25027 7308
rect 25061 7274 25107 7308
rect 25141 7274 25187 7308
rect 25221 7274 25277 7308
rect 24739 7260 25277 7274
rect 25471 7311 26009 7331
rect 25471 7277 25519 7311
rect 25553 7277 25599 7311
rect 25633 7277 25679 7311
rect 25713 7277 25759 7311
rect 25793 7277 25839 7311
rect 25873 7277 25919 7311
rect 25953 7277 26009 7311
rect 25471 7263 26009 7277
rect 26069 7311 26607 7331
rect 26069 7277 26125 7311
rect 26159 7277 26205 7311
rect 26239 7277 26285 7311
rect 26319 7277 26365 7311
rect 26399 7277 26445 7311
rect 26479 7277 26525 7311
rect 26559 7277 26607 7311
rect 26069 7263 26607 7277
rect 26683 7311 27221 7331
rect 26683 7277 26731 7311
rect 26765 7277 26811 7311
rect 26845 7277 26891 7311
rect 26925 7277 26971 7311
rect 27005 7277 27051 7311
rect 27085 7277 27131 7311
rect 27165 7277 27221 7311
rect 26683 7263 27221 7277
rect 27281 7311 27819 7331
rect 27281 7277 27337 7311
rect 27371 7277 27417 7311
rect 27451 7277 27497 7311
rect 27531 7277 27577 7311
rect 27611 7277 27657 7311
rect 27691 7277 27737 7311
rect 27771 7277 27819 7311
rect 27281 7263 27819 7277
rect 27895 7311 28433 7331
rect 27895 7277 27943 7311
rect 27977 7277 28023 7311
rect 28057 7277 28103 7311
rect 28137 7277 28183 7311
rect 28217 7277 28263 7311
rect 28297 7277 28343 7311
rect 28377 7277 28433 7311
rect 27895 7263 28433 7277
rect 28493 7311 29031 7331
rect 28493 7277 28549 7311
rect 28583 7277 28629 7311
rect 28663 7277 28709 7311
rect 28743 7277 28789 7311
rect 28823 7277 28869 7311
rect 28903 7277 28949 7311
rect 28983 7277 29031 7311
rect 28493 7263 29031 7277
rect 29107 7311 29645 7331
rect 29107 7277 29155 7311
rect 29189 7277 29235 7311
rect 29269 7277 29315 7311
rect 29349 7277 29395 7311
rect 29429 7277 29475 7311
rect 29509 7277 29555 7311
rect 29589 7277 29645 7311
rect 29107 7263 29645 7277
rect 29705 7311 30243 7331
rect 29705 7277 29761 7311
rect 29795 7277 29841 7311
rect 29875 7277 29921 7311
rect 29955 7277 30001 7311
rect 30035 7277 30081 7311
rect 30115 7277 30161 7311
rect 30195 7277 30243 7311
rect 29705 7263 30243 7277
rect 30475 7260 30561 7286
rect 30475 7226 30501 7260
rect 30535 7226 30561 7260
rect 30475 7200 30561 7226
rect 11498 7084 11527 7118
rect 11561 7084 11619 7118
rect 11653 7084 11711 7118
rect 11745 7084 11803 7118
rect 11837 7084 11895 7118
rect 11929 7084 11987 7118
rect 12021 7084 12079 7118
rect 12113 7084 12142 7118
rect 12758 7084 12787 7118
rect 12821 7084 12879 7118
rect 12913 7084 12971 7118
rect 13005 7084 13063 7118
rect 13097 7084 13155 7118
rect 13189 7084 13247 7118
rect 13281 7084 13339 7118
rect 13373 7084 13431 7118
rect 13465 7084 13523 7118
rect 13557 7084 13615 7118
rect 13649 7084 13707 7118
rect 13741 7084 13799 7118
rect 13833 7084 13891 7118
rect 13925 7084 13983 7118
rect 14017 7084 14075 7118
rect 14109 7084 14167 7118
rect 14201 7084 14259 7118
rect 14293 7084 14351 7118
rect 14385 7084 14443 7118
rect 14477 7084 14535 7118
rect 14569 7084 14598 7118
rect 24729 7130 24812 7155
rect 24729 7095 24754 7130
rect 24788 7095 24812 7130
rect 24729 7071 24812 7095
rect 30480 7116 30566 7142
rect 30480 7082 30506 7116
rect 30540 7082 30566 7116
rect 30480 7056 30566 7082
rect 30481 6964 30567 6990
rect 30481 6930 30507 6964
rect 30541 6930 30567 6964
rect 30481 6904 30567 6930
rect 30481 6794 30567 6820
rect 30481 6760 30507 6794
rect 30541 6760 30567 6794
rect 24043 6742 24459 6744
rect 24043 6708 24073 6742
rect 24107 6708 24203 6742
rect 24237 6708 24349 6742
rect 24383 6708 24459 6742
rect 24043 6704 24459 6708
rect 30481 6734 30567 6760
rect 30480 6637 30566 6663
rect 30480 6603 30506 6637
rect 30540 6603 30566 6637
rect 30480 6577 30566 6603
rect 30679 6369 31048 6371
rect 30679 6335 30708 6369
rect 30742 6335 30891 6369
rect 30925 6335 31048 6369
rect 11497 6211 11526 6245
rect 11560 6211 11618 6245
rect 11652 6211 11710 6245
rect 11744 6211 11802 6245
rect 11836 6211 11894 6245
rect 11928 6211 11986 6245
rect 12020 6211 12078 6245
rect 12112 6211 12170 6245
rect 12204 6211 12262 6245
rect 12296 6211 12354 6245
rect 12388 6211 12446 6245
rect 12480 6211 12538 6245
rect 12572 6211 12630 6245
rect 12664 6211 12722 6245
rect 12756 6211 12814 6245
rect 12848 6211 12906 6245
rect 12940 6211 12998 6245
rect 13032 6211 13090 6245
rect 13124 6211 13182 6245
rect 13216 6211 13274 6245
rect 13308 6211 13358 6245
rect 13470 6211 13550 6245
rect 13584 6211 13642 6245
rect 13676 6211 13734 6245
rect 13768 6211 13826 6245
rect 13860 6211 13918 6245
rect 13952 6211 14010 6245
rect 14044 6211 14103 6245
rect 14137 6211 14194 6245
rect 14228 6211 14286 6245
rect 14320 6211 14378 6245
rect 14412 6211 14470 6245
rect 14504 6211 14602 6245
rect 14712 6211 14746 6245
rect 14780 6211 14838 6245
rect 14872 6211 14930 6245
rect 14964 6211 15022 6245
rect 15056 6211 15114 6245
rect 15148 6211 15206 6245
rect 15240 6211 15298 6245
rect 15332 6211 15390 6245
rect 15424 6211 15482 6245
rect 15516 6211 15574 6245
rect 15608 6211 15666 6245
rect 15700 6211 15758 6245
rect 15792 6211 15850 6245
rect 15884 6211 15942 6245
rect 15976 6211 16034 6245
rect 16068 6211 16126 6245
rect 16160 6211 16218 6245
rect 16252 6211 16310 6245
rect 16344 6211 16402 6245
rect 16436 6211 16494 6245
rect 16528 6211 16586 6245
rect 16620 6211 16678 6245
rect 16712 6211 16770 6245
rect 16804 6211 16862 6245
rect 16896 6211 16994 6245
rect 17104 6211 17138 6245
rect 17172 6211 17230 6245
rect 17264 6211 17322 6245
rect 17356 6211 17414 6245
rect 17448 6211 17506 6245
rect 17540 6211 17598 6245
rect 17632 6211 17690 6245
rect 17724 6211 17782 6245
rect 17816 6211 17874 6245
rect 17908 6211 17966 6245
rect 18000 6211 18058 6245
rect 18092 6211 18150 6245
rect 18184 6211 18242 6245
rect 18276 6211 18334 6245
rect 18368 6211 18426 6245
rect 18460 6211 18518 6245
rect 18552 6211 18610 6245
rect 18644 6211 18702 6245
rect 18736 6211 18794 6245
rect 18828 6211 18886 6245
rect 18920 6211 18978 6245
rect 19012 6211 19070 6245
rect 19104 6211 19162 6245
rect 19196 6211 19254 6245
rect 19288 6211 19386 6245
rect 19496 6211 19530 6245
rect 19564 6211 19622 6245
rect 19656 6211 19714 6245
rect 19748 6211 19806 6245
rect 19840 6211 19898 6245
rect 19932 6211 19990 6245
rect 20024 6211 20082 6245
rect 20116 6211 20174 6245
rect 20208 6211 20266 6245
rect 20300 6211 20358 6245
rect 20392 6211 20450 6245
rect 20484 6211 20542 6245
rect 20576 6211 20634 6245
rect 20668 6211 20726 6245
rect 20760 6211 20818 6245
rect 20852 6211 20910 6245
rect 20944 6211 21002 6245
rect 21036 6211 21094 6245
rect 21128 6211 21186 6245
rect 21220 6211 21278 6245
rect 21312 6211 21370 6245
rect 21404 6211 21462 6245
rect 21496 6211 21554 6245
rect 21588 6211 21646 6245
rect 21680 6211 21778 6245
rect 21888 6211 21922 6245
rect 21956 6211 22014 6245
rect 22048 6211 22106 6245
rect 22140 6211 22198 6245
rect 22232 6211 22290 6245
rect 22324 6211 22382 6245
rect 22416 6211 22474 6245
rect 22508 6211 22566 6245
rect 22600 6211 22658 6245
rect 22692 6211 22750 6245
rect 22784 6211 22842 6245
rect 22876 6211 22934 6245
rect 22968 6211 23026 6245
rect 23060 6211 23118 6245
rect 23152 6211 23210 6245
rect 23244 6211 23302 6245
rect 23336 6211 23394 6245
rect 23428 6211 23457 6245
rect 11057 5522 11086 5556
rect 11120 5522 11178 5556
rect 11212 5522 11270 5556
rect 11304 5522 11362 5556
rect 11396 5522 11454 5556
rect 11488 5522 11546 5556
rect 11580 5522 11638 5556
rect 11672 5522 11730 5556
rect 11764 5522 11822 5556
rect 11856 5522 11914 5556
rect 11948 5522 12006 5556
rect 12040 5522 12098 5556
rect 12132 5522 12190 5556
rect 12224 5522 12282 5556
rect 12316 5522 12374 5556
rect 12408 5522 12466 5556
rect 12500 5522 12558 5556
rect 12592 5522 12650 5556
rect 12684 5522 12742 5556
rect 12776 5522 12814 5556
rect 12868 5522 12906 5556
rect 12940 5522 12998 5556
rect 13032 5522 13090 5556
rect 13124 5522 13182 5556
rect 13216 5522 13274 5556
rect 13308 5522 13366 5556
rect 13400 5522 13458 5556
rect 13492 5522 13550 5556
rect 13584 5522 13642 5556
rect 13676 5522 13734 5556
rect 13768 5522 13826 5556
rect 13860 5522 13918 5556
rect 13952 5522 14010 5556
rect 14044 5522 14102 5556
rect 14136 5522 14194 5556
rect 14228 5522 14286 5556
rect 14320 5522 14378 5556
rect 14412 5522 14470 5556
rect 14504 5522 14562 5556
rect 14596 5522 14673 5556
rect 14783 5522 14838 5556
rect 14872 5522 14930 5556
rect 14964 5522 15022 5556
rect 15056 5522 15114 5556
rect 15148 5522 15206 5556
rect 15240 5522 15298 5556
rect 15332 5522 15390 5556
rect 15424 5522 15482 5556
rect 15516 5522 15574 5556
rect 15608 5522 15666 5556
rect 15700 5522 15758 5556
rect 15792 5522 15850 5556
rect 15884 5522 15942 5556
rect 15976 5522 16034 5556
rect 16068 5522 16126 5556
rect 16160 5522 16218 5556
rect 16252 5522 16310 5556
rect 16344 5522 16402 5556
rect 16436 5522 16494 5556
rect 16528 5522 16586 5556
rect 16620 5522 16678 5556
rect 16712 5522 16770 5556
rect 16804 5522 16862 5556
rect 16896 5522 16954 5556
rect 16988 5522 17065 5556
rect 17175 5522 17230 5556
rect 17264 5522 17322 5556
rect 17356 5522 17414 5556
rect 17448 5522 17506 5556
rect 17540 5522 17598 5556
rect 17632 5522 17690 5556
rect 17724 5522 17782 5556
rect 17816 5522 17874 5556
rect 17908 5522 17966 5556
rect 18000 5522 18058 5556
rect 18092 5522 18150 5556
rect 18184 5522 18242 5556
rect 18276 5522 18334 5556
rect 18368 5522 18426 5556
rect 18460 5522 18518 5556
rect 18552 5522 18610 5556
rect 18644 5522 18702 5556
rect 18736 5522 18794 5556
rect 18828 5522 18886 5556
rect 18920 5522 18978 5556
rect 19012 5522 19070 5556
rect 19104 5522 19162 5556
rect 19196 5522 19254 5556
rect 19288 5522 19346 5556
rect 19380 5522 19457 5556
rect 19567 5522 19622 5556
rect 19656 5522 19714 5556
rect 19748 5522 19806 5556
rect 19840 5522 19898 5556
rect 19932 5522 19990 5556
rect 20024 5522 20082 5556
rect 20116 5522 20174 5556
rect 20208 5522 20266 5556
rect 20300 5522 20358 5556
rect 20392 5522 20450 5556
rect 20484 5522 20542 5556
rect 20576 5522 20634 5556
rect 20668 5522 20726 5556
rect 20760 5522 20818 5556
rect 20852 5522 20910 5556
rect 20944 5522 21002 5556
rect 21036 5522 21094 5556
rect 21128 5522 21186 5556
rect 21220 5522 21278 5556
rect 21312 5522 21370 5556
rect 21404 5522 21462 5556
rect 21496 5522 21554 5556
rect 21588 5522 21646 5556
rect 21680 5522 21738 5556
rect 21772 5522 21849 5556
rect 21959 5522 22014 5556
rect 22048 5522 22106 5556
rect 22140 5522 22198 5556
rect 22232 5522 22290 5556
rect 22324 5522 22382 5556
rect 22416 5522 22474 5556
rect 22508 5522 22566 5556
rect 22600 5522 22658 5556
rect 22692 5522 22750 5556
rect 22784 5522 22842 5556
rect 22876 5522 22934 5556
rect 22968 5522 23026 5556
rect 23060 5522 23118 5556
rect 23152 5522 23210 5556
rect 23244 5522 23302 5556
rect 23336 5522 23394 5556
rect 23428 5522 23459 5556
rect 11089 4658 11118 4692
rect 11152 4658 11210 4692
rect 11244 4658 11302 4692
rect 11336 4658 11394 4692
rect 11428 4658 11486 4692
rect 11520 4658 11577 4692
rect 11611 4658 11669 4692
rect 11703 4658 11762 4692
rect 11796 4658 11854 4692
rect 11888 4658 11918 4692
rect 11089 4657 11918 4658
rect 13631 4649 13660 4683
rect 13694 4649 13752 4683
rect 13786 4649 13844 4683
rect 13878 4649 13936 4683
rect 13970 4649 14028 4683
rect 14062 4649 14120 4683
rect 14154 4649 14212 4683
rect 14246 4649 14304 4683
rect 14338 4649 14396 4683
rect 14430 4649 14488 4683
rect 14522 4649 14580 4683
rect 14614 4649 14672 4683
rect 14706 4649 14764 4683
rect 14798 4649 14856 4683
rect 14890 4649 14948 4683
rect 14982 4649 15040 4683
rect 15074 4649 15132 4683
rect 15166 4649 15224 4683
rect 15258 4649 15316 4683
rect 15350 4649 15408 4683
rect 15442 4649 15481 4683
rect 15515 4649 15573 4683
rect 15607 4649 15665 4683
rect 15699 4649 15757 4683
rect 15791 4649 15849 4683
rect 15883 4649 15941 4683
rect 15975 4649 16033 4683
rect 16067 4649 16125 4683
rect 16159 4649 16217 4683
rect 16251 4649 16309 4683
rect 16343 4649 16401 4683
rect 16435 4649 16493 4683
rect 16527 4649 16585 4683
rect 16619 4649 16677 4683
rect 16711 4649 16769 4683
rect 16803 4649 16861 4683
rect 16895 4649 16953 4683
rect 16987 4649 17045 4683
rect 17079 4649 17137 4683
rect 17171 4649 17229 4683
rect 17263 4649 17321 4683
rect 17355 4649 17413 4683
rect 17447 4649 17505 4683
rect 17539 4649 17597 4683
rect 17631 4649 17689 4683
rect 17723 4649 17781 4683
rect 17815 4649 17873 4683
rect 17907 4649 17965 4683
rect 17999 4649 18057 4683
rect 18091 4649 18149 4683
rect 18183 4649 18241 4683
rect 18275 4649 18333 4683
rect 18367 4649 18425 4683
rect 18459 4649 18517 4683
rect 18551 4649 18609 4683
rect 18643 4649 18701 4683
rect 18735 4649 18793 4683
rect 18827 4649 18885 4683
rect 18919 4649 18977 4683
rect 19011 4649 19069 4683
rect 19103 4649 19161 4683
rect 19195 4649 19253 4683
rect 19287 4649 19345 4683
rect 19379 4649 19437 4683
rect 19471 4649 19529 4683
rect 19563 4649 19621 4683
rect 19655 4649 19713 4683
rect 19747 4649 19805 4683
rect 19839 4649 19897 4683
rect 19931 4649 19989 4683
rect 20023 4649 20081 4683
rect 20115 4649 20173 4683
rect 20207 4649 20265 4683
rect 20299 4649 20357 4683
rect 20391 4649 20449 4683
rect 20483 4649 20541 4683
rect 20575 4649 20633 4683
rect 20667 4649 20725 4683
rect 20759 4649 20817 4683
rect 20851 4649 20909 4683
rect 20943 4649 21001 4683
rect 21035 4649 21093 4683
rect 21127 4649 21185 4683
rect 21219 4649 21277 4683
rect 21311 4649 21369 4683
rect 21403 4649 21461 4683
rect 21495 4649 21553 4683
rect 21587 4649 21645 4683
rect 21679 4649 21737 4683
rect 21771 4649 21829 4683
rect 21863 4649 21921 4683
rect 21955 4649 22013 4683
rect 22047 4649 22105 4683
rect 22139 4649 22197 4683
rect 22231 4649 22289 4683
rect 22323 4649 22381 4683
rect 22415 4649 22473 4683
rect 22507 4649 22565 4683
rect 22599 4649 22657 4683
rect 22691 4649 22749 4683
rect 22783 4649 22841 4683
rect 22875 4649 22933 4683
rect 22967 4649 23025 4683
rect 23059 4649 23117 4683
rect 23151 4649 23209 4683
rect 23243 4649 23301 4683
rect 23335 4649 23393 4683
rect 23427 4649 23456 4683
rect 11496 3776 11525 3810
rect 11559 3776 11617 3810
rect 11651 3776 11709 3810
rect 11743 3776 11801 3810
rect 11835 3776 11893 3810
rect 11927 3776 11985 3810
rect 12019 3776 12077 3810
rect 12111 3776 12169 3810
rect 12203 3776 12261 3810
rect 12295 3776 12353 3810
rect 12387 3776 12445 3810
rect 12479 3776 12537 3810
rect 12571 3776 12629 3810
rect 12663 3776 12721 3810
rect 12755 3776 12813 3810
rect 12847 3776 12905 3810
rect 12939 3776 12997 3810
rect 13031 3776 13089 3810
rect 13123 3776 13181 3810
rect 13215 3776 13273 3810
rect 13307 3776 13365 3810
rect 13399 3776 13457 3810
rect 13491 3776 13549 3810
rect 13583 3776 13641 3810
rect 13675 3776 13733 3810
rect 13767 3776 13825 3810
rect 13859 3776 13917 3810
rect 13951 3776 14009 3810
rect 14043 3776 14101 3810
rect 14135 3776 14193 3810
rect 14227 3776 14285 3810
rect 14319 3776 14377 3810
rect 14411 3776 14469 3810
rect 14503 3776 14561 3810
rect 14595 3776 14653 3810
rect 14687 3776 14745 3810
rect 14779 3776 14837 3810
rect 14871 3776 14929 3810
rect 14963 3776 15021 3810
rect 15055 3776 15113 3810
rect 15147 3776 15205 3810
rect 15239 3776 15297 3810
rect 15331 3776 15389 3810
rect 15423 3776 15481 3810
rect 15515 3776 15573 3810
rect 15607 3776 15665 3810
rect 15699 3776 15757 3810
rect 15791 3776 15849 3810
rect 15883 3776 15941 3810
rect 15975 3776 16033 3810
rect 16067 3776 16125 3810
rect 16159 3776 16217 3810
rect 16251 3776 16309 3810
rect 16343 3776 16401 3810
rect 16435 3776 16493 3810
rect 16527 3776 16585 3810
rect 16619 3776 16677 3810
rect 16711 3776 16769 3810
rect 16803 3776 16861 3810
rect 16895 3776 16953 3810
rect 16987 3776 17045 3810
rect 17079 3776 17137 3810
rect 17171 3776 17229 3810
rect 17263 3776 17321 3810
rect 17355 3776 17413 3810
rect 17447 3776 17505 3810
rect 17539 3776 17597 3810
rect 17631 3776 17689 3810
rect 17723 3776 17781 3810
rect 17815 3776 17873 3810
rect 17907 3776 17965 3810
rect 17999 3776 18057 3810
rect 18091 3776 18149 3810
rect 18183 3776 18241 3810
rect 18275 3776 18333 3810
rect 18367 3776 18425 3810
rect 18459 3776 18517 3810
rect 18551 3776 18609 3810
rect 18643 3776 18701 3810
rect 18735 3776 18793 3810
rect 18827 3776 18885 3810
rect 18919 3776 18977 3810
rect 19011 3776 19069 3810
rect 19103 3776 19161 3810
rect 19195 3776 19253 3810
rect 19287 3776 19345 3810
rect 19379 3776 19437 3810
rect 19471 3776 19529 3810
rect 19563 3776 19621 3810
rect 19655 3776 19713 3810
rect 19747 3776 19805 3810
rect 19839 3776 19897 3810
rect 19931 3776 19989 3810
rect 20023 3776 20081 3810
rect 20115 3776 20173 3810
rect 20207 3776 20265 3810
rect 20299 3776 20357 3810
rect 20391 3776 20449 3810
rect 20483 3776 20541 3810
rect 20575 3776 20633 3810
rect 20667 3776 20725 3810
rect 20759 3776 20817 3810
rect 20851 3776 20909 3810
rect 20943 3776 21001 3810
rect 21035 3776 21093 3810
rect 21127 3776 21185 3810
rect 21219 3776 21277 3810
rect 21311 3776 21369 3810
rect 21403 3776 21461 3810
rect 21495 3776 21553 3810
rect 21587 3776 21645 3810
rect 21679 3776 21737 3810
rect 21771 3776 21829 3810
rect 21863 3776 21921 3810
rect 21955 3776 22013 3810
rect 22047 3776 22105 3810
rect 22139 3776 22197 3810
rect 22231 3776 22289 3810
rect 22323 3776 22381 3810
rect 22415 3776 22473 3810
rect 22507 3776 22565 3810
rect 22599 3776 22657 3810
rect 22691 3776 22749 3810
rect 22783 3776 22841 3810
rect 22875 3776 22933 3810
rect 22967 3776 23025 3810
rect 23059 3776 23117 3810
rect 23151 3776 23209 3810
rect 23243 3776 23301 3810
rect 23335 3776 23393 3810
rect 23427 3776 23456 3810
rect 25577 3672 25607 3706
rect 25641 3672 25698 3706
rect 25732 3672 25791 3706
rect 25825 3672 25882 3706
rect 25916 3672 25973 3706
rect 26007 3672 26067 3706
rect 26101 3672 26158 3706
rect 26192 3672 26251 3706
rect 26285 3672 26342 3706
rect 26376 3672 26434 3706
rect 26468 3672 26525 3706
rect 26559 3672 26618 3706
rect 26652 3672 26711 3706
rect 26745 3672 26802 3706
rect 26836 3672 26894 3706
rect 26928 3672 26986 3706
rect 27020 3672 27078 3706
rect 27112 3672 27170 3706
rect 27204 3672 27262 3706
rect 27296 3672 27354 3706
rect 27388 3672 27447 3706
rect 27481 3672 27537 3706
rect 27571 3672 27630 3706
rect 27664 3672 27723 3706
rect 27757 3672 27815 3706
rect 27849 3672 27906 3706
rect 27940 3672 27999 3706
rect 28033 3672 28091 3706
rect 28125 3672 28183 3706
rect 28217 3672 28275 3706
rect 28309 3672 28367 3706
rect 28401 3672 28459 3706
rect 28493 3672 28550 3706
rect 28584 3672 28641 3706
rect 28675 3672 28734 3706
rect 28768 3672 28827 3706
rect 28861 3672 28919 3706
rect 28953 3672 29010 3706
rect 29044 3672 29104 3706
rect 29138 3672 29194 3706
rect 29228 3672 29285 3706
rect 29319 3672 29378 3706
rect 29412 3672 29471 3706
rect 29505 3672 29563 3706
rect 29597 3672 29654 3706
rect 29688 3672 29746 3706
rect 29780 3672 29838 3706
rect 29872 3672 29929 3706
rect 29963 3672 30021 3706
rect 30055 3672 30114 3706
rect 30148 3672 30206 3706
rect 30240 3672 30298 3706
rect 30332 3672 30361 3706
rect 25577 2391 25609 2425
rect 25643 2391 25699 2425
rect 25733 2391 25792 2425
rect 25826 2391 25882 2425
rect 25916 2391 25973 2425
rect 26007 2391 26067 2425
rect 26101 2391 26158 2425
rect 26192 2391 26250 2425
rect 26284 2391 26342 2425
rect 26376 2391 26435 2425
rect 26469 2391 26526 2425
rect 26560 2391 26618 2425
rect 26652 2391 26710 2425
rect 26744 2391 26802 2425
rect 26836 2391 26895 2425
rect 26929 2391 26986 2425
rect 27020 2391 27077 2425
rect 27111 2391 27170 2425
rect 27204 2391 27263 2425
rect 27297 2391 27354 2425
rect 27388 2391 27446 2425
rect 27480 2391 27538 2425
rect 27572 2391 27630 2425
rect 27664 2391 27723 2425
rect 27757 2391 27813 2425
rect 27847 2391 27906 2425
rect 27940 2391 27998 2425
rect 28032 2391 28091 2425
rect 28125 2391 28185 2425
rect 28219 2391 28274 2425
rect 28308 2391 28366 2425
rect 28400 2391 28458 2425
rect 28492 2391 28550 2425
rect 28584 2391 28642 2425
rect 28676 2391 28734 2425
rect 28768 2391 28826 2425
rect 28860 2391 28918 2425
rect 28952 2391 29010 2425
rect 29044 2391 29102 2425
rect 29136 2391 29194 2425
rect 29228 2391 29286 2425
rect 29320 2391 29378 2425
rect 29412 2391 29470 2425
rect 29504 2391 29562 2425
rect 29596 2391 29654 2425
rect 29688 2391 29746 2425
rect 29780 2391 29838 2425
rect 29872 2391 29930 2425
rect 29964 2391 30022 2425
rect 30056 2391 30114 2425
rect 30148 2391 30207 2425
rect 30241 2391 30298 2425
rect 30332 2391 30361 2425
rect 8577 1396 8606 1430
rect 8640 1396 8698 1430
rect 8732 1396 8790 1430
rect 8824 1396 8882 1430
rect 8916 1396 8974 1430
rect 9008 1396 9066 1430
rect 9100 1396 9158 1430
rect 9192 1396 9250 1430
rect 9284 1396 9342 1430
rect 9376 1396 9434 1430
rect 9468 1396 9526 1430
rect 9560 1396 9618 1430
rect 9652 1396 9710 1430
rect 9744 1396 9802 1430
rect 9836 1396 9894 1430
rect 9928 1396 9986 1430
rect 10020 1396 10078 1430
rect 10112 1396 10170 1430
rect 10204 1396 10262 1430
rect 10296 1396 10354 1430
rect 10388 1396 10446 1430
rect 10480 1396 10538 1430
rect 10572 1396 10630 1430
rect 10664 1396 10722 1430
rect 10756 1396 10814 1430
rect 10848 1396 10906 1430
rect 10940 1396 10998 1430
rect 11032 1396 11090 1430
rect 11124 1396 11182 1430
rect 11216 1396 11274 1430
rect 11308 1396 11366 1430
rect 11400 1396 11429 1430
rect 12961 1396 12990 1430
rect 13024 1396 13082 1430
rect 13116 1396 13174 1430
rect 13208 1396 13266 1430
rect 13300 1396 13358 1430
rect 13392 1396 13450 1430
rect 13484 1396 13542 1430
rect 13576 1396 13634 1430
rect 13668 1396 13726 1430
rect 13760 1396 13818 1430
rect 13852 1396 13910 1430
rect 13944 1396 14002 1430
rect 14036 1396 14094 1430
rect 14128 1396 14186 1430
rect 14220 1396 14278 1430
rect 14312 1396 14370 1430
rect 14404 1396 14462 1430
rect 14496 1396 14554 1430
rect 14588 1396 14646 1430
rect 14680 1396 14738 1430
rect 14772 1396 14830 1430
rect 14864 1396 14922 1430
rect 14956 1396 15014 1430
rect 15048 1396 15106 1430
rect 15140 1396 15198 1430
rect 15232 1396 15290 1430
rect 15324 1396 15382 1430
rect 15416 1396 15474 1430
rect 15508 1396 15566 1430
rect 15600 1396 15658 1430
rect 15692 1396 15750 1430
rect 15784 1396 15813 1430
rect 8575 254 8604 288
rect 8638 254 8696 288
rect 8730 254 8788 288
rect 8822 254 8880 288
rect 8914 254 8972 288
rect 9006 254 9064 288
rect 9098 254 9156 288
rect 9190 254 9248 288
rect 9282 254 9340 288
rect 9374 254 9432 288
rect 9466 254 9524 288
rect 9558 254 9616 288
rect 9650 254 9708 288
rect 9742 254 9800 288
rect 9834 254 9892 288
rect 9926 254 9984 288
rect 10018 254 10076 288
rect 10110 254 10168 288
rect 10202 254 10260 288
rect 10294 254 10352 288
rect 10386 254 10444 288
rect 10478 254 10536 288
rect 10570 254 10628 288
rect 10662 254 10720 288
rect 10754 254 10812 288
rect 10846 254 10904 288
rect 10938 254 10996 288
rect 11030 254 11088 288
rect 11122 254 11180 288
rect 11214 254 11272 288
rect 11306 254 11364 288
rect 11398 254 11456 288
rect 11490 254 11548 288
rect 11582 254 11640 288
rect 11674 254 11732 288
rect 11766 254 11824 288
rect 11858 254 11916 288
rect 11950 254 12008 288
rect 12042 254 12100 288
rect 12134 254 12192 288
rect 12226 254 12284 288
rect 12318 254 12376 288
rect 12410 254 12468 288
rect 12502 254 12560 288
rect 12594 254 12652 288
rect 12686 254 12744 288
rect 12778 254 12836 288
rect 12870 254 12928 288
rect 12962 254 13020 288
rect 13054 254 13112 288
rect 13146 254 13204 288
rect 13238 254 13296 288
rect 13330 254 13388 288
rect 13422 254 13480 288
rect 13514 254 13572 288
rect 13606 254 13664 288
rect 13698 254 13756 288
rect 13790 254 13848 288
rect 13882 254 13940 288
rect 13974 254 14032 288
rect 14066 254 14124 288
rect 14158 254 14216 288
rect 14250 284 14279 288
rect 14791 284 14820 288
rect 14250 254 14820 284
rect 14854 254 14912 288
rect 14946 254 15004 288
rect 15038 254 15096 288
rect 15130 254 15188 288
rect 15222 254 15280 288
rect 15314 254 15372 288
rect 15406 254 15464 288
rect 15498 254 15556 288
rect 15590 254 15648 288
rect 15682 254 15740 288
rect 15774 254 15832 288
rect 15866 254 15924 288
rect 15958 254 16016 288
rect 16050 254 16108 288
rect 16142 254 16200 288
rect 16234 254 16292 288
rect 16326 254 16384 288
rect 16418 254 16476 288
rect 16510 254 16568 288
rect 16602 254 16660 288
rect 16694 254 16752 288
rect 16786 254 16844 288
rect 16878 254 16936 288
rect 16970 254 17028 288
rect 17062 254 17120 288
rect 17154 254 17212 288
rect 17246 254 17304 288
rect 17338 254 17396 288
rect 17430 254 17488 288
rect 17522 254 17580 288
rect 17614 254 17672 288
rect 17706 254 17764 288
rect 17798 254 17856 288
rect 17890 254 17948 288
rect 17982 254 18040 288
rect 18074 254 18132 288
rect 18166 254 18224 288
rect 18258 254 18316 288
rect 18350 254 18408 288
rect 18442 254 18500 288
rect 18534 254 18592 288
rect 18626 254 18684 288
rect 18718 254 18776 288
rect 18810 254 18868 288
rect 18902 254 18960 288
rect 18994 254 19052 288
rect 19086 254 19144 288
rect 19178 254 19236 288
rect 19270 254 19328 288
rect 19362 254 19420 288
rect 19454 254 19512 288
rect 19546 254 19604 288
rect 19638 254 19696 288
rect 19730 254 19788 288
rect 19822 254 19880 288
rect 19914 254 19972 288
rect 20006 254 20064 288
rect 20098 254 20156 288
rect 20190 254 20248 288
rect 20282 254 20340 288
rect 20374 254 20432 288
rect 20466 284 20495 288
rect 20557 284 20586 288
rect 20466 254 20586 284
rect 20620 254 20678 288
rect 20712 254 20770 288
rect 20804 254 20862 288
rect 20896 254 20954 288
rect 20988 254 21046 288
rect 21080 254 21138 288
rect 21172 254 21230 288
rect 21264 254 21322 288
rect 21356 254 21414 288
rect 21448 254 21506 288
rect 21540 254 21598 288
rect 21632 254 21690 288
rect 21724 254 21782 288
rect 21816 254 21874 288
rect 21908 254 21966 288
rect 22000 254 22058 288
rect 22092 254 22150 288
rect 22184 254 22242 288
rect 22276 254 22334 288
rect 22368 254 22426 288
rect 22460 254 22518 288
rect 22552 254 22610 288
rect 22644 254 22702 288
rect 22736 254 22794 288
rect 22828 254 22886 288
rect 22920 254 22978 288
rect 23012 254 23070 288
rect 23104 254 23162 288
rect 23196 254 23254 288
rect 23288 254 23346 288
rect 23380 254 23438 288
rect 23472 254 23530 288
rect 23564 254 23622 288
rect 23656 254 23714 288
rect 23748 254 23806 288
rect 23840 254 23898 288
rect 23932 254 23990 288
rect 24024 254 24082 288
rect 24116 254 24174 288
rect 24208 254 24266 288
rect 24300 254 24358 288
rect 24392 254 24450 288
rect 24484 254 24542 288
rect 24576 254 24634 288
rect 24668 254 24726 288
rect 24760 254 24818 288
rect 24852 254 24910 288
rect 24944 254 25002 288
rect 25036 254 25094 288
rect 25128 284 25157 288
rect 25128 254 25189 284
rect 12279 239 12332 254
rect 8576 -404 8604 -400
rect 8574 -434 8604 -404
rect 8638 -434 8696 -400
rect 8730 -434 8788 -400
rect 8822 -434 8880 -400
rect 8914 -434 8972 -400
rect 9006 -434 9064 -400
rect 9098 -434 9156 -400
rect 9190 -434 9248 -400
rect 9282 -434 9340 -400
rect 9374 -434 9432 -400
rect 9466 -434 9524 -400
rect 9558 -434 9616 -400
rect 9650 -434 9708 -400
rect 9742 -434 9800 -400
rect 9834 -434 9892 -400
rect 9926 -434 9984 -400
rect 10018 -434 10076 -400
rect 10110 -434 10168 -400
rect 10202 -434 10260 -400
rect 10294 -434 10352 -400
rect 10386 -404 10410 -400
rect 10386 -434 10418 -404
rect 10604 -404 10628 -400
rect 10570 -434 10628 -404
rect 10662 -434 10720 -400
rect 10754 -434 10812 -400
rect 10846 -434 10904 -400
rect 10938 -434 10996 -400
rect 11030 -434 11088 -400
rect 11122 -434 11180 -400
rect 11214 -434 11272 -400
rect 11306 -434 11364 -400
rect 11398 -434 11456 -400
rect 11490 -434 11548 -400
rect 11582 -434 11640 -400
rect 11674 -434 11732 -400
rect 11766 -434 11824 -400
rect 11858 -434 11916 -400
rect 11950 -434 12008 -400
rect 12042 -434 12100 -400
rect 12134 -434 12192 -400
rect 12226 -434 12284 -400
rect 12318 -434 12376 -400
rect 12410 -434 12468 -400
rect 12502 -434 12560 -400
rect 12594 -434 12652 -400
rect 12686 -434 12744 -400
rect 12778 -404 12802 -400
rect 12778 -434 12829 -404
rect 12996 -404 13020 -400
rect 12962 -434 13020 -404
rect 13054 -434 13112 -400
rect 13146 -434 13204 -400
rect 13238 -434 13296 -400
rect 13330 -434 13388 -400
rect 13422 -434 13480 -400
rect 13514 -434 13572 -400
rect 13606 -434 13664 -400
rect 13698 -434 13756 -400
rect 13790 -434 13848 -400
rect 13882 -434 13940 -400
rect 13974 -434 14032 -400
rect 14066 -434 14124 -400
rect 14158 -434 14216 -400
rect 14250 -434 14308 -400
rect 14342 -434 14400 -400
rect 14434 -434 14492 -400
rect 14526 -434 14584 -400
rect 14618 -434 14676 -400
rect 14710 -434 14768 -400
rect 14802 -434 14860 -400
rect 14894 -434 14952 -400
rect 14986 -434 15044 -400
rect 15078 -434 15136 -400
rect 15170 -404 15194 -400
rect 15170 -434 15218 -404
rect 15388 -404 15412 -400
rect 15354 -434 15412 -404
rect 15446 -434 15504 -400
rect 15538 -434 15596 -400
rect 15630 -434 15688 -400
rect 15722 -434 15780 -400
rect 15814 -434 15872 -400
rect 15906 -434 15964 -400
rect 15998 -434 16056 -400
rect 16090 -434 16148 -400
rect 16182 -434 16240 -400
rect 16274 -434 16332 -400
rect 16366 -434 16424 -400
rect 16458 -434 16516 -400
rect 16550 -434 16608 -400
rect 16642 -434 16700 -400
rect 16734 -434 16792 -400
rect 16826 -434 16884 -400
rect 16918 -434 16976 -400
rect 17010 -434 17068 -400
rect 17102 -434 17160 -400
rect 17194 -434 17252 -400
rect 17286 -434 17344 -400
rect 17378 -434 17436 -400
rect 17470 -434 17528 -400
rect 17562 -404 17586 -400
rect 17562 -434 17612 -404
rect 17780 -404 17804 -400
rect 17746 -434 17804 -404
rect 17838 -434 17896 -400
rect 17930 -434 17988 -400
rect 18022 -434 18080 -400
rect 18114 -434 18172 -400
rect 18206 -434 18264 -400
rect 18298 -434 18356 -400
rect 18390 -434 18448 -400
rect 18482 -434 18540 -400
rect 18574 -434 18632 -400
rect 18666 -434 18724 -400
rect 18758 -434 18816 -400
rect 18850 -434 18908 -400
rect 18942 -434 19000 -400
rect 19034 -434 19092 -400
rect 19126 -434 19184 -400
rect 19218 -434 19276 -400
rect 19310 -434 19368 -400
rect 19402 -434 19460 -400
rect 19494 -434 19552 -400
rect 19586 -434 19644 -400
rect 19678 -434 19736 -400
rect 19770 -434 19828 -400
rect 19862 -434 19920 -400
rect 19954 -404 19978 -400
rect 19954 -434 20002 -404
rect 20172 -404 20196 -400
rect 20138 -434 20196 -404
rect 20230 -434 20288 -400
rect 20322 -434 20380 -400
rect 20414 -434 20472 -400
rect 20506 -434 20564 -400
rect 20598 -434 20656 -400
rect 20690 -434 20748 -400
rect 20782 -434 20840 -400
rect 20874 -434 20932 -400
rect 20966 -434 21024 -400
rect 21058 -434 21116 -400
rect 21150 -434 21208 -400
rect 21242 -434 21300 -400
rect 21334 -434 21392 -400
rect 21426 -434 21484 -400
rect 21518 -434 21576 -400
rect 21610 -434 21668 -400
rect 21702 -434 21760 -400
rect 21794 -434 21852 -400
rect 21886 -434 21944 -400
rect 21978 -434 22036 -400
rect 22070 -434 22128 -400
rect 22162 -434 22220 -400
rect 22254 -434 22312 -400
rect 22346 -404 22370 -400
rect 22346 -434 22394 -404
rect 22564 -404 22588 -400
rect 22530 -434 22588 -404
rect 22622 -434 22680 -400
rect 22714 -434 22772 -400
rect 22806 -434 22864 -400
rect 22898 -434 22956 -400
rect 22990 -434 23048 -400
rect 23082 -434 23140 -400
rect 23174 -434 23232 -400
rect 23266 -434 23324 -400
rect 23358 -434 23416 -400
rect 23450 -434 23508 -400
rect 23542 -434 23600 -400
rect 23634 -434 23692 -400
rect 23726 -434 23784 -400
rect 23818 -434 23876 -400
rect 23910 -434 23968 -400
rect 24002 -434 24060 -400
rect 24094 -434 24152 -400
rect 24186 -434 24244 -400
rect 24278 -434 24336 -400
rect 24370 -434 24428 -400
rect 24462 -434 24520 -400
rect 24554 -434 24612 -400
rect 24646 -434 24704 -400
rect 24738 -404 24762 -400
rect 24738 -434 24786 -404
rect 24956 -404 24980 -400
rect 24922 -434 24980 -404
rect 25014 -434 25072 -400
rect 25106 -434 25164 -400
rect 25198 -434 25256 -400
rect 25290 -434 25319 -400
rect 8575 -1089 9146 -1088
rect 8575 -1123 8604 -1089
rect 8638 -1123 8696 -1089
rect 8730 -1123 8788 -1089
rect 8822 -1123 8880 -1089
rect 8914 -1123 8969 -1089
rect 9003 -1123 9071 -1089
rect 9105 -1123 9156 -1089
rect 9190 -1123 9248 -1089
rect 9282 -1123 9340 -1089
rect 9374 -1123 9432 -1089
rect 9466 -1123 9524 -1089
rect 9558 -1123 9616 -1089
rect 9650 -1123 9708 -1089
rect 9742 -1123 9800 -1089
rect 9834 -1123 9892 -1089
rect 9926 -1123 9984 -1089
rect 10018 -1123 10076 -1089
rect 10110 -1123 10134 -1089
rect 10328 -1123 10352 -1089
rect 10386 -1123 10444 -1089
rect 10478 -1123 10536 -1089
rect 10570 -1123 10628 -1089
rect 10662 -1123 10720 -1089
rect 10754 -1123 10812 -1089
rect 10846 -1123 10904 -1089
rect 10938 -1123 10996 -1089
rect 11030 -1123 11088 -1089
rect 11122 -1123 11180 -1089
rect 11214 -1123 11272 -1089
rect 11306 -1123 11366 -1089
rect 11400 -1123 11457 -1089
rect 11491 -1123 11548 -1089
rect 11582 -1123 11640 -1089
rect 11674 -1123 11732 -1089
rect 11766 -1123 11824 -1089
rect 11858 -1123 11916 -1089
rect 11950 -1123 12008 -1089
rect 12042 -1123 12100 -1089
rect 12134 -1123 12192 -1089
rect 12226 -1123 12284 -1089
rect 12318 -1123 12376 -1089
rect 12410 -1123 12468 -1089
rect 12502 -1123 12530 -1089
rect 12720 -1123 12744 -1089
rect 12778 -1123 12836 -1089
rect 12870 -1123 12928 -1089
rect 12962 -1123 13020 -1089
rect 13054 -1123 13112 -1089
rect 13146 -1123 13204 -1089
rect 13238 -1123 13296 -1089
rect 13330 -1123 13388 -1089
rect 13422 -1123 13480 -1089
rect 13514 -1123 13572 -1089
rect 13606 -1123 13664 -1089
rect 13698 -1123 13754 -1089
rect 13788 -1123 13848 -1089
rect 13882 -1123 13940 -1089
rect 13974 -1123 14032 -1089
rect 14066 -1123 14124 -1089
rect 14158 -1123 14216 -1089
rect 14250 -1123 14308 -1089
rect 14342 -1123 14400 -1089
rect 14434 -1123 14492 -1089
rect 14526 -1123 14584 -1089
rect 14618 -1123 14676 -1089
rect 14710 -1123 14768 -1089
rect 14802 -1123 14860 -1089
rect 14894 -1123 14928 -1089
rect 15093 -1123 15136 -1089
rect 15170 -1123 15228 -1089
rect 15262 -1123 15320 -1089
rect 15354 -1123 15412 -1089
rect 15446 -1123 15504 -1089
rect 15538 -1123 15596 -1089
rect 15630 -1123 15688 -1089
rect 15722 -1123 15780 -1089
rect 15814 -1123 15872 -1089
rect 15906 -1123 15964 -1089
rect 15998 -1123 16056 -1089
rect 16090 -1123 16149 -1089
rect 16183 -1123 16240 -1089
rect 16274 -1123 16332 -1089
rect 16366 -1123 16424 -1089
rect 16458 -1123 16516 -1089
rect 16550 -1123 16608 -1089
rect 16642 -1123 16700 -1089
rect 16734 -1123 16792 -1089
rect 16826 -1123 16884 -1089
rect 16918 -1123 16976 -1089
rect 17010 -1123 17068 -1089
rect 17102 -1123 17160 -1089
rect 17194 -1123 17252 -1089
rect 17286 -1123 17320 -1089
rect 17504 -1123 17528 -1089
rect 17562 -1123 17620 -1089
rect 17654 -1123 17712 -1089
rect 17746 -1123 17804 -1089
rect 17838 -1123 17896 -1089
rect 17930 -1123 17988 -1089
rect 18022 -1123 18080 -1089
rect 18114 -1123 18172 -1089
rect 18206 -1123 18264 -1089
rect 18298 -1123 18356 -1089
rect 18390 -1123 18448 -1089
rect 18482 -1123 18538 -1089
rect 18572 -1123 18633 -1089
rect 18667 -1123 18724 -1089
rect 18758 -1123 18816 -1089
rect 18850 -1123 18908 -1089
rect 18942 -1123 19000 -1089
rect 19034 -1123 19092 -1089
rect 19126 -1123 19184 -1089
rect 19218 -1123 19276 -1089
rect 19310 -1123 19368 -1089
rect 19402 -1123 19460 -1089
rect 19494 -1123 19552 -1089
rect 19586 -1123 19644 -1089
rect 19678 -1123 19702 -1089
rect 19890 -1123 19920 -1089
rect 19954 -1123 20012 -1089
rect 20046 -1123 20104 -1089
rect 20138 -1123 20196 -1089
rect 20230 -1123 20288 -1089
rect 20322 -1123 20380 -1089
rect 20414 -1123 20472 -1089
rect 20506 -1123 20564 -1089
rect 20598 -1123 20656 -1089
rect 20690 -1123 20748 -1089
rect 20782 -1123 20840 -1089
rect 20874 -1123 20932 -1089
rect 20966 -1123 21023 -1089
rect 21057 -1123 21116 -1089
rect 21150 -1123 21208 -1089
rect 21242 -1123 21300 -1089
rect 21334 -1123 21392 -1089
rect 21426 -1123 21484 -1089
rect 21518 -1123 21576 -1089
rect 21610 -1123 21668 -1089
rect 21702 -1123 21760 -1089
rect 21794 -1123 21852 -1089
rect 21886 -1123 21944 -1089
rect 21978 -1123 22036 -1089
rect 22070 -1123 22094 -1089
rect 22214 -1123 22312 -1089
rect 22346 -1123 22404 -1089
rect 22438 -1123 22496 -1089
rect 22530 -1123 22588 -1089
rect 22622 -1123 22680 -1089
rect 22714 -1123 22772 -1089
rect 22806 -1123 22864 -1089
rect 22898 -1123 22956 -1089
rect 22990 -1123 23048 -1089
rect 23082 -1123 23140 -1089
rect 23174 -1123 23232 -1089
rect 23266 -1123 23323 -1089
rect 23357 -1123 23417 -1089
rect 23451 -1123 23508 -1089
rect 23542 -1123 23600 -1089
rect 23634 -1123 23692 -1089
rect 23726 -1123 23784 -1089
rect 23818 -1123 23876 -1089
rect 23910 -1123 23968 -1089
rect 24002 -1123 24060 -1089
rect 24094 -1123 24152 -1089
rect 24186 -1123 24244 -1089
rect 24278 -1123 24336 -1089
rect 24370 -1123 24428 -1089
rect 24462 -1123 24496 -1089
rect 24606 -1123 24704 -1089
rect 24738 -1123 24796 -1089
rect 24830 -1123 24888 -1089
rect 24922 -1123 24980 -1089
rect 25014 -1123 25072 -1089
rect 25106 -1123 25164 -1089
rect 25198 -1123 25256 -1089
rect 25290 -1123 25319 -1089
<< psubdiffcont >>
rect 10911 12466 10945 12500
rect 11003 12466 11037 12500
rect 11095 12466 11129 12500
rect 11187 12466 11221 12500
rect 11279 12466 11313 12500
rect 11371 12466 11405 12500
rect 11463 12466 11497 12500
rect 11555 12466 11589 12500
rect 11647 12466 11681 12500
rect 11739 12466 11773 12500
rect 11831 12466 11865 12500
rect 11923 12466 11957 12500
rect 12015 12466 12049 12500
rect 12107 12466 12141 12500
rect 12199 12466 12233 12500
rect 12291 12466 12325 12500
rect 12383 12466 12417 12500
rect 12475 12466 12509 12500
rect 12567 12466 12601 12500
rect 12659 12466 12693 12500
rect 12751 12466 12785 12500
rect 12843 12466 12877 12500
rect 12935 12466 12969 12500
rect 13027 12466 13061 12500
rect 13119 12466 13153 12500
rect 13211 12466 13245 12500
rect 13368 12403 13402 12437
rect 13486 12403 13520 12437
rect 13630 12403 13664 12437
rect 2480 11928 2514 11962
rect 2598 11928 2632 11962
rect 2742 11928 2776 11962
rect 20077 12403 20111 12437
rect 20195 12403 20229 12437
rect 20339 12403 20373 12437
rect 9091 11538 9125 11572
rect 9183 11538 9217 11572
rect 9277 11536 9311 11570
rect 13315 11539 13381 11596
rect 10911 11214 10945 11248
rect 11003 11214 11037 11248
rect 11095 11214 11129 11248
rect 11187 11214 11221 11248
rect 11279 11214 11313 11248
rect 11371 11214 11405 11248
rect 14099 11178 14133 11212
rect 20808 11178 20842 11212
rect 14492 11007 14526 11041
rect 14572 11007 14606 11041
rect 14652 11007 14686 11041
rect 14732 11007 14766 11041
rect 15224 11007 15258 11041
rect 15304 11007 15338 11041
rect 15384 11007 15418 11041
rect 15464 11007 15498 11041
rect 15832 11007 15866 11041
rect 15912 11007 15946 11041
rect 15992 11007 16026 11041
rect 16072 11007 16106 11041
rect 16436 11007 16470 11041
rect 16516 11007 16550 11041
rect 16596 11007 16630 11041
rect 16676 11007 16710 11041
rect 17044 11007 17078 11041
rect 17124 11007 17158 11041
rect 17204 11007 17238 11041
rect 17284 11007 17318 11041
rect 17774 11007 17808 11041
rect 17854 11007 17888 11041
rect 17934 11007 17968 11041
rect 18014 11007 18048 11041
rect 18382 11007 18416 11041
rect 18462 11007 18496 11041
rect 18542 11007 18576 11041
rect 18622 11007 18656 11041
rect 19116 11007 19150 11041
rect 19196 11007 19230 11041
rect 19276 11007 19310 11041
rect 19356 11007 19390 11041
rect 21201 11007 21235 11041
rect 21281 11007 21315 11041
rect 21361 11007 21395 11041
rect 21441 11007 21475 11041
rect 21933 11007 21967 11041
rect 22013 11007 22047 11041
rect 22093 11007 22127 11041
rect 22173 11007 22207 11041
rect 22541 11007 22575 11041
rect 22621 11007 22655 11041
rect 22701 11007 22735 11041
rect 22781 11007 22815 11041
rect 23145 11007 23179 11041
rect 23225 11007 23259 11041
rect 23305 11007 23339 11041
rect 23385 11007 23419 11041
rect 23753 11007 23787 11041
rect 23833 11007 23867 11041
rect 23913 11007 23947 11041
rect 23993 11007 24027 11041
rect 24483 11007 24517 11041
rect 24563 11007 24597 11041
rect 24643 11007 24677 11041
rect 24723 11007 24757 11041
rect 25091 11007 25125 11041
rect 25171 11007 25205 11041
rect 25251 11007 25285 11041
rect 25331 11007 25365 11041
rect 25825 11007 25859 11041
rect 25905 11007 25939 11041
rect 25985 11007 26019 11041
rect 26065 11007 26099 11041
rect 3211 10703 3245 10737
rect 3604 10532 3638 10566
rect 3684 10532 3718 10566
rect 3764 10532 3798 10566
rect 3844 10532 3878 10566
rect 4336 10532 4370 10566
rect 4416 10532 4450 10566
rect 4496 10532 4530 10566
rect 4576 10532 4610 10566
rect 4944 10532 4978 10566
rect 5024 10532 5058 10566
rect 5104 10532 5138 10566
rect 5184 10532 5218 10566
rect 5548 10532 5582 10566
rect 5628 10532 5662 10566
rect 5708 10532 5742 10566
rect 5788 10532 5822 10566
rect 6156 10532 6190 10566
rect 6236 10532 6270 10566
rect 6316 10532 6350 10566
rect 6396 10532 6430 10566
rect 6886 10532 6920 10566
rect 6966 10532 7000 10566
rect 7046 10532 7080 10566
rect 7126 10532 7160 10566
rect 7494 10532 7528 10566
rect 7574 10532 7608 10566
rect 7654 10532 7688 10566
rect 7734 10532 7768 10566
rect 8228 10532 8262 10566
rect 8308 10532 8342 10566
rect 8388 10532 8422 10566
rect 8468 10532 8502 10566
rect 3604 10080 3638 10114
rect 3684 10080 3718 10114
rect 3764 10080 3798 10114
rect 3844 10080 3878 10114
rect 4336 10080 4370 10114
rect 4416 10080 4450 10114
rect 4496 10080 4530 10114
rect 4576 10080 4610 10114
rect 4944 10080 4978 10114
rect 5024 10080 5058 10114
rect 5104 10080 5138 10114
rect 5184 10080 5218 10114
rect 5548 10080 5582 10114
rect 5628 10080 5662 10114
rect 5708 10080 5742 10114
rect 5788 10080 5822 10114
rect 6156 10080 6190 10114
rect 6236 10080 6270 10114
rect 6316 10080 6350 10114
rect 6396 10080 6430 10114
rect 6886 10080 6920 10114
rect 6966 10080 7000 10114
rect 7046 10080 7080 10114
rect 7126 10080 7160 10114
rect 7494 10080 7528 10114
rect 7574 10080 7608 10114
rect 7654 10080 7688 10114
rect 7734 10080 7768 10114
rect 8228 10080 8262 10114
rect 8308 10080 8342 10114
rect 8388 10080 8422 10114
rect 8468 10080 8502 10114
rect 13789 10068 13823 10102
rect 13869 10068 13903 10102
rect 13949 10068 13983 10102
rect 14029 10068 14063 10102
rect 14523 10068 14557 10102
rect 14603 10068 14637 10102
rect 14683 10068 14717 10102
rect 14763 10068 14797 10102
rect 15131 10068 15165 10102
rect 15211 10068 15245 10102
rect 15291 10068 15325 10102
rect 15371 10068 15405 10102
rect 15861 10068 15895 10102
rect 15941 10068 15975 10102
rect 16021 10068 16055 10102
rect 16101 10068 16135 10102
rect 16469 10068 16503 10102
rect 16549 10068 16583 10102
rect 16629 10068 16663 10102
rect 16709 10068 16743 10102
rect 17073 10068 17107 10102
rect 17153 10068 17187 10102
rect 17233 10068 17267 10102
rect 17313 10068 17347 10102
rect 17681 10068 17715 10102
rect 17761 10068 17795 10102
rect 17841 10068 17875 10102
rect 17921 10068 17955 10102
rect 18413 10068 18447 10102
rect 18493 10068 18527 10102
rect 18573 10068 18607 10102
rect 18653 10068 18687 10102
rect 20498 10068 20532 10102
rect 20578 10068 20612 10102
rect 20658 10068 20692 10102
rect 20738 10068 20772 10102
rect 21232 10068 21266 10102
rect 21312 10068 21346 10102
rect 21392 10068 21426 10102
rect 21472 10068 21506 10102
rect 21840 10068 21874 10102
rect 21920 10068 21954 10102
rect 22000 10068 22034 10102
rect 22080 10068 22114 10102
rect 22570 10068 22604 10102
rect 22650 10068 22684 10102
rect 22730 10068 22764 10102
rect 22810 10068 22844 10102
rect 23178 10068 23212 10102
rect 23258 10068 23292 10102
rect 23338 10068 23372 10102
rect 23418 10068 23452 10102
rect 23782 10068 23816 10102
rect 23862 10068 23896 10102
rect 23942 10068 23976 10102
rect 24022 10068 24056 10102
rect 24390 10068 24424 10102
rect 24470 10068 24504 10102
rect 24550 10068 24584 10102
rect 24630 10068 24664 10102
rect 25122 10068 25156 10102
rect 25202 10068 25236 10102
rect 25282 10068 25316 10102
rect 25362 10068 25396 10102
rect 3211 9909 3245 9943
rect 19046 9897 19080 9931
rect 25755 9897 25789 9931
rect 9090 9068 9124 9102
rect 9182 9068 9216 9102
rect 9274 9068 9308 9102
rect 9346 9068 9380 9102
rect 9438 9067 9472 9101
rect 9530 9068 9564 9102
rect 9714 9068 9748 9102
rect 9806 9068 9840 9102
rect 9898 9069 9932 9103
rect 9990 9068 10024 9102
rect 10082 9067 10116 9101
rect 10174 9068 10208 9102
rect 10266 9068 10300 9102
rect 10358 9068 10392 9102
rect 10450 9068 10484 9102
rect 10542 9068 10576 9102
rect 10634 9068 10668 9102
rect 10726 9068 10760 9102
rect 10818 9068 10852 9102
rect 10910 9067 10944 9101
rect 11002 9068 11036 9102
rect 11094 9068 11128 9102
rect 11278 9068 11312 9102
rect 11370 9068 11404 9102
rect 11462 9068 11496 9102
rect 11554 9068 11588 9102
rect 11646 9067 11680 9101
rect 2480 8684 2514 8718
rect 2598 8684 2632 8718
rect 2742 8684 2776 8718
rect 19515 8672 19549 8706
rect 19659 8672 19693 8706
rect 19777 8672 19811 8706
rect 26224 8672 26258 8706
rect 26368 8672 26402 8706
rect 26486 8672 26520 8706
rect 10083 7737 10117 7771
rect 10175 7737 10209 7771
rect 10267 7737 10301 7771
rect 10359 7737 10393 7771
rect 10451 7737 10485 7771
rect 10727 7737 10761 7771
rect 10819 7736 10853 7770
rect 10910 7737 10944 7771
rect 11002 7737 11036 7771
rect 11095 7737 11129 7771
rect 11186 7737 11220 7771
rect 11278 7737 11312 7771
rect 11554 7736 11588 7770
rect 11646 7736 11680 7770
rect 11527 6492 11561 6526
rect 11619 6492 11653 6526
rect 11711 6492 11745 6526
rect 11803 6492 11837 6526
rect 11895 6492 11929 6526
rect 11987 6492 12021 6526
rect 12079 6492 12113 6526
rect 12171 6492 12205 6526
rect 12263 6492 12297 6526
rect 12355 6492 12389 6526
rect 12447 6492 12481 6526
rect 12539 6492 12573 6526
rect 12631 6492 12665 6526
rect 12723 6492 12757 6526
rect 12815 6492 12849 6526
rect 12907 6492 12941 6526
rect 12999 6492 13033 6526
rect 13091 6492 13125 6526
rect 13183 6492 13217 6526
rect 13275 6492 13309 6526
rect 13367 6492 13401 6526
rect 13459 6492 13493 6526
rect 13551 6492 13585 6526
rect 13643 6492 13677 6526
rect 13735 6492 13769 6526
rect 13827 6492 13861 6526
rect 13919 6492 13953 6526
rect 14011 6492 14045 6526
rect 14103 6492 14137 6526
rect 14195 6492 14229 6526
rect 14287 6492 14321 6526
rect 14379 6492 14413 6526
rect 14471 6492 14505 6526
rect 24093 6106 24127 6140
rect 24211 6106 24245 6140
rect 24355 6106 24389 6140
rect 30708 5723 30742 5757
rect 30800 5724 30834 5758
rect 30892 5724 30926 5758
rect 30985 5724 31019 5758
rect 11526 5619 11560 5653
rect 11618 5619 11652 5653
rect 11710 5619 11744 5653
rect 11802 5619 11836 5653
rect 11894 5619 11928 5653
rect 11986 5619 12020 5653
rect 12078 5619 12112 5653
rect 12170 5619 12204 5653
rect 12262 5619 12296 5653
rect 12354 5619 12388 5653
rect 12446 5619 12480 5653
rect 12538 5619 12572 5653
rect 12630 5619 12664 5653
rect 12722 5619 12756 5653
rect 12814 5619 12848 5653
rect 12906 5619 12940 5653
rect 12998 5619 13032 5653
rect 13090 5619 13124 5653
rect 13182 5619 13216 5653
rect 13274 5619 13308 5653
rect 13366 5619 13400 5653
rect 13458 5619 13492 5653
rect 13550 5619 13584 5653
rect 13642 5619 13676 5653
rect 13734 5619 13768 5653
rect 13826 5619 13860 5653
rect 13918 5619 13952 5653
rect 14010 5619 14044 5653
rect 14102 5619 14136 5653
rect 14194 5619 14228 5653
rect 14286 5619 14320 5653
rect 14378 5619 14412 5653
rect 14470 5619 14504 5653
rect 14562 5619 14596 5653
rect 14654 5619 14688 5653
rect 14746 5619 14780 5653
rect 14838 5619 14872 5653
rect 14930 5619 14964 5653
rect 15022 5619 15056 5653
rect 15114 5619 15148 5653
rect 15206 5619 15240 5653
rect 15298 5619 15332 5653
rect 15390 5619 15424 5653
rect 15482 5619 15516 5653
rect 15574 5619 15608 5653
rect 15666 5619 15700 5653
rect 15758 5619 15792 5653
rect 15850 5619 15884 5653
rect 15942 5619 15976 5653
rect 16034 5619 16068 5653
rect 16126 5619 16160 5653
rect 16218 5619 16252 5653
rect 16310 5619 16344 5653
rect 16402 5619 16436 5653
rect 16494 5619 16528 5653
rect 16586 5619 16620 5653
rect 16678 5619 16712 5653
rect 16770 5619 16804 5653
rect 16862 5619 16896 5653
rect 16954 5619 16988 5653
rect 17046 5619 17080 5653
rect 17138 5619 17172 5653
rect 17230 5619 17264 5653
rect 17322 5619 17356 5653
rect 17414 5619 17448 5653
rect 17506 5619 17540 5653
rect 17598 5619 17632 5653
rect 17690 5619 17724 5653
rect 17782 5619 17816 5653
rect 17874 5619 17908 5653
rect 17966 5619 18000 5653
rect 18058 5619 18092 5653
rect 18150 5619 18184 5653
rect 18242 5619 18276 5653
rect 18334 5619 18368 5653
rect 18426 5619 18460 5653
rect 18518 5619 18552 5653
rect 18610 5619 18644 5653
rect 18702 5619 18736 5653
rect 18794 5619 18828 5653
rect 18886 5619 18920 5653
rect 18978 5619 19012 5653
rect 19070 5619 19104 5653
rect 19162 5619 19196 5653
rect 19254 5619 19288 5653
rect 19346 5619 19380 5653
rect 19438 5619 19472 5653
rect 19530 5619 19564 5653
rect 19622 5619 19656 5653
rect 19714 5619 19748 5653
rect 19806 5619 19840 5653
rect 19898 5619 19932 5653
rect 19990 5619 20024 5653
rect 20082 5619 20116 5653
rect 20174 5619 20208 5653
rect 20266 5619 20300 5653
rect 20358 5619 20392 5653
rect 20450 5619 20484 5653
rect 20542 5619 20576 5653
rect 20634 5619 20668 5653
rect 20726 5619 20760 5653
rect 20818 5619 20852 5653
rect 20910 5619 20944 5653
rect 21002 5619 21036 5653
rect 21094 5619 21128 5653
rect 21186 5619 21220 5653
rect 21278 5619 21312 5653
rect 21370 5619 21404 5653
rect 21462 5619 21496 5653
rect 21554 5619 21588 5653
rect 21646 5619 21680 5653
rect 21738 5619 21772 5653
rect 21830 5619 21864 5653
rect 21922 5619 21956 5653
rect 22014 5619 22048 5653
rect 22106 5619 22140 5653
rect 22198 5619 22232 5653
rect 22290 5619 22324 5653
rect 22382 5619 22416 5653
rect 22474 5619 22508 5653
rect 22566 5619 22600 5653
rect 22658 5619 22692 5653
rect 22750 5619 22784 5653
rect 22842 5619 22876 5653
rect 22934 5619 22968 5653
rect 23026 5619 23060 5653
rect 23118 5619 23152 5653
rect 23210 5619 23244 5653
rect 23302 5619 23336 5653
rect 23394 5619 23428 5653
rect 11086 4930 11120 4964
rect 11178 4930 11212 4964
rect 11270 4930 11304 4964
rect 11362 4930 11396 4964
rect 11454 4930 11488 4964
rect 11546 4930 11580 4964
rect 11638 4930 11672 4964
rect 11730 4930 11764 4964
rect 11822 4930 11856 4964
rect 11914 4930 11948 4964
rect 12006 4930 12040 4964
rect 12098 4930 12132 4964
rect 12190 4930 12224 4964
rect 12282 4930 12316 4964
rect 12374 4930 12408 4964
rect 12466 4930 12500 4964
rect 12558 4930 12592 4964
rect 12650 4930 12684 4964
rect 12742 4930 12776 4964
rect 12834 4930 12868 4964
rect 12926 4930 12960 4964
rect 13018 4930 13052 4964
rect 13110 4930 13144 4964
rect 13202 4930 13236 4964
rect 13294 4930 13328 4964
rect 13386 4930 13420 4964
rect 13478 4930 13512 4964
rect 13570 4930 13604 4964
rect 13662 4930 13696 4964
rect 13754 4930 13788 4964
rect 13846 4930 13880 4964
rect 13938 4930 13972 4964
rect 14030 4930 14064 4964
rect 14122 4930 14156 4964
rect 14214 4930 14248 4964
rect 14306 4930 14340 4964
rect 14398 4930 14432 4964
rect 14490 4930 14524 4964
rect 14582 4930 14616 4964
rect 14674 4930 14708 4964
rect 14766 4930 14800 4964
rect 14858 4930 14892 4964
rect 14950 4930 14984 4964
rect 15042 4930 15076 4964
rect 15134 4930 15168 4964
rect 15226 4930 15260 4964
rect 15318 4930 15352 4964
rect 15410 4930 15444 4964
rect 15502 4930 15536 4964
rect 15594 4930 15628 4964
rect 15686 4930 15720 4964
rect 15778 4930 15812 4964
rect 15870 4930 15904 4964
rect 15962 4930 15996 4964
rect 16054 4930 16088 4964
rect 16146 4930 16180 4964
rect 16238 4930 16272 4964
rect 16330 4930 16364 4964
rect 16422 4930 16456 4964
rect 16514 4930 16548 4964
rect 16606 4930 16640 4964
rect 16698 4930 16732 4964
rect 16790 4930 16824 4964
rect 16882 4930 16916 4964
rect 16974 4930 17008 4964
rect 17066 4930 17100 4964
rect 17158 4930 17192 4964
rect 17250 4930 17284 4964
rect 17342 4930 17376 4964
rect 17434 4930 17468 4964
rect 17526 4930 17560 4964
rect 17618 4930 17652 4964
rect 17710 4930 17744 4964
rect 17802 4930 17836 4964
rect 17894 4930 17928 4964
rect 17986 4930 18020 4964
rect 18078 4930 18112 4964
rect 18170 4930 18204 4964
rect 18262 4930 18296 4964
rect 18354 4930 18388 4964
rect 18446 4930 18480 4964
rect 18538 4930 18572 4964
rect 18630 4930 18664 4964
rect 18722 4930 18756 4964
rect 18814 4930 18848 4964
rect 18906 4930 18940 4964
rect 18998 4930 19032 4964
rect 19090 4930 19124 4964
rect 19182 4930 19216 4964
rect 19274 4930 19308 4964
rect 19366 4930 19400 4964
rect 19458 4930 19492 4964
rect 19550 4930 19584 4964
rect 19642 4930 19676 4964
rect 19734 4930 19768 4964
rect 19826 4930 19860 4964
rect 19898 4930 19932 4964
rect 19990 4930 20024 4964
rect 20082 4930 20116 4964
rect 20174 4930 20208 4964
rect 20266 4930 20300 4964
rect 20358 4930 20392 4964
rect 20450 4930 20484 4964
rect 20542 4930 20576 4964
rect 20634 4930 20668 4964
rect 20726 4930 20760 4964
rect 20818 4930 20852 4964
rect 20910 4930 20944 4964
rect 21002 4930 21036 4964
rect 21094 4930 21128 4964
rect 21186 4930 21220 4964
rect 21278 4930 21312 4964
rect 21370 4930 21404 4964
rect 21462 4930 21496 4964
rect 21554 4930 21588 4964
rect 21646 4930 21680 4964
rect 21738 4930 21772 4964
rect 21830 4930 21864 4964
rect 21922 4930 21956 4964
rect 22014 4930 22048 4964
rect 22106 4930 22140 4964
rect 22198 4930 22232 4964
rect 22290 4930 22324 4964
rect 22382 4930 22416 4964
rect 22474 4930 22508 4964
rect 22566 4930 22600 4964
rect 22658 4930 22692 4964
rect 22750 4930 22784 4964
rect 22842 4930 22876 4964
rect 22934 4930 22968 4964
rect 23026 4930 23060 4964
rect 23118 4930 23152 4964
rect 23210 4930 23244 4964
rect 23302 4930 23336 4964
rect 23394 4930 23428 4964
rect 24824 4881 24858 4915
rect 25217 4710 25251 4744
rect 25297 4710 25331 4744
rect 25377 4710 25411 4744
rect 25457 4710 25491 4744
rect 25949 4710 25983 4744
rect 26029 4710 26063 4744
rect 26109 4710 26143 4744
rect 26189 4710 26223 4744
rect 26557 4710 26591 4744
rect 26637 4710 26671 4744
rect 26717 4710 26751 4744
rect 26797 4710 26831 4744
rect 27161 4710 27195 4744
rect 27241 4710 27275 4744
rect 27321 4710 27355 4744
rect 27401 4710 27435 4744
rect 27769 4710 27803 4744
rect 27849 4710 27883 4744
rect 27929 4710 27963 4744
rect 28009 4710 28043 4744
rect 28499 4710 28533 4744
rect 28579 4710 28613 4744
rect 28659 4710 28693 4744
rect 28739 4710 28773 4744
rect 29107 4710 29141 4744
rect 29187 4710 29221 4744
rect 29267 4710 29301 4744
rect 29347 4710 29381 4744
rect 29841 4710 29875 4744
rect 29921 4710 29955 4744
rect 30001 4710 30035 4744
rect 30081 4710 30115 4744
rect 25606 4298 25640 4332
rect 25698 4298 25732 4332
rect 25790 4298 25824 4332
rect 25882 4298 25916 4332
rect 25974 4298 26008 4332
rect 26066 4298 26100 4332
rect 26158 4298 26192 4332
rect 26250 4298 26284 4332
rect 26342 4298 26376 4332
rect 26433 4298 26467 4332
rect 26526 4298 26560 4332
rect 26618 4298 26652 4332
rect 26710 4298 26744 4332
rect 26802 4298 26836 4332
rect 26894 4298 26928 4332
rect 26986 4298 27020 4332
rect 27078 4298 27112 4332
rect 27170 4298 27204 4332
rect 27262 4298 27296 4332
rect 27354 4298 27388 4332
rect 27446 4298 27480 4332
rect 27538 4298 27572 4332
rect 27630 4298 27664 4332
rect 27722 4298 27756 4332
rect 27814 4298 27848 4332
rect 27906 4298 27940 4332
rect 27998 4298 28032 4332
rect 28090 4298 28124 4332
rect 28182 4298 28216 4332
rect 28274 4298 28308 4332
rect 28366 4298 28400 4332
rect 28458 4298 28492 4332
rect 28550 4298 28584 4332
rect 28642 4298 28676 4332
rect 28734 4298 28768 4332
rect 28826 4298 28860 4332
rect 28918 4298 28952 4332
rect 29010 4298 29044 4332
rect 29102 4298 29136 4332
rect 29194 4298 29228 4332
rect 29286 4298 29320 4332
rect 29378 4298 29412 4332
rect 29470 4298 29504 4332
rect 29562 4298 29596 4332
rect 29654 4298 29688 4332
rect 29746 4298 29780 4332
rect 29838 4298 29872 4332
rect 29930 4298 29964 4332
rect 30022 4298 30056 4332
rect 30114 4298 30148 4332
rect 30206 4298 30240 4332
rect 30298 4298 30332 4332
rect 11117 4045 11151 4079
rect 11210 4045 11244 4079
rect 11302 4045 11336 4079
rect 11394 4045 11428 4079
rect 11486 4045 11520 4079
rect 11578 4045 11612 4079
rect 11670 4045 11704 4079
rect 11762 4045 11796 4079
rect 11854 4045 11888 4079
rect 13660 4057 13694 4091
rect 13752 4057 13786 4091
rect 13844 4057 13878 4091
rect 13936 4057 13970 4091
rect 14028 4057 14062 4091
rect 14120 4057 14154 4091
rect 14212 4057 14246 4091
rect 14304 4057 14338 4091
rect 14396 4057 14430 4091
rect 14488 4057 14522 4091
rect 14580 4057 14614 4091
rect 14672 4057 14706 4091
rect 14764 4057 14798 4091
rect 14856 4057 14890 4091
rect 14948 4057 14982 4091
rect 15040 4057 15074 4091
rect 15132 4057 15166 4091
rect 15224 4057 15258 4091
rect 15316 4057 15350 4091
rect 15408 4057 15442 4091
rect 15500 4057 15534 4091
rect 15592 4057 15626 4091
rect 15684 4057 15718 4091
rect 15776 4057 15810 4091
rect 15868 4057 15902 4091
rect 15960 4057 15994 4091
rect 16052 4057 16086 4091
rect 16144 4057 16178 4091
rect 16236 4057 16270 4091
rect 16328 4057 16362 4091
rect 16420 4057 16454 4091
rect 16512 4057 16546 4091
rect 16604 4057 16638 4091
rect 16696 4057 16730 4091
rect 16788 4057 16822 4091
rect 16880 4057 16914 4091
rect 16972 4057 17006 4091
rect 17064 4057 17098 4091
rect 17156 4057 17190 4091
rect 17248 4057 17282 4091
rect 17340 4057 17374 4091
rect 17432 4057 17466 4091
rect 17524 4057 17558 4091
rect 17616 4057 17650 4091
rect 17708 4057 17742 4091
rect 17800 4057 17834 4091
rect 17892 4057 17926 4091
rect 17984 4057 18018 4091
rect 18076 4057 18110 4091
rect 18168 4057 18202 4091
rect 18260 4057 18294 4091
rect 18352 4057 18386 4091
rect 18444 4057 18478 4091
rect 18536 4057 18570 4091
rect 18628 4057 18662 4091
rect 18720 4057 18754 4091
rect 18812 4057 18846 4091
rect 18904 4057 18938 4091
rect 18996 4057 19030 4091
rect 19088 4057 19122 4091
rect 19180 4057 19214 4091
rect 19272 4057 19306 4091
rect 19364 4057 19398 4091
rect 19456 4057 19490 4091
rect 19548 4057 19582 4091
rect 19640 4057 19674 4091
rect 19732 4057 19766 4091
rect 19824 4057 19858 4091
rect 19916 4057 19950 4091
rect 20008 4057 20042 4091
rect 20100 4057 20134 4091
rect 20192 4057 20226 4091
rect 20284 4057 20318 4091
rect 20357 4057 20410 4091
rect 20449 4057 20502 4091
rect 20541 4057 20594 4091
rect 20633 4057 20686 4091
rect 20725 4057 20778 4091
rect 20817 4057 20870 4091
rect 20909 4057 20962 4091
rect 21001 4057 21054 4091
rect 21093 4057 21146 4091
rect 21185 4057 21238 4091
rect 21277 4057 21330 4091
rect 21369 4057 21422 4091
rect 21461 4057 21514 4091
rect 21553 4057 21606 4091
rect 21645 4057 21698 4091
rect 21737 4057 21790 4091
rect 21829 4057 21882 4091
rect 21921 4057 21974 4091
rect 22013 4057 22066 4091
rect 22105 4057 22158 4091
rect 22197 4057 22250 4091
rect 22289 4057 22342 4091
rect 22381 4057 22434 4091
rect 22473 4057 22507 4091
rect 22565 4057 22599 4091
rect 22657 4057 22691 4091
rect 22749 4057 22783 4091
rect 22841 4057 22875 4091
rect 22933 4057 22967 4091
rect 23025 4057 23059 4091
rect 23117 4057 23151 4091
rect 23209 4057 23243 4091
rect 23301 4057 23335 4091
rect 23393 4057 23427 4091
rect 11525 3184 11559 3218
rect 11617 3184 11651 3218
rect 11709 3184 11743 3218
rect 11801 3184 11835 3218
rect 11893 3184 11927 3218
rect 11985 3184 12019 3218
rect 12077 3184 12111 3218
rect 12169 3184 12203 3218
rect 12261 3184 12295 3218
rect 12353 3184 12387 3218
rect 12445 3184 12479 3218
rect 12537 3184 12571 3218
rect 12629 3184 12663 3218
rect 12721 3184 12755 3218
rect 12813 3184 12847 3218
rect 12905 3184 12939 3218
rect 12997 3184 13031 3218
rect 13089 3184 13123 3218
rect 13181 3184 13215 3218
rect 13273 3184 13307 3218
rect 13365 3184 13399 3218
rect 13457 3184 13491 3218
rect 13549 3184 13583 3218
rect 13641 3184 13675 3218
rect 13733 3184 13767 3218
rect 13825 3184 13859 3218
rect 13917 3184 13951 3218
rect 14009 3184 14043 3218
rect 14101 3184 14135 3218
rect 14193 3184 14227 3218
rect 14285 3184 14319 3218
rect 14377 3184 14411 3218
rect 14469 3184 14503 3218
rect 14561 3184 14595 3218
rect 14653 3184 14687 3218
rect 14745 3184 14779 3218
rect 14837 3184 14871 3218
rect 14929 3184 14963 3218
rect 15021 3184 15055 3218
rect 15113 3184 15147 3218
rect 15205 3184 15239 3218
rect 15297 3184 15331 3218
rect 15389 3184 15423 3218
rect 15481 3184 15515 3218
rect 15573 3184 15607 3218
rect 15665 3184 15699 3218
rect 15757 3184 15791 3218
rect 15849 3184 15883 3218
rect 15941 3184 15975 3218
rect 16033 3184 16067 3218
rect 16125 3184 16159 3218
rect 16217 3184 16251 3218
rect 16309 3184 16343 3218
rect 16401 3184 16435 3218
rect 16493 3184 16527 3218
rect 16585 3184 16619 3218
rect 16677 3184 16711 3218
rect 16769 3184 16803 3218
rect 16861 3184 16895 3218
rect 16953 3184 16987 3218
rect 17045 3184 17079 3218
rect 17137 3184 17171 3218
rect 17229 3184 17263 3218
rect 17321 3184 17355 3218
rect 17413 3184 17447 3218
rect 17505 3184 17539 3218
rect 17597 3184 17631 3218
rect 17689 3184 17723 3218
rect 17781 3184 17815 3218
rect 17873 3184 17907 3218
rect 17965 3184 17999 3218
rect 18057 3184 18091 3218
rect 18149 3184 18183 3218
rect 18241 3184 18275 3218
rect 18333 3184 18367 3218
rect 18425 3184 18459 3218
rect 18517 3184 18551 3218
rect 18609 3184 18643 3218
rect 18701 3184 18735 3218
rect 18793 3184 18827 3218
rect 18885 3184 18919 3218
rect 18977 3184 19011 3218
rect 19069 3184 19103 3218
rect 19161 3184 19195 3218
rect 19253 3184 19287 3218
rect 19345 3184 19379 3218
rect 19437 3184 19471 3218
rect 19529 3184 19563 3218
rect 19621 3184 19655 3218
rect 19713 3184 19747 3218
rect 19805 3184 19839 3218
rect 19897 3184 19931 3218
rect 19989 3184 20023 3218
rect 20081 3184 20115 3218
rect 20173 3184 20207 3218
rect 20265 3184 20299 3218
rect 20357 3184 20391 3218
rect 20449 3184 20483 3218
rect 20541 3184 20575 3218
rect 20633 3184 20667 3218
rect 20725 3184 20759 3218
rect 20817 3184 20851 3218
rect 20909 3184 20943 3218
rect 21001 3184 21035 3218
rect 21093 3184 21127 3218
rect 21185 3184 21219 3218
rect 21277 3184 21311 3218
rect 21369 3184 21403 3218
rect 21461 3184 21495 3218
rect 21553 3184 21587 3218
rect 21645 3184 21679 3218
rect 21737 3184 21771 3218
rect 21829 3184 21863 3218
rect 21921 3184 21955 3218
rect 22013 3184 22047 3218
rect 22105 3184 22139 3218
rect 22197 3184 22231 3218
rect 22289 3184 22323 3218
rect 22381 3184 22415 3218
rect 22473 3184 22507 3218
rect 22565 3184 22599 3218
rect 22657 3184 22691 3218
rect 22749 3184 22783 3218
rect 22841 3184 22875 3218
rect 22933 3184 22967 3218
rect 23025 3184 23059 3218
rect 23117 3184 23151 3218
rect 23209 3184 23243 3218
rect 23301 3184 23335 3218
rect 23393 3184 23427 3218
rect 25606 3033 25640 3067
rect 25698 3033 25732 3067
rect 25790 3033 25824 3067
rect 25882 3033 25916 3067
rect 25974 3033 26008 3067
rect 26066 3033 26100 3067
rect 26158 3033 26192 3067
rect 26250 3033 26284 3067
rect 26342 3033 26376 3067
rect 26434 3033 26468 3067
rect 26526 3033 26560 3067
rect 26618 3033 26652 3067
rect 26710 3033 26744 3067
rect 26802 3033 26836 3067
rect 26894 3033 26928 3067
rect 26986 3033 27020 3067
rect 27078 3033 27112 3067
rect 27171 3033 27205 3067
rect 27262 3033 27296 3067
rect 27354 3033 27388 3067
rect 27446 3033 27480 3067
rect 27539 3033 27573 3067
rect 27630 3033 27664 3067
rect 27722 3033 27756 3067
rect 27814 3033 27848 3067
rect 27906 3033 27940 3067
rect 27998 3033 28032 3067
rect 28090 3033 28124 3067
rect 28182 3033 28216 3067
rect 28274 3033 28308 3067
rect 28366 3033 28400 3067
rect 28458 3033 28492 3067
rect 28550 3033 28584 3067
rect 28642 3033 28676 3067
rect 28733 3033 28767 3067
rect 28825 3033 28859 3067
rect 28918 3033 28952 3067
rect 29010 3033 29044 3067
rect 29102 3033 29136 3067
rect 29193 3033 29227 3067
rect 29286 3033 29320 3067
rect 29377 3033 29411 3067
rect 29470 3033 29504 3067
rect 29562 3033 29596 3067
rect 29654 3033 29688 3067
rect 29746 3033 29780 3067
rect 29838 3033 29872 3067
rect 29930 3033 29964 3067
rect 30022 3033 30056 3067
rect 30114 3033 30148 3067
rect 30206 3033 30240 3067
rect 30298 3033 30332 3067
rect 25606 1766 25640 1800
rect 25698 1766 25732 1800
rect 25790 1766 25824 1800
rect 25882 1766 25916 1800
rect 25974 1766 26008 1800
rect 26066 1766 26100 1800
rect 26158 1766 26192 1800
rect 26250 1766 26284 1800
rect 26342 1766 26376 1800
rect 26434 1766 26468 1800
rect 26526 1766 26560 1800
rect 26618 1766 26652 1800
rect 26710 1766 26744 1800
rect 26802 1766 26836 1800
rect 26894 1766 26928 1800
rect 26986 1766 27020 1800
rect 27078 1766 27112 1800
rect 27170 1766 27204 1800
rect 27262 1766 27296 1800
rect 27354 1766 27388 1800
rect 27446 1766 27480 1800
rect 27538 1766 27572 1800
rect 27630 1766 27664 1800
rect 27722 1766 27756 1800
rect 27814 1766 27848 1800
rect 27906 1766 27940 1800
rect 27998 1766 28032 1800
rect 28090 1766 28124 1800
rect 28182 1766 28216 1800
rect 28274 1766 28308 1800
rect 28366 1766 28400 1800
rect 28458 1766 28492 1800
rect 28550 1766 28584 1800
rect 28642 1766 28676 1800
rect 28734 1766 28768 1800
rect 28826 1766 28860 1800
rect 28918 1766 28952 1800
rect 29010 1766 29044 1800
rect 29102 1766 29136 1800
rect 29194 1766 29228 1800
rect 29286 1766 29320 1800
rect 29378 1766 29412 1800
rect 29470 1766 29504 1800
rect 29562 1766 29596 1800
rect 29654 1766 29688 1800
rect 29746 1766 29780 1800
rect 29838 1766 29872 1800
rect 29930 1766 29964 1800
rect 30022 1766 30056 1800
rect 30114 1766 30148 1800
rect 30206 1766 30240 1800
rect 30298 1766 30332 1800
rect 8606 804 8640 838
rect 8698 804 8732 838
rect 8790 804 8824 838
rect 8882 804 8916 838
rect 8974 804 9008 838
rect 9066 804 9100 838
rect 9158 804 9192 838
rect 9250 804 9284 838
rect 9342 804 9376 838
rect 9434 804 9468 838
rect 9526 804 9560 838
rect 9618 804 9652 838
rect 9710 804 9744 838
rect 9802 804 9836 838
rect 9894 804 9928 838
rect 9986 804 10020 838
rect 10078 804 10112 838
rect 10170 804 10204 838
rect 10262 804 10296 838
rect 10354 804 10388 838
rect 10446 804 10480 838
rect 10538 804 10572 838
rect 10630 804 10664 838
rect 10722 804 10756 838
rect 10814 804 10848 838
rect 10906 804 10940 838
rect 10998 804 11032 838
rect 11090 804 11124 838
rect 11182 804 11216 838
rect 11274 804 11308 838
rect 11366 804 11400 838
rect 12990 804 13024 838
rect 13082 804 13116 838
rect 13174 804 13208 838
rect 13266 804 13300 838
rect 13358 804 13392 838
rect 13450 804 13484 838
rect 13542 804 13576 838
rect 13634 804 13668 838
rect 13726 804 13760 838
rect 13818 804 13852 838
rect 13910 804 13944 838
rect 14002 804 14036 838
rect 14094 804 14128 838
rect 14186 804 14220 838
rect 14278 804 14312 838
rect 14370 804 14404 838
rect 14462 804 14496 838
rect 14554 804 14588 838
rect 14646 804 14680 838
rect 14738 804 14772 838
rect 14830 804 14864 838
rect 14922 804 14956 838
rect 15014 804 15048 838
rect 15106 804 15140 838
rect 15198 804 15232 838
rect 15290 804 15324 838
rect 15382 804 15416 838
rect 15474 804 15508 838
rect 15566 804 15600 838
rect 15658 804 15692 838
rect 15750 804 15784 838
rect 8604 -338 8638 -304
rect 8696 -338 8730 -304
rect 8788 -338 8822 -304
rect 8880 -338 8914 -304
rect 8972 -338 9006 -304
rect 9064 -338 9098 -304
rect 9156 -338 9190 -304
rect 9248 -338 9282 -304
rect 9340 -338 9374 -304
rect 9432 -338 9466 -304
rect 9524 -338 9558 -304
rect 9616 -338 9650 -304
rect 9708 -338 9742 -304
rect 9800 -338 9834 -304
rect 9892 -338 9926 -304
rect 9984 -338 10018 -304
rect 10076 -338 10110 -304
rect 10168 -338 10202 -304
rect 10260 -338 10294 -304
rect 10352 -338 10386 -304
rect 10444 -338 10478 -304
rect 10536 -338 10570 -304
rect 10628 -338 10662 -304
rect 10720 -338 10754 -304
rect 10812 -338 10846 -304
rect 10904 -338 10938 -304
rect 10996 -338 11030 -304
rect 11088 -338 11122 -304
rect 11180 -338 11214 -304
rect 11272 -338 11306 -304
rect 11364 -338 11398 -304
rect 11456 -338 11490 -304
rect 11548 -338 11582 -304
rect 11640 -338 11674 -304
rect 11732 -338 11766 -304
rect 11824 -338 11858 -304
rect 11916 -338 11950 -304
rect 12008 -338 12042 -304
rect 12100 -338 12134 -304
rect 12192 -338 12226 -304
rect 12284 -338 12318 -304
rect 12376 -338 12410 -304
rect 12468 -338 12502 -304
rect 12560 -338 12594 -304
rect 12652 -338 12686 -304
rect 12744 -338 12778 -304
rect 12836 -338 12870 -304
rect 12928 -338 12962 -304
rect 13020 -338 13054 -304
rect 13112 -338 13146 -304
rect 13204 -338 13238 -304
rect 13296 -338 13330 -304
rect 13388 -338 13422 -304
rect 13480 -338 13514 -304
rect 13572 -338 13606 -304
rect 13664 -338 13698 -304
rect 13756 -338 13790 -304
rect 13848 -338 13882 -304
rect 13940 -338 13974 -304
rect 14032 -338 14066 -304
rect 14124 -338 14158 -304
rect 14216 -338 14250 -304
rect 14820 -338 14854 -304
rect 14912 -338 14946 -304
rect 15004 -338 15038 -304
rect 15096 -338 15130 -304
rect 15188 -338 15222 -304
rect 15280 -338 15314 -304
rect 15372 -338 15406 -304
rect 15464 -338 15498 -304
rect 15556 -338 15590 -304
rect 15648 -338 15682 -304
rect 15740 -338 15774 -304
rect 15832 -338 15866 -304
rect 15924 -338 15958 -304
rect 16016 -338 16050 -304
rect 16108 -338 16142 -304
rect 16200 -338 16234 -304
rect 16292 -338 16326 -304
rect 16384 -338 16418 -304
rect 16476 -338 16510 -304
rect 16568 -338 16602 -304
rect 16660 -338 16694 -304
rect 16752 -338 16786 -304
rect 16844 -338 16878 -304
rect 16936 -338 16970 -304
rect 17028 -338 17062 -304
rect 17120 -338 17154 -304
rect 17212 -338 17246 -304
rect 17304 -338 17338 -304
rect 17396 -338 17430 -304
rect 17488 -338 17522 -304
rect 17580 -338 17614 -304
rect 17672 -338 17706 -304
rect 17764 -338 17798 -304
rect 17856 -338 17890 -304
rect 17948 -338 17982 -304
rect 18040 -338 18074 -304
rect 18132 -338 18166 -304
rect 18224 -338 18258 -304
rect 18316 -338 18350 -304
rect 18408 -338 18442 -304
rect 18500 -338 18534 -304
rect 18592 -338 18626 -304
rect 18684 -338 18718 -304
rect 18776 -338 18810 -304
rect 18868 -338 18902 -304
rect 18960 -338 18994 -304
rect 19052 -338 19086 -304
rect 19144 -338 19178 -304
rect 19236 -338 19270 -304
rect 19328 -338 19362 -304
rect 19420 -338 19454 -304
rect 19512 -338 19546 -304
rect 19604 -338 19638 -304
rect 19696 -338 19730 -304
rect 19788 -338 19822 -304
rect 19880 -338 19914 -304
rect 19972 -338 20006 -304
rect 20064 -338 20098 -304
rect 20156 -338 20190 -304
rect 20248 -338 20282 -304
rect 20340 -338 20374 -304
rect 20432 -338 20466 -304
rect 20586 -338 20620 -304
rect 20678 -338 20712 -304
rect 20770 -338 20804 -304
rect 20862 -338 20896 -304
rect 20954 -338 20988 -304
rect 21046 -338 21080 -304
rect 21138 -338 21172 -304
rect 21230 -338 21264 -304
rect 21322 -338 21356 -304
rect 21414 -338 21448 -304
rect 21506 -338 21540 -304
rect 21598 -338 21632 -304
rect 21690 -338 21724 -304
rect 21782 -338 21816 -304
rect 21874 -338 21908 -304
rect 21966 -338 22000 -304
rect 22058 -338 22092 -304
rect 22150 -338 22184 -304
rect 22242 -338 22276 -304
rect 22334 -338 22368 -304
rect 22426 -338 22460 -304
rect 22518 -338 22552 -304
rect 22610 -338 22644 -304
rect 22702 -338 22736 -304
rect 22794 -338 22828 -304
rect 22886 -338 22920 -304
rect 22978 -338 23012 -304
rect 23070 -338 23104 -304
rect 23162 -338 23196 -304
rect 23254 -338 23288 -304
rect 23346 -338 23380 -304
rect 23438 -338 23472 -304
rect 23530 -338 23564 -304
rect 23622 -338 23656 -304
rect 23714 -338 23748 -304
rect 23806 -338 23840 -304
rect 23898 -338 23932 -304
rect 23990 -338 24024 -304
rect 24082 -338 24116 -304
rect 24174 -338 24208 -304
rect 24266 -338 24300 -304
rect 24358 -338 24392 -304
rect 24450 -338 24484 -304
rect 24542 -338 24576 -304
rect 24634 -338 24668 -304
rect 24726 -338 24760 -304
rect 24818 -338 24852 -304
rect 24910 -338 24944 -304
rect 25002 -338 25036 -304
rect 25094 -338 25128 -304
rect 8604 -1026 8638 -992
rect 8696 -1026 8730 -992
rect 8788 -1026 8822 -992
rect 8880 -1026 8914 -992
rect 8972 -1026 9006 -992
rect 9064 -1026 9098 -992
rect 9156 -1026 9190 -992
rect 9248 -1026 9282 -992
rect 9340 -1026 9374 -992
rect 9432 -1026 9466 -992
rect 9524 -1026 9558 -992
rect 9616 -1026 9650 -992
rect 9708 -1026 9742 -992
rect 9800 -1026 9834 -992
rect 9892 -1026 9926 -992
rect 9984 -1026 10018 -992
rect 10076 -1026 10110 -992
rect 10168 -1026 10202 -992
rect 10260 -1026 10294 -992
rect 10352 -1026 10386 -992
rect 10444 -1026 10478 -992
rect 10536 -1026 10570 -992
rect 10628 -1026 10662 -992
rect 10720 -1026 10754 -992
rect 10812 -1026 10846 -992
rect 10904 -1026 10938 -992
rect 10996 -1026 11030 -992
rect 11088 -1026 11122 -992
rect 11180 -1026 11214 -992
rect 11272 -1026 11306 -992
rect 11364 -1026 11398 -992
rect 11456 -1026 11490 -992
rect 11548 -1026 11582 -992
rect 11640 -1026 11674 -992
rect 11732 -1026 11766 -992
rect 11824 -1026 11858 -992
rect 11916 -1026 11950 -992
rect 12008 -1026 12042 -992
rect 12100 -1026 12134 -992
rect 12192 -1026 12226 -992
rect 12284 -1026 12318 -992
rect 12376 -1026 12410 -992
rect 12468 -1026 12502 -992
rect 12560 -1026 12594 -992
rect 12652 -1026 12686 -992
rect 12744 -1026 12778 -992
rect 12836 -1026 12870 -992
rect 12928 -1026 12962 -992
rect 13020 -1026 13054 -992
rect 13112 -1026 13146 -992
rect 13204 -1026 13238 -992
rect 13296 -1026 13330 -992
rect 13388 -1026 13422 -992
rect 13480 -1026 13514 -992
rect 13572 -1026 13606 -992
rect 13664 -1026 13698 -992
rect 13756 -1026 13790 -992
rect 13848 -1026 13882 -992
rect 13940 -1026 13974 -992
rect 14032 -1026 14066 -992
rect 14124 -1026 14158 -992
rect 14216 -1026 14250 -992
rect 14308 -1026 14342 -992
rect 14400 -1026 14434 -992
rect 14492 -1026 14526 -992
rect 14584 -1026 14618 -992
rect 14676 -1026 14710 -992
rect 14768 -1026 14802 -992
rect 14860 -1026 14894 -992
rect 14952 -1026 14986 -992
rect 15044 -1026 15078 -992
rect 15136 -1026 15170 -992
rect 15228 -1026 15262 -992
rect 15320 -1026 15354 -992
rect 15412 -1026 15446 -992
rect 15504 -1026 15538 -992
rect 15596 -1026 15630 -992
rect 15688 -1026 15722 -992
rect 15780 -1026 15814 -992
rect 15872 -1026 15906 -992
rect 15964 -1026 15998 -992
rect 16056 -1026 16090 -992
rect 16148 -1026 16182 -992
rect 16240 -1026 16274 -992
rect 16332 -1026 16366 -992
rect 16424 -1026 16458 -992
rect 16516 -1026 16550 -992
rect 16608 -1026 16642 -992
rect 16700 -1026 16734 -992
rect 16792 -1026 16826 -992
rect 16884 -1026 16918 -992
rect 16976 -1026 17010 -992
rect 17068 -1026 17102 -992
rect 17160 -1026 17194 -992
rect 17252 -1026 17286 -992
rect 17344 -1026 17378 -992
rect 17436 -1026 17470 -992
rect 17528 -1026 17562 -992
rect 17620 -1026 17654 -992
rect 17712 -1026 17746 -992
rect 17804 -1026 17838 -992
rect 17896 -1026 17930 -992
rect 17988 -1026 18022 -992
rect 18080 -1026 18114 -992
rect 18172 -1026 18206 -992
rect 18264 -1026 18298 -992
rect 18356 -1026 18390 -992
rect 18448 -1026 18482 -992
rect 18540 -1026 18574 -992
rect 18632 -1026 18666 -992
rect 18724 -1026 18758 -992
rect 18816 -1026 18850 -992
rect 18908 -1026 18942 -992
rect 19000 -1026 19034 -992
rect 19092 -1026 19126 -992
rect 19184 -1026 19218 -992
rect 19276 -1026 19310 -992
rect 19368 -1026 19402 -992
rect 19460 -1026 19494 -992
rect 19552 -1026 19586 -992
rect 19644 -1026 19678 -992
rect 19736 -1026 19770 -992
rect 19828 -1026 19862 -992
rect 19920 -1026 19954 -992
rect 20012 -1026 20046 -992
rect 20104 -1026 20138 -992
rect 20196 -1026 20230 -992
rect 20288 -1026 20322 -992
rect 20380 -1026 20414 -992
rect 20472 -1026 20506 -992
rect 20564 -1026 20598 -992
rect 20656 -1026 20690 -992
rect 20748 -1026 20782 -992
rect 20840 -1026 20874 -992
rect 20932 -1026 20966 -992
rect 21024 -1026 21058 -992
rect 21116 -1026 21150 -992
rect 21208 -1026 21242 -992
rect 21300 -1026 21334 -992
rect 21392 -1026 21426 -992
rect 21484 -1026 21518 -992
rect 21576 -1026 21610 -992
rect 21668 -1026 21702 -992
rect 21760 -1026 21794 -992
rect 21852 -1026 21886 -992
rect 21944 -1026 21978 -992
rect 22036 -1026 22070 -992
rect 22128 -1026 22162 -992
rect 22220 -1026 22254 -992
rect 22312 -1026 22346 -992
rect 22404 -1026 22438 -992
rect 22496 -1026 22530 -992
rect 22588 -1026 22622 -992
rect 22680 -1026 22714 -992
rect 22772 -1026 22806 -992
rect 22864 -1026 22898 -992
rect 22956 -1026 22990 -992
rect 23048 -1026 23082 -992
rect 23140 -1026 23174 -992
rect 23232 -1026 23266 -992
rect 23324 -1026 23358 -992
rect 23416 -1026 23450 -992
rect 23508 -1026 23542 -992
rect 23600 -1026 23634 -992
rect 23692 -1026 23726 -992
rect 23784 -1026 23818 -992
rect 23876 -1026 23910 -992
rect 23968 -1026 24002 -992
rect 24060 -1026 24094 -992
rect 24152 -1026 24186 -992
rect 24244 -1026 24278 -992
rect 24336 -1026 24370 -992
rect 24428 -1026 24462 -992
rect 24520 -1026 24554 -992
rect 24612 -1026 24646 -992
rect 24704 -1026 24738 -992
rect 24796 -1026 24830 -992
rect 24888 -1026 24922 -992
rect 24980 -1026 25014 -992
rect 25072 -1026 25106 -992
rect 25164 -1026 25198 -992
rect 25256 -1026 25290 -992
rect 8604 -1715 8638 -1681
rect 8696 -1715 8730 -1681
rect 8788 -1715 8822 -1681
rect 8880 -1715 8914 -1681
rect 8972 -1715 9006 -1681
rect 9064 -1715 9098 -1681
rect 9156 -1715 9190 -1681
rect 9248 -1715 9282 -1681
rect 9340 -1715 9374 -1681
rect 9432 -1715 9466 -1681
rect 9524 -1715 9558 -1681
rect 9616 -1715 9650 -1681
rect 9708 -1715 9742 -1681
rect 9800 -1715 9834 -1681
rect 9892 -1715 9926 -1681
rect 9984 -1715 10018 -1681
rect 10076 -1715 10110 -1681
rect 10168 -1715 10202 -1681
rect 10260 -1715 10294 -1681
rect 10352 -1715 10386 -1681
rect 10444 -1715 10478 -1681
rect 10536 -1715 10570 -1681
rect 10628 -1715 10662 -1681
rect 10720 -1715 10754 -1681
rect 10812 -1715 10846 -1681
rect 10904 -1715 10938 -1681
rect 10996 -1715 11030 -1681
rect 11088 -1715 11122 -1681
rect 11180 -1715 11214 -1681
rect 11272 -1715 11306 -1681
rect 11364 -1715 11398 -1681
rect 11456 -1715 11490 -1681
rect 11548 -1715 11582 -1681
rect 11640 -1715 11674 -1681
rect 11732 -1715 11766 -1681
rect 11824 -1715 11858 -1681
rect 11916 -1715 11950 -1681
rect 12008 -1715 12042 -1681
rect 12100 -1715 12134 -1681
rect 12192 -1715 12226 -1681
rect 12284 -1715 12318 -1681
rect 12376 -1715 12410 -1681
rect 12468 -1715 12502 -1681
rect 12560 -1715 12594 -1681
rect 12652 -1715 12686 -1681
rect 12744 -1715 12778 -1681
rect 12836 -1715 12870 -1681
rect 12928 -1715 12962 -1681
rect 13020 -1715 13054 -1681
rect 13112 -1715 13146 -1681
rect 13204 -1715 13238 -1681
rect 13296 -1715 13330 -1681
rect 13388 -1715 13422 -1681
rect 13480 -1715 13514 -1681
rect 13572 -1715 13606 -1681
rect 13664 -1715 13698 -1681
rect 13756 -1715 13790 -1681
rect 13848 -1715 13882 -1681
rect 13940 -1715 13974 -1681
rect 14032 -1715 14066 -1681
rect 14124 -1715 14158 -1681
rect 14216 -1715 14250 -1681
rect 14308 -1715 14342 -1681
rect 14400 -1715 14434 -1681
rect 14492 -1715 14526 -1681
rect 14584 -1715 14618 -1681
rect 14676 -1715 14710 -1681
rect 14768 -1715 14802 -1681
rect 14860 -1715 14894 -1681
rect 14952 -1715 14986 -1681
rect 15044 -1715 15078 -1681
rect 15136 -1715 15170 -1681
rect 15228 -1715 15262 -1681
rect 15320 -1715 15354 -1681
rect 15412 -1715 15446 -1681
rect 15504 -1715 15538 -1681
rect 15596 -1715 15630 -1681
rect 15688 -1715 15722 -1681
rect 15780 -1715 15814 -1681
rect 15872 -1715 15906 -1681
rect 15964 -1715 15998 -1681
rect 16056 -1715 16090 -1681
rect 16148 -1715 16182 -1681
rect 16240 -1715 16274 -1681
rect 16332 -1715 16366 -1681
rect 16424 -1715 16458 -1681
rect 16516 -1715 16550 -1681
rect 16608 -1715 16642 -1681
rect 16700 -1715 16734 -1681
rect 16792 -1715 16826 -1681
rect 16884 -1715 16918 -1681
rect 16976 -1715 17010 -1681
rect 17068 -1715 17102 -1681
rect 17160 -1715 17194 -1681
rect 17252 -1715 17286 -1681
rect 17344 -1715 17378 -1681
rect 17436 -1715 17470 -1681
rect 17528 -1715 17562 -1681
rect 17620 -1715 17654 -1681
rect 17712 -1715 17746 -1681
rect 17804 -1715 17838 -1681
rect 17896 -1715 17930 -1681
rect 17988 -1715 18022 -1681
rect 18080 -1715 18114 -1681
rect 18172 -1715 18206 -1681
rect 18264 -1715 18298 -1681
rect 18356 -1715 18390 -1681
rect 18448 -1715 18482 -1681
rect 18540 -1715 18574 -1681
rect 18632 -1715 18666 -1681
rect 18724 -1715 18758 -1681
rect 18816 -1715 18850 -1681
rect 18908 -1715 18942 -1681
rect 19000 -1715 19034 -1681
rect 19092 -1715 19126 -1681
rect 19184 -1715 19218 -1681
rect 19276 -1715 19310 -1681
rect 19368 -1715 19402 -1681
rect 19460 -1715 19494 -1681
rect 19552 -1715 19586 -1681
rect 19644 -1715 19678 -1681
rect 19736 -1715 19770 -1681
rect 19828 -1715 19862 -1681
rect 19920 -1715 19954 -1681
rect 20012 -1715 20046 -1681
rect 20104 -1715 20138 -1681
rect 20196 -1715 20230 -1681
rect 20288 -1715 20322 -1681
rect 20380 -1715 20414 -1681
rect 20472 -1715 20506 -1681
rect 20564 -1715 20598 -1681
rect 20656 -1715 20690 -1681
rect 20748 -1715 20782 -1681
rect 20840 -1715 20874 -1681
rect 20932 -1715 20966 -1681
rect 21024 -1715 21058 -1681
rect 21116 -1715 21150 -1681
rect 21208 -1715 21242 -1681
rect 21300 -1715 21334 -1681
rect 21392 -1715 21426 -1681
rect 21484 -1715 21518 -1681
rect 21576 -1715 21610 -1681
rect 21668 -1715 21702 -1681
rect 21760 -1715 21794 -1681
rect 21852 -1715 21886 -1681
rect 21944 -1715 21978 -1681
rect 22036 -1715 22070 -1681
rect 22128 -1715 22162 -1681
rect 22220 -1715 22254 -1681
rect 22312 -1715 22346 -1681
rect 22404 -1715 22438 -1681
rect 22496 -1715 22530 -1681
rect 22588 -1715 22622 -1681
rect 22680 -1715 22714 -1681
rect 22772 -1715 22806 -1681
rect 22864 -1715 22898 -1681
rect 22956 -1715 22990 -1681
rect 23048 -1715 23082 -1681
rect 23140 -1715 23174 -1681
rect 23232 -1715 23266 -1681
rect 23324 -1715 23358 -1681
rect 23416 -1715 23450 -1681
rect 23508 -1715 23542 -1681
rect 23600 -1715 23634 -1681
rect 23692 -1715 23726 -1681
rect 23784 -1715 23818 -1681
rect 23876 -1715 23910 -1681
rect 23968 -1715 24002 -1681
rect 24060 -1715 24094 -1681
rect 24152 -1715 24186 -1681
rect 24244 -1715 24278 -1681
rect 24336 -1715 24370 -1681
rect 24428 -1715 24462 -1681
rect 24520 -1715 24554 -1681
rect 24612 -1715 24646 -1681
rect 24704 -1715 24738 -1681
rect 24796 -1715 24830 -1681
rect 24888 -1715 24922 -1681
rect 24980 -1715 25014 -1681
rect 25072 -1715 25106 -1681
rect 25164 -1715 25198 -1681
rect 25256 -1715 25290 -1681
<< nsubdiffcont >>
rect 14062 13571 14096 13605
rect 14142 13571 14176 13605
rect 14222 13571 14256 13605
rect 14302 13571 14336 13605
rect 14382 13571 14416 13605
rect 14462 13571 14496 13605
rect 14794 13574 14828 13608
rect 14874 13574 14908 13608
rect 14954 13574 14988 13608
rect 15034 13574 15068 13608
rect 15114 13574 15148 13608
rect 15194 13574 15228 13608
rect 15400 13574 15434 13608
rect 15480 13574 15514 13608
rect 15560 13574 15594 13608
rect 15640 13574 15674 13608
rect 15720 13574 15754 13608
rect 15800 13574 15834 13608
rect 16006 13574 16040 13608
rect 16086 13574 16120 13608
rect 16166 13574 16200 13608
rect 16246 13574 16280 13608
rect 16326 13574 16360 13608
rect 16406 13574 16440 13608
rect 16612 13574 16646 13608
rect 16692 13574 16726 13608
rect 16772 13574 16806 13608
rect 16852 13574 16886 13608
rect 16932 13574 16966 13608
rect 17012 13574 17046 13608
rect 17218 13574 17252 13608
rect 17298 13574 17332 13608
rect 17378 13574 17412 13608
rect 17458 13574 17492 13608
rect 17538 13574 17572 13608
rect 17618 13574 17652 13608
rect 17824 13574 17858 13608
rect 17904 13574 17938 13608
rect 17984 13574 18018 13608
rect 18064 13574 18098 13608
rect 18144 13574 18178 13608
rect 18224 13574 18258 13608
rect 18430 13574 18464 13608
rect 18510 13574 18544 13608
rect 18590 13574 18624 13608
rect 18670 13574 18704 13608
rect 18750 13574 18784 13608
rect 18830 13574 18864 13608
rect 19036 13574 19070 13608
rect 19116 13574 19150 13608
rect 19196 13574 19230 13608
rect 19276 13574 19310 13608
rect 19356 13574 19390 13608
rect 19436 13574 19470 13608
rect 19776 13523 19810 13557
rect 20253 13526 20287 13560
rect 20771 13571 20805 13605
rect 20851 13571 20885 13605
rect 20931 13571 20965 13605
rect 21011 13571 21045 13605
rect 21091 13571 21125 13605
rect 21171 13571 21205 13605
rect 21503 13574 21537 13608
rect 21583 13574 21617 13608
rect 21663 13574 21697 13608
rect 21743 13574 21777 13608
rect 21823 13574 21857 13608
rect 21903 13574 21937 13608
rect 22109 13574 22143 13608
rect 22189 13574 22223 13608
rect 22269 13574 22303 13608
rect 22349 13574 22383 13608
rect 22429 13574 22463 13608
rect 22509 13574 22543 13608
rect 22715 13574 22749 13608
rect 22795 13574 22829 13608
rect 22875 13574 22909 13608
rect 22955 13574 22989 13608
rect 23035 13574 23069 13608
rect 23115 13574 23149 13608
rect 23321 13574 23355 13608
rect 23401 13574 23435 13608
rect 23481 13574 23515 13608
rect 23561 13574 23595 13608
rect 23641 13574 23675 13608
rect 23721 13574 23755 13608
rect 23927 13574 23961 13608
rect 24007 13574 24041 13608
rect 24087 13574 24121 13608
rect 24167 13574 24201 13608
rect 24247 13574 24281 13608
rect 24327 13574 24361 13608
rect 24533 13574 24567 13608
rect 24613 13574 24647 13608
rect 24693 13574 24727 13608
rect 24773 13574 24807 13608
rect 24853 13574 24887 13608
rect 24933 13574 24967 13608
rect 25139 13574 25173 13608
rect 25219 13574 25253 13608
rect 25299 13574 25333 13608
rect 25379 13574 25413 13608
rect 25459 13574 25493 13608
rect 25539 13574 25573 13608
rect 25745 13574 25779 13608
rect 25825 13574 25859 13608
rect 25905 13574 25939 13608
rect 25985 13574 26019 13608
rect 26065 13574 26099 13608
rect 26145 13574 26179 13608
rect 26485 13523 26519 13557
rect 14029 13392 14063 13427
rect 19781 13379 19815 13413
rect 20242 13354 20276 13388
rect 20738 13392 20772 13427
rect 26490 13379 26524 13413
rect 19782 13227 19816 13261
rect 3174 13096 3208 13130
rect 3254 13096 3288 13130
rect 3334 13096 3368 13130
rect 3414 13096 3448 13130
rect 3494 13096 3528 13130
rect 3574 13096 3608 13130
rect 3906 13099 3940 13133
rect 3986 13099 4020 13133
rect 4066 13099 4100 13133
rect 4146 13099 4180 13133
rect 4226 13099 4260 13133
rect 4306 13099 4340 13133
rect 4512 13099 4546 13133
rect 4592 13099 4626 13133
rect 4672 13099 4706 13133
rect 4752 13099 4786 13133
rect 4832 13099 4866 13133
rect 4912 13099 4946 13133
rect 5118 13099 5152 13133
rect 5198 13099 5232 13133
rect 5278 13099 5312 13133
rect 5358 13099 5392 13133
rect 5438 13099 5472 13133
rect 5518 13099 5552 13133
rect 5724 13099 5758 13133
rect 5804 13099 5838 13133
rect 5884 13099 5918 13133
rect 5964 13099 5998 13133
rect 6044 13099 6078 13133
rect 6124 13099 6158 13133
rect 6330 13099 6364 13133
rect 6410 13099 6444 13133
rect 6490 13099 6524 13133
rect 6570 13099 6604 13133
rect 6650 13099 6684 13133
rect 6730 13099 6764 13133
rect 6936 13099 6970 13133
rect 7016 13099 7050 13133
rect 7096 13099 7130 13133
rect 7176 13099 7210 13133
rect 7256 13099 7290 13133
rect 7336 13099 7370 13133
rect 7542 13099 7576 13133
rect 7622 13099 7656 13133
rect 7702 13099 7736 13133
rect 7782 13099 7816 13133
rect 7862 13099 7896 13133
rect 7942 13099 7976 13133
rect 8148 13099 8182 13133
rect 8228 13099 8262 13133
rect 8308 13099 8342 13133
rect 8388 13099 8422 13133
rect 8468 13099 8502 13133
rect 8548 13099 8582 13133
rect 20242 13162 20276 13196
rect 26491 13227 26525 13261
rect 8888 13048 8922 13082
rect 19782 13057 19816 13091
rect 13348 13005 13382 13039
rect 13478 13005 13512 13039
rect 13624 13005 13658 13039
rect 3141 12917 3175 12952
rect 26491 13057 26525 13091
rect 20057 13005 20091 13039
rect 20187 13005 20221 13039
rect 20333 13005 20367 13039
rect 8893 12904 8927 12938
rect 8894 12752 8928 12786
rect 19781 12900 19815 12934
rect 26490 12900 26524 12934
rect 8894 12582 8928 12616
rect 2460 12530 2494 12564
rect 2590 12530 2624 12564
rect 2736 12530 2770 12564
rect 8893 12425 8927 12459
rect 9090 12159 9124 12193
rect 9182 12160 9216 12194
rect 9274 12160 9308 12194
rect 10911 11840 10945 11874
rect 11004 11839 11038 11873
rect 11096 11840 11130 11874
rect 11186 11841 11220 11875
rect 11281 11841 11315 11875
rect 11372 11842 11406 11876
rect 11463 11854 11497 11888
rect 11555 11854 11589 11888
rect 11647 11854 11681 11888
rect 11739 11854 11773 11888
rect 11831 11854 11865 11888
rect 11923 11854 11957 11888
rect 12015 11854 12049 11888
rect 12107 11854 12141 11888
rect 12199 11854 12233 11888
rect 12291 11854 12325 11888
rect 12383 11854 12417 11888
rect 12475 11854 12509 11888
rect 12567 11854 12601 11888
rect 12659 11854 12693 11888
rect 12751 11854 12785 11888
rect 12843 11854 12877 11888
rect 12935 11854 12969 11888
rect 13027 11854 13061 11888
rect 13119 11854 13153 11888
rect 13211 11854 13245 11888
rect 9152 8416 9186 8450
rect 9288 8420 9322 8454
rect 9406 8419 9440 8453
rect 9549 8419 9583 8453
rect 9624 8420 9658 8454
rect 9709 8421 9743 8455
rect 9811 8414 9845 8448
rect 9900 8416 9934 8450
rect 9997 8421 10031 8455
rect 10083 8410 10117 8444
rect 10175 8418 10209 8452
rect 10267 8417 10301 8451
rect 10355 8404 10389 8438
rect 10456 8406 10490 8440
rect 10544 8408 10578 8442
rect 10637 8409 10671 8443
rect 10733 8408 10767 8442
rect 10822 8412 10856 8446
rect 10919 8415 10953 8449
rect 11003 8411 11037 8445
rect 11093 8413 11127 8447
rect 11191 8409 11225 8443
rect 11462 8414 11496 8448
rect 11560 8414 11594 8448
rect 11643 8412 11677 8446
rect 8893 8187 8927 8221
rect 2460 8082 2494 8116
rect 2590 8082 2624 8116
rect 2736 8082 2770 8116
rect 8894 8030 8928 8064
rect 8894 7860 8928 7894
rect 12452 8337 12486 8371
rect 12531 8336 12565 8370
rect 13364 8175 13398 8209
rect 20073 8175 20107 8209
rect 19521 8070 19555 8104
rect 19667 8070 19701 8104
rect 19797 8070 19831 8104
rect 13363 8018 13397 8052
rect 26230 8070 26264 8104
rect 26376 8070 26410 8104
rect 26506 8070 26540 8104
rect 20072 8018 20106 8052
rect 3141 7694 3175 7729
rect 8893 7708 8927 7742
rect 8888 7564 8922 7598
rect 19650 7946 19684 7980
rect 12947 7884 12981 7918
rect 13363 7848 13397 7882
rect 20072 7848 20106 7882
rect 12939 7664 12973 7698
rect 13364 7696 13398 7730
rect 19650 7750 19684 7784
rect 19116 7682 19150 7717
rect 20073 7696 20107 7730
rect 25825 7682 25859 7717
rect 3174 7516 3208 7550
rect 3254 7516 3288 7550
rect 3334 7516 3368 7550
rect 3414 7516 3448 7550
rect 3494 7516 3528 7550
rect 3574 7516 3608 7550
rect 3906 7513 3940 7547
rect 3986 7513 4020 7547
rect 4066 7513 4100 7547
rect 4146 7513 4180 7547
rect 4226 7513 4260 7547
rect 4306 7513 4340 7547
rect 4512 7513 4546 7547
rect 4592 7513 4626 7547
rect 4672 7513 4706 7547
rect 4752 7513 4786 7547
rect 4832 7513 4866 7547
rect 4912 7513 4946 7547
rect 5118 7513 5152 7547
rect 5198 7513 5232 7547
rect 5278 7513 5312 7547
rect 5358 7513 5392 7547
rect 5438 7513 5472 7547
rect 5518 7513 5552 7547
rect 5724 7513 5758 7547
rect 5804 7513 5838 7547
rect 5884 7513 5918 7547
rect 5964 7513 5998 7547
rect 6044 7513 6078 7547
rect 6124 7513 6158 7547
rect 6330 7513 6364 7547
rect 6410 7513 6444 7547
rect 6490 7513 6524 7547
rect 6570 7513 6604 7547
rect 6650 7513 6684 7547
rect 6730 7513 6764 7547
rect 6936 7513 6970 7547
rect 7016 7513 7050 7547
rect 7096 7513 7130 7547
rect 7176 7513 7210 7547
rect 7256 7513 7290 7547
rect 7336 7513 7370 7547
rect 7542 7513 7576 7547
rect 7622 7513 7656 7547
rect 7702 7513 7736 7547
rect 7782 7513 7816 7547
rect 7862 7513 7896 7547
rect 7942 7513 7976 7547
rect 8148 7513 8182 7547
rect 8228 7513 8262 7547
rect 8308 7513 8342 7547
rect 8388 7513 8422 7547
rect 8468 7513 8502 7547
rect 8548 7513 8582 7547
rect 13369 7552 13403 7586
rect 13709 7501 13743 7535
rect 13789 7501 13823 7535
rect 13869 7501 13903 7535
rect 13949 7501 13983 7535
rect 14029 7501 14063 7535
rect 14109 7501 14143 7535
rect 14315 7501 14349 7535
rect 14395 7501 14429 7535
rect 14475 7501 14509 7535
rect 14555 7501 14589 7535
rect 14635 7501 14669 7535
rect 14715 7501 14749 7535
rect 14921 7501 14955 7535
rect 15001 7501 15035 7535
rect 15081 7501 15115 7535
rect 15161 7501 15195 7535
rect 15241 7501 15275 7535
rect 15321 7501 15355 7535
rect 15527 7501 15561 7535
rect 15607 7501 15641 7535
rect 15687 7501 15721 7535
rect 15767 7501 15801 7535
rect 15847 7501 15881 7535
rect 15927 7501 15961 7535
rect 16133 7501 16167 7535
rect 16213 7501 16247 7535
rect 16293 7501 16327 7535
rect 16373 7501 16407 7535
rect 16453 7501 16487 7535
rect 16533 7501 16567 7535
rect 16739 7501 16773 7535
rect 16819 7501 16853 7535
rect 16899 7501 16933 7535
rect 16979 7501 17013 7535
rect 17059 7501 17093 7535
rect 17139 7501 17173 7535
rect 17345 7501 17379 7535
rect 17425 7501 17459 7535
rect 17505 7501 17539 7535
rect 17585 7501 17619 7535
rect 17665 7501 17699 7535
rect 17745 7501 17779 7535
rect 17951 7501 17985 7535
rect 18031 7501 18065 7535
rect 18111 7501 18145 7535
rect 18191 7501 18225 7535
rect 18271 7501 18305 7535
rect 18351 7501 18385 7535
rect 18683 7504 18717 7538
rect 18763 7504 18797 7538
rect 18843 7504 18877 7538
rect 18923 7504 18957 7538
rect 19003 7504 19037 7538
rect 19083 7504 19117 7538
rect 19650 7575 19684 7609
rect 20078 7552 20112 7586
rect 20418 7501 20452 7535
rect 20498 7501 20532 7535
rect 20578 7501 20612 7535
rect 20658 7501 20692 7535
rect 20738 7501 20772 7535
rect 20818 7501 20852 7535
rect 21024 7501 21058 7535
rect 21104 7501 21138 7535
rect 21184 7501 21218 7535
rect 21264 7501 21298 7535
rect 21344 7501 21378 7535
rect 21424 7501 21458 7535
rect 21630 7501 21664 7535
rect 21710 7501 21744 7535
rect 21790 7501 21824 7535
rect 21870 7501 21904 7535
rect 21950 7501 21984 7535
rect 22030 7501 22064 7535
rect 22236 7501 22270 7535
rect 22316 7501 22350 7535
rect 22396 7501 22430 7535
rect 22476 7501 22510 7535
rect 22556 7501 22590 7535
rect 22636 7501 22670 7535
rect 22842 7501 22876 7535
rect 22922 7501 22956 7535
rect 23002 7501 23036 7535
rect 23082 7501 23116 7535
rect 23162 7501 23196 7535
rect 23242 7501 23276 7535
rect 23448 7501 23482 7535
rect 23528 7501 23562 7535
rect 23608 7501 23642 7535
rect 23688 7501 23722 7535
rect 23768 7501 23802 7535
rect 23848 7501 23882 7535
rect 24054 7501 24088 7535
rect 24134 7501 24168 7535
rect 24214 7501 24248 7535
rect 24294 7501 24328 7535
rect 24374 7501 24408 7535
rect 24454 7501 24488 7535
rect 24660 7501 24694 7535
rect 24740 7501 24774 7535
rect 24820 7501 24854 7535
rect 24900 7501 24934 7535
rect 24980 7501 25014 7535
rect 25060 7501 25094 7535
rect 25392 7504 25426 7538
rect 25472 7504 25506 7538
rect 25552 7504 25586 7538
rect 25632 7504 25666 7538
rect 25712 7504 25746 7538
rect 25792 7504 25826 7538
rect 24787 7274 24821 7308
rect 24867 7274 24901 7308
rect 24947 7274 24981 7308
rect 25027 7274 25061 7308
rect 25107 7274 25141 7308
rect 25187 7274 25221 7308
rect 25519 7277 25553 7311
rect 25599 7277 25633 7311
rect 25679 7277 25713 7311
rect 25759 7277 25793 7311
rect 25839 7277 25873 7311
rect 25919 7277 25953 7311
rect 26125 7277 26159 7311
rect 26205 7277 26239 7311
rect 26285 7277 26319 7311
rect 26365 7277 26399 7311
rect 26445 7277 26479 7311
rect 26525 7277 26559 7311
rect 26731 7277 26765 7311
rect 26811 7277 26845 7311
rect 26891 7277 26925 7311
rect 26971 7277 27005 7311
rect 27051 7277 27085 7311
rect 27131 7277 27165 7311
rect 27337 7277 27371 7311
rect 27417 7277 27451 7311
rect 27497 7277 27531 7311
rect 27577 7277 27611 7311
rect 27657 7277 27691 7311
rect 27737 7277 27771 7311
rect 27943 7277 27977 7311
rect 28023 7277 28057 7311
rect 28103 7277 28137 7311
rect 28183 7277 28217 7311
rect 28263 7277 28297 7311
rect 28343 7277 28377 7311
rect 28549 7277 28583 7311
rect 28629 7277 28663 7311
rect 28709 7277 28743 7311
rect 28789 7277 28823 7311
rect 28869 7277 28903 7311
rect 28949 7277 28983 7311
rect 29155 7277 29189 7311
rect 29235 7277 29269 7311
rect 29315 7277 29349 7311
rect 29395 7277 29429 7311
rect 29475 7277 29509 7311
rect 29555 7277 29589 7311
rect 29761 7277 29795 7311
rect 29841 7277 29875 7311
rect 29921 7277 29955 7311
rect 30001 7277 30035 7311
rect 30081 7277 30115 7311
rect 30161 7277 30195 7311
rect 30501 7226 30535 7260
rect 11527 7084 11561 7118
rect 11619 7084 11653 7118
rect 11711 7084 11745 7118
rect 11803 7084 11837 7118
rect 11895 7084 11929 7118
rect 11987 7084 12021 7118
rect 12079 7084 12113 7118
rect 12787 7084 12821 7118
rect 12879 7084 12913 7118
rect 12971 7084 13005 7118
rect 13063 7084 13097 7118
rect 13155 7084 13189 7118
rect 13247 7084 13281 7118
rect 13339 7084 13373 7118
rect 13431 7084 13465 7118
rect 13523 7084 13557 7118
rect 13615 7084 13649 7118
rect 13707 7084 13741 7118
rect 13799 7084 13833 7118
rect 13891 7084 13925 7118
rect 13983 7084 14017 7118
rect 14075 7084 14109 7118
rect 14167 7084 14201 7118
rect 14259 7084 14293 7118
rect 14351 7084 14385 7118
rect 14443 7084 14477 7118
rect 14535 7084 14569 7118
rect 24754 7095 24788 7130
rect 30506 7082 30540 7116
rect 30507 6930 30541 6964
rect 30507 6760 30541 6794
rect 24073 6708 24107 6742
rect 24203 6708 24237 6742
rect 24349 6708 24383 6742
rect 30506 6603 30540 6637
rect 30708 6335 30742 6369
rect 30891 6335 30925 6369
rect 11526 6211 11560 6245
rect 11618 6211 11652 6245
rect 11710 6211 11744 6245
rect 11802 6211 11836 6245
rect 11894 6211 11928 6245
rect 11986 6211 12020 6245
rect 12078 6211 12112 6245
rect 12170 6211 12204 6245
rect 12262 6211 12296 6245
rect 12354 6211 12388 6245
rect 12446 6211 12480 6245
rect 12538 6211 12572 6245
rect 12630 6211 12664 6245
rect 12722 6211 12756 6245
rect 12814 6211 12848 6245
rect 12906 6211 12940 6245
rect 12998 6211 13032 6245
rect 13090 6211 13124 6245
rect 13182 6211 13216 6245
rect 13274 6211 13308 6245
rect 13550 6211 13584 6245
rect 13642 6211 13676 6245
rect 13734 6211 13768 6245
rect 13826 6211 13860 6245
rect 13918 6211 13952 6245
rect 14010 6211 14044 6245
rect 14103 6211 14137 6245
rect 14194 6211 14228 6245
rect 14286 6211 14320 6245
rect 14378 6211 14412 6245
rect 14470 6211 14504 6245
rect 14746 6211 14780 6245
rect 14838 6211 14872 6245
rect 14930 6211 14964 6245
rect 15022 6211 15056 6245
rect 15114 6211 15148 6245
rect 15206 6211 15240 6245
rect 15298 6211 15332 6245
rect 15390 6211 15424 6245
rect 15482 6211 15516 6245
rect 15574 6211 15608 6245
rect 15666 6211 15700 6245
rect 15758 6211 15792 6245
rect 15850 6211 15884 6245
rect 15942 6211 15976 6245
rect 16034 6211 16068 6245
rect 16126 6211 16160 6245
rect 16218 6211 16252 6245
rect 16310 6211 16344 6245
rect 16402 6211 16436 6245
rect 16494 6211 16528 6245
rect 16586 6211 16620 6245
rect 16678 6211 16712 6245
rect 16770 6211 16804 6245
rect 16862 6211 16896 6245
rect 17138 6211 17172 6245
rect 17230 6211 17264 6245
rect 17322 6211 17356 6245
rect 17414 6211 17448 6245
rect 17506 6211 17540 6245
rect 17598 6211 17632 6245
rect 17690 6211 17724 6245
rect 17782 6211 17816 6245
rect 17874 6211 17908 6245
rect 17966 6211 18000 6245
rect 18058 6211 18092 6245
rect 18150 6211 18184 6245
rect 18242 6211 18276 6245
rect 18334 6211 18368 6245
rect 18426 6211 18460 6245
rect 18518 6211 18552 6245
rect 18610 6211 18644 6245
rect 18702 6211 18736 6245
rect 18794 6211 18828 6245
rect 18886 6211 18920 6245
rect 18978 6211 19012 6245
rect 19070 6211 19104 6245
rect 19162 6211 19196 6245
rect 19254 6211 19288 6245
rect 19530 6211 19564 6245
rect 19622 6211 19656 6245
rect 19714 6211 19748 6245
rect 19806 6211 19840 6245
rect 19898 6211 19932 6245
rect 19990 6211 20024 6245
rect 20082 6211 20116 6245
rect 20174 6211 20208 6245
rect 20266 6211 20300 6245
rect 20358 6211 20392 6245
rect 20450 6211 20484 6245
rect 20542 6211 20576 6245
rect 20634 6211 20668 6245
rect 20726 6211 20760 6245
rect 20818 6211 20852 6245
rect 20910 6211 20944 6245
rect 21002 6211 21036 6245
rect 21094 6211 21128 6245
rect 21186 6211 21220 6245
rect 21278 6211 21312 6245
rect 21370 6211 21404 6245
rect 21462 6211 21496 6245
rect 21554 6211 21588 6245
rect 21646 6211 21680 6245
rect 21922 6211 21956 6245
rect 22014 6211 22048 6245
rect 22106 6211 22140 6245
rect 22198 6211 22232 6245
rect 22290 6211 22324 6245
rect 22382 6211 22416 6245
rect 22474 6211 22508 6245
rect 22566 6211 22600 6245
rect 22658 6211 22692 6245
rect 22750 6211 22784 6245
rect 22842 6211 22876 6245
rect 22934 6211 22968 6245
rect 23026 6211 23060 6245
rect 23118 6211 23152 6245
rect 23210 6211 23244 6245
rect 23302 6211 23336 6245
rect 23394 6211 23428 6245
rect 11086 5522 11120 5556
rect 11178 5522 11212 5556
rect 11270 5522 11304 5556
rect 11362 5522 11396 5556
rect 11454 5522 11488 5556
rect 11546 5522 11580 5556
rect 11638 5522 11672 5556
rect 11730 5522 11764 5556
rect 11822 5522 11856 5556
rect 11914 5522 11948 5556
rect 12006 5522 12040 5556
rect 12098 5522 12132 5556
rect 12190 5522 12224 5556
rect 12282 5522 12316 5556
rect 12374 5522 12408 5556
rect 12466 5522 12500 5556
rect 12558 5522 12592 5556
rect 12650 5522 12684 5556
rect 12742 5522 12776 5556
rect 12814 5522 12868 5556
rect 12906 5522 12940 5556
rect 12998 5522 13032 5556
rect 13090 5522 13124 5556
rect 13182 5522 13216 5556
rect 13274 5522 13308 5556
rect 13366 5522 13400 5556
rect 13458 5522 13492 5556
rect 13550 5522 13584 5556
rect 13642 5522 13676 5556
rect 13734 5522 13768 5556
rect 13826 5522 13860 5556
rect 13918 5522 13952 5556
rect 14010 5522 14044 5556
rect 14102 5522 14136 5556
rect 14194 5522 14228 5556
rect 14286 5522 14320 5556
rect 14378 5522 14412 5556
rect 14470 5522 14504 5556
rect 14562 5522 14596 5556
rect 14838 5522 14872 5556
rect 14930 5522 14964 5556
rect 15022 5522 15056 5556
rect 15114 5522 15148 5556
rect 15206 5522 15240 5556
rect 15298 5522 15332 5556
rect 15390 5522 15424 5556
rect 15482 5522 15516 5556
rect 15574 5522 15608 5556
rect 15666 5522 15700 5556
rect 15758 5522 15792 5556
rect 15850 5522 15884 5556
rect 15942 5522 15976 5556
rect 16034 5522 16068 5556
rect 16126 5522 16160 5556
rect 16218 5522 16252 5556
rect 16310 5522 16344 5556
rect 16402 5522 16436 5556
rect 16494 5522 16528 5556
rect 16586 5522 16620 5556
rect 16678 5522 16712 5556
rect 16770 5522 16804 5556
rect 16862 5522 16896 5556
rect 16954 5522 16988 5556
rect 17230 5522 17264 5556
rect 17322 5522 17356 5556
rect 17414 5522 17448 5556
rect 17506 5522 17540 5556
rect 17598 5522 17632 5556
rect 17690 5522 17724 5556
rect 17782 5522 17816 5556
rect 17874 5522 17908 5556
rect 17966 5522 18000 5556
rect 18058 5522 18092 5556
rect 18150 5522 18184 5556
rect 18242 5522 18276 5556
rect 18334 5522 18368 5556
rect 18426 5522 18460 5556
rect 18518 5522 18552 5556
rect 18610 5522 18644 5556
rect 18702 5522 18736 5556
rect 18794 5522 18828 5556
rect 18886 5522 18920 5556
rect 18978 5522 19012 5556
rect 19070 5522 19104 5556
rect 19162 5522 19196 5556
rect 19254 5522 19288 5556
rect 19346 5522 19380 5556
rect 19622 5522 19656 5556
rect 19714 5522 19748 5556
rect 19806 5522 19840 5556
rect 19898 5522 19932 5556
rect 19990 5522 20024 5556
rect 20082 5522 20116 5556
rect 20174 5522 20208 5556
rect 20266 5522 20300 5556
rect 20358 5522 20392 5556
rect 20450 5522 20484 5556
rect 20542 5522 20576 5556
rect 20634 5522 20668 5556
rect 20726 5522 20760 5556
rect 20818 5522 20852 5556
rect 20910 5522 20944 5556
rect 21002 5522 21036 5556
rect 21094 5522 21128 5556
rect 21186 5522 21220 5556
rect 21278 5522 21312 5556
rect 21370 5522 21404 5556
rect 21462 5522 21496 5556
rect 21554 5522 21588 5556
rect 21646 5522 21680 5556
rect 21738 5522 21772 5556
rect 22014 5522 22048 5556
rect 22106 5522 22140 5556
rect 22198 5522 22232 5556
rect 22290 5522 22324 5556
rect 22382 5522 22416 5556
rect 22474 5522 22508 5556
rect 22566 5522 22600 5556
rect 22658 5522 22692 5556
rect 22750 5522 22784 5556
rect 22842 5522 22876 5556
rect 22934 5522 22968 5556
rect 23026 5522 23060 5556
rect 23118 5522 23152 5556
rect 23210 5522 23244 5556
rect 23302 5522 23336 5556
rect 23394 5522 23428 5556
rect 11118 4658 11152 4692
rect 11210 4658 11244 4692
rect 11302 4658 11336 4692
rect 11394 4658 11428 4692
rect 11486 4658 11520 4692
rect 11577 4658 11611 4692
rect 11669 4658 11703 4692
rect 11762 4658 11796 4692
rect 11854 4658 11888 4692
rect 13660 4649 13694 4683
rect 13752 4649 13786 4683
rect 13844 4649 13878 4683
rect 13936 4649 13970 4683
rect 14028 4649 14062 4683
rect 14120 4649 14154 4683
rect 14212 4649 14246 4683
rect 14304 4649 14338 4683
rect 14396 4649 14430 4683
rect 14488 4649 14522 4683
rect 14580 4649 14614 4683
rect 14672 4649 14706 4683
rect 14764 4649 14798 4683
rect 14856 4649 14890 4683
rect 14948 4649 14982 4683
rect 15040 4649 15074 4683
rect 15132 4649 15166 4683
rect 15224 4649 15258 4683
rect 15316 4649 15350 4683
rect 15408 4649 15442 4683
rect 15481 4649 15515 4683
rect 15573 4649 15607 4683
rect 15665 4649 15699 4683
rect 15757 4649 15791 4683
rect 15849 4649 15883 4683
rect 15941 4649 15975 4683
rect 16033 4649 16067 4683
rect 16125 4649 16159 4683
rect 16217 4649 16251 4683
rect 16309 4649 16343 4683
rect 16401 4649 16435 4683
rect 16493 4649 16527 4683
rect 16585 4649 16619 4683
rect 16677 4649 16711 4683
rect 16769 4649 16803 4683
rect 16861 4649 16895 4683
rect 16953 4649 16987 4683
rect 17045 4649 17079 4683
rect 17137 4649 17171 4683
rect 17229 4649 17263 4683
rect 17321 4649 17355 4683
rect 17413 4649 17447 4683
rect 17505 4649 17539 4683
rect 17597 4649 17631 4683
rect 17689 4649 17723 4683
rect 17781 4649 17815 4683
rect 17873 4649 17907 4683
rect 17965 4649 17999 4683
rect 18057 4649 18091 4683
rect 18149 4649 18183 4683
rect 18241 4649 18275 4683
rect 18333 4649 18367 4683
rect 18425 4649 18459 4683
rect 18517 4649 18551 4683
rect 18609 4649 18643 4683
rect 18701 4649 18735 4683
rect 18793 4649 18827 4683
rect 18885 4649 18919 4683
rect 18977 4649 19011 4683
rect 19069 4649 19103 4683
rect 19161 4649 19195 4683
rect 19253 4649 19287 4683
rect 19345 4649 19379 4683
rect 19437 4649 19471 4683
rect 19529 4649 19563 4683
rect 19621 4649 19655 4683
rect 19713 4649 19747 4683
rect 19805 4649 19839 4683
rect 19897 4649 19931 4683
rect 19989 4649 20023 4683
rect 20081 4649 20115 4683
rect 20173 4649 20207 4683
rect 20265 4649 20299 4683
rect 20357 4649 20391 4683
rect 20449 4649 20483 4683
rect 20541 4649 20575 4683
rect 20633 4649 20667 4683
rect 20725 4649 20759 4683
rect 20817 4649 20851 4683
rect 20909 4649 20943 4683
rect 21001 4649 21035 4683
rect 21093 4649 21127 4683
rect 21185 4649 21219 4683
rect 21277 4649 21311 4683
rect 21369 4649 21403 4683
rect 21461 4649 21495 4683
rect 21553 4649 21587 4683
rect 21645 4649 21679 4683
rect 21737 4649 21771 4683
rect 21829 4649 21863 4683
rect 21921 4649 21955 4683
rect 22013 4649 22047 4683
rect 22105 4649 22139 4683
rect 22197 4649 22231 4683
rect 22289 4649 22323 4683
rect 22381 4649 22415 4683
rect 22473 4649 22507 4683
rect 22565 4649 22599 4683
rect 22657 4649 22691 4683
rect 22749 4649 22783 4683
rect 22841 4649 22875 4683
rect 22933 4649 22967 4683
rect 23025 4649 23059 4683
rect 23117 4649 23151 4683
rect 23209 4649 23243 4683
rect 23301 4649 23335 4683
rect 23393 4649 23427 4683
rect 11525 3776 11559 3810
rect 11617 3776 11651 3810
rect 11709 3776 11743 3810
rect 11801 3776 11835 3810
rect 11893 3776 11927 3810
rect 11985 3776 12019 3810
rect 12077 3776 12111 3810
rect 12169 3776 12203 3810
rect 12261 3776 12295 3810
rect 12353 3776 12387 3810
rect 12445 3776 12479 3810
rect 12537 3776 12571 3810
rect 12629 3776 12663 3810
rect 12721 3776 12755 3810
rect 12813 3776 12847 3810
rect 12905 3776 12939 3810
rect 12997 3776 13031 3810
rect 13089 3776 13123 3810
rect 13181 3776 13215 3810
rect 13273 3776 13307 3810
rect 13365 3776 13399 3810
rect 13457 3776 13491 3810
rect 13549 3776 13583 3810
rect 13641 3776 13675 3810
rect 13733 3776 13767 3810
rect 13825 3776 13859 3810
rect 13917 3776 13951 3810
rect 14009 3776 14043 3810
rect 14101 3776 14135 3810
rect 14193 3776 14227 3810
rect 14285 3776 14319 3810
rect 14377 3776 14411 3810
rect 14469 3776 14503 3810
rect 14561 3776 14595 3810
rect 14653 3776 14687 3810
rect 14745 3776 14779 3810
rect 14837 3776 14871 3810
rect 14929 3776 14963 3810
rect 15021 3776 15055 3810
rect 15113 3776 15147 3810
rect 15205 3776 15239 3810
rect 15297 3776 15331 3810
rect 15389 3776 15423 3810
rect 15481 3776 15515 3810
rect 15573 3776 15607 3810
rect 15665 3776 15699 3810
rect 15757 3776 15791 3810
rect 15849 3776 15883 3810
rect 15941 3776 15975 3810
rect 16033 3776 16067 3810
rect 16125 3776 16159 3810
rect 16217 3776 16251 3810
rect 16309 3776 16343 3810
rect 16401 3776 16435 3810
rect 16493 3776 16527 3810
rect 16585 3776 16619 3810
rect 16677 3776 16711 3810
rect 16769 3776 16803 3810
rect 16861 3776 16895 3810
rect 16953 3776 16987 3810
rect 17045 3776 17079 3810
rect 17137 3776 17171 3810
rect 17229 3776 17263 3810
rect 17321 3776 17355 3810
rect 17413 3776 17447 3810
rect 17505 3776 17539 3810
rect 17597 3776 17631 3810
rect 17689 3776 17723 3810
rect 17781 3776 17815 3810
rect 17873 3776 17907 3810
rect 17965 3776 17999 3810
rect 18057 3776 18091 3810
rect 18149 3776 18183 3810
rect 18241 3776 18275 3810
rect 18333 3776 18367 3810
rect 18425 3776 18459 3810
rect 18517 3776 18551 3810
rect 18609 3776 18643 3810
rect 18701 3776 18735 3810
rect 18793 3776 18827 3810
rect 18885 3776 18919 3810
rect 18977 3776 19011 3810
rect 19069 3776 19103 3810
rect 19161 3776 19195 3810
rect 19253 3776 19287 3810
rect 19345 3776 19379 3810
rect 19437 3776 19471 3810
rect 19529 3776 19563 3810
rect 19621 3776 19655 3810
rect 19713 3776 19747 3810
rect 19805 3776 19839 3810
rect 19897 3776 19931 3810
rect 19989 3776 20023 3810
rect 20081 3776 20115 3810
rect 20173 3776 20207 3810
rect 20265 3776 20299 3810
rect 20357 3776 20391 3810
rect 20449 3776 20483 3810
rect 20541 3776 20575 3810
rect 20633 3776 20667 3810
rect 20725 3776 20759 3810
rect 20817 3776 20851 3810
rect 20909 3776 20943 3810
rect 21001 3776 21035 3810
rect 21093 3776 21127 3810
rect 21185 3776 21219 3810
rect 21277 3776 21311 3810
rect 21369 3776 21403 3810
rect 21461 3776 21495 3810
rect 21553 3776 21587 3810
rect 21645 3776 21679 3810
rect 21737 3776 21771 3810
rect 21829 3776 21863 3810
rect 21921 3776 21955 3810
rect 22013 3776 22047 3810
rect 22105 3776 22139 3810
rect 22197 3776 22231 3810
rect 22289 3776 22323 3810
rect 22381 3776 22415 3810
rect 22473 3776 22507 3810
rect 22565 3776 22599 3810
rect 22657 3776 22691 3810
rect 22749 3776 22783 3810
rect 22841 3776 22875 3810
rect 22933 3776 22967 3810
rect 23025 3776 23059 3810
rect 23117 3776 23151 3810
rect 23209 3776 23243 3810
rect 23301 3776 23335 3810
rect 23393 3776 23427 3810
rect 25607 3672 25641 3706
rect 25698 3672 25732 3706
rect 25791 3672 25825 3706
rect 25882 3672 25916 3706
rect 25973 3672 26007 3706
rect 26067 3672 26101 3706
rect 26158 3672 26192 3706
rect 26251 3672 26285 3706
rect 26342 3672 26376 3706
rect 26434 3672 26468 3706
rect 26525 3672 26559 3706
rect 26618 3672 26652 3706
rect 26711 3672 26745 3706
rect 26802 3672 26836 3706
rect 26894 3672 26928 3706
rect 26986 3672 27020 3706
rect 27078 3672 27112 3706
rect 27170 3672 27204 3706
rect 27262 3672 27296 3706
rect 27354 3672 27388 3706
rect 27447 3672 27481 3706
rect 27537 3672 27571 3706
rect 27630 3672 27664 3706
rect 27723 3672 27757 3706
rect 27815 3672 27849 3706
rect 27906 3672 27940 3706
rect 27999 3672 28033 3706
rect 28091 3672 28125 3706
rect 28183 3672 28217 3706
rect 28275 3672 28309 3706
rect 28367 3672 28401 3706
rect 28459 3672 28493 3706
rect 28550 3672 28584 3706
rect 28641 3672 28675 3706
rect 28734 3672 28768 3706
rect 28827 3672 28861 3706
rect 28919 3672 28953 3706
rect 29010 3672 29044 3706
rect 29104 3672 29138 3706
rect 29194 3672 29228 3706
rect 29285 3672 29319 3706
rect 29378 3672 29412 3706
rect 29471 3672 29505 3706
rect 29563 3672 29597 3706
rect 29654 3672 29688 3706
rect 29746 3672 29780 3706
rect 29838 3672 29872 3706
rect 29929 3672 29963 3706
rect 30021 3672 30055 3706
rect 30114 3672 30148 3706
rect 30206 3672 30240 3706
rect 30298 3672 30332 3706
rect 25609 2391 25643 2425
rect 25699 2391 25733 2425
rect 25792 2391 25826 2425
rect 25882 2391 25916 2425
rect 25973 2391 26007 2425
rect 26067 2391 26101 2425
rect 26158 2391 26192 2425
rect 26250 2391 26284 2425
rect 26342 2391 26376 2425
rect 26435 2391 26469 2425
rect 26526 2391 26560 2425
rect 26618 2391 26652 2425
rect 26710 2391 26744 2425
rect 26802 2391 26836 2425
rect 26895 2391 26929 2425
rect 26986 2391 27020 2425
rect 27077 2391 27111 2425
rect 27170 2391 27204 2425
rect 27263 2391 27297 2425
rect 27354 2391 27388 2425
rect 27446 2391 27480 2425
rect 27538 2391 27572 2425
rect 27630 2391 27664 2425
rect 27723 2391 27757 2425
rect 27813 2391 27847 2425
rect 27906 2391 27940 2425
rect 27998 2391 28032 2425
rect 28091 2391 28125 2425
rect 28185 2391 28219 2425
rect 28274 2391 28308 2425
rect 28366 2391 28400 2425
rect 28458 2391 28492 2425
rect 28550 2391 28584 2425
rect 28642 2391 28676 2425
rect 28734 2391 28768 2425
rect 28826 2391 28860 2425
rect 28918 2391 28952 2425
rect 29010 2391 29044 2425
rect 29102 2391 29136 2425
rect 29194 2391 29228 2425
rect 29286 2391 29320 2425
rect 29378 2391 29412 2425
rect 29470 2391 29504 2425
rect 29562 2391 29596 2425
rect 29654 2391 29688 2425
rect 29746 2391 29780 2425
rect 29838 2391 29872 2425
rect 29930 2391 29964 2425
rect 30022 2391 30056 2425
rect 30114 2391 30148 2425
rect 30207 2391 30241 2425
rect 30298 2391 30332 2425
rect 8606 1396 8640 1430
rect 8698 1396 8732 1430
rect 8790 1396 8824 1430
rect 8882 1396 8916 1430
rect 8974 1396 9008 1430
rect 9066 1396 9100 1430
rect 9158 1396 9192 1430
rect 9250 1396 9284 1430
rect 9342 1396 9376 1430
rect 9434 1396 9468 1430
rect 9526 1396 9560 1430
rect 9618 1396 9652 1430
rect 9710 1396 9744 1430
rect 9802 1396 9836 1430
rect 9894 1396 9928 1430
rect 9986 1396 10020 1430
rect 10078 1396 10112 1430
rect 10170 1396 10204 1430
rect 10262 1396 10296 1430
rect 10354 1396 10388 1430
rect 10446 1396 10480 1430
rect 10538 1396 10572 1430
rect 10630 1396 10664 1430
rect 10722 1396 10756 1430
rect 10814 1396 10848 1430
rect 10906 1396 10940 1430
rect 10998 1396 11032 1430
rect 11090 1396 11124 1430
rect 11182 1396 11216 1430
rect 11274 1396 11308 1430
rect 11366 1396 11400 1430
rect 12990 1396 13024 1430
rect 13082 1396 13116 1430
rect 13174 1396 13208 1430
rect 13266 1396 13300 1430
rect 13358 1396 13392 1430
rect 13450 1396 13484 1430
rect 13542 1396 13576 1430
rect 13634 1396 13668 1430
rect 13726 1396 13760 1430
rect 13818 1396 13852 1430
rect 13910 1396 13944 1430
rect 14002 1396 14036 1430
rect 14094 1396 14128 1430
rect 14186 1396 14220 1430
rect 14278 1396 14312 1430
rect 14370 1396 14404 1430
rect 14462 1396 14496 1430
rect 14554 1396 14588 1430
rect 14646 1396 14680 1430
rect 14738 1396 14772 1430
rect 14830 1396 14864 1430
rect 14922 1396 14956 1430
rect 15014 1396 15048 1430
rect 15106 1396 15140 1430
rect 15198 1396 15232 1430
rect 15290 1396 15324 1430
rect 15382 1396 15416 1430
rect 15474 1396 15508 1430
rect 15566 1396 15600 1430
rect 15658 1396 15692 1430
rect 15750 1396 15784 1430
rect 8604 254 8638 288
rect 8696 254 8730 288
rect 8788 254 8822 288
rect 8880 254 8914 288
rect 8972 254 9006 288
rect 9064 254 9098 288
rect 9156 254 9190 288
rect 9248 254 9282 288
rect 9340 254 9374 288
rect 9432 254 9466 288
rect 9524 254 9558 288
rect 9616 254 9650 288
rect 9708 254 9742 288
rect 9800 254 9834 288
rect 9892 254 9926 288
rect 9984 254 10018 288
rect 10076 254 10110 288
rect 10168 254 10202 288
rect 10260 254 10294 288
rect 10352 254 10386 288
rect 10444 254 10478 288
rect 10536 254 10570 288
rect 10628 254 10662 288
rect 10720 254 10754 288
rect 10812 254 10846 288
rect 10904 254 10938 288
rect 10996 254 11030 288
rect 11088 254 11122 288
rect 11180 254 11214 288
rect 11272 254 11306 288
rect 11364 254 11398 288
rect 11456 254 11490 288
rect 11548 254 11582 288
rect 11640 254 11674 288
rect 11732 254 11766 288
rect 11824 254 11858 288
rect 11916 254 11950 288
rect 12008 254 12042 288
rect 12100 254 12134 288
rect 12192 254 12226 288
rect 12284 254 12318 288
rect 12376 254 12410 288
rect 12468 254 12502 288
rect 12560 254 12594 288
rect 12652 254 12686 288
rect 12744 254 12778 288
rect 12836 254 12870 288
rect 12928 254 12962 288
rect 13020 254 13054 288
rect 13112 254 13146 288
rect 13204 254 13238 288
rect 13296 254 13330 288
rect 13388 254 13422 288
rect 13480 254 13514 288
rect 13572 254 13606 288
rect 13664 254 13698 288
rect 13756 254 13790 288
rect 13848 254 13882 288
rect 13940 254 13974 288
rect 14032 254 14066 288
rect 14124 254 14158 288
rect 14216 254 14250 288
rect 14820 254 14854 288
rect 14912 254 14946 288
rect 15004 254 15038 288
rect 15096 254 15130 288
rect 15188 254 15222 288
rect 15280 254 15314 288
rect 15372 254 15406 288
rect 15464 254 15498 288
rect 15556 254 15590 288
rect 15648 254 15682 288
rect 15740 254 15774 288
rect 15832 254 15866 288
rect 15924 254 15958 288
rect 16016 254 16050 288
rect 16108 254 16142 288
rect 16200 254 16234 288
rect 16292 254 16326 288
rect 16384 254 16418 288
rect 16476 254 16510 288
rect 16568 254 16602 288
rect 16660 254 16694 288
rect 16752 254 16786 288
rect 16844 254 16878 288
rect 16936 254 16970 288
rect 17028 254 17062 288
rect 17120 254 17154 288
rect 17212 254 17246 288
rect 17304 254 17338 288
rect 17396 254 17430 288
rect 17488 254 17522 288
rect 17580 254 17614 288
rect 17672 254 17706 288
rect 17764 254 17798 288
rect 17856 254 17890 288
rect 17948 254 17982 288
rect 18040 254 18074 288
rect 18132 254 18166 288
rect 18224 254 18258 288
rect 18316 254 18350 288
rect 18408 254 18442 288
rect 18500 254 18534 288
rect 18592 254 18626 288
rect 18684 254 18718 288
rect 18776 254 18810 288
rect 18868 254 18902 288
rect 18960 254 18994 288
rect 19052 254 19086 288
rect 19144 254 19178 288
rect 19236 254 19270 288
rect 19328 254 19362 288
rect 19420 254 19454 288
rect 19512 254 19546 288
rect 19604 254 19638 288
rect 19696 254 19730 288
rect 19788 254 19822 288
rect 19880 254 19914 288
rect 19972 254 20006 288
rect 20064 254 20098 288
rect 20156 254 20190 288
rect 20248 254 20282 288
rect 20340 254 20374 288
rect 20432 254 20466 288
rect 20586 254 20620 288
rect 20678 254 20712 288
rect 20770 254 20804 288
rect 20862 254 20896 288
rect 20954 254 20988 288
rect 21046 254 21080 288
rect 21138 254 21172 288
rect 21230 254 21264 288
rect 21322 254 21356 288
rect 21414 254 21448 288
rect 21506 254 21540 288
rect 21598 254 21632 288
rect 21690 254 21724 288
rect 21782 254 21816 288
rect 21874 254 21908 288
rect 21966 254 22000 288
rect 22058 254 22092 288
rect 22150 254 22184 288
rect 22242 254 22276 288
rect 22334 254 22368 288
rect 22426 254 22460 288
rect 22518 254 22552 288
rect 22610 254 22644 288
rect 22702 254 22736 288
rect 22794 254 22828 288
rect 22886 254 22920 288
rect 22978 254 23012 288
rect 23070 254 23104 288
rect 23162 254 23196 288
rect 23254 254 23288 288
rect 23346 254 23380 288
rect 23438 254 23472 288
rect 23530 254 23564 288
rect 23622 254 23656 288
rect 23714 254 23748 288
rect 23806 254 23840 288
rect 23898 254 23932 288
rect 23990 254 24024 288
rect 24082 254 24116 288
rect 24174 254 24208 288
rect 24266 254 24300 288
rect 24358 254 24392 288
rect 24450 254 24484 288
rect 24542 254 24576 288
rect 24634 254 24668 288
rect 24726 254 24760 288
rect 24818 254 24852 288
rect 24910 254 24944 288
rect 25002 254 25036 288
rect 25094 254 25128 288
rect 8604 -434 8638 -400
rect 8696 -434 8730 -400
rect 8788 -434 8822 -400
rect 8880 -434 8914 -400
rect 8972 -434 9006 -400
rect 9064 -434 9098 -400
rect 9156 -434 9190 -400
rect 9248 -434 9282 -400
rect 9340 -434 9374 -400
rect 9432 -434 9466 -400
rect 9524 -434 9558 -400
rect 9616 -434 9650 -400
rect 9708 -434 9742 -400
rect 9800 -434 9834 -400
rect 9892 -434 9926 -400
rect 9984 -434 10018 -400
rect 10076 -434 10110 -400
rect 10168 -434 10202 -400
rect 10260 -434 10294 -400
rect 10352 -434 10386 -400
rect 10628 -434 10662 -400
rect 10720 -434 10754 -400
rect 10812 -434 10846 -400
rect 10904 -434 10938 -400
rect 10996 -434 11030 -400
rect 11088 -434 11122 -400
rect 11180 -434 11214 -400
rect 11272 -434 11306 -400
rect 11364 -434 11398 -400
rect 11456 -434 11490 -400
rect 11548 -434 11582 -400
rect 11640 -434 11674 -400
rect 11732 -434 11766 -400
rect 11824 -434 11858 -400
rect 11916 -434 11950 -400
rect 12008 -434 12042 -400
rect 12100 -434 12134 -400
rect 12192 -434 12226 -400
rect 12284 -434 12318 -400
rect 12376 -434 12410 -400
rect 12468 -434 12502 -400
rect 12560 -434 12594 -400
rect 12652 -434 12686 -400
rect 12744 -434 12778 -400
rect 13020 -434 13054 -400
rect 13112 -434 13146 -400
rect 13204 -434 13238 -400
rect 13296 -434 13330 -400
rect 13388 -434 13422 -400
rect 13480 -434 13514 -400
rect 13572 -434 13606 -400
rect 13664 -434 13698 -400
rect 13756 -434 13790 -400
rect 13848 -434 13882 -400
rect 13940 -434 13974 -400
rect 14032 -434 14066 -400
rect 14124 -434 14158 -400
rect 14216 -434 14250 -400
rect 14308 -434 14342 -400
rect 14400 -434 14434 -400
rect 14492 -434 14526 -400
rect 14584 -434 14618 -400
rect 14676 -434 14710 -400
rect 14768 -434 14802 -400
rect 14860 -434 14894 -400
rect 14952 -434 14986 -400
rect 15044 -434 15078 -400
rect 15136 -434 15170 -400
rect 15412 -434 15446 -400
rect 15504 -434 15538 -400
rect 15596 -434 15630 -400
rect 15688 -434 15722 -400
rect 15780 -434 15814 -400
rect 15872 -434 15906 -400
rect 15964 -434 15998 -400
rect 16056 -434 16090 -400
rect 16148 -434 16182 -400
rect 16240 -434 16274 -400
rect 16332 -434 16366 -400
rect 16424 -434 16458 -400
rect 16516 -434 16550 -400
rect 16608 -434 16642 -400
rect 16700 -434 16734 -400
rect 16792 -434 16826 -400
rect 16884 -434 16918 -400
rect 16976 -434 17010 -400
rect 17068 -434 17102 -400
rect 17160 -434 17194 -400
rect 17252 -434 17286 -400
rect 17344 -434 17378 -400
rect 17436 -434 17470 -400
rect 17528 -434 17562 -400
rect 17804 -434 17838 -400
rect 17896 -434 17930 -400
rect 17988 -434 18022 -400
rect 18080 -434 18114 -400
rect 18172 -434 18206 -400
rect 18264 -434 18298 -400
rect 18356 -434 18390 -400
rect 18448 -434 18482 -400
rect 18540 -434 18574 -400
rect 18632 -434 18666 -400
rect 18724 -434 18758 -400
rect 18816 -434 18850 -400
rect 18908 -434 18942 -400
rect 19000 -434 19034 -400
rect 19092 -434 19126 -400
rect 19184 -434 19218 -400
rect 19276 -434 19310 -400
rect 19368 -434 19402 -400
rect 19460 -434 19494 -400
rect 19552 -434 19586 -400
rect 19644 -434 19678 -400
rect 19736 -434 19770 -400
rect 19828 -434 19862 -400
rect 19920 -434 19954 -400
rect 20196 -434 20230 -400
rect 20288 -434 20322 -400
rect 20380 -434 20414 -400
rect 20472 -434 20506 -400
rect 20564 -434 20598 -400
rect 20656 -434 20690 -400
rect 20748 -434 20782 -400
rect 20840 -434 20874 -400
rect 20932 -434 20966 -400
rect 21024 -434 21058 -400
rect 21116 -434 21150 -400
rect 21208 -434 21242 -400
rect 21300 -434 21334 -400
rect 21392 -434 21426 -400
rect 21484 -434 21518 -400
rect 21576 -434 21610 -400
rect 21668 -434 21702 -400
rect 21760 -434 21794 -400
rect 21852 -434 21886 -400
rect 21944 -434 21978 -400
rect 22036 -434 22070 -400
rect 22128 -434 22162 -400
rect 22220 -434 22254 -400
rect 22312 -434 22346 -400
rect 22588 -434 22622 -400
rect 22680 -434 22714 -400
rect 22772 -434 22806 -400
rect 22864 -434 22898 -400
rect 22956 -434 22990 -400
rect 23048 -434 23082 -400
rect 23140 -434 23174 -400
rect 23232 -434 23266 -400
rect 23324 -434 23358 -400
rect 23416 -434 23450 -400
rect 23508 -434 23542 -400
rect 23600 -434 23634 -400
rect 23692 -434 23726 -400
rect 23784 -434 23818 -400
rect 23876 -434 23910 -400
rect 23968 -434 24002 -400
rect 24060 -434 24094 -400
rect 24152 -434 24186 -400
rect 24244 -434 24278 -400
rect 24336 -434 24370 -400
rect 24428 -434 24462 -400
rect 24520 -434 24554 -400
rect 24612 -434 24646 -400
rect 24704 -434 24738 -400
rect 24980 -434 25014 -400
rect 25072 -434 25106 -400
rect 25164 -434 25198 -400
rect 25256 -434 25290 -400
rect 8604 -1123 8638 -1089
rect 8696 -1123 8730 -1089
rect 8788 -1123 8822 -1089
rect 8880 -1123 8914 -1089
rect 8969 -1123 9003 -1089
rect 9071 -1123 9105 -1089
rect 9156 -1123 9190 -1089
rect 9248 -1123 9282 -1089
rect 9340 -1123 9374 -1089
rect 9432 -1123 9466 -1089
rect 9524 -1123 9558 -1089
rect 9616 -1123 9650 -1089
rect 9708 -1123 9742 -1089
rect 9800 -1123 9834 -1089
rect 9892 -1123 9926 -1089
rect 9984 -1123 10018 -1089
rect 10076 -1123 10110 -1089
rect 10352 -1123 10386 -1089
rect 10444 -1123 10478 -1089
rect 10536 -1123 10570 -1089
rect 10628 -1123 10662 -1089
rect 10720 -1123 10754 -1089
rect 10812 -1123 10846 -1089
rect 10904 -1123 10938 -1089
rect 10996 -1123 11030 -1089
rect 11088 -1123 11122 -1089
rect 11180 -1123 11214 -1089
rect 11272 -1123 11306 -1089
rect 11366 -1123 11400 -1089
rect 11457 -1123 11491 -1089
rect 11548 -1123 11582 -1089
rect 11640 -1123 11674 -1089
rect 11732 -1123 11766 -1089
rect 11824 -1123 11858 -1089
rect 11916 -1123 11950 -1089
rect 12008 -1123 12042 -1089
rect 12100 -1123 12134 -1089
rect 12192 -1123 12226 -1089
rect 12284 -1123 12318 -1089
rect 12376 -1123 12410 -1089
rect 12468 -1123 12502 -1089
rect 12744 -1123 12778 -1089
rect 12836 -1123 12870 -1089
rect 12928 -1123 12962 -1089
rect 13020 -1123 13054 -1089
rect 13112 -1123 13146 -1089
rect 13204 -1123 13238 -1089
rect 13296 -1123 13330 -1089
rect 13388 -1123 13422 -1089
rect 13480 -1123 13514 -1089
rect 13572 -1123 13606 -1089
rect 13664 -1123 13698 -1089
rect 13754 -1123 13788 -1089
rect 13848 -1123 13882 -1089
rect 13940 -1123 13974 -1089
rect 14032 -1123 14066 -1089
rect 14124 -1123 14158 -1089
rect 14216 -1123 14250 -1089
rect 14308 -1123 14342 -1089
rect 14400 -1123 14434 -1089
rect 14492 -1123 14526 -1089
rect 14584 -1123 14618 -1089
rect 14676 -1123 14710 -1089
rect 14768 -1123 14802 -1089
rect 14860 -1123 14894 -1089
rect 15136 -1123 15170 -1089
rect 15228 -1123 15262 -1089
rect 15320 -1123 15354 -1089
rect 15412 -1123 15446 -1089
rect 15504 -1123 15538 -1089
rect 15596 -1123 15630 -1089
rect 15688 -1123 15722 -1089
rect 15780 -1123 15814 -1089
rect 15872 -1123 15906 -1089
rect 15964 -1123 15998 -1089
rect 16056 -1123 16090 -1089
rect 16149 -1123 16183 -1089
rect 16240 -1123 16274 -1089
rect 16332 -1123 16366 -1089
rect 16424 -1123 16458 -1089
rect 16516 -1123 16550 -1089
rect 16608 -1123 16642 -1089
rect 16700 -1123 16734 -1089
rect 16792 -1123 16826 -1089
rect 16884 -1123 16918 -1089
rect 16976 -1123 17010 -1089
rect 17068 -1123 17102 -1089
rect 17160 -1123 17194 -1089
rect 17252 -1123 17286 -1089
rect 17528 -1123 17562 -1089
rect 17620 -1123 17654 -1089
rect 17712 -1123 17746 -1089
rect 17804 -1123 17838 -1089
rect 17896 -1123 17930 -1089
rect 17988 -1123 18022 -1089
rect 18080 -1123 18114 -1089
rect 18172 -1123 18206 -1089
rect 18264 -1123 18298 -1089
rect 18356 -1123 18390 -1089
rect 18448 -1123 18482 -1089
rect 18538 -1123 18572 -1089
rect 18633 -1123 18667 -1089
rect 18724 -1123 18758 -1089
rect 18816 -1123 18850 -1089
rect 18908 -1123 18942 -1089
rect 19000 -1123 19034 -1089
rect 19092 -1123 19126 -1089
rect 19184 -1123 19218 -1089
rect 19276 -1123 19310 -1089
rect 19368 -1123 19402 -1089
rect 19460 -1123 19494 -1089
rect 19552 -1123 19586 -1089
rect 19644 -1123 19678 -1089
rect 19920 -1123 19954 -1089
rect 20012 -1123 20046 -1089
rect 20104 -1123 20138 -1089
rect 20196 -1123 20230 -1089
rect 20288 -1123 20322 -1089
rect 20380 -1123 20414 -1089
rect 20472 -1123 20506 -1089
rect 20564 -1123 20598 -1089
rect 20656 -1123 20690 -1089
rect 20748 -1123 20782 -1089
rect 20840 -1123 20874 -1089
rect 20932 -1123 20966 -1089
rect 21023 -1123 21057 -1089
rect 21116 -1123 21150 -1089
rect 21208 -1123 21242 -1089
rect 21300 -1123 21334 -1089
rect 21392 -1123 21426 -1089
rect 21484 -1123 21518 -1089
rect 21576 -1123 21610 -1089
rect 21668 -1123 21702 -1089
rect 21760 -1123 21794 -1089
rect 21852 -1123 21886 -1089
rect 21944 -1123 21978 -1089
rect 22036 -1123 22070 -1089
rect 22312 -1123 22346 -1089
rect 22404 -1123 22438 -1089
rect 22496 -1123 22530 -1089
rect 22588 -1123 22622 -1089
rect 22680 -1123 22714 -1089
rect 22772 -1123 22806 -1089
rect 22864 -1123 22898 -1089
rect 22956 -1123 22990 -1089
rect 23048 -1123 23082 -1089
rect 23140 -1123 23174 -1089
rect 23232 -1123 23266 -1089
rect 23323 -1123 23357 -1089
rect 23417 -1123 23451 -1089
rect 23508 -1123 23542 -1089
rect 23600 -1123 23634 -1089
rect 23692 -1123 23726 -1089
rect 23784 -1123 23818 -1089
rect 23876 -1123 23910 -1089
rect 23968 -1123 24002 -1089
rect 24060 -1123 24094 -1089
rect 24152 -1123 24186 -1089
rect 24244 -1123 24278 -1089
rect 24336 -1123 24370 -1089
rect 24428 -1123 24462 -1089
rect 24704 -1123 24738 -1089
rect 24796 -1123 24830 -1089
rect 24888 -1123 24922 -1089
rect 24980 -1123 25014 -1089
rect 25072 -1123 25106 -1089
rect 25164 -1123 25198 -1089
rect 25256 -1123 25290 -1089
<< poly >>
rect 13862 13593 13892 13623
rect 20571 13593 20601 13623
rect 13862 13455 13892 13509
rect 20571 13455 20601 13509
rect 13862 13317 13892 13371
rect 20571 13317 20601 13371
rect 13862 13179 13892 13233
rect 2974 13118 3004 13148
rect 20571 13179 20601 13233
rect 2974 12980 3004 13034
rect 13862 13041 13892 13095
rect 2974 12842 3004 12896
rect 13394 12946 13424 12972
rect 13584 12946 13614 12972
rect 20571 13041 20601 13095
rect 2974 12704 3004 12758
rect 13862 12903 13892 12957
rect 20103 12946 20133 12972
rect 20293 12946 20323 12972
rect 13862 12788 13892 12819
rect 13844 12772 13910 12788
rect 13394 12714 13424 12746
rect 13338 12698 13424 12714
rect 13338 12664 13354 12698
rect 13388 12664 13424 12698
rect 13338 12648 13424 12664
rect 2974 12566 3004 12620
rect 13394 12626 13424 12648
rect 13584 12714 13614 12746
rect 13844 12738 13860 12772
rect 13894 12738 13910 12772
rect 20571 12903 20601 12957
rect 20571 12788 20601 12819
rect 20553 12772 20619 12788
rect 13844 12722 13910 12738
rect 20103 12714 20133 12746
rect 13584 12698 13670 12714
rect 13584 12664 13620 12698
rect 13654 12664 13670 12698
rect 13584 12648 13670 12664
rect 20047 12698 20133 12714
rect 20047 12664 20063 12698
rect 20097 12664 20133 12698
rect 20047 12648 20133 12664
rect 13584 12626 13614 12648
rect 20103 12626 20133 12648
rect 20293 12714 20323 12746
rect 20553 12738 20569 12772
rect 20603 12738 20619 12772
rect 20553 12722 20619 12738
rect 20293 12698 20379 12714
rect 20293 12664 20329 12698
rect 20363 12664 20379 12698
rect 20293 12648 20379 12664
rect 20293 12626 20323 12648
rect 2506 12471 2536 12497
rect 2696 12471 2726 12497
rect 2974 12428 3004 12482
rect 19647 12592 19677 12623
rect 14486 12529 14552 12545
rect 13394 12470 13424 12496
rect 13584 12470 13614 12496
rect 14486 12495 14502 12529
rect 14536 12495 14552 12529
rect 14486 12479 14552 12495
rect 15218 12532 15284 12548
rect 15218 12498 15234 12532
rect 15268 12498 15284 12532
rect 15218 12482 15284 12498
rect 15344 12532 15410 12548
rect 15344 12498 15360 12532
rect 15394 12498 15410 12532
rect 15344 12482 15410 12498
rect 16430 12532 16496 12548
rect 16430 12498 16446 12532
rect 16480 12498 16496 12532
rect 16430 12482 16496 12498
rect 16556 12532 16622 12548
rect 16556 12498 16572 12532
rect 16606 12498 16622 12532
rect 16556 12482 16622 12498
rect 17642 12532 17708 12548
rect 17642 12498 17658 12532
rect 17692 12498 17708 12532
rect 17642 12482 17708 12498
rect 17768 12532 17834 12548
rect 17768 12498 17784 12532
rect 17818 12498 17834 12532
rect 17768 12482 17834 12498
rect 18854 12532 18920 12548
rect 18854 12498 18870 12532
rect 18904 12498 18920 12532
rect 18854 12482 18920 12498
rect 18980 12532 19046 12548
rect 18980 12498 18996 12532
rect 19030 12498 19046 12532
rect 18980 12482 19046 12498
rect 14504 12448 14534 12479
rect 15236 12451 15266 12482
rect 15362 12451 15392 12482
rect 16448 12451 16478 12482
rect 16574 12451 16604 12482
rect 17660 12451 17690 12482
rect 17786 12451 17816 12482
rect 18872 12451 18902 12482
rect 18998 12451 19028 12482
rect 19647 12454 19677 12508
rect 26356 12592 26386 12623
rect 21195 12529 21261 12545
rect 19739 12454 19769 12480
rect 19835 12454 19865 12485
rect 20103 12470 20133 12496
rect 20293 12470 20323 12496
rect 21195 12495 21211 12529
rect 21245 12495 21261 12529
rect 21195 12479 21261 12495
rect 21927 12532 21993 12548
rect 21927 12498 21943 12532
rect 21977 12498 21993 12532
rect 21927 12482 21993 12498
rect 22053 12532 22119 12548
rect 22053 12498 22069 12532
rect 22103 12498 22119 12532
rect 22053 12482 22119 12498
rect 23139 12532 23205 12548
rect 23139 12498 23155 12532
rect 23189 12498 23205 12532
rect 23139 12482 23205 12498
rect 23265 12532 23331 12548
rect 23265 12498 23281 12532
rect 23315 12498 23331 12532
rect 23265 12482 23331 12498
rect 24351 12532 24417 12548
rect 24351 12498 24367 12532
rect 24401 12498 24417 12532
rect 24351 12482 24417 12498
rect 24477 12532 24543 12548
rect 24477 12498 24493 12532
rect 24527 12498 24543 12532
rect 24477 12482 24543 12498
rect 25563 12532 25629 12548
rect 25563 12498 25579 12532
rect 25613 12498 25629 12532
rect 25563 12482 25629 12498
rect 25689 12532 25755 12548
rect 25689 12498 25705 12532
rect 25739 12498 25755 12532
rect 25689 12482 25755 12498
rect 10961 12402 10991 12428
rect 11045 12402 11075 12428
rect 11233 12402 11263 12428
rect 11328 12402 11358 12428
rect 11434 12402 11464 12428
rect 11530 12402 11560 12428
rect 11640 12402 11670 12428
rect 11740 12402 11770 12428
rect 11824 12402 11854 12428
rect 12012 12402 12042 12428
rect 12107 12402 12137 12428
rect 12216 12402 12246 12428
rect 12311 12402 12341 12428
rect 12397 12402 12427 12428
rect 12515 12402 12545 12428
rect 12599 12402 12629 12428
rect 12787 12402 12817 12428
rect 12882 12402 12912 12428
rect 13070 12402 13100 12428
rect 13165 12402 13195 12428
rect 2974 12313 3004 12344
rect 2956 12297 3022 12313
rect 10961 12303 10991 12318
rect 2506 12239 2536 12271
rect 2450 12223 2536 12239
rect 2450 12189 2466 12223
rect 2500 12189 2536 12223
rect 2450 12173 2536 12189
rect 2506 12151 2536 12173
rect 2696 12239 2726 12271
rect 2956 12263 2972 12297
rect 3006 12263 3022 12297
rect 2956 12247 3022 12263
rect 10928 12273 10991 12303
rect 2696 12223 2782 12239
rect 10928 12235 10958 12273
rect 2696 12189 2732 12223
rect 2766 12189 2782 12223
rect 10903 12219 10958 12235
rect 11045 12229 11075 12318
rect 11233 12248 11263 12318
rect 11328 12308 11358 12330
rect 11328 12292 11392 12308
rect 11328 12258 11348 12292
rect 11382 12258 11392 12292
rect 2696 12173 2782 12189
rect 2696 12151 2726 12173
rect 10903 12185 10914 12219
rect 10948 12185 10958 12219
rect 10903 12169 10958 12185
rect 11000 12219 11075 12229
rect 11000 12185 11016 12219
rect 11050 12185 11075 12219
rect 11000 12175 11075 12185
rect 11222 12232 11276 12248
rect 11328 12242 11392 12258
rect 11434 12296 11464 12330
rect 11434 12280 11488 12296
rect 11434 12246 11444 12280
rect 11478 12246 11488 12280
rect 11222 12198 11232 12232
rect 11266 12198 11276 12232
rect 11434 12230 11488 12246
rect 11434 12200 11464 12230
rect 11222 12182 11276 12198
rect 8759 12117 8789 12148
rect 10928 12131 10958 12169
rect 3598 12054 3664 12070
rect 2506 11995 2536 12021
rect 2696 11995 2726 12021
rect 3598 12020 3614 12054
rect 3648 12020 3664 12054
rect 3598 12004 3664 12020
rect 4330 12057 4396 12073
rect 4330 12023 4346 12057
rect 4380 12023 4396 12057
rect 4330 12007 4396 12023
rect 4456 12057 4522 12073
rect 4456 12023 4472 12057
rect 4506 12023 4522 12057
rect 4456 12007 4522 12023
rect 5542 12057 5608 12073
rect 5542 12023 5558 12057
rect 5592 12023 5608 12057
rect 5542 12007 5608 12023
rect 5668 12057 5734 12073
rect 5668 12023 5684 12057
rect 5718 12023 5734 12057
rect 5668 12007 5734 12023
rect 6754 12057 6820 12073
rect 6754 12023 6770 12057
rect 6804 12023 6820 12057
rect 6754 12007 6820 12023
rect 6880 12057 6946 12073
rect 6880 12023 6896 12057
rect 6930 12023 6946 12057
rect 6880 12007 6946 12023
rect 7966 12057 8032 12073
rect 7966 12023 7982 12057
rect 8016 12023 8032 12057
rect 7966 12007 8032 12023
rect 8092 12057 8158 12073
rect 8092 12023 8108 12057
rect 8142 12023 8158 12057
rect 9181 12094 9211 12120
rect 10928 12101 10991 12131
rect 8092 12007 8158 12023
rect 3616 11973 3646 12004
rect 4348 11976 4378 12007
rect 4474 11976 4504 12007
rect 5560 11976 5590 12007
rect 5686 11976 5716 12007
rect 6772 11976 6802 12007
rect 6898 11976 6928 12007
rect 7984 11976 8014 12007
rect 8110 11976 8140 12007
rect 8759 11979 8789 12033
rect 8851 11979 8881 12005
rect 8947 11979 8977 12010
rect 3616 11861 3646 11889
rect 4348 11864 4378 11892
rect 4474 11864 4504 11892
rect 5560 11864 5590 11892
rect 5686 11864 5716 11892
rect 6772 11864 6802 11892
rect 6898 11864 6928 11892
rect 7984 11864 8014 11892
rect 8110 11864 8140 11892
rect 8759 11870 8789 11895
rect 8630 11850 8789 11870
rect 8851 11870 8881 11895
rect 8947 11870 8977 11895
rect 10961 12086 10991 12101
rect 11045 12086 11075 12175
rect 11233 12036 11263 12182
rect 11326 12170 11464 12200
rect 11326 12036 11356 12170
rect 11530 12134 11560 12318
rect 11640 12286 11670 12318
rect 11606 12270 11670 12286
rect 12107 12308 12137 12330
rect 12107 12292 12174 12308
rect 11606 12236 11616 12270
rect 11650 12256 11670 12270
rect 11650 12236 11666 12256
rect 11606 12220 11666 12236
rect 11398 12118 11464 12128
rect 11398 12084 11414 12118
rect 11448 12084 11464 12118
rect 11398 12074 11464 12084
rect 11530 12118 11594 12134
rect 11530 12084 11550 12118
rect 11584 12084 11594 12118
rect 11410 12036 11440 12074
rect 11530 12068 11594 12084
rect 11530 12036 11560 12068
rect 11636 12036 11666 12220
rect 11740 12218 11770 12274
rect 11824 12218 11854 12274
rect 12012 12252 12042 12274
rect 11988 12236 12042 12252
rect 12107 12258 12130 12292
rect 12164 12258 12174 12292
rect 12107 12242 12174 12258
rect 11708 12202 11774 12218
rect 11708 12168 11718 12202
rect 11752 12168 11774 12202
rect 11708 12152 11774 12168
rect 11824 12202 11914 12218
rect 11988 12216 11998 12236
rect 11824 12168 11870 12202
rect 11904 12168 11914 12202
rect 11824 12152 11914 12168
rect 11965 12202 11998 12216
rect 12032 12202 12042 12236
rect 11965 12186 12042 12202
rect 12216 12200 12246 12330
rect 11744 12120 11774 12152
rect 11828 12120 11858 12152
rect 11965 12120 11995 12186
rect 12109 12170 12246 12200
rect 12109 12134 12139 12170
rect 10961 11932 10991 11958
rect 11045 11932 11075 11958
rect 12085 12118 12139 12134
rect 12311 12134 12341 12318
rect 12397 12286 12427 12318
rect 12383 12270 12449 12286
rect 12383 12236 12393 12270
rect 12427 12236 12449 12270
rect 12383 12220 12449 12236
rect 12515 12234 12545 12274
rect 12085 12084 12095 12118
rect 12129 12084 12139 12118
rect 12085 12068 12139 12084
rect 12181 12118 12247 12128
rect 12181 12084 12197 12118
rect 12231 12084 12247 12118
rect 12181 12074 12247 12084
rect 12311 12118 12377 12134
rect 12311 12084 12333 12118
rect 12367 12084 12377 12118
rect 12109 12036 12139 12068
rect 12193 12036 12223 12074
rect 12311 12068 12377 12084
rect 12311 12036 12341 12068
rect 12419 12036 12449 12220
rect 12491 12218 12545 12234
rect 12491 12184 12501 12218
rect 12535 12184 12545 12218
rect 12491 12168 12545 12184
rect 12599 12218 12629 12274
rect 12787 12246 12817 12318
rect 13070 12303 13100 12318
rect 13044 12273 13100 12303
rect 12882 12250 12912 12272
rect 12754 12230 12818 12246
rect 12599 12202 12683 12218
rect 12599 12182 12639 12202
rect 12515 12120 12545 12168
rect 12587 12168 12639 12182
rect 12673 12168 12683 12202
rect 12754 12196 12770 12230
rect 12804 12196 12818 12230
rect 12754 12180 12818 12196
rect 12860 12244 12912 12250
rect 13044 12244 13074 12273
rect 21213 12448 21243 12479
rect 21945 12451 21975 12482
rect 22071 12451 22101 12482
rect 23157 12451 23187 12482
rect 23283 12451 23313 12482
rect 24369 12451 24399 12482
rect 24495 12451 24525 12482
rect 25581 12451 25611 12482
rect 25707 12451 25737 12482
rect 26356 12454 26386 12508
rect 26448 12454 26478 12480
rect 26544 12454 26574 12485
rect 14504 12336 14534 12364
rect 15236 12339 15266 12367
rect 15362 12339 15392 12367
rect 16448 12339 16478 12367
rect 16574 12339 16604 12367
rect 17660 12339 17690 12367
rect 17786 12339 17816 12367
rect 18872 12339 18902 12367
rect 18998 12339 19028 12367
rect 19647 12345 19677 12370
rect 19518 12325 19677 12345
rect 19739 12345 19769 12370
rect 19835 12345 19865 12370
rect 19739 12339 19865 12345
rect 19518 12291 19530 12325
rect 19564 12291 19677 12325
rect 13165 12250 13195 12272
rect 14857 12250 14887 12276
rect 15589 12250 15619 12276
rect 15711 12250 15741 12276
rect 16801 12250 16831 12276
rect 16923 12250 16953 12276
rect 18139 12250 18169 12276
rect 18261 12250 18291 12276
rect 18995 12250 19025 12276
rect 19518 12272 19677 12291
rect 19721 12323 19865 12339
rect 21213 12336 21243 12364
rect 21945 12339 21975 12367
rect 22071 12339 22101 12367
rect 23157 12339 23187 12367
rect 23283 12339 23313 12367
rect 24369 12339 24399 12367
rect 24495 12339 24525 12367
rect 25581 12339 25611 12367
rect 25707 12339 25737 12367
rect 26356 12345 26386 12370
rect 19721 12289 19737 12323
rect 19771 12289 19865 12323
rect 19721 12273 19865 12289
rect 26227 12325 26386 12345
rect 26448 12345 26478 12370
rect 26544 12345 26574 12370
rect 26448 12339 26574 12345
rect 26227 12291 26239 12325
rect 26273 12291 26386 12325
rect 19647 12251 19677 12272
rect 19739 12266 19865 12273
rect 19739 12251 19769 12266
rect 19835 12251 19865 12266
rect 12860 12234 13074 12244
rect 12860 12200 12870 12234
rect 12904 12200 13074 12234
rect 12860 12190 13074 12200
rect 12860 12184 12912 12190
rect 12587 12152 12683 12168
rect 12587 12120 12617 12152
rect 12785 12148 12815 12180
rect 12882 12152 12912 12184
rect 12785 11994 12815 12020
rect 13044 12142 13074 12190
rect 13136 12234 13195 12250
rect 13136 12200 13146 12234
rect 13180 12200 13195 12234
rect 13136 12184 13195 12200
rect 13165 12152 13195 12184
rect 21566 12250 21596 12276
rect 22298 12250 22328 12276
rect 22420 12250 22450 12276
rect 23510 12250 23540 12276
rect 23632 12250 23662 12276
rect 24848 12250 24878 12276
rect 24970 12250 25000 12276
rect 25704 12250 25734 12276
rect 26227 12272 26386 12291
rect 26430 12323 26574 12339
rect 26430 12289 26446 12323
rect 26480 12289 26574 12323
rect 26430 12273 26574 12289
rect 26356 12251 26386 12272
rect 26448 12266 26574 12273
rect 26448 12251 26478 12266
rect 26544 12251 26574 12266
rect 13044 12112 13100 12142
rect 13070 12096 13100 12112
rect 11233 11926 11263 11952
rect 11326 11926 11356 11952
rect 11410 11926 11440 11952
rect 11530 11926 11560 11952
rect 11636 11926 11666 11952
rect 11744 11926 11774 11952
rect 11828 11926 11858 11952
rect 11965 11926 11995 11952
rect 12109 11926 12139 11952
rect 12193 11926 12223 11952
rect 12311 11926 12341 11952
rect 12419 11926 12449 11952
rect 12515 11926 12545 11952
rect 12587 11926 12617 11952
rect 12882 11926 12912 11952
rect 13070 11942 13100 11968
rect 13855 12138 13921 12154
rect 14857 12144 14887 12166
rect 15589 12144 15619 12166
rect 15711 12144 15741 12166
rect 16801 12144 16831 12166
rect 16923 12144 16953 12166
rect 18139 12144 18169 12166
rect 18261 12144 18291 12166
rect 18995 12144 19025 12166
rect 13855 12111 13871 12138
rect 13837 12104 13871 12111
rect 13905 12111 13921 12138
rect 14839 12128 14905 12144
rect 13905 12104 13939 12111
rect 13837 12081 13939 12104
rect 13837 12066 13867 12081
rect 13909 12066 13939 12081
rect 14839 12094 14855 12128
rect 14889 12094 14905 12128
rect 14839 12078 14905 12094
rect 15571 12128 15637 12144
rect 15571 12094 15587 12128
rect 15621 12094 15637 12128
rect 15571 12078 15637 12094
rect 15693 12128 15759 12144
rect 15693 12094 15709 12128
rect 15743 12094 15759 12128
rect 15693 12078 15759 12094
rect 16783 12128 16849 12144
rect 16783 12094 16799 12128
rect 16833 12094 16849 12128
rect 16783 12078 16849 12094
rect 16905 12128 16971 12144
rect 16905 12094 16921 12128
rect 16955 12094 16971 12128
rect 16905 12078 16971 12094
rect 18121 12128 18187 12144
rect 18121 12094 18137 12128
rect 18171 12094 18187 12128
rect 18121 12078 18187 12094
rect 18243 12128 18309 12144
rect 18243 12094 18259 12128
rect 18293 12094 18309 12128
rect 18243 12078 18309 12094
rect 18977 12128 19043 12144
rect 18977 12094 18993 12128
rect 19027 12094 19043 12128
rect 19647 12113 19677 12167
rect 19739 12141 19769 12167
rect 19835 12141 19865 12167
rect 20564 12138 20630 12154
rect 21566 12144 21596 12166
rect 22298 12144 22328 12166
rect 22420 12144 22450 12166
rect 23510 12144 23540 12166
rect 23632 12144 23662 12166
rect 24848 12144 24878 12166
rect 24970 12144 25000 12166
rect 25704 12144 25734 12166
rect 18977 12078 19043 12094
rect 20564 12111 20580 12138
rect 20546 12104 20580 12111
rect 20614 12111 20630 12138
rect 21548 12128 21614 12144
rect 20614 12104 20648 12111
rect 20546 12081 20648 12104
rect 20546 12066 20576 12081
rect 20618 12066 20648 12081
rect 21548 12094 21564 12128
rect 21598 12094 21614 12128
rect 21548 12078 21614 12094
rect 22280 12128 22346 12144
rect 22280 12094 22296 12128
rect 22330 12094 22346 12128
rect 22280 12078 22346 12094
rect 22402 12128 22468 12144
rect 22402 12094 22418 12128
rect 22452 12094 22468 12128
rect 22402 12078 22468 12094
rect 23492 12128 23558 12144
rect 23492 12094 23508 12128
rect 23542 12094 23558 12128
rect 23492 12078 23558 12094
rect 23614 12128 23680 12144
rect 23614 12094 23630 12128
rect 23664 12094 23680 12128
rect 23614 12078 23680 12094
rect 24830 12128 24896 12144
rect 24830 12094 24846 12128
rect 24880 12094 24896 12128
rect 24830 12078 24896 12094
rect 24952 12128 25018 12144
rect 24952 12094 24968 12128
rect 25002 12094 25018 12128
rect 24952 12078 25018 12094
rect 25686 12128 25752 12144
rect 25686 12094 25702 12128
rect 25736 12094 25752 12128
rect 26356 12113 26386 12167
rect 26448 12141 26478 12167
rect 26544 12141 26574 12167
rect 25686 12078 25752 12094
rect 19647 12002 19677 12029
rect 26356 12002 26386 12029
rect 13165 11926 13195 11952
rect 13837 11928 13867 11982
rect 13909 11928 13939 11982
rect 20546 11928 20576 11982
rect 20618 11928 20648 11982
rect 8851 11864 8977 11870
rect 8630 11816 8642 11850
rect 8676 11816 8789 11850
rect 3969 11775 3999 11801
rect 4701 11775 4731 11801
rect 4823 11775 4853 11801
rect 5913 11775 5943 11801
rect 6035 11775 6065 11801
rect 7251 11775 7281 11801
rect 7373 11775 7403 11801
rect 8107 11775 8137 11801
rect 8630 11797 8789 11816
rect 8833 11848 8977 11864
rect 9181 11862 9211 11894
rect 8833 11814 8849 11848
rect 8883 11814 8977 11848
rect 8833 11798 8977 11814
rect 8759 11776 8789 11797
rect 8851 11791 8977 11798
rect 9125 11846 9211 11862
rect 9125 11812 9141 11846
rect 9175 11812 9211 11846
rect 9125 11796 9211 11812
rect 8851 11776 8881 11791
rect 8947 11776 8977 11791
rect 9181 11774 9211 11796
rect 13837 11790 13867 11844
rect 13909 11790 13939 11844
rect 20546 11790 20576 11844
rect 20618 11790 20648 11844
rect 2967 11663 3033 11679
rect 3969 11669 3999 11691
rect 4701 11669 4731 11691
rect 4823 11669 4853 11691
rect 5913 11669 5943 11691
rect 6035 11669 6065 11691
rect 7251 11669 7281 11691
rect 7373 11669 7403 11691
rect 8107 11669 8137 11691
rect 2967 11636 2983 11663
rect 2949 11629 2983 11636
rect 3017 11636 3033 11663
rect 3951 11653 4017 11669
rect 3017 11629 3051 11636
rect 2949 11606 3051 11629
rect 2949 11591 2979 11606
rect 3021 11591 3051 11606
rect 3951 11619 3967 11653
rect 4001 11619 4017 11653
rect 3951 11603 4017 11619
rect 4683 11653 4749 11669
rect 4683 11619 4699 11653
rect 4733 11619 4749 11653
rect 4683 11603 4749 11619
rect 4805 11653 4871 11669
rect 4805 11619 4821 11653
rect 4855 11619 4871 11653
rect 4805 11603 4871 11619
rect 5895 11653 5961 11669
rect 5895 11619 5911 11653
rect 5945 11619 5961 11653
rect 5895 11603 5961 11619
rect 6017 11653 6083 11669
rect 6017 11619 6033 11653
rect 6067 11619 6083 11653
rect 6017 11603 6083 11619
rect 7233 11653 7299 11669
rect 7233 11619 7249 11653
rect 7283 11619 7299 11653
rect 7233 11603 7299 11619
rect 7355 11653 7421 11669
rect 7355 11619 7371 11653
rect 7405 11619 7421 11653
rect 7355 11603 7421 11619
rect 8089 11653 8155 11669
rect 8089 11619 8105 11653
rect 8139 11619 8155 11653
rect 8759 11638 8789 11692
rect 8851 11666 8881 11692
rect 8947 11666 8977 11692
rect 11002 11762 11032 11788
rect 11278 11762 11308 11788
rect 8089 11603 8155 11619
rect 9181 11618 9211 11644
rect 8759 11527 8789 11554
rect 13837 11652 13867 11706
rect 13909 11652 13939 11706
rect 20546 11652 20576 11706
rect 20618 11652 20648 11706
rect 11002 11530 11032 11562
rect 11278 11530 11308 11562
rect 10946 11514 11032 11530
rect 2949 11453 2979 11507
rect 3021 11453 3051 11507
rect 10946 11480 10962 11514
rect 10996 11480 11032 11514
rect 10946 11464 11032 11480
rect 11222 11514 11308 11530
rect 13837 11514 13867 11568
rect 13909 11514 13939 11568
rect 20546 11514 20576 11568
rect 20618 11514 20648 11568
rect 11222 11480 11238 11514
rect 11272 11480 11308 11514
rect 11222 11464 11308 11480
rect 11002 11442 11032 11464
rect 11278 11442 11308 11464
rect 2949 11315 2979 11369
rect 3021 11315 3051 11369
rect 13837 11376 13867 11430
rect 13909 11376 13939 11430
rect 20546 11376 20576 11430
rect 20618 11376 20648 11430
rect 11002 11286 11032 11312
rect 11278 11286 11308 11312
rect 2949 11177 2979 11231
rect 3021 11177 3051 11231
rect 13837 11238 13867 11292
rect 13909 11238 13939 11292
rect 20546 11238 20576 11292
rect 20618 11238 20648 11292
rect 13837 11100 13867 11154
rect 13909 11100 13939 11154
rect 20546 11100 20576 11154
rect 20618 11100 20648 11154
rect 2949 11039 2979 11093
rect 3021 11039 3051 11093
rect 13837 10990 13867 11016
rect 13909 10990 13939 11016
rect 20546 10990 20576 11016
rect 20618 10990 20648 11016
rect 2949 10901 2979 10955
rect 3021 10901 3051 10955
rect 2949 10763 2979 10817
rect 3021 10763 3051 10817
rect 2949 10625 2979 10679
rect 3021 10625 3051 10679
rect 2949 10515 2979 10541
rect 3021 10515 3051 10541
rect 2949 10105 2979 10131
rect 3021 10105 3051 10131
rect 19240 10093 19270 10119
rect 19312 10093 19342 10119
rect 2949 9967 2979 10021
rect 3021 9967 3051 10021
rect 25949 10093 25979 10119
rect 26021 10093 26051 10119
rect 2949 9829 2979 9883
rect 3021 9829 3051 9883
rect 19240 9955 19270 10009
rect 19312 9955 19342 10009
rect 25949 9955 25979 10009
rect 26021 9955 26051 10009
rect 19240 9817 19270 9871
rect 19312 9817 19342 9871
rect 25949 9817 25979 9871
rect 26021 9817 26051 9871
rect 2949 9691 2979 9745
rect 3021 9691 3051 9745
rect 19240 9679 19270 9733
rect 19312 9679 19342 9733
rect 25949 9679 25979 9733
rect 26021 9679 26051 9733
rect 2949 9553 2979 9607
rect 3021 9553 3051 9607
rect 19240 9541 19270 9595
rect 19312 9541 19342 9595
rect 25949 9541 25979 9595
rect 26021 9541 26051 9595
rect 2949 9415 2979 9469
rect 3021 9415 3051 9469
rect 19240 9403 19270 9457
rect 19312 9403 19342 9457
rect 25949 9403 25979 9457
rect 26021 9403 26051 9457
rect 2949 9277 2979 9331
rect 3021 9277 3051 9331
rect 19240 9265 19270 9319
rect 19312 9265 19342 9319
rect 25949 9265 25979 9319
rect 26021 9265 26051 9319
rect 2949 9139 2979 9193
rect 3021 9139 3051 9193
rect 19240 9127 19270 9181
rect 19312 9127 19342 9181
rect 25949 9127 25979 9181
rect 26021 9127 26051 9181
rect 8759 9092 8789 9119
rect 2949 9040 2979 9055
rect 3021 9040 3051 9055
rect 2949 9017 3051 9040
rect 2949 9010 2983 9017
rect 2967 8983 2983 9010
rect 3017 9010 3051 9017
rect 3951 9027 4017 9043
rect 3017 8983 3033 9010
rect 2967 8967 3033 8983
rect 3951 8993 3967 9027
rect 4001 8993 4017 9027
rect 3951 8977 4017 8993
rect 4683 9027 4749 9043
rect 4683 8993 4699 9027
rect 4733 8993 4749 9027
rect 4683 8977 4749 8993
rect 4805 9027 4871 9043
rect 4805 8993 4821 9027
rect 4855 8993 4871 9027
rect 4805 8977 4871 8993
rect 5895 9027 5961 9043
rect 5895 8993 5911 9027
rect 5945 8993 5961 9027
rect 5895 8977 5961 8993
rect 6017 9027 6083 9043
rect 6017 8993 6033 9027
rect 6067 8993 6083 9027
rect 6017 8977 6083 8993
rect 7233 9027 7299 9043
rect 7233 8993 7249 9027
rect 7283 8993 7299 9027
rect 7233 8977 7299 8993
rect 7355 9027 7421 9043
rect 7355 8993 7371 9027
rect 7405 8993 7421 9027
rect 7355 8977 7421 8993
rect 8089 9027 8155 9043
rect 8089 8993 8105 9027
rect 8139 8993 8155 9027
rect 13502 9080 13532 9107
rect 8089 8977 8155 8993
rect 3969 8955 3999 8977
rect 4701 8955 4731 8977
rect 4823 8955 4853 8977
rect 5913 8955 5943 8977
rect 6035 8955 6065 8977
rect 7251 8955 7281 8977
rect 7373 8955 7403 8977
rect 8107 8955 8137 8977
rect 8759 8954 8789 9008
rect 9181 9004 9211 9030
rect 9396 9004 9426 9030
rect 9491 9004 9521 9030
rect 9679 9004 9709 9030
rect 9774 9004 9804 9030
rect 9962 9004 9992 9030
rect 10046 9004 10076 9030
rect 10164 9004 10194 9030
rect 10250 9004 10280 9030
rect 10345 9004 10375 9030
rect 10454 9004 10484 9030
rect 10549 9004 10579 9030
rect 10737 9004 10767 9030
rect 10821 9004 10851 9030
rect 10921 9004 10951 9030
rect 11031 9004 11061 9030
rect 11127 9004 11157 9030
rect 11233 9004 11263 9030
rect 11328 9004 11358 9030
rect 11516 9004 11546 9030
rect 11600 9004 11630 9030
rect 8851 8954 8881 8980
rect 8947 8954 8977 8980
rect 3969 8845 3999 8871
rect 4701 8845 4731 8871
rect 4823 8845 4853 8871
rect 5913 8845 5943 8871
rect 6035 8845 6065 8871
rect 7251 8845 7281 8871
rect 7373 8845 7403 8871
rect 8107 8845 8137 8871
rect 9491 8905 9521 8920
rect 9491 8875 9547 8905
rect 8759 8849 8789 8870
rect 8630 8830 8789 8849
rect 8851 8855 8881 8870
rect 8947 8855 8977 8870
rect 8851 8848 8977 8855
rect 9181 8852 9211 8874
rect 8630 8796 8642 8830
rect 8676 8796 8789 8830
rect 3616 8757 3646 8785
rect 4348 8754 4378 8782
rect 4474 8754 4504 8782
rect 5560 8754 5590 8782
rect 5686 8754 5716 8782
rect 6772 8754 6802 8782
rect 6898 8754 6928 8782
rect 7984 8754 8014 8782
rect 8110 8754 8140 8782
rect 8630 8776 8789 8796
rect 8833 8832 8977 8848
rect 8833 8798 8849 8832
rect 8883 8798 8977 8832
rect 8833 8782 8977 8798
rect 9125 8836 9211 8852
rect 9125 8802 9141 8836
rect 9175 8802 9211 8836
rect 9125 8786 9211 8802
rect 2506 8625 2536 8651
rect 2696 8625 2726 8651
rect 3616 8642 3646 8673
rect 8759 8751 8789 8776
rect 8851 8776 8977 8782
rect 8851 8751 8881 8776
rect 8947 8751 8977 8776
rect 9181 8754 9211 8786
rect 9396 8852 9426 8874
rect 9396 8836 9455 8852
rect 9396 8802 9411 8836
rect 9445 8802 9455 8836
rect 9396 8786 9455 8802
rect 9517 8846 9547 8875
rect 9679 8852 9709 8874
rect 9679 8846 9731 8852
rect 9774 8848 9804 8920
rect 10164 8888 10194 8920
rect 9517 8836 9731 8846
rect 9517 8802 9687 8836
rect 9721 8802 9731 8836
rect 9517 8792 9731 8802
rect 9396 8754 9426 8786
rect 3598 8626 3664 8642
rect 4348 8639 4378 8670
rect 4474 8639 4504 8670
rect 5560 8639 5590 8670
rect 5686 8639 5716 8670
rect 6772 8639 6802 8670
rect 6898 8639 6928 8670
rect 7984 8639 8014 8670
rect 8110 8639 8140 8670
rect 3598 8592 3614 8626
rect 3648 8592 3664 8626
rect 3598 8576 3664 8592
rect 4330 8623 4396 8639
rect 4330 8589 4346 8623
rect 4380 8589 4396 8623
rect 4330 8573 4396 8589
rect 4456 8623 4522 8639
rect 4456 8589 4472 8623
rect 4506 8589 4522 8623
rect 4456 8573 4522 8589
rect 5542 8623 5608 8639
rect 5542 8589 5558 8623
rect 5592 8589 5608 8623
rect 5542 8573 5608 8589
rect 5668 8623 5734 8639
rect 5668 8589 5684 8623
rect 5718 8589 5734 8623
rect 5668 8573 5734 8589
rect 6754 8623 6820 8639
rect 6754 8589 6770 8623
rect 6804 8589 6820 8623
rect 6754 8573 6820 8589
rect 6880 8623 6946 8639
rect 6880 8589 6896 8623
rect 6930 8589 6946 8623
rect 6880 8573 6946 8589
rect 7966 8623 8032 8639
rect 7966 8589 7982 8623
rect 8016 8589 8032 8623
rect 7966 8573 8032 8589
rect 8092 8623 8158 8639
rect 8092 8589 8108 8623
rect 8142 8589 8158 8623
rect 8759 8613 8789 8667
rect 8851 8641 8881 8667
rect 8947 8636 8977 8667
rect 8092 8573 8158 8589
rect 9517 8744 9547 8792
rect 9679 8786 9731 8792
rect 9773 8832 9837 8848
rect 9773 8798 9787 8832
rect 9821 8798 9837 8832
rect 9962 8820 9992 8876
rect 9679 8754 9709 8786
rect 9773 8782 9837 8798
rect 9908 8804 9992 8820
rect 9491 8714 9547 8744
rect 9491 8698 9521 8714
rect 8759 8498 8789 8529
rect 9181 8528 9211 8554
rect 9396 8528 9426 8554
rect 9491 8544 9521 8570
rect 9776 8750 9806 8782
rect 9908 8770 9918 8804
rect 9952 8784 9992 8804
rect 10046 8836 10076 8876
rect 10142 8872 10208 8888
rect 10142 8838 10164 8872
rect 10198 8838 10208 8872
rect 10046 8820 10100 8836
rect 10046 8786 10056 8820
rect 10090 8786 10100 8820
rect 9952 8770 10004 8784
rect 9908 8754 10004 8770
rect 9974 8722 10004 8754
rect 10046 8770 10100 8786
rect 10142 8822 10208 8838
rect 10046 8722 10076 8770
rect 9776 8596 9806 8622
rect 10142 8638 10172 8822
rect 10250 8736 10280 8920
rect 10345 8802 10375 8932
rect 10454 8910 10484 8932
rect 10417 8894 10484 8910
rect 10417 8860 10427 8894
rect 10461 8860 10484 8894
rect 10921 8888 10951 8920
rect 10417 8844 10484 8860
rect 10549 8854 10579 8876
rect 10549 8838 10603 8854
rect 10549 8804 10559 8838
rect 10593 8818 10603 8838
rect 10737 8820 10767 8876
rect 10821 8820 10851 8876
rect 10921 8872 10985 8888
rect 10921 8858 10941 8872
rect 10925 8838 10941 8858
rect 10975 8838 10985 8872
rect 10925 8822 10985 8838
rect 10593 8804 10626 8818
rect 10345 8772 10482 8802
rect 10549 8788 10626 8804
rect 10214 8720 10280 8736
rect 10452 8736 10482 8772
rect 10214 8686 10224 8720
rect 10258 8686 10280 8720
rect 10214 8670 10280 8686
rect 10344 8720 10410 8730
rect 10344 8686 10360 8720
rect 10394 8686 10410 8720
rect 10344 8676 10410 8686
rect 10452 8720 10506 8736
rect 10596 8722 10626 8788
rect 10677 8804 10767 8820
rect 10677 8770 10687 8804
rect 10721 8770 10767 8804
rect 10677 8754 10767 8770
rect 10817 8804 10883 8820
rect 10817 8770 10839 8804
rect 10873 8770 10883 8804
rect 10817 8754 10883 8770
rect 10733 8722 10763 8754
rect 10817 8722 10847 8754
rect 10452 8686 10462 8720
rect 10496 8686 10506 8720
rect 10250 8638 10280 8670
rect 10368 8638 10398 8676
rect 10452 8670 10506 8686
rect 10452 8638 10482 8670
rect 10925 8638 10955 8822
rect 11031 8736 11061 8920
rect 11127 8898 11157 8932
rect 11233 8910 11263 8932
rect 12728 8991 12758 9017
rect 12812 8991 12842 9017
rect 13051 8991 13081 9017
rect 20211 9080 20241 9107
rect 14136 9015 14202 9031
rect 11883 8956 11913 8982
rect 11979 8956 12009 8982
rect 12075 8956 12105 8982
rect 11103 8882 11157 8898
rect 11103 8848 11113 8882
rect 11147 8848 11157 8882
rect 11103 8832 11157 8848
rect 11199 8894 11263 8910
rect 11199 8860 11209 8894
rect 11243 8860 11263 8894
rect 11199 8844 11263 8860
rect 11328 8850 11358 8920
rect 11127 8802 11157 8832
rect 11315 8834 11369 8850
rect 11127 8772 11265 8802
rect 11315 8800 11325 8834
rect 11359 8800 11369 8834
rect 11315 8784 11369 8800
rect 11516 8831 11546 8920
rect 11600 8905 11630 8920
rect 11600 8875 11663 8905
rect 11633 8837 11663 8875
rect 12279 8944 12309 8970
rect 11883 8857 11913 8872
rect 11979 8857 12009 8872
rect 12075 8857 12105 8872
rect 12480 8943 12510 8969
rect 11883 8850 12105 8857
rect 11516 8821 11591 8831
rect 11516 8787 11541 8821
rect 11575 8787 11591 8821
rect 10997 8720 11061 8736
rect 10997 8686 11007 8720
rect 11041 8686 11061 8720
rect 10997 8670 11061 8686
rect 11127 8720 11193 8730
rect 11127 8686 11143 8720
rect 11177 8686 11193 8720
rect 11127 8676 11193 8686
rect 11031 8638 11061 8670
rect 11151 8638 11181 8676
rect 11235 8638 11265 8772
rect 11328 8638 11358 8784
rect 11516 8777 11591 8787
rect 11633 8821 11688 8837
rect 11883 8827 12123 8850
rect 12279 8838 12309 8860
rect 13314 8942 13344 8968
rect 13410 8942 13440 8968
rect 13502 8942 13532 8996
rect 14136 8981 14152 9015
rect 14186 8981 14202 9015
rect 14136 8965 14202 8981
rect 14870 9015 14936 9031
rect 14870 8981 14886 9015
rect 14920 8981 14936 9015
rect 14870 8965 14936 8981
rect 14992 9015 15058 9031
rect 14992 8981 15008 9015
rect 15042 8981 15058 9015
rect 14992 8965 15058 8981
rect 16208 9015 16274 9031
rect 16208 8981 16224 9015
rect 16258 8981 16274 9015
rect 16208 8965 16274 8981
rect 16330 9015 16396 9031
rect 16330 8981 16346 9015
rect 16380 8981 16396 9015
rect 16330 8965 16396 8981
rect 17420 9015 17486 9031
rect 17420 8981 17436 9015
rect 17470 8981 17486 9015
rect 17420 8965 17486 8981
rect 17542 9015 17608 9031
rect 17542 8981 17558 9015
rect 17592 8981 17608 9015
rect 17542 8965 17608 8981
rect 18274 9015 18340 9031
rect 18274 8981 18290 9015
rect 18324 8981 18340 9015
rect 19240 9028 19270 9043
rect 19312 9028 19342 9043
rect 19240 9005 19342 9028
rect 19240 8998 19274 9005
rect 18274 8965 18340 8981
rect 19258 8971 19274 8998
rect 19308 8998 19342 9005
rect 19308 8971 19324 8998
rect 20845 9015 20911 9031
rect 14154 8943 14184 8965
rect 14888 8943 14918 8965
rect 15010 8943 15040 8965
rect 16226 8943 16256 8965
rect 16348 8943 16378 8965
rect 17438 8943 17468 8965
rect 17560 8943 17590 8965
rect 18292 8943 18322 8965
rect 19258 8955 19324 8971
rect 11633 8787 11643 8821
rect 11677 8787 11688 8821
rect 11516 8688 11546 8777
rect 11633 8771 11688 8787
rect 12057 8821 12123 8827
rect 12057 8787 12073 8821
rect 12107 8787 12123 8821
rect 12057 8785 12123 8787
rect 11883 8771 12123 8785
rect 12261 8822 12327 8838
rect 12480 8837 12510 8859
rect 12728 8839 12758 8861
rect 12261 8788 12277 8822
rect 12311 8788 12327 8822
rect 12261 8772 12327 8788
rect 12462 8821 12528 8837
rect 12462 8787 12478 8821
rect 12512 8787 12528 8821
rect 11633 8733 11663 8771
rect 11883 8755 12105 8771
rect 11883 8740 11913 8755
rect 11979 8740 12009 8755
rect 12075 8740 12105 8755
rect 12279 8741 12309 8772
rect 12462 8771 12528 8787
rect 12670 8823 12758 8839
rect 12670 8789 12687 8823
rect 12721 8789 12758 8823
rect 12670 8773 12758 8789
rect 11600 8703 11663 8733
rect 11600 8688 11630 8703
rect 9679 8528 9709 8554
rect 9974 8528 10004 8554
rect 10046 8528 10076 8554
rect 10142 8528 10172 8554
rect 10250 8528 10280 8554
rect 10368 8528 10398 8554
rect 10452 8528 10482 8554
rect 10596 8528 10626 8554
rect 10733 8528 10763 8554
rect 10817 8528 10847 8554
rect 10925 8528 10955 8554
rect 11031 8528 11061 8554
rect 11151 8528 11181 8554
rect 11235 8528 11265 8554
rect 11328 8528 11358 8554
rect 11516 8534 11546 8560
rect 11600 8534 11630 8560
rect 11316 8507 11388 8528
rect 2506 8473 2536 8495
rect 2450 8457 2536 8473
rect 2450 8423 2466 8457
rect 2500 8423 2536 8457
rect 2450 8407 2536 8423
rect 2506 8375 2536 8407
rect 2696 8473 2726 8495
rect 11316 8473 11332 8507
rect 11366 8473 11388 8507
rect 12480 8740 12510 8771
rect 12728 8741 12758 8773
rect 12812 8839 12842 8861
rect 13051 8839 13081 8861
rect 20023 8942 20053 8968
rect 20119 8942 20149 8968
rect 20211 8942 20241 8996
rect 20845 8981 20861 9015
rect 20895 8981 20911 9015
rect 20845 8965 20911 8981
rect 21579 9015 21645 9031
rect 21579 8981 21595 9015
rect 21629 8981 21645 9015
rect 21579 8965 21645 8981
rect 21701 9015 21767 9031
rect 21701 8981 21717 9015
rect 21751 8981 21767 9015
rect 21701 8965 21767 8981
rect 22917 9015 22983 9031
rect 22917 8981 22933 9015
rect 22967 8981 22983 9015
rect 22917 8965 22983 8981
rect 23039 9015 23105 9031
rect 23039 8981 23055 9015
rect 23089 8981 23105 9015
rect 23039 8965 23105 8981
rect 24129 9015 24195 9031
rect 24129 8981 24145 9015
rect 24179 8981 24195 9015
rect 24129 8965 24195 8981
rect 24251 9015 24317 9031
rect 24251 8981 24267 9015
rect 24301 8981 24317 9015
rect 24251 8965 24317 8981
rect 24983 9015 25049 9031
rect 24983 8981 24999 9015
rect 25033 8981 25049 9015
rect 25949 9028 25979 9043
rect 26021 9028 26051 9043
rect 25949 9005 26051 9028
rect 25949 8998 25983 9005
rect 24983 8965 25049 8981
rect 25967 8971 25983 8998
rect 26017 8998 26051 9005
rect 26017 8971 26033 8998
rect 20863 8943 20893 8965
rect 21597 8943 21627 8965
rect 21719 8943 21749 8965
rect 22935 8943 22965 8965
rect 23057 8943 23087 8965
rect 24147 8943 24177 8965
rect 24269 8943 24299 8965
rect 25001 8943 25031 8965
rect 25967 8955 26033 8971
rect 13314 8843 13344 8858
rect 13410 8843 13440 8858
rect 12812 8823 12904 8839
rect 12812 8789 12855 8823
rect 12889 8789 12904 8823
rect 12812 8773 12904 8789
rect 13051 8823 13137 8839
rect 13051 8789 13087 8823
rect 13121 8789 13137 8823
rect 13051 8773 13137 8789
rect 13314 8836 13440 8843
rect 13502 8837 13532 8858
rect 13314 8820 13458 8836
rect 13314 8786 13408 8820
rect 13442 8786 13458 8820
rect 12812 8741 12842 8773
rect 13051 8741 13081 8773
rect 13314 8770 13458 8786
rect 13502 8818 13661 8837
rect 14154 8833 14184 8859
rect 14888 8833 14918 8859
rect 15010 8833 15040 8859
rect 16226 8833 16256 8859
rect 16348 8833 16378 8859
rect 17438 8833 17468 8859
rect 17560 8833 17590 8859
rect 18292 8833 18322 8859
rect 20023 8843 20053 8858
rect 20119 8843 20149 8858
rect 20023 8836 20149 8843
rect 20211 8837 20241 8858
rect 13502 8784 13615 8818
rect 13649 8784 13661 8818
rect 13314 8764 13440 8770
rect 2696 8457 2782 8473
rect 11316 8458 11388 8473
rect 11883 8462 11913 8488
rect 11979 8458 12009 8488
rect 12075 8462 12105 8488
rect 12279 8460 12309 8489
rect 13314 8739 13344 8764
rect 13410 8739 13440 8764
rect 13502 8764 13661 8784
rect 20023 8820 20167 8836
rect 20023 8786 20117 8820
rect 20151 8786 20167 8820
rect 13502 8739 13532 8764
rect 14151 8742 14181 8770
rect 14277 8742 14307 8770
rect 15363 8742 15393 8770
rect 15489 8742 15519 8770
rect 16575 8742 16605 8770
rect 16701 8742 16731 8770
rect 17787 8742 17817 8770
rect 17913 8742 17943 8770
rect 18645 8745 18675 8773
rect 20023 8770 20167 8786
rect 20211 8818 20370 8837
rect 20863 8833 20893 8859
rect 21597 8833 21627 8859
rect 21719 8833 21749 8859
rect 22935 8833 22965 8859
rect 23057 8833 23087 8859
rect 24147 8833 24177 8859
rect 24269 8833 24299 8859
rect 25001 8833 25031 8859
rect 20211 8784 20324 8818
rect 20358 8784 20370 8818
rect 20023 8764 20149 8770
rect 20023 8739 20053 8764
rect 20119 8739 20149 8764
rect 20211 8764 20370 8784
rect 20211 8739 20241 8764
rect 20860 8742 20890 8770
rect 20986 8742 21016 8770
rect 22072 8742 22102 8770
rect 22198 8742 22228 8770
rect 23284 8742 23314 8770
rect 23410 8742 23440 8770
rect 24496 8742 24526 8770
rect 24622 8742 24652 8770
rect 25354 8745 25384 8773
rect 13314 8624 13344 8655
rect 13410 8629 13440 8655
rect 13502 8601 13532 8655
rect 14151 8627 14181 8658
rect 14277 8627 14307 8658
rect 15363 8627 15393 8658
rect 15489 8627 15519 8658
rect 16575 8627 16605 8658
rect 16701 8627 16731 8658
rect 17787 8627 17817 8658
rect 17913 8627 17943 8658
rect 18645 8630 18675 8661
rect 14133 8611 14199 8627
rect 12728 8515 12758 8541
rect 12812 8515 12842 8541
rect 13051 8515 13081 8541
rect 14133 8577 14149 8611
rect 14183 8577 14199 8611
rect 14133 8561 14199 8577
rect 14259 8611 14325 8627
rect 14259 8577 14275 8611
rect 14309 8577 14325 8611
rect 14259 8561 14325 8577
rect 15345 8611 15411 8627
rect 15345 8577 15361 8611
rect 15395 8577 15411 8611
rect 15345 8561 15411 8577
rect 15471 8611 15537 8627
rect 15471 8577 15487 8611
rect 15521 8577 15537 8611
rect 15471 8561 15537 8577
rect 16557 8611 16623 8627
rect 16557 8577 16573 8611
rect 16607 8577 16623 8611
rect 16557 8561 16623 8577
rect 16683 8611 16749 8627
rect 16683 8577 16699 8611
rect 16733 8577 16749 8611
rect 16683 8561 16749 8577
rect 17769 8611 17835 8627
rect 17769 8577 17785 8611
rect 17819 8577 17835 8611
rect 17769 8561 17835 8577
rect 17895 8611 17961 8627
rect 17895 8577 17911 8611
rect 17945 8577 17961 8611
rect 17895 8561 17961 8577
rect 18627 8614 18693 8630
rect 18627 8580 18643 8614
rect 18677 8580 18693 8614
rect 19565 8613 19595 8639
rect 19755 8613 19785 8639
rect 20023 8624 20053 8655
rect 20119 8629 20149 8655
rect 18627 8564 18693 8580
rect 13502 8486 13532 8517
rect 20211 8601 20241 8655
rect 20860 8627 20890 8658
rect 20986 8627 21016 8658
rect 22072 8627 22102 8658
rect 22198 8627 22228 8658
rect 23284 8627 23314 8658
rect 23410 8627 23440 8658
rect 24496 8627 24526 8658
rect 24622 8627 24652 8658
rect 25354 8630 25384 8661
rect 20842 8611 20908 8627
rect 20842 8577 20858 8611
rect 20892 8577 20908 8611
rect 20842 8561 20908 8577
rect 20968 8611 21034 8627
rect 20968 8577 20984 8611
rect 21018 8577 21034 8611
rect 20968 8561 21034 8577
rect 22054 8611 22120 8627
rect 22054 8577 22070 8611
rect 22104 8577 22120 8611
rect 22054 8561 22120 8577
rect 22180 8611 22246 8627
rect 22180 8577 22196 8611
rect 22230 8577 22246 8611
rect 22180 8561 22246 8577
rect 23266 8611 23332 8627
rect 23266 8577 23282 8611
rect 23316 8577 23332 8611
rect 23266 8561 23332 8577
rect 23392 8611 23458 8627
rect 23392 8577 23408 8611
rect 23442 8577 23458 8611
rect 23392 8561 23458 8577
rect 24478 8611 24544 8627
rect 24478 8577 24494 8611
rect 24528 8577 24544 8611
rect 24478 8561 24544 8577
rect 24604 8611 24670 8627
rect 24604 8577 24620 8611
rect 24654 8577 24670 8611
rect 24604 8561 24670 8577
rect 25336 8614 25402 8630
rect 25336 8580 25352 8614
rect 25386 8580 25402 8614
rect 26274 8613 26304 8639
rect 26464 8613 26494 8639
rect 25336 8564 25402 8580
rect 20211 8486 20241 8517
rect 19565 8461 19595 8483
rect 2696 8423 2732 8457
rect 2766 8423 2782 8457
rect 2696 8407 2782 8423
rect 2696 8375 2726 8407
rect 12480 8432 12510 8460
rect 19509 8445 19595 8461
rect 2956 8383 3022 8399
rect 19509 8411 19525 8445
rect 19559 8411 19595 8445
rect 19509 8395 19595 8411
rect 2956 8349 2972 8383
rect 3006 8349 3022 8383
rect 2956 8333 3022 8349
rect 11883 8336 11913 8362
rect 11979 8336 12009 8366
rect 12075 8336 12105 8362
rect 2974 8302 3004 8333
rect 10133 8285 10163 8311
rect 10960 8285 10990 8311
rect 2506 8149 2536 8175
rect 2696 8149 2726 8175
rect 2974 8164 3004 8218
rect 2974 8026 3004 8080
rect 10242 8246 10272 8272
rect 10345 8246 10375 8272
rect 10559 8246 10589 8272
rect 10631 8246 10661 8272
rect 10727 8246 10757 8272
rect 10133 8053 10163 8085
rect 10242 8053 10272 8162
rect 10345 8147 10375 8162
rect 10345 8117 10493 8147
rect 10559 8130 10589 8162
rect 10130 8037 10184 8053
rect 10130 8003 10140 8037
rect 10174 8003 10184 8037
rect 10130 7987 10184 8003
rect 10226 8037 10280 8053
rect 10226 8003 10236 8037
rect 10270 8003 10280 8037
rect 10463 8017 10493 8117
rect 10535 8114 10589 8130
rect 10535 8080 10545 8114
rect 10579 8080 10589 8114
rect 10535 8064 10589 8080
rect 10226 7987 10280 8003
rect 10338 8001 10421 8017
rect 10133 7965 10163 7987
rect 2974 7888 3004 7942
rect 10242 7919 10272 7987
rect 10338 7967 10377 8001
rect 10411 7967 10421 8001
rect 10338 7951 10421 7967
rect 10463 8001 10517 8017
rect 10631 8011 10661 8162
rect 10727 8130 10757 8162
rect 10703 8114 10757 8130
rect 10703 8080 10713 8114
rect 10747 8080 10757 8114
rect 11069 8246 11099 8272
rect 11172 8246 11202 8272
rect 11386 8246 11416 8272
rect 11458 8246 11488 8272
rect 11554 8246 11584 8272
rect 10703 8064 10757 8080
rect 10463 7967 10473 8001
rect 10507 7967 10517 8001
rect 10619 8001 10685 8011
rect 10619 7987 10635 8001
rect 10463 7951 10517 7967
rect 10559 7967 10635 7987
rect 10669 7967 10685 8001
rect 10559 7957 10685 7967
rect 10338 7919 10368 7951
rect 10463 7919 10493 7951
rect 10559 7919 10589 7957
rect 10727 7919 10757 8064
rect 10960 8053 10990 8085
rect 11069 8053 11099 8162
rect 11172 8147 11202 8162
rect 11172 8117 11320 8147
rect 11386 8130 11416 8162
rect 10957 8037 11011 8053
rect 10957 8003 10967 8037
rect 11001 8003 11011 8037
rect 10957 7987 11011 8003
rect 11053 8037 11107 8053
rect 11053 8003 11063 8037
rect 11097 8003 11107 8037
rect 11290 8017 11320 8117
rect 11362 8114 11416 8130
rect 11362 8080 11372 8114
rect 11406 8080 11416 8114
rect 11362 8064 11416 8080
rect 11053 7987 11107 8003
rect 11165 8001 11248 8017
rect 10960 7965 10990 7987
rect 11069 7919 11099 7987
rect 11165 7967 11204 8001
rect 11238 7967 11248 8001
rect 11165 7951 11248 7967
rect 11290 8001 11344 8017
rect 11458 8011 11488 8162
rect 11554 8130 11584 8162
rect 11530 8114 11584 8130
rect 11530 8080 11540 8114
rect 11574 8080 11584 8114
rect 12279 8335 12309 8364
rect 11530 8064 11584 8080
rect 11290 7967 11300 8001
rect 11334 7967 11344 8001
rect 11446 8001 11512 8011
rect 11446 7987 11462 8001
rect 11290 7951 11344 7967
rect 11386 7967 11462 7987
rect 11496 7967 11512 8001
rect 11386 7957 11512 7967
rect 11165 7919 11195 7951
rect 11290 7919 11320 7951
rect 11386 7919 11416 7957
rect 11554 7919 11584 8064
rect 11883 8069 11913 8084
rect 11979 8069 12009 8084
rect 12075 8069 12105 8084
rect 19269 8371 19335 8387
rect 19269 8337 19285 8371
rect 19319 8337 19335 8371
rect 19565 8363 19595 8395
rect 19755 8461 19785 8483
rect 26274 8461 26304 8483
rect 19755 8445 19841 8461
rect 19755 8411 19791 8445
rect 19825 8411 19841 8445
rect 19755 8395 19841 8411
rect 26218 8445 26304 8461
rect 26218 8411 26234 8445
rect 26268 8411 26304 8445
rect 26218 8395 26304 8411
rect 19755 8363 19785 8395
rect 25978 8371 26044 8387
rect 19269 8321 19335 8337
rect 19287 8290 19317 8321
rect 12730 8224 12796 8240
rect 12730 8190 12746 8224
rect 12780 8190 12796 8224
rect 12730 8174 12796 8190
rect 12748 8152 12778 8174
rect 11883 8053 12105 8069
rect 11883 8039 12123 8053
rect 12279 8052 12309 8083
rect 19287 8152 19317 8206
rect 25978 8337 25994 8371
rect 26028 8337 26044 8371
rect 26274 8363 26304 8395
rect 26464 8461 26494 8483
rect 26464 8445 26550 8461
rect 26464 8411 26500 8445
rect 26534 8411 26550 8445
rect 26464 8395 26550 8411
rect 26464 8363 26494 8395
rect 25978 8321 26044 8337
rect 25996 8290 26026 8321
rect 12057 8037 12123 8039
rect 12057 8003 12073 8037
rect 12107 8003 12123 8037
rect 12057 7997 12123 8003
rect 11883 7974 12123 7997
rect 12261 8036 12327 8052
rect 12748 8042 12778 8068
rect 19565 8137 19595 8163
rect 19755 8137 19785 8163
rect 25996 8152 26026 8206
rect 12261 8002 12277 8036
rect 12311 8002 12327 8036
rect 12261 7986 12327 8002
rect 11883 7967 12105 7974
rect 11883 7952 11913 7967
rect 11979 7952 12009 7967
rect 12075 7952 12105 7967
rect 12279 7964 12309 7986
rect 12748 7964 12778 7994
rect 19287 8014 19317 8068
rect 26274 8137 26304 8163
rect 26464 8137 26494 8163
rect 11883 7842 11913 7868
rect 11979 7842 12009 7868
rect 12075 7842 12105 7868
rect 12279 7854 12309 7880
rect 10133 7809 10163 7835
rect 10242 7809 10272 7835
rect 10338 7809 10368 7835
rect 10463 7809 10493 7835
rect 10559 7809 10589 7835
rect 10727 7809 10757 7835
rect 10960 7809 10990 7835
rect 11069 7809 11099 7835
rect 11165 7809 11195 7835
rect 11290 7809 11320 7835
rect 11386 7809 11416 7835
rect 11554 7809 11584 7835
rect 2974 7750 3004 7804
rect 2974 7612 3004 7666
rect 25996 8014 26026 8068
rect 19287 7876 19317 7930
rect 25996 7876 26026 7930
rect 19287 7738 19317 7792
rect 25996 7738 26026 7792
rect 19287 7600 19317 7654
rect 2974 7498 3004 7528
rect 12748 7553 12778 7584
rect 12730 7537 12796 7553
rect 12730 7503 12746 7537
rect 12780 7503 12796 7537
rect 12730 7487 12796 7503
rect 25996 7600 26026 7654
rect 19287 7486 19317 7516
rect 25996 7486 26026 7516
rect 24587 7296 24617 7326
rect 24587 7158 24617 7212
rect 11577 7030 11607 7056
rect 11665 7030 11695 7056
rect 11853 7030 11883 7056
rect 11937 7030 11967 7056
rect 12021 7030 12051 7056
rect 12105 7030 12135 7056
rect 12189 7030 12219 7056
rect 12852 7030 12882 7056
rect 12936 7030 12966 7056
rect 13036 7030 13066 7056
rect 13120 7030 13150 7056
rect 13217 7030 13247 7056
rect 13318 7030 13348 7056
rect 13402 7030 13432 7056
rect 13537 7030 13567 7056
rect 11577 6857 11607 6872
rect 11571 6833 11607 6857
rect 11571 6798 11601 6833
rect 11665 6811 11695 6872
rect 11525 6782 11601 6798
rect 11525 6748 11535 6782
rect 11569 6748 11601 6782
rect 11525 6732 11601 6748
rect 11643 6795 11697 6811
rect 11643 6761 11653 6795
rect 11687 6761 11697 6795
rect 11853 6794 11883 6830
rect 11643 6745 11697 6761
rect 11802 6782 11883 6794
rect 11937 6792 11967 6830
rect 12021 6792 12051 6830
rect 12105 6792 12135 6830
rect 12189 6792 12219 6830
rect 11802 6748 11818 6782
rect 11852 6748 11883 6782
rect 11571 6723 11601 6732
rect 11571 6699 11607 6723
rect 11577 6684 11607 6699
rect 11665 6684 11695 6745
rect 11802 6736 11883 6748
rect 11936 6782 12219 6792
rect 11936 6748 11952 6782
rect 11986 6748 12219 6782
rect 11936 6738 12219 6748
rect 11853 6710 11883 6736
rect 11937 6710 11967 6738
rect 12021 6710 12051 6738
rect 12105 6710 12135 6738
rect 12189 6710 12219 6738
rect 12852 6798 12882 6830
rect 12936 6798 12966 6830
rect 13036 6798 13066 6830
rect 13120 6798 13150 6830
rect 13217 6798 13247 6902
rect 13318 6848 13348 6946
rect 13402 6908 13432 6946
rect 13390 6898 13456 6908
rect 13725 7026 14027 7056
rect 13725 6957 13755 7026
rect 13997 7006 14027 7026
rect 14081 7006 14111 7056
rect 14225 7030 14255 7056
rect 14309 7030 14339 7056
rect 14405 7030 14435 7056
rect 14489 7030 14519 7056
rect 13809 6957 13839 6983
rect 13390 6864 13406 6898
rect 13440 6864 13456 6898
rect 13390 6854 13456 6864
rect 13294 6832 13348 6848
rect 13294 6798 13304 6832
rect 13338 6812 13348 6832
rect 13537 6812 13567 6902
rect 14225 6908 14255 6946
rect 14201 6898 14267 6908
rect 13725 6823 13755 6849
rect 13338 6798 13456 6812
rect 12852 6782 13156 6798
rect 12852 6748 13112 6782
rect 13146 6748 13156 6782
rect 12852 6732 13156 6748
rect 13198 6782 13252 6798
rect 13294 6782 13456 6798
rect 13198 6748 13208 6782
rect 13242 6748 13252 6782
rect 13198 6732 13252 6748
rect 12852 6710 12882 6732
rect 12936 6710 12966 6732
rect 13036 6710 13066 6732
rect 13120 6710 13150 6732
rect 13221 6664 13251 6732
rect 13316 6724 13384 6740
rect 13316 6690 13340 6724
rect 13374 6690 13384 6724
rect 13316 6674 13384 6690
rect 13316 6652 13346 6674
rect 13426 6652 13456 6782
rect 13537 6796 13618 6812
rect 13537 6776 13574 6796
rect 13533 6762 13574 6776
rect 13608 6762 13618 6796
rect 13809 6805 13839 6849
rect 13809 6795 13951 6805
rect 13809 6781 13901 6795
rect 13533 6746 13618 6762
rect 13721 6761 13901 6781
rect 13935 6761 13951 6795
rect 13721 6751 13951 6761
rect 13997 6752 14027 6878
rect 14081 6863 14111 6878
rect 14201 6864 14217 6898
rect 14251 6864 14267 6898
rect 14081 6833 14134 6863
rect 14201 6854 14267 6864
rect 14309 6856 14339 6946
rect 24587 7020 24617 7074
rect 14104 6752 14134 6833
rect 14309 6840 14363 6856
rect 14309 6812 14319 6840
rect 14200 6806 14319 6812
rect 14353 6806 14363 6840
rect 14200 6790 14363 6806
rect 14200 6782 14339 6790
rect 13533 6664 13563 6746
rect 13721 6664 13751 6751
rect 13993 6736 14047 6752
rect 13993 6709 14003 6736
rect 13806 6702 14003 6709
rect 14037 6702 14047 6736
rect 13806 6686 14047 6702
rect 14089 6736 14143 6752
rect 14089 6702 14099 6736
rect 14133 6702 14143 6736
rect 14089 6686 14143 6702
rect 13806 6679 14028 6686
rect 13806 6664 13836 6679
rect 13996 6664 14026 6679
rect 14104 6664 14134 6686
rect 14200 6652 14230 6782
rect 14405 6752 14435 6902
rect 14489 6798 14519 6902
rect 24587 6882 24617 6936
rect 14489 6782 14577 6798
rect 14272 6724 14340 6740
rect 14272 6690 14282 6724
rect 14316 6690 14340 6724
rect 14272 6674 14340 6690
rect 14386 6736 14440 6752
rect 14386 6702 14396 6736
rect 14430 6702 14440 6736
rect 14386 6686 14440 6702
rect 14489 6748 14532 6782
rect 14566 6748 14577 6782
rect 14489 6732 14577 6748
rect 24587 6744 24617 6798
rect 14310 6652 14340 6674
rect 14405 6664 14435 6686
rect 14489 6664 14519 6732
rect 24119 6649 24149 6675
rect 24309 6649 24339 6675
rect 11577 6554 11607 6580
rect 11665 6554 11695 6580
rect 11853 6554 11883 6580
rect 11937 6554 11967 6580
rect 12021 6554 12051 6580
rect 12105 6554 12135 6580
rect 12189 6554 12219 6580
rect 12852 6554 12882 6580
rect 12936 6554 12966 6580
rect 13036 6554 13066 6580
rect 13120 6554 13150 6580
rect 13221 6554 13251 6580
rect 13316 6554 13346 6580
rect 13426 6554 13456 6580
rect 13533 6554 13563 6580
rect 13721 6554 13751 6580
rect 13806 6554 13836 6580
rect 13996 6554 14026 6580
rect 14104 6554 14134 6580
rect 14200 6554 14230 6580
rect 14310 6554 14340 6580
rect 14405 6554 14435 6580
rect 14489 6554 14519 6580
rect 24587 6606 24617 6660
rect 24587 6491 24617 6522
rect 24569 6475 24635 6491
rect 24119 6417 24149 6449
rect 24063 6401 24149 6417
rect 24063 6367 24079 6401
rect 24113 6367 24149 6401
rect 24063 6351 24149 6367
rect 24119 6329 24149 6351
rect 24309 6417 24339 6449
rect 24569 6441 24585 6475
rect 24619 6441 24635 6475
rect 24569 6425 24635 6441
rect 24309 6401 24395 6417
rect 24309 6367 24345 6401
rect 24379 6367 24395 6401
rect 24309 6351 24395 6367
rect 24309 6329 24339 6351
rect 13381 6236 13447 6246
rect 13381 6202 13397 6236
rect 13431 6202 13447 6236
rect 14624 6239 14690 6249
rect 13381 6192 13447 6202
rect 14624 6205 14640 6239
rect 14674 6205 14690 6239
rect 17016 6241 17082 6251
rect 14624 6195 14690 6205
rect 17016 6207 17032 6241
rect 17066 6207 17082 6241
rect 19408 6241 19474 6251
rect 17016 6197 17082 6207
rect 19408 6207 19424 6241
rect 19458 6207 19474 6241
rect 21800 6242 21866 6252
rect 19408 6197 19474 6207
rect 21800 6208 21816 6242
rect 21850 6208 21866 6242
rect 21800 6198 21866 6208
rect 30372 6295 30402 6326
rect 25211 6232 25277 6248
rect 11576 6151 11606 6177
rect 11660 6151 11690 6177
rect 11848 6157 11878 6183
rect 11941 6157 11971 6183
rect 12025 6157 12055 6183
rect 12145 6157 12175 6183
rect 12251 6157 12281 6183
rect 12359 6157 12389 6183
rect 12443 6157 12473 6183
rect 12580 6157 12610 6183
rect 12724 6157 12754 6183
rect 12808 6157 12838 6183
rect 12926 6157 12956 6183
rect 13034 6157 13064 6183
rect 13130 6157 13160 6183
rect 13202 6157 13232 6183
rect 11576 6008 11606 6023
rect 11543 5978 11606 6008
rect 11543 5940 11573 5978
rect 11518 5924 11573 5940
rect 11660 5934 11690 6023
rect 11518 5890 11529 5924
rect 11563 5890 11573 5924
rect 11518 5874 11573 5890
rect 11615 5924 11690 5934
rect 11848 5927 11878 6073
rect 11941 5939 11971 6073
rect 12025 6035 12055 6073
rect 12145 6041 12175 6073
rect 12013 6025 12079 6035
rect 12013 5991 12029 6025
rect 12063 5991 12079 6025
rect 12013 5981 12079 5991
rect 12145 6025 12209 6041
rect 12145 5991 12165 6025
rect 12199 5991 12209 6025
rect 12145 5975 12209 5991
rect 11615 5890 11631 5924
rect 11665 5890 11690 5924
rect 11615 5880 11690 5890
rect 11543 5836 11573 5874
rect 11543 5806 11606 5836
rect 11576 5791 11606 5806
rect 11660 5791 11690 5880
rect 11837 5911 11891 5927
rect 11837 5877 11847 5911
rect 11881 5877 11891 5911
rect 11941 5909 12079 5939
rect 11837 5861 11891 5877
rect 12049 5879 12079 5909
rect 11848 5791 11878 5861
rect 11943 5851 12007 5867
rect 11943 5817 11963 5851
rect 11997 5817 12007 5851
rect 11943 5801 12007 5817
rect 12049 5863 12103 5879
rect 12049 5829 12059 5863
rect 12093 5829 12103 5863
rect 12049 5813 12103 5829
rect 11943 5779 11973 5801
rect 12049 5779 12079 5813
rect 12145 5791 12175 5975
rect 12251 5889 12281 6073
rect 12724 6041 12754 6073
rect 12700 6025 12754 6041
rect 12808 6035 12838 6073
rect 12926 6041 12956 6073
rect 12700 5991 12710 6025
rect 12744 5991 12754 6025
rect 12359 5957 12389 5989
rect 12443 5957 12473 5989
rect 12323 5941 12389 5957
rect 12323 5907 12333 5941
rect 12367 5907 12389 5941
rect 12323 5891 12389 5907
rect 12439 5941 12529 5957
rect 12439 5907 12485 5941
rect 12519 5907 12529 5941
rect 12439 5891 12529 5907
rect 12580 5923 12610 5989
rect 12700 5975 12754 5991
rect 12796 6025 12862 6035
rect 12796 5991 12812 6025
rect 12846 5991 12862 6025
rect 12796 5981 12862 5991
rect 12926 6025 12992 6041
rect 12926 5991 12948 6025
rect 12982 5991 12992 6025
rect 12724 5939 12754 5975
rect 12926 5975 12992 5991
rect 12580 5907 12657 5923
rect 12724 5909 12861 5939
rect 12580 5893 12613 5907
rect 12221 5873 12281 5889
rect 12221 5839 12231 5873
rect 12265 5853 12281 5873
rect 12265 5839 12285 5853
rect 12221 5823 12285 5839
rect 12355 5835 12385 5891
rect 12439 5835 12469 5891
rect 12603 5873 12613 5893
rect 12647 5873 12657 5907
rect 12603 5857 12657 5873
rect 12627 5835 12657 5857
rect 12722 5851 12789 5867
rect 12255 5791 12285 5823
rect 12722 5817 12745 5851
rect 12779 5817 12789 5851
rect 12722 5801 12789 5817
rect 12722 5779 12752 5801
rect 12831 5779 12861 5909
rect 12926 5791 12956 5975
rect 13034 5889 13064 6073
rect 13400 6089 13430 6192
rect 13497 6157 13527 6183
rect 13130 5941 13160 5989
rect 12998 5873 13064 5889
rect 13106 5925 13160 5941
rect 13202 5957 13232 5989
rect 13202 5941 13298 5957
rect 13202 5927 13254 5941
rect 13106 5891 13116 5925
rect 13150 5891 13160 5925
rect 13106 5875 13160 5891
rect 12998 5839 13008 5873
rect 13042 5839 13064 5873
rect 12998 5823 13064 5839
rect 13130 5835 13160 5875
rect 13214 5907 13254 5927
rect 13288 5907 13298 5941
rect 13400 5929 13430 5961
rect 13685 6141 13715 6167
rect 13780 6157 13810 6183
rect 13685 5997 13715 6013
rect 13659 5967 13715 5997
rect 13214 5891 13298 5907
rect 13369 5913 13433 5929
rect 13497 5925 13527 5957
rect 13214 5835 13244 5891
rect 13369 5879 13385 5913
rect 13419 5879 13433 5913
rect 13369 5863 13433 5879
rect 13475 5919 13527 5925
rect 13659 5919 13689 5967
rect 13968 6151 13998 6177
rect 14052 6151 14082 6177
rect 14240 6157 14270 6183
rect 14333 6157 14363 6183
rect 14417 6157 14447 6183
rect 14537 6157 14567 6183
rect 14643 6157 14673 6195
rect 14751 6157 14781 6183
rect 14835 6157 14865 6183
rect 14972 6157 15002 6183
rect 15116 6157 15146 6183
rect 15200 6157 15230 6183
rect 15318 6157 15348 6183
rect 15426 6157 15456 6183
rect 15522 6157 15552 6183
rect 15594 6157 15624 6183
rect 15889 6157 15919 6183
rect 13968 6008 13998 6023
rect 13935 5978 13998 6008
rect 13780 5925 13810 5957
rect 13935 5940 13965 5978
rect 13475 5909 13689 5919
rect 13475 5875 13485 5909
rect 13519 5875 13689 5909
rect 13475 5865 13689 5875
rect 13012 5791 13042 5823
rect 13402 5791 13432 5863
rect 13475 5859 13527 5865
rect 13497 5837 13527 5859
rect 13659 5836 13689 5865
rect 13751 5909 13810 5925
rect 13751 5875 13761 5909
rect 13795 5875 13810 5909
rect 13751 5859 13810 5875
rect 13910 5924 13965 5940
rect 14052 5934 14082 6023
rect 13910 5890 13921 5924
rect 13955 5890 13965 5924
rect 13910 5874 13965 5890
rect 14007 5924 14082 5934
rect 14240 5927 14270 6073
rect 14333 5939 14363 6073
rect 14417 6035 14447 6073
rect 14537 6041 14567 6073
rect 14405 6025 14471 6035
rect 14405 5991 14421 6025
rect 14455 5991 14471 6025
rect 14405 5981 14471 5991
rect 14537 6025 14601 6041
rect 14537 5991 14557 6025
rect 14591 5991 14601 6025
rect 14537 5975 14601 5991
rect 14007 5890 14023 5924
rect 14057 5890 14082 5924
rect 14007 5880 14082 5890
rect 13780 5837 13810 5859
rect 13659 5806 13715 5836
rect 13685 5791 13715 5806
rect 13935 5836 13965 5874
rect 13935 5806 13998 5836
rect 13968 5791 13998 5806
rect 14052 5791 14082 5880
rect 14229 5911 14283 5927
rect 14229 5877 14239 5911
rect 14273 5877 14283 5911
rect 14333 5909 14471 5939
rect 14229 5861 14283 5877
rect 14441 5879 14471 5909
rect 14240 5791 14270 5861
rect 14335 5851 14399 5867
rect 14335 5817 14355 5851
rect 14389 5817 14399 5851
rect 14335 5801 14399 5817
rect 14441 5863 14495 5879
rect 14441 5829 14451 5863
rect 14485 5829 14495 5863
rect 14441 5813 14495 5829
rect 14335 5779 14365 5801
rect 14441 5779 14471 5813
rect 14537 5791 14567 5975
rect 14643 5889 14673 6073
rect 15116 6041 15146 6073
rect 15092 6025 15146 6041
rect 15200 6035 15230 6073
rect 15318 6041 15348 6073
rect 15092 5991 15102 6025
rect 15136 5991 15146 6025
rect 14751 5957 14781 5989
rect 14835 5957 14865 5989
rect 14715 5941 14781 5957
rect 14715 5907 14725 5941
rect 14759 5907 14781 5941
rect 14715 5891 14781 5907
rect 14831 5941 14921 5957
rect 14831 5907 14877 5941
rect 14911 5907 14921 5941
rect 14831 5891 14921 5907
rect 14972 5923 15002 5989
rect 15092 5975 15146 5991
rect 15188 6025 15254 6035
rect 15188 5991 15204 6025
rect 15238 5991 15254 6025
rect 15188 5981 15254 5991
rect 15318 6025 15384 6041
rect 15318 5991 15340 6025
rect 15374 5991 15384 6025
rect 15116 5939 15146 5975
rect 15318 5975 15384 5991
rect 14972 5907 15049 5923
rect 15116 5909 15253 5939
rect 14972 5893 15005 5907
rect 14613 5873 14673 5889
rect 14613 5839 14623 5873
rect 14657 5853 14673 5873
rect 14657 5839 14677 5853
rect 14613 5823 14677 5839
rect 14747 5835 14777 5891
rect 14831 5835 14861 5891
rect 14995 5873 15005 5893
rect 15039 5873 15049 5907
rect 14995 5857 15049 5873
rect 15019 5835 15049 5857
rect 15114 5851 15181 5867
rect 14647 5791 14677 5823
rect 15114 5817 15137 5851
rect 15171 5817 15181 5851
rect 15114 5801 15181 5817
rect 15114 5779 15144 5801
rect 15223 5779 15253 5909
rect 15318 5791 15348 5975
rect 15426 5889 15456 6073
rect 15792 6089 15822 6115
rect 15522 5941 15552 5989
rect 15390 5873 15456 5889
rect 15498 5925 15552 5941
rect 15594 5957 15624 5989
rect 15594 5941 15690 5957
rect 15594 5927 15646 5941
rect 15498 5891 15508 5925
rect 15542 5891 15552 5925
rect 15498 5875 15552 5891
rect 15390 5839 15400 5873
rect 15434 5839 15456 5873
rect 15390 5823 15456 5839
rect 15522 5835 15552 5875
rect 15606 5907 15646 5927
rect 15680 5907 15690 5941
rect 15792 5929 15822 5961
rect 16077 6141 16107 6167
rect 16172 6157 16202 6183
rect 16077 5997 16107 6013
rect 16051 5967 16107 5997
rect 15606 5891 15690 5907
rect 15761 5913 15825 5929
rect 15889 5925 15919 5957
rect 15606 5835 15636 5891
rect 15761 5879 15777 5913
rect 15811 5879 15825 5913
rect 15761 5863 15825 5879
rect 15867 5919 15919 5925
rect 16051 5919 16081 5967
rect 16360 6151 16390 6177
rect 16444 6151 16474 6177
rect 16632 6157 16662 6183
rect 16725 6157 16755 6183
rect 16809 6157 16839 6183
rect 16929 6157 16959 6183
rect 17035 6157 17065 6197
rect 17143 6157 17173 6183
rect 17227 6157 17257 6183
rect 17364 6157 17394 6183
rect 17508 6157 17538 6183
rect 17592 6157 17622 6183
rect 17710 6157 17740 6183
rect 17818 6157 17848 6183
rect 17914 6157 17944 6183
rect 17986 6157 18016 6183
rect 18281 6157 18311 6183
rect 16360 6008 16390 6023
rect 16327 5978 16390 6008
rect 16172 5925 16202 5957
rect 16327 5940 16357 5978
rect 15867 5909 16081 5919
rect 15867 5875 15877 5909
rect 15911 5875 16081 5909
rect 15867 5865 16081 5875
rect 15404 5791 15434 5823
rect 15794 5791 15824 5863
rect 15867 5859 15919 5865
rect 15889 5837 15919 5859
rect 16051 5836 16081 5865
rect 16143 5909 16202 5925
rect 16143 5875 16153 5909
rect 16187 5875 16202 5909
rect 16143 5859 16202 5875
rect 16302 5924 16357 5940
rect 16444 5934 16474 6023
rect 16302 5890 16313 5924
rect 16347 5890 16357 5924
rect 16302 5874 16357 5890
rect 16399 5924 16474 5934
rect 16632 5927 16662 6073
rect 16725 5939 16755 6073
rect 16809 6035 16839 6073
rect 16929 6041 16959 6073
rect 16797 6025 16863 6035
rect 16797 5991 16813 6025
rect 16847 5991 16863 6025
rect 16797 5981 16863 5991
rect 16929 6025 16993 6041
rect 16929 5991 16949 6025
rect 16983 5991 16993 6025
rect 16929 5975 16993 5991
rect 16399 5890 16415 5924
rect 16449 5890 16474 5924
rect 16399 5880 16474 5890
rect 16172 5837 16202 5859
rect 16051 5806 16107 5836
rect 16077 5791 16107 5806
rect 16327 5836 16357 5874
rect 16327 5806 16390 5836
rect 16360 5791 16390 5806
rect 16444 5791 16474 5880
rect 16621 5911 16675 5927
rect 16621 5877 16631 5911
rect 16665 5877 16675 5911
rect 16725 5909 16863 5939
rect 16621 5861 16675 5877
rect 16833 5879 16863 5909
rect 16632 5791 16662 5861
rect 16727 5851 16791 5867
rect 16727 5817 16747 5851
rect 16781 5817 16791 5851
rect 16727 5801 16791 5817
rect 16833 5863 16887 5879
rect 16833 5829 16843 5863
rect 16877 5829 16887 5863
rect 16833 5813 16887 5829
rect 16727 5779 16757 5801
rect 16833 5779 16863 5813
rect 16929 5791 16959 5975
rect 17035 5889 17065 6073
rect 17508 6041 17538 6073
rect 17484 6025 17538 6041
rect 17592 6035 17622 6073
rect 17710 6041 17740 6073
rect 17484 5991 17494 6025
rect 17528 5991 17538 6025
rect 17143 5957 17173 5989
rect 17227 5957 17257 5989
rect 17107 5941 17173 5957
rect 17107 5907 17117 5941
rect 17151 5907 17173 5941
rect 17107 5891 17173 5907
rect 17223 5941 17313 5957
rect 17223 5907 17269 5941
rect 17303 5907 17313 5941
rect 17223 5891 17313 5907
rect 17364 5923 17394 5989
rect 17484 5975 17538 5991
rect 17580 6025 17646 6035
rect 17580 5991 17596 6025
rect 17630 5991 17646 6025
rect 17580 5981 17646 5991
rect 17710 6025 17776 6041
rect 17710 5991 17732 6025
rect 17766 5991 17776 6025
rect 17508 5939 17538 5975
rect 17710 5975 17776 5991
rect 17364 5907 17441 5923
rect 17508 5909 17645 5939
rect 17364 5893 17397 5907
rect 17005 5873 17065 5889
rect 17005 5839 17015 5873
rect 17049 5853 17065 5873
rect 17049 5839 17069 5853
rect 17005 5823 17069 5839
rect 17139 5835 17169 5891
rect 17223 5835 17253 5891
rect 17387 5873 17397 5893
rect 17431 5873 17441 5907
rect 17387 5857 17441 5873
rect 17411 5835 17441 5857
rect 17506 5851 17573 5867
rect 17039 5791 17069 5823
rect 17506 5817 17529 5851
rect 17563 5817 17573 5851
rect 17506 5801 17573 5817
rect 17506 5779 17536 5801
rect 17615 5779 17645 5909
rect 17710 5791 17740 5975
rect 17818 5889 17848 6073
rect 18184 6089 18214 6115
rect 17914 5941 17944 5989
rect 17782 5873 17848 5889
rect 17890 5925 17944 5941
rect 17986 5957 18016 5989
rect 17986 5941 18082 5957
rect 17986 5927 18038 5941
rect 17890 5891 17900 5925
rect 17934 5891 17944 5925
rect 17890 5875 17944 5891
rect 17782 5839 17792 5873
rect 17826 5839 17848 5873
rect 17782 5823 17848 5839
rect 17914 5835 17944 5875
rect 17998 5907 18038 5927
rect 18072 5907 18082 5941
rect 18184 5929 18214 5961
rect 18469 6141 18499 6167
rect 18564 6157 18594 6183
rect 18469 5997 18499 6013
rect 18443 5967 18499 5997
rect 17998 5891 18082 5907
rect 18153 5913 18217 5929
rect 18281 5925 18311 5957
rect 17998 5835 18028 5891
rect 18153 5879 18169 5913
rect 18203 5879 18217 5913
rect 18153 5863 18217 5879
rect 18259 5919 18311 5925
rect 18443 5919 18473 5967
rect 18752 6151 18782 6177
rect 18836 6151 18866 6177
rect 19024 6157 19054 6183
rect 19117 6157 19147 6183
rect 19201 6157 19231 6183
rect 19321 6157 19351 6183
rect 19427 6157 19457 6197
rect 19535 6157 19565 6183
rect 19619 6157 19649 6183
rect 19756 6157 19786 6183
rect 19900 6157 19930 6183
rect 19984 6157 20014 6183
rect 20102 6157 20132 6183
rect 20210 6157 20240 6183
rect 20306 6157 20336 6183
rect 20378 6157 20408 6183
rect 20673 6157 20703 6183
rect 18752 6008 18782 6023
rect 18719 5978 18782 6008
rect 18564 5925 18594 5957
rect 18719 5940 18749 5978
rect 18259 5909 18473 5919
rect 18259 5875 18269 5909
rect 18303 5875 18473 5909
rect 18259 5865 18473 5875
rect 17796 5791 17826 5823
rect 18186 5791 18216 5863
rect 18259 5859 18311 5865
rect 18281 5837 18311 5859
rect 18443 5836 18473 5865
rect 18535 5909 18594 5925
rect 18535 5875 18545 5909
rect 18579 5875 18594 5909
rect 18535 5859 18594 5875
rect 18694 5924 18749 5940
rect 18836 5934 18866 6023
rect 18694 5890 18705 5924
rect 18739 5890 18749 5924
rect 18694 5874 18749 5890
rect 18791 5924 18866 5934
rect 19024 5927 19054 6073
rect 19117 5939 19147 6073
rect 19201 6035 19231 6073
rect 19321 6041 19351 6073
rect 19189 6025 19255 6035
rect 19189 5991 19205 6025
rect 19239 5991 19255 6025
rect 19189 5981 19255 5991
rect 19321 6025 19385 6041
rect 19321 5991 19341 6025
rect 19375 5991 19385 6025
rect 19321 5975 19385 5991
rect 18791 5890 18807 5924
rect 18841 5890 18866 5924
rect 18791 5880 18866 5890
rect 18564 5837 18594 5859
rect 18443 5806 18499 5836
rect 18469 5791 18499 5806
rect 18719 5836 18749 5874
rect 18719 5806 18782 5836
rect 18752 5791 18782 5806
rect 18836 5791 18866 5880
rect 19013 5911 19067 5927
rect 19013 5877 19023 5911
rect 19057 5877 19067 5911
rect 19117 5909 19255 5939
rect 19013 5861 19067 5877
rect 19225 5879 19255 5909
rect 19024 5791 19054 5861
rect 19119 5851 19183 5867
rect 19119 5817 19139 5851
rect 19173 5817 19183 5851
rect 19119 5801 19183 5817
rect 19225 5863 19279 5879
rect 19225 5829 19235 5863
rect 19269 5829 19279 5863
rect 19225 5813 19279 5829
rect 19119 5779 19149 5801
rect 19225 5779 19255 5813
rect 19321 5791 19351 5975
rect 19427 5889 19457 6073
rect 19900 6041 19930 6073
rect 19876 6025 19930 6041
rect 19984 6035 20014 6073
rect 20102 6041 20132 6073
rect 19876 5991 19886 6025
rect 19920 5991 19930 6025
rect 19535 5957 19565 5989
rect 19619 5957 19649 5989
rect 19499 5941 19565 5957
rect 19499 5907 19509 5941
rect 19543 5907 19565 5941
rect 19499 5891 19565 5907
rect 19615 5941 19705 5957
rect 19615 5907 19661 5941
rect 19695 5907 19705 5941
rect 19615 5891 19705 5907
rect 19756 5923 19786 5989
rect 19876 5975 19930 5991
rect 19972 6025 20038 6035
rect 19972 5991 19988 6025
rect 20022 5991 20038 6025
rect 19972 5981 20038 5991
rect 20102 6025 20168 6041
rect 20102 5991 20124 6025
rect 20158 5991 20168 6025
rect 19900 5939 19930 5975
rect 20102 5975 20168 5991
rect 19756 5907 19833 5923
rect 19900 5909 20037 5939
rect 19756 5893 19789 5907
rect 19397 5873 19457 5889
rect 19397 5839 19407 5873
rect 19441 5853 19457 5873
rect 19441 5839 19461 5853
rect 19397 5823 19461 5839
rect 19531 5835 19561 5891
rect 19615 5835 19645 5891
rect 19779 5873 19789 5893
rect 19823 5873 19833 5907
rect 19779 5857 19833 5873
rect 19803 5835 19833 5857
rect 19898 5851 19965 5867
rect 19431 5791 19461 5823
rect 19898 5817 19921 5851
rect 19955 5817 19965 5851
rect 19898 5801 19965 5817
rect 19898 5779 19928 5801
rect 20007 5779 20037 5909
rect 20102 5791 20132 5975
rect 20210 5889 20240 6073
rect 20576 6089 20606 6115
rect 20306 5941 20336 5989
rect 20174 5873 20240 5889
rect 20282 5925 20336 5941
rect 20378 5957 20408 5989
rect 20378 5941 20474 5957
rect 20378 5927 20430 5941
rect 20282 5891 20292 5925
rect 20326 5891 20336 5925
rect 20282 5875 20336 5891
rect 20174 5839 20184 5873
rect 20218 5839 20240 5873
rect 20174 5823 20240 5839
rect 20306 5835 20336 5875
rect 20390 5907 20430 5927
rect 20464 5907 20474 5941
rect 20576 5929 20606 5961
rect 20861 6141 20891 6167
rect 20956 6157 20986 6183
rect 20861 5997 20891 6013
rect 20835 5967 20891 5997
rect 20390 5891 20474 5907
rect 20545 5913 20609 5929
rect 20673 5925 20703 5957
rect 20390 5835 20420 5891
rect 20545 5879 20561 5913
rect 20595 5879 20609 5913
rect 20545 5863 20609 5879
rect 20651 5919 20703 5925
rect 20835 5919 20865 5967
rect 21144 6151 21174 6177
rect 21228 6151 21258 6177
rect 21416 6157 21446 6183
rect 21509 6157 21539 6183
rect 21593 6157 21623 6183
rect 21713 6157 21743 6183
rect 21819 6157 21849 6198
rect 21927 6157 21957 6183
rect 22011 6157 22041 6183
rect 22148 6157 22178 6183
rect 22292 6157 22322 6183
rect 22376 6157 22406 6183
rect 22494 6157 22524 6183
rect 22602 6157 22632 6183
rect 22698 6157 22728 6183
rect 22770 6157 22800 6183
rect 23065 6157 23095 6183
rect 21144 6008 21174 6023
rect 21111 5978 21174 6008
rect 20956 5925 20986 5957
rect 21111 5940 21141 5978
rect 20651 5909 20865 5919
rect 20651 5875 20661 5909
rect 20695 5875 20865 5909
rect 20651 5865 20865 5875
rect 20188 5791 20218 5823
rect 20578 5791 20608 5863
rect 20651 5859 20703 5865
rect 20673 5837 20703 5859
rect 20835 5836 20865 5865
rect 20927 5909 20986 5925
rect 20927 5875 20937 5909
rect 20971 5875 20986 5909
rect 20927 5859 20986 5875
rect 21086 5924 21141 5940
rect 21228 5934 21258 6023
rect 21086 5890 21097 5924
rect 21131 5890 21141 5924
rect 21086 5874 21141 5890
rect 21183 5924 21258 5934
rect 21416 5927 21446 6073
rect 21509 5939 21539 6073
rect 21593 6035 21623 6073
rect 21713 6041 21743 6073
rect 21581 6025 21647 6035
rect 21581 5991 21597 6025
rect 21631 5991 21647 6025
rect 21581 5981 21647 5991
rect 21713 6025 21777 6041
rect 21713 5991 21733 6025
rect 21767 5991 21777 6025
rect 21713 5975 21777 5991
rect 21183 5890 21199 5924
rect 21233 5890 21258 5924
rect 21183 5880 21258 5890
rect 20956 5837 20986 5859
rect 20835 5806 20891 5836
rect 20861 5791 20891 5806
rect 21111 5836 21141 5874
rect 21111 5806 21174 5836
rect 21144 5791 21174 5806
rect 21228 5791 21258 5880
rect 21405 5911 21459 5927
rect 21405 5877 21415 5911
rect 21449 5877 21459 5911
rect 21509 5909 21647 5939
rect 21405 5861 21459 5877
rect 21617 5879 21647 5909
rect 21416 5791 21446 5861
rect 21511 5851 21575 5867
rect 21511 5817 21531 5851
rect 21565 5817 21575 5851
rect 21511 5801 21575 5817
rect 21617 5863 21671 5879
rect 21617 5829 21627 5863
rect 21661 5829 21671 5863
rect 21617 5813 21671 5829
rect 21511 5779 21541 5801
rect 21617 5779 21647 5813
rect 21713 5791 21743 5975
rect 21819 5889 21849 6073
rect 22292 6041 22322 6073
rect 22268 6025 22322 6041
rect 22376 6035 22406 6073
rect 22494 6041 22524 6073
rect 22268 5991 22278 6025
rect 22312 5991 22322 6025
rect 21927 5957 21957 5989
rect 22011 5957 22041 5989
rect 21891 5941 21957 5957
rect 21891 5907 21901 5941
rect 21935 5907 21957 5941
rect 21891 5891 21957 5907
rect 22007 5941 22097 5957
rect 22007 5907 22053 5941
rect 22087 5907 22097 5941
rect 22007 5891 22097 5907
rect 22148 5923 22178 5989
rect 22268 5975 22322 5991
rect 22364 6025 22430 6035
rect 22364 5991 22380 6025
rect 22414 5991 22430 6025
rect 22364 5981 22430 5991
rect 22494 6025 22560 6041
rect 22494 5991 22516 6025
rect 22550 5991 22560 6025
rect 22292 5939 22322 5975
rect 22494 5975 22560 5991
rect 22148 5907 22225 5923
rect 22292 5909 22429 5939
rect 22148 5893 22181 5907
rect 21789 5873 21849 5889
rect 21789 5839 21799 5873
rect 21833 5853 21849 5873
rect 21833 5839 21853 5853
rect 21789 5823 21853 5839
rect 21923 5835 21953 5891
rect 22007 5835 22037 5891
rect 22171 5873 22181 5893
rect 22215 5873 22225 5907
rect 22171 5857 22225 5873
rect 22195 5835 22225 5857
rect 22290 5851 22357 5867
rect 21823 5791 21853 5823
rect 22290 5817 22313 5851
rect 22347 5817 22357 5851
rect 22290 5801 22357 5817
rect 22290 5779 22320 5801
rect 22399 5779 22429 5909
rect 22494 5791 22524 5975
rect 22602 5889 22632 6073
rect 22968 6089 22998 6115
rect 22698 5941 22728 5989
rect 22566 5873 22632 5889
rect 22674 5925 22728 5941
rect 22770 5957 22800 5989
rect 22770 5941 22866 5957
rect 22770 5927 22822 5941
rect 22674 5891 22684 5925
rect 22718 5891 22728 5925
rect 22674 5875 22728 5891
rect 22566 5839 22576 5873
rect 22610 5839 22632 5873
rect 22566 5823 22632 5839
rect 22698 5835 22728 5875
rect 22782 5907 22822 5927
rect 22856 5907 22866 5941
rect 22968 5929 22998 5961
rect 23253 6141 23283 6167
rect 23348 6157 23378 6183
rect 24119 6173 24149 6199
rect 24309 6173 24339 6199
rect 25211 6198 25227 6232
rect 25261 6198 25277 6232
rect 25211 6182 25277 6198
rect 25943 6235 26009 6251
rect 25943 6201 25959 6235
rect 25993 6201 26009 6235
rect 25943 6185 26009 6201
rect 26069 6235 26135 6251
rect 26069 6201 26085 6235
rect 26119 6201 26135 6235
rect 26069 6185 26135 6201
rect 27155 6235 27221 6251
rect 27155 6201 27171 6235
rect 27205 6201 27221 6235
rect 27155 6185 27221 6201
rect 27281 6235 27347 6251
rect 27281 6201 27297 6235
rect 27331 6201 27347 6235
rect 27281 6185 27347 6201
rect 28367 6235 28433 6251
rect 28367 6201 28383 6235
rect 28417 6201 28433 6235
rect 28367 6185 28433 6201
rect 28493 6235 28559 6251
rect 28493 6201 28509 6235
rect 28543 6201 28559 6235
rect 28493 6185 28559 6201
rect 29579 6235 29645 6251
rect 29579 6201 29595 6235
rect 29629 6201 29645 6235
rect 29579 6185 29645 6201
rect 29705 6235 29771 6251
rect 29705 6201 29721 6235
rect 29755 6201 29771 6235
rect 30758 6264 30788 6290
rect 30853 6272 30883 6298
rect 30937 6272 30967 6298
rect 29705 6185 29771 6201
rect 23253 5997 23283 6013
rect 23227 5967 23283 5997
rect 22782 5891 22866 5907
rect 22937 5913 23001 5929
rect 23065 5925 23095 5957
rect 22782 5835 22812 5891
rect 22937 5879 22953 5913
rect 22987 5879 23001 5913
rect 22937 5863 23001 5879
rect 23043 5919 23095 5925
rect 23227 5919 23257 5967
rect 25229 6151 25259 6182
rect 25961 6154 25991 6185
rect 26087 6154 26117 6185
rect 27173 6154 27203 6185
rect 27299 6154 27329 6185
rect 28385 6154 28415 6185
rect 28511 6154 28541 6185
rect 29597 6154 29627 6185
rect 29723 6154 29753 6185
rect 30372 6157 30402 6211
rect 30464 6157 30494 6183
rect 30560 6157 30590 6188
rect 25229 6039 25259 6067
rect 25961 6042 25991 6070
rect 26087 6042 26117 6070
rect 27173 6042 27203 6070
rect 27299 6042 27329 6070
rect 28385 6042 28415 6070
rect 28511 6042 28541 6070
rect 29597 6042 29627 6070
rect 29723 6042 29753 6070
rect 30372 6048 30402 6073
rect 30243 6028 30402 6048
rect 30464 6048 30494 6073
rect 30560 6048 30590 6073
rect 30464 6042 30590 6048
rect 30243 5994 30255 6028
rect 30289 5994 30402 6028
rect 23348 5925 23378 5957
rect 25582 5953 25612 5979
rect 26314 5953 26344 5979
rect 26436 5953 26466 5979
rect 27526 5953 27556 5979
rect 27648 5953 27678 5979
rect 28864 5953 28894 5979
rect 28986 5953 29016 5979
rect 29720 5953 29750 5979
rect 30243 5975 30402 5994
rect 30446 6026 30590 6042
rect 30758 6040 30788 6136
rect 30853 6040 30883 6072
rect 30937 6040 30967 6072
rect 30446 5992 30462 6026
rect 30496 5992 30590 6026
rect 30446 5976 30590 5992
rect 30372 5954 30402 5975
rect 30464 5969 30590 5976
rect 30706 6024 30788 6040
rect 30706 5990 30716 6024
rect 30750 5990 30788 6024
rect 30706 5974 30788 5990
rect 30830 6024 30967 6040
rect 30830 5990 30840 6024
rect 30874 5990 30967 6024
rect 30830 5974 30967 5990
rect 30464 5954 30494 5969
rect 30560 5954 30590 5969
rect 23043 5909 23257 5919
rect 23043 5875 23053 5909
rect 23087 5875 23257 5909
rect 23043 5865 23257 5875
rect 22580 5791 22610 5823
rect 22970 5791 23000 5863
rect 23043 5859 23095 5865
rect 23065 5837 23095 5859
rect 23227 5836 23257 5865
rect 23319 5909 23378 5925
rect 23319 5875 23329 5909
rect 23363 5875 23378 5909
rect 23319 5859 23378 5875
rect 30758 5906 30788 5974
rect 30853 5952 30883 5974
rect 30937 5952 30967 5974
rect 23348 5837 23378 5859
rect 24580 5841 24646 5857
rect 25582 5847 25612 5869
rect 26314 5847 26344 5869
rect 26436 5847 26466 5869
rect 27526 5847 27556 5869
rect 27648 5847 27678 5869
rect 28864 5847 28894 5869
rect 28986 5847 29016 5869
rect 29720 5847 29750 5869
rect 23227 5806 23283 5836
rect 23253 5791 23283 5806
rect 24580 5814 24596 5841
rect 24562 5807 24596 5814
rect 24630 5814 24646 5841
rect 25564 5831 25630 5847
rect 24630 5807 24664 5814
rect 24562 5784 24664 5807
rect 24562 5769 24592 5784
rect 24634 5769 24664 5784
rect 25564 5797 25580 5831
rect 25614 5797 25630 5831
rect 25564 5781 25630 5797
rect 26296 5831 26362 5847
rect 26296 5797 26312 5831
rect 26346 5797 26362 5831
rect 26296 5781 26362 5797
rect 26418 5831 26484 5847
rect 26418 5797 26434 5831
rect 26468 5797 26484 5831
rect 26418 5781 26484 5797
rect 27508 5831 27574 5847
rect 27508 5797 27524 5831
rect 27558 5797 27574 5831
rect 27508 5781 27574 5797
rect 27630 5831 27696 5847
rect 27630 5797 27646 5831
rect 27680 5797 27696 5831
rect 27630 5781 27696 5797
rect 28846 5831 28912 5847
rect 28846 5797 28862 5831
rect 28896 5797 28912 5831
rect 28846 5781 28912 5797
rect 28968 5831 29034 5847
rect 28968 5797 28984 5831
rect 29018 5797 29034 5831
rect 28968 5781 29034 5797
rect 29702 5831 29768 5847
rect 29702 5797 29718 5831
rect 29752 5797 29768 5831
rect 30372 5816 30402 5870
rect 30464 5844 30494 5870
rect 30560 5844 30590 5870
rect 29702 5781 29768 5797
rect 11576 5681 11606 5707
rect 11660 5681 11690 5707
rect 11848 5681 11878 5707
rect 11943 5681 11973 5707
rect 12049 5681 12079 5707
rect 12145 5681 12175 5707
rect 12255 5681 12285 5707
rect 12355 5681 12385 5707
rect 12439 5681 12469 5707
rect 12627 5681 12657 5707
rect 12722 5681 12752 5707
rect 12831 5681 12861 5707
rect 12926 5681 12956 5707
rect 13012 5681 13042 5707
rect 13130 5681 13160 5707
rect 13214 5681 13244 5707
rect 13402 5681 13432 5707
rect 13497 5681 13527 5707
rect 13685 5681 13715 5707
rect 13780 5681 13810 5707
rect 13968 5681 13998 5707
rect 14052 5681 14082 5707
rect 14240 5681 14270 5707
rect 14335 5681 14365 5707
rect 14441 5681 14471 5707
rect 14537 5681 14567 5707
rect 14647 5681 14677 5707
rect 14747 5681 14777 5707
rect 14831 5681 14861 5707
rect 15019 5681 15049 5707
rect 15114 5681 15144 5707
rect 15223 5681 15253 5707
rect 15318 5681 15348 5707
rect 15404 5681 15434 5707
rect 15522 5681 15552 5707
rect 15606 5681 15636 5707
rect 15794 5681 15824 5707
rect 15889 5681 15919 5707
rect 16077 5681 16107 5707
rect 16172 5681 16202 5707
rect 16360 5681 16390 5707
rect 16444 5681 16474 5707
rect 16632 5681 16662 5707
rect 16727 5681 16757 5707
rect 16833 5681 16863 5707
rect 16929 5681 16959 5707
rect 17039 5681 17069 5707
rect 17139 5681 17169 5707
rect 17223 5681 17253 5707
rect 17411 5681 17441 5707
rect 17506 5681 17536 5707
rect 17615 5681 17645 5707
rect 17710 5681 17740 5707
rect 17796 5681 17826 5707
rect 17914 5681 17944 5707
rect 17998 5681 18028 5707
rect 18186 5681 18216 5707
rect 18281 5681 18311 5707
rect 18469 5681 18499 5707
rect 18564 5681 18594 5707
rect 18752 5681 18782 5707
rect 18836 5681 18866 5707
rect 19024 5681 19054 5707
rect 19119 5681 19149 5707
rect 19225 5681 19255 5707
rect 19321 5681 19351 5707
rect 19431 5681 19461 5707
rect 19531 5681 19561 5707
rect 19615 5681 19645 5707
rect 19803 5681 19833 5707
rect 19898 5681 19928 5707
rect 20007 5681 20037 5707
rect 20102 5681 20132 5707
rect 20188 5681 20218 5707
rect 20306 5681 20336 5707
rect 20390 5681 20420 5707
rect 20578 5681 20608 5707
rect 20673 5681 20703 5707
rect 20861 5681 20891 5707
rect 20956 5681 20986 5707
rect 21144 5681 21174 5707
rect 21228 5681 21258 5707
rect 21416 5681 21446 5707
rect 21511 5681 21541 5707
rect 21617 5681 21647 5707
rect 21713 5681 21743 5707
rect 21823 5681 21853 5707
rect 21923 5681 21953 5707
rect 22007 5681 22037 5707
rect 22195 5681 22225 5707
rect 22290 5681 22320 5707
rect 22399 5681 22429 5707
rect 22494 5681 22524 5707
rect 22580 5681 22610 5707
rect 22698 5681 22728 5707
rect 22782 5681 22812 5707
rect 22970 5681 23000 5707
rect 23065 5681 23095 5707
rect 23253 5681 23283 5707
rect 23348 5681 23378 5707
rect 30758 5796 30788 5822
rect 30853 5796 30883 5822
rect 30937 5796 30967 5822
rect 30372 5705 30402 5732
rect 24562 5631 24592 5685
rect 24634 5631 24664 5685
rect 14695 5553 14761 5563
rect 14695 5519 14711 5553
rect 14745 5519 14761 5553
rect 17087 5553 17153 5563
rect 14695 5509 14761 5519
rect 17087 5519 17103 5553
rect 17137 5519 17153 5553
rect 19479 5553 19545 5563
rect 17087 5509 17153 5519
rect 19479 5519 19495 5553
rect 19529 5519 19545 5553
rect 21871 5553 21937 5563
rect 19479 5509 19545 5519
rect 21871 5519 21887 5553
rect 21921 5519 21937 5553
rect 21871 5509 21937 5519
rect 11136 5468 11166 5494
rect 11224 5468 11254 5494
rect 11412 5468 11442 5494
rect 11496 5468 11526 5494
rect 11580 5468 11610 5494
rect 11664 5468 11694 5494
rect 11748 5468 11778 5494
rect 11944 5468 11974 5494
rect 12028 5468 12058 5494
rect 12112 5468 12142 5494
rect 12196 5468 12226 5494
rect 12280 5468 12310 5494
rect 12364 5468 12394 5494
rect 12448 5468 12478 5494
rect 12532 5468 12562 5494
rect 12616 5468 12646 5494
rect 12700 5468 12730 5494
rect 12784 5468 12814 5494
rect 12868 5468 12898 5494
rect 12952 5468 12982 5494
rect 13036 5468 13066 5494
rect 13120 5468 13150 5494
rect 13204 5468 13234 5494
rect 13288 5468 13318 5494
rect 13372 5468 13402 5494
rect 13456 5468 13486 5494
rect 13540 5468 13570 5494
rect 13624 5468 13654 5494
rect 13708 5468 13738 5494
rect 13968 5468 13998 5494
rect 11136 5295 11166 5310
rect 11130 5271 11166 5295
rect 11130 5236 11160 5271
rect 11224 5249 11254 5310
rect 14063 5452 14093 5478
rect 14251 5468 14281 5494
rect 14546 5468 14576 5494
rect 14618 5468 14648 5494
rect 14714 5468 14744 5509
rect 14822 5468 14852 5494
rect 14940 5468 14970 5494
rect 15024 5468 15054 5494
rect 15168 5468 15198 5494
rect 15305 5468 15335 5494
rect 15389 5468 15419 5494
rect 15497 5468 15527 5494
rect 15603 5468 15633 5494
rect 15723 5468 15753 5494
rect 15807 5468 15837 5494
rect 15900 5468 15930 5494
rect 14063 5308 14093 5324
rect 14063 5278 14119 5308
rect 11084 5220 11160 5236
rect 11084 5186 11094 5220
rect 11128 5186 11160 5220
rect 11084 5170 11160 5186
rect 11202 5233 11256 5249
rect 11202 5199 11212 5233
rect 11246 5199 11256 5233
rect 11412 5232 11442 5268
rect 11202 5183 11256 5199
rect 11361 5220 11442 5232
rect 11496 5230 11526 5268
rect 11580 5230 11610 5268
rect 11664 5230 11694 5268
rect 11748 5230 11778 5268
rect 11361 5186 11377 5220
rect 11411 5186 11442 5220
rect 11130 5161 11160 5170
rect 11130 5137 11166 5161
rect 11136 5122 11166 5137
rect 11224 5122 11254 5183
rect 11361 5174 11442 5186
rect 11495 5220 11778 5230
rect 11495 5186 11511 5220
rect 11545 5186 11778 5220
rect 11495 5176 11778 5186
rect 11412 5148 11442 5174
rect 11496 5148 11526 5176
rect 11580 5148 11610 5176
rect 11664 5148 11694 5176
rect 11748 5148 11778 5176
rect 11944 5230 11974 5268
rect 12028 5230 12058 5268
rect 12112 5230 12142 5268
rect 12196 5230 12226 5268
rect 12280 5230 12310 5268
rect 12364 5230 12394 5268
rect 11944 5220 12394 5230
rect 11944 5186 11968 5220
rect 12002 5186 12036 5220
rect 12070 5186 12104 5220
rect 12138 5186 12172 5220
rect 12206 5186 12240 5220
rect 12274 5186 12308 5220
rect 12342 5186 12394 5220
rect 11944 5176 12394 5186
rect 11944 5148 11974 5176
rect 12028 5148 12058 5176
rect 12112 5148 12142 5176
rect 12196 5148 12226 5176
rect 12280 5148 12310 5176
rect 12364 5148 12394 5176
rect 12448 5230 12478 5268
rect 12532 5230 12562 5268
rect 12616 5230 12646 5268
rect 12700 5230 12730 5268
rect 12784 5230 12814 5268
rect 12868 5230 12898 5268
rect 12952 5230 12982 5268
rect 13036 5230 13066 5268
rect 13120 5230 13150 5268
rect 13204 5230 13234 5268
rect 13288 5230 13318 5268
rect 13372 5230 13402 5268
rect 13456 5230 13486 5268
rect 13540 5230 13570 5268
rect 13624 5230 13654 5268
rect 13708 5230 13738 5268
rect 13968 5236 13998 5268
rect 12448 5220 13742 5230
rect 12448 5186 12468 5220
rect 12502 5186 12536 5220
rect 12570 5186 12604 5220
rect 12638 5186 12672 5220
rect 12706 5186 12740 5220
rect 12774 5186 12808 5220
rect 12842 5186 12876 5220
rect 12910 5186 12944 5220
rect 12978 5186 13012 5220
rect 13046 5186 13080 5220
rect 13114 5186 13148 5220
rect 13182 5186 13216 5220
rect 13250 5186 13284 5220
rect 13318 5186 13352 5220
rect 13386 5186 13420 5220
rect 13454 5186 13488 5220
rect 13522 5186 13556 5220
rect 13590 5186 13624 5220
rect 13658 5186 13692 5220
rect 13726 5186 13742 5220
rect 12448 5176 13742 5186
rect 13968 5220 14027 5236
rect 13968 5186 13983 5220
rect 14017 5186 14027 5220
rect 12448 5148 12478 5176
rect 12532 5148 12562 5176
rect 12616 5148 12646 5176
rect 12700 5148 12730 5176
rect 12784 5148 12814 5176
rect 12868 5148 12898 5176
rect 12952 5148 12982 5176
rect 13036 5148 13066 5176
rect 13120 5148 13150 5176
rect 13204 5148 13234 5176
rect 13288 5148 13318 5176
rect 13372 5148 13402 5176
rect 13456 5148 13486 5176
rect 13540 5148 13570 5176
rect 13624 5148 13654 5176
rect 13708 5148 13738 5176
rect 13968 5170 14027 5186
rect 14089 5230 14119 5278
rect 14348 5400 14378 5426
rect 14251 5236 14281 5268
rect 14348 5240 14378 5272
rect 14546 5268 14576 5300
rect 14480 5252 14576 5268
rect 14251 5230 14303 5236
rect 14089 5220 14303 5230
rect 14089 5186 14259 5220
rect 14293 5186 14303 5220
rect 14089 5176 14303 5186
rect 13968 5148 13998 5170
rect 14089 5147 14119 5176
rect 14251 5170 14303 5176
rect 14345 5224 14409 5240
rect 14345 5190 14359 5224
rect 14393 5190 14409 5224
rect 14480 5218 14490 5252
rect 14524 5238 14576 5252
rect 14618 5252 14648 5300
rect 14524 5218 14564 5238
rect 14480 5202 14564 5218
rect 14345 5174 14409 5190
rect 14251 5148 14281 5170
rect 14063 5117 14119 5147
rect 14063 5102 14093 5117
rect 14346 5102 14376 5174
rect 14534 5146 14564 5202
rect 14618 5236 14672 5252
rect 14618 5202 14628 5236
rect 14662 5202 14672 5236
rect 14618 5186 14672 5202
rect 14714 5200 14744 5384
rect 14822 5352 14852 5384
rect 14786 5336 14852 5352
rect 14940 5346 14970 5384
rect 15024 5352 15054 5384
rect 14786 5302 14796 5336
rect 14830 5302 14852 5336
rect 14786 5286 14852 5302
rect 14916 5336 14982 5346
rect 14916 5302 14932 5336
rect 14966 5302 14982 5336
rect 14916 5292 14982 5302
rect 15024 5336 15078 5352
rect 15024 5302 15034 5336
rect 15068 5302 15078 5336
rect 14618 5146 14648 5186
rect 14714 5184 14780 5200
rect 14714 5150 14736 5184
rect 14770 5150 14780 5184
rect 14714 5134 14780 5150
rect 14736 5102 14766 5134
rect 14822 5102 14852 5286
rect 15024 5286 15078 5302
rect 16088 5462 16118 5488
rect 16172 5462 16202 5488
rect 16360 5468 16390 5494
rect 15024 5250 15054 5286
rect 14917 5220 15054 5250
rect 15168 5234 15198 5300
rect 15305 5268 15335 5300
rect 15389 5268 15419 5300
rect 14917 5090 14947 5220
rect 15121 5218 15198 5234
rect 15121 5184 15131 5218
rect 15165 5204 15198 5218
rect 15249 5252 15339 5268
rect 15249 5218 15259 5252
rect 15293 5218 15339 5252
rect 15165 5184 15175 5204
rect 15249 5202 15339 5218
rect 15389 5252 15455 5268
rect 15389 5218 15411 5252
rect 15445 5218 15455 5252
rect 15389 5202 15455 5218
rect 14989 5162 15056 5178
rect 14989 5128 14999 5162
rect 15033 5128 15056 5162
rect 15121 5168 15175 5184
rect 15121 5146 15151 5168
rect 15309 5146 15339 5202
rect 15393 5146 15423 5202
rect 15497 5200 15527 5384
rect 15603 5352 15633 5384
rect 15569 5336 15633 5352
rect 15723 5346 15753 5384
rect 15569 5302 15579 5336
rect 15613 5302 15633 5336
rect 15569 5286 15633 5302
rect 15699 5336 15765 5346
rect 15699 5302 15715 5336
rect 15749 5302 15765 5336
rect 15699 5292 15765 5302
rect 15497 5184 15557 5200
rect 15497 5164 15513 5184
rect 15493 5150 15513 5164
rect 15547 5150 15557 5184
rect 14989 5112 15056 5128
rect 15026 5090 15056 5112
rect 15493 5134 15557 5150
rect 15493 5102 15523 5134
rect 15603 5102 15633 5286
rect 15807 5250 15837 5384
rect 15699 5220 15837 5250
rect 15900 5238 15930 5384
rect 16088 5245 16118 5334
rect 16172 5319 16202 5334
rect 16172 5289 16235 5319
rect 16205 5251 16235 5289
rect 16455 5452 16485 5478
rect 16643 5468 16673 5494
rect 16938 5468 16968 5494
rect 17010 5468 17040 5494
rect 17106 5468 17136 5509
rect 17214 5468 17244 5494
rect 17332 5468 17362 5494
rect 17416 5468 17446 5494
rect 17560 5468 17590 5494
rect 17697 5468 17727 5494
rect 17781 5468 17811 5494
rect 17889 5468 17919 5494
rect 17995 5468 18025 5494
rect 18115 5468 18145 5494
rect 18199 5468 18229 5494
rect 18292 5468 18322 5494
rect 16455 5308 16485 5324
rect 16455 5278 16511 5308
rect 15887 5222 15941 5238
rect 15699 5190 15729 5220
rect 15675 5174 15729 5190
rect 15887 5188 15897 5222
rect 15931 5188 15941 5222
rect 15675 5140 15685 5174
rect 15719 5140 15729 5174
rect 15675 5124 15729 5140
rect 15699 5090 15729 5124
rect 15771 5162 15835 5178
rect 15887 5172 15941 5188
rect 16088 5235 16163 5245
rect 16088 5201 16113 5235
rect 16147 5201 16163 5235
rect 16088 5191 16163 5201
rect 16205 5235 16260 5251
rect 16205 5201 16215 5235
rect 16249 5201 16260 5235
rect 15771 5128 15781 5162
rect 15815 5128 15835 5162
rect 15771 5112 15835 5128
rect 15805 5090 15835 5112
rect 15900 5102 15930 5172
rect 16088 5102 16118 5191
rect 16205 5185 16260 5201
rect 16360 5236 16390 5268
rect 16360 5220 16419 5236
rect 16360 5186 16375 5220
rect 16409 5186 16419 5220
rect 16205 5147 16235 5185
rect 16360 5170 16419 5186
rect 16481 5230 16511 5278
rect 16740 5400 16770 5426
rect 16643 5236 16673 5268
rect 16740 5240 16770 5272
rect 16938 5268 16968 5300
rect 16872 5252 16968 5268
rect 16643 5230 16695 5236
rect 16481 5220 16695 5230
rect 16481 5186 16651 5220
rect 16685 5186 16695 5220
rect 16481 5176 16695 5186
rect 16360 5148 16390 5170
rect 16172 5117 16235 5147
rect 16172 5102 16202 5117
rect 16481 5147 16511 5176
rect 16643 5170 16695 5176
rect 16737 5224 16801 5240
rect 16737 5190 16751 5224
rect 16785 5190 16801 5224
rect 16872 5218 16882 5252
rect 16916 5238 16968 5252
rect 17010 5252 17040 5300
rect 16916 5218 16956 5238
rect 16872 5202 16956 5218
rect 16737 5174 16801 5190
rect 16643 5148 16673 5170
rect 16455 5117 16511 5147
rect 16455 5102 16485 5117
rect 16738 5102 16768 5174
rect 16926 5146 16956 5202
rect 17010 5236 17064 5252
rect 17010 5202 17020 5236
rect 17054 5202 17064 5236
rect 17010 5186 17064 5202
rect 17106 5200 17136 5384
rect 17214 5352 17244 5384
rect 17178 5336 17244 5352
rect 17332 5346 17362 5384
rect 17416 5352 17446 5384
rect 17178 5302 17188 5336
rect 17222 5302 17244 5336
rect 17178 5286 17244 5302
rect 17308 5336 17374 5346
rect 17308 5302 17324 5336
rect 17358 5302 17374 5336
rect 17308 5292 17374 5302
rect 17416 5336 17470 5352
rect 17416 5302 17426 5336
rect 17460 5302 17470 5336
rect 17010 5146 17040 5186
rect 17106 5184 17172 5200
rect 17106 5150 17128 5184
rect 17162 5150 17172 5184
rect 17106 5134 17172 5150
rect 17128 5102 17158 5134
rect 17214 5102 17244 5286
rect 17416 5286 17470 5302
rect 18480 5462 18510 5488
rect 18564 5462 18594 5488
rect 18752 5468 18782 5494
rect 17416 5250 17446 5286
rect 17309 5220 17446 5250
rect 17560 5234 17590 5300
rect 17697 5268 17727 5300
rect 17781 5268 17811 5300
rect 17309 5090 17339 5220
rect 17513 5218 17590 5234
rect 17513 5184 17523 5218
rect 17557 5204 17590 5218
rect 17641 5252 17731 5268
rect 17641 5218 17651 5252
rect 17685 5218 17731 5252
rect 17557 5184 17567 5204
rect 17641 5202 17731 5218
rect 17781 5252 17847 5268
rect 17781 5218 17803 5252
rect 17837 5218 17847 5252
rect 17781 5202 17847 5218
rect 17381 5162 17448 5178
rect 17381 5128 17391 5162
rect 17425 5128 17448 5162
rect 17513 5168 17567 5184
rect 17513 5146 17543 5168
rect 17701 5146 17731 5202
rect 17785 5146 17815 5202
rect 17889 5200 17919 5384
rect 17995 5352 18025 5384
rect 17961 5336 18025 5352
rect 18115 5346 18145 5384
rect 17961 5302 17971 5336
rect 18005 5302 18025 5336
rect 17961 5286 18025 5302
rect 18091 5336 18157 5346
rect 18091 5302 18107 5336
rect 18141 5302 18157 5336
rect 18091 5292 18157 5302
rect 17889 5184 17949 5200
rect 17889 5164 17905 5184
rect 17885 5150 17905 5164
rect 17939 5150 17949 5184
rect 17381 5112 17448 5128
rect 17418 5090 17448 5112
rect 17885 5134 17949 5150
rect 17885 5102 17915 5134
rect 17995 5102 18025 5286
rect 18199 5250 18229 5384
rect 18091 5220 18229 5250
rect 18292 5238 18322 5384
rect 18480 5245 18510 5334
rect 18564 5319 18594 5334
rect 18564 5289 18627 5319
rect 18597 5251 18627 5289
rect 18847 5452 18877 5478
rect 19035 5468 19065 5494
rect 19330 5468 19360 5494
rect 19402 5468 19432 5494
rect 19498 5468 19528 5509
rect 19606 5468 19636 5494
rect 19724 5468 19754 5494
rect 19808 5468 19838 5494
rect 19952 5468 19982 5494
rect 20089 5468 20119 5494
rect 20173 5468 20203 5494
rect 20281 5468 20311 5494
rect 20387 5468 20417 5494
rect 20507 5468 20537 5494
rect 20591 5468 20621 5494
rect 20684 5468 20714 5494
rect 18847 5308 18877 5324
rect 18847 5278 18903 5308
rect 18279 5222 18333 5238
rect 18091 5190 18121 5220
rect 18067 5174 18121 5190
rect 18279 5188 18289 5222
rect 18323 5188 18333 5222
rect 18067 5140 18077 5174
rect 18111 5140 18121 5174
rect 18067 5124 18121 5140
rect 18091 5090 18121 5124
rect 18163 5162 18227 5178
rect 18279 5172 18333 5188
rect 18480 5235 18555 5245
rect 18480 5201 18505 5235
rect 18539 5201 18555 5235
rect 18480 5191 18555 5201
rect 18597 5235 18652 5251
rect 18597 5201 18607 5235
rect 18641 5201 18652 5235
rect 18163 5128 18173 5162
rect 18207 5128 18227 5162
rect 18163 5112 18227 5128
rect 18197 5090 18227 5112
rect 18292 5102 18322 5172
rect 18480 5102 18510 5191
rect 18597 5185 18652 5201
rect 18752 5236 18782 5268
rect 18752 5220 18811 5236
rect 18752 5186 18767 5220
rect 18801 5186 18811 5220
rect 18597 5147 18627 5185
rect 18752 5170 18811 5186
rect 18873 5230 18903 5278
rect 19132 5400 19162 5426
rect 19035 5236 19065 5268
rect 19132 5240 19162 5272
rect 19330 5268 19360 5300
rect 19264 5252 19360 5268
rect 19035 5230 19087 5236
rect 18873 5220 19087 5230
rect 18873 5186 19043 5220
rect 19077 5186 19087 5220
rect 18873 5176 19087 5186
rect 18752 5148 18782 5170
rect 18564 5117 18627 5147
rect 18564 5102 18594 5117
rect 18873 5147 18903 5176
rect 19035 5170 19087 5176
rect 19129 5224 19193 5240
rect 19129 5190 19143 5224
rect 19177 5190 19193 5224
rect 19264 5218 19274 5252
rect 19308 5238 19360 5252
rect 19402 5252 19432 5300
rect 19308 5218 19348 5238
rect 19264 5202 19348 5218
rect 19129 5174 19193 5190
rect 19035 5148 19065 5170
rect 18847 5117 18903 5147
rect 18847 5102 18877 5117
rect 19130 5102 19160 5174
rect 19318 5146 19348 5202
rect 19402 5236 19456 5252
rect 19402 5202 19412 5236
rect 19446 5202 19456 5236
rect 19402 5186 19456 5202
rect 19498 5200 19528 5384
rect 19606 5352 19636 5384
rect 19570 5336 19636 5352
rect 19724 5346 19754 5384
rect 19808 5352 19838 5384
rect 19570 5302 19580 5336
rect 19614 5302 19636 5336
rect 19570 5286 19636 5302
rect 19700 5336 19766 5346
rect 19700 5302 19716 5336
rect 19750 5302 19766 5336
rect 19700 5292 19766 5302
rect 19808 5336 19862 5352
rect 19808 5302 19818 5336
rect 19852 5302 19862 5336
rect 19402 5146 19432 5186
rect 19498 5184 19564 5200
rect 19498 5150 19520 5184
rect 19554 5150 19564 5184
rect 19498 5134 19564 5150
rect 19520 5102 19550 5134
rect 19606 5102 19636 5286
rect 19808 5286 19862 5302
rect 20872 5462 20902 5488
rect 20956 5462 20986 5488
rect 21144 5468 21174 5494
rect 19808 5250 19838 5286
rect 19701 5220 19838 5250
rect 19952 5234 19982 5300
rect 20089 5268 20119 5300
rect 20173 5268 20203 5300
rect 19701 5090 19731 5220
rect 19905 5218 19982 5234
rect 19905 5184 19915 5218
rect 19949 5204 19982 5218
rect 20033 5252 20123 5268
rect 20033 5218 20043 5252
rect 20077 5218 20123 5252
rect 19949 5184 19959 5204
rect 20033 5202 20123 5218
rect 20173 5252 20239 5268
rect 20173 5218 20195 5252
rect 20229 5218 20239 5252
rect 20173 5202 20239 5218
rect 19773 5162 19840 5178
rect 19773 5128 19783 5162
rect 19817 5128 19840 5162
rect 19905 5168 19959 5184
rect 19905 5146 19935 5168
rect 20093 5146 20123 5202
rect 20177 5146 20207 5202
rect 20281 5200 20311 5384
rect 20387 5352 20417 5384
rect 20353 5336 20417 5352
rect 20507 5346 20537 5384
rect 20353 5302 20363 5336
rect 20397 5302 20417 5336
rect 20353 5286 20417 5302
rect 20483 5336 20549 5346
rect 20483 5302 20499 5336
rect 20533 5302 20549 5336
rect 20483 5292 20549 5302
rect 20281 5184 20341 5200
rect 20281 5164 20297 5184
rect 20277 5150 20297 5164
rect 20331 5150 20341 5184
rect 19773 5112 19840 5128
rect 19810 5090 19840 5112
rect 20277 5134 20341 5150
rect 20277 5102 20307 5134
rect 20387 5102 20417 5286
rect 20591 5250 20621 5384
rect 20483 5220 20621 5250
rect 20684 5238 20714 5384
rect 20872 5245 20902 5334
rect 20956 5319 20986 5334
rect 20956 5289 21019 5319
rect 20989 5251 21019 5289
rect 21239 5452 21269 5478
rect 21427 5468 21457 5494
rect 21722 5468 21752 5494
rect 21794 5468 21824 5494
rect 21890 5468 21920 5509
rect 21998 5468 22028 5494
rect 22116 5468 22146 5494
rect 22200 5468 22230 5494
rect 22344 5468 22374 5494
rect 22481 5468 22511 5494
rect 22565 5468 22595 5494
rect 22673 5468 22703 5494
rect 22779 5468 22809 5494
rect 22899 5468 22929 5494
rect 22983 5468 23013 5494
rect 23076 5468 23106 5494
rect 24562 5493 24592 5547
rect 24634 5493 24664 5547
rect 21239 5308 21269 5324
rect 21239 5278 21295 5308
rect 20671 5222 20725 5238
rect 20483 5190 20513 5220
rect 20459 5174 20513 5190
rect 20671 5188 20681 5222
rect 20715 5188 20725 5222
rect 20459 5140 20469 5174
rect 20503 5140 20513 5174
rect 20459 5124 20513 5140
rect 20483 5090 20513 5124
rect 20555 5162 20619 5178
rect 20671 5172 20725 5188
rect 20872 5235 20947 5245
rect 20872 5201 20897 5235
rect 20931 5201 20947 5235
rect 20872 5191 20947 5201
rect 20989 5235 21044 5251
rect 20989 5201 20999 5235
rect 21033 5201 21044 5235
rect 20555 5128 20565 5162
rect 20599 5128 20619 5162
rect 20555 5112 20619 5128
rect 20589 5090 20619 5112
rect 20684 5102 20714 5172
rect 20872 5102 20902 5191
rect 20989 5185 21044 5201
rect 21144 5236 21174 5268
rect 21144 5220 21203 5236
rect 21144 5186 21159 5220
rect 21193 5186 21203 5220
rect 20989 5147 21019 5185
rect 21144 5170 21203 5186
rect 21265 5230 21295 5278
rect 21524 5400 21554 5426
rect 21427 5236 21457 5268
rect 21524 5240 21554 5272
rect 21722 5268 21752 5300
rect 21656 5252 21752 5268
rect 21427 5230 21479 5236
rect 21265 5220 21479 5230
rect 21265 5186 21435 5220
rect 21469 5186 21479 5220
rect 21265 5176 21479 5186
rect 21144 5148 21174 5170
rect 20956 5117 21019 5147
rect 20956 5102 20986 5117
rect 21265 5147 21295 5176
rect 21427 5170 21479 5176
rect 21521 5224 21585 5240
rect 21521 5190 21535 5224
rect 21569 5190 21585 5224
rect 21656 5218 21666 5252
rect 21700 5238 21752 5252
rect 21794 5252 21824 5300
rect 21700 5218 21740 5238
rect 21656 5202 21740 5218
rect 21521 5174 21585 5190
rect 21427 5148 21457 5170
rect 21239 5117 21295 5147
rect 21239 5102 21269 5117
rect 21522 5102 21552 5174
rect 21710 5146 21740 5202
rect 21794 5236 21848 5252
rect 21794 5202 21804 5236
rect 21838 5202 21848 5236
rect 21794 5186 21848 5202
rect 21890 5200 21920 5384
rect 21998 5352 22028 5384
rect 21962 5336 22028 5352
rect 22116 5346 22146 5384
rect 22200 5352 22230 5384
rect 21962 5302 21972 5336
rect 22006 5302 22028 5336
rect 21962 5286 22028 5302
rect 22092 5336 22158 5346
rect 22092 5302 22108 5336
rect 22142 5302 22158 5336
rect 22092 5292 22158 5302
rect 22200 5336 22254 5352
rect 22200 5302 22210 5336
rect 22244 5302 22254 5336
rect 21794 5146 21824 5186
rect 21890 5184 21956 5200
rect 21890 5150 21912 5184
rect 21946 5150 21956 5184
rect 21890 5134 21956 5150
rect 21912 5102 21942 5134
rect 21998 5102 22028 5286
rect 22200 5286 22254 5302
rect 23264 5462 23294 5488
rect 23348 5462 23378 5488
rect 22200 5250 22230 5286
rect 22093 5220 22230 5250
rect 22344 5234 22374 5300
rect 22481 5268 22511 5300
rect 22565 5268 22595 5300
rect 22093 5090 22123 5220
rect 22297 5218 22374 5234
rect 22297 5184 22307 5218
rect 22341 5204 22374 5218
rect 22425 5252 22515 5268
rect 22425 5218 22435 5252
rect 22469 5218 22515 5252
rect 22341 5184 22351 5204
rect 22425 5202 22515 5218
rect 22565 5252 22631 5268
rect 22565 5218 22587 5252
rect 22621 5218 22631 5252
rect 22565 5202 22631 5218
rect 22165 5162 22232 5178
rect 22165 5128 22175 5162
rect 22209 5128 22232 5162
rect 22297 5168 22351 5184
rect 22297 5146 22327 5168
rect 22485 5146 22515 5202
rect 22569 5146 22599 5202
rect 22673 5200 22703 5384
rect 22779 5352 22809 5384
rect 22745 5336 22809 5352
rect 22899 5346 22929 5384
rect 22745 5302 22755 5336
rect 22789 5302 22809 5336
rect 22745 5286 22809 5302
rect 22875 5336 22941 5346
rect 22875 5302 22891 5336
rect 22925 5302 22941 5336
rect 22875 5292 22941 5302
rect 22673 5184 22733 5200
rect 22673 5164 22689 5184
rect 22669 5150 22689 5164
rect 22723 5150 22733 5184
rect 22165 5112 22232 5128
rect 22202 5090 22232 5112
rect 22669 5134 22733 5150
rect 22669 5102 22699 5134
rect 22779 5102 22809 5286
rect 22983 5250 23013 5384
rect 22875 5220 23013 5250
rect 23076 5238 23106 5384
rect 24562 5355 24592 5409
rect 24634 5355 24664 5409
rect 23264 5245 23294 5334
rect 23348 5319 23378 5334
rect 23348 5289 23411 5319
rect 23381 5251 23411 5289
rect 23063 5222 23117 5238
rect 22875 5190 22905 5220
rect 22851 5174 22905 5190
rect 23063 5188 23073 5222
rect 23107 5188 23117 5222
rect 22851 5140 22861 5174
rect 22895 5140 22905 5174
rect 22851 5124 22905 5140
rect 22875 5090 22905 5124
rect 22947 5162 23011 5178
rect 23063 5172 23117 5188
rect 23264 5235 23339 5245
rect 23264 5201 23289 5235
rect 23323 5201 23339 5235
rect 23264 5191 23339 5201
rect 23381 5235 23436 5251
rect 23381 5201 23391 5235
rect 23425 5201 23436 5235
rect 24562 5217 24592 5271
rect 24634 5217 24664 5271
rect 22947 5128 22957 5162
rect 22991 5128 23011 5162
rect 22947 5112 23011 5128
rect 22981 5090 23011 5112
rect 23076 5102 23106 5172
rect 23264 5102 23294 5191
rect 23381 5185 23436 5201
rect 23381 5147 23411 5185
rect 23348 5117 23411 5147
rect 23348 5102 23378 5117
rect 24562 5079 24592 5133
rect 24634 5079 24664 5133
rect 11136 4992 11166 5018
rect 11224 4992 11254 5018
rect 11412 4992 11442 5018
rect 11496 4992 11526 5018
rect 11580 4992 11610 5018
rect 11664 4992 11694 5018
rect 11748 4992 11778 5018
rect 11944 4992 11974 5018
rect 12028 4992 12058 5018
rect 12112 4992 12142 5018
rect 12196 4992 12226 5018
rect 12280 4992 12310 5018
rect 12364 4992 12394 5018
rect 12448 4992 12478 5018
rect 12532 4992 12562 5018
rect 12616 4992 12646 5018
rect 12700 4992 12730 5018
rect 12784 4992 12814 5018
rect 12868 4992 12898 5018
rect 12952 4992 12982 5018
rect 13036 4992 13066 5018
rect 13120 4992 13150 5018
rect 13204 4992 13234 5018
rect 13288 4992 13318 5018
rect 13372 4992 13402 5018
rect 13456 4992 13486 5018
rect 13540 4992 13570 5018
rect 13624 4992 13654 5018
rect 13708 4992 13738 5018
rect 13968 4992 13998 5018
rect 14063 4992 14093 5018
rect 14251 4992 14281 5018
rect 14346 4992 14376 5018
rect 14534 4992 14564 5018
rect 14618 4992 14648 5018
rect 14736 4992 14766 5018
rect 14822 4992 14852 5018
rect 14917 4992 14947 5018
rect 15026 4992 15056 5018
rect 15121 4992 15151 5018
rect 15309 4992 15339 5018
rect 15393 4992 15423 5018
rect 15493 4992 15523 5018
rect 15603 4992 15633 5018
rect 15699 4992 15729 5018
rect 15805 4992 15835 5018
rect 15900 4992 15930 5018
rect 16088 4992 16118 5018
rect 16172 4992 16202 5018
rect 16360 4992 16390 5018
rect 16455 4992 16485 5018
rect 16643 4992 16673 5018
rect 16738 4992 16768 5018
rect 16926 4992 16956 5018
rect 17010 4992 17040 5018
rect 17128 4992 17158 5018
rect 17214 4992 17244 5018
rect 17309 4992 17339 5018
rect 17418 4992 17448 5018
rect 17513 4992 17543 5018
rect 17701 4992 17731 5018
rect 17785 4992 17815 5018
rect 17885 4992 17915 5018
rect 17995 4992 18025 5018
rect 18091 4992 18121 5018
rect 18197 4992 18227 5018
rect 18292 4992 18322 5018
rect 18480 4992 18510 5018
rect 18564 4992 18594 5018
rect 18752 4992 18782 5018
rect 18847 4992 18877 5018
rect 19035 4992 19065 5018
rect 19130 4992 19160 5018
rect 19318 4992 19348 5018
rect 19402 4992 19432 5018
rect 19520 4992 19550 5018
rect 19606 4992 19636 5018
rect 19701 4992 19731 5018
rect 19810 4992 19840 5018
rect 19905 4992 19935 5018
rect 20093 4992 20123 5018
rect 20177 4992 20207 5018
rect 20277 4992 20307 5018
rect 20387 4992 20417 5018
rect 20483 4992 20513 5018
rect 20589 4992 20619 5018
rect 20684 4992 20714 5018
rect 20872 4992 20902 5018
rect 20956 4992 20986 5018
rect 21144 4992 21174 5018
rect 21239 4992 21269 5018
rect 21427 4992 21457 5018
rect 21522 4992 21552 5018
rect 21710 4992 21740 5018
rect 21794 4992 21824 5018
rect 21912 4992 21942 5018
rect 21998 4992 22028 5018
rect 22093 4992 22123 5018
rect 22202 4992 22232 5018
rect 22297 4992 22327 5018
rect 22485 4992 22515 5018
rect 22569 4992 22599 5018
rect 22669 4992 22699 5018
rect 22779 4992 22809 5018
rect 22875 4992 22905 5018
rect 22981 4992 23011 5018
rect 23076 4992 23106 5018
rect 23264 4992 23294 5018
rect 23348 4992 23378 5018
rect 24562 4941 24592 4995
rect 24634 4941 24664 4995
rect 24562 4803 24592 4857
rect 24634 4803 24664 4857
rect 24562 4693 24592 4719
rect 24634 4693 24664 4719
rect 11168 4594 11198 4620
rect 11256 4594 11286 4620
rect 11444 4594 11474 4620
rect 11528 4594 11558 4620
rect 11612 4594 11642 4620
rect 11696 4594 11726 4620
rect 11780 4594 11810 4620
rect 13751 4595 13781 4621
rect 11168 4421 11198 4436
rect 11162 4397 11198 4421
rect 11162 4362 11192 4397
rect 11256 4375 11286 4436
rect 13967 4589 13997 4615
rect 14051 4589 14081 4615
rect 14239 4595 14269 4621
rect 14332 4595 14362 4621
rect 14416 4595 14446 4621
rect 14536 4595 14566 4621
rect 14642 4595 14672 4621
rect 14750 4595 14780 4621
rect 14834 4595 14864 4621
rect 14971 4595 15001 4621
rect 15115 4595 15145 4621
rect 15199 4595 15229 4621
rect 15317 4595 15347 4621
rect 15425 4595 15455 4621
rect 15521 4595 15551 4621
rect 15593 4595 15623 4621
rect 15888 4595 15918 4621
rect 13967 4446 13997 4461
rect 13934 4416 13997 4446
rect 11116 4346 11192 4362
rect 11116 4312 11126 4346
rect 11160 4312 11192 4346
rect 11116 4296 11192 4312
rect 11234 4359 11288 4375
rect 11234 4325 11244 4359
rect 11278 4325 11288 4359
rect 11444 4358 11474 4394
rect 11234 4309 11288 4325
rect 11393 4346 11474 4358
rect 11528 4356 11558 4394
rect 11612 4356 11642 4394
rect 11696 4356 11726 4394
rect 11780 4356 11810 4394
rect 13751 4363 13781 4395
rect 13934 4378 13964 4416
rect 11393 4312 11409 4346
rect 11443 4312 11474 4346
rect 11162 4287 11192 4296
rect 11162 4263 11198 4287
rect 11168 4248 11198 4263
rect 11256 4248 11286 4309
rect 11393 4300 11474 4312
rect 11527 4346 11810 4356
rect 11527 4312 11543 4346
rect 11577 4312 11810 4346
rect 11527 4302 11810 4312
rect 11444 4274 11474 4300
rect 11528 4274 11558 4302
rect 11612 4274 11642 4302
rect 11696 4274 11726 4302
rect 11780 4274 11810 4302
rect 13695 4347 13781 4363
rect 13695 4313 13711 4347
rect 13745 4313 13781 4347
rect 13695 4297 13781 4313
rect 13909 4362 13964 4378
rect 14051 4372 14081 4461
rect 13909 4328 13920 4362
rect 13954 4328 13964 4362
rect 13909 4312 13964 4328
rect 14006 4362 14081 4372
rect 14239 4365 14269 4511
rect 14332 4377 14362 4511
rect 14416 4473 14446 4511
rect 14536 4479 14566 4511
rect 14404 4463 14470 4473
rect 14404 4429 14420 4463
rect 14454 4429 14470 4463
rect 14404 4419 14470 4429
rect 14536 4463 14600 4479
rect 14536 4429 14556 4463
rect 14590 4429 14600 4463
rect 14536 4413 14600 4429
rect 14006 4328 14022 4362
rect 14056 4328 14081 4362
rect 14006 4318 14081 4328
rect 13751 4275 13781 4297
rect 13934 4274 13964 4312
rect 13934 4244 13997 4274
rect 13967 4229 13997 4244
rect 14051 4229 14081 4318
rect 14228 4349 14282 4365
rect 14228 4315 14238 4349
rect 14272 4315 14282 4349
rect 14332 4347 14470 4377
rect 14228 4299 14282 4315
rect 14440 4317 14470 4347
rect 14239 4229 14269 4299
rect 14334 4289 14398 4305
rect 14334 4255 14354 4289
rect 14388 4255 14398 4289
rect 14334 4239 14398 4255
rect 14440 4301 14494 4317
rect 14440 4267 14450 4301
rect 14484 4267 14494 4301
rect 14440 4251 14494 4267
rect 14334 4217 14364 4239
rect 14440 4217 14470 4251
rect 14536 4229 14566 4413
rect 14642 4327 14672 4511
rect 15115 4479 15145 4511
rect 15091 4463 15145 4479
rect 15199 4473 15229 4511
rect 15317 4479 15347 4511
rect 15091 4429 15101 4463
rect 15135 4429 15145 4463
rect 14750 4395 14780 4427
rect 14834 4395 14864 4427
rect 14714 4379 14780 4395
rect 14714 4345 14724 4379
rect 14758 4345 14780 4379
rect 14714 4329 14780 4345
rect 14830 4379 14920 4395
rect 14830 4345 14876 4379
rect 14910 4345 14920 4379
rect 14830 4329 14920 4345
rect 14971 4361 15001 4427
rect 15091 4413 15145 4429
rect 15187 4463 15253 4473
rect 15187 4429 15203 4463
rect 15237 4429 15253 4463
rect 15187 4419 15253 4429
rect 15317 4463 15383 4479
rect 15317 4429 15339 4463
rect 15373 4429 15383 4463
rect 15115 4377 15145 4413
rect 15317 4413 15383 4429
rect 14971 4345 15048 4361
rect 15115 4347 15252 4377
rect 14971 4331 15004 4345
rect 14612 4311 14672 4327
rect 14612 4277 14622 4311
rect 14656 4291 14672 4311
rect 14656 4277 14676 4291
rect 14612 4261 14676 4277
rect 14746 4273 14776 4329
rect 14830 4273 14860 4329
rect 14994 4311 15004 4331
rect 15038 4311 15048 4345
rect 14994 4295 15048 4311
rect 15018 4273 15048 4295
rect 15113 4289 15180 4305
rect 14646 4229 14676 4261
rect 15113 4255 15136 4289
rect 15170 4255 15180 4289
rect 15113 4239 15180 4255
rect 15113 4217 15143 4239
rect 15222 4217 15252 4347
rect 15317 4229 15347 4413
rect 15425 4327 15455 4511
rect 15791 4527 15821 4553
rect 15521 4379 15551 4427
rect 15389 4311 15455 4327
rect 15497 4363 15551 4379
rect 15593 4395 15623 4427
rect 15593 4379 15689 4395
rect 15593 4365 15645 4379
rect 15497 4329 15507 4363
rect 15541 4329 15551 4363
rect 15497 4313 15551 4329
rect 15389 4277 15399 4311
rect 15433 4277 15455 4311
rect 15389 4261 15455 4277
rect 15521 4273 15551 4313
rect 15605 4345 15645 4365
rect 15679 4345 15689 4379
rect 15791 4367 15821 4399
rect 16076 4579 16106 4605
rect 16171 4595 16201 4621
rect 16076 4435 16106 4451
rect 16050 4405 16106 4435
rect 15605 4329 15689 4345
rect 15760 4351 15824 4367
rect 15888 4363 15918 4395
rect 15605 4273 15635 4329
rect 15760 4317 15776 4351
rect 15810 4317 15824 4351
rect 15760 4301 15824 4317
rect 15866 4357 15918 4363
rect 16050 4357 16080 4405
rect 16359 4589 16389 4615
rect 16443 4589 16473 4615
rect 16631 4595 16661 4621
rect 16724 4595 16754 4621
rect 16808 4595 16838 4621
rect 16928 4595 16958 4621
rect 17034 4595 17064 4621
rect 17142 4595 17172 4621
rect 17226 4595 17256 4621
rect 17363 4595 17393 4621
rect 17507 4595 17537 4621
rect 17591 4595 17621 4621
rect 17709 4595 17739 4621
rect 17817 4595 17847 4621
rect 17913 4595 17943 4621
rect 17985 4595 18015 4621
rect 18280 4595 18310 4621
rect 16359 4446 16389 4461
rect 16326 4416 16389 4446
rect 16171 4363 16201 4395
rect 16326 4378 16356 4416
rect 15866 4347 16080 4357
rect 15866 4313 15876 4347
rect 15910 4313 16080 4347
rect 15866 4303 16080 4313
rect 15403 4229 15433 4261
rect 15793 4229 15823 4301
rect 15866 4297 15918 4303
rect 15888 4275 15918 4297
rect 16050 4274 16080 4303
rect 16142 4347 16201 4363
rect 16142 4313 16152 4347
rect 16186 4313 16201 4347
rect 16142 4297 16201 4313
rect 16301 4362 16356 4378
rect 16443 4372 16473 4461
rect 16301 4328 16312 4362
rect 16346 4328 16356 4362
rect 16301 4312 16356 4328
rect 16398 4362 16473 4372
rect 16631 4365 16661 4511
rect 16724 4377 16754 4511
rect 16808 4473 16838 4511
rect 16928 4479 16958 4511
rect 16796 4463 16862 4473
rect 16796 4429 16812 4463
rect 16846 4429 16862 4463
rect 16796 4419 16862 4429
rect 16928 4463 16992 4479
rect 16928 4429 16948 4463
rect 16982 4429 16992 4463
rect 16928 4413 16992 4429
rect 16398 4328 16414 4362
rect 16448 4328 16473 4362
rect 16398 4318 16473 4328
rect 16171 4275 16201 4297
rect 16050 4244 16106 4274
rect 16076 4229 16106 4244
rect 16326 4274 16356 4312
rect 16326 4244 16389 4274
rect 16359 4229 16389 4244
rect 16443 4229 16473 4318
rect 16620 4349 16674 4365
rect 16620 4315 16630 4349
rect 16664 4315 16674 4349
rect 16724 4347 16862 4377
rect 16620 4299 16674 4315
rect 16832 4317 16862 4347
rect 16631 4229 16661 4299
rect 16726 4289 16790 4305
rect 16726 4255 16746 4289
rect 16780 4255 16790 4289
rect 16726 4239 16790 4255
rect 16832 4301 16886 4317
rect 16832 4267 16842 4301
rect 16876 4267 16886 4301
rect 16832 4251 16886 4267
rect 16726 4217 16756 4239
rect 16832 4217 16862 4251
rect 16928 4229 16958 4413
rect 17034 4327 17064 4511
rect 17507 4479 17537 4511
rect 17483 4463 17537 4479
rect 17591 4473 17621 4511
rect 17709 4479 17739 4511
rect 17483 4429 17493 4463
rect 17527 4429 17537 4463
rect 17142 4395 17172 4427
rect 17226 4395 17256 4427
rect 17106 4379 17172 4395
rect 17106 4345 17116 4379
rect 17150 4345 17172 4379
rect 17106 4329 17172 4345
rect 17222 4379 17312 4395
rect 17222 4345 17268 4379
rect 17302 4345 17312 4379
rect 17222 4329 17312 4345
rect 17363 4361 17393 4427
rect 17483 4413 17537 4429
rect 17579 4463 17645 4473
rect 17579 4429 17595 4463
rect 17629 4429 17645 4463
rect 17579 4419 17645 4429
rect 17709 4463 17775 4479
rect 17709 4429 17731 4463
rect 17765 4429 17775 4463
rect 17507 4377 17537 4413
rect 17709 4413 17775 4429
rect 17363 4345 17440 4361
rect 17507 4347 17644 4377
rect 17363 4331 17396 4345
rect 17004 4311 17064 4327
rect 17004 4277 17014 4311
rect 17048 4291 17064 4311
rect 17048 4277 17068 4291
rect 17004 4261 17068 4277
rect 17138 4273 17168 4329
rect 17222 4273 17252 4329
rect 17386 4311 17396 4331
rect 17430 4311 17440 4345
rect 17386 4295 17440 4311
rect 17410 4273 17440 4295
rect 17505 4289 17572 4305
rect 17038 4229 17068 4261
rect 17505 4255 17528 4289
rect 17562 4255 17572 4289
rect 17505 4239 17572 4255
rect 17505 4217 17535 4239
rect 17614 4217 17644 4347
rect 17709 4229 17739 4413
rect 17817 4327 17847 4511
rect 18183 4527 18213 4553
rect 17913 4379 17943 4427
rect 17781 4311 17847 4327
rect 17889 4363 17943 4379
rect 17985 4395 18015 4427
rect 17985 4379 18081 4395
rect 17985 4365 18037 4379
rect 17889 4329 17899 4363
rect 17933 4329 17943 4363
rect 17889 4313 17943 4329
rect 17781 4277 17791 4311
rect 17825 4277 17847 4311
rect 17781 4261 17847 4277
rect 17913 4273 17943 4313
rect 17997 4345 18037 4365
rect 18071 4345 18081 4379
rect 18183 4367 18213 4399
rect 18468 4579 18498 4605
rect 18563 4595 18593 4621
rect 18468 4435 18498 4451
rect 18442 4405 18498 4435
rect 17997 4329 18081 4345
rect 18152 4351 18216 4367
rect 18280 4363 18310 4395
rect 17997 4273 18027 4329
rect 18152 4317 18168 4351
rect 18202 4317 18216 4351
rect 18152 4301 18216 4317
rect 18258 4357 18310 4363
rect 18442 4357 18472 4405
rect 18751 4589 18781 4615
rect 18835 4589 18865 4615
rect 19023 4595 19053 4621
rect 19116 4595 19146 4621
rect 19200 4595 19230 4621
rect 19320 4595 19350 4621
rect 19426 4595 19456 4621
rect 19534 4595 19564 4621
rect 19618 4595 19648 4621
rect 19755 4595 19785 4621
rect 19899 4595 19929 4621
rect 19983 4595 20013 4621
rect 20101 4595 20131 4621
rect 20209 4595 20239 4621
rect 20305 4595 20335 4621
rect 20377 4595 20407 4621
rect 20672 4595 20702 4621
rect 18751 4446 18781 4461
rect 18718 4416 18781 4446
rect 18563 4363 18593 4395
rect 18718 4378 18748 4416
rect 18258 4347 18472 4357
rect 18258 4313 18268 4347
rect 18302 4313 18472 4347
rect 18258 4303 18472 4313
rect 17795 4229 17825 4261
rect 18185 4229 18215 4301
rect 18258 4297 18310 4303
rect 18280 4275 18310 4297
rect 18442 4274 18472 4303
rect 18534 4347 18593 4363
rect 18534 4313 18544 4347
rect 18578 4313 18593 4347
rect 18534 4297 18593 4313
rect 18693 4362 18748 4378
rect 18835 4372 18865 4461
rect 18693 4328 18704 4362
rect 18738 4328 18748 4362
rect 18693 4312 18748 4328
rect 18790 4362 18865 4372
rect 19023 4365 19053 4511
rect 19116 4377 19146 4511
rect 19200 4473 19230 4511
rect 19320 4479 19350 4511
rect 19188 4463 19254 4473
rect 19188 4429 19204 4463
rect 19238 4429 19254 4463
rect 19188 4419 19254 4429
rect 19320 4463 19384 4479
rect 19320 4429 19340 4463
rect 19374 4429 19384 4463
rect 19320 4413 19384 4429
rect 18790 4328 18806 4362
rect 18840 4328 18865 4362
rect 18790 4318 18865 4328
rect 18563 4275 18593 4297
rect 18442 4244 18498 4274
rect 18468 4229 18498 4244
rect 18718 4274 18748 4312
rect 18718 4244 18781 4274
rect 18751 4229 18781 4244
rect 18835 4229 18865 4318
rect 19012 4349 19066 4365
rect 19012 4315 19022 4349
rect 19056 4315 19066 4349
rect 19116 4347 19254 4377
rect 19012 4299 19066 4315
rect 19224 4317 19254 4347
rect 19023 4229 19053 4299
rect 19118 4289 19182 4305
rect 19118 4255 19138 4289
rect 19172 4255 19182 4289
rect 19118 4239 19182 4255
rect 19224 4301 19278 4317
rect 19224 4267 19234 4301
rect 19268 4267 19278 4301
rect 19224 4251 19278 4267
rect 19118 4217 19148 4239
rect 19224 4217 19254 4251
rect 19320 4229 19350 4413
rect 19426 4327 19456 4511
rect 19899 4479 19929 4511
rect 19875 4463 19929 4479
rect 19983 4473 20013 4511
rect 20101 4479 20131 4511
rect 19875 4429 19885 4463
rect 19919 4429 19929 4463
rect 19534 4395 19564 4427
rect 19618 4395 19648 4427
rect 19498 4379 19564 4395
rect 19498 4345 19508 4379
rect 19542 4345 19564 4379
rect 19498 4329 19564 4345
rect 19614 4379 19704 4395
rect 19614 4345 19660 4379
rect 19694 4345 19704 4379
rect 19614 4329 19704 4345
rect 19755 4361 19785 4427
rect 19875 4413 19929 4429
rect 19971 4463 20037 4473
rect 19971 4429 19987 4463
rect 20021 4429 20037 4463
rect 19971 4419 20037 4429
rect 20101 4463 20167 4479
rect 20101 4429 20123 4463
rect 20157 4429 20167 4463
rect 19899 4377 19929 4413
rect 20101 4413 20167 4429
rect 19755 4345 19832 4361
rect 19899 4347 20036 4377
rect 19755 4331 19788 4345
rect 19396 4311 19456 4327
rect 19396 4277 19406 4311
rect 19440 4291 19456 4311
rect 19440 4277 19460 4291
rect 19396 4261 19460 4277
rect 19530 4273 19560 4329
rect 19614 4273 19644 4329
rect 19778 4311 19788 4331
rect 19822 4311 19832 4345
rect 19778 4295 19832 4311
rect 19802 4273 19832 4295
rect 19897 4289 19964 4305
rect 19430 4229 19460 4261
rect 19897 4255 19920 4289
rect 19954 4255 19964 4289
rect 19897 4239 19964 4255
rect 19897 4217 19927 4239
rect 20006 4217 20036 4347
rect 20101 4229 20131 4413
rect 20209 4327 20239 4511
rect 20575 4527 20605 4553
rect 20305 4379 20335 4427
rect 20173 4311 20239 4327
rect 20281 4363 20335 4379
rect 20377 4395 20407 4427
rect 20377 4379 20473 4395
rect 20377 4365 20429 4379
rect 20281 4329 20291 4363
rect 20325 4329 20335 4363
rect 20281 4313 20335 4329
rect 20173 4277 20183 4311
rect 20217 4277 20239 4311
rect 20173 4261 20239 4277
rect 20305 4273 20335 4313
rect 20389 4345 20429 4365
rect 20463 4345 20473 4379
rect 20575 4367 20605 4399
rect 20860 4579 20890 4605
rect 20955 4595 20985 4621
rect 20860 4435 20890 4451
rect 20834 4405 20890 4435
rect 20389 4329 20473 4345
rect 20544 4351 20608 4367
rect 20672 4363 20702 4395
rect 20389 4273 20419 4329
rect 20544 4317 20560 4351
rect 20594 4317 20608 4351
rect 20544 4301 20608 4317
rect 20650 4357 20702 4363
rect 20834 4357 20864 4405
rect 21143 4589 21173 4615
rect 21227 4589 21257 4615
rect 21415 4595 21445 4621
rect 21508 4595 21538 4621
rect 21592 4595 21622 4621
rect 21712 4595 21742 4621
rect 21818 4595 21848 4621
rect 21926 4595 21956 4621
rect 22010 4595 22040 4621
rect 22147 4595 22177 4621
rect 22291 4595 22321 4621
rect 22375 4595 22405 4621
rect 22493 4595 22523 4621
rect 22601 4595 22631 4621
rect 22697 4595 22727 4621
rect 22769 4595 22799 4621
rect 23064 4595 23094 4621
rect 21143 4446 21173 4461
rect 21110 4416 21173 4446
rect 20955 4363 20985 4395
rect 21110 4378 21140 4416
rect 20650 4347 20864 4357
rect 20650 4313 20660 4347
rect 20694 4313 20864 4347
rect 20650 4303 20864 4313
rect 20187 4229 20217 4261
rect 20577 4229 20607 4301
rect 20650 4297 20702 4303
rect 20672 4275 20702 4297
rect 20834 4274 20864 4303
rect 20926 4347 20985 4363
rect 20926 4313 20936 4347
rect 20970 4313 20985 4347
rect 20926 4297 20985 4313
rect 21085 4362 21140 4378
rect 21227 4372 21257 4461
rect 21085 4328 21096 4362
rect 21130 4328 21140 4362
rect 21085 4312 21140 4328
rect 21182 4362 21257 4372
rect 21415 4365 21445 4511
rect 21508 4377 21538 4511
rect 21592 4473 21622 4511
rect 21712 4479 21742 4511
rect 21580 4463 21646 4473
rect 21580 4429 21596 4463
rect 21630 4429 21646 4463
rect 21580 4419 21646 4429
rect 21712 4463 21776 4479
rect 21712 4429 21732 4463
rect 21766 4429 21776 4463
rect 21712 4413 21776 4429
rect 21182 4328 21198 4362
rect 21232 4328 21257 4362
rect 21182 4318 21257 4328
rect 20955 4275 20985 4297
rect 20834 4244 20890 4274
rect 20860 4229 20890 4244
rect 21110 4274 21140 4312
rect 21110 4244 21173 4274
rect 21143 4229 21173 4244
rect 21227 4229 21257 4318
rect 21404 4349 21458 4365
rect 21404 4315 21414 4349
rect 21448 4315 21458 4349
rect 21508 4347 21646 4377
rect 21404 4299 21458 4315
rect 21616 4317 21646 4347
rect 21415 4229 21445 4299
rect 21510 4289 21574 4305
rect 21510 4255 21530 4289
rect 21564 4255 21574 4289
rect 21510 4239 21574 4255
rect 21616 4301 21670 4317
rect 21616 4267 21626 4301
rect 21660 4267 21670 4301
rect 21616 4251 21670 4267
rect 21510 4217 21540 4239
rect 21616 4217 21646 4251
rect 21712 4229 21742 4413
rect 21818 4327 21848 4511
rect 22291 4479 22321 4511
rect 22267 4463 22321 4479
rect 22375 4473 22405 4511
rect 22493 4479 22523 4511
rect 22267 4429 22277 4463
rect 22311 4429 22321 4463
rect 21926 4395 21956 4427
rect 22010 4395 22040 4427
rect 21890 4379 21956 4395
rect 21890 4345 21900 4379
rect 21934 4345 21956 4379
rect 21890 4329 21956 4345
rect 22006 4379 22096 4395
rect 22006 4345 22052 4379
rect 22086 4345 22096 4379
rect 22006 4329 22096 4345
rect 22147 4361 22177 4427
rect 22267 4413 22321 4429
rect 22363 4463 22429 4473
rect 22363 4429 22379 4463
rect 22413 4429 22429 4463
rect 22363 4419 22429 4429
rect 22493 4463 22559 4479
rect 22493 4429 22515 4463
rect 22549 4429 22559 4463
rect 22291 4377 22321 4413
rect 22493 4413 22559 4429
rect 22147 4345 22224 4361
rect 22291 4347 22428 4377
rect 22147 4331 22180 4345
rect 21788 4311 21848 4327
rect 21788 4277 21798 4311
rect 21832 4291 21848 4311
rect 21832 4277 21852 4291
rect 21788 4261 21852 4277
rect 21922 4273 21952 4329
rect 22006 4273 22036 4329
rect 22170 4311 22180 4331
rect 22214 4311 22224 4345
rect 22170 4295 22224 4311
rect 22194 4273 22224 4295
rect 22289 4289 22356 4305
rect 21822 4229 21852 4261
rect 22289 4255 22312 4289
rect 22346 4255 22356 4289
rect 22289 4239 22356 4255
rect 22289 4217 22319 4239
rect 22398 4217 22428 4347
rect 22493 4229 22523 4413
rect 22601 4327 22631 4511
rect 22967 4527 22997 4553
rect 22697 4379 22727 4427
rect 22565 4311 22631 4327
rect 22673 4363 22727 4379
rect 22769 4395 22799 4427
rect 22769 4379 22865 4395
rect 22769 4365 22821 4379
rect 22673 4329 22683 4363
rect 22717 4329 22727 4363
rect 22673 4313 22727 4329
rect 22565 4277 22575 4311
rect 22609 4277 22631 4311
rect 22565 4261 22631 4277
rect 22697 4273 22727 4313
rect 22781 4345 22821 4365
rect 22855 4345 22865 4379
rect 22967 4367 22997 4399
rect 23252 4579 23282 4605
rect 23347 4595 23377 4621
rect 23252 4435 23282 4451
rect 23226 4405 23282 4435
rect 22781 4329 22865 4345
rect 22936 4351 23000 4367
rect 23064 4363 23094 4395
rect 22781 4273 22811 4329
rect 22936 4317 22952 4351
rect 22986 4317 23000 4351
rect 22936 4301 23000 4317
rect 23042 4357 23094 4363
rect 23226 4357 23256 4405
rect 23347 4363 23377 4395
rect 23042 4347 23256 4357
rect 23042 4313 23052 4347
rect 23086 4313 23256 4347
rect 23042 4303 23256 4313
rect 22579 4229 22609 4261
rect 22969 4229 22999 4301
rect 23042 4297 23094 4303
rect 23064 4275 23094 4297
rect 23226 4274 23256 4303
rect 23318 4347 23377 4363
rect 23318 4313 23328 4347
rect 23362 4313 23377 4347
rect 23318 4297 23377 4313
rect 23347 4275 23377 4297
rect 23226 4244 23282 4274
rect 23252 4229 23282 4244
rect 25656 4234 25686 4260
rect 25740 4234 25770 4260
rect 25928 4234 25958 4260
rect 26023 4234 26053 4260
rect 26129 4234 26159 4260
rect 26225 4234 26255 4260
rect 26335 4234 26365 4260
rect 26435 4234 26465 4260
rect 26519 4234 26549 4260
rect 26707 4234 26737 4260
rect 26802 4234 26832 4260
rect 26911 4234 26941 4260
rect 27006 4234 27036 4260
rect 27092 4234 27122 4260
rect 27210 4234 27240 4260
rect 27294 4234 27324 4260
rect 27482 4234 27512 4260
rect 27577 4234 27607 4260
rect 27765 4234 27795 4260
rect 27860 4234 27890 4260
rect 28048 4234 28078 4260
rect 28132 4234 28162 4260
rect 28320 4234 28350 4260
rect 28415 4234 28445 4260
rect 28521 4234 28551 4260
rect 28617 4234 28647 4260
rect 28727 4234 28757 4260
rect 28827 4234 28857 4260
rect 28911 4234 28941 4260
rect 29099 4234 29129 4260
rect 29194 4234 29224 4260
rect 29303 4234 29333 4260
rect 29398 4234 29428 4260
rect 29484 4234 29514 4260
rect 29602 4234 29632 4260
rect 29686 4234 29716 4260
rect 29874 4234 29904 4260
rect 29969 4234 29999 4260
rect 30157 4234 30187 4260
rect 30252 4234 30282 4260
rect 11168 4118 11198 4144
rect 11256 4118 11286 4144
rect 11444 4118 11474 4144
rect 11528 4118 11558 4144
rect 11612 4118 11642 4144
rect 11696 4118 11726 4144
rect 11780 4118 11810 4144
rect 13751 4119 13781 4145
rect 13967 4119 13997 4145
rect 14051 4119 14081 4145
rect 14239 4119 14269 4145
rect 14334 4119 14364 4145
rect 14440 4119 14470 4145
rect 14536 4119 14566 4145
rect 14646 4119 14676 4145
rect 14746 4119 14776 4145
rect 14830 4119 14860 4145
rect 15018 4119 15048 4145
rect 15113 4119 15143 4145
rect 15222 4119 15252 4145
rect 15317 4119 15347 4145
rect 15403 4119 15433 4145
rect 15521 4119 15551 4145
rect 15605 4119 15635 4145
rect 15793 4119 15823 4145
rect 15888 4119 15918 4145
rect 16076 4119 16106 4145
rect 16171 4119 16201 4145
rect 16359 4119 16389 4145
rect 16443 4119 16473 4145
rect 16631 4119 16661 4145
rect 16726 4119 16756 4145
rect 16832 4119 16862 4145
rect 16928 4119 16958 4145
rect 17038 4119 17068 4145
rect 17138 4119 17168 4145
rect 17222 4119 17252 4145
rect 17410 4119 17440 4145
rect 17505 4119 17535 4145
rect 17614 4119 17644 4145
rect 17709 4119 17739 4145
rect 17795 4119 17825 4145
rect 17913 4119 17943 4145
rect 17997 4119 18027 4145
rect 18185 4119 18215 4145
rect 18280 4119 18310 4145
rect 18468 4119 18498 4145
rect 18563 4119 18593 4145
rect 18751 4119 18781 4145
rect 18835 4119 18865 4145
rect 19023 4119 19053 4145
rect 19118 4119 19148 4145
rect 19224 4119 19254 4145
rect 19320 4119 19350 4145
rect 19430 4119 19460 4145
rect 19530 4119 19560 4145
rect 19614 4119 19644 4145
rect 19802 4119 19832 4145
rect 19897 4119 19927 4145
rect 20006 4119 20036 4145
rect 20101 4119 20131 4145
rect 20187 4119 20217 4145
rect 20305 4119 20335 4145
rect 20389 4119 20419 4145
rect 20577 4119 20607 4145
rect 20672 4119 20702 4145
rect 20860 4119 20890 4145
rect 20955 4119 20985 4145
rect 21143 4119 21173 4145
rect 21227 4119 21257 4145
rect 21415 4119 21445 4145
rect 21510 4119 21540 4145
rect 21616 4119 21646 4145
rect 21712 4119 21742 4145
rect 21822 4119 21852 4145
rect 21922 4119 21952 4145
rect 22006 4119 22036 4145
rect 22194 4119 22224 4145
rect 22289 4119 22319 4145
rect 22398 4119 22428 4145
rect 22493 4119 22523 4145
rect 22579 4119 22609 4145
rect 22697 4119 22727 4145
rect 22781 4119 22811 4145
rect 22969 4119 22999 4145
rect 23064 4119 23094 4145
rect 23252 4119 23282 4145
rect 23347 4119 23377 4145
rect 25656 4135 25686 4150
rect 25623 4105 25686 4135
rect 25623 4067 25653 4105
rect 25598 4051 25653 4067
rect 25740 4061 25770 4150
rect 25928 4080 25958 4150
rect 26023 4140 26053 4162
rect 26023 4124 26087 4140
rect 26023 4090 26043 4124
rect 26077 4090 26087 4124
rect 25598 4017 25609 4051
rect 25643 4017 25653 4051
rect 25598 4001 25653 4017
rect 25695 4051 25770 4061
rect 25695 4017 25711 4051
rect 25745 4017 25770 4051
rect 25695 4007 25770 4017
rect 25917 4064 25971 4080
rect 26023 4074 26087 4090
rect 26129 4128 26159 4162
rect 26129 4112 26183 4128
rect 26129 4078 26139 4112
rect 26173 4078 26183 4112
rect 25917 4030 25927 4064
rect 25961 4030 25971 4064
rect 26129 4062 26183 4078
rect 26129 4032 26159 4062
rect 25917 4014 25971 4030
rect 25623 3963 25653 4001
rect 25623 3933 25686 3963
rect 25656 3918 25686 3933
rect 25740 3918 25770 4007
rect 25928 3868 25958 4014
rect 26021 4002 26159 4032
rect 26021 3868 26051 4002
rect 26225 3966 26255 4150
rect 26335 4118 26365 4150
rect 26301 4102 26365 4118
rect 26802 4140 26832 4162
rect 26802 4124 26869 4140
rect 26301 4068 26311 4102
rect 26345 4088 26365 4102
rect 26345 4068 26361 4088
rect 26301 4052 26361 4068
rect 26093 3950 26159 3960
rect 26093 3916 26109 3950
rect 26143 3916 26159 3950
rect 26093 3906 26159 3916
rect 26225 3950 26289 3966
rect 26225 3916 26245 3950
rect 26279 3916 26289 3950
rect 26105 3868 26135 3906
rect 26225 3900 26289 3916
rect 26225 3868 26255 3900
rect 26331 3868 26361 4052
rect 26435 4050 26465 4106
rect 26519 4050 26549 4106
rect 26707 4084 26737 4106
rect 26683 4068 26737 4084
rect 26802 4090 26825 4124
rect 26859 4090 26869 4124
rect 26802 4074 26869 4090
rect 26403 4034 26469 4050
rect 26403 4000 26413 4034
rect 26447 4000 26469 4034
rect 26403 3984 26469 4000
rect 26519 4034 26609 4050
rect 26683 4048 26693 4068
rect 26519 4000 26565 4034
rect 26599 4000 26609 4034
rect 26519 3984 26609 4000
rect 26660 4034 26693 4048
rect 26727 4034 26737 4068
rect 26660 4018 26737 4034
rect 26911 4032 26941 4162
rect 26439 3952 26469 3984
rect 26523 3952 26553 3984
rect 26660 3952 26690 4018
rect 26804 4002 26941 4032
rect 26804 3966 26834 4002
rect 25656 3764 25686 3790
rect 25740 3764 25770 3790
rect 26780 3950 26834 3966
rect 27006 3966 27036 4150
rect 27092 4118 27122 4150
rect 27078 4102 27144 4118
rect 27078 4068 27088 4102
rect 27122 4068 27144 4102
rect 27078 4052 27144 4068
rect 27210 4066 27240 4106
rect 26780 3916 26790 3950
rect 26824 3916 26834 3950
rect 26780 3900 26834 3916
rect 26876 3950 26942 3960
rect 26876 3916 26892 3950
rect 26926 3916 26942 3950
rect 26876 3906 26942 3916
rect 27006 3950 27072 3966
rect 27006 3916 27028 3950
rect 27062 3916 27072 3950
rect 26804 3868 26834 3900
rect 26888 3868 26918 3906
rect 27006 3900 27072 3916
rect 27006 3868 27036 3900
rect 27114 3868 27144 4052
rect 27186 4050 27240 4066
rect 27186 4016 27196 4050
rect 27230 4016 27240 4050
rect 27186 4000 27240 4016
rect 27294 4050 27324 4106
rect 27482 4078 27512 4150
rect 27765 4135 27795 4150
rect 27739 4105 27795 4135
rect 27577 4082 27607 4104
rect 27449 4062 27513 4078
rect 27294 4034 27378 4050
rect 27294 4014 27334 4034
rect 27210 3952 27240 4000
rect 27282 4000 27334 4014
rect 27368 4000 27378 4034
rect 27449 4028 27465 4062
rect 27499 4028 27513 4062
rect 27449 4012 27513 4028
rect 27555 4076 27607 4082
rect 27739 4076 27769 4105
rect 28048 4135 28078 4150
rect 28015 4105 28078 4135
rect 27860 4082 27890 4104
rect 27555 4066 27769 4076
rect 27555 4032 27565 4066
rect 27599 4032 27769 4066
rect 27555 4022 27769 4032
rect 27555 4016 27607 4022
rect 27282 3984 27378 4000
rect 27282 3952 27312 3984
rect 27480 3980 27510 4012
rect 27577 3984 27607 4016
rect 27480 3826 27510 3852
rect 27739 3974 27769 4022
rect 27831 4066 27890 4082
rect 28015 4067 28045 4105
rect 27831 4032 27841 4066
rect 27875 4032 27890 4066
rect 27831 4016 27890 4032
rect 27860 3984 27890 4016
rect 27990 4051 28045 4067
rect 28132 4061 28162 4150
rect 28320 4080 28350 4150
rect 28415 4140 28445 4162
rect 28415 4124 28479 4140
rect 28415 4090 28435 4124
rect 28469 4090 28479 4124
rect 27990 4017 28001 4051
rect 28035 4017 28045 4051
rect 27990 4001 28045 4017
rect 28087 4051 28162 4061
rect 28087 4017 28103 4051
rect 28137 4017 28162 4051
rect 28087 4007 28162 4017
rect 28309 4064 28363 4080
rect 28415 4074 28479 4090
rect 28521 4128 28551 4162
rect 28521 4112 28575 4128
rect 28521 4078 28531 4112
rect 28565 4078 28575 4112
rect 28309 4030 28319 4064
rect 28353 4030 28363 4064
rect 28521 4062 28575 4078
rect 28521 4032 28551 4062
rect 28309 4014 28363 4030
rect 27739 3944 27795 3974
rect 27765 3928 27795 3944
rect 25928 3758 25958 3784
rect 26021 3758 26051 3784
rect 26105 3758 26135 3784
rect 26225 3758 26255 3784
rect 26331 3758 26361 3784
rect 26439 3758 26469 3784
rect 26523 3758 26553 3784
rect 26660 3758 26690 3784
rect 26804 3758 26834 3784
rect 26888 3758 26918 3784
rect 27006 3758 27036 3784
rect 27114 3758 27144 3784
rect 27210 3758 27240 3784
rect 27282 3758 27312 3784
rect 27577 3758 27607 3784
rect 27765 3774 27795 3800
rect 28015 3963 28045 4001
rect 28015 3933 28078 3963
rect 28048 3918 28078 3933
rect 28132 3918 28162 4007
rect 28320 3868 28350 4014
rect 28413 4002 28551 4032
rect 28413 3868 28443 4002
rect 28617 3966 28647 4150
rect 28727 4118 28757 4150
rect 28693 4102 28757 4118
rect 29194 4140 29224 4162
rect 29194 4124 29261 4140
rect 28693 4068 28703 4102
rect 28737 4088 28757 4102
rect 28737 4068 28753 4088
rect 28693 4052 28753 4068
rect 28485 3950 28551 3960
rect 28485 3916 28501 3950
rect 28535 3916 28551 3950
rect 28485 3906 28551 3916
rect 28617 3950 28681 3966
rect 28617 3916 28637 3950
rect 28671 3916 28681 3950
rect 28497 3868 28527 3906
rect 28617 3900 28681 3916
rect 28617 3868 28647 3900
rect 28723 3868 28753 4052
rect 28827 4050 28857 4106
rect 28911 4050 28941 4106
rect 29099 4084 29129 4106
rect 29075 4068 29129 4084
rect 29194 4090 29217 4124
rect 29251 4090 29261 4124
rect 29194 4074 29261 4090
rect 28795 4034 28861 4050
rect 28795 4000 28805 4034
rect 28839 4000 28861 4034
rect 28795 3984 28861 4000
rect 28911 4034 29001 4050
rect 29075 4048 29085 4068
rect 28911 4000 28957 4034
rect 28991 4000 29001 4034
rect 28911 3984 29001 4000
rect 29052 4034 29085 4048
rect 29119 4034 29129 4068
rect 29052 4018 29129 4034
rect 29303 4032 29333 4162
rect 28831 3952 28861 3984
rect 28915 3952 28945 3984
rect 29052 3952 29082 4018
rect 29196 4002 29333 4032
rect 29196 3966 29226 4002
rect 27860 3758 27890 3784
rect 28048 3764 28078 3790
rect 28132 3764 28162 3790
rect 29172 3950 29226 3966
rect 29398 3966 29428 4150
rect 29484 4118 29514 4150
rect 29470 4102 29536 4118
rect 29470 4068 29480 4102
rect 29514 4068 29536 4102
rect 29470 4052 29536 4068
rect 29602 4066 29632 4106
rect 29172 3916 29182 3950
rect 29216 3916 29226 3950
rect 29172 3900 29226 3916
rect 29268 3950 29334 3960
rect 29268 3916 29284 3950
rect 29318 3916 29334 3950
rect 29268 3906 29334 3916
rect 29398 3950 29464 3966
rect 29398 3916 29420 3950
rect 29454 3916 29464 3950
rect 29196 3868 29226 3900
rect 29280 3868 29310 3906
rect 29398 3900 29464 3916
rect 29398 3868 29428 3900
rect 29506 3868 29536 4052
rect 29578 4050 29632 4066
rect 29578 4016 29588 4050
rect 29622 4016 29632 4050
rect 29578 4000 29632 4016
rect 29686 4050 29716 4106
rect 29874 4078 29904 4150
rect 30157 4135 30187 4150
rect 30131 4105 30187 4135
rect 29969 4082 29999 4104
rect 29841 4062 29905 4078
rect 29686 4034 29770 4050
rect 29686 4014 29726 4034
rect 29602 3952 29632 4000
rect 29674 4000 29726 4014
rect 29760 4000 29770 4034
rect 29841 4028 29857 4062
rect 29891 4028 29905 4062
rect 29841 4012 29905 4028
rect 29947 4076 29999 4082
rect 30131 4076 30161 4105
rect 30252 4082 30282 4104
rect 29947 4066 30161 4076
rect 29947 4032 29957 4066
rect 29991 4032 30161 4066
rect 29947 4022 30161 4032
rect 29947 4016 29999 4022
rect 29674 3984 29770 4000
rect 29674 3952 29704 3984
rect 29872 3980 29902 4012
rect 29969 3984 29999 4016
rect 29872 3826 29902 3852
rect 30131 3974 30161 4022
rect 30223 4066 30282 4082
rect 30223 4032 30233 4066
rect 30267 4032 30282 4066
rect 30223 4016 30282 4032
rect 30252 3984 30282 4016
rect 30131 3944 30187 3974
rect 30157 3928 30187 3944
rect 28320 3758 28350 3784
rect 28413 3758 28443 3784
rect 28497 3758 28527 3784
rect 28617 3758 28647 3784
rect 28723 3758 28753 3784
rect 28831 3758 28861 3784
rect 28915 3758 28945 3784
rect 29052 3758 29082 3784
rect 29196 3758 29226 3784
rect 29280 3758 29310 3784
rect 29398 3758 29428 3784
rect 29506 3758 29536 3784
rect 29602 3758 29632 3784
rect 29674 3758 29704 3784
rect 29969 3758 29999 3784
rect 30157 3774 30187 3800
rect 30252 3758 30282 3784
rect 11575 3722 11605 3748
rect 11670 3706 11700 3732
rect 11858 3722 11888 3748
rect 12153 3722 12183 3748
rect 12225 3722 12255 3748
rect 12321 3722 12351 3748
rect 12429 3722 12459 3748
rect 12547 3722 12577 3748
rect 12631 3722 12661 3748
rect 12775 3722 12805 3748
rect 12912 3722 12942 3748
rect 12996 3722 13026 3748
rect 13104 3722 13134 3748
rect 13210 3722 13240 3748
rect 13330 3722 13360 3748
rect 13414 3722 13444 3748
rect 13507 3722 13537 3748
rect 11670 3562 11700 3578
rect 11670 3532 11726 3562
rect 11575 3490 11605 3522
rect 11575 3474 11634 3490
rect 11575 3440 11590 3474
rect 11624 3440 11634 3474
rect 11575 3424 11634 3440
rect 11696 3484 11726 3532
rect 11955 3654 11985 3680
rect 11858 3490 11888 3522
rect 11955 3494 11985 3526
rect 12153 3522 12183 3554
rect 12087 3506 12183 3522
rect 11858 3484 11910 3490
rect 11696 3474 11910 3484
rect 11696 3440 11866 3474
rect 11900 3440 11910 3474
rect 11696 3430 11910 3440
rect 11575 3402 11605 3424
rect 11696 3401 11726 3430
rect 11858 3424 11910 3430
rect 11952 3478 12016 3494
rect 11952 3444 11966 3478
rect 12000 3444 12016 3478
rect 12087 3472 12097 3506
rect 12131 3492 12183 3506
rect 12225 3506 12255 3554
rect 12131 3472 12171 3492
rect 12087 3456 12171 3472
rect 11952 3428 12016 3444
rect 11858 3402 11888 3424
rect 11670 3371 11726 3401
rect 11670 3356 11700 3371
rect 11953 3356 11983 3428
rect 12141 3400 12171 3456
rect 12225 3490 12279 3506
rect 12225 3456 12235 3490
rect 12269 3456 12279 3490
rect 12225 3440 12279 3456
rect 12321 3454 12351 3638
rect 12429 3606 12459 3638
rect 12393 3590 12459 3606
rect 12547 3600 12577 3638
rect 12631 3606 12661 3638
rect 12393 3556 12403 3590
rect 12437 3556 12459 3590
rect 12393 3540 12459 3556
rect 12523 3590 12589 3600
rect 12523 3556 12539 3590
rect 12573 3556 12589 3590
rect 12523 3546 12589 3556
rect 12631 3590 12685 3606
rect 12631 3556 12641 3590
rect 12675 3556 12685 3590
rect 12225 3400 12255 3440
rect 12321 3438 12387 3454
rect 12321 3404 12343 3438
rect 12377 3404 12387 3438
rect 12321 3388 12387 3404
rect 12343 3356 12373 3388
rect 12429 3356 12459 3540
rect 12631 3540 12685 3556
rect 13695 3716 13725 3742
rect 13779 3716 13809 3742
rect 13967 3722 13997 3748
rect 12631 3504 12661 3540
rect 12524 3474 12661 3504
rect 12775 3488 12805 3554
rect 12912 3522 12942 3554
rect 12996 3522 13026 3554
rect 12524 3344 12554 3474
rect 12728 3472 12805 3488
rect 12728 3438 12738 3472
rect 12772 3458 12805 3472
rect 12856 3506 12946 3522
rect 12856 3472 12866 3506
rect 12900 3472 12946 3506
rect 12772 3438 12782 3458
rect 12856 3456 12946 3472
rect 12996 3506 13062 3522
rect 12996 3472 13018 3506
rect 13052 3472 13062 3506
rect 12996 3456 13062 3472
rect 12596 3416 12663 3432
rect 12596 3382 12606 3416
rect 12640 3382 12663 3416
rect 12728 3422 12782 3438
rect 12728 3400 12758 3422
rect 12916 3400 12946 3456
rect 13000 3400 13030 3456
rect 13104 3454 13134 3638
rect 13210 3606 13240 3638
rect 13176 3590 13240 3606
rect 13330 3600 13360 3638
rect 13176 3556 13186 3590
rect 13220 3556 13240 3590
rect 13176 3540 13240 3556
rect 13306 3590 13372 3600
rect 13306 3556 13322 3590
rect 13356 3556 13372 3590
rect 13306 3546 13372 3556
rect 13104 3438 13164 3454
rect 13104 3418 13120 3438
rect 13100 3404 13120 3418
rect 13154 3404 13164 3438
rect 12596 3366 12663 3382
rect 12633 3344 12663 3366
rect 13100 3388 13164 3404
rect 13100 3356 13130 3388
rect 13210 3356 13240 3540
rect 13414 3504 13444 3638
rect 13306 3474 13444 3504
rect 13507 3492 13537 3638
rect 13695 3499 13725 3588
rect 13779 3573 13809 3588
rect 13779 3543 13842 3573
rect 13812 3505 13842 3543
rect 14062 3706 14092 3732
rect 14250 3722 14280 3748
rect 14545 3722 14575 3748
rect 14617 3722 14647 3748
rect 14713 3722 14743 3748
rect 14821 3722 14851 3748
rect 14939 3722 14969 3748
rect 15023 3722 15053 3748
rect 15167 3722 15197 3748
rect 15304 3722 15334 3748
rect 15388 3722 15418 3748
rect 15496 3722 15526 3748
rect 15602 3722 15632 3748
rect 15722 3722 15752 3748
rect 15806 3722 15836 3748
rect 15899 3722 15929 3748
rect 14062 3562 14092 3578
rect 14062 3532 14118 3562
rect 13494 3476 13548 3492
rect 13306 3444 13336 3474
rect 13282 3428 13336 3444
rect 13494 3442 13504 3476
rect 13538 3442 13548 3476
rect 13282 3394 13292 3428
rect 13326 3394 13336 3428
rect 13282 3378 13336 3394
rect 13306 3344 13336 3378
rect 13378 3416 13442 3432
rect 13494 3426 13548 3442
rect 13695 3489 13770 3499
rect 13695 3455 13720 3489
rect 13754 3455 13770 3489
rect 13695 3445 13770 3455
rect 13812 3489 13867 3505
rect 13812 3455 13822 3489
rect 13856 3455 13867 3489
rect 13378 3382 13388 3416
rect 13422 3382 13442 3416
rect 13378 3366 13442 3382
rect 13412 3344 13442 3366
rect 13507 3356 13537 3426
rect 13695 3356 13725 3445
rect 13812 3439 13867 3455
rect 13967 3490 13997 3522
rect 13967 3474 14026 3490
rect 13967 3440 13982 3474
rect 14016 3440 14026 3474
rect 13812 3401 13842 3439
rect 13967 3424 14026 3440
rect 14088 3484 14118 3532
rect 14347 3654 14377 3680
rect 14250 3490 14280 3522
rect 14347 3494 14377 3526
rect 14545 3522 14575 3554
rect 14479 3506 14575 3522
rect 14250 3484 14302 3490
rect 14088 3474 14302 3484
rect 14088 3440 14258 3474
rect 14292 3440 14302 3474
rect 14088 3430 14302 3440
rect 13967 3402 13997 3424
rect 13779 3371 13842 3401
rect 13779 3356 13809 3371
rect 14088 3401 14118 3430
rect 14250 3424 14302 3430
rect 14344 3478 14408 3494
rect 14344 3444 14358 3478
rect 14392 3444 14408 3478
rect 14479 3472 14489 3506
rect 14523 3492 14575 3506
rect 14617 3506 14647 3554
rect 14523 3472 14563 3492
rect 14479 3456 14563 3472
rect 14344 3428 14408 3444
rect 14250 3402 14280 3424
rect 14062 3371 14118 3401
rect 14062 3356 14092 3371
rect 14345 3356 14375 3428
rect 14533 3400 14563 3456
rect 14617 3490 14671 3506
rect 14617 3456 14627 3490
rect 14661 3456 14671 3490
rect 14617 3440 14671 3456
rect 14713 3454 14743 3638
rect 14821 3606 14851 3638
rect 14785 3590 14851 3606
rect 14939 3600 14969 3638
rect 15023 3606 15053 3638
rect 14785 3556 14795 3590
rect 14829 3556 14851 3590
rect 14785 3540 14851 3556
rect 14915 3590 14981 3600
rect 14915 3556 14931 3590
rect 14965 3556 14981 3590
rect 14915 3546 14981 3556
rect 15023 3590 15077 3606
rect 15023 3556 15033 3590
rect 15067 3556 15077 3590
rect 14617 3400 14647 3440
rect 14713 3438 14779 3454
rect 14713 3404 14735 3438
rect 14769 3404 14779 3438
rect 14713 3388 14779 3404
rect 14735 3356 14765 3388
rect 14821 3356 14851 3540
rect 15023 3540 15077 3556
rect 16087 3716 16117 3742
rect 16171 3716 16201 3742
rect 16359 3722 16389 3748
rect 15023 3504 15053 3540
rect 14916 3474 15053 3504
rect 15167 3488 15197 3554
rect 15304 3522 15334 3554
rect 15388 3522 15418 3554
rect 14916 3344 14946 3474
rect 15120 3472 15197 3488
rect 15120 3438 15130 3472
rect 15164 3458 15197 3472
rect 15248 3506 15338 3522
rect 15248 3472 15258 3506
rect 15292 3472 15338 3506
rect 15164 3438 15174 3458
rect 15248 3456 15338 3472
rect 15388 3506 15454 3522
rect 15388 3472 15410 3506
rect 15444 3472 15454 3506
rect 15388 3456 15454 3472
rect 14988 3416 15055 3432
rect 14988 3382 14998 3416
rect 15032 3382 15055 3416
rect 15120 3422 15174 3438
rect 15120 3400 15150 3422
rect 15308 3400 15338 3456
rect 15392 3400 15422 3456
rect 15496 3454 15526 3638
rect 15602 3606 15632 3638
rect 15568 3590 15632 3606
rect 15722 3600 15752 3638
rect 15568 3556 15578 3590
rect 15612 3556 15632 3590
rect 15568 3540 15632 3556
rect 15698 3590 15764 3600
rect 15698 3556 15714 3590
rect 15748 3556 15764 3590
rect 15698 3546 15764 3556
rect 15496 3438 15556 3454
rect 15496 3418 15512 3438
rect 15492 3404 15512 3418
rect 15546 3404 15556 3438
rect 14988 3366 15055 3382
rect 15025 3344 15055 3366
rect 15492 3388 15556 3404
rect 15492 3356 15522 3388
rect 15602 3356 15632 3540
rect 15806 3504 15836 3638
rect 15698 3474 15836 3504
rect 15899 3492 15929 3638
rect 16087 3499 16117 3588
rect 16171 3573 16201 3588
rect 16171 3543 16234 3573
rect 16204 3505 16234 3543
rect 16454 3706 16484 3732
rect 16642 3722 16672 3748
rect 16937 3722 16967 3748
rect 17009 3722 17039 3748
rect 17105 3722 17135 3748
rect 17213 3722 17243 3748
rect 17331 3722 17361 3748
rect 17415 3722 17445 3748
rect 17559 3722 17589 3748
rect 17696 3722 17726 3748
rect 17780 3722 17810 3748
rect 17888 3722 17918 3748
rect 17994 3722 18024 3748
rect 18114 3722 18144 3748
rect 18198 3722 18228 3748
rect 18291 3722 18321 3748
rect 16454 3562 16484 3578
rect 16454 3532 16510 3562
rect 15886 3476 15940 3492
rect 15698 3444 15728 3474
rect 15674 3428 15728 3444
rect 15886 3442 15896 3476
rect 15930 3442 15940 3476
rect 15674 3394 15684 3428
rect 15718 3394 15728 3428
rect 15674 3378 15728 3394
rect 15698 3344 15728 3378
rect 15770 3416 15834 3432
rect 15886 3426 15940 3442
rect 16087 3489 16162 3499
rect 16087 3455 16112 3489
rect 16146 3455 16162 3489
rect 16087 3445 16162 3455
rect 16204 3489 16259 3505
rect 16204 3455 16214 3489
rect 16248 3455 16259 3489
rect 15770 3382 15780 3416
rect 15814 3382 15834 3416
rect 15770 3366 15834 3382
rect 15804 3344 15834 3366
rect 15899 3356 15929 3426
rect 16087 3356 16117 3445
rect 16204 3439 16259 3455
rect 16359 3490 16389 3522
rect 16359 3474 16418 3490
rect 16359 3440 16374 3474
rect 16408 3440 16418 3474
rect 16204 3401 16234 3439
rect 16359 3424 16418 3440
rect 16480 3484 16510 3532
rect 16739 3654 16769 3680
rect 16642 3490 16672 3522
rect 16739 3494 16769 3526
rect 16937 3522 16967 3554
rect 16871 3506 16967 3522
rect 16642 3484 16694 3490
rect 16480 3474 16694 3484
rect 16480 3440 16650 3474
rect 16684 3440 16694 3474
rect 16480 3430 16694 3440
rect 16359 3402 16389 3424
rect 16171 3371 16234 3401
rect 16171 3356 16201 3371
rect 16480 3401 16510 3430
rect 16642 3424 16694 3430
rect 16736 3478 16800 3494
rect 16736 3444 16750 3478
rect 16784 3444 16800 3478
rect 16871 3472 16881 3506
rect 16915 3492 16967 3506
rect 17009 3506 17039 3554
rect 16915 3472 16955 3492
rect 16871 3456 16955 3472
rect 16736 3428 16800 3444
rect 16642 3402 16672 3424
rect 16454 3371 16510 3401
rect 16454 3356 16484 3371
rect 16737 3356 16767 3428
rect 16925 3400 16955 3456
rect 17009 3490 17063 3506
rect 17009 3456 17019 3490
rect 17053 3456 17063 3490
rect 17009 3440 17063 3456
rect 17105 3454 17135 3638
rect 17213 3606 17243 3638
rect 17177 3590 17243 3606
rect 17331 3600 17361 3638
rect 17415 3606 17445 3638
rect 17177 3556 17187 3590
rect 17221 3556 17243 3590
rect 17177 3540 17243 3556
rect 17307 3590 17373 3600
rect 17307 3556 17323 3590
rect 17357 3556 17373 3590
rect 17307 3546 17373 3556
rect 17415 3590 17469 3606
rect 17415 3556 17425 3590
rect 17459 3556 17469 3590
rect 17009 3400 17039 3440
rect 17105 3438 17171 3454
rect 17105 3404 17127 3438
rect 17161 3404 17171 3438
rect 17105 3388 17171 3404
rect 17127 3356 17157 3388
rect 17213 3356 17243 3540
rect 17415 3540 17469 3556
rect 18479 3716 18509 3742
rect 18563 3716 18593 3742
rect 18751 3722 18781 3748
rect 17415 3504 17445 3540
rect 17308 3474 17445 3504
rect 17559 3488 17589 3554
rect 17696 3522 17726 3554
rect 17780 3522 17810 3554
rect 17308 3344 17338 3474
rect 17512 3472 17589 3488
rect 17512 3438 17522 3472
rect 17556 3458 17589 3472
rect 17640 3506 17730 3522
rect 17640 3472 17650 3506
rect 17684 3472 17730 3506
rect 17556 3438 17566 3458
rect 17640 3456 17730 3472
rect 17780 3506 17846 3522
rect 17780 3472 17802 3506
rect 17836 3472 17846 3506
rect 17780 3456 17846 3472
rect 17380 3416 17447 3432
rect 17380 3382 17390 3416
rect 17424 3382 17447 3416
rect 17512 3422 17566 3438
rect 17512 3400 17542 3422
rect 17700 3400 17730 3456
rect 17784 3400 17814 3456
rect 17888 3454 17918 3638
rect 17994 3606 18024 3638
rect 17960 3590 18024 3606
rect 18114 3600 18144 3638
rect 17960 3556 17970 3590
rect 18004 3556 18024 3590
rect 17960 3540 18024 3556
rect 18090 3590 18156 3600
rect 18090 3556 18106 3590
rect 18140 3556 18156 3590
rect 18090 3546 18156 3556
rect 17888 3438 17948 3454
rect 17888 3418 17904 3438
rect 17884 3404 17904 3418
rect 17938 3404 17948 3438
rect 17380 3366 17447 3382
rect 17417 3344 17447 3366
rect 17884 3388 17948 3404
rect 17884 3356 17914 3388
rect 17994 3356 18024 3540
rect 18198 3504 18228 3638
rect 18090 3474 18228 3504
rect 18291 3492 18321 3638
rect 18479 3499 18509 3588
rect 18563 3573 18593 3588
rect 18563 3543 18626 3573
rect 18596 3505 18626 3543
rect 18846 3706 18876 3732
rect 19034 3722 19064 3748
rect 19329 3722 19359 3748
rect 19401 3722 19431 3748
rect 19497 3722 19527 3748
rect 19605 3722 19635 3748
rect 19723 3722 19753 3748
rect 19807 3722 19837 3748
rect 19951 3722 19981 3748
rect 20088 3722 20118 3748
rect 20172 3722 20202 3748
rect 20280 3722 20310 3748
rect 20386 3722 20416 3748
rect 20506 3722 20536 3748
rect 20590 3722 20620 3748
rect 20683 3722 20713 3748
rect 18846 3562 18876 3578
rect 18846 3532 18902 3562
rect 18278 3476 18332 3492
rect 18090 3444 18120 3474
rect 18066 3428 18120 3444
rect 18278 3442 18288 3476
rect 18322 3442 18332 3476
rect 18066 3394 18076 3428
rect 18110 3394 18120 3428
rect 18066 3378 18120 3394
rect 18090 3344 18120 3378
rect 18162 3416 18226 3432
rect 18278 3426 18332 3442
rect 18479 3489 18554 3499
rect 18479 3455 18504 3489
rect 18538 3455 18554 3489
rect 18479 3445 18554 3455
rect 18596 3489 18651 3505
rect 18596 3455 18606 3489
rect 18640 3455 18651 3489
rect 18162 3382 18172 3416
rect 18206 3382 18226 3416
rect 18162 3366 18226 3382
rect 18196 3344 18226 3366
rect 18291 3356 18321 3426
rect 18479 3356 18509 3445
rect 18596 3439 18651 3455
rect 18751 3490 18781 3522
rect 18751 3474 18810 3490
rect 18751 3440 18766 3474
rect 18800 3440 18810 3474
rect 18596 3401 18626 3439
rect 18751 3424 18810 3440
rect 18872 3484 18902 3532
rect 19131 3654 19161 3680
rect 19034 3490 19064 3522
rect 19131 3494 19161 3526
rect 19329 3522 19359 3554
rect 19263 3506 19359 3522
rect 19034 3484 19086 3490
rect 18872 3474 19086 3484
rect 18872 3440 19042 3474
rect 19076 3440 19086 3474
rect 18872 3430 19086 3440
rect 18751 3402 18781 3424
rect 18563 3371 18626 3401
rect 18563 3356 18593 3371
rect 18872 3401 18902 3430
rect 19034 3424 19086 3430
rect 19128 3478 19192 3494
rect 19128 3444 19142 3478
rect 19176 3444 19192 3478
rect 19263 3472 19273 3506
rect 19307 3492 19359 3506
rect 19401 3506 19431 3554
rect 19307 3472 19347 3492
rect 19263 3456 19347 3472
rect 19128 3428 19192 3444
rect 19034 3402 19064 3424
rect 18846 3371 18902 3401
rect 18846 3356 18876 3371
rect 19129 3356 19159 3428
rect 19317 3400 19347 3456
rect 19401 3490 19455 3506
rect 19401 3456 19411 3490
rect 19445 3456 19455 3490
rect 19401 3440 19455 3456
rect 19497 3454 19527 3638
rect 19605 3606 19635 3638
rect 19569 3590 19635 3606
rect 19723 3600 19753 3638
rect 19807 3606 19837 3638
rect 19569 3556 19579 3590
rect 19613 3556 19635 3590
rect 19569 3540 19635 3556
rect 19699 3590 19765 3600
rect 19699 3556 19715 3590
rect 19749 3556 19765 3590
rect 19699 3546 19765 3556
rect 19807 3590 19861 3606
rect 19807 3556 19817 3590
rect 19851 3556 19861 3590
rect 19401 3400 19431 3440
rect 19497 3438 19563 3454
rect 19497 3404 19519 3438
rect 19553 3404 19563 3438
rect 19497 3388 19563 3404
rect 19519 3356 19549 3388
rect 19605 3356 19635 3540
rect 19807 3540 19861 3556
rect 20871 3716 20901 3742
rect 20955 3716 20985 3742
rect 21143 3722 21173 3748
rect 19807 3504 19837 3540
rect 19700 3474 19837 3504
rect 19951 3488 19981 3554
rect 20088 3522 20118 3554
rect 20172 3522 20202 3554
rect 19700 3344 19730 3474
rect 19904 3472 19981 3488
rect 19904 3438 19914 3472
rect 19948 3458 19981 3472
rect 20032 3506 20122 3522
rect 20032 3472 20042 3506
rect 20076 3472 20122 3506
rect 19948 3438 19958 3458
rect 20032 3456 20122 3472
rect 20172 3506 20238 3522
rect 20172 3472 20194 3506
rect 20228 3472 20238 3506
rect 20172 3456 20238 3472
rect 19772 3416 19839 3432
rect 19772 3382 19782 3416
rect 19816 3382 19839 3416
rect 19904 3422 19958 3438
rect 19904 3400 19934 3422
rect 20092 3400 20122 3456
rect 20176 3400 20206 3456
rect 20280 3454 20310 3638
rect 20386 3606 20416 3638
rect 20352 3590 20416 3606
rect 20506 3600 20536 3638
rect 20352 3556 20362 3590
rect 20396 3556 20416 3590
rect 20352 3540 20416 3556
rect 20482 3590 20548 3600
rect 20482 3556 20498 3590
rect 20532 3556 20548 3590
rect 20482 3546 20548 3556
rect 20280 3438 20340 3454
rect 20280 3418 20296 3438
rect 20276 3404 20296 3418
rect 20330 3404 20340 3438
rect 19772 3366 19839 3382
rect 19809 3344 19839 3366
rect 20276 3388 20340 3404
rect 20276 3356 20306 3388
rect 20386 3356 20416 3540
rect 20590 3504 20620 3638
rect 20482 3474 20620 3504
rect 20683 3492 20713 3638
rect 20871 3499 20901 3588
rect 20955 3573 20985 3588
rect 20955 3543 21018 3573
rect 20988 3505 21018 3543
rect 21238 3706 21268 3732
rect 21426 3722 21456 3748
rect 21721 3722 21751 3748
rect 21793 3722 21823 3748
rect 21889 3722 21919 3748
rect 21997 3722 22027 3748
rect 22115 3722 22145 3748
rect 22199 3722 22229 3748
rect 22343 3722 22373 3748
rect 22480 3722 22510 3748
rect 22564 3722 22594 3748
rect 22672 3722 22702 3748
rect 22778 3722 22808 3748
rect 22898 3722 22928 3748
rect 22982 3722 23012 3748
rect 23075 3722 23105 3748
rect 21238 3562 21268 3578
rect 21238 3532 21294 3562
rect 20670 3476 20724 3492
rect 20482 3444 20512 3474
rect 20458 3428 20512 3444
rect 20670 3442 20680 3476
rect 20714 3442 20724 3476
rect 20458 3394 20468 3428
rect 20502 3394 20512 3428
rect 20458 3378 20512 3394
rect 20482 3344 20512 3378
rect 20554 3416 20618 3432
rect 20670 3426 20724 3442
rect 20871 3489 20946 3499
rect 20871 3455 20896 3489
rect 20930 3455 20946 3489
rect 20871 3445 20946 3455
rect 20988 3489 21043 3505
rect 20988 3455 20998 3489
rect 21032 3455 21043 3489
rect 20554 3382 20564 3416
rect 20598 3382 20618 3416
rect 20554 3366 20618 3382
rect 20588 3344 20618 3366
rect 20683 3356 20713 3426
rect 20871 3356 20901 3445
rect 20988 3439 21043 3455
rect 21143 3490 21173 3522
rect 21143 3474 21202 3490
rect 21143 3440 21158 3474
rect 21192 3440 21202 3474
rect 20988 3401 21018 3439
rect 21143 3424 21202 3440
rect 21264 3484 21294 3532
rect 21523 3654 21553 3680
rect 21426 3490 21456 3522
rect 21523 3494 21553 3526
rect 21721 3522 21751 3554
rect 21655 3506 21751 3522
rect 21426 3484 21478 3490
rect 21264 3474 21478 3484
rect 21264 3440 21434 3474
rect 21468 3440 21478 3474
rect 21264 3430 21478 3440
rect 21143 3402 21173 3424
rect 20955 3371 21018 3401
rect 20955 3356 20985 3371
rect 21264 3401 21294 3430
rect 21426 3424 21478 3430
rect 21520 3478 21584 3494
rect 21520 3444 21534 3478
rect 21568 3444 21584 3478
rect 21655 3472 21665 3506
rect 21699 3492 21751 3506
rect 21793 3506 21823 3554
rect 21699 3472 21739 3492
rect 21655 3456 21739 3472
rect 21520 3428 21584 3444
rect 21426 3402 21456 3424
rect 21238 3371 21294 3401
rect 21238 3356 21268 3371
rect 21521 3356 21551 3428
rect 21709 3400 21739 3456
rect 21793 3490 21847 3506
rect 21793 3456 21803 3490
rect 21837 3456 21847 3490
rect 21793 3440 21847 3456
rect 21889 3454 21919 3638
rect 21997 3606 22027 3638
rect 21961 3590 22027 3606
rect 22115 3600 22145 3638
rect 22199 3606 22229 3638
rect 21961 3556 21971 3590
rect 22005 3556 22027 3590
rect 21961 3540 22027 3556
rect 22091 3590 22157 3600
rect 22091 3556 22107 3590
rect 22141 3556 22157 3590
rect 22091 3546 22157 3556
rect 22199 3590 22253 3606
rect 22199 3556 22209 3590
rect 22243 3556 22253 3590
rect 21793 3400 21823 3440
rect 21889 3438 21955 3454
rect 21889 3404 21911 3438
rect 21945 3404 21955 3438
rect 21889 3388 21955 3404
rect 21911 3356 21941 3388
rect 21997 3356 22027 3540
rect 22199 3540 22253 3556
rect 23263 3716 23293 3742
rect 23347 3716 23377 3742
rect 22199 3504 22229 3540
rect 22092 3474 22229 3504
rect 22343 3488 22373 3554
rect 22480 3522 22510 3554
rect 22564 3522 22594 3554
rect 22092 3344 22122 3474
rect 22296 3472 22373 3488
rect 22296 3438 22306 3472
rect 22340 3458 22373 3472
rect 22424 3506 22514 3522
rect 22424 3472 22434 3506
rect 22468 3472 22514 3506
rect 22340 3438 22350 3458
rect 22424 3456 22514 3472
rect 22564 3506 22630 3522
rect 22564 3472 22586 3506
rect 22620 3472 22630 3506
rect 22564 3456 22630 3472
rect 22164 3416 22231 3432
rect 22164 3382 22174 3416
rect 22208 3382 22231 3416
rect 22296 3422 22350 3438
rect 22296 3400 22326 3422
rect 22484 3400 22514 3456
rect 22568 3400 22598 3456
rect 22672 3454 22702 3638
rect 22778 3606 22808 3638
rect 22744 3590 22808 3606
rect 22898 3600 22928 3638
rect 22744 3556 22754 3590
rect 22788 3556 22808 3590
rect 22744 3540 22808 3556
rect 22874 3590 22940 3600
rect 22874 3556 22890 3590
rect 22924 3556 22940 3590
rect 22874 3546 22940 3556
rect 22672 3438 22732 3454
rect 22672 3418 22688 3438
rect 22668 3404 22688 3418
rect 22722 3404 22732 3438
rect 22164 3366 22231 3382
rect 22201 3344 22231 3366
rect 22668 3388 22732 3404
rect 22668 3356 22698 3388
rect 22778 3356 22808 3540
rect 22982 3504 23012 3638
rect 22874 3474 23012 3504
rect 23075 3492 23105 3638
rect 25656 3588 25686 3614
rect 25740 3588 25770 3614
rect 25928 3594 25958 3620
rect 26021 3594 26051 3620
rect 26105 3594 26135 3620
rect 26225 3594 26255 3620
rect 26331 3594 26361 3620
rect 26439 3594 26469 3620
rect 26523 3594 26553 3620
rect 26660 3594 26690 3620
rect 26804 3594 26834 3620
rect 26888 3594 26918 3620
rect 27006 3594 27036 3620
rect 27114 3594 27144 3620
rect 27210 3594 27240 3620
rect 27282 3594 27312 3620
rect 27577 3594 27607 3620
rect 23263 3499 23293 3588
rect 23347 3573 23377 3588
rect 23347 3543 23410 3573
rect 23380 3505 23410 3543
rect 23062 3476 23116 3492
rect 22874 3444 22904 3474
rect 22850 3428 22904 3444
rect 23062 3442 23072 3476
rect 23106 3442 23116 3476
rect 22850 3394 22860 3428
rect 22894 3394 22904 3428
rect 22850 3378 22904 3394
rect 22874 3344 22904 3378
rect 22946 3416 23010 3432
rect 23062 3426 23116 3442
rect 23263 3489 23338 3499
rect 23263 3455 23288 3489
rect 23322 3455 23338 3489
rect 23263 3445 23338 3455
rect 23380 3489 23435 3505
rect 23380 3455 23390 3489
rect 23424 3455 23435 3489
rect 22946 3382 22956 3416
rect 22990 3382 23010 3416
rect 22946 3366 23010 3382
rect 22980 3344 23010 3366
rect 23075 3356 23105 3426
rect 23263 3356 23293 3445
rect 23380 3439 23435 3455
rect 25656 3445 25686 3460
rect 23380 3401 23410 3439
rect 23347 3371 23410 3401
rect 25623 3415 25686 3445
rect 25623 3377 25653 3415
rect 23347 3356 23377 3371
rect 25598 3361 25653 3377
rect 25740 3371 25770 3460
rect 25598 3327 25609 3361
rect 25643 3327 25653 3361
rect 25598 3311 25653 3327
rect 25695 3361 25770 3371
rect 25928 3364 25958 3510
rect 26021 3376 26051 3510
rect 26105 3472 26135 3510
rect 26225 3478 26255 3510
rect 26093 3462 26159 3472
rect 26093 3428 26109 3462
rect 26143 3428 26159 3462
rect 26093 3418 26159 3428
rect 26225 3462 26289 3478
rect 26225 3428 26245 3462
rect 26279 3428 26289 3462
rect 26225 3412 26289 3428
rect 25695 3327 25711 3361
rect 25745 3327 25770 3361
rect 25695 3317 25770 3327
rect 25623 3273 25653 3311
rect 11575 3246 11605 3272
rect 11670 3246 11700 3272
rect 11858 3246 11888 3272
rect 11953 3246 11983 3272
rect 12141 3246 12171 3272
rect 12225 3246 12255 3272
rect 12343 3246 12373 3272
rect 12429 3246 12459 3272
rect 12524 3246 12554 3272
rect 12633 3246 12663 3272
rect 12728 3246 12758 3272
rect 12916 3246 12946 3272
rect 13000 3246 13030 3272
rect 13100 3246 13130 3272
rect 13210 3246 13240 3272
rect 13306 3246 13336 3272
rect 13412 3246 13442 3272
rect 13507 3246 13537 3272
rect 13695 3246 13725 3272
rect 13779 3246 13809 3272
rect 13967 3246 13997 3272
rect 14062 3246 14092 3272
rect 14250 3246 14280 3272
rect 14345 3246 14375 3272
rect 14533 3246 14563 3272
rect 14617 3246 14647 3272
rect 14735 3246 14765 3272
rect 14821 3246 14851 3272
rect 14916 3246 14946 3272
rect 15025 3246 15055 3272
rect 15120 3246 15150 3272
rect 15308 3246 15338 3272
rect 15392 3246 15422 3272
rect 15492 3246 15522 3272
rect 15602 3246 15632 3272
rect 15698 3246 15728 3272
rect 15804 3246 15834 3272
rect 15899 3246 15929 3272
rect 16087 3246 16117 3272
rect 16171 3246 16201 3272
rect 16359 3246 16389 3272
rect 16454 3246 16484 3272
rect 16642 3246 16672 3272
rect 16737 3246 16767 3272
rect 16925 3246 16955 3272
rect 17009 3246 17039 3272
rect 17127 3246 17157 3272
rect 17213 3246 17243 3272
rect 17308 3246 17338 3272
rect 17417 3246 17447 3272
rect 17512 3246 17542 3272
rect 17700 3246 17730 3272
rect 17784 3246 17814 3272
rect 17884 3246 17914 3272
rect 17994 3246 18024 3272
rect 18090 3246 18120 3272
rect 18196 3246 18226 3272
rect 18291 3246 18321 3272
rect 18479 3246 18509 3272
rect 18563 3246 18593 3272
rect 18751 3246 18781 3272
rect 18846 3246 18876 3272
rect 19034 3246 19064 3272
rect 19129 3246 19159 3272
rect 19317 3246 19347 3272
rect 19401 3246 19431 3272
rect 19519 3246 19549 3272
rect 19605 3246 19635 3272
rect 19700 3246 19730 3272
rect 19809 3246 19839 3272
rect 19904 3246 19934 3272
rect 20092 3246 20122 3272
rect 20176 3246 20206 3272
rect 20276 3246 20306 3272
rect 20386 3246 20416 3272
rect 20482 3246 20512 3272
rect 20588 3246 20618 3272
rect 20683 3246 20713 3272
rect 20871 3246 20901 3272
rect 20955 3246 20985 3272
rect 21143 3246 21173 3272
rect 21238 3246 21268 3272
rect 21426 3246 21456 3272
rect 21521 3246 21551 3272
rect 21709 3246 21739 3272
rect 21793 3246 21823 3272
rect 21911 3246 21941 3272
rect 21997 3246 22027 3272
rect 22092 3246 22122 3272
rect 22201 3246 22231 3272
rect 22296 3246 22326 3272
rect 22484 3246 22514 3272
rect 22568 3246 22598 3272
rect 22668 3246 22698 3272
rect 22778 3246 22808 3272
rect 22874 3246 22904 3272
rect 22980 3246 23010 3272
rect 23075 3246 23105 3272
rect 23263 3246 23293 3272
rect 23347 3246 23377 3272
rect 25623 3243 25686 3273
rect 25656 3228 25686 3243
rect 25740 3228 25770 3317
rect 25917 3348 25971 3364
rect 25917 3314 25927 3348
rect 25961 3314 25971 3348
rect 26021 3346 26159 3376
rect 25917 3298 25971 3314
rect 26129 3316 26159 3346
rect 25928 3228 25958 3298
rect 26023 3288 26087 3304
rect 26023 3254 26043 3288
rect 26077 3254 26087 3288
rect 26023 3238 26087 3254
rect 26129 3300 26183 3316
rect 26129 3266 26139 3300
rect 26173 3266 26183 3300
rect 26129 3250 26183 3266
rect 26023 3216 26053 3238
rect 26129 3216 26159 3250
rect 26225 3228 26255 3412
rect 26331 3326 26361 3510
rect 26804 3478 26834 3510
rect 26780 3462 26834 3478
rect 26888 3472 26918 3510
rect 27006 3478 27036 3510
rect 26780 3428 26790 3462
rect 26824 3428 26834 3462
rect 26439 3394 26469 3426
rect 26523 3394 26553 3426
rect 26403 3378 26469 3394
rect 26403 3344 26413 3378
rect 26447 3344 26469 3378
rect 26403 3328 26469 3344
rect 26519 3378 26609 3394
rect 26519 3344 26565 3378
rect 26599 3344 26609 3378
rect 26519 3328 26609 3344
rect 26660 3360 26690 3426
rect 26780 3412 26834 3428
rect 26876 3462 26942 3472
rect 26876 3428 26892 3462
rect 26926 3428 26942 3462
rect 26876 3418 26942 3428
rect 27006 3462 27072 3478
rect 27006 3428 27028 3462
rect 27062 3428 27072 3462
rect 26804 3376 26834 3412
rect 27006 3412 27072 3428
rect 26660 3344 26737 3360
rect 26804 3346 26941 3376
rect 26660 3330 26693 3344
rect 26301 3310 26361 3326
rect 26301 3276 26311 3310
rect 26345 3290 26361 3310
rect 26345 3276 26365 3290
rect 26301 3260 26365 3276
rect 26435 3272 26465 3328
rect 26519 3272 26549 3328
rect 26683 3310 26693 3330
rect 26727 3310 26737 3344
rect 26683 3294 26737 3310
rect 26707 3272 26737 3294
rect 26802 3288 26869 3304
rect 26335 3228 26365 3260
rect 26802 3254 26825 3288
rect 26859 3254 26869 3288
rect 26802 3238 26869 3254
rect 26802 3216 26832 3238
rect 26911 3216 26941 3346
rect 27006 3228 27036 3412
rect 27114 3326 27144 3510
rect 27480 3526 27510 3552
rect 27210 3378 27240 3426
rect 27078 3310 27144 3326
rect 27186 3362 27240 3378
rect 27282 3394 27312 3426
rect 27282 3378 27378 3394
rect 27282 3364 27334 3378
rect 27186 3328 27196 3362
rect 27230 3328 27240 3362
rect 27186 3312 27240 3328
rect 27078 3276 27088 3310
rect 27122 3276 27144 3310
rect 27078 3260 27144 3276
rect 27210 3272 27240 3312
rect 27294 3344 27334 3364
rect 27368 3344 27378 3378
rect 27480 3366 27510 3398
rect 27765 3578 27795 3604
rect 27860 3594 27890 3620
rect 27765 3434 27795 3450
rect 27739 3404 27795 3434
rect 27294 3328 27378 3344
rect 27449 3350 27513 3366
rect 27577 3362 27607 3394
rect 27294 3272 27324 3328
rect 27449 3316 27465 3350
rect 27499 3316 27513 3350
rect 27449 3300 27513 3316
rect 27555 3356 27607 3362
rect 27739 3356 27769 3404
rect 28048 3588 28078 3614
rect 28132 3588 28162 3614
rect 28320 3594 28350 3620
rect 28413 3594 28443 3620
rect 28497 3594 28527 3620
rect 28617 3594 28647 3620
rect 28723 3594 28753 3620
rect 28831 3594 28861 3620
rect 28915 3594 28945 3620
rect 29052 3594 29082 3620
rect 29196 3594 29226 3620
rect 29280 3594 29310 3620
rect 29398 3594 29428 3620
rect 29506 3594 29536 3620
rect 29602 3594 29632 3620
rect 29674 3594 29704 3620
rect 29969 3594 29999 3620
rect 28048 3445 28078 3460
rect 28015 3415 28078 3445
rect 27860 3362 27890 3394
rect 28015 3377 28045 3415
rect 27555 3346 27769 3356
rect 27555 3312 27565 3346
rect 27599 3312 27769 3346
rect 27555 3302 27769 3312
rect 27092 3228 27122 3260
rect 27482 3228 27512 3300
rect 27555 3296 27607 3302
rect 27577 3274 27607 3296
rect 27739 3273 27769 3302
rect 27831 3346 27890 3362
rect 27831 3312 27841 3346
rect 27875 3312 27890 3346
rect 27831 3296 27890 3312
rect 27990 3361 28045 3377
rect 28132 3371 28162 3460
rect 27990 3327 28001 3361
rect 28035 3327 28045 3361
rect 27990 3311 28045 3327
rect 28087 3361 28162 3371
rect 28320 3364 28350 3510
rect 28413 3376 28443 3510
rect 28497 3472 28527 3510
rect 28617 3478 28647 3510
rect 28485 3462 28551 3472
rect 28485 3428 28501 3462
rect 28535 3428 28551 3462
rect 28485 3418 28551 3428
rect 28617 3462 28681 3478
rect 28617 3428 28637 3462
rect 28671 3428 28681 3462
rect 28617 3412 28681 3428
rect 28087 3327 28103 3361
rect 28137 3327 28162 3361
rect 28087 3317 28162 3327
rect 27860 3274 27890 3296
rect 27739 3243 27795 3273
rect 27765 3228 27795 3243
rect 28015 3273 28045 3311
rect 28015 3243 28078 3273
rect 28048 3228 28078 3243
rect 28132 3228 28162 3317
rect 28309 3348 28363 3364
rect 28309 3314 28319 3348
rect 28353 3314 28363 3348
rect 28413 3346 28551 3376
rect 28309 3298 28363 3314
rect 28521 3316 28551 3346
rect 28320 3228 28350 3298
rect 28415 3288 28479 3304
rect 28415 3254 28435 3288
rect 28469 3254 28479 3288
rect 28415 3238 28479 3254
rect 28521 3300 28575 3316
rect 28521 3266 28531 3300
rect 28565 3266 28575 3300
rect 28521 3250 28575 3266
rect 28415 3216 28445 3238
rect 28521 3216 28551 3250
rect 28617 3228 28647 3412
rect 28723 3326 28753 3510
rect 29196 3478 29226 3510
rect 29172 3462 29226 3478
rect 29280 3472 29310 3510
rect 29398 3478 29428 3510
rect 29172 3428 29182 3462
rect 29216 3428 29226 3462
rect 28831 3394 28861 3426
rect 28915 3394 28945 3426
rect 28795 3378 28861 3394
rect 28795 3344 28805 3378
rect 28839 3344 28861 3378
rect 28795 3328 28861 3344
rect 28911 3378 29001 3394
rect 28911 3344 28957 3378
rect 28991 3344 29001 3378
rect 28911 3328 29001 3344
rect 29052 3360 29082 3426
rect 29172 3412 29226 3428
rect 29268 3462 29334 3472
rect 29268 3428 29284 3462
rect 29318 3428 29334 3462
rect 29268 3418 29334 3428
rect 29398 3462 29464 3478
rect 29398 3428 29420 3462
rect 29454 3428 29464 3462
rect 29196 3376 29226 3412
rect 29398 3412 29464 3428
rect 29052 3344 29129 3360
rect 29196 3346 29333 3376
rect 29052 3330 29085 3344
rect 28693 3310 28753 3326
rect 28693 3276 28703 3310
rect 28737 3290 28753 3310
rect 28737 3276 28757 3290
rect 28693 3260 28757 3276
rect 28827 3272 28857 3328
rect 28911 3272 28941 3328
rect 29075 3310 29085 3330
rect 29119 3310 29129 3344
rect 29075 3294 29129 3310
rect 29099 3272 29129 3294
rect 29194 3288 29261 3304
rect 28727 3228 28757 3260
rect 29194 3254 29217 3288
rect 29251 3254 29261 3288
rect 29194 3238 29261 3254
rect 29194 3216 29224 3238
rect 29303 3216 29333 3346
rect 29398 3228 29428 3412
rect 29506 3326 29536 3510
rect 29872 3526 29902 3552
rect 29602 3378 29632 3426
rect 29470 3310 29536 3326
rect 29578 3362 29632 3378
rect 29674 3394 29704 3426
rect 29674 3378 29770 3394
rect 29674 3364 29726 3378
rect 29578 3328 29588 3362
rect 29622 3328 29632 3362
rect 29578 3312 29632 3328
rect 29470 3276 29480 3310
rect 29514 3276 29536 3310
rect 29470 3260 29536 3276
rect 29602 3272 29632 3312
rect 29686 3344 29726 3364
rect 29760 3344 29770 3378
rect 29872 3366 29902 3398
rect 30157 3578 30187 3604
rect 30252 3594 30282 3620
rect 30157 3434 30187 3450
rect 30131 3404 30187 3434
rect 29686 3328 29770 3344
rect 29841 3350 29905 3366
rect 29969 3362 29999 3394
rect 29686 3272 29716 3328
rect 29841 3316 29857 3350
rect 29891 3316 29905 3350
rect 29841 3300 29905 3316
rect 29947 3356 29999 3362
rect 30131 3356 30161 3404
rect 30252 3362 30282 3394
rect 29947 3346 30161 3356
rect 29947 3312 29957 3346
rect 29991 3312 30161 3346
rect 29947 3302 30161 3312
rect 29484 3228 29514 3260
rect 29874 3228 29904 3300
rect 29947 3296 29999 3302
rect 29969 3274 29999 3296
rect 30131 3273 30161 3302
rect 30223 3346 30282 3362
rect 30223 3312 30233 3346
rect 30267 3312 30282 3346
rect 30223 3296 30282 3312
rect 30252 3274 30282 3296
rect 30131 3243 30187 3273
rect 30157 3228 30187 3243
rect 25656 3118 25686 3144
rect 25740 3118 25770 3144
rect 25928 3118 25958 3144
rect 26023 3118 26053 3144
rect 26129 3118 26159 3144
rect 26225 3118 26255 3144
rect 26335 3118 26365 3144
rect 26435 3118 26465 3144
rect 26519 3118 26549 3144
rect 26707 3118 26737 3144
rect 26802 3118 26832 3144
rect 26911 3118 26941 3144
rect 27006 3118 27036 3144
rect 27092 3118 27122 3144
rect 27210 3118 27240 3144
rect 27294 3118 27324 3144
rect 27482 3118 27512 3144
rect 27577 3118 27607 3144
rect 27765 3118 27795 3144
rect 27860 3118 27890 3144
rect 28048 3118 28078 3144
rect 28132 3118 28162 3144
rect 28320 3118 28350 3144
rect 28415 3118 28445 3144
rect 28521 3118 28551 3144
rect 28617 3118 28647 3144
rect 28727 3118 28757 3144
rect 28827 3118 28857 3144
rect 28911 3118 28941 3144
rect 29099 3118 29129 3144
rect 29194 3118 29224 3144
rect 29303 3118 29333 3144
rect 29398 3118 29428 3144
rect 29484 3118 29514 3144
rect 29602 3118 29632 3144
rect 29686 3118 29716 3144
rect 29874 3118 29904 3144
rect 29969 3118 29999 3144
rect 30157 3118 30187 3144
rect 30252 3118 30282 3144
rect 25656 2954 25686 2980
rect 25740 2954 25770 2980
rect 25928 2954 25958 2980
rect 26023 2954 26053 2980
rect 26129 2954 26159 2980
rect 26225 2954 26255 2980
rect 26335 2954 26365 2980
rect 26435 2954 26465 2980
rect 26519 2954 26549 2980
rect 26707 2954 26737 2980
rect 26802 2954 26832 2980
rect 26911 2954 26941 2980
rect 27006 2954 27036 2980
rect 27092 2954 27122 2980
rect 27210 2954 27240 2980
rect 27294 2954 27324 2980
rect 27482 2954 27512 2980
rect 27577 2954 27607 2980
rect 27765 2954 27795 2980
rect 27860 2954 27890 2980
rect 28048 2954 28078 2980
rect 28132 2954 28162 2980
rect 28320 2954 28350 2980
rect 28415 2954 28445 2980
rect 28521 2954 28551 2980
rect 28617 2954 28647 2980
rect 28727 2954 28757 2980
rect 28827 2954 28857 2980
rect 28911 2954 28941 2980
rect 29099 2954 29129 2980
rect 29194 2954 29224 2980
rect 29303 2954 29333 2980
rect 29398 2954 29428 2980
rect 29484 2954 29514 2980
rect 29602 2954 29632 2980
rect 29686 2954 29716 2980
rect 29874 2954 29904 2980
rect 29969 2954 29999 2980
rect 30157 2954 30187 2980
rect 30252 2954 30282 2980
rect 25656 2855 25686 2870
rect 25623 2825 25686 2855
rect 25623 2787 25653 2825
rect 25598 2771 25653 2787
rect 25740 2781 25770 2870
rect 25928 2800 25958 2870
rect 26023 2860 26053 2882
rect 26023 2844 26087 2860
rect 26023 2810 26043 2844
rect 26077 2810 26087 2844
rect 25598 2737 25609 2771
rect 25643 2737 25653 2771
rect 25598 2721 25653 2737
rect 25695 2771 25770 2781
rect 25695 2737 25711 2771
rect 25745 2737 25770 2771
rect 25695 2727 25770 2737
rect 25917 2784 25971 2800
rect 26023 2794 26087 2810
rect 26129 2848 26159 2882
rect 26129 2832 26183 2848
rect 26129 2798 26139 2832
rect 26173 2798 26183 2832
rect 25917 2750 25927 2784
rect 25961 2750 25971 2784
rect 26129 2782 26183 2798
rect 26129 2752 26159 2782
rect 25917 2734 25971 2750
rect 25623 2683 25653 2721
rect 25623 2653 25686 2683
rect 25656 2638 25686 2653
rect 25740 2638 25770 2727
rect 25928 2588 25958 2734
rect 26021 2722 26159 2752
rect 26021 2588 26051 2722
rect 26225 2686 26255 2870
rect 26335 2838 26365 2870
rect 26301 2822 26365 2838
rect 26802 2860 26832 2882
rect 26802 2844 26869 2860
rect 26301 2788 26311 2822
rect 26345 2808 26365 2822
rect 26345 2788 26361 2808
rect 26301 2772 26361 2788
rect 26093 2670 26159 2680
rect 26093 2636 26109 2670
rect 26143 2636 26159 2670
rect 26093 2626 26159 2636
rect 26225 2670 26289 2686
rect 26225 2636 26245 2670
rect 26279 2636 26289 2670
rect 26105 2588 26135 2626
rect 26225 2620 26289 2636
rect 26225 2588 26255 2620
rect 26331 2588 26361 2772
rect 26435 2770 26465 2826
rect 26519 2770 26549 2826
rect 26707 2804 26737 2826
rect 26683 2788 26737 2804
rect 26802 2810 26825 2844
rect 26859 2810 26869 2844
rect 26802 2794 26869 2810
rect 26403 2754 26469 2770
rect 26403 2720 26413 2754
rect 26447 2720 26469 2754
rect 26403 2704 26469 2720
rect 26519 2754 26609 2770
rect 26683 2768 26693 2788
rect 26519 2720 26565 2754
rect 26599 2720 26609 2754
rect 26519 2704 26609 2720
rect 26660 2754 26693 2768
rect 26727 2754 26737 2788
rect 26660 2738 26737 2754
rect 26911 2752 26941 2882
rect 26439 2672 26469 2704
rect 26523 2672 26553 2704
rect 26660 2672 26690 2738
rect 26804 2722 26941 2752
rect 26804 2686 26834 2722
rect 25656 2484 25686 2510
rect 25740 2484 25770 2510
rect 26780 2670 26834 2686
rect 27006 2686 27036 2870
rect 27092 2838 27122 2870
rect 27078 2822 27144 2838
rect 27078 2788 27088 2822
rect 27122 2788 27144 2822
rect 27078 2772 27144 2788
rect 27210 2786 27240 2826
rect 26780 2636 26790 2670
rect 26824 2636 26834 2670
rect 26780 2620 26834 2636
rect 26876 2670 26942 2680
rect 26876 2636 26892 2670
rect 26926 2636 26942 2670
rect 26876 2626 26942 2636
rect 27006 2670 27072 2686
rect 27006 2636 27028 2670
rect 27062 2636 27072 2670
rect 26804 2588 26834 2620
rect 26888 2588 26918 2626
rect 27006 2620 27072 2636
rect 27006 2588 27036 2620
rect 27114 2588 27144 2772
rect 27186 2770 27240 2786
rect 27186 2736 27196 2770
rect 27230 2736 27240 2770
rect 27186 2720 27240 2736
rect 27294 2770 27324 2826
rect 27482 2798 27512 2870
rect 27765 2855 27795 2870
rect 27739 2825 27795 2855
rect 27577 2802 27607 2824
rect 27449 2782 27513 2798
rect 27294 2754 27378 2770
rect 27294 2734 27334 2754
rect 27210 2672 27240 2720
rect 27282 2720 27334 2734
rect 27368 2720 27378 2754
rect 27449 2748 27465 2782
rect 27499 2748 27513 2782
rect 27449 2732 27513 2748
rect 27555 2796 27607 2802
rect 27739 2796 27769 2825
rect 28048 2855 28078 2870
rect 28015 2825 28078 2855
rect 27860 2802 27890 2824
rect 27555 2786 27769 2796
rect 27555 2752 27565 2786
rect 27599 2752 27769 2786
rect 27555 2742 27769 2752
rect 27555 2736 27607 2742
rect 27282 2704 27378 2720
rect 27282 2672 27312 2704
rect 27480 2700 27510 2732
rect 27577 2704 27607 2736
rect 27480 2546 27510 2572
rect 27739 2694 27769 2742
rect 27831 2786 27890 2802
rect 28015 2787 28045 2825
rect 27831 2752 27841 2786
rect 27875 2752 27890 2786
rect 27831 2736 27890 2752
rect 27860 2704 27890 2736
rect 27990 2771 28045 2787
rect 28132 2781 28162 2870
rect 28320 2800 28350 2870
rect 28415 2860 28445 2882
rect 28415 2844 28479 2860
rect 28415 2810 28435 2844
rect 28469 2810 28479 2844
rect 27990 2737 28001 2771
rect 28035 2737 28045 2771
rect 27990 2721 28045 2737
rect 28087 2771 28162 2781
rect 28087 2737 28103 2771
rect 28137 2737 28162 2771
rect 28087 2727 28162 2737
rect 28309 2784 28363 2800
rect 28415 2794 28479 2810
rect 28521 2848 28551 2882
rect 28521 2832 28575 2848
rect 28521 2798 28531 2832
rect 28565 2798 28575 2832
rect 28309 2750 28319 2784
rect 28353 2750 28363 2784
rect 28521 2782 28575 2798
rect 28521 2752 28551 2782
rect 28309 2734 28363 2750
rect 27739 2664 27795 2694
rect 27765 2648 27795 2664
rect 25928 2478 25958 2504
rect 26021 2478 26051 2504
rect 26105 2478 26135 2504
rect 26225 2478 26255 2504
rect 26331 2478 26361 2504
rect 26439 2478 26469 2504
rect 26523 2478 26553 2504
rect 26660 2478 26690 2504
rect 26804 2478 26834 2504
rect 26888 2478 26918 2504
rect 27006 2478 27036 2504
rect 27114 2478 27144 2504
rect 27210 2478 27240 2504
rect 27282 2478 27312 2504
rect 27577 2478 27607 2504
rect 27765 2494 27795 2520
rect 28015 2683 28045 2721
rect 28015 2653 28078 2683
rect 28048 2638 28078 2653
rect 28132 2638 28162 2727
rect 28320 2588 28350 2734
rect 28413 2722 28551 2752
rect 28413 2588 28443 2722
rect 28617 2686 28647 2870
rect 28727 2838 28757 2870
rect 28693 2822 28757 2838
rect 29194 2860 29224 2882
rect 29194 2844 29261 2860
rect 28693 2788 28703 2822
rect 28737 2808 28757 2822
rect 28737 2788 28753 2808
rect 28693 2772 28753 2788
rect 28485 2670 28551 2680
rect 28485 2636 28501 2670
rect 28535 2636 28551 2670
rect 28485 2626 28551 2636
rect 28617 2670 28681 2686
rect 28617 2636 28637 2670
rect 28671 2636 28681 2670
rect 28497 2588 28527 2626
rect 28617 2620 28681 2636
rect 28617 2588 28647 2620
rect 28723 2588 28753 2772
rect 28827 2770 28857 2826
rect 28911 2770 28941 2826
rect 29099 2804 29129 2826
rect 29075 2788 29129 2804
rect 29194 2810 29217 2844
rect 29251 2810 29261 2844
rect 29194 2794 29261 2810
rect 28795 2754 28861 2770
rect 28795 2720 28805 2754
rect 28839 2720 28861 2754
rect 28795 2704 28861 2720
rect 28911 2754 29001 2770
rect 29075 2768 29085 2788
rect 28911 2720 28957 2754
rect 28991 2720 29001 2754
rect 28911 2704 29001 2720
rect 29052 2754 29085 2768
rect 29119 2754 29129 2788
rect 29052 2738 29129 2754
rect 29303 2752 29333 2882
rect 28831 2672 28861 2704
rect 28915 2672 28945 2704
rect 29052 2672 29082 2738
rect 29196 2722 29333 2752
rect 29196 2686 29226 2722
rect 27860 2478 27890 2504
rect 28048 2484 28078 2510
rect 28132 2484 28162 2510
rect 29172 2670 29226 2686
rect 29398 2686 29428 2870
rect 29484 2838 29514 2870
rect 29470 2822 29536 2838
rect 29470 2788 29480 2822
rect 29514 2788 29536 2822
rect 29470 2772 29536 2788
rect 29602 2786 29632 2826
rect 29172 2636 29182 2670
rect 29216 2636 29226 2670
rect 29172 2620 29226 2636
rect 29268 2670 29334 2680
rect 29268 2636 29284 2670
rect 29318 2636 29334 2670
rect 29268 2626 29334 2636
rect 29398 2670 29464 2686
rect 29398 2636 29420 2670
rect 29454 2636 29464 2670
rect 29196 2588 29226 2620
rect 29280 2588 29310 2626
rect 29398 2620 29464 2636
rect 29398 2588 29428 2620
rect 29506 2588 29536 2772
rect 29578 2770 29632 2786
rect 29578 2736 29588 2770
rect 29622 2736 29632 2770
rect 29578 2720 29632 2736
rect 29686 2770 29716 2826
rect 29874 2798 29904 2870
rect 30157 2855 30187 2870
rect 30131 2825 30187 2855
rect 29969 2802 29999 2824
rect 29841 2782 29905 2798
rect 29686 2754 29770 2770
rect 29686 2734 29726 2754
rect 29602 2672 29632 2720
rect 29674 2720 29726 2734
rect 29760 2720 29770 2754
rect 29841 2748 29857 2782
rect 29891 2748 29905 2782
rect 29841 2732 29905 2748
rect 29947 2796 29999 2802
rect 30131 2796 30161 2825
rect 30252 2802 30282 2824
rect 29947 2786 30161 2796
rect 29947 2752 29957 2786
rect 29991 2752 30161 2786
rect 29947 2742 30161 2752
rect 29947 2736 29999 2742
rect 29674 2704 29770 2720
rect 29674 2672 29704 2704
rect 29872 2700 29902 2732
rect 29969 2704 29999 2736
rect 29872 2546 29902 2572
rect 30131 2694 30161 2742
rect 30223 2786 30282 2802
rect 30223 2752 30233 2786
rect 30267 2752 30282 2786
rect 30223 2736 30282 2752
rect 30252 2704 30282 2736
rect 30131 2664 30187 2694
rect 30157 2648 30187 2664
rect 28320 2478 28350 2504
rect 28413 2478 28443 2504
rect 28497 2478 28527 2504
rect 28617 2478 28647 2504
rect 28723 2478 28753 2504
rect 28831 2478 28861 2504
rect 28915 2478 28945 2504
rect 29052 2478 29082 2504
rect 29196 2478 29226 2504
rect 29280 2478 29310 2504
rect 29398 2478 29428 2504
rect 29506 2478 29536 2504
rect 29602 2478 29632 2504
rect 29674 2478 29704 2504
rect 29969 2478 29999 2504
rect 30157 2494 30187 2520
rect 30252 2478 30282 2504
rect 25656 2308 25686 2334
rect 25740 2308 25770 2334
rect 25928 2314 25958 2340
rect 26021 2314 26051 2340
rect 26105 2314 26135 2340
rect 26225 2314 26255 2340
rect 26331 2314 26361 2340
rect 26439 2314 26469 2340
rect 26523 2314 26553 2340
rect 26660 2314 26690 2340
rect 26804 2314 26834 2340
rect 26888 2314 26918 2340
rect 27006 2314 27036 2340
rect 27114 2314 27144 2340
rect 27210 2314 27240 2340
rect 27282 2314 27312 2340
rect 27577 2314 27607 2340
rect 25656 2165 25686 2180
rect 25623 2135 25686 2165
rect 25623 2097 25653 2135
rect 25598 2081 25653 2097
rect 25740 2091 25770 2180
rect 25598 2047 25609 2081
rect 25643 2047 25653 2081
rect 25598 2031 25653 2047
rect 25695 2081 25770 2091
rect 25928 2084 25958 2230
rect 26021 2096 26051 2230
rect 26105 2192 26135 2230
rect 26225 2198 26255 2230
rect 26093 2182 26159 2192
rect 26093 2148 26109 2182
rect 26143 2148 26159 2182
rect 26093 2138 26159 2148
rect 26225 2182 26289 2198
rect 26225 2148 26245 2182
rect 26279 2148 26289 2182
rect 26225 2132 26289 2148
rect 25695 2047 25711 2081
rect 25745 2047 25770 2081
rect 25695 2037 25770 2047
rect 25623 1993 25653 2031
rect 25623 1963 25686 1993
rect 25656 1948 25686 1963
rect 25740 1948 25770 2037
rect 25917 2068 25971 2084
rect 25917 2034 25927 2068
rect 25961 2034 25971 2068
rect 26021 2066 26159 2096
rect 25917 2018 25971 2034
rect 26129 2036 26159 2066
rect 25928 1948 25958 2018
rect 26023 2008 26087 2024
rect 26023 1974 26043 2008
rect 26077 1974 26087 2008
rect 26023 1958 26087 1974
rect 26129 2020 26183 2036
rect 26129 1986 26139 2020
rect 26173 1986 26183 2020
rect 26129 1970 26183 1986
rect 26023 1936 26053 1958
rect 26129 1936 26159 1970
rect 26225 1948 26255 2132
rect 26331 2046 26361 2230
rect 26804 2198 26834 2230
rect 26780 2182 26834 2198
rect 26888 2192 26918 2230
rect 27006 2198 27036 2230
rect 26780 2148 26790 2182
rect 26824 2148 26834 2182
rect 26439 2114 26469 2146
rect 26523 2114 26553 2146
rect 26403 2098 26469 2114
rect 26403 2064 26413 2098
rect 26447 2064 26469 2098
rect 26403 2048 26469 2064
rect 26519 2098 26609 2114
rect 26519 2064 26565 2098
rect 26599 2064 26609 2098
rect 26519 2048 26609 2064
rect 26660 2080 26690 2146
rect 26780 2132 26834 2148
rect 26876 2182 26942 2192
rect 26876 2148 26892 2182
rect 26926 2148 26942 2182
rect 26876 2138 26942 2148
rect 27006 2182 27072 2198
rect 27006 2148 27028 2182
rect 27062 2148 27072 2182
rect 26804 2096 26834 2132
rect 27006 2132 27072 2148
rect 26660 2064 26737 2080
rect 26804 2066 26941 2096
rect 26660 2050 26693 2064
rect 26301 2030 26361 2046
rect 26301 1996 26311 2030
rect 26345 2010 26361 2030
rect 26345 1996 26365 2010
rect 26301 1980 26365 1996
rect 26435 1992 26465 2048
rect 26519 1992 26549 2048
rect 26683 2030 26693 2050
rect 26727 2030 26737 2064
rect 26683 2014 26737 2030
rect 26707 1992 26737 2014
rect 26802 2008 26869 2024
rect 26335 1948 26365 1980
rect 26802 1974 26825 2008
rect 26859 1974 26869 2008
rect 26802 1958 26869 1974
rect 26802 1936 26832 1958
rect 26911 1936 26941 2066
rect 27006 1948 27036 2132
rect 27114 2046 27144 2230
rect 27480 2246 27510 2272
rect 27210 2098 27240 2146
rect 27078 2030 27144 2046
rect 27186 2082 27240 2098
rect 27282 2114 27312 2146
rect 27282 2098 27378 2114
rect 27282 2084 27334 2098
rect 27186 2048 27196 2082
rect 27230 2048 27240 2082
rect 27186 2032 27240 2048
rect 27078 1996 27088 2030
rect 27122 1996 27144 2030
rect 27078 1980 27144 1996
rect 27210 1992 27240 2032
rect 27294 2064 27334 2084
rect 27368 2064 27378 2098
rect 27480 2086 27510 2118
rect 27765 2298 27795 2324
rect 27860 2314 27890 2340
rect 27765 2154 27795 2170
rect 27739 2124 27795 2154
rect 27294 2048 27378 2064
rect 27449 2070 27513 2086
rect 27577 2082 27607 2114
rect 27294 1992 27324 2048
rect 27449 2036 27465 2070
rect 27499 2036 27513 2070
rect 27449 2020 27513 2036
rect 27555 2076 27607 2082
rect 27739 2076 27769 2124
rect 28048 2308 28078 2334
rect 28132 2308 28162 2334
rect 28320 2314 28350 2340
rect 28413 2314 28443 2340
rect 28497 2314 28527 2340
rect 28617 2314 28647 2340
rect 28723 2314 28753 2340
rect 28831 2314 28861 2340
rect 28915 2314 28945 2340
rect 29052 2314 29082 2340
rect 29196 2314 29226 2340
rect 29280 2314 29310 2340
rect 29398 2314 29428 2340
rect 29506 2314 29536 2340
rect 29602 2314 29632 2340
rect 29674 2314 29704 2340
rect 29969 2314 29999 2340
rect 28048 2165 28078 2180
rect 28015 2135 28078 2165
rect 27860 2082 27890 2114
rect 28015 2097 28045 2135
rect 27555 2066 27769 2076
rect 27555 2032 27565 2066
rect 27599 2032 27769 2066
rect 27555 2022 27769 2032
rect 27092 1948 27122 1980
rect 27482 1948 27512 2020
rect 27555 2016 27607 2022
rect 27577 1994 27607 2016
rect 27739 1993 27769 2022
rect 27831 2066 27890 2082
rect 27831 2032 27841 2066
rect 27875 2032 27890 2066
rect 27831 2016 27890 2032
rect 27990 2081 28045 2097
rect 28132 2091 28162 2180
rect 27990 2047 28001 2081
rect 28035 2047 28045 2081
rect 27990 2031 28045 2047
rect 28087 2081 28162 2091
rect 28320 2084 28350 2230
rect 28413 2096 28443 2230
rect 28497 2192 28527 2230
rect 28617 2198 28647 2230
rect 28485 2182 28551 2192
rect 28485 2148 28501 2182
rect 28535 2148 28551 2182
rect 28485 2138 28551 2148
rect 28617 2182 28681 2198
rect 28617 2148 28637 2182
rect 28671 2148 28681 2182
rect 28617 2132 28681 2148
rect 28087 2047 28103 2081
rect 28137 2047 28162 2081
rect 28087 2037 28162 2047
rect 27860 1994 27890 2016
rect 27739 1963 27795 1993
rect 27765 1948 27795 1963
rect 28015 1993 28045 2031
rect 28015 1963 28078 1993
rect 28048 1948 28078 1963
rect 28132 1948 28162 2037
rect 28309 2068 28363 2084
rect 28309 2034 28319 2068
rect 28353 2034 28363 2068
rect 28413 2066 28551 2096
rect 28309 2018 28363 2034
rect 28521 2036 28551 2066
rect 28320 1948 28350 2018
rect 28415 2008 28479 2024
rect 28415 1974 28435 2008
rect 28469 1974 28479 2008
rect 28415 1958 28479 1974
rect 28521 2020 28575 2036
rect 28521 1986 28531 2020
rect 28565 1986 28575 2020
rect 28521 1970 28575 1986
rect 28415 1936 28445 1958
rect 28521 1936 28551 1970
rect 28617 1948 28647 2132
rect 28723 2046 28753 2230
rect 29196 2198 29226 2230
rect 29172 2182 29226 2198
rect 29280 2192 29310 2230
rect 29398 2198 29428 2230
rect 29172 2148 29182 2182
rect 29216 2148 29226 2182
rect 28831 2114 28861 2146
rect 28915 2114 28945 2146
rect 28795 2098 28861 2114
rect 28795 2064 28805 2098
rect 28839 2064 28861 2098
rect 28795 2048 28861 2064
rect 28911 2098 29001 2114
rect 28911 2064 28957 2098
rect 28991 2064 29001 2098
rect 28911 2048 29001 2064
rect 29052 2080 29082 2146
rect 29172 2132 29226 2148
rect 29268 2182 29334 2192
rect 29268 2148 29284 2182
rect 29318 2148 29334 2182
rect 29268 2138 29334 2148
rect 29398 2182 29464 2198
rect 29398 2148 29420 2182
rect 29454 2148 29464 2182
rect 29196 2096 29226 2132
rect 29398 2132 29464 2148
rect 29052 2064 29129 2080
rect 29196 2066 29333 2096
rect 29052 2050 29085 2064
rect 28693 2030 28753 2046
rect 28693 1996 28703 2030
rect 28737 2010 28753 2030
rect 28737 1996 28757 2010
rect 28693 1980 28757 1996
rect 28827 1992 28857 2048
rect 28911 1992 28941 2048
rect 29075 2030 29085 2050
rect 29119 2030 29129 2064
rect 29075 2014 29129 2030
rect 29099 1992 29129 2014
rect 29194 2008 29261 2024
rect 28727 1948 28757 1980
rect 29194 1974 29217 2008
rect 29251 1974 29261 2008
rect 29194 1958 29261 1974
rect 29194 1936 29224 1958
rect 29303 1936 29333 2066
rect 29398 1948 29428 2132
rect 29506 2046 29536 2230
rect 29872 2246 29902 2272
rect 29602 2098 29632 2146
rect 29470 2030 29536 2046
rect 29578 2082 29632 2098
rect 29674 2114 29704 2146
rect 29674 2098 29770 2114
rect 29674 2084 29726 2098
rect 29578 2048 29588 2082
rect 29622 2048 29632 2082
rect 29578 2032 29632 2048
rect 29470 1996 29480 2030
rect 29514 1996 29536 2030
rect 29470 1980 29536 1996
rect 29602 1992 29632 2032
rect 29686 2064 29726 2084
rect 29760 2064 29770 2098
rect 29872 2086 29902 2118
rect 30157 2298 30187 2324
rect 30252 2314 30282 2340
rect 30157 2154 30187 2170
rect 30131 2124 30187 2154
rect 29686 2048 29770 2064
rect 29841 2070 29905 2086
rect 29969 2082 29999 2114
rect 29686 1992 29716 2048
rect 29841 2036 29857 2070
rect 29891 2036 29905 2070
rect 29841 2020 29905 2036
rect 29947 2076 29999 2082
rect 30131 2076 30161 2124
rect 30252 2082 30282 2114
rect 29947 2066 30161 2076
rect 29947 2032 29957 2066
rect 29991 2032 30161 2066
rect 29947 2022 30161 2032
rect 29484 1948 29514 1980
rect 29874 1948 29904 2020
rect 29947 2016 29999 2022
rect 29969 1994 29999 2016
rect 30131 1993 30161 2022
rect 30223 2066 30282 2082
rect 30223 2032 30233 2066
rect 30267 2032 30282 2066
rect 30223 2016 30282 2032
rect 30252 1994 30282 2016
rect 30131 1963 30187 1993
rect 30157 1948 30187 1963
rect 25656 1838 25686 1864
rect 25740 1838 25770 1864
rect 25928 1838 25958 1864
rect 26023 1838 26053 1864
rect 26129 1838 26159 1864
rect 26225 1838 26255 1864
rect 26335 1838 26365 1864
rect 26435 1838 26465 1864
rect 26519 1838 26549 1864
rect 26707 1838 26737 1864
rect 26802 1838 26832 1864
rect 26911 1838 26941 1864
rect 27006 1838 27036 1864
rect 27092 1838 27122 1864
rect 27210 1838 27240 1864
rect 27294 1838 27324 1864
rect 27482 1838 27512 1864
rect 27577 1838 27607 1864
rect 27765 1838 27795 1864
rect 27860 1838 27890 1864
rect 28048 1838 28078 1864
rect 28132 1838 28162 1864
rect 28320 1838 28350 1864
rect 28415 1838 28445 1864
rect 28521 1838 28551 1864
rect 28617 1838 28647 1864
rect 28727 1838 28757 1864
rect 28827 1838 28857 1864
rect 28911 1838 28941 1864
rect 29099 1838 29129 1864
rect 29194 1838 29224 1864
rect 29303 1838 29333 1864
rect 29398 1838 29428 1864
rect 29484 1838 29514 1864
rect 29602 1838 29632 1864
rect 29686 1838 29716 1864
rect 29874 1838 29904 1864
rect 29969 1838 29999 1864
rect 30157 1838 30187 1864
rect 30252 1838 30282 1864
rect 8656 1342 8686 1368
rect 8744 1342 8774 1368
rect 8932 1342 8962 1368
rect 9016 1342 9046 1368
rect 9100 1342 9130 1368
rect 9184 1342 9214 1368
rect 9268 1342 9298 1368
rect 9484 1342 9514 1368
rect 9568 1342 9598 1368
rect 9652 1342 9682 1368
rect 9736 1342 9766 1368
rect 9820 1342 9850 1368
rect 9904 1342 9934 1368
rect 9988 1342 10018 1368
rect 10072 1342 10102 1368
rect 10156 1342 10186 1368
rect 10240 1342 10270 1368
rect 10324 1342 10354 1368
rect 10408 1342 10438 1368
rect 10492 1342 10522 1368
rect 10576 1342 10606 1368
rect 10660 1342 10690 1368
rect 10744 1342 10774 1368
rect 10828 1342 10858 1368
rect 10912 1342 10942 1368
rect 10996 1342 11026 1368
rect 11080 1342 11110 1368
rect 11164 1342 11194 1368
rect 11248 1342 11278 1368
rect 13040 1342 13070 1368
rect 13128 1342 13158 1368
rect 13316 1342 13346 1368
rect 13400 1342 13430 1368
rect 13484 1342 13514 1368
rect 13568 1342 13598 1368
rect 13652 1342 13682 1368
rect 13868 1342 13898 1368
rect 13952 1342 13982 1368
rect 14036 1342 14066 1368
rect 14120 1342 14150 1368
rect 14204 1342 14234 1368
rect 14288 1342 14318 1368
rect 14372 1342 14402 1368
rect 14456 1342 14486 1368
rect 14540 1342 14570 1368
rect 14624 1342 14654 1368
rect 14708 1342 14738 1368
rect 14792 1342 14822 1368
rect 14876 1342 14906 1368
rect 14960 1342 14990 1368
rect 15044 1342 15074 1368
rect 15128 1342 15158 1368
rect 15212 1342 15242 1368
rect 15296 1342 15326 1368
rect 15380 1342 15410 1368
rect 15464 1342 15494 1368
rect 15548 1342 15578 1368
rect 15632 1342 15662 1368
rect 8656 1169 8686 1184
rect 8650 1145 8686 1169
rect 8650 1110 8680 1145
rect 8744 1123 8774 1184
rect 13040 1169 13070 1184
rect 13034 1145 13070 1169
rect 8604 1094 8680 1110
rect 8604 1060 8614 1094
rect 8648 1060 8680 1094
rect 8604 1044 8680 1060
rect 8722 1107 8776 1123
rect 8722 1073 8732 1107
rect 8766 1073 8776 1107
rect 8932 1106 8962 1142
rect 8722 1057 8776 1073
rect 8881 1094 8962 1106
rect 9016 1104 9046 1142
rect 9100 1104 9130 1142
rect 9184 1104 9214 1142
rect 9268 1104 9298 1142
rect 8881 1060 8897 1094
rect 8931 1060 8962 1094
rect 8650 1035 8680 1044
rect 8650 1011 8686 1035
rect 8656 996 8686 1011
rect 8744 996 8774 1057
rect 8881 1048 8962 1060
rect 9015 1094 9298 1104
rect 9015 1060 9031 1094
rect 9065 1060 9298 1094
rect 9015 1050 9298 1060
rect 8932 1022 8962 1048
rect 9016 1022 9046 1050
rect 9100 1022 9130 1050
rect 9184 1022 9214 1050
rect 9268 1022 9298 1050
rect 9484 1104 9514 1142
rect 9568 1104 9598 1142
rect 9652 1104 9682 1142
rect 9736 1104 9766 1142
rect 9820 1104 9850 1142
rect 9904 1104 9934 1142
rect 9484 1094 9934 1104
rect 9484 1060 9508 1094
rect 9542 1060 9576 1094
rect 9610 1060 9644 1094
rect 9678 1060 9712 1094
rect 9746 1060 9780 1094
rect 9814 1060 9848 1094
rect 9882 1060 9934 1094
rect 9484 1050 9934 1060
rect 9484 1022 9514 1050
rect 9568 1022 9598 1050
rect 9652 1022 9682 1050
rect 9736 1022 9766 1050
rect 9820 1022 9850 1050
rect 9904 1022 9934 1050
rect 9988 1104 10018 1142
rect 10072 1104 10102 1142
rect 10156 1104 10186 1142
rect 10240 1104 10270 1142
rect 10324 1104 10354 1142
rect 10408 1104 10438 1142
rect 10492 1104 10522 1142
rect 10576 1104 10606 1142
rect 10660 1104 10690 1142
rect 10744 1104 10774 1142
rect 10828 1104 10858 1142
rect 10912 1104 10942 1142
rect 10996 1104 11026 1142
rect 11080 1104 11110 1142
rect 11164 1104 11194 1142
rect 11248 1104 11278 1142
rect 13034 1110 13064 1145
rect 13128 1123 13158 1184
rect 9988 1094 11282 1104
rect 9988 1060 10008 1094
rect 10042 1060 10076 1094
rect 10110 1060 10144 1094
rect 10178 1060 10212 1094
rect 10246 1060 10280 1094
rect 10314 1060 10348 1094
rect 10382 1060 10416 1094
rect 10450 1060 10484 1094
rect 10518 1060 10552 1094
rect 10586 1060 10620 1094
rect 10654 1060 10688 1094
rect 10722 1060 10756 1094
rect 10790 1060 10824 1094
rect 10858 1060 10892 1094
rect 10926 1060 10960 1094
rect 10994 1060 11028 1094
rect 11062 1060 11096 1094
rect 11130 1060 11164 1094
rect 11198 1060 11232 1094
rect 11266 1060 11282 1094
rect 9988 1050 11282 1060
rect 12988 1094 13064 1110
rect 12988 1060 12998 1094
rect 13032 1060 13064 1094
rect 9988 1022 10018 1050
rect 10072 1022 10102 1050
rect 10156 1022 10186 1050
rect 10240 1022 10270 1050
rect 10324 1022 10354 1050
rect 10408 1022 10438 1050
rect 10492 1022 10522 1050
rect 10576 1022 10606 1050
rect 10660 1022 10690 1050
rect 10744 1022 10774 1050
rect 10828 1022 10858 1050
rect 10912 1022 10942 1050
rect 10996 1022 11026 1050
rect 11080 1022 11110 1050
rect 11164 1022 11194 1050
rect 11248 1022 11278 1050
rect 12988 1044 13064 1060
rect 13106 1107 13160 1123
rect 13106 1073 13116 1107
rect 13150 1073 13160 1107
rect 13316 1106 13346 1142
rect 13106 1057 13160 1073
rect 13265 1094 13346 1106
rect 13400 1104 13430 1142
rect 13484 1104 13514 1142
rect 13568 1104 13598 1142
rect 13652 1104 13682 1142
rect 13265 1060 13281 1094
rect 13315 1060 13346 1094
rect 13034 1035 13064 1044
rect 13034 1011 13070 1035
rect 13040 996 13070 1011
rect 13128 996 13158 1057
rect 13265 1048 13346 1060
rect 13399 1094 13682 1104
rect 13399 1060 13415 1094
rect 13449 1060 13682 1094
rect 13399 1050 13682 1060
rect 13316 1022 13346 1048
rect 13400 1022 13430 1050
rect 13484 1022 13514 1050
rect 13568 1022 13598 1050
rect 13652 1022 13682 1050
rect 13868 1104 13898 1142
rect 13952 1104 13982 1142
rect 14036 1104 14066 1142
rect 14120 1104 14150 1142
rect 14204 1104 14234 1142
rect 14288 1104 14318 1142
rect 13868 1094 14318 1104
rect 13868 1060 13892 1094
rect 13926 1060 13960 1094
rect 13994 1060 14028 1094
rect 14062 1060 14096 1094
rect 14130 1060 14164 1094
rect 14198 1060 14232 1094
rect 14266 1060 14318 1094
rect 13868 1050 14318 1060
rect 13868 1022 13898 1050
rect 13952 1022 13982 1050
rect 14036 1022 14066 1050
rect 14120 1022 14150 1050
rect 14204 1022 14234 1050
rect 14288 1022 14318 1050
rect 14372 1104 14402 1142
rect 14456 1104 14486 1142
rect 14540 1104 14570 1142
rect 14624 1104 14654 1142
rect 14708 1104 14738 1142
rect 14792 1104 14822 1142
rect 14876 1104 14906 1142
rect 14960 1104 14990 1142
rect 15044 1104 15074 1142
rect 15128 1104 15158 1142
rect 15212 1104 15242 1142
rect 15296 1104 15326 1142
rect 15380 1104 15410 1142
rect 15464 1104 15494 1142
rect 15548 1104 15578 1142
rect 15632 1104 15662 1142
rect 14372 1094 15666 1104
rect 14372 1060 14392 1094
rect 14426 1060 14460 1094
rect 14494 1060 14528 1094
rect 14562 1060 14596 1094
rect 14630 1060 14664 1094
rect 14698 1060 14732 1094
rect 14766 1060 14800 1094
rect 14834 1060 14868 1094
rect 14902 1060 14936 1094
rect 14970 1060 15004 1094
rect 15038 1060 15072 1094
rect 15106 1060 15140 1094
rect 15174 1060 15208 1094
rect 15242 1060 15276 1094
rect 15310 1060 15344 1094
rect 15378 1060 15412 1094
rect 15446 1060 15480 1094
rect 15514 1060 15548 1094
rect 15582 1060 15616 1094
rect 15650 1060 15666 1094
rect 14372 1050 15666 1060
rect 14372 1022 14402 1050
rect 14456 1022 14486 1050
rect 14540 1022 14570 1050
rect 14624 1022 14654 1050
rect 14708 1022 14738 1050
rect 14792 1022 14822 1050
rect 14876 1022 14906 1050
rect 14960 1022 14990 1050
rect 15044 1022 15074 1050
rect 15128 1022 15158 1050
rect 15212 1022 15242 1050
rect 15296 1022 15326 1050
rect 15380 1022 15410 1050
rect 15464 1022 15494 1050
rect 15548 1022 15578 1050
rect 15632 1022 15662 1050
rect 8656 866 8686 892
rect 8744 866 8774 892
rect 8932 866 8962 892
rect 9016 866 9046 892
rect 9100 866 9130 892
rect 9184 866 9214 892
rect 9268 866 9298 892
rect 9484 866 9514 892
rect 9568 866 9598 892
rect 9652 866 9682 892
rect 9736 866 9766 892
rect 9820 866 9850 892
rect 9904 866 9934 892
rect 9988 866 10018 892
rect 10072 866 10102 892
rect 10156 866 10186 892
rect 10240 866 10270 892
rect 10324 866 10354 892
rect 10408 866 10438 892
rect 10492 866 10522 892
rect 10576 866 10606 892
rect 10660 866 10690 892
rect 10744 866 10774 892
rect 10828 866 10858 892
rect 10912 866 10942 892
rect 10996 866 11026 892
rect 11080 866 11110 892
rect 11164 866 11194 892
rect 11248 866 11278 892
rect 13040 866 13070 892
rect 13128 866 13158 892
rect 13316 866 13346 892
rect 13400 866 13430 892
rect 13484 866 13514 892
rect 13568 866 13598 892
rect 13652 866 13682 892
rect 13868 866 13898 892
rect 13952 866 13982 892
rect 14036 866 14066 892
rect 14120 866 14150 892
rect 14204 866 14234 892
rect 14288 866 14318 892
rect 14372 866 14402 892
rect 14456 866 14486 892
rect 14540 866 14570 892
rect 14624 866 14654 892
rect 14708 866 14738 892
rect 14792 866 14822 892
rect 14876 866 14906 892
rect 14960 866 14990 892
rect 15044 866 15074 892
rect 15128 866 15158 892
rect 15212 866 15242 892
rect 15296 866 15326 892
rect 15380 866 15410 892
rect 15464 866 15494 892
rect 15548 866 15578 892
rect 15632 866 15662 892
rect 8654 200 8684 226
rect 10728 200 10758 226
rect 11046 200 11076 226
rect 13120 200 13150 226
rect 13438 200 13468 226
rect 15510 200 15540 226
rect 15830 200 15860 226
rect 17904 200 17934 226
rect 18222 200 18252 226
rect 20296 200 20326 226
rect 20614 200 20644 226
rect 22686 200 22716 226
rect 23006 200 23036 226
rect 25080 200 25110 226
rect 8763 161 8793 187
rect 8866 161 8896 187
rect 9080 161 9110 187
rect 9152 161 9182 187
rect 9248 161 9278 187
rect 10134 161 10164 187
rect 10230 161 10260 187
rect 10302 161 10332 187
rect 10516 161 10546 187
rect 10619 161 10649 187
rect 8654 -32 8684 0
rect 8763 -32 8793 77
rect 8866 62 8896 77
rect 8866 32 9014 62
rect 9080 45 9110 77
rect 8651 -48 8705 -32
rect 8651 -82 8661 -48
rect 8695 -82 8705 -48
rect 8651 -98 8705 -82
rect 8747 -48 8801 -32
rect 8747 -82 8757 -48
rect 8791 -82 8801 -48
rect 8984 -68 9014 32
rect 9056 29 9110 45
rect 9056 -5 9066 29
rect 9100 -5 9110 29
rect 9056 -21 9110 -5
rect 8747 -98 8801 -82
rect 8859 -84 8942 -68
rect 8654 -120 8684 -98
rect 8763 -166 8793 -98
rect 8859 -118 8898 -84
rect 8932 -118 8942 -84
rect 8859 -134 8942 -118
rect 8984 -84 9038 -68
rect 9152 -74 9182 77
rect 9248 45 9278 77
rect 9224 29 9278 45
rect 9224 -5 9234 29
rect 9268 -5 9278 29
rect 9224 -21 9278 -5
rect 8984 -118 8994 -84
rect 9028 -118 9038 -84
rect 9140 -84 9206 -74
rect 9140 -98 9156 -84
rect 8984 -134 9038 -118
rect 9080 -118 9156 -98
rect 9190 -118 9206 -84
rect 9080 -128 9206 -118
rect 8859 -166 8889 -134
rect 8984 -166 9014 -134
rect 9080 -166 9110 -128
rect 9248 -166 9278 -21
rect 10134 45 10164 77
rect 10134 29 10188 45
rect 10134 -5 10144 29
rect 10178 -5 10188 29
rect 10134 -21 10188 -5
rect 10134 -166 10164 -21
rect 10230 -74 10260 77
rect 10302 45 10332 77
rect 10516 62 10546 77
rect 10302 29 10356 45
rect 10302 -5 10312 29
rect 10346 -5 10356 29
rect 10302 -21 10356 -5
rect 10398 32 10546 62
rect 10398 -68 10428 32
rect 10619 -32 10649 77
rect 11155 161 11185 187
rect 11258 161 11288 187
rect 11472 161 11502 187
rect 11544 161 11574 187
rect 11640 161 11670 187
rect 12526 161 12556 187
rect 12622 161 12652 187
rect 12694 161 12724 187
rect 12908 161 12938 187
rect 13011 161 13041 187
rect 10728 -32 10758 0
rect 11046 -32 11076 0
rect 11155 -32 11185 77
rect 11258 62 11288 77
rect 11258 32 11406 62
rect 11472 45 11502 77
rect 10611 -48 10665 -32
rect 10206 -84 10272 -74
rect 10206 -118 10222 -84
rect 10256 -98 10272 -84
rect 10374 -84 10428 -68
rect 10256 -118 10332 -98
rect 10206 -128 10332 -118
rect 10302 -166 10332 -128
rect 10374 -118 10384 -84
rect 10418 -118 10428 -84
rect 10374 -134 10428 -118
rect 10470 -84 10553 -68
rect 10470 -118 10480 -84
rect 10514 -118 10553 -84
rect 10611 -82 10621 -48
rect 10655 -82 10665 -48
rect 10611 -98 10665 -82
rect 10707 -48 10761 -32
rect 10707 -82 10717 -48
rect 10751 -82 10761 -48
rect 10707 -98 10761 -82
rect 11043 -48 11097 -32
rect 11043 -82 11053 -48
rect 11087 -82 11097 -48
rect 11043 -98 11097 -82
rect 11139 -48 11193 -32
rect 11139 -82 11149 -48
rect 11183 -82 11193 -48
rect 11376 -68 11406 32
rect 11448 29 11502 45
rect 11448 -5 11458 29
rect 11492 -5 11502 29
rect 11448 -21 11502 -5
rect 11139 -98 11193 -82
rect 11251 -84 11334 -68
rect 10470 -134 10553 -118
rect 10398 -166 10428 -134
rect 10523 -166 10553 -134
rect 10619 -166 10649 -98
rect 10728 -120 10758 -98
rect 11046 -120 11076 -98
rect 11155 -166 11185 -98
rect 11251 -118 11290 -84
rect 11324 -118 11334 -84
rect 11251 -134 11334 -118
rect 11376 -84 11430 -68
rect 11544 -74 11574 77
rect 11640 45 11670 77
rect 11616 29 11670 45
rect 11616 -5 11626 29
rect 11660 -5 11670 29
rect 11616 -21 11670 -5
rect 11376 -118 11386 -84
rect 11420 -118 11430 -84
rect 11532 -84 11598 -74
rect 11532 -98 11548 -84
rect 11376 -134 11430 -118
rect 11472 -118 11548 -98
rect 11582 -118 11598 -84
rect 11472 -128 11598 -118
rect 11251 -166 11281 -134
rect 11376 -166 11406 -134
rect 11472 -166 11502 -128
rect 11640 -166 11670 -21
rect 12526 45 12556 77
rect 12526 29 12580 45
rect 12526 -5 12536 29
rect 12570 -5 12580 29
rect 12526 -21 12580 -5
rect 12526 -166 12556 -21
rect 12622 -74 12652 77
rect 12694 45 12724 77
rect 12908 62 12938 77
rect 12694 29 12748 45
rect 12694 -5 12704 29
rect 12738 -5 12748 29
rect 12694 -21 12748 -5
rect 12790 32 12938 62
rect 12790 -68 12820 32
rect 13011 -32 13041 77
rect 13547 161 13577 187
rect 13650 161 13680 187
rect 13864 161 13894 187
rect 13936 161 13966 187
rect 14032 161 14062 187
rect 14916 161 14946 187
rect 15012 161 15042 187
rect 15084 161 15114 187
rect 15298 161 15328 187
rect 15401 161 15431 187
rect 13120 -32 13150 0
rect 13438 -32 13468 0
rect 13547 -32 13577 77
rect 13650 62 13680 77
rect 13650 32 13798 62
rect 13864 45 13894 77
rect 13003 -48 13057 -32
rect 12598 -84 12664 -74
rect 12598 -118 12614 -84
rect 12648 -98 12664 -84
rect 12766 -84 12820 -68
rect 12648 -118 12724 -98
rect 12598 -128 12724 -118
rect 12694 -166 12724 -128
rect 12766 -118 12776 -84
rect 12810 -118 12820 -84
rect 12766 -134 12820 -118
rect 12862 -84 12945 -68
rect 12862 -118 12872 -84
rect 12906 -118 12945 -84
rect 13003 -82 13013 -48
rect 13047 -82 13057 -48
rect 13003 -98 13057 -82
rect 13099 -48 13153 -32
rect 13099 -82 13109 -48
rect 13143 -82 13153 -48
rect 13099 -98 13153 -82
rect 13435 -48 13489 -32
rect 13435 -82 13445 -48
rect 13479 -82 13489 -48
rect 13435 -98 13489 -82
rect 13531 -48 13585 -32
rect 13531 -82 13541 -48
rect 13575 -82 13585 -48
rect 13768 -68 13798 32
rect 13840 29 13894 45
rect 13840 -5 13850 29
rect 13884 -5 13894 29
rect 13840 -21 13894 -5
rect 13531 -98 13585 -82
rect 13643 -84 13726 -68
rect 12862 -134 12945 -118
rect 12790 -166 12820 -134
rect 12915 -166 12945 -134
rect 13011 -166 13041 -98
rect 13120 -120 13150 -98
rect 13438 -120 13468 -98
rect 13547 -166 13577 -98
rect 13643 -118 13682 -84
rect 13716 -118 13726 -84
rect 13643 -134 13726 -118
rect 13768 -84 13822 -68
rect 13936 -74 13966 77
rect 14032 45 14062 77
rect 14008 29 14062 45
rect 14008 -5 14018 29
rect 14052 -5 14062 29
rect 14008 -21 14062 -5
rect 13768 -118 13778 -84
rect 13812 -118 13822 -84
rect 13924 -84 13990 -74
rect 13924 -98 13940 -84
rect 13768 -134 13822 -118
rect 13864 -118 13940 -98
rect 13974 -118 13990 -84
rect 13864 -128 13990 -118
rect 13643 -166 13673 -134
rect 13768 -166 13798 -134
rect 13864 -166 13894 -128
rect 14032 -166 14062 -21
rect 14916 45 14946 77
rect 14916 29 14970 45
rect 14916 -5 14926 29
rect 14960 -5 14970 29
rect 14916 -21 14970 -5
rect 14916 -166 14946 -21
rect 15012 -74 15042 77
rect 15084 45 15114 77
rect 15298 62 15328 77
rect 15084 29 15138 45
rect 15084 -5 15094 29
rect 15128 -5 15138 29
rect 15084 -21 15138 -5
rect 15180 32 15328 62
rect 15180 -68 15210 32
rect 15401 -32 15431 77
rect 15939 161 15969 187
rect 16042 161 16072 187
rect 16256 161 16286 187
rect 16328 161 16358 187
rect 16424 161 16454 187
rect 17310 161 17340 187
rect 17406 161 17436 187
rect 17478 161 17508 187
rect 17692 161 17722 187
rect 17795 161 17825 187
rect 15510 -32 15540 0
rect 15830 -32 15860 0
rect 15939 -32 15969 77
rect 16042 62 16072 77
rect 16042 32 16190 62
rect 16256 45 16286 77
rect 15393 -48 15447 -32
rect 14988 -84 15054 -74
rect 14988 -118 15004 -84
rect 15038 -98 15054 -84
rect 15156 -84 15210 -68
rect 15038 -118 15114 -98
rect 14988 -128 15114 -118
rect 15084 -166 15114 -128
rect 15156 -118 15166 -84
rect 15200 -118 15210 -84
rect 15156 -134 15210 -118
rect 15252 -84 15335 -68
rect 15252 -118 15262 -84
rect 15296 -118 15335 -84
rect 15393 -82 15403 -48
rect 15437 -82 15447 -48
rect 15393 -98 15447 -82
rect 15489 -48 15543 -32
rect 15489 -82 15499 -48
rect 15533 -82 15543 -48
rect 15489 -98 15543 -82
rect 15827 -48 15881 -32
rect 15827 -82 15837 -48
rect 15871 -82 15881 -48
rect 15827 -98 15881 -82
rect 15923 -48 15977 -32
rect 15923 -82 15933 -48
rect 15967 -82 15977 -48
rect 16160 -68 16190 32
rect 16232 29 16286 45
rect 16232 -5 16242 29
rect 16276 -5 16286 29
rect 16232 -21 16286 -5
rect 15923 -98 15977 -82
rect 16035 -84 16118 -68
rect 15252 -134 15335 -118
rect 15180 -166 15210 -134
rect 15305 -166 15335 -134
rect 15401 -166 15431 -98
rect 15510 -120 15540 -98
rect 15830 -120 15860 -98
rect 15939 -166 15969 -98
rect 16035 -118 16074 -84
rect 16108 -118 16118 -84
rect 16035 -134 16118 -118
rect 16160 -84 16214 -68
rect 16328 -74 16358 77
rect 16424 45 16454 77
rect 16400 29 16454 45
rect 16400 -5 16410 29
rect 16444 -5 16454 29
rect 16400 -21 16454 -5
rect 16160 -118 16170 -84
rect 16204 -118 16214 -84
rect 16316 -84 16382 -74
rect 16316 -98 16332 -84
rect 16160 -134 16214 -118
rect 16256 -118 16332 -98
rect 16366 -118 16382 -84
rect 16256 -128 16382 -118
rect 16035 -166 16065 -134
rect 16160 -166 16190 -134
rect 16256 -166 16286 -128
rect 16424 -166 16454 -21
rect 17310 45 17340 77
rect 17310 29 17364 45
rect 17310 -5 17320 29
rect 17354 -5 17364 29
rect 17310 -21 17364 -5
rect 17310 -166 17340 -21
rect 17406 -74 17436 77
rect 17478 45 17508 77
rect 17692 62 17722 77
rect 17478 29 17532 45
rect 17478 -5 17488 29
rect 17522 -5 17532 29
rect 17478 -21 17532 -5
rect 17574 32 17722 62
rect 17574 -68 17604 32
rect 17795 -32 17825 77
rect 18331 161 18361 187
rect 18434 161 18464 187
rect 18648 161 18678 187
rect 18720 161 18750 187
rect 18816 161 18846 187
rect 19702 161 19732 187
rect 19798 161 19828 187
rect 19870 161 19900 187
rect 20084 161 20114 187
rect 20187 161 20217 187
rect 17904 -32 17934 0
rect 18222 -32 18252 0
rect 18331 -32 18361 77
rect 18434 62 18464 77
rect 18434 32 18582 62
rect 18648 45 18678 77
rect 17787 -48 17841 -32
rect 17382 -84 17448 -74
rect 17382 -118 17398 -84
rect 17432 -98 17448 -84
rect 17550 -84 17604 -68
rect 17432 -118 17508 -98
rect 17382 -128 17508 -118
rect 17478 -166 17508 -128
rect 17550 -118 17560 -84
rect 17594 -118 17604 -84
rect 17550 -134 17604 -118
rect 17646 -84 17729 -68
rect 17646 -118 17656 -84
rect 17690 -118 17729 -84
rect 17787 -82 17797 -48
rect 17831 -82 17841 -48
rect 17787 -98 17841 -82
rect 17883 -48 17937 -32
rect 17883 -82 17893 -48
rect 17927 -82 17937 -48
rect 17883 -98 17937 -82
rect 18219 -48 18273 -32
rect 18219 -82 18229 -48
rect 18263 -82 18273 -48
rect 18219 -98 18273 -82
rect 18315 -48 18369 -32
rect 18315 -82 18325 -48
rect 18359 -82 18369 -48
rect 18552 -68 18582 32
rect 18624 29 18678 45
rect 18624 -5 18634 29
rect 18668 -5 18678 29
rect 18624 -21 18678 -5
rect 18315 -98 18369 -82
rect 18427 -84 18510 -68
rect 17646 -134 17729 -118
rect 17574 -166 17604 -134
rect 17699 -166 17729 -134
rect 17795 -166 17825 -98
rect 17904 -120 17934 -98
rect 18222 -120 18252 -98
rect 18331 -166 18361 -98
rect 18427 -118 18466 -84
rect 18500 -118 18510 -84
rect 18427 -134 18510 -118
rect 18552 -84 18606 -68
rect 18720 -74 18750 77
rect 18816 45 18846 77
rect 18792 29 18846 45
rect 18792 -5 18802 29
rect 18836 -5 18846 29
rect 18792 -21 18846 -5
rect 18552 -118 18562 -84
rect 18596 -118 18606 -84
rect 18708 -84 18774 -74
rect 18708 -98 18724 -84
rect 18552 -134 18606 -118
rect 18648 -118 18724 -98
rect 18758 -118 18774 -84
rect 18648 -128 18774 -118
rect 18427 -166 18457 -134
rect 18552 -166 18582 -134
rect 18648 -166 18678 -128
rect 18816 -166 18846 -21
rect 19702 45 19732 77
rect 19702 29 19756 45
rect 19702 -5 19712 29
rect 19746 -5 19756 29
rect 19702 -21 19756 -5
rect 19702 -166 19732 -21
rect 19798 -74 19828 77
rect 19870 45 19900 77
rect 20084 62 20114 77
rect 19870 29 19924 45
rect 19870 -5 19880 29
rect 19914 -5 19924 29
rect 19870 -21 19924 -5
rect 19966 32 20114 62
rect 19966 -68 19996 32
rect 20187 -32 20217 77
rect 20723 161 20753 187
rect 20826 161 20856 187
rect 21040 161 21070 187
rect 21112 161 21142 187
rect 21208 161 21238 187
rect 22092 161 22122 187
rect 22188 161 22218 187
rect 22260 161 22290 187
rect 22474 161 22504 187
rect 22577 161 22607 187
rect 20296 -32 20326 0
rect 20614 -32 20644 0
rect 20723 -32 20753 77
rect 20826 62 20856 77
rect 20826 32 20974 62
rect 21040 45 21070 77
rect 20179 -48 20233 -32
rect 19774 -84 19840 -74
rect 19774 -118 19790 -84
rect 19824 -98 19840 -84
rect 19942 -84 19996 -68
rect 19824 -118 19900 -98
rect 19774 -128 19900 -118
rect 19870 -166 19900 -128
rect 19942 -118 19952 -84
rect 19986 -118 19996 -84
rect 19942 -134 19996 -118
rect 20038 -84 20121 -68
rect 20038 -118 20048 -84
rect 20082 -118 20121 -84
rect 20179 -82 20189 -48
rect 20223 -82 20233 -48
rect 20179 -98 20233 -82
rect 20275 -48 20329 -32
rect 20275 -82 20285 -48
rect 20319 -82 20329 -48
rect 20275 -98 20329 -82
rect 20611 -48 20665 -32
rect 20611 -82 20621 -48
rect 20655 -82 20665 -48
rect 20611 -98 20665 -82
rect 20707 -48 20761 -32
rect 20707 -82 20717 -48
rect 20751 -82 20761 -48
rect 20944 -68 20974 32
rect 21016 29 21070 45
rect 21016 -5 21026 29
rect 21060 -5 21070 29
rect 21016 -21 21070 -5
rect 20707 -98 20761 -82
rect 20819 -84 20902 -68
rect 20038 -134 20121 -118
rect 19966 -166 19996 -134
rect 20091 -166 20121 -134
rect 20187 -166 20217 -98
rect 20296 -120 20326 -98
rect 20614 -120 20644 -98
rect 20723 -166 20753 -98
rect 20819 -118 20858 -84
rect 20892 -118 20902 -84
rect 20819 -134 20902 -118
rect 20944 -84 20998 -68
rect 21112 -74 21142 77
rect 21208 45 21238 77
rect 21184 29 21238 45
rect 21184 -5 21194 29
rect 21228 -5 21238 29
rect 21184 -21 21238 -5
rect 20944 -118 20954 -84
rect 20988 -118 20998 -84
rect 21100 -84 21166 -74
rect 21100 -98 21116 -84
rect 20944 -134 20998 -118
rect 21040 -118 21116 -98
rect 21150 -118 21166 -84
rect 21040 -128 21166 -118
rect 20819 -166 20849 -134
rect 20944 -166 20974 -134
rect 21040 -166 21070 -128
rect 21208 -166 21238 -21
rect 22092 45 22122 77
rect 22092 29 22146 45
rect 22092 -5 22102 29
rect 22136 -5 22146 29
rect 22092 -21 22146 -5
rect 22092 -166 22122 -21
rect 22188 -74 22218 77
rect 22260 45 22290 77
rect 22474 62 22504 77
rect 22260 29 22314 45
rect 22260 -5 22270 29
rect 22304 -5 22314 29
rect 22260 -21 22314 -5
rect 22356 32 22504 62
rect 22356 -68 22386 32
rect 22577 -32 22607 77
rect 23115 161 23145 187
rect 23218 161 23248 187
rect 23432 161 23462 187
rect 23504 161 23534 187
rect 23600 161 23630 187
rect 24486 161 24516 187
rect 24582 161 24612 187
rect 24654 161 24684 187
rect 24868 161 24898 187
rect 24971 161 25001 187
rect 22686 -32 22716 0
rect 23006 -32 23036 0
rect 23115 -32 23145 77
rect 23218 62 23248 77
rect 23218 32 23366 62
rect 23432 45 23462 77
rect 22569 -48 22623 -32
rect 22164 -84 22230 -74
rect 22164 -118 22180 -84
rect 22214 -98 22230 -84
rect 22332 -84 22386 -68
rect 22214 -118 22290 -98
rect 22164 -128 22290 -118
rect 22260 -166 22290 -128
rect 22332 -118 22342 -84
rect 22376 -118 22386 -84
rect 22332 -134 22386 -118
rect 22428 -84 22511 -68
rect 22428 -118 22438 -84
rect 22472 -118 22511 -84
rect 22569 -82 22579 -48
rect 22613 -82 22623 -48
rect 22569 -98 22623 -82
rect 22665 -48 22719 -32
rect 22665 -82 22675 -48
rect 22709 -82 22719 -48
rect 22665 -98 22719 -82
rect 23003 -48 23057 -32
rect 23003 -82 23013 -48
rect 23047 -82 23057 -48
rect 23003 -98 23057 -82
rect 23099 -48 23153 -32
rect 23099 -82 23109 -48
rect 23143 -82 23153 -48
rect 23336 -68 23366 32
rect 23408 29 23462 45
rect 23408 -5 23418 29
rect 23452 -5 23462 29
rect 23408 -21 23462 -5
rect 23099 -98 23153 -82
rect 23211 -84 23294 -68
rect 22428 -134 22511 -118
rect 22356 -166 22386 -134
rect 22481 -166 22511 -134
rect 22577 -166 22607 -98
rect 22686 -120 22716 -98
rect 23006 -120 23036 -98
rect 23115 -166 23145 -98
rect 23211 -118 23250 -84
rect 23284 -118 23294 -84
rect 23211 -134 23294 -118
rect 23336 -84 23390 -68
rect 23504 -74 23534 77
rect 23600 45 23630 77
rect 23576 29 23630 45
rect 23576 -5 23586 29
rect 23620 -5 23630 29
rect 23576 -21 23630 -5
rect 23336 -118 23346 -84
rect 23380 -118 23390 -84
rect 23492 -84 23558 -74
rect 23492 -98 23508 -84
rect 23336 -134 23390 -118
rect 23432 -118 23508 -98
rect 23542 -118 23558 -84
rect 23432 -128 23558 -118
rect 23211 -166 23241 -134
rect 23336 -166 23366 -134
rect 23432 -166 23462 -128
rect 23600 -166 23630 -21
rect 24486 45 24516 77
rect 24486 29 24540 45
rect 24486 -5 24496 29
rect 24530 -5 24540 29
rect 24486 -21 24540 -5
rect 24486 -166 24516 -21
rect 24582 -74 24612 77
rect 24654 45 24684 77
rect 24868 62 24898 77
rect 24654 29 24708 45
rect 24654 -5 24664 29
rect 24698 -5 24708 29
rect 24654 -21 24708 -5
rect 24750 32 24898 62
rect 24750 -68 24780 32
rect 24971 -32 25001 77
rect 25080 -32 25110 0
rect 24963 -48 25017 -32
rect 24558 -84 24624 -74
rect 24558 -118 24574 -84
rect 24608 -98 24624 -84
rect 24726 -84 24780 -68
rect 24608 -118 24684 -98
rect 24558 -128 24684 -118
rect 24654 -166 24684 -128
rect 24726 -118 24736 -84
rect 24770 -118 24780 -84
rect 24726 -134 24780 -118
rect 24822 -84 24905 -68
rect 24822 -118 24832 -84
rect 24866 -118 24905 -84
rect 24963 -82 24973 -48
rect 25007 -82 25017 -48
rect 24963 -98 25017 -82
rect 25059 -48 25113 -32
rect 25059 -82 25069 -48
rect 25103 -82 25113 -48
rect 25059 -98 25113 -82
rect 24822 -134 24905 -118
rect 24750 -166 24780 -134
rect 24875 -166 24905 -134
rect 24971 -166 25001 -98
rect 25080 -120 25110 -98
rect 8654 -276 8684 -250
rect 8763 -276 8793 -250
rect 8859 -276 8889 -250
rect 8984 -276 9014 -250
rect 9080 -276 9110 -250
rect 9248 -276 9278 -250
rect 10134 -276 10164 -250
rect 10302 -276 10332 -250
rect 10398 -276 10428 -250
rect 10523 -276 10553 -250
rect 10619 -276 10649 -250
rect 10728 -276 10758 -250
rect 11046 -276 11076 -250
rect 11155 -276 11185 -250
rect 11251 -276 11281 -250
rect 11376 -276 11406 -250
rect 11472 -276 11502 -250
rect 11640 -276 11670 -250
rect 12526 -276 12556 -250
rect 12694 -276 12724 -250
rect 12790 -276 12820 -250
rect 12915 -276 12945 -250
rect 13011 -276 13041 -250
rect 13120 -276 13150 -250
rect 13438 -276 13468 -250
rect 13547 -276 13577 -250
rect 13643 -276 13673 -250
rect 13768 -276 13798 -250
rect 13864 -276 13894 -250
rect 14032 -276 14062 -250
rect 14916 -276 14946 -250
rect 15084 -276 15114 -250
rect 15180 -276 15210 -250
rect 15305 -276 15335 -250
rect 15401 -276 15431 -250
rect 15510 -276 15540 -250
rect 15830 -276 15860 -250
rect 15939 -276 15969 -250
rect 16035 -276 16065 -250
rect 16160 -276 16190 -250
rect 16256 -276 16286 -250
rect 16424 -276 16454 -250
rect 17310 -276 17340 -250
rect 17478 -276 17508 -250
rect 17574 -276 17604 -250
rect 17699 -276 17729 -250
rect 17795 -276 17825 -250
rect 17904 -276 17934 -250
rect 18222 -276 18252 -250
rect 18331 -276 18361 -250
rect 18427 -276 18457 -250
rect 18552 -276 18582 -250
rect 18648 -276 18678 -250
rect 18816 -276 18846 -250
rect 19702 -276 19732 -250
rect 19870 -276 19900 -250
rect 19966 -276 19996 -250
rect 20091 -276 20121 -250
rect 20187 -276 20217 -250
rect 20296 -276 20326 -250
rect 20614 -276 20644 -250
rect 20723 -276 20753 -250
rect 20819 -276 20849 -250
rect 20944 -276 20974 -250
rect 21040 -276 21070 -250
rect 21208 -276 21238 -250
rect 22092 -276 22122 -250
rect 22260 -276 22290 -250
rect 22356 -276 22386 -250
rect 22481 -276 22511 -250
rect 22577 -276 22607 -250
rect 22686 -276 22716 -250
rect 23006 -276 23036 -250
rect 23115 -276 23145 -250
rect 23211 -276 23241 -250
rect 23336 -276 23366 -250
rect 23432 -276 23462 -250
rect 23600 -276 23630 -250
rect 24486 -276 24516 -250
rect 24654 -276 24684 -250
rect 24750 -276 24780 -250
rect 24875 -276 24905 -250
rect 24971 -276 25001 -250
rect 25080 -276 25110 -250
rect 10460 -407 10526 -391
rect 10460 -441 10476 -407
rect 10510 -441 10526 -407
rect 12852 -408 12918 -392
rect 10460 -457 10526 -441
rect 12852 -442 12868 -408
rect 12902 -442 12918 -408
rect 15244 -408 15310 -392
rect 8654 -494 8684 -468
rect 8738 -494 8768 -468
rect 8926 -488 8956 -462
rect 9018 -488 9048 -462
rect 9102 -488 9132 -462
rect 9222 -488 9252 -462
rect 9328 -488 9358 -462
rect 9436 -488 9466 -462
rect 9520 -488 9550 -462
rect 9657 -488 9687 -462
rect 9801 -488 9831 -462
rect 9885 -488 9915 -462
rect 9990 -488 10020 -462
rect 10111 -488 10141 -462
rect 10217 -488 10247 -462
rect 10289 -488 10319 -462
rect 8654 -637 8684 -622
rect 8620 -667 8684 -637
rect 8620 -705 8650 -667
rect 8596 -721 8650 -705
rect 8738 -711 8768 -622
rect 8596 -755 8606 -721
rect 8640 -755 8650 -721
rect 8596 -771 8650 -755
rect 8692 -721 8768 -711
rect 8926 -718 8956 -572
rect 9018 -706 9048 -572
rect 9102 -610 9132 -572
rect 9222 -604 9252 -572
rect 9090 -620 9156 -610
rect 9090 -654 9106 -620
rect 9140 -654 9156 -620
rect 9090 -664 9156 -654
rect 9222 -620 9286 -604
rect 9222 -654 9242 -620
rect 9276 -654 9286 -620
rect 9222 -670 9286 -654
rect 8692 -755 8708 -721
rect 8742 -755 8768 -721
rect 8692 -765 8768 -755
rect 8620 -809 8650 -771
rect 8620 -839 8684 -809
rect 8654 -854 8684 -839
rect 8738 -854 8768 -765
rect 8914 -734 8968 -718
rect 8914 -768 8924 -734
rect 8958 -768 8968 -734
rect 9018 -736 9156 -706
rect 8914 -784 8968 -768
rect 9126 -766 9156 -736
rect 8926 -854 8956 -784
rect 9021 -794 9084 -778
rect 9021 -828 9040 -794
rect 9074 -828 9084 -794
rect 9021 -844 9084 -828
rect 9126 -782 9180 -766
rect 9126 -816 9136 -782
rect 9170 -816 9180 -782
rect 9126 -832 9180 -816
rect 9021 -866 9051 -844
rect 9126 -866 9156 -832
rect 9222 -854 9252 -670
rect 9328 -756 9358 -572
rect 9801 -604 9831 -572
rect 9777 -620 9831 -604
rect 9885 -610 9915 -572
rect 9990 -604 10020 -572
rect 9777 -654 9787 -620
rect 9821 -654 9831 -620
rect 9436 -688 9466 -656
rect 9520 -688 9550 -656
rect 9400 -704 9466 -688
rect 9400 -738 9410 -704
rect 9444 -738 9466 -704
rect 9400 -754 9466 -738
rect 9516 -704 9606 -688
rect 9516 -738 9562 -704
rect 9596 -738 9606 -704
rect 9516 -754 9606 -738
rect 9657 -722 9687 -656
rect 9777 -670 9831 -654
rect 9873 -620 9939 -610
rect 9873 -654 9889 -620
rect 9923 -654 9939 -620
rect 9873 -664 9939 -654
rect 9990 -620 10069 -604
rect 9990 -654 10025 -620
rect 10059 -654 10069 -620
rect 9990 -670 10069 -654
rect 9801 -706 9831 -670
rect 9657 -738 9734 -722
rect 9801 -736 9938 -706
rect 9657 -752 9690 -738
rect 9298 -772 9358 -756
rect 9298 -806 9308 -772
rect 9342 -792 9358 -772
rect 9342 -806 9366 -792
rect 9298 -822 9366 -806
rect 9432 -810 9462 -754
rect 9516 -810 9546 -754
rect 9680 -772 9690 -752
rect 9724 -772 9734 -738
rect 9680 -788 9734 -772
rect 9704 -810 9734 -788
rect 9812 -794 9866 -778
rect 9336 -854 9366 -822
rect 9812 -828 9822 -794
rect 9856 -828 9866 -794
rect 9812 -844 9866 -828
rect 9824 -866 9854 -844
rect 9908 -866 9938 -736
rect 10003 -854 10033 -670
rect 10111 -749 10141 -572
rect 10478 -556 10508 -457
rect 12852 -458 12918 -442
rect 15244 -442 15260 -408
rect 15294 -442 15310 -408
rect 17636 -407 17702 -391
rect 15244 -458 15310 -442
rect 17636 -441 17652 -407
rect 17686 -441 17702 -407
rect 20028 -407 20094 -391
rect 17636 -457 17702 -441
rect 20028 -441 20044 -407
rect 20078 -441 20094 -407
rect 22420 -408 22486 -392
rect 20028 -457 20094 -441
rect 22420 -442 22436 -408
rect 22470 -442 22486 -408
rect 24812 -408 24878 -392
rect 10575 -488 10605 -462
rect 10217 -704 10247 -656
rect 10076 -772 10141 -749
rect 10183 -720 10247 -704
rect 10183 -754 10193 -720
rect 10227 -754 10247 -720
rect 10289 -688 10319 -656
rect 10289 -704 10373 -688
rect 10289 -738 10329 -704
rect 10363 -738 10373 -704
rect 10478 -716 10508 -684
rect 10763 -504 10793 -478
rect 10858 -488 10888 -462
rect 10763 -648 10793 -632
rect 10738 -678 10793 -648
rect 10289 -754 10373 -738
rect 10428 -732 10510 -716
rect 10575 -720 10605 -688
rect 10183 -770 10247 -754
rect 10076 -806 10086 -772
rect 10120 -779 10141 -772
rect 10120 -806 10130 -779
rect 10076 -822 10130 -806
rect 10208 -810 10238 -770
rect 10292 -810 10322 -754
rect 10428 -766 10438 -732
rect 10472 -766 10510 -732
rect 10428 -782 10510 -766
rect 10100 -854 10130 -822
rect 10480 -854 10510 -782
rect 10556 -726 10610 -720
rect 10738 -726 10768 -678
rect 11046 -494 11076 -468
rect 11130 -494 11160 -468
rect 11318 -488 11348 -462
rect 11410 -488 11440 -462
rect 11494 -488 11524 -462
rect 11614 -488 11644 -462
rect 11720 -488 11750 -462
rect 11828 -488 11858 -462
rect 11912 -488 11942 -462
rect 12049 -488 12079 -462
rect 12193 -488 12223 -462
rect 12277 -488 12307 -462
rect 12382 -488 12412 -462
rect 12503 -488 12533 -462
rect 12609 -488 12639 -462
rect 12681 -488 12711 -462
rect 11046 -637 11076 -622
rect 11012 -667 11076 -637
rect 10858 -720 10888 -688
rect 11012 -705 11042 -667
rect 10556 -736 10768 -726
rect 10556 -770 10566 -736
rect 10600 -770 10768 -736
rect 10556 -780 10768 -770
rect 10556 -786 10605 -780
rect 10575 -808 10605 -786
rect 10738 -809 10768 -780
rect 10830 -736 10889 -720
rect 10830 -770 10840 -736
rect 10874 -770 10889 -736
rect 10830 -786 10889 -770
rect 10988 -721 11042 -705
rect 11130 -711 11160 -622
rect 10988 -755 10998 -721
rect 11032 -755 11042 -721
rect 10988 -771 11042 -755
rect 11084 -721 11160 -711
rect 11318 -718 11348 -572
rect 11410 -706 11440 -572
rect 11494 -610 11524 -572
rect 11614 -604 11644 -572
rect 11482 -620 11548 -610
rect 11482 -654 11498 -620
rect 11532 -654 11548 -620
rect 11482 -664 11548 -654
rect 11614 -620 11678 -604
rect 11614 -654 11634 -620
rect 11668 -654 11678 -620
rect 11614 -670 11678 -654
rect 11084 -755 11100 -721
rect 11134 -755 11160 -721
rect 11084 -765 11160 -755
rect 10858 -808 10888 -786
rect 10738 -839 10793 -809
rect 10763 -854 10793 -839
rect 11012 -809 11042 -771
rect 11012 -839 11076 -809
rect 11046 -854 11076 -839
rect 11130 -854 11160 -765
rect 11306 -734 11360 -718
rect 11306 -768 11316 -734
rect 11350 -768 11360 -734
rect 11410 -736 11548 -706
rect 11306 -784 11360 -768
rect 11518 -766 11548 -736
rect 11318 -854 11348 -784
rect 11413 -794 11476 -778
rect 11413 -828 11432 -794
rect 11466 -828 11476 -794
rect 11413 -844 11476 -828
rect 11518 -782 11572 -766
rect 11518 -816 11528 -782
rect 11562 -816 11572 -782
rect 11518 -832 11572 -816
rect 11413 -866 11443 -844
rect 11518 -866 11548 -832
rect 11614 -854 11644 -670
rect 11720 -756 11750 -572
rect 12193 -604 12223 -572
rect 12169 -620 12223 -604
rect 12277 -610 12307 -572
rect 12382 -604 12412 -572
rect 12169 -654 12179 -620
rect 12213 -654 12223 -620
rect 11828 -688 11858 -656
rect 11912 -688 11942 -656
rect 11792 -704 11858 -688
rect 11792 -738 11802 -704
rect 11836 -738 11858 -704
rect 11792 -754 11858 -738
rect 11908 -704 11998 -688
rect 11908 -738 11954 -704
rect 11988 -738 11998 -704
rect 11908 -754 11998 -738
rect 12049 -722 12079 -656
rect 12169 -670 12223 -654
rect 12265 -620 12331 -610
rect 12265 -654 12281 -620
rect 12315 -654 12331 -620
rect 12265 -664 12331 -654
rect 12382 -620 12461 -604
rect 12382 -654 12417 -620
rect 12451 -654 12461 -620
rect 12382 -670 12461 -654
rect 12193 -706 12223 -670
rect 12049 -738 12126 -722
rect 12193 -736 12330 -706
rect 12049 -752 12082 -738
rect 11690 -772 11750 -756
rect 11690 -806 11700 -772
rect 11734 -792 11750 -772
rect 11734 -806 11758 -792
rect 11690 -822 11758 -806
rect 11824 -810 11854 -754
rect 11908 -810 11938 -754
rect 12072 -772 12082 -752
rect 12116 -772 12126 -738
rect 12072 -788 12126 -772
rect 12096 -810 12126 -788
rect 12204 -794 12258 -778
rect 11728 -854 11758 -822
rect 12204 -828 12214 -794
rect 12248 -828 12258 -794
rect 12204 -844 12258 -828
rect 12216 -866 12246 -844
rect 12300 -866 12330 -736
rect 12395 -854 12425 -670
rect 12503 -749 12533 -572
rect 12870 -556 12900 -458
rect 12967 -488 12997 -462
rect 12609 -704 12639 -656
rect 12468 -772 12533 -749
rect 12575 -720 12639 -704
rect 12575 -754 12585 -720
rect 12619 -754 12639 -720
rect 12681 -688 12711 -656
rect 12681 -704 12765 -688
rect 12681 -738 12721 -704
rect 12755 -738 12765 -704
rect 12870 -716 12900 -684
rect 13155 -504 13185 -478
rect 13250 -488 13280 -462
rect 13155 -648 13185 -632
rect 13130 -678 13185 -648
rect 12681 -754 12765 -738
rect 12820 -732 12902 -716
rect 12967 -720 12997 -688
rect 12575 -770 12639 -754
rect 12468 -806 12478 -772
rect 12512 -779 12533 -772
rect 12512 -806 12522 -779
rect 12468 -822 12522 -806
rect 12600 -810 12630 -770
rect 12684 -810 12714 -754
rect 12820 -766 12830 -732
rect 12864 -766 12902 -732
rect 12820 -782 12902 -766
rect 12492 -854 12522 -822
rect 12872 -854 12902 -782
rect 12948 -726 13002 -720
rect 13130 -726 13160 -678
rect 13438 -494 13468 -468
rect 13522 -494 13552 -468
rect 13710 -488 13740 -462
rect 13802 -488 13832 -462
rect 13886 -488 13916 -462
rect 14006 -488 14036 -462
rect 14112 -488 14142 -462
rect 14220 -488 14250 -462
rect 14304 -488 14334 -462
rect 14441 -488 14471 -462
rect 14585 -488 14615 -462
rect 14669 -488 14699 -462
rect 14774 -488 14804 -462
rect 14895 -488 14925 -462
rect 15001 -488 15031 -462
rect 15073 -488 15103 -462
rect 13438 -637 13468 -622
rect 13404 -667 13468 -637
rect 13250 -720 13280 -688
rect 13404 -705 13434 -667
rect 12948 -736 13160 -726
rect 12948 -770 12958 -736
rect 12992 -770 13160 -736
rect 12948 -780 13160 -770
rect 12948 -786 12997 -780
rect 12967 -808 12997 -786
rect 13130 -809 13160 -780
rect 13222 -736 13281 -720
rect 13222 -770 13232 -736
rect 13266 -770 13281 -736
rect 13222 -786 13281 -770
rect 13380 -721 13434 -705
rect 13522 -711 13552 -622
rect 13380 -755 13390 -721
rect 13424 -755 13434 -721
rect 13380 -771 13434 -755
rect 13476 -721 13552 -711
rect 13710 -718 13740 -572
rect 13802 -706 13832 -572
rect 13886 -610 13916 -572
rect 14006 -604 14036 -572
rect 13874 -620 13940 -610
rect 13874 -654 13890 -620
rect 13924 -654 13940 -620
rect 13874 -664 13940 -654
rect 14006 -620 14070 -604
rect 14006 -654 14026 -620
rect 14060 -654 14070 -620
rect 14006 -670 14070 -654
rect 13476 -755 13492 -721
rect 13526 -755 13552 -721
rect 13476 -765 13552 -755
rect 13250 -808 13280 -786
rect 13130 -839 13185 -809
rect 13155 -854 13185 -839
rect 13404 -809 13434 -771
rect 13404 -839 13468 -809
rect 13438 -854 13468 -839
rect 13522 -854 13552 -765
rect 13698 -734 13752 -718
rect 13698 -768 13708 -734
rect 13742 -768 13752 -734
rect 13802 -736 13940 -706
rect 13698 -784 13752 -768
rect 13910 -766 13940 -736
rect 13710 -854 13740 -784
rect 13805 -794 13868 -778
rect 13805 -828 13824 -794
rect 13858 -828 13868 -794
rect 13805 -844 13868 -828
rect 13910 -782 13964 -766
rect 13910 -816 13920 -782
rect 13954 -816 13964 -782
rect 13910 -832 13964 -816
rect 13805 -866 13835 -844
rect 13910 -866 13940 -832
rect 14006 -854 14036 -670
rect 14112 -756 14142 -572
rect 14585 -604 14615 -572
rect 14561 -620 14615 -604
rect 14669 -610 14699 -572
rect 14774 -604 14804 -572
rect 14561 -654 14571 -620
rect 14605 -654 14615 -620
rect 14220 -688 14250 -656
rect 14304 -688 14334 -656
rect 14184 -704 14250 -688
rect 14184 -738 14194 -704
rect 14228 -738 14250 -704
rect 14184 -754 14250 -738
rect 14300 -704 14390 -688
rect 14300 -738 14346 -704
rect 14380 -738 14390 -704
rect 14300 -754 14390 -738
rect 14441 -722 14471 -656
rect 14561 -670 14615 -654
rect 14657 -620 14723 -610
rect 14657 -654 14673 -620
rect 14707 -654 14723 -620
rect 14657 -664 14723 -654
rect 14774 -620 14853 -604
rect 14774 -654 14809 -620
rect 14843 -654 14853 -620
rect 14774 -670 14853 -654
rect 14585 -706 14615 -670
rect 14441 -738 14518 -722
rect 14585 -736 14722 -706
rect 14441 -752 14474 -738
rect 14082 -772 14142 -756
rect 14082 -806 14092 -772
rect 14126 -792 14142 -772
rect 14126 -806 14150 -792
rect 14082 -822 14150 -806
rect 14216 -810 14246 -754
rect 14300 -810 14330 -754
rect 14464 -772 14474 -752
rect 14508 -772 14518 -738
rect 14464 -788 14518 -772
rect 14488 -810 14518 -788
rect 14596 -794 14650 -778
rect 14120 -854 14150 -822
rect 14596 -828 14606 -794
rect 14640 -828 14650 -794
rect 14596 -844 14650 -828
rect 14608 -866 14638 -844
rect 14692 -866 14722 -736
rect 14787 -854 14817 -670
rect 14895 -749 14925 -572
rect 15262 -556 15292 -458
rect 15359 -488 15389 -462
rect 15001 -704 15031 -656
rect 14860 -772 14925 -749
rect 14967 -720 15031 -704
rect 14967 -754 14977 -720
rect 15011 -754 15031 -720
rect 15073 -688 15103 -656
rect 15073 -704 15157 -688
rect 15073 -738 15113 -704
rect 15147 -738 15157 -704
rect 15262 -716 15292 -684
rect 15547 -504 15577 -478
rect 15642 -488 15672 -462
rect 15547 -648 15577 -632
rect 15522 -678 15577 -648
rect 15073 -754 15157 -738
rect 15212 -732 15294 -716
rect 15359 -720 15389 -688
rect 14967 -770 15031 -754
rect 14860 -806 14870 -772
rect 14904 -779 14925 -772
rect 14904 -806 14914 -779
rect 14860 -822 14914 -806
rect 14992 -810 15022 -770
rect 15076 -810 15106 -754
rect 15212 -766 15222 -732
rect 15256 -766 15294 -732
rect 15212 -782 15294 -766
rect 14884 -854 14914 -822
rect 15264 -854 15294 -782
rect 15340 -726 15394 -720
rect 15522 -726 15552 -678
rect 15830 -494 15860 -468
rect 15914 -494 15944 -468
rect 16102 -488 16132 -462
rect 16194 -488 16224 -462
rect 16278 -488 16308 -462
rect 16398 -488 16428 -462
rect 16504 -488 16534 -462
rect 16612 -488 16642 -462
rect 16696 -488 16726 -462
rect 16833 -488 16863 -462
rect 16977 -488 17007 -462
rect 17061 -488 17091 -462
rect 17166 -488 17196 -462
rect 17287 -488 17317 -462
rect 17393 -488 17423 -462
rect 17465 -488 17495 -462
rect 15830 -637 15860 -622
rect 15796 -667 15860 -637
rect 15642 -720 15672 -688
rect 15796 -705 15826 -667
rect 15340 -736 15552 -726
rect 15340 -770 15350 -736
rect 15384 -770 15552 -736
rect 15340 -780 15552 -770
rect 15340 -786 15389 -780
rect 15359 -808 15389 -786
rect 15522 -809 15552 -780
rect 15614 -736 15673 -720
rect 15614 -770 15624 -736
rect 15658 -770 15673 -736
rect 15614 -786 15673 -770
rect 15772 -721 15826 -705
rect 15914 -711 15944 -622
rect 15772 -755 15782 -721
rect 15816 -755 15826 -721
rect 15772 -771 15826 -755
rect 15868 -721 15944 -711
rect 16102 -718 16132 -572
rect 16194 -706 16224 -572
rect 16278 -610 16308 -572
rect 16398 -604 16428 -572
rect 16266 -620 16332 -610
rect 16266 -654 16282 -620
rect 16316 -654 16332 -620
rect 16266 -664 16332 -654
rect 16398 -620 16462 -604
rect 16398 -654 16418 -620
rect 16452 -654 16462 -620
rect 16398 -670 16462 -654
rect 15868 -755 15884 -721
rect 15918 -755 15944 -721
rect 15868 -765 15944 -755
rect 15642 -808 15672 -786
rect 15522 -839 15577 -809
rect 15547 -854 15577 -839
rect 15796 -809 15826 -771
rect 15796 -839 15860 -809
rect 15830 -854 15860 -839
rect 15914 -854 15944 -765
rect 16090 -734 16144 -718
rect 16090 -768 16100 -734
rect 16134 -768 16144 -734
rect 16194 -736 16332 -706
rect 16090 -784 16144 -768
rect 16302 -766 16332 -736
rect 16102 -854 16132 -784
rect 16197 -794 16260 -778
rect 16197 -828 16216 -794
rect 16250 -828 16260 -794
rect 16197 -844 16260 -828
rect 16302 -782 16356 -766
rect 16302 -816 16312 -782
rect 16346 -816 16356 -782
rect 16302 -832 16356 -816
rect 16197 -866 16227 -844
rect 16302 -866 16332 -832
rect 16398 -854 16428 -670
rect 16504 -756 16534 -572
rect 16977 -604 17007 -572
rect 16953 -620 17007 -604
rect 17061 -610 17091 -572
rect 17166 -604 17196 -572
rect 16953 -654 16963 -620
rect 16997 -654 17007 -620
rect 16612 -688 16642 -656
rect 16696 -688 16726 -656
rect 16576 -704 16642 -688
rect 16576 -738 16586 -704
rect 16620 -738 16642 -704
rect 16576 -754 16642 -738
rect 16692 -704 16782 -688
rect 16692 -738 16738 -704
rect 16772 -738 16782 -704
rect 16692 -754 16782 -738
rect 16833 -722 16863 -656
rect 16953 -670 17007 -654
rect 17049 -620 17115 -610
rect 17049 -654 17065 -620
rect 17099 -654 17115 -620
rect 17049 -664 17115 -654
rect 17166 -620 17245 -604
rect 17166 -654 17201 -620
rect 17235 -654 17245 -620
rect 17166 -670 17245 -654
rect 16977 -706 17007 -670
rect 16833 -738 16910 -722
rect 16977 -736 17114 -706
rect 16833 -752 16866 -738
rect 16474 -772 16534 -756
rect 16474 -806 16484 -772
rect 16518 -792 16534 -772
rect 16518 -806 16542 -792
rect 16474 -822 16542 -806
rect 16608 -810 16638 -754
rect 16692 -810 16722 -754
rect 16856 -772 16866 -752
rect 16900 -772 16910 -738
rect 16856 -788 16910 -772
rect 16880 -810 16910 -788
rect 16988 -794 17042 -778
rect 16512 -854 16542 -822
rect 16988 -828 16998 -794
rect 17032 -828 17042 -794
rect 16988 -844 17042 -828
rect 17000 -866 17030 -844
rect 17084 -866 17114 -736
rect 17179 -854 17209 -670
rect 17287 -749 17317 -572
rect 17654 -556 17684 -457
rect 17751 -488 17781 -462
rect 17393 -704 17423 -656
rect 17252 -772 17317 -749
rect 17359 -720 17423 -704
rect 17359 -754 17369 -720
rect 17403 -754 17423 -720
rect 17465 -688 17495 -656
rect 17465 -704 17549 -688
rect 17465 -738 17505 -704
rect 17539 -738 17549 -704
rect 17654 -716 17684 -684
rect 17939 -504 17969 -478
rect 18034 -488 18064 -462
rect 17939 -648 17969 -632
rect 17914 -678 17969 -648
rect 17465 -754 17549 -738
rect 17604 -732 17686 -716
rect 17751 -720 17781 -688
rect 17359 -770 17423 -754
rect 17252 -806 17262 -772
rect 17296 -779 17317 -772
rect 17296 -806 17306 -779
rect 17252 -822 17306 -806
rect 17384 -810 17414 -770
rect 17468 -810 17498 -754
rect 17604 -766 17614 -732
rect 17648 -766 17686 -732
rect 17604 -782 17686 -766
rect 17276 -854 17306 -822
rect 17656 -854 17686 -782
rect 17732 -726 17786 -720
rect 17914 -726 17944 -678
rect 18222 -494 18252 -468
rect 18306 -494 18336 -468
rect 18494 -488 18524 -462
rect 18586 -488 18616 -462
rect 18670 -488 18700 -462
rect 18790 -488 18820 -462
rect 18896 -488 18926 -462
rect 19004 -488 19034 -462
rect 19088 -488 19118 -462
rect 19225 -488 19255 -462
rect 19369 -488 19399 -462
rect 19453 -488 19483 -462
rect 19558 -488 19588 -462
rect 19679 -488 19709 -462
rect 19785 -488 19815 -462
rect 19857 -488 19887 -462
rect 18222 -637 18252 -622
rect 18188 -667 18252 -637
rect 18034 -720 18064 -688
rect 18188 -705 18218 -667
rect 17732 -736 17944 -726
rect 17732 -770 17742 -736
rect 17776 -770 17944 -736
rect 17732 -780 17944 -770
rect 17732 -786 17781 -780
rect 17751 -808 17781 -786
rect 17914 -809 17944 -780
rect 18006 -736 18065 -720
rect 18006 -770 18016 -736
rect 18050 -770 18065 -736
rect 18006 -786 18065 -770
rect 18164 -721 18218 -705
rect 18306 -711 18336 -622
rect 18164 -755 18174 -721
rect 18208 -755 18218 -721
rect 18164 -771 18218 -755
rect 18260 -721 18336 -711
rect 18494 -718 18524 -572
rect 18586 -706 18616 -572
rect 18670 -610 18700 -572
rect 18790 -604 18820 -572
rect 18658 -620 18724 -610
rect 18658 -654 18674 -620
rect 18708 -654 18724 -620
rect 18658 -664 18724 -654
rect 18790 -620 18854 -604
rect 18790 -654 18810 -620
rect 18844 -654 18854 -620
rect 18790 -670 18854 -654
rect 18260 -755 18276 -721
rect 18310 -755 18336 -721
rect 18260 -765 18336 -755
rect 18034 -808 18064 -786
rect 17914 -839 17969 -809
rect 17939 -854 17969 -839
rect 18188 -809 18218 -771
rect 18188 -839 18252 -809
rect 18222 -854 18252 -839
rect 18306 -854 18336 -765
rect 18482 -734 18536 -718
rect 18482 -768 18492 -734
rect 18526 -768 18536 -734
rect 18586 -736 18724 -706
rect 18482 -784 18536 -768
rect 18694 -766 18724 -736
rect 18494 -854 18524 -784
rect 18589 -794 18652 -778
rect 18589 -828 18608 -794
rect 18642 -828 18652 -794
rect 18589 -844 18652 -828
rect 18694 -782 18748 -766
rect 18694 -816 18704 -782
rect 18738 -816 18748 -782
rect 18694 -832 18748 -816
rect 18589 -866 18619 -844
rect 18694 -866 18724 -832
rect 18790 -854 18820 -670
rect 18896 -756 18926 -572
rect 19369 -604 19399 -572
rect 19345 -620 19399 -604
rect 19453 -610 19483 -572
rect 19558 -604 19588 -572
rect 19345 -654 19355 -620
rect 19389 -654 19399 -620
rect 19004 -688 19034 -656
rect 19088 -688 19118 -656
rect 18968 -704 19034 -688
rect 18968 -738 18978 -704
rect 19012 -738 19034 -704
rect 18968 -754 19034 -738
rect 19084 -704 19174 -688
rect 19084 -738 19130 -704
rect 19164 -738 19174 -704
rect 19084 -754 19174 -738
rect 19225 -722 19255 -656
rect 19345 -670 19399 -654
rect 19441 -620 19507 -610
rect 19441 -654 19457 -620
rect 19491 -654 19507 -620
rect 19441 -664 19507 -654
rect 19558 -620 19637 -604
rect 19558 -654 19593 -620
rect 19627 -654 19637 -620
rect 19558 -670 19637 -654
rect 19369 -706 19399 -670
rect 19225 -738 19302 -722
rect 19369 -736 19506 -706
rect 19225 -752 19258 -738
rect 18866 -772 18926 -756
rect 18866 -806 18876 -772
rect 18910 -792 18926 -772
rect 18910 -806 18934 -792
rect 18866 -822 18934 -806
rect 19000 -810 19030 -754
rect 19084 -810 19114 -754
rect 19248 -772 19258 -752
rect 19292 -772 19302 -738
rect 19248 -788 19302 -772
rect 19272 -810 19302 -788
rect 19380 -794 19434 -778
rect 18904 -854 18934 -822
rect 19380 -828 19390 -794
rect 19424 -828 19434 -794
rect 19380 -844 19434 -828
rect 19392 -866 19422 -844
rect 19476 -866 19506 -736
rect 19571 -854 19601 -670
rect 19679 -749 19709 -572
rect 20046 -556 20076 -457
rect 22420 -458 22486 -442
rect 24812 -442 24828 -408
rect 24862 -442 24878 -408
rect 24812 -458 24878 -442
rect 20143 -488 20173 -462
rect 19785 -704 19815 -656
rect 19644 -772 19709 -749
rect 19751 -720 19815 -704
rect 19751 -754 19761 -720
rect 19795 -754 19815 -720
rect 19857 -688 19887 -656
rect 19857 -704 19941 -688
rect 19857 -738 19897 -704
rect 19931 -738 19941 -704
rect 20046 -716 20076 -684
rect 20331 -504 20361 -478
rect 20426 -488 20456 -462
rect 20331 -648 20361 -632
rect 20306 -678 20361 -648
rect 19857 -754 19941 -738
rect 19996 -732 20078 -716
rect 20143 -720 20173 -688
rect 19751 -770 19815 -754
rect 19644 -806 19654 -772
rect 19688 -779 19709 -772
rect 19688 -806 19698 -779
rect 19644 -822 19698 -806
rect 19776 -810 19806 -770
rect 19860 -810 19890 -754
rect 19996 -766 20006 -732
rect 20040 -766 20078 -732
rect 19996 -782 20078 -766
rect 19668 -854 19698 -822
rect 20048 -854 20078 -782
rect 20124 -726 20178 -720
rect 20306 -726 20336 -678
rect 20614 -494 20644 -468
rect 20698 -494 20728 -468
rect 20886 -488 20916 -462
rect 20978 -488 21008 -462
rect 21062 -488 21092 -462
rect 21182 -488 21212 -462
rect 21288 -488 21318 -462
rect 21396 -488 21426 -462
rect 21480 -488 21510 -462
rect 21617 -488 21647 -462
rect 21761 -488 21791 -462
rect 21845 -488 21875 -462
rect 21950 -488 21980 -462
rect 22071 -488 22101 -462
rect 22177 -488 22207 -462
rect 22249 -488 22279 -462
rect 20614 -637 20644 -622
rect 20580 -667 20644 -637
rect 20426 -720 20456 -688
rect 20580 -705 20610 -667
rect 20124 -736 20336 -726
rect 20124 -770 20134 -736
rect 20168 -770 20336 -736
rect 20124 -780 20336 -770
rect 20124 -786 20173 -780
rect 20143 -808 20173 -786
rect 20306 -809 20336 -780
rect 20398 -736 20457 -720
rect 20398 -770 20408 -736
rect 20442 -770 20457 -736
rect 20398 -786 20457 -770
rect 20556 -721 20610 -705
rect 20698 -711 20728 -622
rect 20556 -755 20566 -721
rect 20600 -755 20610 -721
rect 20556 -771 20610 -755
rect 20652 -721 20728 -711
rect 20886 -718 20916 -572
rect 20978 -706 21008 -572
rect 21062 -610 21092 -572
rect 21182 -604 21212 -572
rect 21050 -620 21116 -610
rect 21050 -654 21066 -620
rect 21100 -654 21116 -620
rect 21050 -664 21116 -654
rect 21182 -620 21246 -604
rect 21182 -654 21202 -620
rect 21236 -654 21246 -620
rect 21182 -670 21246 -654
rect 20652 -755 20668 -721
rect 20702 -755 20728 -721
rect 20652 -765 20728 -755
rect 20426 -808 20456 -786
rect 20306 -839 20361 -809
rect 20331 -854 20361 -839
rect 20580 -809 20610 -771
rect 20580 -839 20644 -809
rect 20614 -854 20644 -839
rect 20698 -854 20728 -765
rect 20874 -734 20928 -718
rect 20874 -768 20884 -734
rect 20918 -768 20928 -734
rect 20978 -736 21116 -706
rect 20874 -784 20928 -768
rect 21086 -766 21116 -736
rect 20886 -854 20916 -784
rect 20981 -794 21044 -778
rect 20981 -828 21000 -794
rect 21034 -828 21044 -794
rect 20981 -844 21044 -828
rect 21086 -782 21140 -766
rect 21086 -816 21096 -782
rect 21130 -816 21140 -782
rect 21086 -832 21140 -816
rect 20981 -866 21011 -844
rect 21086 -866 21116 -832
rect 21182 -854 21212 -670
rect 21288 -756 21318 -572
rect 21761 -604 21791 -572
rect 21737 -620 21791 -604
rect 21845 -610 21875 -572
rect 21950 -604 21980 -572
rect 21737 -654 21747 -620
rect 21781 -654 21791 -620
rect 21396 -688 21426 -656
rect 21480 -688 21510 -656
rect 21360 -704 21426 -688
rect 21360 -738 21370 -704
rect 21404 -738 21426 -704
rect 21360 -754 21426 -738
rect 21476 -704 21566 -688
rect 21476 -738 21522 -704
rect 21556 -738 21566 -704
rect 21476 -754 21566 -738
rect 21617 -722 21647 -656
rect 21737 -670 21791 -654
rect 21833 -620 21899 -610
rect 21833 -654 21849 -620
rect 21883 -654 21899 -620
rect 21833 -664 21899 -654
rect 21950 -620 22029 -604
rect 21950 -654 21985 -620
rect 22019 -654 22029 -620
rect 21950 -670 22029 -654
rect 21761 -706 21791 -670
rect 21617 -738 21694 -722
rect 21761 -736 21898 -706
rect 21617 -752 21650 -738
rect 21258 -772 21318 -756
rect 21258 -806 21268 -772
rect 21302 -792 21318 -772
rect 21302 -806 21326 -792
rect 21258 -822 21326 -806
rect 21392 -810 21422 -754
rect 21476 -810 21506 -754
rect 21640 -772 21650 -752
rect 21684 -772 21694 -738
rect 21640 -788 21694 -772
rect 21664 -810 21694 -788
rect 21772 -794 21826 -778
rect 21296 -854 21326 -822
rect 21772 -828 21782 -794
rect 21816 -828 21826 -794
rect 21772 -844 21826 -828
rect 21784 -866 21814 -844
rect 21868 -866 21898 -736
rect 21963 -854 21993 -670
rect 22071 -749 22101 -572
rect 22438 -556 22468 -458
rect 22535 -488 22565 -462
rect 22177 -704 22207 -656
rect 22036 -772 22101 -749
rect 22143 -720 22207 -704
rect 22143 -754 22153 -720
rect 22187 -754 22207 -720
rect 22249 -688 22279 -656
rect 22249 -704 22333 -688
rect 22249 -738 22289 -704
rect 22323 -738 22333 -704
rect 22438 -716 22468 -684
rect 22723 -504 22753 -478
rect 22818 -488 22848 -462
rect 22723 -648 22753 -632
rect 22698 -678 22753 -648
rect 22249 -754 22333 -738
rect 22388 -732 22470 -716
rect 22535 -720 22565 -688
rect 22143 -770 22207 -754
rect 22036 -806 22046 -772
rect 22080 -779 22101 -772
rect 22080 -806 22090 -779
rect 22036 -822 22090 -806
rect 22168 -810 22198 -770
rect 22252 -810 22282 -754
rect 22388 -766 22398 -732
rect 22432 -766 22470 -732
rect 22388 -782 22470 -766
rect 22060 -854 22090 -822
rect 22440 -854 22470 -782
rect 22516 -726 22570 -720
rect 22698 -726 22728 -678
rect 23006 -494 23036 -468
rect 23090 -494 23120 -468
rect 23278 -488 23308 -462
rect 23370 -488 23400 -462
rect 23454 -488 23484 -462
rect 23574 -488 23604 -462
rect 23680 -488 23710 -462
rect 23788 -488 23818 -462
rect 23872 -488 23902 -462
rect 24009 -488 24039 -462
rect 24153 -488 24183 -462
rect 24237 -488 24267 -462
rect 24342 -488 24372 -462
rect 24463 -488 24493 -462
rect 24569 -488 24599 -462
rect 24641 -488 24671 -462
rect 23006 -637 23036 -622
rect 22972 -667 23036 -637
rect 22818 -720 22848 -688
rect 22972 -705 23002 -667
rect 22516 -736 22728 -726
rect 22516 -770 22526 -736
rect 22560 -770 22728 -736
rect 22516 -780 22728 -770
rect 22516 -786 22565 -780
rect 22535 -808 22565 -786
rect 22698 -809 22728 -780
rect 22790 -736 22849 -720
rect 22790 -770 22800 -736
rect 22834 -770 22849 -736
rect 22790 -786 22849 -770
rect 22948 -721 23002 -705
rect 23090 -711 23120 -622
rect 22948 -755 22958 -721
rect 22992 -755 23002 -721
rect 22948 -771 23002 -755
rect 23044 -721 23120 -711
rect 23278 -718 23308 -572
rect 23370 -706 23400 -572
rect 23454 -610 23484 -572
rect 23574 -604 23604 -572
rect 23442 -620 23508 -610
rect 23442 -654 23458 -620
rect 23492 -654 23508 -620
rect 23442 -664 23508 -654
rect 23574 -620 23638 -604
rect 23574 -654 23594 -620
rect 23628 -654 23638 -620
rect 23574 -670 23638 -654
rect 23044 -755 23060 -721
rect 23094 -755 23120 -721
rect 23044 -765 23120 -755
rect 22818 -808 22848 -786
rect 22698 -839 22753 -809
rect 22723 -854 22753 -839
rect 22972 -809 23002 -771
rect 22972 -839 23036 -809
rect 23006 -854 23036 -839
rect 23090 -854 23120 -765
rect 23266 -734 23320 -718
rect 23266 -768 23276 -734
rect 23310 -768 23320 -734
rect 23370 -736 23508 -706
rect 23266 -784 23320 -768
rect 23478 -766 23508 -736
rect 23278 -854 23308 -784
rect 23373 -794 23436 -778
rect 23373 -828 23392 -794
rect 23426 -828 23436 -794
rect 23373 -844 23436 -828
rect 23478 -782 23532 -766
rect 23478 -816 23488 -782
rect 23522 -816 23532 -782
rect 23478 -832 23532 -816
rect 23373 -866 23403 -844
rect 23478 -866 23508 -832
rect 23574 -854 23604 -670
rect 23680 -756 23710 -572
rect 24153 -604 24183 -572
rect 24129 -620 24183 -604
rect 24237 -610 24267 -572
rect 24342 -604 24372 -572
rect 24129 -654 24139 -620
rect 24173 -654 24183 -620
rect 23788 -688 23818 -656
rect 23872 -688 23902 -656
rect 23752 -704 23818 -688
rect 23752 -738 23762 -704
rect 23796 -738 23818 -704
rect 23752 -754 23818 -738
rect 23868 -704 23958 -688
rect 23868 -738 23914 -704
rect 23948 -738 23958 -704
rect 23868 -754 23958 -738
rect 24009 -722 24039 -656
rect 24129 -670 24183 -654
rect 24225 -620 24291 -610
rect 24225 -654 24241 -620
rect 24275 -654 24291 -620
rect 24225 -664 24291 -654
rect 24342 -620 24421 -604
rect 24342 -654 24377 -620
rect 24411 -654 24421 -620
rect 24342 -670 24421 -654
rect 24153 -706 24183 -670
rect 24009 -738 24086 -722
rect 24153 -736 24290 -706
rect 24009 -752 24042 -738
rect 23650 -772 23710 -756
rect 23650 -806 23660 -772
rect 23694 -792 23710 -772
rect 23694 -806 23718 -792
rect 23650 -822 23718 -806
rect 23784 -810 23814 -754
rect 23868 -810 23898 -754
rect 24032 -772 24042 -752
rect 24076 -772 24086 -738
rect 24032 -788 24086 -772
rect 24056 -810 24086 -788
rect 24164 -794 24218 -778
rect 23688 -854 23718 -822
rect 24164 -828 24174 -794
rect 24208 -828 24218 -794
rect 24164 -844 24218 -828
rect 24176 -866 24206 -844
rect 24260 -866 24290 -736
rect 24355 -854 24385 -670
rect 24463 -749 24493 -572
rect 24830 -556 24860 -458
rect 24927 -488 24957 -462
rect 24569 -704 24599 -656
rect 24428 -772 24493 -749
rect 24535 -720 24599 -704
rect 24535 -754 24545 -720
rect 24579 -754 24599 -720
rect 24641 -688 24671 -656
rect 24641 -704 24725 -688
rect 24641 -738 24681 -704
rect 24715 -738 24725 -704
rect 24830 -716 24860 -684
rect 25115 -504 25145 -478
rect 25210 -488 25240 -462
rect 25115 -648 25145 -632
rect 25090 -678 25145 -648
rect 24641 -754 24725 -738
rect 24780 -732 24862 -716
rect 24927 -720 24957 -688
rect 24535 -770 24599 -754
rect 24428 -806 24438 -772
rect 24472 -779 24493 -772
rect 24472 -806 24482 -779
rect 24428 -822 24482 -806
rect 24560 -810 24590 -770
rect 24644 -810 24674 -754
rect 24780 -766 24790 -732
rect 24824 -766 24862 -732
rect 24780 -782 24862 -766
rect 24452 -854 24482 -822
rect 24832 -854 24862 -782
rect 24908 -726 24962 -720
rect 25090 -726 25120 -678
rect 25210 -720 25240 -688
rect 24908 -736 25120 -726
rect 24908 -770 24918 -736
rect 24952 -770 25120 -736
rect 24908 -780 25120 -770
rect 24908 -786 24957 -780
rect 24927 -808 24957 -786
rect 25090 -809 25120 -780
rect 25182 -736 25241 -720
rect 25182 -770 25192 -736
rect 25226 -770 25241 -736
rect 25182 -786 25241 -770
rect 25210 -808 25240 -786
rect 25090 -839 25145 -809
rect 25115 -854 25145 -839
rect 8654 -964 8684 -938
rect 8738 -964 8768 -938
rect 8926 -964 8956 -938
rect 9021 -964 9051 -938
rect 9126 -964 9156 -938
rect 9222 -964 9252 -938
rect 9336 -964 9366 -938
rect 9432 -964 9462 -938
rect 9516 -964 9546 -938
rect 9704 -964 9734 -938
rect 9824 -964 9854 -938
rect 9908 -964 9938 -938
rect 10003 -964 10033 -938
rect 10100 -964 10130 -938
rect 10208 -964 10238 -938
rect 10292 -964 10322 -938
rect 10480 -964 10510 -938
rect 10575 -964 10605 -938
rect 10763 -964 10793 -938
rect 10858 -964 10888 -938
rect 11046 -964 11076 -938
rect 11130 -964 11160 -938
rect 11318 -964 11348 -938
rect 11413 -964 11443 -938
rect 11518 -964 11548 -938
rect 11614 -964 11644 -938
rect 11728 -964 11758 -938
rect 11824 -964 11854 -938
rect 11908 -964 11938 -938
rect 12096 -964 12126 -938
rect 12216 -964 12246 -938
rect 12300 -964 12330 -938
rect 12395 -964 12425 -938
rect 12492 -964 12522 -938
rect 12600 -964 12630 -938
rect 12684 -964 12714 -938
rect 12872 -964 12902 -938
rect 12967 -964 12997 -938
rect 13155 -964 13185 -938
rect 13250 -964 13280 -938
rect 13438 -964 13468 -938
rect 13522 -964 13552 -938
rect 13710 -964 13740 -938
rect 13805 -964 13835 -938
rect 13910 -964 13940 -938
rect 14006 -964 14036 -938
rect 14120 -964 14150 -938
rect 14216 -964 14246 -938
rect 14300 -964 14330 -938
rect 14488 -964 14518 -938
rect 14608 -964 14638 -938
rect 14692 -964 14722 -938
rect 14787 -964 14817 -938
rect 14884 -964 14914 -938
rect 14992 -964 15022 -938
rect 15076 -964 15106 -938
rect 15264 -964 15294 -938
rect 15359 -964 15389 -938
rect 15547 -964 15577 -938
rect 15642 -964 15672 -938
rect 15830 -964 15860 -938
rect 15914 -964 15944 -938
rect 16102 -964 16132 -938
rect 16197 -964 16227 -938
rect 16302 -964 16332 -938
rect 16398 -964 16428 -938
rect 16512 -964 16542 -938
rect 16608 -964 16638 -938
rect 16692 -964 16722 -938
rect 16880 -964 16910 -938
rect 17000 -964 17030 -938
rect 17084 -964 17114 -938
rect 17179 -964 17209 -938
rect 17276 -964 17306 -938
rect 17384 -964 17414 -938
rect 17468 -964 17498 -938
rect 17656 -964 17686 -938
rect 17751 -964 17781 -938
rect 17939 -964 17969 -938
rect 18034 -964 18064 -938
rect 18222 -964 18252 -938
rect 18306 -964 18336 -938
rect 18494 -964 18524 -938
rect 18589 -964 18619 -938
rect 18694 -964 18724 -938
rect 18790 -964 18820 -938
rect 18904 -964 18934 -938
rect 19000 -964 19030 -938
rect 19084 -964 19114 -938
rect 19272 -964 19302 -938
rect 19392 -964 19422 -938
rect 19476 -964 19506 -938
rect 19571 -964 19601 -938
rect 19668 -964 19698 -938
rect 19776 -964 19806 -938
rect 19860 -964 19890 -938
rect 20048 -964 20078 -938
rect 20143 -964 20173 -938
rect 20331 -964 20361 -938
rect 20426 -964 20456 -938
rect 20614 -964 20644 -938
rect 20698 -964 20728 -938
rect 20886 -964 20916 -938
rect 20981 -964 21011 -938
rect 21086 -964 21116 -938
rect 21182 -964 21212 -938
rect 21296 -964 21326 -938
rect 21392 -964 21422 -938
rect 21476 -964 21506 -938
rect 21664 -964 21694 -938
rect 21784 -964 21814 -938
rect 21868 -964 21898 -938
rect 21963 -964 21993 -938
rect 22060 -964 22090 -938
rect 22168 -964 22198 -938
rect 22252 -964 22282 -938
rect 22440 -964 22470 -938
rect 22535 -964 22565 -938
rect 22723 -964 22753 -938
rect 22818 -964 22848 -938
rect 23006 -964 23036 -938
rect 23090 -964 23120 -938
rect 23278 -964 23308 -938
rect 23373 -964 23403 -938
rect 23478 -964 23508 -938
rect 23574 -964 23604 -938
rect 23688 -964 23718 -938
rect 23784 -964 23814 -938
rect 23868 -964 23898 -938
rect 24056 -964 24086 -938
rect 24176 -964 24206 -938
rect 24260 -964 24290 -938
rect 24355 -964 24385 -938
rect 24452 -964 24482 -938
rect 24560 -964 24590 -938
rect 24644 -964 24674 -938
rect 24832 -964 24862 -938
rect 24927 -964 24957 -938
rect 25115 -964 25145 -938
rect 25210 -964 25240 -938
rect 10166 -1093 10232 -1077
rect 10166 -1127 10182 -1093
rect 10216 -1127 10232 -1093
rect 12558 -1093 12624 -1077
rect 10166 -1143 10232 -1127
rect 12558 -1127 12574 -1093
rect 12608 -1127 12624 -1093
rect 14950 -1093 15016 -1077
rect 12558 -1143 12624 -1127
rect 14950 -1127 14966 -1093
rect 15000 -1127 15016 -1093
rect 17342 -1093 17408 -1077
rect 14950 -1143 15016 -1127
rect 17342 -1127 17358 -1093
rect 17392 -1127 17408 -1093
rect 19734 -1093 19800 -1077
rect 17342 -1143 17408 -1127
rect 19734 -1127 19750 -1093
rect 19784 -1127 19800 -1093
rect 22126 -1093 22192 -1077
rect 19734 -1143 19800 -1127
rect 22126 -1127 22142 -1093
rect 22176 -1127 22192 -1093
rect 24518 -1096 24584 -1080
rect 22126 -1143 22192 -1127
rect 24518 -1130 24534 -1096
rect 24568 -1130 24584 -1096
rect 8654 -1177 8684 -1151
rect 8749 -1193 8779 -1167
rect 8937 -1177 8967 -1151
rect 9223 -1177 9253 -1151
rect 9295 -1177 9325 -1151
rect 9401 -1177 9431 -1151
rect 9522 -1177 9552 -1151
rect 9627 -1177 9657 -1151
rect 9711 -1177 9741 -1151
rect 9855 -1177 9885 -1151
rect 9992 -1177 10022 -1151
rect 10076 -1177 10106 -1151
rect 10184 -1177 10214 -1143
rect 10290 -1177 10320 -1151
rect 10410 -1177 10440 -1151
rect 10494 -1177 10524 -1151
rect 10586 -1177 10616 -1151
rect 8749 -1337 8779 -1321
rect 8749 -1367 8804 -1337
rect 8654 -1409 8684 -1377
rect 8653 -1425 8712 -1409
rect 8653 -1459 8668 -1425
rect 8702 -1459 8712 -1425
rect 8653 -1475 8712 -1459
rect 8774 -1415 8804 -1367
rect 9034 -1245 9064 -1219
rect 8937 -1409 8967 -1377
rect 9034 -1405 9064 -1373
rect 9223 -1377 9253 -1345
rect 9169 -1393 9253 -1377
rect 8932 -1415 8986 -1409
rect 8774 -1425 8986 -1415
rect 8774 -1459 8942 -1425
rect 8976 -1459 8986 -1425
rect 8774 -1469 8986 -1459
rect 8654 -1497 8684 -1475
rect 8774 -1498 8804 -1469
rect 8937 -1475 8986 -1469
rect 9032 -1421 9114 -1405
rect 9032 -1455 9070 -1421
rect 9104 -1455 9114 -1421
rect 9169 -1427 9179 -1393
rect 9213 -1427 9253 -1393
rect 9169 -1443 9253 -1427
rect 9295 -1393 9325 -1345
rect 9295 -1409 9359 -1393
rect 9295 -1443 9315 -1409
rect 9349 -1443 9359 -1409
rect 9032 -1471 9114 -1455
rect 8937 -1497 8967 -1475
rect 8749 -1528 8804 -1498
rect 8749 -1543 8779 -1528
rect 9032 -1543 9062 -1471
rect 9220 -1499 9250 -1443
rect 9295 -1459 9359 -1443
rect 9401 -1438 9431 -1261
rect 9522 -1293 9552 -1261
rect 9473 -1309 9552 -1293
rect 9627 -1299 9657 -1261
rect 9711 -1293 9741 -1261
rect 9473 -1343 9483 -1309
rect 9517 -1343 9552 -1309
rect 9473 -1359 9552 -1343
rect 9603 -1309 9669 -1299
rect 9603 -1343 9619 -1309
rect 9653 -1343 9669 -1309
rect 9603 -1353 9669 -1343
rect 9711 -1309 9765 -1293
rect 9711 -1343 9721 -1309
rect 9755 -1343 9765 -1309
rect 9711 -1359 9765 -1343
rect 10774 -1183 10804 -1157
rect 10858 -1183 10888 -1157
rect 11046 -1177 11076 -1151
rect 9304 -1499 9334 -1459
rect 9401 -1461 9466 -1438
rect 9401 -1468 9422 -1461
rect 9412 -1495 9422 -1468
rect 9456 -1495 9466 -1461
rect 9412 -1511 9466 -1495
rect 9412 -1543 9442 -1511
rect 9509 -1543 9539 -1359
rect 9711 -1395 9741 -1359
rect 9604 -1425 9741 -1395
rect 9855 -1411 9885 -1345
rect 9992 -1377 10022 -1345
rect 10076 -1377 10106 -1345
rect 9604 -1555 9634 -1425
rect 9808 -1427 9885 -1411
rect 9808 -1461 9818 -1427
rect 9852 -1441 9885 -1427
rect 9936 -1393 10026 -1377
rect 9936 -1427 9946 -1393
rect 9980 -1427 10026 -1393
rect 9852 -1461 9862 -1441
rect 9936 -1443 10026 -1427
rect 10076 -1393 10142 -1377
rect 10076 -1427 10098 -1393
rect 10132 -1427 10142 -1393
rect 10076 -1443 10142 -1427
rect 9676 -1483 9730 -1467
rect 9676 -1517 9686 -1483
rect 9720 -1517 9730 -1483
rect 9808 -1477 9862 -1461
rect 9808 -1499 9838 -1477
rect 9996 -1499 10026 -1443
rect 10080 -1499 10110 -1443
rect 10184 -1445 10214 -1261
rect 10290 -1293 10320 -1261
rect 10256 -1309 10320 -1293
rect 10410 -1299 10440 -1261
rect 10256 -1343 10266 -1309
rect 10300 -1343 10320 -1309
rect 10256 -1359 10320 -1343
rect 10386 -1309 10452 -1299
rect 10386 -1343 10402 -1309
rect 10436 -1343 10452 -1309
rect 10386 -1353 10452 -1343
rect 10184 -1461 10244 -1445
rect 10184 -1481 10200 -1461
rect 10176 -1495 10200 -1481
rect 10234 -1495 10244 -1461
rect 9676 -1533 9730 -1517
rect 9688 -1555 9718 -1533
rect 10176 -1511 10244 -1495
rect 10176 -1543 10206 -1511
rect 10290 -1543 10320 -1359
rect 10494 -1395 10524 -1261
rect 10386 -1425 10524 -1395
rect 10586 -1407 10616 -1261
rect 10774 -1400 10804 -1311
rect 10858 -1326 10888 -1311
rect 10858 -1356 10922 -1326
rect 10892 -1394 10922 -1356
rect 11141 -1193 11171 -1167
rect 11329 -1177 11359 -1151
rect 11615 -1177 11645 -1151
rect 11687 -1177 11717 -1151
rect 11793 -1177 11823 -1151
rect 11914 -1177 11944 -1151
rect 12019 -1177 12049 -1151
rect 12103 -1177 12133 -1151
rect 12247 -1177 12277 -1151
rect 12384 -1177 12414 -1151
rect 12468 -1177 12498 -1151
rect 12576 -1177 12606 -1143
rect 12682 -1177 12712 -1151
rect 12802 -1177 12832 -1151
rect 12886 -1177 12916 -1151
rect 12978 -1177 13008 -1151
rect 11141 -1337 11171 -1321
rect 11141 -1367 11196 -1337
rect 10574 -1423 10628 -1407
rect 10386 -1455 10416 -1425
rect 10362 -1471 10416 -1455
rect 10574 -1457 10584 -1423
rect 10618 -1457 10628 -1423
rect 10362 -1505 10372 -1471
rect 10406 -1505 10416 -1471
rect 10362 -1521 10416 -1505
rect 10386 -1555 10416 -1521
rect 10458 -1483 10521 -1467
rect 10574 -1473 10628 -1457
rect 10774 -1410 10850 -1400
rect 10774 -1444 10800 -1410
rect 10834 -1444 10850 -1410
rect 10774 -1454 10850 -1444
rect 10892 -1410 10946 -1394
rect 11046 -1409 11076 -1377
rect 10892 -1444 10902 -1410
rect 10936 -1444 10946 -1410
rect 10458 -1517 10468 -1483
rect 10502 -1517 10521 -1483
rect 10458 -1533 10521 -1517
rect 10491 -1555 10521 -1533
rect 10586 -1543 10616 -1473
rect 10774 -1543 10804 -1454
rect 10892 -1460 10946 -1444
rect 11045 -1425 11104 -1409
rect 11045 -1459 11060 -1425
rect 11094 -1459 11104 -1425
rect 10892 -1498 10922 -1460
rect 11045 -1475 11104 -1459
rect 11166 -1415 11196 -1367
rect 11426 -1245 11456 -1219
rect 11329 -1409 11359 -1377
rect 11426 -1405 11456 -1373
rect 11615 -1377 11645 -1345
rect 11561 -1393 11645 -1377
rect 11324 -1415 11378 -1409
rect 11166 -1425 11378 -1415
rect 11166 -1459 11334 -1425
rect 11368 -1459 11378 -1425
rect 11166 -1469 11378 -1459
rect 11046 -1497 11076 -1475
rect 10858 -1528 10922 -1498
rect 10858 -1543 10888 -1528
rect 11166 -1498 11196 -1469
rect 11329 -1475 11378 -1469
rect 11424 -1421 11506 -1405
rect 11424 -1455 11462 -1421
rect 11496 -1455 11506 -1421
rect 11561 -1427 11571 -1393
rect 11605 -1427 11645 -1393
rect 11561 -1443 11645 -1427
rect 11687 -1393 11717 -1345
rect 11687 -1409 11751 -1393
rect 11687 -1443 11707 -1409
rect 11741 -1443 11751 -1409
rect 11424 -1471 11506 -1455
rect 11329 -1497 11359 -1475
rect 11141 -1528 11196 -1498
rect 11141 -1543 11171 -1528
rect 11424 -1543 11454 -1471
rect 11612 -1499 11642 -1443
rect 11687 -1459 11751 -1443
rect 11793 -1438 11823 -1261
rect 11914 -1293 11944 -1261
rect 11865 -1309 11944 -1293
rect 12019 -1299 12049 -1261
rect 12103 -1293 12133 -1261
rect 11865 -1343 11875 -1309
rect 11909 -1343 11944 -1309
rect 11865 -1359 11944 -1343
rect 11995 -1309 12061 -1299
rect 11995 -1343 12011 -1309
rect 12045 -1343 12061 -1309
rect 11995 -1353 12061 -1343
rect 12103 -1309 12157 -1293
rect 12103 -1343 12113 -1309
rect 12147 -1343 12157 -1309
rect 12103 -1359 12157 -1343
rect 13166 -1183 13196 -1157
rect 13250 -1183 13280 -1157
rect 13438 -1177 13468 -1151
rect 11696 -1499 11726 -1459
rect 11793 -1461 11858 -1438
rect 11793 -1468 11814 -1461
rect 11804 -1495 11814 -1468
rect 11848 -1495 11858 -1461
rect 11804 -1511 11858 -1495
rect 11804 -1543 11834 -1511
rect 11901 -1543 11931 -1359
rect 12103 -1395 12133 -1359
rect 11996 -1425 12133 -1395
rect 12247 -1411 12277 -1345
rect 12384 -1377 12414 -1345
rect 12468 -1377 12498 -1345
rect 11996 -1555 12026 -1425
rect 12200 -1427 12277 -1411
rect 12200 -1461 12210 -1427
rect 12244 -1441 12277 -1427
rect 12328 -1393 12418 -1377
rect 12328 -1427 12338 -1393
rect 12372 -1427 12418 -1393
rect 12244 -1461 12254 -1441
rect 12328 -1443 12418 -1427
rect 12468 -1393 12534 -1377
rect 12468 -1427 12490 -1393
rect 12524 -1427 12534 -1393
rect 12468 -1443 12534 -1427
rect 12068 -1483 12122 -1467
rect 12068 -1517 12078 -1483
rect 12112 -1517 12122 -1483
rect 12200 -1477 12254 -1461
rect 12200 -1499 12230 -1477
rect 12388 -1499 12418 -1443
rect 12472 -1499 12502 -1443
rect 12576 -1445 12606 -1261
rect 12682 -1293 12712 -1261
rect 12648 -1309 12712 -1293
rect 12802 -1299 12832 -1261
rect 12648 -1343 12658 -1309
rect 12692 -1343 12712 -1309
rect 12648 -1359 12712 -1343
rect 12778 -1309 12844 -1299
rect 12778 -1343 12794 -1309
rect 12828 -1343 12844 -1309
rect 12778 -1353 12844 -1343
rect 12576 -1461 12636 -1445
rect 12576 -1481 12592 -1461
rect 12568 -1495 12592 -1481
rect 12626 -1495 12636 -1461
rect 12068 -1533 12122 -1517
rect 12080 -1555 12110 -1533
rect 12568 -1511 12636 -1495
rect 12568 -1543 12598 -1511
rect 12682 -1543 12712 -1359
rect 12886 -1395 12916 -1261
rect 12778 -1425 12916 -1395
rect 12978 -1407 13008 -1261
rect 13166 -1400 13196 -1311
rect 13250 -1326 13280 -1311
rect 13250 -1356 13314 -1326
rect 13284 -1394 13314 -1356
rect 13533 -1193 13563 -1167
rect 13721 -1177 13751 -1151
rect 14007 -1177 14037 -1151
rect 14079 -1177 14109 -1151
rect 14185 -1177 14215 -1151
rect 14306 -1177 14336 -1151
rect 14411 -1177 14441 -1151
rect 14495 -1177 14525 -1151
rect 14639 -1177 14669 -1151
rect 14776 -1177 14806 -1151
rect 14860 -1177 14890 -1151
rect 14968 -1177 14998 -1143
rect 15074 -1177 15104 -1151
rect 15194 -1177 15224 -1151
rect 15278 -1177 15308 -1151
rect 15370 -1177 15400 -1151
rect 13533 -1337 13563 -1321
rect 13533 -1367 13588 -1337
rect 12966 -1423 13020 -1407
rect 12778 -1455 12808 -1425
rect 12754 -1471 12808 -1455
rect 12966 -1457 12976 -1423
rect 13010 -1457 13020 -1423
rect 12754 -1505 12764 -1471
rect 12798 -1505 12808 -1471
rect 12754 -1521 12808 -1505
rect 12778 -1555 12808 -1521
rect 12850 -1483 12913 -1467
rect 12966 -1473 13020 -1457
rect 13166 -1410 13242 -1400
rect 13166 -1444 13192 -1410
rect 13226 -1444 13242 -1410
rect 13166 -1454 13242 -1444
rect 13284 -1410 13338 -1394
rect 13438 -1409 13468 -1377
rect 13284 -1444 13294 -1410
rect 13328 -1444 13338 -1410
rect 12850 -1517 12860 -1483
rect 12894 -1517 12913 -1483
rect 12850 -1533 12913 -1517
rect 12883 -1555 12913 -1533
rect 12978 -1543 13008 -1473
rect 13166 -1543 13196 -1454
rect 13284 -1460 13338 -1444
rect 13437 -1425 13496 -1409
rect 13437 -1459 13452 -1425
rect 13486 -1459 13496 -1425
rect 13284 -1498 13314 -1460
rect 13437 -1475 13496 -1459
rect 13558 -1415 13588 -1367
rect 13818 -1245 13848 -1219
rect 13721 -1409 13751 -1377
rect 13818 -1405 13848 -1373
rect 14007 -1377 14037 -1345
rect 13953 -1393 14037 -1377
rect 13716 -1415 13770 -1409
rect 13558 -1425 13770 -1415
rect 13558 -1459 13726 -1425
rect 13760 -1459 13770 -1425
rect 13558 -1469 13770 -1459
rect 13438 -1497 13468 -1475
rect 13250 -1528 13314 -1498
rect 13250 -1543 13280 -1528
rect 13558 -1498 13588 -1469
rect 13721 -1475 13770 -1469
rect 13816 -1421 13898 -1405
rect 13816 -1455 13854 -1421
rect 13888 -1455 13898 -1421
rect 13953 -1427 13963 -1393
rect 13997 -1427 14037 -1393
rect 13953 -1443 14037 -1427
rect 14079 -1393 14109 -1345
rect 14079 -1409 14143 -1393
rect 14079 -1443 14099 -1409
rect 14133 -1443 14143 -1409
rect 13816 -1471 13898 -1455
rect 13721 -1497 13751 -1475
rect 13533 -1528 13588 -1498
rect 13533 -1543 13563 -1528
rect 13816 -1543 13846 -1471
rect 14004 -1499 14034 -1443
rect 14079 -1459 14143 -1443
rect 14185 -1438 14215 -1261
rect 14306 -1293 14336 -1261
rect 14257 -1309 14336 -1293
rect 14411 -1299 14441 -1261
rect 14495 -1293 14525 -1261
rect 14257 -1343 14267 -1309
rect 14301 -1343 14336 -1309
rect 14257 -1359 14336 -1343
rect 14387 -1309 14453 -1299
rect 14387 -1343 14403 -1309
rect 14437 -1343 14453 -1309
rect 14387 -1353 14453 -1343
rect 14495 -1309 14549 -1293
rect 14495 -1343 14505 -1309
rect 14539 -1343 14549 -1309
rect 14495 -1359 14549 -1343
rect 15558 -1183 15588 -1157
rect 15642 -1183 15672 -1157
rect 15830 -1177 15860 -1151
rect 14088 -1499 14118 -1459
rect 14185 -1461 14250 -1438
rect 14185 -1468 14206 -1461
rect 14196 -1495 14206 -1468
rect 14240 -1495 14250 -1461
rect 14196 -1511 14250 -1495
rect 14196 -1543 14226 -1511
rect 14293 -1543 14323 -1359
rect 14495 -1395 14525 -1359
rect 14388 -1425 14525 -1395
rect 14639 -1411 14669 -1345
rect 14776 -1377 14806 -1345
rect 14860 -1377 14890 -1345
rect 14388 -1555 14418 -1425
rect 14592 -1427 14669 -1411
rect 14592 -1461 14602 -1427
rect 14636 -1441 14669 -1427
rect 14720 -1393 14810 -1377
rect 14720 -1427 14730 -1393
rect 14764 -1427 14810 -1393
rect 14636 -1461 14646 -1441
rect 14720 -1443 14810 -1427
rect 14860 -1393 14926 -1377
rect 14860 -1427 14882 -1393
rect 14916 -1427 14926 -1393
rect 14860 -1443 14926 -1427
rect 14460 -1483 14514 -1467
rect 14460 -1517 14470 -1483
rect 14504 -1517 14514 -1483
rect 14592 -1477 14646 -1461
rect 14592 -1499 14622 -1477
rect 14780 -1499 14810 -1443
rect 14864 -1499 14894 -1443
rect 14968 -1445 14998 -1261
rect 15074 -1293 15104 -1261
rect 15040 -1309 15104 -1293
rect 15194 -1299 15224 -1261
rect 15040 -1343 15050 -1309
rect 15084 -1343 15104 -1309
rect 15040 -1359 15104 -1343
rect 15170 -1309 15236 -1299
rect 15170 -1343 15186 -1309
rect 15220 -1343 15236 -1309
rect 15170 -1353 15236 -1343
rect 14968 -1461 15028 -1445
rect 14968 -1481 14984 -1461
rect 14960 -1495 14984 -1481
rect 15018 -1495 15028 -1461
rect 14460 -1533 14514 -1517
rect 14472 -1555 14502 -1533
rect 14960 -1511 15028 -1495
rect 14960 -1543 14990 -1511
rect 15074 -1543 15104 -1359
rect 15278 -1395 15308 -1261
rect 15170 -1425 15308 -1395
rect 15370 -1407 15400 -1261
rect 15558 -1400 15588 -1311
rect 15642 -1326 15672 -1311
rect 15642 -1356 15706 -1326
rect 15676 -1394 15706 -1356
rect 15925 -1193 15955 -1167
rect 16113 -1177 16143 -1151
rect 16399 -1177 16429 -1151
rect 16471 -1177 16501 -1151
rect 16577 -1177 16607 -1151
rect 16698 -1177 16728 -1151
rect 16803 -1177 16833 -1151
rect 16887 -1177 16917 -1151
rect 17031 -1177 17061 -1151
rect 17168 -1177 17198 -1151
rect 17252 -1177 17282 -1151
rect 17360 -1177 17390 -1143
rect 17466 -1177 17496 -1151
rect 17586 -1177 17616 -1151
rect 17670 -1177 17700 -1151
rect 17762 -1177 17792 -1151
rect 15925 -1337 15955 -1321
rect 15925 -1367 15980 -1337
rect 15358 -1423 15412 -1407
rect 15170 -1455 15200 -1425
rect 15146 -1471 15200 -1455
rect 15358 -1457 15368 -1423
rect 15402 -1457 15412 -1423
rect 15146 -1505 15156 -1471
rect 15190 -1505 15200 -1471
rect 15146 -1521 15200 -1505
rect 15170 -1555 15200 -1521
rect 15242 -1483 15305 -1467
rect 15358 -1473 15412 -1457
rect 15558 -1410 15634 -1400
rect 15558 -1444 15584 -1410
rect 15618 -1444 15634 -1410
rect 15558 -1454 15634 -1444
rect 15676 -1410 15730 -1394
rect 15830 -1409 15860 -1377
rect 15676 -1444 15686 -1410
rect 15720 -1444 15730 -1410
rect 15242 -1517 15252 -1483
rect 15286 -1517 15305 -1483
rect 15242 -1533 15305 -1517
rect 15275 -1555 15305 -1533
rect 15370 -1543 15400 -1473
rect 15558 -1543 15588 -1454
rect 15676 -1460 15730 -1444
rect 15829 -1425 15888 -1409
rect 15829 -1459 15844 -1425
rect 15878 -1459 15888 -1425
rect 15676 -1498 15706 -1460
rect 15829 -1475 15888 -1459
rect 15950 -1415 15980 -1367
rect 16210 -1245 16240 -1219
rect 16113 -1409 16143 -1377
rect 16210 -1405 16240 -1373
rect 16399 -1377 16429 -1345
rect 16345 -1393 16429 -1377
rect 16108 -1415 16162 -1409
rect 15950 -1425 16162 -1415
rect 15950 -1459 16118 -1425
rect 16152 -1459 16162 -1425
rect 15950 -1469 16162 -1459
rect 15830 -1497 15860 -1475
rect 15642 -1528 15706 -1498
rect 15642 -1543 15672 -1528
rect 15950 -1498 15980 -1469
rect 16113 -1475 16162 -1469
rect 16208 -1421 16290 -1405
rect 16208 -1455 16246 -1421
rect 16280 -1455 16290 -1421
rect 16345 -1427 16355 -1393
rect 16389 -1427 16429 -1393
rect 16345 -1443 16429 -1427
rect 16471 -1393 16501 -1345
rect 16471 -1409 16535 -1393
rect 16471 -1443 16491 -1409
rect 16525 -1443 16535 -1409
rect 16208 -1471 16290 -1455
rect 16113 -1497 16143 -1475
rect 15925 -1528 15980 -1498
rect 15925 -1543 15955 -1528
rect 16208 -1543 16238 -1471
rect 16396 -1499 16426 -1443
rect 16471 -1459 16535 -1443
rect 16577 -1438 16607 -1261
rect 16698 -1293 16728 -1261
rect 16649 -1309 16728 -1293
rect 16803 -1299 16833 -1261
rect 16887 -1293 16917 -1261
rect 16649 -1343 16659 -1309
rect 16693 -1343 16728 -1309
rect 16649 -1359 16728 -1343
rect 16779 -1309 16845 -1299
rect 16779 -1343 16795 -1309
rect 16829 -1343 16845 -1309
rect 16779 -1353 16845 -1343
rect 16887 -1309 16941 -1293
rect 16887 -1343 16897 -1309
rect 16931 -1343 16941 -1309
rect 16887 -1359 16941 -1343
rect 17950 -1183 17980 -1157
rect 18034 -1183 18064 -1157
rect 18222 -1177 18252 -1151
rect 16480 -1499 16510 -1459
rect 16577 -1461 16642 -1438
rect 16577 -1468 16598 -1461
rect 16588 -1495 16598 -1468
rect 16632 -1495 16642 -1461
rect 16588 -1511 16642 -1495
rect 16588 -1543 16618 -1511
rect 16685 -1543 16715 -1359
rect 16887 -1395 16917 -1359
rect 16780 -1425 16917 -1395
rect 17031 -1411 17061 -1345
rect 17168 -1377 17198 -1345
rect 17252 -1377 17282 -1345
rect 16780 -1555 16810 -1425
rect 16984 -1427 17061 -1411
rect 16984 -1461 16994 -1427
rect 17028 -1441 17061 -1427
rect 17112 -1393 17202 -1377
rect 17112 -1427 17122 -1393
rect 17156 -1427 17202 -1393
rect 17028 -1461 17038 -1441
rect 17112 -1443 17202 -1427
rect 17252 -1393 17318 -1377
rect 17252 -1427 17274 -1393
rect 17308 -1427 17318 -1393
rect 17252 -1443 17318 -1427
rect 16852 -1483 16906 -1467
rect 16852 -1517 16862 -1483
rect 16896 -1517 16906 -1483
rect 16984 -1477 17038 -1461
rect 16984 -1499 17014 -1477
rect 17172 -1499 17202 -1443
rect 17256 -1499 17286 -1443
rect 17360 -1445 17390 -1261
rect 17466 -1293 17496 -1261
rect 17432 -1309 17496 -1293
rect 17586 -1299 17616 -1261
rect 17432 -1343 17442 -1309
rect 17476 -1343 17496 -1309
rect 17432 -1359 17496 -1343
rect 17562 -1309 17628 -1299
rect 17562 -1343 17578 -1309
rect 17612 -1343 17628 -1309
rect 17562 -1353 17628 -1343
rect 17360 -1461 17420 -1445
rect 17360 -1481 17376 -1461
rect 17352 -1495 17376 -1481
rect 17410 -1495 17420 -1461
rect 16852 -1533 16906 -1517
rect 16864 -1555 16894 -1533
rect 17352 -1511 17420 -1495
rect 17352 -1543 17382 -1511
rect 17466 -1543 17496 -1359
rect 17670 -1395 17700 -1261
rect 17562 -1425 17700 -1395
rect 17762 -1407 17792 -1261
rect 17950 -1400 17980 -1311
rect 18034 -1326 18064 -1311
rect 18034 -1356 18098 -1326
rect 18068 -1394 18098 -1356
rect 18317 -1193 18347 -1167
rect 18505 -1177 18535 -1151
rect 18791 -1177 18821 -1151
rect 18863 -1177 18893 -1151
rect 18969 -1177 18999 -1151
rect 19090 -1177 19120 -1151
rect 19195 -1177 19225 -1151
rect 19279 -1177 19309 -1151
rect 19423 -1177 19453 -1151
rect 19560 -1177 19590 -1151
rect 19644 -1177 19674 -1151
rect 19752 -1177 19782 -1143
rect 19858 -1177 19888 -1151
rect 19978 -1177 20008 -1151
rect 20062 -1177 20092 -1151
rect 20154 -1177 20184 -1151
rect 18317 -1337 18347 -1321
rect 18317 -1367 18372 -1337
rect 17750 -1423 17804 -1407
rect 17562 -1455 17592 -1425
rect 17538 -1471 17592 -1455
rect 17750 -1457 17760 -1423
rect 17794 -1457 17804 -1423
rect 17538 -1505 17548 -1471
rect 17582 -1505 17592 -1471
rect 17538 -1521 17592 -1505
rect 17562 -1555 17592 -1521
rect 17634 -1483 17697 -1467
rect 17750 -1473 17804 -1457
rect 17950 -1410 18026 -1400
rect 17950 -1444 17976 -1410
rect 18010 -1444 18026 -1410
rect 17950 -1454 18026 -1444
rect 18068 -1410 18122 -1394
rect 18222 -1409 18252 -1377
rect 18068 -1444 18078 -1410
rect 18112 -1444 18122 -1410
rect 17634 -1517 17644 -1483
rect 17678 -1517 17697 -1483
rect 17634 -1533 17697 -1517
rect 17667 -1555 17697 -1533
rect 17762 -1543 17792 -1473
rect 17950 -1543 17980 -1454
rect 18068 -1460 18122 -1444
rect 18221 -1425 18280 -1409
rect 18221 -1459 18236 -1425
rect 18270 -1459 18280 -1425
rect 18068 -1498 18098 -1460
rect 18221 -1475 18280 -1459
rect 18342 -1415 18372 -1367
rect 18602 -1245 18632 -1219
rect 18505 -1409 18535 -1377
rect 18602 -1405 18632 -1373
rect 18791 -1377 18821 -1345
rect 18737 -1393 18821 -1377
rect 18500 -1415 18554 -1409
rect 18342 -1425 18554 -1415
rect 18342 -1459 18510 -1425
rect 18544 -1459 18554 -1425
rect 18342 -1469 18554 -1459
rect 18222 -1497 18252 -1475
rect 18034 -1528 18098 -1498
rect 18034 -1543 18064 -1528
rect 18342 -1498 18372 -1469
rect 18505 -1475 18554 -1469
rect 18600 -1421 18682 -1405
rect 18600 -1455 18638 -1421
rect 18672 -1455 18682 -1421
rect 18737 -1427 18747 -1393
rect 18781 -1427 18821 -1393
rect 18737 -1443 18821 -1427
rect 18863 -1393 18893 -1345
rect 18863 -1409 18927 -1393
rect 18863 -1443 18883 -1409
rect 18917 -1443 18927 -1409
rect 18600 -1471 18682 -1455
rect 18505 -1497 18535 -1475
rect 18317 -1528 18372 -1498
rect 18317 -1543 18347 -1528
rect 18600 -1543 18630 -1471
rect 18788 -1499 18818 -1443
rect 18863 -1459 18927 -1443
rect 18969 -1438 18999 -1261
rect 19090 -1293 19120 -1261
rect 19041 -1309 19120 -1293
rect 19195 -1299 19225 -1261
rect 19279 -1293 19309 -1261
rect 19041 -1343 19051 -1309
rect 19085 -1343 19120 -1309
rect 19041 -1359 19120 -1343
rect 19171 -1309 19237 -1299
rect 19171 -1343 19187 -1309
rect 19221 -1343 19237 -1309
rect 19171 -1353 19237 -1343
rect 19279 -1309 19333 -1293
rect 19279 -1343 19289 -1309
rect 19323 -1343 19333 -1309
rect 19279 -1359 19333 -1343
rect 20342 -1183 20372 -1157
rect 20426 -1183 20456 -1157
rect 20614 -1177 20644 -1151
rect 18872 -1499 18902 -1459
rect 18969 -1461 19034 -1438
rect 18969 -1468 18990 -1461
rect 18980 -1495 18990 -1468
rect 19024 -1495 19034 -1461
rect 18980 -1511 19034 -1495
rect 18980 -1543 19010 -1511
rect 19077 -1543 19107 -1359
rect 19279 -1395 19309 -1359
rect 19172 -1425 19309 -1395
rect 19423 -1411 19453 -1345
rect 19560 -1377 19590 -1345
rect 19644 -1377 19674 -1345
rect 19172 -1555 19202 -1425
rect 19376 -1427 19453 -1411
rect 19376 -1461 19386 -1427
rect 19420 -1441 19453 -1427
rect 19504 -1393 19594 -1377
rect 19504 -1427 19514 -1393
rect 19548 -1427 19594 -1393
rect 19420 -1461 19430 -1441
rect 19504 -1443 19594 -1427
rect 19644 -1393 19710 -1377
rect 19644 -1427 19666 -1393
rect 19700 -1427 19710 -1393
rect 19644 -1443 19710 -1427
rect 19244 -1483 19298 -1467
rect 19244 -1517 19254 -1483
rect 19288 -1517 19298 -1483
rect 19376 -1477 19430 -1461
rect 19376 -1499 19406 -1477
rect 19564 -1499 19594 -1443
rect 19648 -1499 19678 -1443
rect 19752 -1445 19782 -1261
rect 19858 -1293 19888 -1261
rect 19824 -1309 19888 -1293
rect 19978 -1299 20008 -1261
rect 19824 -1343 19834 -1309
rect 19868 -1343 19888 -1309
rect 19824 -1359 19888 -1343
rect 19954 -1309 20020 -1299
rect 19954 -1343 19970 -1309
rect 20004 -1343 20020 -1309
rect 19954 -1353 20020 -1343
rect 19752 -1461 19812 -1445
rect 19752 -1481 19768 -1461
rect 19744 -1495 19768 -1481
rect 19802 -1495 19812 -1461
rect 19244 -1533 19298 -1517
rect 19256 -1555 19286 -1533
rect 19744 -1511 19812 -1495
rect 19744 -1543 19774 -1511
rect 19858 -1543 19888 -1359
rect 20062 -1395 20092 -1261
rect 19954 -1425 20092 -1395
rect 20154 -1407 20184 -1261
rect 20342 -1400 20372 -1311
rect 20426 -1326 20456 -1311
rect 20426 -1356 20490 -1326
rect 20460 -1394 20490 -1356
rect 20709 -1193 20739 -1167
rect 20897 -1177 20927 -1151
rect 21183 -1177 21213 -1151
rect 21255 -1177 21285 -1151
rect 21361 -1177 21391 -1151
rect 21482 -1177 21512 -1151
rect 21587 -1177 21617 -1151
rect 21671 -1177 21701 -1151
rect 21815 -1177 21845 -1151
rect 21952 -1177 21982 -1151
rect 22036 -1177 22066 -1151
rect 22144 -1177 22174 -1143
rect 24518 -1146 24584 -1130
rect 22250 -1177 22280 -1151
rect 22370 -1177 22400 -1151
rect 22454 -1177 22484 -1151
rect 22546 -1177 22576 -1151
rect 20709 -1337 20739 -1321
rect 20709 -1367 20764 -1337
rect 20142 -1423 20196 -1407
rect 19954 -1455 19984 -1425
rect 19930 -1471 19984 -1455
rect 20142 -1457 20152 -1423
rect 20186 -1457 20196 -1423
rect 19930 -1505 19940 -1471
rect 19974 -1505 19984 -1471
rect 19930 -1521 19984 -1505
rect 19954 -1555 19984 -1521
rect 20026 -1483 20089 -1467
rect 20142 -1473 20196 -1457
rect 20342 -1410 20418 -1400
rect 20342 -1444 20368 -1410
rect 20402 -1444 20418 -1410
rect 20342 -1454 20418 -1444
rect 20460 -1410 20514 -1394
rect 20614 -1409 20644 -1377
rect 20460 -1444 20470 -1410
rect 20504 -1444 20514 -1410
rect 20026 -1517 20036 -1483
rect 20070 -1517 20089 -1483
rect 20026 -1533 20089 -1517
rect 20059 -1555 20089 -1533
rect 20154 -1543 20184 -1473
rect 20342 -1543 20372 -1454
rect 20460 -1460 20514 -1444
rect 20613 -1425 20672 -1409
rect 20613 -1459 20628 -1425
rect 20662 -1459 20672 -1425
rect 20460 -1498 20490 -1460
rect 20613 -1475 20672 -1459
rect 20734 -1415 20764 -1367
rect 20994 -1245 21024 -1219
rect 20897 -1409 20927 -1377
rect 20994 -1405 21024 -1373
rect 21183 -1377 21213 -1345
rect 21129 -1393 21213 -1377
rect 20892 -1415 20946 -1409
rect 20734 -1425 20946 -1415
rect 20734 -1459 20902 -1425
rect 20936 -1459 20946 -1425
rect 20734 -1469 20946 -1459
rect 20614 -1497 20644 -1475
rect 20426 -1528 20490 -1498
rect 20426 -1543 20456 -1528
rect 20734 -1498 20764 -1469
rect 20897 -1475 20946 -1469
rect 20992 -1421 21074 -1405
rect 20992 -1455 21030 -1421
rect 21064 -1455 21074 -1421
rect 21129 -1427 21139 -1393
rect 21173 -1427 21213 -1393
rect 21129 -1443 21213 -1427
rect 21255 -1393 21285 -1345
rect 21255 -1409 21319 -1393
rect 21255 -1443 21275 -1409
rect 21309 -1443 21319 -1409
rect 20992 -1471 21074 -1455
rect 20897 -1497 20927 -1475
rect 20709 -1528 20764 -1498
rect 20709 -1543 20739 -1528
rect 20992 -1543 21022 -1471
rect 21180 -1499 21210 -1443
rect 21255 -1459 21319 -1443
rect 21361 -1438 21391 -1261
rect 21482 -1293 21512 -1261
rect 21433 -1309 21512 -1293
rect 21587 -1299 21617 -1261
rect 21671 -1293 21701 -1261
rect 21433 -1343 21443 -1309
rect 21477 -1343 21512 -1309
rect 21433 -1359 21512 -1343
rect 21563 -1309 21629 -1299
rect 21563 -1343 21579 -1309
rect 21613 -1343 21629 -1309
rect 21563 -1353 21629 -1343
rect 21671 -1309 21725 -1293
rect 21671 -1343 21681 -1309
rect 21715 -1343 21725 -1309
rect 21671 -1359 21725 -1343
rect 22734 -1183 22764 -1157
rect 22818 -1183 22848 -1157
rect 23006 -1177 23036 -1151
rect 21264 -1499 21294 -1459
rect 21361 -1461 21426 -1438
rect 21361 -1468 21382 -1461
rect 21372 -1495 21382 -1468
rect 21416 -1495 21426 -1461
rect 21372 -1511 21426 -1495
rect 21372 -1543 21402 -1511
rect 21469 -1543 21499 -1359
rect 21671 -1395 21701 -1359
rect 21564 -1425 21701 -1395
rect 21815 -1411 21845 -1345
rect 21952 -1377 21982 -1345
rect 22036 -1377 22066 -1345
rect 21564 -1555 21594 -1425
rect 21768 -1427 21845 -1411
rect 21768 -1461 21778 -1427
rect 21812 -1441 21845 -1427
rect 21896 -1393 21986 -1377
rect 21896 -1427 21906 -1393
rect 21940 -1427 21986 -1393
rect 21812 -1461 21822 -1441
rect 21896 -1443 21986 -1427
rect 22036 -1393 22102 -1377
rect 22036 -1427 22058 -1393
rect 22092 -1427 22102 -1393
rect 22036 -1443 22102 -1427
rect 21636 -1483 21690 -1467
rect 21636 -1517 21646 -1483
rect 21680 -1517 21690 -1483
rect 21768 -1477 21822 -1461
rect 21768 -1499 21798 -1477
rect 21956 -1499 21986 -1443
rect 22040 -1499 22070 -1443
rect 22144 -1445 22174 -1261
rect 22250 -1293 22280 -1261
rect 22216 -1309 22280 -1293
rect 22370 -1299 22400 -1261
rect 22216 -1343 22226 -1309
rect 22260 -1343 22280 -1309
rect 22216 -1359 22280 -1343
rect 22346 -1309 22412 -1299
rect 22346 -1343 22362 -1309
rect 22396 -1343 22412 -1309
rect 22346 -1353 22412 -1343
rect 22144 -1461 22204 -1445
rect 22144 -1481 22160 -1461
rect 22136 -1495 22160 -1481
rect 22194 -1495 22204 -1461
rect 21636 -1533 21690 -1517
rect 21648 -1555 21678 -1533
rect 22136 -1511 22204 -1495
rect 22136 -1543 22166 -1511
rect 22250 -1543 22280 -1359
rect 22454 -1395 22484 -1261
rect 22346 -1425 22484 -1395
rect 22546 -1407 22576 -1261
rect 22734 -1400 22764 -1311
rect 22818 -1326 22848 -1311
rect 22818 -1356 22882 -1326
rect 22852 -1394 22882 -1356
rect 23101 -1193 23131 -1167
rect 23289 -1177 23319 -1151
rect 23575 -1177 23605 -1151
rect 23647 -1177 23677 -1151
rect 23753 -1177 23783 -1151
rect 23874 -1177 23904 -1151
rect 23979 -1177 24009 -1151
rect 24063 -1177 24093 -1151
rect 24207 -1177 24237 -1151
rect 24344 -1177 24374 -1151
rect 24428 -1177 24458 -1151
rect 24536 -1177 24566 -1146
rect 24642 -1177 24672 -1151
rect 24762 -1177 24792 -1151
rect 24846 -1177 24876 -1151
rect 24938 -1177 24968 -1151
rect 23101 -1337 23131 -1321
rect 23101 -1367 23156 -1337
rect 22534 -1423 22588 -1407
rect 22346 -1455 22376 -1425
rect 22322 -1471 22376 -1455
rect 22534 -1457 22544 -1423
rect 22578 -1457 22588 -1423
rect 22322 -1505 22332 -1471
rect 22366 -1505 22376 -1471
rect 22322 -1521 22376 -1505
rect 22346 -1555 22376 -1521
rect 22418 -1483 22481 -1467
rect 22534 -1473 22588 -1457
rect 22734 -1410 22810 -1400
rect 22734 -1444 22760 -1410
rect 22794 -1444 22810 -1410
rect 22734 -1454 22810 -1444
rect 22852 -1410 22906 -1394
rect 23006 -1409 23036 -1377
rect 22852 -1444 22862 -1410
rect 22896 -1444 22906 -1410
rect 22418 -1517 22428 -1483
rect 22462 -1517 22481 -1483
rect 22418 -1533 22481 -1517
rect 22451 -1555 22481 -1533
rect 22546 -1543 22576 -1473
rect 22734 -1543 22764 -1454
rect 22852 -1460 22906 -1444
rect 23005 -1425 23064 -1409
rect 23005 -1459 23020 -1425
rect 23054 -1459 23064 -1425
rect 22852 -1498 22882 -1460
rect 23005 -1475 23064 -1459
rect 23126 -1415 23156 -1367
rect 23386 -1245 23416 -1219
rect 23289 -1409 23319 -1377
rect 23386 -1405 23416 -1373
rect 23575 -1377 23605 -1345
rect 23521 -1393 23605 -1377
rect 23284 -1415 23338 -1409
rect 23126 -1425 23338 -1415
rect 23126 -1459 23294 -1425
rect 23328 -1459 23338 -1425
rect 23126 -1469 23338 -1459
rect 23006 -1497 23036 -1475
rect 22818 -1528 22882 -1498
rect 22818 -1543 22848 -1528
rect 23126 -1498 23156 -1469
rect 23289 -1475 23338 -1469
rect 23384 -1421 23466 -1405
rect 23384 -1455 23422 -1421
rect 23456 -1455 23466 -1421
rect 23521 -1427 23531 -1393
rect 23565 -1427 23605 -1393
rect 23521 -1443 23605 -1427
rect 23647 -1393 23677 -1345
rect 23647 -1409 23711 -1393
rect 23647 -1443 23667 -1409
rect 23701 -1443 23711 -1409
rect 23384 -1471 23466 -1455
rect 23289 -1497 23319 -1475
rect 23101 -1528 23156 -1498
rect 23101 -1543 23131 -1528
rect 23384 -1543 23414 -1471
rect 23572 -1499 23602 -1443
rect 23647 -1459 23711 -1443
rect 23753 -1438 23783 -1261
rect 23874 -1293 23904 -1261
rect 23825 -1309 23904 -1293
rect 23979 -1299 24009 -1261
rect 24063 -1293 24093 -1261
rect 23825 -1343 23835 -1309
rect 23869 -1343 23904 -1309
rect 23825 -1359 23904 -1343
rect 23955 -1309 24021 -1299
rect 23955 -1343 23971 -1309
rect 24005 -1343 24021 -1309
rect 23955 -1353 24021 -1343
rect 24063 -1309 24117 -1293
rect 24063 -1343 24073 -1309
rect 24107 -1343 24117 -1309
rect 24063 -1359 24117 -1343
rect 25126 -1183 25156 -1157
rect 25210 -1183 25240 -1157
rect 23656 -1499 23686 -1459
rect 23753 -1461 23818 -1438
rect 23753 -1468 23774 -1461
rect 23764 -1495 23774 -1468
rect 23808 -1495 23818 -1461
rect 23764 -1511 23818 -1495
rect 23764 -1543 23794 -1511
rect 23861 -1543 23891 -1359
rect 24063 -1395 24093 -1359
rect 23956 -1425 24093 -1395
rect 24207 -1411 24237 -1345
rect 24344 -1377 24374 -1345
rect 24428 -1377 24458 -1345
rect 23956 -1555 23986 -1425
rect 24160 -1427 24237 -1411
rect 24160 -1461 24170 -1427
rect 24204 -1441 24237 -1427
rect 24288 -1393 24378 -1377
rect 24288 -1427 24298 -1393
rect 24332 -1427 24378 -1393
rect 24204 -1461 24214 -1441
rect 24288 -1443 24378 -1427
rect 24428 -1393 24494 -1377
rect 24428 -1427 24450 -1393
rect 24484 -1427 24494 -1393
rect 24428 -1443 24494 -1427
rect 24028 -1483 24082 -1467
rect 24028 -1517 24038 -1483
rect 24072 -1517 24082 -1483
rect 24160 -1477 24214 -1461
rect 24160 -1499 24190 -1477
rect 24348 -1499 24378 -1443
rect 24432 -1499 24462 -1443
rect 24536 -1445 24566 -1261
rect 24642 -1293 24672 -1261
rect 24608 -1309 24672 -1293
rect 24762 -1299 24792 -1261
rect 24608 -1343 24618 -1309
rect 24652 -1343 24672 -1309
rect 24608 -1359 24672 -1343
rect 24738 -1309 24804 -1299
rect 24738 -1343 24754 -1309
rect 24788 -1343 24804 -1309
rect 24738 -1353 24804 -1343
rect 24536 -1461 24596 -1445
rect 24536 -1481 24552 -1461
rect 24528 -1495 24552 -1481
rect 24586 -1495 24596 -1461
rect 24028 -1533 24082 -1517
rect 24040 -1555 24070 -1533
rect 24528 -1511 24596 -1495
rect 24528 -1543 24558 -1511
rect 24642 -1543 24672 -1359
rect 24846 -1395 24876 -1261
rect 24738 -1425 24876 -1395
rect 24938 -1407 24968 -1261
rect 25126 -1400 25156 -1311
rect 25210 -1326 25240 -1311
rect 25210 -1356 25274 -1326
rect 25244 -1394 25274 -1356
rect 24926 -1423 24980 -1407
rect 24738 -1455 24768 -1425
rect 24714 -1471 24768 -1455
rect 24926 -1457 24936 -1423
rect 24970 -1457 24980 -1423
rect 24714 -1505 24724 -1471
rect 24758 -1505 24768 -1471
rect 24714 -1521 24768 -1505
rect 24738 -1555 24768 -1521
rect 24810 -1483 24873 -1467
rect 24926 -1473 24980 -1457
rect 25126 -1410 25202 -1400
rect 25126 -1444 25152 -1410
rect 25186 -1444 25202 -1410
rect 25126 -1454 25202 -1444
rect 25244 -1410 25298 -1394
rect 25244 -1444 25254 -1410
rect 25288 -1444 25298 -1410
rect 24810 -1517 24820 -1483
rect 24854 -1517 24873 -1483
rect 24810 -1533 24873 -1517
rect 24843 -1555 24873 -1533
rect 24938 -1543 24968 -1473
rect 25126 -1543 25156 -1454
rect 25244 -1460 25298 -1444
rect 25244 -1498 25274 -1460
rect 25210 -1528 25274 -1498
rect 25210 -1543 25240 -1528
rect 8654 -1653 8684 -1627
rect 8749 -1653 8779 -1627
rect 8937 -1653 8967 -1627
rect 9032 -1653 9062 -1627
rect 9220 -1653 9250 -1627
rect 9304 -1653 9334 -1627
rect 9412 -1653 9442 -1627
rect 9509 -1653 9539 -1627
rect 9604 -1653 9634 -1627
rect 9688 -1653 9718 -1627
rect 9808 -1653 9838 -1627
rect 9996 -1653 10026 -1627
rect 10080 -1653 10110 -1627
rect 10176 -1653 10206 -1627
rect 10290 -1653 10320 -1627
rect 10386 -1653 10416 -1627
rect 10491 -1653 10521 -1627
rect 10586 -1653 10616 -1627
rect 10774 -1653 10804 -1627
rect 10858 -1653 10888 -1627
rect 11046 -1653 11076 -1627
rect 11141 -1653 11171 -1627
rect 11329 -1653 11359 -1627
rect 11424 -1653 11454 -1627
rect 11612 -1653 11642 -1627
rect 11696 -1653 11726 -1627
rect 11804 -1653 11834 -1627
rect 11901 -1653 11931 -1627
rect 11996 -1653 12026 -1627
rect 12080 -1653 12110 -1627
rect 12200 -1653 12230 -1627
rect 12388 -1653 12418 -1627
rect 12472 -1653 12502 -1627
rect 12568 -1653 12598 -1627
rect 12682 -1653 12712 -1627
rect 12778 -1653 12808 -1627
rect 12883 -1653 12913 -1627
rect 12978 -1653 13008 -1627
rect 13166 -1653 13196 -1627
rect 13250 -1653 13280 -1627
rect 13438 -1653 13468 -1627
rect 13533 -1653 13563 -1627
rect 13721 -1653 13751 -1627
rect 13816 -1653 13846 -1627
rect 14004 -1653 14034 -1627
rect 14088 -1653 14118 -1627
rect 14196 -1653 14226 -1627
rect 14293 -1653 14323 -1627
rect 14388 -1653 14418 -1627
rect 14472 -1653 14502 -1627
rect 14592 -1653 14622 -1627
rect 14780 -1653 14810 -1627
rect 14864 -1653 14894 -1627
rect 14960 -1653 14990 -1627
rect 15074 -1653 15104 -1627
rect 15170 -1653 15200 -1627
rect 15275 -1653 15305 -1627
rect 15370 -1653 15400 -1627
rect 15558 -1653 15588 -1627
rect 15642 -1653 15672 -1627
rect 15830 -1653 15860 -1627
rect 15925 -1653 15955 -1627
rect 16113 -1653 16143 -1627
rect 16208 -1653 16238 -1627
rect 16396 -1653 16426 -1627
rect 16480 -1653 16510 -1627
rect 16588 -1653 16618 -1627
rect 16685 -1653 16715 -1627
rect 16780 -1653 16810 -1627
rect 16864 -1653 16894 -1627
rect 16984 -1653 17014 -1627
rect 17172 -1653 17202 -1627
rect 17256 -1653 17286 -1627
rect 17352 -1653 17382 -1627
rect 17466 -1653 17496 -1627
rect 17562 -1653 17592 -1627
rect 17667 -1653 17697 -1627
rect 17762 -1653 17792 -1627
rect 17950 -1653 17980 -1627
rect 18034 -1653 18064 -1627
rect 18222 -1653 18252 -1627
rect 18317 -1653 18347 -1627
rect 18505 -1653 18535 -1627
rect 18600 -1653 18630 -1627
rect 18788 -1653 18818 -1627
rect 18872 -1653 18902 -1627
rect 18980 -1653 19010 -1627
rect 19077 -1653 19107 -1627
rect 19172 -1653 19202 -1627
rect 19256 -1653 19286 -1627
rect 19376 -1653 19406 -1627
rect 19564 -1653 19594 -1627
rect 19648 -1653 19678 -1627
rect 19744 -1653 19774 -1627
rect 19858 -1653 19888 -1627
rect 19954 -1653 19984 -1627
rect 20059 -1653 20089 -1627
rect 20154 -1653 20184 -1627
rect 20342 -1653 20372 -1627
rect 20426 -1653 20456 -1627
rect 20614 -1653 20644 -1627
rect 20709 -1653 20739 -1627
rect 20897 -1653 20927 -1627
rect 20992 -1653 21022 -1627
rect 21180 -1653 21210 -1627
rect 21264 -1653 21294 -1627
rect 21372 -1653 21402 -1627
rect 21469 -1653 21499 -1627
rect 21564 -1653 21594 -1627
rect 21648 -1653 21678 -1627
rect 21768 -1653 21798 -1627
rect 21956 -1653 21986 -1627
rect 22040 -1653 22070 -1627
rect 22136 -1653 22166 -1627
rect 22250 -1653 22280 -1627
rect 22346 -1653 22376 -1627
rect 22451 -1653 22481 -1627
rect 22546 -1653 22576 -1627
rect 22734 -1653 22764 -1627
rect 22818 -1653 22848 -1627
rect 23006 -1653 23036 -1627
rect 23101 -1653 23131 -1627
rect 23289 -1653 23319 -1627
rect 23384 -1653 23414 -1627
rect 23572 -1653 23602 -1627
rect 23656 -1653 23686 -1627
rect 23764 -1653 23794 -1627
rect 23861 -1653 23891 -1627
rect 23956 -1653 23986 -1627
rect 24040 -1653 24070 -1627
rect 24160 -1653 24190 -1627
rect 24348 -1653 24378 -1627
rect 24432 -1653 24462 -1627
rect 24528 -1653 24558 -1627
rect 24642 -1653 24672 -1627
rect 24738 -1653 24768 -1627
rect 24843 -1653 24873 -1627
rect 24938 -1653 24968 -1627
rect 25126 -1653 25156 -1627
rect 25210 -1653 25240 -1627
<< polycont >>
rect 13354 12664 13388 12698
rect 13860 12738 13894 12772
rect 13620 12664 13654 12698
rect 20063 12664 20097 12698
rect 20569 12738 20603 12772
rect 20329 12664 20363 12698
rect 14502 12495 14536 12529
rect 15234 12498 15268 12532
rect 15360 12498 15394 12532
rect 16446 12498 16480 12532
rect 16572 12498 16606 12532
rect 17658 12498 17692 12532
rect 17784 12498 17818 12532
rect 18870 12498 18904 12532
rect 18996 12498 19030 12532
rect 21211 12495 21245 12529
rect 21943 12498 21977 12532
rect 22069 12498 22103 12532
rect 23155 12498 23189 12532
rect 23281 12498 23315 12532
rect 24367 12498 24401 12532
rect 24493 12498 24527 12532
rect 25579 12498 25613 12532
rect 25705 12498 25739 12532
rect 2466 12189 2500 12223
rect 2972 12263 3006 12297
rect 2732 12189 2766 12223
rect 11348 12258 11382 12292
rect 10914 12185 10948 12219
rect 11016 12185 11050 12219
rect 11444 12246 11478 12280
rect 11232 12198 11266 12232
rect 3614 12020 3648 12054
rect 4346 12023 4380 12057
rect 4472 12023 4506 12057
rect 5558 12023 5592 12057
rect 5684 12023 5718 12057
rect 6770 12023 6804 12057
rect 6896 12023 6930 12057
rect 7982 12023 8016 12057
rect 8108 12023 8142 12057
rect 11616 12236 11650 12270
rect 11414 12084 11448 12118
rect 11550 12084 11584 12118
rect 12130 12258 12164 12292
rect 11718 12168 11752 12202
rect 11870 12168 11904 12202
rect 11998 12202 12032 12236
rect 12393 12236 12427 12270
rect 12095 12084 12129 12118
rect 12197 12084 12231 12118
rect 12333 12084 12367 12118
rect 12501 12184 12535 12218
rect 12639 12168 12673 12202
rect 12770 12196 12804 12230
rect 19530 12291 19564 12325
rect 19737 12289 19771 12323
rect 26239 12291 26273 12325
rect 12870 12200 12904 12234
rect 13146 12200 13180 12234
rect 26446 12289 26480 12323
rect 13871 12104 13905 12138
rect 14855 12094 14889 12128
rect 15587 12094 15621 12128
rect 15709 12094 15743 12128
rect 16799 12094 16833 12128
rect 16921 12094 16955 12128
rect 18137 12094 18171 12128
rect 18259 12094 18293 12128
rect 18993 12094 19027 12128
rect 20580 12104 20614 12138
rect 21564 12094 21598 12128
rect 22296 12094 22330 12128
rect 22418 12094 22452 12128
rect 23508 12094 23542 12128
rect 23630 12094 23664 12128
rect 24846 12094 24880 12128
rect 24968 12094 25002 12128
rect 25702 12094 25736 12128
rect 8642 11816 8676 11850
rect 8849 11814 8883 11848
rect 9141 11812 9175 11846
rect 2983 11629 3017 11663
rect 3967 11619 4001 11653
rect 4699 11619 4733 11653
rect 4821 11619 4855 11653
rect 5911 11619 5945 11653
rect 6033 11619 6067 11653
rect 7249 11619 7283 11653
rect 7371 11619 7405 11653
rect 8105 11619 8139 11653
rect 10962 11480 10996 11514
rect 11238 11480 11272 11514
rect 2983 8983 3017 9017
rect 3967 8993 4001 9027
rect 4699 8993 4733 9027
rect 4821 8993 4855 9027
rect 5911 8993 5945 9027
rect 6033 8993 6067 9027
rect 7249 8993 7283 9027
rect 7371 8993 7405 9027
rect 8105 8993 8139 9027
rect 8642 8796 8676 8830
rect 8849 8798 8883 8832
rect 9141 8802 9175 8836
rect 9411 8802 9445 8836
rect 9687 8802 9721 8836
rect 3614 8592 3648 8626
rect 4346 8589 4380 8623
rect 4472 8589 4506 8623
rect 5558 8589 5592 8623
rect 5684 8589 5718 8623
rect 6770 8589 6804 8623
rect 6896 8589 6930 8623
rect 7982 8589 8016 8623
rect 8108 8589 8142 8623
rect 9787 8798 9821 8832
rect 9918 8770 9952 8804
rect 10164 8838 10198 8872
rect 10056 8786 10090 8820
rect 10427 8860 10461 8894
rect 10559 8804 10593 8838
rect 10941 8838 10975 8872
rect 10224 8686 10258 8720
rect 10360 8686 10394 8720
rect 10687 8770 10721 8804
rect 10839 8770 10873 8804
rect 10462 8686 10496 8720
rect 11113 8848 11147 8882
rect 11209 8860 11243 8894
rect 11325 8800 11359 8834
rect 11541 8787 11575 8821
rect 11007 8686 11041 8720
rect 11143 8686 11177 8720
rect 14152 8981 14186 9015
rect 14886 8981 14920 9015
rect 15008 8981 15042 9015
rect 16224 8981 16258 9015
rect 16346 8981 16380 9015
rect 17436 8981 17470 9015
rect 17558 8981 17592 9015
rect 18290 8981 18324 9015
rect 19274 8971 19308 9005
rect 11643 8787 11677 8821
rect 12073 8787 12107 8821
rect 12277 8788 12311 8822
rect 12478 8787 12512 8821
rect 12687 8789 12721 8823
rect 2466 8423 2500 8457
rect 11332 8473 11366 8507
rect 20861 8981 20895 9015
rect 21595 8981 21629 9015
rect 21717 8981 21751 9015
rect 22933 8981 22967 9015
rect 23055 8981 23089 9015
rect 24145 8981 24179 9015
rect 24267 8981 24301 9015
rect 24999 8981 25033 9015
rect 25983 8971 26017 9005
rect 12855 8789 12889 8823
rect 13087 8789 13121 8823
rect 13408 8786 13442 8820
rect 13615 8784 13649 8818
rect 20117 8786 20151 8820
rect 20324 8784 20358 8818
rect 14149 8577 14183 8611
rect 14275 8577 14309 8611
rect 15361 8577 15395 8611
rect 15487 8577 15521 8611
rect 16573 8577 16607 8611
rect 16699 8577 16733 8611
rect 17785 8577 17819 8611
rect 17911 8577 17945 8611
rect 18643 8580 18677 8614
rect 20858 8577 20892 8611
rect 20984 8577 21018 8611
rect 22070 8577 22104 8611
rect 22196 8577 22230 8611
rect 23282 8577 23316 8611
rect 23408 8577 23442 8611
rect 24494 8577 24528 8611
rect 24620 8577 24654 8611
rect 25352 8580 25386 8614
rect 2732 8423 2766 8457
rect 19525 8411 19559 8445
rect 2972 8349 3006 8383
rect 10140 8003 10174 8037
rect 10236 8003 10270 8037
rect 10545 8080 10579 8114
rect 10377 7967 10411 8001
rect 10713 8080 10747 8114
rect 10473 7967 10507 8001
rect 10635 7967 10669 8001
rect 10967 8003 11001 8037
rect 11063 8003 11097 8037
rect 11372 8080 11406 8114
rect 11204 7967 11238 8001
rect 11540 8080 11574 8114
rect 11300 7967 11334 8001
rect 11462 7967 11496 8001
rect 19285 8337 19319 8371
rect 19791 8411 19825 8445
rect 26234 8411 26268 8445
rect 12746 8190 12780 8224
rect 25994 8337 26028 8371
rect 26500 8411 26534 8445
rect 12073 8003 12107 8037
rect 12277 8002 12311 8036
rect 12746 7503 12780 7537
rect 11535 6748 11569 6782
rect 11653 6761 11687 6795
rect 11818 6748 11852 6782
rect 11952 6748 11986 6782
rect 13406 6864 13440 6898
rect 13304 6798 13338 6832
rect 13112 6748 13146 6782
rect 13208 6748 13242 6782
rect 13340 6690 13374 6724
rect 13574 6762 13608 6796
rect 13901 6761 13935 6795
rect 14217 6864 14251 6898
rect 14319 6806 14353 6840
rect 14003 6702 14037 6736
rect 14099 6702 14133 6736
rect 14282 6690 14316 6724
rect 14396 6702 14430 6736
rect 14532 6748 14566 6782
rect 24079 6367 24113 6401
rect 24585 6441 24619 6475
rect 24345 6367 24379 6401
rect 13397 6202 13431 6236
rect 14640 6205 14674 6239
rect 17032 6207 17066 6241
rect 19424 6207 19458 6241
rect 21816 6208 21850 6242
rect 11529 5890 11563 5924
rect 12029 5991 12063 6025
rect 12165 5991 12199 6025
rect 11631 5890 11665 5924
rect 11847 5877 11881 5911
rect 11963 5817 11997 5851
rect 12059 5829 12093 5863
rect 12710 5991 12744 6025
rect 12333 5907 12367 5941
rect 12485 5907 12519 5941
rect 12812 5991 12846 6025
rect 12948 5991 12982 6025
rect 12231 5839 12265 5873
rect 12613 5873 12647 5907
rect 12745 5817 12779 5851
rect 13116 5891 13150 5925
rect 13008 5839 13042 5873
rect 13254 5907 13288 5941
rect 13385 5879 13419 5913
rect 13485 5875 13519 5909
rect 13761 5875 13795 5909
rect 13921 5890 13955 5924
rect 14421 5991 14455 6025
rect 14557 5991 14591 6025
rect 14023 5890 14057 5924
rect 14239 5877 14273 5911
rect 14355 5817 14389 5851
rect 14451 5829 14485 5863
rect 15102 5991 15136 6025
rect 14725 5907 14759 5941
rect 14877 5907 14911 5941
rect 15204 5991 15238 6025
rect 15340 5991 15374 6025
rect 14623 5839 14657 5873
rect 15005 5873 15039 5907
rect 15137 5817 15171 5851
rect 15508 5891 15542 5925
rect 15400 5839 15434 5873
rect 15646 5907 15680 5941
rect 15777 5879 15811 5913
rect 15877 5875 15911 5909
rect 16153 5875 16187 5909
rect 16313 5890 16347 5924
rect 16813 5991 16847 6025
rect 16949 5991 16983 6025
rect 16415 5890 16449 5924
rect 16631 5877 16665 5911
rect 16747 5817 16781 5851
rect 16843 5829 16877 5863
rect 17494 5991 17528 6025
rect 17117 5907 17151 5941
rect 17269 5907 17303 5941
rect 17596 5991 17630 6025
rect 17732 5991 17766 6025
rect 17015 5839 17049 5873
rect 17397 5873 17431 5907
rect 17529 5817 17563 5851
rect 17900 5891 17934 5925
rect 17792 5839 17826 5873
rect 18038 5907 18072 5941
rect 18169 5879 18203 5913
rect 18269 5875 18303 5909
rect 18545 5875 18579 5909
rect 18705 5890 18739 5924
rect 19205 5991 19239 6025
rect 19341 5991 19375 6025
rect 18807 5890 18841 5924
rect 19023 5877 19057 5911
rect 19139 5817 19173 5851
rect 19235 5829 19269 5863
rect 19886 5991 19920 6025
rect 19509 5907 19543 5941
rect 19661 5907 19695 5941
rect 19988 5991 20022 6025
rect 20124 5991 20158 6025
rect 19407 5839 19441 5873
rect 19789 5873 19823 5907
rect 19921 5817 19955 5851
rect 20292 5891 20326 5925
rect 20184 5839 20218 5873
rect 20430 5907 20464 5941
rect 20561 5879 20595 5913
rect 20661 5875 20695 5909
rect 20937 5875 20971 5909
rect 21097 5890 21131 5924
rect 21597 5991 21631 6025
rect 21733 5991 21767 6025
rect 21199 5890 21233 5924
rect 21415 5877 21449 5911
rect 21531 5817 21565 5851
rect 21627 5829 21661 5863
rect 22278 5991 22312 6025
rect 21901 5907 21935 5941
rect 22053 5907 22087 5941
rect 22380 5991 22414 6025
rect 22516 5991 22550 6025
rect 21799 5839 21833 5873
rect 22181 5873 22215 5907
rect 22313 5817 22347 5851
rect 22684 5891 22718 5925
rect 22576 5839 22610 5873
rect 22822 5907 22856 5941
rect 25227 6198 25261 6232
rect 25959 6201 25993 6235
rect 26085 6201 26119 6235
rect 27171 6201 27205 6235
rect 27297 6201 27331 6235
rect 28383 6201 28417 6235
rect 28509 6201 28543 6235
rect 29595 6201 29629 6235
rect 29721 6201 29755 6235
rect 22953 5879 22987 5913
rect 30255 5994 30289 6028
rect 30462 5992 30496 6026
rect 30716 5990 30750 6024
rect 30840 5990 30874 6024
rect 23053 5875 23087 5909
rect 23329 5875 23363 5909
rect 24596 5807 24630 5841
rect 25580 5797 25614 5831
rect 26312 5797 26346 5831
rect 26434 5797 26468 5831
rect 27524 5797 27558 5831
rect 27646 5797 27680 5831
rect 28862 5797 28896 5831
rect 28984 5797 29018 5831
rect 29718 5797 29752 5831
rect 14711 5519 14745 5553
rect 17103 5519 17137 5553
rect 19495 5519 19529 5553
rect 21887 5519 21921 5553
rect 11094 5186 11128 5220
rect 11212 5199 11246 5233
rect 11377 5186 11411 5220
rect 11511 5186 11545 5220
rect 11968 5186 12002 5220
rect 12036 5186 12070 5220
rect 12104 5186 12138 5220
rect 12172 5186 12206 5220
rect 12240 5186 12274 5220
rect 12308 5186 12342 5220
rect 12468 5186 12502 5220
rect 12536 5186 12570 5220
rect 12604 5186 12638 5220
rect 12672 5186 12706 5220
rect 12740 5186 12774 5220
rect 12808 5186 12842 5220
rect 12876 5186 12910 5220
rect 12944 5186 12978 5220
rect 13012 5186 13046 5220
rect 13080 5186 13114 5220
rect 13148 5186 13182 5220
rect 13216 5186 13250 5220
rect 13284 5186 13318 5220
rect 13352 5186 13386 5220
rect 13420 5186 13454 5220
rect 13488 5186 13522 5220
rect 13556 5186 13590 5220
rect 13624 5186 13658 5220
rect 13692 5186 13726 5220
rect 13983 5186 14017 5220
rect 14259 5186 14293 5220
rect 14359 5190 14393 5224
rect 14490 5218 14524 5252
rect 14628 5202 14662 5236
rect 14796 5302 14830 5336
rect 14932 5302 14966 5336
rect 15034 5302 15068 5336
rect 14736 5150 14770 5184
rect 15131 5184 15165 5218
rect 15259 5218 15293 5252
rect 15411 5218 15445 5252
rect 14999 5128 15033 5162
rect 15579 5302 15613 5336
rect 15715 5302 15749 5336
rect 15513 5150 15547 5184
rect 15897 5188 15931 5222
rect 15685 5140 15719 5174
rect 16113 5201 16147 5235
rect 16215 5201 16249 5235
rect 15781 5128 15815 5162
rect 16375 5186 16409 5220
rect 16651 5186 16685 5220
rect 16751 5190 16785 5224
rect 16882 5218 16916 5252
rect 17020 5202 17054 5236
rect 17188 5302 17222 5336
rect 17324 5302 17358 5336
rect 17426 5302 17460 5336
rect 17128 5150 17162 5184
rect 17523 5184 17557 5218
rect 17651 5218 17685 5252
rect 17803 5218 17837 5252
rect 17391 5128 17425 5162
rect 17971 5302 18005 5336
rect 18107 5302 18141 5336
rect 17905 5150 17939 5184
rect 18289 5188 18323 5222
rect 18077 5140 18111 5174
rect 18505 5201 18539 5235
rect 18607 5201 18641 5235
rect 18173 5128 18207 5162
rect 18767 5186 18801 5220
rect 19043 5186 19077 5220
rect 19143 5190 19177 5224
rect 19274 5218 19308 5252
rect 19412 5202 19446 5236
rect 19580 5302 19614 5336
rect 19716 5302 19750 5336
rect 19818 5302 19852 5336
rect 19520 5150 19554 5184
rect 19915 5184 19949 5218
rect 20043 5218 20077 5252
rect 20195 5218 20229 5252
rect 19783 5128 19817 5162
rect 20363 5302 20397 5336
rect 20499 5302 20533 5336
rect 20297 5150 20331 5184
rect 20681 5188 20715 5222
rect 20469 5140 20503 5174
rect 20897 5201 20931 5235
rect 20999 5201 21033 5235
rect 20565 5128 20599 5162
rect 21159 5186 21193 5220
rect 21435 5186 21469 5220
rect 21535 5190 21569 5224
rect 21666 5218 21700 5252
rect 21804 5202 21838 5236
rect 21972 5302 22006 5336
rect 22108 5302 22142 5336
rect 22210 5302 22244 5336
rect 21912 5150 21946 5184
rect 22307 5184 22341 5218
rect 22435 5218 22469 5252
rect 22587 5218 22621 5252
rect 22175 5128 22209 5162
rect 22755 5302 22789 5336
rect 22891 5302 22925 5336
rect 22689 5150 22723 5184
rect 23073 5188 23107 5222
rect 22861 5140 22895 5174
rect 23289 5201 23323 5235
rect 23391 5201 23425 5235
rect 22957 5128 22991 5162
rect 11126 4312 11160 4346
rect 11244 4325 11278 4359
rect 11409 4312 11443 4346
rect 11543 4312 11577 4346
rect 13711 4313 13745 4347
rect 13920 4328 13954 4362
rect 14420 4429 14454 4463
rect 14556 4429 14590 4463
rect 14022 4328 14056 4362
rect 14238 4315 14272 4349
rect 14354 4255 14388 4289
rect 14450 4267 14484 4301
rect 15101 4429 15135 4463
rect 14724 4345 14758 4379
rect 14876 4345 14910 4379
rect 15203 4429 15237 4463
rect 15339 4429 15373 4463
rect 14622 4277 14656 4311
rect 15004 4311 15038 4345
rect 15136 4255 15170 4289
rect 15507 4329 15541 4363
rect 15399 4277 15433 4311
rect 15645 4345 15679 4379
rect 15776 4317 15810 4351
rect 15876 4313 15910 4347
rect 16152 4313 16186 4347
rect 16312 4328 16346 4362
rect 16812 4429 16846 4463
rect 16948 4429 16982 4463
rect 16414 4328 16448 4362
rect 16630 4315 16664 4349
rect 16746 4255 16780 4289
rect 16842 4267 16876 4301
rect 17493 4429 17527 4463
rect 17116 4345 17150 4379
rect 17268 4345 17302 4379
rect 17595 4429 17629 4463
rect 17731 4429 17765 4463
rect 17014 4277 17048 4311
rect 17396 4311 17430 4345
rect 17528 4255 17562 4289
rect 17899 4329 17933 4363
rect 17791 4277 17825 4311
rect 18037 4345 18071 4379
rect 18168 4317 18202 4351
rect 18268 4313 18302 4347
rect 18544 4313 18578 4347
rect 18704 4328 18738 4362
rect 19204 4429 19238 4463
rect 19340 4429 19374 4463
rect 18806 4328 18840 4362
rect 19022 4315 19056 4349
rect 19138 4255 19172 4289
rect 19234 4267 19268 4301
rect 19885 4429 19919 4463
rect 19508 4345 19542 4379
rect 19660 4345 19694 4379
rect 19987 4429 20021 4463
rect 20123 4429 20157 4463
rect 19406 4277 19440 4311
rect 19788 4311 19822 4345
rect 19920 4255 19954 4289
rect 20291 4329 20325 4363
rect 20183 4277 20217 4311
rect 20429 4345 20463 4379
rect 20560 4317 20594 4351
rect 20660 4313 20694 4347
rect 20936 4313 20970 4347
rect 21096 4328 21130 4362
rect 21596 4429 21630 4463
rect 21732 4429 21766 4463
rect 21198 4328 21232 4362
rect 21414 4315 21448 4349
rect 21530 4255 21564 4289
rect 21626 4267 21660 4301
rect 22277 4429 22311 4463
rect 21900 4345 21934 4379
rect 22052 4345 22086 4379
rect 22379 4429 22413 4463
rect 22515 4429 22549 4463
rect 21798 4277 21832 4311
rect 22180 4311 22214 4345
rect 22312 4255 22346 4289
rect 22683 4329 22717 4363
rect 22575 4277 22609 4311
rect 22821 4345 22855 4379
rect 22952 4317 22986 4351
rect 23052 4313 23086 4347
rect 23328 4313 23362 4347
rect 26043 4090 26077 4124
rect 25609 4017 25643 4051
rect 25711 4017 25745 4051
rect 26139 4078 26173 4112
rect 25927 4030 25961 4064
rect 26311 4068 26345 4102
rect 26109 3916 26143 3950
rect 26245 3916 26279 3950
rect 26825 4090 26859 4124
rect 26413 4000 26447 4034
rect 26565 4000 26599 4034
rect 26693 4034 26727 4068
rect 27088 4068 27122 4102
rect 26790 3916 26824 3950
rect 26892 3916 26926 3950
rect 27028 3916 27062 3950
rect 27196 4016 27230 4050
rect 27334 4000 27368 4034
rect 27465 4028 27499 4062
rect 27565 4032 27599 4066
rect 27841 4032 27875 4066
rect 28435 4090 28469 4124
rect 28001 4017 28035 4051
rect 28103 4017 28137 4051
rect 28531 4078 28565 4112
rect 28319 4030 28353 4064
rect 28703 4068 28737 4102
rect 28501 3916 28535 3950
rect 28637 3916 28671 3950
rect 29217 4090 29251 4124
rect 28805 4000 28839 4034
rect 28957 4000 28991 4034
rect 29085 4034 29119 4068
rect 29480 4068 29514 4102
rect 29182 3916 29216 3950
rect 29284 3916 29318 3950
rect 29420 3916 29454 3950
rect 29588 4016 29622 4050
rect 29726 4000 29760 4034
rect 29857 4028 29891 4062
rect 29957 4032 29991 4066
rect 30233 4032 30267 4066
rect 11590 3440 11624 3474
rect 11866 3440 11900 3474
rect 11966 3444 12000 3478
rect 12097 3472 12131 3506
rect 12235 3456 12269 3490
rect 12403 3556 12437 3590
rect 12539 3556 12573 3590
rect 12641 3556 12675 3590
rect 12343 3404 12377 3438
rect 12738 3438 12772 3472
rect 12866 3472 12900 3506
rect 13018 3472 13052 3506
rect 12606 3382 12640 3416
rect 13186 3556 13220 3590
rect 13322 3556 13356 3590
rect 13120 3404 13154 3438
rect 13504 3442 13538 3476
rect 13292 3394 13326 3428
rect 13720 3455 13754 3489
rect 13822 3455 13856 3489
rect 13388 3382 13422 3416
rect 13982 3440 14016 3474
rect 14258 3440 14292 3474
rect 14358 3444 14392 3478
rect 14489 3472 14523 3506
rect 14627 3456 14661 3490
rect 14795 3556 14829 3590
rect 14931 3556 14965 3590
rect 15033 3556 15067 3590
rect 14735 3404 14769 3438
rect 15130 3438 15164 3472
rect 15258 3472 15292 3506
rect 15410 3472 15444 3506
rect 14998 3382 15032 3416
rect 15578 3556 15612 3590
rect 15714 3556 15748 3590
rect 15512 3404 15546 3438
rect 15896 3442 15930 3476
rect 15684 3394 15718 3428
rect 16112 3455 16146 3489
rect 16214 3455 16248 3489
rect 15780 3382 15814 3416
rect 16374 3440 16408 3474
rect 16650 3440 16684 3474
rect 16750 3444 16784 3478
rect 16881 3472 16915 3506
rect 17019 3456 17053 3490
rect 17187 3556 17221 3590
rect 17323 3556 17357 3590
rect 17425 3556 17459 3590
rect 17127 3404 17161 3438
rect 17522 3438 17556 3472
rect 17650 3472 17684 3506
rect 17802 3472 17836 3506
rect 17390 3382 17424 3416
rect 17970 3556 18004 3590
rect 18106 3556 18140 3590
rect 17904 3404 17938 3438
rect 18288 3442 18322 3476
rect 18076 3394 18110 3428
rect 18504 3455 18538 3489
rect 18606 3455 18640 3489
rect 18172 3382 18206 3416
rect 18766 3440 18800 3474
rect 19042 3440 19076 3474
rect 19142 3444 19176 3478
rect 19273 3472 19307 3506
rect 19411 3456 19445 3490
rect 19579 3556 19613 3590
rect 19715 3556 19749 3590
rect 19817 3556 19851 3590
rect 19519 3404 19553 3438
rect 19914 3438 19948 3472
rect 20042 3472 20076 3506
rect 20194 3472 20228 3506
rect 19782 3382 19816 3416
rect 20362 3556 20396 3590
rect 20498 3556 20532 3590
rect 20296 3404 20330 3438
rect 20680 3442 20714 3476
rect 20468 3394 20502 3428
rect 20896 3455 20930 3489
rect 20998 3455 21032 3489
rect 20564 3382 20598 3416
rect 21158 3440 21192 3474
rect 21434 3440 21468 3474
rect 21534 3444 21568 3478
rect 21665 3472 21699 3506
rect 21803 3456 21837 3490
rect 21971 3556 22005 3590
rect 22107 3556 22141 3590
rect 22209 3556 22243 3590
rect 21911 3404 21945 3438
rect 22306 3438 22340 3472
rect 22434 3472 22468 3506
rect 22586 3472 22620 3506
rect 22174 3382 22208 3416
rect 22754 3556 22788 3590
rect 22890 3556 22924 3590
rect 22688 3404 22722 3438
rect 23072 3442 23106 3476
rect 22860 3394 22894 3428
rect 23288 3455 23322 3489
rect 23390 3455 23424 3489
rect 22956 3382 22990 3416
rect 25609 3327 25643 3361
rect 26109 3428 26143 3462
rect 26245 3428 26279 3462
rect 25711 3327 25745 3361
rect 25927 3314 25961 3348
rect 26043 3254 26077 3288
rect 26139 3266 26173 3300
rect 26790 3428 26824 3462
rect 26413 3344 26447 3378
rect 26565 3344 26599 3378
rect 26892 3428 26926 3462
rect 27028 3428 27062 3462
rect 26311 3276 26345 3310
rect 26693 3310 26727 3344
rect 26825 3254 26859 3288
rect 27196 3328 27230 3362
rect 27088 3276 27122 3310
rect 27334 3344 27368 3378
rect 27465 3316 27499 3350
rect 27565 3312 27599 3346
rect 27841 3312 27875 3346
rect 28001 3327 28035 3361
rect 28501 3428 28535 3462
rect 28637 3428 28671 3462
rect 28103 3327 28137 3361
rect 28319 3314 28353 3348
rect 28435 3254 28469 3288
rect 28531 3266 28565 3300
rect 29182 3428 29216 3462
rect 28805 3344 28839 3378
rect 28957 3344 28991 3378
rect 29284 3428 29318 3462
rect 29420 3428 29454 3462
rect 28703 3276 28737 3310
rect 29085 3310 29119 3344
rect 29217 3254 29251 3288
rect 29588 3328 29622 3362
rect 29480 3276 29514 3310
rect 29726 3344 29760 3378
rect 29857 3316 29891 3350
rect 29957 3312 29991 3346
rect 30233 3312 30267 3346
rect 26043 2810 26077 2844
rect 25609 2737 25643 2771
rect 25711 2737 25745 2771
rect 26139 2798 26173 2832
rect 25927 2750 25961 2784
rect 26311 2788 26345 2822
rect 26109 2636 26143 2670
rect 26245 2636 26279 2670
rect 26825 2810 26859 2844
rect 26413 2720 26447 2754
rect 26565 2720 26599 2754
rect 26693 2754 26727 2788
rect 27088 2788 27122 2822
rect 26790 2636 26824 2670
rect 26892 2636 26926 2670
rect 27028 2636 27062 2670
rect 27196 2736 27230 2770
rect 27334 2720 27368 2754
rect 27465 2748 27499 2782
rect 27565 2752 27599 2786
rect 27841 2752 27875 2786
rect 28435 2810 28469 2844
rect 28001 2737 28035 2771
rect 28103 2737 28137 2771
rect 28531 2798 28565 2832
rect 28319 2750 28353 2784
rect 28703 2788 28737 2822
rect 28501 2636 28535 2670
rect 28637 2636 28671 2670
rect 29217 2810 29251 2844
rect 28805 2720 28839 2754
rect 28957 2720 28991 2754
rect 29085 2754 29119 2788
rect 29480 2788 29514 2822
rect 29182 2636 29216 2670
rect 29284 2636 29318 2670
rect 29420 2636 29454 2670
rect 29588 2736 29622 2770
rect 29726 2720 29760 2754
rect 29857 2748 29891 2782
rect 29957 2752 29991 2786
rect 30233 2752 30267 2786
rect 25609 2047 25643 2081
rect 26109 2148 26143 2182
rect 26245 2148 26279 2182
rect 25711 2047 25745 2081
rect 25927 2034 25961 2068
rect 26043 1974 26077 2008
rect 26139 1986 26173 2020
rect 26790 2148 26824 2182
rect 26413 2064 26447 2098
rect 26565 2064 26599 2098
rect 26892 2148 26926 2182
rect 27028 2148 27062 2182
rect 26311 1996 26345 2030
rect 26693 2030 26727 2064
rect 26825 1974 26859 2008
rect 27196 2048 27230 2082
rect 27088 1996 27122 2030
rect 27334 2064 27368 2098
rect 27465 2036 27499 2070
rect 27565 2032 27599 2066
rect 27841 2032 27875 2066
rect 28001 2047 28035 2081
rect 28501 2148 28535 2182
rect 28637 2148 28671 2182
rect 28103 2047 28137 2081
rect 28319 2034 28353 2068
rect 28435 1974 28469 2008
rect 28531 1986 28565 2020
rect 29182 2148 29216 2182
rect 28805 2064 28839 2098
rect 28957 2064 28991 2098
rect 29284 2148 29318 2182
rect 29420 2148 29454 2182
rect 28703 1996 28737 2030
rect 29085 2030 29119 2064
rect 29217 1974 29251 2008
rect 29588 2048 29622 2082
rect 29480 1996 29514 2030
rect 29726 2064 29760 2098
rect 29857 2036 29891 2070
rect 29957 2032 29991 2066
rect 30233 2032 30267 2066
rect 8614 1060 8648 1094
rect 8732 1073 8766 1107
rect 8897 1060 8931 1094
rect 9031 1060 9065 1094
rect 9508 1060 9542 1094
rect 9576 1060 9610 1094
rect 9644 1060 9678 1094
rect 9712 1060 9746 1094
rect 9780 1060 9814 1094
rect 9848 1060 9882 1094
rect 10008 1060 10042 1094
rect 10076 1060 10110 1094
rect 10144 1060 10178 1094
rect 10212 1060 10246 1094
rect 10280 1060 10314 1094
rect 10348 1060 10382 1094
rect 10416 1060 10450 1094
rect 10484 1060 10518 1094
rect 10552 1060 10586 1094
rect 10620 1060 10654 1094
rect 10688 1060 10722 1094
rect 10756 1060 10790 1094
rect 10824 1060 10858 1094
rect 10892 1060 10926 1094
rect 10960 1060 10994 1094
rect 11028 1060 11062 1094
rect 11096 1060 11130 1094
rect 11164 1060 11198 1094
rect 11232 1060 11266 1094
rect 12998 1060 13032 1094
rect 13116 1073 13150 1107
rect 13281 1060 13315 1094
rect 13415 1060 13449 1094
rect 13892 1060 13926 1094
rect 13960 1060 13994 1094
rect 14028 1060 14062 1094
rect 14096 1060 14130 1094
rect 14164 1060 14198 1094
rect 14232 1060 14266 1094
rect 14392 1060 14426 1094
rect 14460 1060 14494 1094
rect 14528 1060 14562 1094
rect 14596 1060 14630 1094
rect 14664 1060 14698 1094
rect 14732 1060 14766 1094
rect 14800 1060 14834 1094
rect 14868 1060 14902 1094
rect 14936 1060 14970 1094
rect 15004 1060 15038 1094
rect 15072 1060 15106 1094
rect 15140 1060 15174 1094
rect 15208 1060 15242 1094
rect 15276 1060 15310 1094
rect 15344 1060 15378 1094
rect 15412 1060 15446 1094
rect 15480 1060 15514 1094
rect 15548 1060 15582 1094
rect 15616 1060 15650 1094
rect 8661 -82 8695 -48
rect 8757 -82 8791 -48
rect 9066 -5 9100 29
rect 8898 -118 8932 -84
rect 9234 -5 9268 29
rect 8994 -118 9028 -84
rect 9156 -118 9190 -84
rect 10144 -5 10178 29
rect 10312 -5 10346 29
rect 10222 -118 10256 -84
rect 10384 -118 10418 -84
rect 10480 -118 10514 -84
rect 10621 -82 10655 -48
rect 10717 -82 10751 -48
rect 11053 -82 11087 -48
rect 11149 -82 11183 -48
rect 11458 -5 11492 29
rect 11290 -118 11324 -84
rect 11626 -5 11660 29
rect 11386 -118 11420 -84
rect 11548 -118 11582 -84
rect 12536 -5 12570 29
rect 12704 -5 12738 29
rect 12614 -118 12648 -84
rect 12776 -118 12810 -84
rect 12872 -118 12906 -84
rect 13013 -82 13047 -48
rect 13109 -82 13143 -48
rect 13445 -82 13479 -48
rect 13541 -82 13575 -48
rect 13850 -5 13884 29
rect 13682 -118 13716 -84
rect 14018 -5 14052 29
rect 13778 -118 13812 -84
rect 13940 -118 13974 -84
rect 14926 -5 14960 29
rect 15094 -5 15128 29
rect 15004 -118 15038 -84
rect 15166 -118 15200 -84
rect 15262 -118 15296 -84
rect 15403 -82 15437 -48
rect 15499 -82 15533 -48
rect 15837 -82 15871 -48
rect 15933 -82 15967 -48
rect 16242 -5 16276 29
rect 16074 -118 16108 -84
rect 16410 -5 16444 29
rect 16170 -118 16204 -84
rect 16332 -118 16366 -84
rect 17320 -5 17354 29
rect 17488 -5 17522 29
rect 17398 -118 17432 -84
rect 17560 -118 17594 -84
rect 17656 -118 17690 -84
rect 17797 -82 17831 -48
rect 17893 -82 17927 -48
rect 18229 -82 18263 -48
rect 18325 -82 18359 -48
rect 18634 -5 18668 29
rect 18466 -118 18500 -84
rect 18802 -5 18836 29
rect 18562 -118 18596 -84
rect 18724 -118 18758 -84
rect 19712 -5 19746 29
rect 19880 -5 19914 29
rect 19790 -118 19824 -84
rect 19952 -118 19986 -84
rect 20048 -118 20082 -84
rect 20189 -82 20223 -48
rect 20285 -82 20319 -48
rect 20621 -82 20655 -48
rect 20717 -82 20751 -48
rect 21026 -5 21060 29
rect 20858 -118 20892 -84
rect 21194 -5 21228 29
rect 20954 -118 20988 -84
rect 21116 -118 21150 -84
rect 22102 -5 22136 29
rect 22270 -5 22304 29
rect 22180 -118 22214 -84
rect 22342 -118 22376 -84
rect 22438 -118 22472 -84
rect 22579 -82 22613 -48
rect 22675 -82 22709 -48
rect 23013 -82 23047 -48
rect 23109 -82 23143 -48
rect 23418 -5 23452 29
rect 23250 -118 23284 -84
rect 23586 -5 23620 29
rect 23346 -118 23380 -84
rect 23508 -118 23542 -84
rect 24496 -5 24530 29
rect 24664 -5 24698 29
rect 24574 -118 24608 -84
rect 24736 -118 24770 -84
rect 24832 -118 24866 -84
rect 24973 -82 25007 -48
rect 25069 -82 25103 -48
rect 10476 -441 10510 -407
rect 12868 -442 12902 -408
rect 8606 -755 8640 -721
rect 9106 -654 9140 -620
rect 9242 -654 9276 -620
rect 8708 -755 8742 -721
rect 8924 -768 8958 -734
rect 9040 -828 9074 -794
rect 9136 -816 9170 -782
rect 9787 -654 9821 -620
rect 9410 -738 9444 -704
rect 9562 -738 9596 -704
rect 9889 -654 9923 -620
rect 10025 -654 10059 -620
rect 9308 -806 9342 -772
rect 9690 -772 9724 -738
rect 9822 -828 9856 -794
rect 15260 -442 15294 -408
rect 17652 -441 17686 -407
rect 20044 -441 20078 -407
rect 22436 -442 22470 -408
rect 10193 -754 10227 -720
rect 10329 -738 10363 -704
rect 10086 -806 10120 -772
rect 10438 -766 10472 -732
rect 10566 -770 10600 -736
rect 10840 -770 10874 -736
rect 10998 -755 11032 -721
rect 11498 -654 11532 -620
rect 11634 -654 11668 -620
rect 11100 -755 11134 -721
rect 11316 -768 11350 -734
rect 11432 -828 11466 -794
rect 11528 -816 11562 -782
rect 12179 -654 12213 -620
rect 11802 -738 11836 -704
rect 11954 -738 11988 -704
rect 12281 -654 12315 -620
rect 12417 -654 12451 -620
rect 11700 -806 11734 -772
rect 12082 -772 12116 -738
rect 12214 -828 12248 -794
rect 12585 -754 12619 -720
rect 12721 -738 12755 -704
rect 12478 -806 12512 -772
rect 12830 -766 12864 -732
rect 12958 -770 12992 -736
rect 13232 -770 13266 -736
rect 13390 -755 13424 -721
rect 13890 -654 13924 -620
rect 14026 -654 14060 -620
rect 13492 -755 13526 -721
rect 13708 -768 13742 -734
rect 13824 -828 13858 -794
rect 13920 -816 13954 -782
rect 14571 -654 14605 -620
rect 14194 -738 14228 -704
rect 14346 -738 14380 -704
rect 14673 -654 14707 -620
rect 14809 -654 14843 -620
rect 14092 -806 14126 -772
rect 14474 -772 14508 -738
rect 14606 -828 14640 -794
rect 14977 -754 15011 -720
rect 15113 -738 15147 -704
rect 14870 -806 14904 -772
rect 15222 -766 15256 -732
rect 15350 -770 15384 -736
rect 15624 -770 15658 -736
rect 15782 -755 15816 -721
rect 16282 -654 16316 -620
rect 16418 -654 16452 -620
rect 15884 -755 15918 -721
rect 16100 -768 16134 -734
rect 16216 -828 16250 -794
rect 16312 -816 16346 -782
rect 16963 -654 16997 -620
rect 16586 -738 16620 -704
rect 16738 -738 16772 -704
rect 17065 -654 17099 -620
rect 17201 -654 17235 -620
rect 16484 -806 16518 -772
rect 16866 -772 16900 -738
rect 16998 -828 17032 -794
rect 17369 -754 17403 -720
rect 17505 -738 17539 -704
rect 17262 -806 17296 -772
rect 17614 -766 17648 -732
rect 17742 -770 17776 -736
rect 18016 -770 18050 -736
rect 18174 -755 18208 -721
rect 18674 -654 18708 -620
rect 18810 -654 18844 -620
rect 18276 -755 18310 -721
rect 18492 -768 18526 -734
rect 18608 -828 18642 -794
rect 18704 -816 18738 -782
rect 19355 -654 19389 -620
rect 18978 -738 19012 -704
rect 19130 -738 19164 -704
rect 19457 -654 19491 -620
rect 19593 -654 19627 -620
rect 18876 -806 18910 -772
rect 19258 -772 19292 -738
rect 19390 -828 19424 -794
rect 24828 -442 24862 -408
rect 19761 -754 19795 -720
rect 19897 -738 19931 -704
rect 19654 -806 19688 -772
rect 20006 -766 20040 -732
rect 20134 -770 20168 -736
rect 20408 -770 20442 -736
rect 20566 -755 20600 -721
rect 21066 -654 21100 -620
rect 21202 -654 21236 -620
rect 20668 -755 20702 -721
rect 20884 -768 20918 -734
rect 21000 -828 21034 -794
rect 21096 -816 21130 -782
rect 21747 -654 21781 -620
rect 21370 -738 21404 -704
rect 21522 -738 21556 -704
rect 21849 -654 21883 -620
rect 21985 -654 22019 -620
rect 21268 -806 21302 -772
rect 21650 -772 21684 -738
rect 21782 -828 21816 -794
rect 22153 -754 22187 -720
rect 22289 -738 22323 -704
rect 22046 -806 22080 -772
rect 22398 -766 22432 -732
rect 22526 -770 22560 -736
rect 22800 -770 22834 -736
rect 22958 -755 22992 -721
rect 23458 -654 23492 -620
rect 23594 -654 23628 -620
rect 23060 -755 23094 -721
rect 23276 -768 23310 -734
rect 23392 -828 23426 -794
rect 23488 -816 23522 -782
rect 24139 -654 24173 -620
rect 23762 -738 23796 -704
rect 23914 -738 23948 -704
rect 24241 -654 24275 -620
rect 24377 -654 24411 -620
rect 23660 -806 23694 -772
rect 24042 -772 24076 -738
rect 24174 -828 24208 -794
rect 24545 -754 24579 -720
rect 24681 -738 24715 -704
rect 24438 -806 24472 -772
rect 24790 -766 24824 -732
rect 24918 -770 24952 -736
rect 25192 -770 25226 -736
rect 10182 -1127 10216 -1093
rect 12574 -1127 12608 -1093
rect 14966 -1127 15000 -1093
rect 17358 -1127 17392 -1093
rect 19750 -1127 19784 -1093
rect 22142 -1127 22176 -1093
rect 24534 -1130 24568 -1096
rect 8668 -1459 8702 -1425
rect 8942 -1459 8976 -1425
rect 9070 -1455 9104 -1421
rect 9179 -1427 9213 -1393
rect 9315 -1443 9349 -1409
rect 9483 -1343 9517 -1309
rect 9619 -1343 9653 -1309
rect 9721 -1343 9755 -1309
rect 9422 -1495 9456 -1461
rect 9818 -1461 9852 -1427
rect 9946 -1427 9980 -1393
rect 10098 -1427 10132 -1393
rect 9686 -1517 9720 -1483
rect 10266 -1343 10300 -1309
rect 10402 -1343 10436 -1309
rect 10200 -1495 10234 -1461
rect 10584 -1457 10618 -1423
rect 10372 -1505 10406 -1471
rect 10800 -1444 10834 -1410
rect 10902 -1444 10936 -1410
rect 10468 -1517 10502 -1483
rect 11060 -1459 11094 -1425
rect 11334 -1459 11368 -1425
rect 11462 -1455 11496 -1421
rect 11571 -1427 11605 -1393
rect 11707 -1443 11741 -1409
rect 11875 -1343 11909 -1309
rect 12011 -1343 12045 -1309
rect 12113 -1343 12147 -1309
rect 11814 -1495 11848 -1461
rect 12210 -1461 12244 -1427
rect 12338 -1427 12372 -1393
rect 12490 -1427 12524 -1393
rect 12078 -1517 12112 -1483
rect 12658 -1343 12692 -1309
rect 12794 -1343 12828 -1309
rect 12592 -1495 12626 -1461
rect 12976 -1457 13010 -1423
rect 12764 -1505 12798 -1471
rect 13192 -1444 13226 -1410
rect 13294 -1444 13328 -1410
rect 12860 -1517 12894 -1483
rect 13452 -1459 13486 -1425
rect 13726 -1459 13760 -1425
rect 13854 -1455 13888 -1421
rect 13963 -1427 13997 -1393
rect 14099 -1443 14133 -1409
rect 14267 -1343 14301 -1309
rect 14403 -1343 14437 -1309
rect 14505 -1343 14539 -1309
rect 14206 -1495 14240 -1461
rect 14602 -1461 14636 -1427
rect 14730 -1427 14764 -1393
rect 14882 -1427 14916 -1393
rect 14470 -1517 14504 -1483
rect 15050 -1343 15084 -1309
rect 15186 -1343 15220 -1309
rect 14984 -1495 15018 -1461
rect 15368 -1457 15402 -1423
rect 15156 -1505 15190 -1471
rect 15584 -1444 15618 -1410
rect 15686 -1444 15720 -1410
rect 15252 -1517 15286 -1483
rect 15844 -1459 15878 -1425
rect 16118 -1459 16152 -1425
rect 16246 -1455 16280 -1421
rect 16355 -1427 16389 -1393
rect 16491 -1443 16525 -1409
rect 16659 -1343 16693 -1309
rect 16795 -1343 16829 -1309
rect 16897 -1343 16931 -1309
rect 16598 -1495 16632 -1461
rect 16994 -1461 17028 -1427
rect 17122 -1427 17156 -1393
rect 17274 -1427 17308 -1393
rect 16862 -1517 16896 -1483
rect 17442 -1343 17476 -1309
rect 17578 -1343 17612 -1309
rect 17376 -1495 17410 -1461
rect 17760 -1457 17794 -1423
rect 17548 -1505 17582 -1471
rect 17976 -1444 18010 -1410
rect 18078 -1444 18112 -1410
rect 17644 -1517 17678 -1483
rect 18236 -1459 18270 -1425
rect 18510 -1459 18544 -1425
rect 18638 -1455 18672 -1421
rect 18747 -1427 18781 -1393
rect 18883 -1443 18917 -1409
rect 19051 -1343 19085 -1309
rect 19187 -1343 19221 -1309
rect 19289 -1343 19323 -1309
rect 18990 -1495 19024 -1461
rect 19386 -1461 19420 -1427
rect 19514 -1427 19548 -1393
rect 19666 -1427 19700 -1393
rect 19254 -1517 19288 -1483
rect 19834 -1343 19868 -1309
rect 19970 -1343 20004 -1309
rect 19768 -1495 19802 -1461
rect 20152 -1457 20186 -1423
rect 19940 -1505 19974 -1471
rect 20368 -1444 20402 -1410
rect 20470 -1444 20504 -1410
rect 20036 -1517 20070 -1483
rect 20628 -1459 20662 -1425
rect 20902 -1459 20936 -1425
rect 21030 -1455 21064 -1421
rect 21139 -1427 21173 -1393
rect 21275 -1443 21309 -1409
rect 21443 -1343 21477 -1309
rect 21579 -1343 21613 -1309
rect 21681 -1343 21715 -1309
rect 21382 -1495 21416 -1461
rect 21778 -1461 21812 -1427
rect 21906 -1427 21940 -1393
rect 22058 -1427 22092 -1393
rect 21646 -1517 21680 -1483
rect 22226 -1343 22260 -1309
rect 22362 -1343 22396 -1309
rect 22160 -1495 22194 -1461
rect 22544 -1457 22578 -1423
rect 22332 -1505 22366 -1471
rect 22760 -1444 22794 -1410
rect 22862 -1444 22896 -1410
rect 22428 -1517 22462 -1483
rect 23020 -1459 23054 -1425
rect 23294 -1459 23328 -1425
rect 23422 -1455 23456 -1421
rect 23531 -1427 23565 -1393
rect 23667 -1443 23701 -1409
rect 23835 -1343 23869 -1309
rect 23971 -1343 24005 -1309
rect 24073 -1343 24107 -1309
rect 23774 -1495 23808 -1461
rect 24170 -1461 24204 -1427
rect 24298 -1427 24332 -1393
rect 24450 -1427 24484 -1393
rect 24038 -1517 24072 -1483
rect 24618 -1343 24652 -1309
rect 24754 -1343 24788 -1309
rect 24552 -1495 24586 -1461
rect 24936 -1457 24970 -1423
rect 24724 -1505 24758 -1471
rect 25152 -1444 25186 -1410
rect 25254 -1444 25288 -1410
rect 24820 -1517 24854 -1483
<< locali >>
rect 13946 13605 14616 13623
rect 13946 13597 14062 13605
rect 13816 13581 13850 13597
rect 13816 13505 13850 13521
rect 13904 13581 14062 13597
rect 13938 13571 14062 13581
rect 14098 13571 14142 13605
rect 14178 13571 14222 13605
rect 14258 13571 14302 13605
rect 14338 13571 14382 13605
rect 14418 13571 14462 13605
rect 14498 13571 14616 13605
rect 13938 13557 14616 13571
rect 14678 13608 19586 13626
rect 14678 13574 14794 13608
rect 14830 13574 14874 13608
rect 14910 13574 14954 13608
rect 14990 13574 15034 13608
rect 15070 13574 15114 13608
rect 15150 13574 15194 13608
rect 15230 13574 15398 13608
rect 15434 13574 15478 13608
rect 15514 13574 15558 13608
rect 15594 13574 15638 13608
rect 15674 13574 15718 13608
rect 15754 13574 15798 13608
rect 15834 13574 16006 13608
rect 16042 13574 16086 13608
rect 16122 13574 16166 13608
rect 16202 13574 16246 13608
rect 16282 13574 16326 13608
rect 16362 13574 16406 13608
rect 16442 13574 16610 13608
rect 16646 13574 16690 13608
rect 16726 13574 16770 13608
rect 16806 13574 16850 13608
rect 16886 13574 16930 13608
rect 16966 13574 17010 13608
rect 17046 13574 17218 13608
rect 17254 13574 17298 13608
rect 17334 13574 17378 13608
rect 17414 13574 17458 13608
rect 17494 13574 17538 13608
rect 17574 13574 17618 13608
rect 17654 13574 17822 13608
rect 17858 13574 17902 13608
rect 17938 13574 17982 13608
rect 18018 13574 18062 13608
rect 18098 13574 18142 13608
rect 18178 13574 18222 13608
rect 18258 13574 18430 13608
rect 18466 13574 18510 13608
rect 18546 13574 18590 13608
rect 18626 13574 18670 13608
rect 18706 13574 18750 13608
rect 18786 13574 18830 13608
rect 18866 13574 19034 13608
rect 19070 13574 19114 13608
rect 19150 13574 19194 13608
rect 19230 13574 19274 13608
rect 19310 13574 19354 13608
rect 19390 13574 19434 13608
rect 19470 13574 19586 13608
rect 20655 13605 21325 13623
rect 20655 13597 20771 13605
rect 14678 13560 19586 13574
rect 19750 13557 19836 13583
rect 13938 13521 14074 13557
rect 13904 13516 14074 13521
rect 13904 13505 13938 13516
rect 13816 13443 13850 13459
rect 13816 13367 13850 13383
rect 13904 13443 13938 13459
rect 14017 13452 14074 13516
rect 19750 13523 19776 13557
rect 19810 13523 19836 13557
rect 19750 13497 19836 13523
rect 20227 13560 20313 13586
rect 20227 13526 20253 13560
rect 20287 13526 20313 13560
rect 20227 13500 20313 13526
rect 20525 13581 20559 13597
rect 20525 13505 20559 13521
rect 20613 13581 20771 13597
rect 20647 13571 20771 13581
rect 20807 13571 20851 13605
rect 20887 13571 20931 13605
rect 20967 13571 21011 13605
rect 21047 13571 21091 13605
rect 21127 13571 21171 13605
rect 21207 13571 21325 13605
rect 20647 13557 21325 13571
rect 21387 13608 26295 13626
rect 21387 13574 21503 13608
rect 21539 13574 21583 13608
rect 21619 13574 21663 13608
rect 21699 13574 21743 13608
rect 21779 13574 21823 13608
rect 21859 13574 21903 13608
rect 21939 13574 22107 13608
rect 22143 13574 22187 13608
rect 22223 13574 22267 13608
rect 22303 13574 22347 13608
rect 22383 13574 22427 13608
rect 22463 13574 22507 13608
rect 22543 13574 22715 13608
rect 22751 13574 22795 13608
rect 22831 13574 22875 13608
rect 22911 13574 22955 13608
rect 22991 13574 23035 13608
rect 23071 13574 23115 13608
rect 23151 13574 23319 13608
rect 23355 13574 23399 13608
rect 23435 13574 23479 13608
rect 23515 13574 23559 13608
rect 23595 13574 23639 13608
rect 23675 13574 23719 13608
rect 23755 13574 23927 13608
rect 23963 13574 24007 13608
rect 24043 13574 24087 13608
rect 24123 13574 24167 13608
rect 24203 13574 24247 13608
rect 24283 13574 24327 13608
rect 24363 13574 24531 13608
rect 24567 13574 24611 13608
rect 24647 13574 24691 13608
rect 24727 13574 24771 13608
rect 24807 13574 24851 13608
rect 24887 13574 24931 13608
rect 24967 13574 25139 13608
rect 25175 13574 25219 13608
rect 25255 13574 25299 13608
rect 25335 13574 25379 13608
rect 25415 13574 25459 13608
rect 25495 13574 25539 13608
rect 25575 13574 25743 13608
rect 25779 13574 25823 13608
rect 25859 13574 25903 13608
rect 25939 13574 25983 13608
rect 26019 13574 26063 13608
rect 26099 13574 26143 13608
rect 26179 13574 26295 13608
rect 21387 13560 26295 13574
rect 26459 13557 26545 13583
rect 20647 13521 20783 13557
rect 20613 13516 20783 13521
rect 20613 13505 20647 13516
rect 13904 13367 13938 13383
rect 14004 13427 14087 13452
rect 20525 13443 20559 13459
rect 14004 13392 14029 13427
rect 14063 13392 14087 13427
rect 14004 13368 14087 13392
rect 19755 13413 19841 13439
rect 19755 13379 19781 13413
rect 19815 13379 19841 13413
rect 19755 13353 19841 13379
rect 20216 13388 20302 13414
rect 20216 13354 20242 13388
rect 20276 13354 20302 13388
rect 20525 13367 20559 13383
rect 20613 13443 20647 13459
rect 20726 13452 20783 13516
rect 26459 13523 26485 13557
rect 26519 13523 26545 13557
rect 26459 13497 26545 13523
rect 20613 13367 20647 13383
rect 20713 13427 20796 13452
rect 20713 13392 20738 13427
rect 20772 13392 20796 13427
rect 20713 13368 20796 13392
rect 26464 13413 26550 13439
rect 26464 13379 26490 13413
rect 26524 13379 26550 13413
rect 20216 13328 20302 13354
rect 26464 13353 26550 13379
rect 13816 13305 13850 13321
rect 13816 13229 13850 13245
rect 13904 13305 13938 13321
rect 20525 13305 20559 13321
rect 13904 13229 13938 13245
rect 19756 13261 19842 13287
rect 19756 13227 19782 13261
rect 19816 13227 19842 13261
rect 20525 13229 20559 13245
rect 20613 13305 20647 13321
rect 20613 13229 20647 13245
rect 26465 13261 26551 13287
rect 19756 13201 19842 13227
rect 26465 13227 26491 13261
rect 26525 13227 26551 13261
rect 20216 13196 20302 13222
rect 26465 13201 26551 13227
rect 13816 13167 13850 13183
rect 3058 13130 3728 13148
rect 3058 13122 3174 13130
rect 2928 13106 2962 13122
rect 2928 13030 2962 13046
rect 3016 13106 3174 13122
rect 3050 13096 3174 13106
rect 3210 13096 3254 13130
rect 3290 13096 3334 13130
rect 3370 13096 3414 13130
rect 3450 13096 3494 13130
rect 3530 13096 3574 13130
rect 3610 13096 3728 13130
rect 3050 13082 3728 13096
rect 3790 13133 8698 13151
rect 3790 13099 3906 13133
rect 3942 13099 3986 13133
rect 4022 13099 4066 13133
rect 4102 13099 4146 13133
rect 4182 13099 4226 13133
rect 4262 13099 4306 13133
rect 4342 13099 4510 13133
rect 4546 13099 4590 13133
rect 4626 13099 4670 13133
rect 4706 13099 4750 13133
rect 4786 13099 4830 13133
rect 4866 13099 4910 13133
rect 4946 13099 5118 13133
rect 5154 13099 5198 13133
rect 5234 13099 5278 13133
rect 5314 13099 5358 13133
rect 5394 13099 5438 13133
rect 5474 13099 5518 13133
rect 5554 13099 5722 13133
rect 5758 13099 5802 13133
rect 5838 13099 5882 13133
rect 5918 13099 5962 13133
rect 5998 13099 6042 13133
rect 6078 13099 6122 13133
rect 6158 13099 6330 13133
rect 6366 13099 6410 13133
rect 6446 13099 6490 13133
rect 6526 13099 6570 13133
rect 6606 13099 6650 13133
rect 6686 13099 6730 13133
rect 6766 13099 6934 13133
rect 6970 13099 7014 13133
rect 7050 13099 7094 13133
rect 7130 13099 7174 13133
rect 7210 13099 7254 13133
rect 7290 13099 7334 13133
rect 7370 13099 7542 13133
rect 7578 13099 7622 13133
rect 7658 13099 7702 13133
rect 7738 13099 7782 13133
rect 7818 13099 7862 13133
rect 7898 13099 7942 13133
rect 7978 13099 8146 13133
rect 8182 13099 8226 13133
rect 8262 13099 8306 13133
rect 8342 13099 8386 13133
rect 8422 13099 8466 13133
rect 8502 13099 8546 13133
rect 8582 13099 8698 13133
rect 3790 13085 8698 13099
rect 8862 13082 8948 13108
rect 13816 13091 13850 13107
rect 13904 13167 13938 13183
rect 20216 13162 20242 13196
rect 20276 13162 20302 13196
rect 20216 13136 20302 13162
rect 20525 13167 20559 13183
rect 13904 13091 13938 13107
rect 19756 13091 19842 13117
rect 20525 13091 20559 13107
rect 20613 13167 20647 13183
rect 20613 13091 20647 13107
rect 26465 13091 26551 13117
rect 3050 13046 3186 13082
rect 3016 13041 3186 13046
rect 3016 13030 3050 13041
rect 2928 12968 2962 12984
rect 2928 12892 2962 12908
rect 3016 12968 3050 12984
rect 3129 12977 3186 13041
rect 8862 13048 8888 13082
rect 8922 13048 8948 13082
rect 8862 13022 8948 13048
rect 19756 13057 19782 13091
rect 19816 13057 19842 13091
rect 13332 13010 13348 13039
rect 3016 12892 3050 12908
rect 3116 12952 3199 12977
rect 13274 12976 13303 13010
rect 13337 13005 13348 13010
rect 13382 13010 13398 13039
rect 13462 13010 13478 13039
rect 13512 13010 13532 13039
rect 13608 13010 13624 13039
rect 13382 13005 13395 13010
rect 13337 12976 13395 13005
rect 13429 13005 13478 13010
rect 13429 12976 13487 13005
rect 13521 12976 13579 13010
rect 13613 13005 13624 13010
rect 13658 13010 13678 13039
rect 13816 13029 13850 13045
rect 13658 13005 13671 13010
rect 13613 12976 13671 13005
rect 13705 12976 13734 13010
rect 3116 12917 3141 12952
rect 3175 12917 3199 12952
rect 3116 12893 3199 12917
rect 8867 12938 8953 12964
rect 8867 12904 8893 12938
rect 8927 12904 8953 12938
rect 8867 12878 8953 12904
rect 13342 12934 13384 12976
rect 13342 12900 13350 12934
rect 13342 12866 13384 12900
rect 2928 12830 2962 12846
rect 2928 12754 2962 12770
rect 3016 12830 3050 12846
rect 13342 12832 13350 12866
rect 3016 12754 3050 12770
rect 8868 12786 8954 12812
rect 8868 12752 8894 12786
rect 8928 12752 8954 12786
rect 8868 12726 8954 12752
rect 13342 12798 13384 12832
rect 13342 12764 13350 12798
rect 13342 12748 13384 12764
rect 13418 12934 13484 12942
rect 13418 12900 13434 12934
rect 13468 12900 13484 12934
rect 13418 12867 13484 12900
rect 13418 12833 13431 12867
rect 13465 12866 13484 12867
rect 13418 12832 13434 12833
rect 13468 12832 13484 12866
rect 13418 12798 13484 12832
rect 13418 12764 13434 12798
rect 13468 12764 13484 12798
rect 13418 12746 13484 12764
rect 2928 12692 2962 12708
rect 2928 12616 2962 12632
rect 3016 12692 3050 12708
rect 13338 12702 13404 12712
rect 13338 12668 13350 12702
rect 13384 12698 13404 12702
rect 13338 12664 13354 12668
rect 13388 12664 13404 12698
rect 3016 12616 3050 12632
rect 8868 12616 8954 12642
rect 8868 12582 8894 12616
rect 8928 12582 8954 12616
rect 2444 12535 2460 12564
rect 2386 12501 2415 12535
rect 2449 12530 2460 12535
rect 2494 12535 2510 12564
rect 2574 12535 2590 12564
rect 2624 12535 2644 12564
rect 2720 12535 2736 12564
rect 2494 12530 2507 12535
rect 2449 12501 2507 12530
rect 2541 12530 2590 12535
rect 2541 12501 2599 12530
rect 2633 12501 2691 12535
rect 2725 12530 2736 12535
rect 2770 12535 2790 12564
rect 2928 12554 2962 12570
rect 2770 12530 2783 12535
rect 2725 12501 2783 12530
rect 2817 12501 2846 12535
rect 2454 12459 2496 12501
rect 2454 12425 2462 12459
rect 2454 12391 2496 12425
rect 2454 12357 2462 12391
rect 2454 12323 2496 12357
rect 2454 12289 2462 12323
rect 2454 12273 2496 12289
rect 2530 12459 2596 12467
rect 2530 12425 2546 12459
rect 2580 12425 2596 12459
rect 2530 12392 2596 12425
rect 2530 12358 2543 12392
rect 2577 12391 2596 12392
rect 2530 12357 2546 12358
rect 2580 12357 2596 12391
rect 2530 12323 2596 12357
rect 2530 12289 2546 12323
rect 2580 12289 2596 12323
rect 2530 12271 2596 12289
rect 2450 12227 2516 12237
rect 2450 12193 2462 12227
rect 2496 12223 2516 12227
rect 2450 12189 2466 12193
rect 2500 12189 2516 12223
rect 2450 12139 2496 12155
rect 2550 12151 2596 12271
rect 2450 12105 2462 12139
rect 2450 12071 2496 12105
rect 2450 12037 2462 12071
rect 2450 11991 2496 12037
rect 2530 12139 2596 12151
rect 2530 12105 2546 12139
rect 2580 12105 2596 12139
rect 2530 12071 2596 12105
rect 2530 12037 2546 12071
rect 2580 12037 2596 12071
rect 2530 12025 2596 12037
rect 2636 12459 2702 12467
rect 2636 12425 2652 12459
rect 2686 12425 2702 12459
rect 2636 12391 2702 12425
rect 2636 12357 2652 12391
rect 2686 12357 2702 12391
rect 2636 12337 2702 12357
rect 2636 12289 2652 12337
rect 2686 12289 2702 12337
rect 2636 12271 2702 12289
rect 2736 12459 2778 12501
rect 2928 12478 2962 12494
rect 3016 12554 3050 12570
rect 8868 12556 8954 12582
rect 13338 12614 13384 12630
rect 13438 12626 13484 12746
rect 13338 12580 13350 12614
rect 13338 12546 13384 12580
rect 13338 12512 13350 12546
rect 3016 12478 3050 12494
rect 2770 12425 2778 12459
rect 8867 12459 8953 12485
rect 2736 12391 2778 12425
rect 2770 12357 2778 12391
rect 2736 12323 2778 12357
rect 2928 12416 2962 12432
rect 2928 12340 2962 12356
rect 3016 12416 3050 12432
rect 8867 12425 8893 12459
rect 8927 12425 8953 12459
rect 10882 12432 10911 12500
rect 10945 12432 11003 12500
rect 11037 12432 11095 12500
rect 11129 12432 11187 12500
rect 11221 12432 11279 12500
rect 11313 12432 11371 12500
rect 11405 12432 11463 12500
rect 11497 12432 11555 12500
rect 11589 12432 11647 12500
rect 11681 12432 11739 12500
rect 11773 12432 11831 12500
rect 11865 12432 11923 12500
rect 11957 12432 12015 12500
rect 12049 12432 12107 12500
rect 12141 12432 12199 12500
rect 12233 12432 12291 12500
rect 12325 12432 12383 12500
rect 12417 12432 12475 12500
rect 12509 12432 12567 12500
rect 12601 12432 12659 12500
rect 12693 12432 12751 12500
rect 12785 12432 12843 12500
rect 12877 12432 12935 12500
rect 12969 12432 13027 12500
rect 13061 12432 13119 12500
rect 13153 12432 13211 12500
rect 13245 12466 13274 12500
rect 13338 12466 13384 12512
rect 13418 12614 13484 12626
rect 13418 12580 13434 12614
rect 13468 12580 13484 12614
rect 13418 12546 13484 12580
rect 13418 12512 13434 12546
rect 13468 12512 13484 12546
rect 13418 12500 13484 12512
rect 13524 12934 13590 12942
rect 13524 12900 13540 12934
rect 13574 12900 13590 12934
rect 13524 12866 13590 12900
rect 13524 12832 13540 12866
rect 13574 12832 13590 12866
rect 13524 12812 13590 12832
rect 13524 12764 13540 12812
rect 13574 12764 13590 12812
rect 13524 12746 13590 12764
rect 13624 12934 13666 12976
rect 13816 12953 13850 12969
rect 13904 13029 13938 13045
rect 19756 13031 19842 13057
rect 26465 13057 26491 13091
rect 26525 13057 26551 13091
rect 20041 13010 20057 13039
rect 19983 12976 20012 13010
rect 20046 13005 20057 13010
rect 20091 13010 20107 13039
rect 20171 13010 20187 13039
rect 20221 13010 20241 13039
rect 20317 13010 20333 13039
rect 20091 13005 20104 13010
rect 20046 12976 20104 13005
rect 20138 13005 20187 13010
rect 20138 12976 20196 13005
rect 20230 12976 20288 13010
rect 20322 13005 20333 13010
rect 20367 13010 20387 13039
rect 20525 13029 20559 13045
rect 20367 13005 20380 13010
rect 20322 12976 20380 13005
rect 20414 12976 20443 13010
rect 13904 12953 13938 12969
rect 13658 12900 13666 12934
rect 19755 12934 19841 12960
rect 13624 12866 13666 12900
rect 13658 12832 13666 12866
rect 13624 12798 13666 12832
rect 13816 12891 13850 12907
rect 13816 12815 13850 12831
rect 13904 12891 13938 12907
rect 19755 12900 19781 12934
rect 19815 12900 19841 12934
rect 19755 12874 19841 12900
rect 20051 12934 20093 12976
rect 20051 12900 20059 12934
rect 13904 12815 13938 12831
rect 20051 12866 20093 12900
rect 20051 12832 20059 12866
rect 13658 12764 13666 12798
rect 20051 12798 20093 12832
rect 13624 12748 13666 12764
rect 13524 12626 13570 12746
rect 13844 12738 13860 12772
rect 13894 12738 13910 12772
rect 20051 12764 20059 12798
rect 20051 12748 20093 12764
rect 20127 12934 20193 12942
rect 20127 12900 20143 12934
rect 20177 12900 20193 12934
rect 20127 12867 20193 12900
rect 20127 12833 20140 12867
rect 20174 12866 20193 12867
rect 20127 12832 20143 12833
rect 20177 12832 20193 12866
rect 20127 12798 20193 12832
rect 20127 12764 20143 12798
rect 20177 12764 20193 12798
rect 20127 12746 20193 12764
rect 13604 12701 13670 12712
rect 13604 12698 13624 12701
rect 13604 12664 13620 12698
rect 13658 12667 13670 12701
rect 13654 12664 13670 12667
rect 13754 12702 13803 12714
rect 13754 12668 13763 12702
rect 13797 12697 13803 12702
rect 20047 12702 20113 12712
rect 13797 12668 14086 12697
rect 13754 12662 14086 12668
rect 20047 12668 20059 12702
rect 20093 12698 20113 12702
rect 20047 12664 20063 12668
rect 20097 12664 20113 12698
rect 13754 12655 13803 12662
rect 14051 12639 14086 12662
rect 13524 12614 13590 12626
rect 13524 12580 13540 12614
rect 13574 12580 13590 12614
rect 13524 12546 13590 12580
rect 13524 12512 13540 12546
rect 13574 12512 13590 12546
rect 13524 12500 13590 12512
rect 13624 12614 13670 12630
rect 14051 12627 14100 12639
rect 13658 12580 13670 12614
rect 13624 12546 13670 12580
rect 13792 12609 13841 12621
rect 13792 12575 13801 12609
rect 13835 12575 14002 12609
rect 14051 12593 14060 12627
rect 14094 12593 14100 12627
rect 20047 12614 20093 12630
rect 20147 12626 20193 12746
rect 14051 12580 14100 12593
rect 19601 12580 19635 12596
rect 13792 12562 13841 12575
rect 13658 12512 13670 12546
rect 13624 12466 13670 12512
rect 13961 12533 14002 12575
rect 14052 12534 14101 12546
rect 14052 12533 14061 12534
rect 13961 12500 14061 12533
rect 14095 12500 14101 12534
rect 13961 12499 14101 12500
rect 14052 12487 14101 12499
rect 14486 12495 14502 12529
rect 14536 12495 14552 12529
rect 15218 12498 15234 12532
rect 15268 12498 15284 12532
rect 15344 12498 15360 12532
rect 15394 12498 15410 12532
rect 16430 12498 16446 12532
rect 16480 12498 16496 12532
rect 16556 12498 16572 12532
rect 16606 12498 16622 12532
rect 17642 12498 17658 12532
rect 17692 12498 17708 12532
rect 17768 12498 17784 12532
rect 17818 12498 17834 12532
rect 18854 12498 18870 12532
rect 18904 12498 18920 12532
rect 18980 12498 18996 12532
rect 19030 12498 19046 12532
rect 19601 12504 19635 12520
rect 19689 12580 19723 12596
rect 19689 12504 19723 12520
rect 20047 12580 20059 12614
rect 20047 12546 20093 12580
rect 20047 12512 20059 12546
rect 20047 12466 20093 12512
rect 20127 12614 20193 12626
rect 20127 12580 20143 12614
rect 20177 12580 20193 12614
rect 20127 12546 20193 12580
rect 20127 12512 20143 12546
rect 20177 12512 20193 12546
rect 20127 12500 20193 12512
rect 20233 12934 20299 12942
rect 20233 12900 20249 12934
rect 20283 12900 20299 12934
rect 20233 12866 20299 12900
rect 20233 12832 20249 12866
rect 20283 12832 20299 12866
rect 20233 12812 20299 12832
rect 20233 12764 20249 12812
rect 20283 12764 20299 12812
rect 20233 12746 20299 12764
rect 20333 12934 20375 12976
rect 20525 12953 20559 12969
rect 20613 13029 20647 13045
rect 26465 13031 26551 13057
rect 20613 12953 20647 12969
rect 20367 12900 20375 12934
rect 26464 12934 26550 12960
rect 20333 12866 20375 12900
rect 20367 12832 20375 12866
rect 20333 12798 20375 12832
rect 20525 12891 20559 12907
rect 20525 12815 20559 12831
rect 20613 12891 20647 12907
rect 26464 12900 26490 12934
rect 26524 12900 26550 12934
rect 26464 12874 26550 12900
rect 20613 12815 20647 12831
rect 20367 12764 20375 12798
rect 20333 12748 20375 12764
rect 20233 12626 20279 12746
rect 20553 12738 20569 12772
rect 20603 12738 20619 12772
rect 20313 12701 20379 12712
rect 20313 12698 20333 12701
rect 20313 12664 20329 12698
rect 20367 12667 20379 12701
rect 20363 12664 20379 12667
rect 20463 12702 20512 12714
rect 20463 12668 20472 12702
rect 20506 12697 20512 12702
rect 20506 12668 20795 12697
rect 20463 12662 20795 12668
rect 20463 12655 20512 12662
rect 20760 12639 20795 12662
rect 20233 12614 20299 12626
rect 20233 12580 20249 12614
rect 20283 12580 20299 12614
rect 20233 12546 20299 12580
rect 20233 12512 20249 12546
rect 20283 12512 20299 12546
rect 20233 12500 20299 12512
rect 20333 12614 20379 12630
rect 20760 12627 20809 12639
rect 20367 12580 20379 12614
rect 20333 12546 20379 12580
rect 20501 12609 20550 12621
rect 20501 12575 20510 12609
rect 20544 12575 20711 12609
rect 20760 12593 20769 12627
rect 20803 12593 20809 12627
rect 20760 12580 20809 12593
rect 26310 12580 26344 12596
rect 20501 12562 20550 12575
rect 20367 12512 20379 12546
rect 20333 12466 20379 12512
rect 20670 12533 20711 12575
rect 20761 12534 20810 12546
rect 20761 12533 20770 12534
rect 20670 12500 20770 12533
rect 20804 12500 20810 12534
rect 20670 12499 20810 12500
rect 20761 12487 20810 12499
rect 21195 12495 21211 12529
rect 21245 12495 21261 12529
rect 21927 12498 21943 12532
rect 21977 12498 21993 12532
rect 22053 12498 22069 12532
rect 22103 12498 22119 12532
rect 23139 12498 23155 12532
rect 23189 12498 23205 12532
rect 23265 12498 23281 12532
rect 23315 12498 23331 12532
rect 24351 12498 24367 12532
rect 24401 12498 24417 12532
rect 24477 12498 24493 12532
rect 24527 12498 24543 12532
rect 25563 12498 25579 12532
rect 25613 12498 25629 12532
rect 25689 12498 25705 12532
rect 25739 12498 25755 12532
rect 26310 12504 26344 12520
rect 26398 12580 26432 12596
rect 26398 12504 26432 12520
rect 13245 12432 13303 12466
rect 13337 12437 13395 12466
rect 13429 12437 13487 12466
rect 13337 12432 13368 12437
rect 13429 12432 13486 12437
rect 13521 12432 13579 12466
rect 13613 12437 13671 12466
rect 13613 12432 13630 12437
rect 8867 12399 8953 12425
rect 10985 12390 11051 12432
rect 3016 12340 3050 12356
rect 10899 12364 10951 12380
rect 2770 12289 2778 12323
rect 10899 12330 10917 12364
rect 10985 12356 11001 12390
rect 11035 12356 11051 12390
rect 11169 12390 11239 12432
rect 11085 12364 11130 12380
rect 10899 12322 10951 12330
rect 11119 12330 11130 12364
rect 11169 12356 11189 12390
rect 11223 12356 11239 12390
rect 11363 12390 11562 12396
rect 11273 12372 11307 12388
rect 2736 12273 2778 12289
rect 2636 12151 2682 12271
rect 2956 12263 2972 12297
rect 3006 12263 3022 12297
rect 10899 12288 11050 12322
rect 2716 12226 2782 12237
rect 2716 12223 2736 12226
rect 2716 12189 2732 12223
rect 2770 12192 2782 12226
rect 2766 12189 2782 12192
rect 2866 12227 2915 12239
rect 2866 12193 2875 12227
rect 2909 12222 2915 12227
rect 2909 12193 3198 12222
rect 10899 12219 10970 12254
rect 2866 12187 3198 12193
rect 2866 12180 2915 12187
rect 3163 12164 3198 12187
rect 9061 12194 9337 12218
rect 9061 12193 9182 12194
rect 2636 12139 2702 12151
rect 2636 12105 2652 12139
rect 2686 12105 2702 12139
rect 2636 12071 2702 12105
rect 2636 12037 2652 12071
rect 2686 12037 2702 12071
rect 2636 12025 2702 12037
rect 2736 12139 2782 12155
rect 3163 12152 3212 12164
rect 2770 12105 2782 12139
rect 2736 12071 2782 12105
rect 2904 12134 2953 12146
rect 2904 12100 2913 12134
rect 2947 12100 3114 12134
rect 3163 12118 3172 12152
rect 3206 12118 3212 12152
rect 9061 12159 9090 12193
rect 9124 12160 9182 12193
rect 9216 12160 9274 12194
rect 9308 12160 9337 12194
rect 9124 12159 9337 12160
rect 9061 12158 9337 12159
rect 9061 12124 9090 12158
rect 9124 12124 9182 12158
rect 9216 12124 9274 12158
rect 9308 12124 9337 12158
rect 10899 12217 10914 12219
rect 10899 12183 10912 12217
rect 10948 12185 10970 12219
rect 10946 12183 10970 12185
rect 10899 12124 10970 12183
rect 11004 12219 11050 12288
rect 11004 12185 11016 12219
rect 3163 12105 3212 12118
rect 8713 12105 8747 12121
rect 2904 12087 2953 12100
rect 2770 12037 2782 12071
rect 2736 11991 2782 12037
rect 3073 12058 3114 12100
rect 3164 12059 3213 12071
rect 3164 12058 3173 12059
rect 3073 12025 3173 12058
rect 3207 12025 3213 12059
rect 3073 12024 3213 12025
rect 3164 12012 3213 12024
rect 3598 12020 3614 12054
rect 3648 12020 3664 12054
rect 4330 12023 4346 12057
rect 4380 12023 4396 12057
rect 4456 12023 4472 12057
rect 4506 12023 4522 12057
rect 5542 12023 5558 12057
rect 5592 12023 5608 12057
rect 5668 12023 5684 12057
rect 5718 12023 5734 12057
rect 6754 12023 6770 12057
rect 6804 12023 6820 12057
rect 6880 12023 6896 12057
rect 6930 12023 6946 12057
rect 7966 12023 7982 12057
rect 8016 12023 8032 12057
rect 8092 12023 8108 12057
rect 8142 12023 8158 12057
rect 8713 12029 8747 12045
rect 8801 12105 8835 12121
rect 8801 12029 8835 12045
rect 9129 12082 9171 12124
rect 11004 12092 11050 12185
rect 9129 12048 9137 12082
rect 9129 12014 9171 12048
rect 2386 11957 2415 11991
rect 2449 11962 2507 11991
rect 2541 11962 2599 11991
rect 2449 11957 2480 11962
rect 2541 11957 2598 11962
rect 2633 11957 2691 11991
rect 2725 11962 2783 11991
rect 2725 11957 2742 11962
rect 2464 11928 2480 11957
rect 2514 11928 2540 11957
rect 2582 11928 2598 11957
rect 2632 11928 2658 11957
rect 2724 11928 2742 11957
rect 2776 11957 2783 11962
rect 2817 11957 2846 11991
rect 3570 11961 3604 11977
rect 2776 11928 2792 11957
rect 3570 11885 3604 11901
rect 3658 11964 3692 11980
rect 3658 11888 3692 11904
rect 4302 11964 4336 11980
rect 4302 11888 4336 11904
rect 4407 11964 4441 11980
rect 4407 11888 4441 11904
rect 4516 11964 4550 11980
rect 4516 11888 4550 11904
rect 5514 11964 5548 11980
rect 5514 11888 5548 11904
rect 5618 11964 5652 11980
rect 5618 11888 5652 11904
rect 5728 11964 5762 11980
rect 5728 11888 5762 11904
rect 6726 11964 6760 11980
rect 6726 11888 6760 11904
rect 6831 11964 6865 11980
rect 6831 11888 6865 11904
rect 6940 11964 6974 11980
rect 6940 11888 6974 11904
rect 7938 11964 7972 11980
rect 7938 11888 7972 11904
rect 8045 11964 8079 11980
rect 8045 11888 8079 11904
rect 8152 11964 8186 11980
rect 8152 11888 8186 11904
rect 8713 11967 8747 11983
rect 8713 11891 8747 11907
rect 8801 11967 8835 11983
rect 8801 11891 8835 11907
rect 8897 11967 8931 11983
rect 8897 11891 8931 11907
rect 8993 11967 9027 11983
rect 8993 11891 9027 11907
rect 9129 11980 9137 12014
rect 9129 11946 9171 11980
rect 9129 11912 9137 11946
rect 9129 11896 9171 11912
rect 9205 12082 9271 12090
rect 9205 12048 9221 12082
rect 9255 12048 9271 12082
rect 9205 12014 9271 12048
rect 9205 11980 9221 12014
rect 9255 11980 9271 12014
rect 9205 11946 9271 11980
rect 10899 12074 11004 12090
rect 10899 12040 10917 12074
rect 10951 12058 11004 12074
rect 11038 12058 11050 12092
rect 10951 12056 11050 12058
rect 11085 12296 11130 12330
rect 11363 12356 11379 12390
rect 11413 12356 11562 12390
rect 11273 12322 11307 12338
rect 11085 12262 11096 12296
rect 11085 12074 11130 12262
rect 10899 12006 10951 12040
rect 11119 12040 11130 12074
rect 11164 12284 11307 12322
rect 11348 12292 11392 12308
rect 11164 12090 11198 12284
rect 11382 12258 11392 12292
rect 11232 12232 11314 12248
rect 11266 12198 11314 12232
rect 11232 12189 11314 12198
rect 11232 12155 11263 12189
rect 11297 12155 11314 12189
rect 11232 12124 11314 12155
rect 11348 12134 11392 12258
rect 11428 12296 11494 12320
rect 11428 12280 11460 12296
rect 11428 12246 11444 12280
rect 11478 12246 11494 12262
rect 11528 12210 11562 12356
rect 11596 12394 11630 12432
rect 11596 12344 11630 12360
rect 11664 12374 11898 12398
rect 11664 12340 11680 12374
rect 11714 12364 11898 12374
rect 11714 12340 11730 12364
rect 11864 12356 11898 12364
rect 11952 12390 12018 12432
rect 11952 12356 11968 12390
rect 12002 12356 12018 12390
rect 12146 12390 12299 12396
rect 12146 12356 12162 12390
rect 12196 12356 12299 12390
rect 11600 12296 11682 12302
rect 11764 12296 11780 12330
rect 11814 12296 11830 12330
rect 11864 12306 11898 12322
rect 11600 12270 11648 12296
rect 11600 12236 11616 12270
rect 11650 12256 11682 12262
rect 11786 12270 11830 12296
rect 12107 12292 12164 12308
rect 11650 12236 11666 12256
rect 11786 12236 12048 12270
rect 11482 12202 11562 12210
rect 11708 12202 11752 12218
rect 11482 12168 11718 12202
rect 11348 12118 11448 12134
rect 11348 12092 11414 12118
rect 11164 12056 11307 12090
rect 11348 12058 11372 12092
rect 11406 12084 11414 12092
rect 11406 12058 11448 12084
rect 10899 11972 10917 12006
rect 10899 11956 10951 11972
rect 10985 11988 11001 12022
rect 11035 11988 11051 12022
rect 9205 11912 9221 11946
rect 9255 11912 9271 11946
rect 10985 11922 11051 11988
rect 11085 12006 11130 12040
rect 11119 11972 11130 12006
rect 11085 11956 11130 11972
rect 11169 11988 11189 12022
rect 11223 11988 11239 12022
rect 11169 11922 11239 11988
rect 11273 12006 11307 12056
rect 11482 11999 11516 12168
rect 11702 12152 11752 12168
rect 11550 12118 11600 12134
rect 11584 12092 11600 12118
rect 11786 12092 11820 12236
rect 11982 12202 11998 12236
rect 12032 12202 12048 12236
rect 12107 12258 12130 12292
rect 12107 12228 12164 12258
rect 11854 12168 11870 12202
rect 11904 12168 11920 12202
rect 12107 12194 12108 12228
rect 12142 12224 12164 12228
rect 12142 12194 12231 12224
rect 12107 12188 12231 12194
rect 11854 12166 11920 12168
rect 11854 12160 12055 12166
rect 11854 12126 12016 12160
rect 12050 12126 12055 12160
rect 11854 12118 12055 12126
rect 12095 12118 12142 12134
rect 11584 12084 11700 12092
rect 11550 12058 11700 12084
rect 11734 12058 11820 12092
rect 12129 12092 12142 12118
rect 11550 12042 11820 12058
rect 11700 12024 11734 12042
rect 11273 11956 11307 11972
rect 11350 11965 11366 11999
rect 11400 11965 11516 11999
rect 11564 11974 11580 12008
rect 11614 11974 11640 12008
rect 11700 11974 11734 11990
rect 11858 12032 11874 12066
rect 11908 12032 11924 12066
rect 12095 12058 12108 12084
rect 12190 12118 12231 12188
rect 12190 12084 12197 12118
rect 12190 12068 12231 12084
rect 12265 12202 12299 12356
rect 12335 12394 12387 12432
rect 12335 12360 12353 12394
rect 12335 12344 12387 12360
rect 12439 12382 12673 12398
rect 12439 12374 12639 12382
rect 12439 12340 12455 12374
rect 12489 12364 12639 12374
rect 12489 12340 12505 12364
rect 12639 12332 12673 12348
rect 12730 12380 12777 12396
rect 12730 12346 12743 12380
rect 12374 12296 12449 12302
rect 12374 12262 12384 12296
rect 12418 12270 12449 12296
rect 12539 12296 12555 12330
rect 12589 12296 12605 12330
rect 12730 12298 12777 12346
rect 12539 12293 12605 12296
rect 12374 12236 12393 12262
rect 12427 12236 12449 12270
rect 12491 12218 12535 12234
rect 12491 12202 12501 12218
rect 12265 12184 12501 12202
rect 12265 12168 12535 12184
rect 12095 12052 12142 12058
rect 11858 11998 11924 12032
rect 12265 11999 12299 12168
rect 12333 12118 12383 12134
rect 12367 12084 12383 12118
rect 12333 12066 12383 12084
rect 12569 12066 12605 12293
rect 12639 12264 12777 12298
rect 12822 12390 12888 12432
rect 12822 12356 12838 12390
rect 12872 12356 12888 12390
rect 12822 12288 12888 12356
rect 12922 12356 12979 12398
rect 12956 12322 12979 12356
rect 12922 12306 12979 12322
rect 12639 12202 12694 12264
rect 12854 12234 12904 12250
rect 12673 12168 12694 12202
rect 12745 12225 12770 12230
rect 12745 12191 12768 12225
rect 12804 12196 12820 12230
rect 12802 12191 12820 12196
rect 12745 12184 12820 12191
rect 12854 12200 12870 12234
rect 12854 12184 12904 12200
rect 12639 12160 12694 12168
rect 12639 12126 12660 12160
rect 12694 12126 12741 12134
rect 12639 12100 12741 12126
rect 12775 12100 12791 12134
rect 12854 12066 12888 12184
rect 12938 12123 12979 12306
rect 12333 12032 12888 12066
rect 12922 12103 12979 12123
rect 12956 12069 12979 12103
rect 12922 12035 12979 12069
rect 11564 11922 11640 11974
rect 11858 11964 11874 11998
rect 11908 11964 11924 11998
rect 12133 11965 12149 11999
rect 12183 11965 12299 11999
rect 12471 12024 12505 12032
rect 11858 11922 11924 11964
rect 12347 11964 12363 11998
rect 12397 11964 12423 11998
rect 12956 12026 12979 12035
rect 12471 11974 12505 11990
rect 12347 11922 12423 11964
rect 12611 11964 12627 11998
rect 12661 11964 12838 11998
rect 12872 11964 12888 11998
rect 12611 11922 12888 11964
rect 12922 11992 12935 12001
rect 12969 11992 12979 12026
rect 12922 11956 12979 11992
rect 13013 12364 13076 12398
rect 13013 12330 13026 12364
rect 13060 12330 13076 12364
rect 13112 12390 13171 12432
rect 13352 12403 13368 12432
rect 13402 12403 13428 12432
rect 13470 12403 13486 12432
rect 13520 12403 13546 12432
rect 13612 12403 13630 12432
rect 13664 12432 13671 12437
rect 13705 12432 13734 12466
rect 14458 12436 14492 12452
rect 13664 12403 13680 12432
rect 13112 12356 13121 12390
rect 13155 12356 13171 12390
rect 13112 12340 13171 12356
rect 13205 12354 13257 12398
rect 14458 12360 14492 12376
rect 14546 12439 14580 12455
rect 14546 12363 14580 12379
rect 15190 12439 15224 12455
rect 15190 12363 15224 12379
rect 15295 12439 15329 12455
rect 15295 12363 15329 12379
rect 15404 12439 15438 12455
rect 15404 12363 15438 12379
rect 16402 12439 16436 12455
rect 16402 12363 16436 12379
rect 16506 12439 16540 12455
rect 16506 12363 16540 12379
rect 16616 12439 16650 12455
rect 16616 12363 16650 12379
rect 17614 12439 17648 12455
rect 17614 12363 17648 12379
rect 17719 12439 17753 12455
rect 17719 12363 17753 12379
rect 17828 12439 17862 12455
rect 17828 12363 17862 12379
rect 18826 12439 18860 12455
rect 18826 12363 18860 12379
rect 18933 12439 18967 12455
rect 18933 12363 18967 12379
rect 19040 12439 19074 12455
rect 19040 12363 19074 12379
rect 19601 12442 19635 12458
rect 19601 12366 19635 12382
rect 19689 12442 19723 12458
rect 19689 12366 19723 12382
rect 19785 12442 19819 12458
rect 19785 12366 19819 12382
rect 19881 12442 19915 12458
rect 19983 12432 20012 12466
rect 20046 12437 20104 12466
rect 20138 12437 20196 12466
rect 20046 12432 20077 12437
rect 20138 12432 20195 12437
rect 20230 12432 20288 12466
rect 20322 12437 20380 12466
rect 20322 12432 20339 12437
rect 20061 12403 20077 12432
rect 20111 12403 20137 12432
rect 20179 12403 20195 12432
rect 20229 12403 20255 12432
rect 20321 12403 20339 12432
rect 20373 12432 20380 12437
rect 20414 12432 20443 12466
rect 21167 12436 21201 12452
rect 20373 12403 20389 12432
rect 19881 12366 19915 12382
rect 21167 12360 21201 12376
rect 21255 12439 21289 12455
rect 21255 12363 21289 12379
rect 21899 12439 21933 12455
rect 21899 12363 21933 12379
rect 22004 12439 22038 12455
rect 22004 12363 22038 12379
rect 22113 12439 22147 12455
rect 22113 12363 22147 12379
rect 23111 12439 23145 12455
rect 23111 12363 23145 12379
rect 23215 12439 23249 12455
rect 23215 12363 23249 12379
rect 23325 12439 23359 12455
rect 23325 12363 23359 12379
rect 24323 12439 24357 12455
rect 24323 12363 24357 12379
rect 24428 12439 24462 12455
rect 24428 12363 24462 12379
rect 24537 12439 24571 12455
rect 24537 12363 24571 12379
rect 25535 12439 25569 12455
rect 25535 12363 25569 12379
rect 25642 12439 25676 12455
rect 25642 12363 25676 12379
rect 25749 12439 25783 12455
rect 25749 12363 25783 12379
rect 26310 12442 26344 12458
rect 26310 12366 26344 12382
rect 26398 12442 26432 12458
rect 26398 12366 26432 12382
rect 26494 12442 26528 12458
rect 26494 12366 26528 12382
rect 26590 12442 26624 12458
rect 26590 12366 26624 12382
rect 13013 12250 13076 12330
rect 13239 12324 13257 12354
rect 13205 12290 13221 12320
rect 13255 12290 13257 12324
rect 19514 12291 19530 12325
rect 19564 12291 19580 12325
rect 13205 12284 13257 12290
rect 19721 12289 19737 12323
rect 19771 12289 19787 12323
rect 26223 12291 26239 12325
rect 26273 12291 26289 12325
rect 26430 12289 26446 12323
rect 26480 12289 26496 12323
rect 13013 12234 13180 12250
rect 13013 12200 13146 12234
rect 13013 12184 13180 12200
rect 13013 12084 13076 12184
rect 13214 12160 13257 12284
rect 14811 12238 14845 12254
rect 14811 12162 14845 12178
rect 14901 12238 14935 12254
rect 14901 12162 14935 12178
rect 15543 12238 15577 12254
rect 15543 12162 15577 12178
rect 15650 12238 15684 12254
rect 15650 12162 15684 12178
rect 15753 12238 15787 12254
rect 15753 12162 15787 12178
rect 16755 12238 16789 12254
rect 16755 12162 16789 12178
rect 16861 12238 16895 12254
rect 16861 12162 16895 12178
rect 16965 12238 16999 12254
rect 16965 12162 16999 12178
rect 18093 12238 18127 12254
rect 18093 12162 18127 12178
rect 18201 12238 18235 12254
rect 18201 12162 18235 12178
rect 18303 12238 18337 12254
rect 18303 12162 18337 12178
rect 18948 12238 18982 12254
rect 18948 12162 18982 12178
rect 19037 12238 19071 12254
rect 19037 12162 19071 12178
rect 19601 12239 19635 12255
rect 19601 12163 19635 12179
rect 19689 12239 19723 12255
rect 19689 12163 19723 12179
rect 19785 12239 19819 12255
rect 19785 12163 19819 12179
rect 19881 12239 19915 12255
rect 19881 12163 19915 12179
rect 21520 12238 21554 12254
rect 21520 12162 21554 12178
rect 21610 12238 21644 12254
rect 21610 12162 21644 12178
rect 22252 12238 22286 12254
rect 22252 12162 22286 12178
rect 22359 12238 22393 12254
rect 22359 12162 22393 12178
rect 22462 12238 22496 12254
rect 22462 12162 22496 12178
rect 23464 12238 23498 12254
rect 23464 12162 23498 12178
rect 23570 12238 23604 12254
rect 23570 12162 23604 12178
rect 23674 12238 23708 12254
rect 23674 12162 23708 12178
rect 24802 12238 24836 12254
rect 24802 12162 24836 12178
rect 24910 12238 24944 12254
rect 24910 12162 24944 12178
rect 25012 12238 25046 12254
rect 25012 12162 25046 12178
rect 25657 12238 25691 12254
rect 25657 12162 25691 12178
rect 25746 12238 25780 12254
rect 25746 12162 25780 12178
rect 26310 12239 26344 12255
rect 26310 12163 26344 12179
rect 26398 12239 26432 12255
rect 26398 12163 26432 12179
rect 26494 12239 26528 12255
rect 26494 12163 26528 12179
rect 26590 12239 26624 12255
rect 26590 12163 26624 12179
rect 13205 12102 13257 12160
rect 13855 12104 13871 12138
rect 13905 12104 13921 12138
rect 13013 12050 13026 12084
rect 13060 12050 13076 12084
rect 13013 12016 13076 12050
rect 13013 11982 13026 12016
rect 13060 11982 13076 12016
rect 13013 11966 13076 11982
rect 13112 12078 13171 12096
rect 13112 12044 13121 12078
rect 13155 12044 13171 12078
rect 13112 12010 13171 12044
rect 13112 11976 13121 12010
rect 13155 11976 13171 12010
rect 13112 11922 13171 11976
rect 13239 12068 13257 12102
rect 14839 12094 14855 12128
rect 14889 12094 14905 12128
rect 15571 12094 15587 12128
rect 15621 12094 15637 12128
rect 15693 12094 15709 12128
rect 15743 12094 15759 12128
rect 16783 12094 16799 12128
rect 16833 12094 16849 12128
rect 16905 12094 16921 12128
rect 16955 12094 16971 12128
rect 18121 12094 18137 12128
rect 18171 12094 18187 12128
rect 18243 12094 18259 12128
rect 18293 12094 18309 12128
rect 18977 12094 18993 12128
rect 19027 12094 19043 12128
rect 19601 12101 19635 12117
rect 13205 12044 13257 12068
rect 13205 12034 13215 12044
rect 13249 12010 13257 12044
rect 13239 12000 13257 12010
rect 13205 11956 13257 12000
rect 13791 12054 13825 12070
rect 13791 11978 13825 11994
rect 13951 12054 13985 12070
rect 19601 12025 19635 12041
rect 19689 12101 19723 12117
rect 20564 12104 20580 12138
rect 20614 12104 20630 12138
rect 21548 12094 21564 12128
rect 21598 12094 21614 12128
rect 22280 12094 22296 12128
rect 22330 12094 22346 12128
rect 22402 12094 22418 12128
rect 22452 12094 22468 12128
rect 23492 12094 23508 12128
rect 23542 12094 23558 12128
rect 23614 12094 23630 12128
rect 23664 12094 23680 12128
rect 24830 12094 24846 12128
rect 24880 12094 24896 12128
rect 24952 12094 24968 12128
rect 25002 12094 25018 12128
rect 25686 12094 25702 12128
rect 25736 12094 25752 12128
rect 26310 12101 26344 12117
rect 19689 12025 19723 12041
rect 20500 12054 20534 12070
rect 13951 11978 13985 11994
rect 20500 11978 20534 11994
rect 20660 12054 20694 12070
rect 26310 12025 26344 12041
rect 26398 12101 26432 12117
rect 26398 12025 26432 12041
rect 20660 11978 20694 11994
rect 9205 11894 9271 11912
rect 9125 11850 9191 11860
rect 8626 11816 8642 11850
rect 8676 11816 8692 11850
rect 8833 11814 8849 11848
rect 8883 11814 8899 11848
rect 9125 11816 9134 11850
rect 9168 11846 9191 11850
rect 9125 11812 9141 11816
rect 9175 11812 9191 11846
rect 9225 11849 9271 11894
rect 10882 11888 10911 11922
rect 10945 11888 11003 11922
rect 11037 11888 11095 11922
rect 11129 11888 11187 11922
rect 11221 11888 11279 11922
rect 11313 11888 11371 11922
rect 11405 11888 11463 11922
rect 9225 11815 9236 11849
rect 9270 11815 9271 11849
rect 10883 11876 11463 11888
rect 10883 11875 11372 11876
rect 10883 11874 11186 11875
rect 10883 11840 10911 11874
rect 10945 11873 11096 11874
rect 10945 11840 11004 11873
rect 10883 11839 11004 11840
rect 11038 11840 11096 11873
rect 11130 11841 11186 11874
rect 11220 11841 11281 11875
rect 11315 11842 11372 11875
rect 11406 11854 11463 11876
rect 11497 11854 11555 11922
rect 11589 11854 11647 11922
rect 11681 11854 11739 11922
rect 11773 11854 11831 11922
rect 11865 11854 11923 11922
rect 11957 11854 12015 11922
rect 12049 11854 12107 11922
rect 12141 11854 12199 11922
rect 12233 11854 12291 11922
rect 12325 11854 12383 11922
rect 12417 11854 12475 11922
rect 12509 11854 12567 11922
rect 12601 11854 12659 11922
rect 12693 11854 12751 11922
rect 12785 11854 12843 11922
rect 12877 11854 12935 11922
rect 12969 11854 13027 11922
rect 13061 11854 13119 11922
rect 13153 11854 13211 11922
rect 13245 11854 13274 11922
rect 11406 11842 13274 11854
rect 11315 11841 13274 11842
rect 11130 11840 13274 11841
rect 13791 11916 13825 11932
rect 13791 11840 13825 11856
rect 13951 11916 13985 11932
rect 13951 11840 13985 11856
rect 20500 11916 20534 11932
rect 20500 11840 20534 11856
rect 20660 11916 20694 11932
rect 20660 11840 20694 11856
rect 11038 11839 13274 11840
rect 10883 11826 13274 11839
rect 3923 11763 3957 11779
rect 3923 11687 3957 11703
rect 4013 11763 4047 11779
rect 4013 11687 4047 11703
rect 4655 11763 4689 11779
rect 4655 11687 4689 11703
rect 4762 11763 4796 11779
rect 4762 11687 4796 11703
rect 4865 11763 4899 11779
rect 4865 11687 4899 11703
rect 5867 11763 5901 11779
rect 5867 11687 5901 11703
rect 5973 11763 6007 11779
rect 5973 11687 6007 11703
rect 6077 11763 6111 11779
rect 6077 11687 6111 11703
rect 7205 11763 7239 11779
rect 7205 11687 7239 11703
rect 7313 11763 7347 11779
rect 7313 11687 7347 11703
rect 7415 11763 7449 11779
rect 7415 11687 7449 11703
rect 8060 11763 8094 11779
rect 8060 11687 8094 11703
rect 8149 11763 8183 11779
rect 8149 11687 8183 11703
rect 8713 11764 8747 11780
rect 8713 11688 8747 11704
rect 8801 11764 8835 11780
rect 8801 11688 8835 11704
rect 8897 11764 8931 11780
rect 8897 11688 8931 11704
rect 8993 11764 9027 11780
rect 8993 11688 9027 11704
rect 9125 11762 9171 11778
rect 9225 11774 9271 11815
rect 10882 11792 10911 11826
rect 10945 11792 11003 11826
rect 11037 11792 11095 11826
rect 11129 11792 11187 11826
rect 11221 11792 11279 11826
rect 11313 11792 11371 11826
rect 11405 11825 13274 11826
rect 11405 11792 11434 11825
rect 9125 11728 9137 11762
rect 9125 11694 9171 11728
rect 2967 11629 2983 11663
rect 3017 11629 3033 11663
rect 9125 11660 9137 11694
rect 3951 11619 3967 11653
rect 4001 11619 4017 11653
rect 4683 11619 4699 11653
rect 4733 11619 4749 11653
rect 4805 11619 4821 11653
rect 4855 11619 4871 11653
rect 5895 11619 5911 11653
rect 5945 11619 5961 11653
rect 6017 11619 6033 11653
rect 6067 11619 6083 11653
rect 7233 11619 7249 11653
rect 7283 11619 7299 11653
rect 7355 11619 7371 11653
rect 7405 11619 7421 11653
rect 8089 11619 8105 11653
rect 8139 11619 8155 11653
rect 8713 11626 8747 11642
rect 2903 11579 2937 11595
rect 2903 11503 2937 11519
rect 3063 11579 3097 11595
rect 8713 11550 8747 11566
rect 8801 11626 8835 11642
rect 9125 11614 9171 11660
rect 9205 11762 9271 11774
rect 9205 11728 9221 11762
rect 9255 11728 9271 11762
rect 9205 11694 9271 11728
rect 9205 11660 9221 11694
rect 9255 11660 9271 11694
rect 9205 11648 9271 11660
rect 10950 11750 10992 11792
rect 10950 11716 10958 11750
rect 10950 11682 10992 11716
rect 10950 11648 10958 11682
rect 10950 11614 10992 11648
rect 8801 11550 8835 11566
rect 9061 11580 9090 11614
rect 9124 11580 9182 11614
rect 9216 11580 9274 11614
rect 9308 11580 9337 11614
rect 10950 11580 10958 11614
rect 9061 11572 9336 11580
rect 9061 11538 9091 11572
rect 9125 11538 9183 11572
rect 9217 11570 9336 11572
rect 9217 11538 9277 11570
rect 9061 11536 9277 11538
rect 9311 11536 9336 11570
rect 10950 11564 10992 11580
rect 11026 11750 11092 11758
rect 11026 11716 11042 11750
rect 11076 11716 11092 11750
rect 11026 11682 11092 11716
rect 11026 11648 11042 11682
rect 11076 11651 11092 11682
rect 11026 11617 11044 11648
rect 11078 11617 11092 11651
rect 11026 11614 11092 11617
rect 11026 11580 11042 11614
rect 11076 11580 11092 11614
rect 11026 11562 11092 11580
rect 11226 11750 11268 11792
rect 13791 11778 13825 11794
rect 11226 11716 11234 11750
rect 11226 11682 11268 11716
rect 11226 11648 11234 11682
rect 11226 11614 11268 11648
rect 11226 11580 11234 11614
rect 11226 11564 11268 11580
rect 11302 11750 11368 11758
rect 11302 11716 11318 11750
rect 11352 11727 11368 11750
rect 11302 11693 11319 11716
rect 11353 11693 11368 11727
rect 13791 11702 13825 11718
rect 13951 11778 13985 11794
rect 13951 11702 13985 11718
rect 20500 11778 20534 11794
rect 20500 11702 20534 11718
rect 20660 11778 20694 11794
rect 20660 11702 20694 11718
rect 11302 11682 11368 11693
rect 11302 11648 11318 11682
rect 11352 11648 11368 11682
rect 11302 11614 11368 11648
rect 13791 11640 13825 11656
rect 11302 11580 11318 11614
rect 11352 11580 11368 11614
rect 11302 11562 11368 11580
rect 9061 11531 9336 11536
rect 3063 11503 3097 11519
rect 10946 11522 11012 11528
rect 10946 11488 10957 11522
rect 10991 11514 11012 11522
rect 10946 11480 10962 11488
rect 10996 11480 11012 11514
rect 2903 11441 2937 11457
rect 2903 11365 2937 11381
rect 3063 11441 3097 11457
rect 3063 11365 3097 11381
rect 10946 11430 10992 11446
rect 11046 11442 11092 11562
rect 11222 11517 11288 11528
rect 11222 11483 11228 11517
rect 11262 11514 11288 11517
rect 11222 11480 11238 11483
rect 11272 11480 11288 11514
rect 10946 11396 10958 11430
rect 10946 11362 10992 11396
rect 10946 11328 10958 11362
rect 2903 11303 2937 11319
rect 2903 11227 2937 11243
rect 3063 11303 3097 11319
rect 10946 11282 10992 11328
rect 11026 11430 11092 11442
rect 11026 11396 11042 11430
rect 11076 11396 11092 11430
rect 11026 11362 11092 11396
rect 11026 11328 11042 11362
rect 11076 11328 11092 11362
rect 11026 11316 11092 11328
rect 11222 11430 11268 11446
rect 11322 11442 11368 11562
rect 13289 11596 13407 11615
rect 13289 11539 13315 11596
rect 13381 11539 13407 11596
rect 13791 11564 13825 11580
rect 13951 11640 13985 11656
rect 13951 11564 13985 11580
rect 20500 11640 20534 11656
rect 20500 11564 20534 11580
rect 20660 11640 20694 11656
rect 20660 11564 20694 11580
rect 13289 11516 13407 11539
rect 11222 11396 11234 11430
rect 11222 11362 11268 11396
rect 11222 11328 11234 11362
rect 11222 11282 11268 11328
rect 11302 11430 11368 11442
rect 11302 11396 11318 11430
rect 11352 11396 11368 11430
rect 13791 11502 13825 11518
rect 13791 11426 13825 11442
rect 13951 11502 13985 11518
rect 13951 11426 13985 11442
rect 20500 11502 20534 11518
rect 20500 11426 20534 11442
rect 20660 11502 20694 11518
rect 20660 11426 20694 11442
rect 11302 11362 11368 11396
rect 11302 11328 11318 11362
rect 11352 11328 11368 11362
rect 11302 11316 11368 11328
rect 13791 11364 13825 11380
rect 13791 11288 13825 11304
rect 13951 11364 13985 11380
rect 13951 11288 13985 11304
rect 20500 11364 20534 11380
rect 20500 11288 20534 11304
rect 20660 11364 20694 11380
rect 20660 11288 20694 11304
rect 3063 11227 3097 11243
rect 10882 11214 10911 11282
rect 10945 11214 11003 11282
rect 11037 11214 11095 11282
rect 11129 11214 11187 11282
rect 11221 11214 11279 11282
rect 11313 11214 11371 11282
rect 11405 11214 11434 11282
rect 13791 11226 13825 11242
rect 2903 11165 2937 11181
rect 2903 11089 2937 11105
rect 3063 11165 3097 11181
rect 13791 11150 13825 11166
rect 13951 11226 13985 11242
rect 13951 11150 13985 11166
rect 14067 11212 14172 11247
rect 14067 11178 14099 11212
rect 14133 11178 14172 11212
rect 14067 11149 14172 11178
rect 20500 11226 20534 11242
rect 20500 11150 20534 11166
rect 20660 11226 20694 11242
rect 20660 11150 20694 11166
rect 20776 11212 20881 11247
rect 20776 11178 20808 11212
rect 20842 11178 20881 11212
rect 20776 11149 20881 11178
rect 3063 11089 3097 11105
rect 13791 11088 13825 11104
rect 2903 11027 2937 11043
rect 2903 10951 2937 10967
rect 3063 11027 3097 11043
rect 13791 11012 13825 11028
rect 13951 11094 13985 11104
rect 14081 11094 14158 11149
rect 13951 11088 14158 11094
rect 13985 11028 14158 11088
rect 20500 11088 20534 11104
rect 13951 11025 14158 11028
rect 14466 11041 14798 11057
rect 13951 11012 13985 11025
rect 14466 11007 14492 11041
rect 14526 11007 14572 11041
rect 14606 11007 14652 11041
rect 14686 11007 14732 11041
rect 14766 11007 14798 11041
rect 14466 10989 14798 11007
rect 15198 11041 15530 11057
rect 15198 11007 15224 11041
rect 15258 11007 15304 11041
rect 15338 11007 15384 11041
rect 15418 11007 15464 11041
rect 15498 11007 15530 11041
rect 15198 10989 15530 11007
rect 15800 11041 16132 11057
rect 15800 11007 15832 11041
rect 15866 11007 15912 11041
rect 15946 11007 15992 11041
rect 16026 11007 16072 11041
rect 16106 11007 16132 11041
rect 15800 10989 16132 11007
rect 16410 11041 16742 11057
rect 16410 11007 16436 11041
rect 16470 11007 16516 11041
rect 16550 11007 16596 11041
rect 16630 11007 16676 11041
rect 16710 11007 16742 11041
rect 16410 10989 16742 11007
rect 17012 11041 17344 11057
rect 17012 11007 17044 11041
rect 17078 11007 17124 11041
rect 17158 11007 17204 11041
rect 17238 11007 17284 11041
rect 17318 11007 17344 11041
rect 17012 10989 17344 11007
rect 17748 11041 18080 11057
rect 17748 11007 17774 11041
rect 17808 11007 17854 11041
rect 17888 11007 17934 11041
rect 17968 11007 18014 11041
rect 18048 11007 18080 11041
rect 17748 10989 18080 11007
rect 18350 11041 18682 11057
rect 18350 11007 18382 11041
rect 18416 11007 18462 11041
rect 18496 11007 18542 11041
rect 18576 11007 18622 11041
rect 18656 11007 18682 11041
rect 18350 10989 18682 11007
rect 19084 11041 19416 11057
rect 19084 11007 19116 11041
rect 19150 11007 19196 11041
rect 19230 11007 19276 11041
rect 19310 11007 19356 11041
rect 19390 11007 19416 11041
rect 20500 11012 20534 11028
rect 20660 11094 20694 11104
rect 20790 11094 20867 11149
rect 20660 11088 20867 11094
rect 20694 11028 20867 11088
rect 20660 11025 20867 11028
rect 21175 11041 21507 11057
rect 20660 11012 20694 11025
rect 19084 10989 19416 11007
rect 21175 11007 21201 11041
rect 21235 11007 21281 11041
rect 21315 11007 21361 11041
rect 21395 11007 21441 11041
rect 21475 11007 21507 11041
rect 21175 10989 21507 11007
rect 21907 11041 22239 11057
rect 21907 11007 21933 11041
rect 21967 11007 22013 11041
rect 22047 11007 22093 11041
rect 22127 11007 22173 11041
rect 22207 11007 22239 11041
rect 21907 10989 22239 11007
rect 22509 11041 22841 11057
rect 22509 11007 22541 11041
rect 22575 11007 22621 11041
rect 22655 11007 22701 11041
rect 22735 11007 22781 11041
rect 22815 11007 22841 11041
rect 22509 10989 22841 11007
rect 23119 11041 23451 11057
rect 23119 11007 23145 11041
rect 23179 11007 23225 11041
rect 23259 11007 23305 11041
rect 23339 11007 23385 11041
rect 23419 11007 23451 11041
rect 23119 10989 23451 11007
rect 23721 11041 24053 11057
rect 23721 11007 23753 11041
rect 23787 11007 23833 11041
rect 23867 11007 23913 11041
rect 23947 11007 23993 11041
rect 24027 11007 24053 11041
rect 23721 10989 24053 11007
rect 24457 11041 24789 11057
rect 24457 11007 24483 11041
rect 24517 11007 24563 11041
rect 24597 11007 24643 11041
rect 24677 11007 24723 11041
rect 24757 11007 24789 11041
rect 24457 10989 24789 11007
rect 25059 11041 25391 11057
rect 25059 11007 25091 11041
rect 25125 11007 25171 11041
rect 25205 11007 25251 11041
rect 25285 11007 25331 11041
rect 25365 11007 25391 11041
rect 25059 10989 25391 11007
rect 25793 11041 26125 11057
rect 25793 11007 25825 11041
rect 25859 11007 25905 11041
rect 25939 11007 25985 11041
rect 26019 11007 26065 11041
rect 26099 11007 26125 11041
rect 25793 10989 26125 11007
rect 3063 10951 3097 10967
rect 2903 10889 2937 10905
rect 2903 10813 2937 10829
rect 3063 10889 3097 10905
rect 3063 10813 3097 10829
rect 2903 10751 2937 10767
rect 2903 10675 2937 10691
rect 3063 10751 3097 10767
rect 3063 10675 3097 10691
rect 3179 10737 3284 10772
rect 3179 10703 3211 10737
rect 3245 10703 3284 10737
rect 3179 10674 3284 10703
rect 2903 10613 2937 10629
rect 2903 10537 2937 10553
rect 3063 10619 3097 10629
rect 3193 10619 3270 10674
rect 3063 10613 3270 10619
rect 3097 10553 3270 10613
rect 3063 10550 3270 10553
rect 3578 10566 3910 10582
rect 3063 10537 3097 10550
rect 3578 10532 3604 10566
rect 3638 10532 3684 10566
rect 3718 10532 3764 10566
rect 3798 10532 3844 10566
rect 3878 10532 3910 10566
rect 3578 10514 3910 10532
rect 4310 10566 4642 10582
rect 4310 10532 4336 10566
rect 4370 10532 4416 10566
rect 4450 10532 4496 10566
rect 4530 10532 4576 10566
rect 4610 10532 4642 10566
rect 4310 10514 4642 10532
rect 4912 10566 5244 10582
rect 4912 10532 4944 10566
rect 4978 10532 5024 10566
rect 5058 10532 5104 10566
rect 5138 10532 5184 10566
rect 5218 10532 5244 10566
rect 4912 10514 5244 10532
rect 5522 10566 5854 10582
rect 5522 10532 5548 10566
rect 5582 10532 5628 10566
rect 5662 10532 5708 10566
rect 5742 10532 5788 10566
rect 5822 10532 5854 10566
rect 5522 10514 5854 10532
rect 6124 10566 6456 10582
rect 6124 10532 6156 10566
rect 6190 10532 6236 10566
rect 6270 10532 6316 10566
rect 6350 10532 6396 10566
rect 6430 10532 6456 10566
rect 6124 10514 6456 10532
rect 6860 10566 7192 10582
rect 6860 10532 6886 10566
rect 6920 10532 6966 10566
rect 7000 10532 7046 10566
rect 7080 10532 7126 10566
rect 7160 10532 7192 10566
rect 6860 10514 7192 10532
rect 7462 10566 7794 10582
rect 7462 10532 7494 10566
rect 7528 10532 7574 10566
rect 7608 10532 7654 10566
rect 7688 10532 7734 10566
rect 7768 10532 7794 10566
rect 7462 10514 7794 10532
rect 8196 10566 8528 10582
rect 8196 10532 8228 10566
rect 8262 10532 8308 10566
rect 8342 10532 8388 10566
rect 8422 10532 8468 10566
rect 8502 10532 8528 10566
rect 8196 10514 8528 10532
rect 3578 10114 3910 10132
rect 2903 10093 2937 10109
rect 2903 10017 2937 10033
rect 3063 10096 3097 10109
rect 3063 10093 3270 10096
rect 3097 10033 3270 10093
rect 3578 10080 3604 10114
rect 3638 10080 3684 10114
rect 3718 10080 3764 10114
rect 3798 10080 3844 10114
rect 3878 10080 3910 10114
rect 3578 10064 3910 10080
rect 4310 10114 4642 10132
rect 4310 10080 4336 10114
rect 4370 10080 4416 10114
rect 4450 10080 4496 10114
rect 4530 10080 4576 10114
rect 4610 10080 4642 10114
rect 4310 10064 4642 10080
rect 4912 10114 5244 10132
rect 4912 10080 4944 10114
rect 4978 10080 5024 10114
rect 5058 10080 5104 10114
rect 5138 10080 5184 10114
rect 5218 10080 5244 10114
rect 4912 10064 5244 10080
rect 5522 10114 5854 10132
rect 5522 10080 5548 10114
rect 5582 10080 5628 10114
rect 5662 10080 5708 10114
rect 5742 10080 5788 10114
rect 5822 10080 5854 10114
rect 5522 10064 5854 10080
rect 6124 10114 6456 10132
rect 6124 10080 6156 10114
rect 6190 10080 6236 10114
rect 6270 10080 6316 10114
rect 6350 10080 6396 10114
rect 6430 10080 6456 10114
rect 6124 10064 6456 10080
rect 6860 10114 7192 10132
rect 6860 10080 6886 10114
rect 6920 10080 6966 10114
rect 7000 10080 7046 10114
rect 7080 10080 7126 10114
rect 7160 10080 7192 10114
rect 6860 10064 7192 10080
rect 7462 10114 7794 10132
rect 7462 10080 7494 10114
rect 7528 10080 7574 10114
rect 7608 10080 7654 10114
rect 7688 10080 7734 10114
rect 7768 10080 7794 10114
rect 7462 10064 7794 10080
rect 8196 10114 8528 10132
rect 8196 10080 8228 10114
rect 8262 10080 8308 10114
rect 8342 10080 8388 10114
rect 8422 10080 8468 10114
rect 8502 10080 8528 10114
rect 8196 10064 8528 10080
rect 13763 10102 14095 10120
rect 13763 10068 13789 10102
rect 13823 10068 13869 10102
rect 13903 10068 13949 10102
rect 13983 10068 14029 10102
rect 14063 10068 14095 10102
rect 13763 10052 14095 10068
rect 14497 10102 14829 10120
rect 14497 10068 14523 10102
rect 14557 10068 14603 10102
rect 14637 10068 14683 10102
rect 14717 10068 14763 10102
rect 14797 10068 14829 10102
rect 14497 10052 14829 10068
rect 15099 10102 15431 10120
rect 15099 10068 15131 10102
rect 15165 10068 15211 10102
rect 15245 10068 15291 10102
rect 15325 10068 15371 10102
rect 15405 10068 15431 10102
rect 15099 10052 15431 10068
rect 15835 10102 16167 10120
rect 15835 10068 15861 10102
rect 15895 10068 15941 10102
rect 15975 10068 16021 10102
rect 16055 10068 16101 10102
rect 16135 10068 16167 10102
rect 15835 10052 16167 10068
rect 16437 10102 16769 10120
rect 16437 10068 16469 10102
rect 16503 10068 16549 10102
rect 16583 10068 16629 10102
rect 16663 10068 16709 10102
rect 16743 10068 16769 10102
rect 16437 10052 16769 10068
rect 17047 10102 17379 10120
rect 17047 10068 17073 10102
rect 17107 10068 17153 10102
rect 17187 10068 17233 10102
rect 17267 10068 17313 10102
rect 17347 10068 17379 10102
rect 17047 10052 17379 10068
rect 17649 10102 17981 10120
rect 17649 10068 17681 10102
rect 17715 10068 17761 10102
rect 17795 10068 17841 10102
rect 17875 10068 17921 10102
rect 17955 10068 17981 10102
rect 17649 10052 17981 10068
rect 18381 10102 18713 10120
rect 18381 10068 18413 10102
rect 18447 10068 18493 10102
rect 18527 10068 18573 10102
rect 18607 10068 18653 10102
rect 18687 10068 18713 10102
rect 20472 10102 20804 10120
rect 19194 10084 19228 10097
rect 18381 10052 18713 10068
rect 19021 10081 19228 10084
rect 3063 10027 3270 10033
rect 3063 10017 3097 10027
rect 3193 9972 3270 10027
rect 19021 10021 19194 10081
rect 19021 10015 19228 10021
rect 2903 9955 2937 9971
rect 2903 9879 2937 9895
rect 3063 9955 3097 9971
rect 3063 9879 3097 9895
rect 3179 9943 3284 9972
rect 19021 9960 19098 10015
rect 19194 10005 19228 10015
rect 19354 10081 19388 10097
rect 20472 10068 20498 10102
rect 20532 10068 20578 10102
rect 20612 10068 20658 10102
rect 20692 10068 20738 10102
rect 20772 10068 20804 10102
rect 20472 10052 20804 10068
rect 21206 10102 21538 10120
rect 21206 10068 21232 10102
rect 21266 10068 21312 10102
rect 21346 10068 21392 10102
rect 21426 10068 21472 10102
rect 21506 10068 21538 10102
rect 21206 10052 21538 10068
rect 21808 10102 22140 10120
rect 21808 10068 21840 10102
rect 21874 10068 21920 10102
rect 21954 10068 22000 10102
rect 22034 10068 22080 10102
rect 22114 10068 22140 10102
rect 21808 10052 22140 10068
rect 22544 10102 22876 10120
rect 22544 10068 22570 10102
rect 22604 10068 22650 10102
rect 22684 10068 22730 10102
rect 22764 10068 22810 10102
rect 22844 10068 22876 10102
rect 22544 10052 22876 10068
rect 23146 10102 23478 10120
rect 23146 10068 23178 10102
rect 23212 10068 23258 10102
rect 23292 10068 23338 10102
rect 23372 10068 23418 10102
rect 23452 10068 23478 10102
rect 23146 10052 23478 10068
rect 23756 10102 24088 10120
rect 23756 10068 23782 10102
rect 23816 10068 23862 10102
rect 23896 10068 23942 10102
rect 23976 10068 24022 10102
rect 24056 10068 24088 10102
rect 23756 10052 24088 10068
rect 24358 10102 24690 10120
rect 24358 10068 24390 10102
rect 24424 10068 24470 10102
rect 24504 10068 24550 10102
rect 24584 10068 24630 10102
rect 24664 10068 24690 10102
rect 24358 10052 24690 10068
rect 25090 10102 25422 10120
rect 25090 10068 25122 10102
rect 25156 10068 25202 10102
rect 25236 10068 25282 10102
rect 25316 10068 25362 10102
rect 25396 10068 25422 10102
rect 25903 10084 25937 10097
rect 25090 10052 25422 10068
rect 25730 10081 25937 10084
rect 19354 10005 19388 10021
rect 25730 10021 25903 10081
rect 25730 10015 25937 10021
rect 25730 9960 25807 10015
rect 25903 10005 25937 10015
rect 26063 10081 26097 10097
rect 26063 10005 26097 10021
rect 3179 9909 3211 9943
rect 3245 9909 3284 9943
rect 3179 9874 3284 9909
rect 19007 9931 19112 9960
rect 19007 9897 19046 9931
rect 19080 9897 19112 9931
rect 19007 9862 19112 9897
rect 19194 9943 19228 9959
rect 19194 9867 19228 9883
rect 19354 9943 19388 9959
rect 19354 9867 19388 9883
rect 25716 9931 25821 9960
rect 25716 9897 25755 9931
rect 25789 9897 25821 9931
rect 25716 9862 25821 9897
rect 25903 9943 25937 9959
rect 25903 9867 25937 9883
rect 26063 9943 26097 9959
rect 26063 9867 26097 9883
rect 2903 9817 2937 9833
rect 2903 9741 2937 9757
rect 3063 9817 3097 9833
rect 3063 9741 3097 9757
rect 19194 9805 19228 9821
rect 19194 9729 19228 9745
rect 19354 9805 19388 9821
rect 19354 9729 19388 9745
rect 25903 9805 25937 9821
rect 25903 9729 25937 9745
rect 26063 9805 26097 9821
rect 26063 9729 26097 9745
rect 2903 9679 2937 9695
rect 2903 9603 2937 9619
rect 3063 9679 3097 9695
rect 3063 9603 3097 9619
rect 19194 9667 19228 9683
rect 19194 9591 19228 9607
rect 19354 9667 19388 9683
rect 19354 9591 19388 9607
rect 25903 9667 25937 9683
rect 25903 9591 25937 9607
rect 26063 9667 26097 9683
rect 26063 9591 26097 9607
rect 2903 9541 2937 9557
rect 2903 9465 2937 9481
rect 3063 9541 3097 9557
rect 3063 9465 3097 9481
rect 19194 9529 19228 9545
rect 19194 9453 19228 9469
rect 19354 9529 19388 9545
rect 19354 9453 19388 9469
rect 25903 9529 25937 9545
rect 25903 9453 25937 9469
rect 26063 9529 26097 9545
rect 26063 9453 26097 9469
rect 2903 9403 2937 9419
rect 2903 9327 2937 9343
rect 3063 9403 3097 9419
rect 3063 9327 3097 9343
rect 19194 9391 19228 9407
rect 19194 9315 19228 9331
rect 19354 9391 19388 9407
rect 19354 9315 19388 9331
rect 25903 9391 25937 9407
rect 25903 9315 25937 9331
rect 26063 9391 26097 9407
rect 26063 9315 26097 9331
rect 2903 9265 2937 9281
rect 2903 9189 2937 9205
rect 3063 9265 3097 9281
rect 3063 9189 3097 9205
rect 19194 9253 19228 9269
rect 19194 9177 19228 9193
rect 19354 9253 19388 9269
rect 19354 9177 19388 9193
rect 25903 9253 25937 9269
rect 25903 9177 25937 9193
rect 26063 9253 26097 9269
rect 26063 9177 26097 9193
rect 2903 9127 2937 9143
rect 2903 9051 2937 9067
rect 3063 9127 3097 9143
rect 19194 9115 19228 9131
rect 9061 9103 11710 9106
rect 9061 9102 9898 9103
rect 3063 9051 3097 9067
rect 8713 9080 8747 9096
rect 2967 8983 2983 9017
rect 3017 8983 3033 9017
rect 3951 8993 3967 9027
rect 4001 8993 4017 9027
rect 4683 8993 4699 9027
rect 4733 8993 4749 9027
rect 4805 8993 4821 9027
rect 4855 8993 4871 9027
rect 5895 8993 5911 9027
rect 5945 8993 5961 9027
rect 6017 8993 6033 9027
rect 6067 8993 6083 9027
rect 7233 8993 7249 9027
rect 7283 8993 7299 9027
rect 7355 8993 7371 9027
rect 7405 8993 7421 9027
rect 8089 8993 8105 9027
rect 8139 8993 8155 9027
rect 8713 9004 8747 9020
rect 8801 9080 8835 9096
rect 9061 9034 9090 9102
rect 9124 9034 9182 9102
rect 9216 9034 9274 9102
rect 9308 9034 9346 9102
rect 9380 9101 9530 9102
rect 9380 9034 9438 9101
rect 9472 9034 9530 9101
rect 9564 9068 9714 9102
rect 9564 9034 9622 9068
rect 9656 9034 9714 9068
rect 9748 9034 9806 9102
rect 9840 9069 9898 9102
rect 9932 9102 11710 9103
rect 9932 9069 9990 9102
rect 9840 9068 9990 9069
rect 10024 9101 10174 9102
rect 9840 9034 9898 9068
rect 9932 9034 9990 9068
rect 10024 9034 10082 9101
rect 10116 9034 10174 9101
rect 10208 9034 10266 9102
rect 10300 9034 10358 9102
rect 10392 9034 10450 9102
rect 10484 9034 10542 9102
rect 10576 9034 10634 9102
rect 10668 9034 10726 9102
rect 10760 9034 10818 9102
rect 10852 9101 11002 9102
rect 10852 9034 10910 9101
rect 10944 9034 11002 9101
rect 11036 9034 11094 9102
rect 11128 9068 11278 9102
rect 11128 9034 11186 9068
rect 11220 9034 11278 9068
rect 11312 9034 11370 9102
rect 11404 9034 11462 9102
rect 11496 9034 11554 9102
rect 11588 9101 11710 9102
rect 11588 9034 11646 9101
rect 11680 9067 11710 9101
rect 11680 9034 11709 9067
rect 12117 9052 12557 9088
rect 13456 9068 13490 9084
rect 8801 9004 8835 9020
rect 9125 8988 9171 9034
rect 3923 8943 3957 8959
rect 3923 8867 3957 8883
rect 4013 8943 4047 8959
rect 4013 8867 4047 8883
rect 4655 8943 4689 8959
rect 4655 8867 4689 8883
rect 4762 8943 4796 8959
rect 4762 8867 4796 8883
rect 4865 8943 4899 8959
rect 4865 8867 4899 8883
rect 5867 8943 5901 8959
rect 5867 8867 5901 8883
rect 5973 8943 6007 8959
rect 5973 8867 6007 8883
rect 6077 8943 6111 8959
rect 6077 8867 6111 8883
rect 7205 8943 7239 8959
rect 7205 8867 7239 8883
rect 7313 8943 7347 8959
rect 7313 8867 7347 8883
rect 7415 8943 7449 8959
rect 7415 8867 7449 8883
rect 8060 8943 8094 8959
rect 8060 8867 8094 8883
rect 8149 8943 8183 8959
rect 8149 8867 8183 8883
rect 8713 8942 8747 8958
rect 8713 8866 8747 8882
rect 8801 8942 8835 8958
rect 8801 8866 8835 8882
rect 8897 8942 8931 8958
rect 8897 8866 8931 8882
rect 8993 8942 9027 8958
rect 8993 8866 9027 8882
rect 9125 8954 9137 8988
rect 9125 8920 9171 8954
rect 9125 8886 9137 8920
rect 9125 8870 9171 8886
rect 9205 8988 9271 9000
rect 9205 8954 9221 8988
rect 9255 8954 9271 8988
rect 9205 8920 9271 8954
rect 9205 8886 9221 8920
rect 9255 8886 9271 8920
rect 9205 8874 9271 8886
rect 9125 8833 9141 8836
rect 8626 8796 8642 8830
rect 8676 8796 8692 8830
rect 8833 8798 8849 8832
rect 8883 8798 8899 8832
rect 9125 8799 9136 8833
rect 9175 8802 9191 8836
rect 9170 8799 9191 8802
rect 9125 8788 9191 8799
rect 9225 8828 9271 8874
rect 9225 8794 9236 8828
rect 9270 8794 9271 8828
rect 3570 8745 3604 8761
rect 2464 8689 2480 8718
rect 2514 8689 2540 8718
rect 2582 8689 2598 8718
rect 2632 8689 2658 8718
rect 2724 8689 2742 8718
rect 2386 8655 2415 8689
rect 2449 8684 2480 8689
rect 2541 8684 2598 8689
rect 2449 8655 2507 8684
rect 2541 8655 2599 8684
rect 2633 8655 2691 8689
rect 2725 8684 2742 8689
rect 2776 8689 2792 8718
rect 2776 8684 2783 8689
rect 2725 8655 2783 8684
rect 2817 8655 2846 8689
rect 3570 8669 3604 8685
rect 3658 8742 3692 8758
rect 3658 8666 3692 8682
rect 4302 8742 4336 8758
rect 4302 8666 4336 8682
rect 4407 8742 4441 8758
rect 4407 8666 4441 8682
rect 4516 8742 4550 8758
rect 4516 8666 4550 8682
rect 5514 8742 5548 8758
rect 5514 8666 5548 8682
rect 5618 8742 5652 8758
rect 5618 8666 5652 8682
rect 5728 8742 5762 8758
rect 5728 8666 5762 8682
rect 6726 8742 6760 8758
rect 6726 8666 6760 8682
rect 6831 8742 6865 8758
rect 6831 8666 6865 8682
rect 6940 8742 6974 8758
rect 6940 8666 6974 8682
rect 7938 8742 7972 8758
rect 7938 8666 7972 8682
rect 8045 8742 8079 8758
rect 8045 8666 8079 8682
rect 8152 8742 8186 8758
rect 8152 8666 8186 8682
rect 8713 8739 8747 8755
rect 8713 8663 8747 8679
rect 8801 8739 8835 8755
rect 8801 8663 8835 8679
rect 8897 8739 8931 8755
rect 8897 8663 8931 8679
rect 8993 8739 9027 8755
rect 9225 8754 9271 8794
rect 8993 8663 9027 8679
rect 9129 8736 9171 8752
rect 9129 8702 9137 8736
rect 9129 8668 9171 8702
rect 2450 8609 2496 8655
rect 2450 8575 2462 8609
rect 2450 8541 2496 8575
rect 2450 8507 2462 8541
rect 2450 8491 2496 8507
rect 2530 8609 2596 8621
rect 2530 8575 2546 8609
rect 2580 8575 2596 8609
rect 2530 8541 2596 8575
rect 2530 8507 2546 8541
rect 2580 8507 2596 8541
rect 2530 8495 2596 8507
rect 2450 8453 2466 8457
rect 2450 8419 2462 8453
rect 2500 8423 2516 8457
rect 2496 8419 2516 8423
rect 2450 8409 2516 8419
rect 2550 8375 2596 8495
rect 2454 8357 2496 8373
rect 2454 8323 2462 8357
rect 2454 8289 2496 8323
rect 2454 8255 2462 8289
rect 2454 8221 2496 8255
rect 2454 8187 2462 8221
rect 2454 8145 2496 8187
rect 2530 8357 2596 8375
rect 2530 8323 2546 8357
rect 2580 8323 2596 8357
rect 2530 8289 2596 8323
rect 2530 8288 2546 8289
rect 2530 8254 2543 8288
rect 2580 8255 2596 8289
rect 2577 8254 2596 8255
rect 2530 8221 2596 8254
rect 2530 8187 2546 8221
rect 2580 8187 2596 8221
rect 2530 8179 2596 8187
rect 2636 8609 2702 8621
rect 2636 8575 2652 8609
rect 2686 8575 2702 8609
rect 2636 8541 2702 8575
rect 2636 8507 2652 8541
rect 2686 8507 2702 8541
rect 2636 8495 2702 8507
rect 2736 8609 2782 8655
rect 9129 8634 9137 8668
rect 3164 8622 3213 8634
rect 2770 8575 2782 8609
rect 2736 8541 2782 8575
rect 3073 8621 3213 8622
rect 3073 8588 3173 8621
rect 2770 8507 2782 8541
rect 2636 8375 2682 8495
rect 2736 8491 2782 8507
rect 2904 8546 2953 8559
rect 3073 8546 3114 8588
rect 3164 8587 3173 8588
rect 3207 8587 3213 8621
rect 3598 8592 3614 8626
rect 3648 8592 3664 8626
rect 4330 8589 4346 8623
rect 4380 8589 4396 8623
rect 4456 8589 4472 8623
rect 4506 8589 4522 8623
rect 5542 8589 5558 8623
rect 5592 8589 5608 8623
rect 5668 8589 5684 8623
rect 5718 8589 5734 8623
rect 6754 8589 6770 8623
rect 6804 8589 6820 8623
rect 6880 8589 6896 8623
rect 6930 8589 6946 8623
rect 7966 8589 7982 8623
rect 8016 8589 8032 8623
rect 8092 8589 8108 8623
rect 8142 8589 8158 8623
rect 8713 8601 8747 8617
rect 3164 8575 3213 8587
rect 2904 8512 2913 8546
rect 2947 8512 3114 8546
rect 3163 8528 3212 8541
rect 2904 8500 2953 8512
rect 3163 8494 3172 8528
rect 3206 8494 3212 8528
rect 8713 8525 8747 8541
rect 8801 8601 8835 8617
rect 8801 8525 8835 8541
rect 9129 8600 9171 8634
rect 9129 8566 9137 8600
rect 9129 8524 9171 8566
rect 9205 8736 9271 8754
rect 9205 8702 9221 8736
rect 9255 8702 9271 8736
rect 9205 8668 9271 8702
rect 9205 8634 9221 8668
rect 9255 8634 9271 8668
rect 9205 8600 9271 8634
rect 9205 8566 9221 8600
rect 9255 8566 9271 8600
rect 9205 8558 9271 8566
rect 9334 8956 9386 9000
rect 9334 8922 9352 8956
rect 9420 8992 9479 9034
rect 9420 8958 9436 8992
rect 9470 8958 9479 8992
rect 9420 8942 9479 8958
rect 9515 8966 9578 9000
rect 9334 8886 9386 8922
rect 9515 8932 9531 8966
rect 9565 8932 9578 8966
rect 9334 8762 9377 8886
rect 9515 8852 9578 8932
rect 9411 8836 9578 8852
rect 9445 8802 9578 8836
rect 9411 8786 9578 8802
rect 9334 8704 9386 8762
rect 9334 8670 9352 8704
rect 9334 8636 9386 8670
rect 9334 8635 9352 8636
rect 9334 8601 9343 8635
rect 9377 8601 9386 8602
rect 9334 8558 9386 8601
rect 9420 8680 9479 8698
rect 9420 8646 9436 8680
rect 9470 8646 9479 8680
rect 9420 8612 9479 8646
rect 9420 8578 9436 8612
rect 9470 8578 9479 8612
rect 9420 8524 9479 8578
rect 9515 8686 9578 8786
rect 9515 8652 9531 8686
rect 9565 8652 9578 8686
rect 9515 8618 9578 8652
rect 9515 8584 9531 8618
rect 9565 8584 9578 8618
rect 9515 8568 9578 8584
rect 9612 8958 9669 9000
rect 9612 8924 9635 8958
rect 9612 8908 9669 8924
rect 9703 8992 9769 9034
rect 9703 8958 9719 8992
rect 9753 8958 9769 8992
rect 9612 8725 9653 8908
rect 9703 8890 9769 8958
rect 9814 8982 9861 8998
rect 9848 8948 9861 8982
rect 9814 8900 9861 8948
rect 9918 8984 10152 9000
rect 9952 8976 10152 8984
rect 9952 8966 10102 8976
rect 9918 8934 9952 8950
rect 10086 8942 10102 8966
rect 10136 8942 10152 8976
rect 10204 8996 10256 9034
rect 10238 8962 10256 8996
rect 10204 8946 10256 8962
rect 10292 8992 10445 8998
rect 10292 8958 10395 8992
rect 10429 8958 10445 8992
rect 10573 8992 10639 9034
rect 10573 8958 10589 8992
rect 10623 8958 10639 8992
rect 10693 8976 10927 9000
rect 10693 8966 10877 8976
rect 10693 8958 10727 8966
rect 9814 8866 9952 8900
rect 9687 8836 9737 8852
rect 9721 8802 9737 8836
rect 9687 8786 9737 8802
rect 9771 8798 9787 8832
rect 9821 8827 9846 8832
rect 9771 8793 9789 8798
rect 9823 8793 9846 8827
rect 9771 8786 9846 8793
rect 9897 8804 9952 8866
rect 9612 8705 9669 8725
rect 9612 8671 9635 8705
rect 9612 8637 9669 8671
rect 9612 8603 9635 8637
rect 9703 8668 9737 8786
rect 9897 8770 9918 8804
rect 9897 8762 9952 8770
rect 9800 8702 9816 8736
rect 9850 8728 9897 8736
rect 9931 8728 9952 8762
rect 9850 8702 9952 8728
rect 9986 8898 10002 8932
rect 10036 8898 10052 8932
rect 9986 8895 10052 8898
rect 10142 8898 10217 8904
rect 9986 8668 10022 8895
rect 10142 8872 10173 8898
rect 10142 8838 10164 8872
rect 10207 8864 10217 8898
rect 10198 8838 10217 8864
rect 10056 8820 10100 8836
rect 10090 8804 10100 8820
rect 10292 8804 10326 8958
rect 10861 8942 10877 8966
rect 10911 8942 10927 8976
rect 10961 8996 10995 9034
rect 10961 8946 10995 8962
rect 11029 8992 11228 8998
rect 11029 8958 11178 8992
rect 11212 8958 11228 8992
rect 11352 8992 11422 9034
rect 11284 8974 11318 8990
rect 10427 8894 10484 8910
rect 10693 8908 10727 8924
rect 10461 8860 10484 8894
rect 10761 8898 10777 8932
rect 10811 8898 10827 8932
rect 10909 8898 10991 8904
rect 10761 8872 10805 8898
rect 10427 8830 10484 8860
rect 10427 8826 10449 8830
rect 10090 8786 10326 8804
rect 10056 8770 10326 8786
rect 10208 8720 10258 8736
rect 10208 8686 10224 8720
rect 10208 8668 10258 8686
rect 9703 8634 10258 8668
rect 9612 8558 9669 8603
rect 10086 8626 10120 8634
rect 9703 8566 9719 8600
rect 9753 8566 9930 8600
rect 9964 8566 9980 8600
rect 10292 8601 10326 8770
rect 10360 8796 10449 8826
rect 10483 8796 10484 8830
rect 10543 8838 10805 8872
rect 10943 8872 10991 8898
rect 10909 8858 10941 8864
rect 10925 8838 10941 8858
rect 10975 8838 10991 8872
rect 10543 8804 10559 8838
rect 10593 8804 10609 8838
rect 10360 8790 10484 8796
rect 10360 8720 10401 8790
rect 10671 8770 10687 8804
rect 10721 8770 10737 8804
rect 10671 8768 10737 8770
rect 10536 8762 10737 8768
rect 10394 8686 10401 8720
rect 10360 8670 10401 8686
rect 10449 8720 10496 8736
rect 10536 8728 10541 8762
rect 10575 8728 10737 8762
rect 10536 8720 10737 8728
rect 10449 8694 10462 8720
rect 10483 8660 10496 8686
rect 10771 8694 10805 8838
rect 10839 8804 10883 8820
rect 11029 8812 11063 8958
rect 11352 8958 11368 8992
rect 11402 8958 11422 8992
rect 11540 8992 11606 9034
rect 12117 9028 12150 9052
rect 11461 8966 11506 8982
rect 11284 8924 11318 8940
rect 11461 8932 11472 8966
rect 11540 8958 11556 8992
rect 11590 8958 11606 8992
rect 11929 9018 12150 9028
rect 12184 9018 12222 9052
rect 12256 9018 12295 9052
rect 12329 9018 12367 9052
rect 12401 9051 12557 9052
rect 12401 9018 12440 9051
rect 11929 9017 12440 9018
rect 12474 9017 12512 9051
rect 12546 9017 12557 9051
rect 12649 9021 12678 9055
rect 12712 9021 12770 9055
rect 12804 9021 12862 9055
rect 12896 9021 12954 9055
rect 12988 9021 13046 9055
rect 13080 9021 13138 9055
rect 13172 9021 13201 9055
rect 11929 8994 12557 9017
rect 11640 8966 11692 8982
rect 11097 8898 11163 8922
rect 11131 8882 11163 8898
rect 11097 8848 11113 8864
rect 11147 8848 11163 8882
rect 11199 8894 11243 8910
rect 11199 8860 11209 8894
rect 11284 8886 11427 8924
rect 11029 8804 11109 8812
rect 10873 8770 11109 8804
rect 10839 8754 10889 8770
rect 10991 8720 11041 8736
rect 10991 8694 11007 8720
rect 10449 8654 10496 8660
rect 10667 8634 10683 8668
rect 10717 8634 10733 8668
rect 10771 8660 10857 8694
rect 10891 8686 11007 8694
rect 10891 8660 11041 8686
rect 10771 8644 11041 8660
rect 10086 8576 10120 8592
rect 9703 8524 9980 8566
rect 10168 8566 10194 8600
rect 10228 8566 10244 8600
rect 10292 8567 10408 8601
rect 10442 8567 10458 8601
rect 10667 8600 10733 8634
rect 10168 8524 10244 8566
rect 10667 8566 10683 8600
rect 10717 8566 10733 8600
rect 10857 8626 10891 8644
rect 10857 8576 10891 8592
rect 10951 8576 10977 8610
rect 11011 8576 11027 8610
rect 10667 8524 10733 8566
rect 10951 8524 11027 8576
rect 11075 8601 11109 8770
rect 11199 8736 11243 8860
rect 11143 8720 11243 8736
rect 11277 8834 11359 8850
rect 11277 8800 11325 8834
rect 11277 8726 11359 8800
rect 11177 8694 11243 8720
rect 11177 8686 11185 8694
rect 11143 8660 11185 8686
rect 11219 8660 11243 8694
rect 11393 8692 11427 8886
rect 11284 8658 11427 8692
rect 11461 8898 11506 8932
rect 11674 8932 11692 8966
rect 11640 8924 11692 8932
rect 11495 8864 11506 8898
rect 11461 8676 11506 8864
rect 11284 8608 11318 8658
rect 11461 8642 11472 8676
rect 11541 8890 11692 8924
rect 11833 8944 11867 8960
rect 11541 8821 11587 8890
rect 11833 8868 11867 8884
rect 11929 8944 11963 8994
rect 12117 8993 12557 8994
rect 11929 8868 11963 8884
rect 12025 8944 12059 8960
rect 12025 8868 12059 8884
rect 12121 8944 12155 8993
rect 12121 8868 12155 8884
rect 12233 8932 12267 8948
rect 12233 8856 12267 8872
rect 12321 8932 12355 8993
rect 12321 8856 12355 8872
rect 12434 8931 12468 8947
rect 11575 8787 11587 8821
rect 11541 8694 11587 8787
rect 11621 8821 11692 8856
rect 12434 8855 12468 8871
rect 12522 8931 12556 8993
rect 12522 8855 12556 8871
rect 12666 8979 12805 8987
rect 12666 8945 12684 8979
rect 12718 8945 12805 8979
rect 12666 8911 12805 8945
rect 12666 8877 12684 8911
rect 12718 8877 12805 8911
rect 12666 8861 12805 8877
rect 12846 8979 12908 9021
rect 12846 8945 12852 8979
rect 12886 8945 12908 8979
rect 12846 8911 12908 8945
rect 12846 8877 12852 8911
rect 12886 8877 12908 8911
rect 12846 8861 12908 8877
rect 12991 8975 13057 8987
rect 12991 8941 13007 8975
rect 13041 8941 13057 8975
rect 12991 8907 13057 8941
rect 12991 8873 13007 8907
rect 13041 8873 13057 8907
rect 12991 8861 13057 8873
rect 13091 8975 13137 9021
rect 13456 8992 13490 9008
rect 13544 9068 13578 9084
rect 19194 9039 19228 9055
rect 19354 9115 19388 9131
rect 25903 9115 25937 9131
rect 19354 9039 19388 9055
rect 20165 9068 20199 9084
rect 13544 8992 13578 9008
rect 14136 8981 14152 9015
rect 14186 8981 14202 9015
rect 14870 8981 14886 9015
rect 14920 8981 14936 9015
rect 14992 8981 15008 9015
rect 15042 8981 15058 9015
rect 16208 8981 16224 9015
rect 16258 8981 16274 9015
rect 16330 8981 16346 9015
rect 16380 8981 16396 9015
rect 17420 8981 17436 9015
rect 17470 8981 17486 9015
rect 17542 8981 17558 9015
rect 17592 8981 17608 9015
rect 18274 8981 18290 9015
rect 18324 8981 18340 9015
rect 13125 8941 13137 8975
rect 19258 8971 19274 9005
rect 19308 8971 19324 9005
rect 20165 8992 20199 9008
rect 20253 9068 20287 9084
rect 25903 9039 25937 9055
rect 26063 9115 26097 9131
rect 26063 9039 26097 9055
rect 20253 8992 20287 9008
rect 20845 8981 20861 9015
rect 20895 8981 20911 9015
rect 21579 8981 21595 9015
rect 21629 8981 21645 9015
rect 21701 8981 21717 9015
rect 21751 8981 21767 9015
rect 22917 8981 22933 9015
rect 22967 8981 22983 9015
rect 23039 8981 23055 9015
rect 23089 8981 23105 9015
rect 24129 8981 24145 9015
rect 24179 8981 24195 9015
rect 24251 8981 24267 9015
rect 24301 8981 24317 9015
rect 24983 8981 24999 9015
rect 25033 8981 25049 9015
rect 25967 8971 25983 9005
rect 26017 8971 26033 9005
rect 13091 8907 13137 8941
rect 13125 8873 13137 8907
rect 11621 8787 11643 8821
rect 11677 8787 11692 8821
rect 12057 8787 12073 8821
rect 12107 8787 12123 8821
rect 12261 8788 12277 8822
rect 12311 8788 12327 8822
rect 12462 8787 12478 8821
rect 12512 8787 12528 8821
rect 11621 8762 11692 8787
rect 12670 8782 12687 8823
rect 12721 8782 12737 8823
rect 12670 8773 12737 8782
rect 11621 8728 11652 8762
rect 11686 8728 11692 8762
rect 11621 8726 11692 8728
rect 11833 8728 11867 8744
rect 11541 8660 11553 8694
rect 11587 8676 11692 8692
rect 11587 8660 11640 8676
rect 11541 8658 11640 8660
rect 11075 8567 11191 8601
rect 11225 8567 11241 8601
rect 11284 8558 11318 8574
rect 11352 8590 11368 8624
rect 11402 8590 11422 8624
rect 11352 8524 11422 8590
rect 11461 8608 11506 8642
rect 11674 8642 11692 8676
rect 11461 8574 11472 8608
rect 11461 8558 11506 8574
rect 11540 8590 11556 8624
rect 11590 8590 11606 8624
rect 11540 8524 11606 8590
rect 11640 8608 11692 8642
rect 11674 8574 11692 8608
rect 11640 8558 11692 8574
rect 9061 8510 9090 8524
rect 3163 8482 3212 8494
rect 9060 8490 9090 8510
rect 9124 8490 9182 8524
rect 9216 8490 9274 8524
rect 9308 8490 9346 8524
rect 9380 8490 9438 8524
rect 9472 8490 9530 8524
rect 9564 8490 9622 8524
rect 9656 8490 9714 8524
rect 9748 8490 9806 8524
rect 9840 8490 9898 8524
rect 9932 8490 9990 8524
rect 10024 8490 10082 8524
rect 10116 8490 10174 8524
rect 10208 8490 10266 8524
rect 10300 8490 10358 8524
rect 10392 8490 10450 8524
rect 10484 8490 10542 8524
rect 10576 8490 10634 8524
rect 10668 8490 10726 8524
rect 10760 8490 10818 8524
rect 10852 8490 10910 8524
rect 10944 8490 11002 8524
rect 11036 8490 11094 8524
rect 11128 8490 11186 8524
rect 11220 8490 11278 8524
rect 11312 8507 11370 8524
rect 11312 8490 11332 8507
rect 2866 8459 2915 8466
rect 3163 8459 3198 8482
rect 2716 8423 2732 8457
rect 2766 8454 2782 8457
rect 2716 8420 2736 8423
rect 2770 8420 2782 8454
rect 2716 8409 2782 8420
rect 2866 8453 3198 8459
rect 2866 8419 2875 8453
rect 2909 8424 3198 8453
rect 9060 8473 11332 8490
rect 11366 8490 11370 8507
rect 11404 8490 11462 8524
rect 11496 8490 11554 8524
rect 11588 8490 11646 8524
rect 11680 8490 11709 8524
rect 11366 8473 11707 8490
rect 11833 8484 11867 8500
rect 11929 8728 11963 8744
rect 9060 8455 11707 8473
rect 9060 8454 9709 8455
rect 9060 8450 9288 8454
rect 2909 8419 2915 8424
rect 2866 8407 2915 8419
rect 9060 8416 9152 8450
rect 9186 8420 9288 8450
rect 9322 8453 9624 8454
rect 9322 8420 9406 8453
rect 9186 8419 9406 8420
rect 9440 8419 9549 8453
rect 9583 8420 9624 8453
rect 9658 8421 9709 8454
rect 9743 8450 9997 8455
rect 9743 8448 9900 8450
rect 9743 8421 9811 8448
rect 9658 8420 9811 8421
rect 9583 8419 9811 8420
rect 9186 8416 9811 8419
rect 9060 8414 9811 8416
rect 9845 8416 9900 8448
rect 9934 8421 9997 8450
rect 10031 8452 11707 8455
rect 10031 8444 10175 8452
rect 10031 8421 10083 8444
rect 9934 8416 10083 8421
rect 9845 8414 10083 8416
rect 9060 8410 10083 8414
rect 10117 8418 10175 8444
rect 10209 8451 11707 8452
rect 10209 8418 10267 8451
rect 10117 8417 10267 8418
rect 10301 8449 11707 8451
rect 10301 8446 10919 8449
rect 10301 8443 10822 8446
rect 10301 8442 10637 8443
rect 10301 8440 10544 8442
rect 10301 8438 10456 8440
rect 10301 8417 10355 8438
rect 10117 8410 10355 8417
rect 9060 8404 10355 8410
rect 10389 8406 10456 8438
rect 10490 8408 10544 8440
rect 10578 8409 10637 8442
rect 10671 8442 10822 8443
rect 10671 8409 10733 8442
rect 10578 8408 10733 8409
rect 10767 8412 10822 8442
rect 10856 8415 10919 8446
rect 10953 8448 11707 8449
rect 10953 8447 11462 8448
rect 10953 8445 11093 8447
rect 10953 8415 11003 8445
rect 10856 8412 11003 8415
rect 10767 8411 11003 8412
rect 11037 8413 11093 8445
rect 11127 8443 11462 8447
rect 11127 8413 11191 8443
rect 11037 8411 11191 8413
rect 10767 8409 11191 8411
rect 11225 8414 11462 8443
rect 11496 8414 11560 8448
rect 11594 8446 11707 8448
rect 11594 8414 11643 8446
rect 11225 8412 11643 8414
rect 11677 8412 11707 8446
rect 11225 8409 11707 8412
rect 10767 8408 11707 8409
rect 10490 8406 11707 8408
rect 10389 8404 11707 8406
rect 9060 8393 11707 8404
rect 2636 8357 2702 8375
rect 2636 8309 2652 8357
rect 2686 8309 2702 8357
rect 2636 8289 2702 8309
rect 2636 8255 2652 8289
rect 2686 8255 2702 8289
rect 2636 8221 2702 8255
rect 2636 8187 2652 8221
rect 2686 8187 2702 8221
rect 2636 8179 2702 8187
rect 2736 8357 2778 8373
rect 2770 8323 2778 8357
rect 2956 8349 2972 8383
rect 3006 8349 3022 8383
rect 10059 8349 11707 8393
rect 11929 8450 11963 8500
rect 12025 8728 12059 8744
rect 12025 8484 12059 8500
rect 12121 8728 12155 8744
rect 12121 8450 12155 8500
rect 12233 8729 12267 8745
rect 12233 8485 12267 8501
rect 12321 8729 12355 8745
rect 12321 8450 12355 8501
rect 12434 8728 12468 8744
rect 12434 8456 12468 8472
rect 12522 8728 12556 8744
rect 12771 8741 12805 8861
rect 12839 8826 12906 8827
rect 12991 8826 13037 8861
rect 13091 8857 13137 8873
rect 13264 8930 13298 8946
rect 13264 8854 13298 8870
rect 13360 8930 13394 8946
rect 13360 8854 13394 8870
rect 13456 8930 13490 8946
rect 13456 8854 13490 8870
rect 13544 8930 13578 8946
rect 13544 8854 13578 8870
rect 14108 8931 14142 8947
rect 14108 8855 14142 8871
rect 14197 8931 14231 8947
rect 14197 8855 14231 8871
rect 14842 8931 14876 8947
rect 14842 8855 14876 8871
rect 14944 8931 14978 8947
rect 14944 8855 14978 8871
rect 15052 8931 15086 8947
rect 15052 8855 15086 8871
rect 16180 8931 16214 8947
rect 16180 8855 16214 8871
rect 16284 8931 16318 8947
rect 16284 8855 16318 8871
rect 16390 8931 16424 8947
rect 16390 8855 16424 8871
rect 17392 8931 17426 8947
rect 17392 8855 17426 8871
rect 17495 8931 17529 8947
rect 17495 8855 17529 8871
rect 17602 8931 17636 8947
rect 17602 8855 17636 8871
rect 18244 8931 18278 8947
rect 18244 8855 18278 8871
rect 18334 8931 18368 8947
rect 18334 8855 18368 8871
rect 19973 8930 20007 8946
rect 19973 8854 20007 8870
rect 20069 8930 20103 8946
rect 20069 8854 20103 8870
rect 20165 8930 20199 8946
rect 20165 8854 20199 8870
rect 20253 8930 20287 8946
rect 20253 8854 20287 8870
rect 20817 8931 20851 8947
rect 20817 8855 20851 8871
rect 20906 8931 20940 8947
rect 20906 8855 20940 8871
rect 21551 8931 21585 8947
rect 21551 8855 21585 8871
rect 21653 8931 21687 8947
rect 21653 8855 21687 8871
rect 21761 8931 21795 8947
rect 21761 8855 21795 8871
rect 22889 8931 22923 8947
rect 22889 8855 22923 8871
rect 22993 8931 23027 8947
rect 22993 8855 23027 8871
rect 23099 8931 23133 8947
rect 23099 8855 23133 8871
rect 24101 8931 24135 8947
rect 24101 8855 24135 8871
rect 24204 8931 24238 8947
rect 24204 8855 24238 8871
rect 24311 8931 24345 8947
rect 24311 8855 24345 8871
rect 24953 8931 24987 8947
rect 24953 8855 24987 8871
rect 25043 8931 25077 8947
rect 25043 8855 25077 8871
rect 12839 8823 13037 8826
rect 12839 8789 12855 8823
rect 12889 8789 13037 8823
rect 12839 8774 13037 8789
rect 13071 8820 13087 8823
rect 13071 8786 13085 8820
rect 13121 8789 13137 8823
rect 13119 8786 13137 8789
rect 13392 8786 13408 8820
rect 13442 8786 13458 8820
rect 13071 8775 13137 8786
rect 13599 8784 13615 8818
rect 13649 8784 13665 8818
rect 20101 8786 20117 8820
rect 20151 8786 20167 8820
rect 20308 8784 20324 8818
rect 20358 8784 20374 8818
rect 12839 8773 12906 8774
rect 12991 8741 13037 8774
rect 12666 8723 12718 8739
rect 12666 8689 12684 8723
rect 12666 8655 12718 8689
rect 12666 8621 12684 8655
rect 12666 8587 12718 8621
rect 12666 8553 12684 8587
rect 12666 8511 12718 8553
rect 12752 8723 12818 8741
rect 12752 8689 12768 8723
rect 12802 8689 12818 8723
rect 12752 8655 12818 8689
rect 12752 8630 12768 8655
rect 12752 8596 12767 8630
rect 12802 8621 12818 8655
rect 12801 8596 12818 8621
rect 12752 8587 12818 8596
rect 12752 8553 12768 8587
rect 12802 8553 12818 8587
rect 12752 8545 12818 8553
rect 12852 8723 12908 8739
rect 12886 8689 12908 8723
rect 12852 8655 12908 8689
rect 12886 8621 12908 8655
rect 12852 8587 12908 8621
rect 12886 8553 12908 8587
rect 12852 8511 12908 8553
rect 12991 8723 13057 8741
rect 12991 8689 13007 8723
rect 13041 8689 13057 8723
rect 12991 8655 13057 8689
rect 12991 8621 13007 8655
rect 13041 8621 13057 8655
rect 12991 8587 13057 8621
rect 12991 8553 13007 8587
rect 13041 8553 13057 8587
rect 12991 8545 13057 8553
rect 13091 8723 13133 8739
rect 13125 8689 13133 8723
rect 13091 8655 13133 8689
rect 13125 8621 13133 8655
rect 13264 8727 13298 8743
rect 13264 8651 13298 8667
rect 13360 8727 13394 8743
rect 13360 8651 13394 8667
rect 13456 8727 13490 8743
rect 13456 8651 13490 8667
rect 13544 8727 13578 8743
rect 13544 8651 13578 8667
rect 14105 8730 14139 8746
rect 14105 8654 14139 8670
rect 14212 8730 14246 8746
rect 14212 8654 14246 8670
rect 14319 8730 14353 8746
rect 14319 8654 14353 8670
rect 15317 8730 15351 8746
rect 15317 8654 15351 8670
rect 15426 8730 15460 8746
rect 15426 8654 15460 8670
rect 15531 8730 15565 8746
rect 15531 8654 15565 8670
rect 16529 8730 16563 8746
rect 16529 8654 16563 8670
rect 16639 8730 16673 8746
rect 16639 8654 16673 8670
rect 16743 8730 16777 8746
rect 16743 8654 16777 8670
rect 17741 8730 17775 8746
rect 17741 8654 17775 8670
rect 17850 8730 17884 8746
rect 17850 8654 17884 8670
rect 17955 8730 17989 8746
rect 17955 8654 17989 8670
rect 18599 8730 18633 8746
rect 18599 8654 18633 8670
rect 18687 8733 18721 8749
rect 19973 8727 20007 8743
rect 19499 8677 19515 8706
rect 18687 8657 18721 8673
rect 19445 8643 19474 8677
rect 19508 8672 19515 8677
rect 19549 8677 19567 8706
rect 19633 8677 19659 8706
rect 19693 8677 19709 8706
rect 19751 8677 19777 8706
rect 19811 8677 19827 8706
rect 19549 8672 19566 8677
rect 19508 8643 19566 8672
rect 19600 8643 19658 8677
rect 19693 8672 19750 8677
rect 19811 8672 19842 8677
rect 19692 8643 19750 8672
rect 19784 8643 19842 8672
rect 19876 8643 19905 8677
rect 19973 8651 20007 8667
rect 20069 8727 20103 8743
rect 20069 8651 20103 8667
rect 20165 8727 20199 8743
rect 20165 8651 20199 8667
rect 20253 8727 20287 8743
rect 20253 8651 20287 8667
rect 20814 8730 20848 8746
rect 20814 8654 20848 8670
rect 20921 8730 20955 8746
rect 20921 8654 20955 8670
rect 21028 8730 21062 8746
rect 21028 8654 21062 8670
rect 22026 8730 22060 8746
rect 22026 8654 22060 8670
rect 22135 8730 22169 8746
rect 22135 8654 22169 8670
rect 22240 8730 22274 8746
rect 22240 8654 22274 8670
rect 23238 8730 23272 8746
rect 23238 8654 23272 8670
rect 23348 8730 23382 8746
rect 23348 8654 23382 8670
rect 23452 8730 23486 8746
rect 23452 8654 23486 8670
rect 24450 8730 24484 8746
rect 24450 8654 24484 8670
rect 24559 8730 24593 8746
rect 24559 8654 24593 8670
rect 24664 8730 24698 8746
rect 24664 8654 24698 8670
rect 25308 8730 25342 8746
rect 25308 8654 25342 8670
rect 25396 8733 25430 8749
rect 26208 8677 26224 8706
rect 25396 8657 25430 8673
rect 26154 8643 26183 8677
rect 26217 8672 26224 8677
rect 26258 8677 26276 8706
rect 26342 8677 26368 8706
rect 26402 8677 26418 8706
rect 26460 8677 26486 8706
rect 26520 8677 26536 8706
rect 26258 8672 26275 8677
rect 26217 8643 26275 8672
rect 26309 8643 26367 8677
rect 26402 8672 26459 8677
rect 26520 8672 26551 8677
rect 26401 8643 26459 8672
rect 26493 8643 26551 8672
rect 26585 8643 26614 8677
rect 13091 8587 13133 8621
rect 13125 8553 13133 8587
rect 13091 8511 13133 8553
rect 13456 8589 13490 8605
rect 13456 8513 13490 8529
rect 13544 8589 13578 8605
rect 14133 8577 14149 8611
rect 14183 8577 14199 8611
rect 14259 8577 14275 8611
rect 14309 8577 14325 8611
rect 15345 8577 15361 8611
rect 15395 8577 15411 8611
rect 15471 8577 15487 8611
rect 15521 8577 15537 8611
rect 16557 8577 16573 8611
rect 16607 8577 16623 8611
rect 16683 8577 16699 8611
rect 16733 8577 16749 8611
rect 17769 8577 17785 8611
rect 17819 8577 17835 8611
rect 17895 8577 17911 8611
rect 17945 8577 17961 8611
rect 18627 8580 18643 8614
rect 18677 8580 18693 8614
rect 19078 8610 19127 8622
rect 19078 8609 19218 8610
rect 19078 8575 19084 8609
rect 19118 8576 19218 8609
rect 19118 8575 19127 8576
rect 19078 8563 19127 8575
rect 19177 8534 19218 8576
rect 19509 8597 19555 8643
rect 19509 8563 19521 8597
rect 19338 8534 19387 8547
rect 13544 8513 13578 8529
rect 19079 8516 19128 8529
rect 12649 8477 12678 8511
rect 12712 8477 12770 8511
rect 12804 8477 12862 8511
rect 12896 8477 12954 8511
rect 12988 8477 13046 8511
rect 13080 8477 13138 8511
rect 13172 8477 13201 8511
rect 19079 8482 19085 8516
rect 19119 8482 19128 8516
rect 19177 8500 19344 8534
rect 19378 8500 19387 8534
rect 19338 8488 19387 8500
rect 19509 8529 19555 8563
rect 19509 8495 19521 8529
rect 11929 8427 12355 8450
rect 11929 8393 12200 8427
rect 12234 8393 12274 8427
rect 12308 8422 12355 8427
rect 12522 8422 12556 8472
rect 19079 8470 19128 8482
rect 19509 8479 19555 8495
rect 19589 8597 19655 8609
rect 19589 8563 19605 8597
rect 19639 8563 19655 8597
rect 19589 8529 19655 8563
rect 19589 8495 19605 8529
rect 19639 8495 19655 8529
rect 19589 8483 19655 8495
rect 12308 8393 12556 8422
rect 19093 8447 19128 8470
rect 19376 8447 19425 8454
rect 19093 8441 19425 8447
rect 19093 8412 19382 8441
rect 19376 8407 19382 8412
rect 19416 8407 19425 8441
rect 19376 8395 19425 8407
rect 19509 8442 19525 8445
rect 19509 8408 19521 8442
rect 19559 8411 19575 8445
rect 19555 8408 19575 8411
rect 19509 8397 19575 8408
rect 11929 8374 12589 8393
rect 2736 8289 2778 8323
rect 10054 8315 10083 8349
rect 10117 8315 10175 8349
rect 10209 8315 10267 8349
rect 10301 8315 10359 8349
rect 10393 8315 10451 8349
rect 10485 8315 10543 8349
rect 10577 8315 10635 8349
rect 10669 8315 10727 8349
rect 10761 8315 10819 8349
rect 10853 8315 10910 8349
rect 10944 8315 11002 8349
rect 11036 8315 11094 8349
rect 11128 8315 11186 8349
rect 11220 8315 11278 8349
rect 11312 8315 11370 8349
rect 11404 8315 11462 8349
rect 11496 8315 11554 8349
rect 11588 8315 11646 8349
rect 11680 8315 11709 8349
rect 11833 8324 11867 8340
rect 2770 8255 2778 8289
rect 2736 8221 2778 8255
rect 2770 8187 2778 8221
rect 2928 8290 2962 8306
rect 2928 8214 2962 8230
rect 3016 8290 3050 8306
rect 10072 8273 10139 8281
rect 3016 8214 3050 8230
rect 8867 8221 8953 8247
rect 2736 8145 2778 8187
rect 8867 8187 8893 8221
rect 8927 8187 8953 8221
rect 2928 8152 2962 8168
rect 2386 8111 2415 8145
rect 2449 8116 2507 8145
rect 2449 8111 2460 8116
rect 2444 8082 2460 8111
rect 2494 8111 2507 8116
rect 2541 8116 2599 8145
rect 2541 8111 2590 8116
rect 2633 8111 2691 8145
rect 2725 8116 2783 8145
rect 2725 8111 2736 8116
rect 2494 8082 2510 8111
rect 2574 8082 2590 8111
rect 2624 8082 2644 8111
rect 2720 8082 2736 8111
rect 2770 8111 2783 8116
rect 2817 8111 2846 8145
rect 2770 8082 2790 8111
rect 2928 8076 2962 8092
rect 3016 8152 3050 8168
rect 8867 8161 8953 8187
rect 10072 8239 10089 8273
rect 10123 8239 10139 8273
rect 10072 8205 10139 8239
rect 10072 8171 10089 8205
rect 10123 8171 10139 8205
rect 3016 8076 3050 8092
rect 10072 8137 10139 8171
rect 10072 8103 10089 8137
rect 10123 8103 10139 8137
rect 8868 8064 8954 8090
rect 8868 8030 8894 8064
rect 8928 8030 8954 8064
rect 2928 8014 2962 8030
rect 2928 7938 2962 7954
rect 3016 8014 3050 8030
rect 8868 8004 8954 8030
rect 10072 8087 10139 8103
rect 10173 8273 10207 8315
rect 10173 8205 10207 8239
rect 10173 8137 10207 8171
rect 10173 8087 10207 8103
rect 10241 8247 10647 8281
rect 3016 7938 3050 7954
rect 10072 7953 10106 8087
rect 10241 8053 10275 8247
rect 10140 8037 10191 8053
rect 10174 8003 10191 8037
rect 10140 7987 10191 8003
rect 10236 8037 10275 8053
rect 10270 8003 10275 8037
rect 10236 7987 10275 8003
rect 10309 8179 10409 8213
rect 10443 8179 10484 8213
rect 10518 8179 10534 8213
rect 10157 7953 10191 7987
rect 10309 7953 10343 8179
rect 8868 7894 8954 7920
rect 2928 7876 2962 7892
rect 2928 7800 2962 7816
rect 3016 7876 3050 7892
rect 8868 7860 8894 7894
rect 8928 7860 8954 7894
rect 8868 7834 8954 7860
rect 10072 7905 10123 7953
rect 10157 7919 10343 7953
rect 10377 8114 10579 8145
rect 10377 8111 10545 8114
rect 10377 8001 10411 8111
rect 10541 8080 10545 8111
rect 10377 7951 10411 7967
rect 10452 8001 10507 8071
rect 10452 7967 10473 8001
rect 10072 7871 10078 7905
rect 10112 7900 10123 7905
rect 10308 7912 10343 7919
rect 10308 7896 10414 7912
rect 10072 7866 10089 7871
rect 10072 7839 10123 7866
rect 10157 7881 10223 7885
rect 10157 7847 10173 7881
rect 10207 7847 10223 7881
rect 3016 7800 3050 7816
rect 10157 7805 10223 7847
rect 10308 7862 10380 7896
rect 10308 7839 10414 7862
rect 10452 7908 10507 7967
rect 10452 7874 10465 7908
rect 10499 7874 10507 7908
rect 10452 7839 10507 7874
rect 10541 7843 10579 8080
rect 10613 8114 10647 8247
rect 10681 8213 10715 8315
rect 10899 8273 10966 8281
rect 10681 8163 10715 8179
rect 10762 8213 10865 8245
rect 10762 8179 10767 8213
rect 10801 8179 10865 8213
rect 10762 8163 10865 8179
rect 10613 8080 10713 8114
rect 10747 8112 10763 8114
rect 10613 8078 10715 8080
rect 10749 8078 10763 8112
rect 10613 8076 10763 8078
rect 10797 8001 10865 8163
rect 10619 7967 10635 8001
rect 10669 7967 10865 8001
rect 10899 8239 10916 8273
rect 10950 8239 10966 8273
rect 10899 8205 10966 8239
rect 10899 8171 10916 8205
rect 10950 8171 10966 8205
rect 10899 8137 10966 8171
rect 10899 8103 10916 8137
rect 10950 8103 10966 8137
rect 10899 8087 10966 8103
rect 11000 8273 11034 8315
rect 11000 8205 11034 8239
rect 11000 8137 11034 8171
rect 11000 8087 11034 8103
rect 11068 8247 11474 8281
rect 10615 7896 10717 7912
rect 10649 7862 10683 7896
rect 10541 7805 10580 7843
rect 10615 7805 10717 7862
rect 10761 7896 10810 7967
rect 10761 7862 10767 7896
rect 10801 7862 10810 7896
rect 10761 7846 10810 7862
rect 10899 7953 10933 8087
rect 11068 8053 11102 8247
rect 10967 8037 11018 8053
rect 11001 8003 11018 8037
rect 10967 7987 11018 8003
rect 11063 8037 11102 8053
rect 11097 8003 11102 8037
rect 11063 7987 11102 8003
rect 11136 8179 11236 8213
rect 11270 8179 11311 8213
rect 11345 8179 11361 8213
rect 10984 7953 11018 7987
rect 11136 7953 11170 8179
rect 10899 7908 10950 7953
rect 10984 7919 11170 7953
rect 11204 8114 11406 8145
rect 11204 8111 11372 8114
rect 11204 8001 11238 8111
rect 11368 8080 11372 8111
rect 11204 7951 11238 7967
rect 11279 8042 11334 8071
rect 11279 8008 11286 8042
rect 11320 8008 11334 8042
rect 11279 8001 11334 8008
rect 11279 7967 11300 8001
rect 10899 7874 10910 7908
rect 10944 7900 10950 7908
rect 11135 7912 11170 7919
rect 11135 7896 11241 7912
rect 10899 7866 10916 7874
rect 10899 7839 10950 7866
rect 10984 7881 11050 7885
rect 10984 7847 11000 7881
rect 11034 7847 11050 7881
rect 10984 7805 11050 7847
rect 11135 7862 11207 7896
rect 11135 7839 11241 7862
rect 11279 7839 11334 7967
rect 11368 7841 11406 8080
rect 11440 8114 11474 8247
rect 11508 8213 11542 8315
rect 11508 8163 11542 8179
rect 11589 8213 11692 8245
rect 11589 8179 11594 8213
rect 11628 8179 11692 8213
rect 11589 8163 11692 8179
rect 11440 8112 11540 8114
rect 11440 8078 11538 8112
rect 11574 8080 11590 8114
rect 11572 8078 11590 8080
rect 11440 8076 11590 8078
rect 11624 8001 11692 8163
rect 11833 8080 11867 8096
rect 11929 8324 11963 8374
rect 11929 8080 11963 8096
rect 12025 8324 12059 8340
rect 12025 8080 12059 8096
rect 12121 8324 12155 8374
rect 12321 8371 12589 8374
rect 12121 8080 12155 8096
rect 12233 8323 12267 8339
rect 12233 8079 12267 8095
rect 12321 8338 12452 8371
rect 12486 8370 12589 8371
rect 12321 8323 12355 8338
rect 12426 8335 12452 8338
rect 12486 8336 12531 8370
rect 12566 8336 12589 8370
rect 19269 8337 19285 8371
rect 19319 8337 19335 8371
rect 19609 8363 19655 8483
rect 19513 8345 19555 8361
rect 12486 8335 12589 8336
rect 12426 8309 12589 8335
rect 19513 8311 19521 8345
rect 19241 8278 19275 8294
rect 12730 8190 12746 8224
rect 12780 8190 12796 8224
rect 13338 8209 13424 8235
rect 13338 8175 13364 8209
rect 13398 8175 13424 8209
rect 19241 8202 19275 8218
rect 19329 8278 19363 8294
rect 19329 8202 19363 8218
rect 19513 8277 19555 8311
rect 19513 8243 19521 8277
rect 19513 8209 19555 8243
rect 12321 8079 12355 8095
rect 12702 8140 12736 8156
rect 12702 8064 12736 8080
rect 12790 8140 12824 8156
rect 13338 8149 13424 8175
rect 19513 8175 19521 8209
rect 12790 8064 12824 8080
rect 19241 8140 19275 8156
rect 13337 8052 13423 8078
rect 19241 8064 19275 8080
rect 19329 8140 19363 8156
rect 19513 8133 19555 8175
rect 19589 8345 19655 8363
rect 19589 8297 19605 8345
rect 19639 8297 19655 8345
rect 19589 8277 19655 8297
rect 19589 8243 19605 8277
rect 19639 8243 19655 8277
rect 19589 8209 19655 8243
rect 19589 8175 19605 8209
rect 19639 8175 19655 8209
rect 19589 8167 19655 8175
rect 19695 8597 19761 8609
rect 19695 8563 19711 8597
rect 19745 8563 19761 8597
rect 19695 8529 19761 8563
rect 19695 8495 19711 8529
rect 19745 8495 19761 8529
rect 19695 8483 19761 8495
rect 19795 8597 19841 8643
rect 19829 8563 19841 8597
rect 19795 8529 19841 8563
rect 19829 8495 19841 8529
rect 20165 8589 20199 8605
rect 20165 8513 20199 8529
rect 20253 8589 20287 8605
rect 20842 8577 20858 8611
rect 20892 8577 20908 8611
rect 20968 8577 20984 8611
rect 21018 8577 21034 8611
rect 22054 8577 22070 8611
rect 22104 8577 22120 8611
rect 22180 8577 22196 8611
rect 22230 8577 22246 8611
rect 23266 8577 23282 8611
rect 23316 8577 23332 8611
rect 23392 8577 23408 8611
rect 23442 8577 23458 8611
rect 24478 8577 24494 8611
rect 24528 8577 24544 8611
rect 24604 8577 24620 8611
rect 24654 8577 24670 8611
rect 25336 8580 25352 8614
rect 25386 8580 25402 8614
rect 25787 8610 25836 8622
rect 25787 8609 25927 8610
rect 25787 8575 25793 8609
rect 25827 8576 25927 8609
rect 25827 8575 25836 8576
rect 25787 8563 25836 8575
rect 25886 8534 25927 8576
rect 26218 8597 26264 8643
rect 26218 8563 26230 8597
rect 26047 8534 26096 8547
rect 20253 8513 20287 8529
rect 25788 8516 25837 8529
rect 19695 8363 19741 8483
rect 19795 8479 19841 8495
rect 25788 8482 25794 8516
rect 25828 8482 25837 8516
rect 25886 8500 26053 8534
rect 26087 8500 26096 8534
rect 26047 8488 26096 8500
rect 26218 8529 26264 8563
rect 26218 8495 26230 8529
rect 25788 8470 25837 8482
rect 26218 8479 26264 8495
rect 26298 8597 26364 8609
rect 26298 8563 26314 8597
rect 26348 8563 26364 8597
rect 26298 8529 26364 8563
rect 26298 8495 26314 8529
rect 26348 8495 26364 8529
rect 26298 8483 26364 8495
rect 25802 8447 25837 8470
rect 26085 8447 26134 8454
rect 19775 8411 19791 8445
rect 19825 8441 19841 8445
rect 19775 8407 19795 8411
rect 19829 8407 19841 8441
rect 25802 8441 26134 8447
rect 25802 8412 26091 8441
rect 19775 8397 19841 8407
rect 26085 8407 26091 8412
rect 26125 8407 26134 8441
rect 26085 8395 26134 8407
rect 26218 8442 26234 8445
rect 26218 8408 26230 8442
rect 26268 8411 26284 8445
rect 26264 8408 26284 8411
rect 26218 8397 26284 8408
rect 19695 8345 19761 8363
rect 19695 8311 19711 8345
rect 19745 8311 19761 8345
rect 19695 8277 19761 8311
rect 19695 8243 19711 8277
rect 19745 8276 19761 8277
rect 19695 8242 19714 8243
rect 19748 8242 19761 8276
rect 19695 8209 19761 8242
rect 19695 8175 19711 8209
rect 19745 8175 19761 8209
rect 19695 8167 19761 8175
rect 19795 8345 19837 8361
rect 19829 8311 19837 8345
rect 25978 8337 25994 8371
rect 26028 8337 26044 8371
rect 26318 8363 26364 8483
rect 26222 8345 26264 8361
rect 19795 8277 19837 8311
rect 26222 8311 26230 8345
rect 19829 8243 19837 8277
rect 19795 8209 19837 8243
rect 25950 8278 25984 8294
rect 19829 8175 19837 8209
rect 19795 8133 19837 8175
rect 20047 8209 20133 8235
rect 20047 8175 20073 8209
rect 20107 8175 20133 8209
rect 25950 8202 25984 8218
rect 26038 8278 26072 8294
rect 26038 8202 26072 8218
rect 26222 8277 26264 8311
rect 26222 8243 26230 8277
rect 26222 8209 26264 8243
rect 20047 8149 20133 8175
rect 26222 8175 26230 8209
rect 25950 8140 25984 8156
rect 19445 8099 19474 8133
rect 19508 8104 19566 8133
rect 19508 8099 19521 8104
rect 19329 8064 19363 8080
rect 19501 8070 19521 8099
rect 19555 8099 19566 8104
rect 19600 8099 19658 8133
rect 19692 8104 19750 8133
rect 19701 8099 19750 8104
rect 19784 8104 19842 8133
rect 19784 8099 19797 8104
rect 19555 8070 19571 8099
rect 19647 8070 19667 8099
rect 19701 8070 19717 8099
rect 19781 8070 19797 8099
rect 19831 8099 19842 8104
rect 19876 8099 19905 8133
rect 19831 8070 19847 8099
rect 12057 8003 12073 8037
rect 12107 8003 12123 8037
rect 12261 8002 12277 8036
rect 12311 8002 12327 8036
rect 13337 8018 13363 8052
rect 13397 8018 13423 8052
rect 20046 8052 20132 8078
rect 25950 8064 25984 8080
rect 26038 8140 26072 8156
rect 26222 8133 26264 8175
rect 26298 8345 26364 8363
rect 26298 8297 26314 8345
rect 26348 8297 26364 8345
rect 26298 8277 26364 8297
rect 26298 8243 26314 8277
rect 26348 8243 26364 8277
rect 26298 8209 26364 8243
rect 26298 8175 26314 8209
rect 26348 8175 26364 8209
rect 26298 8167 26364 8175
rect 26404 8597 26470 8609
rect 26404 8563 26420 8597
rect 26454 8563 26470 8597
rect 26404 8529 26470 8563
rect 26404 8495 26420 8529
rect 26454 8495 26470 8529
rect 26404 8483 26470 8495
rect 26504 8597 26550 8643
rect 26538 8563 26550 8597
rect 26504 8529 26550 8563
rect 26538 8495 26550 8529
rect 26404 8363 26450 8483
rect 26504 8479 26550 8495
rect 26484 8411 26500 8445
rect 26534 8441 26550 8445
rect 26484 8407 26504 8411
rect 26538 8407 26550 8441
rect 26484 8397 26550 8407
rect 26404 8345 26470 8363
rect 26404 8311 26420 8345
rect 26454 8311 26470 8345
rect 26404 8277 26470 8311
rect 26404 8243 26420 8277
rect 26454 8276 26470 8277
rect 26404 8242 26423 8243
rect 26457 8242 26470 8276
rect 26404 8209 26470 8242
rect 26404 8175 26420 8209
rect 26454 8175 26470 8209
rect 26404 8167 26470 8175
rect 26504 8345 26546 8361
rect 26538 8311 26546 8345
rect 26504 8277 26546 8311
rect 26538 8243 26546 8277
rect 26504 8209 26546 8243
rect 26538 8175 26546 8209
rect 26504 8133 26546 8175
rect 26154 8099 26183 8133
rect 26217 8104 26275 8133
rect 26217 8099 26230 8104
rect 26038 8064 26072 8080
rect 26210 8070 26230 8099
rect 26264 8099 26275 8104
rect 26309 8099 26367 8133
rect 26401 8104 26459 8133
rect 26410 8099 26459 8104
rect 26493 8104 26551 8133
rect 26493 8099 26506 8104
rect 26264 8070 26280 8099
rect 26356 8070 26376 8099
rect 26410 8070 26426 8099
rect 26490 8070 26506 8099
rect 26540 8099 26551 8104
rect 26585 8099 26614 8133
rect 26540 8070 26556 8099
rect 20046 8018 20072 8052
rect 20106 8018 20132 8052
rect 11446 7967 11462 8001
rect 11496 7967 11692 8001
rect 13337 7992 13423 8018
rect 19241 8002 19275 8018
rect 11442 7896 11544 7912
rect 11476 7862 11510 7896
rect 11368 7805 11407 7841
rect 11442 7805 11544 7862
rect 11588 7896 11637 7967
rect 11588 7862 11594 7896
rect 11628 7862 11637 7896
rect 11833 7940 11867 7956
rect 11833 7864 11867 7880
rect 11929 7940 11963 7956
rect 11588 7846 11637 7862
rect 11929 7830 11963 7880
rect 12025 7940 12059 7956
rect 12025 7864 12059 7880
rect 12121 7940 12155 7956
rect 12121 7830 12155 7880
rect 12233 7952 12267 7968
rect 12233 7876 12267 7892
rect 12321 7952 12355 7968
rect 12321 7830 12355 7892
rect 2928 7738 2962 7754
rect 2928 7662 2962 7678
rect 3016 7738 3050 7754
rect 3016 7662 3050 7678
rect 3116 7729 3199 7753
rect 3116 7694 3141 7729
rect 3175 7694 3199 7729
rect 3116 7669 3199 7694
rect 8867 7742 8953 7768
rect 8867 7708 8893 7742
rect 8927 7708 8953 7742
rect 10054 7737 10083 7805
rect 10117 7737 10175 7805
rect 10209 7737 10267 7805
rect 10301 7737 10359 7805
rect 10393 7737 10451 7805
rect 10485 7771 10543 7805
rect 10577 7771 10635 7805
rect 10669 7771 10727 7805
rect 10761 7771 10819 7805
rect 10853 7771 10910 7805
rect 10485 7737 10534 7771
rect 10054 7734 10534 7737
rect 10668 7737 10727 7771
rect 10761 7770 10910 7771
rect 10761 7737 10819 7770
rect 10668 7736 10819 7737
rect 10853 7737 10910 7770
rect 10944 7737 11002 7805
rect 11036 7771 11094 7805
rect 11128 7771 11186 7805
rect 11036 7737 11095 7771
rect 11129 7737 11186 7771
rect 11220 7737 11278 7805
rect 11312 7771 11370 7805
rect 11404 7771 11462 7805
rect 11496 7771 11554 7805
rect 11588 7771 11646 7805
rect 11680 7771 11709 7805
rect 11312 7737 11336 7771
rect 10853 7736 11336 7737
rect 10668 7732 11336 7736
rect 11494 7770 11707 7771
rect 11494 7736 11554 7770
rect 11588 7736 11646 7770
rect 11680 7736 11707 7770
rect 11929 7768 12355 7830
rect 11494 7732 11707 7736
rect 11928 7762 12355 7768
rect 8867 7682 8953 7708
rect 11928 7728 11942 7762
rect 11976 7728 12014 7762
rect 12048 7728 12087 7762
rect 12121 7728 12159 7762
rect 12193 7761 12355 7762
rect 12193 7728 12232 7761
rect 11928 7727 12232 7728
rect 12266 7727 12304 7761
rect 12338 7760 12355 7761
rect 12702 7952 12736 7968
rect 12338 7727 12356 7760
rect 11928 7690 12356 7727
rect 2928 7600 2962 7616
rect 2928 7524 2962 7540
rect 3016 7605 3050 7616
rect 3129 7605 3186 7669
rect 11928 7656 11941 7690
rect 11975 7656 12013 7690
rect 12047 7656 12086 7690
rect 12120 7656 12158 7690
rect 12192 7689 12356 7690
rect 12192 7656 12231 7689
rect 11928 7655 12231 7656
rect 12265 7655 12303 7689
rect 12337 7655 12356 7689
rect 3016 7600 3186 7605
rect 3050 7564 3186 7600
rect 8862 7598 8948 7624
rect 8862 7564 8888 7598
rect 8922 7564 8948 7598
rect 3050 7550 3728 7564
rect 3050 7540 3174 7550
rect 3016 7524 3174 7540
rect 3058 7516 3174 7524
rect 3210 7516 3254 7550
rect 3290 7516 3334 7550
rect 3370 7516 3414 7550
rect 3450 7516 3494 7550
rect 3530 7516 3574 7550
rect 3610 7516 3728 7550
rect 3058 7498 3728 7516
rect 3790 7547 8698 7561
rect 3790 7513 3906 7547
rect 3942 7513 3986 7547
rect 4022 7513 4066 7547
rect 4102 7513 4146 7547
rect 4182 7513 4226 7547
rect 4262 7513 4306 7547
rect 4342 7513 4510 7547
rect 4546 7513 4590 7547
rect 4626 7513 4670 7547
rect 4706 7513 4750 7547
rect 4786 7513 4830 7547
rect 4866 7513 4910 7547
rect 4946 7513 5118 7547
rect 5154 7513 5198 7547
rect 5234 7513 5278 7547
rect 5314 7513 5358 7547
rect 5394 7513 5438 7547
rect 5474 7513 5518 7547
rect 5554 7513 5722 7547
rect 5758 7513 5802 7547
rect 5838 7513 5882 7547
rect 5918 7513 5962 7547
rect 5998 7513 6042 7547
rect 6078 7513 6122 7547
rect 6158 7513 6330 7547
rect 6366 7513 6410 7547
rect 6446 7513 6490 7547
rect 6526 7513 6570 7547
rect 6606 7513 6650 7547
rect 6686 7513 6730 7547
rect 6766 7513 6934 7547
rect 6970 7513 7014 7547
rect 7050 7513 7094 7547
rect 7130 7513 7174 7547
rect 7210 7513 7254 7547
rect 7290 7513 7334 7547
rect 7370 7513 7542 7547
rect 7578 7513 7622 7547
rect 7658 7513 7702 7547
rect 7738 7513 7782 7547
rect 7818 7513 7862 7547
rect 7898 7513 7942 7547
rect 7978 7513 8146 7547
rect 8182 7513 8226 7547
rect 8262 7513 8306 7547
rect 8342 7513 8386 7547
rect 8422 7513 8466 7547
rect 8502 7513 8546 7547
rect 8582 7513 8698 7547
rect 8862 7538 8948 7564
rect 11928 7618 12356 7655
rect 11928 7584 11941 7618
rect 11975 7584 12013 7618
rect 12047 7584 12086 7618
rect 12120 7584 12158 7618
rect 12192 7617 12356 7618
rect 12192 7584 12231 7617
rect 11928 7583 12231 7584
rect 12265 7583 12303 7617
rect 12337 7583 12356 7617
rect 11928 7546 12356 7583
rect 12702 7580 12736 7596
rect 12790 7952 12824 7968
rect 12921 7918 13007 7944
rect 19241 7926 19275 7942
rect 19329 8002 19363 8018
rect 19329 7926 19363 7942
rect 19624 7980 19710 8006
rect 20046 7992 20132 8018
rect 25950 8002 25984 8018
rect 19624 7946 19650 7980
rect 19684 7946 19710 7980
rect 19624 7920 19710 7946
rect 25950 7926 25984 7942
rect 26038 8002 26072 8018
rect 26038 7926 26072 7942
rect 12921 7884 12947 7918
rect 12981 7884 13007 7918
rect 12921 7858 13007 7884
rect 13337 7882 13423 7908
rect 13337 7848 13363 7882
rect 13397 7848 13423 7882
rect 20046 7882 20132 7908
rect 13337 7822 13423 7848
rect 19241 7864 19275 7880
rect 19241 7788 19275 7804
rect 19329 7864 19363 7880
rect 20046 7848 20072 7882
rect 20106 7848 20132 7882
rect 20046 7822 20132 7848
rect 25950 7864 25984 7880
rect 19329 7788 19363 7804
rect 19624 7784 19710 7810
rect 25950 7788 25984 7804
rect 26038 7864 26072 7880
rect 26038 7788 26072 7804
rect 13338 7730 13424 7756
rect 19624 7750 19650 7784
rect 19684 7750 19710 7784
rect 12913 7698 12999 7724
rect 12913 7664 12939 7698
rect 12973 7664 12999 7698
rect 13338 7696 13364 7730
rect 13398 7696 13424 7730
rect 13338 7670 13424 7696
rect 19092 7717 19175 7741
rect 19092 7682 19116 7717
rect 19150 7682 19175 7717
rect 12913 7638 12999 7664
rect 19092 7657 19175 7682
rect 19241 7726 19275 7742
rect 12790 7580 12824 7596
rect 13343 7586 13429 7612
rect 3790 7495 8698 7513
rect 11928 7512 11940 7546
rect 11974 7512 12012 7546
rect 12046 7512 12085 7546
rect 12119 7512 12157 7546
rect 12191 7545 12356 7546
rect 12191 7512 12230 7545
rect 11928 7511 12230 7512
rect 12264 7511 12302 7545
rect 12336 7511 12356 7545
rect 13343 7552 13369 7586
rect 13403 7552 13429 7586
rect 19105 7593 19162 7657
rect 19241 7650 19275 7666
rect 19329 7726 19363 7742
rect 19624 7724 19710 7750
rect 20047 7730 20133 7756
rect 20047 7696 20073 7730
rect 20107 7696 20133 7730
rect 20047 7670 20133 7696
rect 25801 7717 25884 7741
rect 25801 7682 25825 7717
rect 25859 7682 25884 7717
rect 19329 7650 19363 7666
rect 25801 7657 25884 7682
rect 25950 7726 25984 7742
rect 19624 7609 19710 7635
rect 19241 7593 19275 7604
rect 19105 7588 19275 7593
rect 19105 7552 19241 7588
rect 11928 7492 12356 7511
rect 12730 7503 12746 7537
rect 12780 7503 12796 7537
rect 13343 7526 13429 7552
rect 13593 7535 18501 7549
rect 13593 7501 13709 7535
rect 13745 7501 13789 7535
rect 13825 7501 13869 7535
rect 13905 7501 13949 7535
rect 13985 7501 14029 7535
rect 14065 7501 14109 7535
rect 14145 7501 14313 7535
rect 14349 7501 14393 7535
rect 14429 7501 14473 7535
rect 14509 7501 14553 7535
rect 14589 7501 14633 7535
rect 14669 7501 14713 7535
rect 14749 7501 14921 7535
rect 14957 7501 15001 7535
rect 15037 7501 15081 7535
rect 15117 7501 15161 7535
rect 15197 7501 15241 7535
rect 15277 7501 15321 7535
rect 15357 7501 15525 7535
rect 15561 7501 15605 7535
rect 15641 7501 15685 7535
rect 15721 7501 15765 7535
rect 15801 7501 15845 7535
rect 15881 7501 15925 7535
rect 15961 7501 16133 7535
rect 16169 7501 16213 7535
rect 16249 7501 16293 7535
rect 16329 7501 16373 7535
rect 16409 7501 16453 7535
rect 16489 7501 16533 7535
rect 16569 7501 16737 7535
rect 16773 7501 16817 7535
rect 16853 7501 16897 7535
rect 16933 7501 16977 7535
rect 17013 7501 17057 7535
rect 17093 7501 17137 7535
rect 17173 7501 17345 7535
rect 17381 7501 17425 7535
rect 17461 7501 17505 7535
rect 17541 7501 17585 7535
rect 17621 7501 17665 7535
rect 17701 7501 17745 7535
rect 17781 7501 17949 7535
rect 17985 7501 18029 7535
rect 18065 7501 18109 7535
rect 18145 7501 18189 7535
rect 18225 7501 18269 7535
rect 18305 7501 18349 7535
rect 18385 7501 18501 7535
rect 13593 7483 18501 7501
rect 18563 7538 19241 7552
rect 18563 7504 18681 7538
rect 18717 7504 18761 7538
rect 18797 7504 18841 7538
rect 18877 7504 18921 7538
rect 18957 7504 19001 7538
rect 19037 7504 19081 7538
rect 19117 7528 19241 7538
rect 19117 7512 19275 7528
rect 19329 7588 19363 7604
rect 19624 7575 19650 7609
rect 19684 7575 19710 7609
rect 19624 7549 19710 7575
rect 20052 7586 20138 7612
rect 20052 7552 20078 7586
rect 20112 7552 20138 7586
rect 25814 7593 25871 7657
rect 25950 7650 25984 7666
rect 26038 7726 26072 7742
rect 26038 7650 26072 7666
rect 25950 7593 25984 7604
rect 25814 7588 25984 7593
rect 25814 7552 25950 7588
rect 19329 7512 19363 7528
rect 20052 7526 20138 7552
rect 20302 7535 25210 7549
rect 19117 7504 19233 7512
rect 18563 7486 19233 7504
rect 20302 7501 20418 7535
rect 20454 7501 20498 7535
rect 20534 7501 20578 7535
rect 20614 7501 20658 7535
rect 20694 7501 20738 7535
rect 20774 7501 20818 7535
rect 20854 7501 21022 7535
rect 21058 7501 21102 7535
rect 21138 7501 21182 7535
rect 21218 7501 21262 7535
rect 21298 7501 21342 7535
rect 21378 7501 21422 7535
rect 21458 7501 21630 7535
rect 21666 7501 21710 7535
rect 21746 7501 21790 7535
rect 21826 7501 21870 7535
rect 21906 7501 21950 7535
rect 21986 7501 22030 7535
rect 22066 7501 22234 7535
rect 22270 7501 22314 7535
rect 22350 7501 22394 7535
rect 22430 7501 22474 7535
rect 22510 7501 22554 7535
rect 22590 7501 22634 7535
rect 22670 7501 22842 7535
rect 22878 7501 22922 7535
rect 22958 7501 23002 7535
rect 23038 7501 23082 7535
rect 23118 7501 23162 7535
rect 23198 7501 23242 7535
rect 23278 7501 23446 7535
rect 23482 7501 23526 7535
rect 23562 7501 23606 7535
rect 23642 7501 23686 7535
rect 23722 7501 23766 7535
rect 23802 7501 23846 7535
rect 23882 7501 24054 7535
rect 24090 7501 24134 7535
rect 24170 7501 24214 7535
rect 24250 7501 24294 7535
rect 24330 7501 24374 7535
rect 24410 7501 24454 7535
rect 24490 7501 24658 7535
rect 24694 7501 24738 7535
rect 24774 7501 24818 7535
rect 24854 7501 24898 7535
rect 24934 7501 24978 7535
rect 25014 7501 25058 7535
rect 25094 7501 25210 7535
rect 20302 7483 25210 7501
rect 25272 7538 25950 7552
rect 25272 7504 25390 7538
rect 25426 7504 25470 7538
rect 25506 7504 25550 7538
rect 25586 7504 25630 7538
rect 25666 7504 25710 7538
rect 25746 7504 25790 7538
rect 25826 7528 25950 7538
rect 25826 7512 25984 7528
rect 26038 7588 26072 7604
rect 26038 7512 26072 7528
rect 25826 7504 25942 7512
rect 25272 7486 25942 7504
rect 24671 7308 25341 7326
rect 24671 7300 24787 7308
rect 24541 7284 24575 7300
rect 24541 7208 24575 7224
rect 24629 7284 24787 7300
rect 24663 7274 24787 7284
rect 24823 7274 24867 7308
rect 24903 7274 24947 7308
rect 24983 7274 25027 7308
rect 25063 7274 25107 7308
rect 25143 7274 25187 7308
rect 25223 7274 25341 7308
rect 24663 7260 25341 7274
rect 25403 7311 30311 7329
rect 25403 7277 25519 7311
rect 25555 7277 25599 7311
rect 25635 7277 25679 7311
rect 25715 7277 25759 7311
rect 25795 7277 25839 7311
rect 25875 7277 25919 7311
rect 25955 7277 26123 7311
rect 26159 7277 26203 7311
rect 26239 7277 26283 7311
rect 26319 7277 26363 7311
rect 26399 7277 26443 7311
rect 26479 7277 26523 7311
rect 26559 7277 26731 7311
rect 26767 7277 26811 7311
rect 26847 7277 26891 7311
rect 26927 7277 26971 7311
rect 27007 7277 27051 7311
rect 27087 7277 27131 7311
rect 27167 7277 27335 7311
rect 27371 7277 27415 7311
rect 27451 7277 27495 7311
rect 27531 7277 27575 7311
rect 27611 7277 27655 7311
rect 27691 7277 27735 7311
rect 27771 7277 27943 7311
rect 27979 7277 28023 7311
rect 28059 7277 28103 7311
rect 28139 7277 28183 7311
rect 28219 7277 28263 7311
rect 28299 7277 28343 7311
rect 28379 7277 28547 7311
rect 28583 7277 28627 7311
rect 28663 7277 28707 7311
rect 28743 7277 28787 7311
rect 28823 7277 28867 7311
rect 28903 7277 28947 7311
rect 28983 7277 29155 7311
rect 29191 7277 29235 7311
rect 29271 7277 29315 7311
rect 29351 7277 29395 7311
rect 29431 7277 29475 7311
rect 29511 7277 29555 7311
rect 29591 7277 29759 7311
rect 29795 7277 29839 7311
rect 29875 7277 29919 7311
rect 29955 7277 29999 7311
rect 30035 7277 30079 7311
rect 30115 7277 30159 7311
rect 30195 7277 30311 7311
rect 25403 7263 30311 7277
rect 30475 7260 30561 7286
rect 24663 7224 24799 7260
rect 24629 7219 24799 7224
rect 24629 7208 24663 7219
rect 24541 7146 24575 7162
rect 11498 7060 11527 7118
rect 11561 7060 11619 7118
rect 11653 7060 11711 7118
rect 11745 7060 11803 7118
rect 11837 7060 11895 7118
rect 11929 7060 11987 7118
rect 12021 7060 12079 7118
rect 12113 7094 12142 7118
rect 12113 7060 12171 7094
rect 12205 7060 12263 7094
rect 12297 7060 12326 7094
rect 12758 7060 12787 7118
rect 12821 7060 12879 7118
rect 12913 7060 12971 7118
rect 13005 7060 13063 7118
rect 13097 7060 13155 7118
rect 13189 7060 13247 7118
rect 13281 7060 13339 7118
rect 13373 7060 13431 7118
rect 13465 7060 13523 7118
rect 13557 7060 13615 7118
rect 13649 7060 13707 7118
rect 13741 7060 13799 7118
rect 13833 7060 13891 7118
rect 13925 7060 13983 7118
rect 14017 7060 14075 7118
rect 14109 7060 14167 7118
rect 14201 7060 14259 7118
rect 14293 7060 14351 7118
rect 14385 7060 14443 7118
rect 14477 7060 14535 7118
rect 14569 7060 14598 7118
rect 24541 7070 24575 7086
rect 24629 7146 24663 7162
rect 24742 7155 24799 7219
rect 30475 7226 30501 7260
rect 30535 7226 30561 7260
rect 30475 7200 30561 7226
rect 24629 7070 24663 7086
rect 24729 7130 24812 7155
rect 24729 7095 24754 7130
rect 24788 7095 24812 7130
rect 24729 7071 24812 7095
rect 30480 7116 30566 7142
rect 30480 7082 30506 7116
rect 30540 7082 30566 7116
rect 11531 7010 11567 7026
rect 11531 6976 11533 7010
rect 11531 6942 11567 6976
rect 11531 6908 11533 6942
rect 11603 7010 11669 7060
rect 11603 6976 11619 7010
rect 11653 6976 11669 7010
rect 11603 6942 11669 6976
rect 11603 6908 11619 6942
rect 11653 6908 11669 6942
rect 11703 7010 11757 7026
rect 11703 6976 11705 7010
rect 11739 6976 11757 7010
rect 11703 6929 11757 6976
rect 11531 6874 11567 6908
rect 11703 6895 11705 6929
rect 11739 6895 11757 6929
rect 11531 6840 11666 6874
rect 11703 6845 11757 6895
rect 11632 6811 11666 6840
rect 11519 6789 11587 6804
rect 11519 6755 11531 6789
rect 11565 6782 11587 6789
rect 11519 6748 11535 6755
rect 11569 6748 11587 6782
rect 11519 6730 11587 6748
rect 11632 6795 11687 6811
rect 11632 6761 11653 6795
rect 11632 6745 11687 6761
rect 11721 6790 11757 6845
rect 11793 7012 11859 7026
rect 11793 6978 11809 7012
rect 11843 6978 11859 7012
rect 11793 6944 11859 6978
rect 11793 6910 11809 6944
rect 11843 6910 11859 6944
rect 11793 6876 11859 6910
rect 11893 7018 11941 7060
rect 11927 6984 11941 7018
rect 11893 6950 11941 6984
rect 11927 6916 11941 6950
rect 11893 6900 11941 6916
rect 11977 6996 12011 7026
rect 11977 6901 12011 6962
rect 11793 6842 11809 6876
rect 11843 6864 11859 6876
rect 12045 7018 12111 7060
rect 12045 6984 12061 7018
rect 12095 6984 12111 7018
rect 12045 6950 12111 6984
rect 12045 6916 12061 6950
rect 12095 6916 12111 6950
rect 12045 6900 12111 6916
rect 12145 6996 12179 7026
rect 12145 6901 12179 6962
rect 11843 6842 11936 6864
rect 11793 6830 11936 6842
rect 11792 6790 11868 6796
rect 11721 6782 11868 6790
rect 11721 6752 11818 6782
rect 11632 6694 11666 6745
rect 11533 6660 11666 6694
rect 11721 6685 11757 6752
rect 11792 6748 11818 6752
rect 11852 6748 11868 6782
rect 11902 6782 11936 6830
rect 11977 6856 12011 6867
rect 12145 6856 12179 6867
rect 11977 6822 12179 6856
rect 12213 7018 12279 7060
rect 12213 6984 12229 7018
rect 12263 6984 12279 7018
rect 12213 6950 12279 6984
rect 12213 6916 12229 6950
rect 12263 6916 12279 6950
rect 12213 6882 12279 6916
rect 12213 6848 12229 6882
rect 12263 6848 12279 6882
rect 12213 6830 12279 6848
rect 12777 7018 12827 7060
rect 12777 6984 12793 7018
rect 12777 6950 12827 6984
rect 12777 6916 12793 6950
rect 12777 6882 12827 6916
rect 12777 6848 12793 6882
rect 12777 6832 12827 6848
rect 12861 7008 12926 7024
rect 12861 6974 12892 7008
rect 12861 6882 12926 6974
rect 12861 6848 12892 6882
rect 12080 6789 12179 6822
rect 12861 6794 12926 6848
rect 12960 7018 13010 7060
rect 12960 6984 12976 7018
rect 12960 6950 13010 6984
rect 12960 6916 12976 6950
rect 12960 6882 13010 6916
rect 12960 6848 12976 6882
rect 12960 6832 13010 6848
rect 13044 7008 13126 7024
rect 13044 6974 13076 7008
rect 13110 6974 13126 7008
rect 13044 6934 13126 6974
rect 13044 6900 13076 6934
rect 13110 6900 13126 6934
rect 13160 7018 13194 7060
rect 13160 6950 13194 6984
rect 13160 6900 13194 6916
rect 13228 6958 13246 6992
rect 13280 6958 13292 6992
rect 13342 6964 13358 6998
rect 13392 6964 13532 6998
rect 13044 6832 13106 6900
rect 13228 6866 13262 6958
rect 13140 6832 13262 6866
rect 13406 6924 13464 6930
rect 13406 6898 13430 6924
rect 13440 6864 13464 6890
rect 13304 6856 13372 6862
rect 13304 6832 13338 6856
rect 13044 6794 13078 6832
rect 13140 6798 13174 6832
rect 13338 6798 13372 6822
rect 11902 6748 11952 6782
rect 11986 6748 12002 6782
rect 12080 6755 12175 6789
rect 12209 6755 12219 6789
rect 12861 6786 13078 6794
rect 11902 6714 11936 6748
rect 12080 6714 12179 6755
rect 11533 6639 11567 6660
rect 11705 6656 11757 6685
rect 11533 6584 11567 6605
rect 11603 6592 11619 6626
rect 11653 6592 11669 6626
rect 11603 6550 11669 6592
rect 11739 6622 11757 6656
rect 11705 6584 11757 6622
rect 11809 6680 11936 6714
rect 11977 6680 12179 6714
rect 12861 6752 12873 6786
rect 12907 6752 13078 6786
rect 12861 6746 13078 6752
rect 11809 6662 11843 6680
rect 11977 6662 12011 6680
rect 11809 6584 11843 6628
rect 11879 6630 11927 6646
rect 11879 6596 11893 6630
rect 11879 6550 11927 6596
rect 12145 6662 12179 6680
rect 11977 6584 12011 6628
rect 12045 6630 12111 6646
rect 12045 6596 12061 6630
rect 12095 6596 12111 6630
rect 12045 6550 12111 6596
rect 12145 6584 12179 6628
rect 12213 6694 12279 6710
rect 12213 6660 12229 6694
rect 12263 6660 12279 6694
rect 12213 6626 12279 6660
rect 12213 6592 12229 6626
rect 12263 6592 12279 6626
rect 12213 6550 12279 6592
rect 12777 6694 12827 6710
rect 12777 6660 12793 6694
rect 12777 6626 12827 6660
rect 12777 6592 12793 6626
rect 12777 6550 12827 6592
rect 12861 6662 12926 6746
rect 12861 6628 12892 6662
rect 12861 6586 12926 6628
rect 12960 6694 13010 6710
rect 12960 6660 12976 6694
rect 12960 6626 13010 6660
rect 12960 6592 12976 6626
rect 12960 6550 13010 6592
rect 13044 6678 13078 6746
rect 13112 6782 13174 6798
rect 13146 6748 13174 6782
rect 13112 6732 13174 6748
rect 13208 6782 13270 6798
rect 13304 6782 13372 6798
rect 13242 6748 13270 6782
rect 13208 6732 13290 6748
rect 13406 6740 13464 6864
rect 13044 6662 13110 6678
rect 13044 6628 13076 6662
rect 13044 6586 13110 6628
rect 13144 6652 13194 6696
rect 13144 6618 13160 6652
rect 13144 6550 13194 6618
rect 13228 6649 13290 6732
rect 13340 6724 13464 6740
rect 13374 6690 13464 6724
rect 13340 6674 13464 6690
rect 13498 6880 13532 6964
rect 13577 6984 13646 7060
rect 14032 6994 14078 7060
rect 13611 6950 13646 6984
rect 13694 6958 13706 6992
rect 13740 6958 13799 6992
rect 13577 6934 13646 6950
rect 13680 6896 13718 6912
rect 13680 6880 13681 6896
rect 13498 6862 13681 6880
rect 13715 6862 13718 6896
rect 13498 6846 13718 6862
rect 13228 6615 13241 6649
rect 13275 6615 13290 6649
rect 13498 6626 13532 6846
rect 13574 6796 13648 6812
rect 13608 6790 13648 6796
rect 13574 6756 13601 6762
rect 13635 6756 13648 6790
rect 13574 6676 13648 6756
rect 13684 6650 13718 6846
rect 13228 6608 13290 6615
rect 13353 6592 13369 6626
rect 13403 6592 13532 6626
rect 13572 6626 13638 6642
rect 13572 6592 13573 6626
rect 13607 6592 13638 6626
rect 13572 6550 13638 6592
rect 13677 6634 13718 6650
rect 13711 6600 13718 6634
rect 13761 6895 13799 6958
rect 13761 6861 13765 6895
rect 13761 6652 13799 6861
rect 13795 6618 13799 6652
rect 13761 6602 13799 6618
rect 13833 6958 13890 6992
rect 13924 6958 13936 6992
rect 14032 6960 14037 6994
rect 14071 6960 14078 6994
rect 14429 7018 14495 7060
rect 30480 7056 30566 7082
rect 13833 6945 13883 6958
rect 13833 6911 13849 6945
rect 14032 6944 14078 6960
rect 14149 6958 14166 6992
rect 14200 6958 14265 6992
rect 14299 6958 14315 6992
rect 14429 6984 14445 7018
rect 14479 6984 14495 7018
rect 24541 7008 24575 7024
rect 14529 6992 14571 7008
rect 14563 6958 14571 6992
rect 13833 6895 13883 6911
rect 13833 6668 13867 6895
rect 13934 6890 13953 6924
rect 13987 6890 14003 6924
rect 13934 6865 13968 6890
rect 13914 6831 13968 6865
rect 13914 6811 13948 6831
rect 13901 6795 13948 6811
rect 14149 6814 14183 6958
rect 14529 6950 14571 6958
rect 14464 6924 14571 6950
rect 24541 6932 24575 6948
rect 24629 7008 24663 7024
rect 24629 6932 24663 6948
rect 30481 6964 30567 6990
rect 14217 6898 14258 6924
rect 14251 6890 14258 6898
rect 14292 6916 14571 6924
rect 30481 6930 30507 6964
rect 30541 6930 30567 6964
rect 14292 6890 14498 6916
rect 30481 6904 30567 6930
rect 14251 6864 14285 6890
rect 14217 6848 14285 6864
rect 13935 6761 13948 6795
rect 13901 6745 13948 6761
rect 13833 6652 13880 6668
rect 13833 6618 13846 6652
rect 13833 6602 13880 6618
rect 13914 6626 13948 6745
rect 13982 6736 14040 6797
rect 13982 6719 14003 6736
rect 14037 6702 14040 6736
rect 14016 6685 14040 6702
rect 13982 6676 14040 6685
rect 14074 6736 14115 6797
rect 14149 6780 14217 6814
rect 14074 6719 14099 6736
rect 14074 6685 14076 6719
rect 14133 6702 14149 6736
rect 14110 6685 14149 6702
rect 14074 6676 14149 6685
rect 14041 6626 14107 6642
rect 13677 6584 13718 6600
rect 13914 6592 13950 6626
rect 13984 6592 14000 6626
rect 14041 6592 14049 6626
rect 14083 6592 14107 6626
rect 14183 6640 14217 6780
rect 14251 6740 14285 6848
rect 14319 6840 14350 6856
rect 14384 6822 14396 6856
rect 14319 6790 14353 6806
rect 14251 6724 14316 6740
rect 14251 6690 14282 6724
rect 14251 6674 14316 6690
rect 14350 6736 14430 6752
rect 14350 6702 14396 6736
rect 14350 6686 14430 6702
rect 14464 6694 14498 6890
rect 14532 6856 14568 6882
rect 14532 6822 14534 6856
rect 14532 6782 14568 6822
rect 24541 6870 24575 6886
rect 24541 6794 24575 6810
rect 24629 6870 24663 6886
rect 24629 6794 24663 6810
rect 30481 6794 30567 6820
rect 14566 6748 14568 6782
rect 30481 6760 30507 6794
rect 30541 6760 30567 6794
rect 14532 6728 14568 6748
rect 24057 6713 24073 6742
rect 14350 6658 14393 6686
rect 14464 6660 14571 6694
rect 23999 6679 24028 6713
rect 24062 6708 24073 6713
rect 24107 6713 24123 6742
rect 24187 6713 24203 6742
rect 24237 6713 24257 6742
rect 24333 6713 24349 6742
rect 24107 6708 24120 6713
rect 24062 6679 24120 6708
rect 24154 6708 24203 6713
rect 24154 6679 24212 6708
rect 24246 6679 24304 6713
rect 24338 6708 24349 6713
rect 24383 6713 24403 6742
rect 24541 6732 24575 6748
rect 24383 6708 24396 6713
rect 24338 6679 24396 6708
rect 24430 6679 24459 6713
rect 14183 6606 14253 6640
rect 14287 6606 14303 6640
rect 14350 6624 14354 6658
rect 14388 6624 14393 6658
rect 14529 6652 14571 6660
rect 14350 6612 14393 6624
rect 14041 6550 14107 6592
rect 14429 6592 14445 6626
rect 14479 6592 14495 6626
rect 14563 6618 14571 6652
rect 14529 6602 14571 6618
rect 24067 6637 24109 6679
rect 24067 6603 24075 6637
rect 14429 6550 14495 6592
rect 24067 6569 24109 6603
rect 11498 6492 11527 6550
rect 11561 6492 11619 6550
rect 11653 6492 11711 6550
rect 11745 6492 11803 6550
rect 11837 6492 11895 6550
rect 11929 6492 11987 6550
rect 12021 6492 12079 6550
rect 12113 6492 12171 6550
rect 12205 6492 12263 6550
rect 12297 6531 12326 6550
rect 12758 6531 12787 6550
rect 12297 6526 12787 6531
rect 12821 6526 12879 6550
rect 12913 6526 12971 6550
rect 13005 6526 13063 6550
rect 13097 6526 13155 6550
rect 13189 6526 13247 6550
rect 13281 6526 13339 6550
rect 13373 6526 13431 6550
rect 13465 6526 13523 6550
rect 13557 6526 13615 6550
rect 13649 6526 13707 6550
rect 13741 6526 13799 6550
rect 13833 6526 13891 6550
rect 13925 6526 13983 6550
rect 14017 6526 14075 6550
rect 14109 6526 14167 6550
rect 14201 6526 14259 6550
rect 14293 6526 14351 6550
rect 14385 6526 14443 6550
rect 14477 6526 14535 6550
rect 12297 6492 12355 6526
rect 12389 6492 12447 6526
rect 12481 6492 12539 6526
rect 12573 6492 12631 6526
rect 12665 6492 12723 6526
rect 12757 6516 12787 6526
rect 12849 6516 12879 6526
rect 12941 6516 12971 6526
rect 13033 6516 13063 6526
rect 13125 6516 13155 6526
rect 13217 6516 13247 6526
rect 13309 6516 13339 6526
rect 13401 6516 13431 6526
rect 13493 6516 13523 6526
rect 13585 6516 13615 6526
rect 13677 6516 13707 6526
rect 13769 6516 13799 6526
rect 13861 6516 13891 6526
rect 13953 6516 13983 6526
rect 14045 6516 14075 6526
rect 14137 6516 14167 6526
rect 14229 6516 14259 6526
rect 14321 6516 14351 6526
rect 14413 6516 14443 6526
rect 14505 6516 14535 6526
rect 14569 6516 14599 6550
rect 12757 6492 12815 6516
rect 12849 6492 12907 6516
rect 12941 6492 12999 6516
rect 13033 6492 13091 6516
rect 13125 6492 13183 6516
rect 13217 6492 13275 6516
rect 13309 6492 13367 6516
rect 13401 6492 13459 6516
rect 13493 6492 13551 6516
rect 13585 6492 13643 6516
rect 13677 6492 13735 6516
rect 13769 6492 13827 6516
rect 13861 6492 13919 6516
rect 13953 6492 14011 6516
rect 14045 6492 14103 6516
rect 14137 6492 14195 6516
rect 14229 6492 14287 6516
rect 14321 6492 14379 6516
rect 14413 6492 14471 6516
rect 14505 6492 14599 6516
rect 24067 6535 24075 6569
rect 24067 6501 24109 6535
rect 24067 6467 24075 6501
rect 24067 6451 24109 6467
rect 24143 6637 24209 6645
rect 24143 6603 24159 6637
rect 24193 6603 24209 6637
rect 24143 6570 24209 6603
rect 24143 6536 24156 6570
rect 24190 6569 24209 6570
rect 24143 6535 24159 6536
rect 24193 6535 24209 6569
rect 24143 6501 24209 6535
rect 24143 6467 24159 6501
rect 24193 6467 24209 6501
rect 24143 6449 24209 6467
rect 24063 6405 24129 6415
rect 24063 6371 24075 6405
rect 24109 6401 24129 6405
rect 24063 6367 24079 6371
rect 24113 6367 24129 6401
rect 24063 6317 24109 6333
rect 24163 6329 24209 6449
rect 24063 6283 24075 6317
rect 24063 6249 24109 6283
rect 11497 6187 11526 6245
rect 11560 6187 11618 6245
rect 11652 6187 11710 6245
rect 11744 6187 11802 6245
rect 11836 6187 11894 6245
rect 11928 6187 11986 6245
rect 12020 6187 12078 6245
rect 12112 6187 12170 6245
rect 12204 6187 12262 6245
rect 12296 6187 12354 6245
rect 12388 6187 12446 6245
rect 12480 6187 12538 6245
rect 12572 6187 12630 6245
rect 12664 6187 12722 6245
rect 12756 6187 12814 6245
rect 12848 6187 12906 6245
rect 12940 6187 12998 6245
rect 13032 6187 13090 6245
rect 13124 6187 13182 6245
rect 13216 6187 13274 6245
rect 13308 6236 13550 6245
rect 13308 6221 13397 6236
rect 13431 6221 13550 6236
rect 13308 6187 13366 6221
rect 13431 6202 13458 6221
rect 13400 6187 13458 6202
rect 13492 6187 13550 6221
rect 13584 6187 13642 6245
rect 13676 6187 13734 6245
rect 13768 6187 13826 6245
rect 13860 6187 13918 6245
rect 13952 6187 14010 6245
rect 14044 6221 14103 6245
rect 14044 6187 14102 6221
rect 14137 6211 14194 6245
rect 14136 6187 14194 6211
rect 14228 6187 14286 6245
rect 14320 6187 14378 6245
rect 14412 6187 14470 6245
rect 14504 6239 14746 6245
rect 14504 6221 14640 6239
rect 14674 6221 14746 6239
rect 14504 6187 14562 6221
rect 14596 6205 14640 6221
rect 14596 6187 14654 6205
rect 14688 6187 14746 6221
rect 14780 6187 14838 6245
rect 14872 6187 14930 6245
rect 14964 6187 15022 6245
rect 15056 6187 15114 6245
rect 15148 6187 15206 6245
rect 15240 6187 15298 6245
rect 15332 6187 15390 6245
rect 15424 6187 15482 6245
rect 15516 6187 15574 6245
rect 15608 6187 15666 6245
rect 15700 6187 15758 6245
rect 15792 6187 15850 6245
rect 15884 6187 15942 6245
rect 15976 6187 16034 6245
rect 16068 6187 16126 6245
rect 16160 6187 16218 6245
rect 16252 6187 16310 6245
rect 16344 6187 16402 6245
rect 16436 6187 16494 6245
rect 16528 6187 16586 6245
rect 16620 6187 16678 6245
rect 16712 6187 16770 6245
rect 16804 6187 16862 6245
rect 16896 6241 17138 6245
rect 16896 6221 17032 6241
rect 17066 6221 17138 6241
rect 16896 6187 16954 6221
rect 16988 6207 17032 6221
rect 16988 6187 17046 6207
rect 17080 6187 17138 6221
rect 17172 6187 17230 6245
rect 17264 6187 17322 6245
rect 17356 6187 17414 6245
rect 17448 6187 17506 6245
rect 17540 6187 17598 6245
rect 17632 6187 17690 6245
rect 17724 6187 17782 6245
rect 17816 6187 17874 6245
rect 17908 6187 17966 6245
rect 18000 6187 18058 6245
rect 18092 6187 18150 6245
rect 18184 6187 18242 6245
rect 18276 6187 18334 6245
rect 18368 6187 18426 6245
rect 18460 6187 18518 6245
rect 18552 6187 18610 6245
rect 18644 6187 18702 6245
rect 18736 6187 18794 6245
rect 18828 6187 18886 6245
rect 18920 6187 18978 6245
rect 19012 6187 19070 6245
rect 19104 6187 19162 6245
rect 19196 6187 19254 6245
rect 19288 6241 19530 6245
rect 19288 6221 19424 6241
rect 19458 6221 19530 6241
rect 19288 6187 19346 6221
rect 19380 6207 19424 6221
rect 19380 6187 19438 6207
rect 19472 6187 19530 6221
rect 19564 6187 19622 6245
rect 19656 6187 19714 6245
rect 19748 6187 19806 6245
rect 19840 6187 19898 6245
rect 19932 6187 19990 6245
rect 20024 6187 20082 6245
rect 20116 6187 20174 6245
rect 20208 6187 20266 6245
rect 20300 6187 20358 6245
rect 20392 6187 20450 6245
rect 20484 6187 20542 6245
rect 20576 6187 20634 6245
rect 20668 6187 20726 6245
rect 20760 6187 20818 6245
rect 20852 6187 20910 6245
rect 20944 6187 21002 6245
rect 21036 6187 21094 6245
rect 21128 6187 21186 6245
rect 21220 6187 21278 6245
rect 21312 6187 21370 6245
rect 21404 6187 21462 6245
rect 21496 6187 21554 6245
rect 21588 6187 21646 6245
rect 21680 6242 21922 6245
rect 21680 6221 21816 6242
rect 21850 6221 21922 6242
rect 21680 6187 21738 6221
rect 21772 6208 21816 6221
rect 21772 6187 21830 6208
rect 21864 6187 21922 6221
rect 21956 6187 22014 6245
rect 22048 6187 22106 6245
rect 22140 6187 22198 6245
rect 22232 6187 22290 6245
rect 22324 6187 22382 6245
rect 22416 6187 22474 6245
rect 22508 6187 22566 6245
rect 22600 6187 22658 6245
rect 22692 6187 22750 6245
rect 22784 6187 22842 6245
rect 22876 6187 22934 6245
rect 22968 6187 23026 6245
rect 23060 6187 23118 6245
rect 23152 6187 23210 6245
rect 23244 6187 23302 6245
rect 23336 6187 23394 6245
rect 23428 6187 23457 6245
rect 24063 6215 24075 6249
rect 11514 6137 11566 6153
rect 11514 6103 11532 6137
rect 11514 6069 11566 6103
rect 11600 6121 11666 6187
rect 11600 6087 11616 6121
rect 11650 6087 11666 6121
rect 11700 6137 11745 6153
rect 11734 6103 11745 6137
rect 11514 6035 11532 6069
rect 11700 6069 11745 6103
rect 11784 6121 11854 6187
rect 11784 6087 11804 6121
rect 11838 6087 11854 6121
rect 11888 6137 11922 6153
rect 11965 6110 11981 6144
rect 12015 6110 12131 6144
rect 11566 6051 11665 6053
rect 11566 6035 11619 6051
rect 11514 6019 11619 6035
rect 11653 6017 11665 6051
rect 11514 5924 11585 5985
rect 11514 5890 11529 5924
rect 11563 5900 11585 5924
rect 11514 5866 11530 5890
rect 11564 5866 11585 5900
rect 11514 5855 11585 5866
rect 11619 5924 11665 6017
rect 11619 5890 11631 5924
rect 11619 5821 11665 5890
rect 11514 5787 11665 5821
rect 11734 6035 11745 6069
rect 11888 6053 11922 6103
rect 11700 5847 11745 6035
rect 11700 5813 11711 5847
rect 11514 5779 11566 5787
rect 11514 5745 11532 5779
rect 11700 5779 11745 5813
rect 11779 6019 11922 6053
rect 11779 5825 11813 6019
rect 11963 6017 11987 6051
rect 12021 6025 12063 6051
rect 12021 6017 12029 6025
rect 11963 5991 12029 6017
rect 11847 5980 11929 5985
rect 11847 5946 11891 5980
rect 11925 5946 11929 5980
rect 11847 5911 11929 5946
rect 11881 5877 11929 5911
rect 11847 5861 11929 5877
rect 11963 5975 12063 5991
rect 11963 5851 12007 5975
rect 12097 5941 12131 6110
rect 12179 6135 12255 6187
rect 12473 6145 12539 6187
rect 12179 6101 12195 6135
rect 12229 6101 12255 6135
rect 12315 6119 12349 6135
rect 12315 6067 12349 6085
rect 12473 6111 12489 6145
rect 12523 6111 12539 6145
rect 12962 6145 13038 6187
rect 12473 6077 12539 6111
rect 12748 6110 12764 6144
rect 12798 6110 12914 6144
rect 12962 6111 12978 6145
rect 13012 6111 13038 6145
rect 13226 6145 13503 6187
rect 13086 6119 13120 6135
rect 12165 6051 12435 6067
rect 12165 6025 12315 6051
rect 12199 6017 12315 6025
rect 12349 6017 12435 6051
rect 12473 6043 12489 6077
rect 12523 6043 12539 6077
rect 12710 6051 12757 6057
rect 12199 5991 12215 6017
rect 12165 5975 12215 5991
rect 12317 5941 12367 5957
rect 12097 5907 12333 5941
rect 12097 5899 12177 5907
rect 11779 5787 11922 5825
rect 11997 5817 12007 5851
rect 11963 5801 12007 5817
rect 12043 5829 12059 5863
rect 12093 5847 12109 5863
rect 12043 5813 12075 5829
rect 12043 5789 12109 5813
rect 11514 5729 11566 5745
rect 11600 5719 11616 5753
rect 11650 5719 11666 5753
rect 11734 5745 11745 5779
rect 11888 5771 11922 5787
rect 11700 5729 11745 5745
rect 11600 5677 11666 5719
rect 11784 5719 11804 5753
rect 11838 5719 11854 5753
rect 12143 5753 12177 5899
rect 12323 5891 12367 5907
rect 12401 5873 12435 6017
rect 12710 6025 12723 6051
rect 12744 5991 12757 6017
rect 12469 5983 12670 5991
rect 12469 5949 12631 5983
rect 12665 5949 12670 5983
rect 12710 5975 12757 5991
rect 12805 6025 12846 6041
rect 12805 5991 12812 6025
rect 12469 5943 12670 5949
rect 12469 5941 12535 5943
rect 12469 5907 12485 5941
rect 12519 5907 12535 5941
rect 12805 5921 12846 5991
rect 12722 5915 12846 5921
rect 12597 5873 12613 5907
rect 12647 5873 12663 5907
rect 12215 5839 12231 5873
rect 12265 5853 12281 5873
rect 12265 5847 12297 5853
rect 12215 5813 12263 5839
rect 12401 5839 12663 5873
rect 12722 5881 12723 5915
rect 12757 5885 12846 5915
rect 12880 5941 12914 6110
rect 13226 6111 13242 6145
rect 13276 6111 13453 6145
rect 13487 6111 13503 6145
rect 13086 6077 13120 6085
rect 13537 6108 13594 6153
rect 12948 6043 13503 6077
rect 12948 6025 12998 6043
rect 12982 5991 12998 6025
rect 12948 5975 12998 5991
rect 12880 5925 13150 5941
rect 12880 5907 13116 5925
rect 12757 5881 12779 5885
rect 12722 5851 12779 5881
rect 12401 5813 12445 5839
rect 12215 5807 12297 5813
rect 12379 5779 12395 5813
rect 12429 5779 12445 5813
rect 12722 5817 12745 5851
rect 12479 5787 12513 5803
rect 12722 5801 12779 5817
rect 11888 5721 11922 5737
rect 11784 5677 11854 5719
rect 11978 5719 11994 5753
rect 12028 5719 12177 5753
rect 11978 5713 12177 5719
rect 12211 5749 12245 5765
rect 12211 5677 12245 5715
rect 12279 5735 12295 5769
rect 12329 5745 12345 5769
rect 12880 5753 12914 5907
rect 13106 5891 13116 5907
rect 13106 5875 13150 5891
rect 12989 5847 13008 5873
rect 12989 5813 12999 5847
rect 13042 5839 13064 5873
rect 13033 5813 13064 5839
rect 13184 5816 13220 6043
rect 12989 5807 13064 5813
rect 13154 5813 13220 5816
rect 13154 5779 13170 5813
rect 13204 5779 13220 5813
rect 13254 5983 13356 6009
rect 13254 5949 13275 5983
rect 13309 5975 13356 5983
rect 13390 5975 13406 6009
rect 13254 5941 13309 5949
rect 13288 5907 13309 5941
rect 13469 5925 13503 6043
rect 13571 6074 13594 6108
rect 13537 6040 13594 6074
rect 13571 6006 13594 6040
rect 13537 5986 13594 6006
rect 13254 5845 13309 5907
rect 13360 5913 13435 5925
rect 13360 5879 13385 5913
rect 13419 5879 13435 5913
rect 13469 5909 13519 5925
rect 13469 5875 13485 5909
rect 13469 5859 13519 5875
rect 13254 5811 13392 5845
rect 12479 5745 12513 5753
rect 12329 5735 12513 5745
rect 12279 5711 12513 5735
rect 12567 5719 12583 5753
rect 12617 5719 12633 5753
rect 12567 5677 12633 5719
rect 12761 5719 12777 5753
rect 12811 5719 12914 5753
rect 12761 5713 12914 5719
rect 12950 5749 13002 5765
rect 12950 5715 12968 5749
rect 12950 5677 13002 5715
rect 13054 5735 13070 5769
rect 13104 5745 13120 5769
rect 13254 5761 13288 5777
rect 13104 5735 13254 5745
rect 13054 5727 13254 5735
rect 13054 5711 13288 5727
rect 13345 5763 13392 5811
rect 13345 5729 13358 5763
rect 13345 5713 13392 5729
rect 13437 5753 13503 5821
rect 13553 5803 13594 5986
rect 13437 5719 13453 5753
rect 13487 5719 13503 5753
rect 13437 5677 13503 5719
rect 13537 5789 13594 5803
rect 13537 5787 13550 5789
rect 13584 5755 13594 5789
rect 13571 5753 13594 5755
rect 13537 5711 13594 5753
rect 13628 6127 13691 6143
rect 13628 6093 13641 6127
rect 13675 6093 13691 6127
rect 13628 6059 13691 6093
rect 13628 6025 13641 6059
rect 13675 6025 13691 6059
rect 13628 5925 13691 6025
rect 13727 6133 13786 6187
rect 13727 6099 13736 6133
rect 13770 6099 13786 6133
rect 13727 6065 13786 6099
rect 13727 6031 13736 6065
rect 13770 6031 13786 6065
rect 13727 6013 13786 6031
rect 13820 6109 13872 6153
rect 13854 6075 13872 6109
rect 13820 6041 13872 6075
rect 13854 6007 13872 6041
rect 13906 6137 13958 6153
rect 13906 6103 13924 6137
rect 13906 6069 13958 6103
rect 13992 6121 14058 6187
rect 13992 6087 14008 6121
rect 14042 6087 14058 6121
rect 14092 6137 14137 6153
rect 14126 6103 14137 6137
rect 13906 6035 13924 6069
rect 14092 6069 14137 6103
rect 14176 6121 14246 6187
rect 14176 6087 14196 6121
rect 14230 6087 14246 6121
rect 14280 6137 14314 6153
rect 14357 6110 14373 6144
rect 14407 6110 14523 6144
rect 13958 6051 14057 6053
rect 13958 6035 14011 6051
rect 13906 6019 14011 6035
rect 13820 5987 13872 6007
rect 13820 5953 13831 5987
rect 13865 5953 13872 5987
rect 14045 6017 14057 6051
rect 13820 5949 13872 5953
rect 13628 5909 13795 5925
rect 13628 5875 13761 5909
rect 13628 5859 13795 5875
rect 13628 5779 13691 5859
rect 13829 5825 13872 5949
rect 13906 5924 13977 5985
rect 13906 5900 13921 5924
rect 13906 5866 13920 5900
rect 13955 5890 13977 5924
rect 13954 5866 13977 5890
rect 13906 5855 13977 5866
rect 14011 5924 14057 6017
rect 14011 5890 14023 5924
rect 13628 5745 13641 5779
rect 13675 5745 13691 5779
rect 13820 5789 13872 5825
rect 14011 5821 14057 5890
rect 13628 5711 13691 5745
rect 13727 5753 13786 5769
rect 13727 5719 13736 5753
rect 13770 5719 13786 5753
rect 13727 5677 13786 5719
rect 13854 5755 13872 5789
rect 13820 5711 13872 5755
rect 13906 5787 14057 5821
rect 14126 6035 14137 6069
rect 14280 6053 14314 6103
rect 14092 5847 14137 6035
rect 14092 5813 14103 5847
rect 13906 5779 13958 5787
rect 13906 5745 13924 5779
rect 14092 5779 14137 5813
rect 14171 6019 14314 6053
rect 14171 5825 14205 6019
rect 14355 6017 14379 6051
rect 14413 6025 14455 6051
rect 14413 6017 14421 6025
rect 14355 5991 14421 6017
rect 14239 5983 14321 5985
rect 14239 5949 14242 5983
rect 14276 5949 14321 5983
rect 14239 5911 14321 5949
rect 14273 5877 14321 5911
rect 14239 5861 14321 5877
rect 14355 5975 14455 5991
rect 14355 5851 14399 5975
rect 14489 5941 14523 6110
rect 14571 6135 14647 6187
rect 14865 6145 14931 6187
rect 14571 6101 14587 6135
rect 14621 6101 14647 6135
rect 14707 6119 14741 6135
rect 14707 6067 14741 6085
rect 14865 6111 14881 6145
rect 14915 6111 14931 6145
rect 15354 6145 15430 6187
rect 14865 6077 14931 6111
rect 15140 6110 15156 6144
rect 15190 6110 15306 6144
rect 15354 6111 15370 6145
rect 15404 6111 15430 6145
rect 15618 6145 15895 6187
rect 15478 6119 15512 6135
rect 14557 6051 14827 6067
rect 14557 6025 14707 6051
rect 14591 6017 14707 6025
rect 14741 6017 14827 6051
rect 14865 6043 14881 6077
rect 14915 6043 14931 6077
rect 15102 6051 15149 6057
rect 14591 5991 14607 6017
rect 14557 5975 14607 5991
rect 14709 5941 14759 5957
rect 14489 5907 14725 5941
rect 14489 5899 14569 5907
rect 14171 5787 14314 5825
rect 14389 5817 14399 5851
rect 14355 5801 14399 5817
rect 14435 5829 14451 5863
rect 14485 5847 14501 5863
rect 14435 5813 14467 5829
rect 14435 5789 14501 5813
rect 13906 5729 13958 5745
rect 13992 5719 14008 5753
rect 14042 5719 14058 5753
rect 14126 5745 14137 5779
rect 14280 5771 14314 5787
rect 14092 5729 14137 5745
rect 13992 5677 14058 5719
rect 14176 5719 14196 5753
rect 14230 5719 14246 5753
rect 14535 5753 14569 5899
rect 14715 5891 14759 5907
rect 14793 5873 14827 6017
rect 15102 6025 15115 6051
rect 15136 5991 15149 6017
rect 14861 5983 15062 5991
rect 14861 5949 15023 5983
rect 15057 5949 15062 5983
rect 15102 5975 15149 5991
rect 15197 6025 15238 6041
rect 15197 5991 15204 6025
rect 14861 5943 15062 5949
rect 14861 5941 14927 5943
rect 14861 5907 14877 5941
rect 14911 5907 14927 5941
rect 15197 5921 15238 5991
rect 15114 5915 15238 5921
rect 14989 5873 15005 5907
rect 15039 5873 15055 5907
rect 14607 5839 14623 5873
rect 14657 5853 14673 5873
rect 14657 5847 14689 5853
rect 14607 5813 14655 5839
rect 14793 5839 15055 5873
rect 15114 5881 15115 5915
rect 15149 5885 15238 5915
rect 15272 5941 15306 6110
rect 15618 6111 15634 6145
rect 15668 6111 15845 6145
rect 15879 6111 15895 6145
rect 15478 6077 15512 6085
rect 15929 6108 15986 6153
rect 15340 6043 15895 6077
rect 15340 6025 15390 6043
rect 15374 5991 15390 6025
rect 15340 5975 15390 5991
rect 15272 5925 15542 5941
rect 15272 5907 15508 5925
rect 15149 5881 15171 5885
rect 15114 5851 15171 5881
rect 14793 5813 14837 5839
rect 14607 5807 14689 5813
rect 14771 5779 14787 5813
rect 14821 5779 14837 5813
rect 15114 5817 15137 5851
rect 14871 5787 14905 5803
rect 15114 5801 15171 5817
rect 14280 5721 14314 5737
rect 14176 5677 14246 5719
rect 14370 5719 14386 5753
rect 14420 5719 14569 5753
rect 14370 5713 14569 5719
rect 14603 5749 14637 5765
rect 14603 5677 14637 5715
rect 14671 5735 14687 5769
rect 14721 5745 14737 5769
rect 15272 5753 15306 5907
rect 15498 5891 15508 5907
rect 15498 5875 15542 5891
rect 15381 5847 15400 5873
rect 15381 5813 15391 5847
rect 15434 5839 15456 5873
rect 15425 5813 15456 5839
rect 15576 5816 15612 6043
rect 15381 5807 15456 5813
rect 15546 5813 15612 5816
rect 15546 5779 15562 5813
rect 15596 5779 15612 5813
rect 15646 5983 15748 6009
rect 15646 5949 15667 5983
rect 15701 5975 15748 5983
rect 15782 5975 15798 6009
rect 15646 5941 15701 5949
rect 15680 5907 15701 5941
rect 15861 5925 15895 6043
rect 15963 6074 15986 6108
rect 15929 6040 15986 6074
rect 15963 6006 15986 6040
rect 15929 5986 15986 6006
rect 15646 5845 15701 5907
rect 15752 5917 15827 5925
rect 15752 5883 15768 5917
rect 15802 5913 15827 5917
rect 15752 5879 15777 5883
rect 15811 5879 15827 5913
rect 15861 5909 15911 5925
rect 15861 5875 15877 5909
rect 15861 5859 15911 5875
rect 15646 5811 15784 5845
rect 14871 5745 14905 5753
rect 14721 5735 14905 5745
rect 14671 5711 14905 5735
rect 14959 5719 14975 5753
rect 15009 5719 15025 5753
rect 14959 5677 15025 5719
rect 15153 5719 15169 5753
rect 15203 5719 15306 5753
rect 15153 5713 15306 5719
rect 15342 5749 15394 5765
rect 15342 5715 15360 5749
rect 15342 5677 15394 5715
rect 15446 5735 15462 5769
rect 15496 5745 15512 5769
rect 15646 5761 15680 5777
rect 15496 5735 15646 5745
rect 15446 5727 15646 5735
rect 15446 5711 15680 5727
rect 15737 5763 15784 5811
rect 15737 5729 15750 5763
rect 15737 5713 15784 5729
rect 15829 5753 15895 5821
rect 15945 5803 15986 5986
rect 15829 5719 15845 5753
rect 15879 5719 15895 5753
rect 15829 5677 15895 5719
rect 15929 5800 15986 5803
rect 15929 5787 15939 5800
rect 15973 5766 15986 5800
rect 15963 5753 15986 5766
rect 15929 5711 15986 5753
rect 16020 6127 16083 6143
rect 16020 6093 16033 6127
rect 16067 6093 16083 6127
rect 16020 6059 16083 6093
rect 16020 6025 16033 6059
rect 16067 6025 16083 6059
rect 16020 5925 16083 6025
rect 16119 6133 16178 6187
rect 16119 6099 16128 6133
rect 16162 6099 16178 6133
rect 16119 6065 16178 6099
rect 16119 6031 16128 6065
rect 16162 6031 16178 6065
rect 16119 6013 16178 6031
rect 16212 6109 16264 6153
rect 16246 6075 16264 6109
rect 16212 6041 16264 6075
rect 16246 6007 16264 6041
rect 16298 6137 16350 6153
rect 16298 6103 16316 6137
rect 16298 6069 16350 6103
rect 16384 6121 16450 6187
rect 16384 6087 16400 6121
rect 16434 6087 16450 6121
rect 16484 6137 16529 6153
rect 16518 6103 16529 6137
rect 16298 6035 16316 6069
rect 16484 6069 16529 6103
rect 16568 6121 16638 6187
rect 16568 6087 16588 6121
rect 16622 6087 16638 6121
rect 16672 6137 16706 6153
rect 16749 6110 16765 6144
rect 16799 6110 16915 6144
rect 16350 6051 16449 6053
rect 16350 6035 16403 6051
rect 16298 6019 16403 6035
rect 16212 5986 16264 6007
rect 16212 5952 16220 5986
rect 16254 5952 16264 5986
rect 16437 6017 16449 6051
rect 16212 5949 16264 5952
rect 16020 5909 16187 5925
rect 16020 5875 16153 5909
rect 16020 5859 16187 5875
rect 16020 5779 16083 5859
rect 16221 5825 16264 5949
rect 16298 5924 16369 5985
rect 16298 5867 16313 5924
rect 16347 5867 16369 5924
rect 16298 5855 16369 5867
rect 16403 5924 16449 6017
rect 16403 5890 16415 5924
rect 16212 5812 16264 5825
rect 16403 5821 16449 5890
rect 16020 5745 16033 5779
rect 16067 5745 16083 5779
rect 16245 5789 16264 5812
rect 16020 5711 16083 5745
rect 16119 5753 16178 5769
rect 16119 5719 16128 5753
rect 16162 5719 16178 5753
rect 16119 5677 16178 5719
rect 16246 5755 16264 5789
rect 16212 5711 16264 5755
rect 16298 5787 16449 5821
rect 16518 6035 16529 6069
rect 16672 6053 16706 6103
rect 16484 5847 16529 6035
rect 16484 5813 16495 5847
rect 16298 5779 16350 5787
rect 16298 5745 16316 5779
rect 16484 5779 16529 5813
rect 16563 6019 16706 6053
rect 16563 5825 16597 6019
rect 16747 6017 16771 6051
rect 16805 6025 16847 6051
rect 16805 6017 16813 6025
rect 16747 5991 16813 6017
rect 16631 5982 16713 5985
rect 16665 5948 16713 5982
rect 16631 5911 16713 5948
rect 16665 5877 16713 5911
rect 16631 5861 16713 5877
rect 16747 5975 16847 5991
rect 16747 5851 16791 5975
rect 16881 5941 16915 6110
rect 16963 6135 17039 6187
rect 17257 6145 17323 6187
rect 16963 6101 16979 6135
rect 17013 6101 17039 6135
rect 17099 6119 17133 6135
rect 17099 6067 17133 6085
rect 17257 6111 17273 6145
rect 17307 6111 17323 6145
rect 17746 6145 17822 6187
rect 17257 6077 17323 6111
rect 17532 6110 17548 6144
rect 17582 6110 17698 6144
rect 17746 6111 17762 6145
rect 17796 6111 17822 6145
rect 18010 6145 18287 6187
rect 17870 6119 17904 6135
rect 16949 6051 17219 6067
rect 16949 6025 17099 6051
rect 16983 6017 17099 6025
rect 17133 6017 17219 6051
rect 17257 6043 17273 6077
rect 17307 6043 17323 6077
rect 17494 6051 17541 6057
rect 16983 5991 16999 6017
rect 16949 5975 16999 5991
rect 17101 5941 17151 5957
rect 16881 5907 17117 5941
rect 16881 5899 16961 5907
rect 16563 5787 16706 5825
rect 16781 5817 16791 5851
rect 16747 5801 16791 5817
rect 16827 5829 16843 5863
rect 16877 5847 16893 5863
rect 16827 5813 16859 5829
rect 16827 5789 16893 5813
rect 16298 5729 16350 5745
rect 16384 5719 16400 5753
rect 16434 5719 16450 5753
rect 16518 5745 16529 5779
rect 16672 5771 16706 5787
rect 16484 5729 16529 5745
rect 16384 5677 16450 5719
rect 16568 5719 16588 5753
rect 16622 5719 16638 5753
rect 16927 5753 16961 5899
rect 17107 5891 17151 5907
rect 17185 5873 17219 6017
rect 17494 6025 17507 6051
rect 17528 5991 17541 6017
rect 17253 5983 17454 5991
rect 17253 5949 17415 5983
rect 17449 5949 17454 5983
rect 17494 5975 17541 5991
rect 17589 6025 17630 6041
rect 17589 5991 17596 6025
rect 17253 5943 17454 5949
rect 17253 5941 17319 5943
rect 17253 5907 17269 5941
rect 17303 5907 17319 5941
rect 17589 5921 17630 5991
rect 17506 5915 17630 5921
rect 17381 5873 17397 5907
rect 17431 5873 17447 5907
rect 16999 5839 17015 5873
rect 17049 5853 17065 5873
rect 17049 5847 17081 5853
rect 16999 5813 17047 5839
rect 17185 5839 17447 5873
rect 17506 5881 17507 5915
rect 17541 5885 17630 5915
rect 17664 5941 17698 6110
rect 18010 6111 18026 6145
rect 18060 6111 18237 6145
rect 18271 6111 18287 6145
rect 17870 6077 17904 6085
rect 18321 6108 18378 6153
rect 17732 6043 18287 6077
rect 17732 6025 17782 6043
rect 17766 5991 17782 6025
rect 17732 5975 17782 5991
rect 17664 5925 17934 5941
rect 17664 5907 17900 5925
rect 17541 5881 17563 5885
rect 17506 5851 17563 5881
rect 17185 5813 17229 5839
rect 16999 5807 17081 5813
rect 17163 5779 17179 5813
rect 17213 5779 17229 5813
rect 17506 5817 17529 5851
rect 17263 5787 17297 5803
rect 17506 5801 17563 5817
rect 16672 5721 16706 5737
rect 16568 5677 16638 5719
rect 16762 5719 16778 5753
rect 16812 5719 16961 5753
rect 16762 5713 16961 5719
rect 16995 5749 17029 5765
rect 16995 5677 17029 5715
rect 17063 5735 17079 5769
rect 17113 5745 17129 5769
rect 17664 5753 17698 5907
rect 17890 5891 17900 5907
rect 17890 5875 17934 5891
rect 17773 5847 17792 5873
rect 17773 5813 17783 5847
rect 17826 5839 17848 5873
rect 17817 5813 17848 5839
rect 17968 5816 18004 6043
rect 17773 5807 17848 5813
rect 17938 5813 18004 5816
rect 17938 5779 17954 5813
rect 17988 5779 18004 5813
rect 18038 5983 18140 6009
rect 18038 5949 18059 5983
rect 18093 5975 18140 5983
rect 18174 5975 18190 6009
rect 18038 5941 18093 5949
rect 18072 5907 18093 5941
rect 18253 5925 18287 6043
rect 18355 6074 18378 6108
rect 18321 6040 18378 6074
rect 18355 6006 18378 6040
rect 18321 5986 18378 6006
rect 18038 5845 18093 5907
rect 18144 5918 18219 5925
rect 18144 5884 18158 5918
rect 18192 5913 18219 5918
rect 18144 5879 18169 5884
rect 18203 5879 18219 5913
rect 18253 5909 18303 5925
rect 18253 5875 18269 5909
rect 18253 5859 18303 5875
rect 18038 5811 18176 5845
rect 17263 5745 17297 5753
rect 17113 5735 17297 5745
rect 17063 5711 17297 5735
rect 17351 5719 17367 5753
rect 17401 5719 17417 5753
rect 17351 5677 17417 5719
rect 17545 5719 17561 5753
rect 17595 5719 17698 5753
rect 17545 5713 17698 5719
rect 17734 5749 17786 5765
rect 17734 5715 17752 5749
rect 17734 5677 17786 5715
rect 17838 5735 17854 5769
rect 17888 5745 17904 5769
rect 18038 5761 18072 5777
rect 17888 5735 18038 5745
rect 17838 5727 18038 5735
rect 17838 5711 18072 5727
rect 18129 5763 18176 5811
rect 18129 5729 18142 5763
rect 18129 5713 18176 5729
rect 18221 5753 18287 5821
rect 18337 5803 18378 5986
rect 18221 5719 18237 5753
rect 18271 5719 18287 5753
rect 18221 5677 18287 5719
rect 18321 5787 18327 5803
rect 18361 5769 18378 5803
rect 18355 5753 18378 5769
rect 18321 5711 18378 5753
rect 18412 6127 18475 6143
rect 18412 6093 18425 6127
rect 18459 6093 18475 6127
rect 18412 6059 18475 6093
rect 18412 6025 18425 6059
rect 18459 6025 18475 6059
rect 18412 5925 18475 6025
rect 18511 6133 18570 6187
rect 18511 6099 18520 6133
rect 18554 6099 18570 6133
rect 18511 6065 18570 6099
rect 18511 6031 18520 6065
rect 18554 6031 18570 6065
rect 18511 6013 18570 6031
rect 18604 6109 18656 6153
rect 18638 6075 18656 6109
rect 18604 6041 18656 6075
rect 18638 6007 18656 6041
rect 18690 6137 18742 6153
rect 18690 6103 18708 6137
rect 18690 6069 18742 6103
rect 18776 6121 18842 6187
rect 18776 6087 18792 6121
rect 18826 6087 18842 6121
rect 18876 6137 18921 6153
rect 18910 6103 18921 6137
rect 18690 6035 18708 6069
rect 18876 6069 18921 6103
rect 18960 6121 19030 6187
rect 18960 6087 18980 6121
rect 19014 6087 19030 6121
rect 19064 6137 19098 6153
rect 19141 6110 19157 6144
rect 19191 6110 19307 6144
rect 18742 6051 18841 6053
rect 18742 6035 18795 6051
rect 18690 6019 18795 6035
rect 18604 5984 18656 6007
rect 18829 6017 18841 6051
rect 18604 5950 18615 5984
rect 18649 5950 18656 5984
rect 18604 5949 18656 5950
rect 18412 5909 18579 5925
rect 18412 5875 18545 5909
rect 18412 5859 18579 5875
rect 18412 5779 18475 5859
rect 18613 5825 18656 5949
rect 18690 5924 18761 5985
rect 18690 5866 18705 5924
rect 18739 5866 18761 5924
rect 18690 5855 18761 5866
rect 18795 5924 18841 6017
rect 18795 5890 18807 5924
rect 18412 5745 18425 5779
rect 18459 5745 18475 5779
rect 18604 5801 18656 5825
rect 18795 5821 18841 5890
rect 18604 5789 18607 5801
rect 18412 5711 18475 5745
rect 18511 5753 18570 5769
rect 18511 5719 18520 5753
rect 18554 5719 18570 5753
rect 18511 5677 18570 5719
rect 18641 5767 18656 5801
rect 18638 5755 18656 5767
rect 18604 5711 18656 5755
rect 18690 5787 18841 5821
rect 18910 6035 18921 6069
rect 19064 6053 19098 6103
rect 18876 5847 18921 6035
rect 18876 5813 18887 5847
rect 18690 5779 18742 5787
rect 18690 5745 18708 5779
rect 18876 5779 18921 5813
rect 18955 6019 19098 6053
rect 18955 5825 18989 6019
rect 19139 6017 19163 6051
rect 19197 6025 19239 6051
rect 19197 6017 19205 6025
rect 19139 5991 19205 6017
rect 19023 5980 19105 5985
rect 19023 5946 19026 5980
rect 19060 5946 19105 5980
rect 19023 5911 19105 5946
rect 19057 5877 19105 5911
rect 19023 5861 19105 5877
rect 19139 5975 19239 5991
rect 19139 5851 19183 5975
rect 19273 5941 19307 6110
rect 19355 6135 19431 6187
rect 19649 6145 19715 6187
rect 19355 6101 19371 6135
rect 19405 6101 19431 6135
rect 19491 6119 19525 6135
rect 19491 6067 19525 6085
rect 19649 6111 19665 6145
rect 19699 6111 19715 6145
rect 20138 6145 20214 6187
rect 19649 6077 19715 6111
rect 19924 6110 19940 6144
rect 19974 6110 20090 6144
rect 20138 6111 20154 6145
rect 20188 6111 20214 6145
rect 20402 6145 20679 6187
rect 20262 6119 20296 6135
rect 19341 6051 19611 6067
rect 19341 6025 19491 6051
rect 19375 6017 19491 6025
rect 19525 6017 19611 6051
rect 19649 6043 19665 6077
rect 19699 6043 19715 6077
rect 19886 6051 19933 6057
rect 19375 5991 19391 6017
rect 19341 5975 19391 5991
rect 19493 5941 19543 5957
rect 19273 5907 19509 5941
rect 19273 5899 19353 5907
rect 18955 5787 19098 5825
rect 19173 5817 19183 5851
rect 19139 5801 19183 5817
rect 19219 5829 19235 5863
rect 19269 5847 19285 5863
rect 19219 5813 19251 5829
rect 19219 5789 19285 5813
rect 18690 5729 18742 5745
rect 18776 5719 18792 5753
rect 18826 5719 18842 5753
rect 18910 5745 18921 5779
rect 19064 5771 19098 5787
rect 18876 5729 18921 5745
rect 18776 5677 18842 5719
rect 18960 5719 18980 5753
rect 19014 5719 19030 5753
rect 19319 5753 19353 5899
rect 19499 5891 19543 5907
rect 19577 5873 19611 6017
rect 19886 6025 19899 6051
rect 19920 5991 19933 6017
rect 19645 5983 19846 5991
rect 19645 5949 19807 5983
rect 19841 5949 19846 5983
rect 19886 5975 19933 5991
rect 19981 6025 20022 6041
rect 19981 5991 19988 6025
rect 19645 5943 19846 5949
rect 19645 5941 19711 5943
rect 19645 5907 19661 5941
rect 19695 5907 19711 5941
rect 19981 5921 20022 5991
rect 19898 5915 20022 5921
rect 19773 5873 19789 5907
rect 19823 5873 19839 5907
rect 19391 5839 19407 5873
rect 19441 5853 19457 5873
rect 19441 5847 19473 5853
rect 19391 5813 19439 5839
rect 19577 5839 19839 5873
rect 19898 5881 19899 5915
rect 19933 5885 20022 5915
rect 20056 5941 20090 6110
rect 20402 6111 20418 6145
rect 20452 6111 20629 6145
rect 20663 6111 20679 6145
rect 20262 6077 20296 6085
rect 20713 6108 20770 6153
rect 20124 6043 20679 6077
rect 20124 6025 20174 6043
rect 20158 5991 20174 6025
rect 20124 5975 20174 5991
rect 20056 5925 20326 5941
rect 20056 5907 20292 5925
rect 19933 5881 19955 5885
rect 19898 5851 19955 5881
rect 19577 5813 19621 5839
rect 19391 5807 19473 5813
rect 19555 5779 19571 5813
rect 19605 5779 19621 5813
rect 19898 5817 19921 5851
rect 19655 5787 19689 5803
rect 19898 5801 19955 5817
rect 19064 5721 19098 5737
rect 18960 5677 19030 5719
rect 19154 5719 19170 5753
rect 19204 5719 19353 5753
rect 19154 5713 19353 5719
rect 19387 5749 19421 5765
rect 19387 5677 19421 5715
rect 19455 5735 19471 5769
rect 19505 5745 19521 5769
rect 20056 5753 20090 5907
rect 20282 5891 20292 5907
rect 20282 5875 20326 5891
rect 20165 5847 20184 5873
rect 20165 5813 20175 5847
rect 20218 5839 20240 5873
rect 20209 5813 20240 5839
rect 20360 5816 20396 6043
rect 20165 5807 20240 5813
rect 20330 5813 20396 5816
rect 20330 5779 20346 5813
rect 20380 5779 20396 5813
rect 20430 5983 20532 6009
rect 20430 5949 20451 5983
rect 20485 5975 20532 5983
rect 20566 5975 20582 6009
rect 20430 5941 20485 5949
rect 20464 5907 20485 5941
rect 20645 5925 20679 6043
rect 20747 6074 20770 6108
rect 20713 6040 20770 6074
rect 20747 6006 20770 6040
rect 20713 5986 20770 6006
rect 20430 5845 20485 5907
rect 20536 5920 20611 5925
rect 20536 5886 20549 5920
rect 20583 5913 20611 5920
rect 20536 5879 20561 5886
rect 20595 5879 20611 5913
rect 20645 5909 20695 5925
rect 20645 5875 20661 5909
rect 20645 5859 20695 5875
rect 20430 5811 20568 5845
rect 19655 5745 19689 5753
rect 19505 5735 19689 5745
rect 19455 5711 19689 5735
rect 19743 5719 19759 5753
rect 19793 5719 19809 5753
rect 19743 5677 19809 5719
rect 19937 5719 19953 5753
rect 19987 5719 20090 5753
rect 19937 5713 20090 5719
rect 20126 5749 20178 5765
rect 20126 5715 20144 5749
rect 20126 5677 20178 5715
rect 20230 5735 20246 5769
rect 20280 5745 20296 5769
rect 20430 5761 20464 5777
rect 20280 5735 20430 5745
rect 20230 5727 20430 5735
rect 20230 5711 20464 5727
rect 20521 5763 20568 5811
rect 20521 5729 20534 5763
rect 20521 5713 20568 5729
rect 20613 5753 20679 5821
rect 20729 5803 20770 5986
rect 20613 5719 20629 5753
rect 20663 5719 20679 5753
rect 20613 5677 20679 5719
rect 20713 5787 20770 5803
rect 20747 5786 20770 5787
rect 20713 5752 20724 5753
rect 20758 5752 20770 5786
rect 20713 5711 20770 5752
rect 20804 6127 20867 6143
rect 20804 6093 20817 6127
rect 20851 6093 20867 6127
rect 20804 6059 20867 6093
rect 20804 6025 20817 6059
rect 20851 6025 20867 6059
rect 20804 5925 20867 6025
rect 20903 6133 20962 6187
rect 20903 6099 20912 6133
rect 20946 6099 20962 6133
rect 20903 6065 20962 6099
rect 20903 6031 20912 6065
rect 20946 6031 20962 6065
rect 20903 6013 20962 6031
rect 20996 6109 21048 6153
rect 21030 6075 21048 6109
rect 20996 6041 21048 6075
rect 21030 6007 21048 6041
rect 21082 6137 21134 6153
rect 21082 6103 21100 6137
rect 21082 6069 21134 6103
rect 21168 6121 21234 6187
rect 21168 6087 21184 6121
rect 21218 6087 21234 6121
rect 21268 6137 21313 6153
rect 21302 6103 21313 6137
rect 21082 6035 21100 6069
rect 21268 6069 21313 6103
rect 21352 6121 21422 6187
rect 21352 6087 21372 6121
rect 21406 6087 21422 6121
rect 21456 6137 21490 6153
rect 21533 6110 21549 6144
rect 21583 6110 21699 6144
rect 21134 6051 21233 6053
rect 21134 6035 21187 6051
rect 21082 6019 21187 6035
rect 20996 5983 21048 6007
rect 21221 6017 21233 6051
rect 20996 5949 21006 5983
rect 21040 5949 21048 5983
rect 20804 5909 20971 5925
rect 20804 5875 20937 5909
rect 20804 5859 20971 5875
rect 20804 5779 20867 5859
rect 21005 5825 21048 5949
rect 21082 5924 21153 5985
rect 21082 5890 21097 5924
rect 21131 5902 21153 5924
rect 21082 5868 21100 5890
rect 21134 5868 21153 5902
rect 21082 5855 21153 5868
rect 21187 5924 21233 6017
rect 21187 5890 21199 5924
rect 20804 5745 20817 5779
rect 20851 5745 20867 5779
rect 20996 5817 21048 5825
rect 21187 5821 21233 5890
rect 20996 5789 21007 5817
rect 21041 5783 21048 5817
rect 20804 5711 20867 5745
rect 20903 5753 20962 5769
rect 20903 5719 20912 5753
rect 20946 5719 20962 5753
rect 20903 5677 20962 5719
rect 21030 5755 21048 5783
rect 20996 5711 21048 5755
rect 21082 5787 21233 5821
rect 21302 6035 21313 6069
rect 21456 6053 21490 6103
rect 21268 5847 21313 6035
rect 21268 5813 21279 5847
rect 21082 5779 21134 5787
rect 21082 5745 21100 5779
rect 21268 5779 21313 5813
rect 21347 6019 21490 6053
rect 21347 5825 21381 6019
rect 21531 6017 21555 6051
rect 21589 6025 21631 6051
rect 21589 6017 21597 6025
rect 21531 5991 21597 6017
rect 21415 5979 21497 5985
rect 21415 5945 21417 5979
rect 21451 5945 21497 5979
rect 21415 5911 21497 5945
rect 21449 5877 21497 5911
rect 21415 5861 21497 5877
rect 21531 5975 21631 5991
rect 21531 5851 21575 5975
rect 21665 5941 21699 6110
rect 21747 6135 21823 6187
rect 22041 6145 22107 6187
rect 21747 6101 21763 6135
rect 21797 6101 21823 6135
rect 21883 6119 21917 6135
rect 21883 6067 21917 6085
rect 22041 6111 22057 6145
rect 22091 6111 22107 6145
rect 22530 6145 22606 6187
rect 22041 6077 22107 6111
rect 22316 6110 22332 6144
rect 22366 6110 22482 6144
rect 22530 6111 22546 6145
rect 22580 6111 22606 6145
rect 22794 6145 23071 6187
rect 22654 6119 22688 6135
rect 21733 6051 22003 6067
rect 21733 6025 21883 6051
rect 21767 6017 21883 6025
rect 21917 6017 22003 6051
rect 22041 6043 22057 6077
rect 22091 6043 22107 6077
rect 22278 6051 22325 6057
rect 21767 5991 21783 6017
rect 21733 5975 21783 5991
rect 21885 5941 21935 5957
rect 21665 5907 21901 5941
rect 21665 5899 21745 5907
rect 21347 5787 21490 5825
rect 21565 5817 21575 5851
rect 21531 5801 21575 5817
rect 21611 5829 21627 5863
rect 21661 5847 21677 5863
rect 21611 5813 21643 5829
rect 21611 5789 21677 5813
rect 21082 5729 21134 5745
rect 21168 5719 21184 5753
rect 21218 5719 21234 5753
rect 21302 5745 21313 5779
rect 21456 5771 21490 5787
rect 21268 5729 21313 5745
rect 21168 5677 21234 5719
rect 21352 5719 21372 5753
rect 21406 5719 21422 5753
rect 21711 5753 21745 5899
rect 21891 5891 21935 5907
rect 21969 5873 22003 6017
rect 22278 6025 22291 6051
rect 22312 5991 22325 6017
rect 22037 5983 22238 5991
rect 22037 5949 22199 5983
rect 22233 5949 22238 5983
rect 22278 5975 22325 5991
rect 22373 6025 22414 6041
rect 22373 5991 22380 6025
rect 22037 5943 22238 5949
rect 22037 5941 22103 5943
rect 22037 5907 22053 5941
rect 22087 5907 22103 5941
rect 22373 5921 22414 5991
rect 22290 5915 22414 5921
rect 22165 5873 22181 5907
rect 22215 5873 22231 5907
rect 21783 5839 21799 5873
rect 21833 5853 21849 5873
rect 21833 5847 21865 5853
rect 21783 5813 21831 5839
rect 21969 5839 22231 5873
rect 22290 5881 22291 5915
rect 22325 5885 22414 5915
rect 22448 5941 22482 6110
rect 22794 6111 22810 6145
rect 22844 6111 23021 6145
rect 23055 6111 23071 6145
rect 22654 6077 22688 6085
rect 23105 6108 23162 6153
rect 22516 6043 23071 6077
rect 22516 6025 22566 6043
rect 22550 5991 22566 6025
rect 22516 5975 22566 5991
rect 22448 5925 22718 5941
rect 22448 5907 22684 5925
rect 22325 5881 22347 5885
rect 22290 5851 22347 5881
rect 21969 5813 22013 5839
rect 21783 5807 21865 5813
rect 21947 5779 21963 5813
rect 21997 5779 22013 5813
rect 22290 5817 22313 5851
rect 22047 5787 22081 5803
rect 22290 5801 22347 5817
rect 21456 5721 21490 5737
rect 21352 5677 21422 5719
rect 21546 5719 21562 5753
rect 21596 5719 21745 5753
rect 21546 5713 21745 5719
rect 21779 5749 21813 5765
rect 21779 5677 21813 5715
rect 21847 5735 21863 5769
rect 21897 5745 21913 5769
rect 22448 5753 22482 5907
rect 22674 5891 22684 5907
rect 22674 5875 22718 5891
rect 22557 5847 22576 5873
rect 22557 5813 22567 5847
rect 22610 5839 22632 5873
rect 22601 5813 22632 5839
rect 22752 5816 22788 6043
rect 22557 5807 22632 5813
rect 22722 5813 22788 5816
rect 22722 5779 22738 5813
rect 22772 5779 22788 5813
rect 22822 5983 22924 6009
rect 22822 5949 22843 5983
rect 22877 5975 22924 5983
rect 22958 5975 22974 6009
rect 22822 5941 22877 5949
rect 22856 5907 22877 5941
rect 23037 5925 23071 6043
rect 23139 6074 23162 6108
rect 23105 6040 23162 6074
rect 23139 6006 23162 6040
rect 23105 5986 23162 6006
rect 22822 5845 22877 5907
rect 22928 5918 23003 5925
rect 22928 5884 22940 5918
rect 22974 5913 23003 5918
rect 22928 5879 22953 5884
rect 22987 5879 23003 5913
rect 23037 5909 23087 5925
rect 23037 5875 23053 5909
rect 23037 5859 23087 5875
rect 22822 5811 22960 5845
rect 22047 5745 22081 5753
rect 21897 5735 22081 5745
rect 21847 5711 22081 5735
rect 22135 5719 22151 5753
rect 22185 5719 22201 5753
rect 22135 5677 22201 5719
rect 22329 5719 22345 5753
rect 22379 5719 22482 5753
rect 22329 5713 22482 5719
rect 22518 5749 22570 5765
rect 22518 5715 22536 5749
rect 22518 5677 22570 5715
rect 22622 5735 22638 5769
rect 22672 5745 22688 5769
rect 22822 5761 22856 5777
rect 22672 5735 22822 5745
rect 22622 5727 22822 5735
rect 22622 5711 22856 5727
rect 22913 5763 22960 5811
rect 22913 5729 22926 5763
rect 22913 5713 22960 5729
rect 23005 5753 23071 5821
rect 23121 5803 23162 5986
rect 23005 5719 23021 5753
rect 23055 5719 23071 5753
rect 23005 5677 23071 5719
rect 23105 5787 23162 5803
rect 23149 5753 23162 5787
rect 23105 5711 23162 5753
rect 23196 6127 23259 6143
rect 23196 6093 23209 6127
rect 23243 6093 23259 6127
rect 23196 6059 23259 6093
rect 23196 6025 23209 6059
rect 23243 6025 23259 6059
rect 23196 5925 23259 6025
rect 23295 6133 23354 6187
rect 24063 6169 24109 6215
rect 24143 6317 24209 6329
rect 24143 6283 24159 6317
rect 24193 6283 24209 6317
rect 24143 6249 24209 6283
rect 24143 6215 24159 6249
rect 24193 6215 24209 6249
rect 24143 6203 24209 6215
rect 24249 6637 24315 6645
rect 24249 6603 24265 6637
rect 24299 6603 24315 6637
rect 24249 6569 24315 6603
rect 24249 6535 24265 6569
rect 24299 6535 24315 6569
rect 24249 6515 24315 6535
rect 24249 6467 24265 6515
rect 24299 6467 24315 6515
rect 24249 6449 24315 6467
rect 24349 6637 24391 6679
rect 24541 6656 24575 6672
rect 24629 6732 24663 6748
rect 30481 6734 30567 6760
rect 24629 6656 24663 6672
rect 24383 6603 24391 6637
rect 30480 6637 30566 6663
rect 24349 6569 24391 6603
rect 24383 6535 24391 6569
rect 24349 6501 24391 6535
rect 24541 6594 24575 6610
rect 24541 6518 24575 6534
rect 24629 6594 24663 6610
rect 30480 6603 30506 6637
rect 30540 6603 30566 6637
rect 30480 6577 30566 6603
rect 24629 6518 24663 6534
rect 24383 6467 24391 6501
rect 24349 6451 24391 6467
rect 24249 6329 24295 6449
rect 24569 6441 24585 6475
rect 24619 6441 24635 6475
rect 24329 6404 24395 6415
rect 24329 6401 24349 6404
rect 24329 6367 24345 6401
rect 24383 6370 24395 6404
rect 24379 6367 24395 6370
rect 24479 6405 24528 6417
rect 24479 6371 24488 6405
rect 24522 6400 24528 6405
rect 24522 6371 24811 6400
rect 24479 6365 24811 6371
rect 24479 6358 24528 6365
rect 24776 6342 24811 6365
rect 30679 6369 31048 6371
rect 24249 6317 24315 6329
rect 24249 6283 24265 6317
rect 24299 6283 24315 6317
rect 24249 6249 24315 6283
rect 24249 6215 24265 6249
rect 24299 6215 24315 6249
rect 24249 6203 24315 6215
rect 24349 6317 24395 6333
rect 24776 6330 24825 6342
rect 24383 6283 24395 6317
rect 24349 6249 24395 6283
rect 24517 6312 24566 6324
rect 24517 6278 24526 6312
rect 24560 6278 24727 6312
rect 24776 6296 24785 6330
rect 24819 6296 24825 6330
rect 30679 6302 30708 6369
rect 30742 6336 30891 6369
rect 30925 6336 31048 6369
rect 30742 6302 30800 6336
rect 30834 6335 30891 6336
rect 30834 6302 30892 6335
rect 30926 6302 30984 6336
rect 31018 6335 31048 6336
rect 31018 6302 31047 6335
rect 24776 6283 24825 6296
rect 30326 6283 30360 6299
rect 24517 6265 24566 6278
rect 24383 6215 24395 6249
rect 24349 6169 24395 6215
rect 24686 6236 24727 6278
rect 24777 6237 24826 6249
rect 24777 6236 24786 6237
rect 24686 6203 24786 6236
rect 24820 6203 24826 6237
rect 24686 6202 24826 6203
rect 24777 6190 24826 6202
rect 25211 6198 25227 6232
rect 25261 6198 25277 6232
rect 25943 6201 25959 6235
rect 25993 6201 26009 6235
rect 26069 6201 26085 6235
rect 26119 6201 26135 6235
rect 27155 6201 27171 6235
rect 27205 6201 27221 6235
rect 27281 6201 27297 6235
rect 27331 6201 27347 6235
rect 28367 6201 28383 6235
rect 28417 6201 28433 6235
rect 28493 6201 28509 6235
rect 28543 6201 28559 6235
rect 29579 6201 29595 6235
rect 29629 6201 29645 6235
rect 29705 6201 29721 6235
rect 29755 6201 29771 6235
rect 30326 6207 30360 6223
rect 30414 6283 30448 6299
rect 30414 6207 30448 6223
rect 30714 6252 30748 6268
rect 30714 6184 30748 6218
rect 23295 6099 23304 6133
rect 23338 6099 23354 6133
rect 23295 6065 23354 6099
rect 23295 6031 23304 6065
rect 23338 6031 23354 6065
rect 23295 6013 23354 6031
rect 23388 6109 23440 6153
rect 23999 6135 24028 6169
rect 24062 6140 24120 6169
rect 24154 6140 24212 6169
rect 24062 6135 24093 6140
rect 24154 6135 24211 6140
rect 24246 6135 24304 6169
rect 24338 6140 24396 6169
rect 24338 6135 24355 6140
rect 23422 6107 23440 6109
rect 23388 6073 23394 6075
rect 23428 6073 23440 6107
rect 24077 6106 24093 6135
rect 24127 6106 24153 6135
rect 24195 6106 24211 6135
rect 24245 6106 24271 6135
rect 24337 6106 24355 6135
rect 24389 6135 24396 6140
rect 24430 6135 24459 6169
rect 25183 6139 25217 6155
rect 24389 6106 24405 6135
rect 23388 6041 23440 6073
rect 25183 6063 25217 6079
rect 25271 6142 25305 6158
rect 25271 6066 25305 6082
rect 25915 6142 25949 6158
rect 25915 6066 25949 6082
rect 26020 6142 26054 6158
rect 26020 6066 26054 6082
rect 26129 6142 26163 6158
rect 26129 6066 26163 6082
rect 27127 6142 27161 6158
rect 27127 6066 27161 6082
rect 27231 6142 27265 6158
rect 27231 6066 27265 6082
rect 27341 6142 27375 6158
rect 27341 6066 27375 6082
rect 28339 6142 28373 6158
rect 28339 6066 28373 6082
rect 28444 6142 28478 6158
rect 28444 6066 28478 6082
rect 28553 6142 28587 6158
rect 28553 6066 28587 6082
rect 29551 6142 29585 6158
rect 29551 6066 29585 6082
rect 29658 6142 29692 6158
rect 29658 6066 29692 6082
rect 29765 6142 29799 6158
rect 29765 6066 29799 6082
rect 30326 6145 30360 6161
rect 30326 6069 30360 6085
rect 30414 6145 30448 6161
rect 30414 6069 30448 6085
rect 30510 6145 30544 6161
rect 30510 6069 30544 6085
rect 30606 6145 30640 6161
rect 30606 6069 30640 6085
rect 30791 6252 30857 6302
rect 30791 6218 30807 6252
rect 30841 6218 30857 6252
rect 30791 6184 30857 6218
rect 30791 6150 30807 6184
rect 30841 6150 30857 6184
rect 30891 6236 30942 6268
rect 30891 6202 30893 6236
rect 30927 6202 30942 6236
rect 30891 6155 30942 6202
rect 30714 6116 30748 6150
rect 30891 6121 30893 6155
rect 30927 6121 30942 6155
rect 30714 6082 30857 6116
rect 30891 6087 30942 6121
rect 23422 6007 23440 6041
rect 23388 5949 23440 6007
rect 30239 5994 30255 6028
rect 30289 5994 30305 6028
rect 30696 6026 30767 6046
rect 30446 5992 30462 6026
rect 30496 5992 30512 6026
rect 30696 5992 30702 6026
rect 30736 6024 30767 6026
rect 30696 5990 30716 5992
rect 30750 5990 30767 6024
rect 30696 5972 30767 5990
rect 30823 6040 30857 6082
rect 30823 6024 30874 6040
rect 30823 5990 30840 6024
rect 30823 5974 30874 5990
rect 30908 6026 30942 6087
rect 30977 6260 31029 6302
rect 31011 6226 31029 6260
rect 30977 6192 31029 6226
rect 31011 6158 31029 6192
rect 30977 6124 31029 6158
rect 31011 6090 31029 6124
rect 30977 6072 31029 6090
rect 30908 5992 30909 6026
rect 23196 5909 23363 5925
rect 23196 5875 23329 5909
rect 23196 5859 23363 5875
rect 23196 5779 23259 5859
rect 23397 5825 23440 5949
rect 25536 5941 25570 5957
rect 25536 5865 25570 5881
rect 25626 5941 25660 5957
rect 25626 5865 25660 5881
rect 26268 5941 26302 5957
rect 26268 5865 26302 5881
rect 26375 5941 26409 5957
rect 26375 5865 26409 5881
rect 26478 5941 26512 5957
rect 26478 5865 26512 5881
rect 27480 5941 27514 5957
rect 27480 5865 27514 5881
rect 27586 5941 27620 5957
rect 27586 5865 27620 5881
rect 27690 5941 27724 5957
rect 27690 5865 27724 5881
rect 28818 5941 28852 5957
rect 28818 5865 28852 5881
rect 28926 5941 28960 5957
rect 28926 5865 28960 5881
rect 29028 5941 29062 5957
rect 29028 5865 29062 5881
rect 29673 5941 29707 5957
rect 29673 5865 29707 5881
rect 29762 5941 29796 5957
rect 29762 5865 29796 5881
rect 30326 5942 30360 5958
rect 30326 5866 30360 5882
rect 30414 5942 30448 5958
rect 30414 5866 30448 5882
rect 30510 5942 30544 5958
rect 30510 5866 30544 5882
rect 30606 5942 30640 5958
rect 30823 5936 30857 5974
rect 30908 5941 30942 5992
rect 30606 5866 30640 5882
rect 30714 5902 30857 5936
rect 30714 5881 30748 5902
rect 30891 5898 30942 5941
rect 23196 5745 23209 5779
rect 23243 5745 23259 5779
rect 23388 5817 23440 5825
rect 23388 5789 23402 5817
rect 23436 5783 23440 5817
rect 24580 5807 24596 5841
rect 24630 5807 24646 5841
rect 25564 5797 25580 5831
rect 25614 5797 25630 5831
rect 26296 5797 26312 5831
rect 26346 5797 26362 5831
rect 26418 5797 26434 5831
rect 26468 5797 26484 5831
rect 27508 5797 27524 5831
rect 27558 5797 27574 5831
rect 27630 5797 27646 5831
rect 27680 5797 27696 5831
rect 28846 5797 28862 5831
rect 28896 5797 28912 5831
rect 28968 5797 28984 5831
rect 29018 5797 29034 5831
rect 29702 5797 29718 5831
rect 29752 5797 29768 5831
rect 30714 5826 30748 5847
rect 30791 5834 30807 5868
rect 30841 5834 30857 5868
rect 30326 5804 30360 5820
rect 23196 5711 23259 5745
rect 23295 5753 23354 5769
rect 23295 5719 23304 5753
rect 23338 5719 23354 5753
rect 23295 5677 23354 5719
rect 23422 5755 23440 5783
rect 23388 5711 23440 5755
rect 24516 5757 24550 5773
rect 24516 5681 24550 5697
rect 24676 5757 24710 5773
rect 30326 5728 30360 5744
rect 30414 5804 30448 5820
rect 30791 5792 30857 5834
rect 30891 5864 30893 5898
rect 30927 5864 30942 5898
rect 30891 5826 30942 5864
rect 30977 5940 31029 5960
rect 31011 5906 31029 5940
rect 30977 5872 31029 5906
rect 31011 5838 31029 5872
rect 30977 5792 31029 5838
rect 30679 5758 30708 5792
rect 30742 5758 30800 5792
rect 30414 5728 30448 5744
rect 30680 5757 30800 5758
rect 30680 5723 30708 5757
rect 30742 5724 30800 5757
rect 30834 5724 30892 5792
rect 30926 5758 30984 5792
rect 31018 5758 31047 5792
rect 30926 5724 30985 5758
rect 31019 5724 31049 5758
rect 30742 5723 31049 5724
rect 30680 5722 31049 5723
rect 24676 5681 24710 5697
rect 11497 5619 11526 5677
rect 11560 5619 11618 5677
rect 11652 5619 11710 5677
rect 11744 5619 11802 5677
rect 11836 5619 11894 5677
rect 11928 5619 11986 5677
rect 12020 5619 12078 5677
rect 12112 5619 12170 5677
rect 12204 5619 12262 5677
rect 12296 5619 12354 5677
rect 12388 5619 12446 5677
rect 12480 5619 12538 5677
rect 12572 5619 12630 5677
rect 12664 5619 12722 5677
rect 12756 5619 12814 5677
rect 12848 5619 12906 5677
rect 12940 5619 12998 5677
rect 13032 5619 13090 5677
rect 13124 5619 13182 5677
rect 13216 5619 13274 5677
rect 13308 5619 13366 5677
rect 13400 5619 13458 5677
rect 13492 5619 13550 5677
rect 13584 5619 13642 5677
rect 13676 5619 13734 5677
rect 13768 5619 13826 5677
rect 13860 5619 13918 5677
rect 13952 5619 14010 5677
rect 14044 5619 14102 5677
rect 14136 5619 14194 5677
rect 14228 5619 14286 5677
rect 14320 5619 14378 5677
rect 14412 5619 14470 5677
rect 14504 5619 14562 5677
rect 14596 5619 14654 5677
rect 14688 5619 14746 5677
rect 14780 5619 14838 5677
rect 14872 5619 14930 5677
rect 14964 5619 15022 5677
rect 15056 5619 15114 5677
rect 15148 5619 15206 5677
rect 15240 5619 15298 5677
rect 15332 5619 15390 5677
rect 15424 5619 15482 5677
rect 15516 5619 15574 5677
rect 15608 5619 15666 5677
rect 15700 5619 15758 5677
rect 15792 5619 15850 5677
rect 15884 5619 15942 5677
rect 15976 5619 16034 5677
rect 16068 5619 16126 5677
rect 16160 5619 16218 5677
rect 16252 5619 16310 5677
rect 16344 5619 16402 5677
rect 16436 5619 16494 5677
rect 16528 5619 16586 5677
rect 16620 5619 16678 5677
rect 16712 5619 16770 5677
rect 16804 5619 16862 5677
rect 16896 5619 16954 5677
rect 16988 5619 17046 5677
rect 17080 5619 17138 5677
rect 17172 5619 17230 5677
rect 17264 5619 17322 5677
rect 17356 5619 17414 5677
rect 17448 5619 17506 5677
rect 17540 5619 17598 5677
rect 17632 5619 17690 5677
rect 17724 5619 17782 5677
rect 17816 5619 17874 5677
rect 17908 5619 17966 5677
rect 18000 5619 18058 5677
rect 18092 5619 18150 5677
rect 18184 5619 18242 5677
rect 18276 5619 18334 5677
rect 18368 5619 18426 5677
rect 18460 5619 18518 5677
rect 18552 5619 18610 5677
rect 18644 5619 18702 5677
rect 18736 5619 18794 5677
rect 18828 5619 18886 5677
rect 18920 5619 18978 5677
rect 19012 5619 19070 5677
rect 19104 5619 19162 5677
rect 19196 5619 19254 5677
rect 19288 5619 19346 5677
rect 19380 5619 19438 5677
rect 19472 5619 19530 5677
rect 19564 5619 19622 5677
rect 19656 5619 19714 5677
rect 19748 5619 19806 5677
rect 19840 5619 19898 5677
rect 19932 5619 19990 5677
rect 20024 5619 20082 5677
rect 20116 5619 20174 5677
rect 20208 5619 20266 5677
rect 20300 5619 20358 5677
rect 20392 5619 20450 5677
rect 20484 5619 20542 5677
rect 20576 5619 20634 5677
rect 20668 5619 20726 5677
rect 20760 5619 20818 5677
rect 20852 5619 20910 5677
rect 20944 5619 21002 5677
rect 21036 5619 21094 5677
rect 21128 5619 21186 5677
rect 21220 5619 21278 5677
rect 21312 5619 21370 5677
rect 21404 5619 21462 5677
rect 21496 5619 21554 5677
rect 21588 5619 21646 5677
rect 21680 5619 21738 5677
rect 21772 5619 21830 5677
rect 21864 5619 21922 5677
rect 21956 5619 22014 5677
rect 22048 5619 22106 5677
rect 22140 5619 22198 5677
rect 22232 5619 22290 5677
rect 22324 5619 22382 5677
rect 22416 5619 22474 5677
rect 22508 5619 22566 5677
rect 22600 5619 22658 5677
rect 22692 5619 22750 5677
rect 22784 5619 22842 5677
rect 22876 5619 22934 5677
rect 22968 5619 23026 5677
rect 23060 5619 23118 5677
rect 23152 5619 23210 5677
rect 23244 5619 23302 5677
rect 23336 5619 23394 5677
rect 23428 5619 23457 5677
rect 24516 5619 24550 5635
rect 11057 5498 11086 5556
rect 11120 5498 11178 5556
rect 11212 5498 11270 5556
rect 11304 5498 11362 5556
rect 11396 5498 11454 5556
rect 11488 5498 11546 5556
rect 11580 5498 11638 5556
rect 11672 5498 11730 5556
rect 11764 5498 11822 5556
rect 11856 5532 11914 5556
rect 11948 5532 12006 5556
rect 12040 5532 12098 5556
rect 12132 5532 12190 5556
rect 12224 5532 12282 5556
rect 12316 5532 12374 5556
rect 12408 5532 12466 5556
rect 12500 5532 12558 5556
rect 12592 5532 12650 5556
rect 12684 5532 12742 5556
rect 11856 5498 11894 5532
rect 11948 5522 11986 5532
rect 12040 5522 12078 5532
rect 12132 5522 12170 5532
rect 12224 5522 12262 5532
rect 12316 5522 12354 5532
rect 12408 5522 12446 5532
rect 12500 5522 12538 5532
rect 12592 5522 12630 5532
rect 12684 5522 12722 5532
rect 12776 5522 12814 5556
rect 12868 5522 12906 5556
rect 11928 5498 11986 5522
rect 12020 5498 12078 5522
rect 12112 5498 12170 5522
rect 12204 5498 12262 5522
rect 12296 5498 12354 5522
rect 12388 5498 12446 5522
rect 12480 5498 12538 5522
rect 12572 5498 12630 5522
rect 12664 5498 12722 5522
rect 12756 5498 12814 5522
rect 12848 5498 12906 5522
rect 12940 5498 12998 5556
rect 13032 5498 13090 5556
rect 13124 5498 13182 5556
rect 13216 5498 13274 5556
rect 13308 5498 13366 5556
rect 13400 5498 13458 5556
rect 13492 5498 13550 5556
rect 13584 5498 13642 5556
rect 13676 5498 13734 5556
rect 13768 5498 13826 5556
rect 13860 5498 13918 5556
rect 13952 5498 14010 5556
rect 14044 5498 14102 5556
rect 14136 5498 14194 5556
rect 14228 5498 14286 5556
rect 14320 5498 14378 5556
rect 14412 5498 14470 5556
rect 14504 5498 14562 5556
rect 14596 5553 14838 5556
rect 14596 5532 14711 5553
rect 14596 5498 14654 5532
rect 14688 5519 14711 5532
rect 14745 5532 14838 5553
rect 14745 5519 14746 5532
rect 14688 5498 14746 5519
rect 14780 5498 14838 5532
rect 14872 5498 14930 5556
rect 14964 5498 15022 5556
rect 15056 5498 15114 5556
rect 15148 5498 15206 5556
rect 15240 5498 15298 5556
rect 15332 5498 15390 5556
rect 15424 5498 15482 5556
rect 15516 5498 15574 5556
rect 15608 5498 15666 5556
rect 15700 5498 15758 5556
rect 15792 5498 15850 5556
rect 15884 5498 15942 5556
rect 15976 5498 16034 5556
rect 16068 5498 16126 5556
rect 16160 5498 16218 5556
rect 16252 5498 16310 5556
rect 16344 5498 16402 5556
rect 16436 5498 16494 5556
rect 16528 5498 16586 5556
rect 16620 5498 16678 5556
rect 16712 5498 16770 5556
rect 16804 5498 16862 5556
rect 16896 5498 16954 5556
rect 16988 5553 17230 5556
rect 16988 5532 17103 5553
rect 16988 5498 17046 5532
rect 17080 5519 17103 5532
rect 17137 5532 17230 5553
rect 17137 5519 17138 5532
rect 17080 5498 17138 5519
rect 17172 5498 17230 5532
rect 17264 5498 17322 5556
rect 17356 5498 17414 5556
rect 17448 5498 17506 5556
rect 17540 5498 17598 5556
rect 17632 5498 17690 5556
rect 17724 5498 17782 5556
rect 17816 5498 17874 5556
rect 17908 5498 17966 5556
rect 18000 5498 18058 5556
rect 18092 5498 18150 5556
rect 18184 5498 18242 5556
rect 18276 5498 18334 5556
rect 18368 5498 18426 5556
rect 18460 5498 18518 5556
rect 18552 5498 18610 5556
rect 18644 5498 18702 5556
rect 18736 5498 18794 5556
rect 18828 5498 18886 5556
rect 18920 5498 18978 5556
rect 19012 5498 19070 5556
rect 19104 5498 19162 5556
rect 19196 5498 19254 5556
rect 19288 5498 19346 5556
rect 19380 5553 19622 5556
rect 19380 5532 19495 5553
rect 19380 5498 19438 5532
rect 19472 5519 19495 5532
rect 19529 5532 19622 5553
rect 19529 5519 19530 5532
rect 19472 5498 19530 5519
rect 19564 5498 19622 5532
rect 19656 5498 19714 5556
rect 19748 5498 19806 5556
rect 19840 5498 19898 5556
rect 19932 5498 19990 5556
rect 20024 5498 20082 5556
rect 20116 5498 20174 5556
rect 20208 5498 20266 5556
rect 20300 5498 20358 5556
rect 20392 5498 20450 5556
rect 20484 5498 20542 5556
rect 20576 5498 20634 5556
rect 20668 5498 20726 5556
rect 20760 5498 20818 5556
rect 20852 5498 20910 5556
rect 20944 5498 21002 5556
rect 21036 5498 21094 5556
rect 21128 5498 21186 5556
rect 21220 5498 21278 5556
rect 21312 5498 21370 5556
rect 21404 5498 21462 5556
rect 21496 5498 21554 5556
rect 21588 5498 21646 5556
rect 21680 5498 21738 5556
rect 21772 5553 22014 5556
rect 21772 5532 21887 5553
rect 21772 5498 21830 5532
rect 21864 5519 21887 5532
rect 21921 5532 22014 5553
rect 21921 5519 21922 5532
rect 21864 5498 21922 5519
rect 21956 5498 22014 5532
rect 22048 5498 22106 5556
rect 22140 5498 22198 5556
rect 22232 5498 22290 5556
rect 22324 5498 22382 5556
rect 22416 5498 22474 5556
rect 22508 5498 22566 5556
rect 22600 5498 22658 5556
rect 22692 5498 22750 5556
rect 22784 5498 22842 5556
rect 22876 5498 22934 5556
rect 22968 5498 23026 5556
rect 23060 5498 23118 5556
rect 23152 5498 23210 5556
rect 23244 5498 23302 5556
rect 23336 5498 23394 5556
rect 23428 5498 23457 5556
rect 24516 5543 24550 5559
rect 24676 5619 24710 5635
rect 24676 5543 24710 5559
rect 11090 5448 11126 5464
rect 11090 5414 11092 5448
rect 11090 5380 11126 5414
rect 11090 5346 11092 5380
rect 11162 5448 11228 5498
rect 11162 5414 11178 5448
rect 11212 5414 11228 5448
rect 11162 5380 11228 5414
rect 11162 5346 11178 5380
rect 11212 5346 11228 5380
rect 11262 5448 11316 5464
rect 11262 5414 11264 5448
rect 11298 5414 11316 5448
rect 11262 5367 11316 5414
rect 11090 5312 11126 5346
rect 11262 5333 11264 5367
rect 11298 5333 11316 5367
rect 11090 5278 11225 5312
rect 11262 5283 11316 5333
rect 11191 5249 11225 5278
rect 11078 5224 11146 5242
rect 11078 5190 11088 5224
rect 11122 5220 11146 5224
rect 11078 5186 11094 5190
rect 11128 5186 11146 5220
rect 11078 5168 11146 5186
rect 11191 5233 11246 5249
rect 11191 5199 11212 5233
rect 11191 5183 11246 5199
rect 11280 5233 11316 5283
rect 11352 5450 11418 5464
rect 11352 5416 11368 5450
rect 11402 5416 11418 5450
rect 11352 5382 11418 5416
rect 11352 5348 11368 5382
rect 11402 5348 11418 5382
rect 11352 5314 11418 5348
rect 11452 5456 11500 5498
rect 11486 5422 11500 5456
rect 11452 5388 11500 5422
rect 11486 5354 11500 5388
rect 11452 5338 11500 5354
rect 11536 5434 11570 5464
rect 11536 5339 11570 5400
rect 11352 5280 11368 5314
rect 11402 5302 11418 5314
rect 11604 5456 11670 5498
rect 11604 5422 11620 5456
rect 11654 5422 11670 5456
rect 11604 5388 11670 5422
rect 11604 5354 11620 5388
rect 11654 5354 11670 5388
rect 11604 5338 11670 5354
rect 11704 5434 11738 5464
rect 11704 5339 11738 5400
rect 11402 5280 11495 5302
rect 11352 5268 11495 5280
rect 11351 5233 11427 5234
rect 11280 5220 11427 5233
rect 11280 5188 11377 5220
rect 11191 5132 11225 5183
rect 11092 5098 11225 5132
rect 11280 5123 11316 5188
rect 11351 5186 11377 5188
rect 11411 5186 11427 5220
rect 11461 5220 11495 5268
rect 11536 5294 11570 5305
rect 11704 5294 11738 5305
rect 11536 5260 11738 5294
rect 11772 5456 11838 5498
rect 11772 5422 11788 5456
rect 11822 5422 11838 5456
rect 11772 5388 11838 5422
rect 11772 5354 11788 5388
rect 11822 5354 11838 5388
rect 11772 5320 11838 5354
rect 11772 5286 11788 5320
rect 11822 5286 11838 5320
rect 11772 5268 11838 5286
rect 11900 5456 11934 5498
rect 11900 5388 11934 5422
rect 11900 5320 11934 5354
rect 11900 5260 11934 5286
rect 11968 5450 12034 5464
rect 11968 5416 11984 5450
rect 12018 5416 12034 5450
rect 11968 5382 12034 5416
rect 11968 5348 11984 5382
rect 12018 5348 12034 5382
rect 11968 5314 12034 5348
rect 12068 5456 12102 5498
rect 12068 5388 12102 5422
rect 12068 5338 12102 5354
rect 12136 5450 12202 5464
rect 12136 5416 12152 5450
rect 12186 5416 12202 5450
rect 12136 5382 12202 5416
rect 12136 5348 12152 5382
rect 12186 5348 12202 5382
rect 11968 5280 11984 5314
rect 12018 5294 12034 5314
rect 12136 5314 12202 5348
rect 12236 5456 12270 5498
rect 12236 5388 12270 5422
rect 12236 5338 12270 5354
rect 12304 5450 12370 5464
rect 12304 5416 12320 5450
rect 12354 5416 12370 5450
rect 12304 5382 12370 5416
rect 12304 5348 12320 5382
rect 12354 5348 12370 5382
rect 12136 5294 12152 5314
rect 12018 5280 12152 5294
rect 12186 5294 12202 5314
rect 12304 5314 12370 5348
rect 12404 5456 12438 5498
rect 12404 5388 12438 5422
rect 12404 5338 12438 5354
rect 12472 5450 12538 5464
rect 12472 5416 12488 5450
rect 12522 5416 12538 5450
rect 12472 5382 12538 5416
rect 12472 5348 12488 5382
rect 12522 5348 12538 5382
rect 12304 5294 12320 5314
rect 12186 5280 12320 5294
rect 12354 5294 12370 5314
rect 12472 5314 12538 5348
rect 12572 5456 12606 5498
rect 12572 5388 12606 5422
rect 12572 5338 12606 5354
rect 12640 5450 12706 5464
rect 12640 5416 12656 5450
rect 12690 5416 12706 5450
rect 12640 5382 12706 5416
rect 12640 5348 12656 5382
rect 12690 5348 12706 5382
rect 12354 5280 12438 5294
rect 11968 5260 12438 5280
rect 12472 5280 12488 5314
rect 12522 5294 12538 5314
rect 12640 5314 12706 5348
rect 12740 5456 12774 5498
rect 12740 5388 12774 5422
rect 12740 5338 12774 5354
rect 12808 5450 12874 5464
rect 12808 5416 12824 5450
rect 12858 5416 12874 5450
rect 12808 5382 12874 5416
rect 12808 5348 12824 5382
rect 12858 5348 12874 5382
rect 12640 5294 12656 5314
rect 12522 5280 12656 5294
rect 12690 5294 12706 5314
rect 12808 5314 12874 5348
rect 12908 5456 12942 5498
rect 12908 5388 12942 5422
rect 12908 5338 12942 5354
rect 12976 5450 13042 5464
rect 12976 5416 12992 5450
rect 13026 5416 13042 5450
rect 12976 5394 13042 5416
rect 12976 5382 13001 5394
rect 12976 5348 12992 5382
rect 13035 5360 13042 5394
rect 13026 5348 13042 5360
rect 12808 5294 12824 5314
rect 12690 5280 12824 5294
rect 12858 5294 12874 5314
rect 12976 5314 13042 5348
rect 13076 5456 13110 5498
rect 13076 5388 13110 5422
rect 13076 5338 13110 5354
rect 13144 5450 13210 5464
rect 13144 5416 13160 5450
rect 13194 5416 13210 5450
rect 13144 5382 13210 5416
rect 13144 5348 13160 5382
rect 13194 5348 13210 5382
rect 12976 5294 12992 5314
rect 12858 5280 12992 5294
rect 13026 5294 13042 5314
rect 13144 5314 13210 5348
rect 13244 5456 13278 5498
rect 13244 5388 13278 5422
rect 13244 5338 13278 5354
rect 13312 5450 13378 5464
rect 13312 5416 13328 5450
rect 13362 5416 13378 5450
rect 13312 5382 13378 5416
rect 13312 5348 13328 5382
rect 13362 5348 13378 5382
rect 13144 5294 13160 5314
rect 13026 5280 13160 5294
rect 13194 5294 13210 5314
rect 13312 5314 13378 5348
rect 13412 5456 13446 5498
rect 13412 5388 13446 5422
rect 13412 5338 13446 5354
rect 13480 5450 13546 5464
rect 13480 5416 13496 5450
rect 13530 5416 13546 5450
rect 13480 5382 13546 5416
rect 13480 5348 13496 5382
rect 13530 5348 13546 5382
rect 13312 5294 13328 5314
rect 13194 5280 13328 5294
rect 13362 5294 13378 5314
rect 13480 5314 13546 5348
rect 13580 5456 13614 5498
rect 13580 5388 13614 5422
rect 13580 5338 13614 5354
rect 13648 5450 13714 5464
rect 13648 5416 13664 5450
rect 13698 5416 13714 5450
rect 13648 5382 13714 5416
rect 13648 5348 13664 5382
rect 13698 5348 13714 5382
rect 13480 5294 13496 5314
rect 13362 5280 13496 5294
rect 13530 5294 13546 5314
rect 13648 5314 13714 5348
rect 13748 5456 13782 5498
rect 13748 5388 13782 5422
rect 13748 5338 13782 5354
rect 13648 5294 13664 5314
rect 13530 5280 13664 5294
rect 13698 5294 13714 5314
rect 13817 5294 13872 5443
rect 13698 5280 13872 5294
rect 12472 5260 13872 5280
rect 11639 5226 11738 5260
rect 12403 5226 12438 5260
rect 11639 5220 12362 5226
rect 11461 5186 11511 5220
rect 11545 5186 11561 5220
rect 11639 5186 11968 5220
rect 12002 5186 12036 5220
rect 12070 5186 12104 5220
rect 12138 5186 12172 5220
rect 12206 5186 12240 5220
rect 12274 5186 12308 5220
rect 12342 5186 12362 5220
rect 12403 5220 13747 5226
rect 12403 5186 12468 5220
rect 12502 5186 12536 5220
rect 12570 5186 12604 5220
rect 12638 5186 12672 5220
rect 12706 5186 12740 5220
rect 12774 5186 12808 5220
rect 12842 5186 12876 5220
rect 12910 5186 12944 5220
rect 12978 5186 13012 5220
rect 13046 5186 13080 5220
rect 13114 5186 13148 5220
rect 13182 5186 13216 5220
rect 13250 5186 13284 5220
rect 13318 5186 13352 5220
rect 13386 5186 13420 5220
rect 13454 5186 13488 5220
rect 13522 5186 13556 5220
rect 13590 5186 13624 5220
rect 13658 5186 13692 5220
rect 13726 5186 13747 5220
rect 11461 5152 11495 5186
rect 11639 5152 11738 5186
rect 12403 5152 12438 5186
rect 13796 5152 13872 5260
rect 11092 5077 11126 5098
rect 11264 5094 11316 5123
rect 11092 5022 11126 5043
rect 11162 5030 11178 5064
rect 11212 5030 11228 5064
rect 11162 4988 11228 5030
rect 11298 5060 11316 5094
rect 11264 5022 11316 5060
rect 11368 5118 11495 5152
rect 11536 5118 11738 5152
rect 11368 5100 11402 5118
rect 11536 5100 11570 5118
rect 11368 5022 11402 5066
rect 11438 5068 11486 5084
rect 11438 5034 11452 5068
rect 11438 4988 11486 5034
rect 11704 5100 11738 5118
rect 11536 5022 11570 5066
rect 11604 5068 11670 5084
rect 11604 5034 11620 5068
rect 11654 5034 11670 5068
rect 11604 4988 11670 5034
rect 11704 5022 11738 5066
rect 11772 5132 11838 5148
rect 11772 5098 11788 5132
rect 11822 5098 11838 5132
rect 11772 5064 11838 5098
rect 11772 5030 11788 5064
rect 11822 5030 11838 5064
rect 11772 4988 11838 5030
rect 11900 5136 11934 5152
rect 11900 5068 11934 5102
rect 11900 4988 11934 5034
rect 11968 5136 12438 5152
rect 11968 5102 11984 5136
rect 12018 5118 12152 5136
rect 12018 5102 12034 5118
rect 11968 5068 12034 5102
rect 12136 5102 12152 5118
rect 12186 5118 12320 5136
rect 12186 5102 12202 5118
rect 11968 5034 11984 5068
rect 12018 5034 12034 5068
rect 11968 5023 12034 5034
rect 12068 5068 12102 5084
rect 12068 4988 12102 5034
rect 12136 5068 12202 5102
rect 12304 5102 12320 5118
rect 12354 5118 12438 5136
rect 12472 5136 13872 5152
rect 12354 5102 12370 5118
rect 12136 5034 12152 5068
rect 12186 5034 12202 5068
rect 12136 5023 12202 5034
rect 12236 5068 12270 5084
rect 12236 4988 12270 5034
rect 12304 5068 12370 5102
rect 12472 5102 12488 5136
rect 12522 5118 12656 5136
rect 12522 5102 12538 5118
rect 12304 5034 12320 5068
rect 12354 5034 12370 5068
rect 12304 5023 12370 5034
rect 12404 5068 12438 5084
rect 12404 4988 12438 5034
rect 12472 5068 12538 5102
rect 12640 5102 12656 5118
rect 12690 5118 12824 5136
rect 12690 5102 12706 5118
rect 12472 5034 12488 5068
rect 12522 5034 12538 5068
rect 12472 5023 12538 5034
rect 12572 5068 12606 5084
rect 12472 5022 12522 5023
rect 12572 4988 12606 5034
rect 12640 5068 12706 5102
rect 12808 5102 12824 5118
rect 12858 5118 12992 5136
rect 12858 5102 12874 5118
rect 12640 5034 12656 5068
rect 12690 5034 12706 5068
rect 12640 5023 12706 5034
rect 12740 5068 12774 5084
rect 12656 5022 12690 5023
rect 12740 4988 12774 5034
rect 12808 5068 12874 5102
rect 12976 5102 12992 5118
rect 13026 5118 13160 5136
rect 13026 5102 13042 5118
rect 12808 5034 12824 5068
rect 12858 5034 12874 5068
rect 12808 5023 12874 5034
rect 12908 5068 12942 5084
rect 12824 5022 12858 5023
rect 12908 4988 12942 5034
rect 12976 5068 13042 5102
rect 13144 5102 13160 5118
rect 13194 5118 13328 5136
rect 13194 5102 13210 5118
rect 12976 5034 12992 5068
rect 13026 5034 13042 5068
rect 12976 5023 13042 5034
rect 13076 5068 13110 5084
rect 13076 4988 13110 5034
rect 13144 5068 13210 5102
rect 13312 5102 13328 5118
rect 13362 5118 13496 5136
rect 13362 5102 13378 5118
rect 13144 5034 13160 5068
rect 13194 5034 13210 5068
rect 13144 5023 13210 5034
rect 13244 5068 13278 5084
rect 13244 4988 13278 5034
rect 13312 5068 13378 5102
rect 13480 5102 13496 5118
rect 13530 5118 13664 5136
rect 13530 5102 13546 5118
rect 13312 5034 13328 5068
rect 13362 5034 13378 5068
rect 13312 5023 13378 5034
rect 13412 5068 13446 5084
rect 13412 4988 13446 5034
rect 13480 5068 13546 5102
rect 13648 5102 13664 5118
rect 13698 5118 13872 5136
rect 13698 5102 13714 5118
rect 13480 5034 13496 5068
rect 13530 5034 13546 5068
rect 13480 5023 13546 5034
rect 13580 5068 13614 5084
rect 13580 4988 13614 5034
rect 13648 5068 13714 5102
rect 13817 5093 13872 5118
rect 13648 5034 13664 5068
rect 13698 5034 13714 5068
rect 13648 5023 13714 5034
rect 13748 5068 13782 5084
rect 13817 5059 13829 5093
rect 13863 5059 13872 5093
rect 13817 5044 13872 5059
rect 13906 5430 13958 5464
rect 13906 5396 13915 5430
rect 13949 5420 13958 5430
rect 13906 5386 13924 5396
rect 13906 5352 13958 5386
rect 13906 5318 13924 5352
rect 13992 5444 14051 5498
rect 13992 5410 14008 5444
rect 14042 5410 14051 5444
rect 13992 5376 14051 5410
rect 13992 5342 14008 5376
rect 14042 5342 14051 5376
rect 13992 5324 14051 5342
rect 14087 5438 14150 5454
rect 14087 5404 14103 5438
rect 14137 5404 14150 5438
rect 14087 5370 14150 5404
rect 14087 5336 14103 5370
rect 14137 5336 14150 5370
rect 13906 5260 13958 5318
rect 13906 5136 13949 5260
rect 14087 5236 14150 5336
rect 13983 5220 14150 5236
rect 14017 5186 14150 5220
rect 13983 5170 14150 5186
rect 13906 5100 13958 5136
rect 13906 5066 13924 5100
rect 14087 5090 14150 5170
rect 13748 4988 13782 5034
rect 13906 5022 13958 5066
rect 13992 5064 14051 5080
rect 13992 5030 14008 5064
rect 14042 5030 14051 5064
rect 13992 4988 14051 5030
rect 14087 5056 14103 5090
rect 14137 5056 14150 5090
rect 14087 5022 14150 5056
rect 14184 5419 14241 5464
rect 14275 5456 14552 5498
rect 14275 5422 14291 5456
rect 14325 5422 14502 5456
rect 14536 5422 14552 5456
rect 14740 5456 14816 5498
rect 14658 5430 14692 5446
rect 14184 5385 14207 5419
rect 14740 5422 14766 5456
rect 14800 5422 14816 5456
rect 15239 5456 15305 5498
rect 14658 5388 14692 5396
rect 14864 5421 14980 5455
rect 15014 5421 15030 5455
rect 15239 5422 15255 5456
rect 15289 5422 15305 5456
rect 15523 5446 15599 5498
rect 14184 5351 14241 5385
rect 14184 5317 14207 5351
rect 14184 5297 14241 5317
rect 14275 5354 14830 5388
rect 14184 5114 14225 5297
rect 14275 5236 14309 5354
rect 14372 5286 14388 5320
rect 14422 5294 14524 5320
rect 14422 5286 14469 5294
rect 14503 5260 14524 5294
rect 14469 5252 14524 5260
rect 14259 5220 14309 5236
rect 14293 5186 14309 5220
rect 14343 5228 14418 5236
rect 14343 5224 14361 5228
rect 14343 5190 14359 5224
rect 14395 5194 14418 5228
rect 14393 5190 14418 5194
rect 14469 5218 14490 5252
rect 14259 5170 14309 5186
rect 14469 5156 14524 5218
rect 14184 5098 14241 5114
rect 14184 5064 14207 5098
rect 14184 5022 14241 5064
rect 14275 5064 14341 5132
rect 14275 5030 14291 5064
rect 14325 5030 14341 5064
rect 14275 4988 14341 5030
rect 14386 5122 14524 5156
rect 14558 5127 14594 5354
rect 14780 5336 14830 5354
rect 14780 5302 14796 5336
rect 14780 5286 14830 5302
rect 14864 5252 14898 5421
rect 15239 5388 15305 5422
rect 15021 5362 15068 5368
rect 14628 5236 14898 5252
rect 14662 5218 14898 5236
rect 14662 5202 14672 5218
rect 14628 5186 14672 5202
rect 14714 5150 14736 5184
rect 14770 5158 14789 5184
rect 14558 5124 14624 5127
rect 14386 5074 14433 5122
rect 14558 5090 14574 5124
rect 14608 5090 14624 5124
rect 14714 5124 14745 5150
rect 14779 5124 14789 5158
rect 14714 5118 14789 5124
rect 14420 5040 14433 5074
rect 14386 5024 14433 5040
rect 14490 5072 14524 5088
rect 14658 5056 14674 5080
rect 14524 5046 14674 5056
rect 14708 5046 14724 5080
rect 14524 5038 14724 5046
rect 14490 5022 14724 5038
rect 14776 5060 14828 5076
rect 14810 5026 14828 5060
rect 14776 4988 14828 5026
rect 14864 5064 14898 5218
rect 14932 5336 14973 5352
rect 14966 5302 14973 5336
rect 14932 5232 14973 5302
rect 15055 5336 15068 5362
rect 15239 5354 15255 5388
rect 15289 5354 15305 5388
rect 15429 5430 15463 5446
rect 15523 5412 15549 5446
rect 15583 5412 15599 5446
rect 15647 5421 15763 5455
rect 15797 5421 15813 5455
rect 15856 5448 15890 5464
rect 15429 5378 15463 5396
rect 15343 5362 15613 5378
rect 15021 5302 15034 5328
rect 15343 5328 15429 5362
rect 15463 5336 15613 5362
rect 15463 5328 15579 5336
rect 15021 5286 15068 5302
rect 15108 5294 15309 5302
rect 15108 5260 15113 5294
rect 15147 5260 15309 5294
rect 15108 5254 15309 5260
rect 15243 5252 15309 5254
rect 14932 5226 15056 5232
rect 14932 5196 15021 5226
rect 14999 5192 15021 5196
rect 15055 5192 15056 5226
rect 15243 5218 15259 5252
rect 15293 5218 15309 5252
rect 14999 5162 15056 5192
rect 15033 5128 15056 5162
rect 15115 5184 15131 5218
rect 15165 5184 15181 5218
rect 15343 5184 15377 5328
rect 15563 5302 15579 5328
rect 15563 5286 15613 5302
rect 15411 5252 15461 5268
rect 15647 5252 15681 5421
rect 15856 5364 15890 5414
rect 15924 5432 15994 5498
rect 15924 5398 15940 5432
rect 15974 5398 15994 5432
rect 16033 5448 16078 5464
rect 16033 5414 16044 5448
rect 16033 5380 16078 5414
rect 16112 5432 16178 5498
rect 16112 5398 16128 5432
rect 16162 5398 16178 5432
rect 16212 5448 16264 5464
rect 16246 5414 16264 5448
rect 15715 5336 15757 5362
rect 15749 5328 15757 5336
rect 15791 5328 15815 5362
rect 15856 5330 15999 5364
rect 15749 5302 15815 5328
rect 15715 5286 15815 5302
rect 15445 5218 15681 5252
rect 15411 5202 15455 5218
rect 15601 5210 15681 5218
rect 15115 5150 15377 5184
rect 15497 5164 15513 5184
rect 14999 5112 15056 5128
rect 15333 5124 15377 5150
rect 15481 5158 15513 5164
rect 15547 5150 15563 5184
rect 15515 5124 15563 5150
rect 15265 5098 15299 5114
rect 15333 5090 15349 5124
rect 15383 5090 15399 5124
rect 15481 5118 15563 5124
rect 14864 5030 14967 5064
rect 15001 5030 15017 5064
rect 14864 5024 15017 5030
rect 15145 5030 15161 5064
rect 15195 5030 15211 5064
rect 15145 4988 15211 5030
rect 15265 5056 15299 5064
rect 15433 5056 15449 5080
rect 15265 5046 15449 5056
rect 15483 5046 15499 5080
rect 15265 5022 15499 5046
rect 15533 5060 15567 5076
rect 15533 4988 15567 5026
rect 15601 5064 15635 5210
rect 15669 5158 15685 5174
rect 15719 5140 15735 5174
rect 15703 5124 15735 5140
rect 15669 5100 15735 5124
rect 15771 5162 15815 5286
rect 15849 5292 15931 5296
rect 15849 5258 15893 5292
rect 15927 5258 15931 5292
rect 15849 5222 15931 5258
rect 15849 5188 15897 5222
rect 15849 5172 15931 5188
rect 15771 5128 15781 5162
rect 15965 5136 15999 5330
rect 15771 5112 15815 5128
rect 15856 5098 15999 5136
rect 16033 5346 16044 5380
rect 16212 5380 16264 5414
rect 16033 5158 16078 5346
rect 16067 5124 16078 5158
rect 15856 5082 15890 5098
rect 15601 5030 15750 5064
rect 15784 5030 15800 5064
rect 16033 5090 16078 5124
rect 16113 5362 16212 5364
rect 16113 5328 16125 5362
rect 16159 5346 16212 5362
rect 16246 5346 16264 5380
rect 16159 5330 16264 5346
rect 16298 5420 16350 5464
rect 16298 5386 16316 5420
rect 16298 5352 16350 5386
rect 16113 5235 16159 5328
rect 16298 5318 16316 5352
rect 16384 5444 16443 5498
rect 16384 5410 16400 5444
rect 16434 5410 16443 5444
rect 16384 5376 16443 5410
rect 16384 5342 16400 5376
rect 16434 5342 16443 5376
rect 16384 5324 16443 5342
rect 16479 5438 16542 5454
rect 16479 5404 16495 5438
rect 16529 5404 16542 5438
rect 16479 5370 16542 5404
rect 16479 5336 16495 5370
rect 16529 5336 16542 5370
rect 16298 5296 16350 5318
rect 16147 5201 16159 5235
rect 16113 5132 16159 5201
rect 16193 5235 16264 5296
rect 16193 5207 16215 5235
rect 16193 5173 16213 5207
rect 16249 5201 16264 5235
rect 16247 5173 16264 5201
rect 16193 5166 16264 5173
rect 16298 5262 16304 5296
rect 16338 5262 16350 5296
rect 16298 5260 16350 5262
rect 16298 5136 16341 5260
rect 16479 5236 16542 5336
rect 16375 5220 16542 5236
rect 16409 5186 16542 5220
rect 16375 5170 16542 5186
rect 16113 5098 16264 5132
rect 15856 5032 15890 5048
rect 15601 5024 15800 5030
rect 15924 5030 15940 5064
rect 15974 5030 15994 5064
rect 16033 5056 16044 5090
rect 16212 5090 16264 5098
rect 16033 5040 16078 5056
rect 15924 4988 15994 5030
rect 16112 5030 16128 5064
rect 16162 5030 16178 5064
rect 16246 5056 16264 5090
rect 16212 5040 16264 5056
rect 16298 5128 16350 5136
rect 16298 5094 16308 5128
rect 16342 5100 16350 5128
rect 16298 5066 16316 5094
rect 16479 5090 16542 5170
rect 16112 4988 16178 5030
rect 16298 5022 16350 5066
rect 16384 5064 16443 5080
rect 16384 5030 16400 5064
rect 16434 5030 16443 5064
rect 16384 4988 16443 5030
rect 16479 5056 16495 5090
rect 16529 5056 16542 5090
rect 16479 5022 16542 5056
rect 16576 5419 16633 5464
rect 16667 5456 16944 5498
rect 16667 5422 16683 5456
rect 16717 5422 16894 5456
rect 16928 5422 16944 5456
rect 17132 5456 17208 5498
rect 17050 5430 17084 5446
rect 16576 5385 16599 5419
rect 17132 5422 17158 5456
rect 17192 5422 17208 5456
rect 17631 5456 17697 5498
rect 17050 5388 17084 5396
rect 17256 5421 17372 5455
rect 17406 5421 17422 5455
rect 17631 5422 17647 5456
rect 17681 5422 17697 5456
rect 17915 5446 17991 5498
rect 16576 5351 16633 5385
rect 16576 5317 16599 5351
rect 16576 5297 16633 5317
rect 16667 5354 17222 5388
rect 16576 5114 16617 5297
rect 16667 5236 16701 5354
rect 16764 5286 16780 5320
rect 16814 5294 16916 5320
rect 16814 5286 16861 5294
rect 16895 5260 16916 5294
rect 16861 5252 16916 5260
rect 16651 5220 16701 5236
rect 16685 5186 16701 5220
rect 16735 5230 16810 5236
rect 16735 5224 16755 5230
rect 16735 5190 16751 5224
rect 16789 5196 16810 5230
rect 16785 5190 16810 5196
rect 16861 5218 16882 5252
rect 16651 5170 16701 5186
rect 16861 5156 16916 5218
rect 16576 5098 16633 5114
rect 16576 5089 16599 5098
rect 16576 5055 16594 5089
rect 16628 5055 16633 5064
rect 16576 5022 16633 5055
rect 16667 5064 16733 5132
rect 16667 5030 16683 5064
rect 16717 5030 16733 5064
rect 16667 4988 16733 5030
rect 16778 5122 16916 5156
rect 16950 5127 16986 5354
rect 17172 5336 17222 5354
rect 17172 5302 17188 5336
rect 17172 5286 17222 5302
rect 17256 5252 17290 5421
rect 17631 5388 17697 5422
rect 17413 5362 17460 5368
rect 17020 5236 17290 5252
rect 17054 5218 17290 5236
rect 17054 5202 17064 5218
rect 17020 5186 17064 5202
rect 17106 5150 17128 5184
rect 17162 5158 17181 5184
rect 16950 5124 17016 5127
rect 16778 5074 16825 5122
rect 16950 5090 16966 5124
rect 17000 5090 17016 5124
rect 17106 5124 17137 5150
rect 17171 5124 17181 5158
rect 17106 5118 17181 5124
rect 16812 5040 16825 5074
rect 16778 5024 16825 5040
rect 16882 5072 16916 5088
rect 17050 5056 17066 5080
rect 16916 5046 17066 5056
rect 17100 5046 17116 5080
rect 16916 5038 17116 5046
rect 16882 5022 17116 5038
rect 17168 5060 17220 5076
rect 17202 5026 17220 5060
rect 17168 4988 17220 5026
rect 17256 5064 17290 5218
rect 17324 5336 17365 5352
rect 17358 5302 17365 5336
rect 17324 5232 17365 5302
rect 17447 5336 17460 5362
rect 17631 5354 17647 5388
rect 17681 5354 17697 5388
rect 17821 5430 17855 5446
rect 17915 5412 17941 5446
rect 17975 5412 17991 5446
rect 18039 5421 18155 5455
rect 18189 5421 18205 5455
rect 18248 5448 18282 5464
rect 17821 5378 17855 5396
rect 17735 5362 18005 5378
rect 17413 5302 17426 5328
rect 17735 5328 17821 5362
rect 17855 5336 18005 5362
rect 17855 5328 17971 5336
rect 17413 5286 17460 5302
rect 17500 5294 17701 5302
rect 17500 5260 17505 5294
rect 17539 5260 17701 5294
rect 17500 5254 17701 5260
rect 17635 5252 17701 5254
rect 17324 5226 17448 5232
rect 17324 5196 17413 5226
rect 17391 5192 17413 5196
rect 17447 5192 17448 5226
rect 17635 5218 17651 5252
rect 17685 5218 17701 5252
rect 17391 5162 17448 5192
rect 17425 5128 17448 5162
rect 17507 5184 17523 5218
rect 17557 5184 17573 5218
rect 17735 5184 17769 5328
rect 17955 5302 17971 5328
rect 17955 5286 18005 5302
rect 17803 5252 17853 5268
rect 18039 5252 18073 5421
rect 18248 5364 18282 5414
rect 18316 5432 18386 5498
rect 18316 5398 18332 5432
rect 18366 5398 18386 5432
rect 18425 5448 18470 5464
rect 18425 5414 18436 5448
rect 18425 5380 18470 5414
rect 18504 5432 18570 5498
rect 18504 5398 18520 5432
rect 18554 5398 18570 5432
rect 18604 5448 18656 5464
rect 18638 5414 18656 5448
rect 18107 5336 18149 5362
rect 18141 5328 18149 5336
rect 18183 5328 18207 5362
rect 18248 5330 18391 5364
rect 18141 5302 18207 5328
rect 18107 5286 18207 5302
rect 17837 5218 18073 5252
rect 17803 5202 17847 5218
rect 17993 5210 18073 5218
rect 17507 5150 17769 5184
rect 17889 5164 17905 5184
rect 17391 5112 17448 5128
rect 17725 5124 17769 5150
rect 17873 5158 17905 5164
rect 17939 5150 17955 5184
rect 17907 5124 17955 5150
rect 17657 5098 17691 5114
rect 17725 5090 17741 5124
rect 17775 5090 17791 5124
rect 17873 5118 17955 5124
rect 17256 5030 17359 5064
rect 17393 5030 17409 5064
rect 17256 5024 17409 5030
rect 17537 5030 17553 5064
rect 17587 5030 17603 5064
rect 17537 4988 17603 5030
rect 17657 5056 17691 5064
rect 17825 5056 17841 5080
rect 17657 5046 17841 5056
rect 17875 5046 17891 5080
rect 17657 5022 17891 5046
rect 17925 5060 17959 5076
rect 17925 4988 17959 5026
rect 17993 5064 18027 5210
rect 18061 5158 18077 5174
rect 18111 5140 18127 5174
rect 18095 5124 18127 5140
rect 18061 5100 18127 5124
rect 18163 5162 18207 5286
rect 18241 5292 18323 5296
rect 18241 5258 18285 5292
rect 18319 5258 18323 5292
rect 18241 5222 18323 5258
rect 18241 5188 18289 5222
rect 18241 5172 18323 5188
rect 18163 5128 18173 5162
rect 18357 5136 18391 5330
rect 18163 5112 18207 5128
rect 18248 5098 18391 5136
rect 18425 5346 18436 5380
rect 18604 5380 18656 5414
rect 18425 5158 18470 5346
rect 18459 5124 18470 5158
rect 18248 5082 18282 5098
rect 17993 5030 18142 5064
rect 18176 5030 18192 5064
rect 18425 5090 18470 5124
rect 18505 5362 18604 5364
rect 18505 5328 18517 5362
rect 18551 5346 18604 5362
rect 18638 5346 18656 5380
rect 18551 5330 18656 5346
rect 18690 5420 18742 5464
rect 18690 5386 18708 5420
rect 18690 5352 18742 5386
rect 18505 5235 18551 5328
rect 18690 5318 18708 5352
rect 18776 5444 18835 5498
rect 18776 5410 18792 5444
rect 18826 5410 18835 5444
rect 18776 5376 18835 5410
rect 18776 5342 18792 5376
rect 18826 5342 18835 5376
rect 18776 5324 18835 5342
rect 18871 5438 18934 5454
rect 18871 5404 18887 5438
rect 18921 5404 18934 5438
rect 18871 5370 18934 5404
rect 18871 5336 18887 5370
rect 18921 5336 18934 5370
rect 18690 5296 18742 5318
rect 18539 5201 18551 5235
rect 18505 5132 18551 5201
rect 18585 5235 18656 5296
rect 18585 5201 18607 5235
rect 18641 5208 18656 5235
rect 18585 5174 18610 5201
rect 18644 5174 18656 5208
rect 18585 5166 18656 5174
rect 18690 5262 18696 5296
rect 18730 5262 18742 5296
rect 18690 5260 18742 5262
rect 18690 5136 18733 5260
rect 18871 5236 18934 5336
rect 18767 5220 18934 5236
rect 18801 5186 18934 5220
rect 18767 5170 18934 5186
rect 18505 5098 18656 5132
rect 18248 5032 18282 5048
rect 17993 5024 18192 5030
rect 18316 5030 18332 5064
rect 18366 5030 18386 5064
rect 18425 5056 18436 5090
rect 18604 5090 18656 5098
rect 18425 5040 18470 5056
rect 18316 4988 18386 5030
rect 18504 5030 18520 5064
rect 18554 5030 18570 5064
rect 18638 5056 18656 5090
rect 18604 5040 18656 5056
rect 18690 5115 18742 5136
rect 18690 5066 18708 5115
rect 18871 5090 18934 5170
rect 18504 4988 18570 5030
rect 18690 5022 18742 5066
rect 18776 5064 18835 5080
rect 18776 5030 18792 5064
rect 18826 5030 18835 5064
rect 18776 4988 18835 5030
rect 18871 5056 18887 5090
rect 18921 5056 18934 5090
rect 18871 5022 18934 5056
rect 18968 5419 19025 5464
rect 19059 5456 19336 5498
rect 19059 5422 19075 5456
rect 19109 5422 19286 5456
rect 19320 5422 19336 5456
rect 19524 5456 19600 5498
rect 19442 5430 19476 5446
rect 18968 5385 18991 5419
rect 19524 5422 19550 5456
rect 19584 5422 19600 5456
rect 20023 5456 20089 5498
rect 19442 5388 19476 5396
rect 19648 5421 19764 5455
rect 19798 5421 19814 5455
rect 20023 5422 20039 5456
rect 20073 5422 20089 5456
rect 20307 5446 20383 5498
rect 18968 5351 19025 5385
rect 18968 5317 18991 5351
rect 18968 5297 19025 5317
rect 19059 5354 19614 5388
rect 18968 5114 19009 5297
rect 19059 5236 19093 5354
rect 19156 5286 19172 5320
rect 19206 5294 19308 5320
rect 19206 5286 19253 5294
rect 19287 5260 19308 5294
rect 19253 5252 19308 5260
rect 19043 5220 19093 5236
rect 19077 5186 19093 5220
rect 19127 5231 19202 5236
rect 19127 5224 19145 5231
rect 19127 5190 19143 5224
rect 19179 5197 19202 5231
rect 19177 5190 19202 5197
rect 19253 5218 19274 5252
rect 19043 5170 19093 5186
rect 19253 5156 19308 5218
rect 18968 5098 19025 5114
rect 18968 5088 18991 5098
rect 18968 5054 18982 5088
rect 19016 5054 19025 5064
rect 18968 5022 19025 5054
rect 19059 5064 19125 5132
rect 19059 5030 19075 5064
rect 19109 5030 19125 5064
rect 19059 4988 19125 5030
rect 19170 5122 19308 5156
rect 19342 5127 19378 5354
rect 19564 5336 19614 5354
rect 19564 5302 19580 5336
rect 19564 5286 19614 5302
rect 19648 5252 19682 5421
rect 20023 5388 20089 5422
rect 19805 5362 19852 5368
rect 19412 5236 19682 5252
rect 19446 5218 19682 5236
rect 19446 5202 19456 5218
rect 19412 5186 19456 5202
rect 19498 5150 19520 5184
rect 19554 5158 19573 5184
rect 19342 5124 19408 5127
rect 19170 5074 19217 5122
rect 19342 5090 19358 5124
rect 19392 5090 19408 5124
rect 19498 5124 19529 5150
rect 19563 5124 19573 5158
rect 19498 5118 19573 5124
rect 19204 5040 19217 5074
rect 19170 5024 19217 5040
rect 19274 5072 19308 5088
rect 19442 5056 19458 5080
rect 19308 5046 19458 5056
rect 19492 5046 19508 5080
rect 19308 5038 19508 5046
rect 19274 5022 19508 5038
rect 19560 5060 19612 5076
rect 19594 5026 19612 5060
rect 19560 4988 19612 5026
rect 19648 5064 19682 5218
rect 19716 5336 19757 5352
rect 19750 5302 19757 5336
rect 19716 5232 19757 5302
rect 19839 5336 19852 5362
rect 20023 5354 20039 5388
rect 20073 5354 20089 5388
rect 20213 5430 20247 5446
rect 20307 5412 20333 5446
rect 20367 5412 20383 5446
rect 20431 5421 20547 5455
rect 20581 5421 20597 5455
rect 20640 5448 20674 5464
rect 20213 5378 20247 5396
rect 20127 5362 20397 5378
rect 19805 5302 19818 5328
rect 20127 5328 20213 5362
rect 20247 5336 20397 5362
rect 20247 5328 20363 5336
rect 19805 5286 19852 5302
rect 19892 5294 20093 5302
rect 19892 5260 19897 5294
rect 19931 5260 20093 5294
rect 19892 5254 20093 5260
rect 20027 5252 20093 5254
rect 19716 5226 19840 5232
rect 19716 5196 19805 5226
rect 19783 5192 19805 5196
rect 19839 5192 19840 5226
rect 20027 5218 20043 5252
rect 20077 5218 20093 5252
rect 19783 5162 19840 5192
rect 19817 5128 19840 5162
rect 19899 5184 19915 5218
rect 19949 5184 19965 5218
rect 20127 5184 20161 5328
rect 20347 5302 20363 5328
rect 20347 5286 20397 5302
rect 20195 5252 20245 5268
rect 20431 5252 20465 5421
rect 20640 5364 20674 5414
rect 20708 5432 20778 5498
rect 20708 5398 20724 5432
rect 20758 5398 20778 5432
rect 20817 5448 20862 5464
rect 20817 5414 20828 5448
rect 20817 5380 20862 5414
rect 20896 5432 20962 5498
rect 20896 5398 20912 5432
rect 20946 5398 20962 5432
rect 20996 5448 21048 5464
rect 21030 5414 21048 5448
rect 20499 5336 20541 5362
rect 20533 5328 20541 5336
rect 20575 5328 20599 5362
rect 20640 5330 20783 5364
rect 20533 5302 20599 5328
rect 20499 5286 20599 5302
rect 20229 5218 20465 5252
rect 20195 5202 20239 5218
rect 20385 5210 20465 5218
rect 19899 5150 20161 5184
rect 20281 5164 20297 5184
rect 19783 5112 19840 5128
rect 20117 5124 20161 5150
rect 20265 5158 20297 5164
rect 20331 5150 20347 5184
rect 20299 5124 20347 5150
rect 20049 5098 20083 5114
rect 20117 5090 20133 5124
rect 20167 5090 20183 5124
rect 20265 5118 20347 5124
rect 19648 5030 19751 5064
rect 19785 5030 19801 5064
rect 19648 5024 19801 5030
rect 19929 5030 19945 5064
rect 19979 5030 19995 5064
rect 19929 4988 19995 5030
rect 20049 5056 20083 5064
rect 20217 5056 20233 5080
rect 20049 5046 20233 5056
rect 20267 5046 20283 5080
rect 20049 5022 20283 5046
rect 20317 5060 20351 5076
rect 20317 4988 20351 5026
rect 20385 5064 20419 5210
rect 20453 5158 20469 5174
rect 20503 5140 20519 5174
rect 20487 5124 20519 5140
rect 20453 5100 20519 5124
rect 20555 5162 20599 5286
rect 20633 5293 20715 5296
rect 20633 5259 20677 5293
rect 20711 5259 20715 5293
rect 20633 5222 20715 5259
rect 20633 5188 20681 5222
rect 20633 5172 20715 5188
rect 20555 5128 20565 5162
rect 20749 5136 20783 5330
rect 20555 5112 20599 5128
rect 20640 5098 20783 5136
rect 20817 5346 20828 5380
rect 20996 5380 21048 5414
rect 20817 5158 20862 5346
rect 20851 5124 20862 5158
rect 20640 5082 20674 5098
rect 20385 5030 20534 5064
rect 20568 5030 20584 5064
rect 20817 5090 20862 5124
rect 20897 5362 20996 5364
rect 20897 5328 20909 5362
rect 20943 5346 20996 5362
rect 21030 5346 21048 5380
rect 20943 5330 21048 5346
rect 21082 5420 21134 5464
rect 21082 5386 21100 5420
rect 21082 5352 21134 5386
rect 20897 5235 20943 5328
rect 21082 5318 21100 5352
rect 21168 5444 21227 5498
rect 21168 5410 21184 5444
rect 21218 5410 21227 5444
rect 21168 5376 21227 5410
rect 21168 5342 21184 5376
rect 21218 5342 21227 5376
rect 21168 5324 21227 5342
rect 21263 5438 21326 5454
rect 21263 5404 21279 5438
rect 21313 5404 21326 5438
rect 21263 5370 21326 5404
rect 21263 5336 21279 5370
rect 21313 5336 21326 5370
rect 21082 5297 21134 5318
rect 20931 5201 20943 5235
rect 20897 5132 20943 5201
rect 20977 5235 21048 5296
rect 20977 5201 20999 5235
rect 21033 5208 21048 5235
rect 20977 5174 21001 5201
rect 21035 5174 21048 5208
rect 20977 5166 21048 5174
rect 21082 5263 21088 5297
rect 21122 5263 21134 5297
rect 21082 5260 21134 5263
rect 21082 5136 21125 5260
rect 21263 5236 21326 5336
rect 21159 5220 21326 5236
rect 21193 5186 21326 5220
rect 21159 5170 21326 5186
rect 20897 5098 21048 5132
rect 20640 5032 20674 5048
rect 20385 5024 20584 5030
rect 20708 5030 20724 5064
rect 20758 5030 20778 5064
rect 20817 5056 20828 5090
rect 20996 5090 21048 5098
rect 20817 5040 20862 5056
rect 20708 4988 20778 5030
rect 20896 5030 20912 5064
rect 20946 5030 20962 5064
rect 21030 5056 21048 5090
rect 20996 5040 21048 5056
rect 21082 5123 21134 5136
rect 21082 5089 21096 5123
rect 21130 5100 21134 5123
rect 21082 5066 21100 5089
rect 21263 5090 21326 5170
rect 20896 4988 20962 5030
rect 21082 5022 21134 5066
rect 21168 5064 21227 5080
rect 21168 5030 21184 5064
rect 21218 5030 21227 5064
rect 21168 4988 21227 5030
rect 21263 5056 21279 5090
rect 21313 5056 21326 5090
rect 21263 5022 21326 5056
rect 21360 5419 21417 5464
rect 21451 5456 21728 5498
rect 21451 5422 21467 5456
rect 21501 5422 21678 5456
rect 21712 5422 21728 5456
rect 21916 5456 21992 5498
rect 21834 5430 21868 5446
rect 21360 5385 21383 5419
rect 21916 5422 21942 5456
rect 21976 5422 21992 5456
rect 22415 5456 22481 5498
rect 21834 5388 21868 5396
rect 22040 5421 22156 5455
rect 22190 5421 22206 5455
rect 22415 5422 22431 5456
rect 22465 5422 22481 5456
rect 22699 5446 22775 5498
rect 21360 5351 21417 5385
rect 21360 5317 21383 5351
rect 21360 5297 21417 5317
rect 21451 5354 22006 5388
rect 21360 5114 21401 5297
rect 21451 5236 21485 5354
rect 21548 5286 21564 5320
rect 21598 5294 21700 5320
rect 21598 5286 21645 5294
rect 21679 5260 21700 5294
rect 21645 5252 21700 5260
rect 21435 5220 21485 5236
rect 21469 5186 21485 5220
rect 21519 5228 21594 5236
rect 21519 5224 21539 5228
rect 21519 5190 21535 5224
rect 21573 5194 21594 5228
rect 21569 5190 21594 5194
rect 21645 5218 21666 5252
rect 21435 5170 21485 5186
rect 21645 5156 21700 5218
rect 21360 5098 21417 5114
rect 21360 5094 21383 5098
rect 21360 5060 21376 5094
rect 21410 5060 21417 5064
rect 21360 5022 21417 5060
rect 21451 5064 21517 5132
rect 21451 5030 21467 5064
rect 21501 5030 21517 5064
rect 21451 4988 21517 5030
rect 21562 5122 21700 5156
rect 21734 5127 21770 5354
rect 21956 5336 22006 5354
rect 21956 5302 21972 5336
rect 21956 5286 22006 5302
rect 22040 5252 22074 5421
rect 22415 5388 22481 5422
rect 22197 5362 22244 5368
rect 21804 5236 22074 5252
rect 21838 5218 22074 5236
rect 21838 5202 21848 5218
rect 21804 5186 21848 5202
rect 21890 5150 21912 5184
rect 21946 5158 21965 5184
rect 21734 5124 21800 5127
rect 21562 5074 21609 5122
rect 21734 5090 21750 5124
rect 21784 5090 21800 5124
rect 21890 5124 21921 5150
rect 21955 5124 21965 5158
rect 21890 5118 21965 5124
rect 21596 5040 21609 5074
rect 21562 5024 21609 5040
rect 21666 5072 21700 5088
rect 21834 5056 21850 5080
rect 21700 5046 21850 5056
rect 21884 5046 21900 5080
rect 21700 5038 21900 5046
rect 21666 5022 21900 5038
rect 21952 5060 22004 5076
rect 21986 5026 22004 5060
rect 21952 4988 22004 5026
rect 22040 5064 22074 5218
rect 22108 5336 22149 5352
rect 22142 5302 22149 5336
rect 22108 5232 22149 5302
rect 22231 5336 22244 5362
rect 22415 5354 22431 5388
rect 22465 5354 22481 5388
rect 22605 5430 22639 5446
rect 22699 5412 22725 5446
rect 22759 5412 22775 5446
rect 22823 5421 22939 5455
rect 22973 5421 22989 5455
rect 23032 5448 23066 5464
rect 22605 5378 22639 5396
rect 22519 5362 22789 5378
rect 22197 5302 22210 5328
rect 22519 5328 22605 5362
rect 22639 5336 22789 5362
rect 22639 5328 22755 5336
rect 22197 5286 22244 5302
rect 22284 5294 22485 5302
rect 22284 5260 22289 5294
rect 22323 5260 22485 5294
rect 22284 5254 22485 5260
rect 22419 5252 22485 5254
rect 22108 5226 22232 5232
rect 22108 5196 22197 5226
rect 22175 5192 22197 5196
rect 22231 5192 22232 5226
rect 22419 5218 22435 5252
rect 22469 5218 22485 5252
rect 22175 5162 22232 5192
rect 22209 5128 22232 5162
rect 22291 5184 22307 5218
rect 22341 5184 22357 5218
rect 22519 5184 22553 5328
rect 22739 5302 22755 5328
rect 22739 5286 22789 5302
rect 22587 5252 22637 5268
rect 22823 5252 22857 5421
rect 23032 5364 23066 5414
rect 23100 5432 23170 5498
rect 23100 5398 23116 5432
rect 23150 5398 23170 5432
rect 23209 5448 23254 5464
rect 23209 5414 23220 5448
rect 23209 5380 23254 5414
rect 23288 5432 23354 5498
rect 24516 5481 24550 5497
rect 23288 5398 23304 5432
rect 23338 5398 23354 5432
rect 23388 5448 23440 5464
rect 23422 5414 23440 5448
rect 22891 5336 22933 5362
rect 22925 5328 22933 5336
rect 22967 5328 22991 5362
rect 23032 5330 23175 5364
rect 22925 5302 22991 5328
rect 22891 5286 22991 5302
rect 22621 5218 22857 5252
rect 22587 5202 22631 5218
rect 22777 5210 22857 5218
rect 22291 5150 22553 5184
rect 22673 5164 22689 5184
rect 22175 5112 22232 5128
rect 22509 5124 22553 5150
rect 22657 5158 22689 5164
rect 22723 5150 22739 5184
rect 22691 5124 22739 5150
rect 22441 5098 22475 5114
rect 22509 5090 22525 5124
rect 22559 5090 22575 5124
rect 22657 5118 22739 5124
rect 22040 5030 22143 5064
rect 22177 5030 22193 5064
rect 22040 5024 22193 5030
rect 22321 5030 22337 5064
rect 22371 5030 22387 5064
rect 22321 4988 22387 5030
rect 22441 5056 22475 5064
rect 22609 5056 22625 5080
rect 22441 5046 22625 5056
rect 22659 5046 22675 5080
rect 22441 5022 22675 5046
rect 22709 5060 22743 5076
rect 22709 4988 22743 5026
rect 22777 5064 22811 5210
rect 22845 5158 22861 5174
rect 22895 5140 22911 5174
rect 22879 5124 22911 5140
rect 22845 5100 22911 5124
rect 22947 5162 22991 5286
rect 23025 5289 23107 5296
rect 23025 5255 23038 5289
rect 23072 5255 23107 5289
rect 23025 5222 23107 5255
rect 23025 5188 23073 5222
rect 23025 5172 23107 5188
rect 22947 5128 22957 5162
rect 23141 5136 23175 5330
rect 22947 5112 22991 5128
rect 23032 5098 23175 5136
rect 23209 5346 23220 5380
rect 23388 5380 23440 5414
rect 24516 5405 24550 5421
rect 24676 5481 24710 5497
rect 24676 5405 24710 5421
rect 23209 5158 23254 5346
rect 23243 5124 23254 5158
rect 23032 5082 23066 5098
rect 22777 5030 22926 5064
rect 22960 5030 22976 5064
rect 23209 5090 23254 5124
rect 23289 5362 23388 5364
rect 23289 5328 23301 5362
rect 23335 5346 23388 5362
rect 23422 5346 23440 5380
rect 23335 5330 23440 5346
rect 24516 5343 24550 5359
rect 23289 5235 23335 5328
rect 23323 5201 23335 5235
rect 23289 5132 23335 5201
rect 23369 5281 23440 5296
rect 23369 5247 23393 5281
rect 23427 5247 23440 5281
rect 24516 5267 24550 5283
rect 24676 5343 24710 5359
rect 24676 5267 24710 5283
rect 23369 5235 23440 5247
rect 23369 5201 23391 5235
rect 23425 5201 23440 5235
rect 23369 5166 23440 5201
rect 24516 5205 24550 5221
rect 23289 5098 23440 5132
rect 24516 5129 24550 5145
rect 24676 5205 24710 5221
rect 24676 5129 24710 5145
rect 23032 5032 23066 5048
rect 22777 5024 22976 5030
rect 23100 5030 23116 5064
rect 23150 5030 23170 5064
rect 23209 5056 23220 5090
rect 23388 5090 23440 5098
rect 23209 5040 23254 5056
rect 23100 4988 23170 5030
rect 23288 5030 23304 5064
rect 23338 5030 23354 5064
rect 23422 5056 23440 5090
rect 23388 5040 23440 5056
rect 24516 5067 24550 5083
rect 23288 4988 23354 5030
rect 24516 4991 24550 5007
rect 24676 5067 24710 5083
rect 24676 4991 24710 5007
rect 11057 4930 11086 4988
rect 11120 4930 11178 4988
rect 11212 4930 11270 4988
rect 11304 4930 11362 4988
rect 11396 4930 11454 4988
rect 11488 4930 11546 4988
rect 11580 4930 11638 4988
rect 11672 4930 11730 4988
rect 11764 4930 11822 4988
rect 11856 4954 11894 4988
rect 11928 4964 11986 4988
rect 12020 4964 12078 4988
rect 12112 4964 12170 4988
rect 12204 4964 12262 4988
rect 12296 4964 12354 4988
rect 12388 4964 12446 4988
rect 12480 4964 12538 4988
rect 12572 4964 12630 4988
rect 12664 4964 12722 4988
rect 12756 4964 12814 4988
rect 12848 4964 12906 4988
rect 12940 4964 12998 4988
rect 13032 4964 13090 4988
rect 13124 4964 13182 4988
rect 13216 4964 13274 4988
rect 13308 4964 13366 4988
rect 13400 4964 13458 4988
rect 13492 4964 13550 4988
rect 13584 4964 13642 4988
rect 13676 4964 13734 4988
rect 13768 4964 13826 4988
rect 13860 4964 13918 4988
rect 13952 4964 14010 4988
rect 14044 4964 14102 4988
rect 14136 4964 14194 4988
rect 14228 4964 14286 4988
rect 14320 4964 14378 4988
rect 14412 4964 14470 4988
rect 14504 4964 14562 4988
rect 14596 4964 14654 4988
rect 14688 4964 14746 4988
rect 14780 4964 14838 4988
rect 14872 4964 14930 4988
rect 14964 4964 15022 4988
rect 15056 4964 15114 4988
rect 15148 4964 15206 4988
rect 15240 4964 15298 4988
rect 15332 4964 15390 4988
rect 15424 4964 15482 4988
rect 15516 4964 15574 4988
rect 15608 4964 15666 4988
rect 15700 4964 15758 4988
rect 15792 4964 15850 4988
rect 15884 4964 15942 4988
rect 15976 4964 16034 4988
rect 16068 4964 16126 4988
rect 16160 4964 16218 4988
rect 16252 4964 16310 4988
rect 16344 4964 16402 4988
rect 16436 4964 16494 4988
rect 16528 4964 16586 4988
rect 16620 4964 16678 4988
rect 16712 4964 16770 4988
rect 16804 4964 16862 4988
rect 16896 4964 16954 4988
rect 16988 4964 17046 4988
rect 17080 4964 17138 4988
rect 17172 4964 17230 4988
rect 17264 4964 17322 4988
rect 17356 4964 17414 4988
rect 17448 4964 17506 4988
rect 17540 4964 17598 4988
rect 17632 4964 17690 4988
rect 17724 4964 17782 4988
rect 17816 4964 17874 4988
rect 17908 4964 17966 4988
rect 18000 4964 18058 4988
rect 18092 4964 18150 4988
rect 18184 4964 18242 4988
rect 18276 4964 18334 4988
rect 18368 4964 18426 4988
rect 18460 4964 18518 4988
rect 18552 4964 18610 4988
rect 18644 4964 18702 4988
rect 18736 4964 18794 4988
rect 18828 4964 18886 4988
rect 18920 4964 18978 4988
rect 19012 4964 19070 4988
rect 19104 4964 19162 4988
rect 19196 4964 19254 4988
rect 19288 4964 19346 4988
rect 19380 4964 19438 4988
rect 19472 4964 19530 4988
rect 19564 4964 19622 4988
rect 19656 4964 19714 4988
rect 19748 4964 19806 4988
rect 19840 4964 19898 4988
rect 11948 4954 11986 4964
rect 12040 4954 12078 4964
rect 12132 4954 12170 4964
rect 12224 4954 12262 4964
rect 12316 4954 12354 4964
rect 12408 4954 12446 4964
rect 12500 4954 12538 4964
rect 12592 4954 12630 4964
rect 12684 4954 12722 4964
rect 12776 4954 12814 4964
rect 12868 4954 12906 4964
rect 12960 4954 12998 4964
rect 13052 4954 13090 4964
rect 13144 4954 13182 4964
rect 13236 4954 13274 4964
rect 13328 4954 13366 4964
rect 13420 4954 13458 4964
rect 13512 4954 13550 4964
rect 13604 4954 13642 4964
rect 13696 4954 13734 4964
rect 13788 4954 13826 4964
rect 13880 4954 13918 4964
rect 13972 4954 14010 4964
rect 14064 4954 14102 4964
rect 14156 4954 14194 4964
rect 14248 4954 14286 4964
rect 14340 4954 14378 4964
rect 14432 4954 14470 4964
rect 14524 4954 14562 4964
rect 14616 4954 14654 4964
rect 14708 4954 14746 4964
rect 14800 4954 14838 4964
rect 14892 4954 14930 4964
rect 14984 4954 15022 4964
rect 15076 4954 15114 4964
rect 15168 4954 15206 4964
rect 15260 4954 15298 4964
rect 15352 4954 15390 4964
rect 15444 4954 15482 4964
rect 15536 4954 15574 4964
rect 15628 4954 15666 4964
rect 15720 4954 15758 4964
rect 15812 4954 15850 4964
rect 15904 4954 15942 4964
rect 15996 4954 16034 4964
rect 16088 4954 16126 4964
rect 16180 4954 16218 4964
rect 16272 4954 16310 4964
rect 16364 4954 16402 4964
rect 16456 4954 16494 4964
rect 16548 4954 16586 4964
rect 16640 4954 16678 4964
rect 16732 4954 16770 4964
rect 16824 4954 16862 4964
rect 16916 4954 16954 4964
rect 17008 4954 17046 4964
rect 17100 4954 17138 4964
rect 17192 4954 17230 4964
rect 17284 4954 17322 4964
rect 17376 4954 17414 4964
rect 17468 4954 17506 4964
rect 17560 4954 17598 4964
rect 17652 4954 17690 4964
rect 17744 4954 17782 4964
rect 17836 4954 17874 4964
rect 17928 4954 17966 4964
rect 18020 4954 18058 4964
rect 18112 4954 18150 4964
rect 18204 4954 18242 4964
rect 18296 4954 18334 4964
rect 18388 4954 18426 4964
rect 18480 4954 18518 4964
rect 18572 4954 18610 4964
rect 18664 4954 18702 4964
rect 18756 4954 18794 4964
rect 18848 4954 18886 4964
rect 18940 4954 18978 4964
rect 19032 4954 19070 4964
rect 19124 4954 19162 4964
rect 19216 4954 19254 4964
rect 19308 4954 19346 4964
rect 19400 4954 19438 4964
rect 19492 4954 19530 4964
rect 19584 4954 19622 4964
rect 19676 4954 19714 4964
rect 19768 4954 19806 4964
rect 11856 4930 11914 4954
rect 11948 4930 12006 4954
rect 12040 4930 12098 4954
rect 12132 4930 12190 4954
rect 12224 4930 12282 4954
rect 12316 4930 12374 4954
rect 12408 4930 12466 4954
rect 12500 4930 12558 4954
rect 12592 4930 12650 4954
rect 12684 4930 12742 4954
rect 12776 4930 12834 4954
rect 12868 4930 12926 4954
rect 12960 4930 13018 4954
rect 13052 4930 13110 4954
rect 13144 4930 13202 4954
rect 13236 4930 13294 4954
rect 13328 4930 13386 4954
rect 13420 4930 13478 4954
rect 13512 4930 13570 4954
rect 13604 4930 13662 4954
rect 13696 4930 13754 4954
rect 13788 4930 13846 4954
rect 13880 4930 13938 4954
rect 13972 4930 14030 4954
rect 14064 4930 14122 4954
rect 14156 4930 14214 4954
rect 14248 4930 14306 4954
rect 14340 4930 14398 4954
rect 14432 4930 14490 4954
rect 14524 4930 14582 4954
rect 14616 4930 14674 4954
rect 14708 4930 14766 4954
rect 14800 4930 14858 4954
rect 14892 4930 14950 4954
rect 14984 4930 15042 4954
rect 15076 4930 15134 4954
rect 15168 4930 15226 4954
rect 15260 4930 15318 4954
rect 15352 4930 15410 4954
rect 15444 4930 15502 4954
rect 15536 4930 15594 4954
rect 15628 4930 15686 4954
rect 15720 4930 15778 4954
rect 15812 4930 15870 4954
rect 15904 4930 15962 4954
rect 15996 4930 16054 4954
rect 16088 4930 16146 4954
rect 16180 4930 16238 4954
rect 16272 4930 16330 4954
rect 16364 4930 16422 4954
rect 16456 4930 16514 4954
rect 16548 4930 16606 4954
rect 16640 4930 16698 4954
rect 16732 4930 16790 4954
rect 16824 4930 16882 4954
rect 16916 4930 16974 4954
rect 17008 4930 17066 4954
rect 17100 4930 17158 4954
rect 17192 4930 17250 4954
rect 17284 4930 17342 4954
rect 17376 4930 17434 4954
rect 17468 4930 17526 4954
rect 17560 4930 17618 4954
rect 17652 4930 17710 4954
rect 17744 4930 17802 4954
rect 17836 4930 17894 4954
rect 17928 4930 17986 4954
rect 18020 4930 18078 4954
rect 18112 4930 18170 4954
rect 18204 4930 18262 4954
rect 18296 4930 18354 4954
rect 18388 4930 18446 4954
rect 18480 4930 18538 4954
rect 18572 4930 18630 4954
rect 18664 4930 18722 4954
rect 18756 4930 18814 4954
rect 18848 4930 18906 4954
rect 18940 4930 18998 4954
rect 19032 4930 19090 4954
rect 19124 4930 19182 4954
rect 19216 4930 19274 4954
rect 19308 4930 19366 4954
rect 19400 4930 19458 4954
rect 19492 4930 19550 4954
rect 19584 4930 19642 4954
rect 19676 4930 19734 4954
rect 19768 4930 19826 4954
rect 19860 4930 19898 4964
rect 19932 4930 19990 4988
rect 20024 4930 20082 4988
rect 20116 4930 20174 4988
rect 20208 4930 20266 4988
rect 20300 4930 20358 4988
rect 20392 4930 20450 4988
rect 20484 4930 20542 4988
rect 20576 4930 20634 4988
rect 20668 4930 20726 4988
rect 20760 4930 20818 4988
rect 20852 4930 20910 4988
rect 20944 4930 21002 4988
rect 21036 4930 21094 4988
rect 21128 4930 21186 4988
rect 21220 4930 21278 4988
rect 21312 4930 21370 4988
rect 21404 4930 21462 4988
rect 21496 4930 21554 4988
rect 21588 4930 21646 4988
rect 21680 4930 21738 4988
rect 21772 4930 21830 4988
rect 21864 4930 21922 4988
rect 21956 4930 22014 4988
rect 22048 4930 22106 4988
rect 22140 4930 22198 4988
rect 22232 4930 22290 4988
rect 22324 4930 22382 4988
rect 22416 4930 22474 4988
rect 22508 4930 22566 4988
rect 22600 4930 22658 4988
rect 22692 4930 22750 4988
rect 22784 4930 22842 4988
rect 22876 4930 22934 4988
rect 22968 4930 23026 4988
rect 23060 4930 23118 4988
rect 23152 4930 23210 4988
rect 23244 4930 23302 4988
rect 23336 4930 23394 4988
rect 23428 4930 23457 4988
rect 24516 4929 24550 4945
rect 24516 4853 24550 4869
rect 24676 4929 24710 4945
rect 24676 4853 24710 4869
rect 24792 4915 24897 4950
rect 24792 4881 24824 4915
rect 24858 4881 24897 4915
rect 24792 4852 24897 4881
rect 24516 4791 24550 4807
rect 24516 4715 24550 4731
rect 24676 4797 24710 4807
rect 24806 4797 24883 4852
rect 24676 4791 24883 4797
rect 24710 4731 24883 4791
rect 24676 4728 24883 4731
rect 25191 4744 25523 4760
rect 24676 4715 24710 4728
rect 25191 4710 25217 4744
rect 25251 4710 25297 4744
rect 25331 4710 25377 4744
rect 25411 4710 25457 4744
rect 25491 4710 25523 4744
rect 25191 4692 25523 4710
rect 25923 4744 26255 4760
rect 25923 4710 25949 4744
rect 25983 4710 26029 4744
rect 26063 4710 26109 4744
rect 26143 4710 26189 4744
rect 26223 4710 26255 4744
rect 25923 4692 26255 4710
rect 26525 4744 26857 4760
rect 26525 4710 26557 4744
rect 26591 4710 26637 4744
rect 26671 4710 26717 4744
rect 26751 4710 26797 4744
rect 26831 4710 26857 4744
rect 26525 4692 26857 4710
rect 27135 4744 27467 4760
rect 27135 4710 27161 4744
rect 27195 4710 27241 4744
rect 27275 4710 27321 4744
rect 27355 4710 27401 4744
rect 27435 4710 27467 4744
rect 27135 4692 27467 4710
rect 27737 4744 28069 4760
rect 27737 4710 27769 4744
rect 27803 4710 27849 4744
rect 27883 4710 27929 4744
rect 27963 4710 28009 4744
rect 28043 4710 28069 4744
rect 27737 4692 28069 4710
rect 28473 4744 28805 4760
rect 28473 4710 28499 4744
rect 28533 4710 28579 4744
rect 28613 4710 28659 4744
rect 28693 4710 28739 4744
rect 28773 4710 28805 4744
rect 28473 4692 28805 4710
rect 29075 4744 29407 4760
rect 29075 4710 29107 4744
rect 29141 4710 29187 4744
rect 29221 4710 29267 4744
rect 29301 4710 29347 4744
rect 29381 4710 29407 4744
rect 29075 4692 29407 4710
rect 29809 4744 30141 4760
rect 29809 4710 29841 4744
rect 29875 4710 29921 4744
rect 29955 4710 30001 4744
rect 30035 4710 30081 4744
rect 30115 4710 30141 4744
rect 29809 4692 30141 4710
rect 11089 4624 11118 4692
rect 11152 4624 11210 4692
rect 11244 4624 11302 4692
rect 11336 4624 11394 4692
rect 11428 4624 11486 4692
rect 11520 4658 11577 4692
rect 11611 4658 11669 4692
rect 11703 4658 11762 4692
rect 11520 4624 11578 4658
rect 11612 4624 11670 4658
rect 11704 4624 11762 4658
rect 11796 4624 11854 4692
rect 11888 4657 11918 4692
rect 11888 4624 11917 4657
rect 13631 4625 13660 4683
rect 13694 4625 13752 4683
rect 13786 4625 13844 4683
rect 13878 4659 13936 4683
rect 13970 4659 14028 4683
rect 14062 4659 14120 4683
rect 14154 4659 14212 4683
rect 14246 4659 14304 4683
rect 14338 4659 14396 4683
rect 14430 4659 14488 4683
rect 14522 4659 14580 4683
rect 14614 4659 14672 4683
rect 14706 4659 14764 4683
rect 14798 4659 14856 4683
rect 14890 4659 14948 4683
rect 14982 4659 15040 4683
rect 15074 4659 15132 4683
rect 15166 4659 15224 4683
rect 15258 4659 15316 4683
rect 15350 4659 15408 4683
rect 13878 4625 13917 4659
rect 13970 4649 14009 4659
rect 14062 4649 14101 4659
rect 14154 4649 14193 4659
rect 14246 4649 14285 4659
rect 14338 4649 14377 4659
rect 14430 4649 14469 4659
rect 14522 4649 14561 4659
rect 14614 4649 14653 4659
rect 14706 4649 14745 4659
rect 14798 4649 14837 4659
rect 14890 4649 14929 4659
rect 14982 4649 15021 4659
rect 15074 4649 15113 4659
rect 15166 4649 15205 4659
rect 15258 4649 15297 4659
rect 15350 4649 15389 4659
rect 15442 4649 15481 4683
rect 13951 4625 14009 4649
rect 14043 4625 14101 4649
rect 14135 4625 14193 4649
rect 14227 4625 14285 4649
rect 14319 4625 14377 4649
rect 14411 4625 14469 4649
rect 14503 4625 14561 4649
rect 14595 4625 14653 4649
rect 14687 4625 14745 4649
rect 14779 4625 14837 4649
rect 14871 4625 14929 4649
rect 14963 4625 15021 4649
rect 15055 4625 15113 4649
rect 15147 4625 15205 4649
rect 15239 4625 15297 4649
rect 15331 4625 15389 4649
rect 15423 4625 15481 4649
rect 15515 4625 15573 4683
rect 15607 4625 15665 4683
rect 15699 4625 15757 4683
rect 15791 4625 15849 4683
rect 15883 4625 15941 4683
rect 15975 4625 16033 4683
rect 16067 4625 16125 4683
rect 16159 4625 16217 4683
rect 16251 4625 16309 4683
rect 16343 4625 16401 4683
rect 16435 4625 16493 4683
rect 16527 4625 16585 4683
rect 16619 4625 16677 4683
rect 16711 4625 16769 4683
rect 16803 4625 16861 4683
rect 16895 4625 16953 4683
rect 16987 4625 17045 4683
rect 17079 4625 17137 4683
rect 17171 4625 17229 4683
rect 17263 4625 17321 4683
rect 17355 4625 17413 4683
rect 17447 4625 17505 4683
rect 17539 4625 17597 4683
rect 17631 4625 17689 4683
rect 17723 4625 17781 4683
rect 17815 4625 17873 4683
rect 17907 4625 17965 4683
rect 17999 4625 18057 4683
rect 18091 4625 18149 4683
rect 18183 4625 18241 4683
rect 18275 4625 18333 4683
rect 18367 4625 18425 4683
rect 18459 4625 18517 4683
rect 18551 4625 18609 4683
rect 18643 4625 18701 4683
rect 18735 4625 18793 4683
rect 18827 4625 18885 4683
rect 18919 4625 18977 4683
rect 19011 4625 19069 4683
rect 19103 4625 19161 4683
rect 19195 4625 19253 4683
rect 19287 4625 19345 4683
rect 19379 4625 19437 4683
rect 19471 4625 19529 4683
rect 19563 4625 19621 4683
rect 19655 4625 19713 4683
rect 19747 4625 19805 4683
rect 19839 4625 19897 4683
rect 19931 4625 19989 4683
rect 20023 4625 20081 4683
rect 20115 4625 20173 4683
rect 20207 4625 20265 4683
rect 20299 4625 20357 4683
rect 20391 4625 20449 4683
rect 20483 4625 20541 4683
rect 20575 4625 20633 4683
rect 20667 4625 20725 4683
rect 20759 4625 20817 4683
rect 20851 4625 20909 4683
rect 20943 4625 21001 4683
rect 21035 4625 21093 4683
rect 21127 4625 21185 4683
rect 21219 4625 21277 4683
rect 21311 4625 21369 4683
rect 21403 4625 21461 4683
rect 21495 4625 21553 4683
rect 21587 4625 21645 4683
rect 21679 4625 21737 4683
rect 21771 4625 21829 4683
rect 21863 4625 21921 4683
rect 21955 4625 22013 4683
rect 22047 4625 22105 4683
rect 22139 4625 22197 4683
rect 22231 4625 22289 4683
rect 22323 4625 22381 4683
rect 22415 4625 22473 4683
rect 22507 4625 22565 4683
rect 22599 4625 22657 4683
rect 22691 4625 22749 4683
rect 22783 4625 22841 4683
rect 22875 4625 22933 4683
rect 22967 4625 23025 4683
rect 23059 4625 23117 4683
rect 23151 4625 23209 4683
rect 23243 4625 23301 4683
rect 23335 4625 23393 4683
rect 23427 4625 23456 4683
rect 11122 4574 11158 4590
rect 11122 4540 11124 4574
rect 11122 4506 11158 4540
rect 11122 4472 11124 4506
rect 11194 4574 11260 4624
rect 11194 4540 11210 4574
rect 11244 4540 11260 4574
rect 11194 4506 11260 4540
rect 11194 4472 11210 4506
rect 11244 4472 11260 4506
rect 11294 4574 11348 4590
rect 11294 4540 11296 4574
rect 11330 4540 11348 4574
rect 11294 4493 11348 4540
rect 11122 4438 11158 4472
rect 11294 4459 11296 4493
rect 11330 4459 11348 4493
rect 11122 4404 11257 4438
rect 11294 4409 11348 4459
rect 11223 4375 11257 4404
rect 11110 4346 11178 4368
rect 11110 4312 11126 4346
rect 11160 4345 11178 4346
rect 11110 4311 11128 4312
rect 11162 4311 11178 4345
rect 11110 4294 11178 4311
rect 11223 4359 11278 4375
rect 11223 4325 11244 4359
rect 11223 4309 11278 4325
rect 11312 4360 11348 4409
rect 11384 4576 11450 4590
rect 11384 4542 11400 4576
rect 11434 4542 11450 4576
rect 11384 4508 11450 4542
rect 11384 4474 11400 4508
rect 11434 4474 11450 4508
rect 11384 4440 11450 4474
rect 11484 4582 11532 4624
rect 11518 4548 11532 4582
rect 11484 4514 11532 4548
rect 11518 4480 11532 4514
rect 11484 4464 11532 4480
rect 11568 4560 11602 4590
rect 11568 4465 11602 4526
rect 11384 4406 11400 4440
rect 11434 4428 11450 4440
rect 11636 4582 11702 4624
rect 11636 4548 11652 4582
rect 11686 4548 11702 4582
rect 11636 4514 11702 4548
rect 11636 4480 11652 4514
rect 11686 4480 11702 4514
rect 11636 4464 11702 4480
rect 11736 4560 11770 4590
rect 11736 4465 11770 4526
rect 11434 4406 11527 4428
rect 11384 4394 11527 4406
rect 11312 4346 11459 4360
rect 11312 4312 11409 4346
rect 11443 4312 11459 4346
rect 11493 4346 11527 4394
rect 11568 4420 11602 4431
rect 11736 4420 11770 4431
rect 11568 4386 11770 4420
rect 11804 4582 11870 4624
rect 11804 4548 11820 4582
rect 11854 4548 11870 4582
rect 11804 4514 11870 4548
rect 11804 4480 11820 4514
rect 11854 4480 11870 4514
rect 11804 4446 11870 4480
rect 11804 4412 11820 4446
rect 11854 4412 11870 4446
rect 11804 4394 11870 4412
rect 13699 4583 13741 4625
rect 13699 4549 13707 4583
rect 13699 4515 13741 4549
rect 13699 4481 13707 4515
rect 13699 4447 13741 4481
rect 13699 4413 13707 4447
rect 13699 4397 13741 4413
rect 13775 4583 13841 4591
rect 13775 4549 13791 4583
rect 13825 4549 13841 4583
rect 13775 4515 13841 4549
rect 13775 4481 13791 4515
rect 13825 4481 13841 4515
rect 13775 4447 13841 4481
rect 13905 4575 13957 4591
rect 13905 4541 13923 4575
rect 13905 4507 13957 4541
rect 13991 4559 14057 4625
rect 13991 4525 14007 4559
rect 14041 4525 14057 4559
rect 14091 4575 14136 4591
rect 14125 4541 14136 4575
rect 13905 4473 13923 4507
rect 14091 4507 14136 4541
rect 14175 4559 14245 4625
rect 14175 4525 14195 4559
rect 14229 4525 14245 4559
rect 14279 4575 14313 4591
rect 14356 4548 14372 4582
rect 14406 4548 14522 4582
rect 13957 4489 14056 4491
rect 13957 4473 14010 4489
rect 13905 4457 14010 4473
rect 13775 4413 13791 4447
rect 13825 4426 13841 4447
rect 14044 4455 14056 4489
rect 13775 4395 13810 4413
rect 11671 4346 11770 4386
rect 13795 4392 13810 4395
rect 11493 4312 11543 4346
rect 11577 4312 11593 4346
rect 11671 4312 11733 4346
rect 11767 4312 11770 4346
rect 13623 4352 13761 4361
rect 13623 4318 13625 4352
rect 13659 4347 13761 4352
rect 13659 4318 13711 4347
rect 13623 4313 13711 4318
rect 13745 4313 13761 4347
rect 11223 4258 11257 4309
rect 11124 4224 11257 4258
rect 11312 4249 11348 4312
rect 11493 4278 11527 4312
rect 11671 4278 11770 4312
rect 11124 4203 11158 4224
rect 11296 4220 11348 4249
rect 11124 4148 11158 4169
rect 11194 4156 11210 4190
rect 11244 4156 11260 4190
rect 11194 4114 11260 4156
rect 11330 4186 11348 4220
rect 11296 4148 11348 4186
rect 11400 4244 11527 4278
rect 11568 4244 11770 4278
rect 11400 4226 11434 4244
rect 11568 4226 11602 4244
rect 11400 4148 11434 4192
rect 11470 4194 11518 4210
rect 11470 4160 11484 4194
rect 11470 4114 11518 4160
rect 11736 4226 11770 4244
rect 11568 4148 11602 4192
rect 11636 4194 11702 4210
rect 11636 4160 11652 4194
rect 11686 4160 11702 4194
rect 11636 4114 11702 4160
rect 11736 4148 11770 4192
rect 11804 4258 11870 4274
rect 11804 4224 11820 4258
rect 11854 4224 11870 4258
rect 11804 4190 11870 4224
rect 11804 4156 11820 4190
rect 11854 4156 11870 4190
rect 11804 4114 11870 4156
rect 13695 4263 13741 4279
rect 13795 4275 13841 4392
rect 13905 4362 13976 4423
rect 13905 4351 13920 4362
rect 13905 4317 13918 4351
rect 13954 4328 13976 4362
rect 13952 4317 13976 4328
rect 13905 4293 13976 4317
rect 14010 4362 14056 4455
rect 14010 4328 14022 4362
rect 13695 4229 13707 4263
rect 13695 4195 13741 4229
rect 13695 4161 13707 4195
rect 13695 4115 13741 4161
rect 13775 4263 13841 4275
rect 13775 4229 13791 4263
rect 13825 4229 13841 4263
rect 14010 4259 14056 4328
rect 13775 4195 13841 4229
rect 13775 4161 13791 4195
rect 13825 4161 13841 4195
rect 13905 4225 14056 4259
rect 14125 4473 14136 4507
rect 14279 4491 14313 4541
rect 14091 4285 14136 4473
rect 14091 4251 14102 4285
rect 13905 4217 13957 4225
rect 13905 4183 13923 4217
rect 14091 4217 14136 4251
rect 14170 4457 14313 4491
rect 14170 4263 14204 4457
rect 14354 4455 14378 4489
rect 14412 4463 14454 4489
rect 14412 4455 14420 4463
rect 14354 4429 14420 4455
rect 14238 4359 14320 4423
rect 14238 4349 14247 4359
rect 14281 4325 14320 4359
rect 14272 4315 14320 4325
rect 14238 4299 14320 4315
rect 14354 4413 14454 4429
rect 14354 4289 14398 4413
rect 14488 4379 14522 4548
rect 14570 4573 14646 4625
rect 14864 4583 14930 4625
rect 14570 4539 14586 4573
rect 14620 4539 14646 4573
rect 14706 4557 14740 4573
rect 14706 4505 14740 4523
rect 14864 4549 14880 4583
rect 14914 4549 14930 4583
rect 15353 4583 15429 4625
rect 14864 4515 14930 4549
rect 15139 4548 15155 4582
rect 15189 4548 15305 4582
rect 15353 4549 15369 4583
rect 15403 4549 15429 4583
rect 15617 4583 15894 4625
rect 15477 4557 15511 4573
rect 14556 4489 14826 4505
rect 14556 4463 14706 4489
rect 14590 4455 14706 4463
rect 14740 4455 14826 4489
rect 14864 4481 14880 4515
rect 14914 4481 14930 4515
rect 15101 4489 15148 4495
rect 14590 4429 14606 4455
rect 14556 4413 14606 4429
rect 14708 4379 14758 4395
rect 14488 4345 14724 4379
rect 14488 4337 14568 4345
rect 14170 4225 14313 4263
rect 14388 4255 14398 4289
rect 14354 4239 14398 4255
rect 14434 4267 14450 4301
rect 14484 4285 14500 4301
rect 14434 4251 14466 4267
rect 14434 4227 14500 4251
rect 13905 4167 13957 4183
rect 13775 4149 13841 4161
rect 13991 4157 14007 4191
rect 14041 4157 14057 4191
rect 14125 4183 14136 4217
rect 14279 4209 14313 4225
rect 14091 4167 14136 4183
rect 13991 4115 14057 4157
rect 14175 4157 14195 4191
rect 14229 4157 14245 4191
rect 14534 4191 14568 4337
rect 14714 4329 14758 4345
rect 14792 4311 14826 4455
rect 15101 4463 15114 4489
rect 15135 4429 15148 4455
rect 14860 4421 15061 4429
rect 14860 4387 15022 4421
rect 15056 4387 15061 4421
rect 15101 4413 15148 4429
rect 15196 4463 15237 4479
rect 15196 4429 15203 4463
rect 14860 4381 15061 4387
rect 14860 4379 14926 4381
rect 14860 4345 14876 4379
rect 14910 4345 14926 4379
rect 15196 4359 15237 4429
rect 15113 4353 15237 4359
rect 14988 4311 15004 4345
rect 15038 4311 15054 4345
rect 14606 4277 14622 4311
rect 14656 4291 14672 4311
rect 14656 4285 14688 4291
rect 14606 4251 14654 4277
rect 14792 4277 15054 4311
rect 15113 4319 15114 4353
rect 15148 4323 15237 4353
rect 15271 4379 15305 4548
rect 15617 4549 15633 4583
rect 15667 4549 15844 4583
rect 15878 4549 15894 4583
rect 15477 4515 15511 4523
rect 15928 4546 15985 4591
rect 15339 4481 15894 4515
rect 15339 4463 15389 4481
rect 15373 4429 15389 4463
rect 15339 4413 15389 4429
rect 15271 4363 15541 4379
rect 15271 4345 15507 4363
rect 15148 4319 15170 4323
rect 15113 4289 15170 4319
rect 14792 4251 14836 4277
rect 14606 4245 14688 4251
rect 14770 4217 14786 4251
rect 14820 4217 14836 4251
rect 15113 4255 15136 4289
rect 14870 4225 14904 4241
rect 15113 4239 15170 4255
rect 14279 4159 14313 4175
rect 14175 4115 14245 4157
rect 14369 4157 14385 4191
rect 14419 4157 14568 4191
rect 14369 4151 14568 4157
rect 14602 4187 14636 4203
rect 14602 4115 14636 4153
rect 14670 4173 14686 4207
rect 14720 4183 14736 4207
rect 15271 4191 15305 4345
rect 15497 4329 15507 4345
rect 15497 4313 15541 4329
rect 15380 4285 15399 4311
rect 15380 4251 15390 4285
rect 15433 4277 15455 4311
rect 15424 4251 15455 4277
rect 15575 4254 15611 4481
rect 15380 4245 15455 4251
rect 15545 4251 15611 4254
rect 15545 4217 15561 4251
rect 15595 4217 15611 4251
rect 15645 4421 15747 4447
rect 15645 4387 15666 4421
rect 15700 4413 15747 4421
rect 15781 4413 15797 4447
rect 15645 4379 15700 4387
rect 15679 4345 15700 4379
rect 15860 4363 15894 4481
rect 15962 4512 15985 4546
rect 15928 4478 15985 4512
rect 15962 4444 15985 4478
rect 15928 4424 15985 4444
rect 15645 4283 15700 4345
rect 15751 4352 15826 4363
rect 15751 4318 15766 4352
rect 15800 4351 15826 4352
rect 15751 4317 15776 4318
rect 15810 4317 15826 4351
rect 15860 4347 15910 4363
rect 15860 4313 15876 4347
rect 15860 4297 15910 4313
rect 15645 4249 15783 4283
rect 14870 4183 14904 4191
rect 14720 4173 14904 4183
rect 14670 4149 14904 4173
rect 14958 4157 14974 4191
rect 15008 4157 15024 4191
rect 14958 4115 15024 4157
rect 15152 4157 15168 4191
rect 15202 4157 15305 4191
rect 15152 4151 15305 4157
rect 15341 4187 15393 4203
rect 15341 4153 15359 4187
rect 15341 4115 15393 4153
rect 15445 4173 15461 4207
rect 15495 4183 15511 4207
rect 15645 4199 15679 4215
rect 15495 4173 15645 4183
rect 15445 4165 15645 4173
rect 15445 4149 15679 4165
rect 15736 4201 15783 4249
rect 15736 4167 15749 4201
rect 15736 4151 15783 4167
rect 15828 4191 15894 4259
rect 15944 4241 15985 4424
rect 15828 4157 15844 4191
rect 15878 4157 15894 4191
rect 15828 4115 15894 4157
rect 15928 4225 15985 4241
rect 15962 4191 15985 4225
rect 15928 4149 15985 4191
rect 16019 4565 16082 4581
rect 16019 4531 16032 4565
rect 16066 4531 16082 4565
rect 16019 4497 16082 4531
rect 16019 4463 16032 4497
rect 16066 4463 16082 4497
rect 16019 4363 16082 4463
rect 16118 4571 16177 4625
rect 16118 4537 16127 4571
rect 16161 4537 16177 4571
rect 16118 4503 16177 4537
rect 16118 4469 16127 4503
rect 16161 4469 16177 4503
rect 16118 4451 16177 4469
rect 16211 4547 16263 4591
rect 16245 4513 16263 4547
rect 16211 4479 16263 4513
rect 16245 4445 16263 4479
rect 16297 4575 16349 4591
rect 16297 4541 16315 4575
rect 16297 4507 16349 4541
rect 16383 4559 16449 4625
rect 16383 4525 16399 4559
rect 16433 4525 16449 4559
rect 16483 4575 16528 4591
rect 16517 4541 16528 4575
rect 16297 4473 16315 4507
rect 16483 4507 16528 4541
rect 16567 4559 16637 4625
rect 16567 4525 16587 4559
rect 16621 4525 16637 4559
rect 16671 4575 16705 4591
rect 16748 4548 16764 4582
rect 16798 4548 16914 4582
rect 16349 4489 16448 4491
rect 16349 4473 16402 4489
rect 16297 4457 16402 4473
rect 16211 4387 16263 4445
rect 16436 4455 16448 4489
rect 16220 4377 16263 4387
rect 16297 4377 16368 4423
rect 16019 4347 16186 4363
rect 16019 4313 16152 4347
rect 16019 4297 16186 4313
rect 16220 4362 16368 4377
rect 16220 4329 16312 4362
rect 16019 4217 16082 4297
rect 16220 4263 16263 4329
rect 16297 4328 16312 4329
rect 16346 4328 16368 4362
rect 16297 4293 16368 4328
rect 16402 4362 16448 4455
rect 16402 4328 16414 4362
rect 16019 4183 16032 4217
rect 16066 4183 16082 4217
rect 16211 4227 16263 4263
rect 16402 4259 16448 4328
rect 16019 4149 16082 4183
rect 16118 4191 16177 4207
rect 16118 4157 16127 4191
rect 16161 4157 16177 4191
rect 16118 4115 16177 4157
rect 16245 4193 16263 4227
rect 16211 4149 16263 4193
rect 16297 4225 16448 4259
rect 16517 4473 16528 4507
rect 16671 4491 16705 4541
rect 16483 4285 16528 4473
rect 16483 4251 16494 4285
rect 16297 4217 16349 4225
rect 16297 4183 16315 4217
rect 16483 4217 16528 4251
rect 16562 4457 16705 4491
rect 16562 4263 16596 4457
rect 16746 4455 16770 4489
rect 16804 4463 16846 4489
rect 16804 4455 16812 4463
rect 16746 4429 16812 4455
rect 16630 4355 16712 4423
rect 16630 4349 16663 4355
rect 16697 4321 16712 4355
rect 16664 4315 16712 4321
rect 16630 4299 16712 4315
rect 16746 4413 16846 4429
rect 16746 4289 16790 4413
rect 16880 4379 16914 4548
rect 16962 4573 17038 4625
rect 17256 4583 17322 4625
rect 16962 4539 16978 4573
rect 17012 4539 17038 4573
rect 17098 4557 17132 4573
rect 17098 4505 17132 4523
rect 17256 4549 17272 4583
rect 17306 4549 17322 4583
rect 17745 4583 17821 4625
rect 17256 4515 17322 4549
rect 17531 4548 17547 4582
rect 17581 4548 17697 4582
rect 17745 4549 17761 4583
rect 17795 4549 17821 4583
rect 18009 4583 18286 4625
rect 17869 4557 17903 4573
rect 16948 4489 17218 4505
rect 16948 4463 17098 4489
rect 16982 4455 17098 4463
rect 17132 4455 17218 4489
rect 17256 4481 17272 4515
rect 17306 4481 17322 4515
rect 17493 4489 17540 4495
rect 16982 4429 16998 4455
rect 16948 4413 16998 4429
rect 17100 4379 17150 4395
rect 16880 4345 17116 4379
rect 16880 4337 16960 4345
rect 16562 4225 16705 4263
rect 16780 4255 16790 4289
rect 16746 4239 16790 4255
rect 16826 4267 16842 4301
rect 16876 4285 16892 4301
rect 16826 4251 16858 4267
rect 16826 4227 16892 4251
rect 16297 4167 16349 4183
rect 16383 4157 16399 4191
rect 16433 4157 16449 4191
rect 16517 4183 16528 4217
rect 16671 4209 16705 4225
rect 16483 4167 16528 4183
rect 16383 4115 16449 4157
rect 16567 4157 16587 4191
rect 16621 4157 16637 4191
rect 16926 4191 16960 4337
rect 17106 4329 17150 4345
rect 17184 4311 17218 4455
rect 17493 4463 17506 4489
rect 17527 4429 17540 4455
rect 17252 4421 17453 4429
rect 17252 4387 17414 4421
rect 17448 4387 17453 4421
rect 17493 4413 17540 4429
rect 17588 4463 17629 4479
rect 17588 4429 17595 4463
rect 17252 4381 17453 4387
rect 17252 4379 17318 4381
rect 17252 4345 17268 4379
rect 17302 4345 17318 4379
rect 17588 4359 17629 4429
rect 17505 4353 17629 4359
rect 17380 4311 17396 4345
rect 17430 4311 17446 4345
rect 16998 4277 17014 4311
rect 17048 4291 17064 4311
rect 17048 4285 17080 4291
rect 16998 4251 17046 4277
rect 17184 4277 17446 4311
rect 17505 4319 17506 4353
rect 17540 4323 17629 4353
rect 17663 4379 17697 4548
rect 18009 4549 18025 4583
rect 18059 4549 18236 4583
rect 18270 4549 18286 4583
rect 17869 4515 17903 4523
rect 18320 4546 18377 4591
rect 17731 4481 18286 4515
rect 17731 4463 17781 4481
rect 17765 4429 17781 4463
rect 17731 4413 17781 4429
rect 17663 4363 17933 4379
rect 17663 4345 17899 4363
rect 17540 4319 17562 4323
rect 17505 4289 17562 4319
rect 17184 4251 17228 4277
rect 16998 4245 17080 4251
rect 17162 4217 17178 4251
rect 17212 4217 17228 4251
rect 17505 4255 17528 4289
rect 17262 4225 17296 4241
rect 17505 4239 17562 4255
rect 16671 4159 16705 4175
rect 16567 4115 16637 4157
rect 16761 4157 16777 4191
rect 16811 4157 16960 4191
rect 16761 4151 16960 4157
rect 16994 4187 17028 4203
rect 16994 4115 17028 4153
rect 17062 4173 17078 4207
rect 17112 4183 17128 4207
rect 17663 4191 17697 4345
rect 17889 4329 17899 4345
rect 17889 4313 17933 4329
rect 17772 4285 17791 4311
rect 17772 4251 17782 4285
rect 17825 4277 17847 4311
rect 17816 4251 17847 4277
rect 17967 4254 18003 4481
rect 17772 4245 17847 4251
rect 17937 4251 18003 4254
rect 17937 4217 17953 4251
rect 17987 4217 18003 4251
rect 18037 4421 18139 4447
rect 18037 4387 18058 4421
rect 18092 4413 18139 4421
rect 18173 4413 18189 4447
rect 18037 4379 18092 4387
rect 18071 4345 18092 4379
rect 18252 4363 18286 4481
rect 18354 4512 18377 4546
rect 18320 4478 18377 4512
rect 18354 4444 18377 4478
rect 18320 4424 18377 4444
rect 18037 4283 18092 4345
rect 18143 4360 18218 4363
rect 18143 4326 18156 4360
rect 18190 4351 18218 4360
rect 18143 4317 18168 4326
rect 18202 4317 18218 4351
rect 18252 4347 18302 4363
rect 18252 4313 18268 4347
rect 18252 4297 18302 4313
rect 18037 4249 18175 4283
rect 17262 4183 17296 4191
rect 17112 4173 17296 4183
rect 17062 4149 17296 4173
rect 17350 4157 17366 4191
rect 17400 4157 17416 4191
rect 17350 4115 17416 4157
rect 17544 4157 17560 4191
rect 17594 4157 17697 4191
rect 17544 4151 17697 4157
rect 17733 4187 17785 4203
rect 17733 4153 17751 4187
rect 17733 4115 17785 4153
rect 17837 4173 17853 4207
rect 17887 4183 17903 4207
rect 18037 4199 18071 4215
rect 17887 4173 18037 4183
rect 17837 4165 18037 4173
rect 17837 4149 18071 4165
rect 18128 4201 18175 4249
rect 18128 4167 18141 4201
rect 18128 4151 18175 4167
rect 18220 4191 18286 4259
rect 18336 4241 18377 4424
rect 18220 4157 18236 4191
rect 18270 4157 18286 4191
rect 18220 4115 18286 4157
rect 18320 4225 18377 4241
rect 18354 4191 18377 4225
rect 18320 4149 18377 4191
rect 18411 4565 18474 4581
rect 18411 4531 18424 4565
rect 18458 4531 18474 4565
rect 18411 4497 18474 4531
rect 18411 4463 18424 4497
rect 18458 4463 18474 4497
rect 18411 4363 18474 4463
rect 18510 4571 18569 4625
rect 18510 4537 18519 4571
rect 18553 4537 18569 4571
rect 18510 4503 18569 4537
rect 18510 4469 18519 4503
rect 18553 4469 18569 4503
rect 18510 4451 18569 4469
rect 18603 4547 18655 4591
rect 18637 4513 18655 4547
rect 18603 4479 18655 4513
rect 18637 4445 18655 4479
rect 18689 4575 18741 4591
rect 18689 4541 18707 4575
rect 18689 4507 18741 4541
rect 18775 4559 18841 4625
rect 18775 4525 18791 4559
rect 18825 4525 18841 4559
rect 18875 4575 18920 4591
rect 18909 4541 18920 4575
rect 18689 4473 18707 4507
rect 18875 4507 18920 4541
rect 18959 4559 19029 4625
rect 18959 4525 18979 4559
rect 19013 4525 19029 4559
rect 19063 4575 19097 4591
rect 19140 4548 19156 4582
rect 19190 4548 19306 4582
rect 18741 4489 18840 4491
rect 18741 4473 18794 4489
rect 18689 4457 18794 4473
rect 18603 4387 18655 4445
rect 18828 4455 18840 4489
rect 18612 4378 18655 4387
rect 18689 4378 18760 4423
rect 18411 4347 18578 4363
rect 18411 4313 18544 4347
rect 18411 4297 18578 4313
rect 18612 4362 18760 4378
rect 18612 4330 18704 4362
rect 18411 4217 18474 4297
rect 18612 4263 18655 4330
rect 18689 4328 18704 4330
rect 18738 4328 18760 4362
rect 18689 4293 18760 4328
rect 18794 4362 18840 4455
rect 18794 4328 18806 4362
rect 18411 4183 18424 4217
rect 18458 4183 18474 4217
rect 18603 4253 18655 4263
rect 18794 4259 18840 4328
rect 18603 4227 18612 4253
rect 18646 4219 18655 4253
rect 18411 4149 18474 4183
rect 18510 4191 18569 4207
rect 18510 4157 18519 4191
rect 18553 4157 18569 4191
rect 18510 4115 18569 4157
rect 18637 4193 18655 4219
rect 18603 4149 18655 4193
rect 18689 4225 18840 4259
rect 18909 4473 18920 4507
rect 19063 4491 19097 4541
rect 18875 4285 18920 4473
rect 18875 4251 18886 4285
rect 18689 4217 18741 4225
rect 18689 4183 18707 4217
rect 18875 4217 18920 4251
rect 18954 4457 19097 4491
rect 18954 4263 18988 4457
rect 19138 4455 19162 4489
rect 19196 4463 19238 4489
rect 19196 4455 19204 4463
rect 19138 4429 19204 4455
rect 19022 4355 19104 4423
rect 19022 4349 19050 4355
rect 19084 4321 19104 4355
rect 19056 4315 19104 4321
rect 19022 4299 19104 4315
rect 19138 4413 19238 4429
rect 19138 4289 19182 4413
rect 19272 4379 19306 4548
rect 19354 4573 19430 4625
rect 19648 4583 19714 4625
rect 19354 4539 19370 4573
rect 19404 4539 19430 4573
rect 19490 4557 19524 4573
rect 19490 4505 19524 4523
rect 19648 4549 19664 4583
rect 19698 4549 19714 4583
rect 20137 4583 20213 4625
rect 19648 4515 19714 4549
rect 19923 4548 19939 4582
rect 19973 4548 20089 4582
rect 20137 4549 20153 4583
rect 20187 4549 20213 4583
rect 20401 4583 20678 4625
rect 20261 4557 20295 4573
rect 19340 4489 19610 4505
rect 19340 4463 19490 4489
rect 19374 4455 19490 4463
rect 19524 4455 19610 4489
rect 19648 4481 19664 4515
rect 19698 4481 19714 4515
rect 19885 4489 19932 4495
rect 19374 4429 19390 4455
rect 19340 4413 19390 4429
rect 19492 4379 19542 4395
rect 19272 4345 19508 4379
rect 19272 4337 19352 4345
rect 18954 4225 19097 4263
rect 19172 4255 19182 4289
rect 19138 4239 19182 4255
rect 19218 4267 19234 4301
rect 19268 4285 19284 4301
rect 19218 4251 19250 4267
rect 19218 4227 19284 4251
rect 18689 4167 18741 4183
rect 18775 4157 18791 4191
rect 18825 4157 18841 4191
rect 18909 4183 18920 4217
rect 19063 4209 19097 4225
rect 18875 4167 18920 4183
rect 18775 4115 18841 4157
rect 18959 4157 18979 4191
rect 19013 4157 19029 4191
rect 19318 4191 19352 4337
rect 19498 4329 19542 4345
rect 19576 4311 19610 4455
rect 19885 4463 19898 4489
rect 19919 4429 19932 4455
rect 19644 4421 19845 4429
rect 19644 4387 19806 4421
rect 19840 4387 19845 4421
rect 19885 4413 19932 4429
rect 19980 4463 20021 4479
rect 19980 4429 19987 4463
rect 19644 4381 19845 4387
rect 19644 4379 19710 4381
rect 19644 4345 19660 4379
rect 19694 4345 19710 4379
rect 19980 4359 20021 4429
rect 19897 4353 20021 4359
rect 19772 4311 19788 4345
rect 19822 4311 19838 4345
rect 19390 4277 19406 4311
rect 19440 4291 19456 4311
rect 19440 4285 19472 4291
rect 19390 4251 19438 4277
rect 19576 4277 19838 4311
rect 19897 4319 19898 4353
rect 19932 4323 20021 4353
rect 20055 4379 20089 4548
rect 20401 4549 20417 4583
rect 20451 4549 20628 4583
rect 20662 4549 20678 4583
rect 20261 4515 20295 4523
rect 20712 4546 20769 4591
rect 20123 4481 20678 4515
rect 20123 4463 20173 4481
rect 20157 4429 20173 4463
rect 20123 4413 20173 4429
rect 20055 4363 20325 4379
rect 20055 4345 20291 4363
rect 19932 4319 19954 4323
rect 19897 4289 19954 4319
rect 19576 4251 19620 4277
rect 19390 4245 19472 4251
rect 19554 4217 19570 4251
rect 19604 4217 19620 4251
rect 19897 4255 19920 4289
rect 19654 4225 19688 4241
rect 19897 4239 19954 4255
rect 19063 4159 19097 4175
rect 18959 4115 19029 4157
rect 19153 4157 19169 4191
rect 19203 4157 19352 4191
rect 19153 4151 19352 4157
rect 19386 4187 19420 4203
rect 19386 4115 19420 4153
rect 19454 4173 19470 4207
rect 19504 4183 19520 4207
rect 20055 4191 20089 4345
rect 20281 4329 20291 4345
rect 20281 4313 20325 4329
rect 20164 4285 20183 4311
rect 20164 4251 20174 4285
rect 20217 4277 20239 4311
rect 20208 4251 20239 4277
rect 20359 4254 20395 4481
rect 20164 4245 20239 4251
rect 20329 4251 20395 4254
rect 20329 4217 20345 4251
rect 20379 4217 20395 4251
rect 20429 4421 20531 4447
rect 20429 4387 20450 4421
rect 20484 4413 20531 4421
rect 20565 4413 20581 4447
rect 20429 4379 20484 4387
rect 20463 4345 20484 4379
rect 20644 4363 20678 4481
rect 20746 4512 20769 4546
rect 20712 4478 20769 4512
rect 20746 4444 20769 4478
rect 20712 4424 20769 4444
rect 20429 4283 20484 4345
rect 20535 4356 20610 4363
rect 20535 4322 20547 4356
rect 20581 4351 20610 4356
rect 20535 4317 20560 4322
rect 20594 4317 20610 4351
rect 20644 4347 20694 4363
rect 20644 4313 20660 4347
rect 20644 4297 20694 4313
rect 20429 4249 20567 4283
rect 19654 4183 19688 4191
rect 19504 4173 19688 4183
rect 19454 4149 19688 4173
rect 19742 4157 19758 4191
rect 19792 4157 19808 4191
rect 19742 4115 19808 4157
rect 19936 4157 19952 4191
rect 19986 4157 20089 4191
rect 19936 4151 20089 4157
rect 20125 4187 20177 4203
rect 20125 4153 20143 4187
rect 20125 4115 20177 4153
rect 20229 4173 20245 4207
rect 20279 4183 20295 4207
rect 20429 4199 20463 4215
rect 20279 4173 20429 4183
rect 20229 4165 20429 4173
rect 20229 4149 20463 4165
rect 20520 4201 20567 4249
rect 20520 4167 20533 4201
rect 20520 4151 20567 4167
rect 20612 4191 20678 4259
rect 20728 4241 20769 4424
rect 20612 4157 20628 4191
rect 20662 4157 20678 4191
rect 20612 4115 20678 4157
rect 20712 4225 20769 4241
rect 20746 4191 20769 4225
rect 20712 4149 20769 4191
rect 20803 4565 20866 4581
rect 20803 4531 20816 4565
rect 20850 4531 20866 4565
rect 20803 4497 20866 4531
rect 20803 4463 20816 4497
rect 20850 4463 20866 4497
rect 20803 4363 20866 4463
rect 20902 4571 20961 4625
rect 20902 4537 20911 4571
rect 20945 4537 20961 4571
rect 20902 4503 20961 4537
rect 20902 4469 20911 4503
rect 20945 4469 20961 4503
rect 20902 4451 20961 4469
rect 20995 4547 21047 4591
rect 21029 4513 21047 4547
rect 20995 4479 21047 4513
rect 21029 4445 21047 4479
rect 21081 4575 21133 4591
rect 21081 4541 21099 4575
rect 21081 4507 21133 4541
rect 21167 4559 21233 4625
rect 21167 4525 21183 4559
rect 21217 4525 21233 4559
rect 21267 4575 21312 4591
rect 21301 4541 21312 4575
rect 21081 4473 21099 4507
rect 21267 4507 21312 4541
rect 21351 4559 21421 4625
rect 21351 4525 21371 4559
rect 21405 4525 21421 4559
rect 21455 4575 21489 4591
rect 21532 4548 21548 4582
rect 21582 4548 21698 4582
rect 21133 4489 21232 4491
rect 21133 4473 21186 4489
rect 21081 4457 21186 4473
rect 20995 4387 21047 4445
rect 21220 4455 21232 4489
rect 21004 4369 21047 4387
rect 21081 4369 21152 4423
rect 20803 4347 20970 4363
rect 20803 4313 20936 4347
rect 20803 4297 20970 4313
rect 21004 4362 21152 4369
rect 21004 4328 21096 4362
rect 21130 4328 21152 4362
rect 21004 4321 21152 4328
rect 20803 4217 20866 4297
rect 21004 4263 21047 4321
rect 21081 4293 21152 4321
rect 21186 4362 21232 4455
rect 21186 4328 21198 4362
rect 20803 4183 20816 4217
rect 20850 4183 20866 4217
rect 20995 4254 21047 4263
rect 21186 4259 21232 4328
rect 20995 4227 21004 4254
rect 21038 4220 21047 4254
rect 20803 4149 20866 4183
rect 20902 4191 20961 4207
rect 20902 4157 20911 4191
rect 20945 4157 20961 4191
rect 20902 4115 20961 4157
rect 21029 4193 21047 4220
rect 20995 4149 21047 4193
rect 21081 4225 21232 4259
rect 21301 4473 21312 4507
rect 21455 4491 21489 4541
rect 21267 4285 21312 4473
rect 21267 4251 21278 4285
rect 21081 4217 21133 4225
rect 21081 4183 21099 4217
rect 21267 4217 21312 4251
rect 21346 4457 21489 4491
rect 21346 4263 21380 4457
rect 21530 4455 21554 4489
rect 21588 4463 21630 4489
rect 21588 4455 21596 4463
rect 21530 4429 21596 4455
rect 21414 4354 21496 4423
rect 21414 4349 21453 4354
rect 21448 4320 21453 4349
rect 21487 4320 21496 4354
rect 21448 4315 21496 4320
rect 21414 4299 21496 4315
rect 21530 4413 21630 4429
rect 21530 4289 21574 4413
rect 21664 4379 21698 4548
rect 21746 4573 21822 4625
rect 22040 4583 22106 4625
rect 21746 4539 21762 4573
rect 21796 4539 21822 4573
rect 21882 4557 21916 4573
rect 21882 4505 21916 4523
rect 22040 4549 22056 4583
rect 22090 4549 22106 4583
rect 22529 4583 22605 4625
rect 22040 4515 22106 4549
rect 22315 4548 22331 4582
rect 22365 4548 22481 4582
rect 22529 4549 22545 4583
rect 22579 4549 22605 4583
rect 22793 4583 23070 4625
rect 22653 4557 22687 4573
rect 21732 4489 22002 4505
rect 21732 4463 21882 4489
rect 21766 4455 21882 4463
rect 21916 4455 22002 4489
rect 22040 4481 22056 4515
rect 22090 4481 22106 4515
rect 22277 4489 22324 4495
rect 21766 4429 21782 4455
rect 21732 4413 21782 4429
rect 21884 4379 21934 4395
rect 21664 4345 21900 4379
rect 21664 4337 21744 4345
rect 21346 4225 21489 4263
rect 21564 4255 21574 4289
rect 21530 4239 21574 4255
rect 21610 4267 21626 4301
rect 21660 4285 21676 4301
rect 21610 4251 21642 4267
rect 21610 4227 21676 4251
rect 21081 4167 21133 4183
rect 21167 4157 21183 4191
rect 21217 4157 21233 4191
rect 21301 4183 21312 4217
rect 21455 4209 21489 4225
rect 21267 4167 21312 4183
rect 21167 4115 21233 4157
rect 21351 4157 21371 4191
rect 21405 4157 21421 4191
rect 21710 4191 21744 4337
rect 21890 4329 21934 4345
rect 21968 4311 22002 4455
rect 22277 4463 22290 4489
rect 22311 4429 22324 4455
rect 22036 4421 22237 4429
rect 22036 4387 22198 4421
rect 22232 4387 22237 4421
rect 22277 4413 22324 4429
rect 22372 4463 22413 4479
rect 22372 4429 22379 4463
rect 22036 4381 22237 4387
rect 22036 4379 22102 4381
rect 22036 4345 22052 4379
rect 22086 4345 22102 4379
rect 22372 4359 22413 4429
rect 22289 4353 22413 4359
rect 22164 4311 22180 4345
rect 22214 4311 22230 4345
rect 21782 4277 21798 4311
rect 21832 4291 21848 4311
rect 21832 4285 21864 4291
rect 21782 4251 21830 4277
rect 21968 4277 22230 4311
rect 22289 4319 22290 4353
rect 22324 4323 22413 4353
rect 22447 4379 22481 4548
rect 22793 4549 22809 4583
rect 22843 4549 23020 4583
rect 23054 4549 23070 4583
rect 22653 4515 22687 4523
rect 23104 4546 23161 4591
rect 22515 4481 23070 4515
rect 22515 4463 22565 4481
rect 22549 4429 22565 4463
rect 22515 4413 22565 4429
rect 22447 4363 22717 4379
rect 22447 4345 22683 4363
rect 22324 4319 22346 4323
rect 22289 4289 22346 4319
rect 21968 4251 22012 4277
rect 21782 4245 21864 4251
rect 21946 4217 21962 4251
rect 21996 4217 22012 4251
rect 22289 4255 22312 4289
rect 22046 4225 22080 4241
rect 22289 4239 22346 4255
rect 21455 4159 21489 4175
rect 21351 4115 21421 4157
rect 21545 4157 21561 4191
rect 21595 4157 21744 4191
rect 21545 4151 21744 4157
rect 21778 4187 21812 4203
rect 21778 4115 21812 4153
rect 21846 4173 21862 4207
rect 21896 4183 21912 4207
rect 22447 4191 22481 4345
rect 22673 4329 22683 4345
rect 22673 4313 22717 4329
rect 22556 4285 22575 4311
rect 22556 4251 22566 4285
rect 22609 4277 22631 4311
rect 22600 4251 22631 4277
rect 22751 4254 22787 4481
rect 22556 4245 22631 4251
rect 22721 4251 22787 4254
rect 22721 4217 22737 4251
rect 22771 4217 22787 4251
rect 22821 4421 22923 4447
rect 22821 4387 22842 4421
rect 22876 4413 22923 4421
rect 22957 4413 22973 4447
rect 22821 4379 22876 4387
rect 22855 4345 22876 4379
rect 23036 4363 23070 4481
rect 23138 4512 23161 4546
rect 23104 4478 23161 4512
rect 23138 4444 23161 4478
rect 23104 4424 23161 4444
rect 22821 4283 22876 4345
rect 22927 4355 23002 4363
rect 22927 4321 22939 4355
rect 22973 4351 23002 4355
rect 22927 4317 22952 4321
rect 22986 4317 23002 4351
rect 23036 4347 23086 4363
rect 23036 4313 23052 4347
rect 23036 4297 23086 4313
rect 22821 4249 22959 4283
rect 22046 4183 22080 4191
rect 21896 4173 22080 4183
rect 21846 4149 22080 4173
rect 22134 4157 22150 4191
rect 22184 4157 22200 4191
rect 22134 4115 22200 4157
rect 22328 4157 22344 4191
rect 22378 4157 22481 4191
rect 22328 4151 22481 4157
rect 22517 4187 22569 4203
rect 22517 4153 22535 4187
rect 22517 4115 22569 4153
rect 22621 4173 22637 4207
rect 22671 4183 22687 4207
rect 22821 4199 22855 4215
rect 22671 4173 22821 4183
rect 22621 4165 22821 4173
rect 22621 4149 22855 4165
rect 22912 4201 22959 4249
rect 22912 4167 22925 4201
rect 22912 4151 22959 4167
rect 23004 4191 23070 4259
rect 23120 4241 23161 4424
rect 23004 4157 23020 4191
rect 23054 4157 23070 4191
rect 23004 4115 23070 4157
rect 23104 4225 23161 4241
rect 23138 4191 23161 4225
rect 23104 4149 23161 4191
rect 23195 4565 23258 4581
rect 23195 4531 23208 4565
rect 23242 4531 23258 4565
rect 23195 4497 23258 4531
rect 23195 4463 23208 4497
rect 23242 4463 23258 4497
rect 23195 4363 23258 4463
rect 23294 4571 23353 4625
rect 23294 4537 23303 4571
rect 23337 4537 23353 4571
rect 23294 4503 23353 4537
rect 23294 4469 23303 4503
rect 23337 4469 23353 4503
rect 23294 4451 23353 4469
rect 23387 4547 23439 4591
rect 23421 4513 23439 4547
rect 23387 4479 23439 4513
rect 23421 4445 23439 4479
rect 23387 4387 23439 4445
rect 23195 4347 23362 4363
rect 23195 4313 23328 4347
rect 23195 4297 23362 4313
rect 23195 4217 23258 4297
rect 23396 4263 23439 4387
rect 25577 4264 25606 4332
rect 25640 4264 25698 4332
rect 25732 4264 25790 4332
rect 25824 4264 25882 4332
rect 25916 4264 25974 4332
rect 26008 4264 26066 4332
rect 26100 4264 26158 4332
rect 26192 4264 26250 4332
rect 26284 4264 26342 4332
rect 26376 4298 26433 4332
rect 26467 4298 26526 4332
rect 26376 4264 26434 4298
rect 26468 4264 26526 4298
rect 26560 4264 26618 4332
rect 26652 4264 26710 4332
rect 26744 4264 26802 4332
rect 26836 4264 26894 4332
rect 26928 4264 26986 4332
rect 27020 4264 27078 4332
rect 27112 4264 27170 4332
rect 27204 4264 27262 4332
rect 27296 4264 27354 4332
rect 27388 4264 27446 4332
rect 27480 4264 27538 4332
rect 27572 4264 27630 4332
rect 27664 4264 27722 4332
rect 27756 4264 27814 4332
rect 27848 4264 27906 4332
rect 27940 4264 27998 4332
rect 28032 4264 28090 4332
rect 28124 4264 28182 4332
rect 28216 4264 28274 4332
rect 28308 4264 28366 4332
rect 28400 4264 28458 4332
rect 28492 4264 28550 4332
rect 28584 4264 28642 4332
rect 28676 4264 28734 4332
rect 28768 4264 28826 4332
rect 28860 4264 28918 4332
rect 28952 4264 29010 4332
rect 29044 4264 29102 4332
rect 29136 4264 29194 4332
rect 29228 4264 29286 4332
rect 29320 4264 29378 4332
rect 29412 4264 29470 4332
rect 29504 4264 29562 4332
rect 29596 4264 29654 4332
rect 29688 4264 29746 4332
rect 29780 4264 29838 4332
rect 29872 4264 29930 4332
rect 29964 4264 30022 4332
rect 30056 4264 30114 4332
rect 30148 4264 30206 4332
rect 30240 4264 30298 4332
rect 30332 4264 30361 4332
rect 23195 4183 23208 4217
rect 23242 4183 23258 4217
rect 23387 4257 23439 4263
rect 23387 4227 23394 4257
rect 23428 4223 23439 4257
rect 23195 4149 23258 4183
rect 23294 4191 23353 4207
rect 23294 4157 23303 4191
rect 23337 4157 23353 4191
rect 23294 4115 23353 4157
rect 23421 4193 23439 4223
rect 25680 4222 25746 4264
rect 23387 4149 23439 4193
rect 25594 4196 25646 4212
rect 25594 4162 25612 4196
rect 25680 4188 25696 4222
rect 25730 4188 25746 4222
rect 25864 4222 25934 4264
rect 25780 4196 25825 4212
rect 25594 4154 25646 4162
rect 25814 4162 25825 4196
rect 25864 4188 25884 4222
rect 25918 4188 25934 4222
rect 26058 4222 26257 4228
rect 25968 4204 26002 4220
rect 25594 4120 25745 4154
rect 11089 4080 11118 4114
rect 11152 4080 11210 4114
rect 11244 4080 11302 4114
rect 11336 4080 11394 4114
rect 11428 4080 11486 4114
rect 11520 4080 11578 4114
rect 11612 4080 11670 4114
rect 11704 4080 11762 4114
rect 11796 4080 11854 4114
rect 11888 4080 11917 4114
rect 13631 4091 13660 4115
rect 11089 4079 11917 4080
rect 11089 4045 11117 4079
rect 11151 4045 11210 4079
rect 11244 4045 11302 4079
rect 11336 4045 11394 4079
rect 11428 4045 11486 4079
rect 11520 4045 11578 4079
rect 11612 4045 11670 4079
rect 11704 4045 11762 4079
rect 11796 4045 11854 4079
rect 11888 4045 11917 4079
rect 13630 4057 13660 4091
rect 13694 4057 13752 4115
rect 13786 4057 13844 4115
rect 13878 4081 13917 4115
rect 13951 4091 14009 4115
rect 14043 4091 14101 4115
rect 14135 4091 14193 4115
rect 14227 4091 14285 4115
rect 14319 4091 14377 4115
rect 14411 4091 14469 4115
rect 14503 4091 14561 4115
rect 14595 4091 14653 4115
rect 14687 4091 14745 4115
rect 14779 4091 14837 4115
rect 14871 4091 14929 4115
rect 14963 4091 15021 4115
rect 15055 4091 15113 4115
rect 15147 4091 15205 4115
rect 15239 4091 15297 4115
rect 15331 4091 15389 4115
rect 15423 4091 15481 4115
rect 15515 4091 15573 4115
rect 15607 4091 15665 4115
rect 15699 4091 15757 4115
rect 15791 4091 15849 4115
rect 15883 4091 15941 4115
rect 15975 4091 16033 4115
rect 16067 4091 16125 4115
rect 16159 4091 16217 4115
rect 16251 4091 16309 4115
rect 16343 4091 16401 4115
rect 16435 4091 16493 4115
rect 16527 4091 16585 4115
rect 16619 4091 16677 4115
rect 16711 4091 16769 4115
rect 16803 4091 16861 4115
rect 16895 4091 16953 4115
rect 16987 4091 17045 4115
rect 17079 4091 17137 4115
rect 17171 4091 17229 4115
rect 17263 4091 17321 4115
rect 17355 4091 17413 4115
rect 17447 4091 17505 4115
rect 17539 4091 17597 4115
rect 17631 4091 17689 4115
rect 17723 4091 17781 4115
rect 17815 4091 17873 4115
rect 17907 4091 17965 4115
rect 17999 4091 18057 4115
rect 18091 4091 18149 4115
rect 18183 4091 18241 4115
rect 18275 4091 18333 4115
rect 18367 4091 18425 4115
rect 18459 4091 18517 4115
rect 18551 4091 18609 4115
rect 18643 4091 18701 4115
rect 18735 4091 18793 4115
rect 18827 4091 18885 4115
rect 18919 4091 18977 4115
rect 19011 4091 19069 4115
rect 19103 4091 19161 4115
rect 19195 4091 19253 4115
rect 19287 4091 19345 4115
rect 19379 4091 19437 4115
rect 19471 4091 19529 4115
rect 19563 4091 19621 4115
rect 19655 4091 19713 4115
rect 19747 4091 19805 4115
rect 19839 4091 19897 4115
rect 19931 4091 19989 4115
rect 20023 4091 20081 4115
rect 20115 4091 20173 4115
rect 20207 4091 20265 4115
rect 20299 4091 20357 4115
rect 20391 4091 20449 4115
rect 20483 4091 20541 4115
rect 20575 4091 20633 4115
rect 20667 4091 20725 4115
rect 20759 4091 20817 4115
rect 20851 4091 20909 4115
rect 20943 4091 21001 4115
rect 21035 4091 21093 4115
rect 21127 4091 21185 4115
rect 21219 4091 21277 4115
rect 21311 4091 21369 4115
rect 21403 4091 21461 4115
rect 21495 4091 21553 4115
rect 21587 4091 21645 4115
rect 21679 4091 21737 4115
rect 21771 4091 21829 4115
rect 21863 4091 21921 4115
rect 21955 4091 22013 4115
rect 22047 4091 22105 4115
rect 22139 4091 22197 4115
rect 22231 4091 22289 4115
rect 22323 4091 22381 4115
rect 22415 4091 22473 4115
rect 13970 4081 14009 4091
rect 14062 4081 14101 4091
rect 14154 4081 14193 4091
rect 14246 4081 14285 4091
rect 14338 4081 14377 4091
rect 14430 4081 14469 4091
rect 14522 4081 14561 4091
rect 14614 4081 14653 4091
rect 14706 4081 14745 4091
rect 14798 4081 14837 4091
rect 14890 4081 14929 4091
rect 14982 4081 15021 4091
rect 15074 4081 15113 4091
rect 15166 4081 15205 4091
rect 15258 4081 15297 4091
rect 15350 4081 15389 4091
rect 15442 4081 15481 4091
rect 15534 4081 15573 4091
rect 15626 4081 15665 4091
rect 15718 4081 15757 4091
rect 15810 4081 15849 4091
rect 15902 4081 15941 4091
rect 15994 4081 16033 4091
rect 16086 4081 16125 4091
rect 16178 4081 16217 4091
rect 16270 4081 16309 4091
rect 16362 4081 16401 4091
rect 16454 4081 16493 4091
rect 16546 4081 16585 4091
rect 16638 4081 16677 4091
rect 16730 4081 16769 4091
rect 16822 4081 16861 4091
rect 16914 4081 16953 4091
rect 17006 4081 17045 4091
rect 17098 4081 17137 4091
rect 17190 4081 17229 4091
rect 17282 4081 17321 4091
rect 17374 4081 17413 4091
rect 17466 4081 17505 4091
rect 17558 4081 17597 4091
rect 17650 4081 17689 4091
rect 17742 4081 17781 4091
rect 17834 4081 17873 4091
rect 17926 4081 17965 4091
rect 18018 4081 18057 4091
rect 18110 4081 18149 4091
rect 18202 4081 18241 4091
rect 18294 4081 18333 4091
rect 18386 4081 18425 4091
rect 18478 4081 18517 4091
rect 18570 4081 18609 4091
rect 18662 4081 18701 4091
rect 18754 4081 18793 4091
rect 18846 4081 18885 4091
rect 18938 4081 18977 4091
rect 19030 4081 19069 4091
rect 19122 4081 19161 4091
rect 19214 4081 19253 4091
rect 19306 4081 19345 4091
rect 19398 4081 19437 4091
rect 19490 4081 19529 4091
rect 19582 4081 19621 4091
rect 19674 4081 19713 4091
rect 19766 4081 19805 4091
rect 19858 4081 19897 4091
rect 19950 4081 19989 4091
rect 20042 4081 20081 4091
rect 20134 4081 20173 4091
rect 20226 4081 20265 4091
rect 13878 4057 13936 4081
rect 13970 4057 14028 4081
rect 14062 4057 14120 4081
rect 14154 4057 14212 4081
rect 14246 4057 14304 4081
rect 14338 4057 14396 4081
rect 14430 4057 14488 4081
rect 14522 4057 14580 4081
rect 14614 4057 14672 4081
rect 14706 4057 14764 4081
rect 14798 4057 14856 4081
rect 14890 4057 14948 4081
rect 14982 4057 15040 4081
rect 15074 4057 15132 4081
rect 15166 4057 15224 4081
rect 15258 4057 15316 4081
rect 15350 4057 15408 4081
rect 15442 4057 15500 4081
rect 15534 4057 15592 4081
rect 15626 4057 15684 4081
rect 15718 4057 15776 4081
rect 15810 4057 15868 4081
rect 15902 4057 15960 4081
rect 15994 4057 16052 4081
rect 16086 4057 16144 4081
rect 16178 4057 16236 4081
rect 16270 4057 16328 4081
rect 16362 4057 16420 4081
rect 16454 4057 16512 4081
rect 16546 4057 16604 4081
rect 16638 4057 16696 4081
rect 16730 4057 16788 4081
rect 16822 4057 16880 4081
rect 16914 4057 16972 4081
rect 17006 4057 17064 4081
rect 17098 4057 17156 4081
rect 17190 4057 17248 4081
rect 17282 4057 17340 4081
rect 17374 4057 17432 4081
rect 17466 4057 17524 4081
rect 17558 4057 17616 4081
rect 17650 4057 17708 4081
rect 17742 4057 17800 4081
rect 17834 4057 17892 4081
rect 17926 4057 17984 4081
rect 18018 4057 18076 4081
rect 18110 4057 18168 4081
rect 18202 4057 18260 4081
rect 18294 4057 18352 4081
rect 18386 4057 18444 4081
rect 18478 4057 18536 4081
rect 18570 4057 18628 4081
rect 18662 4057 18720 4081
rect 18754 4057 18812 4081
rect 18846 4057 18904 4081
rect 18938 4057 18996 4081
rect 19030 4057 19088 4081
rect 19122 4057 19180 4081
rect 19214 4057 19272 4081
rect 19306 4057 19364 4081
rect 19398 4057 19456 4081
rect 19490 4057 19548 4081
rect 19582 4057 19640 4081
rect 19674 4057 19732 4081
rect 19766 4057 19824 4081
rect 19858 4057 19916 4081
rect 19950 4057 20008 4081
rect 20042 4057 20100 4081
rect 20134 4057 20192 4081
rect 20226 4057 20284 4081
rect 20318 4057 20357 4091
rect 20410 4057 20449 4091
rect 20502 4057 20541 4091
rect 20594 4057 20633 4091
rect 20686 4057 20725 4091
rect 20778 4057 20817 4091
rect 20870 4057 20909 4091
rect 20962 4057 21001 4091
rect 21054 4057 21093 4091
rect 21146 4057 21185 4091
rect 21238 4057 21277 4091
rect 21330 4057 21369 4091
rect 21422 4057 21461 4091
rect 21514 4057 21553 4091
rect 21606 4057 21645 4091
rect 21698 4057 21737 4091
rect 21790 4057 21829 4091
rect 21882 4057 21921 4091
rect 21974 4057 22013 4091
rect 22066 4057 22105 4091
rect 22158 4057 22197 4091
rect 22250 4057 22289 4091
rect 22342 4057 22381 4091
rect 22434 4057 22473 4091
rect 22507 4057 22565 4115
rect 22599 4057 22657 4115
rect 22691 4057 22749 4115
rect 22783 4057 22841 4115
rect 22875 4057 22933 4115
rect 22967 4057 23025 4115
rect 23059 4057 23117 4115
rect 23151 4057 23209 4115
rect 23243 4057 23301 4115
rect 23335 4057 23393 4115
rect 23427 4081 23456 4115
rect 23427 4057 23455 4081
rect 25594 4072 25665 4086
rect 25594 4051 25623 4072
rect 25594 4017 25609 4051
rect 25657 4038 25665 4072
rect 25643 4017 25665 4038
rect 25594 3956 25665 4017
rect 25699 4051 25745 4120
rect 25699 4017 25711 4051
rect 25699 3924 25745 4017
rect 25594 3906 25699 3922
rect 25594 3872 25612 3906
rect 25646 3890 25699 3906
rect 25733 3890 25745 3924
rect 25646 3888 25745 3890
rect 25780 4128 25825 4162
rect 26058 4188 26074 4222
rect 26108 4188 26257 4222
rect 25968 4154 26002 4170
rect 25780 4094 25791 4128
rect 25780 3906 25825 4094
rect 25594 3838 25646 3872
rect 25814 3872 25825 3906
rect 25859 4116 26002 4154
rect 26043 4124 26087 4140
rect 25859 3922 25893 4116
rect 26077 4090 26087 4124
rect 25927 4064 26009 4080
rect 25961 4030 26009 4064
rect 25927 3998 26009 4030
rect 25927 3964 25943 3998
rect 25977 3964 26009 3998
rect 25927 3956 26009 3964
rect 26043 3966 26087 4090
rect 26123 4128 26189 4152
rect 26123 4112 26155 4128
rect 26123 4078 26139 4112
rect 26173 4078 26189 4094
rect 26223 4042 26257 4188
rect 26291 4226 26325 4264
rect 26291 4176 26325 4192
rect 26359 4206 26593 4230
rect 26359 4172 26375 4206
rect 26409 4196 26593 4206
rect 26409 4172 26425 4196
rect 26559 4188 26593 4196
rect 26647 4222 26713 4264
rect 26647 4188 26663 4222
rect 26697 4188 26713 4222
rect 26841 4222 26994 4228
rect 26841 4188 26857 4222
rect 26891 4188 26994 4222
rect 26295 4128 26377 4134
rect 26459 4128 26475 4162
rect 26509 4128 26525 4162
rect 26559 4138 26593 4154
rect 26295 4102 26343 4128
rect 26295 4068 26311 4102
rect 26345 4088 26377 4094
rect 26481 4102 26525 4128
rect 26802 4124 26859 4140
rect 26345 4068 26361 4088
rect 26481 4068 26743 4102
rect 26177 4034 26257 4042
rect 26403 4034 26447 4050
rect 26177 4000 26413 4034
rect 26043 3950 26143 3966
rect 26043 3924 26109 3950
rect 25859 3888 26002 3922
rect 26043 3890 26067 3924
rect 26101 3916 26109 3924
rect 26101 3890 26143 3916
rect 11496 3752 11525 3810
rect 11559 3752 11617 3810
rect 11651 3752 11709 3810
rect 11743 3752 11801 3810
rect 11835 3752 11893 3810
rect 11927 3752 11985 3810
rect 12019 3752 12077 3810
rect 12111 3752 12169 3810
rect 12203 3752 12261 3810
rect 12295 3752 12353 3810
rect 12387 3752 12445 3810
rect 12479 3752 12537 3810
rect 12571 3752 12629 3810
rect 12663 3752 12721 3810
rect 12755 3752 12813 3810
rect 12847 3752 12905 3810
rect 12939 3752 12997 3810
rect 13031 3752 13089 3810
rect 13123 3752 13181 3810
rect 13215 3752 13273 3810
rect 13307 3752 13365 3810
rect 13399 3752 13457 3810
rect 13491 3752 13549 3810
rect 13583 3752 13641 3810
rect 13675 3752 13733 3810
rect 13767 3752 13825 3810
rect 13859 3752 13917 3810
rect 13951 3752 14009 3810
rect 14043 3752 14101 3810
rect 14135 3752 14193 3810
rect 14227 3752 14285 3810
rect 14319 3752 14377 3810
rect 14411 3752 14469 3810
rect 14503 3752 14561 3810
rect 14595 3752 14653 3810
rect 14687 3752 14745 3810
rect 14779 3752 14837 3810
rect 14871 3752 14929 3810
rect 14963 3752 15021 3810
rect 15055 3752 15113 3810
rect 15147 3752 15205 3810
rect 15239 3752 15297 3810
rect 15331 3752 15389 3810
rect 15423 3752 15481 3810
rect 15515 3752 15573 3810
rect 15607 3752 15665 3810
rect 15699 3752 15757 3810
rect 15791 3752 15849 3810
rect 15883 3752 15941 3810
rect 15975 3752 16033 3810
rect 16067 3752 16125 3810
rect 16159 3752 16217 3810
rect 16251 3752 16309 3810
rect 16343 3752 16401 3810
rect 16435 3752 16493 3810
rect 16527 3752 16585 3810
rect 16619 3752 16677 3810
rect 16711 3752 16769 3810
rect 16803 3752 16861 3810
rect 16895 3752 16953 3810
rect 16987 3752 17045 3810
rect 17079 3752 17137 3810
rect 17171 3752 17229 3810
rect 17263 3752 17321 3810
rect 17355 3752 17413 3810
rect 17447 3752 17505 3810
rect 17539 3752 17597 3810
rect 17631 3752 17689 3810
rect 17723 3752 17781 3810
rect 17815 3752 17873 3810
rect 17907 3752 17965 3810
rect 17999 3752 18057 3810
rect 18091 3752 18149 3810
rect 18183 3752 18241 3810
rect 18275 3752 18333 3810
rect 18367 3752 18425 3810
rect 18459 3752 18517 3810
rect 18551 3752 18609 3810
rect 18643 3752 18701 3810
rect 18735 3752 18793 3810
rect 18827 3752 18885 3810
rect 18919 3752 18977 3810
rect 19011 3752 19069 3810
rect 19103 3752 19161 3810
rect 19195 3752 19253 3810
rect 19287 3752 19345 3810
rect 19379 3752 19437 3810
rect 19471 3752 19529 3810
rect 19563 3752 19621 3810
rect 19655 3752 19713 3810
rect 19747 3752 19805 3810
rect 19839 3752 19897 3810
rect 19931 3752 19989 3810
rect 20023 3752 20081 3810
rect 20115 3752 20173 3810
rect 20207 3752 20265 3810
rect 20299 3752 20357 3810
rect 20391 3752 20449 3810
rect 20483 3752 20541 3810
rect 20575 3752 20633 3810
rect 20667 3752 20725 3810
rect 20759 3752 20817 3810
rect 20851 3752 20909 3810
rect 20943 3752 21001 3810
rect 21035 3752 21093 3810
rect 21127 3752 21185 3810
rect 21219 3752 21277 3810
rect 21311 3752 21369 3810
rect 21403 3752 21461 3810
rect 21495 3752 21553 3810
rect 21587 3752 21645 3810
rect 21679 3752 21737 3810
rect 21771 3752 21829 3810
rect 21863 3752 21921 3810
rect 21955 3752 22013 3810
rect 22047 3752 22105 3810
rect 22139 3752 22197 3810
rect 22231 3752 22289 3810
rect 22323 3752 22381 3810
rect 22415 3752 22473 3810
rect 22507 3752 22565 3810
rect 22599 3752 22657 3810
rect 22691 3752 22749 3810
rect 22783 3752 22841 3810
rect 22875 3752 22933 3810
rect 22967 3752 23025 3810
rect 23059 3752 23117 3810
rect 23151 3752 23209 3810
rect 23243 3752 23301 3810
rect 23335 3752 23393 3810
rect 23427 3752 23456 3810
rect 25594 3804 25612 3838
rect 25594 3788 25646 3804
rect 25680 3820 25696 3854
rect 25730 3820 25746 3854
rect 25680 3754 25746 3820
rect 25780 3838 25825 3872
rect 25814 3804 25825 3838
rect 25780 3788 25825 3804
rect 25864 3820 25884 3854
rect 25918 3820 25934 3854
rect 25864 3754 25934 3820
rect 25968 3838 26002 3888
rect 26177 3831 26211 4000
rect 26397 3984 26447 4000
rect 26245 3950 26295 3966
rect 26279 3924 26295 3950
rect 26481 3924 26515 4068
rect 26677 4034 26693 4068
rect 26727 4034 26743 4068
rect 26802 4090 26825 4124
rect 26802 4060 26859 4090
rect 26549 4000 26565 4034
rect 26599 4000 26615 4034
rect 26802 4026 26803 4060
rect 26837 4056 26859 4060
rect 26837 4026 26926 4056
rect 26802 4020 26926 4026
rect 26549 3998 26615 4000
rect 26549 3992 26750 3998
rect 26549 3958 26711 3992
rect 26745 3958 26750 3992
rect 26549 3950 26750 3958
rect 26790 3950 26837 3966
rect 26279 3916 26395 3924
rect 26245 3890 26395 3916
rect 26429 3890 26515 3924
rect 26824 3924 26837 3950
rect 26245 3874 26515 3890
rect 26395 3856 26429 3874
rect 25968 3788 26002 3804
rect 26045 3797 26061 3831
rect 26095 3797 26211 3831
rect 26259 3806 26275 3840
rect 26309 3806 26335 3840
rect 26395 3806 26429 3822
rect 26553 3864 26569 3898
rect 26603 3864 26619 3898
rect 26790 3890 26803 3916
rect 26885 3950 26926 4020
rect 26885 3916 26892 3950
rect 26885 3900 26926 3916
rect 26960 4034 26994 4188
rect 27030 4226 27082 4264
rect 27030 4192 27048 4226
rect 27030 4176 27082 4192
rect 27134 4214 27368 4230
rect 27134 4206 27334 4214
rect 27134 4172 27150 4206
rect 27184 4196 27334 4206
rect 27184 4172 27200 4196
rect 27334 4164 27368 4180
rect 27425 4212 27472 4228
rect 27425 4178 27438 4212
rect 27069 4128 27144 4134
rect 27069 4094 27079 4128
rect 27113 4102 27144 4128
rect 27234 4128 27250 4162
rect 27284 4128 27300 4162
rect 27425 4130 27472 4178
rect 27234 4125 27300 4128
rect 27069 4068 27088 4094
rect 27122 4068 27144 4102
rect 27186 4050 27230 4066
rect 27186 4034 27196 4050
rect 26960 4016 27196 4034
rect 26960 4000 27230 4016
rect 26790 3884 26837 3890
rect 26553 3830 26619 3864
rect 26960 3831 26994 4000
rect 27028 3950 27078 3966
rect 27062 3916 27078 3950
rect 27028 3898 27078 3916
rect 27264 3898 27300 4125
rect 27334 4096 27472 4130
rect 27517 4222 27583 4264
rect 27517 4188 27533 4222
rect 27567 4188 27583 4222
rect 27517 4120 27583 4188
rect 27617 4188 27674 4230
rect 27651 4154 27674 4188
rect 27617 4138 27674 4154
rect 27334 4034 27389 4096
rect 27549 4066 27599 4082
rect 27368 4000 27389 4034
rect 27440 4057 27465 4062
rect 27440 4023 27462 4057
rect 27499 4028 27515 4062
rect 27496 4023 27515 4028
rect 27440 4016 27515 4023
rect 27549 4032 27565 4066
rect 27549 4016 27599 4032
rect 27334 3992 27389 4000
rect 27334 3958 27355 3992
rect 27389 3958 27436 3966
rect 27334 3932 27436 3958
rect 27470 3932 27486 3966
rect 27549 3898 27583 4016
rect 27633 3955 27674 4138
rect 27028 3864 27583 3898
rect 27617 3935 27674 3955
rect 27651 3901 27674 3935
rect 27617 3867 27674 3901
rect 26259 3754 26335 3806
rect 26553 3796 26569 3830
rect 26603 3796 26619 3830
rect 26828 3797 26844 3831
rect 26878 3797 26994 3831
rect 27166 3856 27200 3864
rect 26553 3754 26619 3796
rect 27042 3796 27058 3830
rect 27092 3796 27118 3830
rect 27651 3833 27674 3867
rect 27166 3806 27200 3822
rect 27042 3754 27118 3796
rect 27306 3796 27322 3830
rect 27356 3796 27533 3830
rect 27567 3796 27583 3830
rect 27306 3754 27583 3796
rect 27617 3788 27674 3833
rect 27708 4196 27771 4230
rect 27708 4162 27721 4196
rect 27755 4162 27771 4196
rect 27807 4222 27866 4264
rect 27807 4188 27816 4222
rect 27850 4188 27866 4222
rect 27807 4172 27866 4188
rect 27900 4186 27952 4230
rect 28072 4222 28138 4264
rect 27708 4082 27771 4162
rect 27934 4152 27952 4186
rect 27900 4116 27952 4152
rect 27986 4196 28038 4212
rect 27986 4162 28004 4196
rect 28072 4188 28088 4222
rect 28122 4188 28138 4222
rect 28256 4222 28326 4264
rect 28172 4196 28217 4212
rect 27986 4154 28038 4162
rect 28206 4162 28217 4196
rect 28256 4188 28276 4222
rect 28310 4188 28326 4222
rect 28450 4222 28649 4228
rect 28360 4204 28394 4220
rect 27986 4120 28137 4154
rect 27708 4066 27875 4082
rect 27708 4032 27841 4066
rect 27708 4016 27875 4032
rect 27708 3916 27771 4016
rect 27909 3992 27952 4116
rect 27900 3934 27952 3992
rect 27986 4051 28057 4086
rect 27986 4017 28001 4051
rect 28035 4027 28057 4051
rect 27986 3993 28012 4017
rect 28046 3993 28057 4027
rect 27986 3956 28057 3993
rect 28091 4051 28137 4120
rect 28091 4017 28103 4051
rect 27708 3882 27721 3916
rect 27755 3882 27771 3916
rect 27708 3848 27771 3882
rect 27708 3814 27721 3848
rect 27755 3814 27771 3848
rect 27708 3798 27771 3814
rect 27807 3910 27866 3928
rect 27807 3876 27816 3910
rect 27850 3876 27866 3910
rect 27807 3842 27866 3876
rect 27807 3808 27816 3842
rect 27850 3808 27866 3842
rect 27807 3754 27866 3808
rect 27934 3900 27952 3934
rect 28091 3924 28137 4017
rect 27900 3866 27952 3900
rect 27934 3860 27952 3866
rect 27900 3826 27910 3832
rect 27944 3826 27952 3860
rect 27900 3788 27952 3826
rect 27986 3906 28091 3922
rect 27986 3872 28004 3906
rect 28038 3890 28091 3906
rect 28125 3890 28137 3924
rect 28038 3888 28137 3890
rect 28172 4128 28217 4162
rect 28450 4188 28466 4222
rect 28500 4188 28649 4222
rect 28360 4154 28394 4170
rect 28172 4094 28183 4128
rect 28172 3906 28217 4094
rect 27986 3838 28038 3872
rect 28206 3872 28217 3906
rect 28251 4116 28394 4154
rect 28435 4124 28479 4140
rect 28251 3922 28285 4116
rect 28469 4090 28479 4124
rect 28319 4064 28401 4080
rect 28353 4060 28401 4064
rect 28319 4026 28345 4030
rect 28379 4026 28401 4060
rect 28319 3956 28401 4026
rect 28435 3966 28479 4090
rect 28515 4128 28581 4152
rect 28515 4112 28547 4128
rect 28515 4078 28531 4112
rect 28565 4078 28581 4094
rect 28615 4042 28649 4188
rect 28683 4226 28717 4264
rect 28683 4176 28717 4192
rect 28751 4206 28985 4230
rect 28751 4172 28767 4206
rect 28801 4196 28985 4206
rect 28801 4172 28817 4196
rect 28951 4188 28985 4196
rect 29039 4222 29105 4264
rect 29039 4188 29055 4222
rect 29089 4188 29105 4222
rect 29233 4222 29386 4228
rect 29233 4188 29249 4222
rect 29283 4188 29386 4222
rect 28687 4128 28769 4134
rect 28851 4128 28867 4162
rect 28901 4128 28917 4162
rect 28951 4138 28985 4154
rect 28687 4102 28735 4128
rect 28687 4068 28703 4102
rect 28737 4088 28769 4094
rect 28873 4102 28917 4128
rect 29194 4124 29251 4140
rect 28737 4068 28753 4088
rect 28873 4068 29135 4102
rect 28569 4034 28649 4042
rect 28795 4034 28839 4050
rect 28569 4000 28805 4034
rect 28435 3950 28535 3966
rect 28435 3924 28501 3950
rect 28251 3888 28394 3922
rect 28435 3890 28459 3924
rect 28493 3916 28501 3924
rect 28493 3890 28535 3916
rect 27986 3804 28004 3838
rect 27986 3788 28038 3804
rect 28072 3820 28088 3854
rect 28122 3820 28138 3854
rect 28072 3754 28138 3820
rect 28172 3838 28217 3872
rect 28206 3804 28217 3838
rect 28172 3788 28217 3804
rect 28256 3820 28276 3854
rect 28310 3820 28326 3854
rect 28256 3754 28326 3820
rect 28360 3838 28394 3888
rect 28569 3831 28603 4000
rect 28789 3984 28839 4000
rect 28637 3950 28687 3966
rect 28671 3924 28687 3950
rect 28873 3924 28907 4068
rect 29069 4034 29085 4068
rect 29119 4034 29135 4068
rect 29194 4090 29217 4124
rect 29194 4060 29251 4090
rect 28941 4000 28957 4034
rect 28991 4000 29007 4034
rect 29194 4026 29195 4060
rect 29229 4056 29251 4060
rect 29229 4026 29318 4056
rect 29194 4020 29318 4026
rect 28941 3998 29007 4000
rect 28941 3992 29142 3998
rect 28941 3958 29103 3992
rect 29137 3958 29142 3992
rect 28941 3950 29142 3958
rect 29182 3950 29229 3966
rect 28671 3916 28787 3924
rect 28637 3890 28787 3916
rect 28821 3890 28907 3924
rect 29216 3924 29229 3950
rect 28637 3874 28907 3890
rect 28787 3856 28821 3874
rect 28360 3788 28394 3804
rect 28437 3797 28453 3831
rect 28487 3797 28603 3831
rect 28651 3806 28667 3840
rect 28701 3806 28727 3840
rect 28787 3806 28821 3822
rect 28945 3864 28961 3898
rect 28995 3864 29011 3898
rect 29182 3890 29195 3916
rect 29277 3950 29318 4020
rect 29277 3916 29284 3950
rect 29277 3900 29318 3916
rect 29352 4034 29386 4188
rect 29422 4226 29474 4264
rect 29422 4192 29440 4226
rect 29422 4176 29474 4192
rect 29526 4214 29760 4230
rect 29526 4206 29726 4214
rect 29526 4172 29542 4206
rect 29576 4196 29726 4206
rect 29576 4172 29592 4196
rect 29726 4164 29760 4180
rect 29817 4212 29864 4228
rect 29817 4178 29830 4212
rect 29461 4128 29536 4134
rect 29461 4094 29471 4128
rect 29505 4102 29536 4128
rect 29626 4128 29642 4162
rect 29676 4128 29692 4162
rect 29817 4130 29864 4178
rect 29626 4125 29692 4128
rect 29461 4068 29480 4094
rect 29514 4068 29536 4102
rect 29578 4050 29622 4066
rect 29578 4034 29588 4050
rect 29352 4016 29588 4034
rect 29352 4000 29622 4016
rect 29182 3884 29229 3890
rect 28945 3830 29011 3864
rect 29352 3831 29386 4000
rect 29420 3950 29470 3966
rect 29454 3916 29470 3950
rect 29420 3898 29470 3916
rect 29656 3898 29692 4125
rect 29726 4096 29864 4130
rect 29909 4222 29975 4264
rect 29909 4188 29925 4222
rect 29959 4188 29975 4222
rect 29909 4120 29975 4188
rect 30009 4188 30066 4230
rect 30043 4154 30066 4188
rect 30009 4138 30066 4154
rect 29726 4034 29781 4096
rect 29941 4066 29991 4082
rect 29760 4000 29781 4034
rect 29832 4028 29857 4062
rect 29891 4061 29907 4062
rect 29832 4027 29861 4028
rect 29895 4027 29907 4061
rect 29832 4016 29907 4027
rect 29941 4032 29957 4066
rect 29941 4016 29991 4032
rect 29726 3992 29781 4000
rect 29726 3958 29747 3992
rect 29781 3958 29828 3966
rect 29726 3932 29828 3958
rect 29862 3932 29878 3966
rect 29941 3898 29975 4016
rect 30025 3955 30066 4138
rect 29420 3864 29975 3898
rect 30009 3935 30066 3955
rect 30043 3901 30066 3935
rect 30009 3867 30066 3901
rect 28651 3754 28727 3806
rect 28945 3796 28961 3830
rect 28995 3796 29011 3830
rect 29220 3797 29236 3831
rect 29270 3797 29386 3831
rect 29558 3856 29592 3864
rect 28945 3754 29011 3796
rect 29434 3796 29450 3830
rect 29484 3796 29510 3830
rect 30043 3833 30066 3867
rect 29558 3806 29592 3822
rect 29434 3754 29510 3796
rect 29698 3796 29714 3830
rect 29748 3796 29925 3830
rect 29959 3796 29975 3830
rect 29698 3754 29975 3796
rect 30009 3788 30066 3833
rect 30100 4196 30163 4230
rect 30100 4162 30113 4196
rect 30147 4162 30163 4196
rect 30199 4222 30258 4264
rect 30199 4188 30208 4222
rect 30242 4188 30258 4222
rect 30199 4172 30258 4188
rect 30292 4186 30344 4230
rect 30326 4177 30344 4186
rect 30100 4082 30163 4162
rect 30292 4143 30298 4152
rect 30332 4143 30344 4177
rect 30292 4116 30344 4143
rect 30100 4066 30267 4082
rect 30100 4032 30233 4066
rect 30100 4016 30267 4032
rect 30100 3916 30163 4016
rect 30301 3992 30344 4116
rect 30292 3934 30344 3992
rect 30100 3882 30113 3916
rect 30147 3882 30163 3916
rect 30100 3848 30163 3882
rect 30100 3814 30113 3848
rect 30147 3814 30163 3848
rect 30100 3798 30163 3814
rect 30199 3910 30258 3928
rect 30199 3876 30208 3910
rect 30242 3876 30258 3910
rect 30199 3842 30258 3876
rect 30199 3808 30208 3842
rect 30242 3808 30258 3842
rect 30199 3754 30258 3808
rect 30326 3900 30344 3934
rect 30292 3866 30344 3900
rect 30326 3832 30344 3866
rect 30292 3788 30344 3832
rect 11513 3674 11565 3718
rect 11513 3640 11531 3674
rect 11513 3606 11565 3640
rect 11513 3572 11531 3606
rect 11599 3698 11658 3752
rect 11599 3664 11615 3698
rect 11649 3664 11658 3698
rect 11599 3630 11658 3664
rect 11599 3596 11615 3630
rect 11649 3596 11658 3630
rect 11599 3578 11658 3596
rect 11694 3692 11757 3708
rect 11694 3658 11710 3692
rect 11744 3658 11757 3692
rect 11694 3624 11757 3658
rect 11694 3590 11710 3624
rect 11744 3590 11757 3624
rect 11513 3514 11565 3572
rect 11513 3390 11556 3514
rect 11694 3490 11757 3590
rect 11590 3474 11757 3490
rect 11624 3440 11757 3474
rect 11590 3424 11757 3440
rect 11513 3354 11565 3390
rect 11513 3353 11531 3354
rect 11513 3319 11522 3353
rect 11694 3344 11757 3424
rect 11556 3319 11565 3320
rect 11513 3276 11565 3319
rect 11599 3318 11658 3334
rect 11599 3284 11615 3318
rect 11649 3284 11658 3318
rect 11599 3242 11658 3284
rect 11694 3310 11710 3344
rect 11744 3310 11757 3344
rect 11694 3276 11757 3310
rect 11791 3673 11848 3718
rect 11882 3710 12159 3752
rect 11882 3676 11898 3710
rect 11932 3676 12109 3710
rect 12143 3676 12159 3710
rect 12347 3710 12423 3752
rect 12265 3684 12299 3700
rect 11791 3639 11814 3673
rect 12347 3676 12373 3710
rect 12407 3676 12423 3710
rect 12846 3710 12912 3752
rect 12265 3642 12299 3650
rect 12471 3675 12587 3709
rect 12621 3675 12637 3709
rect 12846 3676 12862 3710
rect 12896 3676 12912 3710
rect 13130 3700 13206 3752
rect 11791 3605 11848 3639
rect 11791 3571 11814 3605
rect 11791 3551 11848 3571
rect 11882 3608 12437 3642
rect 11791 3368 11832 3551
rect 11882 3490 11916 3608
rect 11979 3540 11995 3574
rect 12029 3548 12131 3574
rect 12029 3540 12076 3548
rect 12110 3514 12131 3548
rect 12076 3506 12131 3514
rect 11866 3474 11916 3490
rect 11900 3440 11916 3474
rect 11950 3478 12025 3490
rect 11950 3444 11966 3478
rect 12000 3444 12025 3478
rect 12076 3472 12097 3506
rect 11866 3424 11916 3440
rect 12076 3410 12131 3472
rect 11791 3352 11848 3368
rect 11791 3318 11814 3352
rect 11791 3276 11848 3318
rect 11882 3318 11948 3386
rect 11882 3284 11898 3318
rect 11932 3284 11948 3318
rect 11882 3242 11948 3284
rect 11993 3376 12131 3410
rect 12165 3381 12201 3608
rect 12387 3590 12437 3608
rect 12387 3556 12403 3590
rect 12387 3540 12437 3556
rect 12471 3506 12505 3675
rect 12846 3642 12912 3676
rect 12628 3616 12675 3622
rect 12235 3490 12505 3506
rect 12269 3472 12505 3490
rect 12269 3456 12279 3472
rect 12235 3440 12279 3456
rect 12321 3404 12343 3438
rect 12377 3412 12396 3438
rect 12165 3378 12231 3381
rect 11993 3328 12040 3376
rect 12165 3344 12181 3378
rect 12215 3344 12231 3378
rect 12321 3378 12352 3404
rect 12386 3378 12396 3412
rect 12321 3372 12396 3378
rect 12027 3294 12040 3328
rect 11993 3278 12040 3294
rect 12097 3326 12131 3342
rect 12265 3310 12281 3334
rect 12131 3300 12281 3310
rect 12315 3300 12331 3334
rect 12131 3292 12331 3300
rect 12097 3276 12331 3292
rect 12383 3314 12435 3330
rect 12417 3280 12435 3314
rect 12383 3242 12435 3280
rect 12471 3318 12505 3472
rect 12539 3590 12580 3606
rect 12573 3556 12580 3590
rect 12539 3486 12580 3556
rect 12662 3590 12675 3616
rect 12846 3608 12862 3642
rect 12896 3608 12912 3642
rect 13036 3684 13070 3700
rect 13130 3666 13156 3700
rect 13190 3666 13206 3700
rect 13254 3675 13370 3709
rect 13404 3675 13420 3709
rect 13463 3702 13497 3718
rect 13036 3632 13070 3650
rect 12950 3616 13220 3632
rect 12628 3556 12641 3582
rect 12950 3582 13036 3616
rect 13070 3590 13220 3616
rect 13070 3582 13186 3590
rect 12628 3540 12675 3556
rect 12715 3548 12916 3556
rect 12715 3514 12720 3548
rect 12754 3514 12916 3548
rect 12715 3508 12916 3514
rect 12850 3506 12916 3508
rect 12539 3480 12663 3486
rect 12539 3450 12628 3480
rect 12606 3446 12628 3450
rect 12662 3446 12663 3480
rect 12850 3472 12866 3506
rect 12900 3472 12916 3506
rect 12606 3416 12663 3446
rect 12640 3382 12663 3416
rect 12722 3438 12738 3472
rect 12772 3438 12788 3472
rect 12950 3438 12984 3582
rect 13170 3556 13186 3582
rect 13170 3540 13220 3556
rect 13018 3506 13068 3522
rect 13254 3506 13288 3675
rect 13463 3618 13497 3668
rect 13531 3686 13601 3752
rect 13531 3652 13547 3686
rect 13581 3652 13601 3686
rect 13640 3702 13685 3718
rect 13640 3668 13651 3702
rect 13640 3634 13685 3668
rect 13719 3686 13785 3752
rect 13719 3652 13735 3686
rect 13769 3652 13785 3686
rect 13819 3702 13871 3718
rect 13853 3668 13871 3702
rect 13322 3590 13364 3616
rect 13356 3582 13364 3590
rect 13398 3582 13422 3616
rect 13463 3584 13606 3618
rect 13356 3556 13422 3582
rect 13322 3540 13422 3556
rect 13052 3472 13288 3506
rect 13018 3456 13062 3472
rect 13208 3464 13288 3472
rect 12722 3404 12984 3438
rect 13104 3418 13120 3438
rect 12606 3366 12663 3382
rect 12940 3378 12984 3404
rect 13088 3412 13120 3418
rect 13154 3404 13170 3438
rect 13122 3378 13170 3404
rect 12872 3352 12906 3368
rect 12940 3344 12956 3378
rect 12990 3344 13006 3378
rect 13088 3372 13170 3378
rect 12471 3284 12574 3318
rect 12608 3284 12624 3318
rect 12471 3278 12624 3284
rect 12752 3284 12768 3318
rect 12802 3284 12818 3318
rect 12752 3242 12818 3284
rect 12872 3310 12906 3318
rect 13040 3310 13056 3334
rect 12872 3300 13056 3310
rect 13090 3300 13106 3334
rect 12872 3276 13106 3300
rect 13140 3314 13174 3330
rect 13140 3242 13174 3280
rect 13208 3318 13242 3464
rect 13276 3412 13292 3428
rect 13326 3394 13342 3428
rect 13310 3378 13342 3394
rect 13276 3354 13342 3378
rect 13378 3416 13422 3540
rect 13456 3538 13538 3550
rect 13456 3504 13478 3538
rect 13512 3504 13538 3538
rect 13456 3476 13538 3504
rect 13456 3442 13504 3476
rect 13456 3426 13538 3442
rect 13378 3382 13388 3416
rect 13572 3390 13606 3584
rect 13378 3366 13422 3382
rect 13463 3352 13606 3390
rect 13640 3600 13651 3634
rect 13819 3634 13871 3668
rect 13640 3412 13685 3600
rect 13674 3378 13685 3412
rect 13463 3336 13497 3352
rect 13208 3284 13357 3318
rect 13391 3284 13407 3318
rect 13640 3344 13685 3378
rect 13720 3616 13819 3618
rect 13720 3582 13732 3616
rect 13766 3600 13819 3616
rect 13853 3600 13871 3634
rect 13766 3584 13871 3600
rect 13905 3674 13957 3718
rect 13905 3640 13923 3674
rect 13905 3606 13957 3640
rect 13720 3489 13766 3582
rect 13905 3572 13923 3606
rect 13991 3698 14050 3752
rect 13991 3664 14007 3698
rect 14041 3664 14050 3698
rect 13991 3630 14050 3664
rect 13991 3596 14007 3630
rect 14041 3596 14050 3630
rect 13991 3578 14050 3596
rect 14086 3692 14149 3708
rect 14086 3658 14102 3692
rect 14136 3658 14149 3692
rect 14086 3624 14149 3658
rect 14086 3590 14102 3624
rect 14136 3590 14149 3624
rect 13754 3455 13766 3489
rect 13720 3386 13766 3455
rect 13800 3489 13871 3550
rect 13800 3455 13822 3489
rect 13856 3488 13871 3489
rect 13905 3514 13957 3572
rect 13905 3488 13948 3514
rect 14086 3490 14149 3590
rect 13856 3455 13948 3488
rect 13800 3440 13948 3455
rect 13800 3420 13871 3440
rect 13905 3390 13948 3440
rect 13982 3474 14149 3490
rect 14016 3440 14149 3474
rect 13982 3424 14149 3440
rect 13720 3352 13871 3386
rect 13463 3286 13497 3302
rect 13208 3278 13407 3284
rect 13531 3284 13547 3318
rect 13581 3284 13601 3318
rect 13640 3310 13651 3344
rect 13819 3344 13871 3352
rect 13640 3294 13685 3310
rect 13531 3242 13601 3284
rect 13719 3284 13735 3318
rect 13769 3284 13785 3318
rect 13853 3310 13871 3344
rect 13819 3294 13871 3310
rect 13905 3376 13957 3390
rect 13905 3342 13913 3376
rect 13947 3354 13957 3376
rect 13905 3320 13923 3342
rect 14086 3344 14149 3424
rect 13719 3242 13785 3284
rect 13905 3276 13957 3320
rect 13991 3318 14050 3334
rect 13991 3284 14007 3318
rect 14041 3284 14050 3318
rect 13991 3242 14050 3284
rect 14086 3310 14102 3344
rect 14136 3310 14149 3344
rect 14086 3276 14149 3310
rect 14183 3673 14240 3718
rect 14274 3710 14551 3752
rect 14274 3676 14290 3710
rect 14324 3676 14501 3710
rect 14535 3676 14551 3710
rect 14739 3710 14815 3752
rect 14657 3684 14691 3700
rect 14183 3639 14206 3673
rect 14739 3676 14765 3710
rect 14799 3676 14815 3710
rect 15238 3710 15304 3752
rect 14657 3642 14691 3650
rect 14863 3675 14979 3709
rect 15013 3675 15029 3709
rect 15238 3676 15254 3710
rect 15288 3676 15304 3710
rect 15522 3700 15598 3752
rect 14183 3605 14240 3639
rect 14183 3571 14206 3605
rect 14183 3551 14240 3571
rect 14274 3608 14829 3642
rect 14183 3368 14224 3551
rect 14274 3490 14308 3608
rect 14371 3540 14387 3574
rect 14421 3548 14523 3574
rect 14421 3540 14468 3548
rect 14502 3514 14523 3548
rect 14468 3506 14523 3514
rect 14258 3474 14308 3490
rect 14292 3440 14308 3474
rect 14342 3483 14417 3490
rect 14342 3478 14359 3483
rect 14342 3444 14358 3478
rect 14393 3449 14417 3483
rect 14392 3444 14417 3449
rect 14468 3472 14489 3506
rect 14258 3424 14308 3440
rect 14468 3410 14523 3472
rect 14183 3352 14240 3368
rect 14183 3318 14206 3352
rect 14183 3276 14240 3318
rect 14274 3318 14340 3386
rect 14274 3284 14290 3318
rect 14324 3284 14340 3318
rect 14274 3242 14340 3284
rect 14385 3376 14523 3410
rect 14557 3381 14593 3608
rect 14779 3590 14829 3608
rect 14779 3556 14795 3590
rect 14779 3540 14829 3556
rect 14863 3506 14897 3675
rect 15238 3642 15304 3676
rect 15020 3616 15067 3622
rect 14627 3490 14897 3506
rect 14661 3472 14897 3490
rect 14661 3456 14671 3472
rect 14627 3440 14671 3456
rect 14713 3404 14735 3438
rect 14769 3412 14788 3438
rect 14557 3378 14623 3381
rect 14385 3328 14432 3376
rect 14557 3344 14573 3378
rect 14607 3344 14623 3378
rect 14713 3378 14744 3404
rect 14778 3378 14788 3412
rect 14713 3372 14788 3378
rect 14419 3294 14432 3328
rect 14385 3278 14432 3294
rect 14489 3326 14523 3342
rect 14657 3310 14673 3334
rect 14523 3300 14673 3310
rect 14707 3300 14723 3334
rect 14523 3292 14723 3300
rect 14489 3276 14723 3292
rect 14775 3314 14827 3330
rect 14809 3280 14827 3314
rect 14775 3242 14827 3280
rect 14863 3318 14897 3472
rect 14931 3590 14972 3606
rect 14965 3556 14972 3590
rect 14931 3486 14972 3556
rect 15054 3590 15067 3616
rect 15238 3608 15254 3642
rect 15288 3608 15304 3642
rect 15428 3684 15462 3700
rect 15522 3666 15548 3700
rect 15582 3666 15598 3700
rect 15646 3675 15762 3709
rect 15796 3675 15812 3709
rect 15855 3702 15889 3718
rect 15428 3632 15462 3650
rect 15342 3616 15612 3632
rect 15020 3556 15033 3582
rect 15342 3582 15428 3616
rect 15462 3590 15612 3616
rect 15462 3582 15578 3590
rect 15020 3540 15067 3556
rect 15107 3548 15308 3556
rect 15107 3514 15112 3548
rect 15146 3514 15308 3548
rect 15107 3508 15308 3514
rect 15242 3506 15308 3508
rect 14931 3480 15055 3486
rect 14931 3450 15020 3480
rect 14998 3446 15020 3450
rect 15054 3446 15055 3480
rect 15242 3472 15258 3506
rect 15292 3472 15308 3506
rect 14998 3416 15055 3446
rect 15032 3382 15055 3416
rect 15114 3438 15130 3472
rect 15164 3438 15180 3472
rect 15342 3438 15376 3582
rect 15562 3556 15578 3582
rect 15562 3540 15612 3556
rect 15410 3506 15460 3522
rect 15646 3506 15680 3675
rect 15855 3618 15889 3668
rect 15923 3686 15993 3752
rect 15923 3652 15939 3686
rect 15973 3652 15993 3686
rect 16032 3702 16077 3718
rect 16032 3668 16043 3702
rect 16032 3634 16077 3668
rect 16111 3686 16177 3752
rect 16111 3652 16127 3686
rect 16161 3652 16177 3686
rect 16211 3702 16263 3718
rect 16245 3668 16263 3702
rect 15714 3590 15756 3616
rect 15748 3582 15756 3590
rect 15790 3582 15814 3616
rect 15855 3584 15998 3618
rect 15748 3556 15814 3582
rect 15714 3540 15814 3556
rect 15444 3472 15680 3506
rect 15410 3456 15454 3472
rect 15600 3464 15680 3472
rect 15114 3404 15376 3438
rect 15496 3418 15512 3438
rect 14998 3366 15055 3382
rect 15332 3378 15376 3404
rect 15480 3412 15512 3418
rect 15546 3404 15562 3438
rect 15514 3378 15562 3404
rect 15264 3352 15298 3368
rect 15332 3344 15348 3378
rect 15382 3344 15398 3378
rect 15480 3372 15562 3378
rect 14863 3284 14966 3318
rect 15000 3284 15016 3318
rect 14863 3278 15016 3284
rect 15144 3284 15160 3318
rect 15194 3284 15210 3318
rect 15144 3242 15210 3284
rect 15264 3310 15298 3318
rect 15432 3310 15448 3334
rect 15264 3300 15448 3310
rect 15482 3300 15498 3334
rect 15264 3276 15498 3300
rect 15532 3314 15566 3330
rect 15532 3242 15566 3280
rect 15600 3318 15634 3464
rect 15668 3412 15684 3428
rect 15718 3394 15734 3428
rect 15702 3378 15734 3394
rect 15668 3354 15734 3378
rect 15770 3416 15814 3540
rect 15848 3535 15930 3550
rect 15848 3501 15859 3535
rect 15893 3501 15930 3535
rect 15848 3476 15930 3501
rect 15848 3442 15896 3476
rect 15848 3426 15930 3442
rect 15770 3382 15780 3416
rect 15964 3390 15998 3584
rect 15770 3366 15814 3382
rect 15855 3352 15998 3390
rect 16032 3600 16043 3634
rect 16211 3634 16263 3668
rect 16032 3412 16077 3600
rect 16066 3378 16077 3412
rect 15855 3336 15889 3352
rect 15600 3284 15749 3318
rect 15783 3284 15799 3318
rect 16032 3344 16077 3378
rect 16112 3616 16211 3618
rect 16112 3582 16124 3616
rect 16158 3600 16211 3616
rect 16245 3600 16263 3634
rect 16158 3584 16263 3600
rect 16297 3674 16349 3718
rect 16297 3640 16315 3674
rect 16297 3606 16349 3640
rect 16112 3489 16158 3582
rect 16297 3572 16315 3606
rect 16383 3698 16442 3752
rect 16383 3664 16399 3698
rect 16433 3664 16442 3698
rect 16383 3630 16442 3664
rect 16383 3596 16399 3630
rect 16433 3596 16442 3630
rect 16383 3578 16442 3596
rect 16478 3692 16541 3708
rect 16478 3658 16494 3692
rect 16528 3658 16541 3692
rect 16478 3624 16541 3658
rect 16478 3590 16494 3624
rect 16528 3590 16541 3624
rect 16146 3455 16158 3489
rect 16112 3386 16158 3455
rect 16192 3491 16263 3550
rect 16297 3514 16349 3572
rect 16297 3491 16340 3514
rect 16192 3489 16340 3491
rect 16478 3490 16541 3590
rect 16192 3455 16214 3489
rect 16248 3455 16340 3489
rect 16192 3443 16340 3455
rect 16192 3420 16263 3443
rect 16297 3390 16340 3443
rect 16374 3474 16541 3490
rect 16408 3440 16541 3474
rect 16374 3424 16541 3440
rect 16112 3352 16263 3386
rect 15855 3286 15889 3302
rect 15600 3278 15799 3284
rect 15923 3284 15939 3318
rect 15973 3284 15993 3318
rect 16032 3310 16043 3344
rect 16211 3344 16263 3352
rect 16032 3294 16077 3310
rect 15923 3242 15993 3284
rect 16111 3284 16127 3318
rect 16161 3284 16177 3318
rect 16245 3310 16263 3344
rect 16211 3294 16263 3310
rect 16297 3375 16349 3390
rect 16297 3341 16304 3375
rect 16338 3354 16349 3375
rect 16297 3320 16315 3341
rect 16478 3344 16541 3424
rect 16111 3242 16177 3284
rect 16297 3276 16349 3320
rect 16383 3318 16442 3334
rect 16383 3284 16399 3318
rect 16433 3284 16442 3318
rect 16383 3242 16442 3284
rect 16478 3310 16494 3344
rect 16528 3310 16541 3344
rect 16478 3276 16541 3310
rect 16575 3673 16632 3718
rect 16666 3710 16943 3752
rect 16666 3676 16682 3710
rect 16716 3676 16893 3710
rect 16927 3676 16943 3710
rect 17131 3710 17207 3752
rect 17049 3684 17083 3700
rect 16575 3639 16598 3673
rect 17131 3676 17157 3710
rect 17191 3676 17207 3710
rect 17630 3710 17696 3752
rect 17049 3642 17083 3650
rect 17255 3675 17371 3709
rect 17405 3675 17421 3709
rect 17630 3676 17646 3710
rect 17680 3676 17696 3710
rect 17914 3700 17990 3752
rect 16575 3605 16632 3639
rect 16575 3571 16598 3605
rect 16575 3551 16632 3571
rect 16666 3608 17221 3642
rect 16575 3368 16616 3551
rect 16666 3490 16700 3608
rect 16763 3540 16779 3574
rect 16813 3548 16915 3574
rect 16813 3540 16860 3548
rect 16894 3514 16915 3548
rect 16860 3506 16915 3514
rect 16650 3474 16700 3490
rect 16684 3440 16700 3474
rect 16734 3483 16809 3490
rect 16734 3478 16753 3483
rect 16734 3444 16750 3478
rect 16787 3449 16809 3483
rect 16784 3444 16809 3449
rect 16860 3472 16881 3506
rect 16650 3424 16700 3440
rect 16860 3410 16915 3472
rect 16575 3352 16632 3368
rect 16575 3318 16598 3352
rect 16575 3276 16632 3318
rect 16666 3318 16732 3386
rect 16666 3284 16682 3318
rect 16716 3284 16732 3318
rect 16666 3242 16732 3284
rect 16777 3376 16915 3410
rect 16949 3381 16985 3608
rect 17171 3590 17221 3608
rect 17171 3556 17187 3590
rect 17171 3540 17221 3556
rect 17255 3506 17289 3675
rect 17630 3642 17696 3676
rect 17412 3616 17459 3622
rect 17019 3490 17289 3506
rect 17053 3472 17289 3490
rect 17053 3456 17063 3472
rect 17019 3440 17063 3456
rect 17105 3404 17127 3438
rect 17161 3412 17180 3438
rect 16949 3378 17015 3381
rect 16777 3328 16824 3376
rect 16949 3344 16965 3378
rect 16999 3344 17015 3378
rect 17105 3378 17136 3404
rect 17170 3378 17180 3412
rect 17105 3372 17180 3378
rect 16811 3294 16824 3328
rect 16777 3278 16824 3294
rect 16881 3326 16915 3342
rect 17049 3310 17065 3334
rect 16915 3300 17065 3310
rect 17099 3300 17115 3334
rect 16915 3292 17115 3300
rect 16881 3276 17115 3292
rect 17167 3314 17219 3330
rect 17201 3280 17219 3314
rect 17167 3242 17219 3280
rect 17255 3318 17289 3472
rect 17323 3590 17364 3606
rect 17357 3556 17364 3590
rect 17323 3486 17364 3556
rect 17446 3590 17459 3616
rect 17630 3608 17646 3642
rect 17680 3608 17696 3642
rect 17820 3684 17854 3700
rect 17914 3666 17940 3700
rect 17974 3666 17990 3700
rect 18038 3675 18154 3709
rect 18188 3675 18204 3709
rect 18247 3702 18281 3718
rect 17820 3632 17854 3650
rect 17734 3616 18004 3632
rect 17412 3556 17425 3582
rect 17734 3582 17820 3616
rect 17854 3590 18004 3616
rect 17854 3582 17970 3590
rect 17412 3540 17459 3556
rect 17499 3548 17700 3556
rect 17499 3514 17504 3548
rect 17538 3514 17700 3548
rect 17499 3508 17700 3514
rect 17634 3506 17700 3508
rect 17323 3480 17447 3486
rect 17323 3450 17412 3480
rect 17390 3446 17412 3450
rect 17446 3446 17447 3480
rect 17634 3472 17650 3506
rect 17684 3472 17700 3506
rect 17390 3416 17447 3446
rect 17424 3382 17447 3416
rect 17506 3438 17522 3472
rect 17556 3438 17572 3472
rect 17734 3438 17768 3582
rect 17954 3556 17970 3582
rect 17954 3540 18004 3556
rect 17802 3506 17852 3522
rect 18038 3506 18072 3675
rect 18247 3618 18281 3668
rect 18315 3686 18385 3752
rect 18315 3652 18331 3686
rect 18365 3652 18385 3686
rect 18424 3702 18469 3718
rect 18424 3668 18435 3702
rect 18424 3634 18469 3668
rect 18503 3686 18569 3752
rect 18503 3652 18519 3686
rect 18553 3652 18569 3686
rect 18603 3702 18655 3718
rect 18637 3668 18655 3702
rect 18106 3590 18148 3616
rect 18140 3582 18148 3590
rect 18182 3582 18206 3616
rect 18247 3584 18390 3618
rect 18140 3556 18206 3582
rect 18106 3540 18206 3556
rect 17836 3472 18072 3506
rect 17802 3456 17846 3472
rect 17992 3464 18072 3472
rect 17506 3404 17768 3438
rect 17888 3418 17904 3438
rect 17390 3366 17447 3382
rect 17724 3378 17768 3404
rect 17872 3412 17904 3418
rect 17938 3404 17954 3438
rect 17906 3378 17954 3404
rect 17656 3352 17690 3368
rect 17724 3344 17740 3378
rect 17774 3344 17790 3378
rect 17872 3372 17954 3378
rect 17255 3284 17358 3318
rect 17392 3284 17408 3318
rect 17255 3278 17408 3284
rect 17536 3284 17552 3318
rect 17586 3284 17602 3318
rect 17536 3242 17602 3284
rect 17656 3310 17690 3318
rect 17824 3310 17840 3334
rect 17656 3300 17840 3310
rect 17874 3300 17890 3334
rect 17656 3276 17890 3300
rect 17924 3314 17958 3330
rect 17924 3242 17958 3280
rect 17992 3318 18026 3464
rect 18060 3412 18076 3428
rect 18110 3394 18126 3428
rect 18094 3378 18126 3394
rect 18060 3354 18126 3378
rect 18162 3416 18206 3540
rect 18240 3539 18322 3550
rect 18240 3505 18250 3539
rect 18284 3505 18322 3539
rect 18240 3476 18322 3505
rect 18240 3442 18288 3476
rect 18240 3426 18322 3442
rect 18162 3382 18172 3416
rect 18356 3390 18390 3584
rect 18162 3366 18206 3382
rect 18247 3352 18390 3390
rect 18424 3600 18435 3634
rect 18603 3634 18655 3668
rect 18424 3412 18469 3600
rect 18458 3378 18469 3412
rect 18247 3336 18281 3352
rect 17992 3284 18141 3318
rect 18175 3284 18191 3318
rect 18424 3344 18469 3378
rect 18504 3616 18603 3618
rect 18504 3582 18516 3616
rect 18550 3600 18603 3616
rect 18637 3600 18655 3634
rect 18550 3584 18655 3600
rect 18689 3674 18741 3718
rect 18689 3640 18707 3674
rect 18689 3606 18741 3640
rect 18504 3489 18550 3582
rect 18689 3572 18707 3606
rect 18775 3698 18834 3752
rect 18775 3664 18791 3698
rect 18825 3664 18834 3698
rect 18775 3630 18834 3664
rect 18775 3596 18791 3630
rect 18825 3596 18834 3630
rect 18775 3578 18834 3596
rect 18870 3692 18933 3708
rect 18870 3658 18886 3692
rect 18920 3658 18933 3692
rect 18870 3624 18933 3658
rect 18870 3590 18886 3624
rect 18920 3590 18933 3624
rect 18538 3455 18550 3489
rect 18504 3386 18550 3455
rect 18584 3492 18655 3550
rect 18689 3514 18741 3572
rect 18689 3492 18732 3514
rect 18584 3489 18732 3492
rect 18870 3490 18933 3590
rect 18584 3455 18606 3489
rect 18640 3455 18732 3489
rect 18584 3444 18732 3455
rect 18584 3420 18655 3444
rect 18689 3390 18732 3444
rect 18766 3474 18933 3490
rect 18800 3440 18933 3474
rect 18766 3424 18933 3440
rect 18504 3352 18655 3386
rect 18247 3286 18281 3302
rect 17992 3278 18191 3284
rect 18315 3284 18331 3318
rect 18365 3284 18385 3318
rect 18424 3310 18435 3344
rect 18603 3344 18655 3352
rect 18424 3294 18469 3310
rect 18315 3242 18385 3284
rect 18503 3284 18519 3318
rect 18553 3284 18569 3318
rect 18637 3310 18655 3344
rect 18603 3294 18655 3310
rect 18689 3378 18741 3390
rect 18689 3344 18699 3378
rect 18733 3354 18741 3378
rect 18689 3320 18707 3344
rect 18870 3344 18933 3424
rect 18503 3242 18569 3284
rect 18689 3276 18741 3320
rect 18775 3318 18834 3334
rect 18775 3284 18791 3318
rect 18825 3284 18834 3318
rect 18775 3242 18834 3284
rect 18870 3310 18886 3344
rect 18920 3310 18933 3344
rect 18870 3276 18933 3310
rect 18967 3673 19024 3718
rect 19058 3710 19335 3752
rect 19058 3676 19074 3710
rect 19108 3676 19285 3710
rect 19319 3676 19335 3710
rect 19523 3710 19599 3752
rect 19441 3684 19475 3700
rect 18967 3639 18990 3673
rect 19523 3676 19549 3710
rect 19583 3676 19599 3710
rect 20022 3710 20088 3752
rect 19441 3642 19475 3650
rect 19647 3675 19763 3709
rect 19797 3675 19813 3709
rect 20022 3676 20038 3710
rect 20072 3676 20088 3710
rect 20306 3700 20382 3752
rect 18967 3605 19024 3639
rect 18967 3571 18990 3605
rect 18967 3551 19024 3571
rect 19058 3608 19613 3642
rect 18967 3368 19008 3551
rect 19058 3490 19092 3608
rect 19155 3540 19171 3574
rect 19205 3548 19307 3574
rect 19205 3540 19252 3548
rect 19286 3514 19307 3548
rect 19252 3506 19307 3514
rect 19042 3474 19092 3490
rect 19076 3440 19092 3474
rect 19126 3484 19201 3490
rect 19126 3478 19145 3484
rect 19126 3444 19142 3478
rect 19179 3450 19201 3484
rect 19176 3444 19201 3450
rect 19252 3472 19273 3506
rect 19042 3424 19092 3440
rect 19252 3410 19307 3472
rect 18967 3352 19024 3368
rect 18967 3318 18990 3352
rect 18967 3276 19024 3318
rect 19058 3318 19124 3386
rect 19058 3284 19074 3318
rect 19108 3284 19124 3318
rect 19058 3242 19124 3284
rect 19169 3376 19307 3410
rect 19341 3381 19377 3608
rect 19563 3590 19613 3608
rect 19563 3556 19579 3590
rect 19563 3540 19613 3556
rect 19647 3506 19681 3675
rect 20022 3642 20088 3676
rect 19804 3616 19851 3622
rect 19411 3490 19681 3506
rect 19445 3472 19681 3490
rect 19445 3456 19455 3472
rect 19411 3440 19455 3456
rect 19497 3404 19519 3438
rect 19553 3412 19572 3438
rect 19341 3378 19407 3381
rect 19169 3328 19216 3376
rect 19341 3344 19357 3378
rect 19391 3344 19407 3378
rect 19497 3378 19528 3404
rect 19562 3378 19572 3412
rect 19497 3372 19572 3378
rect 19203 3294 19216 3328
rect 19169 3278 19216 3294
rect 19273 3326 19307 3342
rect 19441 3310 19457 3334
rect 19307 3300 19457 3310
rect 19491 3300 19507 3334
rect 19307 3292 19507 3300
rect 19273 3276 19507 3292
rect 19559 3314 19611 3330
rect 19593 3280 19611 3314
rect 19559 3242 19611 3280
rect 19647 3318 19681 3472
rect 19715 3590 19756 3606
rect 19749 3556 19756 3590
rect 19715 3486 19756 3556
rect 19838 3590 19851 3616
rect 20022 3608 20038 3642
rect 20072 3608 20088 3642
rect 20212 3684 20246 3700
rect 20306 3666 20332 3700
rect 20366 3666 20382 3700
rect 20430 3675 20546 3709
rect 20580 3675 20596 3709
rect 20639 3702 20673 3718
rect 20212 3632 20246 3650
rect 20126 3616 20396 3632
rect 19804 3556 19817 3582
rect 20126 3582 20212 3616
rect 20246 3590 20396 3616
rect 20246 3582 20362 3590
rect 19804 3540 19851 3556
rect 19891 3548 20092 3556
rect 19891 3514 19896 3548
rect 19930 3514 20092 3548
rect 19891 3508 20092 3514
rect 20026 3506 20092 3508
rect 19715 3480 19839 3486
rect 19715 3450 19804 3480
rect 19782 3446 19804 3450
rect 19838 3446 19839 3480
rect 20026 3472 20042 3506
rect 20076 3472 20092 3506
rect 19782 3416 19839 3446
rect 19816 3382 19839 3416
rect 19898 3438 19914 3472
rect 19948 3438 19964 3472
rect 20126 3438 20160 3582
rect 20346 3556 20362 3582
rect 20346 3540 20396 3556
rect 20194 3506 20244 3522
rect 20430 3506 20464 3675
rect 20639 3618 20673 3668
rect 20707 3686 20777 3752
rect 20707 3652 20723 3686
rect 20757 3652 20777 3686
rect 20816 3702 20861 3718
rect 20816 3668 20827 3702
rect 20816 3634 20861 3668
rect 20895 3686 20961 3752
rect 20895 3652 20911 3686
rect 20945 3652 20961 3686
rect 20995 3702 21047 3718
rect 21029 3668 21047 3702
rect 20498 3590 20540 3616
rect 20532 3582 20540 3590
rect 20574 3582 20598 3616
rect 20639 3584 20782 3618
rect 20532 3556 20598 3582
rect 20498 3540 20598 3556
rect 20228 3472 20464 3506
rect 20194 3456 20238 3472
rect 20384 3464 20464 3472
rect 19898 3404 20160 3438
rect 20280 3418 20296 3438
rect 19782 3366 19839 3382
rect 20116 3378 20160 3404
rect 20264 3412 20296 3418
rect 20330 3404 20346 3438
rect 20298 3378 20346 3404
rect 20048 3352 20082 3368
rect 20116 3344 20132 3378
rect 20166 3344 20182 3378
rect 20264 3372 20346 3378
rect 19647 3284 19750 3318
rect 19784 3284 19800 3318
rect 19647 3278 19800 3284
rect 19928 3284 19944 3318
rect 19978 3284 19994 3318
rect 19928 3242 19994 3284
rect 20048 3310 20082 3318
rect 20216 3310 20232 3334
rect 20048 3300 20232 3310
rect 20266 3300 20282 3334
rect 20048 3276 20282 3300
rect 20316 3314 20350 3330
rect 20316 3242 20350 3280
rect 20384 3318 20418 3464
rect 20452 3412 20468 3428
rect 20502 3394 20518 3428
rect 20486 3378 20518 3394
rect 20452 3354 20518 3378
rect 20554 3416 20598 3540
rect 20632 3540 20714 3550
rect 20632 3506 20639 3540
rect 20673 3506 20714 3540
rect 20632 3476 20714 3506
rect 20632 3442 20680 3476
rect 20632 3426 20714 3442
rect 20554 3382 20564 3416
rect 20748 3390 20782 3584
rect 20554 3366 20598 3382
rect 20639 3352 20782 3390
rect 20816 3600 20827 3634
rect 20995 3634 21047 3668
rect 20816 3412 20861 3600
rect 20850 3378 20861 3412
rect 20639 3336 20673 3352
rect 20384 3284 20533 3318
rect 20567 3284 20583 3318
rect 20816 3344 20861 3378
rect 20896 3616 20995 3618
rect 20896 3582 20908 3616
rect 20942 3600 20995 3616
rect 21029 3600 21047 3634
rect 20942 3584 21047 3600
rect 21081 3674 21133 3718
rect 21081 3640 21099 3674
rect 21081 3606 21133 3640
rect 20896 3489 20942 3582
rect 21081 3572 21099 3606
rect 21167 3698 21226 3752
rect 21167 3664 21183 3698
rect 21217 3664 21226 3698
rect 21167 3630 21226 3664
rect 21167 3596 21183 3630
rect 21217 3596 21226 3630
rect 21167 3578 21226 3596
rect 21262 3692 21325 3708
rect 21262 3658 21278 3692
rect 21312 3658 21325 3692
rect 21262 3624 21325 3658
rect 21262 3590 21278 3624
rect 21312 3590 21325 3624
rect 20930 3455 20942 3489
rect 20896 3386 20942 3455
rect 20976 3489 21047 3550
rect 20976 3455 20998 3489
rect 21032 3481 21047 3489
rect 21081 3514 21133 3572
rect 21081 3481 21124 3514
rect 21262 3490 21325 3590
rect 21032 3455 21124 3481
rect 20976 3433 21124 3455
rect 20976 3420 21047 3433
rect 21081 3390 21124 3433
rect 21158 3474 21325 3490
rect 21192 3440 21325 3474
rect 21158 3424 21325 3440
rect 20896 3352 21047 3386
rect 20639 3286 20673 3302
rect 20384 3278 20583 3284
rect 20707 3284 20723 3318
rect 20757 3284 20777 3318
rect 20816 3310 20827 3344
rect 20995 3344 21047 3352
rect 20816 3294 20861 3310
rect 20707 3242 20777 3284
rect 20895 3284 20911 3318
rect 20945 3284 20961 3318
rect 21029 3310 21047 3344
rect 20995 3294 21047 3310
rect 21081 3376 21133 3390
rect 21081 3342 21088 3376
rect 21122 3354 21133 3376
rect 21081 3320 21099 3342
rect 21262 3344 21325 3424
rect 20895 3242 20961 3284
rect 21081 3276 21133 3320
rect 21167 3318 21226 3334
rect 21167 3284 21183 3318
rect 21217 3284 21226 3318
rect 21167 3242 21226 3284
rect 21262 3310 21278 3344
rect 21312 3310 21325 3344
rect 21262 3276 21325 3310
rect 21359 3673 21416 3718
rect 21450 3710 21727 3752
rect 21450 3676 21466 3710
rect 21500 3676 21677 3710
rect 21711 3676 21727 3710
rect 21915 3710 21991 3752
rect 21833 3684 21867 3700
rect 21359 3639 21382 3673
rect 21915 3676 21941 3710
rect 21975 3676 21991 3710
rect 22414 3710 22480 3752
rect 21833 3642 21867 3650
rect 22039 3675 22155 3709
rect 22189 3675 22205 3709
rect 22414 3676 22430 3710
rect 22464 3676 22480 3710
rect 22698 3700 22774 3752
rect 21359 3605 21416 3639
rect 21359 3571 21382 3605
rect 21359 3551 21416 3571
rect 21450 3608 22005 3642
rect 21359 3368 21400 3551
rect 21450 3490 21484 3608
rect 21547 3540 21563 3574
rect 21597 3548 21699 3574
rect 21597 3540 21644 3548
rect 21678 3514 21699 3548
rect 21644 3506 21699 3514
rect 21434 3474 21484 3490
rect 21468 3440 21484 3474
rect 21518 3485 21593 3490
rect 21518 3478 21538 3485
rect 21518 3444 21534 3478
rect 21572 3451 21593 3485
rect 21568 3444 21593 3451
rect 21644 3472 21665 3506
rect 21434 3424 21484 3440
rect 21644 3410 21699 3472
rect 21359 3352 21416 3368
rect 21359 3318 21382 3352
rect 21359 3276 21416 3318
rect 21450 3318 21516 3386
rect 21450 3284 21466 3318
rect 21500 3284 21516 3318
rect 21450 3242 21516 3284
rect 21561 3376 21699 3410
rect 21733 3381 21769 3608
rect 21955 3590 22005 3608
rect 21955 3556 21971 3590
rect 21955 3540 22005 3556
rect 22039 3506 22073 3675
rect 22414 3642 22480 3676
rect 22196 3616 22243 3622
rect 21803 3490 22073 3506
rect 21837 3472 22073 3490
rect 21837 3456 21847 3472
rect 21803 3440 21847 3456
rect 21889 3404 21911 3438
rect 21945 3412 21964 3438
rect 21733 3378 21799 3381
rect 21561 3328 21608 3376
rect 21733 3344 21749 3378
rect 21783 3344 21799 3378
rect 21889 3378 21920 3404
rect 21954 3378 21964 3412
rect 21889 3372 21964 3378
rect 21595 3294 21608 3328
rect 21561 3278 21608 3294
rect 21665 3326 21699 3342
rect 21833 3310 21849 3334
rect 21699 3300 21849 3310
rect 21883 3300 21899 3334
rect 21699 3292 21899 3300
rect 21665 3276 21899 3292
rect 21951 3314 22003 3330
rect 21985 3280 22003 3314
rect 21951 3242 22003 3280
rect 22039 3318 22073 3472
rect 22107 3590 22148 3606
rect 22141 3556 22148 3590
rect 22107 3486 22148 3556
rect 22230 3590 22243 3616
rect 22414 3608 22430 3642
rect 22464 3608 22480 3642
rect 22604 3684 22638 3700
rect 22698 3666 22724 3700
rect 22758 3666 22774 3700
rect 22822 3675 22938 3709
rect 22972 3675 22988 3709
rect 23031 3702 23065 3718
rect 22604 3632 22638 3650
rect 22518 3616 22788 3632
rect 22196 3556 22209 3582
rect 22518 3582 22604 3616
rect 22638 3590 22788 3616
rect 22638 3582 22754 3590
rect 22196 3540 22243 3556
rect 22283 3548 22484 3556
rect 22283 3514 22288 3548
rect 22322 3514 22484 3548
rect 22283 3508 22484 3514
rect 22418 3506 22484 3508
rect 22107 3480 22231 3486
rect 22107 3450 22196 3480
rect 22174 3446 22196 3450
rect 22230 3446 22231 3480
rect 22418 3472 22434 3506
rect 22468 3472 22484 3506
rect 22174 3416 22231 3446
rect 22208 3382 22231 3416
rect 22290 3438 22306 3472
rect 22340 3438 22356 3472
rect 22518 3438 22552 3582
rect 22738 3556 22754 3582
rect 22738 3540 22788 3556
rect 22586 3506 22636 3522
rect 22822 3506 22856 3675
rect 23031 3618 23065 3668
rect 23099 3686 23169 3752
rect 23099 3652 23115 3686
rect 23149 3652 23169 3686
rect 23208 3702 23253 3718
rect 23208 3668 23219 3702
rect 23208 3634 23253 3668
rect 23287 3686 23353 3752
rect 25577 3720 25606 3754
rect 25640 3720 25698 3754
rect 25732 3720 25790 3754
rect 25824 3720 25882 3754
rect 25916 3720 25974 3754
rect 26008 3720 26066 3754
rect 26100 3720 26158 3754
rect 26192 3720 26250 3754
rect 26284 3720 26342 3754
rect 26376 3720 26434 3754
rect 26468 3720 26526 3754
rect 26560 3720 26618 3754
rect 26652 3720 26710 3754
rect 26744 3720 26802 3754
rect 26836 3720 26894 3754
rect 26928 3720 26986 3754
rect 27020 3720 27078 3754
rect 27112 3720 27170 3754
rect 27204 3720 27262 3754
rect 27296 3720 27354 3754
rect 27388 3720 27446 3754
rect 27480 3720 27538 3754
rect 27572 3720 27630 3754
rect 27664 3720 27722 3754
rect 27756 3720 27814 3754
rect 27848 3720 27906 3754
rect 27940 3720 27998 3754
rect 28032 3720 28090 3754
rect 28124 3720 28182 3754
rect 28216 3720 28274 3754
rect 28308 3720 28366 3754
rect 28400 3720 28458 3754
rect 28492 3720 28550 3754
rect 28584 3720 28642 3754
rect 28676 3720 28734 3754
rect 28768 3720 28826 3754
rect 28860 3720 28918 3754
rect 28952 3720 29010 3754
rect 29044 3720 29102 3754
rect 29136 3720 29194 3754
rect 29228 3720 29286 3754
rect 29320 3720 29378 3754
rect 29412 3720 29470 3754
rect 29504 3720 29562 3754
rect 29596 3720 29654 3754
rect 29688 3720 29746 3754
rect 29780 3720 29838 3754
rect 29872 3720 29930 3754
rect 29964 3720 30022 3754
rect 30056 3720 30114 3754
rect 30148 3720 30206 3754
rect 30240 3720 30298 3754
rect 30332 3720 30361 3754
rect 23287 3652 23303 3686
rect 23337 3652 23353 3686
rect 23387 3702 23439 3718
rect 23421 3668 23439 3702
rect 22890 3590 22932 3616
rect 22924 3582 22932 3590
rect 22966 3582 22990 3616
rect 23031 3584 23174 3618
rect 22924 3556 22990 3582
rect 22890 3540 22990 3556
rect 22620 3472 22856 3506
rect 22586 3456 22630 3472
rect 22776 3464 22856 3472
rect 22290 3404 22552 3438
rect 22672 3418 22688 3438
rect 22174 3366 22231 3382
rect 22508 3378 22552 3404
rect 22656 3412 22688 3418
rect 22722 3404 22738 3438
rect 22690 3378 22738 3404
rect 22440 3352 22474 3368
rect 22508 3344 22524 3378
rect 22558 3344 22574 3378
rect 22656 3372 22738 3378
rect 22039 3284 22142 3318
rect 22176 3284 22192 3318
rect 22039 3278 22192 3284
rect 22320 3284 22336 3318
rect 22370 3284 22386 3318
rect 22320 3242 22386 3284
rect 22440 3310 22474 3318
rect 22608 3310 22624 3334
rect 22440 3300 22624 3310
rect 22658 3300 22674 3334
rect 22440 3276 22674 3300
rect 22708 3314 22742 3330
rect 22708 3242 22742 3280
rect 22776 3318 22810 3464
rect 22844 3412 22860 3428
rect 22894 3394 22910 3428
rect 22878 3378 22910 3394
rect 22844 3354 22910 3378
rect 22946 3416 22990 3540
rect 23024 3540 23106 3550
rect 23024 3506 23033 3540
rect 23067 3506 23106 3540
rect 23024 3476 23106 3506
rect 23024 3442 23072 3476
rect 23024 3426 23106 3442
rect 22946 3382 22956 3416
rect 23140 3390 23174 3584
rect 22946 3366 22990 3382
rect 23031 3352 23174 3390
rect 23208 3600 23219 3634
rect 23387 3634 23439 3668
rect 23208 3412 23253 3600
rect 23242 3378 23253 3412
rect 23031 3336 23065 3352
rect 22776 3284 22925 3318
rect 22959 3284 22975 3318
rect 23208 3344 23253 3378
rect 23288 3616 23387 3618
rect 23288 3582 23300 3616
rect 23334 3600 23387 3616
rect 23421 3600 23439 3634
rect 25577 3706 30361 3720
rect 25577 3672 25607 3706
rect 25641 3672 25698 3706
rect 25732 3672 25791 3706
rect 25825 3672 25882 3706
rect 25916 3672 25973 3706
rect 26007 3672 26067 3706
rect 26101 3672 26158 3706
rect 26192 3672 26251 3706
rect 26285 3672 26342 3706
rect 26376 3672 26434 3706
rect 26468 3672 26525 3706
rect 26559 3672 26618 3706
rect 26652 3672 26711 3706
rect 26745 3672 26802 3706
rect 26836 3672 26894 3706
rect 26928 3672 26986 3706
rect 27020 3672 27078 3706
rect 27112 3672 27170 3706
rect 27204 3672 27262 3706
rect 27296 3672 27354 3706
rect 27388 3672 27447 3706
rect 27481 3672 27537 3706
rect 27571 3672 27630 3706
rect 27664 3672 27723 3706
rect 27757 3672 27815 3706
rect 27849 3672 27906 3706
rect 27940 3672 27999 3706
rect 28033 3672 28091 3706
rect 28125 3672 28183 3706
rect 28217 3672 28275 3706
rect 28309 3672 28367 3706
rect 28401 3672 28459 3706
rect 28493 3672 28550 3706
rect 28584 3672 28641 3706
rect 28675 3672 28734 3706
rect 28768 3672 28827 3706
rect 28861 3672 28919 3706
rect 28953 3672 29010 3706
rect 29044 3672 29104 3706
rect 29138 3672 29194 3706
rect 29228 3672 29285 3706
rect 29319 3672 29378 3706
rect 29412 3672 29471 3706
rect 29505 3672 29563 3706
rect 29597 3672 29654 3706
rect 29688 3672 29746 3706
rect 29780 3672 29838 3706
rect 29872 3672 29929 3706
rect 29963 3672 30021 3706
rect 30055 3672 30114 3706
rect 30148 3672 30206 3706
rect 30240 3672 30298 3706
rect 30332 3672 30361 3706
rect 25577 3658 30361 3672
rect 25577 3624 25606 3658
rect 25640 3624 25698 3658
rect 25732 3624 25790 3658
rect 25824 3624 25882 3658
rect 25916 3624 25974 3658
rect 26008 3624 26066 3658
rect 26100 3624 26158 3658
rect 26192 3624 26250 3658
rect 26284 3624 26342 3658
rect 26376 3624 26434 3658
rect 26468 3624 26526 3658
rect 26560 3624 26618 3658
rect 26652 3624 26710 3658
rect 26744 3624 26802 3658
rect 26836 3624 26894 3658
rect 26928 3624 26986 3658
rect 27020 3624 27078 3658
rect 27112 3624 27170 3658
rect 27204 3624 27262 3658
rect 27296 3624 27354 3658
rect 27388 3624 27446 3658
rect 27480 3624 27538 3658
rect 27572 3624 27630 3658
rect 27664 3624 27722 3658
rect 27756 3624 27814 3658
rect 27848 3624 27906 3658
rect 27940 3624 27998 3658
rect 28032 3624 28090 3658
rect 28124 3624 28182 3658
rect 28216 3624 28274 3658
rect 28308 3624 28366 3658
rect 28400 3624 28458 3658
rect 28492 3624 28550 3658
rect 28584 3624 28642 3658
rect 28676 3624 28734 3658
rect 28768 3624 28826 3658
rect 28860 3624 28918 3658
rect 28952 3624 29010 3658
rect 29044 3624 29102 3658
rect 29136 3624 29194 3658
rect 29228 3624 29286 3658
rect 29320 3624 29378 3658
rect 29412 3624 29470 3658
rect 29504 3624 29562 3658
rect 29596 3624 29654 3658
rect 29688 3624 29746 3658
rect 29780 3624 29838 3658
rect 29872 3624 29930 3658
rect 29964 3624 30022 3658
rect 30056 3624 30114 3658
rect 30148 3624 30206 3658
rect 30240 3624 30298 3658
rect 30332 3624 30361 3658
rect 23334 3584 23439 3600
rect 23288 3489 23334 3582
rect 25594 3574 25646 3590
rect 23322 3455 23334 3489
rect 23288 3386 23334 3455
rect 23368 3489 23439 3550
rect 23368 3455 23390 3489
rect 23424 3455 23439 3489
rect 25594 3540 25612 3574
rect 25594 3506 25646 3540
rect 25680 3558 25746 3624
rect 25680 3524 25696 3558
rect 25730 3524 25746 3558
rect 25780 3574 25825 3590
rect 25814 3540 25825 3574
rect 25594 3472 25612 3506
rect 25780 3506 25825 3540
rect 25864 3558 25934 3624
rect 25864 3524 25884 3558
rect 25918 3524 25934 3558
rect 25968 3574 26002 3590
rect 26045 3547 26061 3581
rect 26095 3547 26211 3581
rect 25646 3488 25745 3490
rect 25646 3472 25699 3488
rect 25594 3456 25699 3472
rect 23368 3420 23439 3455
rect 25733 3454 25745 3488
rect 25594 3388 25618 3422
rect 25652 3388 25665 3422
rect 23288 3352 23439 3386
rect 23031 3286 23065 3302
rect 22776 3278 22975 3284
rect 23099 3284 23115 3318
rect 23149 3284 23169 3318
rect 23208 3310 23219 3344
rect 23387 3344 23439 3352
rect 23208 3294 23253 3310
rect 23099 3242 23169 3284
rect 23287 3284 23303 3318
rect 23337 3284 23353 3318
rect 23421 3310 23439 3344
rect 23387 3294 23439 3310
rect 25594 3361 25665 3388
rect 25594 3327 25609 3361
rect 25643 3327 25665 3361
rect 25594 3292 25665 3327
rect 25699 3361 25745 3454
rect 25699 3327 25711 3361
rect 23287 3242 23353 3284
rect 25699 3258 25745 3327
rect 11496 3184 11525 3242
rect 11559 3184 11617 3242
rect 11651 3184 11709 3242
rect 11743 3184 11801 3242
rect 11835 3184 11893 3242
rect 11927 3184 11985 3242
rect 12019 3184 12077 3242
rect 12111 3184 12169 3242
rect 12203 3184 12261 3242
rect 12295 3184 12353 3242
rect 12387 3184 12445 3242
rect 12479 3184 12537 3242
rect 12571 3184 12629 3242
rect 12663 3184 12721 3242
rect 12755 3184 12813 3242
rect 12847 3184 12905 3242
rect 12939 3184 12997 3242
rect 13031 3184 13089 3242
rect 13123 3184 13181 3242
rect 13215 3184 13273 3242
rect 13307 3184 13365 3242
rect 13399 3184 13457 3242
rect 13491 3184 13549 3242
rect 13583 3184 13641 3242
rect 13675 3184 13733 3242
rect 13767 3184 13825 3242
rect 13859 3184 13917 3242
rect 13951 3184 14009 3242
rect 14043 3184 14101 3242
rect 14135 3184 14193 3242
rect 14227 3184 14285 3242
rect 14319 3184 14377 3242
rect 14411 3184 14469 3242
rect 14503 3184 14561 3242
rect 14595 3184 14653 3242
rect 14687 3184 14745 3242
rect 14779 3184 14837 3242
rect 14871 3184 14929 3242
rect 14963 3184 15021 3242
rect 15055 3184 15113 3242
rect 15147 3184 15205 3242
rect 15239 3184 15297 3242
rect 15331 3184 15389 3242
rect 15423 3184 15481 3242
rect 15515 3184 15573 3242
rect 15607 3184 15665 3242
rect 15699 3184 15757 3242
rect 15791 3184 15849 3242
rect 15883 3184 15941 3242
rect 15975 3184 16033 3242
rect 16067 3184 16125 3242
rect 16159 3184 16217 3242
rect 16251 3184 16309 3242
rect 16343 3184 16401 3242
rect 16435 3184 16493 3242
rect 16527 3184 16585 3242
rect 16619 3184 16677 3242
rect 16711 3184 16769 3242
rect 16803 3184 16861 3242
rect 16895 3184 16953 3242
rect 16987 3184 17045 3242
rect 17079 3184 17137 3242
rect 17171 3184 17229 3242
rect 17263 3184 17321 3242
rect 17355 3184 17413 3242
rect 17447 3184 17505 3242
rect 17539 3184 17597 3242
rect 17631 3184 17689 3242
rect 17723 3184 17781 3242
rect 17815 3184 17873 3242
rect 17907 3184 17965 3242
rect 17999 3184 18057 3242
rect 18091 3184 18149 3242
rect 18183 3184 18241 3242
rect 18275 3184 18333 3242
rect 18367 3184 18425 3242
rect 18459 3184 18517 3242
rect 18551 3184 18609 3242
rect 18643 3184 18701 3242
rect 18735 3184 18793 3242
rect 18827 3184 18885 3242
rect 18919 3184 18977 3242
rect 19011 3184 19069 3242
rect 19103 3184 19161 3242
rect 19195 3184 19253 3242
rect 19287 3184 19345 3242
rect 19379 3184 19437 3242
rect 19471 3184 19529 3242
rect 19563 3184 19621 3242
rect 19655 3184 19713 3242
rect 19747 3184 19805 3242
rect 19839 3184 19897 3242
rect 19931 3184 19989 3242
rect 20023 3184 20081 3242
rect 20115 3184 20173 3242
rect 20207 3184 20265 3242
rect 20299 3184 20357 3242
rect 20391 3184 20449 3242
rect 20483 3184 20541 3242
rect 20575 3184 20633 3242
rect 20667 3184 20725 3242
rect 20759 3184 20817 3242
rect 20851 3184 20909 3242
rect 20943 3184 21001 3242
rect 21035 3184 21093 3242
rect 21127 3184 21185 3242
rect 21219 3184 21277 3242
rect 21311 3184 21369 3242
rect 21403 3184 21461 3242
rect 21495 3184 21553 3242
rect 21587 3184 21645 3242
rect 21679 3184 21737 3242
rect 21771 3184 21829 3242
rect 21863 3184 21921 3242
rect 21955 3184 22013 3242
rect 22047 3184 22105 3242
rect 22139 3184 22197 3242
rect 22231 3184 22289 3242
rect 22323 3184 22381 3242
rect 22415 3184 22473 3242
rect 22507 3184 22565 3242
rect 22599 3184 22657 3242
rect 22691 3184 22749 3242
rect 22783 3184 22841 3242
rect 22875 3184 22933 3242
rect 22967 3184 23025 3242
rect 23059 3184 23117 3242
rect 23151 3184 23209 3242
rect 23243 3184 23301 3242
rect 23335 3184 23393 3242
rect 23427 3184 23456 3242
rect 25594 3224 25745 3258
rect 25814 3472 25825 3506
rect 25968 3490 26002 3540
rect 25780 3284 25825 3472
rect 25780 3250 25791 3284
rect 25594 3216 25646 3224
rect 25594 3182 25612 3216
rect 25780 3216 25825 3250
rect 25859 3456 26002 3490
rect 25859 3262 25893 3456
rect 26043 3454 26067 3488
rect 26101 3462 26143 3488
rect 26101 3454 26109 3462
rect 26043 3428 26109 3454
rect 25927 3352 26009 3422
rect 25927 3348 25948 3352
rect 25982 3318 26009 3352
rect 25961 3314 26009 3318
rect 25927 3298 26009 3314
rect 26043 3412 26143 3428
rect 26043 3288 26087 3412
rect 26177 3378 26211 3547
rect 26259 3572 26335 3624
rect 26553 3582 26619 3624
rect 26259 3538 26275 3572
rect 26309 3538 26335 3572
rect 26395 3556 26429 3572
rect 26395 3504 26429 3522
rect 26553 3548 26569 3582
rect 26603 3548 26619 3582
rect 27042 3582 27118 3624
rect 26553 3514 26619 3548
rect 26828 3547 26844 3581
rect 26878 3547 26994 3581
rect 27042 3548 27058 3582
rect 27092 3548 27118 3582
rect 27306 3582 27583 3624
rect 27166 3556 27200 3572
rect 26245 3488 26515 3504
rect 26245 3462 26395 3488
rect 26279 3454 26395 3462
rect 26429 3454 26515 3488
rect 26553 3480 26569 3514
rect 26603 3480 26619 3514
rect 26790 3488 26837 3494
rect 26279 3428 26295 3454
rect 26245 3412 26295 3428
rect 26397 3378 26447 3394
rect 26177 3344 26413 3378
rect 26177 3336 26257 3344
rect 25859 3224 26002 3262
rect 26077 3254 26087 3288
rect 26043 3238 26087 3254
rect 26123 3266 26139 3300
rect 26173 3284 26189 3300
rect 26123 3250 26155 3266
rect 26123 3226 26189 3250
rect 25594 3166 25646 3182
rect 25680 3156 25696 3190
rect 25730 3156 25746 3190
rect 25814 3182 25825 3216
rect 25968 3208 26002 3224
rect 25780 3166 25825 3182
rect 25680 3114 25746 3156
rect 25864 3156 25884 3190
rect 25918 3156 25934 3190
rect 26223 3190 26257 3336
rect 26403 3328 26447 3344
rect 26481 3310 26515 3454
rect 26790 3462 26803 3488
rect 26824 3428 26837 3454
rect 26549 3420 26750 3428
rect 26549 3386 26711 3420
rect 26745 3386 26750 3420
rect 26790 3412 26837 3428
rect 26885 3462 26926 3478
rect 26885 3428 26892 3462
rect 26549 3380 26750 3386
rect 26549 3378 26615 3380
rect 26549 3344 26565 3378
rect 26599 3344 26615 3378
rect 26885 3358 26926 3428
rect 26802 3352 26926 3358
rect 26677 3310 26693 3344
rect 26727 3310 26743 3344
rect 26295 3276 26311 3310
rect 26345 3290 26361 3310
rect 26345 3284 26377 3290
rect 26295 3250 26343 3276
rect 26481 3276 26743 3310
rect 26802 3318 26803 3352
rect 26837 3322 26926 3352
rect 26960 3378 26994 3547
rect 27306 3548 27322 3582
rect 27356 3548 27533 3582
rect 27567 3548 27583 3582
rect 27166 3514 27200 3522
rect 27617 3545 27674 3590
rect 27028 3480 27583 3514
rect 27028 3462 27078 3480
rect 27062 3428 27078 3462
rect 27028 3412 27078 3428
rect 26960 3362 27230 3378
rect 26960 3344 27196 3362
rect 26837 3318 26859 3322
rect 26802 3288 26859 3318
rect 26481 3250 26525 3276
rect 26295 3244 26377 3250
rect 26459 3216 26475 3250
rect 26509 3216 26525 3250
rect 26802 3254 26825 3288
rect 26559 3224 26593 3240
rect 26802 3238 26859 3254
rect 25968 3158 26002 3174
rect 25864 3114 25934 3156
rect 26058 3156 26074 3190
rect 26108 3156 26257 3190
rect 26058 3150 26257 3156
rect 26291 3186 26325 3202
rect 26291 3114 26325 3152
rect 26359 3172 26375 3206
rect 26409 3182 26425 3206
rect 26960 3190 26994 3344
rect 27186 3328 27196 3344
rect 27186 3312 27230 3328
rect 27069 3284 27088 3310
rect 27069 3250 27079 3284
rect 27122 3276 27144 3310
rect 27113 3250 27144 3276
rect 27264 3253 27300 3480
rect 27069 3244 27144 3250
rect 27234 3250 27300 3253
rect 27234 3216 27250 3250
rect 27284 3216 27300 3250
rect 27334 3420 27436 3446
rect 27334 3386 27355 3420
rect 27389 3412 27436 3420
rect 27470 3412 27486 3446
rect 27334 3378 27389 3386
rect 27368 3344 27389 3378
rect 27549 3362 27583 3480
rect 27651 3511 27674 3545
rect 27617 3477 27674 3511
rect 27651 3443 27674 3477
rect 27617 3423 27674 3443
rect 27334 3282 27389 3344
rect 27440 3350 27515 3362
rect 27440 3316 27463 3350
rect 27499 3316 27515 3350
rect 27549 3346 27599 3362
rect 27549 3312 27565 3346
rect 27549 3296 27599 3312
rect 27334 3248 27472 3282
rect 26559 3182 26593 3190
rect 26409 3172 26593 3182
rect 26359 3148 26593 3172
rect 26647 3156 26663 3190
rect 26697 3156 26713 3190
rect 26647 3114 26713 3156
rect 26841 3156 26857 3190
rect 26891 3156 26994 3190
rect 26841 3150 26994 3156
rect 27030 3186 27082 3202
rect 27030 3152 27048 3186
rect 27030 3114 27082 3152
rect 27134 3172 27150 3206
rect 27184 3182 27200 3206
rect 27334 3198 27368 3214
rect 27184 3172 27334 3182
rect 27134 3164 27334 3172
rect 27134 3148 27368 3164
rect 27425 3200 27472 3248
rect 27425 3166 27438 3200
rect 27425 3150 27472 3166
rect 27517 3190 27583 3258
rect 27633 3240 27674 3423
rect 27517 3156 27533 3190
rect 27567 3156 27583 3190
rect 27517 3114 27583 3156
rect 27617 3224 27674 3240
rect 27651 3190 27674 3224
rect 27617 3148 27674 3190
rect 27708 3564 27771 3580
rect 27708 3530 27721 3564
rect 27755 3530 27771 3564
rect 27708 3496 27771 3530
rect 27708 3462 27721 3496
rect 27755 3462 27771 3496
rect 27708 3362 27771 3462
rect 27807 3570 27866 3624
rect 27807 3536 27816 3570
rect 27850 3536 27866 3570
rect 27807 3502 27866 3536
rect 27807 3468 27816 3502
rect 27850 3468 27866 3502
rect 27807 3450 27866 3468
rect 27900 3548 27952 3590
rect 27900 3546 27909 3548
rect 27943 3514 27952 3548
rect 27934 3512 27952 3514
rect 27900 3478 27952 3512
rect 27934 3444 27952 3478
rect 27986 3574 28038 3590
rect 27986 3540 28004 3574
rect 27986 3506 28038 3540
rect 28072 3558 28138 3624
rect 28072 3524 28088 3558
rect 28122 3524 28138 3558
rect 28172 3574 28217 3590
rect 28206 3540 28217 3574
rect 27986 3472 28004 3506
rect 28172 3506 28217 3540
rect 28256 3558 28326 3624
rect 28256 3524 28276 3558
rect 28310 3524 28326 3558
rect 28360 3574 28394 3590
rect 28437 3547 28453 3581
rect 28487 3547 28603 3581
rect 28038 3488 28137 3490
rect 28038 3472 28091 3488
rect 27986 3456 28091 3472
rect 27900 3386 27952 3444
rect 28125 3454 28137 3488
rect 27708 3346 27875 3362
rect 27708 3312 27841 3346
rect 27708 3296 27875 3312
rect 27708 3216 27771 3296
rect 27909 3262 27952 3386
rect 27986 3379 28057 3422
rect 27986 3361 28013 3379
rect 27986 3327 28001 3361
rect 28047 3345 28057 3379
rect 28035 3327 28057 3345
rect 27986 3292 28057 3327
rect 28091 3361 28137 3454
rect 28091 3327 28103 3361
rect 27708 3182 27721 3216
rect 27755 3182 27771 3216
rect 27900 3226 27952 3262
rect 28091 3258 28137 3327
rect 27708 3148 27771 3182
rect 27807 3190 27866 3206
rect 27807 3156 27816 3190
rect 27850 3156 27866 3190
rect 27807 3114 27866 3156
rect 27934 3192 27952 3226
rect 27900 3148 27952 3192
rect 27986 3224 28137 3258
rect 28206 3472 28217 3506
rect 28360 3490 28394 3540
rect 28172 3284 28217 3472
rect 28172 3250 28183 3284
rect 27986 3216 28038 3224
rect 27986 3182 28004 3216
rect 28172 3216 28217 3250
rect 28251 3456 28394 3490
rect 28251 3262 28285 3456
rect 28435 3454 28459 3488
rect 28493 3462 28535 3488
rect 28493 3454 28501 3462
rect 28435 3428 28501 3454
rect 28319 3351 28401 3422
rect 28319 3348 28346 3351
rect 28380 3317 28401 3351
rect 28353 3314 28401 3317
rect 28319 3298 28401 3314
rect 28435 3412 28535 3428
rect 28435 3288 28479 3412
rect 28569 3378 28603 3547
rect 28651 3572 28727 3624
rect 28945 3582 29011 3624
rect 28651 3538 28667 3572
rect 28701 3538 28727 3572
rect 28787 3556 28821 3572
rect 28787 3504 28821 3522
rect 28945 3548 28961 3582
rect 28995 3548 29011 3582
rect 29434 3582 29510 3624
rect 28945 3514 29011 3548
rect 29220 3547 29236 3581
rect 29270 3547 29386 3581
rect 29434 3548 29450 3582
rect 29484 3548 29510 3582
rect 29698 3582 29975 3624
rect 29558 3556 29592 3572
rect 28637 3488 28907 3504
rect 28637 3462 28787 3488
rect 28671 3454 28787 3462
rect 28821 3454 28907 3488
rect 28945 3480 28961 3514
rect 28995 3480 29011 3514
rect 29182 3488 29229 3494
rect 28671 3428 28687 3454
rect 28637 3412 28687 3428
rect 28789 3378 28839 3394
rect 28569 3344 28805 3378
rect 28569 3336 28649 3344
rect 28251 3224 28394 3262
rect 28469 3254 28479 3288
rect 28435 3238 28479 3254
rect 28515 3266 28531 3300
rect 28565 3284 28581 3300
rect 28515 3250 28547 3266
rect 28515 3226 28581 3250
rect 27986 3166 28038 3182
rect 28072 3156 28088 3190
rect 28122 3156 28138 3190
rect 28206 3182 28217 3216
rect 28360 3208 28394 3224
rect 28172 3166 28217 3182
rect 28072 3114 28138 3156
rect 28256 3156 28276 3190
rect 28310 3156 28326 3190
rect 28615 3190 28649 3336
rect 28795 3328 28839 3344
rect 28873 3310 28907 3454
rect 29182 3462 29195 3488
rect 29216 3428 29229 3454
rect 28941 3420 29142 3428
rect 28941 3386 29103 3420
rect 29137 3386 29142 3420
rect 29182 3412 29229 3428
rect 29277 3462 29318 3478
rect 29277 3428 29284 3462
rect 28941 3380 29142 3386
rect 28941 3378 29007 3380
rect 28941 3344 28957 3378
rect 28991 3344 29007 3378
rect 29277 3358 29318 3428
rect 29194 3352 29318 3358
rect 29069 3310 29085 3344
rect 29119 3310 29135 3344
rect 28687 3276 28703 3310
rect 28737 3290 28753 3310
rect 28737 3284 28769 3290
rect 28687 3250 28735 3276
rect 28873 3276 29135 3310
rect 29194 3318 29195 3352
rect 29229 3322 29318 3352
rect 29352 3378 29386 3547
rect 29698 3548 29714 3582
rect 29748 3548 29925 3582
rect 29959 3548 29975 3582
rect 29558 3514 29592 3522
rect 30009 3545 30066 3590
rect 29420 3480 29975 3514
rect 29420 3462 29470 3480
rect 29454 3428 29470 3462
rect 29420 3412 29470 3428
rect 29352 3362 29622 3378
rect 29352 3344 29588 3362
rect 29229 3318 29251 3322
rect 29194 3288 29251 3318
rect 28873 3250 28917 3276
rect 28687 3244 28769 3250
rect 28851 3216 28867 3250
rect 28901 3216 28917 3250
rect 29194 3254 29217 3288
rect 28951 3224 28985 3240
rect 29194 3238 29251 3254
rect 28360 3158 28394 3174
rect 28256 3114 28326 3156
rect 28450 3156 28466 3190
rect 28500 3156 28649 3190
rect 28450 3150 28649 3156
rect 28683 3186 28717 3202
rect 28683 3114 28717 3152
rect 28751 3172 28767 3206
rect 28801 3182 28817 3206
rect 29352 3190 29386 3344
rect 29578 3328 29588 3344
rect 29578 3312 29622 3328
rect 29461 3284 29480 3310
rect 29461 3250 29471 3284
rect 29514 3276 29536 3310
rect 29505 3250 29536 3276
rect 29656 3253 29692 3480
rect 29461 3244 29536 3250
rect 29626 3250 29692 3253
rect 29626 3216 29642 3250
rect 29676 3216 29692 3250
rect 29726 3420 29828 3446
rect 29726 3386 29747 3420
rect 29781 3412 29828 3420
rect 29862 3412 29878 3446
rect 29726 3378 29781 3386
rect 29760 3344 29781 3378
rect 29941 3362 29975 3480
rect 30043 3511 30066 3545
rect 30009 3477 30066 3511
rect 30043 3443 30066 3477
rect 30009 3423 30066 3443
rect 29726 3282 29781 3344
rect 29832 3351 29907 3362
rect 29832 3317 29856 3351
rect 29890 3350 29907 3351
rect 29832 3316 29857 3317
rect 29891 3316 29907 3350
rect 29941 3346 29991 3362
rect 29941 3312 29957 3346
rect 29941 3296 29991 3312
rect 29726 3248 29864 3282
rect 28951 3182 28985 3190
rect 28801 3172 28985 3182
rect 28751 3148 28985 3172
rect 29039 3156 29055 3190
rect 29089 3156 29105 3190
rect 29039 3114 29105 3156
rect 29233 3156 29249 3190
rect 29283 3156 29386 3190
rect 29233 3150 29386 3156
rect 29422 3186 29474 3202
rect 29422 3152 29440 3186
rect 29422 3114 29474 3152
rect 29526 3172 29542 3206
rect 29576 3182 29592 3206
rect 29726 3198 29760 3214
rect 29576 3172 29726 3182
rect 29526 3164 29726 3172
rect 29526 3148 29760 3164
rect 29817 3200 29864 3248
rect 29817 3166 29830 3200
rect 29817 3150 29864 3166
rect 29909 3190 29975 3258
rect 30025 3240 30066 3423
rect 29909 3156 29925 3190
rect 29959 3156 29975 3190
rect 29909 3114 29975 3156
rect 30009 3224 30066 3240
rect 30043 3190 30066 3224
rect 30009 3148 30066 3190
rect 30100 3564 30163 3580
rect 30100 3530 30113 3564
rect 30147 3530 30163 3564
rect 30100 3496 30163 3530
rect 30100 3462 30113 3496
rect 30147 3462 30163 3496
rect 30100 3362 30163 3462
rect 30199 3570 30258 3624
rect 30199 3536 30208 3570
rect 30242 3536 30258 3570
rect 30199 3502 30258 3536
rect 30199 3468 30208 3502
rect 30242 3468 30258 3502
rect 30199 3450 30258 3468
rect 30292 3546 30344 3590
rect 30326 3512 30344 3546
rect 30292 3478 30344 3512
rect 30326 3444 30344 3478
rect 30292 3386 30344 3444
rect 30100 3346 30267 3362
rect 30100 3312 30233 3346
rect 30100 3296 30267 3312
rect 30100 3216 30163 3296
rect 30301 3262 30344 3386
rect 30100 3182 30113 3216
rect 30147 3182 30163 3216
rect 30292 3226 30344 3262
rect 30326 3219 30344 3226
rect 30100 3148 30163 3182
rect 30199 3190 30258 3206
rect 30199 3156 30208 3190
rect 30242 3156 30258 3190
rect 30199 3114 30258 3156
rect 30292 3185 30299 3192
rect 30333 3185 30344 3219
rect 30292 3148 30344 3185
rect 25577 3080 25606 3114
rect 25640 3080 25698 3114
rect 25732 3080 25790 3114
rect 25824 3080 25882 3114
rect 25916 3080 25974 3114
rect 26008 3080 26066 3114
rect 26100 3080 26158 3114
rect 26192 3080 26250 3114
rect 26284 3080 26342 3114
rect 26376 3080 26434 3114
rect 26468 3080 26526 3114
rect 26560 3080 26618 3114
rect 26652 3080 26710 3114
rect 26744 3080 26802 3114
rect 26836 3080 26894 3114
rect 26928 3080 26986 3114
rect 27020 3080 27078 3114
rect 27112 3080 27170 3114
rect 27204 3080 27262 3114
rect 27296 3080 27354 3114
rect 27388 3080 27446 3114
rect 27480 3080 27538 3114
rect 27572 3080 27630 3114
rect 27664 3080 27722 3114
rect 27756 3080 27814 3114
rect 27848 3080 27906 3114
rect 27940 3080 27998 3114
rect 28032 3080 28090 3114
rect 28124 3080 28182 3114
rect 28216 3080 28274 3114
rect 28308 3080 28366 3114
rect 28400 3080 28458 3114
rect 28492 3080 28550 3114
rect 28584 3080 28642 3114
rect 28676 3080 28734 3114
rect 28768 3080 28826 3114
rect 28860 3080 28918 3114
rect 28952 3080 29010 3114
rect 29044 3080 29102 3114
rect 29136 3080 29194 3114
rect 29228 3080 29286 3114
rect 29320 3080 29378 3114
rect 29412 3080 29470 3114
rect 29504 3080 29562 3114
rect 29596 3080 29654 3114
rect 29688 3080 29746 3114
rect 29780 3080 29838 3114
rect 29872 3080 29930 3114
rect 29964 3080 30022 3114
rect 30056 3080 30114 3114
rect 30148 3080 30206 3114
rect 30240 3080 30298 3114
rect 30332 3080 30361 3114
rect 25577 3067 30361 3080
rect 25577 3033 25606 3067
rect 25640 3033 25698 3067
rect 25732 3033 25790 3067
rect 25824 3033 25882 3067
rect 25916 3033 25974 3067
rect 26008 3033 26066 3067
rect 26100 3033 26158 3067
rect 26192 3033 26250 3067
rect 26284 3033 26342 3067
rect 26376 3033 26434 3067
rect 26468 3033 26526 3067
rect 26560 3033 26618 3067
rect 26652 3033 26710 3067
rect 26744 3033 26802 3067
rect 26836 3033 26894 3067
rect 26928 3033 26986 3067
rect 27020 3033 27078 3067
rect 27112 3033 27171 3067
rect 27205 3033 27262 3067
rect 27296 3033 27354 3067
rect 27388 3033 27446 3067
rect 27480 3033 27539 3067
rect 27573 3033 27630 3067
rect 27664 3033 27722 3067
rect 27756 3033 27814 3067
rect 27848 3033 27906 3067
rect 27940 3033 27998 3067
rect 28032 3033 28090 3067
rect 28124 3033 28182 3067
rect 28216 3033 28274 3067
rect 28308 3033 28366 3067
rect 28400 3033 28458 3067
rect 28492 3033 28550 3067
rect 28584 3033 28642 3067
rect 28676 3033 28733 3067
rect 28767 3033 28825 3067
rect 28859 3033 28918 3067
rect 28952 3033 29010 3067
rect 29044 3033 29102 3067
rect 29136 3033 29193 3067
rect 29227 3033 29286 3067
rect 29320 3033 29377 3067
rect 29411 3033 29470 3067
rect 29504 3033 29562 3067
rect 29596 3033 29654 3067
rect 29688 3033 29746 3067
rect 29780 3033 29838 3067
rect 29872 3033 29930 3067
rect 29964 3033 30022 3067
rect 30056 3033 30114 3067
rect 30148 3033 30206 3067
rect 30240 3033 30298 3067
rect 30332 3033 30361 3067
rect 25577 3018 30361 3033
rect 25577 2984 25606 3018
rect 25640 2984 25698 3018
rect 25732 2984 25790 3018
rect 25824 2984 25882 3018
rect 25916 2984 25974 3018
rect 26008 2984 26066 3018
rect 26100 2984 26158 3018
rect 26192 2984 26250 3018
rect 26284 2984 26342 3018
rect 26376 2984 26434 3018
rect 26468 2984 26526 3018
rect 26560 2984 26618 3018
rect 26652 2984 26710 3018
rect 26744 2984 26802 3018
rect 26836 2984 26894 3018
rect 26928 2984 26986 3018
rect 27020 2984 27078 3018
rect 27112 2984 27170 3018
rect 27204 2984 27262 3018
rect 27296 2984 27354 3018
rect 27388 2984 27446 3018
rect 27480 2984 27538 3018
rect 27572 2984 27630 3018
rect 27664 2984 27722 3018
rect 27756 2984 27814 3018
rect 27848 2984 27906 3018
rect 27940 2984 27998 3018
rect 28032 2984 28090 3018
rect 28124 2984 28182 3018
rect 28216 2984 28274 3018
rect 28308 2984 28366 3018
rect 28400 2984 28458 3018
rect 28492 2984 28550 3018
rect 28584 2984 28642 3018
rect 28676 2984 28734 3018
rect 28768 2984 28826 3018
rect 28860 2984 28918 3018
rect 28952 2984 29010 3018
rect 29044 2984 29102 3018
rect 29136 2984 29194 3018
rect 29228 2984 29286 3018
rect 29320 2984 29378 3018
rect 29412 2984 29470 3018
rect 29504 2984 29562 3018
rect 29596 2984 29654 3018
rect 29688 2984 29746 3018
rect 29780 2984 29838 3018
rect 29872 2984 29930 3018
rect 29964 2984 30022 3018
rect 30056 2984 30114 3018
rect 30148 2984 30206 3018
rect 30240 2984 30298 3018
rect 30332 2984 30361 3018
rect 25680 2942 25746 2984
rect 25594 2916 25646 2932
rect 25594 2882 25612 2916
rect 25680 2908 25696 2942
rect 25730 2908 25746 2942
rect 25864 2942 25934 2984
rect 25780 2916 25825 2932
rect 25594 2874 25646 2882
rect 25814 2882 25825 2916
rect 25864 2908 25884 2942
rect 25918 2908 25934 2942
rect 26058 2942 26257 2948
rect 25968 2924 26002 2940
rect 25594 2840 25745 2874
rect 25594 2772 25626 2806
rect 25660 2772 25665 2806
rect 25594 2771 25665 2772
rect 25594 2737 25609 2771
rect 25643 2737 25665 2771
rect 25594 2676 25665 2737
rect 25699 2771 25745 2840
rect 25699 2737 25711 2771
rect 25699 2644 25745 2737
rect 25594 2626 25699 2642
rect 25594 2592 25612 2626
rect 25646 2610 25699 2626
rect 25733 2610 25745 2644
rect 25646 2608 25745 2610
rect 25780 2848 25825 2882
rect 26058 2908 26074 2942
rect 26108 2908 26257 2942
rect 25968 2874 26002 2890
rect 25780 2814 25791 2848
rect 25780 2626 25825 2814
rect 25594 2558 25646 2592
rect 25814 2592 25825 2626
rect 25859 2836 26002 2874
rect 26043 2844 26087 2860
rect 25859 2642 25893 2836
rect 26077 2810 26087 2844
rect 25927 2784 26009 2800
rect 25961 2750 26009 2784
rect 25927 2722 26009 2750
rect 25927 2688 25953 2722
rect 25987 2688 26009 2722
rect 25927 2676 26009 2688
rect 26043 2686 26087 2810
rect 26123 2848 26189 2872
rect 26123 2832 26155 2848
rect 26123 2798 26139 2832
rect 26173 2798 26189 2814
rect 26223 2762 26257 2908
rect 26291 2946 26325 2984
rect 26291 2896 26325 2912
rect 26359 2926 26593 2950
rect 26359 2892 26375 2926
rect 26409 2916 26593 2926
rect 26409 2892 26425 2916
rect 26559 2908 26593 2916
rect 26647 2942 26713 2984
rect 26647 2908 26663 2942
rect 26697 2908 26713 2942
rect 26841 2942 26994 2948
rect 26841 2908 26857 2942
rect 26891 2908 26994 2942
rect 26295 2848 26377 2854
rect 26459 2848 26475 2882
rect 26509 2848 26525 2882
rect 26559 2858 26593 2874
rect 26295 2822 26343 2848
rect 26295 2788 26311 2822
rect 26345 2808 26377 2814
rect 26481 2822 26525 2848
rect 26802 2844 26859 2860
rect 26345 2788 26361 2808
rect 26481 2788 26743 2822
rect 26177 2754 26257 2762
rect 26403 2754 26447 2770
rect 26177 2720 26413 2754
rect 26043 2670 26143 2686
rect 26043 2644 26109 2670
rect 25859 2608 26002 2642
rect 26043 2610 26067 2644
rect 26101 2636 26109 2644
rect 26101 2610 26143 2636
rect 25594 2524 25612 2558
rect 25594 2508 25646 2524
rect 25680 2540 25696 2574
rect 25730 2540 25746 2574
rect 25680 2474 25746 2540
rect 25780 2558 25825 2592
rect 25814 2524 25825 2558
rect 25780 2508 25825 2524
rect 25864 2540 25884 2574
rect 25918 2540 25934 2574
rect 25864 2474 25934 2540
rect 25968 2558 26002 2608
rect 26177 2551 26211 2720
rect 26397 2704 26447 2720
rect 26245 2670 26295 2686
rect 26279 2644 26295 2670
rect 26481 2644 26515 2788
rect 26677 2754 26693 2788
rect 26727 2754 26743 2788
rect 26802 2810 26825 2844
rect 26802 2780 26859 2810
rect 26549 2720 26565 2754
rect 26599 2720 26615 2754
rect 26802 2746 26803 2780
rect 26837 2776 26859 2780
rect 26837 2746 26926 2776
rect 26802 2740 26926 2746
rect 26549 2718 26615 2720
rect 26549 2712 26750 2718
rect 26549 2678 26711 2712
rect 26745 2678 26750 2712
rect 26549 2670 26750 2678
rect 26790 2670 26837 2686
rect 26279 2636 26395 2644
rect 26245 2610 26395 2636
rect 26429 2610 26515 2644
rect 26824 2644 26837 2670
rect 26245 2594 26515 2610
rect 26395 2576 26429 2594
rect 25968 2508 26002 2524
rect 26045 2517 26061 2551
rect 26095 2517 26211 2551
rect 26259 2526 26275 2560
rect 26309 2526 26335 2560
rect 26395 2526 26429 2542
rect 26553 2584 26569 2618
rect 26603 2584 26619 2618
rect 26790 2610 26803 2636
rect 26885 2670 26926 2740
rect 26885 2636 26892 2670
rect 26885 2620 26926 2636
rect 26960 2754 26994 2908
rect 27030 2946 27082 2984
rect 27030 2912 27048 2946
rect 27030 2896 27082 2912
rect 27134 2934 27368 2950
rect 27134 2926 27334 2934
rect 27134 2892 27150 2926
rect 27184 2916 27334 2926
rect 27184 2892 27200 2916
rect 27334 2884 27368 2900
rect 27425 2932 27472 2948
rect 27425 2898 27438 2932
rect 27069 2848 27144 2854
rect 27069 2814 27079 2848
rect 27113 2822 27144 2848
rect 27234 2848 27250 2882
rect 27284 2848 27300 2882
rect 27425 2850 27472 2898
rect 27234 2845 27300 2848
rect 27069 2788 27088 2814
rect 27122 2788 27144 2822
rect 27186 2770 27230 2786
rect 27186 2754 27196 2770
rect 26960 2736 27196 2754
rect 26960 2720 27230 2736
rect 26790 2604 26837 2610
rect 26553 2550 26619 2584
rect 26960 2551 26994 2720
rect 27028 2670 27078 2686
rect 27062 2636 27078 2670
rect 27028 2618 27078 2636
rect 27264 2618 27300 2845
rect 27334 2816 27472 2850
rect 27517 2942 27583 2984
rect 27517 2908 27533 2942
rect 27567 2908 27583 2942
rect 27517 2840 27583 2908
rect 27617 2908 27674 2950
rect 27651 2874 27674 2908
rect 27617 2858 27674 2874
rect 27334 2754 27389 2816
rect 27549 2786 27599 2802
rect 27368 2720 27389 2754
rect 27440 2748 27465 2782
rect 27499 2780 27515 2782
rect 27440 2746 27472 2748
rect 27506 2746 27515 2780
rect 27440 2736 27515 2746
rect 27549 2752 27565 2786
rect 27549 2736 27599 2752
rect 27334 2712 27389 2720
rect 27334 2678 27355 2712
rect 27389 2678 27436 2686
rect 27334 2652 27436 2678
rect 27470 2652 27486 2686
rect 27549 2618 27583 2736
rect 27633 2675 27674 2858
rect 27028 2584 27583 2618
rect 27617 2655 27674 2675
rect 27651 2621 27674 2655
rect 27617 2587 27674 2621
rect 26259 2474 26335 2526
rect 26553 2516 26569 2550
rect 26603 2516 26619 2550
rect 26828 2517 26844 2551
rect 26878 2517 26994 2551
rect 27166 2576 27200 2584
rect 26553 2474 26619 2516
rect 27042 2516 27058 2550
rect 27092 2516 27118 2550
rect 27651 2553 27674 2587
rect 27166 2526 27200 2542
rect 27042 2474 27118 2516
rect 27306 2516 27322 2550
rect 27356 2516 27533 2550
rect 27567 2516 27583 2550
rect 27306 2474 27583 2516
rect 27617 2508 27674 2553
rect 27708 2916 27771 2950
rect 27708 2882 27721 2916
rect 27755 2882 27771 2916
rect 27807 2942 27866 2984
rect 27807 2908 27816 2942
rect 27850 2908 27866 2942
rect 27807 2892 27866 2908
rect 27900 2906 27952 2950
rect 28072 2942 28138 2984
rect 27708 2802 27771 2882
rect 27934 2872 27952 2906
rect 27900 2836 27952 2872
rect 27986 2916 28038 2932
rect 27986 2882 28004 2916
rect 28072 2908 28088 2942
rect 28122 2908 28138 2942
rect 28256 2942 28326 2984
rect 28172 2916 28217 2932
rect 27986 2874 28038 2882
rect 28206 2882 28217 2916
rect 28256 2908 28276 2942
rect 28310 2908 28326 2942
rect 28450 2942 28649 2948
rect 28360 2924 28394 2940
rect 27986 2840 28137 2874
rect 27708 2786 27875 2802
rect 27708 2752 27841 2786
rect 27708 2736 27875 2752
rect 27708 2636 27771 2736
rect 27909 2712 27952 2836
rect 27900 2654 27952 2712
rect 27986 2771 28057 2806
rect 27986 2737 28001 2771
rect 28035 2762 28057 2771
rect 27986 2728 28010 2737
rect 28044 2728 28057 2762
rect 27986 2676 28057 2728
rect 28091 2771 28137 2840
rect 28091 2737 28103 2771
rect 27708 2602 27721 2636
rect 27755 2602 27771 2636
rect 27708 2568 27771 2602
rect 27708 2534 27721 2568
rect 27755 2534 27771 2568
rect 27708 2518 27771 2534
rect 27807 2630 27866 2648
rect 27807 2596 27816 2630
rect 27850 2596 27866 2630
rect 27807 2562 27866 2596
rect 27807 2528 27816 2562
rect 27850 2528 27866 2562
rect 27807 2474 27866 2528
rect 27934 2620 27952 2654
rect 28091 2644 28137 2737
rect 27900 2586 27952 2620
rect 27934 2585 27952 2586
rect 27900 2551 27906 2552
rect 27940 2551 27952 2585
rect 27900 2508 27952 2551
rect 27986 2626 28091 2642
rect 27986 2592 28004 2626
rect 28038 2610 28091 2626
rect 28125 2610 28137 2644
rect 28038 2608 28137 2610
rect 28172 2848 28217 2882
rect 28450 2908 28466 2942
rect 28500 2908 28649 2942
rect 28360 2874 28394 2890
rect 28172 2814 28183 2848
rect 28172 2626 28217 2814
rect 27986 2558 28038 2592
rect 28206 2592 28217 2626
rect 28251 2836 28394 2874
rect 28435 2844 28479 2860
rect 28251 2642 28285 2836
rect 28469 2810 28479 2844
rect 28319 2784 28401 2800
rect 28353 2779 28401 2784
rect 28319 2745 28347 2750
rect 28381 2745 28401 2779
rect 28319 2676 28401 2745
rect 28435 2686 28479 2810
rect 28515 2848 28581 2872
rect 28515 2832 28547 2848
rect 28515 2798 28531 2832
rect 28565 2798 28581 2814
rect 28615 2762 28649 2908
rect 28683 2946 28717 2984
rect 28683 2896 28717 2912
rect 28751 2926 28985 2950
rect 28751 2892 28767 2926
rect 28801 2916 28985 2926
rect 28801 2892 28817 2916
rect 28951 2908 28985 2916
rect 29039 2942 29105 2984
rect 29039 2908 29055 2942
rect 29089 2908 29105 2942
rect 29233 2942 29386 2948
rect 29233 2908 29249 2942
rect 29283 2908 29386 2942
rect 28687 2848 28769 2854
rect 28851 2848 28867 2882
rect 28901 2848 28917 2882
rect 28951 2858 28985 2874
rect 28687 2822 28735 2848
rect 28687 2788 28703 2822
rect 28737 2808 28769 2814
rect 28873 2822 28917 2848
rect 29194 2844 29251 2860
rect 28737 2788 28753 2808
rect 28873 2788 29135 2822
rect 28569 2754 28649 2762
rect 28795 2754 28839 2770
rect 28569 2720 28805 2754
rect 28435 2670 28535 2686
rect 28435 2644 28501 2670
rect 28251 2608 28394 2642
rect 28435 2610 28459 2644
rect 28493 2636 28501 2644
rect 28493 2610 28535 2636
rect 27986 2524 28004 2558
rect 27986 2508 28038 2524
rect 28072 2540 28088 2574
rect 28122 2540 28138 2574
rect 28072 2474 28138 2540
rect 28172 2558 28217 2592
rect 28206 2524 28217 2558
rect 28172 2508 28217 2524
rect 28256 2540 28276 2574
rect 28310 2540 28326 2574
rect 28256 2474 28326 2540
rect 28360 2558 28394 2608
rect 28569 2551 28603 2720
rect 28789 2704 28839 2720
rect 28637 2670 28687 2686
rect 28671 2644 28687 2670
rect 28873 2644 28907 2788
rect 29069 2754 29085 2788
rect 29119 2754 29135 2788
rect 29194 2810 29217 2844
rect 29194 2780 29251 2810
rect 28941 2720 28957 2754
rect 28991 2720 29007 2754
rect 29194 2746 29195 2780
rect 29229 2776 29251 2780
rect 29229 2746 29318 2776
rect 29194 2740 29318 2746
rect 28941 2718 29007 2720
rect 28941 2712 29142 2718
rect 28941 2678 29103 2712
rect 29137 2678 29142 2712
rect 28941 2670 29142 2678
rect 29182 2670 29229 2686
rect 28671 2636 28787 2644
rect 28637 2610 28787 2636
rect 28821 2610 28907 2644
rect 29216 2644 29229 2670
rect 28637 2594 28907 2610
rect 28787 2576 28821 2594
rect 28360 2508 28394 2524
rect 28437 2517 28453 2551
rect 28487 2517 28603 2551
rect 28651 2526 28667 2560
rect 28701 2526 28727 2560
rect 28787 2526 28821 2542
rect 28945 2584 28961 2618
rect 28995 2584 29011 2618
rect 29182 2610 29195 2636
rect 29277 2670 29318 2740
rect 29277 2636 29284 2670
rect 29277 2620 29318 2636
rect 29352 2754 29386 2908
rect 29422 2946 29474 2984
rect 29422 2912 29440 2946
rect 29422 2896 29474 2912
rect 29526 2934 29760 2950
rect 29526 2926 29726 2934
rect 29526 2892 29542 2926
rect 29576 2916 29726 2926
rect 29576 2892 29592 2916
rect 29726 2884 29760 2900
rect 29817 2932 29864 2948
rect 29817 2898 29830 2932
rect 29461 2848 29536 2854
rect 29461 2814 29471 2848
rect 29505 2822 29536 2848
rect 29626 2848 29642 2882
rect 29676 2848 29692 2882
rect 29817 2850 29864 2898
rect 29626 2845 29692 2848
rect 29461 2788 29480 2814
rect 29514 2788 29536 2822
rect 29578 2770 29622 2786
rect 29578 2754 29588 2770
rect 29352 2736 29588 2754
rect 29352 2720 29622 2736
rect 29182 2604 29229 2610
rect 28945 2550 29011 2584
rect 29352 2551 29386 2720
rect 29420 2670 29470 2686
rect 29454 2636 29470 2670
rect 29420 2618 29470 2636
rect 29656 2618 29692 2845
rect 29726 2816 29864 2850
rect 29909 2942 29975 2984
rect 29909 2908 29925 2942
rect 29959 2908 29975 2942
rect 29909 2840 29975 2908
rect 30009 2908 30066 2950
rect 30043 2874 30066 2908
rect 30009 2858 30066 2874
rect 29726 2754 29781 2816
rect 29941 2786 29991 2802
rect 29760 2720 29781 2754
rect 29832 2748 29856 2782
rect 29891 2748 29907 2782
rect 29832 2736 29907 2748
rect 29941 2752 29957 2786
rect 29941 2736 29991 2752
rect 29726 2712 29781 2720
rect 29726 2678 29747 2712
rect 29781 2678 29828 2686
rect 29726 2652 29828 2678
rect 29862 2652 29878 2686
rect 29941 2618 29975 2736
rect 30025 2675 30066 2858
rect 29420 2584 29975 2618
rect 30009 2655 30066 2675
rect 30043 2621 30066 2655
rect 30009 2587 30066 2621
rect 28651 2474 28727 2526
rect 28945 2516 28961 2550
rect 28995 2516 29011 2550
rect 29220 2517 29236 2551
rect 29270 2517 29386 2551
rect 29558 2576 29592 2584
rect 28945 2474 29011 2516
rect 29434 2516 29450 2550
rect 29484 2516 29510 2550
rect 30043 2553 30066 2587
rect 29558 2526 29592 2542
rect 29434 2474 29510 2516
rect 29698 2516 29714 2550
rect 29748 2516 29925 2550
rect 29959 2516 29975 2550
rect 29698 2474 29975 2516
rect 30009 2508 30066 2553
rect 30100 2916 30163 2950
rect 30100 2882 30113 2916
rect 30147 2882 30163 2916
rect 30199 2942 30258 2984
rect 30199 2908 30208 2942
rect 30242 2908 30258 2942
rect 30199 2892 30258 2908
rect 30292 2906 30344 2950
rect 30326 2896 30344 2906
rect 30100 2802 30163 2882
rect 30292 2862 30293 2872
rect 30327 2862 30344 2896
rect 30292 2836 30344 2862
rect 30100 2786 30267 2802
rect 30100 2752 30233 2786
rect 30100 2736 30267 2752
rect 30100 2636 30163 2736
rect 30301 2712 30344 2836
rect 30292 2654 30344 2712
rect 30100 2602 30113 2636
rect 30147 2602 30163 2636
rect 30100 2568 30163 2602
rect 30100 2534 30113 2568
rect 30147 2534 30163 2568
rect 30100 2518 30163 2534
rect 30199 2630 30258 2648
rect 30199 2596 30208 2630
rect 30242 2596 30258 2630
rect 30199 2562 30258 2596
rect 30199 2528 30208 2562
rect 30242 2528 30258 2562
rect 30199 2474 30258 2528
rect 30326 2620 30344 2654
rect 30292 2586 30344 2620
rect 30326 2552 30344 2586
rect 30292 2508 30344 2552
rect 25577 2440 25606 2474
rect 25640 2440 25698 2474
rect 25732 2440 25790 2474
rect 25824 2440 25882 2474
rect 25916 2440 25974 2474
rect 26008 2440 26066 2474
rect 26100 2440 26158 2474
rect 26192 2440 26250 2474
rect 26284 2440 26342 2474
rect 26376 2440 26434 2474
rect 26468 2440 26526 2474
rect 26560 2440 26618 2474
rect 26652 2440 26710 2474
rect 26744 2440 26802 2474
rect 26836 2440 26894 2474
rect 26928 2440 26986 2474
rect 27020 2440 27078 2474
rect 27112 2440 27170 2474
rect 27204 2440 27262 2474
rect 27296 2440 27354 2474
rect 27388 2440 27446 2474
rect 27480 2440 27538 2474
rect 27572 2440 27630 2474
rect 27664 2440 27722 2474
rect 27756 2440 27814 2474
rect 27848 2440 27906 2474
rect 27940 2440 27998 2474
rect 28032 2440 28090 2474
rect 28124 2440 28182 2474
rect 28216 2440 28274 2474
rect 28308 2440 28366 2474
rect 28400 2440 28458 2474
rect 28492 2440 28550 2474
rect 28584 2440 28642 2474
rect 28676 2440 28734 2474
rect 28768 2440 28826 2474
rect 28860 2440 28918 2474
rect 28952 2440 29010 2474
rect 29044 2440 29102 2474
rect 29136 2440 29194 2474
rect 29228 2440 29286 2474
rect 29320 2440 29378 2474
rect 29412 2440 29470 2474
rect 29504 2440 29562 2474
rect 29596 2440 29654 2474
rect 29688 2440 29746 2474
rect 29780 2440 29838 2474
rect 29872 2440 29930 2474
rect 29964 2440 30022 2474
rect 30056 2440 30114 2474
rect 30148 2440 30206 2474
rect 30240 2440 30298 2474
rect 30332 2440 30361 2474
rect 25577 2425 30361 2440
rect 25577 2391 25609 2425
rect 25643 2391 25699 2425
rect 25733 2391 25792 2425
rect 25826 2391 25882 2425
rect 25916 2391 25973 2425
rect 26007 2391 26067 2425
rect 26101 2391 26158 2425
rect 26192 2391 26250 2425
rect 26284 2391 26342 2425
rect 26376 2391 26435 2425
rect 26469 2391 26526 2425
rect 26560 2391 26618 2425
rect 26652 2391 26710 2425
rect 26744 2391 26802 2425
rect 26836 2391 26895 2425
rect 26929 2391 26986 2425
rect 27020 2391 27077 2425
rect 27111 2391 27170 2425
rect 27204 2391 27263 2425
rect 27297 2391 27354 2425
rect 27388 2391 27446 2425
rect 27480 2391 27538 2425
rect 27572 2391 27630 2425
rect 27664 2391 27723 2425
rect 27757 2391 27813 2425
rect 27847 2391 27906 2425
rect 27940 2391 27998 2425
rect 28032 2391 28091 2425
rect 28125 2391 28185 2425
rect 28219 2391 28274 2425
rect 28308 2391 28366 2425
rect 28400 2391 28458 2425
rect 28492 2391 28550 2425
rect 28584 2391 28642 2425
rect 28676 2391 28734 2425
rect 28768 2391 28826 2425
rect 28860 2391 28918 2425
rect 28952 2391 29010 2425
rect 29044 2391 29102 2425
rect 29136 2391 29194 2425
rect 29228 2391 29286 2425
rect 29320 2391 29378 2425
rect 29412 2391 29470 2425
rect 29504 2391 29562 2425
rect 29596 2391 29654 2425
rect 29688 2391 29746 2425
rect 29780 2391 29838 2425
rect 29872 2391 29930 2425
rect 29964 2391 30022 2425
rect 30056 2391 30114 2425
rect 30148 2391 30207 2425
rect 30241 2391 30298 2425
rect 30332 2391 30361 2425
rect 25577 2378 30361 2391
rect 25577 2344 25606 2378
rect 25640 2344 25698 2378
rect 25732 2344 25790 2378
rect 25824 2344 25882 2378
rect 25916 2344 25974 2378
rect 26008 2344 26066 2378
rect 26100 2344 26158 2378
rect 26192 2344 26250 2378
rect 26284 2344 26342 2378
rect 26376 2344 26434 2378
rect 26468 2344 26526 2378
rect 26560 2344 26618 2378
rect 26652 2344 26710 2378
rect 26744 2344 26802 2378
rect 26836 2344 26894 2378
rect 26928 2344 26986 2378
rect 27020 2344 27078 2378
rect 27112 2344 27170 2378
rect 27204 2344 27262 2378
rect 27296 2344 27354 2378
rect 27388 2344 27446 2378
rect 27480 2344 27538 2378
rect 27572 2344 27630 2378
rect 27664 2344 27722 2378
rect 27756 2344 27814 2378
rect 27848 2344 27906 2378
rect 27940 2344 27998 2378
rect 28032 2344 28090 2378
rect 28124 2344 28182 2378
rect 28216 2344 28274 2378
rect 28308 2344 28366 2378
rect 28400 2344 28458 2378
rect 28492 2344 28550 2378
rect 28584 2344 28642 2378
rect 28676 2344 28734 2378
rect 28768 2344 28826 2378
rect 28860 2344 28918 2378
rect 28952 2344 29010 2378
rect 29044 2344 29102 2378
rect 29136 2344 29194 2378
rect 29228 2344 29286 2378
rect 29320 2344 29378 2378
rect 29412 2344 29470 2378
rect 29504 2344 29562 2378
rect 29596 2344 29654 2378
rect 29688 2344 29746 2378
rect 29780 2344 29838 2378
rect 29872 2344 29930 2378
rect 29964 2344 30022 2378
rect 30056 2344 30114 2378
rect 30148 2344 30206 2378
rect 30240 2344 30298 2378
rect 30332 2344 30361 2378
rect 25594 2294 25646 2310
rect 25594 2260 25612 2294
rect 25594 2226 25646 2260
rect 25680 2278 25746 2344
rect 25680 2244 25696 2278
rect 25730 2244 25746 2278
rect 25780 2294 25825 2310
rect 25814 2260 25825 2294
rect 25594 2192 25612 2226
rect 25780 2226 25825 2260
rect 25864 2278 25934 2344
rect 25864 2244 25884 2278
rect 25918 2244 25934 2278
rect 25968 2294 26002 2310
rect 26045 2267 26061 2301
rect 26095 2267 26211 2301
rect 25646 2208 25745 2210
rect 25646 2192 25699 2208
rect 25594 2176 25699 2192
rect 25733 2174 25745 2208
rect 25594 2081 25665 2142
rect 25594 2047 25609 2081
rect 25643 2047 25665 2081
rect 25594 2046 25665 2047
rect 25594 2012 25622 2046
rect 25656 2012 25665 2046
rect 25699 2081 25745 2174
rect 25699 2047 25711 2081
rect 25699 1978 25745 2047
rect 25594 1944 25745 1978
rect 25814 2192 25825 2226
rect 25968 2210 26002 2260
rect 25780 2004 25825 2192
rect 25780 1970 25791 2004
rect 25594 1936 25646 1944
rect 25594 1902 25612 1936
rect 25780 1936 25825 1970
rect 25859 2176 26002 2210
rect 25859 1982 25893 2176
rect 26043 2174 26067 2208
rect 26101 2182 26143 2208
rect 26101 2174 26109 2182
rect 26043 2148 26109 2174
rect 25927 2130 26009 2142
rect 25927 2096 25950 2130
rect 25984 2096 26009 2130
rect 25927 2068 26009 2096
rect 25961 2034 26009 2068
rect 25927 2018 26009 2034
rect 26043 2132 26143 2148
rect 26043 2008 26087 2132
rect 26177 2098 26211 2267
rect 26259 2292 26335 2344
rect 26553 2302 26619 2344
rect 26259 2258 26275 2292
rect 26309 2258 26335 2292
rect 26395 2276 26429 2292
rect 26395 2224 26429 2242
rect 26553 2268 26569 2302
rect 26603 2268 26619 2302
rect 27042 2302 27118 2344
rect 26553 2234 26619 2268
rect 26828 2267 26844 2301
rect 26878 2267 26994 2301
rect 27042 2268 27058 2302
rect 27092 2268 27118 2302
rect 27306 2302 27583 2344
rect 27166 2276 27200 2292
rect 26245 2208 26515 2224
rect 26245 2182 26395 2208
rect 26279 2174 26395 2182
rect 26429 2174 26515 2208
rect 26553 2200 26569 2234
rect 26603 2200 26619 2234
rect 26790 2208 26837 2214
rect 26279 2148 26295 2174
rect 26245 2132 26295 2148
rect 26397 2098 26447 2114
rect 26177 2064 26413 2098
rect 26177 2056 26257 2064
rect 25859 1944 26002 1982
rect 26077 1974 26087 2008
rect 26043 1958 26087 1974
rect 26123 1986 26139 2020
rect 26173 2004 26189 2020
rect 26123 1970 26155 1986
rect 26123 1946 26189 1970
rect 25594 1886 25646 1902
rect 25680 1876 25696 1910
rect 25730 1876 25746 1910
rect 25814 1902 25825 1936
rect 25968 1928 26002 1944
rect 25780 1886 25825 1902
rect 25680 1834 25746 1876
rect 25864 1876 25884 1910
rect 25918 1876 25934 1910
rect 26223 1910 26257 2056
rect 26403 2048 26447 2064
rect 26481 2030 26515 2174
rect 26790 2182 26803 2208
rect 26824 2148 26837 2174
rect 26549 2140 26750 2148
rect 26549 2106 26711 2140
rect 26745 2106 26750 2140
rect 26790 2132 26837 2148
rect 26885 2182 26926 2198
rect 26885 2148 26892 2182
rect 26549 2100 26750 2106
rect 26549 2098 26615 2100
rect 26549 2064 26565 2098
rect 26599 2064 26615 2098
rect 26885 2078 26926 2148
rect 26802 2072 26926 2078
rect 26677 2030 26693 2064
rect 26727 2030 26743 2064
rect 26295 1996 26311 2030
rect 26345 2010 26361 2030
rect 26345 2004 26377 2010
rect 26295 1970 26343 1996
rect 26481 1996 26743 2030
rect 26802 2038 26803 2072
rect 26837 2042 26926 2072
rect 26960 2098 26994 2267
rect 27306 2268 27322 2302
rect 27356 2268 27533 2302
rect 27567 2268 27583 2302
rect 27166 2234 27200 2242
rect 27617 2265 27674 2310
rect 27028 2200 27583 2234
rect 27028 2182 27078 2200
rect 27062 2148 27078 2182
rect 27028 2132 27078 2148
rect 26960 2082 27230 2098
rect 26960 2064 27196 2082
rect 26837 2038 26859 2042
rect 26802 2008 26859 2038
rect 26481 1970 26525 1996
rect 26295 1964 26377 1970
rect 26459 1936 26475 1970
rect 26509 1936 26525 1970
rect 26802 1974 26825 2008
rect 26559 1944 26593 1960
rect 26802 1958 26859 1974
rect 25968 1878 26002 1894
rect 25864 1834 25934 1876
rect 26058 1876 26074 1910
rect 26108 1876 26257 1910
rect 26058 1870 26257 1876
rect 26291 1906 26325 1922
rect 26291 1834 26325 1872
rect 26359 1892 26375 1926
rect 26409 1902 26425 1926
rect 26960 1910 26994 2064
rect 27186 2048 27196 2064
rect 27186 2032 27230 2048
rect 27069 2004 27088 2030
rect 27069 1970 27079 2004
rect 27122 1996 27144 2030
rect 27113 1970 27144 1996
rect 27264 1973 27300 2200
rect 27069 1964 27144 1970
rect 27234 1970 27300 1973
rect 27234 1936 27250 1970
rect 27284 1936 27300 1970
rect 27334 2140 27436 2166
rect 27334 2106 27355 2140
rect 27389 2132 27436 2140
rect 27470 2132 27486 2166
rect 27334 2098 27389 2106
rect 27368 2064 27389 2098
rect 27549 2082 27583 2200
rect 27651 2231 27674 2265
rect 27617 2197 27674 2231
rect 27651 2163 27674 2197
rect 27617 2143 27674 2163
rect 27334 2002 27389 2064
rect 27440 2070 27515 2082
rect 27440 2036 27464 2070
rect 27499 2036 27515 2070
rect 27549 2066 27599 2082
rect 27549 2032 27565 2066
rect 27549 2016 27599 2032
rect 27334 1968 27472 2002
rect 26559 1902 26593 1910
rect 26409 1892 26593 1902
rect 26359 1868 26593 1892
rect 26647 1876 26663 1910
rect 26697 1876 26713 1910
rect 26647 1834 26713 1876
rect 26841 1876 26857 1910
rect 26891 1876 26994 1910
rect 26841 1870 26994 1876
rect 27030 1906 27082 1922
rect 27030 1872 27048 1906
rect 27030 1834 27082 1872
rect 27134 1892 27150 1926
rect 27184 1902 27200 1926
rect 27334 1918 27368 1934
rect 27184 1892 27334 1902
rect 27134 1884 27334 1892
rect 27134 1868 27368 1884
rect 27425 1920 27472 1968
rect 27425 1886 27438 1920
rect 27425 1870 27472 1886
rect 27517 1910 27583 1978
rect 27633 1960 27674 2143
rect 27517 1876 27533 1910
rect 27567 1876 27583 1910
rect 27517 1834 27583 1876
rect 27617 1944 27674 1960
rect 27651 1910 27674 1944
rect 27617 1868 27674 1910
rect 27708 2284 27771 2300
rect 27708 2250 27721 2284
rect 27755 2250 27771 2284
rect 27708 2216 27771 2250
rect 27708 2182 27721 2216
rect 27755 2182 27771 2216
rect 27708 2082 27771 2182
rect 27807 2290 27866 2344
rect 27807 2256 27816 2290
rect 27850 2256 27866 2290
rect 27807 2222 27866 2256
rect 27807 2188 27816 2222
rect 27850 2188 27866 2222
rect 27807 2170 27866 2188
rect 27900 2270 27952 2310
rect 27900 2266 27906 2270
rect 27940 2236 27952 2270
rect 27934 2232 27952 2236
rect 27900 2198 27952 2232
rect 27934 2164 27952 2198
rect 27986 2294 28038 2310
rect 27986 2260 28004 2294
rect 27986 2226 28038 2260
rect 28072 2278 28138 2344
rect 28072 2244 28088 2278
rect 28122 2244 28138 2278
rect 28172 2294 28217 2310
rect 28206 2260 28217 2294
rect 27986 2192 28004 2226
rect 28172 2226 28217 2260
rect 28256 2278 28326 2344
rect 28256 2244 28276 2278
rect 28310 2244 28326 2278
rect 28360 2294 28394 2310
rect 28437 2267 28453 2301
rect 28487 2267 28603 2301
rect 28038 2208 28137 2210
rect 28038 2192 28091 2208
rect 27986 2176 28091 2192
rect 27900 2106 27952 2164
rect 28125 2174 28137 2208
rect 27708 2066 27875 2082
rect 27708 2032 27841 2066
rect 27708 2016 27875 2032
rect 27708 1936 27771 2016
rect 27909 1982 27952 2106
rect 27986 2081 28057 2142
rect 27986 2047 28001 2081
rect 28035 2076 28057 2081
rect 27986 2042 28011 2047
rect 28045 2042 28057 2076
rect 27986 2012 28057 2042
rect 28091 2081 28137 2174
rect 28091 2047 28103 2081
rect 27708 1902 27721 1936
rect 27755 1902 27771 1936
rect 27900 1946 27952 1982
rect 28091 1978 28137 2047
rect 27708 1868 27771 1902
rect 27807 1910 27866 1926
rect 27807 1876 27816 1910
rect 27850 1876 27866 1910
rect 27807 1834 27866 1876
rect 27934 1912 27952 1946
rect 27900 1868 27952 1912
rect 27986 1944 28137 1978
rect 28206 2192 28217 2226
rect 28360 2210 28394 2260
rect 28172 2004 28217 2192
rect 28172 1970 28183 2004
rect 27986 1936 28038 1944
rect 27986 1902 28004 1936
rect 28172 1936 28217 1970
rect 28251 2176 28394 2210
rect 28251 1982 28285 2176
rect 28435 2174 28459 2208
rect 28493 2182 28535 2208
rect 28493 2174 28501 2182
rect 28435 2148 28501 2174
rect 28319 2071 28401 2142
rect 28319 2068 28348 2071
rect 28382 2037 28401 2071
rect 28353 2034 28401 2037
rect 28319 2018 28401 2034
rect 28435 2132 28535 2148
rect 28435 2008 28479 2132
rect 28569 2098 28603 2267
rect 28651 2292 28727 2344
rect 28945 2302 29011 2344
rect 28651 2258 28667 2292
rect 28701 2258 28727 2292
rect 28787 2276 28821 2292
rect 28787 2224 28821 2242
rect 28945 2268 28961 2302
rect 28995 2268 29011 2302
rect 29434 2302 29510 2344
rect 28945 2234 29011 2268
rect 29220 2267 29236 2301
rect 29270 2267 29386 2301
rect 29434 2268 29450 2302
rect 29484 2268 29510 2302
rect 29698 2302 29975 2344
rect 29558 2276 29592 2292
rect 28637 2208 28907 2224
rect 28637 2182 28787 2208
rect 28671 2174 28787 2182
rect 28821 2174 28907 2208
rect 28945 2200 28961 2234
rect 28995 2200 29011 2234
rect 29182 2208 29229 2214
rect 28671 2148 28687 2174
rect 28637 2132 28687 2148
rect 28789 2098 28839 2114
rect 28569 2064 28805 2098
rect 28569 2056 28649 2064
rect 28251 1944 28394 1982
rect 28469 1974 28479 2008
rect 28435 1958 28479 1974
rect 28515 1986 28531 2020
rect 28565 2004 28581 2020
rect 28515 1970 28547 1986
rect 28515 1946 28581 1970
rect 27986 1886 28038 1902
rect 28072 1876 28088 1910
rect 28122 1876 28138 1910
rect 28206 1902 28217 1936
rect 28360 1928 28394 1944
rect 28172 1886 28217 1902
rect 28072 1834 28138 1876
rect 28256 1876 28276 1910
rect 28310 1876 28326 1910
rect 28615 1910 28649 2056
rect 28795 2048 28839 2064
rect 28873 2030 28907 2174
rect 29182 2182 29195 2208
rect 29216 2148 29229 2174
rect 28941 2140 29142 2148
rect 28941 2106 29103 2140
rect 29137 2106 29142 2140
rect 29182 2132 29229 2148
rect 29277 2182 29318 2198
rect 29277 2148 29284 2182
rect 28941 2100 29142 2106
rect 28941 2098 29007 2100
rect 28941 2064 28957 2098
rect 28991 2064 29007 2098
rect 29277 2078 29318 2148
rect 29194 2072 29318 2078
rect 29069 2030 29085 2064
rect 29119 2030 29135 2064
rect 28687 1996 28703 2030
rect 28737 2010 28753 2030
rect 28737 2004 28769 2010
rect 28687 1970 28735 1996
rect 28873 1996 29135 2030
rect 29194 2038 29195 2072
rect 29229 2042 29318 2072
rect 29352 2098 29386 2267
rect 29698 2268 29714 2302
rect 29748 2268 29925 2302
rect 29959 2268 29975 2302
rect 29558 2234 29592 2242
rect 30009 2265 30066 2310
rect 29420 2200 29975 2234
rect 29420 2182 29470 2200
rect 29454 2148 29470 2182
rect 29420 2132 29470 2148
rect 29352 2082 29622 2098
rect 29352 2064 29588 2082
rect 29229 2038 29251 2042
rect 29194 2008 29251 2038
rect 28873 1970 28917 1996
rect 28687 1964 28769 1970
rect 28851 1936 28867 1970
rect 28901 1936 28917 1970
rect 29194 1974 29217 2008
rect 28951 1944 28985 1960
rect 29194 1958 29251 1974
rect 28360 1878 28394 1894
rect 28256 1834 28326 1876
rect 28450 1876 28466 1910
rect 28500 1876 28649 1910
rect 28450 1870 28649 1876
rect 28683 1906 28717 1922
rect 28683 1834 28717 1872
rect 28751 1892 28767 1926
rect 28801 1902 28817 1926
rect 29352 1910 29386 2064
rect 29578 2048 29588 2064
rect 29578 2032 29622 2048
rect 29461 2004 29480 2030
rect 29461 1970 29471 2004
rect 29514 1996 29536 2030
rect 29505 1970 29536 1996
rect 29656 1973 29692 2200
rect 29461 1964 29536 1970
rect 29626 1970 29692 1973
rect 29626 1936 29642 1970
rect 29676 1936 29692 1970
rect 29726 2140 29828 2166
rect 29726 2106 29747 2140
rect 29781 2132 29828 2140
rect 29862 2132 29878 2166
rect 29726 2098 29781 2106
rect 29760 2064 29781 2098
rect 29941 2082 29975 2200
rect 30043 2231 30066 2265
rect 30009 2197 30066 2231
rect 30043 2163 30066 2197
rect 30009 2143 30066 2163
rect 29726 2002 29781 2064
rect 29832 2071 29907 2082
rect 29832 2037 29856 2071
rect 29890 2070 29907 2071
rect 29832 2036 29857 2037
rect 29891 2036 29907 2070
rect 29941 2066 29991 2082
rect 29941 2032 29957 2066
rect 29941 2016 29991 2032
rect 29726 1968 29864 2002
rect 28951 1902 28985 1910
rect 28801 1892 28985 1902
rect 28751 1868 28985 1892
rect 29039 1876 29055 1910
rect 29089 1876 29105 1910
rect 29039 1834 29105 1876
rect 29233 1876 29249 1910
rect 29283 1876 29386 1910
rect 29233 1870 29386 1876
rect 29422 1906 29474 1922
rect 29422 1872 29440 1906
rect 29422 1834 29474 1872
rect 29526 1892 29542 1926
rect 29576 1902 29592 1926
rect 29726 1918 29760 1934
rect 29576 1892 29726 1902
rect 29526 1884 29726 1892
rect 29526 1868 29760 1884
rect 29817 1920 29864 1968
rect 29817 1886 29830 1920
rect 29817 1870 29864 1886
rect 29909 1910 29975 1978
rect 30025 1960 30066 2143
rect 29909 1876 29925 1910
rect 29959 1876 29975 1910
rect 29909 1834 29975 1876
rect 30009 1944 30066 1960
rect 30043 1910 30066 1944
rect 30009 1868 30066 1910
rect 30100 2284 30163 2300
rect 30100 2250 30113 2284
rect 30147 2250 30163 2284
rect 30100 2216 30163 2250
rect 30100 2182 30113 2216
rect 30147 2182 30163 2216
rect 30100 2082 30163 2182
rect 30199 2290 30258 2344
rect 30199 2256 30208 2290
rect 30242 2256 30258 2290
rect 30199 2222 30258 2256
rect 30199 2188 30208 2222
rect 30242 2188 30258 2222
rect 30199 2170 30258 2188
rect 30292 2266 30344 2310
rect 30326 2232 30344 2266
rect 30292 2198 30344 2232
rect 30326 2164 30344 2198
rect 30292 2106 30344 2164
rect 30100 2066 30267 2082
rect 30100 2032 30233 2066
rect 30100 2016 30267 2032
rect 30100 1936 30163 2016
rect 30301 1982 30344 2106
rect 30100 1902 30113 1936
rect 30147 1902 30163 1936
rect 30292 1946 30344 1982
rect 30326 1937 30344 1946
rect 30100 1868 30163 1902
rect 30199 1910 30258 1926
rect 30199 1876 30208 1910
rect 30242 1876 30258 1910
rect 30199 1834 30258 1876
rect 30292 1903 30294 1912
rect 30328 1903 30344 1937
rect 30292 1868 30344 1903
rect 25577 1766 25606 1834
rect 25640 1766 25698 1834
rect 25732 1766 25790 1834
rect 25824 1766 25882 1834
rect 25916 1766 25974 1834
rect 26008 1766 26066 1834
rect 26100 1766 26158 1834
rect 26192 1766 26250 1834
rect 26284 1766 26342 1834
rect 26376 1766 26434 1834
rect 26468 1766 26526 1834
rect 26560 1766 26618 1834
rect 26652 1766 26710 1834
rect 26744 1766 26802 1834
rect 26836 1766 26894 1834
rect 26928 1766 26986 1834
rect 27020 1766 27078 1834
rect 27112 1766 27170 1834
rect 27204 1766 27262 1834
rect 27296 1766 27354 1834
rect 27388 1766 27446 1834
rect 27480 1766 27538 1834
rect 27572 1766 27630 1834
rect 27664 1766 27722 1834
rect 27756 1766 27814 1834
rect 27848 1766 27906 1834
rect 27940 1766 27998 1834
rect 28032 1766 28090 1834
rect 28124 1766 28182 1834
rect 28216 1766 28274 1834
rect 28308 1766 28366 1834
rect 28400 1766 28458 1834
rect 28492 1766 28550 1834
rect 28584 1766 28642 1834
rect 28676 1766 28734 1834
rect 28768 1766 28826 1834
rect 28860 1766 28918 1834
rect 28952 1766 29010 1834
rect 29044 1766 29102 1834
rect 29136 1766 29194 1834
rect 29228 1766 29286 1834
rect 29320 1766 29378 1834
rect 29412 1766 29470 1834
rect 29504 1766 29562 1834
rect 29596 1766 29654 1834
rect 29688 1766 29746 1834
rect 29780 1766 29838 1834
rect 29872 1766 29930 1834
rect 29964 1766 30022 1834
rect 30056 1766 30114 1834
rect 30148 1766 30206 1834
rect 30240 1766 30298 1834
rect 30332 1766 30361 1834
rect 8577 1372 8606 1430
rect 8640 1372 8698 1430
rect 8732 1372 8790 1430
rect 8824 1372 8882 1430
rect 8916 1372 8974 1430
rect 9008 1372 9066 1430
rect 9100 1372 9158 1430
rect 9192 1372 9250 1430
rect 9284 1372 9342 1430
rect 9376 1372 9434 1430
rect 9468 1372 9526 1430
rect 9560 1372 9618 1430
rect 9652 1372 9710 1430
rect 9744 1372 9802 1430
rect 9836 1372 9894 1430
rect 9928 1372 9986 1430
rect 10020 1372 10078 1430
rect 10112 1372 10170 1430
rect 10204 1372 10262 1430
rect 10296 1372 10354 1430
rect 10388 1372 10446 1430
rect 10480 1372 10538 1430
rect 10572 1372 10630 1430
rect 10664 1372 10722 1430
rect 10756 1372 10814 1430
rect 10848 1372 10906 1430
rect 10940 1372 10998 1430
rect 11032 1372 11090 1430
rect 11124 1372 11182 1430
rect 11216 1372 11274 1430
rect 11308 1372 11366 1430
rect 11400 1372 11429 1430
rect 12961 1372 12990 1430
rect 13024 1372 13082 1430
rect 13116 1372 13174 1430
rect 13208 1372 13266 1430
rect 13300 1372 13358 1430
rect 13392 1372 13450 1430
rect 13484 1372 13542 1430
rect 13576 1372 13634 1430
rect 13668 1372 13726 1430
rect 13760 1372 13818 1430
rect 13852 1372 13910 1430
rect 13944 1372 14002 1430
rect 14036 1372 14094 1430
rect 14128 1372 14186 1430
rect 14220 1372 14278 1430
rect 14312 1372 14370 1430
rect 14404 1372 14462 1430
rect 14496 1372 14554 1430
rect 14588 1372 14646 1430
rect 14680 1372 14738 1430
rect 14772 1372 14830 1430
rect 14864 1372 14922 1430
rect 14956 1372 15014 1430
rect 15048 1372 15106 1430
rect 15140 1372 15198 1430
rect 15232 1372 15290 1430
rect 15324 1372 15382 1430
rect 15416 1372 15474 1430
rect 15508 1372 15566 1430
rect 15600 1372 15658 1430
rect 15692 1372 15750 1430
rect 15784 1372 15813 1430
rect 8610 1322 8646 1338
rect 8610 1288 8612 1322
rect 8610 1254 8646 1288
rect 8610 1220 8612 1254
rect 8682 1322 8748 1372
rect 8682 1288 8698 1322
rect 8732 1288 8748 1322
rect 8682 1254 8748 1288
rect 8682 1220 8698 1254
rect 8732 1220 8748 1254
rect 8782 1322 8836 1338
rect 8782 1288 8784 1322
rect 8818 1288 8836 1322
rect 8782 1241 8836 1288
rect 8610 1186 8646 1220
rect 8782 1207 8784 1241
rect 8818 1207 8836 1241
rect 8610 1152 8745 1186
rect 8782 1157 8836 1207
rect 8711 1123 8745 1152
rect 8598 1110 8666 1116
rect 8598 1060 8614 1110
rect 8648 1060 8666 1110
rect 8598 1042 8666 1060
rect 8711 1107 8766 1123
rect 8711 1073 8732 1107
rect 8711 1057 8766 1073
rect 8800 1105 8836 1157
rect 8872 1324 8938 1338
rect 8872 1290 8888 1324
rect 8922 1290 8938 1324
rect 8872 1256 8938 1290
rect 8872 1222 8888 1256
rect 8922 1222 8938 1256
rect 8872 1188 8938 1222
rect 8972 1330 9020 1372
rect 9006 1296 9020 1330
rect 8972 1262 9020 1296
rect 9006 1228 9020 1262
rect 8972 1212 9020 1228
rect 9056 1308 9090 1338
rect 9056 1213 9090 1274
rect 8872 1154 8888 1188
rect 8922 1176 8938 1188
rect 9124 1330 9190 1372
rect 9124 1296 9140 1330
rect 9174 1296 9190 1330
rect 9124 1262 9190 1296
rect 9124 1228 9140 1262
rect 9174 1228 9190 1262
rect 9124 1212 9190 1228
rect 9224 1308 9258 1338
rect 9224 1213 9258 1274
rect 8922 1154 9015 1176
rect 8872 1142 9015 1154
rect 8871 1105 8947 1108
rect 8800 1094 8947 1105
rect 8800 1061 8897 1094
rect 8711 1006 8745 1057
rect 8612 972 8745 1006
rect 8800 997 8836 1061
rect 8871 1060 8897 1061
rect 8931 1060 8947 1094
rect 8981 1094 9015 1142
rect 9056 1168 9090 1179
rect 9224 1168 9258 1179
rect 9056 1134 9258 1168
rect 9292 1330 9358 1372
rect 9292 1296 9308 1330
rect 9342 1296 9358 1330
rect 9292 1262 9358 1296
rect 9292 1228 9308 1262
rect 9342 1228 9358 1262
rect 9292 1194 9358 1228
rect 9292 1160 9308 1194
rect 9342 1160 9358 1194
rect 9292 1142 9358 1160
rect 9440 1330 9474 1372
rect 9440 1262 9474 1296
rect 9440 1194 9474 1228
rect 9440 1134 9474 1160
rect 9508 1324 9574 1338
rect 9508 1290 9524 1324
rect 9558 1290 9574 1324
rect 9508 1256 9574 1290
rect 9508 1222 9524 1256
rect 9558 1222 9574 1256
rect 9508 1188 9574 1222
rect 9608 1330 9642 1372
rect 9608 1262 9642 1296
rect 9608 1212 9642 1228
rect 9676 1324 9742 1338
rect 9676 1290 9692 1324
rect 9726 1290 9742 1324
rect 9676 1256 9742 1290
rect 9676 1222 9692 1256
rect 9726 1222 9742 1256
rect 9508 1154 9524 1188
rect 9558 1168 9574 1188
rect 9676 1188 9742 1222
rect 9776 1330 9810 1372
rect 9776 1262 9810 1296
rect 9776 1212 9810 1228
rect 9844 1324 9910 1338
rect 9844 1290 9860 1324
rect 9894 1290 9910 1324
rect 9844 1256 9910 1290
rect 9844 1222 9860 1256
rect 9894 1222 9910 1256
rect 9676 1168 9692 1188
rect 9558 1154 9692 1168
rect 9726 1168 9742 1188
rect 9844 1188 9910 1222
rect 9944 1330 9978 1372
rect 9944 1262 9978 1296
rect 9944 1212 9978 1228
rect 10012 1324 10078 1338
rect 10012 1290 10028 1324
rect 10062 1290 10078 1324
rect 10012 1256 10078 1290
rect 10012 1222 10028 1256
rect 10062 1222 10078 1256
rect 9844 1168 9860 1188
rect 9726 1154 9860 1168
rect 9894 1168 9910 1188
rect 10012 1188 10078 1222
rect 10112 1330 10146 1372
rect 10112 1262 10146 1296
rect 10112 1212 10146 1228
rect 10180 1324 10246 1338
rect 10180 1290 10196 1324
rect 10230 1290 10246 1324
rect 10180 1256 10246 1290
rect 10180 1222 10196 1256
rect 10230 1222 10246 1256
rect 9894 1154 9978 1168
rect 9508 1134 9978 1154
rect 10012 1154 10028 1188
rect 10062 1168 10078 1188
rect 10180 1188 10246 1222
rect 10280 1330 10314 1372
rect 10280 1262 10314 1296
rect 10280 1212 10314 1228
rect 10348 1324 10414 1338
rect 10348 1290 10364 1324
rect 10398 1290 10414 1324
rect 10348 1256 10414 1290
rect 10348 1222 10364 1256
rect 10398 1222 10414 1256
rect 10180 1168 10196 1188
rect 10062 1154 10196 1168
rect 10230 1168 10246 1188
rect 10348 1188 10414 1222
rect 10448 1330 10482 1372
rect 10448 1262 10482 1296
rect 10448 1212 10482 1228
rect 10516 1324 10582 1338
rect 10516 1290 10532 1324
rect 10566 1290 10582 1324
rect 10516 1256 10582 1290
rect 10516 1222 10532 1256
rect 10566 1222 10582 1256
rect 10348 1168 10364 1188
rect 10230 1154 10364 1168
rect 10398 1168 10414 1188
rect 10516 1188 10582 1222
rect 10616 1330 10650 1372
rect 10616 1262 10650 1296
rect 10616 1212 10650 1228
rect 10684 1324 10750 1338
rect 10684 1290 10700 1324
rect 10734 1290 10750 1324
rect 10684 1256 10750 1290
rect 10684 1222 10700 1256
rect 10734 1222 10750 1256
rect 10516 1168 10532 1188
rect 10398 1154 10532 1168
rect 10566 1168 10582 1188
rect 10684 1188 10750 1222
rect 10784 1330 10818 1372
rect 10784 1262 10818 1296
rect 10784 1212 10818 1228
rect 10852 1324 10918 1338
rect 10852 1290 10868 1324
rect 10902 1290 10918 1324
rect 10852 1256 10918 1290
rect 10852 1222 10868 1256
rect 10902 1222 10918 1256
rect 10684 1168 10700 1188
rect 10566 1154 10700 1168
rect 10734 1168 10750 1188
rect 10852 1188 10918 1222
rect 10952 1330 10986 1372
rect 10952 1262 10986 1296
rect 10952 1212 10986 1228
rect 11020 1324 11086 1338
rect 11020 1290 11036 1324
rect 11070 1290 11086 1324
rect 11020 1256 11086 1290
rect 11020 1222 11036 1256
rect 11070 1222 11086 1256
rect 10852 1168 10868 1188
rect 10734 1154 10868 1168
rect 10902 1168 10918 1188
rect 11020 1188 11086 1222
rect 11120 1330 11154 1372
rect 11120 1262 11154 1296
rect 11120 1212 11154 1228
rect 11188 1324 11254 1338
rect 11188 1290 11204 1324
rect 11238 1290 11254 1324
rect 11188 1256 11254 1290
rect 11188 1222 11204 1256
rect 11238 1222 11254 1256
rect 11020 1168 11036 1188
rect 10902 1154 11036 1168
rect 11070 1168 11086 1188
rect 11188 1188 11254 1222
rect 11288 1330 11322 1372
rect 12994 1322 13030 1338
rect 11288 1262 11322 1296
rect 11288 1212 11322 1228
rect 11188 1168 11204 1188
rect 11070 1154 11204 1168
rect 11238 1168 11254 1188
rect 11357 1168 11412 1317
rect 11238 1154 11412 1168
rect 10012 1134 11412 1154
rect 12994 1288 12996 1322
rect 12994 1254 13030 1288
rect 12994 1220 12996 1254
rect 13066 1322 13132 1372
rect 13066 1288 13082 1322
rect 13116 1288 13132 1322
rect 13066 1254 13132 1288
rect 13066 1220 13082 1254
rect 13116 1220 13132 1254
rect 13166 1322 13220 1338
rect 13166 1288 13168 1322
rect 13202 1288 13220 1322
rect 13166 1241 13220 1288
rect 12994 1186 13030 1220
rect 13166 1207 13168 1241
rect 13202 1207 13220 1241
rect 12994 1152 13129 1186
rect 13166 1157 13220 1207
rect 9159 1099 9258 1134
rect 9943 1100 9978 1134
rect 11336 1100 11412 1134
rect 13095 1123 13129 1152
rect 9422 1099 9902 1100
rect 9159 1094 9902 1099
rect 8981 1060 9031 1094
rect 9065 1060 9081 1094
rect 9159 1061 9508 1094
rect 8981 1026 9015 1060
rect 9159 1026 9258 1061
rect 9422 1060 9508 1061
rect 9542 1060 9576 1094
rect 9610 1060 9644 1094
rect 9678 1060 9712 1094
rect 9746 1060 9780 1094
rect 9814 1060 9848 1094
rect 9882 1060 9902 1094
rect 9943 1094 11287 1100
rect 9943 1060 10008 1094
rect 10042 1060 10076 1094
rect 10110 1060 10144 1094
rect 10178 1060 10212 1094
rect 10246 1060 10280 1094
rect 10314 1060 10348 1094
rect 10382 1060 10416 1094
rect 10450 1060 10484 1094
rect 10518 1060 10552 1094
rect 10586 1060 10620 1094
rect 10654 1060 10688 1094
rect 10722 1060 10756 1094
rect 10790 1060 10824 1094
rect 10858 1060 10892 1094
rect 10926 1060 10960 1094
rect 10994 1060 11028 1094
rect 11062 1060 11096 1094
rect 11130 1060 11164 1094
rect 11198 1060 11232 1094
rect 11266 1060 11287 1094
rect 11336 1099 11490 1100
rect 11336 1065 11451 1099
rect 11485 1065 11490 1099
rect 11336 1064 11490 1065
rect 12982 1094 13050 1116
rect 9943 1026 9978 1060
rect 11336 1026 11412 1064
rect 12982 1059 12998 1094
rect 13032 1059 13050 1094
rect 12982 1042 13050 1059
rect 13095 1107 13150 1123
rect 13095 1073 13116 1107
rect 13095 1057 13150 1073
rect 13184 1107 13220 1157
rect 13256 1324 13322 1338
rect 13256 1290 13272 1324
rect 13306 1290 13322 1324
rect 13256 1256 13322 1290
rect 13256 1222 13272 1256
rect 13306 1222 13322 1256
rect 13256 1188 13322 1222
rect 13356 1330 13404 1372
rect 13390 1296 13404 1330
rect 13356 1262 13404 1296
rect 13390 1228 13404 1262
rect 13356 1212 13404 1228
rect 13440 1308 13474 1338
rect 13440 1213 13474 1274
rect 13256 1154 13272 1188
rect 13306 1176 13322 1188
rect 13508 1330 13574 1372
rect 13508 1296 13524 1330
rect 13558 1296 13574 1330
rect 13508 1262 13574 1296
rect 13508 1228 13524 1262
rect 13558 1228 13574 1262
rect 13508 1212 13574 1228
rect 13608 1308 13642 1338
rect 13608 1213 13642 1274
rect 13306 1154 13399 1176
rect 13256 1142 13399 1154
rect 13255 1107 13331 1108
rect 13184 1094 13331 1107
rect 13184 1061 13281 1094
rect 8612 951 8646 972
rect 8784 968 8836 997
rect 8612 896 8646 917
rect 8682 904 8698 938
rect 8732 904 8748 938
rect 8682 862 8748 904
rect 8818 934 8836 968
rect 8784 896 8836 934
rect 8888 992 9015 1026
rect 9056 992 9258 1026
rect 8888 974 8922 992
rect 9056 974 9090 992
rect 8888 896 8922 940
rect 8958 942 9006 958
rect 8958 908 8972 942
rect 8958 862 9006 908
rect 9224 974 9258 992
rect 9056 896 9090 940
rect 9124 942 9190 958
rect 9124 908 9140 942
rect 9174 908 9190 942
rect 9124 862 9190 908
rect 9224 896 9258 940
rect 9292 1006 9358 1022
rect 9292 972 9308 1006
rect 9342 972 9358 1006
rect 9292 938 9358 972
rect 9292 904 9308 938
rect 9342 904 9358 938
rect 9292 862 9358 904
rect 9440 1010 9474 1026
rect 9440 942 9474 976
rect 9440 862 9474 908
rect 9508 1010 9978 1026
rect 9508 976 9524 1010
rect 9558 992 9692 1010
rect 9558 976 9574 992
rect 9508 942 9574 976
rect 9676 976 9692 992
rect 9726 992 9860 1010
rect 9726 976 9742 992
rect 9508 908 9524 942
rect 9558 908 9574 942
rect 9508 897 9574 908
rect 9608 942 9642 958
rect 9608 862 9642 908
rect 9676 942 9742 976
rect 9844 976 9860 992
rect 9894 992 9978 1010
rect 10012 1010 11412 1026
rect 9894 976 9910 992
rect 9676 908 9692 942
rect 9726 908 9742 942
rect 9676 897 9742 908
rect 9776 942 9810 958
rect 9776 862 9810 908
rect 9844 942 9910 976
rect 10012 976 10028 1010
rect 10062 992 10196 1010
rect 10062 976 10078 992
rect 9844 908 9860 942
rect 9894 908 9910 942
rect 9844 897 9910 908
rect 9944 942 9978 958
rect 9944 862 9978 908
rect 10012 942 10078 976
rect 10180 976 10196 992
rect 10230 992 10364 1010
rect 10230 976 10246 992
rect 10012 908 10028 942
rect 10062 908 10078 942
rect 10012 897 10078 908
rect 10112 942 10146 958
rect 10012 896 10062 897
rect 10112 862 10146 908
rect 10180 942 10246 976
rect 10348 976 10364 992
rect 10398 992 10532 1010
rect 10398 976 10414 992
rect 10180 908 10196 942
rect 10230 908 10246 942
rect 10180 897 10246 908
rect 10280 942 10314 958
rect 10196 896 10230 897
rect 10280 862 10314 908
rect 10348 942 10414 976
rect 10516 976 10532 992
rect 10566 992 10700 1010
rect 10566 976 10582 992
rect 10348 908 10364 942
rect 10398 908 10414 942
rect 10348 897 10414 908
rect 10448 942 10482 958
rect 10364 896 10398 897
rect 10448 862 10482 908
rect 10516 942 10582 976
rect 10684 976 10700 992
rect 10734 992 10868 1010
rect 10734 976 10750 992
rect 10516 908 10532 942
rect 10566 908 10582 942
rect 10516 897 10582 908
rect 10616 942 10650 958
rect 10616 862 10650 908
rect 10684 942 10750 976
rect 10852 976 10868 992
rect 10902 992 11036 1010
rect 10902 976 10918 992
rect 10684 908 10700 942
rect 10734 908 10750 942
rect 10684 897 10750 908
rect 10784 942 10818 958
rect 10784 862 10818 908
rect 10852 942 10918 976
rect 11020 976 11036 992
rect 11070 992 11204 1010
rect 11070 976 11086 992
rect 10852 908 10868 942
rect 10902 908 10918 942
rect 10852 897 10918 908
rect 10952 942 10986 958
rect 10952 862 10986 908
rect 11020 942 11086 976
rect 11188 976 11204 992
rect 11238 992 11412 1010
rect 13095 1006 13129 1057
rect 11238 976 11254 992
rect 11020 908 11036 942
rect 11070 908 11086 942
rect 11020 897 11086 908
rect 11120 942 11154 958
rect 11120 862 11154 908
rect 11188 942 11254 976
rect 11188 908 11204 942
rect 11238 908 11254 942
rect 11188 897 11254 908
rect 11288 942 11322 958
rect 11357 918 11412 992
rect 12996 972 13129 1006
rect 13184 997 13220 1061
rect 13255 1060 13281 1061
rect 13315 1060 13331 1094
rect 13365 1094 13399 1142
rect 13440 1168 13474 1179
rect 13608 1168 13642 1179
rect 13440 1134 13642 1168
rect 13676 1330 13742 1372
rect 13676 1296 13692 1330
rect 13726 1296 13742 1330
rect 13676 1262 13742 1296
rect 13676 1228 13692 1262
rect 13726 1228 13742 1262
rect 13676 1194 13742 1228
rect 13676 1160 13692 1194
rect 13726 1160 13742 1194
rect 13676 1142 13742 1160
rect 13824 1330 13858 1372
rect 13824 1262 13858 1296
rect 13824 1194 13858 1228
rect 13824 1134 13858 1160
rect 13892 1324 13958 1338
rect 13892 1290 13908 1324
rect 13942 1290 13958 1324
rect 13892 1256 13958 1290
rect 13892 1222 13908 1256
rect 13942 1222 13958 1256
rect 13892 1188 13958 1222
rect 13992 1330 14026 1372
rect 13992 1262 14026 1296
rect 13992 1212 14026 1228
rect 14060 1324 14126 1338
rect 14060 1290 14076 1324
rect 14110 1290 14126 1324
rect 14060 1256 14126 1290
rect 14060 1222 14076 1256
rect 14110 1222 14126 1256
rect 13892 1154 13908 1188
rect 13942 1168 13958 1188
rect 14060 1188 14126 1222
rect 14160 1330 14194 1372
rect 14160 1262 14194 1296
rect 14160 1212 14194 1228
rect 14228 1324 14294 1338
rect 14228 1290 14244 1324
rect 14278 1290 14294 1324
rect 14228 1256 14294 1290
rect 14228 1222 14244 1256
rect 14278 1222 14294 1256
rect 14060 1168 14076 1188
rect 13942 1154 14076 1168
rect 14110 1168 14126 1188
rect 14228 1188 14294 1222
rect 14328 1330 14362 1372
rect 14328 1262 14362 1296
rect 14328 1212 14362 1228
rect 14396 1324 14462 1338
rect 14396 1290 14412 1324
rect 14446 1290 14462 1324
rect 14396 1256 14462 1290
rect 14396 1222 14412 1256
rect 14446 1222 14462 1256
rect 14228 1168 14244 1188
rect 14110 1154 14244 1168
rect 14278 1168 14294 1188
rect 14396 1188 14462 1222
rect 14496 1330 14530 1372
rect 14496 1262 14530 1296
rect 14496 1212 14530 1228
rect 14564 1324 14630 1338
rect 14564 1290 14580 1324
rect 14614 1290 14630 1324
rect 14564 1256 14630 1290
rect 14564 1222 14580 1256
rect 14614 1222 14630 1256
rect 14278 1154 14362 1168
rect 13892 1134 14362 1154
rect 14396 1154 14412 1188
rect 14446 1168 14462 1188
rect 14564 1188 14630 1222
rect 14664 1330 14698 1372
rect 14664 1262 14698 1296
rect 14664 1212 14698 1228
rect 14732 1324 14798 1338
rect 14732 1290 14748 1324
rect 14782 1290 14798 1324
rect 14732 1256 14798 1290
rect 14732 1222 14748 1256
rect 14782 1222 14798 1256
rect 14564 1168 14580 1188
rect 14446 1154 14580 1168
rect 14614 1168 14630 1188
rect 14732 1188 14798 1222
rect 14832 1330 14866 1372
rect 14832 1262 14866 1296
rect 14832 1212 14866 1228
rect 14900 1324 14966 1338
rect 14900 1290 14916 1324
rect 14950 1290 14966 1324
rect 14900 1256 14966 1290
rect 14900 1222 14916 1256
rect 14950 1222 14966 1256
rect 14732 1168 14748 1188
rect 14614 1154 14748 1168
rect 14782 1168 14798 1188
rect 14900 1188 14966 1222
rect 15000 1330 15034 1372
rect 15000 1262 15034 1296
rect 15000 1212 15034 1228
rect 15068 1324 15134 1338
rect 15068 1290 15084 1324
rect 15118 1290 15134 1324
rect 15068 1256 15134 1290
rect 15068 1222 15084 1256
rect 15118 1222 15134 1256
rect 14900 1168 14916 1188
rect 14782 1154 14916 1168
rect 14950 1168 14966 1188
rect 15068 1188 15134 1222
rect 15168 1330 15202 1372
rect 15168 1262 15202 1296
rect 15168 1212 15202 1228
rect 15236 1324 15302 1338
rect 15236 1290 15252 1324
rect 15286 1290 15302 1324
rect 15236 1256 15302 1290
rect 15236 1222 15252 1256
rect 15286 1222 15302 1256
rect 15068 1168 15084 1188
rect 14950 1154 15084 1168
rect 15118 1168 15134 1188
rect 15236 1188 15302 1222
rect 15336 1330 15370 1372
rect 15336 1262 15370 1296
rect 15336 1212 15370 1228
rect 15404 1324 15470 1338
rect 15404 1290 15420 1324
rect 15454 1290 15470 1324
rect 15404 1256 15470 1290
rect 15404 1222 15420 1256
rect 15454 1222 15470 1256
rect 15236 1168 15252 1188
rect 15118 1154 15252 1168
rect 15286 1168 15302 1188
rect 15404 1188 15470 1222
rect 15504 1330 15538 1372
rect 15504 1262 15538 1296
rect 15504 1212 15538 1228
rect 15572 1324 15638 1338
rect 15572 1290 15588 1324
rect 15622 1290 15638 1324
rect 15572 1256 15638 1290
rect 15572 1222 15588 1256
rect 15622 1222 15638 1256
rect 15404 1168 15420 1188
rect 15286 1154 15420 1168
rect 15454 1168 15470 1188
rect 15572 1188 15638 1222
rect 15672 1330 15706 1372
rect 15672 1262 15706 1296
rect 15672 1212 15706 1228
rect 15572 1168 15588 1188
rect 15454 1154 15588 1168
rect 15622 1168 15638 1188
rect 15741 1168 15796 1317
rect 15622 1154 15796 1168
rect 14396 1134 15796 1154
rect 13543 1101 13642 1134
rect 13543 1100 13813 1101
rect 14327 1100 14362 1134
rect 15720 1101 15796 1134
rect 13543 1094 14286 1100
rect 13365 1060 13415 1094
rect 13449 1060 13465 1094
rect 13543 1061 13892 1094
rect 13365 1026 13399 1060
rect 13543 1026 13642 1061
rect 13806 1060 13892 1061
rect 13926 1060 13960 1094
rect 13994 1060 14028 1094
rect 14062 1060 14096 1094
rect 14130 1060 14164 1094
rect 14198 1060 14232 1094
rect 14266 1060 14286 1094
rect 14327 1094 15671 1100
rect 14327 1060 14392 1094
rect 14426 1060 14460 1094
rect 14494 1060 14528 1094
rect 14562 1060 14596 1094
rect 14630 1060 14664 1094
rect 14698 1060 14732 1094
rect 14766 1060 14800 1094
rect 14834 1060 14868 1094
rect 14902 1060 14936 1094
rect 14970 1060 15004 1094
rect 15038 1060 15072 1094
rect 15106 1060 15140 1094
rect 15174 1060 15208 1094
rect 15242 1060 15276 1094
rect 15310 1060 15344 1094
rect 15378 1060 15412 1094
rect 15446 1060 15480 1094
rect 15514 1060 15548 1094
rect 15582 1060 15616 1094
rect 15650 1060 15671 1094
rect 15720 1067 15751 1101
rect 15785 1067 15796 1101
rect 14327 1026 14362 1060
rect 15720 1026 15796 1067
rect 12996 951 13030 972
rect 11288 862 11322 908
rect 13168 968 13220 997
rect 12996 896 13030 917
rect 13066 904 13082 938
rect 13116 904 13132 938
rect 13066 862 13132 904
rect 13202 934 13220 968
rect 13168 896 13220 934
rect 13272 992 13399 1026
rect 13440 992 13642 1026
rect 13272 974 13306 992
rect 13440 974 13474 992
rect 13272 896 13306 940
rect 13342 942 13390 958
rect 13342 908 13356 942
rect 13342 862 13390 908
rect 13608 974 13642 992
rect 13440 896 13474 940
rect 13508 942 13574 958
rect 13508 908 13524 942
rect 13558 908 13574 942
rect 13508 862 13574 908
rect 13608 896 13642 940
rect 13676 1006 13742 1022
rect 13676 972 13692 1006
rect 13726 972 13742 1006
rect 13676 938 13742 972
rect 13676 904 13692 938
rect 13726 904 13742 938
rect 13676 862 13742 904
rect 13824 1010 13858 1026
rect 13824 942 13858 976
rect 13824 862 13858 908
rect 13892 1010 14362 1026
rect 13892 976 13908 1010
rect 13942 992 14076 1010
rect 13942 976 13958 992
rect 13892 942 13958 976
rect 14060 976 14076 992
rect 14110 992 14244 1010
rect 14110 976 14126 992
rect 13892 908 13908 942
rect 13942 908 13958 942
rect 13892 897 13958 908
rect 13992 942 14026 958
rect 13992 862 14026 908
rect 14060 942 14126 976
rect 14228 976 14244 992
rect 14278 992 14362 1010
rect 14396 1010 15796 1026
rect 14278 976 14294 992
rect 14060 908 14076 942
rect 14110 908 14126 942
rect 14060 897 14126 908
rect 14160 942 14194 958
rect 14160 862 14194 908
rect 14228 942 14294 976
rect 14396 976 14412 1010
rect 14446 992 14580 1010
rect 14446 976 14462 992
rect 14228 908 14244 942
rect 14278 908 14294 942
rect 14228 897 14294 908
rect 14328 942 14362 958
rect 14328 862 14362 908
rect 14396 942 14462 976
rect 14564 976 14580 992
rect 14614 992 14748 1010
rect 14614 976 14630 992
rect 14396 908 14412 942
rect 14446 908 14462 942
rect 14396 897 14462 908
rect 14496 942 14530 958
rect 14396 896 14446 897
rect 14496 862 14530 908
rect 14564 942 14630 976
rect 14732 976 14748 992
rect 14782 992 14916 1010
rect 14782 976 14798 992
rect 14564 908 14580 942
rect 14614 908 14630 942
rect 14564 897 14630 908
rect 14664 942 14698 958
rect 14580 896 14614 897
rect 14664 862 14698 908
rect 14732 942 14798 976
rect 14900 976 14916 992
rect 14950 992 15084 1010
rect 14950 976 14966 992
rect 14732 908 14748 942
rect 14782 908 14798 942
rect 14732 897 14798 908
rect 14832 942 14866 958
rect 14748 896 14782 897
rect 14832 862 14866 908
rect 14900 942 14966 976
rect 15068 976 15084 992
rect 15118 992 15252 1010
rect 15118 976 15134 992
rect 14900 908 14916 942
rect 14950 908 14966 942
rect 14900 897 14966 908
rect 15000 942 15034 958
rect 15000 862 15034 908
rect 15068 942 15134 976
rect 15236 976 15252 992
rect 15286 992 15420 1010
rect 15286 976 15302 992
rect 15068 908 15084 942
rect 15118 908 15134 942
rect 15068 897 15134 908
rect 15168 942 15202 958
rect 15168 862 15202 908
rect 15236 942 15302 976
rect 15404 976 15420 992
rect 15454 992 15588 1010
rect 15454 976 15470 992
rect 15236 908 15252 942
rect 15286 908 15302 942
rect 15236 897 15302 908
rect 15336 942 15370 958
rect 15336 862 15370 908
rect 15404 942 15470 976
rect 15572 976 15588 992
rect 15622 992 15796 1010
rect 15622 976 15638 992
rect 15404 908 15420 942
rect 15454 908 15470 942
rect 15404 897 15470 908
rect 15504 942 15538 958
rect 15504 862 15538 908
rect 15572 942 15638 976
rect 15572 908 15588 942
rect 15622 908 15638 942
rect 15572 897 15638 908
rect 15672 942 15706 958
rect 15741 918 15796 992
rect 15672 862 15706 908
rect 8577 804 8606 862
rect 8640 804 8698 862
rect 8732 804 8790 862
rect 8824 804 8882 862
rect 8916 804 8974 862
rect 9008 804 9066 862
rect 9100 804 9158 862
rect 9192 804 9250 862
rect 9284 804 9342 862
rect 9376 804 9434 862
rect 9468 804 9526 862
rect 9560 804 9618 862
rect 9652 804 9710 862
rect 9744 804 9802 862
rect 9836 804 9894 862
rect 9928 804 9986 862
rect 10020 804 10078 862
rect 10112 804 10170 862
rect 10204 804 10262 862
rect 10296 804 10354 862
rect 10388 804 10446 862
rect 10480 804 10538 862
rect 10572 804 10630 862
rect 10664 804 10722 862
rect 10756 804 10814 862
rect 10848 804 10906 862
rect 10940 804 10998 862
rect 11032 804 11090 862
rect 11124 804 11182 862
rect 11216 804 11274 862
rect 11308 804 11366 862
rect 11400 804 11429 862
rect 12961 804 12990 862
rect 13024 804 13082 862
rect 13116 804 13174 862
rect 13208 804 13266 862
rect 13300 804 13358 862
rect 13392 804 13450 862
rect 13484 804 13542 862
rect 13576 804 13634 862
rect 13668 804 13726 862
rect 13760 804 13818 862
rect 13852 804 13910 862
rect 13944 804 14002 862
rect 14036 804 14094 862
rect 14128 804 14186 862
rect 14220 804 14278 862
rect 14312 804 14370 862
rect 14404 804 14462 862
rect 14496 804 14554 862
rect 14588 804 14646 862
rect 14680 804 14738 862
rect 14772 804 14830 862
rect 14864 804 14922 862
rect 14956 804 15014 862
rect 15048 804 15106 862
rect 15140 804 15198 862
rect 15232 804 15290 862
rect 15324 804 15382 862
rect 15416 804 15474 862
rect 15508 804 15566 862
rect 15600 804 15658 862
rect 15692 804 15750 862
rect 15784 804 15813 862
rect 8575 230 8604 288
rect 8638 230 8696 288
rect 8730 230 8788 288
rect 8822 230 8880 288
rect 8914 230 8972 288
rect 9006 230 9064 288
rect 9098 230 9156 288
rect 9190 230 9248 288
rect 9282 230 9340 288
rect 9374 254 9432 288
rect 9466 254 9524 288
rect 9558 254 9616 288
rect 9650 254 9708 288
rect 9742 254 9800 288
rect 9834 254 9892 288
rect 9926 254 9984 288
rect 10018 264 10076 288
rect 10018 254 10038 264
rect 9374 239 10038 254
rect 9374 230 9403 239
rect 10009 230 10038 239
rect 10072 254 10076 264
rect 10110 264 10168 288
rect 10110 254 10130 264
rect 10072 230 10130 254
rect 10164 254 10168 264
rect 10202 264 10260 288
rect 10202 254 10222 264
rect 10164 230 10222 254
rect 10256 254 10260 264
rect 10294 264 10352 288
rect 10294 254 10314 264
rect 10256 230 10314 254
rect 10348 254 10352 264
rect 10386 264 10444 288
rect 10386 254 10406 264
rect 10348 230 10406 254
rect 10440 254 10444 264
rect 10478 264 10536 288
rect 10478 254 10498 264
rect 10440 230 10498 254
rect 10532 254 10536 264
rect 10570 264 10628 288
rect 10570 254 10590 264
rect 10532 230 10590 254
rect 10624 254 10628 264
rect 10662 264 10720 288
rect 10662 254 10682 264
rect 10624 230 10682 254
rect 10716 254 10720 264
rect 10754 264 10812 288
rect 10754 254 10774 264
rect 10716 230 10774 254
rect 10808 254 10812 264
rect 10846 254 10904 288
rect 10938 254 10996 288
rect 10808 239 10996 254
rect 10808 230 10837 239
rect 10967 230 10996 239
rect 11030 230 11088 288
rect 11122 230 11180 288
rect 11214 230 11272 288
rect 11306 230 11364 288
rect 11398 230 11456 288
rect 11490 230 11548 288
rect 11582 230 11640 288
rect 11674 230 11732 288
rect 11766 254 11824 288
rect 11858 254 11916 288
rect 11950 254 12008 288
rect 12042 254 12100 288
rect 12134 254 12192 288
rect 12226 254 12284 288
rect 12318 254 12376 288
rect 12410 264 12468 288
rect 12410 254 12430 264
rect 11766 239 12430 254
rect 11766 230 11795 239
rect 12401 230 12430 239
rect 12464 254 12468 264
rect 12502 264 12560 288
rect 12502 254 12522 264
rect 12464 230 12522 254
rect 12556 254 12560 264
rect 12594 264 12652 288
rect 12594 254 12614 264
rect 12556 230 12614 254
rect 12648 254 12652 264
rect 12686 264 12744 288
rect 12686 254 12706 264
rect 12648 230 12706 254
rect 12740 254 12744 264
rect 12778 264 12836 288
rect 12778 254 12798 264
rect 12740 230 12798 254
rect 12832 254 12836 264
rect 12870 264 12928 288
rect 12870 254 12890 264
rect 12832 230 12890 254
rect 12924 254 12928 264
rect 12962 264 13020 288
rect 12962 254 12982 264
rect 12924 230 12982 254
rect 13016 254 13020 264
rect 13054 264 13112 288
rect 13054 254 13074 264
rect 13016 230 13074 254
rect 13108 254 13112 264
rect 13146 264 13204 288
rect 13146 254 13166 264
rect 13108 230 13166 254
rect 13200 254 13204 264
rect 13238 254 13296 288
rect 13330 254 13388 288
rect 13200 239 13388 254
rect 13200 230 13229 239
rect 13359 230 13388 239
rect 13422 230 13480 288
rect 13514 230 13572 288
rect 13606 230 13664 288
rect 13698 230 13756 288
rect 13790 230 13848 288
rect 13882 230 13940 288
rect 13974 230 14032 288
rect 14066 230 14124 288
rect 14158 254 14216 288
rect 14250 254 14820 288
rect 14158 239 14820 254
rect 14158 230 14187 239
rect 14791 230 14820 239
rect 14854 230 14912 288
rect 14946 230 15004 288
rect 15038 230 15096 288
rect 15130 230 15188 288
rect 15222 230 15280 288
rect 15314 230 15372 288
rect 15406 230 15464 288
rect 15498 230 15556 288
rect 15590 254 15648 288
rect 15682 254 15740 288
rect 15774 264 15832 288
rect 15774 254 15780 264
rect 15590 239 15780 254
rect 15590 230 15619 239
rect 15751 230 15780 239
rect 15814 254 15832 264
rect 15866 264 15924 288
rect 15866 254 15872 264
rect 15814 230 15872 254
rect 15906 254 15924 264
rect 15958 264 16016 288
rect 15958 254 15964 264
rect 15906 230 15964 254
rect 15998 254 16016 264
rect 16050 264 16108 288
rect 16050 254 16056 264
rect 15998 230 16056 254
rect 16090 254 16108 264
rect 16142 264 16200 288
rect 16142 254 16148 264
rect 16090 230 16148 254
rect 16182 254 16200 264
rect 16234 264 16292 288
rect 16234 254 16240 264
rect 16182 230 16240 254
rect 16274 254 16292 264
rect 16326 264 16384 288
rect 16326 254 16332 264
rect 16274 230 16332 254
rect 16366 254 16384 264
rect 16418 264 16476 288
rect 16418 254 16424 264
rect 16366 230 16424 254
rect 16458 254 16476 264
rect 16510 264 16568 288
rect 16510 254 16516 264
rect 16458 230 16516 254
rect 16550 254 16568 264
rect 16602 254 16660 288
rect 16694 254 16752 288
rect 16786 254 16844 288
rect 16878 254 16936 288
rect 16970 254 17028 288
rect 17062 254 17120 288
rect 17154 254 17212 288
rect 17246 264 17304 288
rect 17338 264 17396 288
rect 17430 264 17488 288
rect 17522 264 17580 288
rect 17614 264 17672 288
rect 17706 264 17764 288
rect 17798 264 17856 288
rect 17890 264 17948 288
rect 17982 264 18040 288
rect 17248 254 17304 264
rect 17340 254 17396 264
rect 17432 254 17488 264
rect 17524 254 17580 264
rect 17616 254 17672 264
rect 17708 254 17764 264
rect 17800 254 17856 264
rect 17892 254 17948 264
rect 17984 254 18040 264
rect 18074 254 18132 288
rect 18166 264 18224 288
rect 18166 254 18172 264
rect 16550 239 17214 254
rect 16550 230 16579 239
rect 17185 230 17214 239
rect 17248 230 17306 254
rect 17340 230 17398 254
rect 17432 230 17490 254
rect 17524 230 17582 254
rect 17616 230 17674 254
rect 17708 230 17766 254
rect 17800 230 17858 254
rect 17892 230 17950 254
rect 17984 239 18172 254
rect 17984 230 18013 239
rect 18143 230 18172 239
rect 18206 254 18224 264
rect 18258 264 18316 288
rect 18258 254 18264 264
rect 18206 230 18264 254
rect 18298 254 18316 264
rect 18350 264 18408 288
rect 18350 254 18356 264
rect 18298 230 18356 254
rect 18390 254 18408 264
rect 18442 264 18500 288
rect 18442 254 18448 264
rect 18390 230 18448 254
rect 18482 254 18500 264
rect 18534 264 18592 288
rect 18534 254 18540 264
rect 18482 230 18540 254
rect 18574 254 18592 264
rect 18626 264 18684 288
rect 18626 254 18632 264
rect 18574 230 18632 254
rect 18666 254 18684 264
rect 18718 264 18776 288
rect 18718 254 18724 264
rect 18666 230 18724 254
rect 18758 254 18776 264
rect 18810 264 18868 288
rect 18810 254 18816 264
rect 18758 230 18816 254
rect 18850 254 18868 264
rect 18902 264 18960 288
rect 18902 254 18908 264
rect 18850 230 18908 254
rect 18942 254 18960 264
rect 18994 254 19052 288
rect 19086 254 19144 288
rect 19178 254 19236 288
rect 19270 254 19328 288
rect 19362 254 19420 288
rect 19454 254 19512 288
rect 19546 254 19604 288
rect 19638 264 19696 288
rect 19730 264 19788 288
rect 19822 264 19880 288
rect 19914 264 19972 288
rect 20006 264 20064 288
rect 20098 264 20156 288
rect 20190 264 20248 288
rect 20282 264 20340 288
rect 20374 264 20432 288
rect 19640 254 19696 264
rect 19732 254 19788 264
rect 19824 254 19880 264
rect 19916 254 19972 264
rect 20008 254 20064 264
rect 20100 254 20156 264
rect 20192 254 20248 264
rect 20284 254 20340 264
rect 20376 254 20432 264
rect 20466 264 20586 288
rect 20620 264 20678 288
rect 20712 264 20770 288
rect 20804 264 20862 288
rect 20896 264 20954 288
rect 20988 264 21046 288
rect 21080 264 21138 288
rect 21172 264 21230 288
rect 21264 264 21322 288
rect 20466 254 20564 264
rect 20620 254 20656 264
rect 20712 254 20748 264
rect 20804 254 20840 264
rect 20896 254 20932 264
rect 20988 254 21024 264
rect 21080 254 21116 264
rect 21172 254 21208 264
rect 21264 254 21300 264
rect 21356 254 21414 288
rect 21448 254 21506 288
rect 21540 254 21598 288
rect 21632 254 21690 288
rect 21724 254 21782 288
rect 21816 254 21874 288
rect 21908 254 21966 288
rect 22000 264 22058 288
rect 22092 264 22150 288
rect 22184 264 22242 288
rect 22276 264 22334 288
rect 22368 264 22426 288
rect 22460 264 22518 288
rect 22552 264 22610 288
rect 22644 264 22702 288
rect 22736 264 22794 288
rect 22030 254 22058 264
rect 22122 254 22150 264
rect 22214 254 22242 264
rect 22306 254 22334 264
rect 22398 254 22426 264
rect 22490 254 22518 264
rect 22582 254 22610 264
rect 22674 254 22702 264
rect 22766 254 22794 264
rect 22828 254 22886 288
rect 22920 264 22978 288
rect 23012 264 23070 288
rect 23104 264 23162 288
rect 23196 264 23254 288
rect 23288 264 23346 288
rect 23380 264 23438 288
rect 23472 264 23530 288
rect 23564 264 23622 288
rect 23656 264 23714 288
rect 22920 254 22956 264
rect 23012 254 23048 264
rect 23104 254 23140 264
rect 23196 254 23232 264
rect 23288 254 23324 264
rect 23380 254 23416 264
rect 23472 254 23508 264
rect 23564 254 23600 264
rect 23656 254 23692 264
rect 23748 254 23806 288
rect 23840 254 23898 288
rect 23932 254 23990 288
rect 24024 254 24082 288
rect 24116 254 24174 288
rect 24208 254 24266 288
rect 24300 254 24358 288
rect 24392 264 24450 288
rect 24484 264 24542 288
rect 24576 264 24634 288
rect 24668 264 24726 288
rect 24760 264 24818 288
rect 24852 264 24910 288
rect 24944 264 25002 288
rect 25036 264 25094 288
rect 25128 264 25189 288
rect 24424 254 24450 264
rect 24516 254 24542 264
rect 24608 254 24634 264
rect 24700 254 24726 264
rect 24792 254 24818 264
rect 24884 254 24910 264
rect 24976 254 25002 264
rect 25068 254 25094 264
rect 18942 239 19606 254
rect 18942 230 18971 239
rect 19577 230 19606 239
rect 19640 230 19698 254
rect 19732 230 19790 254
rect 19824 230 19882 254
rect 19916 230 19974 254
rect 20008 230 20066 254
rect 20100 230 20158 254
rect 20192 230 20250 254
rect 20284 230 20342 254
rect 20376 239 20564 254
rect 20376 230 20405 239
rect 20535 230 20564 239
rect 20598 230 20656 254
rect 20690 230 20748 254
rect 20782 230 20840 254
rect 20874 230 20932 254
rect 20966 230 21024 254
rect 21058 230 21116 254
rect 21150 230 21208 254
rect 21242 230 21300 254
rect 21334 239 21996 254
rect 21334 230 21363 239
rect 21967 230 21996 239
rect 22030 230 22088 254
rect 22122 230 22180 254
rect 22214 230 22272 254
rect 22306 230 22364 254
rect 22398 230 22456 254
rect 22490 230 22548 254
rect 22582 230 22640 254
rect 22674 230 22732 254
rect 22766 239 22956 254
rect 22766 230 22795 239
rect 22927 230 22956 239
rect 22990 230 23048 254
rect 23082 230 23140 254
rect 23174 230 23232 254
rect 23266 230 23324 254
rect 23358 230 23416 254
rect 23450 230 23508 254
rect 23542 230 23600 254
rect 23634 230 23692 254
rect 23726 239 24390 254
rect 23726 230 23755 239
rect 24361 230 24390 239
rect 24424 230 24482 254
rect 24516 230 24574 254
rect 24608 230 24666 254
rect 24700 230 24758 254
rect 24792 230 24850 254
rect 24884 230 24942 254
rect 24976 230 25034 254
rect 25068 230 25126 254
rect 25160 230 25189 264
rect 8593 188 8660 196
rect 8593 154 8610 188
rect 8644 154 8660 188
rect 8593 120 8660 154
rect 8593 86 8610 120
rect 8644 86 8660 120
rect 8593 52 8660 86
rect 8593 18 8610 52
rect 8644 18 8660 52
rect 8593 2 8660 18
rect 8694 188 8728 230
rect 8694 120 8728 154
rect 8694 52 8728 86
rect 8694 2 8728 18
rect 8762 162 9168 196
rect 8593 -132 8627 2
rect 8762 -32 8796 162
rect 8661 -48 8712 -32
rect 8695 -82 8712 -48
rect 8661 -98 8712 -82
rect 8757 -48 8796 -32
rect 8791 -82 8796 -48
rect 8757 -98 8796 -82
rect 8830 94 8930 128
rect 8964 94 9005 128
rect 9039 94 9055 128
rect 8678 -132 8712 -98
rect 8830 -132 8864 94
rect 8593 -159 8644 -132
rect 8593 -193 8603 -159
rect 8637 -185 8644 -159
rect 8678 -166 8864 -132
rect 8898 42 9100 60
rect 8898 26 9059 42
rect 9093 29 9100 42
rect 8898 -84 8932 26
rect 9062 -5 9066 8
rect 8898 -134 8932 -118
rect 8973 -84 9028 -14
rect 8973 -118 8994 -84
rect 8593 -219 8610 -193
rect 8829 -173 8864 -166
rect 8829 -189 8935 -173
rect 8593 -246 8644 -219
rect 8678 -204 8744 -200
rect 8678 -238 8694 -204
rect 8728 -238 8744 -204
rect 8678 -280 8744 -238
rect 8829 -223 8901 -189
rect 8829 -246 8935 -223
rect 8973 -280 9028 -118
rect 9062 -246 9100 -5
rect 9134 29 9168 162
rect 9202 128 9236 230
rect 9202 78 9236 94
rect 9283 128 9386 160
rect 9283 94 9288 128
rect 9322 94 9386 128
rect 9283 78 9386 94
rect 9134 26 9234 29
rect 9134 -8 9231 26
rect 9268 -5 9284 29
rect 9265 -8 9284 -5
rect 9134 -9 9284 -8
rect 9318 -84 9386 78
rect 9140 -118 9156 -84
rect 9190 -118 9386 -84
rect 10026 128 10129 160
rect 10026 94 10090 128
rect 10124 94 10129 128
rect 10026 78 10129 94
rect 10176 128 10210 230
rect 10176 78 10210 94
rect 10244 162 10650 196
rect 10026 -84 10094 78
rect 10244 29 10278 162
rect 10357 94 10373 128
rect 10407 94 10448 128
rect 10482 94 10582 128
rect 10128 27 10144 29
rect 10128 -7 10141 27
rect 10178 -5 10278 29
rect 10175 -7 10278 -5
rect 10128 -9 10278 -7
rect 10312 42 10514 60
rect 10312 29 10321 42
rect 10355 26 10514 42
rect 10346 -5 10350 8
rect 10026 -118 10222 -84
rect 10256 -118 10272 -84
rect 9136 -189 9238 -173
rect 9170 -223 9204 -189
rect 9136 -280 9238 -223
rect 9282 -189 9331 -118
rect 9282 -223 9288 -189
rect 9322 -223 9331 -189
rect 9282 -239 9331 -223
rect 10081 -189 10130 -118
rect 10081 -223 10090 -189
rect 10124 -223 10130 -189
rect 10081 -239 10130 -223
rect 10174 -189 10276 -173
rect 10208 -223 10242 -189
rect 10174 -280 10276 -223
rect 10312 -246 10350 -5
rect 10384 -84 10439 -14
rect 10418 -118 10439 -84
rect 10384 -280 10439 -118
rect 10480 -84 10514 26
rect 10480 -134 10514 -118
rect 10548 -132 10582 94
rect 10616 -32 10650 162
rect 10684 188 10718 230
rect 10684 120 10718 154
rect 10684 52 10718 86
rect 10684 2 10718 18
rect 10752 188 10819 196
rect 10752 154 10768 188
rect 10802 154 10819 188
rect 10752 120 10819 154
rect 10752 86 10768 120
rect 10802 86 10819 120
rect 10752 52 10819 86
rect 10752 18 10768 52
rect 10802 18 10819 52
rect 10752 2 10819 18
rect 10616 -48 10655 -32
rect 10616 -82 10621 -48
rect 10616 -98 10655 -82
rect 10700 -48 10751 -32
rect 10700 -82 10717 -48
rect 10700 -98 10751 -82
rect 10700 -132 10734 -98
rect 10785 -132 10819 2
rect 10548 -166 10734 -132
rect 10768 -161 10819 -132
rect 10548 -173 10583 -166
rect 10477 -189 10583 -173
rect 10511 -223 10583 -189
rect 10768 -185 10779 -161
rect 10813 -195 10819 -161
rect 10477 -246 10583 -223
rect 10668 -204 10734 -200
rect 10668 -238 10684 -204
rect 10718 -238 10734 -204
rect 10668 -280 10734 -238
rect 10802 -219 10819 -195
rect 10768 -246 10819 -219
rect 10985 188 11052 196
rect 10985 154 11002 188
rect 11036 154 11052 188
rect 10985 120 11052 154
rect 10985 86 11002 120
rect 11036 86 11052 120
rect 10985 52 11052 86
rect 10985 18 11002 52
rect 11036 18 11052 52
rect 10985 2 11052 18
rect 11086 188 11120 230
rect 11086 120 11120 154
rect 11086 52 11120 86
rect 11086 2 11120 18
rect 11154 162 11560 196
rect 10985 -132 11019 2
rect 11154 -32 11188 162
rect 11053 -48 11104 -32
rect 11087 -82 11104 -48
rect 11053 -98 11104 -82
rect 11149 -48 11188 -32
rect 11183 -82 11188 -48
rect 11149 -98 11188 -82
rect 11222 94 11322 128
rect 11356 94 11397 128
rect 11431 94 11447 128
rect 11070 -132 11104 -98
rect 11222 -132 11256 94
rect 10985 -159 11036 -132
rect 10985 -193 10995 -159
rect 11029 -185 11036 -159
rect 11070 -166 11256 -132
rect 11290 41 11492 60
rect 11290 26 11452 41
rect 11486 29 11492 41
rect 11290 -84 11324 26
rect 11454 -5 11458 7
rect 11290 -134 11324 -118
rect 11365 -84 11420 -14
rect 11365 -118 11386 -84
rect 10985 -219 11002 -193
rect 11221 -173 11256 -166
rect 11221 -189 11327 -173
rect 10985 -246 11036 -219
rect 11070 -204 11136 -200
rect 11070 -238 11086 -204
rect 11120 -238 11136 -204
rect 11070 -280 11136 -238
rect 11221 -223 11293 -189
rect 11221 -246 11327 -223
rect 11365 -280 11420 -118
rect 11454 -246 11492 -5
rect 11526 29 11560 162
rect 11594 128 11628 230
rect 11594 78 11628 94
rect 11675 128 11778 160
rect 11675 94 11680 128
rect 11714 94 11778 128
rect 11675 78 11778 94
rect 11526 25 11626 29
rect 11526 -9 11623 25
rect 11660 -5 11676 29
rect 11657 -9 11676 -5
rect 11710 -84 11778 78
rect 11532 -118 11548 -84
rect 11582 -118 11778 -84
rect 12418 128 12521 160
rect 12418 94 12482 128
rect 12516 94 12521 128
rect 12418 78 12521 94
rect 12568 128 12602 230
rect 12568 78 12602 94
rect 12636 162 13042 196
rect 12418 -84 12486 78
rect 12636 29 12670 162
rect 12749 94 12765 128
rect 12799 94 12840 128
rect 12874 94 12974 128
rect 12520 26 12536 29
rect 12520 -8 12533 26
rect 12570 -5 12670 29
rect 12567 -8 12670 -5
rect 12520 -9 12670 -8
rect 12704 42 12906 60
rect 12704 29 12713 42
rect 12747 26 12906 42
rect 12738 -5 12742 8
rect 12418 -118 12614 -84
rect 12648 -118 12664 -84
rect 11528 -189 11630 -173
rect 11562 -223 11596 -189
rect 11528 -280 11630 -223
rect 11674 -189 11723 -118
rect 11674 -223 11680 -189
rect 11714 -223 11723 -189
rect 11674 -239 11723 -223
rect 12473 -189 12522 -118
rect 12473 -223 12482 -189
rect 12516 -223 12522 -189
rect 12473 -239 12522 -223
rect 12566 -189 12668 -173
rect 12600 -223 12634 -189
rect 12566 -280 12668 -223
rect 12704 -246 12742 -5
rect 12776 -84 12831 -14
rect 12810 -118 12831 -84
rect 12776 -280 12831 -118
rect 12872 -84 12906 26
rect 12872 -134 12906 -118
rect 12940 -132 12974 94
rect 13008 -32 13042 162
rect 13076 188 13110 230
rect 13076 120 13110 154
rect 13076 52 13110 86
rect 13076 2 13110 18
rect 13144 188 13211 196
rect 13144 154 13160 188
rect 13194 154 13211 188
rect 13144 120 13211 154
rect 13144 86 13160 120
rect 13194 86 13211 120
rect 13144 52 13211 86
rect 13144 18 13160 52
rect 13194 18 13211 52
rect 13144 2 13211 18
rect 13008 -48 13047 -32
rect 13008 -82 13013 -48
rect 13008 -98 13047 -82
rect 13092 -48 13143 -32
rect 13092 -82 13109 -48
rect 13092 -98 13143 -82
rect 13092 -132 13126 -98
rect 13177 -132 13211 2
rect 12940 -166 13126 -132
rect 13160 -161 13211 -132
rect 12940 -173 12975 -166
rect 12869 -189 12975 -173
rect 12903 -223 12975 -189
rect 13160 -185 13173 -161
rect 13207 -195 13211 -161
rect 12869 -246 12975 -223
rect 13060 -204 13126 -200
rect 13060 -238 13076 -204
rect 13110 -238 13126 -204
rect 13060 -280 13126 -238
rect 13194 -219 13211 -195
rect 13160 -246 13211 -219
rect 13377 188 13444 196
rect 13377 154 13394 188
rect 13428 154 13444 188
rect 13377 120 13444 154
rect 13377 86 13394 120
rect 13428 86 13444 120
rect 13377 52 13444 86
rect 13377 18 13394 52
rect 13428 18 13444 52
rect 13377 2 13444 18
rect 13478 188 13512 230
rect 13478 120 13512 154
rect 13478 52 13512 86
rect 13478 2 13512 18
rect 13546 162 13952 196
rect 13377 -132 13411 2
rect 13546 -32 13580 162
rect 13445 -48 13496 -32
rect 13479 -82 13496 -48
rect 13445 -98 13496 -82
rect 13541 -48 13580 -32
rect 13575 -82 13580 -48
rect 13541 -98 13580 -82
rect 13614 94 13714 128
rect 13748 94 13789 128
rect 13823 94 13839 128
rect 13462 -132 13496 -98
rect 13614 -132 13648 94
rect 13377 -159 13428 -132
rect 13377 -193 13387 -159
rect 13421 -185 13428 -159
rect 13462 -166 13648 -132
rect 13682 41 13884 60
rect 13682 26 13844 41
rect 13878 29 13884 41
rect 13682 -84 13716 26
rect 13846 -5 13850 7
rect 13682 -134 13716 -118
rect 13757 -84 13812 -14
rect 13757 -118 13778 -84
rect 13377 -219 13394 -193
rect 13613 -173 13648 -166
rect 13613 -189 13719 -173
rect 13377 -246 13428 -219
rect 13462 -204 13528 -200
rect 13462 -238 13478 -204
rect 13512 -238 13528 -204
rect 13462 -280 13528 -238
rect 13613 -223 13685 -189
rect 13613 -246 13719 -223
rect 13757 -280 13812 -118
rect 13846 -246 13884 -5
rect 13918 29 13952 162
rect 13986 128 14020 230
rect 13986 78 14020 94
rect 14067 128 14170 160
rect 14067 94 14072 128
rect 14106 94 14170 128
rect 14067 78 14170 94
rect 13918 26 14018 29
rect 13918 -8 14014 26
rect 14052 -5 14068 29
rect 14048 -8 14068 -5
rect 13918 -9 14068 -8
rect 14102 -84 14170 78
rect 13924 -118 13940 -84
rect 13974 -118 14170 -84
rect 14808 128 14911 160
rect 14808 94 14872 128
rect 14906 94 14911 128
rect 14808 78 14911 94
rect 14958 128 14992 230
rect 14958 78 14992 94
rect 15026 162 15432 196
rect 14808 -84 14876 78
rect 15026 29 15060 162
rect 15139 94 15155 128
rect 15189 94 15230 128
rect 15264 94 15364 128
rect 14910 26 14926 29
rect 14910 -8 14923 26
rect 14960 -5 15060 29
rect 14957 -8 15060 -5
rect 14910 -9 15060 -8
rect 15094 43 15296 60
rect 15094 29 15104 43
rect 15138 26 15296 43
rect 15128 -5 15132 9
rect 14808 -118 15004 -84
rect 15038 -118 15054 -84
rect 13920 -189 14022 -173
rect 13954 -223 13988 -189
rect 13920 -280 14022 -223
rect 14066 -189 14115 -118
rect 14066 -223 14072 -189
rect 14106 -223 14115 -189
rect 14066 -239 14115 -223
rect 14863 -189 14912 -118
rect 14863 -223 14872 -189
rect 14906 -223 14912 -189
rect 14863 -239 14912 -223
rect 14956 -189 15058 -173
rect 14990 -223 15024 -189
rect 14956 -280 15058 -223
rect 15094 -246 15132 -5
rect 15166 -84 15221 -14
rect 15200 -118 15221 -84
rect 15166 -280 15221 -118
rect 15262 -84 15296 26
rect 15262 -134 15296 -118
rect 15330 -132 15364 94
rect 15398 -32 15432 162
rect 15466 188 15500 230
rect 15466 120 15500 154
rect 15466 52 15500 86
rect 15466 2 15500 18
rect 15534 188 15601 196
rect 15534 154 15550 188
rect 15584 154 15601 188
rect 15534 120 15601 154
rect 15534 86 15550 120
rect 15584 86 15601 120
rect 15534 52 15601 86
rect 15534 18 15550 52
rect 15584 18 15601 52
rect 15534 2 15601 18
rect 15398 -48 15437 -32
rect 15398 -82 15403 -48
rect 15398 -98 15437 -82
rect 15482 -48 15533 -32
rect 15482 -82 15499 -48
rect 15482 -98 15533 -82
rect 15482 -132 15516 -98
rect 15567 -132 15601 2
rect 15330 -166 15516 -132
rect 15550 -159 15601 -132
rect 15330 -173 15365 -166
rect 15259 -189 15365 -173
rect 15293 -223 15365 -189
rect 15550 -185 15563 -159
rect 15597 -193 15601 -159
rect 15259 -246 15365 -223
rect 15450 -204 15516 -200
rect 15450 -238 15466 -204
rect 15500 -238 15516 -204
rect 15450 -280 15516 -238
rect 15584 -219 15601 -193
rect 15550 -246 15601 -219
rect 15769 188 15836 196
rect 15769 154 15786 188
rect 15820 154 15836 188
rect 15769 120 15836 154
rect 15769 86 15786 120
rect 15820 86 15836 120
rect 15769 52 15836 86
rect 15769 18 15786 52
rect 15820 18 15836 52
rect 15769 2 15836 18
rect 15870 188 15904 230
rect 15870 120 15904 154
rect 15870 52 15904 86
rect 15870 2 15904 18
rect 15938 162 16344 196
rect 15769 -132 15803 2
rect 15938 -32 15972 162
rect 15837 -48 15888 -32
rect 15871 -82 15888 -48
rect 15837 -98 15888 -82
rect 15933 -48 15972 -32
rect 15967 -82 15972 -48
rect 15933 -98 15972 -82
rect 16006 94 16106 128
rect 16140 94 16181 128
rect 16215 94 16231 128
rect 15854 -132 15888 -98
rect 16006 -132 16040 94
rect 15769 -159 15820 -132
rect 15769 -193 15779 -159
rect 15813 -185 15820 -159
rect 15854 -166 16040 -132
rect 16074 42 16276 60
rect 16074 26 16236 42
rect 16270 29 16276 42
rect 16074 -84 16108 26
rect 16238 -5 16242 8
rect 16074 -134 16108 -118
rect 16149 -84 16204 -14
rect 16149 -118 16170 -84
rect 15769 -219 15786 -193
rect 16005 -173 16040 -166
rect 16005 -189 16111 -173
rect 15769 -246 15820 -219
rect 15854 -204 15920 -200
rect 15854 -238 15870 -204
rect 15904 -238 15920 -204
rect 15854 -280 15920 -238
rect 16005 -223 16077 -189
rect 16005 -246 16111 -223
rect 16149 -280 16204 -118
rect 16238 -246 16276 -5
rect 16310 29 16344 162
rect 16378 128 16412 230
rect 16378 78 16412 94
rect 16459 128 16562 160
rect 16459 94 16464 128
rect 16498 94 16562 128
rect 16459 78 16562 94
rect 16310 26 16410 29
rect 16310 -8 16407 26
rect 16444 -5 16460 29
rect 16441 -8 16460 -5
rect 16310 -9 16460 -8
rect 16494 -84 16562 78
rect 16316 -118 16332 -84
rect 16366 -118 16562 -84
rect 17202 128 17305 160
rect 17202 94 17266 128
rect 17300 94 17305 128
rect 17202 78 17305 94
rect 17352 128 17386 230
rect 17352 78 17386 94
rect 17420 162 17826 196
rect 17202 -84 17270 78
rect 17420 29 17454 162
rect 17533 94 17549 128
rect 17583 94 17624 128
rect 17658 94 17758 128
rect 17304 27 17320 29
rect 17304 -7 17317 27
rect 17354 -5 17454 29
rect 17351 -7 17454 -5
rect 17304 -9 17454 -7
rect 17488 43 17690 60
rect 17488 29 17497 43
rect 17531 26 17690 43
rect 17522 -5 17526 9
rect 17202 -118 17398 -84
rect 17432 -118 17448 -84
rect 16312 -189 16414 -173
rect 16346 -223 16380 -189
rect 16312 -280 16414 -223
rect 16458 -189 16507 -118
rect 16458 -223 16464 -189
rect 16498 -223 16507 -189
rect 16458 -239 16507 -223
rect 17257 -189 17306 -118
rect 17257 -223 17266 -189
rect 17300 -223 17306 -189
rect 17257 -239 17306 -223
rect 17350 -189 17452 -173
rect 17384 -223 17418 -189
rect 17350 -280 17452 -223
rect 17488 -246 17526 -5
rect 17560 -84 17615 -14
rect 17594 -118 17615 -84
rect 17560 -280 17615 -118
rect 17656 -84 17690 26
rect 17656 -134 17690 -118
rect 17724 -132 17758 94
rect 17792 -32 17826 162
rect 17860 188 17894 230
rect 17860 120 17894 154
rect 17860 52 17894 86
rect 17860 2 17894 18
rect 17928 188 17995 196
rect 17928 154 17944 188
rect 17978 154 17995 188
rect 17928 120 17995 154
rect 17928 86 17944 120
rect 17978 86 17995 120
rect 17928 52 17995 86
rect 17928 18 17944 52
rect 17978 18 17995 52
rect 17928 2 17995 18
rect 17792 -48 17831 -32
rect 17792 -82 17797 -48
rect 17792 -98 17831 -82
rect 17876 -48 17927 -32
rect 17876 -82 17893 -48
rect 17876 -98 17927 -82
rect 17876 -132 17910 -98
rect 17961 -132 17995 2
rect 17724 -166 17910 -132
rect 17944 -161 17995 -132
rect 17724 -173 17759 -166
rect 17653 -189 17759 -173
rect 17687 -223 17759 -189
rect 17944 -185 17955 -161
rect 17989 -195 17995 -161
rect 17653 -246 17759 -223
rect 17844 -204 17910 -200
rect 17844 -238 17860 -204
rect 17894 -238 17910 -204
rect 17844 -280 17910 -238
rect 17978 -219 17995 -195
rect 17944 -246 17995 -219
rect 18161 188 18228 196
rect 18161 154 18178 188
rect 18212 154 18228 188
rect 18161 120 18228 154
rect 18161 86 18178 120
rect 18212 86 18228 120
rect 18161 52 18228 86
rect 18161 18 18178 52
rect 18212 18 18228 52
rect 18161 2 18228 18
rect 18262 188 18296 230
rect 18262 120 18296 154
rect 18262 52 18296 86
rect 18262 2 18296 18
rect 18330 162 18736 196
rect 18161 -132 18195 2
rect 18330 -32 18364 162
rect 18229 -48 18280 -32
rect 18263 -82 18280 -48
rect 18229 -98 18280 -82
rect 18325 -48 18364 -32
rect 18359 -82 18364 -48
rect 18325 -98 18364 -82
rect 18398 94 18498 128
rect 18532 94 18573 128
rect 18607 94 18623 128
rect 18246 -132 18280 -98
rect 18398 -132 18432 94
rect 18161 -158 18212 -132
rect 18161 -192 18170 -158
rect 18204 -185 18212 -158
rect 18246 -166 18432 -132
rect 18466 41 18668 60
rect 18466 26 18627 41
rect 18661 29 18668 41
rect 18466 -84 18500 26
rect 18630 -5 18634 7
rect 18466 -134 18500 -118
rect 18541 -84 18596 -14
rect 18541 -118 18562 -84
rect 18161 -219 18178 -192
rect 18397 -173 18432 -166
rect 18397 -189 18503 -173
rect 18161 -246 18212 -219
rect 18246 -204 18312 -200
rect 18246 -238 18262 -204
rect 18296 -238 18312 -204
rect 18246 -280 18312 -238
rect 18397 -223 18469 -189
rect 18397 -246 18503 -223
rect 18541 -280 18596 -118
rect 18630 -246 18668 -5
rect 18702 29 18736 162
rect 18770 128 18804 230
rect 18770 78 18804 94
rect 18851 128 18954 160
rect 18851 94 18856 128
rect 18890 94 18954 128
rect 18851 78 18954 94
rect 18702 27 18802 29
rect 18702 -7 18798 27
rect 18836 -5 18852 29
rect 18832 -7 18852 -5
rect 18702 -9 18852 -7
rect 18886 -84 18954 78
rect 18708 -118 18724 -84
rect 18758 -118 18954 -84
rect 19594 128 19697 160
rect 19594 94 19658 128
rect 19692 94 19697 128
rect 19594 78 19697 94
rect 19744 128 19778 230
rect 19744 78 19778 94
rect 19812 162 20218 196
rect 19594 -84 19662 78
rect 19812 29 19846 162
rect 19925 94 19941 128
rect 19975 94 20016 128
rect 20050 94 20150 128
rect 19696 26 19712 29
rect 19696 -8 19709 26
rect 19746 -5 19846 29
rect 19743 -8 19846 -5
rect 19696 -9 19846 -8
rect 19880 43 20082 60
rect 19880 29 19890 43
rect 19924 26 20082 43
rect 19914 -5 19918 9
rect 19594 -118 19790 -84
rect 19824 -118 19840 -84
rect 18704 -189 18806 -173
rect 18738 -223 18772 -189
rect 18704 -280 18806 -223
rect 18850 -189 18899 -118
rect 18850 -223 18856 -189
rect 18890 -223 18899 -189
rect 18850 -239 18899 -223
rect 19649 -189 19698 -118
rect 19649 -223 19658 -189
rect 19692 -223 19698 -189
rect 19649 -239 19698 -223
rect 19742 -189 19844 -173
rect 19776 -223 19810 -189
rect 19742 -280 19844 -223
rect 19880 -246 19918 -5
rect 19952 -84 20007 -14
rect 19986 -118 20007 -84
rect 19952 -280 20007 -118
rect 20048 -84 20082 26
rect 20048 -134 20082 -118
rect 20116 -132 20150 94
rect 20184 -32 20218 162
rect 20252 188 20286 230
rect 20252 120 20286 154
rect 20252 52 20286 86
rect 20252 2 20286 18
rect 20320 188 20387 196
rect 20320 154 20336 188
rect 20370 154 20387 188
rect 20320 120 20387 154
rect 20320 86 20336 120
rect 20370 86 20387 120
rect 20320 52 20387 86
rect 20320 18 20336 52
rect 20370 18 20387 52
rect 20320 2 20387 18
rect 20184 -48 20223 -32
rect 20184 -82 20189 -48
rect 20184 -98 20223 -82
rect 20268 -48 20319 -32
rect 20268 -82 20285 -48
rect 20268 -98 20319 -82
rect 20268 -132 20302 -98
rect 20353 -132 20387 2
rect 20116 -166 20302 -132
rect 20336 -159 20387 -132
rect 20116 -173 20151 -166
rect 20045 -189 20151 -173
rect 20079 -223 20151 -189
rect 20336 -185 20347 -159
rect 20381 -193 20387 -159
rect 20045 -246 20151 -223
rect 20236 -204 20302 -200
rect 20236 -238 20252 -204
rect 20286 -238 20302 -204
rect 20236 -280 20302 -238
rect 20370 -219 20387 -193
rect 20336 -246 20387 -219
rect 20553 188 20620 196
rect 20553 154 20570 188
rect 20604 154 20620 188
rect 20553 120 20620 154
rect 20553 86 20570 120
rect 20604 86 20620 120
rect 20553 52 20620 86
rect 20553 18 20570 52
rect 20604 18 20620 52
rect 20553 2 20620 18
rect 20654 188 20688 230
rect 20654 120 20688 154
rect 20654 52 20688 86
rect 20654 2 20688 18
rect 20722 162 21128 196
rect 20553 -132 20587 2
rect 20722 -32 20756 162
rect 20621 -48 20672 -32
rect 20655 -82 20672 -48
rect 20621 -98 20672 -82
rect 20717 -48 20756 -32
rect 20751 -82 20756 -48
rect 20717 -98 20756 -82
rect 20790 94 20890 128
rect 20924 94 20965 128
rect 20999 94 21015 128
rect 20638 -132 20672 -98
rect 20790 -132 20824 94
rect 20553 -159 20604 -132
rect 20553 -193 20562 -159
rect 20596 -185 20604 -159
rect 20638 -166 20824 -132
rect 20858 40 21060 60
rect 20858 26 21019 40
rect 21053 29 21060 40
rect 20858 -84 20892 26
rect 21022 -5 21026 6
rect 20858 -134 20892 -118
rect 20933 -84 20988 -14
rect 20933 -118 20954 -84
rect 20553 -219 20570 -193
rect 20789 -173 20824 -166
rect 20789 -189 20895 -173
rect 20553 -246 20604 -219
rect 20638 -204 20704 -200
rect 20638 -238 20654 -204
rect 20688 -238 20704 -204
rect 20638 -280 20704 -238
rect 20789 -223 20861 -189
rect 20789 -246 20895 -223
rect 20933 -280 20988 -118
rect 21022 -246 21060 -5
rect 21094 29 21128 162
rect 21162 128 21196 230
rect 21162 78 21196 94
rect 21243 128 21346 160
rect 21243 94 21248 128
rect 21282 94 21346 128
rect 21243 78 21346 94
rect 21094 27 21194 29
rect 21094 -7 21190 27
rect 21228 -5 21244 29
rect 21224 -7 21244 -5
rect 21094 -9 21244 -7
rect 21278 -84 21346 78
rect 21100 -118 21116 -84
rect 21150 -118 21346 -84
rect 21984 128 22087 160
rect 21984 94 22048 128
rect 22082 94 22087 128
rect 21984 78 22087 94
rect 22134 128 22168 230
rect 22134 78 22168 94
rect 22202 162 22608 196
rect 21984 -84 22052 78
rect 22202 29 22236 162
rect 22315 94 22331 128
rect 22365 94 22406 128
rect 22440 94 22540 128
rect 22086 26 22102 29
rect 22086 -8 22098 26
rect 22136 -5 22236 29
rect 22132 -8 22236 -5
rect 22086 -9 22236 -8
rect 22270 43 22472 60
rect 22270 29 22279 43
rect 22313 26 22472 43
rect 22304 -5 22308 9
rect 21984 -118 22180 -84
rect 22214 -118 22230 -84
rect 21096 -189 21198 -173
rect 21130 -223 21164 -189
rect 21096 -280 21198 -223
rect 21242 -189 21291 -118
rect 21242 -223 21248 -189
rect 21282 -223 21291 -189
rect 21242 -239 21291 -223
rect 22039 -189 22088 -118
rect 22039 -223 22048 -189
rect 22082 -223 22088 -189
rect 22039 -239 22088 -223
rect 22132 -189 22234 -173
rect 22166 -223 22200 -189
rect 22132 -280 22234 -223
rect 22270 -246 22308 -5
rect 22342 -84 22397 -14
rect 22376 -118 22397 -84
rect 22342 -280 22397 -118
rect 22438 -84 22472 26
rect 22438 -134 22472 -118
rect 22506 -132 22540 94
rect 22574 -32 22608 162
rect 22642 188 22676 230
rect 22642 120 22676 154
rect 22642 52 22676 86
rect 22642 2 22676 18
rect 22710 188 22777 196
rect 22710 154 22726 188
rect 22760 154 22777 188
rect 22710 120 22777 154
rect 22710 86 22726 120
rect 22760 86 22777 120
rect 22710 52 22777 86
rect 22710 18 22726 52
rect 22760 18 22777 52
rect 22710 2 22777 18
rect 22574 -48 22613 -32
rect 22574 -82 22579 -48
rect 22574 -98 22613 -82
rect 22658 -48 22709 -32
rect 22658 -82 22675 -48
rect 22658 -98 22709 -82
rect 22658 -132 22692 -98
rect 22743 -132 22777 2
rect 22506 -166 22692 -132
rect 22726 -161 22777 -132
rect 22506 -173 22541 -166
rect 22435 -189 22541 -173
rect 22469 -223 22541 -189
rect 22726 -185 22739 -161
rect 22773 -195 22777 -161
rect 22435 -246 22541 -223
rect 22626 -204 22692 -200
rect 22626 -238 22642 -204
rect 22676 -238 22692 -204
rect 22626 -280 22692 -238
rect 22760 -219 22777 -195
rect 22726 -246 22777 -219
rect 22945 188 23012 196
rect 22945 154 22962 188
rect 22996 154 23012 188
rect 22945 120 23012 154
rect 22945 86 22962 120
rect 22996 86 23012 120
rect 22945 52 23012 86
rect 22945 18 22962 52
rect 22996 18 23012 52
rect 22945 2 23012 18
rect 23046 188 23080 230
rect 23046 120 23080 154
rect 23046 52 23080 86
rect 23046 2 23080 18
rect 23114 162 23520 196
rect 22945 -132 22979 2
rect 23114 -32 23148 162
rect 23013 -48 23064 -32
rect 23047 -82 23064 -48
rect 23013 -98 23064 -82
rect 23109 -48 23148 -32
rect 23143 -82 23148 -48
rect 23109 -98 23148 -82
rect 23182 94 23282 128
rect 23316 94 23357 128
rect 23391 94 23407 128
rect 23030 -132 23064 -98
rect 23182 -132 23216 94
rect 22945 -158 22996 -132
rect 22945 -192 22955 -158
rect 22989 -185 22996 -158
rect 23030 -166 23216 -132
rect 23250 41 23452 60
rect 23250 26 23411 41
rect 23445 29 23452 41
rect 23250 -84 23284 26
rect 23414 -5 23418 7
rect 23250 -134 23284 -118
rect 23325 -84 23380 -14
rect 23325 -118 23346 -84
rect 22945 -219 22962 -192
rect 23181 -173 23216 -166
rect 23181 -189 23287 -173
rect 22945 -246 22996 -219
rect 23030 -204 23096 -200
rect 23030 -238 23046 -204
rect 23080 -238 23096 -204
rect 23030 -280 23096 -238
rect 23181 -223 23253 -189
rect 23181 -246 23287 -223
rect 23325 -280 23380 -118
rect 23414 -246 23452 -5
rect 23486 29 23520 162
rect 23554 128 23588 230
rect 23554 78 23588 94
rect 23635 128 23738 160
rect 23635 94 23640 128
rect 23674 94 23738 128
rect 23635 78 23738 94
rect 23486 27 23586 29
rect 23486 -7 23583 27
rect 23620 -5 23636 29
rect 23617 -7 23636 -5
rect 23486 -9 23636 -7
rect 23670 -84 23738 78
rect 23492 -118 23508 -84
rect 23542 -118 23738 -84
rect 24378 128 24481 160
rect 24378 94 24442 128
rect 24476 94 24481 128
rect 24378 78 24481 94
rect 24528 128 24562 230
rect 24528 78 24562 94
rect 24596 162 25002 196
rect 24378 -84 24446 78
rect 24596 29 24630 162
rect 24709 94 24725 128
rect 24759 94 24800 128
rect 24834 94 24934 128
rect 24480 27 24496 29
rect 24480 -7 24493 27
rect 24530 -5 24630 29
rect 24527 -7 24630 -5
rect 24480 -9 24630 -7
rect 24664 43 24866 60
rect 24664 29 24674 43
rect 24708 26 24866 43
rect 24698 -5 24702 9
rect 24378 -118 24574 -84
rect 24608 -118 24624 -84
rect 23488 -189 23590 -173
rect 23522 -223 23556 -189
rect 23488 -280 23590 -223
rect 23634 -189 23683 -118
rect 23634 -223 23640 -189
rect 23674 -223 23683 -189
rect 23634 -239 23683 -223
rect 24433 -189 24482 -118
rect 24433 -223 24442 -189
rect 24476 -223 24482 -189
rect 24433 -239 24482 -223
rect 24526 -189 24628 -173
rect 24560 -223 24594 -189
rect 24526 -280 24628 -223
rect 24664 -246 24702 -5
rect 24736 -84 24791 -14
rect 24770 -118 24791 -84
rect 24736 -280 24791 -118
rect 24832 -84 24866 26
rect 24832 -134 24866 -118
rect 24900 -132 24934 94
rect 24968 -32 25002 162
rect 25036 188 25070 230
rect 25036 120 25070 154
rect 25036 52 25070 86
rect 25036 2 25070 18
rect 25104 188 25171 196
rect 25104 154 25120 188
rect 25154 154 25171 188
rect 25104 120 25171 154
rect 25104 86 25120 120
rect 25154 86 25171 120
rect 25104 52 25171 86
rect 25104 18 25120 52
rect 25154 18 25171 52
rect 25104 2 25171 18
rect 24968 -48 25007 -32
rect 24968 -82 24973 -48
rect 24968 -98 25007 -82
rect 25052 -48 25103 -32
rect 25052 -82 25069 -48
rect 25052 -98 25103 -82
rect 25052 -132 25086 -98
rect 25137 -132 25171 2
rect 24900 -166 25086 -132
rect 25120 -159 25171 -132
rect 24900 -173 24935 -166
rect 24829 -189 24935 -173
rect 24863 -223 24935 -189
rect 25120 -185 25131 -159
rect 25165 -193 25171 -159
rect 24829 -246 24935 -223
rect 25020 -204 25086 -200
rect 25020 -238 25036 -204
rect 25070 -238 25086 -204
rect 25020 -280 25086 -238
rect 25154 -219 25171 -193
rect 25120 -246 25171 -219
rect 8575 -338 8604 -280
rect 8638 -338 8696 -280
rect 8730 -338 8788 -280
rect 8822 -338 8880 -280
rect 8914 -338 8972 -280
rect 9006 -338 9064 -280
rect 9098 -338 9156 -280
rect 9190 -338 9248 -280
rect 9282 -338 9340 -280
rect 9374 -289 9403 -280
rect 10009 -289 10038 -280
rect 9374 -304 10038 -289
rect 9374 -338 9432 -304
rect 9466 -338 9524 -304
rect 9558 -338 9616 -304
rect 9650 -338 9708 -304
rect 9742 -338 9800 -304
rect 9834 -338 9892 -304
rect 9926 -338 9984 -304
rect 10018 -314 10038 -304
rect 10072 -304 10130 -280
rect 10072 -314 10076 -304
rect 10018 -338 10076 -314
rect 10110 -314 10130 -304
rect 10164 -304 10222 -280
rect 10164 -314 10168 -304
rect 10110 -338 10168 -314
rect 10202 -314 10222 -304
rect 10256 -304 10314 -280
rect 10256 -314 10260 -304
rect 10202 -338 10260 -314
rect 10294 -314 10314 -304
rect 10348 -304 10406 -280
rect 10348 -314 10352 -304
rect 10294 -338 10352 -314
rect 10386 -314 10406 -304
rect 10440 -304 10498 -280
rect 10440 -314 10444 -304
rect 10386 -338 10444 -314
rect 10478 -314 10498 -304
rect 10532 -304 10590 -280
rect 10532 -314 10536 -304
rect 10478 -338 10536 -314
rect 10570 -314 10590 -304
rect 10624 -304 10682 -280
rect 10624 -314 10628 -304
rect 10570 -338 10628 -314
rect 10662 -314 10682 -304
rect 10716 -304 10774 -280
rect 10716 -314 10720 -304
rect 10662 -338 10720 -314
rect 10754 -314 10774 -304
rect 10808 -289 10837 -280
rect 10967 -289 10996 -280
rect 10808 -304 10996 -289
rect 10808 -314 10812 -304
rect 10754 -338 10812 -314
rect 10846 -338 10904 -304
rect 10938 -338 10996 -304
rect 11030 -338 11088 -280
rect 11122 -338 11180 -280
rect 11214 -338 11272 -280
rect 11306 -338 11364 -280
rect 11398 -338 11456 -280
rect 11490 -338 11548 -280
rect 11582 -338 11640 -280
rect 11674 -338 11732 -280
rect 11766 -289 11795 -280
rect 12401 -289 12430 -280
rect 11766 -304 12430 -289
rect 11766 -338 11824 -304
rect 11858 -338 11916 -304
rect 11950 -338 12008 -304
rect 12042 -338 12100 -304
rect 12134 -338 12192 -304
rect 12226 -338 12284 -304
rect 12318 -338 12376 -304
rect 12410 -314 12430 -304
rect 12464 -304 12522 -280
rect 12464 -314 12468 -304
rect 12410 -338 12468 -314
rect 12502 -314 12522 -304
rect 12556 -304 12614 -280
rect 12556 -314 12560 -304
rect 12502 -338 12560 -314
rect 12594 -314 12614 -304
rect 12648 -304 12706 -280
rect 12648 -314 12652 -304
rect 12594 -338 12652 -314
rect 12686 -314 12706 -304
rect 12740 -304 12798 -280
rect 12740 -314 12744 -304
rect 12686 -338 12744 -314
rect 12778 -314 12798 -304
rect 12832 -304 12890 -280
rect 12832 -314 12836 -304
rect 12778 -338 12836 -314
rect 12870 -314 12890 -304
rect 12924 -304 12982 -280
rect 12924 -314 12928 -304
rect 12870 -338 12928 -314
rect 12962 -314 12982 -304
rect 13016 -304 13074 -280
rect 13016 -314 13020 -304
rect 12962 -338 13020 -314
rect 13054 -314 13074 -304
rect 13108 -304 13166 -280
rect 13108 -314 13112 -304
rect 13054 -338 13112 -314
rect 13146 -314 13166 -304
rect 13200 -289 13229 -280
rect 13359 -289 13388 -280
rect 13200 -304 13388 -289
rect 13200 -314 13204 -304
rect 13146 -338 13204 -314
rect 13238 -338 13296 -304
rect 13330 -338 13388 -304
rect 13422 -338 13480 -280
rect 13514 -338 13572 -280
rect 13606 -338 13664 -280
rect 13698 -338 13756 -280
rect 13790 -338 13848 -280
rect 13882 -338 13940 -280
rect 13974 -338 14032 -280
rect 14066 -338 14124 -280
rect 14158 -289 14187 -280
rect 14791 -289 14820 -280
rect 14158 -304 14820 -289
rect 14158 -338 14216 -304
rect 14250 -338 14820 -304
rect 14854 -338 14912 -280
rect 14946 -338 15004 -280
rect 15038 -338 15096 -280
rect 15130 -338 15188 -280
rect 15222 -338 15280 -280
rect 15314 -338 15372 -280
rect 15406 -338 15464 -280
rect 15498 -338 15556 -280
rect 15590 -289 15619 -280
rect 15751 -289 15780 -280
rect 15590 -304 15780 -289
rect 15590 -338 15648 -304
rect 15682 -338 15740 -304
rect 15774 -314 15780 -304
rect 15814 -304 15872 -280
rect 15814 -314 15832 -304
rect 15774 -338 15832 -314
rect 15866 -314 15872 -304
rect 15906 -304 15964 -280
rect 15906 -314 15924 -304
rect 15866 -338 15924 -314
rect 15958 -314 15964 -304
rect 15998 -304 16056 -280
rect 15998 -314 16016 -304
rect 15958 -338 16016 -314
rect 16050 -314 16056 -304
rect 16090 -304 16148 -280
rect 16090 -314 16108 -304
rect 16050 -338 16108 -314
rect 16142 -314 16148 -304
rect 16182 -304 16240 -280
rect 16182 -314 16200 -304
rect 16142 -338 16200 -314
rect 16234 -314 16240 -304
rect 16274 -304 16332 -280
rect 16274 -314 16292 -304
rect 16234 -338 16292 -314
rect 16326 -314 16332 -304
rect 16366 -304 16424 -280
rect 16366 -314 16384 -304
rect 16326 -338 16384 -314
rect 16418 -314 16424 -304
rect 16458 -304 16516 -280
rect 16458 -314 16476 -304
rect 16418 -338 16476 -314
rect 16510 -314 16516 -304
rect 16550 -289 16579 -280
rect 17185 -289 17214 -280
rect 16550 -304 17214 -289
rect 17248 -304 17306 -280
rect 17340 -304 17398 -280
rect 17432 -304 17490 -280
rect 17524 -304 17582 -280
rect 17616 -304 17674 -280
rect 17708 -304 17766 -280
rect 17800 -304 17858 -280
rect 17892 -304 17950 -280
rect 17984 -289 18013 -280
rect 18143 -289 18172 -280
rect 17984 -304 18172 -289
rect 16550 -314 16568 -304
rect 16510 -338 16568 -314
rect 16602 -338 16660 -304
rect 16694 -338 16752 -304
rect 16786 -338 16844 -304
rect 16878 -338 16936 -304
rect 16970 -338 17028 -304
rect 17062 -338 17120 -304
rect 17154 -338 17212 -304
rect 17248 -314 17304 -304
rect 17340 -314 17396 -304
rect 17432 -314 17488 -304
rect 17524 -314 17580 -304
rect 17616 -314 17672 -304
rect 17708 -314 17764 -304
rect 17800 -314 17856 -304
rect 17892 -314 17948 -304
rect 17984 -314 18040 -304
rect 17246 -338 17304 -314
rect 17338 -338 17396 -314
rect 17430 -338 17488 -314
rect 17522 -338 17580 -314
rect 17614 -338 17672 -314
rect 17706 -338 17764 -314
rect 17798 -338 17856 -314
rect 17890 -338 17948 -314
rect 17982 -338 18040 -314
rect 18074 -338 18132 -304
rect 18166 -314 18172 -304
rect 18206 -304 18264 -280
rect 18206 -314 18224 -304
rect 18166 -338 18224 -314
rect 18258 -314 18264 -304
rect 18298 -304 18356 -280
rect 18298 -314 18316 -304
rect 18258 -338 18316 -314
rect 18350 -314 18356 -304
rect 18390 -304 18448 -280
rect 18390 -314 18408 -304
rect 18350 -338 18408 -314
rect 18442 -314 18448 -304
rect 18482 -304 18540 -280
rect 18482 -314 18500 -304
rect 18442 -338 18500 -314
rect 18534 -314 18540 -304
rect 18574 -304 18632 -280
rect 18574 -314 18592 -304
rect 18534 -338 18592 -314
rect 18626 -314 18632 -304
rect 18666 -304 18724 -280
rect 18666 -314 18684 -304
rect 18626 -338 18684 -314
rect 18718 -314 18724 -304
rect 18758 -304 18816 -280
rect 18758 -314 18776 -304
rect 18718 -338 18776 -314
rect 18810 -314 18816 -304
rect 18850 -304 18908 -280
rect 18850 -314 18868 -304
rect 18810 -338 18868 -314
rect 18902 -314 18908 -304
rect 18942 -289 18971 -280
rect 19577 -289 19606 -280
rect 18942 -304 19606 -289
rect 19640 -304 19698 -280
rect 19732 -304 19790 -280
rect 19824 -304 19882 -280
rect 19916 -304 19974 -280
rect 20008 -304 20066 -280
rect 20100 -304 20158 -280
rect 20192 -304 20250 -280
rect 20284 -304 20342 -280
rect 20376 -289 20405 -280
rect 20535 -289 20564 -280
rect 20376 -304 20564 -289
rect 20598 -304 20656 -280
rect 20690 -304 20748 -280
rect 20782 -304 20840 -280
rect 20874 -304 20932 -280
rect 20966 -304 21024 -280
rect 21058 -304 21116 -280
rect 21150 -304 21208 -280
rect 21242 -304 21300 -280
rect 21334 -289 21363 -280
rect 21967 -289 21996 -280
rect 21334 -304 21996 -289
rect 22030 -304 22088 -280
rect 22122 -304 22180 -280
rect 22214 -304 22272 -280
rect 22306 -304 22364 -280
rect 22398 -304 22456 -280
rect 22490 -304 22548 -280
rect 22582 -304 22640 -280
rect 22674 -304 22732 -280
rect 22766 -289 22795 -280
rect 22927 -289 22956 -280
rect 22766 -304 22956 -289
rect 22990 -304 23048 -280
rect 23082 -304 23140 -280
rect 23174 -304 23232 -280
rect 23266 -304 23324 -280
rect 23358 -304 23416 -280
rect 23450 -304 23508 -280
rect 23542 -304 23600 -280
rect 23634 -304 23692 -280
rect 23726 -289 23755 -280
rect 24361 -289 24390 -280
rect 23726 -304 24390 -289
rect 24424 -304 24482 -280
rect 24516 -304 24574 -280
rect 24608 -304 24666 -280
rect 24700 -304 24758 -280
rect 24792 -304 24850 -280
rect 24884 -304 24942 -280
rect 24976 -304 25034 -280
rect 25068 -304 25126 -280
rect 18942 -314 18960 -304
rect 18902 -338 18960 -314
rect 18994 -338 19052 -304
rect 19086 -338 19144 -304
rect 19178 -338 19236 -304
rect 19270 -338 19328 -304
rect 19362 -338 19420 -304
rect 19454 -338 19512 -304
rect 19546 -338 19604 -304
rect 19640 -314 19696 -304
rect 19732 -314 19788 -304
rect 19824 -314 19880 -304
rect 19916 -314 19972 -304
rect 20008 -314 20064 -304
rect 20100 -314 20156 -304
rect 20192 -314 20248 -304
rect 20284 -314 20340 -304
rect 20376 -314 20432 -304
rect 19638 -338 19696 -314
rect 19730 -338 19788 -314
rect 19822 -338 19880 -314
rect 19914 -338 19972 -314
rect 20006 -338 20064 -314
rect 20098 -338 20156 -314
rect 20190 -338 20248 -314
rect 20282 -338 20340 -314
rect 20374 -338 20432 -314
rect 20466 -314 20564 -304
rect 20620 -314 20656 -304
rect 20712 -314 20748 -304
rect 20804 -314 20840 -304
rect 20896 -314 20932 -304
rect 20988 -314 21024 -304
rect 21080 -314 21116 -304
rect 21172 -314 21208 -304
rect 21264 -314 21300 -304
rect 20466 -338 20586 -314
rect 20620 -338 20678 -314
rect 20712 -338 20770 -314
rect 20804 -338 20862 -314
rect 20896 -338 20954 -314
rect 20988 -338 21046 -314
rect 21080 -338 21138 -314
rect 21172 -338 21230 -314
rect 21264 -338 21322 -314
rect 21356 -338 21414 -304
rect 21448 -338 21506 -304
rect 21540 -338 21598 -304
rect 21632 -338 21690 -304
rect 21724 -338 21782 -304
rect 21816 -338 21874 -304
rect 21908 -338 21966 -304
rect 22030 -314 22058 -304
rect 22122 -314 22150 -304
rect 22214 -314 22242 -304
rect 22306 -314 22334 -304
rect 22398 -314 22426 -304
rect 22490 -314 22518 -304
rect 22582 -314 22610 -304
rect 22674 -314 22702 -304
rect 22766 -314 22794 -304
rect 22000 -338 22058 -314
rect 22092 -338 22150 -314
rect 22184 -338 22242 -314
rect 22276 -338 22334 -314
rect 22368 -338 22426 -314
rect 22460 -338 22518 -314
rect 22552 -338 22610 -314
rect 22644 -338 22702 -314
rect 22736 -338 22794 -314
rect 22828 -338 22886 -304
rect 22920 -314 22956 -304
rect 23012 -314 23048 -304
rect 23104 -314 23140 -304
rect 23196 -314 23232 -304
rect 23288 -314 23324 -304
rect 23380 -314 23416 -304
rect 23472 -314 23508 -304
rect 23564 -314 23600 -304
rect 23656 -314 23692 -304
rect 22920 -338 22978 -314
rect 23012 -338 23070 -314
rect 23104 -338 23162 -314
rect 23196 -338 23254 -314
rect 23288 -338 23346 -314
rect 23380 -338 23438 -314
rect 23472 -338 23530 -314
rect 23564 -338 23622 -314
rect 23656 -338 23714 -314
rect 23748 -338 23806 -304
rect 23840 -338 23898 -304
rect 23932 -338 23990 -304
rect 24024 -338 24082 -304
rect 24116 -338 24174 -304
rect 24208 -338 24266 -304
rect 24300 -338 24358 -304
rect 24424 -314 24450 -304
rect 24516 -314 24542 -304
rect 24608 -314 24634 -304
rect 24700 -314 24726 -304
rect 24792 -314 24818 -304
rect 24884 -314 24910 -304
rect 24976 -314 25002 -304
rect 25068 -314 25094 -304
rect 25160 -314 25189 -280
rect 24392 -338 24450 -314
rect 24484 -338 24542 -314
rect 24576 -338 24634 -314
rect 24668 -338 24726 -314
rect 24760 -338 24818 -314
rect 24852 -338 24910 -314
rect 24944 -338 25002 -314
rect 25036 -338 25094 -314
rect 25128 -338 25189 -314
rect 24812 -400 24878 -392
rect 8575 -458 8604 -400
rect 8638 -458 8696 -400
rect 8730 -458 8788 -400
rect 8822 -458 8880 -400
rect 8914 -458 8972 -400
rect 9006 -458 9064 -400
rect 9098 -458 9156 -400
rect 9190 -458 9248 -400
rect 9282 -458 9340 -400
rect 9374 -458 9432 -400
rect 9466 -458 9524 -400
rect 9558 -458 9616 -400
rect 9650 -458 9708 -400
rect 9742 -458 9800 -400
rect 9834 -458 9892 -400
rect 9926 -458 9984 -400
rect 10018 -458 10076 -400
rect 10110 -458 10168 -400
rect 10202 -458 10260 -400
rect 10294 -458 10352 -400
rect 10386 -407 10628 -400
rect 10386 -424 10476 -407
rect 10510 -424 10628 -407
rect 10386 -458 10444 -424
rect 10510 -441 10536 -424
rect 10478 -458 10536 -441
rect 10570 -458 10628 -424
rect 10662 -458 10720 -400
rect 10754 -458 10812 -400
rect 10846 -458 10904 -400
rect 10938 -458 10996 -400
rect 11030 -458 11088 -400
rect 11122 -458 11180 -400
rect 11214 -458 11272 -400
rect 11306 -458 11364 -400
rect 11398 -458 11456 -400
rect 11490 -458 11548 -400
rect 11582 -458 11640 -400
rect 11674 -458 11732 -400
rect 11766 -458 11824 -400
rect 11858 -458 11916 -400
rect 11950 -458 12008 -400
rect 12042 -458 12100 -400
rect 12134 -458 12192 -400
rect 12226 -458 12284 -400
rect 12318 -458 12376 -400
rect 12410 -458 12468 -400
rect 12502 -458 12560 -400
rect 12594 -458 12652 -400
rect 12686 -458 12744 -400
rect 12778 -408 13020 -400
rect 12778 -424 12868 -408
rect 12902 -424 13020 -408
rect 12778 -458 12836 -424
rect 12902 -442 12928 -424
rect 12870 -458 12928 -442
rect 12962 -458 13020 -424
rect 13054 -458 13112 -400
rect 13146 -458 13204 -400
rect 13238 -458 13296 -400
rect 13330 -458 13388 -400
rect 13422 -458 13480 -400
rect 13514 -458 13572 -400
rect 13606 -458 13664 -400
rect 13698 -458 13756 -400
rect 13790 -458 13848 -400
rect 13882 -458 13940 -400
rect 13974 -458 14032 -400
rect 14066 -458 14124 -400
rect 14158 -458 14216 -400
rect 14250 -458 14308 -400
rect 14342 -458 14400 -400
rect 14434 -458 14492 -400
rect 14526 -458 14584 -400
rect 14618 -458 14676 -400
rect 14710 -458 14768 -400
rect 14802 -458 14860 -400
rect 14894 -458 14952 -400
rect 14986 -458 15044 -400
rect 15078 -458 15136 -400
rect 15170 -408 15412 -400
rect 15170 -424 15260 -408
rect 15294 -424 15412 -408
rect 15170 -458 15228 -424
rect 15294 -442 15320 -424
rect 15262 -458 15320 -442
rect 15354 -458 15412 -424
rect 15446 -458 15504 -400
rect 15538 -458 15596 -400
rect 15630 -458 15688 -400
rect 15722 -458 15780 -400
rect 15814 -458 15872 -400
rect 15906 -458 15964 -400
rect 15998 -458 16056 -400
rect 16090 -458 16148 -400
rect 16182 -458 16240 -400
rect 16274 -458 16332 -400
rect 16366 -458 16424 -400
rect 16458 -458 16516 -400
rect 16550 -458 16608 -400
rect 16642 -458 16700 -400
rect 16734 -458 16792 -400
rect 16826 -458 16884 -400
rect 16918 -458 16976 -400
rect 17010 -458 17068 -400
rect 17102 -458 17160 -400
rect 17194 -458 17252 -400
rect 17286 -458 17344 -400
rect 17378 -458 17436 -400
rect 17470 -458 17528 -400
rect 17562 -407 17804 -400
rect 17562 -424 17652 -407
rect 17686 -424 17804 -407
rect 17562 -458 17620 -424
rect 17686 -441 17712 -424
rect 17654 -458 17712 -441
rect 17746 -458 17804 -424
rect 17838 -458 17896 -400
rect 17930 -458 17988 -400
rect 18022 -458 18080 -400
rect 18114 -458 18172 -400
rect 18206 -458 18264 -400
rect 18298 -458 18356 -400
rect 18390 -458 18448 -400
rect 18482 -458 18540 -400
rect 18574 -458 18632 -400
rect 18666 -458 18724 -400
rect 18758 -458 18816 -400
rect 18850 -458 18908 -400
rect 18942 -458 19000 -400
rect 19034 -458 19092 -400
rect 19126 -458 19184 -400
rect 19218 -458 19276 -400
rect 19310 -458 19368 -400
rect 19402 -458 19460 -400
rect 19494 -458 19552 -400
rect 19586 -458 19644 -400
rect 19678 -458 19736 -400
rect 19770 -458 19828 -400
rect 19862 -458 19920 -400
rect 19954 -407 20196 -400
rect 19954 -424 20044 -407
rect 20078 -424 20196 -407
rect 19954 -458 20012 -424
rect 20078 -441 20104 -424
rect 20046 -458 20104 -441
rect 20138 -458 20196 -424
rect 20230 -458 20288 -400
rect 20322 -458 20380 -400
rect 20414 -458 20472 -400
rect 20506 -458 20564 -400
rect 20598 -458 20656 -400
rect 20690 -458 20748 -400
rect 20782 -458 20840 -400
rect 20874 -458 20932 -400
rect 20966 -458 21024 -400
rect 21058 -458 21116 -400
rect 21150 -458 21208 -400
rect 21242 -458 21300 -400
rect 21334 -458 21392 -400
rect 21426 -458 21484 -400
rect 21518 -458 21576 -400
rect 21610 -458 21668 -400
rect 21702 -458 21760 -400
rect 21794 -458 21852 -400
rect 21886 -458 21944 -400
rect 21978 -458 22036 -400
rect 22070 -458 22128 -400
rect 22162 -458 22220 -400
rect 22254 -458 22312 -400
rect 22346 -408 22588 -400
rect 22346 -424 22436 -408
rect 22470 -424 22588 -408
rect 22346 -458 22404 -424
rect 22470 -442 22496 -424
rect 22438 -458 22496 -442
rect 22530 -458 22588 -424
rect 22622 -458 22680 -400
rect 22714 -458 22772 -400
rect 22806 -458 22864 -400
rect 22898 -458 22956 -400
rect 22990 -458 23048 -400
rect 23082 -458 23140 -400
rect 23174 -458 23232 -400
rect 23266 -458 23324 -400
rect 23358 -458 23416 -400
rect 23450 -458 23508 -400
rect 23542 -458 23600 -400
rect 23634 -458 23692 -400
rect 23726 -458 23784 -400
rect 23818 -458 23876 -400
rect 23910 -458 23968 -400
rect 24002 -458 24060 -400
rect 24094 -458 24152 -400
rect 24186 -458 24244 -400
rect 24278 -458 24336 -400
rect 24370 -458 24428 -400
rect 24462 -458 24520 -400
rect 24554 -458 24612 -400
rect 24646 -458 24704 -400
rect 24738 -408 24980 -400
rect 24738 -424 24828 -408
rect 24862 -424 24980 -408
rect 24738 -458 24796 -424
rect 24862 -442 24888 -424
rect 24830 -458 24888 -442
rect 24922 -458 24980 -424
rect 25014 -458 25072 -400
rect 25106 -458 25164 -400
rect 25198 -458 25256 -400
rect 25290 -458 25319 -400
rect 8610 -508 8644 -492
rect 8610 -576 8644 -542
rect 8678 -524 8744 -458
rect 8678 -558 8694 -524
rect 8728 -558 8744 -524
rect 8778 -508 8822 -492
rect 8812 -542 8822 -508
rect 8778 -576 8822 -542
rect 8861 -524 8932 -458
rect 8861 -558 8882 -524
rect 8916 -558 8932 -524
rect 8966 -508 9000 -492
rect 9042 -535 9058 -501
rect 9092 -535 9208 -501
rect 8644 -610 8743 -592
rect 8610 -626 8743 -610
rect 8592 -706 8662 -660
rect 8592 -740 8601 -706
rect 8635 -721 8662 -706
rect 8592 -755 8606 -740
rect 8640 -755 8662 -721
rect 8592 -790 8662 -755
rect 8697 -721 8743 -626
rect 8697 -755 8708 -721
rect 8742 -755 8743 -721
rect 8697 -798 8743 -755
rect 8610 -832 8697 -824
rect 8731 -832 8743 -798
rect 8610 -858 8743 -832
rect 8812 -594 8822 -576
rect 8966 -592 9000 -542
rect 8778 -628 8788 -610
rect 8610 -866 8644 -858
rect 8778 -866 8822 -628
rect 8856 -626 9000 -592
rect 8856 -820 8890 -626
rect 9040 -628 9064 -594
rect 9098 -620 9140 -594
rect 9098 -628 9106 -620
rect 9040 -654 9106 -628
rect 8924 -682 9006 -660
rect 8924 -716 8941 -682
rect 8975 -716 9006 -682
rect 8924 -734 9006 -716
rect 8958 -768 9006 -734
rect 8924 -784 9006 -768
rect 9040 -670 9140 -654
rect 9040 -794 9084 -670
rect 9174 -704 9208 -535
rect 9256 -510 9332 -458
rect 9550 -500 9616 -458
rect 9256 -544 9272 -510
rect 9306 -544 9332 -510
rect 9392 -526 9426 -510
rect 9392 -578 9426 -560
rect 9550 -534 9566 -500
rect 9600 -534 9616 -500
rect 10039 -500 10115 -458
rect 9550 -568 9616 -534
rect 9825 -535 9841 -501
rect 9875 -535 9991 -501
rect 10039 -534 10055 -500
rect 10089 -534 10115 -500
rect 10303 -500 10581 -458
rect 10163 -526 10197 -510
rect 9242 -594 9512 -578
rect 9242 -620 9392 -594
rect 9276 -628 9392 -620
rect 9426 -628 9512 -594
rect 9550 -602 9566 -568
rect 9600 -602 9616 -568
rect 9787 -594 9834 -588
rect 9276 -654 9292 -628
rect 9242 -670 9292 -654
rect 9394 -704 9444 -688
rect 9174 -738 9410 -704
rect 9174 -746 9258 -738
rect 8856 -858 9000 -820
rect 9074 -828 9084 -794
rect 9040 -844 9084 -828
rect 9120 -816 9136 -782
rect 9170 -798 9190 -782
rect 9120 -832 9156 -816
rect 9120 -856 9190 -832
rect 8610 -916 8644 -900
rect 8678 -926 8694 -892
rect 8728 -926 8744 -892
rect 8812 -900 8822 -866
rect 8966 -874 9000 -858
rect 8778 -916 8822 -900
rect 8678 -968 8744 -926
rect 8861 -926 8882 -892
rect 8916 -926 8932 -892
rect 9224 -892 9258 -746
rect 9400 -754 9444 -738
rect 9478 -772 9512 -628
rect 9787 -620 9800 -594
rect 9821 -654 9834 -628
rect 9546 -662 9747 -654
rect 9546 -696 9708 -662
rect 9742 -696 9747 -662
rect 9787 -670 9834 -654
rect 9882 -620 9923 -604
rect 9882 -654 9889 -620
rect 9546 -702 9747 -696
rect 9546 -704 9612 -702
rect 9546 -738 9562 -704
rect 9596 -738 9612 -704
rect 9882 -724 9923 -654
rect 9788 -730 9923 -724
rect 9674 -772 9690 -738
rect 9724 -772 9740 -738
rect 9292 -806 9308 -772
rect 9342 -792 9358 -772
rect 9342 -798 9374 -792
rect 9292 -832 9340 -806
rect 9478 -806 9740 -772
rect 9788 -764 9800 -730
rect 9834 -760 9923 -730
rect 9957 -704 9991 -535
rect 10303 -534 10329 -500
rect 10363 -534 10531 -500
rect 10565 -534 10581 -500
rect 10163 -568 10197 -560
rect 10615 -537 10672 -492
rect 10025 -602 10581 -568
rect 10025 -620 10075 -602
rect 10059 -654 10075 -620
rect 10025 -670 10075 -654
rect 9957 -720 10227 -704
rect 9957 -738 10193 -720
rect 9834 -764 9856 -760
rect 9788 -773 9856 -764
rect 9812 -794 9856 -773
rect 9478 -832 9522 -806
rect 9292 -838 9374 -832
rect 9456 -866 9472 -832
rect 9506 -866 9522 -832
rect 9812 -828 9822 -794
rect 9556 -858 9590 -842
rect 9812 -844 9856 -828
rect 8966 -924 9000 -908
rect 8861 -968 8932 -926
rect 9055 -926 9071 -892
rect 9105 -926 9258 -892
rect 9055 -932 9258 -926
rect 9292 -896 9326 -880
rect 9292 -968 9326 -930
rect 9360 -890 9426 -884
rect 9360 -924 9376 -890
rect 9410 -900 9426 -890
rect 9957 -892 9991 -738
rect 10183 -754 10193 -738
rect 10183 -770 10227 -754
rect 10031 -806 10086 -772
rect 10120 -798 10140 -772
rect 10031 -832 10090 -806
rect 10124 -832 10140 -798
rect 10261 -817 10295 -602
rect 10329 -662 10433 -636
rect 10329 -696 10346 -662
rect 10380 -670 10433 -662
rect 10467 -670 10486 -636
rect 10380 -696 10386 -670
rect 10329 -704 10386 -696
rect 10363 -738 10386 -704
rect 10547 -720 10581 -602
rect 10649 -571 10672 -537
rect 10615 -605 10672 -571
rect 10649 -610 10672 -605
rect 10615 -644 10626 -639
rect 10660 -644 10672 -610
rect 10615 -659 10672 -644
rect 10329 -763 10386 -738
rect 10342 -800 10386 -763
rect 10422 -732 10513 -720
rect 10422 -766 10438 -732
rect 10472 -766 10513 -732
rect 10547 -736 10600 -720
rect 10547 -770 10566 -736
rect 10547 -786 10600 -770
rect 10261 -818 10298 -817
rect 10031 -838 10140 -832
rect 10218 -852 10248 -818
rect 10282 -852 10298 -818
rect 10342 -834 10470 -800
rect 9556 -900 9590 -892
rect 9410 -924 9590 -900
rect 9360 -934 9590 -924
rect 9640 -926 9660 -892
rect 9694 -926 9710 -892
rect 9640 -968 9710 -926
rect 9835 -926 9864 -892
rect 9898 -926 9991 -892
rect 9835 -932 9991 -926
rect 10025 -896 10090 -880
rect 10025 -930 10056 -896
rect 10025 -968 10090 -930
rect 10124 -910 10140 -876
rect 10174 -900 10190 -876
rect 10332 -884 10366 -868
rect 10174 -910 10332 -900
rect 10124 -918 10332 -910
rect 10124 -934 10366 -918
rect 10428 -882 10470 -834
rect 10428 -916 10436 -882
rect 10428 -932 10470 -916
rect 10520 -892 10581 -824
rect 10636 -842 10672 -659
rect 10520 -926 10531 -892
rect 10565 -926 10581 -892
rect 10520 -968 10581 -926
rect 10615 -858 10672 -842
rect 10649 -892 10672 -858
rect 10615 -934 10672 -892
rect 10707 -518 10770 -502
rect 10707 -552 10719 -518
rect 10753 -552 10770 -518
rect 10707 -586 10770 -552
rect 10707 -620 10719 -586
rect 10753 -620 10770 -586
rect 10707 -720 10770 -620
rect 10806 -512 10864 -458
rect 10806 -546 10814 -512
rect 10848 -546 10864 -512
rect 10806 -580 10864 -546
rect 10806 -614 10814 -580
rect 10848 -614 10864 -580
rect 10806 -632 10864 -614
rect 10898 -531 10950 -492
rect 10898 -536 10909 -531
rect 10943 -565 10950 -531
rect 10932 -570 10950 -565
rect 10898 -604 10950 -570
rect 10932 -638 10950 -604
rect 11002 -508 11036 -492
rect 11002 -576 11036 -542
rect 11070 -524 11136 -458
rect 11070 -558 11086 -524
rect 11120 -558 11136 -524
rect 11170 -508 11214 -492
rect 11204 -542 11214 -508
rect 11170 -576 11214 -542
rect 11253 -524 11324 -458
rect 11253 -558 11274 -524
rect 11308 -558 11324 -524
rect 11358 -508 11392 -492
rect 11434 -535 11450 -501
rect 11484 -535 11600 -501
rect 11036 -610 11135 -592
rect 11002 -626 11135 -610
rect 10898 -694 10950 -638
rect 10707 -736 10874 -720
rect 10707 -770 10840 -736
rect 10707 -786 10874 -770
rect 10707 -866 10770 -786
rect 10908 -820 10950 -694
rect 10984 -706 11054 -660
rect 10984 -740 10993 -706
rect 11027 -721 11054 -706
rect 10984 -755 10998 -740
rect 11032 -755 11054 -721
rect 10984 -790 11054 -755
rect 11089 -721 11135 -626
rect 11089 -755 11100 -721
rect 11134 -755 11135 -721
rect 10707 -900 10719 -866
rect 10753 -900 10770 -866
rect 10898 -856 10950 -820
rect 11089 -798 11135 -755
rect 10707 -934 10770 -900
rect 10805 -892 10864 -876
rect 10805 -926 10814 -892
rect 10848 -926 10864 -892
rect 10805 -968 10864 -926
rect 10932 -890 10950 -856
rect 10898 -934 10950 -890
rect 11002 -832 11089 -824
rect 11123 -832 11135 -798
rect 11002 -858 11135 -832
rect 11204 -594 11214 -576
rect 11358 -592 11392 -542
rect 11170 -628 11180 -610
rect 11002 -866 11036 -858
rect 11170 -866 11214 -628
rect 11248 -626 11392 -592
rect 11248 -820 11282 -626
rect 11432 -628 11456 -594
rect 11490 -620 11532 -594
rect 11490 -628 11498 -620
rect 11432 -654 11498 -628
rect 11316 -682 11398 -660
rect 11316 -716 11333 -682
rect 11367 -716 11398 -682
rect 11316 -734 11398 -716
rect 11350 -768 11398 -734
rect 11316 -784 11398 -768
rect 11432 -670 11532 -654
rect 11432 -794 11476 -670
rect 11566 -704 11600 -535
rect 11648 -510 11724 -458
rect 11942 -500 12008 -458
rect 11648 -544 11664 -510
rect 11698 -544 11724 -510
rect 11784 -526 11818 -510
rect 11784 -578 11818 -560
rect 11942 -534 11958 -500
rect 11992 -534 12008 -500
rect 12431 -500 12507 -458
rect 11942 -568 12008 -534
rect 12217 -535 12233 -501
rect 12267 -535 12383 -501
rect 12431 -534 12447 -500
rect 12481 -534 12507 -500
rect 12695 -500 12973 -458
rect 12555 -526 12589 -510
rect 11634 -594 11904 -578
rect 11634 -620 11784 -594
rect 11668 -628 11784 -620
rect 11818 -628 11904 -594
rect 11942 -602 11958 -568
rect 11992 -602 12008 -568
rect 12179 -594 12226 -588
rect 11668 -654 11684 -628
rect 11634 -670 11684 -654
rect 11786 -704 11836 -688
rect 11566 -738 11802 -704
rect 11566 -746 11650 -738
rect 11248 -858 11392 -820
rect 11466 -828 11476 -794
rect 11432 -844 11476 -828
rect 11512 -816 11528 -782
rect 11562 -798 11582 -782
rect 11512 -832 11548 -816
rect 11512 -856 11582 -832
rect 11002 -916 11036 -900
rect 11070 -926 11086 -892
rect 11120 -926 11136 -892
rect 11204 -900 11214 -866
rect 11358 -874 11392 -858
rect 11170 -916 11214 -900
rect 11070 -968 11136 -926
rect 11253 -926 11274 -892
rect 11308 -926 11324 -892
rect 11616 -892 11650 -746
rect 11792 -754 11836 -738
rect 11870 -772 11904 -628
rect 12179 -620 12192 -594
rect 12213 -654 12226 -628
rect 11938 -662 12139 -654
rect 11938 -696 12100 -662
rect 12134 -696 12139 -662
rect 12179 -670 12226 -654
rect 12274 -620 12315 -604
rect 12274 -654 12281 -620
rect 11938 -702 12139 -696
rect 11938 -704 12004 -702
rect 11938 -738 11954 -704
rect 11988 -738 12004 -704
rect 12274 -724 12315 -654
rect 12180 -730 12315 -724
rect 12066 -772 12082 -738
rect 12116 -772 12132 -738
rect 11684 -806 11700 -772
rect 11734 -792 11750 -772
rect 11734 -798 11766 -792
rect 11684 -832 11732 -806
rect 11870 -806 12132 -772
rect 12180 -764 12192 -730
rect 12226 -760 12315 -730
rect 12349 -704 12383 -535
rect 12695 -534 12721 -500
rect 12755 -534 12923 -500
rect 12957 -534 12973 -500
rect 12555 -568 12589 -560
rect 13007 -537 13064 -492
rect 12417 -602 12973 -568
rect 12417 -620 12467 -602
rect 12451 -654 12467 -620
rect 12417 -670 12467 -654
rect 12349 -720 12619 -704
rect 12349 -738 12585 -720
rect 12226 -764 12248 -760
rect 12180 -773 12248 -764
rect 12204 -794 12248 -773
rect 11870 -832 11914 -806
rect 11684 -838 11766 -832
rect 11848 -866 11864 -832
rect 11898 -866 11914 -832
rect 12204 -828 12214 -794
rect 11948 -858 11982 -842
rect 12204 -844 12248 -828
rect 11358 -924 11392 -908
rect 11253 -968 11324 -926
rect 11447 -926 11463 -892
rect 11497 -926 11650 -892
rect 11447 -932 11650 -926
rect 11684 -896 11718 -880
rect 11684 -968 11718 -930
rect 11752 -890 11818 -884
rect 11752 -924 11768 -890
rect 11802 -900 11818 -890
rect 12349 -892 12383 -738
rect 12575 -754 12585 -738
rect 12575 -770 12619 -754
rect 12423 -806 12478 -772
rect 12512 -798 12532 -772
rect 12423 -832 12482 -806
rect 12516 -832 12532 -798
rect 12653 -817 12687 -602
rect 12721 -662 12825 -636
rect 12721 -696 12738 -662
rect 12772 -670 12825 -662
rect 12859 -670 12878 -636
rect 12772 -696 12778 -670
rect 12721 -704 12778 -696
rect 12755 -738 12778 -704
rect 12939 -720 12973 -602
rect 13041 -571 13064 -537
rect 13007 -605 13064 -571
rect 13041 -609 13064 -605
rect 13007 -643 13018 -639
rect 13052 -643 13064 -609
rect 13007 -659 13064 -643
rect 12721 -763 12778 -738
rect 12734 -800 12778 -763
rect 12814 -732 12905 -720
rect 12814 -766 12830 -732
rect 12864 -766 12905 -732
rect 12939 -736 12992 -720
rect 12939 -770 12958 -736
rect 12939 -786 12992 -770
rect 12653 -818 12690 -817
rect 12423 -838 12532 -832
rect 12610 -852 12640 -818
rect 12674 -852 12690 -818
rect 12734 -834 12862 -800
rect 11948 -900 11982 -892
rect 11802 -924 11982 -900
rect 11752 -934 11982 -924
rect 12032 -926 12052 -892
rect 12086 -926 12102 -892
rect 12032 -968 12102 -926
rect 12227 -926 12256 -892
rect 12290 -926 12383 -892
rect 12227 -932 12383 -926
rect 12417 -896 12482 -880
rect 12417 -930 12448 -896
rect 12417 -968 12482 -930
rect 12516 -910 12532 -876
rect 12566 -900 12582 -876
rect 12724 -884 12758 -868
rect 12566 -910 12724 -900
rect 12516 -918 12724 -910
rect 12516 -934 12758 -918
rect 12820 -882 12862 -834
rect 12820 -916 12828 -882
rect 12820 -932 12862 -916
rect 12912 -892 12973 -824
rect 13028 -842 13064 -659
rect 12912 -926 12923 -892
rect 12957 -926 12973 -892
rect 12912 -968 12973 -926
rect 13007 -858 13064 -842
rect 13041 -892 13064 -858
rect 13007 -934 13064 -892
rect 13099 -518 13162 -502
rect 13099 -552 13111 -518
rect 13145 -552 13162 -518
rect 13099 -586 13162 -552
rect 13099 -620 13111 -586
rect 13145 -620 13162 -586
rect 13099 -720 13162 -620
rect 13198 -512 13256 -458
rect 13198 -546 13206 -512
rect 13240 -546 13256 -512
rect 13198 -580 13256 -546
rect 13198 -614 13206 -580
rect 13240 -614 13256 -580
rect 13198 -632 13256 -614
rect 13290 -531 13342 -492
rect 13290 -536 13301 -531
rect 13335 -565 13342 -531
rect 13324 -570 13342 -565
rect 13290 -604 13342 -570
rect 13324 -638 13342 -604
rect 13394 -508 13428 -492
rect 13394 -576 13428 -542
rect 13462 -524 13528 -458
rect 13462 -558 13478 -524
rect 13512 -558 13528 -524
rect 13562 -508 13606 -492
rect 13596 -542 13606 -508
rect 13562 -576 13606 -542
rect 13645 -524 13716 -458
rect 13645 -558 13666 -524
rect 13700 -558 13716 -524
rect 13750 -508 13784 -492
rect 13826 -535 13842 -501
rect 13876 -535 13992 -501
rect 13428 -610 13527 -592
rect 13394 -626 13527 -610
rect 13290 -694 13342 -638
rect 13099 -736 13266 -720
rect 13099 -770 13232 -736
rect 13099 -786 13266 -770
rect 13099 -866 13162 -786
rect 13300 -820 13342 -694
rect 13376 -706 13446 -660
rect 13376 -740 13385 -706
rect 13419 -721 13446 -706
rect 13376 -755 13390 -740
rect 13424 -755 13446 -721
rect 13376 -790 13446 -755
rect 13481 -721 13527 -626
rect 13481 -755 13492 -721
rect 13526 -755 13527 -721
rect 13099 -900 13111 -866
rect 13145 -900 13162 -866
rect 13290 -856 13342 -820
rect 13481 -798 13527 -755
rect 13099 -934 13162 -900
rect 13197 -892 13256 -876
rect 13197 -926 13206 -892
rect 13240 -926 13256 -892
rect 13197 -968 13256 -926
rect 13324 -890 13342 -856
rect 13290 -934 13342 -890
rect 13394 -832 13481 -824
rect 13515 -832 13527 -798
rect 13394 -858 13527 -832
rect 13596 -594 13606 -576
rect 13750 -592 13784 -542
rect 13562 -628 13572 -610
rect 13394 -866 13428 -858
rect 13562 -866 13606 -628
rect 13640 -626 13784 -592
rect 13640 -820 13674 -626
rect 13824 -628 13848 -594
rect 13882 -620 13924 -594
rect 13882 -628 13890 -620
rect 13824 -654 13890 -628
rect 13708 -681 13790 -660
rect 13708 -715 13725 -681
rect 13759 -715 13790 -681
rect 13708 -734 13790 -715
rect 13742 -768 13790 -734
rect 13708 -784 13790 -768
rect 13824 -670 13924 -654
rect 13824 -794 13868 -670
rect 13958 -704 13992 -535
rect 14040 -510 14116 -458
rect 14334 -500 14400 -458
rect 14040 -544 14056 -510
rect 14090 -544 14116 -510
rect 14176 -526 14210 -510
rect 14176 -578 14210 -560
rect 14334 -534 14350 -500
rect 14384 -534 14400 -500
rect 14823 -500 14899 -458
rect 14334 -568 14400 -534
rect 14609 -535 14625 -501
rect 14659 -535 14775 -501
rect 14823 -534 14839 -500
rect 14873 -534 14899 -500
rect 15087 -500 15365 -458
rect 14947 -526 14981 -510
rect 14026 -594 14296 -578
rect 14026 -620 14176 -594
rect 14060 -628 14176 -620
rect 14210 -628 14296 -594
rect 14334 -602 14350 -568
rect 14384 -602 14400 -568
rect 14571 -594 14618 -588
rect 14060 -654 14076 -628
rect 14026 -670 14076 -654
rect 14178 -704 14228 -688
rect 13958 -738 14194 -704
rect 13958 -746 14042 -738
rect 13640 -858 13784 -820
rect 13858 -828 13868 -794
rect 13824 -844 13868 -828
rect 13904 -816 13920 -782
rect 13954 -798 13974 -782
rect 13904 -832 13940 -816
rect 13904 -856 13974 -832
rect 13394 -916 13428 -900
rect 13462 -926 13478 -892
rect 13512 -926 13528 -892
rect 13596 -900 13606 -866
rect 13750 -874 13784 -858
rect 13562 -916 13606 -900
rect 13462 -968 13528 -926
rect 13645 -926 13666 -892
rect 13700 -926 13716 -892
rect 14008 -892 14042 -746
rect 14184 -754 14228 -738
rect 14262 -772 14296 -628
rect 14571 -620 14584 -594
rect 14605 -654 14618 -628
rect 14330 -662 14531 -654
rect 14330 -696 14492 -662
rect 14526 -696 14531 -662
rect 14571 -670 14618 -654
rect 14666 -620 14707 -604
rect 14666 -654 14673 -620
rect 14330 -702 14531 -696
rect 14330 -704 14396 -702
rect 14330 -738 14346 -704
rect 14380 -738 14396 -704
rect 14666 -724 14707 -654
rect 14572 -730 14707 -724
rect 14458 -772 14474 -738
rect 14508 -772 14524 -738
rect 14076 -806 14092 -772
rect 14126 -792 14142 -772
rect 14126 -798 14158 -792
rect 14076 -832 14124 -806
rect 14262 -806 14524 -772
rect 14572 -764 14584 -730
rect 14618 -760 14707 -730
rect 14741 -704 14775 -535
rect 15087 -534 15113 -500
rect 15147 -534 15315 -500
rect 15349 -534 15365 -500
rect 14947 -568 14981 -560
rect 15399 -537 15456 -492
rect 14809 -602 15365 -568
rect 14809 -620 14859 -602
rect 14843 -654 14859 -620
rect 14809 -670 14859 -654
rect 14741 -720 15011 -704
rect 14741 -738 14977 -720
rect 14618 -764 14640 -760
rect 14572 -773 14640 -764
rect 14596 -794 14640 -773
rect 14262 -832 14306 -806
rect 14076 -838 14158 -832
rect 14240 -866 14256 -832
rect 14290 -866 14306 -832
rect 14596 -828 14606 -794
rect 14340 -858 14374 -842
rect 14596 -844 14640 -828
rect 13750 -924 13784 -908
rect 13645 -968 13716 -926
rect 13839 -926 13855 -892
rect 13889 -926 14042 -892
rect 13839 -932 14042 -926
rect 14076 -896 14110 -880
rect 14076 -968 14110 -930
rect 14144 -890 14210 -884
rect 14144 -924 14160 -890
rect 14194 -900 14210 -890
rect 14741 -892 14775 -738
rect 14967 -754 14977 -738
rect 14967 -770 15011 -754
rect 14815 -806 14870 -772
rect 14904 -798 14924 -772
rect 14815 -832 14874 -806
rect 14908 -832 14924 -798
rect 15045 -817 15079 -602
rect 15113 -662 15217 -636
rect 15113 -696 15130 -662
rect 15164 -670 15217 -662
rect 15251 -670 15270 -636
rect 15164 -696 15170 -670
rect 15113 -704 15170 -696
rect 15147 -738 15170 -704
rect 15331 -720 15365 -602
rect 15433 -571 15456 -537
rect 15399 -605 15456 -571
rect 15433 -609 15456 -605
rect 15399 -643 15409 -639
rect 15443 -643 15456 -609
rect 15399 -659 15456 -643
rect 15113 -763 15170 -738
rect 15126 -800 15170 -763
rect 15206 -732 15297 -720
rect 15206 -766 15222 -732
rect 15256 -766 15297 -732
rect 15331 -736 15384 -720
rect 15331 -770 15350 -736
rect 15331 -786 15384 -770
rect 15045 -818 15082 -817
rect 14815 -838 14924 -832
rect 15002 -852 15032 -818
rect 15066 -852 15082 -818
rect 15126 -834 15254 -800
rect 14340 -900 14374 -892
rect 14194 -924 14374 -900
rect 14144 -934 14374 -924
rect 14424 -926 14444 -892
rect 14478 -926 14494 -892
rect 14424 -968 14494 -926
rect 14619 -926 14648 -892
rect 14682 -926 14775 -892
rect 14619 -932 14775 -926
rect 14809 -896 14874 -880
rect 14809 -930 14840 -896
rect 14809 -968 14874 -930
rect 14908 -910 14924 -876
rect 14958 -900 14974 -876
rect 15116 -884 15150 -868
rect 14958 -910 15116 -900
rect 14908 -918 15116 -910
rect 14908 -934 15150 -918
rect 15212 -882 15254 -834
rect 15212 -916 15220 -882
rect 15212 -932 15254 -916
rect 15304 -892 15365 -824
rect 15420 -842 15456 -659
rect 15304 -926 15315 -892
rect 15349 -926 15365 -892
rect 15304 -968 15365 -926
rect 15399 -858 15456 -842
rect 15433 -892 15456 -858
rect 15399 -934 15456 -892
rect 15491 -518 15554 -502
rect 15491 -552 15503 -518
rect 15537 -552 15554 -518
rect 15491 -586 15554 -552
rect 15491 -620 15503 -586
rect 15537 -620 15554 -586
rect 15491 -720 15554 -620
rect 15590 -512 15648 -458
rect 15590 -546 15598 -512
rect 15632 -546 15648 -512
rect 15590 -580 15648 -546
rect 15590 -614 15598 -580
rect 15632 -614 15648 -580
rect 15590 -632 15648 -614
rect 15682 -531 15734 -492
rect 15682 -536 15693 -531
rect 15727 -565 15734 -531
rect 15716 -570 15734 -565
rect 15682 -604 15734 -570
rect 15716 -638 15734 -604
rect 15786 -508 15820 -492
rect 15786 -576 15820 -542
rect 15854 -524 15920 -458
rect 15854 -558 15870 -524
rect 15904 -558 15920 -524
rect 15954 -508 15998 -492
rect 15988 -542 15998 -508
rect 15954 -576 15998 -542
rect 16037 -524 16108 -458
rect 16037 -558 16058 -524
rect 16092 -558 16108 -524
rect 16142 -508 16176 -492
rect 16218 -535 16234 -501
rect 16268 -535 16384 -501
rect 15820 -610 15919 -592
rect 15786 -626 15919 -610
rect 15682 -694 15734 -638
rect 15491 -736 15658 -720
rect 15491 -770 15624 -736
rect 15491 -786 15658 -770
rect 15491 -866 15554 -786
rect 15692 -820 15734 -694
rect 15768 -706 15838 -660
rect 15768 -740 15777 -706
rect 15811 -721 15838 -706
rect 15768 -755 15782 -740
rect 15816 -755 15838 -721
rect 15768 -790 15838 -755
rect 15873 -721 15919 -626
rect 15873 -755 15884 -721
rect 15918 -755 15919 -721
rect 15491 -900 15503 -866
rect 15537 -900 15554 -866
rect 15682 -856 15734 -820
rect 15873 -798 15919 -755
rect 15491 -934 15554 -900
rect 15589 -892 15648 -876
rect 15589 -926 15598 -892
rect 15632 -926 15648 -892
rect 15589 -968 15648 -926
rect 15716 -890 15734 -856
rect 15682 -934 15734 -890
rect 15786 -832 15873 -824
rect 15907 -832 15919 -798
rect 15786 -858 15919 -832
rect 15988 -594 15998 -576
rect 16142 -592 16176 -542
rect 15954 -628 15964 -610
rect 15786 -866 15820 -858
rect 15954 -866 15998 -628
rect 16032 -626 16176 -592
rect 16032 -820 16066 -626
rect 16216 -628 16240 -594
rect 16274 -620 16316 -594
rect 16274 -628 16282 -620
rect 16216 -654 16282 -628
rect 16100 -681 16182 -660
rect 16100 -715 16117 -681
rect 16151 -715 16182 -681
rect 16100 -734 16182 -715
rect 16134 -768 16182 -734
rect 16100 -784 16182 -768
rect 16216 -670 16316 -654
rect 16216 -794 16260 -670
rect 16350 -704 16384 -535
rect 16432 -510 16508 -458
rect 16726 -500 16792 -458
rect 16432 -544 16448 -510
rect 16482 -544 16508 -510
rect 16568 -526 16602 -510
rect 16568 -578 16602 -560
rect 16726 -534 16742 -500
rect 16776 -534 16792 -500
rect 17215 -500 17291 -458
rect 16726 -568 16792 -534
rect 17001 -535 17017 -501
rect 17051 -535 17167 -501
rect 17215 -534 17231 -500
rect 17265 -534 17291 -500
rect 17479 -500 17757 -458
rect 17339 -526 17373 -510
rect 16418 -594 16688 -578
rect 16418 -620 16568 -594
rect 16452 -628 16568 -620
rect 16602 -628 16688 -594
rect 16726 -602 16742 -568
rect 16776 -602 16792 -568
rect 16963 -594 17010 -588
rect 16452 -654 16468 -628
rect 16418 -670 16468 -654
rect 16570 -704 16620 -688
rect 16350 -738 16586 -704
rect 16350 -746 16434 -738
rect 16032 -858 16176 -820
rect 16250 -828 16260 -794
rect 16216 -844 16260 -828
rect 16296 -816 16312 -782
rect 16346 -798 16366 -782
rect 16296 -832 16332 -816
rect 16296 -856 16366 -832
rect 15786 -916 15820 -900
rect 15854 -926 15870 -892
rect 15904 -926 15920 -892
rect 15988 -900 15998 -866
rect 16142 -874 16176 -858
rect 15954 -916 15998 -900
rect 15854 -968 15920 -926
rect 16037 -926 16058 -892
rect 16092 -926 16108 -892
rect 16400 -892 16434 -746
rect 16576 -754 16620 -738
rect 16654 -772 16688 -628
rect 16963 -620 16976 -594
rect 16997 -654 17010 -628
rect 16722 -662 16923 -654
rect 16722 -696 16884 -662
rect 16918 -696 16923 -662
rect 16963 -670 17010 -654
rect 17058 -620 17099 -604
rect 17058 -654 17065 -620
rect 16722 -702 16923 -696
rect 16722 -704 16788 -702
rect 16722 -738 16738 -704
rect 16772 -738 16788 -704
rect 17058 -724 17099 -654
rect 16964 -730 17099 -724
rect 16850 -772 16866 -738
rect 16900 -772 16916 -738
rect 16468 -806 16484 -772
rect 16518 -792 16534 -772
rect 16518 -798 16550 -792
rect 16468 -832 16516 -806
rect 16654 -806 16916 -772
rect 16964 -764 16976 -730
rect 17010 -760 17099 -730
rect 17133 -704 17167 -535
rect 17479 -534 17505 -500
rect 17539 -534 17707 -500
rect 17741 -534 17757 -500
rect 17339 -568 17373 -560
rect 17791 -537 17848 -492
rect 17201 -602 17757 -568
rect 17201 -620 17251 -602
rect 17235 -654 17251 -620
rect 17201 -670 17251 -654
rect 17133 -720 17403 -704
rect 17133 -738 17369 -720
rect 17010 -764 17032 -760
rect 16964 -773 17032 -764
rect 16988 -794 17032 -773
rect 16654 -832 16698 -806
rect 16468 -838 16550 -832
rect 16632 -866 16648 -832
rect 16682 -866 16698 -832
rect 16988 -828 16998 -794
rect 16732 -858 16766 -842
rect 16988 -844 17032 -828
rect 16142 -924 16176 -908
rect 16037 -968 16108 -926
rect 16231 -926 16247 -892
rect 16281 -926 16434 -892
rect 16231 -932 16434 -926
rect 16468 -896 16502 -880
rect 16468 -968 16502 -930
rect 16536 -890 16602 -884
rect 16536 -924 16552 -890
rect 16586 -900 16602 -890
rect 17133 -892 17167 -738
rect 17359 -754 17369 -738
rect 17359 -770 17403 -754
rect 17207 -806 17262 -772
rect 17296 -798 17316 -772
rect 17207 -832 17266 -806
rect 17300 -832 17316 -798
rect 17437 -817 17471 -602
rect 17505 -662 17609 -636
rect 17505 -696 17522 -662
rect 17556 -670 17609 -662
rect 17643 -670 17662 -636
rect 17556 -696 17562 -670
rect 17505 -704 17562 -696
rect 17539 -738 17562 -704
rect 17723 -720 17757 -602
rect 17825 -571 17848 -537
rect 17791 -605 17848 -571
rect 17825 -608 17848 -605
rect 17791 -642 17802 -639
rect 17836 -642 17848 -608
rect 17791 -659 17848 -642
rect 17505 -763 17562 -738
rect 17518 -800 17562 -763
rect 17598 -732 17689 -720
rect 17598 -766 17614 -732
rect 17648 -766 17689 -732
rect 17723 -736 17776 -720
rect 17723 -770 17742 -736
rect 17723 -786 17776 -770
rect 17437 -818 17474 -817
rect 17207 -838 17316 -832
rect 17394 -852 17424 -818
rect 17458 -852 17474 -818
rect 17518 -834 17646 -800
rect 16732 -900 16766 -892
rect 16586 -924 16766 -900
rect 16536 -934 16766 -924
rect 16816 -926 16836 -892
rect 16870 -926 16886 -892
rect 16816 -968 16886 -926
rect 17011 -926 17040 -892
rect 17074 -926 17167 -892
rect 17011 -932 17167 -926
rect 17201 -896 17266 -880
rect 17201 -930 17232 -896
rect 17201 -968 17266 -930
rect 17300 -910 17316 -876
rect 17350 -900 17366 -876
rect 17508 -884 17542 -868
rect 17350 -910 17508 -900
rect 17300 -918 17508 -910
rect 17300 -934 17542 -918
rect 17604 -882 17646 -834
rect 17604 -916 17612 -882
rect 17604 -932 17646 -916
rect 17696 -892 17757 -824
rect 17812 -842 17848 -659
rect 17696 -926 17707 -892
rect 17741 -926 17757 -892
rect 17696 -968 17757 -926
rect 17791 -858 17848 -842
rect 17825 -892 17848 -858
rect 17791 -934 17848 -892
rect 17883 -518 17946 -502
rect 17883 -552 17895 -518
rect 17929 -552 17946 -518
rect 17883 -586 17946 -552
rect 17883 -620 17895 -586
rect 17929 -620 17946 -586
rect 17883 -720 17946 -620
rect 17982 -512 18040 -458
rect 17982 -546 17990 -512
rect 18024 -546 18040 -512
rect 17982 -580 18040 -546
rect 17982 -614 17990 -580
rect 18024 -614 18040 -580
rect 17982 -632 18040 -614
rect 18074 -531 18126 -492
rect 18074 -536 18085 -531
rect 18119 -565 18126 -531
rect 18108 -570 18126 -565
rect 18074 -604 18126 -570
rect 18108 -638 18126 -604
rect 18178 -508 18212 -492
rect 18178 -576 18212 -542
rect 18246 -524 18312 -458
rect 18246 -558 18262 -524
rect 18296 -558 18312 -524
rect 18346 -508 18390 -492
rect 18380 -542 18390 -508
rect 18346 -576 18390 -542
rect 18429 -524 18500 -458
rect 18429 -558 18450 -524
rect 18484 -558 18500 -524
rect 18534 -508 18568 -492
rect 18610 -535 18626 -501
rect 18660 -535 18776 -501
rect 18212 -610 18311 -592
rect 18178 -626 18311 -610
rect 18074 -694 18126 -638
rect 17883 -736 18050 -720
rect 17883 -770 18016 -736
rect 17883 -786 18050 -770
rect 17883 -866 17946 -786
rect 18084 -820 18126 -694
rect 18160 -705 18230 -660
rect 18160 -739 18168 -705
rect 18202 -721 18230 -705
rect 18160 -755 18174 -739
rect 18208 -755 18230 -721
rect 18160 -790 18230 -755
rect 18265 -721 18311 -626
rect 18265 -755 18276 -721
rect 18310 -755 18311 -721
rect 17883 -900 17895 -866
rect 17929 -900 17946 -866
rect 18074 -856 18126 -820
rect 18265 -798 18311 -755
rect 17883 -934 17946 -900
rect 17981 -892 18040 -876
rect 17981 -926 17990 -892
rect 18024 -926 18040 -892
rect 17981 -968 18040 -926
rect 18108 -890 18126 -856
rect 18074 -934 18126 -890
rect 18178 -832 18265 -824
rect 18299 -832 18311 -798
rect 18178 -858 18311 -832
rect 18380 -594 18390 -576
rect 18534 -592 18568 -542
rect 18346 -628 18356 -610
rect 18178 -866 18212 -858
rect 18346 -866 18390 -628
rect 18424 -626 18568 -592
rect 18424 -820 18458 -626
rect 18608 -628 18632 -594
rect 18666 -620 18708 -594
rect 18666 -628 18674 -620
rect 18608 -654 18674 -628
rect 18492 -682 18574 -660
rect 18492 -716 18509 -682
rect 18543 -716 18574 -682
rect 18492 -734 18574 -716
rect 18526 -768 18574 -734
rect 18492 -784 18574 -768
rect 18608 -670 18708 -654
rect 18608 -794 18652 -670
rect 18742 -704 18776 -535
rect 18824 -510 18900 -458
rect 19118 -500 19184 -458
rect 18824 -544 18840 -510
rect 18874 -544 18900 -510
rect 18960 -526 18994 -510
rect 18960 -578 18994 -560
rect 19118 -534 19134 -500
rect 19168 -534 19184 -500
rect 19607 -500 19683 -458
rect 19118 -568 19184 -534
rect 19393 -535 19409 -501
rect 19443 -535 19559 -501
rect 19607 -534 19623 -500
rect 19657 -534 19683 -500
rect 19871 -500 20149 -458
rect 19731 -526 19765 -510
rect 18810 -594 19080 -578
rect 18810 -620 18960 -594
rect 18844 -628 18960 -620
rect 18994 -628 19080 -594
rect 19118 -602 19134 -568
rect 19168 -602 19184 -568
rect 19355 -594 19402 -588
rect 18844 -654 18860 -628
rect 18810 -670 18860 -654
rect 18962 -704 19012 -688
rect 18742 -738 18978 -704
rect 18742 -746 18826 -738
rect 18424 -858 18568 -820
rect 18642 -828 18652 -794
rect 18608 -844 18652 -828
rect 18688 -816 18704 -782
rect 18738 -798 18758 -782
rect 18688 -832 18724 -816
rect 18688 -856 18758 -832
rect 18178 -916 18212 -900
rect 18246 -926 18262 -892
rect 18296 -926 18312 -892
rect 18380 -900 18390 -866
rect 18534 -874 18568 -858
rect 18346 -916 18390 -900
rect 18246 -968 18312 -926
rect 18429 -926 18450 -892
rect 18484 -926 18500 -892
rect 18792 -892 18826 -746
rect 18968 -754 19012 -738
rect 19046 -772 19080 -628
rect 19355 -620 19368 -594
rect 19389 -654 19402 -628
rect 19114 -662 19315 -654
rect 19114 -696 19276 -662
rect 19310 -696 19315 -662
rect 19355 -670 19402 -654
rect 19450 -620 19491 -604
rect 19450 -654 19457 -620
rect 19114 -702 19315 -696
rect 19114 -704 19180 -702
rect 19114 -738 19130 -704
rect 19164 -738 19180 -704
rect 19450 -724 19491 -654
rect 19356 -730 19491 -724
rect 19242 -772 19258 -738
rect 19292 -772 19308 -738
rect 18860 -806 18876 -772
rect 18910 -792 18926 -772
rect 18910 -798 18942 -792
rect 18860 -832 18908 -806
rect 19046 -806 19308 -772
rect 19356 -764 19368 -730
rect 19402 -760 19491 -730
rect 19525 -704 19559 -535
rect 19871 -534 19897 -500
rect 19931 -534 20099 -500
rect 20133 -534 20149 -500
rect 19731 -568 19765 -560
rect 20183 -537 20240 -492
rect 19593 -602 20149 -568
rect 19593 -620 19643 -602
rect 19627 -654 19643 -620
rect 19593 -670 19643 -654
rect 19525 -720 19795 -704
rect 19525 -738 19761 -720
rect 19402 -764 19424 -760
rect 19356 -773 19424 -764
rect 19380 -794 19424 -773
rect 19046 -832 19090 -806
rect 18860 -838 18942 -832
rect 19024 -866 19040 -832
rect 19074 -866 19090 -832
rect 19380 -828 19390 -794
rect 19124 -858 19158 -842
rect 19380 -844 19424 -828
rect 18534 -924 18568 -908
rect 18429 -968 18500 -926
rect 18623 -926 18639 -892
rect 18673 -926 18826 -892
rect 18623 -932 18826 -926
rect 18860 -896 18894 -880
rect 18860 -968 18894 -930
rect 18928 -890 18994 -884
rect 18928 -924 18944 -890
rect 18978 -900 18994 -890
rect 19525 -892 19559 -738
rect 19751 -754 19761 -738
rect 19751 -770 19795 -754
rect 19599 -806 19654 -772
rect 19688 -798 19708 -772
rect 19599 -832 19658 -806
rect 19692 -832 19708 -798
rect 19829 -817 19863 -602
rect 19897 -662 20001 -636
rect 19897 -696 19914 -662
rect 19948 -670 20001 -662
rect 20035 -670 20054 -636
rect 19948 -696 19954 -670
rect 19897 -704 19954 -696
rect 19931 -738 19954 -704
rect 20115 -720 20149 -602
rect 20217 -571 20240 -537
rect 20183 -605 20240 -571
rect 20217 -609 20240 -605
rect 20183 -643 20193 -639
rect 20227 -643 20240 -609
rect 20183 -659 20240 -643
rect 19897 -763 19954 -738
rect 19910 -800 19954 -763
rect 19990 -732 20081 -720
rect 19990 -766 20006 -732
rect 20040 -766 20081 -732
rect 20115 -736 20168 -720
rect 20115 -770 20134 -736
rect 20115 -786 20168 -770
rect 19829 -818 19866 -817
rect 19599 -838 19708 -832
rect 19786 -852 19816 -818
rect 19850 -852 19866 -818
rect 19910 -834 20038 -800
rect 19124 -900 19158 -892
rect 18978 -924 19158 -900
rect 18928 -934 19158 -924
rect 19208 -926 19228 -892
rect 19262 -926 19278 -892
rect 19208 -968 19278 -926
rect 19403 -926 19432 -892
rect 19466 -926 19559 -892
rect 19403 -932 19559 -926
rect 19593 -896 19658 -880
rect 19593 -930 19624 -896
rect 19593 -968 19658 -930
rect 19692 -910 19708 -876
rect 19742 -900 19758 -876
rect 19900 -884 19934 -868
rect 19742 -910 19900 -900
rect 19692 -918 19900 -910
rect 19692 -934 19934 -918
rect 19996 -882 20038 -834
rect 19996 -916 20004 -882
rect 19996 -932 20038 -916
rect 20088 -892 20149 -824
rect 20204 -842 20240 -659
rect 20088 -926 20099 -892
rect 20133 -926 20149 -892
rect 20088 -968 20149 -926
rect 20183 -858 20240 -842
rect 20217 -892 20240 -858
rect 20183 -934 20240 -892
rect 20275 -518 20338 -502
rect 20275 -552 20287 -518
rect 20321 -552 20338 -518
rect 20275 -586 20338 -552
rect 20275 -620 20287 -586
rect 20321 -620 20338 -586
rect 20275 -720 20338 -620
rect 20374 -512 20432 -458
rect 20374 -546 20382 -512
rect 20416 -546 20432 -512
rect 20374 -580 20432 -546
rect 20374 -614 20382 -580
rect 20416 -614 20432 -580
rect 20374 -632 20432 -614
rect 20466 -531 20518 -492
rect 20466 -536 20477 -531
rect 20511 -565 20518 -531
rect 20500 -570 20518 -565
rect 20466 -604 20518 -570
rect 20500 -638 20518 -604
rect 20570 -508 20604 -492
rect 20570 -576 20604 -542
rect 20638 -524 20704 -458
rect 20638 -558 20654 -524
rect 20688 -558 20704 -524
rect 20738 -508 20782 -492
rect 20772 -542 20782 -508
rect 20738 -576 20782 -542
rect 20821 -524 20892 -458
rect 20821 -558 20842 -524
rect 20876 -558 20892 -524
rect 20926 -508 20960 -492
rect 21002 -535 21018 -501
rect 21052 -535 21168 -501
rect 20604 -610 20703 -592
rect 20570 -626 20703 -610
rect 20466 -694 20518 -638
rect 20275 -736 20442 -720
rect 20275 -770 20408 -736
rect 20275 -786 20442 -770
rect 20275 -866 20338 -786
rect 20476 -820 20518 -694
rect 20552 -706 20622 -660
rect 20552 -740 20560 -706
rect 20594 -721 20622 -706
rect 20552 -755 20566 -740
rect 20600 -755 20622 -721
rect 20552 -790 20622 -755
rect 20657 -721 20703 -626
rect 20657 -755 20668 -721
rect 20702 -755 20703 -721
rect 20275 -900 20287 -866
rect 20321 -900 20338 -866
rect 20466 -856 20518 -820
rect 20657 -798 20703 -755
rect 20275 -934 20338 -900
rect 20373 -892 20432 -876
rect 20373 -926 20382 -892
rect 20416 -926 20432 -892
rect 20373 -968 20432 -926
rect 20500 -890 20518 -856
rect 20466 -934 20518 -890
rect 20570 -832 20657 -824
rect 20691 -832 20703 -798
rect 20570 -858 20703 -832
rect 20772 -594 20782 -576
rect 20926 -592 20960 -542
rect 20738 -628 20748 -610
rect 20570 -866 20604 -858
rect 20738 -866 20782 -628
rect 20816 -626 20960 -592
rect 20816 -820 20850 -626
rect 21000 -628 21024 -594
rect 21058 -620 21100 -594
rect 21058 -628 21066 -620
rect 21000 -654 21066 -628
rect 20884 -681 20966 -660
rect 20884 -715 20901 -681
rect 20935 -715 20966 -681
rect 20884 -734 20966 -715
rect 20918 -768 20966 -734
rect 20884 -784 20966 -768
rect 21000 -670 21100 -654
rect 21000 -794 21044 -670
rect 21134 -704 21168 -535
rect 21216 -510 21292 -458
rect 21510 -500 21576 -458
rect 21216 -544 21232 -510
rect 21266 -544 21292 -510
rect 21352 -526 21386 -510
rect 21352 -578 21386 -560
rect 21510 -534 21526 -500
rect 21560 -534 21576 -500
rect 21999 -500 22075 -458
rect 21510 -568 21576 -534
rect 21785 -535 21801 -501
rect 21835 -535 21951 -501
rect 21999 -534 22015 -500
rect 22049 -534 22075 -500
rect 22263 -500 22541 -458
rect 22123 -526 22157 -510
rect 21202 -594 21472 -578
rect 21202 -620 21352 -594
rect 21236 -628 21352 -620
rect 21386 -628 21472 -594
rect 21510 -602 21526 -568
rect 21560 -602 21576 -568
rect 21747 -594 21794 -588
rect 21236 -654 21252 -628
rect 21202 -670 21252 -654
rect 21354 -704 21404 -688
rect 21134 -738 21370 -704
rect 21134 -746 21218 -738
rect 20816 -858 20960 -820
rect 21034 -828 21044 -794
rect 21000 -844 21044 -828
rect 21080 -816 21096 -782
rect 21130 -798 21150 -782
rect 21080 -832 21116 -816
rect 21080 -856 21150 -832
rect 20570 -916 20604 -900
rect 20638 -926 20654 -892
rect 20688 -926 20704 -892
rect 20772 -900 20782 -866
rect 20926 -874 20960 -858
rect 20738 -916 20782 -900
rect 20638 -968 20704 -926
rect 20821 -926 20842 -892
rect 20876 -926 20892 -892
rect 21184 -892 21218 -746
rect 21360 -754 21404 -738
rect 21438 -772 21472 -628
rect 21747 -620 21760 -594
rect 21781 -654 21794 -628
rect 21506 -662 21707 -654
rect 21506 -696 21668 -662
rect 21702 -696 21707 -662
rect 21747 -670 21794 -654
rect 21842 -620 21883 -604
rect 21842 -654 21849 -620
rect 21506 -702 21707 -696
rect 21506 -704 21572 -702
rect 21506 -738 21522 -704
rect 21556 -738 21572 -704
rect 21842 -724 21883 -654
rect 21748 -730 21883 -724
rect 21634 -772 21650 -738
rect 21684 -772 21700 -738
rect 21252 -806 21268 -772
rect 21302 -792 21318 -772
rect 21302 -798 21334 -792
rect 21252 -832 21300 -806
rect 21438 -806 21700 -772
rect 21748 -764 21760 -730
rect 21794 -760 21883 -730
rect 21917 -704 21951 -535
rect 22263 -534 22289 -500
rect 22323 -534 22491 -500
rect 22525 -534 22541 -500
rect 22123 -568 22157 -560
rect 22575 -537 22632 -492
rect 21985 -602 22541 -568
rect 21985 -620 22035 -602
rect 22019 -654 22035 -620
rect 21985 -670 22035 -654
rect 21917 -720 22187 -704
rect 21917 -738 22153 -720
rect 21794 -764 21816 -760
rect 21748 -773 21816 -764
rect 21772 -794 21816 -773
rect 21438 -832 21482 -806
rect 21252 -838 21334 -832
rect 21416 -866 21432 -832
rect 21466 -866 21482 -832
rect 21772 -828 21782 -794
rect 21516 -858 21550 -842
rect 21772 -844 21816 -828
rect 20926 -924 20960 -908
rect 20821 -968 20892 -926
rect 21015 -926 21031 -892
rect 21065 -926 21218 -892
rect 21015 -932 21218 -926
rect 21252 -896 21286 -880
rect 21252 -968 21286 -930
rect 21320 -890 21386 -884
rect 21320 -924 21336 -890
rect 21370 -900 21386 -890
rect 21917 -892 21951 -738
rect 22143 -754 22153 -738
rect 22143 -770 22187 -754
rect 21991 -806 22046 -772
rect 22080 -798 22100 -772
rect 21991 -832 22050 -806
rect 22084 -832 22100 -798
rect 22221 -817 22255 -602
rect 22289 -662 22393 -636
rect 22289 -696 22306 -662
rect 22340 -670 22393 -662
rect 22427 -670 22446 -636
rect 22340 -696 22346 -670
rect 22289 -704 22346 -696
rect 22323 -738 22346 -704
rect 22507 -720 22541 -602
rect 22609 -571 22632 -537
rect 22575 -605 22632 -571
rect 22609 -610 22632 -605
rect 22575 -644 22586 -639
rect 22620 -644 22632 -610
rect 22575 -659 22632 -644
rect 22289 -763 22346 -738
rect 22302 -800 22346 -763
rect 22382 -732 22473 -720
rect 22382 -766 22398 -732
rect 22432 -766 22473 -732
rect 22507 -736 22560 -720
rect 22507 -770 22526 -736
rect 22507 -786 22560 -770
rect 22221 -818 22258 -817
rect 21991 -838 22100 -832
rect 22178 -852 22208 -818
rect 22242 -852 22258 -818
rect 22302 -834 22430 -800
rect 21516 -900 21550 -892
rect 21370 -924 21550 -900
rect 21320 -934 21550 -924
rect 21600 -926 21620 -892
rect 21654 -926 21670 -892
rect 21600 -968 21670 -926
rect 21795 -926 21824 -892
rect 21858 -926 21951 -892
rect 21795 -932 21951 -926
rect 21985 -896 22050 -880
rect 21985 -930 22016 -896
rect 21985 -968 22050 -930
rect 22084 -910 22100 -876
rect 22134 -900 22150 -876
rect 22292 -884 22326 -868
rect 22134 -910 22292 -900
rect 22084 -918 22292 -910
rect 22084 -934 22326 -918
rect 22388 -882 22430 -834
rect 22388 -916 22396 -882
rect 22388 -932 22430 -916
rect 22480 -892 22541 -824
rect 22596 -842 22632 -659
rect 22480 -926 22491 -892
rect 22525 -926 22541 -892
rect 22480 -968 22541 -926
rect 22575 -858 22632 -842
rect 22609 -892 22632 -858
rect 22575 -934 22632 -892
rect 22667 -518 22730 -502
rect 22667 -552 22679 -518
rect 22713 -552 22730 -518
rect 22667 -586 22730 -552
rect 22667 -620 22679 -586
rect 22713 -620 22730 -586
rect 22667 -720 22730 -620
rect 22766 -512 22824 -458
rect 22766 -546 22774 -512
rect 22808 -546 22824 -512
rect 22766 -580 22824 -546
rect 22766 -614 22774 -580
rect 22808 -614 22824 -580
rect 22766 -632 22824 -614
rect 22858 -531 22910 -492
rect 22858 -536 22869 -531
rect 22903 -565 22910 -531
rect 22892 -570 22910 -565
rect 22858 -604 22910 -570
rect 22892 -638 22910 -604
rect 22962 -508 22996 -492
rect 22962 -576 22996 -542
rect 23030 -524 23096 -458
rect 23030 -558 23046 -524
rect 23080 -558 23096 -524
rect 23130 -508 23174 -492
rect 23164 -542 23174 -508
rect 23130 -576 23174 -542
rect 23213 -524 23284 -458
rect 23213 -558 23234 -524
rect 23268 -558 23284 -524
rect 23318 -508 23352 -492
rect 23394 -535 23410 -501
rect 23444 -535 23560 -501
rect 22996 -610 23095 -592
rect 22962 -626 23095 -610
rect 22858 -694 22910 -638
rect 22667 -736 22834 -720
rect 22667 -770 22800 -736
rect 22667 -786 22834 -770
rect 22667 -866 22730 -786
rect 22868 -820 22910 -694
rect 22944 -705 23014 -660
rect 22944 -739 22953 -705
rect 22987 -721 23014 -705
rect 22944 -755 22958 -739
rect 22992 -755 23014 -721
rect 22944 -790 23014 -755
rect 23049 -721 23095 -626
rect 23049 -755 23060 -721
rect 23094 -755 23095 -721
rect 22667 -900 22679 -866
rect 22713 -900 22730 -866
rect 22858 -856 22910 -820
rect 23049 -798 23095 -755
rect 22667 -934 22730 -900
rect 22765 -892 22824 -876
rect 22765 -926 22774 -892
rect 22808 -926 22824 -892
rect 22765 -968 22824 -926
rect 22892 -890 22910 -856
rect 22858 -934 22910 -890
rect 22962 -832 23049 -824
rect 23083 -832 23095 -798
rect 22962 -858 23095 -832
rect 23164 -594 23174 -576
rect 23318 -592 23352 -542
rect 23130 -628 23140 -610
rect 22962 -866 22996 -858
rect 23130 -866 23174 -628
rect 23208 -626 23352 -592
rect 23208 -820 23242 -626
rect 23392 -628 23416 -594
rect 23450 -620 23492 -594
rect 23450 -628 23458 -620
rect 23392 -654 23458 -628
rect 23276 -682 23358 -660
rect 23276 -716 23294 -682
rect 23328 -716 23358 -682
rect 23276 -734 23358 -716
rect 23310 -768 23358 -734
rect 23276 -784 23358 -768
rect 23392 -670 23492 -654
rect 23392 -794 23436 -670
rect 23526 -704 23560 -535
rect 23608 -510 23684 -458
rect 23902 -500 23968 -458
rect 23608 -544 23624 -510
rect 23658 -544 23684 -510
rect 23744 -526 23778 -510
rect 23744 -578 23778 -560
rect 23902 -534 23918 -500
rect 23952 -534 23968 -500
rect 24391 -500 24467 -458
rect 23902 -568 23968 -534
rect 24177 -535 24193 -501
rect 24227 -535 24343 -501
rect 24391 -534 24407 -500
rect 24441 -534 24467 -500
rect 24655 -500 24933 -458
rect 24515 -526 24549 -510
rect 23594 -594 23864 -578
rect 23594 -620 23744 -594
rect 23628 -628 23744 -620
rect 23778 -628 23864 -594
rect 23902 -602 23918 -568
rect 23952 -602 23968 -568
rect 24139 -594 24186 -588
rect 23628 -654 23644 -628
rect 23594 -670 23644 -654
rect 23746 -704 23796 -688
rect 23526 -738 23762 -704
rect 23526 -746 23610 -738
rect 23208 -858 23352 -820
rect 23426 -828 23436 -794
rect 23392 -844 23436 -828
rect 23472 -816 23488 -782
rect 23522 -798 23542 -782
rect 23472 -832 23508 -816
rect 23472 -856 23542 -832
rect 22962 -916 22996 -900
rect 23030 -926 23046 -892
rect 23080 -926 23096 -892
rect 23164 -900 23174 -866
rect 23318 -874 23352 -858
rect 23130 -916 23174 -900
rect 23030 -968 23096 -926
rect 23213 -926 23234 -892
rect 23268 -926 23284 -892
rect 23576 -892 23610 -746
rect 23752 -754 23796 -738
rect 23830 -772 23864 -628
rect 24139 -620 24152 -594
rect 24173 -654 24186 -628
rect 23898 -662 24099 -654
rect 23898 -696 24060 -662
rect 24094 -696 24099 -662
rect 24139 -670 24186 -654
rect 24234 -620 24275 -604
rect 24234 -654 24241 -620
rect 23898 -702 24099 -696
rect 23898 -704 23964 -702
rect 23898 -738 23914 -704
rect 23948 -738 23964 -704
rect 24234 -724 24275 -654
rect 24140 -730 24275 -724
rect 24026 -772 24042 -738
rect 24076 -772 24092 -738
rect 23644 -806 23660 -772
rect 23694 -792 23710 -772
rect 23694 -798 23726 -792
rect 23644 -832 23692 -806
rect 23830 -806 24092 -772
rect 24140 -764 24152 -730
rect 24186 -760 24275 -730
rect 24309 -704 24343 -535
rect 24655 -534 24681 -500
rect 24715 -534 24883 -500
rect 24917 -534 24933 -500
rect 24515 -568 24549 -560
rect 24967 -537 25024 -492
rect 24377 -602 24933 -568
rect 24377 -620 24427 -602
rect 24411 -654 24427 -620
rect 24377 -670 24427 -654
rect 24309 -720 24579 -704
rect 24309 -738 24545 -720
rect 24186 -764 24208 -760
rect 24140 -773 24208 -764
rect 24164 -794 24208 -773
rect 23830 -832 23874 -806
rect 23644 -838 23726 -832
rect 23808 -866 23824 -832
rect 23858 -866 23874 -832
rect 24164 -828 24174 -794
rect 23908 -858 23942 -842
rect 24164 -844 24208 -828
rect 23318 -924 23352 -908
rect 23213 -968 23284 -926
rect 23407 -926 23423 -892
rect 23457 -926 23610 -892
rect 23407 -932 23610 -926
rect 23644 -896 23678 -880
rect 23644 -968 23678 -930
rect 23712 -890 23778 -884
rect 23712 -924 23728 -890
rect 23762 -900 23778 -890
rect 24309 -892 24343 -738
rect 24535 -754 24545 -738
rect 24535 -770 24579 -754
rect 24383 -806 24438 -772
rect 24472 -798 24492 -772
rect 24383 -832 24442 -806
rect 24476 -832 24492 -798
rect 24613 -817 24647 -602
rect 24681 -662 24785 -636
rect 24681 -696 24698 -662
rect 24732 -670 24785 -662
rect 24819 -670 24838 -636
rect 24732 -696 24738 -670
rect 24681 -704 24738 -696
rect 24715 -738 24738 -704
rect 24899 -720 24933 -602
rect 25001 -571 25024 -537
rect 24967 -605 25024 -571
rect 25001 -608 25024 -605
rect 24967 -642 24979 -639
rect 25013 -642 25024 -608
rect 24967 -659 25024 -642
rect 24681 -763 24738 -738
rect 24694 -800 24738 -763
rect 24774 -732 24865 -720
rect 24774 -766 24790 -732
rect 24824 -766 24865 -732
rect 24899 -736 24952 -720
rect 24899 -770 24918 -736
rect 24899 -786 24952 -770
rect 24613 -818 24650 -817
rect 24383 -838 24492 -832
rect 24570 -852 24600 -818
rect 24634 -852 24650 -818
rect 24694 -834 24822 -800
rect 23908 -900 23942 -892
rect 23762 -924 23942 -900
rect 23712 -934 23942 -924
rect 23992 -926 24012 -892
rect 24046 -926 24062 -892
rect 23992 -968 24062 -926
rect 24187 -926 24216 -892
rect 24250 -926 24343 -892
rect 24187 -932 24343 -926
rect 24377 -896 24442 -880
rect 24377 -930 24408 -896
rect 24377 -968 24442 -930
rect 24476 -910 24492 -876
rect 24526 -900 24542 -876
rect 24684 -884 24718 -868
rect 24526 -910 24684 -900
rect 24476 -918 24684 -910
rect 24476 -934 24718 -918
rect 24780 -882 24822 -834
rect 24780 -916 24788 -882
rect 24780 -932 24822 -916
rect 24872 -892 24933 -824
rect 24988 -842 25024 -659
rect 24872 -926 24883 -892
rect 24917 -926 24933 -892
rect 24872 -968 24933 -926
rect 24967 -858 25024 -842
rect 25001 -892 25024 -858
rect 24967 -934 25024 -892
rect 25059 -518 25122 -502
rect 25059 -552 25071 -518
rect 25105 -552 25122 -518
rect 25059 -586 25122 -552
rect 25059 -620 25071 -586
rect 25105 -620 25122 -586
rect 25059 -720 25122 -620
rect 25158 -512 25216 -458
rect 25158 -546 25166 -512
rect 25200 -546 25216 -512
rect 25158 -580 25216 -546
rect 25158 -614 25166 -580
rect 25200 -614 25216 -580
rect 25158 -632 25216 -614
rect 25250 -531 25302 -492
rect 25250 -536 25261 -531
rect 25295 -565 25302 -531
rect 25284 -570 25302 -565
rect 25250 -604 25302 -570
rect 25284 -638 25302 -604
rect 25250 -694 25302 -638
rect 25059 -736 25226 -720
rect 25059 -770 25192 -736
rect 25059 -786 25226 -770
rect 25059 -866 25122 -786
rect 25260 -820 25302 -694
rect 25059 -900 25071 -866
rect 25105 -900 25122 -866
rect 25250 -856 25302 -820
rect 25059 -934 25122 -900
rect 25157 -892 25216 -876
rect 25157 -926 25166 -892
rect 25200 -926 25216 -892
rect 25157 -968 25216 -926
rect 25284 -890 25302 -856
rect 25250 -934 25302 -890
rect 8575 -1026 8604 -968
rect 8638 -1026 8696 -968
rect 8730 -1026 8788 -968
rect 8822 -1026 8880 -968
rect 8914 -1026 8972 -968
rect 9006 -1026 9064 -968
rect 9098 -1026 9156 -968
rect 9190 -1026 9248 -968
rect 9282 -1026 9340 -968
rect 9374 -1026 9432 -968
rect 9466 -1026 9524 -968
rect 9558 -1026 9616 -968
rect 9650 -1026 9708 -968
rect 9742 -1026 9800 -968
rect 9834 -1026 9892 -968
rect 9926 -1026 9984 -968
rect 10018 -1026 10076 -968
rect 10110 -1026 10168 -968
rect 10202 -1026 10260 -968
rect 10294 -1026 10352 -968
rect 10386 -1026 10444 -968
rect 10478 -1026 10536 -968
rect 10570 -1026 10628 -968
rect 10662 -1026 10720 -968
rect 10754 -1026 10812 -968
rect 10846 -1026 10904 -968
rect 10938 -1026 10996 -968
rect 11030 -1026 11088 -968
rect 11122 -1026 11180 -968
rect 11214 -1026 11272 -968
rect 11306 -1026 11364 -968
rect 11398 -1026 11456 -968
rect 11490 -1026 11548 -968
rect 11582 -1026 11640 -968
rect 11674 -1026 11732 -968
rect 11766 -1026 11824 -968
rect 11858 -1026 11916 -968
rect 11950 -1026 12008 -968
rect 12042 -1026 12100 -968
rect 12134 -1026 12192 -968
rect 12226 -1026 12284 -968
rect 12318 -1026 12376 -968
rect 12410 -1026 12468 -968
rect 12502 -1026 12560 -968
rect 12594 -1026 12652 -968
rect 12686 -1026 12744 -968
rect 12778 -1026 12836 -968
rect 12870 -1026 12928 -968
rect 12962 -1026 13020 -968
rect 13054 -1026 13112 -968
rect 13146 -1026 13204 -968
rect 13238 -1026 13296 -968
rect 13330 -1026 13388 -968
rect 13422 -1026 13480 -968
rect 13514 -1026 13572 -968
rect 13606 -1026 13664 -968
rect 13698 -1026 13756 -968
rect 13790 -1026 13848 -968
rect 13882 -1026 13940 -968
rect 13974 -1026 14032 -968
rect 14066 -1026 14124 -968
rect 14158 -1026 14216 -968
rect 14250 -1026 14308 -968
rect 14342 -1026 14400 -968
rect 14434 -1026 14492 -968
rect 14526 -1026 14584 -968
rect 14618 -1026 14676 -968
rect 14710 -1026 14768 -968
rect 14802 -1026 14860 -968
rect 14894 -1026 14952 -968
rect 14986 -1026 15044 -968
rect 15078 -1026 15136 -968
rect 15170 -1026 15228 -968
rect 15262 -1026 15320 -968
rect 15354 -1026 15412 -968
rect 15446 -1026 15504 -968
rect 15538 -1026 15596 -968
rect 15630 -1026 15688 -968
rect 15722 -1026 15780 -968
rect 15814 -1026 15872 -968
rect 15906 -1026 15964 -968
rect 15998 -1026 16056 -968
rect 16090 -1026 16148 -968
rect 16182 -1026 16240 -968
rect 16274 -1026 16332 -968
rect 16366 -1026 16424 -968
rect 16458 -1026 16516 -968
rect 16550 -1026 16608 -968
rect 16642 -1026 16700 -968
rect 16734 -1026 16792 -968
rect 16826 -1026 16884 -968
rect 16918 -1026 16976 -968
rect 17010 -1026 17068 -968
rect 17102 -1026 17160 -968
rect 17194 -1026 17252 -968
rect 17286 -1026 17344 -968
rect 17378 -1026 17436 -968
rect 17470 -1026 17528 -968
rect 17562 -1026 17620 -968
rect 17654 -1026 17712 -968
rect 17746 -1026 17804 -968
rect 17838 -1026 17896 -968
rect 17930 -1026 17988 -968
rect 18022 -1026 18080 -968
rect 18114 -1026 18172 -968
rect 18206 -1026 18264 -968
rect 18298 -1026 18356 -968
rect 18390 -1026 18448 -968
rect 18482 -1026 18540 -968
rect 18574 -1026 18632 -968
rect 18666 -1026 18724 -968
rect 18758 -1026 18816 -968
rect 18850 -1026 18908 -968
rect 18942 -1026 19000 -968
rect 19034 -1026 19092 -968
rect 19126 -1026 19184 -968
rect 19218 -1026 19276 -968
rect 19310 -1026 19368 -968
rect 19402 -1026 19460 -968
rect 19494 -1026 19552 -968
rect 19586 -1026 19644 -968
rect 19678 -1026 19736 -968
rect 19770 -1026 19828 -968
rect 19862 -1026 19920 -968
rect 19954 -1026 20012 -968
rect 20046 -1026 20104 -968
rect 20138 -1026 20196 -968
rect 20230 -1026 20288 -968
rect 20322 -1026 20380 -968
rect 20414 -1026 20472 -968
rect 20506 -1026 20564 -968
rect 20598 -1026 20656 -968
rect 20690 -1026 20748 -968
rect 20782 -1026 20840 -968
rect 20874 -1026 20932 -968
rect 20966 -1026 21024 -968
rect 21058 -1026 21116 -968
rect 21150 -1026 21208 -968
rect 21242 -1026 21300 -968
rect 21334 -1026 21392 -968
rect 21426 -1026 21484 -968
rect 21518 -1026 21576 -968
rect 21610 -1026 21668 -968
rect 21702 -1026 21760 -968
rect 21794 -1026 21852 -968
rect 21886 -1026 21944 -968
rect 21978 -1026 22036 -968
rect 22070 -1026 22128 -968
rect 22162 -1026 22220 -968
rect 22254 -1026 22312 -968
rect 22346 -1026 22404 -968
rect 22438 -1026 22496 -968
rect 22530 -1026 22588 -968
rect 22622 -1026 22680 -968
rect 22714 -1026 22772 -968
rect 22806 -1026 22864 -968
rect 22898 -1026 22956 -968
rect 22990 -1026 23048 -968
rect 23082 -1026 23140 -968
rect 23174 -1026 23232 -968
rect 23266 -1026 23324 -968
rect 23358 -1026 23416 -968
rect 23450 -1026 23508 -968
rect 23542 -1026 23600 -968
rect 23634 -1026 23692 -968
rect 23726 -1026 23784 -968
rect 23818 -1026 23876 -968
rect 23910 -1026 23968 -968
rect 24002 -1026 24060 -968
rect 24094 -1026 24152 -968
rect 24186 -1026 24244 -968
rect 24278 -1026 24336 -968
rect 24370 -1026 24428 -968
rect 24462 -1026 24520 -968
rect 24554 -1026 24612 -968
rect 24646 -1026 24704 -968
rect 24738 -1026 24796 -968
rect 24830 -1026 24888 -968
rect 24922 -1026 24980 -968
rect 25014 -1026 25072 -968
rect 25106 -1026 25164 -968
rect 25198 -1026 25256 -968
rect 25290 -1026 25319 -968
rect 8575 -1089 9146 -1088
rect 8575 -1147 8604 -1089
rect 8638 -1147 8696 -1089
rect 8730 -1147 8788 -1089
rect 8822 -1147 8880 -1089
rect 8914 -1123 8969 -1089
rect 9003 -1113 9071 -1089
rect 8914 -1147 8972 -1123
rect 9006 -1147 9064 -1113
rect 9105 -1123 9156 -1089
rect 9098 -1147 9156 -1123
rect 9190 -1147 9248 -1089
rect 9282 -1147 9340 -1089
rect 9374 -1147 9432 -1089
rect 9466 -1147 9524 -1089
rect 9558 -1147 9616 -1089
rect 9650 -1147 9708 -1089
rect 9742 -1147 9800 -1089
rect 9834 -1147 9892 -1089
rect 9926 -1147 9984 -1089
rect 10018 -1147 10076 -1089
rect 10110 -1093 10352 -1089
rect 10110 -1113 10182 -1093
rect 10216 -1113 10352 -1093
rect 10110 -1147 10168 -1113
rect 10216 -1127 10260 -1113
rect 10202 -1147 10260 -1127
rect 10294 -1147 10352 -1113
rect 10386 -1147 10444 -1089
rect 10478 -1147 10536 -1089
rect 10570 -1147 10628 -1089
rect 10662 -1147 10720 -1089
rect 10754 -1147 10812 -1089
rect 10846 -1147 10904 -1089
rect 10938 -1147 10996 -1089
rect 11030 -1147 11088 -1089
rect 11122 -1147 11180 -1089
rect 11214 -1147 11272 -1089
rect 11306 -1113 11366 -1089
rect 11400 -1113 11457 -1089
rect 11306 -1147 11364 -1113
rect 11400 -1123 11456 -1113
rect 11491 -1123 11548 -1089
rect 11398 -1147 11456 -1123
rect 11490 -1147 11548 -1123
rect 11582 -1147 11640 -1089
rect 11674 -1147 11732 -1089
rect 11766 -1147 11824 -1089
rect 11858 -1147 11916 -1089
rect 11950 -1147 12008 -1089
rect 12042 -1147 12100 -1089
rect 12134 -1147 12192 -1089
rect 12226 -1147 12284 -1089
rect 12318 -1147 12376 -1089
rect 12410 -1147 12468 -1089
rect 12502 -1093 12744 -1089
rect 12502 -1113 12574 -1093
rect 12608 -1113 12744 -1093
rect 12502 -1147 12560 -1113
rect 12608 -1127 12652 -1113
rect 12594 -1147 12652 -1127
rect 12686 -1147 12744 -1113
rect 12778 -1147 12836 -1089
rect 12870 -1147 12928 -1089
rect 12962 -1147 13020 -1089
rect 13054 -1147 13112 -1089
rect 13146 -1147 13204 -1089
rect 13238 -1147 13296 -1089
rect 13330 -1147 13388 -1089
rect 13422 -1147 13480 -1089
rect 13514 -1147 13572 -1089
rect 13606 -1147 13664 -1089
rect 13698 -1123 13754 -1089
rect 13788 -1113 13848 -1089
rect 13698 -1147 13756 -1123
rect 13790 -1147 13848 -1113
rect 13882 -1147 13940 -1089
rect 13974 -1147 14032 -1089
rect 14066 -1147 14124 -1089
rect 14158 -1147 14216 -1089
rect 14250 -1147 14308 -1089
rect 14342 -1147 14400 -1089
rect 14434 -1147 14492 -1089
rect 14526 -1147 14584 -1089
rect 14618 -1147 14676 -1089
rect 14710 -1147 14768 -1089
rect 14802 -1147 14860 -1089
rect 14894 -1093 15136 -1089
rect 14894 -1113 14966 -1093
rect 15000 -1113 15136 -1093
rect 14894 -1147 14952 -1113
rect 15000 -1127 15044 -1113
rect 14986 -1147 15044 -1127
rect 15078 -1147 15136 -1113
rect 15170 -1147 15228 -1089
rect 15262 -1147 15320 -1089
rect 15354 -1147 15412 -1089
rect 15446 -1147 15504 -1089
rect 15538 -1147 15596 -1089
rect 15630 -1147 15688 -1089
rect 15722 -1147 15780 -1089
rect 15814 -1147 15872 -1089
rect 15906 -1147 15964 -1089
rect 15998 -1147 16056 -1089
rect 16090 -1113 16149 -1089
rect 16090 -1147 16148 -1113
rect 16183 -1123 16240 -1089
rect 16182 -1147 16240 -1123
rect 16274 -1147 16332 -1089
rect 16366 -1147 16424 -1089
rect 16458 -1147 16516 -1089
rect 16550 -1147 16608 -1089
rect 16642 -1147 16700 -1089
rect 16734 -1147 16792 -1089
rect 16826 -1147 16884 -1089
rect 16918 -1147 16976 -1089
rect 17010 -1147 17068 -1089
rect 17102 -1147 17160 -1089
rect 17194 -1147 17252 -1089
rect 17286 -1093 17528 -1089
rect 17286 -1113 17358 -1093
rect 17392 -1113 17528 -1093
rect 17286 -1147 17344 -1113
rect 17392 -1127 17436 -1113
rect 17378 -1147 17436 -1127
rect 17470 -1147 17528 -1113
rect 17562 -1147 17620 -1089
rect 17654 -1147 17712 -1089
rect 17746 -1147 17804 -1089
rect 17838 -1147 17896 -1089
rect 17930 -1147 17988 -1089
rect 18022 -1147 18080 -1089
rect 18114 -1147 18172 -1089
rect 18206 -1147 18264 -1089
rect 18298 -1147 18356 -1089
rect 18390 -1147 18448 -1089
rect 18482 -1123 18538 -1089
rect 18572 -1113 18633 -1089
rect 18482 -1147 18540 -1123
rect 18574 -1147 18632 -1113
rect 18667 -1123 18724 -1089
rect 18666 -1147 18724 -1123
rect 18758 -1147 18816 -1089
rect 18850 -1147 18908 -1089
rect 18942 -1147 19000 -1089
rect 19034 -1147 19092 -1089
rect 19126 -1147 19184 -1089
rect 19218 -1147 19276 -1089
rect 19310 -1147 19368 -1089
rect 19402 -1147 19460 -1089
rect 19494 -1147 19552 -1089
rect 19586 -1147 19644 -1089
rect 19678 -1093 19920 -1089
rect 19678 -1113 19750 -1093
rect 19784 -1113 19920 -1093
rect 19678 -1147 19736 -1113
rect 19784 -1127 19828 -1113
rect 19770 -1147 19828 -1127
rect 19862 -1147 19920 -1113
rect 19954 -1147 20012 -1089
rect 20046 -1147 20104 -1089
rect 20138 -1147 20196 -1089
rect 20230 -1147 20288 -1089
rect 20322 -1147 20380 -1089
rect 20414 -1147 20472 -1089
rect 20506 -1147 20564 -1089
rect 20598 -1147 20656 -1089
rect 20690 -1147 20748 -1089
rect 20782 -1147 20840 -1089
rect 20874 -1147 20932 -1089
rect 20966 -1123 21023 -1089
rect 21057 -1113 21116 -1089
rect 20966 -1147 21024 -1123
rect 21058 -1147 21116 -1113
rect 21150 -1147 21208 -1089
rect 21242 -1147 21300 -1089
rect 21334 -1147 21392 -1089
rect 21426 -1147 21484 -1089
rect 21518 -1147 21576 -1089
rect 21610 -1147 21668 -1089
rect 21702 -1147 21760 -1089
rect 21794 -1147 21852 -1089
rect 21886 -1147 21944 -1089
rect 21978 -1147 22036 -1089
rect 22070 -1093 22312 -1089
rect 22070 -1113 22142 -1093
rect 22176 -1113 22312 -1093
rect 22070 -1147 22128 -1113
rect 22176 -1127 22220 -1113
rect 22162 -1147 22220 -1127
rect 22254 -1147 22312 -1113
rect 22346 -1147 22404 -1089
rect 22438 -1147 22496 -1089
rect 22530 -1147 22588 -1089
rect 22622 -1147 22680 -1089
rect 22714 -1147 22772 -1089
rect 22806 -1147 22864 -1089
rect 22898 -1147 22956 -1089
rect 22990 -1147 23048 -1089
rect 23082 -1147 23140 -1089
rect 23174 -1147 23232 -1089
rect 23266 -1123 23323 -1089
rect 23357 -1113 23417 -1089
rect 23266 -1147 23324 -1123
rect 23358 -1147 23416 -1113
rect 23451 -1123 23508 -1089
rect 23450 -1147 23508 -1123
rect 23542 -1147 23600 -1089
rect 23634 -1147 23692 -1089
rect 23726 -1147 23784 -1089
rect 23818 -1147 23876 -1089
rect 23910 -1147 23968 -1089
rect 24002 -1147 24060 -1089
rect 24094 -1147 24152 -1089
rect 24186 -1147 24244 -1089
rect 24278 -1147 24336 -1089
rect 24370 -1147 24428 -1089
rect 24462 -1096 24704 -1089
rect 24462 -1113 24534 -1096
rect 24568 -1113 24704 -1096
rect 24462 -1147 24520 -1113
rect 24568 -1130 24612 -1113
rect 24554 -1147 24612 -1130
rect 24646 -1147 24704 -1113
rect 24738 -1147 24796 -1089
rect 24830 -1147 24888 -1089
rect 24922 -1147 24980 -1089
rect 25014 -1147 25072 -1089
rect 25106 -1147 25164 -1089
rect 25198 -1147 25256 -1089
rect 25290 -1147 25319 -1089
rect 8592 -1223 8644 -1181
rect 8592 -1257 8601 -1223
rect 8635 -1225 8644 -1223
rect 8592 -1259 8610 -1257
rect 8592 -1293 8644 -1259
rect 8592 -1327 8610 -1293
rect 8678 -1201 8736 -1147
rect 8678 -1235 8694 -1201
rect 8728 -1235 8736 -1201
rect 8678 -1269 8736 -1235
rect 8678 -1303 8694 -1269
rect 8728 -1303 8736 -1269
rect 8678 -1321 8736 -1303
rect 8772 -1207 8835 -1191
rect 8772 -1241 8789 -1207
rect 8823 -1241 8835 -1207
rect 8772 -1275 8835 -1241
rect 8772 -1309 8789 -1275
rect 8823 -1309 8835 -1275
rect 8592 -1383 8644 -1327
rect 8592 -1509 8634 -1383
rect 8772 -1409 8835 -1309
rect 8668 -1425 8835 -1409
rect 8702 -1459 8835 -1425
rect 8668 -1475 8835 -1459
rect 8592 -1545 8644 -1509
rect 8592 -1579 8610 -1545
rect 8772 -1555 8835 -1475
rect 8592 -1623 8644 -1579
rect 8678 -1581 8737 -1565
rect 8678 -1615 8694 -1581
rect 8728 -1615 8737 -1581
rect 8678 -1657 8737 -1615
rect 8772 -1589 8789 -1555
rect 8823 -1589 8835 -1555
rect 8772 -1623 8835 -1589
rect 8870 -1226 8927 -1181
rect 8961 -1189 9239 -1147
rect 8961 -1223 8977 -1189
rect 9011 -1223 9179 -1189
rect 9213 -1223 9239 -1189
rect 9427 -1189 9503 -1147
rect 9345 -1215 9379 -1199
rect 8870 -1260 8893 -1226
rect 9427 -1223 9453 -1189
rect 9487 -1223 9503 -1189
rect 9926 -1189 9992 -1147
rect 9345 -1257 9379 -1249
rect 9551 -1224 9667 -1190
rect 9701 -1224 9717 -1190
rect 9926 -1223 9942 -1189
rect 9976 -1223 9992 -1189
rect 10210 -1199 10286 -1147
rect 8870 -1289 8927 -1260
rect 8870 -1323 8881 -1289
rect 8915 -1294 8927 -1289
rect 8870 -1328 8893 -1323
rect 8870 -1348 8927 -1328
rect 8961 -1291 9517 -1257
rect 8870 -1531 8906 -1348
rect 8961 -1409 8995 -1291
rect 9056 -1359 9075 -1325
rect 9109 -1351 9213 -1325
rect 9109 -1359 9162 -1351
rect 9156 -1385 9162 -1359
rect 9196 -1385 9213 -1351
rect 9156 -1393 9213 -1385
rect 8942 -1425 8995 -1409
rect 8976 -1459 8995 -1425
rect 9029 -1417 9120 -1409
rect 9029 -1421 9077 -1417
rect 9029 -1455 9070 -1421
rect 9111 -1451 9120 -1417
rect 9104 -1455 9120 -1451
rect 9156 -1427 9179 -1393
rect 9156 -1452 9213 -1427
rect 8942 -1475 8995 -1459
rect 9156 -1489 9200 -1452
rect 8870 -1547 8927 -1531
rect 8870 -1581 8893 -1547
rect 8870 -1623 8927 -1581
rect 8961 -1581 9022 -1513
rect 8961 -1615 8977 -1581
rect 9011 -1615 9022 -1581
rect 8961 -1657 9022 -1615
rect 9072 -1523 9200 -1489
rect 9247 -1506 9281 -1291
rect 9467 -1309 9517 -1291
rect 9467 -1343 9483 -1309
rect 9467 -1359 9517 -1343
rect 9551 -1393 9585 -1224
rect 9926 -1257 9992 -1223
rect 9708 -1283 9755 -1277
rect 9315 -1409 9585 -1393
rect 9349 -1427 9585 -1409
rect 9349 -1443 9359 -1427
rect 9315 -1459 9359 -1443
rect 9244 -1507 9281 -1506
rect 9402 -1487 9422 -1461
rect 9072 -1571 9114 -1523
rect 9244 -1541 9260 -1507
rect 9294 -1541 9324 -1507
rect 9402 -1521 9418 -1487
rect 9456 -1495 9511 -1461
rect 9452 -1521 9511 -1495
rect 9402 -1527 9511 -1521
rect 9106 -1605 9114 -1571
rect 9072 -1621 9114 -1605
rect 9176 -1573 9210 -1557
rect 9352 -1589 9368 -1565
rect 9210 -1599 9368 -1589
rect 9402 -1599 9418 -1565
rect 9210 -1607 9418 -1599
rect 9176 -1623 9418 -1607
rect 9452 -1585 9517 -1569
rect 9486 -1619 9517 -1585
rect 9452 -1657 9517 -1619
rect 9551 -1581 9585 -1427
rect 9619 -1309 9660 -1293
rect 9653 -1343 9660 -1309
rect 9619 -1413 9660 -1343
rect 9742 -1309 9755 -1283
rect 9926 -1291 9942 -1257
rect 9976 -1291 9992 -1257
rect 10116 -1215 10150 -1199
rect 10210 -1233 10236 -1199
rect 10270 -1233 10286 -1199
rect 10334 -1224 10450 -1190
rect 10484 -1224 10500 -1190
rect 10542 -1197 10576 -1181
rect 10116 -1267 10150 -1249
rect 10030 -1283 10300 -1267
rect 9708 -1343 9721 -1317
rect 10030 -1317 10116 -1283
rect 10150 -1309 10300 -1283
rect 10150 -1317 10266 -1309
rect 9708 -1359 9755 -1343
rect 9795 -1351 9996 -1343
rect 9795 -1385 9800 -1351
rect 9834 -1385 9996 -1351
rect 9795 -1391 9996 -1385
rect 9930 -1393 9996 -1391
rect 9619 -1419 9754 -1413
rect 9619 -1449 9708 -1419
rect 9686 -1453 9708 -1449
rect 9742 -1453 9754 -1419
rect 9930 -1427 9946 -1393
rect 9980 -1427 9996 -1393
rect 9686 -1462 9754 -1453
rect 9802 -1461 9818 -1427
rect 9852 -1461 9868 -1427
rect 10030 -1461 10064 -1317
rect 10250 -1343 10266 -1317
rect 10250 -1359 10300 -1343
rect 10098 -1393 10148 -1377
rect 10334 -1393 10368 -1224
rect 10542 -1281 10576 -1231
rect 10610 -1213 10681 -1147
rect 10610 -1247 10626 -1213
rect 10660 -1247 10681 -1213
rect 10720 -1197 10764 -1181
rect 10720 -1231 10730 -1197
rect 10720 -1265 10764 -1231
rect 10798 -1213 10864 -1147
rect 10798 -1247 10814 -1213
rect 10848 -1247 10864 -1213
rect 10898 -1197 10932 -1181
rect 10402 -1309 10444 -1283
rect 10436 -1317 10444 -1309
rect 10478 -1317 10502 -1283
rect 10542 -1315 10686 -1281
rect 10436 -1343 10502 -1317
rect 10402 -1359 10502 -1343
rect 10132 -1427 10368 -1393
rect 10098 -1443 10142 -1427
rect 10284 -1435 10368 -1427
rect 9686 -1483 9730 -1462
rect 9720 -1517 9730 -1483
rect 9802 -1495 10064 -1461
rect 10184 -1481 10200 -1461
rect 9686 -1533 9730 -1517
rect 10020 -1521 10064 -1495
rect 10168 -1487 10200 -1481
rect 10234 -1495 10250 -1461
rect 10202 -1521 10250 -1495
rect 9952 -1547 9986 -1531
rect 10020 -1555 10036 -1521
rect 10070 -1555 10086 -1521
rect 10168 -1527 10250 -1521
rect 9551 -1615 9644 -1581
rect 9678 -1615 9707 -1581
rect 9551 -1621 9707 -1615
rect 9832 -1615 9848 -1581
rect 9882 -1615 9902 -1581
rect 9832 -1657 9902 -1615
rect 9952 -1589 9986 -1581
rect 10116 -1579 10182 -1573
rect 10116 -1589 10132 -1579
rect 9952 -1613 10132 -1589
rect 10166 -1613 10182 -1579
rect 9952 -1623 10182 -1613
rect 10216 -1585 10250 -1569
rect 10216 -1657 10250 -1619
rect 10284 -1581 10318 -1435
rect 10352 -1487 10372 -1471
rect 10406 -1505 10422 -1471
rect 10386 -1521 10422 -1505
rect 10352 -1545 10422 -1521
rect 10458 -1483 10502 -1359
rect 10536 -1416 10618 -1349
rect 10536 -1450 10543 -1416
rect 10577 -1423 10618 -1416
rect 10577 -1450 10584 -1423
rect 10536 -1457 10584 -1450
rect 10536 -1473 10618 -1457
rect 10458 -1517 10468 -1483
rect 10652 -1509 10686 -1315
rect 10458 -1533 10502 -1517
rect 10542 -1547 10686 -1509
rect 10720 -1283 10730 -1265
rect 10898 -1265 10932 -1231
rect 10754 -1317 10764 -1299
rect 10542 -1563 10576 -1547
rect 10284 -1615 10437 -1581
rect 10471 -1615 10487 -1581
rect 10720 -1555 10764 -1317
rect 10799 -1299 10898 -1281
rect 10799 -1315 10932 -1299
rect 10984 -1223 11036 -1181
rect 10984 -1257 10993 -1223
rect 11027 -1225 11036 -1223
rect 10984 -1259 11002 -1257
rect 10984 -1293 11036 -1259
rect 10799 -1410 10845 -1315
rect 10984 -1327 11002 -1293
rect 11070 -1201 11128 -1147
rect 11070 -1235 11086 -1201
rect 11120 -1235 11128 -1201
rect 11070 -1269 11128 -1235
rect 11070 -1303 11086 -1269
rect 11120 -1303 11128 -1269
rect 11070 -1321 11128 -1303
rect 11164 -1207 11227 -1191
rect 11164 -1241 11181 -1207
rect 11215 -1241 11227 -1207
rect 11164 -1275 11227 -1241
rect 11164 -1309 11181 -1275
rect 11215 -1309 11227 -1275
rect 10799 -1444 10800 -1410
rect 10834 -1444 10845 -1410
rect 10799 -1487 10845 -1444
rect 10880 -1360 10950 -1349
rect 10880 -1394 10889 -1360
rect 10923 -1394 10950 -1360
rect 10880 -1410 10950 -1394
rect 10880 -1444 10902 -1410
rect 10936 -1444 10950 -1410
rect 10880 -1479 10950 -1444
rect 10984 -1383 11036 -1327
rect 10799 -1521 10811 -1487
rect 10984 -1509 11026 -1383
rect 11164 -1409 11227 -1309
rect 11060 -1425 11227 -1409
rect 11094 -1459 11227 -1425
rect 11060 -1475 11227 -1459
rect 10845 -1521 10932 -1513
rect 10799 -1547 10932 -1521
rect 10542 -1613 10576 -1597
rect 10284 -1621 10487 -1615
rect 10610 -1615 10626 -1581
rect 10660 -1615 10681 -1581
rect 10720 -1589 10730 -1555
rect 10898 -1555 10932 -1547
rect 10720 -1605 10764 -1589
rect 10610 -1657 10681 -1615
rect 10798 -1615 10814 -1581
rect 10848 -1615 10864 -1581
rect 10898 -1605 10932 -1589
rect 10984 -1545 11036 -1509
rect 10984 -1579 11002 -1545
rect 11164 -1555 11227 -1475
rect 10798 -1657 10864 -1615
rect 10984 -1623 11036 -1579
rect 11070 -1581 11129 -1565
rect 11070 -1615 11086 -1581
rect 11120 -1615 11129 -1581
rect 11070 -1657 11129 -1615
rect 11164 -1589 11181 -1555
rect 11215 -1589 11227 -1555
rect 11164 -1623 11227 -1589
rect 11262 -1226 11319 -1181
rect 11353 -1189 11631 -1147
rect 11353 -1223 11369 -1189
rect 11403 -1223 11571 -1189
rect 11605 -1223 11631 -1189
rect 11819 -1189 11895 -1147
rect 11737 -1215 11771 -1199
rect 11262 -1260 11285 -1226
rect 11819 -1223 11845 -1189
rect 11879 -1223 11895 -1189
rect 12318 -1189 12384 -1147
rect 11737 -1257 11771 -1249
rect 11943 -1224 12059 -1190
rect 12093 -1224 12109 -1190
rect 12318 -1223 12334 -1189
rect 12368 -1223 12384 -1189
rect 12602 -1199 12678 -1147
rect 11262 -1289 11319 -1260
rect 11262 -1323 11273 -1289
rect 11307 -1294 11319 -1289
rect 11262 -1328 11285 -1323
rect 11262 -1348 11319 -1328
rect 11353 -1291 11909 -1257
rect 11262 -1531 11298 -1348
rect 11353 -1409 11387 -1291
rect 11448 -1359 11467 -1325
rect 11501 -1351 11605 -1325
rect 11501 -1359 11554 -1351
rect 11548 -1385 11554 -1359
rect 11588 -1385 11605 -1351
rect 11548 -1393 11605 -1385
rect 11334 -1425 11387 -1409
rect 11368 -1459 11387 -1425
rect 11421 -1415 11512 -1409
rect 11421 -1421 11466 -1415
rect 11421 -1455 11462 -1421
rect 11500 -1449 11512 -1415
rect 11496 -1455 11512 -1449
rect 11548 -1427 11571 -1393
rect 11548 -1452 11605 -1427
rect 11334 -1475 11387 -1459
rect 11548 -1489 11592 -1452
rect 11262 -1547 11319 -1531
rect 11262 -1581 11285 -1547
rect 11262 -1623 11319 -1581
rect 11353 -1581 11414 -1513
rect 11353 -1615 11369 -1581
rect 11403 -1615 11414 -1581
rect 11353 -1657 11414 -1615
rect 11464 -1523 11592 -1489
rect 11639 -1506 11673 -1291
rect 11859 -1309 11909 -1291
rect 11859 -1343 11875 -1309
rect 11859 -1359 11909 -1343
rect 11943 -1393 11977 -1224
rect 12318 -1257 12384 -1223
rect 12100 -1283 12147 -1277
rect 11707 -1409 11977 -1393
rect 11741 -1427 11977 -1409
rect 11741 -1443 11751 -1427
rect 11707 -1459 11751 -1443
rect 11636 -1507 11673 -1506
rect 11794 -1487 11814 -1461
rect 11464 -1571 11506 -1523
rect 11636 -1541 11652 -1507
rect 11686 -1541 11716 -1507
rect 11794 -1521 11810 -1487
rect 11848 -1495 11903 -1461
rect 11844 -1521 11903 -1495
rect 11794 -1527 11903 -1521
rect 11498 -1605 11506 -1571
rect 11464 -1621 11506 -1605
rect 11568 -1573 11602 -1557
rect 11744 -1589 11760 -1565
rect 11602 -1599 11760 -1589
rect 11794 -1599 11810 -1565
rect 11602 -1607 11810 -1599
rect 11568 -1623 11810 -1607
rect 11844 -1585 11909 -1569
rect 11878 -1619 11909 -1585
rect 11844 -1657 11909 -1619
rect 11943 -1581 11977 -1427
rect 12011 -1309 12052 -1293
rect 12045 -1343 12052 -1309
rect 12011 -1413 12052 -1343
rect 12134 -1309 12147 -1283
rect 12318 -1291 12334 -1257
rect 12368 -1291 12384 -1257
rect 12508 -1215 12542 -1199
rect 12602 -1233 12628 -1199
rect 12662 -1233 12678 -1199
rect 12726 -1224 12842 -1190
rect 12876 -1224 12892 -1190
rect 12934 -1197 12968 -1181
rect 12508 -1267 12542 -1249
rect 12422 -1283 12692 -1267
rect 12100 -1343 12113 -1317
rect 12422 -1317 12508 -1283
rect 12542 -1309 12692 -1283
rect 12542 -1317 12658 -1309
rect 12100 -1359 12147 -1343
rect 12187 -1351 12388 -1343
rect 12187 -1385 12192 -1351
rect 12226 -1385 12388 -1351
rect 12187 -1391 12388 -1385
rect 12322 -1393 12388 -1391
rect 12011 -1419 12146 -1413
rect 12011 -1449 12100 -1419
rect 12078 -1453 12100 -1449
rect 12134 -1453 12146 -1419
rect 12322 -1427 12338 -1393
rect 12372 -1427 12388 -1393
rect 12078 -1462 12146 -1453
rect 12194 -1461 12210 -1427
rect 12244 -1461 12260 -1427
rect 12422 -1461 12456 -1317
rect 12642 -1343 12658 -1317
rect 12642 -1359 12692 -1343
rect 12490 -1393 12540 -1377
rect 12726 -1393 12760 -1224
rect 12934 -1281 12968 -1231
rect 13002 -1213 13073 -1147
rect 13002 -1247 13018 -1213
rect 13052 -1247 13073 -1213
rect 13112 -1197 13156 -1181
rect 13112 -1231 13122 -1197
rect 13112 -1265 13156 -1231
rect 13190 -1213 13256 -1147
rect 13190 -1247 13206 -1213
rect 13240 -1247 13256 -1213
rect 13290 -1197 13324 -1181
rect 12794 -1309 12836 -1283
rect 12828 -1317 12836 -1309
rect 12870 -1317 12894 -1283
rect 12934 -1315 13078 -1281
rect 12828 -1343 12894 -1317
rect 12794 -1359 12894 -1343
rect 12524 -1427 12760 -1393
rect 12490 -1443 12534 -1427
rect 12676 -1435 12760 -1427
rect 12078 -1483 12122 -1462
rect 12112 -1517 12122 -1483
rect 12194 -1495 12456 -1461
rect 12576 -1481 12592 -1461
rect 12078 -1533 12122 -1517
rect 12412 -1521 12456 -1495
rect 12560 -1487 12592 -1481
rect 12626 -1495 12642 -1461
rect 12594 -1521 12642 -1495
rect 12344 -1547 12378 -1531
rect 12412 -1555 12428 -1521
rect 12462 -1555 12478 -1521
rect 12560 -1527 12642 -1521
rect 11943 -1615 12036 -1581
rect 12070 -1615 12099 -1581
rect 11943 -1621 12099 -1615
rect 12224 -1615 12240 -1581
rect 12274 -1615 12294 -1581
rect 12224 -1657 12294 -1615
rect 12344 -1589 12378 -1581
rect 12508 -1579 12574 -1573
rect 12508 -1589 12524 -1579
rect 12344 -1613 12524 -1589
rect 12558 -1613 12574 -1579
rect 12344 -1623 12574 -1613
rect 12608 -1585 12642 -1569
rect 12608 -1657 12642 -1619
rect 12676 -1581 12710 -1435
rect 12744 -1487 12764 -1471
rect 12798 -1505 12814 -1471
rect 12778 -1521 12814 -1505
rect 12744 -1545 12814 -1521
rect 12850 -1483 12894 -1359
rect 12928 -1416 13010 -1349
rect 12928 -1450 12935 -1416
rect 12969 -1423 13010 -1416
rect 12969 -1450 12976 -1423
rect 12928 -1457 12976 -1450
rect 12928 -1473 13010 -1457
rect 12850 -1517 12860 -1483
rect 13044 -1509 13078 -1315
rect 12850 -1533 12894 -1517
rect 12934 -1547 13078 -1509
rect 13112 -1283 13122 -1265
rect 13290 -1265 13324 -1231
rect 13146 -1317 13156 -1299
rect 12934 -1563 12968 -1547
rect 12676 -1615 12829 -1581
rect 12863 -1615 12879 -1581
rect 13112 -1555 13156 -1317
rect 13191 -1299 13290 -1281
rect 13191 -1315 13324 -1299
rect 13376 -1223 13428 -1181
rect 13376 -1257 13386 -1223
rect 13420 -1225 13428 -1223
rect 13376 -1259 13394 -1257
rect 13376 -1293 13428 -1259
rect 13191 -1410 13237 -1315
rect 13376 -1327 13394 -1293
rect 13462 -1201 13520 -1147
rect 13462 -1235 13478 -1201
rect 13512 -1235 13520 -1201
rect 13462 -1269 13520 -1235
rect 13462 -1303 13478 -1269
rect 13512 -1303 13520 -1269
rect 13462 -1321 13520 -1303
rect 13556 -1207 13619 -1191
rect 13556 -1241 13573 -1207
rect 13607 -1241 13619 -1207
rect 13556 -1275 13619 -1241
rect 13556 -1309 13573 -1275
rect 13607 -1309 13619 -1275
rect 13191 -1444 13192 -1410
rect 13226 -1444 13237 -1410
rect 13191 -1487 13237 -1444
rect 13272 -1360 13342 -1349
rect 13272 -1394 13283 -1360
rect 13317 -1394 13342 -1360
rect 13272 -1410 13342 -1394
rect 13272 -1444 13294 -1410
rect 13328 -1444 13342 -1410
rect 13272 -1479 13342 -1444
rect 13376 -1383 13428 -1327
rect 13191 -1521 13203 -1487
rect 13376 -1509 13418 -1383
rect 13556 -1409 13619 -1309
rect 13452 -1425 13619 -1409
rect 13486 -1459 13619 -1425
rect 13452 -1475 13619 -1459
rect 13237 -1521 13324 -1513
rect 13191 -1547 13324 -1521
rect 12934 -1613 12968 -1597
rect 12676 -1621 12879 -1615
rect 13002 -1615 13018 -1581
rect 13052 -1615 13073 -1581
rect 13112 -1589 13122 -1555
rect 13290 -1555 13324 -1547
rect 13112 -1605 13156 -1589
rect 13002 -1657 13073 -1615
rect 13190 -1615 13206 -1581
rect 13240 -1615 13256 -1581
rect 13290 -1605 13324 -1589
rect 13376 -1545 13428 -1509
rect 13376 -1579 13394 -1545
rect 13556 -1555 13619 -1475
rect 13190 -1657 13256 -1615
rect 13376 -1623 13428 -1579
rect 13462 -1581 13521 -1565
rect 13462 -1615 13478 -1581
rect 13512 -1615 13521 -1581
rect 13462 -1657 13521 -1615
rect 13556 -1589 13573 -1555
rect 13607 -1589 13619 -1555
rect 13556 -1623 13619 -1589
rect 13654 -1226 13711 -1181
rect 13745 -1189 14023 -1147
rect 13745 -1223 13761 -1189
rect 13795 -1223 13963 -1189
rect 13997 -1223 14023 -1189
rect 14211 -1189 14287 -1147
rect 14129 -1215 14163 -1199
rect 13654 -1260 13677 -1226
rect 14211 -1223 14237 -1189
rect 14271 -1223 14287 -1189
rect 14710 -1189 14776 -1147
rect 14129 -1257 14163 -1249
rect 14335 -1224 14451 -1190
rect 14485 -1224 14501 -1190
rect 14710 -1223 14726 -1189
rect 14760 -1223 14776 -1189
rect 14994 -1199 15070 -1147
rect 13654 -1289 13711 -1260
rect 13654 -1323 13664 -1289
rect 13698 -1294 13711 -1289
rect 13654 -1328 13677 -1323
rect 13654 -1348 13711 -1328
rect 13745 -1291 14301 -1257
rect 13654 -1531 13690 -1348
rect 13745 -1409 13779 -1291
rect 13840 -1359 13859 -1325
rect 13893 -1351 13997 -1325
rect 13893 -1359 13946 -1351
rect 13940 -1385 13946 -1359
rect 13980 -1385 13997 -1351
rect 13940 -1393 13997 -1385
rect 13726 -1425 13779 -1409
rect 13760 -1459 13779 -1425
rect 13813 -1415 13904 -1409
rect 13813 -1421 13859 -1415
rect 13813 -1455 13854 -1421
rect 13893 -1449 13904 -1415
rect 13888 -1455 13904 -1449
rect 13940 -1427 13963 -1393
rect 13940 -1452 13997 -1427
rect 13726 -1475 13779 -1459
rect 13940 -1489 13984 -1452
rect 13654 -1547 13711 -1531
rect 13654 -1581 13677 -1547
rect 13654 -1623 13711 -1581
rect 13745 -1581 13806 -1513
rect 13745 -1615 13761 -1581
rect 13795 -1615 13806 -1581
rect 13745 -1657 13806 -1615
rect 13856 -1523 13984 -1489
rect 14031 -1506 14065 -1291
rect 14251 -1309 14301 -1291
rect 14251 -1343 14267 -1309
rect 14251 -1359 14301 -1343
rect 14335 -1393 14369 -1224
rect 14710 -1257 14776 -1223
rect 14492 -1283 14539 -1277
rect 14099 -1409 14369 -1393
rect 14133 -1427 14369 -1409
rect 14133 -1443 14143 -1427
rect 14099 -1459 14143 -1443
rect 14028 -1507 14065 -1506
rect 14186 -1487 14206 -1461
rect 13856 -1571 13898 -1523
rect 14028 -1541 14044 -1507
rect 14078 -1541 14108 -1507
rect 14186 -1521 14202 -1487
rect 14240 -1495 14295 -1461
rect 14236 -1521 14295 -1495
rect 14186 -1527 14295 -1521
rect 13890 -1605 13898 -1571
rect 13856 -1621 13898 -1605
rect 13960 -1573 13994 -1557
rect 14136 -1589 14152 -1565
rect 13994 -1599 14152 -1589
rect 14186 -1599 14202 -1565
rect 13994 -1607 14202 -1599
rect 13960 -1623 14202 -1607
rect 14236 -1585 14301 -1569
rect 14270 -1619 14301 -1585
rect 14236 -1657 14301 -1619
rect 14335 -1581 14369 -1427
rect 14403 -1309 14444 -1293
rect 14437 -1343 14444 -1309
rect 14403 -1413 14444 -1343
rect 14526 -1309 14539 -1283
rect 14710 -1291 14726 -1257
rect 14760 -1291 14776 -1257
rect 14900 -1215 14934 -1199
rect 14994 -1233 15020 -1199
rect 15054 -1233 15070 -1199
rect 15118 -1224 15234 -1190
rect 15268 -1224 15284 -1190
rect 15326 -1197 15360 -1181
rect 14900 -1267 14934 -1249
rect 14814 -1283 15084 -1267
rect 14492 -1343 14505 -1317
rect 14814 -1317 14900 -1283
rect 14934 -1309 15084 -1283
rect 14934 -1317 15050 -1309
rect 14492 -1359 14539 -1343
rect 14579 -1351 14780 -1343
rect 14579 -1385 14584 -1351
rect 14618 -1385 14780 -1351
rect 14579 -1391 14780 -1385
rect 14714 -1393 14780 -1391
rect 14403 -1419 14538 -1413
rect 14403 -1449 14492 -1419
rect 14470 -1453 14492 -1449
rect 14526 -1453 14538 -1419
rect 14714 -1427 14730 -1393
rect 14764 -1427 14780 -1393
rect 14470 -1462 14538 -1453
rect 14586 -1461 14602 -1427
rect 14636 -1461 14652 -1427
rect 14814 -1461 14848 -1317
rect 15034 -1343 15050 -1317
rect 15034 -1359 15084 -1343
rect 14882 -1393 14932 -1377
rect 15118 -1393 15152 -1224
rect 15326 -1281 15360 -1231
rect 15394 -1213 15465 -1147
rect 15394 -1247 15410 -1213
rect 15444 -1247 15465 -1213
rect 15504 -1197 15548 -1181
rect 15504 -1231 15514 -1197
rect 15504 -1265 15548 -1231
rect 15582 -1213 15648 -1147
rect 15582 -1247 15598 -1213
rect 15632 -1247 15648 -1213
rect 15682 -1197 15716 -1181
rect 15186 -1309 15228 -1283
rect 15220 -1317 15228 -1309
rect 15262 -1317 15286 -1283
rect 15326 -1315 15470 -1281
rect 15220 -1343 15286 -1317
rect 15186 -1359 15286 -1343
rect 14916 -1427 15152 -1393
rect 14882 -1443 14926 -1427
rect 15068 -1435 15152 -1427
rect 14470 -1483 14514 -1462
rect 14504 -1517 14514 -1483
rect 14586 -1495 14848 -1461
rect 14968 -1481 14984 -1461
rect 14470 -1533 14514 -1517
rect 14804 -1521 14848 -1495
rect 14952 -1487 14984 -1481
rect 15018 -1495 15034 -1461
rect 14986 -1521 15034 -1495
rect 14736 -1547 14770 -1531
rect 14804 -1555 14820 -1521
rect 14854 -1555 14870 -1521
rect 14952 -1527 15034 -1521
rect 14335 -1615 14428 -1581
rect 14462 -1615 14491 -1581
rect 14335 -1621 14491 -1615
rect 14616 -1615 14632 -1581
rect 14666 -1615 14686 -1581
rect 14616 -1657 14686 -1615
rect 14736 -1589 14770 -1581
rect 14900 -1579 14966 -1573
rect 14900 -1589 14916 -1579
rect 14736 -1613 14916 -1589
rect 14950 -1613 14966 -1579
rect 14736 -1623 14966 -1613
rect 15000 -1585 15034 -1569
rect 15000 -1657 15034 -1619
rect 15068 -1581 15102 -1435
rect 15136 -1487 15156 -1471
rect 15190 -1505 15206 -1471
rect 15170 -1521 15206 -1505
rect 15136 -1545 15206 -1521
rect 15242 -1483 15286 -1359
rect 15320 -1415 15402 -1349
rect 15320 -1449 15326 -1415
rect 15360 -1423 15402 -1415
rect 15360 -1449 15368 -1423
rect 15320 -1457 15368 -1449
rect 15320 -1473 15402 -1457
rect 15242 -1517 15252 -1483
rect 15436 -1509 15470 -1315
rect 15242 -1533 15286 -1517
rect 15326 -1547 15470 -1509
rect 15504 -1283 15514 -1265
rect 15682 -1265 15716 -1231
rect 15538 -1317 15548 -1299
rect 15326 -1563 15360 -1547
rect 15068 -1615 15221 -1581
rect 15255 -1615 15271 -1581
rect 15504 -1555 15548 -1317
rect 15583 -1299 15682 -1281
rect 15583 -1315 15716 -1299
rect 15768 -1223 15820 -1181
rect 15768 -1257 15777 -1223
rect 15811 -1225 15820 -1223
rect 15768 -1259 15786 -1257
rect 15768 -1293 15820 -1259
rect 15583 -1410 15629 -1315
rect 15768 -1327 15786 -1293
rect 15854 -1201 15912 -1147
rect 15854 -1235 15870 -1201
rect 15904 -1235 15912 -1201
rect 15854 -1269 15912 -1235
rect 15854 -1303 15870 -1269
rect 15904 -1303 15912 -1269
rect 15854 -1321 15912 -1303
rect 15948 -1207 16011 -1191
rect 15948 -1241 15965 -1207
rect 15999 -1241 16011 -1207
rect 15948 -1275 16011 -1241
rect 15948 -1309 15965 -1275
rect 15999 -1309 16011 -1275
rect 15583 -1444 15584 -1410
rect 15618 -1444 15629 -1410
rect 15583 -1487 15629 -1444
rect 15664 -1358 15734 -1349
rect 15664 -1392 15673 -1358
rect 15707 -1392 15734 -1358
rect 15664 -1410 15734 -1392
rect 15664 -1444 15686 -1410
rect 15720 -1444 15734 -1410
rect 15664 -1479 15734 -1444
rect 15768 -1383 15820 -1327
rect 15583 -1521 15595 -1487
rect 15768 -1509 15810 -1383
rect 15948 -1409 16011 -1309
rect 15844 -1425 16011 -1409
rect 15878 -1459 16011 -1425
rect 15844 -1475 16011 -1459
rect 15629 -1521 15716 -1513
rect 15583 -1547 15716 -1521
rect 15326 -1613 15360 -1597
rect 15068 -1621 15271 -1615
rect 15394 -1615 15410 -1581
rect 15444 -1615 15465 -1581
rect 15504 -1589 15514 -1555
rect 15682 -1555 15716 -1547
rect 15504 -1605 15548 -1589
rect 15394 -1657 15465 -1615
rect 15582 -1615 15598 -1581
rect 15632 -1615 15648 -1581
rect 15682 -1605 15716 -1589
rect 15768 -1545 15820 -1509
rect 15768 -1579 15786 -1545
rect 15948 -1555 16011 -1475
rect 15582 -1657 15648 -1615
rect 15768 -1623 15820 -1579
rect 15854 -1581 15913 -1565
rect 15854 -1615 15870 -1581
rect 15904 -1615 15913 -1581
rect 15854 -1657 15913 -1615
rect 15948 -1589 15965 -1555
rect 15999 -1589 16011 -1555
rect 15948 -1623 16011 -1589
rect 16046 -1226 16103 -1181
rect 16137 -1189 16415 -1147
rect 16137 -1223 16153 -1189
rect 16187 -1223 16355 -1189
rect 16389 -1223 16415 -1189
rect 16603 -1189 16679 -1147
rect 16521 -1215 16555 -1199
rect 16046 -1260 16069 -1226
rect 16603 -1223 16629 -1189
rect 16663 -1223 16679 -1189
rect 17102 -1189 17168 -1147
rect 16521 -1257 16555 -1249
rect 16727 -1224 16843 -1190
rect 16877 -1224 16893 -1190
rect 17102 -1223 17118 -1189
rect 17152 -1223 17168 -1189
rect 17386 -1199 17462 -1147
rect 16046 -1289 16103 -1260
rect 16046 -1323 16057 -1289
rect 16091 -1294 16103 -1289
rect 16046 -1328 16069 -1323
rect 16046 -1348 16103 -1328
rect 16137 -1291 16693 -1257
rect 16046 -1531 16082 -1348
rect 16137 -1409 16171 -1291
rect 16232 -1359 16251 -1325
rect 16285 -1351 16389 -1325
rect 16285 -1359 16338 -1351
rect 16332 -1385 16338 -1359
rect 16372 -1385 16389 -1351
rect 16332 -1393 16389 -1385
rect 16118 -1425 16171 -1409
rect 16152 -1459 16171 -1425
rect 16205 -1415 16296 -1409
rect 16205 -1421 16252 -1415
rect 16205 -1455 16246 -1421
rect 16286 -1449 16296 -1415
rect 16280 -1455 16296 -1449
rect 16332 -1427 16355 -1393
rect 16332 -1452 16389 -1427
rect 16118 -1475 16171 -1459
rect 16332 -1489 16376 -1452
rect 16046 -1547 16103 -1531
rect 16046 -1581 16069 -1547
rect 16046 -1623 16103 -1581
rect 16137 -1581 16198 -1513
rect 16137 -1615 16153 -1581
rect 16187 -1615 16198 -1581
rect 16137 -1657 16198 -1615
rect 16248 -1523 16376 -1489
rect 16423 -1506 16457 -1291
rect 16643 -1309 16693 -1291
rect 16643 -1343 16659 -1309
rect 16643 -1359 16693 -1343
rect 16727 -1393 16761 -1224
rect 17102 -1257 17168 -1223
rect 16884 -1283 16931 -1277
rect 16491 -1409 16761 -1393
rect 16525 -1427 16761 -1409
rect 16525 -1443 16535 -1427
rect 16491 -1459 16535 -1443
rect 16420 -1507 16457 -1506
rect 16578 -1487 16598 -1461
rect 16248 -1571 16290 -1523
rect 16420 -1541 16436 -1507
rect 16470 -1541 16500 -1507
rect 16578 -1521 16594 -1487
rect 16632 -1495 16687 -1461
rect 16628 -1521 16687 -1495
rect 16578 -1527 16687 -1521
rect 16282 -1605 16290 -1571
rect 16248 -1621 16290 -1605
rect 16352 -1573 16386 -1557
rect 16528 -1589 16544 -1565
rect 16386 -1599 16544 -1589
rect 16578 -1599 16594 -1565
rect 16386 -1607 16594 -1599
rect 16352 -1623 16594 -1607
rect 16628 -1585 16693 -1569
rect 16662 -1619 16693 -1585
rect 16628 -1657 16693 -1619
rect 16727 -1581 16761 -1427
rect 16795 -1309 16836 -1293
rect 16829 -1343 16836 -1309
rect 16795 -1413 16836 -1343
rect 16918 -1309 16931 -1283
rect 17102 -1291 17118 -1257
rect 17152 -1291 17168 -1257
rect 17292 -1215 17326 -1199
rect 17386 -1233 17412 -1199
rect 17446 -1233 17462 -1199
rect 17510 -1224 17626 -1190
rect 17660 -1224 17676 -1190
rect 17718 -1197 17752 -1181
rect 17292 -1267 17326 -1249
rect 17206 -1283 17476 -1267
rect 16884 -1343 16897 -1317
rect 17206 -1317 17292 -1283
rect 17326 -1309 17476 -1283
rect 17326 -1317 17442 -1309
rect 16884 -1359 16931 -1343
rect 16971 -1351 17172 -1343
rect 16971 -1385 16976 -1351
rect 17010 -1385 17172 -1351
rect 16971 -1391 17172 -1385
rect 17106 -1393 17172 -1391
rect 16795 -1419 16930 -1413
rect 16795 -1449 16884 -1419
rect 16862 -1453 16884 -1449
rect 16918 -1453 16930 -1419
rect 17106 -1427 17122 -1393
rect 17156 -1427 17172 -1393
rect 16862 -1462 16930 -1453
rect 16978 -1461 16994 -1427
rect 17028 -1461 17044 -1427
rect 17206 -1461 17240 -1317
rect 17426 -1343 17442 -1317
rect 17426 -1359 17476 -1343
rect 17274 -1393 17324 -1377
rect 17510 -1393 17544 -1224
rect 17718 -1281 17752 -1231
rect 17786 -1213 17857 -1147
rect 17786 -1247 17802 -1213
rect 17836 -1247 17857 -1213
rect 17896 -1197 17940 -1181
rect 17896 -1231 17906 -1197
rect 17896 -1265 17940 -1231
rect 17974 -1213 18040 -1147
rect 17974 -1247 17990 -1213
rect 18024 -1247 18040 -1213
rect 18074 -1197 18108 -1181
rect 17578 -1309 17620 -1283
rect 17612 -1317 17620 -1309
rect 17654 -1317 17678 -1283
rect 17718 -1315 17862 -1281
rect 17612 -1343 17678 -1317
rect 17578 -1359 17678 -1343
rect 17308 -1427 17544 -1393
rect 17274 -1443 17318 -1427
rect 17460 -1435 17544 -1427
rect 16862 -1483 16906 -1462
rect 16896 -1517 16906 -1483
rect 16978 -1495 17240 -1461
rect 17360 -1481 17376 -1461
rect 16862 -1533 16906 -1517
rect 17196 -1521 17240 -1495
rect 17344 -1487 17376 -1481
rect 17410 -1495 17426 -1461
rect 17378 -1521 17426 -1495
rect 17128 -1547 17162 -1531
rect 17196 -1555 17212 -1521
rect 17246 -1555 17262 -1521
rect 17344 -1527 17426 -1521
rect 16727 -1615 16820 -1581
rect 16854 -1615 16883 -1581
rect 16727 -1621 16883 -1615
rect 17008 -1615 17024 -1581
rect 17058 -1615 17078 -1581
rect 17008 -1657 17078 -1615
rect 17128 -1589 17162 -1581
rect 17292 -1579 17358 -1573
rect 17292 -1589 17308 -1579
rect 17128 -1613 17308 -1589
rect 17342 -1613 17358 -1579
rect 17128 -1623 17358 -1613
rect 17392 -1585 17426 -1569
rect 17392 -1657 17426 -1619
rect 17460 -1581 17494 -1435
rect 17528 -1487 17548 -1471
rect 17582 -1505 17598 -1471
rect 17562 -1521 17598 -1505
rect 17528 -1545 17598 -1521
rect 17634 -1483 17678 -1359
rect 17712 -1416 17794 -1349
rect 17712 -1450 17719 -1416
rect 17753 -1423 17794 -1416
rect 17753 -1450 17760 -1423
rect 17712 -1457 17760 -1450
rect 17712 -1473 17794 -1457
rect 17634 -1517 17644 -1483
rect 17828 -1509 17862 -1315
rect 17634 -1533 17678 -1517
rect 17718 -1547 17862 -1509
rect 17896 -1283 17906 -1265
rect 18074 -1265 18108 -1231
rect 17930 -1317 17940 -1299
rect 17718 -1563 17752 -1547
rect 17460 -1615 17613 -1581
rect 17647 -1615 17663 -1581
rect 17896 -1555 17940 -1317
rect 17975 -1299 18074 -1281
rect 17975 -1315 18108 -1299
rect 18160 -1224 18212 -1181
rect 18160 -1258 18169 -1224
rect 18203 -1225 18212 -1224
rect 18160 -1259 18178 -1258
rect 18160 -1293 18212 -1259
rect 17975 -1410 18021 -1315
rect 18160 -1327 18178 -1293
rect 18246 -1201 18304 -1147
rect 18246 -1235 18262 -1201
rect 18296 -1235 18304 -1201
rect 18246 -1269 18304 -1235
rect 18246 -1303 18262 -1269
rect 18296 -1303 18304 -1269
rect 18246 -1321 18304 -1303
rect 18340 -1207 18403 -1191
rect 18340 -1241 18357 -1207
rect 18391 -1241 18403 -1207
rect 18340 -1275 18403 -1241
rect 18340 -1309 18357 -1275
rect 18391 -1309 18403 -1275
rect 17975 -1444 17976 -1410
rect 18010 -1444 18021 -1410
rect 17975 -1487 18021 -1444
rect 18056 -1360 18126 -1349
rect 18056 -1394 18065 -1360
rect 18099 -1394 18126 -1360
rect 18056 -1410 18126 -1394
rect 18056 -1444 18078 -1410
rect 18112 -1444 18126 -1410
rect 18056 -1479 18126 -1444
rect 18160 -1383 18212 -1327
rect 17975 -1521 17987 -1487
rect 18160 -1509 18202 -1383
rect 18340 -1409 18403 -1309
rect 18236 -1425 18403 -1409
rect 18270 -1459 18403 -1425
rect 18236 -1475 18403 -1459
rect 18021 -1521 18108 -1513
rect 17975 -1547 18108 -1521
rect 17718 -1613 17752 -1597
rect 17460 -1621 17663 -1615
rect 17786 -1615 17802 -1581
rect 17836 -1615 17857 -1581
rect 17896 -1589 17906 -1555
rect 18074 -1555 18108 -1547
rect 17896 -1605 17940 -1589
rect 17786 -1657 17857 -1615
rect 17974 -1615 17990 -1581
rect 18024 -1615 18040 -1581
rect 18074 -1605 18108 -1589
rect 18160 -1545 18212 -1509
rect 18160 -1579 18178 -1545
rect 18340 -1555 18403 -1475
rect 17974 -1657 18040 -1615
rect 18160 -1623 18212 -1579
rect 18246 -1581 18305 -1565
rect 18246 -1615 18262 -1581
rect 18296 -1615 18305 -1581
rect 18246 -1657 18305 -1615
rect 18340 -1589 18357 -1555
rect 18391 -1589 18403 -1555
rect 18340 -1623 18403 -1589
rect 18438 -1226 18495 -1181
rect 18529 -1189 18807 -1147
rect 18529 -1223 18545 -1189
rect 18579 -1223 18747 -1189
rect 18781 -1223 18807 -1189
rect 18995 -1189 19071 -1147
rect 18913 -1215 18947 -1199
rect 18438 -1260 18461 -1226
rect 18995 -1223 19021 -1189
rect 19055 -1223 19071 -1189
rect 19494 -1189 19560 -1147
rect 18913 -1257 18947 -1249
rect 19119 -1224 19235 -1190
rect 19269 -1224 19285 -1190
rect 19494 -1223 19510 -1189
rect 19544 -1223 19560 -1189
rect 19778 -1199 19854 -1147
rect 18438 -1289 18495 -1260
rect 18438 -1323 18449 -1289
rect 18483 -1294 18495 -1289
rect 18438 -1328 18461 -1323
rect 18438 -1348 18495 -1328
rect 18529 -1291 19085 -1257
rect 18438 -1531 18474 -1348
rect 18529 -1409 18563 -1291
rect 18624 -1359 18643 -1325
rect 18677 -1351 18781 -1325
rect 18677 -1359 18730 -1351
rect 18724 -1385 18730 -1359
rect 18764 -1385 18781 -1351
rect 18724 -1393 18781 -1385
rect 18510 -1425 18563 -1409
rect 18544 -1459 18563 -1425
rect 18597 -1415 18688 -1409
rect 18597 -1421 18643 -1415
rect 18597 -1455 18638 -1421
rect 18677 -1449 18688 -1415
rect 18672 -1455 18688 -1449
rect 18724 -1427 18747 -1393
rect 18724 -1452 18781 -1427
rect 18510 -1475 18563 -1459
rect 18724 -1489 18768 -1452
rect 18438 -1547 18495 -1531
rect 18438 -1581 18461 -1547
rect 18438 -1623 18495 -1581
rect 18529 -1581 18590 -1513
rect 18529 -1615 18545 -1581
rect 18579 -1615 18590 -1581
rect 18529 -1657 18590 -1615
rect 18640 -1523 18768 -1489
rect 18815 -1506 18849 -1291
rect 19035 -1309 19085 -1291
rect 19035 -1343 19051 -1309
rect 19035 -1359 19085 -1343
rect 19119 -1393 19153 -1224
rect 19494 -1257 19560 -1223
rect 19276 -1283 19323 -1277
rect 18883 -1409 19153 -1393
rect 18917 -1427 19153 -1409
rect 18917 -1443 18927 -1427
rect 18883 -1459 18927 -1443
rect 18812 -1507 18849 -1506
rect 18970 -1487 18990 -1461
rect 18640 -1571 18682 -1523
rect 18812 -1541 18828 -1507
rect 18862 -1541 18892 -1507
rect 18970 -1521 18986 -1487
rect 19024 -1495 19079 -1461
rect 19020 -1521 19079 -1495
rect 18970 -1527 19079 -1521
rect 18674 -1605 18682 -1571
rect 18640 -1621 18682 -1605
rect 18744 -1573 18778 -1557
rect 18920 -1589 18936 -1565
rect 18778 -1599 18936 -1589
rect 18970 -1599 18986 -1565
rect 18778 -1607 18986 -1599
rect 18744 -1623 18986 -1607
rect 19020 -1585 19085 -1569
rect 19054 -1619 19085 -1585
rect 19020 -1657 19085 -1619
rect 19119 -1581 19153 -1427
rect 19187 -1309 19228 -1293
rect 19221 -1343 19228 -1309
rect 19187 -1413 19228 -1343
rect 19310 -1309 19323 -1283
rect 19494 -1291 19510 -1257
rect 19544 -1291 19560 -1257
rect 19684 -1215 19718 -1199
rect 19778 -1233 19804 -1199
rect 19838 -1233 19854 -1199
rect 19902 -1224 20018 -1190
rect 20052 -1224 20068 -1190
rect 20110 -1197 20144 -1181
rect 19684 -1267 19718 -1249
rect 19598 -1283 19868 -1267
rect 19276 -1343 19289 -1317
rect 19598 -1317 19684 -1283
rect 19718 -1309 19868 -1283
rect 19718 -1317 19834 -1309
rect 19276 -1359 19323 -1343
rect 19363 -1351 19564 -1343
rect 19363 -1385 19368 -1351
rect 19402 -1385 19564 -1351
rect 19363 -1391 19564 -1385
rect 19498 -1393 19564 -1391
rect 19187 -1419 19322 -1413
rect 19187 -1449 19276 -1419
rect 19254 -1453 19276 -1449
rect 19310 -1453 19322 -1419
rect 19498 -1427 19514 -1393
rect 19548 -1427 19564 -1393
rect 19254 -1462 19322 -1453
rect 19370 -1461 19386 -1427
rect 19420 -1461 19436 -1427
rect 19598 -1461 19632 -1317
rect 19818 -1343 19834 -1317
rect 19818 -1359 19868 -1343
rect 19666 -1393 19716 -1377
rect 19902 -1393 19936 -1224
rect 20110 -1281 20144 -1231
rect 20178 -1213 20249 -1147
rect 20178 -1247 20194 -1213
rect 20228 -1247 20249 -1213
rect 20288 -1197 20332 -1181
rect 20288 -1231 20298 -1197
rect 20288 -1265 20332 -1231
rect 20366 -1213 20432 -1147
rect 20366 -1247 20382 -1213
rect 20416 -1247 20432 -1213
rect 20466 -1197 20500 -1181
rect 19970 -1309 20012 -1283
rect 20004 -1317 20012 -1309
rect 20046 -1317 20070 -1283
rect 20110 -1315 20254 -1281
rect 20004 -1343 20070 -1317
rect 19970 -1359 20070 -1343
rect 19700 -1427 19936 -1393
rect 19666 -1443 19710 -1427
rect 19852 -1435 19936 -1427
rect 19254 -1483 19298 -1462
rect 19288 -1517 19298 -1483
rect 19370 -1495 19632 -1461
rect 19752 -1481 19768 -1461
rect 19254 -1533 19298 -1517
rect 19588 -1521 19632 -1495
rect 19736 -1487 19768 -1481
rect 19802 -1495 19818 -1461
rect 19770 -1521 19818 -1495
rect 19520 -1547 19554 -1531
rect 19588 -1555 19604 -1521
rect 19638 -1555 19654 -1521
rect 19736 -1527 19818 -1521
rect 19119 -1615 19212 -1581
rect 19246 -1615 19275 -1581
rect 19119 -1621 19275 -1615
rect 19400 -1615 19416 -1581
rect 19450 -1615 19470 -1581
rect 19400 -1657 19470 -1615
rect 19520 -1589 19554 -1581
rect 19684 -1579 19750 -1573
rect 19684 -1589 19700 -1579
rect 19520 -1613 19700 -1589
rect 19734 -1613 19750 -1579
rect 19520 -1623 19750 -1613
rect 19784 -1585 19818 -1569
rect 19784 -1657 19818 -1619
rect 19852 -1581 19886 -1435
rect 19920 -1487 19940 -1471
rect 19974 -1505 19990 -1471
rect 19954 -1521 19990 -1505
rect 19920 -1545 19990 -1521
rect 20026 -1483 20070 -1359
rect 20104 -1416 20186 -1349
rect 20104 -1450 20110 -1416
rect 20144 -1423 20186 -1416
rect 20144 -1450 20152 -1423
rect 20104 -1457 20152 -1450
rect 20104 -1473 20186 -1457
rect 20026 -1517 20036 -1483
rect 20220 -1509 20254 -1315
rect 20026 -1533 20070 -1517
rect 20110 -1547 20254 -1509
rect 20288 -1283 20298 -1265
rect 20466 -1265 20500 -1231
rect 20322 -1317 20332 -1299
rect 20110 -1563 20144 -1547
rect 19852 -1615 20005 -1581
rect 20039 -1615 20055 -1581
rect 20288 -1555 20332 -1317
rect 20367 -1299 20466 -1281
rect 20367 -1315 20500 -1299
rect 20552 -1222 20604 -1181
rect 20552 -1256 20562 -1222
rect 20596 -1225 20604 -1222
rect 20552 -1259 20570 -1256
rect 20552 -1293 20604 -1259
rect 20367 -1410 20413 -1315
rect 20552 -1327 20570 -1293
rect 20638 -1201 20696 -1147
rect 20638 -1235 20654 -1201
rect 20688 -1235 20696 -1201
rect 20638 -1269 20696 -1235
rect 20638 -1303 20654 -1269
rect 20688 -1303 20696 -1269
rect 20638 -1321 20696 -1303
rect 20732 -1207 20795 -1191
rect 20732 -1241 20749 -1207
rect 20783 -1241 20795 -1207
rect 20732 -1275 20795 -1241
rect 20732 -1309 20749 -1275
rect 20783 -1309 20795 -1275
rect 20367 -1444 20368 -1410
rect 20402 -1444 20413 -1410
rect 20367 -1487 20413 -1444
rect 20448 -1358 20518 -1349
rect 20448 -1392 20457 -1358
rect 20491 -1392 20518 -1358
rect 20448 -1410 20518 -1392
rect 20448 -1444 20470 -1410
rect 20504 -1444 20518 -1410
rect 20448 -1479 20518 -1444
rect 20552 -1383 20604 -1327
rect 20367 -1521 20379 -1487
rect 20552 -1509 20594 -1383
rect 20732 -1409 20795 -1309
rect 20628 -1425 20795 -1409
rect 20662 -1459 20795 -1425
rect 20628 -1475 20795 -1459
rect 20413 -1521 20500 -1513
rect 20367 -1547 20500 -1521
rect 20110 -1613 20144 -1597
rect 19852 -1621 20055 -1615
rect 20178 -1615 20194 -1581
rect 20228 -1615 20249 -1581
rect 20288 -1589 20298 -1555
rect 20466 -1555 20500 -1547
rect 20288 -1605 20332 -1589
rect 20178 -1657 20249 -1615
rect 20366 -1615 20382 -1581
rect 20416 -1615 20432 -1581
rect 20466 -1605 20500 -1589
rect 20552 -1545 20604 -1509
rect 20552 -1579 20570 -1545
rect 20732 -1555 20795 -1475
rect 20366 -1657 20432 -1615
rect 20552 -1623 20604 -1579
rect 20638 -1581 20697 -1565
rect 20638 -1615 20654 -1581
rect 20688 -1615 20697 -1581
rect 20638 -1657 20697 -1615
rect 20732 -1589 20749 -1555
rect 20783 -1589 20795 -1555
rect 20732 -1623 20795 -1589
rect 20830 -1226 20887 -1181
rect 20921 -1189 21199 -1147
rect 20921 -1223 20937 -1189
rect 20971 -1223 21139 -1189
rect 21173 -1223 21199 -1189
rect 21387 -1189 21463 -1147
rect 21305 -1215 21339 -1199
rect 20830 -1260 20853 -1226
rect 21387 -1223 21413 -1189
rect 21447 -1223 21463 -1189
rect 21886 -1189 21952 -1147
rect 21305 -1257 21339 -1249
rect 21511 -1224 21627 -1190
rect 21661 -1224 21677 -1190
rect 21886 -1223 21902 -1189
rect 21936 -1223 21952 -1189
rect 22170 -1199 22246 -1147
rect 20830 -1288 20887 -1260
rect 20830 -1322 20840 -1288
rect 20874 -1294 20887 -1288
rect 20830 -1328 20853 -1322
rect 20830 -1348 20887 -1328
rect 20921 -1291 21477 -1257
rect 20830 -1531 20866 -1348
rect 20921 -1409 20955 -1291
rect 21016 -1359 21035 -1325
rect 21069 -1351 21173 -1325
rect 21069 -1359 21122 -1351
rect 21116 -1385 21122 -1359
rect 21156 -1385 21173 -1351
rect 21116 -1393 21173 -1385
rect 20902 -1425 20955 -1409
rect 20936 -1459 20955 -1425
rect 20989 -1415 21080 -1409
rect 20989 -1421 21036 -1415
rect 20989 -1455 21030 -1421
rect 21070 -1449 21080 -1415
rect 21064 -1455 21080 -1449
rect 21116 -1427 21139 -1393
rect 21116 -1452 21173 -1427
rect 20902 -1475 20955 -1459
rect 21116 -1489 21160 -1452
rect 20830 -1547 20887 -1531
rect 20830 -1581 20853 -1547
rect 20830 -1623 20887 -1581
rect 20921 -1581 20982 -1513
rect 20921 -1615 20937 -1581
rect 20971 -1615 20982 -1581
rect 20921 -1657 20982 -1615
rect 21032 -1523 21160 -1489
rect 21207 -1506 21241 -1291
rect 21427 -1309 21477 -1291
rect 21427 -1343 21443 -1309
rect 21427 -1359 21477 -1343
rect 21511 -1393 21545 -1224
rect 21886 -1257 21952 -1223
rect 21668 -1283 21715 -1277
rect 21275 -1409 21545 -1393
rect 21309 -1427 21545 -1409
rect 21309 -1443 21319 -1427
rect 21275 -1459 21319 -1443
rect 21204 -1507 21241 -1506
rect 21362 -1487 21382 -1461
rect 21032 -1571 21074 -1523
rect 21204 -1541 21220 -1507
rect 21254 -1541 21284 -1507
rect 21362 -1521 21378 -1487
rect 21416 -1495 21471 -1461
rect 21412 -1521 21471 -1495
rect 21362 -1527 21471 -1521
rect 21066 -1605 21074 -1571
rect 21032 -1621 21074 -1605
rect 21136 -1573 21170 -1557
rect 21312 -1589 21328 -1565
rect 21170 -1599 21328 -1589
rect 21362 -1599 21378 -1565
rect 21170 -1607 21378 -1599
rect 21136 -1623 21378 -1607
rect 21412 -1585 21477 -1569
rect 21446 -1619 21477 -1585
rect 21412 -1657 21477 -1619
rect 21511 -1581 21545 -1427
rect 21579 -1309 21620 -1293
rect 21613 -1343 21620 -1309
rect 21579 -1413 21620 -1343
rect 21702 -1309 21715 -1283
rect 21886 -1291 21902 -1257
rect 21936 -1291 21952 -1257
rect 22076 -1215 22110 -1199
rect 22170 -1233 22196 -1199
rect 22230 -1233 22246 -1199
rect 22294 -1224 22410 -1190
rect 22444 -1224 22460 -1190
rect 22502 -1197 22536 -1181
rect 22076 -1267 22110 -1249
rect 21990 -1283 22260 -1267
rect 21668 -1343 21681 -1317
rect 21990 -1317 22076 -1283
rect 22110 -1309 22260 -1283
rect 22110 -1317 22226 -1309
rect 21668 -1359 21715 -1343
rect 21755 -1351 21956 -1343
rect 21755 -1385 21760 -1351
rect 21794 -1385 21956 -1351
rect 21755 -1391 21956 -1385
rect 21890 -1393 21956 -1391
rect 21579 -1419 21714 -1413
rect 21579 -1449 21668 -1419
rect 21646 -1453 21668 -1449
rect 21702 -1453 21714 -1419
rect 21890 -1427 21906 -1393
rect 21940 -1427 21956 -1393
rect 21646 -1462 21714 -1453
rect 21762 -1461 21778 -1427
rect 21812 -1461 21828 -1427
rect 21990 -1461 22024 -1317
rect 22210 -1343 22226 -1317
rect 22210 -1359 22260 -1343
rect 22058 -1393 22108 -1377
rect 22294 -1393 22328 -1224
rect 22502 -1281 22536 -1231
rect 22570 -1213 22641 -1147
rect 22570 -1247 22586 -1213
rect 22620 -1247 22641 -1213
rect 22680 -1197 22724 -1181
rect 22680 -1231 22690 -1197
rect 22680 -1265 22724 -1231
rect 22758 -1213 22824 -1147
rect 22758 -1247 22774 -1213
rect 22808 -1247 22824 -1213
rect 22858 -1197 22892 -1181
rect 22362 -1309 22404 -1283
rect 22396 -1317 22404 -1309
rect 22438 -1317 22462 -1283
rect 22502 -1315 22646 -1281
rect 22396 -1343 22462 -1317
rect 22362 -1359 22462 -1343
rect 22092 -1427 22328 -1393
rect 22058 -1443 22102 -1427
rect 22244 -1435 22328 -1427
rect 21646 -1483 21690 -1462
rect 21680 -1517 21690 -1483
rect 21762 -1495 22024 -1461
rect 22144 -1481 22160 -1461
rect 21646 -1533 21690 -1517
rect 21980 -1521 22024 -1495
rect 22128 -1487 22160 -1481
rect 22194 -1495 22210 -1461
rect 22162 -1521 22210 -1495
rect 21912 -1547 21946 -1531
rect 21980 -1555 21996 -1521
rect 22030 -1555 22046 -1521
rect 22128 -1527 22210 -1521
rect 21511 -1615 21604 -1581
rect 21638 -1615 21667 -1581
rect 21511 -1621 21667 -1615
rect 21792 -1615 21808 -1581
rect 21842 -1615 21862 -1581
rect 21792 -1657 21862 -1615
rect 21912 -1589 21946 -1581
rect 22076 -1579 22142 -1573
rect 22076 -1589 22092 -1579
rect 21912 -1613 22092 -1589
rect 22126 -1613 22142 -1579
rect 21912 -1623 22142 -1613
rect 22176 -1585 22210 -1569
rect 22176 -1657 22210 -1619
rect 22244 -1581 22278 -1435
rect 22312 -1487 22332 -1471
rect 22366 -1505 22382 -1471
rect 22346 -1521 22382 -1505
rect 22312 -1545 22382 -1521
rect 22418 -1483 22462 -1359
rect 22496 -1416 22578 -1349
rect 22496 -1450 22503 -1416
rect 22537 -1423 22578 -1416
rect 22537 -1450 22544 -1423
rect 22496 -1457 22544 -1450
rect 22496 -1473 22578 -1457
rect 22418 -1517 22428 -1483
rect 22612 -1509 22646 -1315
rect 22418 -1533 22462 -1517
rect 22502 -1547 22646 -1509
rect 22680 -1283 22690 -1265
rect 22858 -1265 22892 -1231
rect 22714 -1317 22724 -1299
rect 22502 -1563 22536 -1547
rect 22244 -1615 22397 -1581
rect 22431 -1615 22447 -1581
rect 22680 -1555 22724 -1317
rect 22759 -1299 22858 -1281
rect 22759 -1315 22892 -1299
rect 22944 -1222 22996 -1181
rect 22944 -1256 22953 -1222
rect 22987 -1225 22996 -1222
rect 22944 -1259 22962 -1256
rect 22944 -1293 22996 -1259
rect 22759 -1410 22805 -1315
rect 22944 -1327 22962 -1293
rect 23030 -1201 23088 -1147
rect 23030 -1235 23046 -1201
rect 23080 -1235 23088 -1201
rect 23030 -1269 23088 -1235
rect 23030 -1303 23046 -1269
rect 23080 -1303 23088 -1269
rect 23030 -1321 23088 -1303
rect 23124 -1207 23187 -1191
rect 23124 -1241 23141 -1207
rect 23175 -1241 23187 -1207
rect 23124 -1275 23187 -1241
rect 23124 -1309 23141 -1275
rect 23175 -1309 23187 -1275
rect 22759 -1444 22760 -1410
rect 22794 -1444 22805 -1410
rect 22759 -1487 22805 -1444
rect 22840 -1360 22910 -1349
rect 22840 -1394 22849 -1360
rect 22883 -1394 22910 -1360
rect 22840 -1410 22910 -1394
rect 22840 -1444 22862 -1410
rect 22896 -1444 22910 -1410
rect 22840 -1479 22910 -1444
rect 22944 -1383 22996 -1327
rect 22759 -1521 22771 -1487
rect 22944 -1509 22986 -1383
rect 23124 -1409 23187 -1309
rect 23020 -1425 23187 -1409
rect 23054 -1459 23187 -1425
rect 23020 -1475 23187 -1459
rect 22805 -1521 22892 -1513
rect 22759 -1547 22892 -1521
rect 22502 -1613 22536 -1597
rect 22244 -1621 22447 -1615
rect 22570 -1615 22586 -1581
rect 22620 -1615 22641 -1581
rect 22680 -1589 22690 -1555
rect 22858 -1555 22892 -1547
rect 22680 -1605 22724 -1589
rect 22570 -1657 22641 -1615
rect 22758 -1615 22774 -1581
rect 22808 -1615 22824 -1581
rect 22858 -1605 22892 -1589
rect 22944 -1545 22996 -1509
rect 22944 -1579 22962 -1545
rect 23124 -1555 23187 -1475
rect 22758 -1657 22824 -1615
rect 22944 -1623 22996 -1579
rect 23030 -1581 23089 -1565
rect 23030 -1615 23046 -1581
rect 23080 -1615 23089 -1581
rect 23030 -1657 23089 -1615
rect 23124 -1589 23141 -1555
rect 23175 -1589 23187 -1555
rect 23124 -1623 23187 -1589
rect 23222 -1226 23279 -1181
rect 23313 -1189 23591 -1147
rect 23313 -1223 23329 -1189
rect 23363 -1223 23531 -1189
rect 23565 -1223 23591 -1189
rect 23779 -1189 23855 -1147
rect 23697 -1215 23731 -1199
rect 23222 -1260 23245 -1226
rect 23779 -1223 23805 -1189
rect 23839 -1223 23855 -1189
rect 24278 -1189 24344 -1147
rect 23697 -1257 23731 -1249
rect 23903 -1224 24019 -1190
rect 24053 -1224 24069 -1190
rect 24278 -1223 24294 -1189
rect 24328 -1223 24344 -1189
rect 24562 -1199 24638 -1147
rect 23222 -1289 23279 -1260
rect 23222 -1323 23233 -1289
rect 23267 -1294 23279 -1289
rect 23222 -1328 23245 -1323
rect 23222 -1348 23279 -1328
rect 23313 -1291 23869 -1257
rect 23222 -1531 23258 -1348
rect 23313 -1409 23347 -1291
rect 23408 -1359 23427 -1325
rect 23461 -1351 23565 -1325
rect 23461 -1359 23514 -1351
rect 23508 -1385 23514 -1359
rect 23548 -1385 23565 -1351
rect 23508 -1393 23565 -1385
rect 23294 -1425 23347 -1409
rect 23328 -1459 23347 -1425
rect 23381 -1415 23472 -1409
rect 23381 -1421 23427 -1415
rect 23381 -1455 23422 -1421
rect 23461 -1449 23472 -1415
rect 23456 -1455 23472 -1449
rect 23508 -1427 23531 -1393
rect 23508 -1452 23565 -1427
rect 23294 -1475 23347 -1459
rect 23508 -1489 23552 -1452
rect 23222 -1547 23279 -1531
rect 23222 -1581 23245 -1547
rect 23222 -1623 23279 -1581
rect 23313 -1581 23374 -1513
rect 23313 -1615 23329 -1581
rect 23363 -1615 23374 -1581
rect 23313 -1657 23374 -1615
rect 23424 -1523 23552 -1489
rect 23599 -1506 23633 -1291
rect 23819 -1309 23869 -1291
rect 23819 -1343 23835 -1309
rect 23819 -1359 23869 -1343
rect 23903 -1393 23937 -1224
rect 24278 -1257 24344 -1223
rect 24060 -1283 24107 -1277
rect 23667 -1409 23937 -1393
rect 23701 -1427 23937 -1409
rect 23701 -1443 23711 -1427
rect 23667 -1459 23711 -1443
rect 23596 -1507 23633 -1506
rect 23754 -1487 23774 -1461
rect 23424 -1571 23466 -1523
rect 23596 -1541 23612 -1507
rect 23646 -1541 23676 -1507
rect 23754 -1521 23770 -1487
rect 23808 -1495 23863 -1461
rect 23804 -1521 23863 -1495
rect 23754 -1527 23863 -1521
rect 23458 -1605 23466 -1571
rect 23424 -1621 23466 -1605
rect 23528 -1573 23562 -1557
rect 23704 -1589 23720 -1565
rect 23562 -1599 23720 -1589
rect 23754 -1599 23770 -1565
rect 23562 -1607 23770 -1599
rect 23528 -1623 23770 -1607
rect 23804 -1585 23869 -1569
rect 23838 -1619 23869 -1585
rect 23804 -1657 23869 -1619
rect 23903 -1581 23937 -1427
rect 23971 -1309 24012 -1293
rect 24005 -1343 24012 -1309
rect 23971 -1413 24012 -1343
rect 24094 -1309 24107 -1283
rect 24278 -1291 24294 -1257
rect 24328 -1291 24344 -1257
rect 24468 -1215 24502 -1199
rect 24562 -1233 24588 -1199
rect 24622 -1233 24638 -1199
rect 24686 -1224 24802 -1190
rect 24836 -1224 24852 -1190
rect 24894 -1197 24928 -1181
rect 24468 -1267 24502 -1249
rect 24382 -1283 24652 -1267
rect 24060 -1343 24073 -1317
rect 24382 -1317 24468 -1283
rect 24502 -1309 24652 -1283
rect 24502 -1317 24618 -1309
rect 24060 -1359 24107 -1343
rect 24147 -1351 24348 -1343
rect 24147 -1385 24152 -1351
rect 24186 -1385 24348 -1351
rect 24147 -1391 24348 -1385
rect 24282 -1393 24348 -1391
rect 23971 -1419 24106 -1413
rect 23971 -1449 24060 -1419
rect 24038 -1453 24060 -1449
rect 24094 -1453 24106 -1419
rect 24282 -1427 24298 -1393
rect 24332 -1427 24348 -1393
rect 24038 -1462 24106 -1453
rect 24154 -1461 24170 -1427
rect 24204 -1461 24220 -1427
rect 24382 -1461 24416 -1317
rect 24602 -1343 24618 -1317
rect 24602 -1359 24652 -1343
rect 24450 -1393 24500 -1377
rect 24686 -1393 24720 -1224
rect 24894 -1281 24928 -1231
rect 24962 -1213 25033 -1147
rect 24962 -1247 24978 -1213
rect 25012 -1247 25033 -1213
rect 25072 -1197 25116 -1181
rect 25072 -1231 25082 -1197
rect 25072 -1265 25116 -1231
rect 25150 -1213 25216 -1147
rect 25150 -1247 25166 -1213
rect 25200 -1247 25216 -1213
rect 25250 -1197 25284 -1181
rect 24754 -1309 24796 -1283
rect 24788 -1317 24796 -1309
rect 24830 -1317 24854 -1283
rect 24894 -1315 25038 -1281
rect 24788 -1343 24854 -1317
rect 24754 -1359 24854 -1343
rect 24484 -1427 24720 -1393
rect 24450 -1443 24494 -1427
rect 24636 -1435 24720 -1427
rect 24038 -1483 24082 -1462
rect 24072 -1517 24082 -1483
rect 24154 -1495 24416 -1461
rect 24536 -1481 24552 -1461
rect 24038 -1533 24082 -1517
rect 24372 -1521 24416 -1495
rect 24520 -1487 24552 -1481
rect 24586 -1495 24602 -1461
rect 24554 -1521 24602 -1495
rect 24304 -1547 24338 -1531
rect 24372 -1555 24388 -1521
rect 24422 -1555 24438 -1521
rect 24520 -1527 24602 -1521
rect 23903 -1615 23996 -1581
rect 24030 -1615 24059 -1581
rect 23903 -1621 24059 -1615
rect 24184 -1615 24200 -1581
rect 24234 -1615 24254 -1581
rect 24184 -1657 24254 -1615
rect 24304 -1589 24338 -1581
rect 24468 -1579 24534 -1573
rect 24468 -1589 24484 -1579
rect 24304 -1613 24484 -1589
rect 24518 -1613 24534 -1579
rect 24304 -1623 24534 -1613
rect 24568 -1585 24602 -1569
rect 24568 -1657 24602 -1619
rect 24636 -1581 24670 -1435
rect 24704 -1487 24724 -1471
rect 24758 -1505 24774 -1471
rect 24738 -1521 24774 -1505
rect 24704 -1545 24774 -1521
rect 24810 -1483 24854 -1359
rect 24888 -1416 24970 -1349
rect 24888 -1450 24896 -1416
rect 24930 -1423 24970 -1416
rect 24930 -1450 24936 -1423
rect 24888 -1457 24936 -1450
rect 24888 -1473 24970 -1457
rect 24810 -1517 24820 -1483
rect 25004 -1509 25038 -1315
rect 24810 -1533 24854 -1517
rect 24894 -1547 25038 -1509
rect 25072 -1283 25082 -1265
rect 25250 -1265 25284 -1231
rect 25106 -1317 25116 -1299
rect 24894 -1563 24928 -1547
rect 24636 -1615 24789 -1581
rect 24823 -1615 24839 -1581
rect 25072 -1555 25116 -1317
rect 25151 -1299 25250 -1281
rect 25151 -1315 25284 -1299
rect 25151 -1410 25197 -1315
rect 25151 -1444 25152 -1410
rect 25186 -1444 25197 -1410
rect 25151 -1487 25197 -1444
rect 25232 -1358 25302 -1349
rect 25232 -1392 25241 -1358
rect 25275 -1392 25302 -1358
rect 25232 -1410 25302 -1392
rect 25232 -1444 25254 -1410
rect 25288 -1444 25302 -1410
rect 25232 -1479 25302 -1444
rect 25151 -1521 25163 -1487
rect 25197 -1521 25284 -1513
rect 25151 -1547 25284 -1521
rect 24894 -1613 24928 -1597
rect 24636 -1621 24839 -1615
rect 24962 -1615 24978 -1581
rect 25012 -1615 25033 -1581
rect 25072 -1589 25082 -1555
rect 25250 -1555 25284 -1547
rect 25072 -1605 25116 -1589
rect 24962 -1657 25033 -1615
rect 25150 -1615 25166 -1581
rect 25200 -1615 25216 -1581
rect 25250 -1605 25284 -1589
rect 25150 -1657 25216 -1615
rect 8575 -1715 8604 -1657
rect 8638 -1715 8696 -1657
rect 8730 -1715 8788 -1657
rect 8822 -1715 8880 -1657
rect 8914 -1715 8972 -1657
rect 9006 -1715 9064 -1657
rect 9098 -1715 9156 -1657
rect 9190 -1715 9248 -1657
rect 9282 -1715 9340 -1657
rect 9374 -1715 9432 -1657
rect 9466 -1715 9524 -1657
rect 9558 -1715 9616 -1657
rect 9650 -1715 9708 -1657
rect 9742 -1715 9800 -1657
rect 9834 -1715 9892 -1657
rect 9926 -1715 9984 -1657
rect 10018 -1715 10076 -1657
rect 10110 -1715 10168 -1657
rect 10202 -1715 10260 -1657
rect 10294 -1715 10352 -1657
rect 10386 -1715 10444 -1657
rect 10478 -1715 10536 -1657
rect 10570 -1715 10628 -1657
rect 10662 -1715 10720 -1657
rect 10754 -1715 10812 -1657
rect 10846 -1715 10904 -1657
rect 10938 -1715 10996 -1657
rect 11030 -1715 11088 -1657
rect 11122 -1715 11180 -1657
rect 11214 -1715 11272 -1657
rect 11306 -1715 11364 -1657
rect 11398 -1715 11456 -1657
rect 11490 -1715 11548 -1657
rect 11582 -1715 11640 -1657
rect 11674 -1715 11732 -1657
rect 11766 -1715 11824 -1657
rect 11858 -1715 11916 -1657
rect 11950 -1715 12008 -1657
rect 12042 -1715 12100 -1657
rect 12134 -1715 12192 -1657
rect 12226 -1715 12284 -1657
rect 12318 -1715 12376 -1657
rect 12410 -1715 12468 -1657
rect 12502 -1715 12560 -1657
rect 12594 -1715 12652 -1657
rect 12686 -1715 12744 -1657
rect 12778 -1715 12836 -1657
rect 12870 -1715 12928 -1657
rect 12962 -1715 13020 -1657
rect 13054 -1715 13112 -1657
rect 13146 -1715 13204 -1657
rect 13238 -1715 13296 -1657
rect 13330 -1715 13388 -1657
rect 13422 -1715 13480 -1657
rect 13514 -1715 13572 -1657
rect 13606 -1715 13664 -1657
rect 13698 -1715 13756 -1657
rect 13790 -1715 13848 -1657
rect 13882 -1715 13940 -1657
rect 13974 -1715 14032 -1657
rect 14066 -1715 14124 -1657
rect 14158 -1715 14216 -1657
rect 14250 -1715 14308 -1657
rect 14342 -1715 14400 -1657
rect 14434 -1715 14492 -1657
rect 14526 -1715 14584 -1657
rect 14618 -1715 14676 -1657
rect 14710 -1715 14768 -1657
rect 14802 -1715 14860 -1657
rect 14894 -1715 14952 -1657
rect 14986 -1715 15044 -1657
rect 15078 -1715 15136 -1657
rect 15170 -1715 15228 -1657
rect 15262 -1715 15320 -1657
rect 15354 -1715 15412 -1657
rect 15446 -1715 15504 -1657
rect 15538 -1715 15596 -1657
rect 15630 -1715 15688 -1657
rect 15722 -1715 15780 -1657
rect 15814 -1715 15872 -1657
rect 15906 -1715 15964 -1657
rect 15998 -1715 16056 -1657
rect 16090 -1715 16148 -1657
rect 16182 -1715 16240 -1657
rect 16274 -1715 16332 -1657
rect 16366 -1715 16424 -1657
rect 16458 -1715 16516 -1657
rect 16550 -1715 16608 -1657
rect 16642 -1715 16700 -1657
rect 16734 -1715 16792 -1657
rect 16826 -1715 16884 -1657
rect 16918 -1715 16976 -1657
rect 17010 -1715 17068 -1657
rect 17102 -1715 17160 -1657
rect 17194 -1715 17252 -1657
rect 17286 -1715 17344 -1657
rect 17378 -1715 17436 -1657
rect 17470 -1715 17528 -1657
rect 17562 -1715 17620 -1657
rect 17654 -1715 17712 -1657
rect 17746 -1715 17804 -1657
rect 17838 -1715 17896 -1657
rect 17930 -1715 17988 -1657
rect 18022 -1715 18080 -1657
rect 18114 -1715 18172 -1657
rect 18206 -1715 18264 -1657
rect 18298 -1715 18356 -1657
rect 18390 -1715 18448 -1657
rect 18482 -1715 18540 -1657
rect 18574 -1715 18632 -1657
rect 18666 -1715 18724 -1657
rect 18758 -1715 18816 -1657
rect 18850 -1715 18908 -1657
rect 18942 -1715 19000 -1657
rect 19034 -1715 19092 -1657
rect 19126 -1715 19184 -1657
rect 19218 -1715 19276 -1657
rect 19310 -1715 19368 -1657
rect 19402 -1715 19460 -1657
rect 19494 -1715 19552 -1657
rect 19586 -1715 19644 -1657
rect 19678 -1715 19736 -1657
rect 19770 -1715 19828 -1657
rect 19862 -1715 19920 -1657
rect 19954 -1715 20012 -1657
rect 20046 -1715 20104 -1657
rect 20138 -1715 20196 -1657
rect 20230 -1715 20288 -1657
rect 20322 -1715 20380 -1657
rect 20414 -1715 20472 -1657
rect 20506 -1715 20564 -1657
rect 20598 -1715 20656 -1657
rect 20690 -1715 20748 -1657
rect 20782 -1715 20840 -1657
rect 20874 -1715 20932 -1657
rect 20966 -1715 21024 -1657
rect 21058 -1715 21116 -1657
rect 21150 -1715 21208 -1657
rect 21242 -1715 21300 -1657
rect 21334 -1715 21392 -1657
rect 21426 -1715 21484 -1657
rect 21518 -1715 21576 -1657
rect 21610 -1715 21668 -1657
rect 21702 -1715 21760 -1657
rect 21794 -1715 21852 -1657
rect 21886 -1715 21944 -1657
rect 21978 -1715 22036 -1657
rect 22070 -1715 22128 -1657
rect 22162 -1715 22220 -1657
rect 22254 -1715 22312 -1657
rect 22346 -1715 22404 -1657
rect 22438 -1715 22496 -1657
rect 22530 -1715 22588 -1657
rect 22622 -1715 22680 -1657
rect 22714 -1715 22772 -1657
rect 22806 -1715 22864 -1657
rect 22898 -1715 22956 -1657
rect 22990 -1715 23048 -1657
rect 23082 -1715 23140 -1657
rect 23174 -1715 23232 -1657
rect 23266 -1715 23324 -1657
rect 23358 -1715 23416 -1657
rect 23450 -1715 23508 -1657
rect 23542 -1715 23600 -1657
rect 23634 -1715 23692 -1657
rect 23726 -1715 23784 -1657
rect 23818 -1715 23876 -1657
rect 23910 -1715 23968 -1657
rect 24002 -1715 24060 -1657
rect 24094 -1715 24152 -1657
rect 24186 -1715 24244 -1657
rect 24278 -1715 24336 -1657
rect 24370 -1715 24428 -1657
rect 24462 -1715 24520 -1657
rect 24554 -1715 24612 -1657
rect 24646 -1715 24704 -1657
rect 24738 -1715 24796 -1657
rect 24830 -1715 24888 -1657
rect 24922 -1715 24980 -1657
rect 25014 -1715 25072 -1657
rect 25106 -1715 25164 -1657
rect 25198 -1715 25256 -1657
rect 25290 -1715 25319 -1657
<< viali >>
rect 13816 13521 13850 13581
rect 13904 13521 13938 13581
rect 14064 13571 14096 13605
rect 14096 13571 14098 13605
rect 14144 13571 14176 13605
rect 14176 13571 14178 13605
rect 14224 13571 14256 13605
rect 14256 13571 14258 13605
rect 14304 13571 14336 13605
rect 14336 13571 14338 13605
rect 14384 13571 14416 13605
rect 14416 13571 14418 13605
rect 14464 13571 14496 13605
rect 14496 13571 14498 13605
rect 14796 13574 14828 13608
rect 14828 13574 14830 13608
rect 14876 13574 14908 13608
rect 14908 13574 14910 13608
rect 14956 13574 14988 13608
rect 14988 13574 14990 13608
rect 15036 13574 15068 13608
rect 15068 13574 15070 13608
rect 15116 13574 15148 13608
rect 15148 13574 15150 13608
rect 15196 13574 15228 13608
rect 15228 13574 15230 13608
rect 15398 13574 15400 13608
rect 15400 13574 15432 13608
rect 15478 13574 15480 13608
rect 15480 13574 15512 13608
rect 15558 13574 15560 13608
rect 15560 13574 15592 13608
rect 15638 13574 15640 13608
rect 15640 13574 15672 13608
rect 15718 13574 15720 13608
rect 15720 13574 15752 13608
rect 15798 13574 15800 13608
rect 15800 13574 15832 13608
rect 16008 13574 16040 13608
rect 16040 13574 16042 13608
rect 16088 13574 16120 13608
rect 16120 13574 16122 13608
rect 16168 13574 16200 13608
rect 16200 13574 16202 13608
rect 16248 13574 16280 13608
rect 16280 13574 16282 13608
rect 16328 13574 16360 13608
rect 16360 13574 16362 13608
rect 16408 13574 16440 13608
rect 16440 13574 16442 13608
rect 16610 13574 16612 13608
rect 16612 13574 16644 13608
rect 16690 13574 16692 13608
rect 16692 13574 16724 13608
rect 16770 13574 16772 13608
rect 16772 13574 16804 13608
rect 16850 13574 16852 13608
rect 16852 13574 16884 13608
rect 16930 13574 16932 13608
rect 16932 13574 16964 13608
rect 17010 13574 17012 13608
rect 17012 13574 17044 13608
rect 17220 13574 17252 13608
rect 17252 13574 17254 13608
rect 17300 13574 17332 13608
rect 17332 13574 17334 13608
rect 17380 13574 17412 13608
rect 17412 13574 17414 13608
rect 17460 13574 17492 13608
rect 17492 13574 17494 13608
rect 17540 13574 17572 13608
rect 17572 13574 17574 13608
rect 17620 13574 17652 13608
rect 17652 13574 17654 13608
rect 17822 13574 17824 13608
rect 17824 13574 17856 13608
rect 17902 13574 17904 13608
rect 17904 13574 17936 13608
rect 17982 13574 17984 13608
rect 17984 13574 18016 13608
rect 18062 13574 18064 13608
rect 18064 13574 18096 13608
rect 18142 13574 18144 13608
rect 18144 13574 18176 13608
rect 18222 13574 18224 13608
rect 18224 13574 18256 13608
rect 18432 13574 18464 13608
rect 18464 13574 18466 13608
rect 18512 13574 18544 13608
rect 18544 13574 18546 13608
rect 18592 13574 18624 13608
rect 18624 13574 18626 13608
rect 18672 13574 18704 13608
rect 18704 13574 18706 13608
rect 18752 13574 18784 13608
rect 18784 13574 18786 13608
rect 18832 13574 18864 13608
rect 18864 13574 18866 13608
rect 19034 13574 19036 13608
rect 19036 13574 19068 13608
rect 19114 13574 19116 13608
rect 19116 13574 19148 13608
rect 19194 13574 19196 13608
rect 19196 13574 19228 13608
rect 19274 13574 19276 13608
rect 19276 13574 19308 13608
rect 19354 13574 19356 13608
rect 19356 13574 19388 13608
rect 19434 13574 19436 13608
rect 19436 13574 19468 13608
rect 13816 13383 13850 13443
rect 19776 13523 19810 13557
rect 20253 13526 20287 13560
rect 20525 13521 20559 13581
rect 20613 13521 20647 13581
rect 20773 13571 20805 13605
rect 20805 13571 20807 13605
rect 20853 13571 20885 13605
rect 20885 13571 20887 13605
rect 20933 13571 20965 13605
rect 20965 13571 20967 13605
rect 21013 13571 21045 13605
rect 21045 13571 21047 13605
rect 21093 13571 21125 13605
rect 21125 13571 21127 13605
rect 21173 13571 21205 13605
rect 21205 13571 21207 13605
rect 21505 13574 21537 13608
rect 21537 13574 21539 13608
rect 21585 13574 21617 13608
rect 21617 13574 21619 13608
rect 21665 13574 21697 13608
rect 21697 13574 21699 13608
rect 21745 13574 21777 13608
rect 21777 13574 21779 13608
rect 21825 13574 21857 13608
rect 21857 13574 21859 13608
rect 21905 13574 21937 13608
rect 21937 13574 21939 13608
rect 22107 13574 22109 13608
rect 22109 13574 22141 13608
rect 22187 13574 22189 13608
rect 22189 13574 22221 13608
rect 22267 13574 22269 13608
rect 22269 13574 22301 13608
rect 22347 13574 22349 13608
rect 22349 13574 22381 13608
rect 22427 13574 22429 13608
rect 22429 13574 22461 13608
rect 22507 13574 22509 13608
rect 22509 13574 22541 13608
rect 22717 13574 22749 13608
rect 22749 13574 22751 13608
rect 22797 13574 22829 13608
rect 22829 13574 22831 13608
rect 22877 13574 22909 13608
rect 22909 13574 22911 13608
rect 22957 13574 22989 13608
rect 22989 13574 22991 13608
rect 23037 13574 23069 13608
rect 23069 13574 23071 13608
rect 23117 13574 23149 13608
rect 23149 13574 23151 13608
rect 23319 13574 23321 13608
rect 23321 13574 23353 13608
rect 23399 13574 23401 13608
rect 23401 13574 23433 13608
rect 23479 13574 23481 13608
rect 23481 13574 23513 13608
rect 23559 13574 23561 13608
rect 23561 13574 23593 13608
rect 23639 13574 23641 13608
rect 23641 13574 23673 13608
rect 23719 13574 23721 13608
rect 23721 13574 23753 13608
rect 23929 13574 23961 13608
rect 23961 13574 23963 13608
rect 24009 13574 24041 13608
rect 24041 13574 24043 13608
rect 24089 13574 24121 13608
rect 24121 13574 24123 13608
rect 24169 13574 24201 13608
rect 24201 13574 24203 13608
rect 24249 13574 24281 13608
rect 24281 13574 24283 13608
rect 24329 13574 24361 13608
rect 24361 13574 24363 13608
rect 24531 13574 24533 13608
rect 24533 13574 24565 13608
rect 24611 13574 24613 13608
rect 24613 13574 24645 13608
rect 24691 13574 24693 13608
rect 24693 13574 24725 13608
rect 24771 13574 24773 13608
rect 24773 13574 24805 13608
rect 24851 13574 24853 13608
rect 24853 13574 24885 13608
rect 24931 13574 24933 13608
rect 24933 13574 24965 13608
rect 25141 13574 25173 13608
rect 25173 13574 25175 13608
rect 25221 13574 25253 13608
rect 25253 13574 25255 13608
rect 25301 13574 25333 13608
rect 25333 13574 25335 13608
rect 25381 13574 25413 13608
rect 25413 13574 25415 13608
rect 25461 13574 25493 13608
rect 25493 13574 25495 13608
rect 25541 13574 25573 13608
rect 25573 13574 25575 13608
rect 25743 13574 25745 13608
rect 25745 13574 25777 13608
rect 25823 13574 25825 13608
rect 25825 13574 25857 13608
rect 25903 13574 25905 13608
rect 25905 13574 25937 13608
rect 25983 13574 25985 13608
rect 25985 13574 26017 13608
rect 26063 13574 26065 13608
rect 26065 13574 26097 13608
rect 26143 13574 26145 13608
rect 26145 13574 26177 13608
rect 13904 13383 13938 13443
rect 19781 13379 19815 13413
rect 20242 13354 20276 13388
rect 20525 13383 20559 13443
rect 26485 13523 26519 13557
rect 20613 13383 20647 13443
rect 26490 13379 26524 13413
rect 13816 13245 13850 13305
rect 13904 13245 13938 13305
rect 19782 13227 19816 13261
rect 20525 13245 20559 13305
rect 20613 13245 20647 13305
rect 26491 13227 26525 13261
rect 2928 13046 2962 13106
rect 3016 13046 3050 13106
rect 3176 13096 3208 13130
rect 3208 13096 3210 13130
rect 3256 13096 3288 13130
rect 3288 13096 3290 13130
rect 3336 13096 3368 13130
rect 3368 13096 3370 13130
rect 3416 13096 3448 13130
rect 3448 13096 3450 13130
rect 3496 13096 3528 13130
rect 3528 13096 3530 13130
rect 3576 13096 3608 13130
rect 3608 13096 3610 13130
rect 3908 13099 3940 13133
rect 3940 13099 3942 13133
rect 3988 13099 4020 13133
rect 4020 13099 4022 13133
rect 4068 13099 4100 13133
rect 4100 13099 4102 13133
rect 4148 13099 4180 13133
rect 4180 13099 4182 13133
rect 4228 13099 4260 13133
rect 4260 13099 4262 13133
rect 4308 13099 4340 13133
rect 4340 13099 4342 13133
rect 4510 13099 4512 13133
rect 4512 13099 4544 13133
rect 4590 13099 4592 13133
rect 4592 13099 4624 13133
rect 4670 13099 4672 13133
rect 4672 13099 4704 13133
rect 4750 13099 4752 13133
rect 4752 13099 4784 13133
rect 4830 13099 4832 13133
rect 4832 13099 4864 13133
rect 4910 13099 4912 13133
rect 4912 13099 4944 13133
rect 5120 13099 5152 13133
rect 5152 13099 5154 13133
rect 5200 13099 5232 13133
rect 5232 13099 5234 13133
rect 5280 13099 5312 13133
rect 5312 13099 5314 13133
rect 5360 13099 5392 13133
rect 5392 13099 5394 13133
rect 5440 13099 5472 13133
rect 5472 13099 5474 13133
rect 5520 13099 5552 13133
rect 5552 13099 5554 13133
rect 5722 13099 5724 13133
rect 5724 13099 5756 13133
rect 5802 13099 5804 13133
rect 5804 13099 5836 13133
rect 5882 13099 5884 13133
rect 5884 13099 5916 13133
rect 5962 13099 5964 13133
rect 5964 13099 5996 13133
rect 6042 13099 6044 13133
rect 6044 13099 6076 13133
rect 6122 13099 6124 13133
rect 6124 13099 6156 13133
rect 6332 13099 6364 13133
rect 6364 13099 6366 13133
rect 6412 13099 6444 13133
rect 6444 13099 6446 13133
rect 6492 13099 6524 13133
rect 6524 13099 6526 13133
rect 6572 13099 6604 13133
rect 6604 13099 6606 13133
rect 6652 13099 6684 13133
rect 6684 13099 6686 13133
rect 6732 13099 6764 13133
rect 6764 13099 6766 13133
rect 6934 13099 6936 13133
rect 6936 13099 6968 13133
rect 7014 13099 7016 13133
rect 7016 13099 7048 13133
rect 7094 13099 7096 13133
rect 7096 13099 7128 13133
rect 7174 13099 7176 13133
rect 7176 13099 7208 13133
rect 7254 13099 7256 13133
rect 7256 13099 7288 13133
rect 7334 13099 7336 13133
rect 7336 13099 7368 13133
rect 7544 13099 7576 13133
rect 7576 13099 7578 13133
rect 7624 13099 7656 13133
rect 7656 13099 7658 13133
rect 7704 13099 7736 13133
rect 7736 13099 7738 13133
rect 7784 13099 7816 13133
rect 7816 13099 7818 13133
rect 7864 13099 7896 13133
rect 7896 13099 7898 13133
rect 7944 13099 7976 13133
rect 7976 13099 7978 13133
rect 8146 13099 8148 13133
rect 8148 13099 8180 13133
rect 8226 13099 8228 13133
rect 8228 13099 8260 13133
rect 8306 13099 8308 13133
rect 8308 13099 8340 13133
rect 8386 13099 8388 13133
rect 8388 13099 8420 13133
rect 8466 13099 8468 13133
rect 8468 13099 8500 13133
rect 8546 13099 8548 13133
rect 8548 13099 8580 13133
rect 13816 13107 13850 13167
rect 13904 13107 13938 13167
rect 20242 13162 20276 13196
rect 20525 13107 20559 13167
rect 20613 13107 20647 13167
rect 2928 12908 2962 12968
rect 8888 13048 8922 13082
rect 19782 13057 19816 13091
rect 3016 12908 3050 12968
rect 13303 12976 13337 13010
rect 13395 12976 13429 13010
rect 13487 13005 13512 13010
rect 13512 13005 13521 13010
rect 13487 12976 13521 13005
rect 13579 12976 13613 13010
rect 13671 12976 13705 13010
rect 8893 12904 8927 12938
rect 2928 12770 2962 12830
rect 3016 12770 3050 12830
rect 8894 12752 8928 12786
rect 13431 12866 13465 12867
rect 13431 12833 13434 12866
rect 13434 12833 13465 12866
rect 2928 12632 2962 12692
rect 3016 12632 3050 12692
rect 13350 12698 13384 12702
rect 13350 12668 13354 12698
rect 13354 12668 13384 12698
rect 8894 12582 8928 12616
rect 2415 12501 2449 12535
rect 2507 12501 2541 12535
rect 2599 12530 2624 12535
rect 2624 12530 2633 12535
rect 2599 12501 2633 12530
rect 2691 12501 2725 12535
rect 2783 12501 2817 12535
rect 2543 12391 2577 12392
rect 2543 12358 2546 12391
rect 2546 12358 2577 12391
rect 2462 12223 2496 12227
rect 2462 12193 2466 12223
rect 2466 12193 2496 12223
rect 2652 12323 2686 12337
rect 2652 12303 2686 12323
rect 2928 12494 2962 12554
rect 3016 12494 3050 12554
rect 2928 12356 2962 12416
rect 3016 12356 3050 12416
rect 8893 12425 8927 12459
rect 10911 12432 10945 12466
rect 11003 12432 11037 12466
rect 11095 12432 11129 12466
rect 11187 12432 11221 12466
rect 11279 12432 11313 12466
rect 11371 12432 11405 12466
rect 11463 12432 11497 12466
rect 11555 12432 11589 12466
rect 11647 12432 11681 12466
rect 11739 12432 11773 12466
rect 11831 12432 11865 12466
rect 11923 12432 11957 12466
rect 12015 12432 12049 12466
rect 12107 12432 12141 12466
rect 12199 12432 12233 12466
rect 12291 12432 12325 12466
rect 12383 12432 12417 12466
rect 12475 12432 12509 12466
rect 12567 12432 12601 12466
rect 12659 12432 12693 12466
rect 12751 12432 12785 12466
rect 12843 12432 12877 12466
rect 12935 12432 12969 12466
rect 13027 12432 13061 12466
rect 13119 12432 13153 12466
rect 13540 12798 13574 12812
rect 13540 12778 13574 12798
rect 13816 12969 13850 13029
rect 26491 13057 26525 13091
rect 13904 12969 13938 13029
rect 20012 12976 20046 13010
rect 20104 12976 20138 13010
rect 20196 13005 20221 13010
rect 20221 13005 20230 13010
rect 20196 12976 20230 13005
rect 20288 12976 20322 13010
rect 20380 12976 20414 13010
rect 13816 12831 13850 12891
rect 13904 12831 13938 12891
rect 19781 12900 19815 12934
rect 13860 12738 13894 12772
rect 20140 12866 20174 12867
rect 20140 12833 20143 12866
rect 20143 12833 20174 12866
rect 13624 12698 13658 12701
rect 13624 12667 13654 12698
rect 13654 12667 13658 12698
rect 13763 12668 13797 12702
rect 20059 12698 20093 12702
rect 20059 12668 20063 12698
rect 20063 12668 20093 12698
rect 13801 12575 13835 12609
rect 14060 12593 14094 12627
rect 14061 12500 14095 12534
rect 14502 12495 14536 12529
rect 15234 12498 15268 12532
rect 15360 12498 15394 12532
rect 16446 12498 16480 12532
rect 16572 12498 16606 12532
rect 17658 12498 17692 12532
rect 17784 12498 17818 12532
rect 18870 12498 18904 12532
rect 18996 12498 19030 12532
rect 19601 12520 19635 12580
rect 19689 12520 19723 12580
rect 20249 12798 20283 12812
rect 20249 12778 20283 12798
rect 20525 12969 20559 13029
rect 20613 12969 20647 13029
rect 20525 12831 20559 12891
rect 20613 12831 20647 12891
rect 26490 12900 26524 12934
rect 20569 12738 20603 12772
rect 20333 12698 20367 12701
rect 20333 12667 20363 12698
rect 20363 12667 20367 12698
rect 20472 12668 20506 12702
rect 20510 12575 20544 12609
rect 20769 12593 20803 12627
rect 20770 12500 20804 12534
rect 21211 12495 21245 12529
rect 21943 12498 21977 12532
rect 22069 12498 22103 12532
rect 23155 12498 23189 12532
rect 23281 12498 23315 12532
rect 24367 12498 24401 12532
rect 24493 12498 24527 12532
rect 25579 12498 25613 12532
rect 25705 12498 25739 12532
rect 26310 12520 26344 12580
rect 26398 12520 26432 12580
rect 13211 12432 13245 12466
rect 13303 12432 13337 12466
rect 13395 12437 13429 12466
rect 13487 12437 13521 12466
rect 13395 12432 13402 12437
rect 13402 12432 13429 12437
rect 13487 12432 13520 12437
rect 13520 12432 13521 12437
rect 13579 12432 13613 12466
rect 2972 12263 3006 12297
rect 2736 12223 2770 12226
rect 2736 12192 2766 12223
rect 2766 12192 2770 12223
rect 2875 12193 2909 12227
rect 2913 12100 2947 12134
rect 3172 12118 3206 12152
rect 9090 12124 9124 12158
rect 9182 12124 9216 12158
rect 9274 12124 9308 12158
rect 10912 12185 10914 12217
rect 10914 12185 10946 12217
rect 10912 12183 10946 12185
rect 3173 12025 3207 12059
rect 3614 12020 3648 12054
rect 4346 12023 4380 12057
rect 4472 12023 4506 12057
rect 5558 12023 5592 12057
rect 5684 12023 5718 12057
rect 6770 12023 6804 12057
rect 6896 12023 6930 12057
rect 7982 12023 8016 12057
rect 8108 12023 8142 12057
rect 8713 12045 8747 12105
rect 8801 12045 8835 12105
rect 2415 11957 2449 11991
rect 2507 11962 2541 11991
rect 2599 11962 2633 11991
rect 2507 11957 2514 11962
rect 2514 11957 2541 11962
rect 2599 11957 2632 11962
rect 2632 11957 2633 11962
rect 2691 11957 2725 11991
rect 2783 11957 2817 11991
rect 3570 11901 3604 11961
rect 3658 11904 3692 11964
rect 4302 11904 4336 11964
rect 4407 11904 4441 11964
rect 4516 11904 4550 11964
rect 5514 11904 5548 11964
rect 5618 11904 5652 11964
rect 5728 11904 5762 11964
rect 6726 11904 6760 11964
rect 6831 11904 6865 11964
rect 6940 11904 6974 11964
rect 7938 11904 7972 11964
rect 8045 11904 8079 11964
rect 8152 11904 8186 11964
rect 8713 11907 8747 11967
rect 8801 11907 8835 11967
rect 8897 11907 8931 11967
rect 8993 11907 9027 11967
rect 11004 12058 11038 12092
rect 11096 12262 11130 12296
rect 11263 12155 11297 12189
rect 11460 12280 11494 12296
rect 11460 12262 11478 12280
rect 11478 12262 11494 12280
rect 11648 12270 11682 12296
rect 11648 12262 11650 12270
rect 11650 12262 11682 12270
rect 11372 12058 11406 12092
rect 12108 12194 12142 12228
rect 12016 12126 12050 12160
rect 12108 12084 12129 12092
rect 12129 12084 12142 12092
rect 12108 12058 12142 12084
rect 12384 12270 12418 12296
rect 12384 12262 12393 12270
rect 12393 12262 12418 12270
rect 12768 12196 12770 12225
rect 12770 12196 12802 12225
rect 12768 12191 12802 12196
rect 12660 12126 12694 12160
rect 12935 12001 12956 12026
rect 12956 12001 12969 12026
rect 12935 11992 12969 12001
rect 13671 12432 13705 12466
rect 14458 12376 14492 12436
rect 14546 12379 14580 12439
rect 15190 12379 15224 12439
rect 15295 12379 15329 12439
rect 15404 12379 15438 12439
rect 16402 12379 16436 12439
rect 16506 12379 16540 12439
rect 16616 12379 16650 12439
rect 17614 12379 17648 12439
rect 17719 12379 17753 12439
rect 17828 12379 17862 12439
rect 18826 12379 18860 12439
rect 18933 12379 18967 12439
rect 19040 12379 19074 12439
rect 19601 12382 19635 12442
rect 19689 12382 19723 12442
rect 19785 12382 19819 12442
rect 19881 12382 19915 12442
rect 20012 12432 20046 12466
rect 20104 12437 20138 12466
rect 20196 12437 20230 12466
rect 20104 12432 20111 12437
rect 20111 12432 20138 12437
rect 20196 12432 20229 12437
rect 20229 12432 20230 12437
rect 20288 12432 20322 12466
rect 20380 12432 20414 12466
rect 21167 12376 21201 12436
rect 21255 12379 21289 12439
rect 21899 12379 21933 12439
rect 22004 12379 22038 12439
rect 22113 12379 22147 12439
rect 23111 12379 23145 12439
rect 23215 12379 23249 12439
rect 23325 12379 23359 12439
rect 24323 12379 24357 12439
rect 24428 12379 24462 12439
rect 24537 12379 24571 12439
rect 25535 12379 25569 12439
rect 25642 12379 25676 12439
rect 25749 12379 25783 12439
rect 26310 12382 26344 12442
rect 26398 12382 26432 12442
rect 26494 12382 26528 12442
rect 26590 12382 26624 12442
rect 13221 12320 13239 12324
rect 13239 12320 13255 12324
rect 13221 12290 13255 12320
rect 19530 12291 19564 12325
rect 19737 12289 19771 12323
rect 26239 12291 26273 12325
rect 26446 12289 26480 12323
rect 14811 12178 14845 12238
rect 14901 12178 14935 12238
rect 15543 12178 15577 12238
rect 15650 12178 15684 12238
rect 15753 12178 15787 12238
rect 16755 12178 16789 12238
rect 16861 12178 16895 12238
rect 16965 12178 16999 12238
rect 18093 12178 18127 12238
rect 18201 12178 18235 12238
rect 18303 12178 18337 12238
rect 18948 12178 18982 12238
rect 19037 12178 19071 12238
rect 19601 12179 19635 12239
rect 19689 12179 19723 12239
rect 19785 12179 19819 12239
rect 19881 12179 19915 12239
rect 21520 12178 21554 12238
rect 21610 12178 21644 12238
rect 22252 12178 22286 12238
rect 22359 12178 22393 12238
rect 22462 12178 22496 12238
rect 23464 12178 23498 12238
rect 23570 12178 23604 12238
rect 23674 12178 23708 12238
rect 24802 12178 24836 12238
rect 24910 12178 24944 12238
rect 25012 12178 25046 12238
rect 25657 12178 25691 12238
rect 25746 12178 25780 12238
rect 26310 12179 26344 12239
rect 26398 12179 26432 12239
rect 26494 12179 26528 12239
rect 26590 12179 26624 12239
rect 13871 12104 13905 12138
rect 14855 12094 14889 12128
rect 15587 12094 15621 12128
rect 15709 12094 15743 12128
rect 16799 12094 16833 12128
rect 16921 12094 16955 12128
rect 18137 12094 18171 12128
rect 18259 12094 18293 12128
rect 18993 12094 19027 12128
rect 13215 12034 13249 12044
rect 13215 12010 13239 12034
rect 13239 12010 13249 12034
rect 13791 11994 13825 12054
rect 13951 11994 13985 12054
rect 19601 12041 19635 12101
rect 20580 12104 20614 12138
rect 19689 12041 19723 12101
rect 21564 12094 21598 12128
rect 22296 12094 22330 12128
rect 22418 12094 22452 12128
rect 23508 12094 23542 12128
rect 23630 12094 23664 12128
rect 24846 12094 24880 12128
rect 24968 12094 25002 12128
rect 25702 12094 25736 12128
rect 20500 11994 20534 12054
rect 20660 11994 20694 12054
rect 26310 12041 26344 12101
rect 26398 12041 26432 12101
rect 8642 11816 8676 11850
rect 8849 11814 8883 11848
rect 9134 11846 9168 11850
rect 9134 11816 9141 11846
rect 9141 11816 9168 11846
rect 10911 11888 10945 11922
rect 11003 11888 11037 11922
rect 11095 11888 11129 11922
rect 11187 11888 11221 11922
rect 11279 11888 11313 11922
rect 11371 11888 11405 11922
rect 11463 11888 11497 11922
rect 9236 11815 9270 11849
rect 11555 11888 11589 11922
rect 11647 11888 11681 11922
rect 11739 11888 11773 11922
rect 11831 11888 11865 11922
rect 11923 11888 11957 11922
rect 12015 11888 12049 11922
rect 12107 11888 12141 11922
rect 12199 11888 12233 11922
rect 12291 11888 12325 11922
rect 12383 11888 12417 11922
rect 12475 11888 12509 11922
rect 12567 11888 12601 11922
rect 12659 11888 12693 11922
rect 12751 11888 12785 11922
rect 12843 11888 12877 11922
rect 12935 11888 12969 11922
rect 13027 11888 13061 11922
rect 13119 11888 13153 11922
rect 13211 11888 13245 11922
rect 13791 11856 13825 11916
rect 13951 11856 13985 11916
rect 20500 11856 20534 11916
rect 20660 11856 20694 11916
rect 3923 11703 3957 11763
rect 4013 11703 4047 11763
rect 4655 11703 4689 11763
rect 4762 11703 4796 11763
rect 4865 11703 4899 11763
rect 5867 11703 5901 11763
rect 5973 11703 6007 11763
rect 6077 11703 6111 11763
rect 7205 11703 7239 11763
rect 7313 11703 7347 11763
rect 7415 11703 7449 11763
rect 8060 11703 8094 11763
rect 8149 11703 8183 11763
rect 8713 11704 8747 11764
rect 8801 11704 8835 11764
rect 8897 11704 8931 11764
rect 8993 11704 9027 11764
rect 10911 11792 10945 11826
rect 11003 11792 11037 11826
rect 11095 11792 11129 11826
rect 11187 11792 11221 11826
rect 11279 11792 11313 11826
rect 11371 11792 11405 11826
rect 2983 11629 3017 11663
rect 3967 11619 4001 11653
rect 4699 11619 4733 11653
rect 4821 11619 4855 11653
rect 5911 11619 5945 11653
rect 6033 11619 6067 11653
rect 7249 11619 7283 11653
rect 7371 11619 7405 11653
rect 8105 11619 8139 11653
rect 2903 11519 2937 11579
rect 3063 11519 3097 11579
rect 8713 11566 8747 11626
rect 8801 11566 8835 11626
rect 9090 11580 9124 11614
rect 9182 11580 9216 11614
rect 9274 11580 9308 11614
rect 11044 11648 11076 11651
rect 11076 11648 11078 11651
rect 11044 11617 11078 11648
rect 11319 11716 11352 11727
rect 11352 11716 11353 11727
rect 11319 11693 11353 11716
rect 13791 11718 13825 11778
rect 13951 11718 13985 11778
rect 20500 11718 20534 11778
rect 20660 11718 20694 11778
rect 10957 11514 10991 11522
rect 10957 11488 10962 11514
rect 10962 11488 10991 11514
rect 2903 11381 2937 11441
rect 3063 11381 3097 11441
rect 11228 11514 11262 11517
rect 11228 11483 11238 11514
rect 11238 11483 11262 11514
rect 2903 11243 2937 11303
rect 3063 11243 3097 11303
rect 13317 11543 13375 11594
rect 13791 11580 13825 11640
rect 13951 11580 13985 11640
rect 20500 11580 20534 11640
rect 20660 11580 20694 11640
rect 13791 11442 13825 11502
rect 13951 11442 13985 11502
rect 20500 11442 20534 11502
rect 20660 11442 20694 11502
rect 13791 11304 13825 11364
rect 13951 11304 13985 11364
rect 20500 11304 20534 11364
rect 20660 11304 20694 11364
rect 10911 11248 10945 11282
rect 11003 11248 11037 11282
rect 11095 11248 11129 11282
rect 11187 11248 11221 11282
rect 11279 11248 11313 11282
rect 11371 11248 11405 11282
rect 2903 11105 2937 11165
rect 3063 11105 3097 11165
rect 13791 11166 13825 11226
rect 13951 11166 13985 11226
rect 20500 11166 20534 11226
rect 20660 11166 20694 11226
rect 2903 10967 2937 11027
rect 3063 10967 3097 11027
rect 13791 11028 13825 11088
rect 13951 11028 13985 11088
rect 14492 11007 14526 11041
rect 14572 11007 14606 11041
rect 14652 11007 14686 11041
rect 14732 11007 14766 11041
rect 15224 11007 15258 11041
rect 15304 11007 15338 11041
rect 15384 11007 15418 11041
rect 15464 11007 15498 11041
rect 15832 11007 15866 11041
rect 15912 11007 15946 11041
rect 15992 11007 16026 11041
rect 16072 11007 16106 11041
rect 16436 11007 16470 11041
rect 16516 11007 16550 11041
rect 16596 11007 16630 11041
rect 16676 11007 16710 11041
rect 17044 11007 17078 11041
rect 17124 11007 17158 11041
rect 17204 11007 17238 11041
rect 17284 11007 17318 11041
rect 17774 11007 17808 11041
rect 17854 11007 17888 11041
rect 17934 11007 17968 11041
rect 18014 11007 18048 11041
rect 18382 11007 18416 11041
rect 18462 11007 18496 11041
rect 18542 11007 18576 11041
rect 18622 11007 18656 11041
rect 19116 11007 19150 11041
rect 19196 11007 19230 11041
rect 19276 11007 19310 11041
rect 19356 11007 19390 11041
rect 20500 11028 20534 11088
rect 20660 11028 20694 11088
rect 21201 11007 21235 11041
rect 21281 11007 21315 11041
rect 21361 11007 21395 11041
rect 21441 11007 21475 11041
rect 21933 11007 21967 11041
rect 22013 11007 22047 11041
rect 22093 11007 22127 11041
rect 22173 11007 22207 11041
rect 22541 11007 22575 11041
rect 22621 11007 22655 11041
rect 22701 11007 22735 11041
rect 22781 11007 22815 11041
rect 23145 11007 23179 11041
rect 23225 11007 23259 11041
rect 23305 11007 23339 11041
rect 23385 11007 23419 11041
rect 23753 11007 23787 11041
rect 23833 11007 23867 11041
rect 23913 11007 23947 11041
rect 23993 11007 24027 11041
rect 24483 11007 24517 11041
rect 24563 11007 24597 11041
rect 24643 11007 24677 11041
rect 24723 11007 24757 11041
rect 25091 11007 25125 11041
rect 25171 11007 25205 11041
rect 25251 11007 25285 11041
rect 25331 11007 25365 11041
rect 25825 11007 25859 11041
rect 25905 11007 25939 11041
rect 25985 11007 26019 11041
rect 26065 11007 26099 11041
rect 2903 10829 2937 10889
rect 3063 10829 3097 10889
rect 2903 10691 2937 10751
rect 3063 10691 3097 10751
rect 2903 10553 2937 10613
rect 3063 10553 3097 10613
rect 3604 10532 3638 10566
rect 3684 10532 3718 10566
rect 3764 10532 3798 10566
rect 3844 10532 3878 10566
rect 4336 10532 4370 10566
rect 4416 10532 4450 10566
rect 4496 10532 4530 10566
rect 4576 10532 4610 10566
rect 4944 10532 4978 10566
rect 5024 10532 5058 10566
rect 5104 10532 5138 10566
rect 5184 10532 5218 10566
rect 5548 10532 5582 10566
rect 5628 10532 5662 10566
rect 5708 10532 5742 10566
rect 5788 10532 5822 10566
rect 6156 10532 6190 10566
rect 6236 10532 6270 10566
rect 6316 10532 6350 10566
rect 6396 10532 6430 10566
rect 6886 10532 6920 10566
rect 6966 10532 7000 10566
rect 7046 10532 7080 10566
rect 7126 10532 7160 10566
rect 7494 10532 7528 10566
rect 7574 10532 7608 10566
rect 7654 10532 7688 10566
rect 7734 10532 7768 10566
rect 8228 10532 8262 10566
rect 8308 10532 8342 10566
rect 8388 10532 8422 10566
rect 8468 10532 8502 10566
rect 2903 10033 2937 10093
rect 3063 10033 3097 10093
rect 3604 10080 3638 10114
rect 3684 10080 3718 10114
rect 3764 10080 3798 10114
rect 3844 10080 3878 10114
rect 4336 10080 4370 10114
rect 4416 10080 4450 10114
rect 4496 10080 4530 10114
rect 4576 10080 4610 10114
rect 4944 10080 4978 10114
rect 5024 10080 5058 10114
rect 5104 10080 5138 10114
rect 5184 10080 5218 10114
rect 5548 10080 5582 10114
rect 5628 10080 5662 10114
rect 5708 10080 5742 10114
rect 5788 10080 5822 10114
rect 6156 10080 6190 10114
rect 6236 10080 6270 10114
rect 6316 10080 6350 10114
rect 6396 10080 6430 10114
rect 6886 10080 6920 10114
rect 6966 10080 7000 10114
rect 7046 10080 7080 10114
rect 7126 10080 7160 10114
rect 7494 10080 7528 10114
rect 7574 10080 7608 10114
rect 7654 10080 7688 10114
rect 7734 10080 7768 10114
rect 8228 10080 8262 10114
rect 8308 10080 8342 10114
rect 8388 10080 8422 10114
rect 8468 10080 8502 10114
rect 13789 10068 13823 10102
rect 13869 10068 13903 10102
rect 13949 10068 13983 10102
rect 14029 10068 14063 10102
rect 14523 10068 14557 10102
rect 14603 10068 14637 10102
rect 14683 10068 14717 10102
rect 14763 10068 14797 10102
rect 15131 10068 15165 10102
rect 15211 10068 15245 10102
rect 15291 10068 15325 10102
rect 15371 10068 15405 10102
rect 15861 10068 15895 10102
rect 15941 10068 15975 10102
rect 16021 10068 16055 10102
rect 16101 10068 16135 10102
rect 16469 10068 16503 10102
rect 16549 10068 16583 10102
rect 16629 10068 16663 10102
rect 16709 10068 16743 10102
rect 17073 10068 17107 10102
rect 17153 10068 17187 10102
rect 17233 10068 17267 10102
rect 17313 10068 17347 10102
rect 17681 10068 17715 10102
rect 17761 10068 17795 10102
rect 17841 10068 17875 10102
rect 17921 10068 17955 10102
rect 18413 10068 18447 10102
rect 18493 10068 18527 10102
rect 18573 10068 18607 10102
rect 18653 10068 18687 10102
rect 19194 10021 19228 10081
rect 2903 9895 2937 9955
rect 3063 9895 3097 9955
rect 19354 10021 19388 10081
rect 20498 10068 20532 10102
rect 20578 10068 20612 10102
rect 20658 10068 20692 10102
rect 20738 10068 20772 10102
rect 21232 10068 21266 10102
rect 21312 10068 21346 10102
rect 21392 10068 21426 10102
rect 21472 10068 21506 10102
rect 21840 10068 21874 10102
rect 21920 10068 21954 10102
rect 22000 10068 22034 10102
rect 22080 10068 22114 10102
rect 22570 10068 22604 10102
rect 22650 10068 22684 10102
rect 22730 10068 22764 10102
rect 22810 10068 22844 10102
rect 23178 10068 23212 10102
rect 23258 10068 23292 10102
rect 23338 10068 23372 10102
rect 23418 10068 23452 10102
rect 23782 10068 23816 10102
rect 23862 10068 23896 10102
rect 23942 10068 23976 10102
rect 24022 10068 24056 10102
rect 24390 10068 24424 10102
rect 24470 10068 24504 10102
rect 24550 10068 24584 10102
rect 24630 10068 24664 10102
rect 25122 10068 25156 10102
rect 25202 10068 25236 10102
rect 25282 10068 25316 10102
rect 25362 10068 25396 10102
rect 25903 10021 25937 10081
rect 26063 10021 26097 10081
rect 19194 9883 19228 9943
rect 19354 9883 19388 9943
rect 25903 9883 25937 9943
rect 26063 9883 26097 9943
rect 2903 9757 2937 9817
rect 3063 9757 3097 9817
rect 19194 9745 19228 9805
rect 19354 9745 19388 9805
rect 25903 9745 25937 9805
rect 26063 9745 26097 9805
rect 2903 9619 2937 9679
rect 3063 9619 3097 9679
rect 19194 9607 19228 9667
rect 19354 9607 19388 9667
rect 25903 9607 25937 9667
rect 26063 9607 26097 9667
rect 2903 9481 2937 9541
rect 3063 9481 3097 9541
rect 19194 9469 19228 9529
rect 19354 9469 19388 9529
rect 25903 9469 25937 9529
rect 26063 9469 26097 9529
rect 2903 9343 2937 9403
rect 3063 9343 3097 9403
rect 19194 9331 19228 9391
rect 19354 9331 19388 9391
rect 25903 9331 25937 9391
rect 26063 9331 26097 9391
rect 2903 9205 2937 9265
rect 3063 9205 3097 9265
rect 19194 9193 19228 9253
rect 19354 9193 19388 9253
rect 25903 9193 25937 9253
rect 26063 9193 26097 9253
rect 2903 9067 2937 9127
rect 3063 9067 3097 9127
rect 2983 8983 3017 9017
rect 3967 8993 4001 9027
rect 4699 8993 4733 9027
rect 4821 8993 4855 9027
rect 5911 8993 5945 9027
rect 6033 8993 6067 9027
rect 7249 8993 7283 9027
rect 7371 8993 7405 9027
rect 8105 8993 8139 9027
rect 8713 9020 8747 9080
rect 8801 9020 8835 9080
rect 9090 9034 9124 9068
rect 9182 9034 9216 9068
rect 9274 9034 9308 9068
rect 9346 9034 9380 9068
rect 9438 9067 9472 9068
rect 9438 9034 9472 9067
rect 9530 9034 9564 9068
rect 9622 9034 9656 9068
rect 9714 9034 9748 9068
rect 9806 9034 9840 9068
rect 9898 9034 9932 9068
rect 9990 9034 10024 9068
rect 10082 9067 10116 9068
rect 10082 9034 10116 9067
rect 10174 9034 10208 9068
rect 10266 9034 10300 9068
rect 10358 9034 10392 9068
rect 10450 9034 10484 9068
rect 10542 9034 10576 9068
rect 10634 9034 10668 9068
rect 10726 9034 10760 9068
rect 10818 9034 10852 9068
rect 10910 9067 10944 9068
rect 10910 9034 10944 9067
rect 11002 9034 11036 9068
rect 11094 9034 11128 9068
rect 11186 9034 11220 9068
rect 11278 9034 11312 9068
rect 11370 9034 11404 9068
rect 11462 9034 11496 9068
rect 11554 9034 11588 9068
rect 11646 9067 11680 9068
rect 11646 9034 11680 9067
rect 3923 8883 3957 8943
rect 4013 8883 4047 8943
rect 4655 8883 4689 8943
rect 4762 8883 4796 8943
rect 4865 8883 4899 8943
rect 5867 8883 5901 8943
rect 5973 8883 6007 8943
rect 6077 8883 6111 8943
rect 7205 8883 7239 8943
rect 7313 8883 7347 8943
rect 7415 8883 7449 8943
rect 8060 8883 8094 8943
rect 8149 8883 8183 8943
rect 8713 8882 8747 8942
rect 8801 8882 8835 8942
rect 8897 8882 8931 8942
rect 8993 8882 9027 8942
rect 8642 8796 8676 8830
rect 8849 8798 8883 8832
rect 9136 8802 9141 8833
rect 9141 8802 9170 8833
rect 9136 8799 9170 8802
rect 9236 8794 9270 8828
rect 2415 8655 2449 8689
rect 2507 8684 2514 8689
rect 2514 8684 2541 8689
rect 2599 8684 2632 8689
rect 2632 8684 2633 8689
rect 2507 8655 2541 8684
rect 2599 8655 2633 8684
rect 2691 8655 2725 8689
rect 2783 8655 2817 8689
rect 3570 8685 3604 8745
rect 3658 8682 3692 8742
rect 4302 8682 4336 8742
rect 4407 8682 4441 8742
rect 4516 8682 4550 8742
rect 5514 8682 5548 8742
rect 5618 8682 5652 8742
rect 5728 8682 5762 8742
rect 6726 8682 6760 8742
rect 6831 8682 6865 8742
rect 6940 8682 6974 8742
rect 7938 8682 7972 8742
rect 8045 8682 8079 8742
rect 8152 8682 8186 8742
rect 8713 8679 8747 8739
rect 8801 8679 8835 8739
rect 8897 8679 8931 8739
rect 8993 8679 9027 8739
rect 2462 8423 2466 8453
rect 2466 8423 2496 8453
rect 2462 8419 2496 8423
rect 2543 8255 2546 8288
rect 2546 8255 2577 8288
rect 2543 8254 2577 8255
rect 3173 8587 3207 8621
rect 3614 8592 3648 8626
rect 4346 8589 4380 8623
rect 4472 8589 4506 8623
rect 5558 8589 5592 8623
rect 5684 8589 5718 8623
rect 6770 8589 6804 8623
rect 6896 8589 6930 8623
rect 7982 8589 8016 8623
rect 8108 8589 8142 8623
rect 2913 8512 2947 8546
rect 8713 8541 8747 8601
rect 3172 8494 3206 8528
rect 8801 8541 8835 8601
rect 9343 8602 9352 8635
rect 9352 8602 9377 8635
rect 9343 8601 9377 8602
rect 9789 8798 9821 8827
rect 9821 8798 9823 8827
rect 9789 8793 9823 8798
rect 9897 8728 9931 8762
rect 10173 8872 10207 8898
rect 10173 8864 10198 8872
rect 10198 8864 10207 8872
rect 10449 8796 10483 8830
rect 10909 8872 10943 8898
rect 10909 8864 10941 8872
rect 10941 8864 10943 8872
rect 10541 8728 10575 8762
rect 10449 8686 10462 8694
rect 10462 8686 10483 8694
rect 10449 8660 10483 8686
rect 12150 9018 12184 9052
rect 12222 9018 12256 9052
rect 12295 9018 12329 9052
rect 12367 9018 12401 9052
rect 12440 9017 12474 9051
rect 12512 9017 12546 9051
rect 12678 9021 12712 9055
rect 12770 9021 12804 9055
rect 12862 9021 12896 9055
rect 12954 9021 12988 9055
rect 13046 9021 13080 9055
rect 13138 9021 13172 9055
rect 11097 8882 11131 8898
rect 11097 8864 11113 8882
rect 11113 8864 11131 8882
rect 11185 8660 11219 8694
rect 11461 8864 11495 8898
rect 11833 8884 11867 8944
rect 11929 8884 11963 8944
rect 12025 8884 12059 8944
rect 12121 8884 12155 8944
rect 12233 8872 12267 8932
rect 12321 8872 12355 8932
rect 12434 8871 12468 8931
rect 12522 8871 12556 8931
rect 13456 9008 13490 9068
rect 13544 9008 13578 9068
rect 19194 9055 19228 9115
rect 19354 9055 19388 9115
rect 14152 8981 14186 9015
rect 14886 8981 14920 9015
rect 15008 8981 15042 9015
rect 16224 8981 16258 9015
rect 16346 8981 16380 9015
rect 17436 8981 17470 9015
rect 17558 8981 17592 9015
rect 18290 8981 18324 9015
rect 20165 9008 20199 9068
rect 19274 8971 19308 9005
rect 20253 9008 20287 9068
rect 25903 9055 25937 9115
rect 26063 9055 26097 9115
rect 20861 8981 20895 9015
rect 21595 8981 21629 9015
rect 21717 8981 21751 9015
rect 22933 8981 22967 9015
rect 23055 8981 23089 9015
rect 24145 8981 24179 9015
rect 24267 8981 24301 9015
rect 24999 8981 25033 9015
rect 25983 8971 26017 9005
rect 12073 8787 12107 8821
rect 12277 8788 12311 8822
rect 12478 8787 12512 8821
rect 12687 8789 12721 8816
rect 12687 8782 12721 8789
rect 11652 8728 11686 8762
rect 11553 8660 11587 8694
rect 9090 8490 9124 8524
rect 9182 8490 9216 8524
rect 9274 8490 9308 8524
rect 9346 8490 9380 8524
rect 9438 8490 9472 8524
rect 9530 8490 9564 8524
rect 9622 8490 9656 8524
rect 9714 8490 9748 8524
rect 9806 8490 9840 8524
rect 9898 8490 9932 8524
rect 9990 8490 10024 8524
rect 10082 8490 10116 8524
rect 10174 8490 10208 8524
rect 10266 8490 10300 8524
rect 10358 8490 10392 8524
rect 10450 8490 10484 8524
rect 10542 8490 10576 8524
rect 10634 8490 10668 8524
rect 10726 8490 10760 8524
rect 10818 8490 10852 8524
rect 10910 8490 10944 8524
rect 11002 8490 11036 8524
rect 11094 8490 11128 8524
rect 11186 8490 11220 8524
rect 11278 8490 11312 8524
rect 2736 8423 2766 8454
rect 2766 8423 2770 8454
rect 2736 8420 2770 8423
rect 2875 8419 2909 8453
rect 11370 8490 11404 8524
rect 11462 8490 11496 8524
rect 11554 8490 11588 8524
rect 11646 8490 11680 8524
rect 11833 8500 11867 8728
rect 11929 8500 11963 8728
rect 2652 8323 2686 8343
rect 2652 8309 2686 8323
rect 2972 8349 3006 8383
rect 12025 8500 12059 8728
rect 12121 8500 12155 8728
rect 12233 8501 12267 8729
rect 12321 8501 12355 8729
rect 12434 8472 12468 8728
rect 13264 8870 13298 8930
rect 13360 8870 13394 8930
rect 13456 8870 13490 8930
rect 13544 8870 13578 8930
rect 14108 8871 14142 8931
rect 14197 8871 14231 8931
rect 14842 8871 14876 8931
rect 14944 8871 14978 8931
rect 15052 8871 15086 8931
rect 16180 8871 16214 8931
rect 16284 8871 16318 8931
rect 16390 8871 16424 8931
rect 17392 8871 17426 8931
rect 17495 8871 17529 8931
rect 17602 8871 17636 8931
rect 18244 8871 18278 8931
rect 18334 8871 18368 8931
rect 19973 8870 20007 8930
rect 20069 8870 20103 8930
rect 20165 8870 20199 8930
rect 20253 8870 20287 8930
rect 20817 8871 20851 8931
rect 20906 8871 20940 8931
rect 21551 8871 21585 8931
rect 21653 8871 21687 8931
rect 21761 8871 21795 8931
rect 22889 8871 22923 8931
rect 22993 8871 23027 8931
rect 23099 8871 23133 8931
rect 24101 8871 24135 8931
rect 24204 8871 24238 8931
rect 24311 8871 24345 8931
rect 24953 8871 24987 8931
rect 25043 8871 25077 8931
rect 13085 8789 13087 8820
rect 13087 8789 13119 8820
rect 13085 8786 13119 8789
rect 13408 8786 13442 8820
rect 13615 8784 13649 8818
rect 20117 8786 20151 8820
rect 20324 8784 20358 8818
rect 12522 8472 12556 8728
rect 12767 8621 12768 8630
rect 12768 8621 12801 8630
rect 12767 8596 12801 8621
rect 13264 8667 13298 8727
rect 13360 8667 13394 8727
rect 13456 8667 13490 8727
rect 13544 8667 13578 8727
rect 14105 8670 14139 8730
rect 14212 8670 14246 8730
rect 14319 8670 14353 8730
rect 15317 8670 15351 8730
rect 15426 8670 15460 8730
rect 15531 8670 15565 8730
rect 16529 8670 16563 8730
rect 16639 8670 16673 8730
rect 16743 8670 16777 8730
rect 17741 8670 17775 8730
rect 17850 8670 17884 8730
rect 17955 8670 17989 8730
rect 18599 8670 18633 8730
rect 18687 8673 18721 8733
rect 19474 8643 19508 8677
rect 19566 8643 19600 8677
rect 19658 8672 19659 8677
rect 19659 8672 19692 8677
rect 19750 8672 19777 8677
rect 19777 8672 19784 8677
rect 19658 8643 19692 8672
rect 19750 8643 19784 8672
rect 19842 8643 19876 8677
rect 19973 8667 20007 8727
rect 20069 8667 20103 8727
rect 20165 8667 20199 8727
rect 20253 8667 20287 8727
rect 20814 8670 20848 8730
rect 20921 8670 20955 8730
rect 21028 8670 21062 8730
rect 22026 8670 22060 8730
rect 22135 8670 22169 8730
rect 22240 8670 22274 8730
rect 23238 8670 23272 8730
rect 23348 8670 23382 8730
rect 23452 8670 23486 8730
rect 24450 8670 24484 8730
rect 24559 8670 24593 8730
rect 24664 8670 24698 8730
rect 25308 8670 25342 8730
rect 25396 8673 25430 8733
rect 26183 8643 26217 8677
rect 26275 8643 26309 8677
rect 26367 8672 26368 8677
rect 26368 8672 26401 8677
rect 26459 8672 26486 8677
rect 26486 8672 26493 8677
rect 26367 8643 26401 8672
rect 26459 8643 26493 8672
rect 26551 8643 26585 8677
rect 13456 8529 13490 8589
rect 13544 8529 13578 8589
rect 14149 8577 14183 8611
rect 14275 8577 14309 8611
rect 15361 8577 15395 8611
rect 15487 8577 15521 8611
rect 16573 8577 16607 8611
rect 16699 8577 16733 8611
rect 17785 8577 17819 8611
rect 17911 8577 17945 8611
rect 18643 8580 18677 8614
rect 19084 8575 19118 8609
rect 12678 8477 12712 8511
rect 12770 8477 12804 8511
rect 12862 8477 12896 8511
rect 12954 8477 12988 8511
rect 13046 8477 13080 8511
rect 13138 8477 13172 8511
rect 19085 8482 19119 8516
rect 19344 8500 19378 8534
rect 12200 8393 12234 8427
rect 12274 8393 12308 8427
rect 19382 8407 19416 8441
rect 19521 8411 19525 8442
rect 19525 8411 19555 8442
rect 19521 8408 19555 8411
rect 10083 8315 10117 8349
rect 10175 8315 10209 8349
rect 10267 8315 10301 8349
rect 10359 8315 10393 8349
rect 10451 8315 10485 8349
rect 10543 8315 10577 8349
rect 10635 8315 10669 8349
rect 10727 8315 10761 8349
rect 10819 8315 10853 8349
rect 10910 8315 10944 8349
rect 11002 8315 11036 8349
rect 11094 8315 11128 8349
rect 11186 8315 11220 8349
rect 11278 8315 11312 8349
rect 11370 8315 11404 8349
rect 11462 8315 11496 8349
rect 11554 8315 11588 8349
rect 11646 8315 11680 8349
rect 2928 8230 2962 8290
rect 3016 8230 3050 8290
rect 8893 8187 8927 8221
rect 2415 8111 2449 8145
rect 2507 8111 2541 8145
rect 2599 8116 2633 8145
rect 2599 8111 2624 8116
rect 2624 8111 2633 8116
rect 2691 8111 2725 8145
rect 2783 8111 2817 8145
rect 2928 8092 2962 8152
rect 3016 8092 3050 8152
rect 8894 8030 8928 8064
rect 2928 7954 2962 8014
rect 3016 7954 3050 8014
rect 2928 7816 2962 7876
rect 3016 7816 3050 7876
rect 8894 7860 8928 7894
rect 10078 7900 10112 7905
rect 10078 7871 10089 7900
rect 10089 7871 10112 7900
rect 10465 7874 10499 7908
rect 10715 8080 10747 8112
rect 10747 8080 10749 8112
rect 10715 8078 10749 8080
rect 11286 8008 11320 8042
rect 10910 7900 10944 7908
rect 10910 7874 10916 7900
rect 10916 7874 10944 7900
rect 11538 8080 11540 8112
rect 11540 8080 11572 8112
rect 11538 8078 11572 8080
rect 11833 8096 11867 8324
rect 11929 8096 11963 8324
rect 12025 8096 12059 8324
rect 12121 8096 12155 8324
rect 12233 8095 12267 8323
rect 12321 8095 12355 8323
rect 12452 8337 12486 8369
rect 12452 8335 12486 8337
rect 12532 8336 12565 8370
rect 12565 8336 12566 8370
rect 19285 8337 19319 8371
rect 12746 8190 12780 8224
rect 13364 8175 13398 8209
rect 19241 8218 19275 8278
rect 19329 8218 19363 8278
rect 12702 8080 12736 8140
rect 12790 8080 12824 8140
rect 19241 8080 19275 8140
rect 19329 8080 19363 8140
rect 19605 8311 19639 8331
rect 19605 8297 19639 8311
rect 20165 8529 20199 8589
rect 20253 8529 20287 8589
rect 20858 8577 20892 8611
rect 20984 8577 21018 8611
rect 22070 8577 22104 8611
rect 22196 8577 22230 8611
rect 23282 8577 23316 8611
rect 23408 8577 23442 8611
rect 24494 8577 24528 8611
rect 24620 8577 24654 8611
rect 25352 8580 25386 8614
rect 25793 8575 25827 8609
rect 25794 8482 25828 8516
rect 26053 8500 26087 8534
rect 19795 8411 19825 8441
rect 19825 8411 19829 8441
rect 19795 8407 19829 8411
rect 26091 8407 26125 8441
rect 26230 8411 26234 8442
rect 26234 8411 26264 8442
rect 26230 8408 26264 8411
rect 19714 8243 19745 8276
rect 19745 8243 19748 8276
rect 19714 8242 19748 8243
rect 25994 8337 26028 8371
rect 20073 8175 20107 8209
rect 25950 8218 25984 8278
rect 26038 8218 26072 8278
rect 19474 8099 19508 8133
rect 19566 8099 19600 8133
rect 19658 8104 19692 8133
rect 19658 8099 19667 8104
rect 19667 8099 19692 8104
rect 19750 8099 19784 8133
rect 19842 8099 19876 8133
rect 25950 8080 25984 8140
rect 12073 8003 12107 8037
rect 12277 8002 12311 8036
rect 13363 8018 13397 8052
rect 26038 8080 26072 8140
rect 26314 8311 26348 8331
rect 26314 8297 26348 8311
rect 26504 8411 26534 8441
rect 26534 8411 26538 8441
rect 26504 8407 26538 8411
rect 26423 8243 26454 8276
rect 26454 8243 26457 8276
rect 26423 8242 26457 8243
rect 26183 8099 26217 8133
rect 26275 8099 26309 8133
rect 26367 8104 26401 8133
rect 26367 8099 26376 8104
rect 26376 8099 26401 8104
rect 26459 8099 26493 8133
rect 26551 8099 26585 8133
rect 20072 8018 20106 8052
rect 11833 7880 11867 7940
rect 11929 7880 11963 7940
rect 12025 7880 12059 7940
rect 12121 7880 12155 7940
rect 12233 7892 12267 7952
rect 12321 7892 12355 7952
rect 2928 7678 2962 7738
rect 3016 7678 3050 7738
rect 8893 7708 8927 7742
rect 10083 7771 10117 7805
rect 10175 7771 10209 7805
rect 10267 7771 10301 7805
rect 10359 7771 10393 7805
rect 10451 7771 10485 7805
rect 10543 7771 10577 7805
rect 10635 7771 10669 7805
rect 10727 7771 10761 7805
rect 10819 7771 10853 7805
rect 10910 7771 10944 7805
rect 11002 7771 11036 7805
rect 11094 7771 11128 7805
rect 11186 7771 11220 7805
rect 11278 7771 11312 7805
rect 11370 7771 11404 7805
rect 11462 7771 11496 7805
rect 11554 7771 11588 7805
rect 11646 7771 11680 7805
rect 11942 7728 11976 7762
rect 12014 7728 12048 7762
rect 12087 7728 12121 7762
rect 12159 7728 12193 7762
rect 12232 7727 12266 7761
rect 12304 7727 12338 7761
rect 2928 7540 2962 7600
rect 11941 7656 11975 7690
rect 12013 7656 12047 7690
rect 12086 7656 12120 7690
rect 12158 7656 12192 7690
rect 12231 7655 12265 7689
rect 12303 7655 12337 7689
rect 3016 7540 3050 7600
rect 8888 7564 8922 7598
rect 3176 7516 3208 7550
rect 3208 7516 3210 7550
rect 3256 7516 3288 7550
rect 3288 7516 3290 7550
rect 3336 7516 3368 7550
rect 3368 7516 3370 7550
rect 3416 7516 3448 7550
rect 3448 7516 3450 7550
rect 3496 7516 3528 7550
rect 3528 7516 3530 7550
rect 3576 7516 3608 7550
rect 3608 7516 3610 7550
rect 3908 7513 3940 7547
rect 3940 7513 3942 7547
rect 3988 7513 4020 7547
rect 4020 7513 4022 7547
rect 4068 7513 4100 7547
rect 4100 7513 4102 7547
rect 4148 7513 4180 7547
rect 4180 7513 4182 7547
rect 4228 7513 4260 7547
rect 4260 7513 4262 7547
rect 4308 7513 4340 7547
rect 4340 7513 4342 7547
rect 4510 7513 4512 7547
rect 4512 7513 4544 7547
rect 4590 7513 4592 7547
rect 4592 7513 4624 7547
rect 4670 7513 4672 7547
rect 4672 7513 4704 7547
rect 4750 7513 4752 7547
rect 4752 7513 4784 7547
rect 4830 7513 4832 7547
rect 4832 7513 4864 7547
rect 4910 7513 4912 7547
rect 4912 7513 4944 7547
rect 5120 7513 5152 7547
rect 5152 7513 5154 7547
rect 5200 7513 5232 7547
rect 5232 7513 5234 7547
rect 5280 7513 5312 7547
rect 5312 7513 5314 7547
rect 5360 7513 5392 7547
rect 5392 7513 5394 7547
rect 5440 7513 5472 7547
rect 5472 7513 5474 7547
rect 5520 7513 5552 7547
rect 5552 7513 5554 7547
rect 5722 7513 5724 7547
rect 5724 7513 5756 7547
rect 5802 7513 5804 7547
rect 5804 7513 5836 7547
rect 5882 7513 5884 7547
rect 5884 7513 5916 7547
rect 5962 7513 5964 7547
rect 5964 7513 5996 7547
rect 6042 7513 6044 7547
rect 6044 7513 6076 7547
rect 6122 7513 6124 7547
rect 6124 7513 6156 7547
rect 6332 7513 6364 7547
rect 6364 7513 6366 7547
rect 6412 7513 6444 7547
rect 6444 7513 6446 7547
rect 6492 7513 6524 7547
rect 6524 7513 6526 7547
rect 6572 7513 6604 7547
rect 6604 7513 6606 7547
rect 6652 7513 6684 7547
rect 6684 7513 6686 7547
rect 6732 7513 6764 7547
rect 6764 7513 6766 7547
rect 6934 7513 6936 7547
rect 6936 7513 6968 7547
rect 7014 7513 7016 7547
rect 7016 7513 7048 7547
rect 7094 7513 7096 7547
rect 7096 7513 7128 7547
rect 7174 7513 7176 7547
rect 7176 7513 7208 7547
rect 7254 7513 7256 7547
rect 7256 7513 7288 7547
rect 7334 7513 7336 7547
rect 7336 7513 7368 7547
rect 7544 7513 7576 7547
rect 7576 7513 7578 7547
rect 7624 7513 7656 7547
rect 7656 7513 7658 7547
rect 7704 7513 7736 7547
rect 7736 7513 7738 7547
rect 7784 7513 7816 7547
rect 7816 7513 7818 7547
rect 7864 7513 7896 7547
rect 7896 7513 7898 7547
rect 7944 7513 7976 7547
rect 7976 7513 7978 7547
rect 8146 7513 8148 7547
rect 8148 7513 8180 7547
rect 8226 7513 8228 7547
rect 8228 7513 8260 7547
rect 8306 7513 8308 7547
rect 8308 7513 8340 7547
rect 8386 7513 8388 7547
rect 8388 7513 8420 7547
rect 8466 7513 8468 7547
rect 8468 7513 8500 7547
rect 8546 7513 8548 7547
rect 8548 7513 8580 7547
rect 11941 7584 11975 7618
rect 12013 7584 12047 7618
rect 12086 7584 12120 7618
rect 12158 7584 12192 7618
rect 12231 7583 12265 7617
rect 12303 7583 12337 7617
rect 12702 7596 12736 7952
rect 12790 7596 12824 7952
rect 19241 7942 19275 8002
rect 19329 7942 19363 8002
rect 19650 7946 19684 7980
rect 25950 7942 25984 8002
rect 26038 7942 26072 8002
rect 12947 7884 12981 7918
rect 13363 7848 13397 7882
rect 19241 7804 19275 7864
rect 19329 7804 19363 7864
rect 20072 7848 20106 7882
rect 25950 7804 25984 7864
rect 26038 7804 26072 7864
rect 19650 7750 19684 7784
rect 12939 7664 12973 7698
rect 13364 7696 13398 7730
rect 19241 7666 19275 7726
rect 11940 7512 11974 7546
rect 12012 7512 12046 7546
rect 12085 7512 12119 7546
rect 12157 7512 12191 7546
rect 12230 7511 12264 7545
rect 12302 7511 12336 7545
rect 13369 7552 13403 7586
rect 19329 7666 19363 7726
rect 20073 7696 20107 7730
rect 25950 7666 25984 7726
rect 12746 7503 12780 7537
rect 13711 7501 13743 7535
rect 13743 7501 13745 7535
rect 13791 7501 13823 7535
rect 13823 7501 13825 7535
rect 13871 7501 13903 7535
rect 13903 7501 13905 7535
rect 13951 7501 13983 7535
rect 13983 7501 13985 7535
rect 14031 7501 14063 7535
rect 14063 7501 14065 7535
rect 14111 7501 14143 7535
rect 14143 7501 14145 7535
rect 14313 7501 14315 7535
rect 14315 7501 14347 7535
rect 14393 7501 14395 7535
rect 14395 7501 14427 7535
rect 14473 7501 14475 7535
rect 14475 7501 14507 7535
rect 14553 7501 14555 7535
rect 14555 7501 14587 7535
rect 14633 7501 14635 7535
rect 14635 7501 14667 7535
rect 14713 7501 14715 7535
rect 14715 7501 14747 7535
rect 14923 7501 14955 7535
rect 14955 7501 14957 7535
rect 15003 7501 15035 7535
rect 15035 7501 15037 7535
rect 15083 7501 15115 7535
rect 15115 7501 15117 7535
rect 15163 7501 15195 7535
rect 15195 7501 15197 7535
rect 15243 7501 15275 7535
rect 15275 7501 15277 7535
rect 15323 7501 15355 7535
rect 15355 7501 15357 7535
rect 15525 7501 15527 7535
rect 15527 7501 15559 7535
rect 15605 7501 15607 7535
rect 15607 7501 15639 7535
rect 15685 7501 15687 7535
rect 15687 7501 15719 7535
rect 15765 7501 15767 7535
rect 15767 7501 15799 7535
rect 15845 7501 15847 7535
rect 15847 7501 15879 7535
rect 15925 7501 15927 7535
rect 15927 7501 15959 7535
rect 16135 7501 16167 7535
rect 16167 7501 16169 7535
rect 16215 7501 16247 7535
rect 16247 7501 16249 7535
rect 16295 7501 16327 7535
rect 16327 7501 16329 7535
rect 16375 7501 16407 7535
rect 16407 7501 16409 7535
rect 16455 7501 16487 7535
rect 16487 7501 16489 7535
rect 16535 7501 16567 7535
rect 16567 7501 16569 7535
rect 16737 7501 16739 7535
rect 16739 7501 16771 7535
rect 16817 7501 16819 7535
rect 16819 7501 16851 7535
rect 16897 7501 16899 7535
rect 16899 7501 16931 7535
rect 16977 7501 16979 7535
rect 16979 7501 17011 7535
rect 17057 7501 17059 7535
rect 17059 7501 17091 7535
rect 17137 7501 17139 7535
rect 17139 7501 17171 7535
rect 17347 7501 17379 7535
rect 17379 7501 17381 7535
rect 17427 7501 17459 7535
rect 17459 7501 17461 7535
rect 17507 7501 17539 7535
rect 17539 7501 17541 7535
rect 17587 7501 17619 7535
rect 17619 7501 17621 7535
rect 17667 7501 17699 7535
rect 17699 7501 17701 7535
rect 17747 7501 17779 7535
rect 17779 7501 17781 7535
rect 17949 7501 17951 7535
rect 17951 7501 17983 7535
rect 18029 7501 18031 7535
rect 18031 7501 18063 7535
rect 18109 7501 18111 7535
rect 18111 7501 18143 7535
rect 18189 7501 18191 7535
rect 18191 7501 18223 7535
rect 18269 7501 18271 7535
rect 18271 7501 18303 7535
rect 18349 7501 18351 7535
rect 18351 7501 18383 7535
rect 18681 7504 18683 7538
rect 18683 7504 18715 7538
rect 18761 7504 18763 7538
rect 18763 7504 18795 7538
rect 18841 7504 18843 7538
rect 18843 7504 18875 7538
rect 18921 7504 18923 7538
rect 18923 7504 18955 7538
rect 19001 7504 19003 7538
rect 19003 7504 19035 7538
rect 19081 7504 19083 7538
rect 19083 7504 19115 7538
rect 19241 7528 19275 7588
rect 19329 7528 19363 7588
rect 19650 7575 19684 7609
rect 20078 7552 20112 7586
rect 26038 7666 26072 7726
rect 20420 7501 20452 7535
rect 20452 7501 20454 7535
rect 20500 7501 20532 7535
rect 20532 7501 20534 7535
rect 20580 7501 20612 7535
rect 20612 7501 20614 7535
rect 20660 7501 20692 7535
rect 20692 7501 20694 7535
rect 20740 7501 20772 7535
rect 20772 7501 20774 7535
rect 20820 7501 20852 7535
rect 20852 7501 20854 7535
rect 21022 7501 21024 7535
rect 21024 7501 21056 7535
rect 21102 7501 21104 7535
rect 21104 7501 21136 7535
rect 21182 7501 21184 7535
rect 21184 7501 21216 7535
rect 21262 7501 21264 7535
rect 21264 7501 21296 7535
rect 21342 7501 21344 7535
rect 21344 7501 21376 7535
rect 21422 7501 21424 7535
rect 21424 7501 21456 7535
rect 21632 7501 21664 7535
rect 21664 7501 21666 7535
rect 21712 7501 21744 7535
rect 21744 7501 21746 7535
rect 21792 7501 21824 7535
rect 21824 7501 21826 7535
rect 21872 7501 21904 7535
rect 21904 7501 21906 7535
rect 21952 7501 21984 7535
rect 21984 7501 21986 7535
rect 22032 7501 22064 7535
rect 22064 7501 22066 7535
rect 22234 7501 22236 7535
rect 22236 7501 22268 7535
rect 22314 7501 22316 7535
rect 22316 7501 22348 7535
rect 22394 7501 22396 7535
rect 22396 7501 22428 7535
rect 22474 7501 22476 7535
rect 22476 7501 22508 7535
rect 22554 7501 22556 7535
rect 22556 7501 22588 7535
rect 22634 7501 22636 7535
rect 22636 7501 22668 7535
rect 22844 7501 22876 7535
rect 22876 7501 22878 7535
rect 22924 7501 22956 7535
rect 22956 7501 22958 7535
rect 23004 7501 23036 7535
rect 23036 7501 23038 7535
rect 23084 7501 23116 7535
rect 23116 7501 23118 7535
rect 23164 7501 23196 7535
rect 23196 7501 23198 7535
rect 23244 7501 23276 7535
rect 23276 7501 23278 7535
rect 23446 7501 23448 7535
rect 23448 7501 23480 7535
rect 23526 7501 23528 7535
rect 23528 7501 23560 7535
rect 23606 7501 23608 7535
rect 23608 7501 23640 7535
rect 23686 7501 23688 7535
rect 23688 7501 23720 7535
rect 23766 7501 23768 7535
rect 23768 7501 23800 7535
rect 23846 7501 23848 7535
rect 23848 7501 23880 7535
rect 24056 7501 24088 7535
rect 24088 7501 24090 7535
rect 24136 7501 24168 7535
rect 24168 7501 24170 7535
rect 24216 7501 24248 7535
rect 24248 7501 24250 7535
rect 24296 7501 24328 7535
rect 24328 7501 24330 7535
rect 24376 7501 24408 7535
rect 24408 7501 24410 7535
rect 24456 7501 24488 7535
rect 24488 7501 24490 7535
rect 24658 7501 24660 7535
rect 24660 7501 24692 7535
rect 24738 7501 24740 7535
rect 24740 7501 24772 7535
rect 24818 7501 24820 7535
rect 24820 7501 24852 7535
rect 24898 7501 24900 7535
rect 24900 7501 24932 7535
rect 24978 7501 24980 7535
rect 24980 7501 25012 7535
rect 25058 7501 25060 7535
rect 25060 7501 25092 7535
rect 25390 7504 25392 7538
rect 25392 7504 25424 7538
rect 25470 7504 25472 7538
rect 25472 7504 25504 7538
rect 25550 7504 25552 7538
rect 25552 7504 25584 7538
rect 25630 7504 25632 7538
rect 25632 7504 25664 7538
rect 25710 7504 25712 7538
rect 25712 7504 25744 7538
rect 25790 7504 25792 7538
rect 25792 7504 25824 7538
rect 25950 7528 25984 7588
rect 26038 7528 26072 7588
rect 24541 7224 24575 7284
rect 24629 7224 24663 7284
rect 24789 7274 24821 7308
rect 24821 7274 24823 7308
rect 24869 7274 24901 7308
rect 24901 7274 24903 7308
rect 24949 7274 24981 7308
rect 24981 7274 24983 7308
rect 25029 7274 25061 7308
rect 25061 7274 25063 7308
rect 25109 7274 25141 7308
rect 25141 7274 25143 7308
rect 25189 7274 25221 7308
rect 25221 7274 25223 7308
rect 25521 7277 25553 7311
rect 25553 7277 25555 7311
rect 25601 7277 25633 7311
rect 25633 7277 25635 7311
rect 25681 7277 25713 7311
rect 25713 7277 25715 7311
rect 25761 7277 25793 7311
rect 25793 7277 25795 7311
rect 25841 7277 25873 7311
rect 25873 7277 25875 7311
rect 25921 7277 25953 7311
rect 25953 7277 25955 7311
rect 26123 7277 26125 7311
rect 26125 7277 26157 7311
rect 26203 7277 26205 7311
rect 26205 7277 26237 7311
rect 26283 7277 26285 7311
rect 26285 7277 26317 7311
rect 26363 7277 26365 7311
rect 26365 7277 26397 7311
rect 26443 7277 26445 7311
rect 26445 7277 26477 7311
rect 26523 7277 26525 7311
rect 26525 7277 26557 7311
rect 26733 7277 26765 7311
rect 26765 7277 26767 7311
rect 26813 7277 26845 7311
rect 26845 7277 26847 7311
rect 26893 7277 26925 7311
rect 26925 7277 26927 7311
rect 26973 7277 27005 7311
rect 27005 7277 27007 7311
rect 27053 7277 27085 7311
rect 27085 7277 27087 7311
rect 27133 7277 27165 7311
rect 27165 7277 27167 7311
rect 27335 7277 27337 7311
rect 27337 7277 27369 7311
rect 27415 7277 27417 7311
rect 27417 7277 27449 7311
rect 27495 7277 27497 7311
rect 27497 7277 27529 7311
rect 27575 7277 27577 7311
rect 27577 7277 27609 7311
rect 27655 7277 27657 7311
rect 27657 7277 27689 7311
rect 27735 7277 27737 7311
rect 27737 7277 27769 7311
rect 27945 7277 27977 7311
rect 27977 7277 27979 7311
rect 28025 7277 28057 7311
rect 28057 7277 28059 7311
rect 28105 7277 28137 7311
rect 28137 7277 28139 7311
rect 28185 7277 28217 7311
rect 28217 7277 28219 7311
rect 28265 7277 28297 7311
rect 28297 7277 28299 7311
rect 28345 7277 28377 7311
rect 28377 7277 28379 7311
rect 28547 7277 28549 7311
rect 28549 7277 28581 7311
rect 28627 7277 28629 7311
rect 28629 7277 28661 7311
rect 28707 7277 28709 7311
rect 28709 7277 28741 7311
rect 28787 7277 28789 7311
rect 28789 7277 28821 7311
rect 28867 7277 28869 7311
rect 28869 7277 28901 7311
rect 28947 7277 28949 7311
rect 28949 7277 28981 7311
rect 29157 7277 29189 7311
rect 29189 7277 29191 7311
rect 29237 7277 29269 7311
rect 29269 7277 29271 7311
rect 29317 7277 29349 7311
rect 29349 7277 29351 7311
rect 29397 7277 29429 7311
rect 29429 7277 29431 7311
rect 29477 7277 29509 7311
rect 29509 7277 29511 7311
rect 29557 7277 29589 7311
rect 29589 7277 29591 7311
rect 29759 7277 29761 7311
rect 29761 7277 29793 7311
rect 29839 7277 29841 7311
rect 29841 7277 29873 7311
rect 29919 7277 29921 7311
rect 29921 7277 29953 7311
rect 29999 7277 30001 7311
rect 30001 7277 30033 7311
rect 30079 7277 30081 7311
rect 30081 7277 30113 7311
rect 30159 7277 30161 7311
rect 30161 7277 30193 7311
rect 11527 7084 11561 7094
rect 11527 7060 11561 7084
rect 11619 7084 11653 7094
rect 11619 7060 11653 7084
rect 11711 7084 11745 7094
rect 11711 7060 11745 7084
rect 11803 7084 11837 7094
rect 11803 7060 11837 7084
rect 11895 7084 11929 7094
rect 11895 7060 11929 7084
rect 11987 7084 12021 7094
rect 11987 7060 12021 7084
rect 12079 7084 12113 7094
rect 12079 7060 12113 7084
rect 12171 7060 12205 7094
rect 12263 7060 12297 7094
rect 12787 7084 12821 7094
rect 12787 7060 12821 7084
rect 12879 7084 12913 7094
rect 12879 7060 12913 7084
rect 12971 7084 13005 7094
rect 12971 7060 13005 7084
rect 13063 7084 13097 7094
rect 13063 7060 13097 7084
rect 13155 7084 13189 7094
rect 13155 7060 13189 7084
rect 13247 7084 13281 7094
rect 13247 7060 13281 7084
rect 13339 7084 13373 7094
rect 13339 7060 13373 7084
rect 13431 7084 13465 7094
rect 13431 7060 13465 7084
rect 13523 7084 13557 7094
rect 13523 7060 13557 7084
rect 13615 7084 13649 7094
rect 13615 7060 13649 7084
rect 13707 7084 13741 7094
rect 13707 7060 13741 7084
rect 13799 7084 13833 7094
rect 13799 7060 13833 7084
rect 13891 7084 13925 7094
rect 13891 7060 13925 7084
rect 13983 7084 14017 7094
rect 13983 7060 14017 7084
rect 14075 7084 14109 7094
rect 14075 7060 14109 7084
rect 14167 7084 14201 7094
rect 14167 7060 14201 7084
rect 14259 7084 14293 7094
rect 14259 7060 14293 7084
rect 14351 7084 14385 7094
rect 14351 7060 14385 7084
rect 14443 7084 14477 7094
rect 14443 7060 14477 7084
rect 14535 7084 14569 7094
rect 14535 7060 14569 7084
rect 24541 7086 24575 7146
rect 30501 7226 30535 7260
rect 24629 7086 24663 7146
rect 30506 7082 30540 7116
rect 11531 6782 11565 6789
rect 11531 6755 11535 6782
rect 11535 6755 11565 6782
rect 13246 6958 13280 6992
rect 13430 6898 13464 6924
rect 13430 6890 13440 6898
rect 13440 6890 13464 6898
rect 13338 6822 13372 6856
rect 12175 6755 12209 6789
rect 12873 6752 12907 6786
rect 13706 6958 13740 6992
rect 13241 6615 13275 6649
rect 13601 6762 13608 6790
rect 13608 6762 13635 6790
rect 13601 6756 13635 6762
rect 13890 6958 13924 6992
rect 14166 6958 14200 6992
rect 24541 6948 24575 7008
rect 24629 6948 24663 7008
rect 14258 6890 14292 6924
rect 30507 6930 30541 6964
rect 13982 6702 14003 6719
rect 14003 6702 14016 6719
rect 13982 6685 14016 6702
rect 14076 6702 14099 6719
rect 14099 6702 14110 6719
rect 14076 6685 14110 6702
rect 14350 6840 14384 6856
rect 14350 6822 14353 6840
rect 14353 6822 14384 6840
rect 14534 6822 14568 6856
rect 24541 6810 24575 6870
rect 24629 6810 24663 6870
rect 30507 6760 30541 6794
rect 24028 6679 24062 6713
rect 24120 6679 24154 6713
rect 24212 6708 24237 6713
rect 24237 6708 24246 6713
rect 24212 6679 24246 6708
rect 24304 6679 24338 6713
rect 24396 6679 24430 6713
rect 14354 6624 14388 6658
rect 11527 6526 11561 6550
rect 11527 6516 11561 6526
rect 11619 6526 11653 6550
rect 11619 6516 11653 6526
rect 11711 6526 11745 6550
rect 11711 6516 11745 6526
rect 11803 6526 11837 6550
rect 11803 6516 11837 6526
rect 11895 6526 11929 6550
rect 11895 6516 11929 6526
rect 11987 6526 12021 6550
rect 11987 6516 12021 6526
rect 12079 6526 12113 6550
rect 12079 6516 12113 6526
rect 12171 6526 12205 6550
rect 12171 6516 12205 6526
rect 12263 6526 12297 6550
rect 12787 6526 12821 6550
rect 12879 6526 12913 6550
rect 12971 6526 13005 6550
rect 13063 6526 13097 6550
rect 13155 6526 13189 6550
rect 13247 6526 13281 6550
rect 13339 6526 13373 6550
rect 13431 6526 13465 6550
rect 13523 6526 13557 6550
rect 13615 6526 13649 6550
rect 13707 6526 13741 6550
rect 13799 6526 13833 6550
rect 13891 6526 13925 6550
rect 13983 6526 14017 6550
rect 14075 6526 14109 6550
rect 14167 6526 14201 6550
rect 14259 6526 14293 6550
rect 14351 6526 14385 6550
rect 14443 6526 14477 6550
rect 12263 6516 12297 6526
rect 12787 6516 12815 6526
rect 12815 6516 12821 6526
rect 12879 6516 12907 6526
rect 12907 6516 12913 6526
rect 12971 6516 12999 6526
rect 12999 6516 13005 6526
rect 13063 6516 13091 6526
rect 13091 6516 13097 6526
rect 13155 6516 13183 6526
rect 13183 6516 13189 6526
rect 13247 6516 13275 6526
rect 13275 6516 13281 6526
rect 13339 6516 13367 6526
rect 13367 6516 13373 6526
rect 13431 6516 13459 6526
rect 13459 6516 13465 6526
rect 13523 6516 13551 6526
rect 13551 6516 13557 6526
rect 13615 6516 13643 6526
rect 13643 6516 13649 6526
rect 13707 6516 13735 6526
rect 13735 6516 13741 6526
rect 13799 6516 13827 6526
rect 13827 6516 13833 6526
rect 13891 6516 13919 6526
rect 13919 6516 13925 6526
rect 13983 6516 14011 6526
rect 14011 6516 14017 6526
rect 14075 6516 14103 6526
rect 14103 6516 14109 6526
rect 14167 6516 14195 6526
rect 14195 6516 14201 6526
rect 14259 6516 14287 6526
rect 14287 6516 14293 6526
rect 14351 6516 14379 6526
rect 14379 6516 14385 6526
rect 14443 6516 14471 6526
rect 14471 6516 14477 6526
rect 14535 6516 14569 6550
rect 24156 6569 24190 6570
rect 24156 6536 24159 6569
rect 24159 6536 24190 6569
rect 24075 6401 24109 6405
rect 24075 6371 24079 6401
rect 24079 6371 24109 6401
rect 11526 6211 11560 6221
rect 11526 6187 11560 6211
rect 11618 6211 11652 6221
rect 11618 6187 11652 6211
rect 11710 6211 11744 6221
rect 11710 6187 11744 6211
rect 11802 6211 11836 6221
rect 11802 6187 11836 6211
rect 11894 6211 11928 6221
rect 11894 6187 11928 6211
rect 11986 6211 12020 6221
rect 11986 6187 12020 6211
rect 12078 6211 12112 6221
rect 12078 6187 12112 6211
rect 12170 6211 12204 6221
rect 12170 6187 12204 6211
rect 12262 6211 12296 6221
rect 12262 6187 12296 6211
rect 12354 6211 12388 6221
rect 12354 6187 12388 6211
rect 12446 6211 12480 6221
rect 12446 6187 12480 6211
rect 12538 6211 12572 6221
rect 12538 6187 12572 6211
rect 12630 6211 12664 6221
rect 12630 6187 12664 6211
rect 12722 6211 12756 6221
rect 12722 6187 12756 6211
rect 12814 6211 12848 6221
rect 12814 6187 12848 6211
rect 12906 6211 12940 6221
rect 12906 6187 12940 6211
rect 12998 6211 13032 6221
rect 12998 6187 13032 6211
rect 13090 6211 13124 6221
rect 13090 6187 13124 6211
rect 13182 6211 13216 6221
rect 13182 6187 13216 6211
rect 13274 6211 13308 6221
rect 13274 6187 13308 6211
rect 13366 6202 13397 6221
rect 13397 6202 13400 6221
rect 13366 6187 13400 6202
rect 13458 6187 13492 6221
rect 13550 6211 13584 6221
rect 13550 6187 13584 6211
rect 13642 6211 13676 6221
rect 13642 6187 13676 6211
rect 13734 6211 13768 6221
rect 13734 6187 13768 6211
rect 13826 6211 13860 6221
rect 13826 6187 13860 6211
rect 13918 6211 13952 6221
rect 13918 6187 13952 6211
rect 14010 6211 14044 6221
rect 14010 6187 14044 6211
rect 14102 6211 14103 6221
rect 14103 6211 14136 6221
rect 14194 6211 14228 6221
rect 14102 6187 14136 6211
rect 14194 6187 14228 6211
rect 14286 6211 14320 6221
rect 14286 6187 14320 6211
rect 14378 6211 14412 6221
rect 14378 6187 14412 6211
rect 14470 6211 14504 6221
rect 14470 6187 14504 6211
rect 14562 6187 14596 6221
rect 14654 6205 14674 6221
rect 14674 6205 14688 6221
rect 14654 6187 14688 6205
rect 14746 6211 14780 6221
rect 14746 6187 14780 6211
rect 14838 6211 14872 6221
rect 14838 6187 14872 6211
rect 14930 6211 14964 6221
rect 14930 6187 14964 6211
rect 15022 6211 15056 6221
rect 15022 6187 15056 6211
rect 15114 6211 15148 6221
rect 15114 6187 15148 6211
rect 15206 6211 15240 6221
rect 15206 6187 15240 6211
rect 15298 6211 15332 6221
rect 15298 6187 15332 6211
rect 15390 6211 15424 6221
rect 15390 6187 15424 6211
rect 15482 6211 15516 6221
rect 15482 6187 15516 6211
rect 15574 6211 15608 6221
rect 15574 6187 15608 6211
rect 15666 6211 15700 6221
rect 15666 6187 15700 6211
rect 15758 6211 15792 6221
rect 15758 6187 15792 6211
rect 15850 6211 15884 6221
rect 15850 6187 15884 6211
rect 15942 6211 15976 6221
rect 15942 6187 15976 6211
rect 16034 6211 16068 6221
rect 16034 6187 16068 6211
rect 16126 6211 16160 6221
rect 16126 6187 16160 6211
rect 16218 6211 16252 6221
rect 16218 6187 16252 6211
rect 16310 6211 16344 6221
rect 16310 6187 16344 6211
rect 16402 6211 16436 6221
rect 16402 6187 16436 6211
rect 16494 6211 16528 6221
rect 16494 6187 16528 6211
rect 16586 6211 16620 6221
rect 16586 6187 16620 6211
rect 16678 6211 16712 6221
rect 16678 6187 16712 6211
rect 16770 6211 16804 6221
rect 16770 6187 16804 6211
rect 16862 6211 16896 6221
rect 16862 6187 16896 6211
rect 16954 6187 16988 6221
rect 17046 6207 17066 6221
rect 17066 6207 17080 6221
rect 17046 6187 17080 6207
rect 17138 6211 17172 6221
rect 17138 6187 17172 6211
rect 17230 6211 17264 6221
rect 17230 6187 17264 6211
rect 17322 6211 17356 6221
rect 17322 6187 17356 6211
rect 17414 6211 17448 6221
rect 17414 6187 17448 6211
rect 17506 6211 17540 6221
rect 17506 6187 17540 6211
rect 17598 6211 17632 6221
rect 17598 6187 17632 6211
rect 17690 6211 17724 6221
rect 17690 6187 17724 6211
rect 17782 6211 17816 6221
rect 17782 6187 17816 6211
rect 17874 6211 17908 6221
rect 17874 6187 17908 6211
rect 17966 6211 18000 6221
rect 17966 6187 18000 6211
rect 18058 6211 18092 6221
rect 18058 6187 18092 6211
rect 18150 6211 18184 6221
rect 18150 6187 18184 6211
rect 18242 6211 18276 6221
rect 18242 6187 18276 6211
rect 18334 6211 18368 6221
rect 18334 6187 18368 6211
rect 18426 6211 18460 6221
rect 18426 6187 18460 6211
rect 18518 6211 18552 6221
rect 18518 6187 18552 6211
rect 18610 6211 18644 6221
rect 18610 6187 18644 6211
rect 18702 6211 18736 6221
rect 18702 6187 18736 6211
rect 18794 6211 18828 6221
rect 18794 6187 18828 6211
rect 18886 6211 18920 6221
rect 18886 6187 18920 6211
rect 18978 6211 19012 6221
rect 18978 6187 19012 6211
rect 19070 6211 19104 6221
rect 19070 6187 19104 6211
rect 19162 6211 19196 6221
rect 19162 6187 19196 6211
rect 19254 6211 19288 6221
rect 19254 6187 19288 6211
rect 19346 6187 19380 6221
rect 19438 6207 19458 6221
rect 19458 6207 19472 6221
rect 19438 6187 19472 6207
rect 19530 6211 19564 6221
rect 19530 6187 19564 6211
rect 19622 6211 19656 6221
rect 19622 6187 19656 6211
rect 19714 6211 19748 6221
rect 19714 6187 19748 6211
rect 19806 6211 19840 6221
rect 19806 6187 19840 6211
rect 19898 6211 19932 6221
rect 19898 6187 19932 6211
rect 19990 6211 20024 6221
rect 19990 6187 20024 6211
rect 20082 6211 20116 6221
rect 20082 6187 20116 6211
rect 20174 6211 20208 6221
rect 20174 6187 20208 6211
rect 20266 6211 20300 6221
rect 20266 6187 20300 6211
rect 20358 6211 20392 6221
rect 20358 6187 20392 6211
rect 20450 6211 20484 6221
rect 20450 6187 20484 6211
rect 20542 6211 20576 6221
rect 20542 6187 20576 6211
rect 20634 6211 20668 6221
rect 20634 6187 20668 6211
rect 20726 6211 20760 6221
rect 20726 6187 20760 6211
rect 20818 6211 20852 6221
rect 20818 6187 20852 6211
rect 20910 6211 20944 6221
rect 20910 6187 20944 6211
rect 21002 6211 21036 6221
rect 21002 6187 21036 6211
rect 21094 6211 21128 6221
rect 21094 6187 21128 6211
rect 21186 6211 21220 6221
rect 21186 6187 21220 6211
rect 21278 6211 21312 6221
rect 21278 6187 21312 6211
rect 21370 6211 21404 6221
rect 21370 6187 21404 6211
rect 21462 6211 21496 6221
rect 21462 6187 21496 6211
rect 21554 6211 21588 6221
rect 21554 6187 21588 6211
rect 21646 6211 21680 6221
rect 21646 6187 21680 6211
rect 21738 6187 21772 6221
rect 21830 6208 21850 6221
rect 21850 6208 21864 6221
rect 21830 6187 21864 6208
rect 21922 6211 21956 6221
rect 21922 6187 21956 6211
rect 22014 6211 22048 6221
rect 22014 6187 22048 6211
rect 22106 6211 22140 6221
rect 22106 6187 22140 6211
rect 22198 6211 22232 6221
rect 22198 6187 22232 6211
rect 22290 6211 22324 6221
rect 22290 6187 22324 6211
rect 22382 6211 22416 6221
rect 22382 6187 22416 6211
rect 22474 6211 22508 6221
rect 22474 6187 22508 6211
rect 22566 6211 22600 6221
rect 22566 6187 22600 6211
rect 22658 6211 22692 6221
rect 22658 6187 22692 6211
rect 22750 6211 22784 6221
rect 22750 6187 22784 6211
rect 22842 6211 22876 6221
rect 22842 6187 22876 6211
rect 22934 6211 22968 6221
rect 22934 6187 22968 6211
rect 23026 6211 23060 6221
rect 23026 6187 23060 6211
rect 23118 6211 23152 6221
rect 23118 6187 23152 6211
rect 23210 6211 23244 6221
rect 23210 6187 23244 6211
rect 23302 6211 23336 6221
rect 23302 6187 23336 6211
rect 23394 6211 23428 6221
rect 23394 6187 23428 6211
rect 11619 6017 11653 6051
rect 11530 5890 11563 5900
rect 11563 5890 11564 5900
rect 11530 5866 11564 5890
rect 11711 5813 11745 5847
rect 11987 6017 12021 6051
rect 11891 5946 11925 5980
rect 12075 5829 12093 5847
rect 12093 5829 12109 5847
rect 12075 5813 12109 5829
rect 12723 6025 12757 6051
rect 12723 6017 12744 6025
rect 12744 6017 12757 6025
rect 12631 5949 12665 5983
rect 12263 5839 12265 5847
rect 12265 5839 12297 5847
rect 12263 5813 12297 5839
rect 12723 5881 12757 5915
rect 12999 5839 13008 5847
rect 13008 5839 13033 5847
rect 12999 5813 13033 5839
rect 13275 5949 13309 5983
rect 13550 5787 13584 5789
rect 13550 5755 13571 5787
rect 13571 5755 13584 5787
rect 13831 5953 13865 5987
rect 14011 6017 14045 6051
rect 13920 5890 13921 5900
rect 13921 5890 13954 5900
rect 13920 5866 13954 5890
rect 14103 5813 14137 5847
rect 14379 6017 14413 6051
rect 14242 5949 14276 5983
rect 14467 5829 14485 5847
rect 14485 5829 14501 5847
rect 14467 5813 14501 5829
rect 15115 6025 15149 6051
rect 15115 6017 15136 6025
rect 15136 6017 15149 6025
rect 15023 5949 15057 5983
rect 14655 5839 14657 5847
rect 14657 5839 14689 5847
rect 14655 5813 14689 5839
rect 15115 5881 15149 5915
rect 15391 5839 15400 5847
rect 15400 5839 15425 5847
rect 15391 5813 15425 5839
rect 15667 5949 15701 5983
rect 15768 5913 15802 5917
rect 15768 5883 15777 5913
rect 15777 5883 15802 5913
rect 15939 5787 15973 5800
rect 15939 5766 15963 5787
rect 15963 5766 15973 5787
rect 16220 5952 16254 5986
rect 16403 6017 16437 6051
rect 16313 5890 16347 5901
rect 16313 5867 16347 5890
rect 16211 5789 16245 5812
rect 16211 5778 16212 5789
rect 16212 5778 16245 5789
rect 16495 5813 16529 5847
rect 16771 6017 16805 6051
rect 16631 5948 16665 5982
rect 16859 5829 16877 5847
rect 16877 5829 16893 5847
rect 16859 5813 16893 5829
rect 17507 6025 17541 6051
rect 17507 6017 17528 6025
rect 17528 6017 17541 6025
rect 17415 5949 17449 5983
rect 17047 5839 17049 5847
rect 17049 5839 17081 5847
rect 17047 5813 17081 5839
rect 17507 5881 17541 5915
rect 17783 5839 17792 5847
rect 17792 5839 17817 5847
rect 17783 5813 17817 5839
rect 18059 5949 18093 5983
rect 18158 5913 18192 5918
rect 18158 5884 18169 5913
rect 18169 5884 18192 5913
rect 18327 5787 18361 5803
rect 18327 5769 18355 5787
rect 18355 5769 18361 5787
rect 18795 6017 18829 6051
rect 18615 5950 18649 5984
rect 18705 5890 18739 5900
rect 18705 5866 18739 5890
rect 18607 5789 18641 5801
rect 18607 5767 18638 5789
rect 18638 5767 18641 5789
rect 18887 5813 18921 5847
rect 19163 6017 19197 6051
rect 19026 5946 19060 5980
rect 19251 5829 19269 5847
rect 19269 5829 19285 5847
rect 19251 5813 19285 5829
rect 19899 6025 19933 6051
rect 19899 6017 19920 6025
rect 19920 6017 19933 6025
rect 19807 5949 19841 5983
rect 19439 5839 19441 5847
rect 19441 5839 19473 5847
rect 19439 5813 19473 5839
rect 19899 5881 19933 5915
rect 20175 5839 20184 5847
rect 20184 5839 20209 5847
rect 20175 5813 20209 5839
rect 20451 5949 20485 5983
rect 20549 5913 20583 5920
rect 20549 5886 20561 5913
rect 20561 5886 20583 5913
rect 20724 5753 20747 5786
rect 20747 5753 20758 5786
rect 20724 5752 20758 5753
rect 21187 6017 21221 6051
rect 21006 5949 21040 5983
rect 21100 5890 21131 5902
rect 21131 5890 21134 5902
rect 21100 5868 21134 5890
rect 21007 5789 21041 5817
rect 21007 5783 21030 5789
rect 21030 5783 21041 5789
rect 21279 5813 21313 5847
rect 21555 6017 21589 6051
rect 21417 5945 21451 5979
rect 21643 5829 21661 5847
rect 21661 5829 21677 5847
rect 21643 5813 21677 5829
rect 22291 6025 22325 6051
rect 22291 6017 22312 6025
rect 22312 6017 22325 6025
rect 22199 5949 22233 5983
rect 21831 5839 21833 5847
rect 21833 5839 21865 5847
rect 21831 5813 21865 5839
rect 22291 5881 22325 5915
rect 22567 5839 22576 5847
rect 22576 5839 22601 5847
rect 22567 5813 22601 5839
rect 22843 5949 22877 5983
rect 22940 5913 22974 5918
rect 22940 5884 22953 5913
rect 22953 5884 22974 5913
rect 23115 5753 23139 5787
rect 23139 5753 23149 5787
rect 24265 6501 24299 6515
rect 24265 6481 24299 6501
rect 24541 6672 24575 6732
rect 24629 6672 24663 6732
rect 24541 6534 24575 6594
rect 24629 6534 24663 6594
rect 30506 6603 30540 6637
rect 24585 6441 24619 6475
rect 24349 6401 24383 6404
rect 24349 6370 24379 6401
rect 24379 6370 24383 6401
rect 24488 6371 24522 6405
rect 24526 6278 24560 6312
rect 24785 6296 24819 6330
rect 30708 6335 30742 6336
rect 30708 6302 30742 6335
rect 30800 6302 30834 6336
rect 30892 6335 30925 6336
rect 30925 6335 30926 6336
rect 30892 6302 30926 6335
rect 30984 6302 31018 6336
rect 24786 6203 24820 6237
rect 25227 6198 25261 6232
rect 25959 6201 25993 6235
rect 26085 6201 26119 6235
rect 27171 6201 27205 6235
rect 27297 6201 27331 6235
rect 28383 6201 28417 6235
rect 28509 6201 28543 6235
rect 29595 6201 29629 6235
rect 29721 6201 29755 6235
rect 30326 6223 30360 6283
rect 30414 6223 30448 6283
rect 24028 6135 24062 6169
rect 24120 6140 24154 6169
rect 24212 6140 24246 6169
rect 24120 6135 24127 6140
rect 24127 6135 24154 6140
rect 24212 6135 24245 6140
rect 24245 6135 24246 6140
rect 24304 6135 24338 6169
rect 23394 6075 23422 6107
rect 23422 6075 23428 6107
rect 23394 6073 23428 6075
rect 24396 6135 24430 6169
rect 25183 6079 25217 6139
rect 25271 6082 25305 6142
rect 25915 6082 25949 6142
rect 26020 6082 26054 6142
rect 26129 6082 26163 6142
rect 27127 6082 27161 6142
rect 27231 6082 27265 6142
rect 27341 6082 27375 6142
rect 28339 6082 28373 6142
rect 28444 6082 28478 6142
rect 28553 6082 28587 6142
rect 29551 6082 29585 6142
rect 29658 6082 29692 6142
rect 29765 6082 29799 6142
rect 30326 6085 30360 6145
rect 30414 6085 30448 6145
rect 30510 6085 30544 6145
rect 30606 6085 30640 6145
rect 30255 5994 30289 6028
rect 30462 5992 30496 6026
rect 30702 6024 30736 6026
rect 30702 5992 30716 6024
rect 30716 5992 30736 6024
rect 30909 5992 30943 6026
rect 25536 5881 25570 5941
rect 25626 5881 25660 5941
rect 26268 5881 26302 5941
rect 26375 5881 26409 5941
rect 26478 5881 26512 5941
rect 27480 5881 27514 5941
rect 27586 5881 27620 5941
rect 27690 5881 27724 5941
rect 28818 5881 28852 5941
rect 28926 5881 28960 5941
rect 29028 5881 29062 5941
rect 29673 5881 29707 5941
rect 29762 5881 29796 5941
rect 30326 5882 30360 5942
rect 30414 5882 30448 5942
rect 30510 5882 30544 5942
rect 30606 5882 30640 5942
rect 23402 5789 23436 5817
rect 23402 5783 23422 5789
rect 23422 5783 23436 5789
rect 24596 5807 24630 5841
rect 25580 5797 25614 5831
rect 26312 5797 26346 5831
rect 26434 5797 26468 5831
rect 27524 5797 27558 5831
rect 27646 5797 27680 5831
rect 28862 5797 28896 5831
rect 28984 5797 29018 5831
rect 29718 5797 29752 5831
rect 24516 5697 24550 5757
rect 24676 5697 24710 5757
rect 30326 5744 30360 5804
rect 30414 5744 30448 5804
rect 30708 5758 30742 5792
rect 30800 5758 30834 5792
rect 30892 5758 30926 5792
rect 30984 5758 31018 5792
rect 11526 5653 11560 5677
rect 11526 5643 11560 5653
rect 11618 5653 11652 5677
rect 11618 5643 11652 5653
rect 11710 5653 11744 5677
rect 11710 5643 11744 5653
rect 11802 5653 11836 5677
rect 11802 5643 11836 5653
rect 11894 5653 11928 5677
rect 11894 5643 11928 5653
rect 11986 5653 12020 5677
rect 11986 5643 12020 5653
rect 12078 5653 12112 5677
rect 12078 5643 12112 5653
rect 12170 5653 12204 5677
rect 12170 5643 12204 5653
rect 12262 5653 12296 5677
rect 12262 5643 12296 5653
rect 12354 5653 12388 5677
rect 12354 5643 12388 5653
rect 12446 5653 12480 5677
rect 12446 5643 12480 5653
rect 12538 5653 12572 5677
rect 12538 5643 12572 5653
rect 12630 5653 12664 5677
rect 12630 5643 12664 5653
rect 12722 5653 12756 5677
rect 12722 5643 12756 5653
rect 12814 5653 12848 5677
rect 12814 5643 12848 5653
rect 12906 5653 12940 5677
rect 12906 5643 12940 5653
rect 12998 5653 13032 5677
rect 12998 5643 13032 5653
rect 13090 5653 13124 5677
rect 13090 5643 13124 5653
rect 13182 5653 13216 5677
rect 13182 5643 13216 5653
rect 13274 5653 13308 5677
rect 13274 5643 13308 5653
rect 13366 5653 13400 5677
rect 13366 5643 13400 5653
rect 13458 5653 13492 5677
rect 13458 5643 13492 5653
rect 13550 5653 13584 5677
rect 13550 5643 13584 5653
rect 13642 5653 13676 5677
rect 13642 5643 13676 5653
rect 13734 5653 13768 5677
rect 13734 5643 13768 5653
rect 13826 5653 13860 5677
rect 13826 5643 13860 5653
rect 13918 5653 13952 5677
rect 13918 5643 13952 5653
rect 14010 5653 14044 5677
rect 14010 5643 14044 5653
rect 14102 5653 14136 5677
rect 14102 5643 14136 5653
rect 14194 5653 14228 5677
rect 14194 5643 14228 5653
rect 14286 5653 14320 5677
rect 14286 5643 14320 5653
rect 14378 5653 14412 5677
rect 14378 5643 14412 5653
rect 14470 5653 14504 5677
rect 14470 5643 14504 5653
rect 14562 5653 14596 5677
rect 14562 5643 14596 5653
rect 14654 5653 14688 5677
rect 14654 5643 14688 5653
rect 14746 5653 14780 5677
rect 14746 5643 14780 5653
rect 14838 5653 14872 5677
rect 14838 5643 14872 5653
rect 14930 5653 14964 5677
rect 14930 5643 14964 5653
rect 15022 5653 15056 5677
rect 15022 5643 15056 5653
rect 15114 5653 15148 5677
rect 15114 5643 15148 5653
rect 15206 5653 15240 5677
rect 15206 5643 15240 5653
rect 15298 5653 15332 5677
rect 15298 5643 15332 5653
rect 15390 5653 15424 5677
rect 15390 5643 15424 5653
rect 15482 5653 15516 5677
rect 15482 5643 15516 5653
rect 15574 5653 15608 5677
rect 15574 5643 15608 5653
rect 15666 5653 15700 5677
rect 15666 5643 15700 5653
rect 15758 5653 15792 5677
rect 15758 5643 15792 5653
rect 15850 5653 15884 5677
rect 15850 5643 15884 5653
rect 15942 5653 15976 5677
rect 15942 5643 15976 5653
rect 16034 5653 16068 5677
rect 16034 5643 16068 5653
rect 16126 5653 16160 5677
rect 16126 5643 16160 5653
rect 16218 5653 16252 5677
rect 16218 5643 16252 5653
rect 16310 5653 16344 5677
rect 16310 5643 16344 5653
rect 16402 5653 16436 5677
rect 16402 5643 16436 5653
rect 16494 5653 16528 5677
rect 16494 5643 16528 5653
rect 16586 5653 16620 5677
rect 16586 5643 16620 5653
rect 16678 5653 16712 5677
rect 16678 5643 16712 5653
rect 16770 5653 16804 5677
rect 16770 5643 16804 5653
rect 16862 5653 16896 5677
rect 16862 5643 16896 5653
rect 16954 5653 16988 5677
rect 16954 5643 16988 5653
rect 17046 5653 17080 5677
rect 17046 5643 17080 5653
rect 17138 5653 17172 5677
rect 17138 5643 17172 5653
rect 17230 5653 17264 5677
rect 17230 5643 17264 5653
rect 17322 5653 17356 5677
rect 17322 5643 17356 5653
rect 17414 5653 17448 5677
rect 17414 5643 17448 5653
rect 17506 5653 17540 5677
rect 17506 5643 17540 5653
rect 17598 5653 17632 5677
rect 17598 5643 17632 5653
rect 17690 5653 17724 5677
rect 17690 5643 17724 5653
rect 17782 5653 17816 5677
rect 17782 5643 17816 5653
rect 17874 5653 17908 5677
rect 17874 5643 17908 5653
rect 17966 5653 18000 5677
rect 17966 5643 18000 5653
rect 18058 5653 18092 5677
rect 18058 5643 18092 5653
rect 18150 5653 18184 5677
rect 18150 5643 18184 5653
rect 18242 5653 18276 5677
rect 18242 5643 18276 5653
rect 18334 5653 18368 5677
rect 18334 5643 18368 5653
rect 18426 5653 18460 5677
rect 18426 5643 18460 5653
rect 18518 5653 18552 5677
rect 18518 5643 18552 5653
rect 18610 5653 18644 5677
rect 18610 5643 18644 5653
rect 18702 5653 18736 5677
rect 18702 5643 18736 5653
rect 18794 5653 18828 5677
rect 18794 5643 18828 5653
rect 18886 5653 18920 5677
rect 18886 5643 18920 5653
rect 18978 5653 19012 5677
rect 18978 5643 19012 5653
rect 19070 5653 19104 5677
rect 19070 5643 19104 5653
rect 19162 5653 19196 5677
rect 19162 5643 19196 5653
rect 19254 5653 19288 5677
rect 19254 5643 19288 5653
rect 19346 5653 19380 5677
rect 19346 5643 19380 5653
rect 19438 5653 19472 5677
rect 19438 5643 19472 5653
rect 19530 5653 19564 5677
rect 19530 5643 19564 5653
rect 19622 5653 19656 5677
rect 19622 5643 19656 5653
rect 19714 5653 19748 5677
rect 19714 5643 19748 5653
rect 19806 5653 19840 5677
rect 19806 5643 19840 5653
rect 19898 5653 19932 5677
rect 19898 5643 19932 5653
rect 19990 5653 20024 5677
rect 19990 5643 20024 5653
rect 20082 5653 20116 5677
rect 20082 5643 20116 5653
rect 20174 5653 20208 5677
rect 20174 5643 20208 5653
rect 20266 5653 20300 5677
rect 20266 5643 20300 5653
rect 20358 5653 20392 5677
rect 20358 5643 20392 5653
rect 20450 5653 20484 5677
rect 20450 5643 20484 5653
rect 20542 5653 20576 5677
rect 20542 5643 20576 5653
rect 20634 5653 20668 5677
rect 20634 5643 20668 5653
rect 20726 5653 20760 5677
rect 20726 5643 20760 5653
rect 20818 5653 20852 5677
rect 20818 5643 20852 5653
rect 20910 5653 20944 5677
rect 20910 5643 20944 5653
rect 21002 5653 21036 5677
rect 21002 5643 21036 5653
rect 21094 5653 21128 5677
rect 21094 5643 21128 5653
rect 21186 5653 21220 5677
rect 21186 5643 21220 5653
rect 21278 5653 21312 5677
rect 21278 5643 21312 5653
rect 21370 5653 21404 5677
rect 21370 5643 21404 5653
rect 21462 5653 21496 5677
rect 21462 5643 21496 5653
rect 21554 5653 21588 5677
rect 21554 5643 21588 5653
rect 21646 5653 21680 5677
rect 21646 5643 21680 5653
rect 21738 5653 21772 5677
rect 21738 5643 21772 5653
rect 21830 5653 21864 5677
rect 21830 5643 21864 5653
rect 21922 5653 21956 5677
rect 21922 5643 21956 5653
rect 22014 5653 22048 5677
rect 22014 5643 22048 5653
rect 22106 5653 22140 5677
rect 22106 5643 22140 5653
rect 22198 5653 22232 5677
rect 22198 5643 22232 5653
rect 22290 5653 22324 5677
rect 22290 5643 22324 5653
rect 22382 5653 22416 5677
rect 22382 5643 22416 5653
rect 22474 5653 22508 5677
rect 22474 5643 22508 5653
rect 22566 5653 22600 5677
rect 22566 5643 22600 5653
rect 22658 5653 22692 5677
rect 22658 5643 22692 5653
rect 22750 5653 22784 5677
rect 22750 5643 22784 5653
rect 22842 5653 22876 5677
rect 22842 5643 22876 5653
rect 22934 5653 22968 5677
rect 22934 5643 22968 5653
rect 23026 5653 23060 5677
rect 23026 5643 23060 5653
rect 23118 5653 23152 5677
rect 23118 5643 23152 5653
rect 23210 5653 23244 5677
rect 23210 5643 23244 5653
rect 23302 5653 23336 5677
rect 23302 5643 23336 5653
rect 23394 5653 23428 5677
rect 23394 5643 23428 5653
rect 24516 5559 24550 5619
rect 11086 5522 11120 5532
rect 11086 5498 11120 5522
rect 11178 5522 11212 5532
rect 11178 5498 11212 5522
rect 11270 5522 11304 5532
rect 11270 5498 11304 5522
rect 11362 5522 11396 5532
rect 11362 5498 11396 5522
rect 11454 5522 11488 5532
rect 11454 5498 11488 5522
rect 11546 5522 11580 5532
rect 11546 5498 11580 5522
rect 11638 5522 11672 5532
rect 11638 5498 11672 5522
rect 11730 5522 11764 5532
rect 11730 5498 11764 5522
rect 11822 5522 11856 5532
rect 11822 5498 11856 5522
rect 11894 5522 11914 5532
rect 11914 5522 11928 5532
rect 11986 5522 12006 5532
rect 12006 5522 12020 5532
rect 12078 5522 12098 5532
rect 12098 5522 12112 5532
rect 12170 5522 12190 5532
rect 12190 5522 12204 5532
rect 12262 5522 12282 5532
rect 12282 5522 12296 5532
rect 12354 5522 12374 5532
rect 12374 5522 12388 5532
rect 12446 5522 12466 5532
rect 12466 5522 12480 5532
rect 12538 5522 12558 5532
rect 12558 5522 12572 5532
rect 12630 5522 12650 5532
rect 12650 5522 12664 5532
rect 12722 5522 12742 5532
rect 12742 5522 12756 5532
rect 12814 5522 12848 5532
rect 12906 5522 12940 5532
rect 11894 5498 11928 5522
rect 11986 5498 12020 5522
rect 12078 5498 12112 5522
rect 12170 5498 12204 5522
rect 12262 5498 12296 5522
rect 12354 5498 12388 5522
rect 12446 5498 12480 5522
rect 12538 5498 12572 5522
rect 12630 5498 12664 5522
rect 12722 5498 12756 5522
rect 12814 5498 12848 5522
rect 12906 5498 12940 5522
rect 12998 5522 13032 5532
rect 12998 5498 13032 5522
rect 13090 5522 13124 5532
rect 13090 5498 13124 5522
rect 13182 5522 13216 5532
rect 13182 5498 13216 5522
rect 13274 5522 13308 5532
rect 13274 5498 13308 5522
rect 13366 5522 13400 5532
rect 13366 5498 13400 5522
rect 13458 5522 13492 5532
rect 13458 5498 13492 5522
rect 13550 5522 13584 5532
rect 13550 5498 13584 5522
rect 13642 5522 13676 5532
rect 13642 5498 13676 5522
rect 13734 5522 13768 5532
rect 13734 5498 13768 5522
rect 13826 5522 13860 5532
rect 13826 5498 13860 5522
rect 13918 5522 13952 5532
rect 13918 5498 13952 5522
rect 14010 5522 14044 5532
rect 14010 5498 14044 5522
rect 14102 5522 14136 5532
rect 14102 5498 14136 5522
rect 14194 5522 14228 5532
rect 14194 5498 14228 5522
rect 14286 5522 14320 5532
rect 14286 5498 14320 5522
rect 14378 5522 14412 5532
rect 14378 5498 14412 5522
rect 14470 5522 14504 5532
rect 14470 5498 14504 5522
rect 14562 5522 14596 5532
rect 14562 5498 14596 5522
rect 14654 5498 14688 5532
rect 14746 5498 14780 5532
rect 14838 5522 14872 5532
rect 14838 5498 14872 5522
rect 14930 5522 14964 5532
rect 14930 5498 14964 5522
rect 15022 5522 15056 5532
rect 15022 5498 15056 5522
rect 15114 5522 15148 5532
rect 15114 5498 15148 5522
rect 15206 5522 15240 5532
rect 15206 5498 15240 5522
rect 15298 5522 15332 5532
rect 15298 5498 15332 5522
rect 15390 5522 15424 5532
rect 15390 5498 15424 5522
rect 15482 5522 15516 5532
rect 15482 5498 15516 5522
rect 15574 5522 15608 5532
rect 15574 5498 15608 5522
rect 15666 5522 15700 5532
rect 15666 5498 15700 5522
rect 15758 5522 15792 5532
rect 15758 5498 15792 5522
rect 15850 5522 15884 5532
rect 15850 5498 15884 5522
rect 15942 5522 15976 5532
rect 15942 5498 15976 5522
rect 16034 5522 16068 5532
rect 16034 5498 16068 5522
rect 16126 5522 16160 5532
rect 16126 5498 16160 5522
rect 16218 5522 16252 5532
rect 16218 5498 16252 5522
rect 16310 5522 16344 5532
rect 16310 5498 16344 5522
rect 16402 5522 16436 5532
rect 16402 5498 16436 5522
rect 16494 5522 16528 5532
rect 16494 5498 16528 5522
rect 16586 5522 16620 5532
rect 16586 5498 16620 5522
rect 16678 5522 16712 5532
rect 16678 5498 16712 5522
rect 16770 5522 16804 5532
rect 16770 5498 16804 5522
rect 16862 5522 16896 5532
rect 16862 5498 16896 5522
rect 16954 5522 16988 5532
rect 16954 5498 16988 5522
rect 17046 5498 17080 5532
rect 17138 5498 17172 5532
rect 17230 5522 17264 5532
rect 17230 5498 17264 5522
rect 17322 5522 17356 5532
rect 17322 5498 17356 5522
rect 17414 5522 17448 5532
rect 17414 5498 17448 5522
rect 17506 5522 17540 5532
rect 17506 5498 17540 5522
rect 17598 5522 17632 5532
rect 17598 5498 17632 5522
rect 17690 5522 17724 5532
rect 17690 5498 17724 5522
rect 17782 5522 17816 5532
rect 17782 5498 17816 5522
rect 17874 5522 17908 5532
rect 17874 5498 17908 5522
rect 17966 5522 18000 5532
rect 17966 5498 18000 5522
rect 18058 5522 18092 5532
rect 18058 5498 18092 5522
rect 18150 5522 18184 5532
rect 18150 5498 18184 5522
rect 18242 5522 18276 5532
rect 18242 5498 18276 5522
rect 18334 5522 18368 5532
rect 18334 5498 18368 5522
rect 18426 5522 18460 5532
rect 18426 5498 18460 5522
rect 18518 5522 18552 5532
rect 18518 5498 18552 5522
rect 18610 5522 18644 5532
rect 18610 5498 18644 5522
rect 18702 5522 18736 5532
rect 18702 5498 18736 5522
rect 18794 5522 18828 5532
rect 18794 5498 18828 5522
rect 18886 5522 18920 5532
rect 18886 5498 18920 5522
rect 18978 5522 19012 5532
rect 18978 5498 19012 5522
rect 19070 5522 19104 5532
rect 19070 5498 19104 5522
rect 19162 5522 19196 5532
rect 19162 5498 19196 5522
rect 19254 5522 19288 5532
rect 19254 5498 19288 5522
rect 19346 5522 19380 5532
rect 19346 5498 19380 5522
rect 19438 5498 19472 5532
rect 19530 5498 19564 5532
rect 19622 5522 19656 5532
rect 19622 5498 19656 5522
rect 19714 5522 19748 5532
rect 19714 5498 19748 5522
rect 19806 5522 19840 5532
rect 19806 5498 19840 5522
rect 19898 5522 19932 5532
rect 19898 5498 19932 5522
rect 19990 5522 20024 5532
rect 19990 5498 20024 5522
rect 20082 5522 20116 5532
rect 20082 5498 20116 5522
rect 20174 5522 20208 5532
rect 20174 5498 20208 5522
rect 20266 5522 20300 5532
rect 20266 5498 20300 5522
rect 20358 5522 20392 5532
rect 20358 5498 20392 5522
rect 20450 5522 20484 5532
rect 20450 5498 20484 5522
rect 20542 5522 20576 5532
rect 20542 5498 20576 5522
rect 20634 5522 20668 5532
rect 20634 5498 20668 5522
rect 20726 5522 20760 5532
rect 20726 5498 20760 5522
rect 20818 5522 20852 5532
rect 20818 5498 20852 5522
rect 20910 5522 20944 5532
rect 20910 5498 20944 5522
rect 21002 5522 21036 5532
rect 21002 5498 21036 5522
rect 21094 5522 21128 5532
rect 21094 5498 21128 5522
rect 21186 5522 21220 5532
rect 21186 5498 21220 5522
rect 21278 5522 21312 5532
rect 21278 5498 21312 5522
rect 21370 5522 21404 5532
rect 21370 5498 21404 5522
rect 21462 5522 21496 5532
rect 21462 5498 21496 5522
rect 21554 5522 21588 5532
rect 21554 5498 21588 5522
rect 21646 5522 21680 5532
rect 21646 5498 21680 5522
rect 21738 5522 21772 5532
rect 21738 5498 21772 5522
rect 21830 5498 21864 5532
rect 21922 5498 21956 5532
rect 22014 5522 22048 5532
rect 22014 5498 22048 5522
rect 22106 5522 22140 5532
rect 22106 5498 22140 5522
rect 22198 5522 22232 5532
rect 22198 5498 22232 5522
rect 22290 5522 22324 5532
rect 22290 5498 22324 5522
rect 22382 5522 22416 5532
rect 22382 5498 22416 5522
rect 22474 5522 22508 5532
rect 22474 5498 22508 5522
rect 22566 5522 22600 5532
rect 22566 5498 22600 5522
rect 22658 5522 22692 5532
rect 22658 5498 22692 5522
rect 22750 5522 22784 5532
rect 22750 5498 22784 5522
rect 22842 5522 22876 5532
rect 22842 5498 22876 5522
rect 22934 5522 22968 5532
rect 22934 5498 22968 5522
rect 23026 5522 23060 5532
rect 23026 5498 23060 5522
rect 23118 5522 23152 5532
rect 23118 5498 23152 5522
rect 23210 5522 23244 5532
rect 23210 5498 23244 5522
rect 23302 5522 23336 5532
rect 23302 5498 23336 5522
rect 23394 5522 23428 5532
rect 23394 5498 23428 5522
rect 24676 5559 24710 5619
rect 11088 5220 11122 5224
rect 11088 5190 11094 5220
rect 11094 5190 11122 5220
rect 13001 5382 13035 5394
rect 13001 5360 13026 5382
rect 13026 5360 13035 5382
rect 13829 5059 13863 5093
rect 13915 5420 13949 5430
rect 13915 5396 13924 5420
rect 13924 5396 13949 5420
rect 14469 5260 14503 5294
rect 14361 5224 14395 5228
rect 14361 5194 14393 5224
rect 14393 5194 14395 5224
rect 14745 5150 14770 5158
rect 14770 5150 14779 5158
rect 14745 5124 14779 5150
rect 15021 5336 15055 5362
rect 15021 5328 15034 5336
rect 15034 5328 15055 5336
rect 15113 5260 15147 5294
rect 15021 5192 15055 5226
rect 15757 5328 15791 5362
rect 15481 5150 15513 5158
rect 15513 5150 15515 5158
rect 15481 5124 15515 5150
rect 15669 5140 15685 5158
rect 15685 5140 15703 5158
rect 15669 5124 15703 5140
rect 15893 5258 15927 5292
rect 16033 5124 16067 5158
rect 16125 5328 16159 5362
rect 16213 5201 16215 5207
rect 16215 5201 16247 5207
rect 16213 5173 16247 5201
rect 16304 5262 16338 5296
rect 16308 5100 16342 5128
rect 16308 5094 16316 5100
rect 16316 5094 16342 5100
rect 16861 5260 16895 5294
rect 16755 5224 16789 5230
rect 16755 5196 16785 5224
rect 16785 5196 16789 5224
rect 16594 5064 16599 5089
rect 16599 5064 16628 5089
rect 16594 5055 16628 5064
rect 17137 5150 17162 5158
rect 17162 5150 17171 5158
rect 17137 5124 17171 5150
rect 17413 5336 17447 5362
rect 17413 5328 17426 5336
rect 17426 5328 17447 5336
rect 17505 5260 17539 5294
rect 17413 5192 17447 5226
rect 18149 5328 18183 5362
rect 17873 5150 17905 5158
rect 17905 5150 17907 5158
rect 17873 5124 17907 5150
rect 18061 5140 18077 5158
rect 18077 5140 18095 5158
rect 18061 5124 18095 5140
rect 18285 5258 18319 5292
rect 18425 5124 18459 5158
rect 18517 5328 18551 5362
rect 18610 5201 18641 5208
rect 18641 5201 18644 5208
rect 18610 5174 18644 5201
rect 18696 5262 18730 5296
rect 18708 5100 18742 5115
rect 18708 5081 18742 5100
rect 19253 5260 19287 5294
rect 19145 5224 19179 5231
rect 19145 5197 19177 5224
rect 19177 5197 19179 5224
rect 18982 5064 18991 5088
rect 18991 5064 19016 5088
rect 18982 5054 19016 5064
rect 19529 5150 19554 5158
rect 19554 5150 19563 5158
rect 19529 5124 19563 5150
rect 19805 5336 19839 5362
rect 19805 5328 19818 5336
rect 19818 5328 19839 5336
rect 19897 5260 19931 5294
rect 19805 5192 19839 5226
rect 20541 5328 20575 5362
rect 20265 5150 20297 5158
rect 20297 5150 20299 5158
rect 20265 5124 20299 5150
rect 20453 5140 20469 5158
rect 20469 5140 20487 5158
rect 20453 5124 20487 5140
rect 20677 5259 20711 5293
rect 20817 5124 20851 5158
rect 20909 5328 20943 5362
rect 21001 5201 21033 5208
rect 21033 5201 21035 5208
rect 21001 5174 21035 5201
rect 21088 5263 21122 5297
rect 21096 5100 21130 5123
rect 21096 5089 21100 5100
rect 21100 5089 21130 5100
rect 21645 5260 21679 5294
rect 21539 5224 21573 5228
rect 21539 5194 21569 5224
rect 21569 5194 21573 5224
rect 21376 5064 21383 5094
rect 21383 5064 21410 5094
rect 21376 5060 21410 5064
rect 21921 5150 21946 5158
rect 21946 5150 21955 5158
rect 21921 5124 21955 5150
rect 22197 5336 22231 5362
rect 22197 5328 22210 5336
rect 22210 5328 22231 5336
rect 22289 5260 22323 5294
rect 22197 5192 22231 5226
rect 22933 5328 22967 5362
rect 22657 5150 22689 5158
rect 22689 5150 22691 5158
rect 22657 5124 22691 5150
rect 22845 5140 22861 5158
rect 22861 5140 22879 5158
rect 22845 5124 22879 5140
rect 23038 5255 23072 5289
rect 24516 5421 24550 5481
rect 24676 5421 24710 5481
rect 23209 5124 23243 5158
rect 23301 5328 23335 5362
rect 23393 5247 23427 5281
rect 24516 5283 24550 5343
rect 24676 5283 24710 5343
rect 24516 5145 24550 5205
rect 24676 5145 24710 5205
rect 24516 5007 24550 5067
rect 24676 5007 24710 5067
rect 11086 4964 11120 4988
rect 11086 4954 11120 4964
rect 11178 4964 11212 4988
rect 11178 4954 11212 4964
rect 11270 4964 11304 4988
rect 11270 4954 11304 4964
rect 11362 4964 11396 4988
rect 11362 4954 11396 4964
rect 11454 4964 11488 4988
rect 11454 4954 11488 4964
rect 11546 4964 11580 4988
rect 11546 4954 11580 4964
rect 11638 4964 11672 4988
rect 11638 4954 11672 4964
rect 11730 4964 11764 4988
rect 11730 4954 11764 4964
rect 11822 4964 11856 4988
rect 11822 4954 11856 4964
rect 11894 4964 11928 4988
rect 11986 4964 12020 4988
rect 12078 4964 12112 4988
rect 12170 4964 12204 4988
rect 12262 4964 12296 4988
rect 12354 4964 12388 4988
rect 12446 4964 12480 4988
rect 12538 4964 12572 4988
rect 12630 4964 12664 4988
rect 12722 4964 12756 4988
rect 12814 4964 12848 4988
rect 12906 4964 12940 4988
rect 12998 4964 13032 4988
rect 13090 4964 13124 4988
rect 13182 4964 13216 4988
rect 13274 4964 13308 4988
rect 13366 4964 13400 4988
rect 13458 4964 13492 4988
rect 13550 4964 13584 4988
rect 13642 4964 13676 4988
rect 13734 4964 13768 4988
rect 13826 4964 13860 4988
rect 13918 4964 13952 4988
rect 14010 4964 14044 4988
rect 14102 4964 14136 4988
rect 14194 4964 14228 4988
rect 14286 4964 14320 4988
rect 14378 4964 14412 4988
rect 14470 4964 14504 4988
rect 14562 4964 14596 4988
rect 14654 4964 14688 4988
rect 14746 4964 14780 4988
rect 14838 4964 14872 4988
rect 14930 4964 14964 4988
rect 15022 4964 15056 4988
rect 15114 4964 15148 4988
rect 15206 4964 15240 4988
rect 15298 4964 15332 4988
rect 15390 4964 15424 4988
rect 15482 4964 15516 4988
rect 15574 4964 15608 4988
rect 15666 4964 15700 4988
rect 15758 4964 15792 4988
rect 15850 4964 15884 4988
rect 15942 4964 15976 4988
rect 16034 4964 16068 4988
rect 16126 4964 16160 4988
rect 16218 4964 16252 4988
rect 16310 4964 16344 4988
rect 16402 4964 16436 4988
rect 16494 4964 16528 4988
rect 16586 4964 16620 4988
rect 16678 4964 16712 4988
rect 16770 4964 16804 4988
rect 16862 4964 16896 4988
rect 16954 4964 16988 4988
rect 17046 4964 17080 4988
rect 17138 4964 17172 4988
rect 17230 4964 17264 4988
rect 17322 4964 17356 4988
rect 17414 4964 17448 4988
rect 17506 4964 17540 4988
rect 17598 4964 17632 4988
rect 17690 4964 17724 4988
rect 17782 4964 17816 4988
rect 17874 4964 17908 4988
rect 17966 4964 18000 4988
rect 18058 4964 18092 4988
rect 18150 4964 18184 4988
rect 18242 4964 18276 4988
rect 18334 4964 18368 4988
rect 18426 4964 18460 4988
rect 18518 4964 18552 4988
rect 18610 4964 18644 4988
rect 18702 4964 18736 4988
rect 18794 4964 18828 4988
rect 18886 4964 18920 4988
rect 18978 4964 19012 4988
rect 19070 4964 19104 4988
rect 19162 4964 19196 4988
rect 19254 4964 19288 4988
rect 19346 4964 19380 4988
rect 19438 4964 19472 4988
rect 19530 4964 19564 4988
rect 19622 4964 19656 4988
rect 19714 4964 19748 4988
rect 19806 4964 19840 4988
rect 19898 4964 19932 4988
rect 11894 4954 11914 4964
rect 11914 4954 11928 4964
rect 11986 4954 12006 4964
rect 12006 4954 12020 4964
rect 12078 4954 12098 4964
rect 12098 4954 12112 4964
rect 12170 4954 12190 4964
rect 12190 4954 12204 4964
rect 12262 4954 12282 4964
rect 12282 4954 12296 4964
rect 12354 4954 12374 4964
rect 12374 4954 12388 4964
rect 12446 4954 12466 4964
rect 12466 4954 12480 4964
rect 12538 4954 12558 4964
rect 12558 4954 12572 4964
rect 12630 4954 12650 4964
rect 12650 4954 12664 4964
rect 12722 4954 12742 4964
rect 12742 4954 12756 4964
rect 12814 4954 12834 4964
rect 12834 4954 12848 4964
rect 12906 4954 12926 4964
rect 12926 4954 12940 4964
rect 12998 4954 13018 4964
rect 13018 4954 13032 4964
rect 13090 4954 13110 4964
rect 13110 4954 13124 4964
rect 13182 4954 13202 4964
rect 13202 4954 13216 4964
rect 13274 4954 13294 4964
rect 13294 4954 13308 4964
rect 13366 4954 13386 4964
rect 13386 4954 13400 4964
rect 13458 4954 13478 4964
rect 13478 4954 13492 4964
rect 13550 4954 13570 4964
rect 13570 4954 13584 4964
rect 13642 4954 13662 4964
rect 13662 4954 13676 4964
rect 13734 4954 13754 4964
rect 13754 4954 13768 4964
rect 13826 4954 13846 4964
rect 13846 4954 13860 4964
rect 13918 4954 13938 4964
rect 13938 4954 13952 4964
rect 14010 4954 14030 4964
rect 14030 4954 14044 4964
rect 14102 4954 14122 4964
rect 14122 4954 14136 4964
rect 14194 4954 14214 4964
rect 14214 4954 14228 4964
rect 14286 4954 14306 4964
rect 14306 4954 14320 4964
rect 14378 4954 14398 4964
rect 14398 4954 14412 4964
rect 14470 4954 14490 4964
rect 14490 4954 14504 4964
rect 14562 4954 14582 4964
rect 14582 4954 14596 4964
rect 14654 4954 14674 4964
rect 14674 4954 14688 4964
rect 14746 4954 14766 4964
rect 14766 4954 14780 4964
rect 14838 4954 14858 4964
rect 14858 4954 14872 4964
rect 14930 4954 14950 4964
rect 14950 4954 14964 4964
rect 15022 4954 15042 4964
rect 15042 4954 15056 4964
rect 15114 4954 15134 4964
rect 15134 4954 15148 4964
rect 15206 4954 15226 4964
rect 15226 4954 15240 4964
rect 15298 4954 15318 4964
rect 15318 4954 15332 4964
rect 15390 4954 15410 4964
rect 15410 4954 15424 4964
rect 15482 4954 15502 4964
rect 15502 4954 15516 4964
rect 15574 4954 15594 4964
rect 15594 4954 15608 4964
rect 15666 4954 15686 4964
rect 15686 4954 15700 4964
rect 15758 4954 15778 4964
rect 15778 4954 15792 4964
rect 15850 4954 15870 4964
rect 15870 4954 15884 4964
rect 15942 4954 15962 4964
rect 15962 4954 15976 4964
rect 16034 4954 16054 4964
rect 16054 4954 16068 4964
rect 16126 4954 16146 4964
rect 16146 4954 16160 4964
rect 16218 4954 16238 4964
rect 16238 4954 16252 4964
rect 16310 4954 16330 4964
rect 16330 4954 16344 4964
rect 16402 4954 16422 4964
rect 16422 4954 16436 4964
rect 16494 4954 16514 4964
rect 16514 4954 16528 4964
rect 16586 4954 16606 4964
rect 16606 4954 16620 4964
rect 16678 4954 16698 4964
rect 16698 4954 16712 4964
rect 16770 4954 16790 4964
rect 16790 4954 16804 4964
rect 16862 4954 16882 4964
rect 16882 4954 16896 4964
rect 16954 4954 16974 4964
rect 16974 4954 16988 4964
rect 17046 4954 17066 4964
rect 17066 4954 17080 4964
rect 17138 4954 17158 4964
rect 17158 4954 17172 4964
rect 17230 4954 17250 4964
rect 17250 4954 17264 4964
rect 17322 4954 17342 4964
rect 17342 4954 17356 4964
rect 17414 4954 17434 4964
rect 17434 4954 17448 4964
rect 17506 4954 17526 4964
rect 17526 4954 17540 4964
rect 17598 4954 17618 4964
rect 17618 4954 17632 4964
rect 17690 4954 17710 4964
rect 17710 4954 17724 4964
rect 17782 4954 17802 4964
rect 17802 4954 17816 4964
rect 17874 4954 17894 4964
rect 17894 4954 17908 4964
rect 17966 4954 17986 4964
rect 17986 4954 18000 4964
rect 18058 4954 18078 4964
rect 18078 4954 18092 4964
rect 18150 4954 18170 4964
rect 18170 4954 18184 4964
rect 18242 4954 18262 4964
rect 18262 4954 18276 4964
rect 18334 4954 18354 4964
rect 18354 4954 18368 4964
rect 18426 4954 18446 4964
rect 18446 4954 18460 4964
rect 18518 4954 18538 4964
rect 18538 4954 18552 4964
rect 18610 4954 18630 4964
rect 18630 4954 18644 4964
rect 18702 4954 18722 4964
rect 18722 4954 18736 4964
rect 18794 4954 18814 4964
rect 18814 4954 18828 4964
rect 18886 4954 18906 4964
rect 18906 4954 18920 4964
rect 18978 4954 18998 4964
rect 18998 4954 19012 4964
rect 19070 4954 19090 4964
rect 19090 4954 19104 4964
rect 19162 4954 19182 4964
rect 19182 4954 19196 4964
rect 19254 4954 19274 4964
rect 19274 4954 19288 4964
rect 19346 4954 19366 4964
rect 19366 4954 19380 4964
rect 19438 4954 19458 4964
rect 19458 4954 19472 4964
rect 19530 4954 19550 4964
rect 19550 4954 19564 4964
rect 19622 4954 19642 4964
rect 19642 4954 19656 4964
rect 19714 4954 19734 4964
rect 19734 4954 19748 4964
rect 19806 4954 19826 4964
rect 19826 4954 19840 4964
rect 19898 4954 19932 4964
rect 19990 4964 20024 4988
rect 19990 4954 20024 4964
rect 20082 4964 20116 4988
rect 20082 4954 20116 4964
rect 20174 4964 20208 4988
rect 20174 4954 20208 4964
rect 20266 4964 20300 4988
rect 20266 4954 20300 4964
rect 20358 4964 20392 4988
rect 20358 4954 20392 4964
rect 20450 4964 20484 4988
rect 20450 4954 20484 4964
rect 20542 4964 20576 4988
rect 20542 4954 20576 4964
rect 20634 4964 20668 4988
rect 20634 4954 20668 4964
rect 20726 4964 20760 4988
rect 20726 4954 20760 4964
rect 20818 4964 20852 4988
rect 20818 4954 20852 4964
rect 20910 4964 20944 4988
rect 20910 4954 20944 4964
rect 21002 4964 21036 4988
rect 21002 4954 21036 4964
rect 21094 4964 21128 4988
rect 21094 4954 21128 4964
rect 21186 4964 21220 4988
rect 21186 4954 21220 4964
rect 21278 4964 21312 4988
rect 21278 4954 21312 4964
rect 21370 4964 21404 4988
rect 21370 4954 21404 4964
rect 21462 4964 21496 4988
rect 21462 4954 21496 4964
rect 21554 4964 21588 4988
rect 21554 4954 21588 4964
rect 21646 4964 21680 4988
rect 21646 4954 21680 4964
rect 21738 4964 21772 4988
rect 21738 4954 21772 4964
rect 21830 4964 21864 4988
rect 21830 4954 21864 4964
rect 21922 4964 21956 4988
rect 21922 4954 21956 4964
rect 22014 4964 22048 4988
rect 22014 4954 22048 4964
rect 22106 4964 22140 4988
rect 22106 4954 22140 4964
rect 22198 4964 22232 4988
rect 22198 4954 22232 4964
rect 22290 4964 22324 4988
rect 22290 4954 22324 4964
rect 22382 4964 22416 4988
rect 22382 4954 22416 4964
rect 22474 4964 22508 4988
rect 22474 4954 22508 4964
rect 22566 4964 22600 4988
rect 22566 4954 22600 4964
rect 22658 4964 22692 4988
rect 22658 4954 22692 4964
rect 22750 4964 22784 4988
rect 22750 4954 22784 4964
rect 22842 4964 22876 4988
rect 22842 4954 22876 4964
rect 22934 4964 22968 4988
rect 22934 4954 22968 4964
rect 23026 4964 23060 4988
rect 23026 4954 23060 4964
rect 23118 4964 23152 4988
rect 23118 4954 23152 4964
rect 23210 4964 23244 4988
rect 23210 4954 23244 4964
rect 23302 4964 23336 4988
rect 23302 4954 23336 4964
rect 23394 4964 23428 4988
rect 23394 4954 23428 4964
rect 24516 4869 24550 4929
rect 24676 4869 24710 4929
rect 24516 4731 24550 4791
rect 24676 4731 24710 4791
rect 25217 4710 25251 4744
rect 25297 4710 25331 4744
rect 25377 4710 25411 4744
rect 25457 4710 25491 4744
rect 25949 4710 25983 4744
rect 26029 4710 26063 4744
rect 26109 4710 26143 4744
rect 26189 4710 26223 4744
rect 26557 4710 26591 4744
rect 26637 4710 26671 4744
rect 26717 4710 26751 4744
rect 26797 4710 26831 4744
rect 27161 4710 27195 4744
rect 27241 4710 27275 4744
rect 27321 4710 27355 4744
rect 27401 4710 27435 4744
rect 27769 4710 27803 4744
rect 27849 4710 27883 4744
rect 27929 4710 27963 4744
rect 28009 4710 28043 4744
rect 28499 4710 28533 4744
rect 28579 4710 28613 4744
rect 28659 4710 28693 4744
rect 28739 4710 28773 4744
rect 29107 4710 29141 4744
rect 29187 4710 29221 4744
rect 29267 4710 29301 4744
rect 29347 4710 29381 4744
rect 29841 4710 29875 4744
rect 29921 4710 29955 4744
rect 30001 4710 30035 4744
rect 30081 4710 30115 4744
rect 11118 4624 11152 4658
rect 11210 4624 11244 4658
rect 11302 4624 11336 4658
rect 11394 4624 11428 4658
rect 11486 4624 11520 4658
rect 11578 4624 11612 4658
rect 11670 4624 11704 4658
rect 11762 4624 11796 4658
rect 11854 4624 11888 4658
rect 13660 4649 13694 4659
rect 13660 4625 13694 4649
rect 13752 4649 13786 4659
rect 13752 4625 13786 4649
rect 13844 4649 13878 4659
rect 13844 4625 13878 4649
rect 13917 4649 13936 4659
rect 13936 4649 13951 4659
rect 14009 4649 14028 4659
rect 14028 4649 14043 4659
rect 14101 4649 14120 4659
rect 14120 4649 14135 4659
rect 14193 4649 14212 4659
rect 14212 4649 14227 4659
rect 14285 4649 14304 4659
rect 14304 4649 14319 4659
rect 14377 4649 14396 4659
rect 14396 4649 14411 4659
rect 14469 4649 14488 4659
rect 14488 4649 14503 4659
rect 14561 4649 14580 4659
rect 14580 4649 14595 4659
rect 14653 4649 14672 4659
rect 14672 4649 14687 4659
rect 14745 4649 14764 4659
rect 14764 4649 14779 4659
rect 14837 4649 14856 4659
rect 14856 4649 14871 4659
rect 14929 4649 14948 4659
rect 14948 4649 14963 4659
rect 15021 4649 15040 4659
rect 15040 4649 15055 4659
rect 15113 4649 15132 4659
rect 15132 4649 15147 4659
rect 15205 4649 15224 4659
rect 15224 4649 15239 4659
rect 15297 4649 15316 4659
rect 15316 4649 15331 4659
rect 15389 4649 15408 4659
rect 15408 4649 15423 4659
rect 15481 4649 15515 4659
rect 13917 4625 13951 4649
rect 14009 4625 14043 4649
rect 14101 4625 14135 4649
rect 14193 4625 14227 4649
rect 14285 4625 14319 4649
rect 14377 4625 14411 4649
rect 14469 4625 14503 4649
rect 14561 4625 14595 4649
rect 14653 4625 14687 4649
rect 14745 4625 14779 4649
rect 14837 4625 14871 4649
rect 14929 4625 14963 4649
rect 15021 4625 15055 4649
rect 15113 4625 15147 4649
rect 15205 4625 15239 4649
rect 15297 4625 15331 4649
rect 15389 4625 15423 4649
rect 15481 4625 15515 4649
rect 15573 4649 15607 4659
rect 15573 4625 15607 4649
rect 15665 4649 15699 4659
rect 15665 4625 15699 4649
rect 15757 4649 15791 4659
rect 15757 4625 15791 4649
rect 15849 4649 15883 4659
rect 15849 4625 15883 4649
rect 15941 4649 15975 4659
rect 15941 4625 15975 4649
rect 16033 4649 16067 4659
rect 16033 4625 16067 4649
rect 16125 4649 16159 4659
rect 16125 4625 16159 4649
rect 16217 4649 16251 4659
rect 16217 4625 16251 4649
rect 16309 4649 16343 4659
rect 16309 4625 16343 4649
rect 16401 4649 16435 4659
rect 16401 4625 16435 4649
rect 16493 4649 16527 4659
rect 16493 4625 16527 4649
rect 16585 4649 16619 4659
rect 16585 4625 16619 4649
rect 16677 4649 16711 4659
rect 16677 4625 16711 4649
rect 16769 4649 16803 4659
rect 16769 4625 16803 4649
rect 16861 4649 16895 4659
rect 16861 4625 16895 4649
rect 16953 4649 16987 4659
rect 16953 4625 16987 4649
rect 17045 4649 17079 4659
rect 17045 4625 17079 4649
rect 17137 4649 17171 4659
rect 17137 4625 17171 4649
rect 17229 4649 17263 4659
rect 17229 4625 17263 4649
rect 17321 4649 17355 4659
rect 17321 4625 17355 4649
rect 17413 4649 17447 4659
rect 17413 4625 17447 4649
rect 17505 4649 17539 4659
rect 17505 4625 17539 4649
rect 17597 4649 17631 4659
rect 17597 4625 17631 4649
rect 17689 4649 17723 4659
rect 17689 4625 17723 4649
rect 17781 4649 17815 4659
rect 17781 4625 17815 4649
rect 17873 4649 17907 4659
rect 17873 4625 17907 4649
rect 17965 4649 17999 4659
rect 17965 4625 17999 4649
rect 18057 4649 18091 4659
rect 18057 4625 18091 4649
rect 18149 4649 18183 4659
rect 18149 4625 18183 4649
rect 18241 4649 18275 4659
rect 18241 4625 18275 4649
rect 18333 4649 18367 4659
rect 18333 4625 18367 4649
rect 18425 4649 18459 4659
rect 18425 4625 18459 4649
rect 18517 4649 18551 4659
rect 18517 4625 18551 4649
rect 18609 4649 18643 4659
rect 18609 4625 18643 4649
rect 18701 4649 18735 4659
rect 18701 4625 18735 4649
rect 18793 4649 18827 4659
rect 18793 4625 18827 4649
rect 18885 4649 18919 4659
rect 18885 4625 18919 4649
rect 18977 4649 19011 4659
rect 18977 4625 19011 4649
rect 19069 4649 19103 4659
rect 19069 4625 19103 4649
rect 19161 4649 19195 4659
rect 19161 4625 19195 4649
rect 19253 4649 19287 4659
rect 19253 4625 19287 4649
rect 19345 4649 19379 4659
rect 19345 4625 19379 4649
rect 19437 4649 19471 4659
rect 19437 4625 19471 4649
rect 19529 4649 19563 4659
rect 19529 4625 19563 4649
rect 19621 4649 19655 4659
rect 19621 4625 19655 4649
rect 19713 4649 19747 4659
rect 19713 4625 19747 4649
rect 19805 4649 19839 4659
rect 19805 4625 19839 4649
rect 19897 4649 19931 4659
rect 19897 4625 19931 4649
rect 19989 4649 20023 4659
rect 19989 4625 20023 4649
rect 20081 4649 20115 4659
rect 20081 4625 20115 4649
rect 20173 4649 20207 4659
rect 20173 4625 20207 4649
rect 20265 4649 20299 4659
rect 20265 4625 20299 4649
rect 20357 4649 20391 4659
rect 20357 4625 20391 4649
rect 20449 4649 20483 4659
rect 20449 4625 20483 4649
rect 20541 4649 20575 4659
rect 20541 4625 20575 4649
rect 20633 4649 20667 4659
rect 20633 4625 20667 4649
rect 20725 4649 20759 4659
rect 20725 4625 20759 4649
rect 20817 4649 20851 4659
rect 20817 4625 20851 4649
rect 20909 4649 20943 4659
rect 20909 4625 20943 4649
rect 21001 4649 21035 4659
rect 21001 4625 21035 4649
rect 21093 4649 21127 4659
rect 21093 4625 21127 4649
rect 21185 4649 21219 4659
rect 21185 4625 21219 4649
rect 21277 4649 21311 4659
rect 21277 4625 21311 4649
rect 21369 4649 21403 4659
rect 21369 4625 21403 4649
rect 21461 4649 21495 4659
rect 21461 4625 21495 4649
rect 21553 4649 21587 4659
rect 21553 4625 21587 4649
rect 21645 4649 21679 4659
rect 21645 4625 21679 4649
rect 21737 4649 21771 4659
rect 21737 4625 21771 4649
rect 21829 4649 21863 4659
rect 21829 4625 21863 4649
rect 21921 4649 21955 4659
rect 21921 4625 21955 4649
rect 22013 4649 22047 4659
rect 22013 4625 22047 4649
rect 22105 4649 22139 4659
rect 22105 4625 22139 4649
rect 22197 4649 22231 4659
rect 22197 4625 22231 4649
rect 22289 4649 22323 4659
rect 22289 4625 22323 4649
rect 22381 4649 22415 4659
rect 22381 4625 22415 4649
rect 22473 4649 22507 4659
rect 22473 4625 22507 4649
rect 22565 4649 22599 4659
rect 22565 4625 22599 4649
rect 22657 4649 22691 4659
rect 22657 4625 22691 4649
rect 22749 4649 22783 4659
rect 22749 4625 22783 4649
rect 22841 4649 22875 4659
rect 22841 4625 22875 4649
rect 22933 4649 22967 4659
rect 22933 4625 22967 4649
rect 23025 4649 23059 4659
rect 23025 4625 23059 4649
rect 23117 4649 23151 4659
rect 23117 4625 23151 4649
rect 23209 4649 23243 4659
rect 23209 4625 23243 4649
rect 23301 4649 23335 4659
rect 23301 4625 23335 4649
rect 23393 4649 23427 4659
rect 23393 4625 23427 4649
rect 11128 4312 11160 4345
rect 11160 4312 11162 4345
rect 11128 4311 11162 4312
rect 14010 4455 14044 4489
rect 13810 4413 13825 4426
rect 13825 4413 13844 4426
rect 13810 4392 13844 4413
rect 11733 4312 11767 4346
rect 13625 4318 13659 4352
rect 13918 4328 13920 4351
rect 13920 4328 13952 4351
rect 13918 4317 13952 4328
rect 14102 4251 14136 4285
rect 14378 4455 14412 4489
rect 14247 4349 14281 4359
rect 14247 4325 14272 4349
rect 14272 4325 14281 4349
rect 14466 4267 14484 4285
rect 14484 4267 14500 4285
rect 14466 4251 14500 4267
rect 15114 4463 15148 4489
rect 15114 4455 15135 4463
rect 15135 4455 15148 4463
rect 15022 4387 15056 4421
rect 14654 4277 14656 4285
rect 14656 4277 14688 4285
rect 14654 4251 14688 4277
rect 15114 4319 15148 4353
rect 15390 4277 15399 4285
rect 15399 4277 15424 4285
rect 15390 4251 15424 4277
rect 15666 4387 15700 4421
rect 15766 4351 15800 4352
rect 15766 4318 15776 4351
rect 15776 4318 15800 4351
rect 16402 4455 16436 4489
rect 16494 4251 16528 4285
rect 16770 4455 16804 4489
rect 16663 4349 16697 4355
rect 16663 4321 16664 4349
rect 16664 4321 16697 4349
rect 16858 4267 16876 4285
rect 16876 4267 16892 4285
rect 16858 4251 16892 4267
rect 17506 4463 17540 4489
rect 17506 4455 17527 4463
rect 17527 4455 17540 4463
rect 17414 4387 17448 4421
rect 17046 4277 17048 4285
rect 17048 4277 17080 4285
rect 17046 4251 17080 4277
rect 17506 4319 17540 4353
rect 17782 4277 17791 4285
rect 17791 4277 17816 4285
rect 17782 4251 17816 4277
rect 18058 4387 18092 4421
rect 18156 4351 18190 4360
rect 18156 4326 18168 4351
rect 18168 4326 18190 4351
rect 18794 4455 18828 4489
rect 18612 4227 18646 4253
rect 18612 4219 18637 4227
rect 18637 4219 18646 4227
rect 18886 4251 18920 4285
rect 19162 4455 19196 4489
rect 19050 4349 19084 4355
rect 19050 4321 19056 4349
rect 19056 4321 19084 4349
rect 19250 4267 19268 4285
rect 19268 4267 19284 4285
rect 19250 4251 19284 4267
rect 19898 4463 19932 4489
rect 19898 4455 19919 4463
rect 19919 4455 19932 4463
rect 19806 4387 19840 4421
rect 19438 4277 19440 4285
rect 19440 4277 19472 4285
rect 19438 4251 19472 4277
rect 19898 4319 19932 4353
rect 20174 4277 20183 4285
rect 20183 4277 20208 4285
rect 20174 4251 20208 4277
rect 20450 4387 20484 4421
rect 20547 4351 20581 4356
rect 20547 4322 20560 4351
rect 20560 4322 20581 4351
rect 21186 4455 21220 4489
rect 21004 4227 21038 4254
rect 21004 4220 21029 4227
rect 21029 4220 21038 4227
rect 21278 4251 21312 4285
rect 21554 4455 21588 4489
rect 21453 4320 21487 4354
rect 21642 4267 21660 4285
rect 21660 4267 21676 4285
rect 21642 4251 21676 4267
rect 22290 4463 22324 4489
rect 22290 4455 22311 4463
rect 22311 4455 22324 4463
rect 22198 4387 22232 4421
rect 21830 4277 21832 4285
rect 21832 4277 21864 4285
rect 21830 4251 21864 4277
rect 22290 4319 22324 4353
rect 22566 4277 22575 4285
rect 22575 4277 22600 4285
rect 22566 4251 22600 4277
rect 22842 4387 22876 4421
rect 22939 4351 22973 4355
rect 22939 4321 22952 4351
rect 22952 4321 22973 4351
rect 25606 4264 25640 4298
rect 25698 4264 25732 4298
rect 25790 4264 25824 4298
rect 25882 4264 25916 4298
rect 25974 4264 26008 4298
rect 26066 4264 26100 4298
rect 26158 4264 26192 4298
rect 26250 4264 26284 4298
rect 26342 4264 26376 4298
rect 26434 4264 26468 4298
rect 26526 4264 26560 4298
rect 26618 4264 26652 4298
rect 26710 4264 26744 4298
rect 26802 4264 26836 4298
rect 26894 4264 26928 4298
rect 26986 4264 27020 4298
rect 27078 4264 27112 4298
rect 27170 4264 27204 4298
rect 27262 4264 27296 4298
rect 27354 4264 27388 4298
rect 27446 4264 27480 4298
rect 27538 4264 27572 4298
rect 27630 4264 27664 4298
rect 27722 4264 27756 4298
rect 27814 4264 27848 4298
rect 27906 4264 27940 4298
rect 27998 4264 28032 4298
rect 28090 4264 28124 4298
rect 28182 4264 28216 4298
rect 28274 4264 28308 4298
rect 28366 4264 28400 4298
rect 28458 4264 28492 4298
rect 28550 4264 28584 4298
rect 28642 4264 28676 4298
rect 28734 4264 28768 4298
rect 28826 4264 28860 4298
rect 28918 4264 28952 4298
rect 29010 4264 29044 4298
rect 29102 4264 29136 4298
rect 29194 4264 29228 4298
rect 29286 4264 29320 4298
rect 29378 4264 29412 4298
rect 29470 4264 29504 4298
rect 29562 4264 29596 4298
rect 29654 4264 29688 4298
rect 29746 4264 29780 4298
rect 29838 4264 29872 4298
rect 29930 4264 29964 4298
rect 30022 4264 30056 4298
rect 30114 4264 30148 4298
rect 30206 4264 30240 4298
rect 30298 4264 30332 4298
rect 23394 4227 23428 4257
rect 23394 4223 23421 4227
rect 23421 4223 23428 4227
rect 11118 4080 11152 4114
rect 11210 4080 11244 4114
rect 11302 4080 11336 4114
rect 11394 4080 11428 4114
rect 11486 4080 11520 4114
rect 11578 4080 11612 4114
rect 11670 4080 11704 4114
rect 11762 4080 11796 4114
rect 11854 4080 11888 4114
rect 13660 4091 13694 4115
rect 13660 4081 13694 4091
rect 13752 4091 13786 4115
rect 13752 4081 13786 4091
rect 13844 4091 13878 4115
rect 13844 4081 13878 4091
rect 13917 4091 13951 4115
rect 14009 4091 14043 4115
rect 14101 4091 14135 4115
rect 14193 4091 14227 4115
rect 14285 4091 14319 4115
rect 14377 4091 14411 4115
rect 14469 4091 14503 4115
rect 14561 4091 14595 4115
rect 14653 4091 14687 4115
rect 14745 4091 14779 4115
rect 14837 4091 14871 4115
rect 14929 4091 14963 4115
rect 15021 4091 15055 4115
rect 15113 4091 15147 4115
rect 15205 4091 15239 4115
rect 15297 4091 15331 4115
rect 15389 4091 15423 4115
rect 15481 4091 15515 4115
rect 15573 4091 15607 4115
rect 15665 4091 15699 4115
rect 15757 4091 15791 4115
rect 15849 4091 15883 4115
rect 15941 4091 15975 4115
rect 16033 4091 16067 4115
rect 16125 4091 16159 4115
rect 16217 4091 16251 4115
rect 16309 4091 16343 4115
rect 16401 4091 16435 4115
rect 16493 4091 16527 4115
rect 16585 4091 16619 4115
rect 16677 4091 16711 4115
rect 16769 4091 16803 4115
rect 16861 4091 16895 4115
rect 16953 4091 16987 4115
rect 17045 4091 17079 4115
rect 17137 4091 17171 4115
rect 17229 4091 17263 4115
rect 17321 4091 17355 4115
rect 17413 4091 17447 4115
rect 17505 4091 17539 4115
rect 17597 4091 17631 4115
rect 17689 4091 17723 4115
rect 17781 4091 17815 4115
rect 17873 4091 17907 4115
rect 17965 4091 17999 4115
rect 18057 4091 18091 4115
rect 18149 4091 18183 4115
rect 18241 4091 18275 4115
rect 18333 4091 18367 4115
rect 18425 4091 18459 4115
rect 18517 4091 18551 4115
rect 18609 4091 18643 4115
rect 18701 4091 18735 4115
rect 18793 4091 18827 4115
rect 18885 4091 18919 4115
rect 18977 4091 19011 4115
rect 19069 4091 19103 4115
rect 19161 4091 19195 4115
rect 19253 4091 19287 4115
rect 19345 4091 19379 4115
rect 19437 4091 19471 4115
rect 19529 4091 19563 4115
rect 19621 4091 19655 4115
rect 19713 4091 19747 4115
rect 19805 4091 19839 4115
rect 19897 4091 19931 4115
rect 19989 4091 20023 4115
rect 20081 4091 20115 4115
rect 20173 4091 20207 4115
rect 20265 4091 20299 4115
rect 20357 4091 20391 4115
rect 20449 4091 20483 4115
rect 20541 4091 20575 4115
rect 20633 4091 20667 4115
rect 20725 4091 20759 4115
rect 20817 4091 20851 4115
rect 20909 4091 20943 4115
rect 21001 4091 21035 4115
rect 21093 4091 21127 4115
rect 21185 4091 21219 4115
rect 21277 4091 21311 4115
rect 21369 4091 21403 4115
rect 21461 4091 21495 4115
rect 21553 4091 21587 4115
rect 21645 4091 21679 4115
rect 21737 4091 21771 4115
rect 21829 4091 21863 4115
rect 21921 4091 21955 4115
rect 22013 4091 22047 4115
rect 22105 4091 22139 4115
rect 22197 4091 22231 4115
rect 22289 4091 22323 4115
rect 22381 4091 22415 4115
rect 22473 4091 22507 4115
rect 13917 4081 13936 4091
rect 13936 4081 13951 4091
rect 14009 4081 14028 4091
rect 14028 4081 14043 4091
rect 14101 4081 14120 4091
rect 14120 4081 14135 4091
rect 14193 4081 14212 4091
rect 14212 4081 14227 4091
rect 14285 4081 14304 4091
rect 14304 4081 14319 4091
rect 14377 4081 14396 4091
rect 14396 4081 14411 4091
rect 14469 4081 14488 4091
rect 14488 4081 14503 4091
rect 14561 4081 14580 4091
rect 14580 4081 14595 4091
rect 14653 4081 14672 4091
rect 14672 4081 14687 4091
rect 14745 4081 14764 4091
rect 14764 4081 14779 4091
rect 14837 4081 14856 4091
rect 14856 4081 14871 4091
rect 14929 4081 14948 4091
rect 14948 4081 14963 4091
rect 15021 4081 15040 4091
rect 15040 4081 15055 4091
rect 15113 4081 15132 4091
rect 15132 4081 15147 4091
rect 15205 4081 15224 4091
rect 15224 4081 15239 4091
rect 15297 4081 15316 4091
rect 15316 4081 15331 4091
rect 15389 4081 15408 4091
rect 15408 4081 15423 4091
rect 15481 4081 15500 4091
rect 15500 4081 15515 4091
rect 15573 4081 15592 4091
rect 15592 4081 15607 4091
rect 15665 4081 15684 4091
rect 15684 4081 15699 4091
rect 15757 4081 15776 4091
rect 15776 4081 15791 4091
rect 15849 4081 15868 4091
rect 15868 4081 15883 4091
rect 15941 4081 15960 4091
rect 15960 4081 15975 4091
rect 16033 4081 16052 4091
rect 16052 4081 16067 4091
rect 16125 4081 16144 4091
rect 16144 4081 16159 4091
rect 16217 4081 16236 4091
rect 16236 4081 16251 4091
rect 16309 4081 16328 4091
rect 16328 4081 16343 4091
rect 16401 4081 16420 4091
rect 16420 4081 16435 4091
rect 16493 4081 16512 4091
rect 16512 4081 16527 4091
rect 16585 4081 16604 4091
rect 16604 4081 16619 4091
rect 16677 4081 16696 4091
rect 16696 4081 16711 4091
rect 16769 4081 16788 4091
rect 16788 4081 16803 4091
rect 16861 4081 16880 4091
rect 16880 4081 16895 4091
rect 16953 4081 16972 4091
rect 16972 4081 16987 4091
rect 17045 4081 17064 4091
rect 17064 4081 17079 4091
rect 17137 4081 17156 4091
rect 17156 4081 17171 4091
rect 17229 4081 17248 4091
rect 17248 4081 17263 4091
rect 17321 4081 17340 4091
rect 17340 4081 17355 4091
rect 17413 4081 17432 4091
rect 17432 4081 17447 4091
rect 17505 4081 17524 4091
rect 17524 4081 17539 4091
rect 17597 4081 17616 4091
rect 17616 4081 17631 4091
rect 17689 4081 17708 4091
rect 17708 4081 17723 4091
rect 17781 4081 17800 4091
rect 17800 4081 17815 4091
rect 17873 4081 17892 4091
rect 17892 4081 17907 4091
rect 17965 4081 17984 4091
rect 17984 4081 17999 4091
rect 18057 4081 18076 4091
rect 18076 4081 18091 4091
rect 18149 4081 18168 4091
rect 18168 4081 18183 4091
rect 18241 4081 18260 4091
rect 18260 4081 18275 4091
rect 18333 4081 18352 4091
rect 18352 4081 18367 4091
rect 18425 4081 18444 4091
rect 18444 4081 18459 4091
rect 18517 4081 18536 4091
rect 18536 4081 18551 4091
rect 18609 4081 18628 4091
rect 18628 4081 18643 4091
rect 18701 4081 18720 4091
rect 18720 4081 18735 4091
rect 18793 4081 18812 4091
rect 18812 4081 18827 4091
rect 18885 4081 18904 4091
rect 18904 4081 18919 4091
rect 18977 4081 18996 4091
rect 18996 4081 19011 4091
rect 19069 4081 19088 4091
rect 19088 4081 19103 4091
rect 19161 4081 19180 4091
rect 19180 4081 19195 4091
rect 19253 4081 19272 4091
rect 19272 4081 19287 4091
rect 19345 4081 19364 4091
rect 19364 4081 19379 4091
rect 19437 4081 19456 4091
rect 19456 4081 19471 4091
rect 19529 4081 19548 4091
rect 19548 4081 19563 4091
rect 19621 4081 19640 4091
rect 19640 4081 19655 4091
rect 19713 4081 19732 4091
rect 19732 4081 19747 4091
rect 19805 4081 19824 4091
rect 19824 4081 19839 4091
rect 19897 4081 19916 4091
rect 19916 4081 19931 4091
rect 19989 4081 20008 4091
rect 20008 4081 20023 4091
rect 20081 4081 20100 4091
rect 20100 4081 20115 4091
rect 20173 4081 20192 4091
rect 20192 4081 20207 4091
rect 20265 4081 20284 4091
rect 20284 4081 20299 4091
rect 20357 4081 20391 4091
rect 20449 4081 20483 4091
rect 20541 4081 20575 4091
rect 20633 4081 20667 4091
rect 20725 4081 20759 4091
rect 20817 4081 20851 4091
rect 20909 4081 20943 4091
rect 21001 4081 21035 4091
rect 21093 4081 21127 4091
rect 21185 4081 21219 4091
rect 21277 4081 21311 4091
rect 21369 4081 21403 4091
rect 21461 4081 21495 4091
rect 21553 4081 21587 4091
rect 21645 4081 21679 4091
rect 21737 4081 21771 4091
rect 21829 4081 21863 4091
rect 21921 4081 21955 4091
rect 22013 4081 22047 4091
rect 22105 4081 22139 4091
rect 22197 4081 22231 4091
rect 22289 4081 22323 4091
rect 22381 4081 22415 4091
rect 22473 4081 22507 4091
rect 22565 4091 22599 4115
rect 22565 4081 22599 4091
rect 22657 4091 22691 4115
rect 22657 4081 22691 4091
rect 22749 4091 22783 4115
rect 22749 4081 22783 4091
rect 22841 4091 22875 4115
rect 22841 4081 22875 4091
rect 22933 4091 22967 4115
rect 22933 4081 22967 4091
rect 23025 4091 23059 4115
rect 23025 4081 23059 4091
rect 23117 4091 23151 4115
rect 23117 4081 23151 4091
rect 23209 4091 23243 4115
rect 23209 4081 23243 4091
rect 23301 4091 23335 4115
rect 23301 4081 23335 4091
rect 23393 4091 23427 4115
rect 23393 4081 23427 4091
rect 25623 4051 25657 4072
rect 25623 4038 25643 4051
rect 25643 4038 25657 4051
rect 25699 3890 25733 3924
rect 25791 4094 25825 4128
rect 25943 3964 25977 3998
rect 26155 4112 26189 4128
rect 26155 4094 26173 4112
rect 26173 4094 26189 4112
rect 26343 4102 26377 4128
rect 26343 4094 26345 4102
rect 26345 4094 26377 4102
rect 26067 3890 26101 3924
rect 11525 3776 11559 3786
rect 11525 3752 11559 3776
rect 11617 3776 11651 3786
rect 11617 3752 11651 3776
rect 11709 3776 11743 3786
rect 11709 3752 11743 3776
rect 11801 3776 11835 3786
rect 11801 3752 11835 3776
rect 11893 3776 11927 3786
rect 11893 3752 11927 3776
rect 11985 3776 12019 3786
rect 11985 3752 12019 3776
rect 12077 3776 12111 3786
rect 12077 3752 12111 3776
rect 12169 3776 12203 3786
rect 12169 3752 12203 3776
rect 12261 3776 12295 3786
rect 12261 3752 12295 3776
rect 12353 3776 12387 3786
rect 12353 3752 12387 3776
rect 12445 3776 12479 3786
rect 12445 3752 12479 3776
rect 12537 3776 12571 3786
rect 12537 3752 12571 3776
rect 12629 3776 12663 3786
rect 12629 3752 12663 3776
rect 12721 3776 12755 3786
rect 12721 3752 12755 3776
rect 12813 3776 12847 3786
rect 12813 3752 12847 3776
rect 12905 3776 12939 3786
rect 12905 3752 12939 3776
rect 12997 3776 13031 3786
rect 12997 3752 13031 3776
rect 13089 3776 13123 3786
rect 13089 3752 13123 3776
rect 13181 3776 13215 3786
rect 13181 3752 13215 3776
rect 13273 3776 13307 3786
rect 13273 3752 13307 3776
rect 13365 3776 13399 3786
rect 13365 3752 13399 3776
rect 13457 3776 13491 3786
rect 13457 3752 13491 3776
rect 13549 3776 13583 3786
rect 13549 3752 13583 3776
rect 13641 3776 13675 3786
rect 13641 3752 13675 3776
rect 13733 3776 13767 3786
rect 13733 3752 13767 3776
rect 13825 3776 13859 3786
rect 13825 3752 13859 3776
rect 13917 3776 13951 3786
rect 13917 3752 13951 3776
rect 14009 3776 14043 3786
rect 14009 3752 14043 3776
rect 14101 3776 14135 3786
rect 14101 3752 14135 3776
rect 14193 3776 14227 3786
rect 14193 3752 14227 3776
rect 14285 3776 14319 3786
rect 14285 3752 14319 3776
rect 14377 3776 14411 3786
rect 14377 3752 14411 3776
rect 14469 3776 14503 3786
rect 14469 3752 14503 3776
rect 14561 3776 14595 3786
rect 14561 3752 14595 3776
rect 14653 3776 14687 3786
rect 14653 3752 14687 3776
rect 14745 3776 14779 3786
rect 14745 3752 14779 3776
rect 14837 3776 14871 3786
rect 14837 3752 14871 3776
rect 14929 3776 14963 3786
rect 14929 3752 14963 3776
rect 15021 3776 15055 3786
rect 15021 3752 15055 3776
rect 15113 3776 15147 3786
rect 15113 3752 15147 3776
rect 15205 3776 15239 3786
rect 15205 3752 15239 3776
rect 15297 3776 15331 3786
rect 15297 3752 15331 3776
rect 15389 3776 15423 3786
rect 15389 3752 15423 3776
rect 15481 3776 15515 3786
rect 15481 3752 15515 3776
rect 15573 3776 15607 3786
rect 15573 3752 15607 3776
rect 15665 3776 15699 3786
rect 15665 3752 15699 3776
rect 15757 3776 15791 3786
rect 15757 3752 15791 3776
rect 15849 3776 15883 3786
rect 15849 3752 15883 3776
rect 15941 3776 15975 3786
rect 15941 3752 15975 3776
rect 16033 3776 16067 3786
rect 16033 3752 16067 3776
rect 16125 3776 16159 3786
rect 16125 3752 16159 3776
rect 16217 3776 16251 3786
rect 16217 3752 16251 3776
rect 16309 3776 16343 3786
rect 16309 3752 16343 3776
rect 16401 3776 16435 3786
rect 16401 3752 16435 3776
rect 16493 3776 16527 3786
rect 16493 3752 16527 3776
rect 16585 3776 16619 3786
rect 16585 3752 16619 3776
rect 16677 3776 16711 3786
rect 16677 3752 16711 3776
rect 16769 3776 16803 3786
rect 16769 3752 16803 3776
rect 16861 3776 16895 3786
rect 16861 3752 16895 3776
rect 16953 3776 16987 3786
rect 16953 3752 16987 3776
rect 17045 3776 17079 3786
rect 17045 3752 17079 3776
rect 17137 3776 17171 3786
rect 17137 3752 17171 3776
rect 17229 3776 17263 3786
rect 17229 3752 17263 3776
rect 17321 3776 17355 3786
rect 17321 3752 17355 3776
rect 17413 3776 17447 3786
rect 17413 3752 17447 3776
rect 17505 3776 17539 3786
rect 17505 3752 17539 3776
rect 17597 3776 17631 3786
rect 17597 3752 17631 3776
rect 17689 3776 17723 3786
rect 17689 3752 17723 3776
rect 17781 3776 17815 3786
rect 17781 3752 17815 3776
rect 17873 3776 17907 3786
rect 17873 3752 17907 3776
rect 17965 3776 17999 3786
rect 17965 3752 17999 3776
rect 18057 3776 18091 3786
rect 18057 3752 18091 3776
rect 18149 3776 18183 3786
rect 18149 3752 18183 3776
rect 18241 3776 18275 3786
rect 18241 3752 18275 3776
rect 18333 3776 18367 3786
rect 18333 3752 18367 3776
rect 18425 3776 18459 3786
rect 18425 3752 18459 3776
rect 18517 3776 18551 3786
rect 18517 3752 18551 3776
rect 18609 3776 18643 3786
rect 18609 3752 18643 3776
rect 18701 3776 18735 3786
rect 18701 3752 18735 3776
rect 18793 3776 18827 3786
rect 18793 3752 18827 3776
rect 18885 3776 18919 3786
rect 18885 3752 18919 3776
rect 18977 3776 19011 3786
rect 18977 3752 19011 3776
rect 19069 3776 19103 3786
rect 19069 3752 19103 3776
rect 19161 3776 19195 3786
rect 19161 3752 19195 3776
rect 19253 3776 19287 3786
rect 19253 3752 19287 3776
rect 19345 3776 19379 3786
rect 19345 3752 19379 3776
rect 19437 3776 19471 3786
rect 19437 3752 19471 3776
rect 19529 3776 19563 3786
rect 19529 3752 19563 3776
rect 19621 3776 19655 3786
rect 19621 3752 19655 3776
rect 19713 3776 19747 3786
rect 19713 3752 19747 3776
rect 19805 3776 19839 3786
rect 19805 3752 19839 3776
rect 19897 3776 19931 3786
rect 19897 3752 19931 3776
rect 19989 3776 20023 3786
rect 19989 3752 20023 3776
rect 20081 3776 20115 3786
rect 20081 3752 20115 3776
rect 20173 3776 20207 3786
rect 20173 3752 20207 3776
rect 20265 3776 20299 3786
rect 20265 3752 20299 3776
rect 20357 3776 20391 3786
rect 20357 3752 20391 3776
rect 20449 3776 20483 3786
rect 20449 3752 20483 3776
rect 20541 3776 20575 3786
rect 20541 3752 20575 3776
rect 20633 3776 20667 3786
rect 20633 3752 20667 3776
rect 20725 3776 20759 3786
rect 20725 3752 20759 3776
rect 20817 3776 20851 3786
rect 20817 3752 20851 3776
rect 20909 3776 20943 3786
rect 20909 3752 20943 3776
rect 21001 3776 21035 3786
rect 21001 3752 21035 3776
rect 21093 3776 21127 3786
rect 21093 3752 21127 3776
rect 21185 3776 21219 3786
rect 21185 3752 21219 3776
rect 21277 3776 21311 3786
rect 21277 3752 21311 3776
rect 21369 3776 21403 3786
rect 21369 3752 21403 3776
rect 21461 3776 21495 3786
rect 21461 3752 21495 3776
rect 21553 3776 21587 3786
rect 21553 3752 21587 3776
rect 21645 3776 21679 3786
rect 21645 3752 21679 3776
rect 21737 3776 21771 3786
rect 21737 3752 21771 3776
rect 21829 3776 21863 3786
rect 21829 3752 21863 3776
rect 21921 3776 21955 3786
rect 21921 3752 21955 3776
rect 22013 3776 22047 3786
rect 22013 3752 22047 3776
rect 22105 3776 22139 3786
rect 22105 3752 22139 3776
rect 22197 3776 22231 3786
rect 22197 3752 22231 3776
rect 22289 3776 22323 3786
rect 22289 3752 22323 3776
rect 22381 3776 22415 3786
rect 22381 3752 22415 3776
rect 22473 3776 22507 3786
rect 22473 3752 22507 3776
rect 22565 3776 22599 3786
rect 22565 3752 22599 3776
rect 22657 3776 22691 3786
rect 22657 3752 22691 3776
rect 22749 3776 22783 3786
rect 22749 3752 22783 3776
rect 22841 3776 22875 3786
rect 22841 3752 22875 3776
rect 22933 3776 22967 3786
rect 22933 3752 22967 3776
rect 23025 3776 23059 3786
rect 23025 3752 23059 3776
rect 23117 3776 23151 3786
rect 23117 3752 23151 3776
rect 23209 3776 23243 3786
rect 23209 3752 23243 3776
rect 23301 3776 23335 3786
rect 23301 3752 23335 3776
rect 23393 3776 23427 3786
rect 23393 3752 23427 3776
rect 26803 4026 26837 4060
rect 26711 3958 26745 3992
rect 26803 3916 26824 3924
rect 26824 3916 26837 3924
rect 26803 3890 26837 3916
rect 27079 4102 27113 4128
rect 27079 4094 27088 4102
rect 27088 4094 27113 4102
rect 27462 4028 27465 4057
rect 27465 4028 27496 4057
rect 27462 4023 27496 4028
rect 27355 3958 27389 3992
rect 28012 4017 28035 4027
rect 28035 4017 28046 4027
rect 28012 3993 28046 4017
rect 27910 3832 27934 3860
rect 27934 3832 27944 3860
rect 27910 3826 27944 3832
rect 28091 3890 28125 3924
rect 28183 4094 28217 4128
rect 28345 4030 28353 4060
rect 28353 4030 28379 4060
rect 28345 4026 28379 4030
rect 28547 4112 28581 4128
rect 28547 4094 28565 4112
rect 28565 4094 28581 4112
rect 28735 4102 28769 4128
rect 28735 4094 28737 4102
rect 28737 4094 28769 4102
rect 28459 3890 28493 3924
rect 29195 4026 29229 4060
rect 29103 3958 29137 3992
rect 29195 3916 29216 3924
rect 29216 3916 29229 3924
rect 29195 3890 29229 3916
rect 29471 4102 29505 4128
rect 29471 4094 29480 4102
rect 29480 4094 29505 4102
rect 29861 4028 29891 4061
rect 29891 4028 29895 4061
rect 29861 4027 29895 4028
rect 29747 3958 29781 3992
rect 30298 4152 30326 4177
rect 30326 4152 30332 4177
rect 30298 4143 30332 4152
rect 11522 3320 11531 3353
rect 11531 3320 11556 3353
rect 11522 3319 11556 3320
rect 12076 3514 12110 3548
rect 11966 3444 12000 3478
rect 12352 3404 12377 3412
rect 12377 3404 12386 3412
rect 12352 3378 12386 3404
rect 12628 3590 12662 3616
rect 12628 3582 12641 3590
rect 12641 3582 12662 3590
rect 12720 3514 12754 3548
rect 12628 3446 12662 3480
rect 13364 3582 13398 3616
rect 13088 3404 13120 3412
rect 13120 3404 13122 3412
rect 13088 3378 13122 3404
rect 13276 3394 13292 3412
rect 13292 3394 13310 3412
rect 13276 3378 13310 3394
rect 13478 3504 13512 3538
rect 13640 3378 13674 3412
rect 13732 3582 13766 3616
rect 13913 3354 13947 3376
rect 13913 3342 13923 3354
rect 13923 3342 13947 3354
rect 14468 3514 14502 3548
rect 14359 3478 14393 3483
rect 14359 3449 14392 3478
rect 14392 3449 14393 3478
rect 14744 3404 14769 3412
rect 14769 3404 14778 3412
rect 14744 3378 14778 3404
rect 15020 3590 15054 3616
rect 15020 3582 15033 3590
rect 15033 3582 15054 3590
rect 15112 3514 15146 3548
rect 15020 3446 15054 3480
rect 15756 3582 15790 3616
rect 15480 3404 15512 3412
rect 15512 3404 15514 3412
rect 15480 3378 15514 3404
rect 15668 3394 15684 3412
rect 15684 3394 15702 3412
rect 15668 3378 15702 3394
rect 15859 3501 15893 3535
rect 16032 3378 16066 3412
rect 16124 3582 16158 3616
rect 16304 3354 16338 3375
rect 16304 3341 16315 3354
rect 16315 3341 16338 3354
rect 16860 3514 16894 3548
rect 16753 3478 16787 3483
rect 16753 3449 16784 3478
rect 16784 3449 16787 3478
rect 17136 3404 17161 3412
rect 17161 3404 17170 3412
rect 17136 3378 17170 3404
rect 17412 3590 17446 3616
rect 17412 3582 17425 3590
rect 17425 3582 17446 3590
rect 17504 3514 17538 3548
rect 17412 3446 17446 3480
rect 18148 3582 18182 3616
rect 17872 3404 17904 3412
rect 17904 3404 17906 3412
rect 17872 3378 17906 3404
rect 18060 3394 18076 3412
rect 18076 3394 18094 3412
rect 18060 3378 18094 3394
rect 18250 3505 18284 3539
rect 18424 3378 18458 3412
rect 18516 3582 18550 3616
rect 18699 3354 18733 3378
rect 18699 3344 18707 3354
rect 18707 3344 18733 3354
rect 19252 3514 19286 3548
rect 19145 3478 19179 3484
rect 19145 3450 19176 3478
rect 19176 3450 19179 3478
rect 19528 3404 19553 3412
rect 19553 3404 19562 3412
rect 19528 3378 19562 3404
rect 19804 3590 19838 3616
rect 19804 3582 19817 3590
rect 19817 3582 19838 3590
rect 19896 3514 19930 3548
rect 19804 3446 19838 3480
rect 20540 3582 20574 3616
rect 20264 3404 20296 3412
rect 20296 3404 20298 3412
rect 20264 3378 20298 3404
rect 20452 3394 20468 3412
rect 20468 3394 20486 3412
rect 20452 3378 20486 3394
rect 20639 3506 20673 3540
rect 20816 3378 20850 3412
rect 20908 3582 20942 3616
rect 21088 3354 21122 3376
rect 21088 3342 21099 3354
rect 21099 3342 21122 3354
rect 21644 3514 21678 3548
rect 21538 3478 21572 3485
rect 21538 3451 21568 3478
rect 21568 3451 21572 3478
rect 21920 3404 21945 3412
rect 21945 3404 21954 3412
rect 21920 3378 21954 3404
rect 22196 3590 22230 3616
rect 22196 3582 22209 3590
rect 22209 3582 22230 3590
rect 22288 3514 22322 3548
rect 22196 3446 22230 3480
rect 25606 3720 25640 3754
rect 25698 3720 25732 3754
rect 25790 3720 25824 3754
rect 25882 3720 25916 3754
rect 25974 3720 26008 3754
rect 26066 3720 26100 3754
rect 26158 3720 26192 3754
rect 26250 3720 26284 3754
rect 26342 3720 26376 3754
rect 26434 3720 26468 3754
rect 26526 3720 26560 3754
rect 26618 3720 26652 3754
rect 26710 3720 26744 3754
rect 26802 3720 26836 3754
rect 26894 3720 26928 3754
rect 26986 3720 27020 3754
rect 27078 3720 27112 3754
rect 27170 3720 27204 3754
rect 27262 3720 27296 3754
rect 27354 3720 27388 3754
rect 27446 3720 27480 3754
rect 27538 3720 27572 3754
rect 27630 3720 27664 3754
rect 27722 3720 27756 3754
rect 27814 3720 27848 3754
rect 27906 3720 27940 3754
rect 27998 3720 28032 3754
rect 28090 3720 28124 3754
rect 28182 3720 28216 3754
rect 28274 3720 28308 3754
rect 28366 3720 28400 3754
rect 28458 3720 28492 3754
rect 28550 3720 28584 3754
rect 28642 3720 28676 3754
rect 28734 3720 28768 3754
rect 28826 3720 28860 3754
rect 28918 3720 28952 3754
rect 29010 3720 29044 3754
rect 29102 3720 29136 3754
rect 29194 3720 29228 3754
rect 29286 3720 29320 3754
rect 29378 3720 29412 3754
rect 29470 3720 29504 3754
rect 29562 3720 29596 3754
rect 29654 3720 29688 3754
rect 29746 3720 29780 3754
rect 29838 3720 29872 3754
rect 29930 3720 29964 3754
rect 30022 3720 30056 3754
rect 30114 3720 30148 3754
rect 30206 3720 30240 3754
rect 30298 3720 30332 3754
rect 22932 3582 22966 3616
rect 22656 3404 22688 3412
rect 22688 3404 22690 3412
rect 22656 3378 22690 3404
rect 22844 3394 22860 3412
rect 22860 3394 22878 3412
rect 22844 3378 22878 3394
rect 23033 3506 23067 3540
rect 23208 3378 23242 3412
rect 23300 3582 23334 3616
rect 25606 3624 25640 3658
rect 25698 3624 25732 3658
rect 25790 3624 25824 3658
rect 25882 3624 25916 3658
rect 25974 3624 26008 3658
rect 26066 3624 26100 3658
rect 26158 3624 26192 3658
rect 26250 3624 26284 3658
rect 26342 3624 26376 3658
rect 26434 3624 26468 3658
rect 26526 3624 26560 3658
rect 26618 3624 26652 3658
rect 26710 3624 26744 3658
rect 26802 3624 26836 3658
rect 26894 3624 26928 3658
rect 26986 3624 27020 3658
rect 27078 3624 27112 3658
rect 27170 3624 27204 3658
rect 27262 3624 27296 3658
rect 27354 3624 27388 3658
rect 27446 3624 27480 3658
rect 27538 3624 27572 3658
rect 27630 3624 27664 3658
rect 27722 3624 27756 3658
rect 27814 3624 27848 3658
rect 27906 3624 27940 3658
rect 27998 3624 28032 3658
rect 28090 3624 28124 3658
rect 28182 3624 28216 3658
rect 28274 3624 28308 3658
rect 28366 3624 28400 3658
rect 28458 3624 28492 3658
rect 28550 3624 28584 3658
rect 28642 3624 28676 3658
rect 28734 3624 28768 3658
rect 28826 3624 28860 3658
rect 28918 3624 28952 3658
rect 29010 3624 29044 3658
rect 29102 3624 29136 3658
rect 29194 3624 29228 3658
rect 29286 3624 29320 3658
rect 29378 3624 29412 3658
rect 29470 3624 29504 3658
rect 29562 3624 29596 3658
rect 29654 3624 29688 3658
rect 29746 3624 29780 3658
rect 29838 3624 29872 3658
rect 29930 3624 29964 3658
rect 30022 3624 30056 3658
rect 30114 3624 30148 3658
rect 30206 3624 30240 3658
rect 30298 3624 30332 3658
rect 23390 3455 23424 3489
rect 25699 3454 25733 3488
rect 25618 3388 25652 3422
rect 11525 3218 11559 3242
rect 11525 3208 11559 3218
rect 11617 3218 11651 3242
rect 11617 3208 11651 3218
rect 11709 3218 11743 3242
rect 11709 3208 11743 3218
rect 11801 3218 11835 3242
rect 11801 3208 11835 3218
rect 11893 3218 11927 3242
rect 11893 3208 11927 3218
rect 11985 3218 12019 3242
rect 11985 3208 12019 3218
rect 12077 3218 12111 3242
rect 12077 3208 12111 3218
rect 12169 3218 12203 3242
rect 12169 3208 12203 3218
rect 12261 3218 12295 3242
rect 12261 3208 12295 3218
rect 12353 3218 12387 3242
rect 12353 3208 12387 3218
rect 12445 3218 12479 3242
rect 12445 3208 12479 3218
rect 12537 3218 12571 3242
rect 12537 3208 12571 3218
rect 12629 3218 12663 3242
rect 12629 3208 12663 3218
rect 12721 3218 12755 3242
rect 12721 3208 12755 3218
rect 12813 3218 12847 3242
rect 12813 3208 12847 3218
rect 12905 3218 12939 3242
rect 12905 3208 12939 3218
rect 12997 3218 13031 3242
rect 12997 3208 13031 3218
rect 13089 3218 13123 3242
rect 13089 3208 13123 3218
rect 13181 3218 13215 3242
rect 13181 3208 13215 3218
rect 13273 3218 13307 3242
rect 13273 3208 13307 3218
rect 13365 3218 13399 3242
rect 13365 3208 13399 3218
rect 13457 3218 13491 3242
rect 13457 3208 13491 3218
rect 13549 3218 13583 3242
rect 13549 3208 13583 3218
rect 13641 3218 13675 3242
rect 13641 3208 13675 3218
rect 13733 3218 13767 3242
rect 13733 3208 13767 3218
rect 13825 3218 13859 3242
rect 13825 3208 13859 3218
rect 13917 3218 13951 3242
rect 13917 3208 13951 3218
rect 14009 3218 14043 3242
rect 14009 3208 14043 3218
rect 14101 3218 14135 3242
rect 14101 3208 14135 3218
rect 14193 3218 14227 3242
rect 14193 3208 14227 3218
rect 14285 3218 14319 3242
rect 14285 3208 14319 3218
rect 14377 3218 14411 3242
rect 14377 3208 14411 3218
rect 14469 3218 14503 3242
rect 14469 3208 14503 3218
rect 14561 3218 14595 3242
rect 14561 3208 14595 3218
rect 14653 3218 14687 3242
rect 14653 3208 14687 3218
rect 14745 3218 14779 3242
rect 14745 3208 14779 3218
rect 14837 3218 14871 3242
rect 14837 3208 14871 3218
rect 14929 3218 14963 3242
rect 14929 3208 14963 3218
rect 15021 3218 15055 3242
rect 15021 3208 15055 3218
rect 15113 3218 15147 3242
rect 15113 3208 15147 3218
rect 15205 3218 15239 3242
rect 15205 3208 15239 3218
rect 15297 3218 15331 3242
rect 15297 3208 15331 3218
rect 15389 3218 15423 3242
rect 15389 3208 15423 3218
rect 15481 3218 15515 3242
rect 15481 3208 15515 3218
rect 15573 3218 15607 3242
rect 15573 3208 15607 3218
rect 15665 3218 15699 3242
rect 15665 3208 15699 3218
rect 15757 3218 15791 3242
rect 15757 3208 15791 3218
rect 15849 3218 15883 3242
rect 15849 3208 15883 3218
rect 15941 3218 15975 3242
rect 15941 3208 15975 3218
rect 16033 3218 16067 3242
rect 16033 3208 16067 3218
rect 16125 3218 16159 3242
rect 16125 3208 16159 3218
rect 16217 3218 16251 3242
rect 16217 3208 16251 3218
rect 16309 3218 16343 3242
rect 16309 3208 16343 3218
rect 16401 3218 16435 3242
rect 16401 3208 16435 3218
rect 16493 3218 16527 3242
rect 16493 3208 16527 3218
rect 16585 3218 16619 3242
rect 16585 3208 16619 3218
rect 16677 3218 16711 3242
rect 16677 3208 16711 3218
rect 16769 3218 16803 3242
rect 16769 3208 16803 3218
rect 16861 3218 16895 3242
rect 16861 3208 16895 3218
rect 16953 3218 16987 3242
rect 16953 3208 16987 3218
rect 17045 3218 17079 3242
rect 17045 3208 17079 3218
rect 17137 3218 17171 3242
rect 17137 3208 17171 3218
rect 17229 3218 17263 3242
rect 17229 3208 17263 3218
rect 17321 3218 17355 3242
rect 17321 3208 17355 3218
rect 17413 3218 17447 3242
rect 17413 3208 17447 3218
rect 17505 3218 17539 3242
rect 17505 3208 17539 3218
rect 17597 3218 17631 3242
rect 17597 3208 17631 3218
rect 17689 3218 17723 3242
rect 17689 3208 17723 3218
rect 17781 3218 17815 3242
rect 17781 3208 17815 3218
rect 17873 3218 17907 3242
rect 17873 3208 17907 3218
rect 17965 3218 17999 3242
rect 17965 3208 17999 3218
rect 18057 3218 18091 3242
rect 18057 3208 18091 3218
rect 18149 3218 18183 3242
rect 18149 3208 18183 3218
rect 18241 3218 18275 3242
rect 18241 3208 18275 3218
rect 18333 3218 18367 3242
rect 18333 3208 18367 3218
rect 18425 3218 18459 3242
rect 18425 3208 18459 3218
rect 18517 3218 18551 3242
rect 18517 3208 18551 3218
rect 18609 3218 18643 3242
rect 18609 3208 18643 3218
rect 18701 3218 18735 3242
rect 18701 3208 18735 3218
rect 18793 3218 18827 3242
rect 18793 3208 18827 3218
rect 18885 3218 18919 3242
rect 18885 3208 18919 3218
rect 18977 3218 19011 3242
rect 18977 3208 19011 3218
rect 19069 3218 19103 3242
rect 19069 3208 19103 3218
rect 19161 3218 19195 3242
rect 19161 3208 19195 3218
rect 19253 3218 19287 3242
rect 19253 3208 19287 3218
rect 19345 3218 19379 3242
rect 19345 3208 19379 3218
rect 19437 3218 19471 3242
rect 19437 3208 19471 3218
rect 19529 3218 19563 3242
rect 19529 3208 19563 3218
rect 19621 3218 19655 3242
rect 19621 3208 19655 3218
rect 19713 3218 19747 3242
rect 19713 3208 19747 3218
rect 19805 3218 19839 3242
rect 19805 3208 19839 3218
rect 19897 3218 19931 3242
rect 19897 3208 19931 3218
rect 19989 3218 20023 3242
rect 19989 3208 20023 3218
rect 20081 3218 20115 3242
rect 20081 3208 20115 3218
rect 20173 3218 20207 3242
rect 20173 3208 20207 3218
rect 20265 3218 20299 3242
rect 20265 3208 20299 3218
rect 20357 3218 20391 3242
rect 20357 3208 20391 3218
rect 20449 3218 20483 3242
rect 20449 3208 20483 3218
rect 20541 3218 20575 3242
rect 20541 3208 20575 3218
rect 20633 3218 20667 3242
rect 20633 3208 20667 3218
rect 20725 3218 20759 3242
rect 20725 3208 20759 3218
rect 20817 3218 20851 3242
rect 20817 3208 20851 3218
rect 20909 3218 20943 3242
rect 20909 3208 20943 3218
rect 21001 3218 21035 3242
rect 21001 3208 21035 3218
rect 21093 3218 21127 3242
rect 21093 3208 21127 3218
rect 21185 3218 21219 3242
rect 21185 3208 21219 3218
rect 21277 3218 21311 3242
rect 21277 3208 21311 3218
rect 21369 3218 21403 3242
rect 21369 3208 21403 3218
rect 21461 3218 21495 3242
rect 21461 3208 21495 3218
rect 21553 3218 21587 3242
rect 21553 3208 21587 3218
rect 21645 3218 21679 3242
rect 21645 3208 21679 3218
rect 21737 3218 21771 3242
rect 21737 3208 21771 3218
rect 21829 3218 21863 3242
rect 21829 3208 21863 3218
rect 21921 3218 21955 3242
rect 21921 3208 21955 3218
rect 22013 3218 22047 3242
rect 22013 3208 22047 3218
rect 22105 3218 22139 3242
rect 22105 3208 22139 3218
rect 22197 3218 22231 3242
rect 22197 3208 22231 3218
rect 22289 3218 22323 3242
rect 22289 3208 22323 3218
rect 22381 3218 22415 3242
rect 22381 3208 22415 3218
rect 22473 3218 22507 3242
rect 22473 3208 22507 3218
rect 22565 3218 22599 3242
rect 22565 3208 22599 3218
rect 22657 3218 22691 3242
rect 22657 3208 22691 3218
rect 22749 3218 22783 3242
rect 22749 3208 22783 3218
rect 22841 3218 22875 3242
rect 22841 3208 22875 3218
rect 22933 3218 22967 3242
rect 22933 3208 22967 3218
rect 23025 3218 23059 3242
rect 23025 3208 23059 3218
rect 23117 3218 23151 3242
rect 23117 3208 23151 3218
rect 23209 3218 23243 3242
rect 23209 3208 23243 3218
rect 23301 3218 23335 3242
rect 23301 3208 23335 3218
rect 23393 3218 23427 3242
rect 23393 3208 23427 3218
rect 25791 3250 25825 3284
rect 26067 3454 26101 3488
rect 25948 3348 25982 3352
rect 25948 3318 25961 3348
rect 25961 3318 25982 3348
rect 26155 3266 26173 3284
rect 26173 3266 26189 3284
rect 26155 3250 26189 3266
rect 26803 3462 26837 3488
rect 26803 3454 26824 3462
rect 26824 3454 26837 3462
rect 26711 3386 26745 3420
rect 26343 3276 26345 3284
rect 26345 3276 26377 3284
rect 26343 3250 26377 3276
rect 26803 3318 26837 3352
rect 27079 3276 27088 3284
rect 27088 3276 27113 3284
rect 27079 3250 27113 3276
rect 27355 3386 27389 3420
rect 27463 3316 27465 3350
rect 27465 3316 27497 3350
rect 27909 3546 27943 3548
rect 27909 3514 27934 3546
rect 27934 3514 27943 3546
rect 28091 3454 28125 3488
rect 28013 3361 28047 3379
rect 28013 3345 28035 3361
rect 28035 3345 28047 3361
rect 28183 3250 28217 3284
rect 28459 3454 28493 3488
rect 28346 3348 28380 3351
rect 28346 3317 28353 3348
rect 28353 3317 28380 3348
rect 28547 3266 28565 3284
rect 28565 3266 28581 3284
rect 28547 3250 28581 3266
rect 29195 3462 29229 3488
rect 29195 3454 29216 3462
rect 29216 3454 29229 3462
rect 29103 3386 29137 3420
rect 28735 3276 28737 3284
rect 28737 3276 28769 3284
rect 28735 3250 28769 3276
rect 29195 3318 29229 3352
rect 29471 3276 29480 3284
rect 29480 3276 29505 3284
rect 29471 3250 29505 3276
rect 29747 3386 29781 3420
rect 29856 3350 29890 3351
rect 29856 3317 29857 3350
rect 29857 3317 29890 3350
rect 30299 3192 30326 3219
rect 30326 3192 30333 3219
rect 30299 3185 30333 3192
rect 25606 3080 25640 3114
rect 25698 3080 25732 3114
rect 25790 3080 25824 3114
rect 25882 3080 25916 3114
rect 25974 3080 26008 3114
rect 26066 3080 26100 3114
rect 26158 3080 26192 3114
rect 26250 3080 26284 3114
rect 26342 3080 26376 3114
rect 26434 3080 26468 3114
rect 26526 3080 26560 3114
rect 26618 3080 26652 3114
rect 26710 3080 26744 3114
rect 26802 3080 26836 3114
rect 26894 3080 26928 3114
rect 26986 3080 27020 3114
rect 27078 3080 27112 3114
rect 27170 3080 27204 3114
rect 27262 3080 27296 3114
rect 27354 3080 27388 3114
rect 27446 3080 27480 3114
rect 27538 3080 27572 3114
rect 27630 3080 27664 3114
rect 27722 3080 27756 3114
rect 27814 3080 27848 3114
rect 27906 3080 27940 3114
rect 27998 3080 28032 3114
rect 28090 3080 28124 3114
rect 28182 3080 28216 3114
rect 28274 3080 28308 3114
rect 28366 3080 28400 3114
rect 28458 3080 28492 3114
rect 28550 3080 28584 3114
rect 28642 3080 28676 3114
rect 28734 3080 28768 3114
rect 28826 3080 28860 3114
rect 28918 3080 28952 3114
rect 29010 3080 29044 3114
rect 29102 3080 29136 3114
rect 29194 3080 29228 3114
rect 29286 3080 29320 3114
rect 29378 3080 29412 3114
rect 29470 3080 29504 3114
rect 29562 3080 29596 3114
rect 29654 3080 29688 3114
rect 29746 3080 29780 3114
rect 29838 3080 29872 3114
rect 29930 3080 29964 3114
rect 30022 3080 30056 3114
rect 30114 3080 30148 3114
rect 30206 3080 30240 3114
rect 30298 3080 30332 3114
rect 25606 2984 25640 3018
rect 25698 2984 25732 3018
rect 25790 2984 25824 3018
rect 25882 2984 25916 3018
rect 25974 2984 26008 3018
rect 26066 2984 26100 3018
rect 26158 2984 26192 3018
rect 26250 2984 26284 3018
rect 26342 2984 26376 3018
rect 26434 2984 26468 3018
rect 26526 2984 26560 3018
rect 26618 2984 26652 3018
rect 26710 2984 26744 3018
rect 26802 2984 26836 3018
rect 26894 2984 26928 3018
rect 26986 2984 27020 3018
rect 27078 2984 27112 3018
rect 27170 2984 27204 3018
rect 27262 2984 27296 3018
rect 27354 2984 27388 3018
rect 27446 2984 27480 3018
rect 27538 2984 27572 3018
rect 27630 2984 27664 3018
rect 27722 2984 27756 3018
rect 27814 2984 27848 3018
rect 27906 2984 27940 3018
rect 27998 2984 28032 3018
rect 28090 2984 28124 3018
rect 28182 2984 28216 3018
rect 28274 2984 28308 3018
rect 28366 2984 28400 3018
rect 28458 2984 28492 3018
rect 28550 2984 28584 3018
rect 28642 2984 28676 3018
rect 28734 2984 28768 3018
rect 28826 2984 28860 3018
rect 28918 2984 28952 3018
rect 29010 2984 29044 3018
rect 29102 2984 29136 3018
rect 29194 2984 29228 3018
rect 29286 2984 29320 3018
rect 29378 2984 29412 3018
rect 29470 2984 29504 3018
rect 29562 2984 29596 3018
rect 29654 2984 29688 3018
rect 29746 2984 29780 3018
rect 29838 2984 29872 3018
rect 29930 2984 29964 3018
rect 30022 2984 30056 3018
rect 30114 2984 30148 3018
rect 30206 2984 30240 3018
rect 30298 2984 30332 3018
rect 25626 2772 25660 2806
rect 25699 2610 25733 2644
rect 25791 2814 25825 2848
rect 25953 2688 25987 2722
rect 26155 2832 26189 2848
rect 26155 2814 26173 2832
rect 26173 2814 26189 2832
rect 26343 2822 26377 2848
rect 26343 2814 26345 2822
rect 26345 2814 26377 2822
rect 26067 2610 26101 2644
rect 26803 2746 26837 2780
rect 26711 2678 26745 2712
rect 26803 2636 26824 2644
rect 26824 2636 26837 2644
rect 26803 2610 26837 2636
rect 27079 2822 27113 2848
rect 27079 2814 27088 2822
rect 27088 2814 27113 2822
rect 27472 2748 27499 2780
rect 27499 2748 27506 2780
rect 27472 2746 27506 2748
rect 27355 2678 27389 2712
rect 28010 2737 28035 2762
rect 28035 2737 28044 2762
rect 28010 2728 28044 2737
rect 27906 2552 27934 2585
rect 27934 2552 27940 2585
rect 27906 2551 27940 2552
rect 28091 2610 28125 2644
rect 28183 2814 28217 2848
rect 28347 2750 28353 2779
rect 28353 2750 28381 2779
rect 28347 2745 28381 2750
rect 28547 2832 28581 2848
rect 28547 2814 28565 2832
rect 28565 2814 28581 2832
rect 28735 2822 28769 2848
rect 28735 2814 28737 2822
rect 28737 2814 28769 2822
rect 28459 2610 28493 2644
rect 29195 2746 29229 2780
rect 29103 2678 29137 2712
rect 29195 2636 29216 2644
rect 29216 2636 29229 2644
rect 29195 2610 29229 2636
rect 29471 2822 29505 2848
rect 29471 2814 29480 2822
rect 29480 2814 29505 2822
rect 29856 2748 29857 2782
rect 29857 2748 29890 2782
rect 29747 2678 29781 2712
rect 30293 2872 30326 2896
rect 30326 2872 30327 2896
rect 30293 2862 30327 2872
rect 25606 2440 25640 2474
rect 25698 2440 25732 2474
rect 25790 2440 25824 2474
rect 25882 2440 25916 2474
rect 25974 2440 26008 2474
rect 26066 2440 26100 2474
rect 26158 2440 26192 2474
rect 26250 2440 26284 2474
rect 26342 2440 26376 2474
rect 26434 2440 26468 2474
rect 26526 2440 26560 2474
rect 26618 2440 26652 2474
rect 26710 2440 26744 2474
rect 26802 2440 26836 2474
rect 26894 2440 26928 2474
rect 26986 2440 27020 2474
rect 27078 2440 27112 2474
rect 27170 2440 27204 2474
rect 27262 2440 27296 2474
rect 27354 2440 27388 2474
rect 27446 2440 27480 2474
rect 27538 2440 27572 2474
rect 27630 2440 27664 2474
rect 27722 2440 27756 2474
rect 27814 2440 27848 2474
rect 27906 2440 27940 2474
rect 27998 2440 28032 2474
rect 28090 2440 28124 2474
rect 28182 2440 28216 2474
rect 28274 2440 28308 2474
rect 28366 2440 28400 2474
rect 28458 2440 28492 2474
rect 28550 2440 28584 2474
rect 28642 2440 28676 2474
rect 28734 2440 28768 2474
rect 28826 2440 28860 2474
rect 28918 2440 28952 2474
rect 29010 2440 29044 2474
rect 29102 2440 29136 2474
rect 29194 2440 29228 2474
rect 29286 2440 29320 2474
rect 29378 2440 29412 2474
rect 29470 2440 29504 2474
rect 29562 2440 29596 2474
rect 29654 2440 29688 2474
rect 29746 2440 29780 2474
rect 29838 2440 29872 2474
rect 29930 2440 29964 2474
rect 30022 2440 30056 2474
rect 30114 2440 30148 2474
rect 30206 2440 30240 2474
rect 30298 2440 30332 2474
rect 25606 2344 25640 2378
rect 25698 2344 25732 2378
rect 25790 2344 25824 2378
rect 25882 2344 25916 2378
rect 25974 2344 26008 2378
rect 26066 2344 26100 2378
rect 26158 2344 26192 2378
rect 26250 2344 26284 2378
rect 26342 2344 26376 2378
rect 26434 2344 26468 2378
rect 26526 2344 26560 2378
rect 26618 2344 26652 2378
rect 26710 2344 26744 2378
rect 26802 2344 26836 2378
rect 26894 2344 26928 2378
rect 26986 2344 27020 2378
rect 27078 2344 27112 2378
rect 27170 2344 27204 2378
rect 27262 2344 27296 2378
rect 27354 2344 27388 2378
rect 27446 2344 27480 2378
rect 27538 2344 27572 2378
rect 27630 2344 27664 2378
rect 27722 2344 27756 2378
rect 27814 2344 27848 2378
rect 27906 2344 27940 2378
rect 27998 2344 28032 2378
rect 28090 2344 28124 2378
rect 28182 2344 28216 2378
rect 28274 2344 28308 2378
rect 28366 2344 28400 2378
rect 28458 2344 28492 2378
rect 28550 2344 28584 2378
rect 28642 2344 28676 2378
rect 28734 2344 28768 2378
rect 28826 2344 28860 2378
rect 28918 2344 28952 2378
rect 29010 2344 29044 2378
rect 29102 2344 29136 2378
rect 29194 2344 29228 2378
rect 29286 2344 29320 2378
rect 29378 2344 29412 2378
rect 29470 2344 29504 2378
rect 29562 2344 29596 2378
rect 29654 2344 29688 2378
rect 29746 2344 29780 2378
rect 29838 2344 29872 2378
rect 29930 2344 29964 2378
rect 30022 2344 30056 2378
rect 30114 2344 30148 2378
rect 30206 2344 30240 2378
rect 30298 2344 30332 2378
rect 25699 2174 25733 2208
rect 25622 2012 25656 2046
rect 25791 1970 25825 2004
rect 26067 2174 26101 2208
rect 25950 2096 25984 2130
rect 26155 1986 26173 2004
rect 26173 1986 26189 2004
rect 26155 1970 26189 1986
rect 26803 2182 26837 2208
rect 26803 2174 26824 2182
rect 26824 2174 26837 2182
rect 26711 2106 26745 2140
rect 26343 1996 26345 2004
rect 26345 1996 26377 2004
rect 26343 1970 26377 1996
rect 26803 2038 26837 2072
rect 27079 1996 27088 2004
rect 27088 1996 27113 2004
rect 27079 1970 27113 1996
rect 27355 2106 27389 2140
rect 27464 2036 27465 2070
rect 27465 2036 27498 2070
rect 27906 2266 27940 2270
rect 27906 2236 27934 2266
rect 27934 2236 27940 2266
rect 28091 2174 28125 2208
rect 28011 2047 28035 2076
rect 28035 2047 28045 2076
rect 28011 2042 28045 2047
rect 28183 1970 28217 2004
rect 28459 2174 28493 2208
rect 28348 2068 28382 2071
rect 28348 2037 28353 2068
rect 28353 2037 28382 2068
rect 28547 1986 28565 2004
rect 28565 1986 28581 2004
rect 28547 1970 28581 1986
rect 29195 2182 29229 2208
rect 29195 2174 29216 2182
rect 29216 2174 29229 2182
rect 29103 2106 29137 2140
rect 28735 1996 28737 2004
rect 28737 1996 28769 2004
rect 28735 1970 28769 1996
rect 29195 2038 29229 2072
rect 29471 1996 29480 2004
rect 29480 1996 29505 2004
rect 29471 1970 29505 1996
rect 29747 2106 29781 2140
rect 29856 2070 29890 2071
rect 29856 2037 29857 2070
rect 29857 2037 29890 2070
rect 30294 1912 30326 1937
rect 30326 1912 30328 1937
rect 30294 1903 30328 1912
rect 25606 1800 25640 1834
rect 25698 1800 25732 1834
rect 25790 1800 25824 1834
rect 25882 1800 25916 1834
rect 25974 1800 26008 1834
rect 26066 1800 26100 1834
rect 26158 1800 26192 1834
rect 26250 1800 26284 1834
rect 26342 1800 26376 1834
rect 26434 1800 26468 1834
rect 26526 1800 26560 1834
rect 26618 1800 26652 1834
rect 26710 1800 26744 1834
rect 26802 1800 26836 1834
rect 26894 1800 26928 1834
rect 26986 1800 27020 1834
rect 27078 1800 27112 1834
rect 27170 1800 27204 1834
rect 27262 1800 27296 1834
rect 27354 1800 27388 1834
rect 27446 1800 27480 1834
rect 27538 1800 27572 1834
rect 27630 1800 27664 1834
rect 27722 1800 27756 1834
rect 27814 1800 27848 1834
rect 27906 1800 27940 1834
rect 27998 1800 28032 1834
rect 28090 1800 28124 1834
rect 28182 1800 28216 1834
rect 28274 1800 28308 1834
rect 28366 1800 28400 1834
rect 28458 1800 28492 1834
rect 28550 1800 28584 1834
rect 28642 1800 28676 1834
rect 28734 1800 28768 1834
rect 28826 1800 28860 1834
rect 28918 1800 28952 1834
rect 29010 1800 29044 1834
rect 29102 1800 29136 1834
rect 29194 1800 29228 1834
rect 29286 1800 29320 1834
rect 29378 1800 29412 1834
rect 29470 1800 29504 1834
rect 29562 1800 29596 1834
rect 29654 1800 29688 1834
rect 29746 1800 29780 1834
rect 29838 1800 29872 1834
rect 29930 1800 29964 1834
rect 30022 1800 30056 1834
rect 30114 1800 30148 1834
rect 30206 1800 30240 1834
rect 30298 1800 30332 1834
rect 8606 1396 8640 1406
rect 8606 1372 8640 1396
rect 8698 1396 8732 1406
rect 8698 1372 8732 1396
rect 8790 1396 8824 1406
rect 8790 1372 8824 1396
rect 8882 1396 8916 1406
rect 8882 1372 8916 1396
rect 8974 1396 9008 1406
rect 8974 1372 9008 1396
rect 9066 1396 9100 1406
rect 9066 1372 9100 1396
rect 9158 1396 9192 1406
rect 9158 1372 9192 1396
rect 9250 1396 9284 1406
rect 9250 1372 9284 1396
rect 9342 1396 9376 1406
rect 9342 1372 9376 1396
rect 9434 1396 9468 1406
rect 9434 1372 9468 1396
rect 9526 1396 9560 1406
rect 9526 1372 9560 1396
rect 9618 1396 9652 1406
rect 9618 1372 9652 1396
rect 9710 1396 9744 1406
rect 9710 1372 9744 1396
rect 9802 1396 9836 1406
rect 9802 1372 9836 1396
rect 9894 1396 9928 1406
rect 9894 1372 9928 1396
rect 9986 1396 10020 1406
rect 9986 1372 10020 1396
rect 10078 1396 10112 1406
rect 10078 1372 10112 1396
rect 10170 1396 10204 1406
rect 10170 1372 10204 1396
rect 10262 1396 10296 1406
rect 10262 1372 10296 1396
rect 10354 1396 10388 1406
rect 10354 1372 10388 1396
rect 10446 1396 10480 1406
rect 10446 1372 10480 1396
rect 10538 1396 10572 1406
rect 10538 1372 10572 1396
rect 10630 1396 10664 1406
rect 10630 1372 10664 1396
rect 10722 1396 10756 1406
rect 10722 1372 10756 1396
rect 10814 1396 10848 1406
rect 10814 1372 10848 1396
rect 10906 1396 10940 1406
rect 10906 1372 10940 1396
rect 10998 1396 11032 1406
rect 10998 1372 11032 1396
rect 11090 1396 11124 1406
rect 11090 1372 11124 1396
rect 11182 1396 11216 1406
rect 11182 1372 11216 1396
rect 11274 1396 11308 1406
rect 11274 1372 11308 1396
rect 11366 1396 11400 1406
rect 11366 1372 11400 1396
rect 12990 1396 13024 1406
rect 12990 1372 13024 1396
rect 13082 1396 13116 1406
rect 13082 1372 13116 1396
rect 13174 1396 13208 1406
rect 13174 1372 13208 1396
rect 13266 1396 13300 1406
rect 13266 1372 13300 1396
rect 13358 1396 13392 1406
rect 13358 1372 13392 1396
rect 13450 1396 13484 1406
rect 13450 1372 13484 1396
rect 13542 1396 13576 1406
rect 13542 1372 13576 1396
rect 13634 1396 13668 1406
rect 13634 1372 13668 1396
rect 13726 1396 13760 1406
rect 13726 1372 13760 1396
rect 13818 1396 13852 1406
rect 13818 1372 13852 1396
rect 13910 1396 13944 1406
rect 13910 1372 13944 1396
rect 14002 1396 14036 1406
rect 14002 1372 14036 1396
rect 14094 1396 14128 1406
rect 14094 1372 14128 1396
rect 14186 1396 14220 1406
rect 14186 1372 14220 1396
rect 14278 1396 14312 1406
rect 14278 1372 14312 1396
rect 14370 1396 14404 1406
rect 14370 1372 14404 1396
rect 14462 1396 14496 1406
rect 14462 1372 14496 1396
rect 14554 1396 14588 1406
rect 14554 1372 14588 1396
rect 14646 1396 14680 1406
rect 14646 1372 14680 1396
rect 14738 1396 14772 1406
rect 14738 1372 14772 1396
rect 14830 1396 14864 1406
rect 14830 1372 14864 1396
rect 14922 1396 14956 1406
rect 14922 1372 14956 1396
rect 15014 1396 15048 1406
rect 15014 1372 15048 1396
rect 15106 1396 15140 1406
rect 15106 1372 15140 1396
rect 15198 1396 15232 1406
rect 15198 1372 15232 1396
rect 15290 1396 15324 1406
rect 15290 1372 15324 1396
rect 15382 1396 15416 1406
rect 15382 1372 15416 1396
rect 15474 1396 15508 1406
rect 15474 1372 15508 1396
rect 15566 1396 15600 1406
rect 15566 1372 15600 1396
rect 15658 1396 15692 1406
rect 15658 1372 15692 1396
rect 15750 1396 15784 1406
rect 15750 1372 15784 1396
rect 8614 1094 8648 1110
rect 8614 1076 8648 1094
rect 11451 1065 11485 1099
rect 12998 1060 13032 1093
rect 12998 1059 13032 1060
rect 15751 1067 15785 1101
rect 8606 838 8640 862
rect 8606 828 8640 838
rect 8698 838 8732 862
rect 8698 828 8732 838
rect 8790 838 8824 862
rect 8790 828 8824 838
rect 8882 838 8916 862
rect 8882 828 8916 838
rect 8974 838 9008 862
rect 8974 828 9008 838
rect 9066 838 9100 862
rect 9066 828 9100 838
rect 9158 838 9192 862
rect 9158 828 9192 838
rect 9250 838 9284 862
rect 9250 828 9284 838
rect 9342 838 9376 862
rect 9342 828 9376 838
rect 9434 838 9468 862
rect 9434 828 9468 838
rect 9526 838 9560 862
rect 9526 828 9560 838
rect 9618 838 9652 862
rect 9618 828 9652 838
rect 9710 838 9744 862
rect 9710 828 9744 838
rect 9802 838 9836 862
rect 9802 828 9836 838
rect 9894 838 9928 862
rect 9894 828 9928 838
rect 9986 838 10020 862
rect 9986 828 10020 838
rect 10078 838 10112 862
rect 10078 828 10112 838
rect 10170 838 10204 862
rect 10170 828 10204 838
rect 10262 838 10296 862
rect 10262 828 10296 838
rect 10354 838 10388 862
rect 10354 828 10388 838
rect 10446 838 10480 862
rect 10446 828 10480 838
rect 10538 838 10572 862
rect 10538 828 10572 838
rect 10630 838 10664 862
rect 10630 828 10664 838
rect 10722 838 10756 862
rect 10722 828 10756 838
rect 10814 838 10848 862
rect 10814 828 10848 838
rect 10906 838 10940 862
rect 10906 828 10940 838
rect 10998 838 11032 862
rect 10998 828 11032 838
rect 11090 838 11124 862
rect 11090 828 11124 838
rect 11182 838 11216 862
rect 11182 828 11216 838
rect 11274 838 11308 862
rect 11274 828 11308 838
rect 11366 838 11400 862
rect 11366 828 11400 838
rect 12990 838 13024 862
rect 12990 828 13024 838
rect 13082 838 13116 862
rect 13082 828 13116 838
rect 13174 838 13208 862
rect 13174 828 13208 838
rect 13266 838 13300 862
rect 13266 828 13300 838
rect 13358 838 13392 862
rect 13358 828 13392 838
rect 13450 838 13484 862
rect 13450 828 13484 838
rect 13542 838 13576 862
rect 13542 828 13576 838
rect 13634 838 13668 862
rect 13634 828 13668 838
rect 13726 838 13760 862
rect 13726 828 13760 838
rect 13818 838 13852 862
rect 13818 828 13852 838
rect 13910 838 13944 862
rect 13910 828 13944 838
rect 14002 838 14036 862
rect 14002 828 14036 838
rect 14094 838 14128 862
rect 14094 828 14128 838
rect 14186 838 14220 862
rect 14186 828 14220 838
rect 14278 838 14312 862
rect 14278 828 14312 838
rect 14370 838 14404 862
rect 14370 828 14404 838
rect 14462 838 14496 862
rect 14462 828 14496 838
rect 14554 838 14588 862
rect 14554 828 14588 838
rect 14646 838 14680 862
rect 14646 828 14680 838
rect 14738 838 14772 862
rect 14738 828 14772 838
rect 14830 838 14864 862
rect 14830 828 14864 838
rect 14922 838 14956 862
rect 14922 828 14956 838
rect 15014 838 15048 862
rect 15014 828 15048 838
rect 15106 838 15140 862
rect 15106 828 15140 838
rect 15198 838 15232 862
rect 15198 828 15232 838
rect 15290 838 15324 862
rect 15290 828 15324 838
rect 15382 838 15416 862
rect 15382 828 15416 838
rect 15474 838 15508 862
rect 15474 828 15508 838
rect 15566 838 15600 862
rect 15566 828 15600 838
rect 15658 838 15692 862
rect 15658 828 15692 838
rect 15750 838 15784 862
rect 15750 828 15784 838
rect 8604 254 8638 264
rect 8604 230 8638 254
rect 8696 254 8730 264
rect 8696 230 8730 254
rect 8788 254 8822 264
rect 8788 230 8822 254
rect 8880 254 8914 264
rect 8880 230 8914 254
rect 8972 254 9006 264
rect 8972 230 9006 254
rect 9064 254 9098 264
rect 9064 230 9098 254
rect 9156 254 9190 264
rect 9156 230 9190 254
rect 9248 254 9282 264
rect 9248 230 9282 254
rect 9340 254 9374 264
rect 9340 230 9374 254
rect 10038 230 10072 264
rect 10130 230 10164 264
rect 10222 230 10256 264
rect 10314 230 10348 264
rect 10406 230 10440 264
rect 10498 230 10532 264
rect 10590 230 10624 264
rect 10682 230 10716 264
rect 10774 230 10808 264
rect 10996 254 11030 264
rect 10996 230 11030 254
rect 11088 254 11122 264
rect 11088 230 11122 254
rect 11180 254 11214 264
rect 11180 230 11214 254
rect 11272 254 11306 264
rect 11272 230 11306 254
rect 11364 254 11398 264
rect 11364 230 11398 254
rect 11456 254 11490 264
rect 11456 230 11490 254
rect 11548 254 11582 264
rect 11548 230 11582 254
rect 11640 254 11674 264
rect 11640 230 11674 254
rect 11732 254 11766 264
rect 11732 230 11766 254
rect 12430 230 12464 264
rect 12522 230 12556 264
rect 12614 230 12648 264
rect 12706 230 12740 264
rect 12798 230 12832 264
rect 12890 230 12924 264
rect 12982 230 13016 264
rect 13074 230 13108 264
rect 13166 230 13200 264
rect 13388 254 13422 264
rect 13388 230 13422 254
rect 13480 254 13514 264
rect 13480 230 13514 254
rect 13572 254 13606 264
rect 13572 230 13606 254
rect 13664 254 13698 264
rect 13664 230 13698 254
rect 13756 254 13790 264
rect 13756 230 13790 254
rect 13848 254 13882 264
rect 13848 230 13882 254
rect 13940 254 13974 264
rect 13940 230 13974 254
rect 14032 254 14066 264
rect 14032 230 14066 254
rect 14124 254 14158 264
rect 14820 254 14854 264
rect 14124 230 14158 254
rect 14820 230 14854 254
rect 14912 254 14946 264
rect 14912 230 14946 254
rect 15004 254 15038 264
rect 15004 230 15038 254
rect 15096 254 15130 264
rect 15096 230 15130 254
rect 15188 254 15222 264
rect 15188 230 15222 254
rect 15280 254 15314 264
rect 15280 230 15314 254
rect 15372 254 15406 264
rect 15372 230 15406 254
rect 15464 254 15498 264
rect 15464 230 15498 254
rect 15556 254 15590 264
rect 15556 230 15590 254
rect 15780 230 15814 264
rect 15872 230 15906 264
rect 15964 230 15998 264
rect 16056 230 16090 264
rect 16148 230 16182 264
rect 16240 230 16274 264
rect 16332 230 16366 264
rect 16424 230 16458 264
rect 16516 230 16550 264
rect 17214 254 17246 264
rect 17246 254 17248 264
rect 17306 254 17338 264
rect 17338 254 17340 264
rect 17398 254 17430 264
rect 17430 254 17432 264
rect 17490 254 17522 264
rect 17522 254 17524 264
rect 17582 254 17614 264
rect 17614 254 17616 264
rect 17674 254 17706 264
rect 17706 254 17708 264
rect 17766 254 17798 264
rect 17798 254 17800 264
rect 17858 254 17890 264
rect 17890 254 17892 264
rect 17950 254 17982 264
rect 17982 254 17984 264
rect 17214 230 17248 254
rect 17306 230 17340 254
rect 17398 230 17432 254
rect 17490 230 17524 254
rect 17582 230 17616 254
rect 17674 230 17708 254
rect 17766 230 17800 254
rect 17858 230 17892 254
rect 17950 230 17984 254
rect 18172 230 18206 264
rect 18264 230 18298 264
rect 18356 230 18390 264
rect 18448 230 18482 264
rect 18540 230 18574 264
rect 18632 230 18666 264
rect 18724 230 18758 264
rect 18816 230 18850 264
rect 18908 230 18942 264
rect 19606 254 19638 264
rect 19638 254 19640 264
rect 19698 254 19730 264
rect 19730 254 19732 264
rect 19790 254 19822 264
rect 19822 254 19824 264
rect 19882 254 19914 264
rect 19914 254 19916 264
rect 19974 254 20006 264
rect 20006 254 20008 264
rect 20066 254 20098 264
rect 20098 254 20100 264
rect 20158 254 20190 264
rect 20190 254 20192 264
rect 20250 254 20282 264
rect 20282 254 20284 264
rect 20342 254 20374 264
rect 20374 254 20376 264
rect 20564 254 20586 264
rect 20586 254 20598 264
rect 20656 254 20678 264
rect 20678 254 20690 264
rect 20748 254 20770 264
rect 20770 254 20782 264
rect 20840 254 20862 264
rect 20862 254 20874 264
rect 20932 254 20954 264
rect 20954 254 20966 264
rect 21024 254 21046 264
rect 21046 254 21058 264
rect 21116 254 21138 264
rect 21138 254 21150 264
rect 21208 254 21230 264
rect 21230 254 21242 264
rect 21300 254 21322 264
rect 21322 254 21334 264
rect 21996 254 22000 264
rect 22000 254 22030 264
rect 22088 254 22092 264
rect 22092 254 22122 264
rect 22180 254 22184 264
rect 22184 254 22214 264
rect 22272 254 22276 264
rect 22276 254 22306 264
rect 22364 254 22368 264
rect 22368 254 22398 264
rect 22456 254 22460 264
rect 22460 254 22490 264
rect 22548 254 22552 264
rect 22552 254 22582 264
rect 22640 254 22644 264
rect 22644 254 22674 264
rect 22732 254 22736 264
rect 22736 254 22766 264
rect 22956 254 22978 264
rect 22978 254 22990 264
rect 23048 254 23070 264
rect 23070 254 23082 264
rect 23140 254 23162 264
rect 23162 254 23174 264
rect 23232 254 23254 264
rect 23254 254 23266 264
rect 23324 254 23346 264
rect 23346 254 23358 264
rect 23416 254 23438 264
rect 23438 254 23450 264
rect 23508 254 23530 264
rect 23530 254 23542 264
rect 23600 254 23622 264
rect 23622 254 23634 264
rect 23692 254 23714 264
rect 23714 254 23726 264
rect 24390 254 24392 264
rect 24392 254 24424 264
rect 24482 254 24484 264
rect 24484 254 24516 264
rect 24574 254 24576 264
rect 24576 254 24608 264
rect 24666 254 24668 264
rect 24668 254 24700 264
rect 24758 254 24760 264
rect 24760 254 24792 264
rect 24850 254 24852 264
rect 24852 254 24884 264
rect 24942 254 24944 264
rect 24944 254 24976 264
rect 25034 254 25036 264
rect 25036 254 25068 264
rect 25126 254 25128 264
rect 25128 254 25160 264
rect 19606 230 19640 254
rect 19698 230 19732 254
rect 19790 230 19824 254
rect 19882 230 19916 254
rect 19974 230 20008 254
rect 20066 230 20100 254
rect 20158 230 20192 254
rect 20250 230 20284 254
rect 20342 230 20376 254
rect 20564 230 20598 254
rect 20656 230 20690 254
rect 20748 230 20782 254
rect 20840 230 20874 254
rect 20932 230 20966 254
rect 21024 230 21058 254
rect 21116 230 21150 254
rect 21208 230 21242 254
rect 21300 230 21334 254
rect 21996 230 22030 254
rect 22088 230 22122 254
rect 22180 230 22214 254
rect 22272 230 22306 254
rect 22364 230 22398 254
rect 22456 230 22490 254
rect 22548 230 22582 254
rect 22640 230 22674 254
rect 22732 230 22766 254
rect 22956 230 22990 254
rect 23048 230 23082 254
rect 23140 230 23174 254
rect 23232 230 23266 254
rect 23324 230 23358 254
rect 23416 230 23450 254
rect 23508 230 23542 254
rect 23600 230 23634 254
rect 23692 230 23726 254
rect 24390 230 24424 254
rect 24482 230 24516 254
rect 24574 230 24608 254
rect 24666 230 24700 254
rect 24758 230 24792 254
rect 24850 230 24884 254
rect 24942 230 24976 254
rect 25034 230 25068 254
rect 25126 230 25160 254
rect 8603 -185 8637 -159
rect 9059 29 9093 42
rect 9059 8 9066 29
rect 9066 8 9093 29
rect 8603 -193 8610 -185
rect 8610 -193 8637 -185
rect 9231 -5 9234 26
rect 9234 -5 9265 26
rect 9231 -8 9265 -5
rect 10141 -5 10144 27
rect 10144 -5 10175 27
rect 10141 -7 10175 -5
rect 10321 29 10355 42
rect 10321 8 10346 29
rect 10346 8 10355 29
rect 10779 -185 10813 -161
rect 10779 -195 10802 -185
rect 10802 -195 10813 -185
rect 10995 -185 11029 -159
rect 11452 29 11486 41
rect 11452 7 11458 29
rect 11458 7 11486 29
rect 10995 -193 11002 -185
rect 11002 -193 11029 -185
rect 11623 -5 11626 25
rect 11626 -5 11657 25
rect 11623 -9 11657 -5
rect 12533 -5 12536 26
rect 12536 -5 12567 26
rect 12533 -8 12567 -5
rect 12713 29 12747 42
rect 12713 8 12738 29
rect 12738 8 12747 29
rect 13173 -185 13207 -161
rect 13173 -195 13194 -185
rect 13194 -195 13207 -185
rect 13387 -185 13421 -159
rect 13844 29 13878 41
rect 13844 7 13850 29
rect 13850 7 13878 29
rect 13387 -193 13394 -185
rect 13394 -193 13421 -185
rect 14014 -5 14018 26
rect 14018 -5 14048 26
rect 14014 -8 14048 -5
rect 14923 -5 14926 26
rect 14926 -5 14957 26
rect 14923 -8 14957 -5
rect 15104 29 15138 43
rect 15104 9 15128 29
rect 15128 9 15138 29
rect 15563 -185 15597 -159
rect 15563 -193 15584 -185
rect 15584 -193 15597 -185
rect 15779 -185 15813 -159
rect 16236 29 16270 42
rect 16236 8 16242 29
rect 16242 8 16270 29
rect 15779 -193 15786 -185
rect 15786 -193 15813 -185
rect 16407 -5 16410 26
rect 16410 -5 16441 26
rect 16407 -8 16441 -5
rect 17317 -5 17320 27
rect 17320 -5 17351 27
rect 17317 -7 17351 -5
rect 17497 29 17531 43
rect 17497 9 17522 29
rect 17522 9 17531 29
rect 17955 -185 17989 -161
rect 17955 -195 17978 -185
rect 17978 -195 17989 -185
rect 18170 -185 18204 -158
rect 18627 29 18661 41
rect 18627 7 18634 29
rect 18634 7 18661 29
rect 18170 -192 18178 -185
rect 18178 -192 18204 -185
rect 18798 -5 18802 27
rect 18802 -5 18832 27
rect 18798 -7 18832 -5
rect 19709 -5 19712 26
rect 19712 -5 19743 26
rect 19709 -8 19743 -5
rect 19890 29 19924 43
rect 19890 9 19914 29
rect 19914 9 19924 29
rect 20347 -185 20381 -159
rect 20347 -193 20370 -185
rect 20370 -193 20381 -185
rect 20562 -185 20596 -159
rect 21019 29 21053 40
rect 21019 6 21026 29
rect 21026 6 21053 29
rect 20562 -193 20570 -185
rect 20570 -193 20596 -185
rect 21190 -5 21194 27
rect 21194 -5 21224 27
rect 21190 -7 21224 -5
rect 22098 -5 22102 26
rect 22102 -5 22132 26
rect 22098 -8 22132 -5
rect 22279 29 22313 43
rect 22279 9 22304 29
rect 22304 9 22313 29
rect 22739 -185 22773 -161
rect 22739 -195 22760 -185
rect 22760 -195 22773 -185
rect 22955 -185 22989 -158
rect 23411 29 23445 41
rect 23411 7 23418 29
rect 23418 7 23445 29
rect 22955 -192 22962 -185
rect 22962 -192 22989 -185
rect 23583 -5 23586 27
rect 23586 -5 23617 27
rect 23583 -7 23617 -5
rect 24493 -5 24496 27
rect 24496 -5 24527 27
rect 24493 -7 24527 -5
rect 24674 29 24708 43
rect 24674 9 24698 29
rect 24698 9 24708 29
rect 25131 -185 25165 -159
rect 25131 -193 25154 -185
rect 25154 -193 25165 -185
rect 8604 -304 8638 -280
rect 8604 -314 8638 -304
rect 8696 -304 8730 -280
rect 8696 -314 8730 -304
rect 8788 -304 8822 -280
rect 8788 -314 8822 -304
rect 8880 -304 8914 -280
rect 8880 -314 8914 -304
rect 8972 -304 9006 -280
rect 8972 -314 9006 -304
rect 9064 -304 9098 -280
rect 9064 -314 9098 -304
rect 9156 -304 9190 -280
rect 9156 -314 9190 -304
rect 9248 -304 9282 -280
rect 9248 -314 9282 -304
rect 9340 -304 9374 -280
rect 9340 -314 9374 -304
rect 10038 -314 10072 -280
rect 10130 -314 10164 -280
rect 10222 -314 10256 -280
rect 10314 -314 10348 -280
rect 10406 -314 10440 -280
rect 10498 -314 10532 -280
rect 10590 -314 10624 -280
rect 10682 -314 10716 -280
rect 10774 -314 10808 -280
rect 10996 -304 11030 -280
rect 10996 -314 11030 -304
rect 11088 -304 11122 -280
rect 11088 -314 11122 -304
rect 11180 -304 11214 -280
rect 11180 -314 11214 -304
rect 11272 -304 11306 -280
rect 11272 -314 11306 -304
rect 11364 -304 11398 -280
rect 11364 -314 11398 -304
rect 11456 -304 11490 -280
rect 11456 -314 11490 -304
rect 11548 -304 11582 -280
rect 11548 -314 11582 -304
rect 11640 -304 11674 -280
rect 11640 -314 11674 -304
rect 11732 -304 11766 -280
rect 11732 -314 11766 -304
rect 12430 -314 12464 -280
rect 12522 -314 12556 -280
rect 12614 -314 12648 -280
rect 12706 -314 12740 -280
rect 12798 -314 12832 -280
rect 12890 -314 12924 -280
rect 12982 -314 13016 -280
rect 13074 -314 13108 -280
rect 13166 -314 13200 -280
rect 13388 -304 13422 -280
rect 13388 -314 13422 -304
rect 13480 -304 13514 -280
rect 13480 -314 13514 -304
rect 13572 -304 13606 -280
rect 13572 -314 13606 -304
rect 13664 -304 13698 -280
rect 13664 -314 13698 -304
rect 13756 -304 13790 -280
rect 13756 -314 13790 -304
rect 13848 -304 13882 -280
rect 13848 -314 13882 -304
rect 13940 -304 13974 -280
rect 13940 -314 13974 -304
rect 14032 -304 14066 -280
rect 14032 -314 14066 -304
rect 14124 -304 14158 -280
rect 14820 -304 14854 -280
rect 14124 -314 14158 -304
rect 14820 -314 14854 -304
rect 14912 -304 14946 -280
rect 14912 -314 14946 -304
rect 15004 -304 15038 -280
rect 15004 -314 15038 -304
rect 15096 -304 15130 -280
rect 15096 -314 15130 -304
rect 15188 -304 15222 -280
rect 15188 -314 15222 -304
rect 15280 -304 15314 -280
rect 15280 -314 15314 -304
rect 15372 -304 15406 -280
rect 15372 -314 15406 -304
rect 15464 -304 15498 -280
rect 15464 -314 15498 -304
rect 15556 -304 15590 -280
rect 15556 -314 15590 -304
rect 15780 -314 15814 -280
rect 15872 -314 15906 -280
rect 15964 -314 15998 -280
rect 16056 -314 16090 -280
rect 16148 -314 16182 -280
rect 16240 -314 16274 -280
rect 16332 -314 16366 -280
rect 16424 -314 16458 -280
rect 16516 -314 16550 -280
rect 17214 -304 17248 -280
rect 17306 -304 17340 -280
rect 17398 -304 17432 -280
rect 17490 -304 17524 -280
rect 17582 -304 17616 -280
rect 17674 -304 17708 -280
rect 17766 -304 17800 -280
rect 17858 -304 17892 -280
rect 17950 -304 17984 -280
rect 17214 -314 17246 -304
rect 17246 -314 17248 -304
rect 17306 -314 17338 -304
rect 17338 -314 17340 -304
rect 17398 -314 17430 -304
rect 17430 -314 17432 -304
rect 17490 -314 17522 -304
rect 17522 -314 17524 -304
rect 17582 -314 17614 -304
rect 17614 -314 17616 -304
rect 17674 -314 17706 -304
rect 17706 -314 17708 -304
rect 17766 -314 17798 -304
rect 17798 -314 17800 -304
rect 17858 -314 17890 -304
rect 17890 -314 17892 -304
rect 17950 -314 17982 -304
rect 17982 -314 17984 -304
rect 18172 -314 18206 -280
rect 18264 -314 18298 -280
rect 18356 -314 18390 -280
rect 18448 -314 18482 -280
rect 18540 -314 18574 -280
rect 18632 -314 18666 -280
rect 18724 -314 18758 -280
rect 18816 -314 18850 -280
rect 18908 -314 18942 -280
rect 19606 -304 19640 -280
rect 19698 -304 19732 -280
rect 19790 -304 19824 -280
rect 19882 -304 19916 -280
rect 19974 -304 20008 -280
rect 20066 -304 20100 -280
rect 20158 -304 20192 -280
rect 20250 -304 20284 -280
rect 20342 -304 20376 -280
rect 20564 -304 20598 -280
rect 20656 -304 20690 -280
rect 20748 -304 20782 -280
rect 20840 -304 20874 -280
rect 20932 -304 20966 -280
rect 21024 -304 21058 -280
rect 21116 -304 21150 -280
rect 21208 -304 21242 -280
rect 21300 -304 21334 -280
rect 21996 -304 22030 -280
rect 22088 -304 22122 -280
rect 22180 -304 22214 -280
rect 22272 -304 22306 -280
rect 22364 -304 22398 -280
rect 22456 -304 22490 -280
rect 22548 -304 22582 -280
rect 22640 -304 22674 -280
rect 22732 -304 22766 -280
rect 22956 -304 22990 -280
rect 23048 -304 23082 -280
rect 23140 -304 23174 -280
rect 23232 -304 23266 -280
rect 23324 -304 23358 -280
rect 23416 -304 23450 -280
rect 23508 -304 23542 -280
rect 23600 -304 23634 -280
rect 23692 -304 23726 -280
rect 24390 -304 24424 -280
rect 24482 -304 24516 -280
rect 24574 -304 24608 -280
rect 24666 -304 24700 -280
rect 24758 -304 24792 -280
rect 24850 -304 24884 -280
rect 24942 -304 24976 -280
rect 25034 -304 25068 -280
rect 25126 -304 25160 -280
rect 19606 -314 19638 -304
rect 19638 -314 19640 -304
rect 19698 -314 19730 -304
rect 19730 -314 19732 -304
rect 19790 -314 19822 -304
rect 19822 -314 19824 -304
rect 19882 -314 19914 -304
rect 19914 -314 19916 -304
rect 19974 -314 20006 -304
rect 20006 -314 20008 -304
rect 20066 -314 20098 -304
rect 20098 -314 20100 -304
rect 20158 -314 20190 -304
rect 20190 -314 20192 -304
rect 20250 -314 20282 -304
rect 20282 -314 20284 -304
rect 20342 -314 20374 -304
rect 20374 -314 20376 -304
rect 20564 -314 20586 -304
rect 20586 -314 20598 -304
rect 20656 -314 20678 -304
rect 20678 -314 20690 -304
rect 20748 -314 20770 -304
rect 20770 -314 20782 -304
rect 20840 -314 20862 -304
rect 20862 -314 20874 -304
rect 20932 -314 20954 -304
rect 20954 -314 20966 -304
rect 21024 -314 21046 -304
rect 21046 -314 21058 -304
rect 21116 -314 21138 -304
rect 21138 -314 21150 -304
rect 21208 -314 21230 -304
rect 21230 -314 21242 -304
rect 21300 -314 21322 -304
rect 21322 -314 21334 -304
rect 21996 -314 22000 -304
rect 22000 -314 22030 -304
rect 22088 -314 22092 -304
rect 22092 -314 22122 -304
rect 22180 -314 22184 -304
rect 22184 -314 22214 -304
rect 22272 -314 22276 -304
rect 22276 -314 22306 -304
rect 22364 -314 22368 -304
rect 22368 -314 22398 -304
rect 22456 -314 22460 -304
rect 22460 -314 22490 -304
rect 22548 -314 22552 -304
rect 22552 -314 22582 -304
rect 22640 -314 22644 -304
rect 22644 -314 22674 -304
rect 22732 -314 22736 -304
rect 22736 -314 22766 -304
rect 22956 -314 22978 -304
rect 22978 -314 22990 -304
rect 23048 -314 23070 -304
rect 23070 -314 23082 -304
rect 23140 -314 23162 -304
rect 23162 -314 23174 -304
rect 23232 -314 23254 -304
rect 23254 -314 23266 -304
rect 23324 -314 23346 -304
rect 23346 -314 23358 -304
rect 23416 -314 23438 -304
rect 23438 -314 23450 -304
rect 23508 -314 23530 -304
rect 23530 -314 23542 -304
rect 23600 -314 23622 -304
rect 23622 -314 23634 -304
rect 23692 -314 23714 -304
rect 23714 -314 23726 -304
rect 24390 -314 24392 -304
rect 24392 -314 24424 -304
rect 24482 -314 24484 -304
rect 24484 -314 24516 -304
rect 24574 -314 24576 -304
rect 24576 -314 24608 -304
rect 24666 -314 24668 -304
rect 24668 -314 24700 -304
rect 24758 -314 24760 -304
rect 24760 -314 24792 -304
rect 24850 -314 24852 -304
rect 24852 -314 24884 -304
rect 24942 -314 24944 -304
rect 24944 -314 24976 -304
rect 25034 -314 25036 -304
rect 25036 -314 25068 -304
rect 25126 -314 25128 -304
rect 25128 -314 25160 -304
rect 8604 -434 8638 -424
rect 8604 -458 8638 -434
rect 8696 -434 8730 -424
rect 8696 -458 8730 -434
rect 8788 -434 8822 -424
rect 8788 -458 8822 -434
rect 8880 -434 8914 -424
rect 8880 -458 8914 -434
rect 8972 -434 9006 -424
rect 8972 -458 9006 -434
rect 9064 -434 9098 -424
rect 9064 -458 9098 -434
rect 9156 -434 9190 -424
rect 9156 -458 9190 -434
rect 9248 -434 9282 -424
rect 9248 -458 9282 -434
rect 9340 -434 9374 -424
rect 9340 -458 9374 -434
rect 9432 -434 9466 -424
rect 9432 -458 9466 -434
rect 9524 -434 9558 -424
rect 9524 -458 9558 -434
rect 9616 -434 9650 -424
rect 9616 -458 9650 -434
rect 9708 -434 9742 -424
rect 9708 -458 9742 -434
rect 9800 -434 9834 -424
rect 9800 -458 9834 -434
rect 9892 -434 9926 -424
rect 9892 -458 9926 -434
rect 9984 -434 10018 -424
rect 9984 -458 10018 -434
rect 10076 -434 10110 -424
rect 10076 -458 10110 -434
rect 10168 -434 10202 -424
rect 10168 -458 10202 -434
rect 10260 -434 10294 -424
rect 10260 -458 10294 -434
rect 10352 -434 10386 -424
rect 10352 -458 10386 -434
rect 10444 -441 10476 -424
rect 10476 -441 10478 -424
rect 10444 -458 10478 -441
rect 10536 -458 10570 -424
rect 10628 -434 10662 -424
rect 10628 -458 10662 -434
rect 10720 -434 10754 -424
rect 10720 -458 10754 -434
rect 10812 -434 10846 -424
rect 10812 -458 10846 -434
rect 10904 -434 10938 -424
rect 10904 -458 10938 -434
rect 10996 -434 11030 -424
rect 10996 -458 11030 -434
rect 11088 -434 11122 -424
rect 11088 -458 11122 -434
rect 11180 -434 11214 -424
rect 11180 -458 11214 -434
rect 11272 -434 11306 -424
rect 11272 -458 11306 -434
rect 11364 -434 11398 -424
rect 11364 -458 11398 -434
rect 11456 -434 11490 -424
rect 11456 -458 11490 -434
rect 11548 -434 11582 -424
rect 11548 -458 11582 -434
rect 11640 -434 11674 -424
rect 11640 -458 11674 -434
rect 11732 -434 11766 -424
rect 11732 -458 11766 -434
rect 11824 -434 11858 -424
rect 11824 -458 11858 -434
rect 11916 -434 11950 -424
rect 11916 -458 11950 -434
rect 12008 -434 12042 -424
rect 12008 -458 12042 -434
rect 12100 -434 12134 -424
rect 12100 -458 12134 -434
rect 12192 -434 12226 -424
rect 12192 -458 12226 -434
rect 12284 -434 12318 -424
rect 12284 -458 12318 -434
rect 12376 -434 12410 -424
rect 12376 -458 12410 -434
rect 12468 -434 12502 -424
rect 12468 -458 12502 -434
rect 12560 -434 12594 -424
rect 12560 -458 12594 -434
rect 12652 -434 12686 -424
rect 12652 -458 12686 -434
rect 12744 -434 12778 -424
rect 12744 -458 12778 -434
rect 12836 -442 12868 -424
rect 12868 -442 12870 -424
rect 12836 -458 12870 -442
rect 12928 -458 12962 -424
rect 13020 -434 13054 -424
rect 13020 -458 13054 -434
rect 13112 -434 13146 -424
rect 13112 -458 13146 -434
rect 13204 -434 13238 -424
rect 13204 -458 13238 -434
rect 13296 -434 13330 -424
rect 13296 -458 13330 -434
rect 13388 -434 13422 -424
rect 13388 -458 13422 -434
rect 13480 -434 13514 -424
rect 13480 -458 13514 -434
rect 13572 -434 13606 -424
rect 13572 -458 13606 -434
rect 13664 -434 13698 -424
rect 13664 -458 13698 -434
rect 13756 -434 13790 -424
rect 13756 -458 13790 -434
rect 13848 -434 13882 -424
rect 13848 -458 13882 -434
rect 13940 -434 13974 -424
rect 13940 -458 13974 -434
rect 14032 -434 14066 -424
rect 14032 -458 14066 -434
rect 14124 -434 14158 -424
rect 14124 -458 14158 -434
rect 14216 -434 14250 -424
rect 14216 -458 14250 -434
rect 14308 -434 14342 -424
rect 14308 -458 14342 -434
rect 14400 -434 14434 -424
rect 14400 -458 14434 -434
rect 14492 -434 14526 -424
rect 14492 -458 14526 -434
rect 14584 -434 14618 -424
rect 14584 -458 14618 -434
rect 14676 -434 14710 -424
rect 14676 -458 14710 -434
rect 14768 -434 14802 -424
rect 14768 -458 14802 -434
rect 14860 -434 14894 -424
rect 14860 -458 14894 -434
rect 14952 -434 14986 -424
rect 14952 -458 14986 -434
rect 15044 -434 15078 -424
rect 15044 -458 15078 -434
rect 15136 -434 15170 -424
rect 15136 -458 15170 -434
rect 15228 -442 15260 -424
rect 15260 -442 15262 -424
rect 15228 -458 15262 -442
rect 15320 -458 15354 -424
rect 15412 -434 15446 -424
rect 15412 -458 15446 -434
rect 15504 -434 15538 -424
rect 15504 -458 15538 -434
rect 15596 -434 15630 -424
rect 15596 -458 15630 -434
rect 15688 -434 15722 -424
rect 15688 -458 15722 -434
rect 15780 -434 15814 -424
rect 15780 -458 15814 -434
rect 15872 -434 15906 -424
rect 15872 -458 15906 -434
rect 15964 -434 15998 -424
rect 15964 -458 15998 -434
rect 16056 -434 16090 -424
rect 16056 -458 16090 -434
rect 16148 -434 16182 -424
rect 16148 -458 16182 -434
rect 16240 -434 16274 -424
rect 16240 -458 16274 -434
rect 16332 -434 16366 -424
rect 16332 -458 16366 -434
rect 16424 -434 16458 -424
rect 16424 -458 16458 -434
rect 16516 -434 16550 -424
rect 16516 -458 16550 -434
rect 16608 -434 16642 -424
rect 16608 -458 16642 -434
rect 16700 -434 16734 -424
rect 16700 -458 16734 -434
rect 16792 -434 16826 -424
rect 16792 -458 16826 -434
rect 16884 -434 16918 -424
rect 16884 -458 16918 -434
rect 16976 -434 17010 -424
rect 16976 -458 17010 -434
rect 17068 -434 17102 -424
rect 17068 -458 17102 -434
rect 17160 -434 17194 -424
rect 17160 -458 17194 -434
rect 17252 -434 17286 -424
rect 17252 -458 17286 -434
rect 17344 -434 17378 -424
rect 17344 -458 17378 -434
rect 17436 -434 17470 -424
rect 17436 -458 17470 -434
rect 17528 -434 17562 -424
rect 17528 -458 17562 -434
rect 17620 -441 17652 -424
rect 17652 -441 17654 -424
rect 17620 -458 17654 -441
rect 17712 -458 17746 -424
rect 17804 -434 17838 -424
rect 17804 -458 17838 -434
rect 17896 -434 17930 -424
rect 17896 -458 17930 -434
rect 17988 -434 18022 -424
rect 17988 -458 18022 -434
rect 18080 -434 18114 -424
rect 18080 -458 18114 -434
rect 18172 -434 18206 -424
rect 18172 -458 18206 -434
rect 18264 -434 18298 -424
rect 18264 -458 18298 -434
rect 18356 -434 18390 -424
rect 18356 -458 18390 -434
rect 18448 -434 18482 -424
rect 18448 -458 18482 -434
rect 18540 -434 18574 -424
rect 18540 -458 18574 -434
rect 18632 -434 18666 -424
rect 18632 -458 18666 -434
rect 18724 -434 18758 -424
rect 18724 -458 18758 -434
rect 18816 -434 18850 -424
rect 18816 -458 18850 -434
rect 18908 -434 18942 -424
rect 18908 -458 18942 -434
rect 19000 -434 19034 -424
rect 19000 -458 19034 -434
rect 19092 -434 19126 -424
rect 19092 -458 19126 -434
rect 19184 -434 19218 -424
rect 19184 -458 19218 -434
rect 19276 -434 19310 -424
rect 19276 -458 19310 -434
rect 19368 -434 19402 -424
rect 19368 -458 19402 -434
rect 19460 -434 19494 -424
rect 19460 -458 19494 -434
rect 19552 -434 19586 -424
rect 19552 -458 19586 -434
rect 19644 -434 19678 -424
rect 19644 -458 19678 -434
rect 19736 -434 19770 -424
rect 19736 -458 19770 -434
rect 19828 -434 19862 -424
rect 19828 -458 19862 -434
rect 19920 -434 19954 -424
rect 19920 -458 19954 -434
rect 20012 -441 20044 -424
rect 20044 -441 20046 -424
rect 20012 -458 20046 -441
rect 20104 -458 20138 -424
rect 20196 -434 20230 -424
rect 20196 -458 20230 -434
rect 20288 -434 20322 -424
rect 20288 -458 20322 -434
rect 20380 -434 20414 -424
rect 20380 -458 20414 -434
rect 20472 -434 20506 -424
rect 20472 -458 20506 -434
rect 20564 -434 20598 -424
rect 20564 -458 20598 -434
rect 20656 -434 20690 -424
rect 20656 -458 20690 -434
rect 20748 -434 20782 -424
rect 20748 -458 20782 -434
rect 20840 -434 20874 -424
rect 20840 -458 20874 -434
rect 20932 -434 20966 -424
rect 20932 -458 20966 -434
rect 21024 -434 21058 -424
rect 21024 -458 21058 -434
rect 21116 -434 21150 -424
rect 21116 -458 21150 -434
rect 21208 -434 21242 -424
rect 21208 -458 21242 -434
rect 21300 -434 21334 -424
rect 21300 -458 21334 -434
rect 21392 -434 21426 -424
rect 21392 -458 21426 -434
rect 21484 -434 21518 -424
rect 21484 -458 21518 -434
rect 21576 -434 21610 -424
rect 21576 -458 21610 -434
rect 21668 -434 21702 -424
rect 21668 -458 21702 -434
rect 21760 -434 21794 -424
rect 21760 -458 21794 -434
rect 21852 -434 21886 -424
rect 21852 -458 21886 -434
rect 21944 -434 21978 -424
rect 21944 -458 21978 -434
rect 22036 -434 22070 -424
rect 22036 -458 22070 -434
rect 22128 -434 22162 -424
rect 22128 -458 22162 -434
rect 22220 -434 22254 -424
rect 22220 -458 22254 -434
rect 22312 -434 22346 -424
rect 22312 -458 22346 -434
rect 22404 -442 22436 -424
rect 22436 -442 22438 -424
rect 22404 -458 22438 -442
rect 22496 -458 22530 -424
rect 22588 -434 22622 -424
rect 22588 -458 22622 -434
rect 22680 -434 22714 -424
rect 22680 -458 22714 -434
rect 22772 -434 22806 -424
rect 22772 -458 22806 -434
rect 22864 -434 22898 -424
rect 22864 -458 22898 -434
rect 22956 -434 22990 -424
rect 22956 -458 22990 -434
rect 23048 -434 23082 -424
rect 23048 -458 23082 -434
rect 23140 -434 23174 -424
rect 23140 -458 23174 -434
rect 23232 -434 23266 -424
rect 23232 -458 23266 -434
rect 23324 -434 23358 -424
rect 23324 -458 23358 -434
rect 23416 -434 23450 -424
rect 23416 -458 23450 -434
rect 23508 -434 23542 -424
rect 23508 -458 23542 -434
rect 23600 -434 23634 -424
rect 23600 -458 23634 -434
rect 23692 -434 23726 -424
rect 23692 -458 23726 -434
rect 23784 -434 23818 -424
rect 23784 -458 23818 -434
rect 23876 -434 23910 -424
rect 23876 -458 23910 -434
rect 23968 -434 24002 -424
rect 23968 -458 24002 -434
rect 24060 -434 24094 -424
rect 24060 -458 24094 -434
rect 24152 -434 24186 -424
rect 24152 -458 24186 -434
rect 24244 -434 24278 -424
rect 24244 -458 24278 -434
rect 24336 -434 24370 -424
rect 24336 -458 24370 -434
rect 24428 -434 24462 -424
rect 24428 -458 24462 -434
rect 24520 -434 24554 -424
rect 24520 -458 24554 -434
rect 24612 -434 24646 -424
rect 24612 -458 24646 -434
rect 24704 -434 24738 -424
rect 24704 -458 24738 -434
rect 24796 -442 24828 -424
rect 24828 -442 24830 -424
rect 24796 -458 24830 -442
rect 24888 -458 24922 -424
rect 24980 -434 25014 -424
rect 24980 -458 25014 -434
rect 25072 -434 25106 -424
rect 25072 -458 25106 -434
rect 25164 -434 25198 -424
rect 25164 -458 25198 -434
rect 25256 -434 25290 -424
rect 25256 -458 25290 -434
rect 8601 -721 8635 -706
rect 8601 -740 8606 -721
rect 8606 -740 8635 -721
rect 8697 -832 8731 -798
rect 8788 -610 8812 -594
rect 8812 -610 8822 -594
rect 8788 -628 8822 -610
rect 9064 -628 9098 -594
rect 8941 -716 8975 -682
rect 9156 -816 9170 -798
rect 9170 -816 9190 -798
rect 9156 -832 9190 -816
rect 9800 -620 9834 -594
rect 9800 -628 9821 -620
rect 9821 -628 9834 -620
rect 9708 -696 9742 -662
rect 9340 -806 9342 -798
rect 9342 -806 9374 -798
rect 9340 -832 9374 -806
rect 9800 -764 9834 -730
rect 10090 -806 10120 -798
rect 10120 -806 10124 -798
rect 10090 -832 10124 -806
rect 10346 -696 10380 -662
rect 10626 -639 10649 -610
rect 10649 -639 10660 -610
rect 10626 -644 10660 -639
rect 10909 -536 10943 -531
rect 10909 -565 10932 -536
rect 10932 -565 10943 -536
rect 10993 -721 11027 -706
rect 10993 -740 10998 -721
rect 10998 -740 11027 -721
rect 11089 -832 11123 -798
rect 11180 -610 11204 -594
rect 11204 -610 11214 -594
rect 11180 -628 11214 -610
rect 11456 -628 11490 -594
rect 11333 -716 11367 -682
rect 11548 -816 11562 -798
rect 11562 -816 11582 -798
rect 11548 -832 11582 -816
rect 12192 -620 12226 -594
rect 12192 -628 12213 -620
rect 12213 -628 12226 -620
rect 12100 -696 12134 -662
rect 11732 -806 11734 -798
rect 11734 -806 11766 -798
rect 11732 -832 11766 -806
rect 12192 -764 12226 -730
rect 12482 -806 12512 -798
rect 12512 -806 12516 -798
rect 12482 -832 12516 -806
rect 12738 -696 12772 -662
rect 13018 -639 13041 -609
rect 13041 -639 13052 -609
rect 13018 -643 13052 -639
rect 13301 -536 13335 -531
rect 13301 -565 13324 -536
rect 13324 -565 13335 -536
rect 13385 -721 13419 -706
rect 13385 -740 13390 -721
rect 13390 -740 13419 -721
rect 13481 -832 13515 -798
rect 13572 -610 13596 -594
rect 13596 -610 13606 -594
rect 13572 -628 13606 -610
rect 13848 -628 13882 -594
rect 13725 -715 13759 -681
rect 13940 -816 13954 -798
rect 13954 -816 13974 -798
rect 13940 -832 13974 -816
rect 14584 -620 14618 -594
rect 14584 -628 14605 -620
rect 14605 -628 14618 -620
rect 14492 -696 14526 -662
rect 14124 -806 14126 -798
rect 14126 -806 14158 -798
rect 14124 -832 14158 -806
rect 14584 -764 14618 -730
rect 14874 -806 14904 -798
rect 14904 -806 14908 -798
rect 14874 -832 14908 -806
rect 15130 -696 15164 -662
rect 15409 -639 15433 -609
rect 15433 -639 15443 -609
rect 15409 -643 15443 -639
rect 15693 -536 15727 -531
rect 15693 -565 15716 -536
rect 15716 -565 15727 -536
rect 15777 -721 15811 -706
rect 15777 -740 15782 -721
rect 15782 -740 15811 -721
rect 15873 -832 15907 -798
rect 15964 -610 15988 -594
rect 15988 -610 15998 -594
rect 15964 -628 15998 -610
rect 16240 -628 16274 -594
rect 16117 -715 16151 -681
rect 16332 -816 16346 -798
rect 16346 -816 16366 -798
rect 16332 -832 16366 -816
rect 16976 -620 17010 -594
rect 16976 -628 16997 -620
rect 16997 -628 17010 -620
rect 16884 -696 16918 -662
rect 16516 -806 16518 -798
rect 16518 -806 16550 -798
rect 16516 -832 16550 -806
rect 16976 -764 17010 -730
rect 17266 -806 17296 -798
rect 17296 -806 17300 -798
rect 17266 -832 17300 -806
rect 17522 -696 17556 -662
rect 17802 -639 17825 -608
rect 17825 -639 17836 -608
rect 17802 -642 17836 -639
rect 18085 -536 18119 -531
rect 18085 -565 18108 -536
rect 18108 -565 18119 -536
rect 18168 -721 18202 -705
rect 18168 -739 18174 -721
rect 18174 -739 18202 -721
rect 18265 -832 18299 -798
rect 18356 -610 18380 -594
rect 18380 -610 18390 -594
rect 18356 -628 18390 -610
rect 18632 -628 18666 -594
rect 18509 -716 18543 -682
rect 18724 -816 18738 -798
rect 18738 -816 18758 -798
rect 18724 -832 18758 -816
rect 19368 -620 19402 -594
rect 19368 -628 19389 -620
rect 19389 -628 19402 -620
rect 19276 -696 19310 -662
rect 18908 -806 18910 -798
rect 18910 -806 18942 -798
rect 18908 -832 18942 -806
rect 19368 -764 19402 -730
rect 19658 -806 19688 -798
rect 19688 -806 19692 -798
rect 19658 -832 19692 -806
rect 19914 -696 19948 -662
rect 20193 -639 20217 -609
rect 20217 -639 20227 -609
rect 20193 -643 20227 -639
rect 20477 -536 20511 -531
rect 20477 -565 20500 -536
rect 20500 -565 20511 -536
rect 20560 -721 20594 -706
rect 20560 -740 20566 -721
rect 20566 -740 20594 -721
rect 20657 -832 20691 -798
rect 20748 -610 20772 -594
rect 20772 -610 20782 -594
rect 20748 -628 20782 -610
rect 21024 -628 21058 -594
rect 20901 -715 20935 -681
rect 21116 -816 21130 -798
rect 21130 -816 21150 -798
rect 21116 -832 21150 -816
rect 21760 -620 21794 -594
rect 21760 -628 21781 -620
rect 21781 -628 21794 -620
rect 21668 -696 21702 -662
rect 21300 -806 21302 -798
rect 21302 -806 21334 -798
rect 21300 -832 21334 -806
rect 21760 -764 21794 -730
rect 22050 -806 22080 -798
rect 22080 -806 22084 -798
rect 22050 -832 22084 -806
rect 22306 -696 22340 -662
rect 22586 -639 22609 -610
rect 22609 -639 22620 -610
rect 22586 -644 22620 -639
rect 22869 -536 22903 -531
rect 22869 -565 22892 -536
rect 22892 -565 22903 -536
rect 22953 -721 22987 -705
rect 22953 -739 22958 -721
rect 22958 -739 22987 -721
rect 23049 -832 23083 -798
rect 23140 -610 23164 -594
rect 23164 -610 23174 -594
rect 23140 -628 23174 -610
rect 23416 -628 23450 -594
rect 23294 -716 23328 -682
rect 23508 -816 23522 -798
rect 23522 -816 23542 -798
rect 23508 -832 23542 -816
rect 24152 -620 24186 -594
rect 24152 -628 24173 -620
rect 24173 -628 24186 -620
rect 24060 -696 24094 -662
rect 23692 -806 23694 -798
rect 23694 -806 23726 -798
rect 23692 -832 23726 -806
rect 24152 -764 24186 -730
rect 24442 -806 24472 -798
rect 24472 -806 24476 -798
rect 24442 -832 24476 -806
rect 24698 -696 24732 -662
rect 24979 -639 25001 -608
rect 25001 -639 25013 -608
rect 24979 -642 25013 -639
rect 25261 -536 25295 -531
rect 25261 -565 25284 -536
rect 25284 -565 25295 -536
rect 8604 -992 8638 -968
rect 8604 -1002 8638 -992
rect 8696 -992 8730 -968
rect 8696 -1002 8730 -992
rect 8788 -992 8822 -968
rect 8788 -1002 8822 -992
rect 8880 -992 8914 -968
rect 8880 -1002 8914 -992
rect 8972 -992 9006 -968
rect 8972 -1002 9006 -992
rect 9064 -992 9098 -968
rect 9064 -1002 9098 -992
rect 9156 -992 9190 -968
rect 9156 -1002 9190 -992
rect 9248 -992 9282 -968
rect 9248 -1002 9282 -992
rect 9340 -992 9374 -968
rect 9340 -1002 9374 -992
rect 9432 -992 9466 -968
rect 9432 -1002 9466 -992
rect 9524 -992 9558 -968
rect 9524 -1002 9558 -992
rect 9616 -992 9650 -968
rect 9616 -1002 9650 -992
rect 9708 -992 9742 -968
rect 9708 -1002 9742 -992
rect 9800 -992 9834 -968
rect 9800 -1002 9834 -992
rect 9892 -992 9926 -968
rect 9892 -1002 9926 -992
rect 9984 -992 10018 -968
rect 9984 -1002 10018 -992
rect 10076 -992 10110 -968
rect 10076 -1002 10110 -992
rect 10168 -992 10202 -968
rect 10168 -1002 10202 -992
rect 10260 -992 10294 -968
rect 10260 -1002 10294 -992
rect 10352 -992 10386 -968
rect 10352 -1002 10386 -992
rect 10444 -992 10478 -968
rect 10444 -1002 10478 -992
rect 10536 -992 10570 -968
rect 10536 -1002 10570 -992
rect 10628 -992 10662 -968
rect 10628 -1002 10662 -992
rect 10720 -992 10754 -968
rect 10720 -1002 10754 -992
rect 10812 -992 10846 -968
rect 10812 -1002 10846 -992
rect 10904 -992 10938 -968
rect 10904 -1002 10938 -992
rect 10996 -992 11030 -968
rect 10996 -1002 11030 -992
rect 11088 -992 11122 -968
rect 11088 -1002 11122 -992
rect 11180 -992 11214 -968
rect 11180 -1002 11214 -992
rect 11272 -992 11306 -968
rect 11272 -1002 11306 -992
rect 11364 -992 11398 -968
rect 11364 -1002 11398 -992
rect 11456 -992 11490 -968
rect 11456 -1002 11490 -992
rect 11548 -992 11582 -968
rect 11548 -1002 11582 -992
rect 11640 -992 11674 -968
rect 11640 -1002 11674 -992
rect 11732 -992 11766 -968
rect 11732 -1002 11766 -992
rect 11824 -992 11858 -968
rect 11824 -1002 11858 -992
rect 11916 -992 11950 -968
rect 11916 -1002 11950 -992
rect 12008 -992 12042 -968
rect 12008 -1002 12042 -992
rect 12100 -992 12134 -968
rect 12100 -1002 12134 -992
rect 12192 -992 12226 -968
rect 12192 -1002 12226 -992
rect 12284 -992 12318 -968
rect 12284 -1002 12318 -992
rect 12376 -992 12410 -968
rect 12376 -1002 12410 -992
rect 12468 -992 12502 -968
rect 12468 -1002 12502 -992
rect 12560 -992 12594 -968
rect 12560 -1002 12594 -992
rect 12652 -992 12686 -968
rect 12652 -1002 12686 -992
rect 12744 -992 12778 -968
rect 12744 -1002 12778 -992
rect 12836 -992 12870 -968
rect 12836 -1002 12870 -992
rect 12928 -992 12962 -968
rect 12928 -1002 12962 -992
rect 13020 -992 13054 -968
rect 13020 -1002 13054 -992
rect 13112 -992 13146 -968
rect 13112 -1002 13146 -992
rect 13204 -992 13238 -968
rect 13204 -1002 13238 -992
rect 13296 -992 13330 -968
rect 13296 -1002 13330 -992
rect 13388 -992 13422 -968
rect 13388 -1002 13422 -992
rect 13480 -992 13514 -968
rect 13480 -1002 13514 -992
rect 13572 -992 13606 -968
rect 13572 -1002 13606 -992
rect 13664 -992 13698 -968
rect 13664 -1002 13698 -992
rect 13756 -992 13790 -968
rect 13756 -1002 13790 -992
rect 13848 -992 13882 -968
rect 13848 -1002 13882 -992
rect 13940 -992 13974 -968
rect 13940 -1002 13974 -992
rect 14032 -992 14066 -968
rect 14032 -1002 14066 -992
rect 14124 -992 14158 -968
rect 14124 -1002 14158 -992
rect 14216 -992 14250 -968
rect 14216 -1002 14250 -992
rect 14308 -992 14342 -968
rect 14308 -1002 14342 -992
rect 14400 -992 14434 -968
rect 14400 -1002 14434 -992
rect 14492 -992 14526 -968
rect 14492 -1002 14526 -992
rect 14584 -992 14618 -968
rect 14584 -1002 14618 -992
rect 14676 -992 14710 -968
rect 14676 -1002 14710 -992
rect 14768 -992 14802 -968
rect 14768 -1002 14802 -992
rect 14860 -992 14894 -968
rect 14860 -1002 14894 -992
rect 14952 -992 14986 -968
rect 14952 -1002 14986 -992
rect 15044 -992 15078 -968
rect 15044 -1002 15078 -992
rect 15136 -992 15170 -968
rect 15136 -1002 15170 -992
rect 15228 -992 15262 -968
rect 15228 -1002 15262 -992
rect 15320 -992 15354 -968
rect 15320 -1002 15354 -992
rect 15412 -992 15446 -968
rect 15412 -1002 15446 -992
rect 15504 -992 15538 -968
rect 15504 -1002 15538 -992
rect 15596 -992 15630 -968
rect 15596 -1002 15630 -992
rect 15688 -992 15722 -968
rect 15688 -1002 15722 -992
rect 15780 -992 15814 -968
rect 15780 -1002 15814 -992
rect 15872 -992 15906 -968
rect 15872 -1002 15906 -992
rect 15964 -992 15998 -968
rect 15964 -1002 15998 -992
rect 16056 -992 16090 -968
rect 16056 -1002 16090 -992
rect 16148 -992 16182 -968
rect 16148 -1002 16182 -992
rect 16240 -992 16274 -968
rect 16240 -1002 16274 -992
rect 16332 -992 16366 -968
rect 16332 -1002 16366 -992
rect 16424 -992 16458 -968
rect 16424 -1002 16458 -992
rect 16516 -992 16550 -968
rect 16516 -1002 16550 -992
rect 16608 -992 16642 -968
rect 16608 -1002 16642 -992
rect 16700 -992 16734 -968
rect 16700 -1002 16734 -992
rect 16792 -992 16826 -968
rect 16792 -1002 16826 -992
rect 16884 -992 16918 -968
rect 16884 -1002 16918 -992
rect 16976 -992 17010 -968
rect 16976 -1002 17010 -992
rect 17068 -992 17102 -968
rect 17068 -1002 17102 -992
rect 17160 -992 17194 -968
rect 17160 -1002 17194 -992
rect 17252 -992 17286 -968
rect 17252 -1002 17286 -992
rect 17344 -992 17378 -968
rect 17344 -1002 17378 -992
rect 17436 -992 17470 -968
rect 17436 -1002 17470 -992
rect 17528 -992 17562 -968
rect 17528 -1002 17562 -992
rect 17620 -992 17654 -968
rect 17620 -1002 17654 -992
rect 17712 -992 17746 -968
rect 17712 -1002 17746 -992
rect 17804 -992 17838 -968
rect 17804 -1002 17838 -992
rect 17896 -992 17930 -968
rect 17896 -1002 17930 -992
rect 17988 -992 18022 -968
rect 17988 -1002 18022 -992
rect 18080 -992 18114 -968
rect 18080 -1002 18114 -992
rect 18172 -992 18206 -968
rect 18172 -1002 18206 -992
rect 18264 -992 18298 -968
rect 18264 -1002 18298 -992
rect 18356 -992 18390 -968
rect 18356 -1002 18390 -992
rect 18448 -992 18482 -968
rect 18448 -1002 18482 -992
rect 18540 -992 18574 -968
rect 18540 -1002 18574 -992
rect 18632 -992 18666 -968
rect 18632 -1002 18666 -992
rect 18724 -992 18758 -968
rect 18724 -1002 18758 -992
rect 18816 -992 18850 -968
rect 18816 -1002 18850 -992
rect 18908 -992 18942 -968
rect 18908 -1002 18942 -992
rect 19000 -992 19034 -968
rect 19000 -1002 19034 -992
rect 19092 -992 19126 -968
rect 19092 -1002 19126 -992
rect 19184 -992 19218 -968
rect 19184 -1002 19218 -992
rect 19276 -992 19310 -968
rect 19276 -1002 19310 -992
rect 19368 -992 19402 -968
rect 19368 -1002 19402 -992
rect 19460 -992 19494 -968
rect 19460 -1002 19494 -992
rect 19552 -992 19586 -968
rect 19552 -1002 19586 -992
rect 19644 -992 19678 -968
rect 19644 -1002 19678 -992
rect 19736 -992 19770 -968
rect 19736 -1002 19770 -992
rect 19828 -992 19862 -968
rect 19828 -1002 19862 -992
rect 19920 -992 19954 -968
rect 19920 -1002 19954 -992
rect 20012 -992 20046 -968
rect 20012 -1002 20046 -992
rect 20104 -992 20138 -968
rect 20104 -1002 20138 -992
rect 20196 -992 20230 -968
rect 20196 -1002 20230 -992
rect 20288 -992 20322 -968
rect 20288 -1002 20322 -992
rect 20380 -992 20414 -968
rect 20380 -1002 20414 -992
rect 20472 -992 20506 -968
rect 20472 -1002 20506 -992
rect 20564 -992 20598 -968
rect 20564 -1002 20598 -992
rect 20656 -992 20690 -968
rect 20656 -1002 20690 -992
rect 20748 -992 20782 -968
rect 20748 -1002 20782 -992
rect 20840 -992 20874 -968
rect 20840 -1002 20874 -992
rect 20932 -992 20966 -968
rect 20932 -1002 20966 -992
rect 21024 -992 21058 -968
rect 21024 -1002 21058 -992
rect 21116 -992 21150 -968
rect 21116 -1002 21150 -992
rect 21208 -992 21242 -968
rect 21208 -1002 21242 -992
rect 21300 -992 21334 -968
rect 21300 -1002 21334 -992
rect 21392 -992 21426 -968
rect 21392 -1002 21426 -992
rect 21484 -992 21518 -968
rect 21484 -1002 21518 -992
rect 21576 -992 21610 -968
rect 21576 -1002 21610 -992
rect 21668 -992 21702 -968
rect 21668 -1002 21702 -992
rect 21760 -992 21794 -968
rect 21760 -1002 21794 -992
rect 21852 -992 21886 -968
rect 21852 -1002 21886 -992
rect 21944 -992 21978 -968
rect 21944 -1002 21978 -992
rect 22036 -992 22070 -968
rect 22036 -1002 22070 -992
rect 22128 -992 22162 -968
rect 22128 -1002 22162 -992
rect 22220 -992 22254 -968
rect 22220 -1002 22254 -992
rect 22312 -992 22346 -968
rect 22312 -1002 22346 -992
rect 22404 -992 22438 -968
rect 22404 -1002 22438 -992
rect 22496 -992 22530 -968
rect 22496 -1002 22530 -992
rect 22588 -992 22622 -968
rect 22588 -1002 22622 -992
rect 22680 -992 22714 -968
rect 22680 -1002 22714 -992
rect 22772 -992 22806 -968
rect 22772 -1002 22806 -992
rect 22864 -992 22898 -968
rect 22864 -1002 22898 -992
rect 22956 -992 22990 -968
rect 22956 -1002 22990 -992
rect 23048 -992 23082 -968
rect 23048 -1002 23082 -992
rect 23140 -992 23174 -968
rect 23140 -1002 23174 -992
rect 23232 -992 23266 -968
rect 23232 -1002 23266 -992
rect 23324 -992 23358 -968
rect 23324 -1002 23358 -992
rect 23416 -992 23450 -968
rect 23416 -1002 23450 -992
rect 23508 -992 23542 -968
rect 23508 -1002 23542 -992
rect 23600 -992 23634 -968
rect 23600 -1002 23634 -992
rect 23692 -992 23726 -968
rect 23692 -1002 23726 -992
rect 23784 -992 23818 -968
rect 23784 -1002 23818 -992
rect 23876 -992 23910 -968
rect 23876 -1002 23910 -992
rect 23968 -992 24002 -968
rect 23968 -1002 24002 -992
rect 24060 -992 24094 -968
rect 24060 -1002 24094 -992
rect 24152 -992 24186 -968
rect 24152 -1002 24186 -992
rect 24244 -992 24278 -968
rect 24244 -1002 24278 -992
rect 24336 -992 24370 -968
rect 24336 -1002 24370 -992
rect 24428 -992 24462 -968
rect 24428 -1002 24462 -992
rect 24520 -992 24554 -968
rect 24520 -1002 24554 -992
rect 24612 -992 24646 -968
rect 24612 -1002 24646 -992
rect 24704 -992 24738 -968
rect 24704 -1002 24738 -992
rect 24796 -992 24830 -968
rect 24796 -1002 24830 -992
rect 24888 -992 24922 -968
rect 24888 -1002 24922 -992
rect 24980 -992 25014 -968
rect 24980 -1002 25014 -992
rect 25072 -992 25106 -968
rect 25072 -1002 25106 -992
rect 25164 -992 25198 -968
rect 25164 -1002 25198 -992
rect 25256 -992 25290 -968
rect 25256 -1002 25290 -992
rect 8604 -1123 8638 -1113
rect 8604 -1147 8638 -1123
rect 8696 -1123 8730 -1113
rect 8696 -1147 8730 -1123
rect 8788 -1123 8822 -1113
rect 8788 -1147 8822 -1123
rect 8880 -1123 8914 -1113
rect 8972 -1123 9003 -1113
rect 9003 -1123 9006 -1113
rect 8880 -1147 8914 -1123
rect 8972 -1147 9006 -1123
rect 9064 -1123 9071 -1113
rect 9071 -1123 9098 -1113
rect 9156 -1123 9190 -1113
rect 9064 -1147 9098 -1123
rect 9156 -1147 9190 -1123
rect 9248 -1123 9282 -1113
rect 9248 -1147 9282 -1123
rect 9340 -1123 9374 -1113
rect 9340 -1147 9374 -1123
rect 9432 -1123 9466 -1113
rect 9432 -1147 9466 -1123
rect 9524 -1123 9558 -1113
rect 9524 -1147 9558 -1123
rect 9616 -1123 9650 -1113
rect 9616 -1147 9650 -1123
rect 9708 -1123 9742 -1113
rect 9708 -1147 9742 -1123
rect 9800 -1123 9834 -1113
rect 9800 -1147 9834 -1123
rect 9892 -1123 9926 -1113
rect 9892 -1147 9926 -1123
rect 9984 -1123 10018 -1113
rect 9984 -1147 10018 -1123
rect 10076 -1123 10110 -1113
rect 10076 -1147 10110 -1123
rect 10168 -1127 10182 -1113
rect 10182 -1127 10202 -1113
rect 10168 -1147 10202 -1127
rect 10260 -1147 10294 -1113
rect 10352 -1123 10386 -1113
rect 10352 -1147 10386 -1123
rect 10444 -1123 10478 -1113
rect 10444 -1147 10478 -1123
rect 10536 -1123 10570 -1113
rect 10536 -1147 10570 -1123
rect 10628 -1123 10662 -1113
rect 10628 -1147 10662 -1123
rect 10720 -1123 10754 -1113
rect 10720 -1147 10754 -1123
rect 10812 -1123 10846 -1113
rect 10812 -1147 10846 -1123
rect 10904 -1123 10938 -1113
rect 10904 -1147 10938 -1123
rect 10996 -1123 11030 -1113
rect 10996 -1147 11030 -1123
rect 11088 -1123 11122 -1113
rect 11088 -1147 11122 -1123
rect 11180 -1123 11214 -1113
rect 11180 -1147 11214 -1123
rect 11272 -1123 11306 -1113
rect 11272 -1147 11306 -1123
rect 11364 -1123 11366 -1113
rect 11366 -1123 11398 -1113
rect 11456 -1123 11457 -1113
rect 11457 -1123 11490 -1113
rect 11548 -1123 11582 -1113
rect 11364 -1147 11398 -1123
rect 11456 -1147 11490 -1123
rect 11548 -1147 11582 -1123
rect 11640 -1123 11674 -1113
rect 11640 -1147 11674 -1123
rect 11732 -1123 11766 -1113
rect 11732 -1147 11766 -1123
rect 11824 -1123 11858 -1113
rect 11824 -1147 11858 -1123
rect 11916 -1123 11950 -1113
rect 11916 -1147 11950 -1123
rect 12008 -1123 12042 -1113
rect 12008 -1147 12042 -1123
rect 12100 -1123 12134 -1113
rect 12100 -1147 12134 -1123
rect 12192 -1123 12226 -1113
rect 12192 -1147 12226 -1123
rect 12284 -1123 12318 -1113
rect 12284 -1147 12318 -1123
rect 12376 -1123 12410 -1113
rect 12376 -1147 12410 -1123
rect 12468 -1123 12502 -1113
rect 12468 -1147 12502 -1123
rect 12560 -1127 12574 -1113
rect 12574 -1127 12594 -1113
rect 12560 -1147 12594 -1127
rect 12652 -1147 12686 -1113
rect 12744 -1123 12778 -1113
rect 12744 -1147 12778 -1123
rect 12836 -1123 12870 -1113
rect 12836 -1147 12870 -1123
rect 12928 -1123 12962 -1113
rect 12928 -1147 12962 -1123
rect 13020 -1123 13054 -1113
rect 13020 -1147 13054 -1123
rect 13112 -1123 13146 -1113
rect 13112 -1147 13146 -1123
rect 13204 -1123 13238 -1113
rect 13204 -1147 13238 -1123
rect 13296 -1123 13330 -1113
rect 13296 -1147 13330 -1123
rect 13388 -1123 13422 -1113
rect 13388 -1147 13422 -1123
rect 13480 -1123 13514 -1113
rect 13480 -1147 13514 -1123
rect 13572 -1123 13606 -1113
rect 13572 -1147 13606 -1123
rect 13664 -1123 13698 -1113
rect 13756 -1123 13788 -1113
rect 13788 -1123 13790 -1113
rect 13664 -1147 13698 -1123
rect 13756 -1147 13790 -1123
rect 13848 -1123 13882 -1113
rect 13848 -1147 13882 -1123
rect 13940 -1123 13974 -1113
rect 13940 -1147 13974 -1123
rect 14032 -1123 14066 -1113
rect 14032 -1147 14066 -1123
rect 14124 -1123 14158 -1113
rect 14124 -1147 14158 -1123
rect 14216 -1123 14250 -1113
rect 14216 -1147 14250 -1123
rect 14308 -1123 14342 -1113
rect 14308 -1147 14342 -1123
rect 14400 -1123 14434 -1113
rect 14400 -1147 14434 -1123
rect 14492 -1123 14526 -1113
rect 14492 -1147 14526 -1123
rect 14584 -1123 14618 -1113
rect 14584 -1147 14618 -1123
rect 14676 -1123 14710 -1113
rect 14676 -1147 14710 -1123
rect 14768 -1123 14802 -1113
rect 14768 -1147 14802 -1123
rect 14860 -1123 14894 -1113
rect 14860 -1147 14894 -1123
rect 14952 -1127 14966 -1113
rect 14966 -1127 14986 -1113
rect 14952 -1147 14986 -1127
rect 15044 -1147 15078 -1113
rect 15136 -1123 15170 -1113
rect 15136 -1147 15170 -1123
rect 15228 -1123 15262 -1113
rect 15228 -1147 15262 -1123
rect 15320 -1123 15354 -1113
rect 15320 -1147 15354 -1123
rect 15412 -1123 15446 -1113
rect 15412 -1147 15446 -1123
rect 15504 -1123 15538 -1113
rect 15504 -1147 15538 -1123
rect 15596 -1123 15630 -1113
rect 15596 -1147 15630 -1123
rect 15688 -1123 15722 -1113
rect 15688 -1147 15722 -1123
rect 15780 -1123 15814 -1113
rect 15780 -1147 15814 -1123
rect 15872 -1123 15906 -1113
rect 15872 -1147 15906 -1123
rect 15964 -1123 15998 -1113
rect 15964 -1147 15998 -1123
rect 16056 -1123 16090 -1113
rect 16056 -1147 16090 -1123
rect 16148 -1123 16149 -1113
rect 16149 -1123 16182 -1113
rect 16240 -1123 16274 -1113
rect 16148 -1147 16182 -1123
rect 16240 -1147 16274 -1123
rect 16332 -1123 16366 -1113
rect 16332 -1147 16366 -1123
rect 16424 -1123 16458 -1113
rect 16424 -1147 16458 -1123
rect 16516 -1123 16550 -1113
rect 16516 -1147 16550 -1123
rect 16608 -1123 16642 -1113
rect 16608 -1147 16642 -1123
rect 16700 -1123 16734 -1113
rect 16700 -1147 16734 -1123
rect 16792 -1123 16826 -1113
rect 16792 -1147 16826 -1123
rect 16884 -1123 16918 -1113
rect 16884 -1147 16918 -1123
rect 16976 -1123 17010 -1113
rect 16976 -1147 17010 -1123
rect 17068 -1123 17102 -1113
rect 17068 -1147 17102 -1123
rect 17160 -1123 17194 -1113
rect 17160 -1147 17194 -1123
rect 17252 -1123 17286 -1113
rect 17252 -1147 17286 -1123
rect 17344 -1127 17358 -1113
rect 17358 -1127 17378 -1113
rect 17344 -1147 17378 -1127
rect 17436 -1147 17470 -1113
rect 17528 -1123 17562 -1113
rect 17528 -1147 17562 -1123
rect 17620 -1123 17654 -1113
rect 17620 -1147 17654 -1123
rect 17712 -1123 17746 -1113
rect 17712 -1147 17746 -1123
rect 17804 -1123 17838 -1113
rect 17804 -1147 17838 -1123
rect 17896 -1123 17930 -1113
rect 17896 -1147 17930 -1123
rect 17988 -1123 18022 -1113
rect 17988 -1147 18022 -1123
rect 18080 -1123 18114 -1113
rect 18080 -1147 18114 -1123
rect 18172 -1123 18206 -1113
rect 18172 -1147 18206 -1123
rect 18264 -1123 18298 -1113
rect 18264 -1147 18298 -1123
rect 18356 -1123 18390 -1113
rect 18356 -1147 18390 -1123
rect 18448 -1123 18482 -1113
rect 18540 -1123 18572 -1113
rect 18572 -1123 18574 -1113
rect 18448 -1147 18482 -1123
rect 18540 -1147 18574 -1123
rect 18632 -1123 18633 -1113
rect 18633 -1123 18666 -1113
rect 18724 -1123 18758 -1113
rect 18632 -1147 18666 -1123
rect 18724 -1147 18758 -1123
rect 18816 -1123 18850 -1113
rect 18816 -1147 18850 -1123
rect 18908 -1123 18942 -1113
rect 18908 -1147 18942 -1123
rect 19000 -1123 19034 -1113
rect 19000 -1147 19034 -1123
rect 19092 -1123 19126 -1113
rect 19092 -1147 19126 -1123
rect 19184 -1123 19218 -1113
rect 19184 -1147 19218 -1123
rect 19276 -1123 19310 -1113
rect 19276 -1147 19310 -1123
rect 19368 -1123 19402 -1113
rect 19368 -1147 19402 -1123
rect 19460 -1123 19494 -1113
rect 19460 -1147 19494 -1123
rect 19552 -1123 19586 -1113
rect 19552 -1147 19586 -1123
rect 19644 -1123 19678 -1113
rect 19644 -1147 19678 -1123
rect 19736 -1127 19750 -1113
rect 19750 -1127 19770 -1113
rect 19736 -1147 19770 -1127
rect 19828 -1147 19862 -1113
rect 19920 -1123 19954 -1113
rect 19920 -1147 19954 -1123
rect 20012 -1123 20046 -1113
rect 20012 -1147 20046 -1123
rect 20104 -1123 20138 -1113
rect 20104 -1147 20138 -1123
rect 20196 -1123 20230 -1113
rect 20196 -1147 20230 -1123
rect 20288 -1123 20322 -1113
rect 20288 -1147 20322 -1123
rect 20380 -1123 20414 -1113
rect 20380 -1147 20414 -1123
rect 20472 -1123 20506 -1113
rect 20472 -1147 20506 -1123
rect 20564 -1123 20598 -1113
rect 20564 -1147 20598 -1123
rect 20656 -1123 20690 -1113
rect 20656 -1147 20690 -1123
rect 20748 -1123 20782 -1113
rect 20748 -1147 20782 -1123
rect 20840 -1123 20874 -1113
rect 20840 -1147 20874 -1123
rect 20932 -1123 20966 -1113
rect 21024 -1123 21057 -1113
rect 21057 -1123 21058 -1113
rect 20932 -1147 20966 -1123
rect 21024 -1147 21058 -1123
rect 21116 -1123 21150 -1113
rect 21116 -1147 21150 -1123
rect 21208 -1123 21242 -1113
rect 21208 -1147 21242 -1123
rect 21300 -1123 21334 -1113
rect 21300 -1147 21334 -1123
rect 21392 -1123 21426 -1113
rect 21392 -1147 21426 -1123
rect 21484 -1123 21518 -1113
rect 21484 -1147 21518 -1123
rect 21576 -1123 21610 -1113
rect 21576 -1147 21610 -1123
rect 21668 -1123 21702 -1113
rect 21668 -1147 21702 -1123
rect 21760 -1123 21794 -1113
rect 21760 -1147 21794 -1123
rect 21852 -1123 21886 -1113
rect 21852 -1147 21886 -1123
rect 21944 -1123 21978 -1113
rect 21944 -1147 21978 -1123
rect 22036 -1123 22070 -1113
rect 22036 -1147 22070 -1123
rect 22128 -1127 22142 -1113
rect 22142 -1127 22162 -1113
rect 22128 -1147 22162 -1127
rect 22220 -1147 22254 -1113
rect 22312 -1123 22346 -1113
rect 22312 -1147 22346 -1123
rect 22404 -1123 22438 -1113
rect 22404 -1147 22438 -1123
rect 22496 -1123 22530 -1113
rect 22496 -1147 22530 -1123
rect 22588 -1123 22622 -1113
rect 22588 -1147 22622 -1123
rect 22680 -1123 22714 -1113
rect 22680 -1147 22714 -1123
rect 22772 -1123 22806 -1113
rect 22772 -1147 22806 -1123
rect 22864 -1123 22898 -1113
rect 22864 -1147 22898 -1123
rect 22956 -1123 22990 -1113
rect 22956 -1147 22990 -1123
rect 23048 -1123 23082 -1113
rect 23048 -1147 23082 -1123
rect 23140 -1123 23174 -1113
rect 23140 -1147 23174 -1123
rect 23232 -1123 23266 -1113
rect 23324 -1123 23357 -1113
rect 23357 -1123 23358 -1113
rect 23232 -1147 23266 -1123
rect 23324 -1147 23358 -1123
rect 23416 -1123 23417 -1113
rect 23417 -1123 23450 -1113
rect 23508 -1123 23542 -1113
rect 23416 -1147 23450 -1123
rect 23508 -1147 23542 -1123
rect 23600 -1123 23634 -1113
rect 23600 -1147 23634 -1123
rect 23692 -1123 23726 -1113
rect 23692 -1147 23726 -1123
rect 23784 -1123 23818 -1113
rect 23784 -1147 23818 -1123
rect 23876 -1123 23910 -1113
rect 23876 -1147 23910 -1123
rect 23968 -1123 24002 -1113
rect 23968 -1147 24002 -1123
rect 24060 -1123 24094 -1113
rect 24060 -1147 24094 -1123
rect 24152 -1123 24186 -1113
rect 24152 -1147 24186 -1123
rect 24244 -1123 24278 -1113
rect 24244 -1147 24278 -1123
rect 24336 -1123 24370 -1113
rect 24336 -1147 24370 -1123
rect 24428 -1123 24462 -1113
rect 24428 -1147 24462 -1123
rect 24520 -1130 24534 -1113
rect 24534 -1130 24554 -1113
rect 24520 -1147 24554 -1130
rect 24612 -1147 24646 -1113
rect 24704 -1123 24738 -1113
rect 24704 -1147 24738 -1123
rect 24796 -1123 24830 -1113
rect 24796 -1147 24830 -1123
rect 24888 -1123 24922 -1113
rect 24888 -1147 24922 -1123
rect 24980 -1123 25014 -1113
rect 24980 -1147 25014 -1123
rect 25072 -1123 25106 -1113
rect 25072 -1147 25106 -1123
rect 25164 -1123 25198 -1113
rect 25164 -1147 25198 -1123
rect 25256 -1123 25290 -1113
rect 25256 -1147 25290 -1123
rect 8601 -1225 8635 -1223
rect 8601 -1257 8610 -1225
rect 8610 -1257 8635 -1225
rect 8881 -1294 8915 -1289
rect 8881 -1323 8893 -1294
rect 8893 -1323 8915 -1294
rect 9162 -1385 9196 -1351
rect 9077 -1421 9111 -1417
rect 9077 -1451 9104 -1421
rect 9104 -1451 9111 -1421
rect 9418 -1495 9422 -1487
rect 9422 -1495 9452 -1487
rect 9418 -1521 9452 -1495
rect 9708 -1309 9742 -1283
rect 9708 -1317 9721 -1309
rect 9721 -1317 9742 -1309
rect 9800 -1385 9834 -1351
rect 9708 -1453 9742 -1419
rect 10444 -1317 10478 -1283
rect 10168 -1495 10200 -1487
rect 10200 -1495 10202 -1487
rect 10168 -1521 10202 -1495
rect 10352 -1505 10372 -1487
rect 10372 -1505 10386 -1487
rect 10352 -1521 10386 -1505
rect 10543 -1450 10577 -1416
rect 10720 -1299 10730 -1283
rect 10730 -1299 10754 -1283
rect 10720 -1317 10754 -1299
rect 10993 -1225 11027 -1223
rect 10993 -1257 11002 -1225
rect 11002 -1257 11027 -1225
rect 10889 -1394 10923 -1360
rect 10811 -1521 10845 -1487
rect 11273 -1294 11307 -1289
rect 11273 -1323 11285 -1294
rect 11285 -1323 11307 -1294
rect 11554 -1385 11588 -1351
rect 11466 -1421 11500 -1415
rect 11466 -1449 11496 -1421
rect 11496 -1449 11500 -1421
rect 11810 -1495 11814 -1487
rect 11814 -1495 11844 -1487
rect 11810 -1521 11844 -1495
rect 12100 -1309 12134 -1283
rect 12100 -1317 12113 -1309
rect 12113 -1317 12134 -1309
rect 12192 -1385 12226 -1351
rect 12100 -1453 12134 -1419
rect 12836 -1317 12870 -1283
rect 12560 -1495 12592 -1487
rect 12592 -1495 12594 -1487
rect 12560 -1521 12594 -1495
rect 12744 -1505 12764 -1487
rect 12764 -1505 12778 -1487
rect 12744 -1521 12778 -1505
rect 12935 -1450 12969 -1416
rect 13112 -1299 13122 -1283
rect 13122 -1299 13146 -1283
rect 13112 -1317 13146 -1299
rect 13386 -1225 13420 -1223
rect 13386 -1257 13394 -1225
rect 13394 -1257 13420 -1225
rect 13283 -1394 13317 -1360
rect 13203 -1521 13237 -1487
rect 13664 -1294 13698 -1289
rect 13664 -1323 13677 -1294
rect 13677 -1323 13698 -1294
rect 13946 -1385 13980 -1351
rect 13859 -1421 13893 -1415
rect 13859 -1449 13888 -1421
rect 13888 -1449 13893 -1421
rect 14202 -1495 14206 -1487
rect 14206 -1495 14236 -1487
rect 14202 -1521 14236 -1495
rect 14492 -1309 14526 -1283
rect 14492 -1317 14505 -1309
rect 14505 -1317 14526 -1309
rect 14584 -1385 14618 -1351
rect 14492 -1453 14526 -1419
rect 15228 -1317 15262 -1283
rect 14952 -1495 14984 -1487
rect 14984 -1495 14986 -1487
rect 14952 -1521 14986 -1495
rect 15136 -1505 15156 -1487
rect 15156 -1505 15170 -1487
rect 15136 -1521 15170 -1505
rect 15326 -1449 15360 -1415
rect 15504 -1299 15514 -1283
rect 15514 -1299 15538 -1283
rect 15504 -1317 15538 -1299
rect 15777 -1225 15811 -1223
rect 15777 -1257 15786 -1225
rect 15786 -1257 15811 -1225
rect 15673 -1392 15707 -1358
rect 15595 -1521 15629 -1487
rect 16057 -1294 16091 -1289
rect 16057 -1323 16069 -1294
rect 16069 -1323 16091 -1294
rect 16338 -1385 16372 -1351
rect 16252 -1421 16286 -1415
rect 16252 -1449 16280 -1421
rect 16280 -1449 16286 -1421
rect 16594 -1495 16598 -1487
rect 16598 -1495 16628 -1487
rect 16594 -1521 16628 -1495
rect 16884 -1309 16918 -1283
rect 16884 -1317 16897 -1309
rect 16897 -1317 16918 -1309
rect 16976 -1385 17010 -1351
rect 16884 -1453 16918 -1419
rect 17620 -1317 17654 -1283
rect 17344 -1495 17376 -1487
rect 17376 -1495 17378 -1487
rect 17344 -1521 17378 -1495
rect 17528 -1505 17548 -1487
rect 17548 -1505 17562 -1487
rect 17528 -1521 17562 -1505
rect 17719 -1450 17753 -1416
rect 17896 -1299 17906 -1283
rect 17906 -1299 17930 -1283
rect 17896 -1317 17930 -1299
rect 18169 -1225 18203 -1224
rect 18169 -1258 18178 -1225
rect 18178 -1258 18203 -1225
rect 18065 -1394 18099 -1360
rect 17987 -1521 18021 -1487
rect 18449 -1294 18483 -1289
rect 18449 -1323 18461 -1294
rect 18461 -1323 18483 -1294
rect 18730 -1385 18764 -1351
rect 18643 -1421 18677 -1415
rect 18643 -1449 18672 -1421
rect 18672 -1449 18677 -1421
rect 18986 -1495 18990 -1487
rect 18990 -1495 19020 -1487
rect 18986 -1521 19020 -1495
rect 19276 -1309 19310 -1283
rect 19276 -1317 19289 -1309
rect 19289 -1317 19310 -1309
rect 19368 -1385 19402 -1351
rect 19276 -1453 19310 -1419
rect 20012 -1317 20046 -1283
rect 19736 -1495 19768 -1487
rect 19768 -1495 19770 -1487
rect 19736 -1521 19770 -1495
rect 19920 -1505 19940 -1487
rect 19940 -1505 19954 -1487
rect 19920 -1521 19954 -1505
rect 20110 -1450 20144 -1416
rect 20288 -1299 20298 -1283
rect 20298 -1299 20322 -1283
rect 20288 -1317 20322 -1299
rect 20562 -1225 20596 -1222
rect 20562 -1256 20570 -1225
rect 20570 -1256 20596 -1225
rect 20457 -1392 20491 -1358
rect 20379 -1521 20413 -1487
rect 20840 -1294 20874 -1288
rect 20840 -1322 20853 -1294
rect 20853 -1322 20874 -1294
rect 21122 -1385 21156 -1351
rect 21036 -1421 21070 -1415
rect 21036 -1449 21064 -1421
rect 21064 -1449 21070 -1421
rect 21378 -1495 21382 -1487
rect 21382 -1495 21412 -1487
rect 21378 -1521 21412 -1495
rect 21668 -1309 21702 -1283
rect 21668 -1317 21681 -1309
rect 21681 -1317 21702 -1309
rect 21760 -1385 21794 -1351
rect 21668 -1453 21702 -1419
rect 22404 -1317 22438 -1283
rect 22128 -1495 22160 -1487
rect 22160 -1495 22162 -1487
rect 22128 -1521 22162 -1495
rect 22312 -1505 22332 -1487
rect 22332 -1505 22346 -1487
rect 22312 -1521 22346 -1505
rect 22503 -1450 22537 -1416
rect 22680 -1299 22690 -1283
rect 22690 -1299 22714 -1283
rect 22680 -1317 22714 -1299
rect 22953 -1225 22987 -1222
rect 22953 -1256 22962 -1225
rect 22962 -1256 22987 -1225
rect 22849 -1394 22883 -1360
rect 22771 -1521 22805 -1487
rect 23233 -1294 23267 -1289
rect 23233 -1323 23245 -1294
rect 23245 -1323 23267 -1294
rect 23514 -1385 23548 -1351
rect 23427 -1421 23461 -1415
rect 23427 -1449 23456 -1421
rect 23456 -1449 23461 -1421
rect 23770 -1495 23774 -1487
rect 23774 -1495 23804 -1487
rect 23770 -1521 23804 -1495
rect 24060 -1309 24094 -1283
rect 24060 -1317 24073 -1309
rect 24073 -1317 24094 -1309
rect 24152 -1385 24186 -1351
rect 24060 -1453 24094 -1419
rect 24796 -1317 24830 -1283
rect 24520 -1495 24552 -1487
rect 24552 -1495 24554 -1487
rect 24520 -1521 24554 -1495
rect 24704 -1505 24724 -1487
rect 24724 -1505 24738 -1487
rect 24704 -1521 24738 -1505
rect 24896 -1450 24930 -1416
rect 25072 -1299 25082 -1283
rect 25082 -1299 25106 -1283
rect 25072 -1317 25106 -1299
rect 25241 -1392 25275 -1358
rect 25163 -1521 25197 -1487
rect 8604 -1681 8638 -1657
rect 8604 -1691 8638 -1681
rect 8696 -1681 8730 -1657
rect 8696 -1691 8730 -1681
rect 8788 -1681 8822 -1657
rect 8788 -1691 8822 -1681
rect 8880 -1681 8914 -1657
rect 8880 -1691 8914 -1681
rect 8972 -1681 9006 -1657
rect 8972 -1691 9006 -1681
rect 9064 -1681 9098 -1657
rect 9064 -1691 9098 -1681
rect 9156 -1681 9190 -1657
rect 9156 -1691 9190 -1681
rect 9248 -1681 9282 -1657
rect 9248 -1691 9282 -1681
rect 9340 -1681 9374 -1657
rect 9340 -1691 9374 -1681
rect 9432 -1681 9466 -1657
rect 9432 -1691 9466 -1681
rect 9524 -1681 9558 -1657
rect 9524 -1691 9558 -1681
rect 9616 -1681 9650 -1657
rect 9616 -1691 9650 -1681
rect 9708 -1681 9742 -1657
rect 9708 -1691 9742 -1681
rect 9800 -1681 9834 -1657
rect 9800 -1691 9834 -1681
rect 9892 -1681 9926 -1657
rect 9892 -1691 9926 -1681
rect 9984 -1681 10018 -1657
rect 9984 -1691 10018 -1681
rect 10076 -1681 10110 -1657
rect 10076 -1691 10110 -1681
rect 10168 -1681 10202 -1657
rect 10168 -1691 10202 -1681
rect 10260 -1681 10294 -1657
rect 10260 -1691 10294 -1681
rect 10352 -1681 10386 -1657
rect 10352 -1691 10386 -1681
rect 10444 -1681 10478 -1657
rect 10444 -1691 10478 -1681
rect 10536 -1681 10570 -1657
rect 10536 -1691 10570 -1681
rect 10628 -1681 10662 -1657
rect 10628 -1691 10662 -1681
rect 10720 -1681 10754 -1657
rect 10720 -1691 10754 -1681
rect 10812 -1681 10846 -1657
rect 10812 -1691 10846 -1681
rect 10904 -1681 10938 -1657
rect 10904 -1691 10938 -1681
rect 10996 -1681 11030 -1657
rect 10996 -1691 11030 -1681
rect 11088 -1681 11122 -1657
rect 11088 -1691 11122 -1681
rect 11180 -1681 11214 -1657
rect 11180 -1691 11214 -1681
rect 11272 -1681 11306 -1657
rect 11272 -1691 11306 -1681
rect 11364 -1681 11398 -1657
rect 11364 -1691 11398 -1681
rect 11456 -1681 11490 -1657
rect 11456 -1691 11490 -1681
rect 11548 -1681 11582 -1657
rect 11548 -1691 11582 -1681
rect 11640 -1681 11674 -1657
rect 11640 -1691 11674 -1681
rect 11732 -1681 11766 -1657
rect 11732 -1691 11766 -1681
rect 11824 -1681 11858 -1657
rect 11824 -1691 11858 -1681
rect 11916 -1681 11950 -1657
rect 11916 -1691 11950 -1681
rect 12008 -1681 12042 -1657
rect 12008 -1691 12042 -1681
rect 12100 -1681 12134 -1657
rect 12100 -1691 12134 -1681
rect 12192 -1681 12226 -1657
rect 12192 -1691 12226 -1681
rect 12284 -1681 12318 -1657
rect 12284 -1691 12318 -1681
rect 12376 -1681 12410 -1657
rect 12376 -1691 12410 -1681
rect 12468 -1681 12502 -1657
rect 12468 -1691 12502 -1681
rect 12560 -1681 12594 -1657
rect 12560 -1691 12594 -1681
rect 12652 -1681 12686 -1657
rect 12652 -1691 12686 -1681
rect 12744 -1681 12778 -1657
rect 12744 -1691 12778 -1681
rect 12836 -1681 12870 -1657
rect 12836 -1691 12870 -1681
rect 12928 -1681 12962 -1657
rect 12928 -1691 12962 -1681
rect 13020 -1681 13054 -1657
rect 13020 -1691 13054 -1681
rect 13112 -1681 13146 -1657
rect 13112 -1691 13146 -1681
rect 13204 -1681 13238 -1657
rect 13204 -1691 13238 -1681
rect 13296 -1681 13330 -1657
rect 13296 -1691 13330 -1681
rect 13388 -1681 13422 -1657
rect 13388 -1691 13422 -1681
rect 13480 -1681 13514 -1657
rect 13480 -1691 13514 -1681
rect 13572 -1681 13606 -1657
rect 13572 -1691 13606 -1681
rect 13664 -1681 13698 -1657
rect 13664 -1691 13698 -1681
rect 13756 -1681 13790 -1657
rect 13756 -1691 13790 -1681
rect 13848 -1681 13882 -1657
rect 13848 -1691 13882 -1681
rect 13940 -1681 13974 -1657
rect 13940 -1691 13974 -1681
rect 14032 -1681 14066 -1657
rect 14032 -1691 14066 -1681
rect 14124 -1681 14158 -1657
rect 14124 -1691 14158 -1681
rect 14216 -1681 14250 -1657
rect 14216 -1691 14250 -1681
rect 14308 -1681 14342 -1657
rect 14308 -1691 14342 -1681
rect 14400 -1681 14434 -1657
rect 14400 -1691 14434 -1681
rect 14492 -1681 14526 -1657
rect 14492 -1691 14526 -1681
rect 14584 -1681 14618 -1657
rect 14584 -1691 14618 -1681
rect 14676 -1681 14710 -1657
rect 14676 -1691 14710 -1681
rect 14768 -1681 14802 -1657
rect 14768 -1691 14802 -1681
rect 14860 -1681 14894 -1657
rect 14860 -1691 14894 -1681
rect 14952 -1681 14986 -1657
rect 14952 -1691 14986 -1681
rect 15044 -1681 15078 -1657
rect 15044 -1691 15078 -1681
rect 15136 -1681 15170 -1657
rect 15136 -1691 15170 -1681
rect 15228 -1681 15262 -1657
rect 15228 -1691 15262 -1681
rect 15320 -1681 15354 -1657
rect 15320 -1691 15354 -1681
rect 15412 -1681 15446 -1657
rect 15412 -1691 15446 -1681
rect 15504 -1681 15538 -1657
rect 15504 -1691 15538 -1681
rect 15596 -1681 15630 -1657
rect 15596 -1691 15630 -1681
rect 15688 -1681 15722 -1657
rect 15688 -1691 15722 -1681
rect 15780 -1681 15814 -1657
rect 15780 -1691 15814 -1681
rect 15872 -1681 15906 -1657
rect 15872 -1691 15906 -1681
rect 15964 -1681 15998 -1657
rect 15964 -1691 15998 -1681
rect 16056 -1681 16090 -1657
rect 16056 -1691 16090 -1681
rect 16148 -1681 16182 -1657
rect 16148 -1691 16182 -1681
rect 16240 -1681 16274 -1657
rect 16240 -1691 16274 -1681
rect 16332 -1681 16366 -1657
rect 16332 -1691 16366 -1681
rect 16424 -1681 16458 -1657
rect 16424 -1691 16458 -1681
rect 16516 -1681 16550 -1657
rect 16516 -1691 16550 -1681
rect 16608 -1681 16642 -1657
rect 16608 -1691 16642 -1681
rect 16700 -1681 16734 -1657
rect 16700 -1691 16734 -1681
rect 16792 -1681 16826 -1657
rect 16792 -1691 16826 -1681
rect 16884 -1681 16918 -1657
rect 16884 -1691 16918 -1681
rect 16976 -1681 17010 -1657
rect 16976 -1691 17010 -1681
rect 17068 -1681 17102 -1657
rect 17068 -1691 17102 -1681
rect 17160 -1681 17194 -1657
rect 17160 -1691 17194 -1681
rect 17252 -1681 17286 -1657
rect 17252 -1691 17286 -1681
rect 17344 -1681 17378 -1657
rect 17344 -1691 17378 -1681
rect 17436 -1681 17470 -1657
rect 17436 -1691 17470 -1681
rect 17528 -1681 17562 -1657
rect 17528 -1691 17562 -1681
rect 17620 -1681 17654 -1657
rect 17620 -1691 17654 -1681
rect 17712 -1681 17746 -1657
rect 17712 -1691 17746 -1681
rect 17804 -1681 17838 -1657
rect 17804 -1691 17838 -1681
rect 17896 -1681 17930 -1657
rect 17896 -1691 17930 -1681
rect 17988 -1681 18022 -1657
rect 17988 -1691 18022 -1681
rect 18080 -1681 18114 -1657
rect 18080 -1691 18114 -1681
rect 18172 -1681 18206 -1657
rect 18172 -1691 18206 -1681
rect 18264 -1681 18298 -1657
rect 18264 -1691 18298 -1681
rect 18356 -1681 18390 -1657
rect 18356 -1691 18390 -1681
rect 18448 -1681 18482 -1657
rect 18448 -1691 18482 -1681
rect 18540 -1681 18574 -1657
rect 18540 -1691 18574 -1681
rect 18632 -1681 18666 -1657
rect 18632 -1691 18666 -1681
rect 18724 -1681 18758 -1657
rect 18724 -1691 18758 -1681
rect 18816 -1681 18850 -1657
rect 18816 -1691 18850 -1681
rect 18908 -1681 18942 -1657
rect 18908 -1691 18942 -1681
rect 19000 -1681 19034 -1657
rect 19000 -1691 19034 -1681
rect 19092 -1681 19126 -1657
rect 19092 -1691 19126 -1681
rect 19184 -1681 19218 -1657
rect 19184 -1691 19218 -1681
rect 19276 -1681 19310 -1657
rect 19276 -1691 19310 -1681
rect 19368 -1681 19402 -1657
rect 19368 -1691 19402 -1681
rect 19460 -1681 19494 -1657
rect 19460 -1691 19494 -1681
rect 19552 -1681 19586 -1657
rect 19552 -1691 19586 -1681
rect 19644 -1681 19678 -1657
rect 19644 -1691 19678 -1681
rect 19736 -1681 19770 -1657
rect 19736 -1691 19770 -1681
rect 19828 -1681 19862 -1657
rect 19828 -1691 19862 -1681
rect 19920 -1681 19954 -1657
rect 19920 -1691 19954 -1681
rect 20012 -1681 20046 -1657
rect 20012 -1691 20046 -1681
rect 20104 -1681 20138 -1657
rect 20104 -1691 20138 -1681
rect 20196 -1681 20230 -1657
rect 20196 -1691 20230 -1681
rect 20288 -1681 20322 -1657
rect 20288 -1691 20322 -1681
rect 20380 -1681 20414 -1657
rect 20380 -1691 20414 -1681
rect 20472 -1681 20506 -1657
rect 20472 -1691 20506 -1681
rect 20564 -1681 20598 -1657
rect 20564 -1691 20598 -1681
rect 20656 -1681 20690 -1657
rect 20656 -1691 20690 -1681
rect 20748 -1681 20782 -1657
rect 20748 -1691 20782 -1681
rect 20840 -1681 20874 -1657
rect 20840 -1691 20874 -1681
rect 20932 -1681 20966 -1657
rect 20932 -1691 20966 -1681
rect 21024 -1681 21058 -1657
rect 21024 -1691 21058 -1681
rect 21116 -1681 21150 -1657
rect 21116 -1691 21150 -1681
rect 21208 -1681 21242 -1657
rect 21208 -1691 21242 -1681
rect 21300 -1681 21334 -1657
rect 21300 -1691 21334 -1681
rect 21392 -1681 21426 -1657
rect 21392 -1691 21426 -1681
rect 21484 -1681 21518 -1657
rect 21484 -1691 21518 -1681
rect 21576 -1681 21610 -1657
rect 21576 -1691 21610 -1681
rect 21668 -1681 21702 -1657
rect 21668 -1691 21702 -1681
rect 21760 -1681 21794 -1657
rect 21760 -1691 21794 -1681
rect 21852 -1681 21886 -1657
rect 21852 -1691 21886 -1681
rect 21944 -1681 21978 -1657
rect 21944 -1691 21978 -1681
rect 22036 -1681 22070 -1657
rect 22036 -1691 22070 -1681
rect 22128 -1681 22162 -1657
rect 22128 -1691 22162 -1681
rect 22220 -1681 22254 -1657
rect 22220 -1691 22254 -1681
rect 22312 -1681 22346 -1657
rect 22312 -1691 22346 -1681
rect 22404 -1681 22438 -1657
rect 22404 -1691 22438 -1681
rect 22496 -1681 22530 -1657
rect 22496 -1691 22530 -1681
rect 22588 -1681 22622 -1657
rect 22588 -1691 22622 -1681
rect 22680 -1681 22714 -1657
rect 22680 -1691 22714 -1681
rect 22772 -1681 22806 -1657
rect 22772 -1691 22806 -1681
rect 22864 -1681 22898 -1657
rect 22864 -1691 22898 -1681
rect 22956 -1681 22990 -1657
rect 22956 -1691 22990 -1681
rect 23048 -1681 23082 -1657
rect 23048 -1691 23082 -1681
rect 23140 -1681 23174 -1657
rect 23140 -1691 23174 -1681
rect 23232 -1681 23266 -1657
rect 23232 -1691 23266 -1681
rect 23324 -1681 23358 -1657
rect 23324 -1691 23358 -1681
rect 23416 -1681 23450 -1657
rect 23416 -1691 23450 -1681
rect 23508 -1681 23542 -1657
rect 23508 -1691 23542 -1681
rect 23600 -1681 23634 -1657
rect 23600 -1691 23634 -1681
rect 23692 -1681 23726 -1657
rect 23692 -1691 23726 -1681
rect 23784 -1681 23818 -1657
rect 23784 -1691 23818 -1681
rect 23876 -1681 23910 -1657
rect 23876 -1691 23910 -1681
rect 23968 -1681 24002 -1657
rect 23968 -1691 24002 -1681
rect 24060 -1681 24094 -1657
rect 24060 -1691 24094 -1681
rect 24152 -1681 24186 -1657
rect 24152 -1691 24186 -1681
rect 24244 -1681 24278 -1657
rect 24244 -1691 24278 -1681
rect 24336 -1681 24370 -1657
rect 24336 -1691 24370 -1681
rect 24428 -1681 24462 -1657
rect 24428 -1691 24462 -1681
rect 24520 -1681 24554 -1657
rect 24520 -1691 24554 -1681
rect 24612 -1681 24646 -1657
rect 24612 -1691 24646 -1681
rect 24704 -1681 24738 -1657
rect 24704 -1691 24738 -1681
rect 24796 -1681 24830 -1657
rect 24796 -1691 24830 -1681
rect 24888 -1681 24922 -1657
rect 24888 -1691 24922 -1681
rect 24980 -1681 25014 -1657
rect 24980 -1691 25014 -1681
rect 25072 -1681 25106 -1657
rect 25072 -1691 25106 -1681
rect 25164 -1681 25198 -1657
rect 25164 -1691 25198 -1681
rect 25256 -1681 25290 -1657
rect 25256 -1691 25290 -1681
<< metal1 >>
rect 13937 13626 14027 13642
rect 20646 13626 20736 13642
rect 13937 13615 13956 13626
rect 13919 13593 13956 13615
rect 13810 13581 13856 13593
rect 13810 13521 13816 13581
rect 13850 13521 13856 13581
rect 13810 13443 13856 13521
rect 13898 13581 13956 13593
rect 13898 13521 13904 13581
rect 13938 13574 13956 13581
rect 14008 13623 14027 13626
rect 14008 13617 14616 13623
rect 14008 13574 14054 13617
rect 13938 13565 14054 13574
rect 14106 13565 14134 13617
rect 14186 13565 14214 13617
rect 14266 13565 14294 13617
rect 14346 13565 14374 13617
rect 14426 13565 14454 13617
rect 14506 13565 14616 13617
rect 13938 13557 14616 13565
rect 14678 13620 19586 13626
rect 14678 13568 14786 13620
rect 14838 13568 14866 13620
rect 14918 13568 14946 13620
rect 14998 13568 15026 13620
rect 15078 13568 15106 13620
rect 15158 13568 15186 13620
rect 15238 13568 15390 13620
rect 15442 13568 15470 13620
rect 15522 13568 15550 13620
rect 15602 13568 15630 13620
rect 15682 13568 15710 13620
rect 15762 13568 15790 13620
rect 15842 13568 15998 13620
rect 16050 13568 16078 13620
rect 16130 13568 16158 13620
rect 16210 13568 16238 13620
rect 16290 13568 16318 13620
rect 16370 13568 16398 13620
rect 16450 13568 16602 13620
rect 16654 13568 16682 13620
rect 16734 13568 16762 13620
rect 16814 13568 16842 13620
rect 16894 13568 16922 13620
rect 16974 13568 17002 13620
rect 17054 13568 17210 13620
rect 17262 13568 17290 13620
rect 17342 13568 17370 13620
rect 17422 13568 17450 13620
rect 17502 13568 17530 13620
rect 17582 13568 17610 13620
rect 17662 13568 17814 13620
rect 17866 13568 17894 13620
rect 17946 13568 17974 13620
rect 18026 13568 18054 13620
rect 18106 13568 18134 13620
rect 18186 13568 18214 13620
rect 18266 13568 18422 13620
rect 18474 13568 18502 13620
rect 18554 13568 18582 13620
rect 18634 13568 18662 13620
rect 18714 13568 18742 13620
rect 18794 13568 18822 13620
rect 18874 13568 19026 13620
rect 19078 13568 19106 13620
rect 19158 13568 19186 13620
rect 19238 13568 19266 13620
rect 19318 13568 19346 13620
rect 19398 13568 19426 13620
rect 19478 13568 19586 13620
rect 20646 13615 20665 13626
rect 20628 13593 20665 13615
rect 14678 13560 19586 13568
rect 19746 13564 19836 13580
rect 13938 13527 13972 13557
rect 13938 13521 13944 13527
rect 13898 13509 13944 13521
rect 19746 13512 19765 13564
rect 19817 13512 19836 13564
rect 19746 13496 19836 13512
rect 20223 13567 20313 13583
rect 20223 13515 20242 13567
rect 20294 13515 20313 13567
rect 20223 13499 20313 13515
rect 20519 13581 20565 13593
rect 20519 13521 20525 13581
rect 20559 13521 20565 13581
rect 13810 13383 13816 13443
rect 13850 13383 13856 13443
rect 13810 13371 13856 13383
rect 13898 13443 13944 13455
rect 13898 13383 13904 13443
rect 13938 13383 13944 13443
rect 20519 13443 20565 13521
rect 20607 13581 20665 13593
rect 20607 13521 20613 13581
rect 20647 13574 20665 13581
rect 20717 13623 20736 13626
rect 20717 13617 21325 13623
rect 20717 13574 20763 13617
rect 20647 13565 20763 13574
rect 20815 13565 20843 13617
rect 20895 13565 20923 13617
rect 20975 13565 21003 13617
rect 21055 13565 21083 13617
rect 21135 13565 21163 13617
rect 21215 13565 21325 13617
rect 20647 13557 21325 13565
rect 21387 13620 26295 13626
rect 21387 13568 21495 13620
rect 21547 13568 21575 13620
rect 21627 13568 21655 13620
rect 21707 13568 21735 13620
rect 21787 13568 21815 13620
rect 21867 13568 21895 13620
rect 21947 13568 22099 13620
rect 22151 13568 22179 13620
rect 22231 13568 22259 13620
rect 22311 13568 22339 13620
rect 22391 13568 22419 13620
rect 22471 13568 22499 13620
rect 22551 13568 22707 13620
rect 22759 13568 22787 13620
rect 22839 13568 22867 13620
rect 22919 13568 22947 13620
rect 22999 13568 23027 13620
rect 23079 13568 23107 13620
rect 23159 13568 23311 13620
rect 23363 13568 23391 13620
rect 23443 13568 23471 13620
rect 23523 13568 23551 13620
rect 23603 13568 23631 13620
rect 23683 13568 23711 13620
rect 23763 13568 23919 13620
rect 23971 13568 23999 13620
rect 24051 13568 24079 13620
rect 24131 13568 24159 13620
rect 24211 13568 24239 13620
rect 24291 13568 24319 13620
rect 24371 13568 24523 13620
rect 24575 13568 24603 13620
rect 24655 13568 24683 13620
rect 24735 13568 24763 13620
rect 24815 13568 24843 13620
rect 24895 13568 24923 13620
rect 24975 13568 25131 13620
rect 25183 13568 25211 13620
rect 25263 13568 25291 13620
rect 25343 13568 25371 13620
rect 25423 13568 25451 13620
rect 25503 13568 25531 13620
rect 25583 13568 25735 13620
rect 25787 13568 25815 13620
rect 25867 13568 25895 13620
rect 25947 13568 25975 13620
rect 26027 13568 26055 13620
rect 26107 13568 26135 13620
rect 26187 13568 26295 13620
rect 21387 13560 26295 13568
rect 26455 13564 26545 13580
rect 20647 13527 20681 13557
rect 20647 13521 20653 13527
rect 20607 13509 20653 13521
rect 26455 13512 26474 13564
rect 26526 13512 26545 13564
rect 26455 13496 26545 13512
rect 13810 13305 13856 13317
rect 13810 13245 13816 13305
rect 13850 13245 13856 13305
rect 13810 13167 13856 13245
rect 13898 13305 13944 13383
rect 19751 13420 19841 13436
rect 19751 13368 19770 13420
rect 19822 13368 19841 13420
rect 19751 13352 19841 13368
rect 20212 13395 20302 13411
rect 20212 13343 20231 13395
rect 20283 13343 20302 13395
rect 20519 13383 20525 13443
rect 20559 13383 20565 13443
rect 20519 13371 20565 13383
rect 20607 13443 20653 13455
rect 20607 13383 20613 13443
rect 20647 13383 20653 13443
rect 20212 13327 20302 13343
rect 13898 13245 13904 13305
rect 13938 13245 13944 13305
rect 20519 13305 20565 13317
rect 13898 13233 13944 13245
rect 19752 13268 19842 13284
rect 19752 13216 19771 13268
rect 19823 13216 19842 13268
rect 20519 13245 20525 13305
rect 20559 13245 20565 13305
rect 19752 13200 19842 13216
rect 20212 13203 20302 13219
rect 3049 13151 3139 13167
rect 3049 13140 3068 13151
rect 3031 13118 3068 13140
rect 2922 13106 2968 13118
rect 2922 13046 2928 13106
rect 2962 13046 2968 13106
rect 2922 12968 2968 13046
rect 3010 13106 3068 13118
rect 3010 13046 3016 13106
rect 3050 13099 3068 13106
rect 3120 13148 3139 13151
rect 3120 13142 3728 13148
rect 3120 13099 3166 13142
rect 3050 13090 3166 13099
rect 3218 13090 3246 13142
rect 3298 13090 3326 13142
rect 3378 13090 3406 13142
rect 3458 13090 3486 13142
rect 3538 13090 3566 13142
rect 3618 13090 3728 13142
rect 3050 13082 3728 13090
rect 3790 13145 8698 13151
rect 3790 13093 3898 13145
rect 3950 13093 3978 13145
rect 4030 13093 4058 13145
rect 4110 13093 4138 13145
rect 4190 13093 4218 13145
rect 4270 13093 4298 13145
rect 4350 13093 4502 13145
rect 4554 13093 4582 13145
rect 4634 13093 4662 13145
rect 4714 13093 4742 13145
rect 4794 13093 4822 13145
rect 4874 13093 4902 13145
rect 4954 13093 5110 13145
rect 5162 13093 5190 13145
rect 5242 13093 5270 13145
rect 5322 13093 5350 13145
rect 5402 13093 5430 13145
rect 5482 13093 5510 13145
rect 5562 13093 5714 13145
rect 5766 13093 5794 13145
rect 5846 13093 5874 13145
rect 5926 13093 5954 13145
rect 6006 13093 6034 13145
rect 6086 13093 6114 13145
rect 6166 13093 6322 13145
rect 6374 13093 6402 13145
rect 6454 13093 6482 13145
rect 6534 13093 6562 13145
rect 6614 13093 6642 13145
rect 6694 13093 6722 13145
rect 6774 13093 6926 13145
rect 6978 13093 7006 13145
rect 7058 13093 7086 13145
rect 7138 13093 7166 13145
rect 7218 13093 7246 13145
rect 7298 13093 7326 13145
rect 7378 13093 7534 13145
rect 7586 13093 7614 13145
rect 7666 13093 7694 13145
rect 7746 13093 7774 13145
rect 7826 13093 7854 13145
rect 7906 13093 7934 13145
rect 7986 13093 8138 13145
rect 8190 13093 8218 13145
rect 8270 13093 8298 13145
rect 8350 13093 8378 13145
rect 8430 13093 8458 13145
rect 8510 13093 8538 13145
rect 8590 13093 8698 13145
rect 13810 13107 13816 13167
rect 13850 13107 13856 13167
rect 3790 13085 8698 13093
rect 8858 13089 8948 13105
rect 13810 13095 13856 13107
rect 13898 13167 13944 13179
rect 13898 13107 13904 13167
rect 13938 13107 13944 13167
rect 20212 13151 20231 13203
rect 20283 13151 20302 13203
rect 20212 13135 20302 13151
rect 20519 13167 20565 13245
rect 20607 13305 20653 13383
rect 26460 13420 26550 13436
rect 26460 13368 26479 13420
rect 26531 13368 26550 13420
rect 26460 13352 26550 13368
rect 20607 13245 20613 13305
rect 20647 13245 20653 13305
rect 20607 13233 20653 13245
rect 26461 13268 26551 13284
rect 26461 13216 26480 13268
rect 26532 13216 26551 13268
rect 26461 13200 26551 13216
rect 3050 13052 3084 13082
rect 3050 13046 3056 13052
rect 3010 13034 3056 13046
rect 8858 13037 8877 13089
rect 8929 13037 8948 13089
rect 8858 13021 8948 13037
rect 13274 13021 13734 13041
rect 13274 13010 13339 13021
rect 2922 12908 2928 12968
rect 2962 12908 2968 12968
rect 2922 12896 2968 12908
rect 3010 12968 3056 12980
rect 3010 12908 3016 12968
rect 3050 12908 3056 12968
rect 13274 12976 13303 13010
rect 13337 12976 13339 13010
rect 13274 12969 13339 12976
rect 13391 13020 13614 13021
rect 13391 13010 13470 13020
rect 13522 13010 13614 13020
rect 13391 12976 13395 13010
rect 13429 12976 13470 13010
rect 13522 12976 13579 13010
rect 13613 12976 13614 13010
rect 13391 12969 13470 12976
rect 13274 12968 13470 12969
rect 13522 12969 13614 12976
rect 13666 13010 13734 13021
rect 13666 12976 13671 13010
rect 13705 12976 13734 13010
rect 13666 12969 13734 12976
rect 13522 12968 13734 12969
rect 2922 12830 2968 12842
rect 2922 12770 2928 12830
rect 2962 12770 2968 12830
rect 2922 12692 2968 12770
rect 3010 12830 3056 12908
rect 8863 12945 8953 12961
rect 13274 12945 13734 12968
rect 13810 13029 13856 13041
rect 13810 12969 13816 13029
rect 13850 12969 13856 13029
rect 8863 12893 8882 12945
rect 8934 12893 8953 12945
rect 8863 12877 8953 12893
rect 13810 12891 13856 12969
rect 13898 13029 13944 13107
rect 19752 13098 19842 13114
rect 19752 13046 19771 13098
rect 19823 13046 19842 13098
rect 20519 13107 20525 13167
rect 20559 13107 20565 13167
rect 20519 13095 20565 13107
rect 20607 13167 20653 13179
rect 20607 13107 20613 13167
rect 20647 13107 20653 13167
rect 19752 13030 19842 13046
rect 13898 12969 13904 13029
rect 13938 12969 13944 13029
rect 13898 12957 13944 12969
rect 19983 13021 20443 13041
rect 19983 13010 20048 13021
rect 19983 12976 20012 13010
rect 20046 12976 20048 13010
rect 19983 12969 20048 12976
rect 20100 13020 20323 13021
rect 20100 13010 20179 13020
rect 20231 13010 20323 13020
rect 20100 12976 20104 13010
rect 20138 12976 20179 13010
rect 20231 12976 20288 13010
rect 20322 12976 20323 13010
rect 20100 12969 20179 12976
rect 19983 12968 20179 12969
rect 20231 12969 20323 12976
rect 20375 13010 20443 13021
rect 20375 12976 20380 13010
rect 20414 12976 20443 13010
rect 20375 12969 20443 12976
rect 20231 12968 20443 12969
rect 19751 12941 19841 12957
rect 19983 12945 20443 12968
rect 20519 13029 20565 13041
rect 20519 12969 20525 13029
rect 20559 12969 20565 13029
rect 3010 12770 3016 12830
rect 3050 12770 3056 12830
rect 13419 12867 13782 12874
rect 13419 12833 13431 12867
rect 13465 12846 13782 12867
rect 13465 12833 13477 12846
rect 13419 12826 13477 12833
rect 13524 12812 13591 12818
rect 3010 12758 3056 12770
rect 8864 12793 8954 12809
rect 8864 12741 8883 12793
rect 8935 12741 8954 12793
rect 13524 12778 13540 12812
rect 13574 12799 13591 12812
rect 13574 12778 13726 12799
rect 13524 12771 13726 12778
rect 8864 12725 8954 12741
rect 13604 12710 13670 12712
rect 13342 12705 13396 12709
rect 2922 12632 2928 12692
rect 2962 12632 2968 12692
rect 2922 12620 2968 12632
rect 3010 12692 3056 12704
rect 13341 12702 13396 12705
rect 3010 12632 3016 12692
rect 3050 12632 3056 12692
rect 13198 12668 13350 12702
rect 13384 12668 13396 12702
rect 13341 12665 13396 12668
rect 13341 12661 13395 12665
rect 13604 12658 13612 12710
rect 13664 12658 13670 12710
rect 13604 12657 13670 12658
rect 2386 12546 2846 12566
rect 2386 12535 2451 12546
rect 2386 12501 2415 12535
rect 2449 12501 2451 12535
rect 2386 12494 2451 12501
rect 2503 12545 2726 12546
rect 2503 12535 2582 12545
rect 2634 12535 2726 12545
rect 2503 12501 2507 12535
rect 2541 12501 2582 12535
rect 2634 12501 2691 12535
rect 2725 12501 2726 12535
rect 2503 12494 2582 12501
rect 2386 12493 2582 12494
rect 2634 12494 2726 12501
rect 2778 12535 2846 12546
rect 2778 12501 2783 12535
rect 2817 12501 2846 12535
rect 2778 12494 2846 12501
rect 2634 12493 2846 12494
rect 2386 12470 2846 12493
rect 2922 12554 2968 12566
rect 2922 12494 2928 12554
rect 2962 12494 2968 12554
rect 2922 12416 2968 12494
rect 3010 12554 3056 12632
rect 8864 12623 8954 12639
rect 8864 12571 8883 12623
rect 8935 12571 8954 12623
rect 13698 12627 13726 12771
rect 13754 12714 13782 12846
rect 13810 12831 13816 12891
rect 13850 12831 13856 12891
rect 13810 12819 13856 12831
rect 13898 12891 14001 12903
rect 13898 12831 13904 12891
rect 13938 12831 14001 12891
rect 19751 12889 19770 12941
rect 19822 12889 19841 12941
rect 19751 12873 19841 12889
rect 20519 12891 20565 12969
rect 20607 13029 20653 13107
rect 26461 13098 26551 13114
rect 26461 13046 26480 13098
rect 26532 13046 26551 13098
rect 26461 13030 26551 13046
rect 20607 12969 20613 13029
rect 20647 12969 20653 13029
rect 20607 12957 20653 12969
rect 26460 12941 26550 12957
rect 13898 12819 14001 12831
rect 20128 12867 20491 12874
rect 20128 12833 20140 12867
rect 20174 12846 20491 12867
rect 20174 12833 20186 12846
rect 20128 12826 20186 12833
rect 13848 12772 13917 12778
rect 13848 12738 13860 12772
rect 13894 12738 13917 12772
rect 13848 12732 13917 12738
rect 13754 12702 13803 12714
rect 13754 12668 13763 12702
rect 13797 12668 13803 12702
rect 13754 12655 13803 12668
rect 13698 12609 13841 12627
rect 13698 12599 13801 12609
rect 8864 12555 8954 12571
rect 10951 12556 11058 12570
rect 11138 12556 11245 12572
rect 11323 12558 11430 12574
rect 11323 12556 11359 12558
rect 3010 12494 3016 12554
rect 3050 12494 3056 12554
rect 10885 12554 11174 12556
rect 10885 12502 10987 12554
rect 11039 12504 11174 12554
rect 11226 12506 11359 12556
rect 11411 12556 11430 12558
rect 11508 12559 11615 12575
rect 11508 12556 11544 12559
rect 11411 12507 11544 12556
rect 11596 12556 11615 12559
rect 11711 12561 11818 12577
rect 11711 12556 11747 12561
rect 11596 12509 11747 12556
rect 11799 12556 11818 12561
rect 11896 12563 12003 12579
rect 11896 12556 11932 12563
rect 11799 12511 11932 12556
rect 11984 12556 12003 12563
rect 12095 12565 12202 12581
rect 12095 12556 12131 12565
rect 11984 12513 12131 12556
rect 12183 12556 12202 12565
rect 12297 12564 12404 12580
rect 12297 12556 12333 12564
rect 12183 12513 12333 12556
rect 11984 12512 12333 12513
rect 12385 12556 12404 12564
rect 12507 12567 12614 12583
rect 12507 12556 12543 12567
rect 12385 12515 12543 12556
rect 12595 12556 12614 12567
rect 12731 12567 12838 12583
rect 12731 12556 12767 12567
rect 12595 12515 12767 12556
rect 12819 12556 12838 12567
rect 12937 12566 13044 12582
rect 12937 12556 12973 12566
rect 12819 12515 12973 12556
rect 12385 12514 12973 12515
rect 13025 12556 13044 12566
rect 13158 12565 13265 12581
rect 13158 12556 13194 12565
rect 13025 12514 13194 12556
rect 12385 12513 13194 12514
rect 13246 12556 13265 12565
rect 13792 12575 13801 12599
rect 13835 12575 13841 12609
rect 13792 12562 13841 12575
rect 13246 12513 13272 12556
rect 12385 12512 13272 12513
rect 11984 12511 13272 12512
rect 11799 12509 13272 12511
rect 11596 12507 13272 12509
rect 11411 12506 13272 12507
rect 11226 12504 13272 12506
rect 11039 12502 13272 12504
rect 10885 12500 13272 12502
rect 3010 12482 3056 12494
rect 10882 12497 13274 12500
rect 8863 12466 8953 12482
rect 2531 12392 2894 12399
rect 2531 12358 2543 12392
rect 2577 12371 2894 12392
rect 2577 12358 2589 12371
rect 2531 12351 2589 12358
rect 2636 12337 2703 12343
rect 2636 12303 2652 12337
rect 2686 12324 2703 12337
rect 2686 12303 2838 12324
rect 2636 12296 2838 12303
rect 2716 12235 2782 12237
rect 2454 12230 2508 12234
rect 2453 12227 2508 12230
rect 2324 12193 2462 12227
rect 2496 12193 2508 12227
rect 2453 12190 2508 12193
rect 2453 12186 2507 12190
rect 2716 12183 2724 12235
rect 2776 12183 2782 12235
rect 2716 12182 2782 12183
rect 2810 12152 2838 12296
rect 2866 12239 2894 12371
rect 2922 12356 2928 12416
rect 2962 12356 2968 12416
rect 2922 12344 2968 12356
rect 3010 12416 3113 12428
rect 3010 12356 3016 12416
rect 3050 12356 3113 12416
rect 8863 12414 8882 12466
rect 8934 12414 8953 12466
rect 8863 12398 8953 12414
rect 10882 12475 13734 12497
rect 10882 12466 13357 12475
rect 13409 12466 13477 12475
rect 13529 12466 13620 12475
rect 13672 12466 13734 12475
rect 10882 12432 10911 12466
rect 10945 12432 11003 12466
rect 11037 12432 11095 12466
rect 11129 12432 11187 12466
rect 11221 12432 11279 12466
rect 11313 12432 11371 12466
rect 11405 12432 11463 12466
rect 11497 12432 11555 12466
rect 11589 12432 11647 12466
rect 11681 12432 11739 12466
rect 11773 12432 11831 12466
rect 11865 12432 11923 12466
rect 11957 12432 12015 12466
rect 12049 12432 12107 12466
rect 12141 12432 12199 12466
rect 12233 12432 12291 12466
rect 12325 12432 12383 12466
rect 12417 12432 12475 12466
rect 12509 12432 12567 12466
rect 12601 12432 12659 12466
rect 12693 12432 12751 12466
rect 12785 12432 12843 12466
rect 12877 12432 12935 12466
rect 12969 12432 13027 12466
rect 13061 12432 13119 12466
rect 13153 12432 13211 12466
rect 13245 12432 13303 12466
rect 13337 12432 13357 12466
rect 13429 12432 13477 12466
rect 13529 12432 13579 12466
rect 13613 12432 13620 12466
rect 13705 12432 13734 12466
rect 10882 12423 13357 12432
rect 13409 12423 13477 12432
rect 13529 12423 13620 12432
rect 13672 12423 13734 12432
rect 10882 12401 13734 12423
rect 3010 12344 3113 12356
rect 2960 12297 3029 12303
rect 2960 12263 2972 12297
rect 3006 12263 3029 12297
rect 2960 12257 3029 12263
rect 2866 12227 2915 12239
rect 2866 12193 2875 12227
rect 2909 12193 2915 12227
rect 2866 12180 2915 12193
rect 2810 12134 2953 12152
rect 2810 12124 2913 12134
rect 2904 12100 2913 12124
rect 2947 12100 2953 12134
rect 2904 12087 2953 12100
rect 2386 12000 2846 12022
rect 2386 11991 2469 12000
rect 2521 11991 2589 12000
rect 2641 11991 2732 12000
rect 2784 11991 2846 12000
rect 2386 11957 2415 11991
rect 2449 11957 2469 11991
rect 2541 11957 2589 11991
rect 2641 11957 2691 11991
rect 2725 11957 2732 11991
rect 2817 11957 2846 11991
rect 2386 11948 2469 11957
rect 2521 11948 2589 11957
rect 2641 11948 2732 11957
rect 2784 11948 2846 11957
rect 2386 11926 2846 11948
rect 2981 11857 3029 12257
rect 2330 11810 3029 11857
rect 2981 11669 3029 11810
rect 2971 11663 3029 11669
rect 2730 11657 2795 11658
rect 2730 11656 2736 11657
rect 2634 11654 2736 11656
rect 2632 11608 2736 11654
rect 2730 11605 2736 11608
rect 2788 11605 2795 11657
rect 2971 11629 2983 11663
rect 3017 11629 3029 11663
rect 2971 11623 3029 11629
rect 3067 11854 3113 12344
rect 13205 12332 13269 12340
rect 13869 12332 13917 12732
rect 13205 12324 13917 12332
rect 11632 12311 11696 12312
rect 9061 12276 9338 12299
rect 8781 12224 8871 12240
rect 8781 12213 8800 12224
rect 8706 12172 8800 12213
rect 8852 12172 8871 12224
rect 3163 12157 3212 12164
rect 3163 12152 3782 12157
rect 3163 12118 3172 12152
rect 3206 12118 3782 12152
rect 3163 12110 3782 12118
rect 3163 12105 3212 12110
rect 3164 12063 3213 12071
rect 3733 12063 3782 12110
rect 8706 12154 8871 12172
rect 9061 12224 9177 12276
rect 9229 12224 9338 12276
rect 11084 12296 11142 12302
rect 11084 12262 11096 12296
rect 11130 12293 11142 12296
rect 11448 12296 11506 12302
rect 11448 12293 11460 12296
rect 11130 12265 11460 12293
rect 11130 12262 11142 12265
rect 11084 12256 11142 12262
rect 11448 12262 11460 12265
rect 11494 12262 11506 12296
rect 11448 12256 11506 12262
rect 11632 12259 11638 12311
rect 11690 12293 11696 12311
rect 12372 12296 12430 12302
rect 12372 12293 12384 12296
rect 11690 12265 12384 12293
rect 11690 12259 11696 12265
rect 12372 12262 12384 12265
rect 12418 12262 12430 12296
rect 13205 12290 13221 12324
rect 13255 12290 13917 12324
rect 13205 12285 13917 12290
rect 13205 12276 13269 12285
rect 11636 12256 11694 12259
rect 12372 12256 12430 12262
rect 10876 12233 10964 12234
rect 9061 12175 9338 12224
rect 10869 12217 10964 12233
rect 10869 12183 10912 12217
rect 10946 12183 10964 12217
rect 11467 12225 11506 12256
rect 12096 12228 12154 12234
rect 12096 12225 12108 12228
rect 11467 12197 12108 12225
rect 9061 12158 9337 12175
rect 10869 12169 10964 12183
rect 8706 12108 8753 12154
rect 9061 12124 9090 12158
rect 9124 12124 9182 12158
rect 9216 12124 9274 12158
rect 9308 12124 9337 12158
rect 11248 12145 11256 12197
rect 11308 12145 11314 12197
rect 12096 12194 12108 12197
rect 12142 12194 12154 12228
rect 12096 12188 12154 12194
rect 12753 12186 12759 12239
rect 12811 12186 12817 12239
rect 12753 12185 12817 12186
rect 12004 12160 12062 12166
rect 8707 12105 8753 12108
rect 3164 12059 3665 12063
rect 3164 12025 3173 12059
rect 3207 12054 3665 12059
rect 3207 12025 3614 12054
rect 3164 12020 3614 12025
rect 3648 12020 3665 12054
rect 3164 12017 3665 12020
rect 3733 12057 8154 12063
rect 3733 12023 4346 12057
rect 4380 12023 4472 12057
rect 4506 12023 5558 12057
rect 5592 12023 5684 12057
rect 5718 12023 6770 12057
rect 6804 12023 6896 12057
rect 6930 12023 7982 12057
rect 8016 12023 8108 12057
rect 8142 12023 8154 12057
rect 8707 12045 8713 12105
rect 8747 12045 8753 12105
rect 8707 12033 8753 12045
rect 8795 12105 8841 12117
rect 8795 12045 8801 12105
rect 8835 12045 8841 12105
rect 9061 12093 9337 12124
rect 12004 12126 12016 12160
rect 12050 12157 12062 12160
rect 12648 12160 12706 12166
rect 12648 12157 12660 12160
rect 12050 12129 12660 12157
rect 12050 12126 12062 12129
rect 12004 12120 12062 12126
rect 12648 12126 12660 12129
rect 12694 12126 12706 12160
rect 13869 12144 13917 12285
rect 13859 12138 13917 12144
rect 13618 12132 13683 12133
rect 13618 12131 13624 12132
rect 13522 12129 13624 12131
rect 12648 12120 12706 12126
rect 10992 12092 11050 12098
rect 10992 12058 11004 12092
rect 11038 12089 11050 12092
rect 11360 12092 11418 12098
rect 11360 12089 11372 12092
rect 11038 12061 11372 12089
rect 11038 12058 11050 12061
rect 10992 12052 11050 12058
rect 11360 12058 11372 12061
rect 11406 12089 11418 12092
rect 12096 12092 12154 12098
rect 12096 12089 12108 12092
rect 11406 12061 12108 12089
rect 11406 12058 11418 12061
rect 11360 12052 11418 12058
rect 12096 12058 12108 12061
rect 12142 12058 12154 12092
rect 13520 12083 13624 12129
rect 13618 12080 13624 12083
rect 13676 12080 13683 12132
rect 13859 12104 13871 12138
rect 13905 12104 13917 12138
rect 13859 12098 13917 12104
rect 13955 12329 14001 12819
rect 20233 12812 20300 12818
rect 20233 12778 20249 12812
rect 20283 12799 20300 12812
rect 20283 12778 20435 12799
rect 20233 12771 20435 12778
rect 19669 12699 19759 12715
rect 20313 12710 20379 12712
rect 20051 12705 20105 12709
rect 20050 12702 20105 12705
rect 19669 12688 19688 12699
rect 19594 12647 19688 12688
rect 19740 12647 19759 12699
rect 19914 12668 20059 12702
rect 20093 12668 20105 12702
rect 20050 12665 20105 12668
rect 20050 12661 20104 12665
rect 20313 12658 20321 12710
rect 20373 12658 20379 12710
rect 20313 12657 20379 12658
rect 14051 12632 14100 12639
rect 14051 12627 14670 12632
rect 14051 12593 14060 12627
rect 14094 12593 14670 12627
rect 14051 12585 14670 12593
rect 14051 12580 14100 12585
rect 14052 12538 14101 12546
rect 14621 12538 14670 12585
rect 19594 12629 19759 12647
rect 19594 12583 19641 12629
rect 20407 12627 20435 12771
rect 20463 12714 20491 12846
rect 20519 12831 20525 12891
rect 20559 12831 20565 12891
rect 20519 12819 20565 12831
rect 20607 12891 20710 12903
rect 20607 12831 20613 12891
rect 20647 12831 20710 12891
rect 26460 12889 26479 12941
rect 26531 12889 26550 12941
rect 26460 12873 26550 12889
rect 20607 12819 20710 12831
rect 20557 12772 20626 12778
rect 20557 12738 20569 12772
rect 20603 12738 20626 12772
rect 20557 12732 20626 12738
rect 20463 12702 20512 12714
rect 20463 12668 20472 12702
rect 20506 12668 20512 12702
rect 20463 12655 20512 12668
rect 20407 12609 20550 12627
rect 20407 12599 20510 12609
rect 19595 12580 19641 12583
rect 14052 12534 14553 12538
rect 14052 12500 14061 12534
rect 14095 12529 14553 12534
rect 14095 12500 14502 12529
rect 14052 12495 14502 12500
rect 14536 12495 14553 12529
rect 14052 12492 14553 12495
rect 14621 12532 19042 12538
rect 14621 12498 15234 12532
rect 15268 12498 15360 12532
rect 15394 12498 16446 12532
rect 16480 12498 16572 12532
rect 16606 12498 17658 12532
rect 17692 12498 17784 12532
rect 17818 12498 18870 12532
rect 18904 12498 18996 12532
rect 19030 12498 19042 12532
rect 19595 12520 19601 12580
rect 19635 12520 19641 12580
rect 19595 12508 19641 12520
rect 19683 12580 19729 12592
rect 19683 12520 19689 12580
rect 19723 12520 19729 12580
rect 20501 12575 20510 12599
rect 20544 12575 20550 12609
rect 20501 12562 20550 12575
rect 19683 12511 19729 12520
rect 14621 12492 19042 12498
rect 14052 12491 14548 12492
rect 14621 12491 15067 12492
rect 14052 12487 14101 12491
rect 14490 12489 14548 12491
rect 19683 12482 19921 12511
rect 14452 12440 14498 12448
rect 14429 12439 14508 12440
rect 14429 12375 14436 12439
rect 14500 12375 14508 12439
rect 14540 12439 14586 12451
rect 15184 12443 15230 12451
rect 14540 12379 14546 12439
rect 14580 12379 14586 12439
rect 14452 12364 14498 12375
rect 14540 12329 14586 12379
rect 15161 12442 15240 12443
rect 15161 12378 15168 12442
rect 15232 12378 15240 12442
rect 15289 12439 15335 12451
rect 15398 12443 15444 12451
rect 16396 12443 16442 12451
rect 15289 12379 15295 12439
rect 15329 12379 15335 12439
rect 15184 12367 15230 12378
rect 15289 12329 15335 12379
rect 15388 12442 15467 12443
rect 15388 12378 15396 12442
rect 15460 12378 15467 12442
rect 16373 12442 16452 12443
rect 16373 12378 16380 12442
rect 16444 12378 16452 12442
rect 16500 12439 16546 12451
rect 16610 12443 16656 12451
rect 17608 12443 17654 12451
rect 16500 12379 16506 12439
rect 16540 12379 16546 12439
rect 15398 12367 15444 12378
rect 16396 12367 16442 12378
rect 16500 12329 16546 12379
rect 16600 12442 16679 12443
rect 16600 12378 16608 12442
rect 16672 12378 16679 12442
rect 17585 12442 17664 12443
rect 17585 12378 17592 12442
rect 17656 12378 17664 12442
rect 17713 12439 17759 12451
rect 17822 12443 17868 12451
rect 18820 12443 18866 12451
rect 17713 12379 17719 12439
rect 17753 12379 17759 12439
rect 16610 12367 16656 12378
rect 17608 12367 17654 12378
rect 17713 12329 17759 12379
rect 17812 12442 17891 12443
rect 17812 12378 17820 12442
rect 17884 12378 17891 12442
rect 18797 12442 18876 12443
rect 18797 12378 18804 12442
rect 18868 12378 18876 12442
rect 18927 12439 18973 12451
rect 19034 12443 19080 12451
rect 18927 12379 18933 12439
rect 18967 12379 18973 12439
rect 17822 12367 17868 12378
rect 18820 12367 18866 12378
rect 18927 12329 18973 12379
rect 19024 12442 19103 12443
rect 19024 12378 19032 12442
rect 19096 12378 19103 12442
rect 19595 12442 19641 12454
rect 19595 12382 19601 12442
rect 19635 12382 19641 12442
rect 19034 12367 19080 12378
rect 19595 12370 19641 12382
rect 19683 12442 19729 12482
rect 19683 12382 19689 12442
rect 19723 12382 19729 12442
rect 19683 12370 19729 12382
rect 19757 12442 19847 12454
rect 19757 12438 19785 12442
rect 19819 12438 19847 12442
rect 19757 12386 19776 12438
rect 19828 12386 19847 12438
rect 19757 12382 19785 12386
rect 19819 12382 19847 12386
rect 19757 12370 19847 12382
rect 19875 12442 19921 12482
rect 19875 12382 19881 12442
rect 19915 12382 19921 12442
rect 19983 12475 20443 12497
rect 19983 12466 20066 12475
rect 20118 12466 20186 12475
rect 20238 12466 20329 12475
rect 20381 12466 20443 12475
rect 19983 12432 20012 12466
rect 20046 12432 20066 12466
rect 20138 12432 20186 12466
rect 20238 12432 20288 12466
rect 20322 12432 20329 12466
rect 20414 12432 20443 12466
rect 19983 12423 20066 12432
rect 20118 12423 20186 12432
rect 20238 12423 20329 12432
rect 20381 12423 20443 12432
rect 19983 12401 20443 12423
rect 19875 12370 19921 12382
rect 19514 12329 19580 12331
rect 13955 12325 19580 12329
rect 13955 12291 19530 12325
rect 19564 12291 19580 12325
rect 13955 12287 19580 12291
rect 13955 12066 14001 12287
rect 14805 12240 14851 12250
rect 14783 12176 14792 12240
rect 14856 12176 14865 12240
rect 14783 12175 14865 12176
rect 14895 12238 14941 12287
rect 15537 12240 15583 12250
rect 14895 12178 14901 12238
rect 14935 12178 14941 12238
rect 14805 12166 14851 12175
rect 14895 12166 14941 12178
rect 15515 12176 15524 12240
rect 15588 12176 15597 12240
rect 15515 12175 15597 12176
rect 15644 12238 15690 12287
rect 15747 12240 15793 12250
rect 16749 12240 16795 12250
rect 15644 12178 15650 12238
rect 15684 12178 15690 12238
rect 15537 12166 15583 12175
rect 15644 12166 15690 12178
rect 15733 12176 15742 12240
rect 15806 12176 15815 12240
rect 15733 12175 15815 12176
rect 16727 12176 16736 12240
rect 16800 12176 16809 12240
rect 16727 12175 16809 12176
rect 16855 12238 16901 12287
rect 16959 12240 17005 12250
rect 18087 12240 18133 12250
rect 16855 12178 16861 12238
rect 16895 12178 16901 12238
rect 15747 12166 15793 12175
rect 16749 12166 16795 12175
rect 16855 12166 16901 12178
rect 16945 12176 16954 12240
rect 17018 12176 17027 12240
rect 16945 12175 17027 12176
rect 18065 12176 18074 12240
rect 18138 12176 18147 12240
rect 18065 12175 18147 12176
rect 18195 12238 18241 12287
rect 18297 12240 18343 12250
rect 18195 12178 18201 12238
rect 18235 12178 18241 12238
rect 16959 12166 17005 12175
rect 18087 12166 18133 12175
rect 18195 12166 18241 12178
rect 18283 12176 18292 12240
rect 18356 12176 18365 12240
rect 18283 12175 18365 12176
rect 18942 12238 18988 12287
rect 19518 12285 19580 12287
rect 19613 12322 19641 12370
rect 20578 12332 20626 12732
rect 19897 12329 20626 12332
rect 19725 12323 20626 12329
rect 19725 12322 19737 12323
rect 19613 12293 19737 12322
rect 19613 12251 19641 12293
rect 19725 12289 19737 12293
rect 19771 12289 20626 12323
rect 19725 12285 20626 12289
rect 19725 12283 19967 12285
rect 19897 12280 19967 12283
rect 19031 12240 19077 12250
rect 18942 12178 18948 12238
rect 18982 12178 18988 12238
rect 18297 12166 18343 12175
rect 18942 12166 18988 12178
rect 19017 12176 19026 12240
rect 19090 12176 19099 12240
rect 19017 12175 19099 12176
rect 19595 12239 19641 12251
rect 19595 12179 19601 12239
rect 19635 12179 19641 12239
rect 19031 12166 19077 12175
rect 19595 12167 19641 12179
rect 19683 12239 19729 12251
rect 19683 12179 19689 12239
rect 19723 12179 19729 12239
rect 19683 12139 19729 12179
rect 19757 12239 19847 12251
rect 19757 12235 19785 12239
rect 19819 12235 19847 12239
rect 19757 12183 19776 12235
rect 19828 12183 19847 12235
rect 19757 12179 19785 12183
rect 19819 12179 19847 12183
rect 19757 12167 19847 12179
rect 19875 12239 19921 12251
rect 19875 12179 19881 12239
rect 19915 12179 19921 12239
rect 19875 12139 19921 12179
rect 20578 12144 20626 12285
rect 18983 12134 19042 12137
rect 14105 12080 14112 12132
rect 14164 12130 14170 12132
rect 14843 12130 14901 12134
rect 14164 12128 14901 12130
rect 14164 12094 14855 12128
rect 14889 12113 14901 12128
rect 15575 12128 16971 12134
rect 14889 12094 14903 12113
rect 14164 12083 14903 12094
rect 15575 12094 15587 12128
rect 15621 12094 15709 12128
rect 15743 12094 16799 12128
rect 16833 12094 16921 12128
rect 16955 12094 16971 12128
rect 15575 12088 16971 12094
rect 18125 12128 18309 12134
rect 18125 12094 18137 12128
rect 18171 12094 18259 12128
rect 18293 12094 18309 12128
rect 18125 12088 18309 12094
rect 18981 12128 19042 12134
rect 18981 12094 18993 12128
rect 19027 12094 19042 12128
rect 18981 12088 19042 12094
rect 14164 12080 14170 12083
rect 14105 12079 14170 12080
rect 14845 12078 14903 12083
rect 12096 12052 12154 12058
rect 13785 12054 13831 12066
rect 8795 12036 8841 12045
rect 3733 12017 8154 12023
rect 3164 12016 3660 12017
rect 3733 12016 4179 12017
rect 3164 12012 3213 12016
rect 3602 12014 3660 12016
rect 8795 12007 9033 12036
rect 3564 11965 3610 11973
rect 3541 11964 3620 11965
rect 3541 11900 3548 11964
rect 3612 11900 3620 11964
rect 3652 11964 3698 11976
rect 4296 11968 4342 11976
rect 3652 11904 3658 11964
rect 3692 11904 3698 11964
rect 3564 11889 3610 11900
rect 3652 11854 3698 11904
rect 4273 11967 4352 11968
rect 4273 11903 4280 11967
rect 4344 11903 4352 11967
rect 4401 11964 4447 11976
rect 4510 11968 4556 11976
rect 5508 11968 5554 11976
rect 4401 11904 4407 11964
rect 4441 11904 4447 11964
rect 4296 11892 4342 11903
rect 4401 11854 4447 11904
rect 4500 11967 4579 11968
rect 4500 11903 4508 11967
rect 4572 11903 4579 11967
rect 5485 11967 5564 11968
rect 5485 11903 5492 11967
rect 5556 11903 5564 11967
rect 5612 11964 5658 11976
rect 5722 11968 5768 11976
rect 6720 11968 6766 11976
rect 5612 11904 5618 11964
rect 5652 11904 5658 11964
rect 4510 11892 4556 11903
rect 5508 11892 5554 11903
rect 5612 11854 5658 11904
rect 5712 11967 5791 11968
rect 5712 11903 5720 11967
rect 5784 11903 5791 11967
rect 6697 11967 6776 11968
rect 6697 11903 6704 11967
rect 6768 11903 6776 11967
rect 6825 11964 6871 11976
rect 6934 11968 6980 11976
rect 7932 11968 7978 11976
rect 6825 11904 6831 11964
rect 6865 11904 6871 11964
rect 5722 11892 5768 11903
rect 6720 11892 6766 11903
rect 6825 11854 6871 11904
rect 6924 11967 7003 11968
rect 6924 11903 6932 11967
rect 6996 11903 7003 11967
rect 7909 11967 7988 11968
rect 7909 11903 7916 11967
rect 7980 11903 7988 11967
rect 8039 11964 8085 11976
rect 8146 11968 8192 11976
rect 8039 11904 8045 11964
rect 8079 11904 8085 11964
rect 6934 11892 6980 11903
rect 7932 11892 7978 11903
rect 8039 11854 8085 11904
rect 8136 11967 8215 11968
rect 8136 11903 8144 11967
rect 8208 11903 8215 11967
rect 8707 11967 8753 11979
rect 8707 11907 8713 11967
rect 8747 11907 8753 11967
rect 8146 11892 8192 11903
rect 8707 11895 8753 11907
rect 8795 11967 8841 12007
rect 8795 11907 8801 11967
rect 8835 11907 8841 11967
rect 8795 11895 8841 11907
rect 8869 11967 8959 11979
rect 8869 11963 8897 11967
rect 8931 11963 8959 11967
rect 8869 11911 8888 11963
rect 8940 11911 8959 11963
rect 8869 11907 8897 11911
rect 8931 11907 8959 11911
rect 8869 11895 8959 11907
rect 8987 11967 9033 12007
rect 11258 11981 11264 12033
rect 11317 12022 11324 12033
rect 12922 12026 12983 12037
rect 12922 12022 12935 12026
rect 11317 11994 12935 12022
rect 11317 11981 11324 11994
rect 12922 11992 12935 11994
rect 12969 11992 12983 12026
rect 13199 12002 13205 12054
rect 13257 12002 13263 12054
rect 12922 11985 12983 11992
rect 13785 11994 13791 12054
rect 13825 11994 13831 12054
rect 8987 11907 8993 11967
rect 9027 11907 9033 11967
rect 8987 11895 9033 11907
rect 10882 11922 13274 11953
rect 8626 11854 8692 11856
rect 3067 11850 8692 11854
rect 3067 11816 8642 11850
rect 8676 11816 8692 11850
rect 3067 11812 8692 11816
rect 3067 11591 3113 11812
rect 3917 11765 3963 11775
rect 3895 11701 3904 11765
rect 3968 11701 3977 11765
rect 3895 11700 3977 11701
rect 4007 11763 4053 11812
rect 4649 11765 4695 11775
rect 4007 11703 4013 11763
rect 4047 11703 4053 11763
rect 3917 11691 3963 11700
rect 4007 11691 4053 11703
rect 4627 11701 4636 11765
rect 4700 11701 4709 11765
rect 4627 11700 4709 11701
rect 4756 11763 4802 11812
rect 4859 11765 4905 11775
rect 5861 11765 5907 11775
rect 4756 11703 4762 11763
rect 4796 11703 4802 11763
rect 4649 11691 4695 11700
rect 4756 11691 4802 11703
rect 4845 11701 4854 11765
rect 4918 11701 4927 11765
rect 4845 11700 4927 11701
rect 5839 11701 5848 11765
rect 5912 11701 5921 11765
rect 5839 11700 5921 11701
rect 5967 11763 6013 11812
rect 6071 11765 6117 11775
rect 7199 11765 7245 11775
rect 5967 11703 5973 11763
rect 6007 11703 6013 11763
rect 4859 11691 4905 11700
rect 5861 11691 5907 11700
rect 5967 11691 6013 11703
rect 6057 11701 6066 11765
rect 6130 11701 6139 11765
rect 6057 11700 6139 11701
rect 7177 11701 7186 11765
rect 7250 11701 7259 11765
rect 7177 11700 7259 11701
rect 7307 11763 7353 11812
rect 7409 11765 7455 11775
rect 7307 11703 7313 11763
rect 7347 11703 7353 11763
rect 6071 11691 6117 11700
rect 7199 11691 7245 11700
rect 7307 11691 7353 11703
rect 7395 11701 7404 11765
rect 7468 11701 7477 11765
rect 7395 11700 7477 11701
rect 8054 11763 8100 11812
rect 8630 11810 8692 11812
rect 8725 11847 8753 11895
rect 10882 11888 10911 11922
rect 10945 11888 11003 11922
rect 11037 11888 11095 11922
rect 11129 11888 11187 11922
rect 11221 11888 11279 11922
rect 11313 11888 11371 11922
rect 11405 11888 11463 11922
rect 11497 11888 11555 11922
rect 11589 11888 11647 11922
rect 11681 11888 11739 11922
rect 11773 11888 11831 11922
rect 11865 11888 11923 11922
rect 11957 11888 12015 11922
rect 12049 11888 12107 11922
rect 12141 11888 12199 11922
rect 12233 11888 12291 11922
rect 12325 11888 12383 11922
rect 12417 11888 12475 11922
rect 12509 11888 12567 11922
rect 12601 11888 12659 11922
rect 12693 11888 12751 11922
rect 12785 11888 12843 11922
rect 12877 11888 12935 11922
rect 12969 11888 13027 11922
rect 13061 11888 13119 11922
rect 13153 11888 13211 11922
rect 13245 11888 13274 11922
rect 10882 11885 13274 11888
rect 10882 11882 11117 11885
rect 9030 11854 9180 11856
rect 8837 11850 9180 11854
rect 8837 11848 9134 11850
rect 8837 11847 8849 11848
rect 8725 11818 8849 11847
rect 8725 11776 8753 11818
rect 8837 11814 8849 11818
rect 8883 11816 9134 11848
rect 9168 11816 9180 11850
rect 8883 11814 9180 11816
rect 8837 11808 9180 11814
rect 9224 11854 9276 11857
rect 10291 11854 10298 11862
rect 9224 11849 10298 11854
rect 9224 11815 9236 11849
rect 9270 11815 10298 11849
rect 9224 11812 10298 11815
rect 9224 11809 9276 11812
rect 10291 11808 10298 11812
rect 10352 11808 10359 11862
rect 10882 11829 10917 11882
rect 10970 11832 11117 11882
rect 11170 11883 13274 11885
rect 11170 11832 11353 11883
rect 10970 11830 11353 11832
rect 11406 11879 13274 11883
rect 11406 11878 12364 11879
rect 11406 11877 11987 11878
rect 11406 11830 11786 11877
rect 10970 11829 11786 11830
rect 10882 11826 11786 11829
rect 10882 11792 10911 11826
rect 10945 11792 11003 11826
rect 11037 11792 11095 11826
rect 11129 11792 11187 11826
rect 11221 11792 11279 11826
rect 11313 11792 11371 11826
rect 11405 11824 11786 11826
rect 11839 11825 11987 11877
rect 12040 11876 12364 11878
rect 12040 11825 12173 11876
rect 11839 11824 12173 11825
rect 11405 11823 12173 11824
rect 12226 11826 12364 11876
rect 12417 11878 13274 11879
rect 12417 11826 12577 11878
rect 12226 11825 12577 11826
rect 12630 11857 13274 11878
rect 13785 11916 13831 11994
rect 13945 12054 14001 12066
rect 13945 11994 13951 12054
rect 13985 11994 14001 12054
rect 13945 11982 14001 11994
rect 12630 11825 12723 11857
rect 13785 11856 13791 11916
rect 13825 11856 13831 11916
rect 13785 11844 13831 11856
rect 13945 11916 13991 11928
rect 13945 11856 13951 11916
rect 13985 11856 13991 11916
rect 12226 11823 12723 11825
rect 11405 11792 12723 11823
rect 8143 11765 8189 11775
rect 8054 11703 8060 11763
rect 8094 11703 8100 11763
rect 7409 11691 7455 11700
rect 8054 11691 8100 11703
rect 8129 11701 8138 11765
rect 8202 11701 8211 11765
rect 8129 11700 8211 11701
rect 8707 11764 8753 11776
rect 8707 11704 8713 11764
rect 8747 11704 8753 11764
rect 8143 11691 8189 11700
rect 8707 11692 8753 11704
rect 8795 11764 8841 11776
rect 8795 11704 8801 11764
rect 8835 11704 8841 11764
rect 8795 11664 8841 11704
rect 8869 11764 8959 11776
rect 8869 11760 8897 11764
rect 8931 11760 8959 11764
rect 8869 11708 8888 11760
rect 8940 11708 8959 11760
rect 8869 11704 8897 11708
rect 8931 11704 8959 11708
rect 8869 11692 8959 11704
rect 8987 11764 9033 11776
rect 8987 11704 8993 11764
rect 9027 11704 9033 11764
rect 10882 11761 12723 11792
rect 13785 11778 13831 11790
rect 12755 11733 12761 11745
rect 8987 11664 9033 11704
rect 11307 11727 12761 11733
rect 11307 11693 11319 11727
rect 11353 11705 12761 11727
rect 11353 11693 11366 11705
rect 12755 11693 12761 11705
rect 12813 11693 12819 11745
rect 13785 11718 13791 11778
rect 13825 11718 13831 11778
rect 11307 11685 11366 11693
rect 8095 11659 8154 11662
rect 3217 11605 3224 11657
rect 3276 11655 3282 11657
rect 3955 11655 4013 11659
rect 3276 11653 4013 11655
rect 3276 11619 3967 11653
rect 4001 11638 4013 11653
rect 4687 11653 6083 11659
rect 4001 11619 4015 11638
rect 3276 11608 4015 11619
rect 4687 11619 4699 11653
rect 4733 11619 4821 11653
rect 4855 11619 5911 11653
rect 5945 11619 6033 11653
rect 6067 11619 6083 11653
rect 4687 11613 6083 11619
rect 7237 11653 7421 11659
rect 7237 11619 7249 11653
rect 7283 11619 7371 11653
rect 7405 11619 7421 11653
rect 7237 11613 7421 11619
rect 8093 11653 8154 11659
rect 8093 11619 8105 11653
rect 8139 11619 8154 11653
rect 8093 11613 8154 11619
rect 3276 11605 3282 11608
rect 3217 11604 3282 11605
rect 3957 11603 4015 11608
rect 2897 11579 2943 11591
rect 2897 11519 2903 11579
rect 2937 11519 2943 11579
rect 2897 11441 2943 11519
rect 3057 11579 3113 11591
rect 3057 11519 3063 11579
rect 3097 11519 3113 11579
rect 3057 11507 3113 11519
rect 2897 11381 2903 11441
rect 2937 11381 2943 11441
rect 2897 11369 2943 11381
rect 3057 11441 3103 11453
rect 3057 11381 3063 11441
rect 3097 11381 3103 11441
rect 2897 11303 2943 11315
rect 2897 11243 2903 11303
rect 2937 11243 2943 11303
rect 2897 11165 2943 11243
rect 3057 11303 3103 11381
rect 3057 11243 3063 11303
rect 3097 11243 3103 11303
rect 3057 11231 3103 11243
rect 2897 11105 2903 11165
rect 2937 11105 2943 11165
rect 2897 11093 2943 11105
rect 3057 11165 3103 11177
rect 3057 11105 3063 11165
rect 3097 11105 3103 11165
rect 2897 11027 2943 11039
rect 2897 10967 2903 11027
rect 2937 10967 2943 11027
rect 2897 10889 2943 10967
rect 3057 11027 3103 11105
rect 3057 10967 3063 11027
rect 3097 10967 3103 11027
rect 3057 10955 3103 10967
rect 2897 10829 2903 10889
rect 2937 10829 2943 10889
rect 2897 10817 2943 10829
rect 3057 10889 3103 10901
rect 3057 10829 3063 10889
rect 3097 10829 3103 10889
rect 2897 10751 2943 10763
rect 2897 10691 2903 10751
rect 2937 10691 2943 10751
rect 2897 10613 2943 10691
rect 3057 10751 3103 10829
rect 3057 10691 3063 10751
rect 3097 10691 3103 10751
rect 3057 10679 3103 10691
rect 2897 10553 2903 10613
rect 2937 10553 2943 10613
rect 3057 10613 3103 10625
rect 3057 10589 3063 10613
rect 2897 10541 2943 10553
rect 3018 10573 3063 10589
rect 3097 10589 3103 10613
rect 3097 10573 3125 10589
rect 3018 10521 3054 10573
rect 3106 10521 3125 10573
rect 3018 10505 3125 10521
rect 3578 10576 3910 10582
rect 3578 10524 3596 10576
rect 3648 10524 3676 10576
rect 3728 10524 3756 10576
rect 3808 10524 3836 10576
rect 3888 10524 3910 10576
rect 3578 10514 3910 10524
rect 4310 10576 4642 10582
rect 4310 10524 4328 10576
rect 4380 10524 4408 10576
rect 4460 10524 4488 10576
rect 4540 10524 4568 10576
rect 4620 10524 4642 10576
rect 4310 10514 4642 10524
rect 4813 10477 4871 11613
rect 4912 10576 5244 10582
rect 4912 10524 4934 10576
rect 4986 10524 5014 10576
rect 5066 10524 5094 10576
rect 5146 10524 5174 10576
rect 5226 10524 5244 10576
rect 4912 10514 5244 10524
rect 5522 10576 5854 10582
rect 5522 10524 5540 10576
rect 5592 10524 5620 10576
rect 5672 10524 5700 10576
rect 5752 10524 5780 10576
rect 5832 10524 5854 10576
rect 5522 10514 5854 10524
rect 6124 10576 6456 10582
rect 6124 10524 6146 10576
rect 6198 10524 6226 10576
rect 6278 10524 6306 10576
rect 6358 10524 6386 10576
rect 6438 10524 6456 10576
rect 6124 10514 6456 10524
rect 6860 10576 7192 10582
rect 6860 10524 6878 10576
rect 6930 10524 6958 10576
rect 7010 10524 7038 10576
rect 7090 10524 7118 10576
rect 7170 10524 7192 10576
rect 6860 10514 7192 10524
rect 2930 10449 4871 10477
rect 7239 10421 7297 11613
rect 7462 10576 7794 10582
rect 7462 10524 7484 10576
rect 7536 10524 7564 10576
rect 7616 10524 7644 10576
rect 7696 10524 7724 10576
rect 7776 10524 7794 10576
rect 7462 10514 7794 10524
rect 2931 10393 7297 10421
rect 8095 10365 8154 11613
rect 8707 11626 8753 11638
rect 8707 11566 8713 11626
rect 8747 11566 8753 11626
rect 8707 11514 8753 11566
rect 8795 11635 9033 11664
rect 11030 11651 11090 11658
rect 8795 11626 8841 11635
rect 8795 11566 8801 11626
rect 8835 11566 8841 11626
rect 8795 11554 8841 11566
rect 9061 11614 9337 11645
rect 9061 11580 9090 11614
rect 9124 11580 9182 11614
rect 9216 11580 9274 11614
rect 9308 11580 9337 11614
rect 11030 11617 11044 11651
rect 11078 11648 11090 11651
rect 11628 11648 11634 11672
rect 11078 11620 11634 11648
rect 11686 11620 11692 11672
rect 13785 11640 13831 11718
rect 13945 11778 13991 11856
rect 13945 11718 13951 11778
rect 13985 11718 13991 11778
rect 13945 11706 13991 11718
rect 11078 11617 11090 11620
rect 11030 11603 11090 11617
rect 9061 11561 9337 11580
rect 13300 11594 13398 11609
rect 9061 11549 9340 11561
rect 9063 11519 9340 11549
rect 13300 11538 13317 11594
rect 13377 11538 13398 11594
rect 13785 11580 13791 11640
rect 13825 11580 13831 11640
rect 13785 11568 13831 11580
rect 13945 11640 13991 11652
rect 13945 11580 13951 11640
rect 13985 11580 13991 11640
rect 8707 11498 8868 11514
rect 8707 11446 8797 11498
rect 8849 11446 8868 11498
rect 8707 11430 8868 11446
rect 9063 11467 9200 11519
rect 9252 11467 9340 11519
rect 9063 11437 9340 11467
rect 10914 11530 11009 11531
rect 10914 11529 11232 11530
rect 10914 11522 11283 11529
rect 10914 11488 10957 11522
rect 10991 11517 11283 11522
rect 13300 11519 13398 11538
rect 10991 11488 11228 11517
rect 10914 11483 11228 11488
rect 11262 11483 11283 11517
rect 10914 11471 11283 11483
rect 13785 11502 13831 11514
rect 10914 11313 11232 11471
rect 13785 11442 13791 11502
rect 13825 11442 13831 11502
rect 13785 11364 13831 11442
rect 13945 11502 13991 11580
rect 13945 11442 13951 11502
rect 13985 11442 13991 11502
rect 13945 11430 13991 11442
rect 10882 11282 11434 11313
rect 13785 11304 13791 11364
rect 13825 11304 13831 11364
rect 13785 11292 13831 11304
rect 13945 11364 13991 11376
rect 13945 11304 13951 11364
rect 13985 11304 13991 11364
rect 10882 11248 10911 11282
rect 10945 11257 11003 11282
rect 10987 11248 11003 11257
rect 11037 11248 11095 11282
rect 11129 11254 11187 11282
rect 11175 11248 11187 11254
rect 11221 11248 11279 11282
rect 11313 11252 11371 11282
rect 11313 11248 11320 11252
rect 11405 11248 11434 11282
rect 10882 11217 10935 11248
rect 10899 11205 10935 11217
rect 10987 11217 11123 11248
rect 10987 11214 11037 11217
rect 10987 11205 11006 11214
rect 10899 11189 11006 11205
rect 11087 11202 11123 11217
rect 11175 11217 11320 11248
rect 11175 11214 11221 11217
rect 11279 11214 11320 11217
rect 11175 11202 11194 11214
rect 11087 11186 11194 11202
rect 11284 11200 11320 11214
rect 11372 11217 11434 11248
rect 13785 11226 13831 11238
rect 11372 11214 11405 11217
rect 11372 11200 11391 11214
rect 11284 11184 11391 11200
rect 13785 11166 13791 11226
rect 13825 11166 13831 11226
rect 13785 11088 13831 11166
rect 13945 11226 13991 11304
rect 13945 11166 13951 11226
rect 13985 11166 13991 11226
rect 13945 11154 13991 11166
rect 13785 11028 13791 11088
rect 13825 11028 13831 11088
rect 13945 11088 13991 11100
rect 13945 11064 13951 11088
rect 13785 11016 13831 11028
rect 13906 11048 13951 11064
rect 13985 11064 13991 11088
rect 13985 11048 14013 11064
rect 13906 10996 13942 11048
rect 13994 10996 14013 11048
rect 13906 10980 14013 10996
rect 14466 11051 14798 11057
rect 14466 10999 14484 11051
rect 14536 10999 14564 11051
rect 14616 10999 14644 11051
rect 14696 10999 14724 11051
rect 14776 10999 14798 11051
rect 14466 10989 14798 10999
rect 15198 11051 15530 11057
rect 15198 10999 15216 11051
rect 15268 10999 15296 11051
rect 15348 10999 15376 11051
rect 15428 10999 15456 11051
rect 15508 10999 15530 11051
rect 15198 10989 15530 10999
rect 15701 10941 15759 12088
rect 15800 11051 16132 11057
rect 15800 10999 15822 11051
rect 15874 10999 15902 11051
rect 15954 10999 15982 11051
rect 16034 10999 16062 11051
rect 16114 10999 16132 11051
rect 15800 10989 16132 10999
rect 16410 11051 16742 11057
rect 16410 10999 16428 11051
rect 16480 10999 16508 11051
rect 16560 10999 16588 11051
rect 16640 10999 16668 11051
rect 16720 10999 16742 11051
rect 16410 10989 16742 10999
rect 17012 11051 17344 11057
rect 17012 10999 17034 11051
rect 17086 10999 17114 11051
rect 17166 10999 17194 11051
rect 17246 10999 17274 11051
rect 17326 10999 17344 11051
rect 17012 10989 17344 10999
rect 17748 11051 18080 11057
rect 17748 10999 17766 11051
rect 17818 10999 17846 11051
rect 17898 10999 17926 11051
rect 17978 10999 18006 11051
rect 18058 10999 18080 11051
rect 17748 10989 18080 10999
rect 13479 10913 15759 10941
rect 18127 10885 18185 12088
rect 18350 11051 18682 11057
rect 18350 10999 18372 11051
rect 18424 10999 18452 11051
rect 18504 10999 18532 11051
rect 18584 10999 18612 11051
rect 18664 10999 18682 11051
rect 18350 10989 18682 10999
rect 13481 10857 18185 10885
rect 18983 10956 19042 12088
rect 19595 12101 19641 12113
rect 19595 12041 19601 12101
rect 19635 12041 19641 12101
rect 19595 11989 19641 12041
rect 19683 12110 19921 12139
rect 20568 12138 20626 12144
rect 20327 12132 20392 12133
rect 20327 12131 20333 12132
rect 20231 12129 20333 12131
rect 19683 12101 19729 12110
rect 19683 12041 19689 12101
rect 19723 12041 19729 12101
rect 20229 12083 20333 12129
rect 20327 12080 20333 12083
rect 20385 12080 20392 12132
rect 20568 12104 20580 12138
rect 20614 12104 20626 12138
rect 20568 12098 20626 12104
rect 20664 12329 20710 12819
rect 26378 12699 26468 12715
rect 26378 12688 26397 12699
rect 26303 12647 26397 12688
rect 26449 12647 26468 12699
rect 20760 12632 20809 12639
rect 20760 12627 21379 12632
rect 20760 12593 20769 12627
rect 20803 12593 21379 12627
rect 20760 12585 21379 12593
rect 20760 12580 20809 12585
rect 20761 12538 20810 12546
rect 21330 12538 21379 12585
rect 26303 12629 26468 12647
rect 26303 12583 26350 12629
rect 26304 12580 26350 12583
rect 20761 12534 21262 12538
rect 20761 12500 20770 12534
rect 20804 12529 21262 12534
rect 20804 12500 21211 12529
rect 20761 12495 21211 12500
rect 21245 12495 21262 12529
rect 20761 12492 21262 12495
rect 21330 12532 25751 12538
rect 21330 12498 21943 12532
rect 21977 12498 22069 12532
rect 22103 12498 23155 12532
rect 23189 12498 23281 12532
rect 23315 12498 24367 12532
rect 24401 12498 24493 12532
rect 24527 12498 25579 12532
rect 25613 12498 25705 12532
rect 25739 12498 25751 12532
rect 26304 12520 26310 12580
rect 26344 12520 26350 12580
rect 26304 12508 26350 12520
rect 26392 12580 26438 12592
rect 26392 12520 26398 12580
rect 26432 12520 26438 12580
rect 26392 12511 26438 12520
rect 21330 12492 25751 12498
rect 20761 12491 21257 12492
rect 21330 12491 21776 12492
rect 20761 12487 20810 12491
rect 21199 12489 21257 12491
rect 26392 12482 26630 12511
rect 21161 12440 21207 12448
rect 21138 12439 21217 12440
rect 21138 12375 21145 12439
rect 21209 12375 21217 12439
rect 21249 12439 21295 12451
rect 21893 12443 21939 12451
rect 21249 12379 21255 12439
rect 21289 12379 21295 12439
rect 21161 12364 21207 12375
rect 21249 12329 21295 12379
rect 21870 12442 21949 12443
rect 21870 12378 21877 12442
rect 21941 12378 21949 12442
rect 21998 12439 22044 12451
rect 22107 12443 22153 12451
rect 23105 12443 23151 12451
rect 21998 12379 22004 12439
rect 22038 12379 22044 12439
rect 21893 12367 21939 12378
rect 21998 12329 22044 12379
rect 22097 12442 22176 12443
rect 22097 12378 22105 12442
rect 22169 12378 22176 12442
rect 23082 12442 23161 12443
rect 23082 12378 23089 12442
rect 23153 12378 23161 12442
rect 23209 12439 23255 12451
rect 23319 12443 23365 12451
rect 24317 12443 24363 12451
rect 23209 12379 23215 12439
rect 23249 12379 23255 12439
rect 22107 12367 22153 12378
rect 23105 12367 23151 12378
rect 23209 12329 23255 12379
rect 23309 12442 23388 12443
rect 23309 12378 23317 12442
rect 23381 12378 23388 12442
rect 24294 12442 24373 12443
rect 24294 12378 24301 12442
rect 24365 12378 24373 12442
rect 24422 12439 24468 12451
rect 24531 12443 24577 12451
rect 25529 12443 25575 12451
rect 24422 12379 24428 12439
rect 24462 12379 24468 12439
rect 23319 12367 23365 12378
rect 24317 12367 24363 12378
rect 24422 12329 24468 12379
rect 24521 12442 24600 12443
rect 24521 12378 24529 12442
rect 24593 12378 24600 12442
rect 25506 12442 25585 12443
rect 25506 12378 25513 12442
rect 25577 12378 25585 12442
rect 25636 12439 25682 12451
rect 25743 12443 25789 12451
rect 25636 12379 25642 12439
rect 25676 12379 25682 12439
rect 24531 12367 24577 12378
rect 25529 12367 25575 12378
rect 25636 12329 25682 12379
rect 25733 12442 25812 12443
rect 25733 12378 25741 12442
rect 25805 12378 25812 12442
rect 26304 12442 26350 12454
rect 26304 12382 26310 12442
rect 26344 12382 26350 12442
rect 25743 12367 25789 12378
rect 26304 12370 26350 12382
rect 26392 12442 26438 12482
rect 26392 12382 26398 12442
rect 26432 12382 26438 12442
rect 26392 12370 26438 12382
rect 26466 12442 26556 12454
rect 26466 12438 26494 12442
rect 26528 12438 26556 12442
rect 26466 12386 26485 12438
rect 26537 12386 26556 12438
rect 26466 12382 26494 12386
rect 26528 12382 26556 12386
rect 26466 12370 26556 12382
rect 26584 12442 26630 12482
rect 26584 12382 26590 12442
rect 26624 12382 26630 12442
rect 26584 12370 26630 12382
rect 26223 12329 26289 12331
rect 20664 12325 26289 12329
rect 20664 12291 26239 12325
rect 26273 12291 26289 12325
rect 20664 12287 26289 12291
rect 20664 12066 20710 12287
rect 21514 12240 21560 12250
rect 21492 12176 21501 12240
rect 21565 12176 21574 12240
rect 21492 12175 21574 12176
rect 21604 12238 21650 12287
rect 22246 12240 22292 12250
rect 21604 12178 21610 12238
rect 21644 12178 21650 12238
rect 21514 12166 21560 12175
rect 21604 12166 21650 12178
rect 22224 12176 22233 12240
rect 22297 12176 22306 12240
rect 22224 12175 22306 12176
rect 22353 12238 22399 12287
rect 22456 12240 22502 12250
rect 23458 12240 23504 12250
rect 22353 12178 22359 12238
rect 22393 12178 22399 12238
rect 22246 12166 22292 12175
rect 22353 12166 22399 12178
rect 22442 12176 22451 12240
rect 22515 12176 22524 12240
rect 22442 12175 22524 12176
rect 23436 12176 23445 12240
rect 23509 12176 23518 12240
rect 23436 12175 23518 12176
rect 23564 12238 23610 12287
rect 23668 12240 23714 12250
rect 24796 12240 24842 12250
rect 23564 12178 23570 12238
rect 23604 12178 23610 12238
rect 22456 12166 22502 12175
rect 23458 12166 23504 12175
rect 23564 12166 23610 12178
rect 23654 12176 23663 12240
rect 23727 12176 23736 12240
rect 23654 12175 23736 12176
rect 24774 12176 24783 12240
rect 24847 12176 24856 12240
rect 24774 12175 24856 12176
rect 24904 12238 24950 12287
rect 25006 12240 25052 12250
rect 24904 12178 24910 12238
rect 24944 12178 24950 12238
rect 23668 12166 23714 12175
rect 24796 12166 24842 12175
rect 24904 12166 24950 12178
rect 24992 12176 25001 12240
rect 25065 12176 25074 12240
rect 24992 12175 25074 12176
rect 25651 12238 25697 12287
rect 26227 12285 26289 12287
rect 26322 12322 26350 12370
rect 26434 12323 26704 12329
rect 26434 12322 26446 12323
rect 26322 12293 26446 12322
rect 26322 12251 26350 12293
rect 26434 12289 26446 12293
rect 26480 12289 26704 12323
rect 26434 12283 26704 12289
rect 25740 12240 25786 12250
rect 25651 12178 25657 12238
rect 25691 12178 25697 12238
rect 25006 12166 25052 12175
rect 25651 12166 25697 12178
rect 25726 12176 25735 12240
rect 25799 12176 25808 12240
rect 25726 12175 25808 12176
rect 26304 12239 26350 12251
rect 26304 12179 26310 12239
rect 26344 12179 26350 12239
rect 25740 12166 25786 12175
rect 26304 12167 26350 12179
rect 26392 12239 26438 12251
rect 26392 12179 26398 12239
rect 26432 12179 26438 12239
rect 26392 12139 26438 12179
rect 26466 12239 26556 12251
rect 26466 12235 26494 12239
rect 26528 12235 26556 12239
rect 26466 12183 26485 12235
rect 26537 12183 26556 12235
rect 26466 12179 26494 12183
rect 26528 12179 26556 12183
rect 26466 12167 26556 12179
rect 26584 12239 26630 12251
rect 26584 12179 26590 12239
rect 26624 12179 26630 12239
rect 26584 12139 26630 12179
rect 25692 12134 25751 12137
rect 20814 12080 20821 12132
rect 20873 12130 20879 12132
rect 21552 12130 21610 12134
rect 20873 12128 21610 12130
rect 20873 12094 21564 12128
rect 21598 12113 21610 12128
rect 22284 12128 23680 12134
rect 21598 12094 21612 12113
rect 20873 12083 21612 12094
rect 22284 12094 22296 12128
rect 22330 12094 22418 12128
rect 22452 12094 23508 12128
rect 23542 12094 23630 12128
rect 23664 12094 23680 12128
rect 22284 12088 23680 12094
rect 24834 12128 25018 12134
rect 24834 12094 24846 12128
rect 24880 12094 24968 12128
rect 25002 12094 25018 12128
rect 24834 12088 25018 12094
rect 25690 12128 25751 12134
rect 25690 12094 25702 12128
rect 25736 12094 25751 12128
rect 25690 12088 25751 12094
rect 20873 12080 20879 12083
rect 20814 12079 20879 12080
rect 21554 12078 21612 12083
rect 19683 12029 19729 12041
rect 20494 12054 20540 12066
rect 20494 11994 20500 12054
rect 20534 11994 20540 12054
rect 19595 11973 19756 11989
rect 19595 11921 19685 11973
rect 19737 11921 19756 11973
rect 19595 11905 19756 11921
rect 20494 11916 20540 11994
rect 20654 12054 20710 12066
rect 20654 11994 20660 12054
rect 20694 11994 20710 12054
rect 20654 11982 20710 11994
rect 20494 11856 20500 11916
rect 20534 11856 20540 11916
rect 20494 11844 20540 11856
rect 20654 11916 20700 11928
rect 20654 11856 20660 11916
rect 20694 11856 20700 11916
rect 20494 11778 20540 11790
rect 20494 11718 20500 11778
rect 20534 11718 20540 11778
rect 20494 11640 20540 11718
rect 20654 11778 20700 11856
rect 20654 11718 20660 11778
rect 20694 11718 20700 11778
rect 20654 11706 20700 11718
rect 20494 11580 20500 11640
rect 20534 11580 20540 11640
rect 20494 11568 20540 11580
rect 20654 11640 20700 11652
rect 20654 11580 20660 11640
rect 20694 11580 20700 11640
rect 20494 11502 20540 11514
rect 20494 11442 20500 11502
rect 20534 11442 20540 11502
rect 20494 11364 20540 11442
rect 20654 11502 20700 11580
rect 20654 11442 20660 11502
rect 20694 11442 20700 11502
rect 20654 11430 20700 11442
rect 20494 11304 20500 11364
rect 20534 11304 20540 11364
rect 20494 11292 20540 11304
rect 20654 11364 20700 11376
rect 20654 11304 20660 11364
rect 20694 11304 20700 11364
rect 20494 11226 20540 11238
rect 20494 11166 20500 11226
rect 20534 11166 20540 11226
rect 20494 11088 20540 11166
rect 20654 11226 20700 11304
rect 20654 11166 20660 11226
rect 20694 11166 20700 11226
rect 20654 11154 20700 11166
rect 19084 11051 19416 11057
rect 19084 10999 19106 11051
rect 19158 10999 19186 11051
rect 19238 10999 19266 11051
rect 19318 10999 19346 11051
rect 19398 10999 19416 11051
rect 20494 11028 20500 11088
rect 20534 11028 20540 11088
rect 20654 11088 20700 11100
rect 20654 11064 20660 11088
rect 20494 11016 20540 11028
rect 20615 11048 20660 11064
rect 20694 11064 20700 11088
rect 20694 11048 20722 11064
rect 19084 10989 19416 10999
rect 20615 10996 20651 11048
rect 20703 10996 20722 11048
rect 20615 10980 20722 10996
rect 21175 11051 21507 11057
rect 21175 10999 21193 11051
rect 21245 10999 21273 11051
rect 21325 10999 21353 11051
rect 21405 10999 21433 11051
rect 21485 10999 21507 11051
rect 21175 10989 21507 10999
rect 21907 11051 22239 11057
rect 21907 10999 21925 11051
rect 21977 10999 22005 11051
rect 22057 10999 22085 11051
rect 22137 10999 22165 11051
rect 22217 10999 22239 11051
rect 21907 10989 22239 10999
rect 18983 10829 19041 10956
rect 13483 10801 19041 10829
rect 22410 10773 22468 12088
rect 22509 11051 22841 11057
rect 22509 10999 22531 11051
rect 22583 10999 22611 11051
rect 22663 10999 22691 11051
rect 22743 10999 22771 11051
rect 22823 10999 22841 11051
rect 22509 10989 22841 10999
rect 23119 11051 23451 11057
rect 23119 10999 23137 11051
rect 23189 10999 23217 11051
rect 23269 10999 23297 11051
rect 23349 10999 23377 11051
rect 23429 10999 23451 11051
rect 23119 10989 23451 10999
rect 23721 11051 24053 11057
rect 23721 10999 23743 11051
rect 23795 10999 23823 11051
rect 23875 10999 23903 11051
rect 23955 10999 23983 11051
rect 24035 10999 24053 11051
rect 23721 10989 24053 10999
rect 24457 11051 24789 11057
rect 24457 10999 24475 11051
rect 24527 10999 24555 11051
rect 24607 10999 24635 11051
rect 24687 10999 24715 11051
rect 24767 10999 24789 11051
rect 24457 10989 24789 10999
rect 13484 10745 22468 10773
rect 24836 10717 24894 12088
rect 25059 11051 25391 11057
rect 25059 10999 25081 11051
rect 25133 10999 25161 11051
rect 25213 10999 25241 11051
rect 25293 10999 25321 11051
rect 25373 10999 25391 11051
rect 25059 10989 25391 10999
rect 13486 10689 24894 10717
rect 25692 10956 25751 12088
rect 26304 12101 26350 12113
rect 26304 12041 26310 12101
rect 26344 12041 26350 12101
rect 26304 11989 26350 12041
rect 26392 12110 26630 12139
rect 26392 12101 26438 12110
rect 26392 12041 26398 12101
rect 26432 12041 26438 12101
rect 26392 12029 26438 12041
rect 26304 11973 26465 11989
rect 26304 11921 26394 11973
rect 26446 11921 26465 11973
rect 26304 11905 26465 11921
rect 25793 11051 26125 11057
rect 25793 10999 25815 11051
rect 25867 10999 25895 11051
rect 25947 10999 25975 11051
rect 26027 10999 26055 11051
rect 26107 10999 26125 11051
rect 25793 10989 26125 10999
rect 25692 10661 25750 10956
rect 13485 10633 25750 10661
rect 8196 10576 8528 10582
rect 8196 10524 8218 10576
rect 8270 10524 8298 10576
rect 8350 10524 8378 10576
rect 8430 10524 8458 10576
rect 8510 10524 8528 10576
rect 8196 10514 8528 10524
rect 13473 10579 25786 10605
rect 13473 10578 25716 10579
rect 13473 10526 14112 10578
rect 14164 10571 25716 10578
rect 14164 10568 20821 10571
rect 14164 10526 19012 10568
rect 13473 10516 19012 10526
rect 19065 10518 20821 10568
rect 20873 10518 25716 10571
rect 19065 10516 25716 10518
rect 13473 10515 25716 10516
rect 25780 10515 25786 10579
rect 13473 10493 25786 10515
rect 13481 10437 24187 10465
rect 13484 10381 21761 10409
rect 2929 10337 8154 10365
rect 13486 10325 20905 10353
rect 2928 10281 8154 10309
rect 2932 10225 7297 10253
rect 2930 10169 4871 10197
rect 3018 10125 3125 10141
rect 2897 10093 2943 10105
rect 2897 10033 2903 10093
rect 2937 10033 2943 10093
rect 3018 10073 3054 10125
rect 3106 10073 3125 10125
rect 3018 10057 3063 10073
rect 2897 9955 2943 10033
rect 3057 10033 3063 10057
rect 3097 10057 3125 10073
rect 3578 10122 3910 10132
rect 3578 10070 3596 10122
rect 3648 10070 3676 10122
rect 3728 10070 3756 10122
rect 3808 10070 3836 10122
rect 3888 10070 3910 10122
rect 3578 10064 3910 10070
rect 4310 10122 4642 10132
rect 4310 10070 4328 10122
rect 4380 10070 4408 10122
rect 4460 10070 4488 10122
rect 4540 10070 4568 10122
rect 4620 10070 4642 10122
rect 4310 10064 4642 10070
rect 3097 10033 3103 10057
rect 3057 10021 3103 10033
rect 2897 9895 2903 9955
rect 2937 9895 2943 9955
rect 2897 9883 2943 9895
rect 3057 9955 3103 9967
rect 3057 9895 3063 9955
rect 3097 9895 3103 9955
rect 2897 9817 2943 9829
rect 2897 9757 2903 9817
rect 2937 9757 2943 9817
rect 2897 9679 2943 9757
rect 3057 9817 3103 9895
rect 3057 9757 3063 9817
rect 3097 9757 3103 9817
rect 3057 9745 3103 9757
rect 2897 9619 2903 9679
rect 2937 9619 2943 9679
rect 2897 9607 2943 9619
rect 3057 9679 3103 9691
rect 3057 9619 3063 9679
rect 3097 9619 3103 9679
rect 2897 9541 2943 9553
rect 2897 9481 2903 9541
rect 2937 9481 2943 9541
rect 2897 9403 2943 9481
rect 3057 9541 3103 9619
rect 3057 9481 3063 9541
rect 3097 9481 3103 9541
rect 3057 9469 3103 9481
rect 2897 9343 2903 9403
rect 2937 9343 2943 9403
rect 2897 9331 2943 9343
rect 3057 9403 3103 9415
rect 3057 9343 3063 9403
rect 3097 9343 3103 9403
rect 2897 9265 2943 9277
rect 2897 9205 2903 9265
rect 2937 9205 2943 9265
rect 2897 9127 2943 9205
rect 3057 9265 3103 9343
rect 3057 9205 3063 9265
rect 3097 9205 3103 9265
rect 3057 9193 3103 9205
rect 2897 9067 2903 9127
rect 2937 9067 2943 9127
rect 2897 9055 2943 9067
rect 3057 9127 3113 9139
rect 3057 9067 3063 9127
rect 3097 9067 3113 9127
rect 3057 9055 3113 9067
rect 2730 9038 2736 9041
rect 2632 8992 2736 9038
rect 2634 8990 2736 8992
rect 2730 8989 2736 8990
rect 2788 8989 2795 9041
rect 2730 8988 2795 8989
rect 2971 9017 3029 9023
rect 2971 8983 2983 9017
rect 3017 8983 3029 9017
rect 2971 8977 3029 8983
rect 2981 8836 3029 8977
rect 2361 8789 3029 8836
rect 2386 8698 2846 8720
rect 2386 8689 2469 8698
rect 2521 8689 2589 8698
rect 2641 8689 2732 8698
rect 2784 8689 2846 8698
rect 2386 8655 2415 8689
rect 2449 8655 2469 8689
rect 2541 8655 2589 8689
rect 2641 8655 2691 8689
rect 2725 8655 2732 8689
rect 2817 8655 2846 8689
rect 2386 8646 2469 8655
rect 2521 8646 2589 8655
rect 2641 8646 2732 8655
rect 2784 8646 2846 8655
rect 2386 8624 2846 8646
rect 2904 8546 2953 8559
rect 2904 8522 2913 8546
rect 2810 8512 2913 8522
rect 2947 8512 2953 8546
rect 2810 8494 2953 8512
rect 2716 8463 2782 8464
rect 2453 8456 2507 8460
rect 2453 8453 2508 8456
rect 2324 8419 2462 8453
rect 2496 8419 2508 8453
rect 2453 8416 2508 8419
rect 2454 8412 2508 8416
rect 2716 8411 2724 8463
rect 2776 8411 2782 8463
rect 2716 8409 2782 8411
rect 2810 8350 2838 8494
rect 2636 8343 2838 8350
rect 2636 8309 2652 8343
rect 2686 8322 2838 8343
rect 2866 8453 2915 8466
rect 2866 8419 2875 8453
rect 2909 8419 2915 8453
rect 2866 8407 2915 8419
rect 2686 8309 2703 8322
rect 2636 8303 2703 8309
rect 2531 8288 2589 8295
rect 2531 8254 2543 8288
rect 2577 8275 2589 8288
rect 2866 8275 2894 8407
rect 2981 8399 3029 8789
rect 3067 8834 3113 9055
rect 3217 9041 3282 9042
rect 3217 8989 3224 9041
rect 3276 9038 3282 9041
rect 3957 9038 4015 9043
rect 3276 9027 4015 9038
rect 4813 9033 4871 10169
rect 4912 10122 5244 10132
rect 4912 10070 4934 10122
rect 4986 10070 5014 10122
rect 5066 10070 5094 10122
rect 5146 10070 5174 10122
rect 5226 10070 5244 10122
rect 4912 10064 5244 10070
rect 5522 10122 5854 10132
rect 5522 10070 5540 10122
rect 5592 10070 5620 10122
rect 5672 10070 5700 10122
rect 5752 10070 5780 10122
rect 5832 10070 5854 10122
rect 5522 10064 5854 10070
rect 6124 10122 6456 10132
rect 6124 10070 6146 10122
rect 6198 10070 6226 10122
rect 6278 10070 6306 10122
rect 6358 10070 6386 10122
rect 6438 10070 6456 10122
rect 6124 10064 6456 10070
rect 6860 10122 7192 10132
rect 6860 10070 6878 10122
rect 6930 10070 6958 10122
rect 7010 10070 7038 10122
rect 7090 10070 7118 10122
rect 7170 10070 7192 10122
rect 6860 10064 7192 10070
rect 7239 9033 7297 10225
rect 7462 10122 7794 10132
rect 7462 10070 7484 10122
rect 7536 10070 7564 10122
rect 7616 10070 7644 10122
rect 7696 10070 7724 10122
rect 7776 10070 7794 10122
rect 7462 10064 7794 10070
rect 8095 9033 8154 10281
rect 13481 10269 17478 10297
rect 13484 10213 15052 10241
rect 13484 10157 14196 10185
rect 8196 10122 8528 10132
rect 8196 10070 8218 10122
rect 8270 10070 8298 10122
rect 8350 10070 8378 10122
rect 8430 10070 8458 10122
rect 8510 10070 8528 10122
rect 8196 10064 8528 10070
rect 13763 10110 14095 10120
rect 13763 10058 13781 10110
rect 13833 10058 13861 10110
rect 13913 10058 13941 10110
rect 13993 10058 14021 10110
rect 14073 10058 14095 10110
rect 13763 10052 14095 10058
rect 12671 9976 12677 10028
rect 12729 10024 12735 10028
rect 13199 10024 13205 10030
rect 12729 9984 13205 10024
rect 12729 9976 12735 9984
rect 13199 9978 13205 9984
rect 13257 9978 13263 10030
rect 3276 8993 3967 9027
rect 4001 9008 4015 9027
rect 4687 9027 6083 9033
rect 4001 8993 4013 9008
rect 3276 8991 4013 8993
rect 3276 8989 3282 8991
rect 3955 8987 4013 8991
rect 4687 8993 4699 9027
rect 4733 8993 4821 9027
rect 4855 8993 5911 9027
rect 5945 8993 6033 9027
rect 6067 8993 6083 9027
rect 4687 8987 6083 8993
rect 7237 9027 7421 9033
rect 7237 8993 7249 9027
rect 7283 8993 7371 9027
rect 7405 8993 7421 9027
rect 7237 8987 7421 8993
rect 8093 9027 8154 9033
rect 8093 8993 8105 9027
rect 8139 8993 8154 9027
rect 8707 9200 8868 9216
rect 8707 9148 8797 9200
rect 8849 9148 8868 9200
rect 13423 9188 13584 9204
rect 8707 9132 8868 9148
rect 9189 9159 9296 9175
rect 8707 9080 8753 9132
rect 9189 9107 9225 9159
rect 9277 9107 9296 9159
rect 9189 9099 9296 9107
rect 9666 9159 9773 9175
rect 9666 9107 9702 9159
rect 9754 9107 9773 9159
rect 9666 9099 9773 9107
rect 10086 9148 10193 9164
rect 9806 9099 9840 9102
rect 9898 9099 9932 9103
rect 9990 9099 10024 9102
rect 10086 9101 10122 9148
rect 10082 9099 10122 9101
rect 9061 9096 10122 9099
rect 10174 9102 10193 9148
rect 10462 9156 10569 9172
rect 10462 9104 10498 9156
rect 10550 9104 10569 9156
rect 10462 9102 10569 9104
rect 10810 9156 10917 9172
rect 10810 9104 10846 9156
rect 10898 9104 10917 9156
rect 10174 9099 10208 9102
rect 10266 9099 10300 9102
rect 10358 9099 10392 9102
rect 10450 9099 10576 9102
rect 10634 9099 10668 9102
rect 10726 9099 10760 9102
rect 10810 9101 10917 9104
rect 11068 9162 11175 9178
rect 11068 9110 11104 9162
rect 11156 9110 11175 9162
rect 10810 9099 10944 9101
rect 11002 9099 11036 9102
rect 11068 9099 11175 9110
rect 11294 9162 11401 9178
rect 11294 9110 11330 9162
rect 11382 9110 11401 9162
rect 11294 9102 11401 9110
rect 11553 9165 11660 9181
rect 11553 9113 11589 9165
rect 11641 9113 11660 9165
rect 11278 9099 11404 9102
rect 11462 9099 11496 9102
rect 11553 9101 11660 9113
rect 12160 9127 12267 9143
rect 11553 9099 11680 9101
rect 10174 9096 11709 9099
rect 8707 9020 8713 9080
rect 8747 9020 8753 9080
rect 8707 9008 8753 9020
rect 8795 9080 8841 9092
rect 8795 9020 8801 9080
rect 8835 9020 8841 9080
rect 8795 9011 8841 9020
rect 9061 9068 11709 9096
rect 12160 9088 12196 9127
rect 12117 9085 12196 9088
rect 9061 9034 9090 9068
rect 9124 9034 9182 9068
rect 9216 9034 9274 9068
rect 9308 9034 9346 9068
rect 9380 9034 9438 9068
rect 9472 9034 9530 9068
rect 9564 9034 9622 9068
rect 9656 9034 9714 9068
rect 9748 9034 9806 9068
rect 9840 9034 9898 9068
rect 9932 9034 9990 9068
rect 10024 9034 10082 9068
rect 10116 9034 10174 9068
rect 10208 9034 10266 9068
rect 10300 9034 10358 9068
rect 10392 9034 10450 9068
rect 10484 9034 10542 9068
rect 10576 9034 10634 9068
rect 10668 9034 10726 9068
rect 10760 9034 10818 9068
rect 10852 9034 10910 9068
rect 10944 9034 11002 9068
rect 11036 9034 11094 9068
rect 11128 9034 11186 9068
rect 11220 9034 11278 9068
rect 11312 9034 11370 9068
rect 11404 9034 11462 9068
rect 11496 9034 11554 9068
rect 11588 9034 11646 9068
rect 11680 9034 11709 9068
rect 8093 8987 8154 8993
rect 8095 8984 8154 8987
rect 8795 8982 9033 9011
rect 9061 9003 11709 9034
rect 12114 9075 12196 9085
rect 12248 9088 12267 9127
rect 12392 9128 12499 9144
rect 12392 9088 12428 9128
rect 12248 9076 12428 9088
rect 12480 9088 12499 9128
rect 12828 9134 12935 9150
rect 12480 9086 12557 9088
rect 12828 9086 12864 9134
rect 12480 9082 12864 9086
rect 12916 9086 12935 9134
rect 13063 9136 13170 9152
rect 13063 9086 13099 9136
rect 12916 9084 13099 9086
rect 13151 9086 13170 9136
rect 13423 9136 13442 9188
rect 13494 9136 13584 9188
rect 13423 9120 13584 9136
rect 13151 9084 13201 9086
rect 12916 9082 13201 9084
rect 12480 9076 13201 9082
rect 12248 9075 13201 9076
rect 12114 9055 13201 9075
rect 12114 9052 12678 9055
rect 12114 9018 12150 9052
rect 12184 9018 12222 9052
rect 12256 9018 12295 9052
rect 12329 9018 12367 9052
rect 12401 9051 12678 9052
rect 12401 9018 12440 9051
rect 3917 8946 3963 8955
rect 3895 8945 3977 8946
rect 3895 8881 3904 8945
rect 3968 8881 3977 8945
rect 4007 8943 4053 8955
rect 4649 8946 4695 8955
rect 4007 8883 4013 8943
rect 4047 8883 4053 8943
rect 3917 8871 3963 8881
rect 4007 8834 4053 8883
rect 4627 8945 4709 8946
rect 4627 8881 4636 8945
rect 4700 8881 4709 8945
rect 4756 8943 4802 8955
rect 4859 8946 4905 8955
rect 5861 8946 5907 8955
rect 4756 8883 4762 8943
rect 4796 8883 4802 8943
rect 4649 8871 4695 8881
rect 4756 8834 4802 8883
rect 4845 8945 4927 8946
rect 4845 8881 4854 8945
rect 4918 8881 4927 8945
rect 5839 8945 5921 8946
rect 5839 8881 5848 8945
rect 5912 8881 5921 8945
rect 5967 8943 6013 8955
rect 6071 8946 6117 8955
rect 7199 8946 7245 8955
rect 5967 8883 5973 8943
rect 6007 8883 6013 8943
rect 4859 8871 4905 8881
rect 5861 8871 5907 8881
rect 5967 8834 6013 8883
rect 6057 8945 6139 8946
rect 6057 8881 6066 8945
rect 6130 8881 6139 8945
rect 7177 8945 7259 8946
rect 7177 8881 7186 8945
rect 7250 8881 7259 8945
rect 7307 8943 7353 8955
rect 7409 8946 7455 8955
rect 7307 8883 7313 8943
rect 7347 8883 7353 8943
rect 6071 8871 6117 8881
rect 7199 8871 7245 8881
rect 7307 8834 7353 8883
rect 7395 8945 7477 8946
rect 7395 8881 7404 8945
rect 7468 8881 7477 8945
rect 8054 8943 8100 8955
rect 8143 8946 8189 8955
rect 8054 8883 8060 8943
rect 8094 8883 8100 8943
rect 7409 8871 7455 8881
rect 8054 8834 8100 8883
rect 8129 8945 8211 8946
rect 8129 8881 8138 8945
rect 8202 8881 8211 8945
rect 8707 8942 8753 8954
rect 8707 8882 8713 8942
rect 8747 8882 8753 8942
rect 8143 8871 8189 8881
rect 8707 8870 8753 8882
rect 8795 8942 8841 8982
rect 8795 8882 8801 8942
rect 8835 8882 8841 8942
rect 8795 8870 8841 8882
rect 8869 8942 8959 8954
rect 8869 8938 8897 8942
rect 8931 8938 8959 8942
rect 8869 8886 8888 8938
rect 8940 8886 8959 8938
rect 8869 8882 8897 8886
rect 8931 8882 8959 8886
rect 8869 8870 8959 8882
rect 8987 8942 9033 8982
rect 8987 8882 8993 8942
rect 9027 8882 9033 8942
rect 11827 8984 12065 9018
rect 12114 9017 12440 9018
rect 12474 9017 12512 9051
rect 12546 9021 12678 9051
rect 12712 9021 12770 9055
rect 12804 9021 12862 9055
rect 12896 9021 12954 9055
rect 12988 9021 13046 9055
rect 13080 9021 13138 9055
rect 13172 9021 13201 9055
rect 12546 9017 13201 9021
rect 12114 8990 13201 9017
rect 13450 9068 13496 9080
rect 13450 9008 13456 9068
rect 13490 9008 13496 9068
rect 13450 8999 13496 9008
rect 12114 8989 12191 8990
rect 11827 8944 11873 8984
rect 10302 8913 10357 8923
rect 8987 8870 9033 8882
rect 10161 8898 10219 8904
rect 8630 8834 8692 8836
rect 3067 8830 8692 8834
rect 3067 8796 8642 8830
rect 8676 8796 8692 8830
rect 3067 8792 8692 8796
rect 2981 8392 3036 8399
rect 2981 8389 2984 8392
rect 2960 8383 2984 8389
rect 2960 8349 2972 8383
rect 2960 8343 2984 8349
rect 2984 8334 3036 8340
rect 3067 8302 3113 8792
rect 3564 8746 3610 8757
rect 3541 8682 3548 8746
rect 3612 8682 3620 8746
rect 3541 8681 3620 8682
rect 3652 8742 3698 8792
rect 4296 8743 4342 8754
rect 3652 8682 3658 8742
rect 3692 8682 3698 8742
rect 3564 8673 3610 8681
rect 3652 8670 3698 8682
rect 4273 8679 4280 8743
rect 4344 8679 4352 8743
rect 4273 8678 4352 8679
rect 4401 8742 4447 8792
rect 4510 8743 4556 8754
rect 5508 8743 5554 8754
rect 4401 8682 4407 8742
rect 4441 8682 4447 8742
rect 4296 8670 4342 8678
rect 4401 8670 4447 8682
rect 4500 8679 4508 8743
rect 4572 8679 4579 8743
rect 4500 8678 4579 8679
rect 5485 8679 5492 8743
rect 5556 8679 5564 8743
rect 5485 8678 5564 8679
rect 5612 8742 5658 8792
rect 5722 8743 5768 8754
rect 6720 8743 6766 8754
rect 5612 8682 5618 8742
rect 5652 8682 5658 8742
rect 4510 8670 4556 8678
rect 5508 8670 5554 8678
rect 5612 8670 5658 8682
rect 5712 8679 5720 8743
rect 5784 8679 5791 8743
rect 5712 8678 5791 8679
rect 6697 8679 6704 8743
rect 6768 8679 6776 8743
rect 6697 8678 6776 8679
rect 6825 8742 6871 8792
rect 6934 8743 6980 8754
rect 7932 8743 7978 8754
rect 6825 8682 6831 8742
rect 6865 8682 6871 8742
rect 5722 8670 5768 8678
rect 6720 8670 6766 8678
rect 6825 8670 6871 8682
rect 6924 8679 6932 8743
rect 6996 8679 7003 8743
rect 6924 8678 7003 8679
rect 7909 8679 7916 8743
rect 7980 8679 7988 8743
rect 7909 8678 7988 8679
rect 8039 8742 8085 8792
rect 8626 8790 8692 8792
rect 8725 8828 8753 8870
rect 10161 8864 10173 8898
rect 10207 8895 10219 8898
rect 10302 8895 10303 8913
rect 10207 8867 10303 8895
rect 10207 8864 10219 8867
rect 10161 8858 10219 8864
rect 10302 8859 10303 8867
rect 10897 8898 10955 8904
rect 10897 8895 10909 8898
rect 10357 8867 10909 8895
rect 10302 8852 10357 8859
rect 10897 8864 10909 8867
rect 10943 8864 10955 8898
rect 10897 8858 10955 8864
rect 11085 8898 11143 8904
rect 11085 8864 11097 8898
rect 11131 8895 11143 8898
rect 11449 8898 11507 8904
rect 11449 8895 11461 8898
rect 11131 8867 11461 8895
rect 11131 8864 11143 8867
rect 11085 8858 11143 8864
rect 11449 8864 11461 8867
rect 11495 8864 11507 8898
rect 11827 8888 11833 8944
rect 11449 8858 11507 8864
rect 11826 8884 11833 8888
rect 11867 8888 11873 8944
rect 11923 8944 11969 8956
rect 11867 8884 11874 8888
rect 9004 8838 9183 8839
rect 8837 8833 9183 8838
rect 8837 8832 9136 8833
rect 8837 8828 8849 8832
rect 8725 8799 8849 8828
rect 8146 8743 8192 8754
rect 8725 8751 8753 8799
rect 8837 8798 8849 8799
rect 8883 8799 9136 8832
rect 9170 8799 9183 8833
rect 8883 8798 9183 8799
rect 8837 8793 9183 8798
rect 9224 8828 9845 8834
rect 9224 8794 9236 8828
rect 9270 8827 9845 8828
rect 9270 8794 9789 8827
rect 9224 8793 9789 8794
rect 9823 8793 9845 8827
rect 8837 8792 9019 8793
rect 9224 8786 9845 8793
rect 10437 8830 10495 8836
rect 10437 8796 10449 8830
rect 10483 8827 10495 8830
rect 11085 8827 11124 8858
rect 10483 8799 11124 8827
rect 10483 8796 10495 8799
rect 10437 8790 10495 8796
rect 9885 8762 9943 8768
rect 8039 8682 8045 8742
rect 8079 8682 8085 8742
rect 6934 8670 6980 8678
rect 7932 8670 7978 8678
rect 8039 8670 8085 8682
rect 8136 8679 8144 8743
rect 8208 8679 8215 8743
rect 8136 8678 8215 8679
rect 8707 8739 8753 8751
rect 8707 8679 8713 8739
rect 8747 8679 8753 8739
rect 8146 8670 8192 8678
rect 8707 8667 8753 8679
rect 8795 8739 8841 8751
rect 8795 8679 8801 8739
rect 8835 8679 8841 8739
rect 8795 8639 8841 8679
rect 8869 8739 8959 8751
rect 8869 8735 8897 8739
rect 8931 8735 8959 8739
rect 8869 8683 8888 8735
rect 8940 8683 8959 8735
rect 8869 8679 8897 8683
rect 8931 8679 8959 8683
rect 8869 8667 8959 8679
rect 8987 8739 9033 8751
rect 8987 8679 8993 8739
rect 9027 8679 9033 8739
rect 9885 8728 9897 8762
rect 9931 8759 9943 8762
rect 10529 8762 10587 8768
rect 10529 8759 10541 8762
rect 9931 8731 10541 8759
rect 9931 8728 9943 8731
rect 9885 8722 9943 8728
rect 10529 8728 10541 8731
rect 10575 8728 10587 8762
rect 11538 8728 11544 8780
rect 11596 8760 11602 8780
rect 11638 8762 11692 8774
rect 11638 8760 11652 8762
rect 11596 8730 11652 8760
rect 11596 8728 11602 8730
rect 11638 8728 11652 8730
rect 11686 8728 11692 8762
rect 10529 8722 10587 8728
rect 11638 8716 11692 8728
rect 11826 8728 11874 8884
rect 11923 8884 11929 8944
rect 11963 8884 11969 8944
rect 11923 8872 11969 8884
rect 12019 8944 12065 8984
rect 13258 8970 13496 8999
rect 13538 9068 13584 9120
rect 13538 9008 13544 9068
rect 13578 9008 13584 9068
rect 13538 8996 13584 9008
rect 14137 9021 14196 10157
rect 14497 10110 14829 10120
rect 14497 10058 14515 10110
rect 14567 10058 14595 10110
rect 14647 10058 14675 10110
rect 14727 10058 14755 10110
rect 14807 10058 14829 10110
rect 14497 10052 14829 10058
rect 14994 9021 15052 10213
rect 15099 10110 15431 10120
rect 15099 10058 15121 10110
rect 15173 10058 15201 10110
rect 15253 10058 15281 10110
rect 15333 10058 15361 10110
rect 15413 10058 15431 10110
rect 15099 10052 15431 10058
rect 15835 10110 16167 10120
rect 15835 10058 15853 10110
rect 15905 10058 15933 10110
rect 15985 10058 16013 10110
rect 16065 10058 16093 10110
rect 16145 10058 16167 10110
rect 15835 10052 16167 10058
rect 16437 10110 16769 10120
rect 16437 10058 16459 10110
rect 16511 10058 16539 10110
rect 16591 10058 16619 10110
rect 16671 10058 16699 10110
rect 16751 10058 16769 10110
rect 16437 10052 16769 10058
rect 17047 10110 17379 10120
rect 17047 10058 17065 10110
rect 17117 10058 17145 10110
rect 17197 10058 17225 10110
rect 17277 10058 17305 10110
rect 17357 10058 17379 10110
rect 17047 10052 17379 10058
rect 17420 9021 17478 10269
rect 20847 10153 20905 10325
rect 17649 10110 17981 10120
rect 17649 10058 17671 10110
rect 17723 10058 17751 10110
rect 17803 10058 17831 10110
rect 17883 10058 17911 10110
rect 17963 10058 17981 10110
rect 17649 10052 17981 10058
rect 18381 10110 18713 10120
rect 18381 10058 18403 10110
rect 18455 10058 18483 10110
rect 18535 10058 18563 10110
rect 18615 10058 18643 10110
rect 18695 10058 18713 10110
rect 18381 10052 18713 10058
rect 19166 10113 19273 10129
rect 19166 10061 19185 10113
rect 19237 10061 19273 10113
rect 20472 10110 20804 10120
rect 19166 10045 19194 10061
rect 19188 10021 19194 10045
rect 19228 10045 19273 10061
rect 19348 10081 19394 10093
rect 19228 10021 19234 10045
rect 19188 10009 19234 10021
rect 19348 10021 19354 10081
rect 19388 10021 19394 10081
rect 20472 10058 20490 10110
rect 20542 10058 20570 10110
rect 20622 10058 20650 10110
rect 20702 10058 20730 10110
rect 20782 10058 20804 10110
rect 20472 10052 20804 10058
rect 19188 9943 19234 9955
rect 19188 9883 19194 9943
rect 19228 9883 19234 9943
rect 19188 9805 19234 9883
rect 19348 9943 19394 10021
rect 19348 9883 19354 9943
rect 19388 9883 19394 9943
rect 19348 9871 19394 9883
rect 19188 9745 19194 9805
rect 19228 9745 19234 9805
rect 19188 9733 19234 9745
rect 19348 9805 19394 9817
rect 19348 9745 19354 9805
rect 19388 9745 19394 9805
rect 19188 9667 19234 9679
rect 19188 9607 19194 9667
rect 19228 9607 19234 9667
rect 19188 9529 19234 9607
rect 19348 9667 19394 9745
rect 19348 9607 19354 9667
rect 19388 9607 19394 9667
rect 19348 9595 19394 9607
rect 19188 9469 19194 9529
rect 19228 9469 19234 9529
rect 19188 9457 19234 9469
rect 19348 9529 19394 9541
rect 19348 9469 19354 9529
rect 19388 9469 19394 9529
rect 19188 9391 19234 9403
rect 19188 9331 19194 9391
rect 19228 9331 19234 9391
rect 19188 9253 19234 9331
rect 19348 9391 19394 9469
rect 19348 9331 19354 9391
rect 19388 9331 19394 9391
rect 19348 9319 19394 9331
rect 19188 9193 19194 9253
rect 19228 9193 19234 9253
rect 19188 9181 19234 9193
rect 19348 9253 19394 9265
rect 19348 9193 19354 9253
rect 19388 9193 19394 9253
rect 19178 9115 19234 9127
rect 19178 9055 19194 9115
rect 19228 9055 19234 9115
rect 19178 9043 19234 9055
rect 19348 9115 19394 9193
rect 20132 9188 20293 9204
rect 20132 9136 20151 9188
rect 20203 9136 20293 9188
rect 20132 9120 20293 9136
rect 19348 9055 19354 9115
rect 19388 9055 19394 9115
rect 19348 9043 19394 9055
rect 20159 9068 20205 9080
rect 18276 9026 18334 9031
rect 19009 9029 19074 9030
rect 19009 9026 19015 9029
rect 14137 9015 14198 9021
rect 14137 8981 14152 9015
rect 14186 8981 14198 9015
rect 14137 8975 14198 8981
rect 14870 9015 15054 9021
rect 14870 8981 14886 9015
rect 14920 8981 15008 9015
rect 15042 8981 15054 9015
rect 14870 8975 15054 8981
rect 16208 9015 17604 9021
rect 16208 8981 16224 9015
rect 16258 8981 16346 9015
rect 16380 8981 17436 9015
rect 17470 8981 17558 9015
rect 17592 8981 17604 9015
rect 18276 9015 19015 9026
rect 18276 8996 18290 9015
rect 16208 8975 17604 8981
rect 18278 8981 18290 8996
rect 18324 8981 19015 9015
rect 18278 8979 19015 8981
rect 18278 8975 18336 8979
rect 19009 8977 19015 8979
rect 19067 8977 19074 9029
rect 14137 8972 14196 8975
rect 12019 8884 12025 8944
rect 12059 8884 12065 8944
rect 12019 8872 12065 8884
rect 12115 8944 12161 8956
rect 12115 8884 12121 8944
rect 12155 8884 12161 8944
rect 12115 8872 12161 8884
rect 12209 8944 12237 8945
rect 12209 8932 12273 8944
rect 12209 8872 12233 8932
rect 12267 8872 12273 8932
rect 12209 8860 12273 8872
rect 12315 8932 12361 8944
rect 12315 8872 12321 8932
rect 12355 8872 12361 8932
rect 12315 8860 12361 8872
rect 12410 8931 12474 8943
rect 12410 8871 12434 8931
rect 12468 8871 12474 8931
rect 12209 8827 12237 8860
rect 12410 8859 12474 8871
rect 12516 8931 12562 8943
rect 12516 8871 12522 8931
rect 12556 8871 12562 8931
rect 12516 8859 12562 8871
rect 13258 8930 13304 8970
rect 13258 8870 13264 8930
rect 13298 8870 13304 8930
rect 12410 8828 12438 8859
rect 13258 8858 13304 8870
rect 13332 8930 13422 8942
rect 13332 8926 13360 8930
rect 13394 8926 13422 8930
rect 13332 8874 13351 8926
rect 13403 8874 13422 8926
rect 13332 8870 13360 8874
rect 13394 8870 13422 8874
rect 13332 8858 13422 8870
rect 13450 8930 13496 8970
rect 13450 8870 13456 8930
rect 13490 8870 13496 8930
rect 13450 8858 13496 8870
rect 13538 8930 13584 8942
rect 14102 8934 14148 8943
rect 13538 8870 13544 8930
rect 13578 8870 13584 8930
rect 13538 8858 13584 8870
rect 14080 8933 14162 8934
rect 14080 8869 14089 8933
rect 14153 8869 14162 8933
rect 14191 8931 14237 8943
rect 14836 8934 14882 8943
rect 14191 8871 14197 8931
rect 14231 8871 14237 8931
rect 14102 8859 14148 8869
rect 12061 8821 12237 8827
rect 12061 8787 12073 8821
rect 12107 8787 12237 8821
rect 12061 8781 12237 8787
rect 12265 8822 12438 8828
rect 12579 8834 12643 8835
rect 12579 8827 12585 8834
rect 12265 8788 12277 8822
rect 12311 8788 12438 8822
rect 12265 8782 12438 8788
rect 12209 8741 12237 8781
rect 11826 8724 11833 8728
rect 8987 8639 9033 8679
rect 10437 8694 10495 8700
rect 3164 8630 3213 8634
rect 3602 8630 3660 8632
rect 3164 8629 3660 8630
rect 3733 8629 4179 8630
rect 3164 8626 3665 8629
rect 3164 8621 3614 8626
rect 3164 8587 3173 8621
rect 3207 8592 3614 8621
rect 3648 8592 3665 8626
rect 3207 8587 3665 8592
rect 3164 8583 3665 8587
rect 3733 8623 8154 8629
rect 3733 8589 4346 8623
rect 4380 8589 4472 8623
rect 4506 8589 5558 8623
rect 5592 8589 5684 8623
rect 5718 8589 6770 8623
rect 6804 8589 6896 8623
rect 6930 8589 7982 8623
rect 8016 8589 8108 8623
rect 8142 8589 8154 8623
rect 3733 8583 8154 8589
rect 8707 8601 8753 8613
rect 3164 8575 3213 8583
rect 3163 8536 3212 8541
rect 3733 8536 3782 8583
rect 8707 8541 8713 8601
rect 8747 8541 8753 8601
rect 8707 8538 8753 8541
rect 3163 8528 3782 8536
rect 3163 8494 3172 8528
rect 3206 8494 3782 8528
rect 3163 8489 3782 8494
rect 8706 8492 8753 8538
rect 8795 8610 9033 8639
rect 9333 8654 9386 8666
rect 10437 8660 10449 8694
rect 10483 8691 10495 8694
rect 11173 8694 11231 8700
rect 11173 8691 11185 8694
rect 10483 8663 11185 8691
rect 10483 8660 10495 8663
rect 10437 8654 10495 8660
rect 11173 8660 11185 8663
rect 11219 8691 11231 8694
rect 11541 8694 11599 8700
rect 11541 8691 11553 8694
rect 11219 8663 11553 8691
rect 11219 8660 11231 8663
rect 11173 8654 11231 8660
rect 11541 8660 11553 8663
rect 11587 8660 11599 8694
rect 11541 8654 11599 8660
rect 8795 8601 8841 8610
rect 8795 8541 8801 8601
rect 8835 8541 8841 8601
rect 9385 8601 9386 8654
rect 9333 8589 9386 8601
rect 8795 8529 8841 8541
rect 9061 8524 11709 8555
rect 3163 8482 3212 8489
rect 8706 8474 8871 8492
rect 8706 8433 8800 8474
rect 8781 8422 8800 8433
rect 8852 8422 8871 8474
rect 8781 8406 8871 8422
rect 9061 8490 9090 8524
rect 9124 8490 9182 8524
rect 9216 8490 9274 8524
rect 9308 8490 9346 8524
rect 9380 8490 9438 8524
rect 9472 8490 9530 8524
rect 9564 8490 9622 8524
rect 9656 8490 9714 8524
rect 9748 8490 9806 8524
rect 9840 8490 9898 8524
rect 9932 8490 9990 8524
rect 10024 8490 10082 8524
rect 10116 8490 10174 8524
rect 10208 8490 10266 8524
rect 10300 8490 10358 8524
rect 10392 8490 10450 8524
rect 10484 8490 10542 8524
rect 10576 8490 10634 8524
rect 10668 8490 10726 8524
rect 10760 8490 10818 8524
rect 10852 8490 10910 8524
rect 10944 8490 11002 8524
rect 11036 8490 11094 8524
rect 11128 8490 11186 8524
rect 11220 8490 11278 8524
rect 11312 8490 11370 8524
rect 11404 8490 11462 8524
rect 11496 8490 11554 8524
rect 11588 8490 11646 8524
rect 11680 8490 11709 8524
rect 9061 8459 11709 8490
rect 11827 8500 11833 8724
rect 11867 8724 11874 8728
rect 11923 8728 11969 8740
rect 11867 8500 11873 8724
rect 11827 8460 11873 8500
rect 11923 8500 11929 8728
rect 11963 8500 11969 8728
rect 11923 8488 11969 8500
rect 12019 8728 12065 8740
rect 12019 8500 12025 8728
rect 12059 8500 12065 8728
rect 12019 8460 12065 8500
rect 12115 8728 12161 8740
rect 12115 8500 12121 8728
rect 12155 8500 12161 8728
rect 12115 8488 12161 8500
rect 12209 8729 12273 8741
rect 12209 8501 12233 8729
rect 12267 8501 12273 8729
rect 12209 8489 12273 8501
rect 12315 8729 12361 8741
rect 12315 8501 12321 8729
rect 12355 8501 12361 8729
rect 12315 8489 12361 8501
rect 12410 8740 12438 8782
rect 12466 8821 12585 8827
rect 12466 8787 12478 8821
rect 12512 8787 12585 8821
rect 12466 8781 12585 8787
rect 12637 8781 12643 8834
rect 12671 8772 12677 8824
rect 12729 8772 12735 8824
rect 13071 8820 13454 8826
rect 13071 8786 13085 8820
rect 13119 8786 13408 8820
rect 13442 8816 13454 8820
rect 13538 8816 13566 8858
rect 13442 8787 13566 8816
rect 13442 8786 13454 8787
rect 13071 8780 13454 8786
rect 12410 8728 12474 8740
rect 12410 8472 12434 8728
rect 12468 8472 12474 8728
rect 12410 8460 12474 8472
rect 12516 8728 12562 8740
rect 13538 8739 13566 8787
rect 13599 8822 13661 8824
rect 14191 8822 14237 8871
rect 14814 8933 14896 8934
rect 14814 8869 14823 8933
rect 14887 8869 14896 8933
rect 14938 8931 14984 8943
rect 15046 8934 15092 8943
rect 16174 8934 16220 8943
rect 14938 8871 14944 8931
rect 14978 8871 14984 8931
rect 14836 8859 14882 8869
rect 14938 8822 14984 8871
rect 15032 8933 15114 8934
rect 15032 8869 15041 8933
rect 15105 8869 15114 8933
rect 16152 8933 16234 8934
rect 16152 8869 16161 8933
rect 16225 8869 16234 8933
rect 16278 8931 16324 8943
rect 16384 8934 16430 8943
rect 17386 8934 17432 8943
rect 16278 8871 16284 8931
rect 16318 8871 16324 8931
rect 15046 8859 15092 8869
rect 16174 8859 16220 8869
rect 16278 8822 16324 8871
rect 16370 8933 16452 8934
rect 16370 8869 16379 8933
rect 16443 8869 16452 8933
rect 17364 8933 17446 8934
rect 17364 8869 17373 8933
rect 17437 8869 17446 8933
rect 17489 8931 17535 8943
rect 17596 8934 17642 8943
rect 17489 8871 17495 8931
rect 17529 8871 17535 8931
rect 16384 8859 16430 8869
rect 17386 8859 17432 8869
rect 17489 8822 17535 8871
rect 17582 8933 17664 8934
rect 17582 8869 17591 8933
rect 17655 8869 17664 8933
rect 18238 8931 18284 8943
rect 18328 8934 18374 8943
rect 18238 8871 18244 8931
rect 18278 8871 18284 8931
rect 17596 8859 17642 8869
rect 18238 8822 18284 8871
rect 18314 8933 18396 8934
rect 18314 8869 18323 8933
rect 18387 8869 18396 8933
rect 18328 8859 18374 8869
rect 19178 8822 19224 9043
rect 13599 8818 19224 8822
rect 13599 8784 13615 8818
rect 13649 8784 19224 8818
rect 13599 8780 19224 8784
rect 13599 8778 13665 8780
rect 12516 8472 12522 8728
rect 12556 8542 12562 8728
rect 13258 8727 13304 8739
rect 13258 8667 13264 8727
rect 13298 8667 13304 8727
rect 12594 8642 12646 8648
rect 12593 8590 12594 8634
rect 12752 8634 12818 8640
rect 12923 8639 12975 8645
rect 12646 8630 12923 8634
rect 12646 8596 12767 8630
rect 12801 8596 12923 8630
rect 12646 8590 12923 8596
rect 12594 8584 12646 8590
rect 12922 8587 12923 8590
rect 12975 8587 12976 8631
rect 13258 8627 13304 8667
rect 13332 8727 13422 8739
rect 13332 8723 13360 8727
rect 13394 8723 13422 8727
rect 13332 8671 13351 8723
rect 13403 8671 13422 8723
rect 13332 8667 13360 8671
rect 13394 8667 13422 8671
rect 13332 8655 13422 8667
rect 13450 8727 13496 8739
rect 13450 8667 13456 8727
rect 13490 8667 13496 8727
rect 13450 8627 13496 8667
rect 13538 8727 13584 8739
rect 14099 8731 14145 8742
rect 13538 8667 13544 8727
rect 13578 8667 13584 8727
rect 13538 8655 13584 8667
rect 14076 8667 14083 8731
rect 14147 8667 14155 8731
rect 14076 8666 14155 8667
rect 14206 8730 14252 8780
rect 14313 8731 14359 8742
rect 15311 8731 15357 8742
rect 14206 8670 14212 8730
rect 14246 8670 14252 8730
rect 14099 8658 14145 8666
rect 14206 8658 14252 8670
rect 14303 8667 14311 8731
rect 14375 8667 14382 8731
rect 14303 8666 14382 8667
rect 15288 8667 15295 8731
rect 15359 8667 15367 8731
rect 15288 8666 15367 8667
rect 15420 8730 15466 8780
rect 15525 8731 15571 8742
rect 16523 8731 16569 8742
rect 15420 8670 15426 8730
rect 15460 8670 15466 8730
rect 14313 8658 14359 8666
rect 15311 8658 15357 8666
rect 15420 8658 15466 8670
rect 15515 8667 15523 8731
rect 15587 8667 15594 8731
rect 15515 8666 15594 8667
rect 16500 8667 16507 8731
rect 16571 8667 16579 8731
rect 16500 8666 16579 8667
rect 16633 8730 16679 8780
rect 16737 8731 16783 8742
rect 17735 8731 17781 8742
rect 16633 8670 16639 8730
rect 16673 8670 16679 8730
rect 15525 8658 15571 8666
rect 16523 8658 16569 8666
rect 16633 8658 16679 8670
rect 16727 8667 16735 8731
rect 16799 8667 16806 8731
rect 16727 8666 16806 8667
rect 17712 8667 17719 8731
rect 17783 8667 17791 8731
rect 17712 8666 17791 8667
rect 17844 8730 17890 8780
rect 17949 8731 17995 8742
rect 17844 8670 17850 8730
rect 17884 8670 17890 8730
rect 16737 8658 16783 8666
rect 17735 8658 17781 8666
rect 17844 8658 17890 8670
rect 17939 8667 17947 8731
rect 18011 8667 18018 8731
rect 17939 8666 18018 8667
rect 18593 8730 18639 8780
rect 18681 8734 18727 8745
rect 18593 8670 18599 8730
rect 18633 8670 18639 8730
rect 17949 8658 17995 8666
rect 18593 8658 18639 8670
rect 18671 8670 18679 8734
rect 18743 8670 18750 8734
rect 18671 8669 18750 8670
rect 18681 8661 18727 8669
rect 13258 8598 13496 8627
rect 18631 8618 18689 8620
rect 19078 8618 19127 8622
rect 18112 8617 18558 8618
rect 18631 8617 19127 8618
rect 14137 8611 18558 8617
rect 13450 8589 13496 8598
rect 12923 8581 12975 8587
rect 12556 8511 13201 8542
rect 13450 8529 13456 8589
rect 13490 8529 13496 8589
rect 13450 8517 13496 8529
rect 13538 8589 13584 8601
rect 13538 8529 13544 8589
rect 13578 8529 13584 8589
rect 14137 8577 14149 8611
rect 14183 8577 14275 8611
rect 14309 8577 15361 8611
rect 15395 8577 15487 8611
rect 15521 8577 16573 8611
rect 16607 8577 16699 8611
rect 16733 8577 17785 8611
rect 17819 8577 17911 8611
rect 17945 8577 18558 8611
rect 14137 8571 18558 8577
rect 18626 8614 19127 8617
rect 18626 8580 18643 8614
rect 18677 8609 19127 8614
rect 18677 8580 19084 8609
rect 18626 8575 19084 8580
rect 19118 8575 19127 8609
rect 18626 8571 19127 8575
rect 13538 8526 13584 8529
rect 12556 8477 12678 8511
rect 12712 8509 12770 8511
rect 12712 8477 12723 8509
rect 12804 8477 12862 8511
rect 12896 8477 12954 8511
rect 12988 8477 13046 8511
rect 13080 8509 13138 8511
rect 13080 8477 13097 8509
rect 13172 8477 13201 8511
rect 13538 8480 13585 8526
rect 12556 8472 12723 8477
rect 12516 8460 12723 8472
rect 9061 8449 10955 8459
rect 9061 8448 9472 8449
rect 9061 8396 9210 8448
rect 9262 8397 9472 8448
rect 9524 8397 9744 8449
rect 9796 8397 10071 8449
rect 10123 8397 10452 8449
rect 10504 8397 10829 8449
rect 10881 8397 10955 8449
rect 9262 8396 10955 8397
rect 9061 8380 10955 8396
rect 11771 8426 12065 8460
rect 12517 8456 12723 8460
rect 12776 8456 13097 8477
rect 13150 8469 13201 8477
rect 13150 8456 13202 8469
rect 12165 8439 12337 8449
rect 12517 8446 13202 8456
rect 12165 8427 12228 8439
rect 12281 8427 12337 8439
rect 9061 8377 11709 8380
rect 2577 8254 2894 8275
rect 2531 8247 2894 8254
rect 2922 8290 2968 8302
rect 2922 8230 2928 8290
rect 2962 8230 2968 8290
rect 2386 8153 2846 8176
rect 2386 8152 2582 8153
rect 2386 8145 2451 8152
rect 2386 8111 2415 8145
rect 2449 8111 2451 8145
rect 2386 8100 2451 8111
rect 2503 8145 2582 8152
rect 2634 8152 2846 8153
rect 2634 8145 2726 8152
rect 2503 8111 2507 8145
rect 2541 8111 2582 8145
rect 2634 8111 2691 8145
rect 2725 8111 2726 8145
rect 2503 8101 2582 8111
rect 2634 8101 2726 8111
rect 2503 8100 2726 8101
rect 2778 8145 2846 8152
rect 2778 8111 2783 8145
rect 2817 8111 2846 8145
rect 2778 8100 2846 8111
rect 2386 8080 2846 8100
rect 2922 8152 2968 8230
rect 3010 8290 3113 8302
rect 3010 8230 3016 8290
rect 3050 8230 3113 8290
rect 10054 8349 11709 8377
rect 10054 8315 10083 8349
rect 10117 8315 10175 8349
rect 10209 8315 10267 8349
rect 10301 8315 10359 8349
rect 10393 8315 10451 8349
rect 10485 8315 10543 8349
rect 10577 8315 10635 8349
rect 10669 8315 10727 8349
rect 10761 8315 10819 8349
rect 10853 8315 10910 8349
rect 10944 8315 11002 8349
rect 11036 8315 11094 8349
rect 11128 8315 11186 8349
rect 11220 8315 11278 8349
rect 11312 8315 11370 8349
rect 11404 8315 11462 8349
rect 11496 8315 11554 8349
rect 11588 8315 11646 8349
rect 11680 8315 11709 8349
rect 10054 8284 11709 8315
rect 3010 8218 3113 8230
rect 8863 8232 8953 8248
rect 8863 8180 8882 8232
rect 8934 8180 8953 8232
rect 8863 8164 8953 8180
rect 2922 8092 2928 8152
rect 2962 8092 2968 8152
rect 2922 8080 2968 8092
rect 3010 8152 3056 8164
rect 3010 8092 3016 8152
rect 3050 8092 3056 8152
rect 2922 8014 2968 8026
rect 2922 7954 2928 8014
rect 2962 7954 2968 8014
rect 2922 7876 2968 7954
rect 3010 8014 3056 8092
rect 10700 8121 10765 8124
rect 3010 7954 3016 8014
rect 3050 7954 3056 8014
rect 8864 8075 8954 8091
rect 8864 8023 8883 8075
rect 8935 8023 8954 8075
rect 10700 8069 10706 8121
rect 10758 8069 10765 8121
rect 10700 8067 10765 8069
rect 11518 8122 11590 8130
rect 11771 8122 11799 8426
rect 11518 8070 11524 8122
rect 11576 8070 11799 8122
rect 11518 8066 11799 8070
rect 11827 8364 12065 8398
rect 12165 8393 12200 8427
rect 12308 8393 12337 8427
rect 12165 8386 12228 8393
rect 12281 8386 12337 8393
rect 12518 8389 13202 8446
rect 13420 8462 13585 8480
rect 18509 8524 18558 8571
rect 19078 8563 19127 8571
rect 19079 8524 19128 8529
rect 18509 8516 19128 8524
rect 18509 8482 19085 8516
rect 19119 8482 19128 8516
rect 18509 8477 19128 8482
rect 19079 8470 19128 8477
rect 13420 8410 13439 8462
rect 13491 8421 13585 8462
rect 13491 8410 13510 8421
rect 13420 8394 13510 8410
rect 12165 8373 12337 8386
rect 11827 8324 11873 8364
rect 11827 8096 11833 8324
rect 11867 8096 11873 8324
rect 11518 8064 11590 8066
rect 8864 8007 8954 8023
rect 9333 8049 9398 8050
rect 9333 7996 9340 8049
rect 9392 8039 9398 8049
rect 11274 8042 11334 8049
rect 11274 8039 11286 8042
rect 9392 8011 11286 8039
rect 9392 7996 9398 8011
rect 11274 8008 11286 8011
rect 11320 8008 11334 8042
rect 11274 8003 11334 8008
rect 11279 8002 11333 8003
rect 3010 7942 3056 7954
rect 11827 7940 11873 8096
rect 11923 8324 11969 8336
rect 11923 8096 11929 8324
rect 11963 8096 11969 8324
rect 11923 8084 11969 8096
rect 12019 8324 12065 8364
rect 12425 8370 13202 8389
rect 12425 8369 12532 8370
rect 12019 8096 12025 8324
rect 12059 8096 12065 8324
rect 12019 8084 12065 8096
rect 12115 8324 12161 8336
rect 12425 8335 12452 8369
rect 12486 8336 12532 8369
rect 12566 8366 13202 8370
rect 12566 8336 12585 8366
rect 12486 8335 12585 8336
rect 12115 8096 12121 8324
rect 12155 8096 12161 8324
rect 12115 8084 12161 8096
rect 12209 8323 12273 8335
rect 12209 8095 12233 8323
rect 12267 8095 12273 8323
rect 12209 8083 12273 8095
rect 12315 8323 12361 8335
rect 12315 8095 12321 8323
rect 12355 8095 12361 8323
rect 12425 8313 12585 8335
rect 12638 8363 13202 8366
rect 12638 8313 12769 8363
rect 12425 8310 12769 8313
rect 12822 8357 13202 8363
rect 12822 8310 13071 8357
rect 12425 8304 13071 8310
rect 13124 8304 13202 8357
rect 12425 8231 13202 8304
rect 19178 8290 19224 8780
rect 19262 9005 19320 9011
rect 19262 8971 19274 9005
rect 19308 8971 19320 9005
rect 19496 8977 19503 9029
rect 19555 9026 19561 9029
rect 19555 8980 19659 9026
rect 20159 9008 20165 9068
rect 20199 9008 20205 9068
rect 20159 8999 20205 9008
rect 19555 8978 19657 8980
rect 19555 8977 19561 8978
rect 19496 8976 19561 8977
rect 19262 8965 19320 8971
rect 19967 8970 20205 8999
rect 20247 9068 20293 9120
rect 20247 9008 20253 9068
rect 20287 9008 20293 9068
rect 20247 8996 20293 9008
rect 20846 9021 20905 10153
rect 21206 10110 21538 10120
rect 21206 10058 21224 10110
rect 21276 10058 21304 10110
rect 21356 10058 21384 10110
rect 21436 10058 21464 10110
rect 21516 10058 21538 10110
rect 21206 10052 21538 10058
rect 21703 9021 21761 10381
rect 21808 10110 22140 10120
rect 21808 10058 21830 10110
rect 21882 10058 21910 10110
rect 21962 10058 21990 10110
rect 22042 10058 22070 10110
rect 22122 10058 22140 10110
rect 21808 10052 22140 10058
rect 22544 10110 22876 10120
rect 22544 10058 22562 10110
rect 22614 10058 22642 10110
rect 22694 10058 22722 10110
rect 22774 10058 22802 10110
rect 22854 10058 22876 10110
rect 22544 10052 22876 10058
rect 23146 10110 23478 10120
rect 23146 10058 23168 10110
rect 23220 10058 23248 10110
rect 23300 10058 23328 10110
rect 23380 10058 23408 10110
rect 23460 10058 23478 10110
rect 23146 10052 23478 10058
rect 23756 10110 24088 10120
rect 23756 10058 23774 10110
rect 23826 10058 23854 10110
rect 23906 10058 23934 10110
rect 23986 10058 24014 10110
rect 24066 10058 24088 10110
rect 23756 10052 24088 10058
rect 24129 9021 24187 10437
rect 24358 10110 24690 10120
rect 24358 10058 24380 10110
rect 24432 10058 24460 10110
rect 24512 10058 24540 10110
rect 24592 10058 24620 10110
rect 24672 10058 24690 10110
rect 24358 10052 24690 10058
rect 25090 10110 25422 10120
rect 25090 10058 25112 10110
rect 25164 10058 25192 10110
rect 25244 10058 25272 10110
rect 25324 10058 25352 10110
rect 25404 10058 25422 10110
rect 25090 10052 25422 10058
rect 25875 10113 25982 10129
rect 25875 10061 25894 10113
rect 25946 10061 25982 10113
rect 25875 10045 25903 10061
rect 25897 10021 25903 10045
rect 25937 10045 25982 10061
rect 26057 10081 26103 10093
rect 25937 10021 25943 10045
rect 25897 10009 25943 10021
rect 26057 10021 26063 10081
rect 26097 10021 26103 10081
rect 25897 9943 25943 9955
rect 25897 9883 25903 9943
rect 25937 9883 25943 9943
rect 25897 9805 25943 9883
rect 26057 9943 26103 10021
rect 26057 9883 26063 9943
rect 26097 9883 26103 9943
rect 26057 9871 26103 9883
rect 25897 9745 25903 9805
rect 25937 9745 25943 9805
rect 25897 9733 25943 9745
rect 26057 9805 26103 9817
rect 26057 9745 26063 9805
rect 26097 9745 26103 9805
rect 25897 9667 25943 9679
rect 25897 9607 25903 9667
rect 25937 9607 25943 9667
rect 25897 9529 25943 9607
rect 26057 9667 26103 9745
rect 26057 9607 26063 9667
rect 26097 9607 26103 9667
rect 26057 9595 26103 9607
rect 25897 9469 25903 9529
rect 25937 9469 25943 9529
rect 25897 9457 25943 9469
rect 26057 9529 26103 9541
rect 26057 9469 26063 9529
rect 26097 9469 26103 9529
rect 25897 9391 25943 9403
rect 25897 9331 25903 9391
rect 25937 9331 25943 9391
rect 25897 9253 25943 9331
rect 26057 9391 26103 9469
rect 26057 9331 26063 9391
rect 26097 9331 26103 9391
rect 26057 9319 26103 9331
rect 25897 9193 25903 9253
rect 25937 9193 25943 9253
rect 25897 9181 25943 9193
rect 26057 9253 26103 9265
rect 26057 9193 26063 9253
rect 26097 9193 26103 9253
rect 25887 9115 25943 9127
rect 25887 9055 25903 9115
rect 25937 9055 25943 9115
rect 25887 9043 25943 9055
rect 26057 9115 26103 9193
rect 26057 9055 26063 9115
rect 26097 9055 26103 9115
rect 26057 9043 26103 9055
rect 24985 9026 25043 9031
rect 25718 9029 25783 9030
rect 25718 9026 25724 9029
rect 20846 9015 20907 9021
rect 20846 8981 20861 9015
rect 20895 8981 20907 9015
rect 20846 8975 20907 8981
rect 21579 9015 21763 9021
rect 21579 8981 21595 9015
rect 21629 8981 21717 9015
rect 21751 8981 21763 9015
rect 21579 8975 21763 8981
rect 22917 9015 24313 9021
rect 22917 8981 22933 9015
rect 22967 8981 23055 9015
rect 23089 8981 24145 9015
rect 24179 8981 24267 9015
rect 24301 8981 24313 9015
rect 24985 9015 25724 9026
rect 24985 8996 24999 9015
rect 22917 8975 24313 8981
rect 24987 8981 24999 8996
rect 25033 8981 25724 9015
rect 24987 8979 25724 8981
rect 24987 8975 25045 8979
rect 25718 8977 25724 8979
rect 25776 8977 25783 9029
rect 20846 8972 20905 8975
rect 19262 8824 19310 8965
rect 19967 8930 20013 8970
rect 19967 8870 19973 8930
rect 20007 8870 20013 8930
rect 19967 8858 20013 8870
rect 20041 8930 20131 8942
rect 20041 8926 20069 8930
rect 20103 8926 20131 8930
rect 20041 8874 20060 8926
rect 20112 8874 20131 8926
rect 20041 8870 20069 8874
rect 20103 8870 20131 8874
rect 20041 8858 20131 8870
rect 20159 8930 20205 8970
rect 20159 8870 20165 8930
rect 20199 8870 20205 8930
rect 20159 8858 20205 8870
rect 20247 8930 20293 8942
rect 20811 8934 20857 8943
rect 20247 8870 20253 8930
rect 20287 8870 20293 8930
rect 20247 8858 20293 8870
rect 20789 8933 20871 8934
rect 20789 8869 20798 8933
rect 20862 8869 20871 8933
rect 20900 8931 20946 8943
rect 21545 8934 21591 8943
rect 20900 8871 20906 8931
rect 20940 8871 20946 8931
rect 20811 8859 20857 8869
rect 19920 8824 20163 8826
rect 19262 8820 20163 8824
rect 19262 8786 20117 8820
rect 20151 8816 20163 8820
rect 20247 8816 20275 8858
rect 20151 8787 20275 8816
rect 20151 8786 20163 8787
rect 19262 8780 20163 8786
rect 19262 8777 19982 8780
rect 19262 8377 19310 8777
rect 20247 8739 20275 8787
rect 20308 8822 20370 8824
rect 20900 8822 20946 8871
rect 21523 8933 21605 8934
rect 21523 8869 21532 8933
rect 21596 8869 21605 8933
rect 21647 8931 21693 8943
rect 21755 8934 21801 8943
rect 22883 8934 22929 8943
rect 21647 8871 21653 8931
rect 21687 8871 21693 8931
rect 21545 8859 21591 8869
rect 21647 8822 21693 8871
rect 21741 8933 21823 8934
rect 21741 8869 21750 8933
rect 21814 8869 21823 8933
rect 22861 8933 22943 8934
rect 22861 8869 22870 8933
rect 22934 8869 22943 8933
rect 22987 8931 23033 8943
rect 23093 8934 23139 8943
rect 24095 8934 24141 8943
rect 22987 8871 22993 8931
rect 23027 8871 23033 8931
rect 21755 8859 21801 8869
rect 22883 8859 22929 8869
rect 22987 8822 23033 8871
rect 23079 8933 23161 8934
rect 23079 8869 23088 8933
rect 23152 8869 23161 8933
rect 24073 8933 24155 8934
rect 24073 8869 24082 8933
rect 24146 8869 24155 8933
rect 24198 8931 24244 8943
rect 24305 8934 24351 8943
rect 24198 8871 24204 8931
rect 24238 8871 24244 8931
rect 23093 8859 23139 8869
rect 24095 8859 24141 8869
rect 24198 8822 24244 8871
rect 24291 8933 24373 8934
rect 24291 8869 24300 8933
rect 24364 8869 24373 8933
rect 24947 8931 24993 8943
rect 25037 8934 25083 8943
rect 24947 8871 24953 8931
rect 24987 8871 24993 8931
rect 24305 8859 24351 8869
rect 24947 8822 24993 8871
rect 25023 8933 25105 8934
rect 25023 8869 25032 8933
rect 25096 8869 25105 8933
rect 25037 8859 25083 8869
rect 25887 8822 25933 9043
rect 20308 8818 25933 8822
rect 20308 8784 20324 8818
rect 20358 8784 25933 8818
rect 20308 8780 25933 8784
rect 20308 8778 20374 8780
rect 19967 8727 20013 8739
rect 19445 8686 19905 8708
rect 19445 8677 19507 8686
rect 19559 8677 19650 8686
rect 19702 8677 19770 8686
rect 19822 8677 19905 8686
rect 19445 8643 19474 8677
rect 19559 8643 19566 8677
rect 19600 8643 19650 8677
rect 19702 8643 19750 8677
rect 19822 8643 19842 8677
rect 19876 8643 19905 8677
rect 19445 8634 19507 8643
rect 19559 8634 19650 8643
rect 19702 8634 19770 8643
rect 19822 8634 19905 8643
rect 19445 8612 19905 8634
rect 19967 8667 19973 8727
rect 20007 8667 20013 8727
rect 19967 8627 20013 8667
rect 20041 8727 20131 8739
rect 20041 8723 20069 8727
rect 20103 8723 20131 8727
rect 20041 8671 20060 8723
rect 20112 8671 20131 8723
rect 20041 8667 20069 8671
rect 20103 8667 20131 8671
rect 20041 8655 20131 8667
rect 20159 8727 20205 8739
rect 20159 8667 20165 8727
rect 20199 8667 20205 8727
rect 20159 8627 20205 8667
rect 20247 8727 20293 8739
rect 20808 8731 20854 8742
rect 20247 8667 20253 8727
rect 20287 8667 20293 8727
rect 20247 8655 20293 8667
rect 20785 8667 20792 8731
rect 20856 8667 20864 8731
rect 20785 8666 20864 8667
rect 20915 8730 20961 8780
rect 21022 8731 21068 8742
rect 22020 8731 22066 8742
rect 20915 8670 20921 8730
rect 20955 8670 20961 8730
rect 20808 8658 20854 8666
rect 20915 8658 20961 8670
rect 21012 8667 21020 8731
rect 21084 8667 21091 8731
rect 21012 8666 21091 8667
rect 21997 8667 22004 8731
rect 22068 8667 22076 8731
rect 21997 8666 22076 8667
rect 22129 8730 22175 8780
rect 22234 8731 22280 8742
rect 23232 8731 23278 8742
rect 22129 8670 22135 8730
rect 22169 8670 22175 8730
rect 21022 8658 21068 8666
rect 22020 8658 22066 8666
rect 22129 8658 22175 8670
rect 22224 8667 22232 8731
rect 22296 8667 22303 8731
rect 22224 8666 22303 8667
rect 23209 8667 23216 8731
rect 23280 8667 23288 8731
rect 23209 8666 23288 8667
rect 23342 8730 23388 8780
rect 23446 8731 23492 8742
rect 24444 8731 24490 8742
rect 23342 8670 23348 8730
rect 23382 8670 23388 8730
rect 22234 8658 22280 8666
rect 23232 8658 23278 8666
rect 23342 8658 23388 8670
rect 23436 8667 23444 8731
rect 23508 8667 23515 8731
rect 23436 8666 23515 8667
rect 24421 8667 24428 8731
rect 24492 8667 24500 8731
rect 24421 8666 24500 8667
rect 24553 8730 24599 8780
rect 24658 8731 24704 8742
rect 24553 8670 24559 8730
rect 24593 8670 24599 8730
rect 23446 8658 23492 8666
rect 24444 8658 24490 8666
rect 24553 8658 24599 8670
rect 24648 8667 24656 8731
rect 24720 8667 24727 8731
rect 24648 8666 24727 8667
rect 25302 8730 25348 8780
rect 25390 8734 25436 8745
rect 25302 8670 25308 8730
rect 25342 8670 25348 8730
rect 24658 8658 24704 8666
rect 25302 8658 25348 8670
rect 25380 8670 25388 8734
rect 25452 8670 25459 8734
rect 25380 8669 25459 8670
rect 25390 8661 25436 8669
rect 19967 8598 20205 8627
rect 25340 8618 25398 8620
rect 25787 8618 25836 8622
rect 24821 8617 25267 8618
rect 25340 8617 25836 8618
rect 20846 8611 25267 8617
rect 20159 8589 20205 8598
rect 19338 8534 19387 8547
rect 19338 8500 19344 8534
rect 19378 8510 19387 8534
rect 20159 8529 20165 8589
rect 20199 8529 20205 8589
rect 20159 8517 20205 8529
rect 20247 8589 20293 8601
rect 20247 8529 20253 8589
rect 20287 8529 20293 8589
rect 20846 8577 20858 8611
rect 20892 8577 20984 8611
rect 21018 8577 22070 8611
rect 22104 8577 22196 8611
rect 22230 8577 23282 8611
rect 23316 8577 23408 8611
rect 23442 8577 24494 8611
rect 24528 8577 24620 8611
rect 24654 8577 25267 8611
rect 20846 8571 25267 8577
rect 25335 8614 25836 8617
rect 25335 8580 25352 8614
rect 25386 8609 25836 8614
rect 25386 8580 25793 8609
rect 25335 8575 25793 8580
rect 25827 8575 25836 8609
rect 25335 8571 25836 8575
rect 20247 8526 20293 8529
rect 19378 8500 19481 8510
rect 19338 8482 19481 8500
rect 19376 8441 19425 8454
rect 19376 8407 19382 8441
rect 19416 8407 19425 8441
rect 19376 8395 19425 8407
rect 19262 8371 19331 8377
rect 19262 8337 19285 8371
rect 19319 8337 19331 8371
rect 19262 8331 19331 8337
rect 19178 8278 19281 8290
rect 12520 8230 13202 8231
rect 12709 8224 12793 8230
rect 12709 8190 12746 8224
rect 12780 8190 12793 8224
rect 12709 8184 12793 8190
rect 13338 8220 13428 8236
rect 13338 8168 13357 8220
rect 13409 8168 13428 8220
rect 19178 8218 19241 8278
rect 19275 8218 19281 8278
rect 19178 8206 19281 8218
rect 19323 8278 19369 8290
rect 19323 8218 19329 8278
rect 19363 8218 19369 8278
rect 19397 8263 19425 8395
rect 19453 8338 19481 8482
rect 20247 8480 20294 8526
rect 20129 8462 20294 8480
rect 25218 8524 25267 8571
rect 25787 8563 25836 8571
rect 25788 8524 25837 8529
rect 25218 8516 25837 8524
rect 25218 8482 25794 8516
rect 25828 8482 25837 8516
rect 25218 8477 25837 8482
rect 25788 8470 25837 8477
rect 19509 8451 19575 8452
rect 19509 8399 19515 8451
rect 19567 8399 19575 8451
rect 19784 8444 19838 8448
rect 19783 8441 19838 8444
rect 19783 8407 19795 8441
rect 19829 8407 19982 8441
rect 20129 8410 20148 8462
rect 20200 8421 20294 8462
rect 20200 8410 20219 8421
rect 19783 8404 19838 8407
rect 19783 8400 19837 8404
rect 19509 8397 19575 8399
rect 20129 8394 20219 8410
rect 19453 8331 19655 8338
rect 19453 8310 19605 8331
rect 19588 8297 19605 8310
rect 19639 8297 19655 8331
rect 19588 8291 19655 8297
rect 25887 8290 25933 8780
rect 25971 9005 26029 9011
rect 25971 8971 25983 9005
rect 26017 8971 26029 9005
rect 26205 8977 26212 9029
rect 26264 9026 26270 9029
rect 26264 8980 26368 9026
rect 26264 8978 26366 8980
rect 26264 8977 26270 8978
rect 26205 8976 26270 8977
rect 25971 8965 26029 8971
rect 25971 8824 26019 8965
rect 26658 8824 26704 12283
rect 25971 8777 26704 8824
rect 25971 8377 26019 8777
rect 26154 8686 26614 8708
rect 26154 8677 26216 8686
rect 26268 8677 26359 8686
rect 26411 8677 26479 8686
rect 26531 8677 26614 8686
rect 26154 8643 26183 8677
rect 26268 8643 26275 8677
rect 26309 8643 26359 8677
rect 26411 8643 26459 8677
rect 26531 8643 26551 8677
rect 26585 8643 26614 8677
rect 26154 8634 26216 8643
rect 26268 8634 26359 8643
rect 26411 8634 26479 8643
rect 26531 8634 26614 8643
rect 26154 8612 26614 8634
rect 26047 8534 26096 8547
rect 26047 8500 26053 8534
rect 26087 8510 26096 8534
rect 26087 8500 26190 8510
rect 26047 8482 26190 8500
rect 26085 8441 26134 8454
rect 26085 8407 26091 8441
rect 26125 8407 26134 8441
rect 26085 8395 26134 8407
rect 25971 8371 26040 8377
rect 25971 8337 25994 8371
rect 26028 8337 26040 8371
rect 25971 8331 26040 8337
rect 19702 8276 19760 8283
rect 19702 8263 19714 8276
rect 19397 8242 19714 8263
rect 19748 8242 19760 8276
rect 19397 8235 19760 8242
rect 25887 8278 25990 8290
rect 13338 8152 13428 8168
rect 12315 8083 12361 8095
rect 12696 8140 12742 8152
rect 12209 8043 12237 8083
rect 12696 8080 12702 8140
rect 12736 8080 12742 8140
rect 12696 8043 12742 8080
rect 12061 8037 12237 8043
rect 12061 8003 12073 8037
rect 12107 8003 12237 8037
rect 12061 7995 12237 8003
rect 12265 8036 12742 8043
rect 12265 8002 12277 8036
rect 12311 8002 12742 8036
rect 12265 7995 12742 8002
rect 12209 7964 12237 7995
rect 12209 7952 12273 7964
rect 8864 7905 8954 7921
rect 10451 7911 10506 7914
rect 10905 7912 10957 7914
rect 10902 7911 10957 7912
rect 2922 7816 2928 7876
rect 2962 7816 2968 7876
rect 2922 7804 2968 7816
rect 3010 7876 3056 7888
rect 3010 7816 3016 7876
rect 3050 7816 3056 7876
rect 8864 7853 8883 7905
rect 8935 7853 8954 7905
rect 8864 7837 8954 7853
rect 9961 7905 10125 7911
rect 9961 7871 10078 7905
rect 10112 7871 10125 7905
rect 9961 7865 10125 7871
rect 10451 7908 10957 7911
rect 10451 7874 10465 7908
rect 10499 7874 10910 7908
rect 10944 7874 10957 7908
rect 10451 7872 10957 7874
rect 10451 7869 10506 7872
rect 10451 7866 10505 7869
rect 10902 7867 10957 7872
rect 11827 7880 11833 7940
rect 11867 7880 11873 7940
rect 2922 7738 2968 7750
rect 2922 7678 2928 7738
rect 2962 7678 2968 7738
rect 2922 7600 2968 7678
rect 3010 7738 3056 7816
rect 3010 7678 3016 7738
rect 3050 7678 3056 7738
rect 8863 7753 8953 7769
rect 8863 7701 8882 7753
rect 8934 7701 8953 7753
rect 8863 7685 8953 7701
rect 3010 7666 3056 7678
rect 2922 7540 2928 7600
rect 2962 7540 2968 7600
rect 2922 7528 2968 7540
rect 3010 7600 3056 7612
rect 3010 7540 3016 7600
rect 3050 7594 3056 7600
rect 8858 7609 8948 7625
rect 3050 7564 3084 7594
rect 3050 7556 3728 7564
rect 3050 7547 3166 7556
rect 3050 7540 3068 7547
rect 3010 7528 3068 7540
rect 3031 7506 3068 7528
rect 3049 7495 3068 7506
rect 3120 7504 3166 7547
rect 3218 7504 3246 7556
rect 3298 7504 3326 7556
rect 3378 7504 3406 7556
rect 3458 7504 3486 7556
rect 3538 7504 3566 7556
rect 3618 7504 3728 7556
rect 3120 7498 3728 7504
rect 3790 7553 8698 7561
rect 3790 7501 3898 7553
rect 3950 7501 3978 7553
rect 4030 7501 4058 7553
rect 4110 7501 4138 7553
rect 4190 7501 4218 7553
rect 4270 7501 4298 7553
rect 4350 7501 4502 7553
rect 4554 7501 4582 7553
rect 4634 7501 4662 7553
rect 4714 7501 4742 7553
rect 4794 7501 4822 7553
rect 4874 7501 4902 7553
rect 4954 7501 5110 7553
rect 5162 7501 5190 7553
rect 5242 7501 5270 7553
rect 5322 7501 5350 7553
rect 5402 7501 5430 7553
rect 5482 7501 5510 7553
rect 5562 7501 5714 7553
rect 5766 7501 5794 7553
rect 5846 7501 5874 7553
rect 5926 7501 5954 7553
rect 6006 7501 6034 7553
rect 6086 7501 6114 7553
rect 6166 7501 6322 7553
rect 6374 7501 6402 7553
rect 6454 7501 6482 7553
rect 6534 7501 6562 7553
rect 6614 7501 6642 7553
rect 6694 7501 6722 7553
rect 6774 7501 6926 7553
rect 6978 7501 7006 7553
rect 7058 7501 7086 7553
rect 7138 7501 7166 7553
rect 7218 7501 7246 7553
rect 7298 7501 7326 7553
rect 7378 7501 7534 7553
rect 7586 7501 7614 7553
rect 7666 7501 7694 7553
rect 7746 7501 7774 7553
rect 7826 7501 7854 7553
rect 7906 7501 7934 7553
rect 7986 7501 8138 7553
rect 8190 7501 8218 7553
rect 8270 7501 8298 7553
rect 8350 7501 8378 7553
rect 8430 7501 8458 7553
rect 8510 7501 8538 7553
rect 8590 7501 8698 7553
rect 8858 7557 8877 7609
rect 8929 7557 8948 7609
rect 8858 7541 8948 7557
rect 3120 7495 3139 7498
rect 3790 7495 8698 7501
rect 3049 7479 3139 7495
rect 9961 7410 9995 7865
rect 11827 7855 11873 7880
rect 11923 7940 11969 7952
rect 11923 7880 11929 7940
rect 11963 7880 11969 7940
rect 11923 7868 11969 7880
rect 12019 7940 12065 7952
rect 12019 7880 12025 7940
rect 12059 7880 12065 7940
rect 11750 7849 11873 7855
rect 11368 7836 11407 7841
rect 10054 7805 11709 7836
rect 10054 7771 10083 7805
rect 10117 7771 10175 7805
rect 10209 7771 10267 7805
rect 10301 7771 10359 7805
rect 10393 7771 10451 7805
rect 10485 7771 10543 7805
rect 10577 7771 10635 7805
rect 10669 7771 10727 7805
rect 10761 7771 10819 7805
rect 10853 7771 10910 7805
rect 10944 7771 11002 7805
rect 11036 7771 11094 7805
rect 11128 7771 11186 7805
rect 11220 7771 11278 7805
rect 11312 7771 11370 7805
rect 11404 7771 11462 7805
rect 11496 7771 11554 7805
rect 11588 7771 11646 7805
rect 11680 7771 11709 7805
rect 11802 7840 11873 7849
rect 12019 7840 12065 7880
rect 12115 7940 12161 7952
rect 12115 7880 12121 7940
rect 12155 7880 12161 7940
rect 12209 7892 12233 7952
rect 12267 7892 12273 7952
rect 12209 7880 12273 7892
rect 12315 7952 12361 7964
rect 12315 7892 12321 7952
rect 12355 7892 12361 7952
rect 12315 7880 12361 7892
rect 12696 7952 12742 7995
rect 12115 7868 12161 7880
rect 11802 7806 12065 7840
rect 11750 7790 11802 7797
rect 10054 7725 11710 7771
rect 10054 7723 11035 7725
rect 10054 7691 10146 7723
rect 10110 7671 10146 7691
rect 10198 7691 10394 7723
rect 10198 7671 10217 7691
rect 10110 7655 10217 7671
rect 10358 7671 10394 7691
rect 10446 7691 10691 7723
rect 10446 7671 10465 7691
rect 10358 7655 10465 7671
rect 10655 7671 10691 7691
rect 10743 7691 11035 7723
rect 10743 7671 10762 7691
rect 10655 7655 10762 7671
rect 10999 7673 11035 7691
rect 11087 7691 11354 7725
rect 11087 7673 11106 7691
rect 10999 7657 11106 7673
rect 11318 7673 11354 7691
rect 11406 7691 11710 7725
rect 11928 7762 12355 7768
rect 11928 7728 11942 7762
rect 11976 7734 12014 7762
rect 12048 7728 12087 7762
rect 12121 7728 12159 7762
rect 12193 7761 12355 7762
rect 12193 7738 12232 7761
rect 12266 7738 12304 7761
rect 12193 7728 12220 7738
rect 11406 7673 11425 7691
rect 11318 7657 11425 7673
rect 11928 7690 11966 7728
rect 12018 7690 12220 7728
rect 12272 7727 12304 7738
rect 12338 7727 12355 7761
rect 11928 7656 11941 7690
rect 11975 7656 12013 7682
rect 12047 7656 12086 7690
rect 12120 7656 12158 7690
rect 12192 7686 12220 7690
rect 12272 7689 12355 7727
rect 12272 7686 12303 7689
rect 12192 7656 12231 7686
rect 11928 7655 12231 7656
rect 12265 7655 12303 7686
rect 12337 7655 12355 7689
rect 11928 7618 12355 7655
rect 11928 7584 11941 7618
rect 11975 7589 12013 7618
rect 11975 7584 11976 7589
rect 12047 7584 12086 7618
rect 12120 7584 12158 7618
rect 12192 7617 12355 7618
rect 12192 7592 12231 7617
rect 12265 7592 12303 7617
rect 12192 7584 12228 7592
rect 11928 7546 11976 7584
rect 12028 7546 12228 7584
rect 12280 7583 12303 7592
rect 12337 7583 12355 7617
rect 12696 7596 12702 7952
rect 12736 7596 12742 7952
rect 12696 7584 12742 7596
rect 12784 8140 12830 8152
rect 12784 8080 12790 8140
rect 12824 8080 12830 8140
rect 12784 8040 12830 8080
rect 19235 8140 19281 8152
rect 19235 8080 19241 8140
rect 19275 8080 19281 8140
rect 13337 8063 13427 8079
rect 12784 7990 12919 8040
rect 12784 7952 12830 7990
rect 12911 7987 12919 7990
rect 12971 7987 12977 8040
rect 13337 8011 13356 8063
rect 13408 8011 13427 8063
rect 13337 7995 13427 8011
rect 19235 8002 19281 8080
rect 19323 8140 19369 8218
rect 20047 8220 20137 8236
rect 20047 8168 20066 8220
rect 20118 8168 20137 8220
rect 25887 8218 25950 8278
rect 25984 8218 25990 8278
rect 25887 8206 25990 8218
rect 26032 8278 26078 8290
rect 26032 8218 26038 8278
rect 26072 8218 26078 8278
rect 26106 8263 26134 8395
rect 26162 8338 26190 8482
rect 26218 8451 26284 8452
rect 26218 8399 26224 8451
rect 26276 8399 26284 8451
rect 26493 8444 26547 8448
rect 26492 8441 26547 8444
rect 26492 8407 26504 8441
rect 26538 8407 26685 8441
rect 26492 8404 26547 8407
rect 26492 8400 26546 8404
rect 26218 8397 26284 8399
rect 26162 8331 26364 8338
rect 26162 8310 26314 8331
rect 26297 8297 26314 8310
rect 26348 8297 26364 8331
rect 26297 8291 26364 8297
rect 26411 8276 26469 8283
rect 26411 8263 26423 8276
rect 26106 8242 26423 8263
rect 26457 8242 26469 8276
rect 26106 8235 26469 8242
rect 19323 8080 19329 8140
rect 19363 8080 19369 8140
rect 19323 8068 19369 8080
rect 19445 8141 19905 8164
rect 20047 8152 20137 8168
rect 19445 8140 19657 8141
rect 19445 8133 19513 8140
rect 19445 8099 19474 8133
rect 19508 8099 19513 8133
rect 19445 8088 19513 8099
rect 19565 8133 19657 8140
rect 19709 8140 19905 8141
rect 19709 8133 19788 8140
rect 19565 8099 19566 8133
rect 19600 8099 19657 8133
rect 19709 8099 19750 8133
rect 19784 8099 19788 8133
rect 19565 8089 19657 8099
rect 19709 8089 19788 8099
rect 19565 8088 19788 8089
rect 19840 8133 19905 8140
rect 19840 8099 19842 8133
rect 19876 8099 19905 8133
rect 19840 8088 19905 8099
rect 19445 8068 19905 8088
rect 25944 8140 25990 8152
rect 25944 8080 25950 8140
rect 25984 8080 25990 8140
rect 20046 8063 20136 8079
rect 12911 7986 12977 7987
rect 12784 7596 12790 7952
rect 12824 7596 12830 7952
rect 12921 7929 13011 7945
rect 19235 7942 19241 8002
rect 19275 7942 19281 8002
rect 19235 7930 19281 7942
rect 19323 8002 19369 8014
rect 20046 8011 20065 8063
rect 20117 8011 20136 8063
rect 19323 7942 19329 8002
rect 19363 7942 19369 8002
rect 12921 7877 12940 7929
rect 12992 7877 13011 7929
rect 12921 7861 13011 7877
rect 13337 7893 13427 7909
rect 13337 7841 13356 7893
rect 13408 7841 13427 7893
rect 13337 7825 13427 7841
rect 19235 7864 19281 7876
rect 19235 7804 19241 7864
rect 19275 7804 19281 7864
rect 13338 7741 13428 7757
rect 12913 7709 13003 7725
rect 12913 7657 12932 7709
rect 12984 7657 13003 7709
rect 13338 7689 13357 7741
rect 13409 7689 13428 7741
rect 13338 7673 13428 7689
rect 19235 7726 19281 7804
rect 19323 7864 19369 7942
rect 19624 7991 19714 8007
rect 20046 7995 20136 8011
rect 25944 8002 25990 8080
rect 26032 8140 26078 8218
rect 26032 8080 26038 8140
rect 26072 8080 26078 8140
rect 26032 8068 26078 8080
rect 26154 8141 26614 8164
rect 26154 8140 26366 8141
rect 26154 8133 26222 8140
rect 26154 8099 26183 8133
rect 26217 8099 26222 8133
rect 26154 8088 26222 8099
rect 26274 8133 26366 8140
rect 26418 8140 26614 8141
rect 26418 8133 26497 8140
rect 26274 8099 26275 8133
rect 26309 8099 26366 8133
rect 26418 8099 26459 8133
rect 26493 8099 26497 8133
rect 26274 8089 26366 8099
rect 26418 8089 26497 8099
rect 26274 8088 26497 8089
rect 26549 8133 26614 8140
rect 26549 8099 26551 8133
rect 26585 8099 26614 8133
rect 26549 8088 26614 8099
rect 26154 8068 26614 8088
rect 19624 7939 19643 7991
rect 19695 7939 19714 7991
rect 19624 7923 19714 7939
rect 25944 7942 25950 8002
rect 25984 7942 25990 8002
rect 25944 7930 25990 7942
rect 26032 8002 26078 8014
rect 26032 7942 26038 8002
rect 26072 7942 26078 8002
rect 19323 7804 19329 7864
rect 19363 7804 19369 7864
rect 20046 7893 20136 7909
rect 20046 7841 20065 7893
rect 20117 7841 20136 7893
rect 20046 7825 20136 7841
rect 25944 7864 25990 7876
rect 19323 7792 19369 7804
rect 19624 7795 19714 7811
rect 19624 7743 19643 7795
rect 19695 7743 19714 7795
rect 25944 7804 25950 7864
rect 25984 7804 25990 7864
rect 12913 7641 13003 7657
rect 19235 7666 19241 7726
rect 19275 7666 19281 7726
rect 19235 7654 19281 7666
rect 19323 7726 19369 7738
rect 19624 7727 19714 7743
rect 20047 7741 20137 7757
rect 19323 7666 19329 7726
rect 19363 7666 19369 7726
rect 20047 7689 20066 7741
rect 20118 7689 20137 7741
rect 20047 7673 20137 7689
rect 25944 7726 25990 7804
rect 26032 7864 26078 7942
rect 26032 7804 26038 7864
rect 26072 7804 26078 7864
rect 26032 7792 26078 7804
rect 12784 7584 12830 7596
rect 13343 7597 13433 7613
rect 10305 7481 10311 7533
rect 10363 7522 10369 7533
rect 11743 7522 11749 7532
rect 10363 7494 11749 7522
rect 10363 7481 10369 7494
rect 11743 7480 11749 7494
rect 11801 7480 11807 7532
rect 11928 7512 11940 7546
rect 11974 7537 11976 7546
rect 11974 7512 12012 7537
rect 12046 7512 12085 7546
rect 12119 7512 12157 7546
rect 12191 7540 12228 7546
rect 12280 7548 12355 7583
rect 12280 7545 12790 7548
rect 12280 7540 12302 7545
rect 12191 7512 12230 7540
rect 11928 7511 12230 7512
rect 12264 7511 12302 7540
rect 12336 7543 12790 7545
rect 13343 7545 13362 7597
rect 13414 7545 13433 7597
rect 19235 7588 19281 7600
rect 19235 7582 19241 7588
rect 19207 7552 19241 7582
rect 12336 7537 12792 7543
rect 12336 7511 12746 7537
rect 11928 7503 12746 7511
rect 12780 7503 12792 7537
rect 13343 7529 13433 7545
rect 13593 7541 18501 7549
rect 11928 7497 12792 7503
rect 11928 7492 12790 7497
rect 13593 7489 13701 7541
rect 13753 7489 13781 7541
rect 13833 7489 13861 7541
rect 13913 7489 13941 7541
rect 13993 7489 14021 7541
rect 14073 7489 14101 7541
rect 14153 7489 14305 7541
rect 14357 7489 14385 7541
rect 14437 7489 14465 7541
rect 14517 7489 14545 7541
rect 14597 7489 14625 7541
rect 14677 7489 14705 7541
rect 14757 7489 14913 7541
rect 14965 7489 14993 7541
rect 15045 7489 15073 7541
rect 15125 7489 15153 7541
rect 15205 7489 15233 7541
rect 15285 7489 15313 7541
rect 15365 7489 15517 7541
rect 15569 7489 15597 7541
rect 15649 7489 15677 7541
rect 15729 7489 15757 7541
rect 15809 7489 15837 7541
rect 15889 7489 15917 7541
rect 15969 7489 16125 7541
rect 16177 7489 16205 7541
rect 16257 7489 16285 7541
rect 16337 7489 16365 7541
rect 16417 7489 16445 7541
rect 16497 7489 16525 7541
rect 16577 7489 16729 7541
rect 16781 7489 16809 7541
rect 16861 7489 16889 7541
rect 16941 7489 16969 7541
rect 17021 7489 17049 7541
rect 17101 7489 17129 7541
rect 17181 7489 17337 7541
rect 17389 7489 17417 7541
rect 17469 7489 17497 7541
rect 17549 7489 17577 7541
rect 17629 7489 17657 7541
rect 17709 7489 17737 7541
rect 17789 7489 17941 7541
rect 17993 7489 18021 7541
rect 18073 7489 18101 7541
rect 18153 7489 18181 7541
rect 18233 7489 18261 7541
rect 18313 7489 18341 7541
rect 18393 7489 18501 7541
rect 13593 7483 18501 7489
rect 18563 7544 19241 7552
rect 18563 7492 18673 7544
rect 18725 7492 18753 7544
rect 18805 7492 18833 7544
rect 18885 7492 18913 7544
rect 18965 7492 18993 7544
rect 19045 7492 19073 7544
rect 19125 7535 19241 7544
rect 19125 7492 19171 7535
rect 18563 7486 19171 7492
rect 19152 7483 19171 7486
rect 19223 7528 19241 7535
rect 19275 7528 19281 7588
rect 19223 7516 19281 7528
rect 19323 7588 19369 7666
rect 25944 7666 25950 7726
rect 25984 7666 25990 7726
rect 25944 7654 25990 7666
rect 26032 7726 26078 7738
rect 26032 7666 26038 7726
rect 26072 7666 26078 7726
rect 19323 7528 19329 7588
rect 19363 7528 19369 7588
rect 19624 7620 19714 7636
rect 19624 7568 19643 7620
rect 19695 7568 19714 7620
rect 19624 7552 19714 7568
rect 20052 7597 20142 7613
rect 20052 7545 20071 7597
rect 20123 7545 20142 7597
rect 25944 7588 25990 7600
rect 25944 7582 25950 7588
rect 25916 7552 25950 7582
rect 20052 7529 20142 7545
rect 20302 7541 25210 7549
rect 19323 7516 19369 7528
rect 19223 7494 19260 7516
rect 19223 7483 19242 7494
rect 20302 7489 20410 7541
rect 20462 7489 20490 7541
rect 20542 7489 20570 7541
rect 20622 7489 20650 7541
rect 20702 7489 20730 7541
rect 20782 7489 20810 7541
rect 20862 7489 21014 7541
rect 21066 7489 21094 7541
rect 21146 7489 21174 7541
rect 21226 7489 21254 7541
rect 21306 7489 21334 7541
rect 21386 7489 21414 7541
rect 21466 7489 21622 7541
rect 21674 7489 21702 7541
rect 21754 7489 21782 7541
rect 21834 7489 21862 7541
rect 21914 7489 21942 7541
rect 21994 7489 22022 7541
rect 22074 7489 22226 7541
rect 22278 7489 22306 7541
rect 22358 7489 22386 7541
rect 22438 7489 22466 7541
rect 22518 7489 22546 7541
rect 22598 7489 22626 7541
rect 22678 7489 22834 7541
rect 22886 7489 22914 7541
rect 22966 7489 22994 7541
rect 23046 7489 23074 7541
rect 23126 7489 23154 7541
rect 23206 7489 23234 7541
rect 23286 7489 23438 7541
rect 23490 7489 23518 7541
rect 23570 7489 23598 7541
rect 23650 7489 23678 7541
rect 23730 7489 23758 7541
rect 23810 7489 23838 7541
rect 23890 7489 24046 7541
rect 24098 7489 24126 7541
rect 24178 7489 24206 7541
rect 24258 7489 24286 7541
rect 24338 7489 24366 7541
rect 24418 7489 24446 7541
rect 24498 7489 24650 7541
rect 24702 7489 24730 7541
rect 24782 7489 24810 7541
rect 24862 7489 24890 7541
rect 24942 7489 24970 7541
rect 25022 7489 25050 7541
rect 25102 7489 25210 7541
rect 20302 7483 25210 7489
rect 25272 7544 25950 7552
rect 25272 7492 25382 7544
rect 25434 7492 25462 7544
rect 25514 7492 25542 7544
rect 25594 7492 25622 7544
rect 25674 7492 25702 7544
rect 25754 7492 25782 7544
rect 25834 7535 25950 7544
rect 25834 7492 25880 7535
rect 25272 7486 25880 7492
rect 25861 7483 25880 7486
rect 25932 7528 25950 7535
rect 25984 7528 25990 7588
rect 25932 7516 25990 7528
rect 26032 7588 26078 7666
rect 26032 7528 26038 7588
rect 26072 7528 26078 7588
rect 26032 7516 26078 7528
rect 25932 7494 25969 7516
rect 25932 7483 25951 7494
rect 19152 7467 19242 7483
rect 25861 7467 25951 7483
rect 2978 7358 2985 7410
rect 3038 7401 3044 7410
rect 9945 7401 9951 7410
rect 3038 7367 9951 7401
rect 3038 7358 3044 7367
rect 9945 7358 9951 7367
rect 10003 7358 10009 7410
rect 10623 7282 10629 7334
rect 10681 7323 10687 7334
rect 23915 7323 23921 7333
rect 10681 7295 23921 7323
rect 10681 7282 10687 7295
rect 10623 7281 10687 7282
rect 23915 7281 23921 7295
rect 23973 7281 23979 7333
rect 24662 7329 24752 7345
rect 24662 7318 24681 7329
rect 24644 7296 24681 7318
rect 23915 7280 23979 7281
rect 24535 7284 24581 7296
rect 24535 7224 24541 7284
rect 24575 7224 24581 7284
rect 24535 7146 24581 7224
rect 24623 7284 24681 7296
rect 24623 7224 24629 7284
rect 24663 7277 24681 7284
rect 24733 7326 24752 7329
rect 24733 7320 25341 7326
rect 24733 7277 24779 7320
rect 24663 7268 24779 7277
rect 24831 7268 24859 7320
rect 24911 7268 24939 7320
rect 24991 7268 25019 7320
rect 25071 7268 25099 7320
rect 25151 7268 25179 7320
rect 25231 7268 25341 7320
rect 24663 7260 25341 7268
rect 25403 7323 30311 7329
rect 25403 7271 25511 7323
rect 25563 7271 25591 7323
rect 25643 7271 25671 7323
rect 25723 7271 25751 7323
rect 25803 7271 25831 7323
rect 25883 7271 25911 7323
rect 25963 7271 26115 7323
rect 26167 7271 26195 7323
rect 26247 7271 26275 7323
rect 26327 7271 26355 7323
rect 26407 7271 26435 7323
rect 26487 7271 26515 7323
rect 26567 7271 26723 7323
rect 26775 7271 26803 7323
rect 26855 7271 26883 7323
rect 26935 7271 26963 7323
rect 27015 7271 27043 7323
rect 27095 7271 27123 7323
rect 27175 7271 27327 7323
rect 27379 7271 27407 7323
rect 27459 7271 27487 7323
rect 27539 7271 27567 7323
rect 27619 7271 27647 7323
rect 27699 7271 27727 7323
rect 27779 7271 27935 7323
rect 27987 7271 28015 7323
rect 28067 7271 28095 7323
rect 28147 7271 28175 7323
rect 28227 7271 28255 7323
rect 28307 7271 28335 7323
rect 28387 7271 28539 7323
rect 28591 7271 28619 7323
rect 28671 7271 28699 7323
rect 28751 7271 28779 7323
rect 28831 7271 28859 7323
rect 28911 7271 28939 7323
rect 28991 7271 29147 7323
rect 29199 7271 29227 7323
rect 29279 7271 29307 7323
rect 29359 7271 29387 7323
rect 29439 7271 29467 7323
rect 29519 7271 29547 7323
rect 29599 7271 29751 7323
rect 29803 7271 29831 7323
rect 29883 7271 29911 7323
rect 29963 7271 29991 7323
rect 30043 7271 30071 7323
rect 30123 7271 30151 7323
rect 30203 7271 30311 7323
rect 25403 7263 30311 7271
rect 30471 7267 30561 7283
rect 24663 7230 24697 7260
rect 24663 7224 24669 7230
rect 24623 7212 24669 7224
rect 30471 7215 30490 7267
rect 30542 7215 30561 7267
rect 30471 7199 30561 7215
rect 11075 7124 14777 7125
rect 10753 7094 14777 7124
rect 10753 7080 11527 7094
rect 10753 6934 10891 7080
rect 11041 7064 11527 7080
rect 11041 6934 11203 7064
rect 10753 6918 11203 6934
rect 11353 7060 11527 7064
rect 11561 7060 11619 7094
rect 11653 7060 11711 7094
rect 11745 7060 11803 7094
rect 11837 7060 11895 7094
rect 11929 7060 11987 7094
rect 12021 7060 12079 7094
rect 12113 7060 12171 7094
rect 12205 7060 12263 7094
rect 12297 7060 12787 7094
rect 12821 7060 12879 7094
rect 12913 7060 12971 7094
rect 13005 7060 13063 7094
rect 13097 7060 13155 7094
rect 13189 7060 13247 7094
rect 13281 7060 13339 7094
rect 13373 7060 13431 7094
rect 13465 7060 13523 7094
rect 13557 7060 13615 7094
rect 13649 7060 13707 7094
rect 13741 7060 13799 7094
rect 13833 7060 13891 7094
rect 13925 7060 13983 7094
rect 14017 7060 14075 7094
rect 14109 7060 14167 7094
rect 14201 7060 14259 7094
rect 14293 7060 14351 7094
rect 14385 7060 14443 7094
rect 14477 7060 14535 7094
rect 14569 7060 14777 7094
rect 24535 7086 24541 7146
rect 24575 7086 24581 7146
rect 24535 7074 24581 7086
rect 24623 7146 24669 7158
rect 24623 7086 24629 7146
rect 24663 7086 24669 7146
rect 11353 7029 14777 7060
rect 11353 6918 11417 7029
rect 24535 7008 24581 7020
rect 13234 6992 13292 6998
rect 13234 6958 13246 6992
rect 13280 6989 13292 6992
rect 13694 6992 13752 6998
rect 13694 6989 13706 6992
rect 13280 6961 13706 6989
rect 13280 6958 13292 6961
rect 13234 6952 13292 6958
rect 13694 6958 13706 6961
rect 13740 6958 13752 6992
rect 13694 6952 13752 6958
rect 13878 6992 13936 6998
rect 13878 6958 13890 6992
rect 13924 6989 13936 6992
rect 14154 6992 14212 6998
rect 14154 6989 14166 6992
rect 13924 6961 14166 6989
rect 13924 6958 13936 6961
rect 13878 6952 13936 6958
rect 14154 6958 14166 6961
rect 14200 6958 14212 6992
rect 14154 6952 14212 6958
rect 24535 6948 24541 7008
rect 24575 6948 24581 7008
rect 10753 6894 11417 6918
rect 13418 6924 13476 6930
rect 13418 6890 13430 6924
rect 13464 6921 13476 6924
rect 14246 6924 14304 6930
rect 14246 6921 14258 6924
rect 13464 6893 14258 6921
rect 13464 6890 13476 6893
rect 13418 6884 13476 6890
rect 14246 6890 14258 6893
rect 14292 6890 14304 6924
rect 14246 6884 14304 6890
rect 24535 6870 24581 6948
rect 24623 7008 24669 7086
rect 30476 7123 30566 7139
rect 30476 7071 30495 7123
rect 30547 7071 30566 7123
rect 30476 7055 30566 7071
rect 24623 6948 24629 7008
rect 24663 6948 24669 7008
rect 24623 6936 24669 6948
rect 30477 6971 30567 6987
rect 30477 6919 30496 6971
rect 30548 6919 30567 6971
rect 30477 6903 30567 6919
rect 10922 6853 10956 6858
rect 13326 6856 13384 6862
rect 13326 6853 13338 6856
rect 10922 6825 13338 6853
rect 10922 6824 10956 6825
rect 13326 6822 13338 6825
rect 13372 6853 13384 6856
rect 14338 6856 14396 6862
rect 14338 6853 14350 6856
rect 13372 6825 14350 6853
rect 13372 6822 13384 6825
rect 13326 6816 13384 6822
rect 14338 6822 14350 6825
rect 14384 6853 14396 6856
rect 14522 6856 14581 6862
rect 14522 6853 14534 6856
rect 14384 6825 14534 6853
rect 14384 6822 14396 6825
rect 14338 6816 14396 6822
rect 14522 6822 14534 6825
rect 14568 6822 14581 6856
rect 14522 6816 14581 6822
rect 18583 6809 18636 6816
rect 9982 6744 9988 6796
rect 10040 6788 10046 6796
rect 11519 6789 11585 6796
rect 10040 6787 10959 6788
rect 11519 6787 11531 6789
rect 10040 6759 11531 6787
rect 10040 6754 10959 6759
rect 11519 6755 11531 6759
rect 11565 6755 11585 6789
rect 10040 6744 10046 6754
rect 11519 6744 11585 6755
rect 12153 6745 12160 6797
rect 12212 6745 12221 6797
rect 12476 6796 12542 6797
rect 12476 6744 12483 6796
rect 12535 6782 12542 6796
rect 12860 6787 12918 6792
rect 13587 6790 13647 6796
rect 12860 6786 12920 6787
rect 12860 6782 12873 6786
rect 12535 6754 12873 6782
rect 12535 6744 12542 6754
rect 12860 6752 12873 6754
rect 12907 6752 12920 6786
rect 12860 6751 12920 6752
rect 13587 6756 13601 6790
rect 13635 6787 13647 6790
rect 13635 6759 18583 6787
rect 13635 6756 13647 6759
rect 12860 6746 12918 6751
rect 13587 6746 13647 6756
rect 18635 6757 18636 6809
rect 24535 6810 24541 6870
rect 24575 6810 24581 6870
rect 24535 6798 24581 6810
rect 24623 6870 24669 6882
rect 24623 6810 24629 6870
rect 24663 6810 24669 6870
rect 18583 6750 18636 6757
rect 20991 6733 21044 6740
rect 10927 6716 10962 6722
rect 13966 6719 14029 6726
rect 13966 6716 13982 6719
rect 10926 6688 13982 6716
rect 10927 6687 10962 6688
rect 13966 6685 13982 6688
rect 14016 6685 14029 6719
rect 13966 6678 14029 6685
rect 14059 6675 14065 6727
rect 14117 6675 14123 6727
rect 14190 6693 20991 6721
rect 13229 6649 13288 6656
rect 13229 6615 13241 6649
rect 13275 6637 13288 6649
rect 14190 6647 14219 6693
rect 21043 6681 21044 6733
rect 20991 6674 21044 6681
rect 23999 6724 24459 6744
rect 23999 6713 24064 6724
rect 23999 6679 24028 6713
rect 24062 6679 24064 6713
rect 23999 6672 24064 6679
rect 24116 6723 24339 6724
rect 24116 6713 24195 6723
rect 24247 6713 24339 6723
rect 24116 6679 24120 6713
rect 24154 6679 24195 6713
rect 24247 6679 24304 6713
rect 24338 6679 24339 6713
rect 24116 6672 24195 6679
rect 23999 6671 24195 6672
rect 24247 6672 24339 6679
rect 24391 6713 24459 6724
rect 24391 6679 24396 6713
rect 24430 6679 24459 6713
rect 24391 6672 24459 6679
rect 24247 6671 24459 6672
rect 14190 6637 14218 6647
rect 13275 6615 14218 6637
rect 13229 6609 14218 6615
rect 14338 6613 14345 6665
rect 14397 6640 14404 6665
rect 16187 6640 16194 6665
rect 14397 6613 16194 6640
rect 16246 6613 16253 6665
rect 23999 6648 24459 6671
rect 24535 6732 24581 6744
rect 24535 6672 24541 6732
rect 24575 6672 24581 6732
rect 14338 6612 16253 6613
rect 24535 6594 24581 6672
rect 24623 6732 24669 6810
rect 30477 6801 30567 6817
rect 30477 6749 30496 6801
rect 30548 6749 30567 6801
rect 30477 6733 30567 6749
rect 24623 6672 24629 6732
rect 24663 6672 24669 6732
rect 24623 6660 24669 6672
rect 30476 6644 30566 6660
rect 10965 6581 11045 6582
rect 10883 6571 22502 6581
rect 22741 6571 23795 6578
rect 10883 6550 23795 6571
rect 10883 6546 11527 6550
rect 10879 6516 11527 6546
rect 11561 6516 11619 6550
rect 11653 6516 11711 6550
rect 11745 6516 11803 6550
rect 11837 6516 11895 6550
rect 11929 6516 11987 6550
rect 12021 6516 12079 6550
rect 12113 6516 12171 6550
rect 12205 6516 12263 6550
rect 12297 6516 12787 6550
rect 12821 6516 12879 6550
rect 12913 6516 12971 6550
rect 13005 6516 13063 6550
rect 13097 6516 13155 6550
rect 13189 6516 13247 6550
rect 13281 6516 13339 6550
rect 13373 6516 13431 6550
rect 13465 6516 13523 6550
rect 13557 6516 13615 6550
rect 13649 6516 13707 6550
rect 13741 6516 13799 6550
rect 13833 6516 13891 6550
rect 13925 6516 13983 6550
rect 14017 6516 14075 6550
rect 14109 6516 14167 6550
rect 14201 6516 14259 6550
rect 14293 6516 14351 6550
rect 14385 6516 14443 6550
rect 14477 6516 14535 6550
rect 14569 6516 23795 6550
rect 24144 6570 24507 6577
rect 24144 6536 24156 6570
rect 24190 6549 24507 6570
rect 24190 6536 24202 6549
rect 24144 6529 24202 6536
rect 10879 6508 23795 6516
rect 10883 6495 23795 6508
rect 10883 6485 22502 6495
rect 23545 6466 23795 6495
rect 24249 6515 24316 6521
rect 24249 6481 24265 6515
rect 24299 6502 24316 6515
rect 24299 6481 24451 6502
rect 24249 6474 24451 6481
rect 11516 6422 11582 6423
rect 11516 6411 11523 6422
rect 11502 6383 11523 6411
rect 11516 6370 11523 6383
rect 11575 6411 11582 6422
rect 12177 6422 12243 6423
rect 12177 6411 12184 6422
rect 11575 6383 12184 6411
rect 11575 6370 11582 6383
rect 12177 6370 12184 6383
rect 12236 6411 12243 6422
rect 13907 6422 13973 6423
rect 13907 6411 13914 6422
rect 12236 6383 13914 6411
rect 12236 6370 12243 6383
rect 13907 6370 13914 6383
rect 13966 6411 13973 6422
rect 16290 6422 16356 6423
rect 16290 6411 16297 6422
rect 13966 6383 16297 6411
rect 13966 6370 13973 6383
rect 16290 6370 16297 6383
rect 16349 6411 16356 6422
rect 18685 6422 18751 6423
rect 18685 6411 18692 6422
rect 16349 6383 18692 6411
rect 16349 6370 16356 6383
rect 18685 6370 18692 6383
rect 18744 6411 18751 6422
rect 21080 6422 21146 6423
rect 21080 6411 21087 6422
rect 18744 6383 21087 6411
rect 18744 6370 18751 6383
rect 21080 6370 21087 6383
rect 21139 6411 21146 6422
rect 23376 6422 23442 6423
rect 23376 6411 23383 6422
rect 21139 6383 23383 6411
rect 21139 6370 21146 6383
rect 23376 6370 23383 6383
rect 23435 6370 23442 6422
rect 23545 6320 23609 6466
rect 23759 6320 23795 6466
rect 24329 6413 24395 6415
rect 24067 6408 24121 6412
rect 24066 6405 24121 6408
rect 23937 6371 24075 6405
rect 24109 6371 24121 6405
rect 24066 6368 24121 6371
rect 24066 6364 24120 6368
rect 24329 6361 24337 6413
rect 24389 6361 24395 6413
rect 24329 6360 24395 6361
rect 23545 6308 23795 6320
rect 10875 6280 23795 6308
rect 24423 6330 24451 6474
rect 24479 6417 24507 6549
rect 24535 6534 24541 6594
rect 24575 6534 24581 6594
rect 24535 6522 24581 6534
rect 24623 6594 24726 6606
rect 24623 6534 24629 6594
rect 24663 6534 24726 6594
rect 30476 6592 30495 6644
rect 30547 6592 30566 6644
rect 30476 6576 30566 6592
rect 24623 6522 24726 6534
rect 24573 6475 24642 6481
rect 24573 6441 24585 6475
rect 24619 6441 24642 6475
rect 24573 6435 24642 6441
rect 24479 6405 24528 6417
rect 24479 6371 24488 6405
rect 24522 6371 24528 6405
rect 24479 6358 24528 6371
rect 24423 6312 24566 6330
rect 24423 6302 24526 6312
rect 24517 6278 24526 6302
rect 24560 6278 24566 6312
rect 24517 6265 24566 6278
rect 10875 6251 23493 6252
rect 10753 6221 23493 6251
rect 10753 6187 11526 6221
rect 11560 6187 11618 6221
rect 11652 6187 11710 6221
rect 11744 6187 11802 6221
rect 11836 6187 11894 6221
rect 11928 6187 11986 6221
rect 12020 6187 12078 6221
rect 12112 6187 12170 6221
rect 12204 6187 12262 6221
rect 12296 6187 12354 6221
rect 12388 6187 12446 6221
rect 12480 6187 12538 6221
rect 12572 6187 12630 6221
rect 12664 6187 12722 6221
rect 12756 6187 12814 6221
rect 12848 6187 12906 6221
rect 12940 6187 12998 6221
rect 13032 6187 13090 6221
rect 13124 6187 13182 6221
rect 13216 6187 13274 6221
rect 13308 6187 13366 6221
rect 13400 6187 13458 6221
rect 13492 6187 13550 6221
rect 13584 6187 13642 6221
rect 13676 6187 13734 6221
rect 13768 6187 13826 6221
rect 13860 6187 13918 6221
rect 13952 6187 14010 6221
rect 14044 6187 14102 6221
rect 14136 6187 14194 6221
rect 14228 6187 14286 6221
rect 14320 6187 14378 6221
rect 14412 6187 14470 6221
rect 14504 6187 14562 6221
rect 14596 6187 14654 6221
rect 14688 6187 14746 6221
rect 14780 6187 14838 6221
rect 14872 6187 14930 6221
rect 14964 6187 15022 6221
rect 15056 6187 15114 6221
rect 15148 6187 15206 6221
rect 15240 6187 15298 6221
rect 15332 6187 15390 6221
rect 15424 6187 15482 6221
rect 15516 6187 15574 6221
rect 15608 6187 15666 6221
rect 15700 6187 15758 6221
rect 15792 6187 15850 6221
rect 15884 6187 15942 6221
rect 15976 6187 16034 6221
rect 16068 6187 16126 6221
rect 16160 6187 16218 6221
rect 16252 6187 16310 6221
rect 16344 6187 16402 6221
rect 16436 6187 16494 6221
rect 16528 6187 16586 6221
rect 16620 6187 16678 6221
rect 16712 6187 16770 6221
rect 16804 6187 16862 6221
rect 16896 6187 16954 6221
rect 16988 6187 17046 6221
rect 17080 6187 17138 6221
rect 17172 6187 17230 6221
rect 17264 6187 17322 6221
rect 17356 6187 17414 6221
rect 17448 6187 17506 6221
rect 17540 6187 17598 6221
rect 17632 6187 17690 6221
rect 17724 6187 17782 6221
rect 17816 6187 17874 6221
rect 17908 6187 17966 6221
rect 18000 6187 18058 6221
rect 18092 6187 18150 6221
rect 18184 6187 18242 6221
rect 18276 6187 18334 6221
rect 18368 6187 18426 6221
rect 18460 6187 18518 6221
rect 18552 6187 18610 6221
rect 18644 6187 18702 6221
rect 18736 6187 18794 6221
rect 18828 6187 18886 6221
rect 18920 6187 18978 6221
rect 19012 6187 19070 6221
rect 19104 6187 19162 6221
rect 19196 6187 19254 6221
rect 19288 6187 19346 6221
rect 19380 6187 19438 6221
rect 19472 6187 19530 6221
rect 19564 6187 19622 6221
rect 19656 6187 19714 6221
rect 19748 6187 19806 6221
rect 19840 6187 19898 6221
rect 19932 6187 19990 6221
rect 20024 6187 20082 6221
rect 20116 6187 20174 6221
rect 20208 6187 20266 6221
rect 20300 6187 20358 6221
rect 20392 6187 20450 6221
rect 20484 6187 20542 6221
rect 20576 6187 20634 6221
rect 20668 6187 20726 6221
rect 20760 6187 20818 6221
rect 20852 6187 20910 6221
rect 20944 6187 21002 6221
rect 21036 6187 21094 6221
rect 21128 6187 21186 6221
rect 21220 6187 21278 6221
rect 21312 6187 21370 6221
rect 21404 6187 21462 6221
rect 21496 6187 21554 6221
rect 21588 6187 21646 6221
rect 21680 6187 21738 6221
rect 21772 6187 21830 6221
rect 21864 6187 21922 6221
rect 21956 6187 22014 6221
rect 22048 6187 22106 6221
rect 22140 6187 22198 6221
rect 22232 6187 22290 6221
rect 22324 6187 22382 6221
rect 22416 6187 22474 6221
rect 22508 6187 22566 6221
rect 22600 6187 22658 6221
rect 22692 6187 22750 6221
rect 22784 6187 22842 6221
rect 22876 6187 22934 6221
rect 22968 6187 23026 6221
rect 23060 6187 23118 6221
rect 23152 6187 23210 6221
rect 23244 6187 23302 6221
rect 23336 6187 23394 6221
rect 23428 6199 23493 6221
rect 23428 6187 23494 6199
rect 10753 6156 23494 6187
rect 23999 6178 24459 6200
rect 23999 6169 24082 6178
rect 24134 6169 24202 6178
rect 24254 6169 24345 6178
rect 24397 6169 24459 6178
rect 10753 6132 11429 6156
rect 23999 6135 24028 6169
rect 24062 6135 24082 6169
rect 24154 6135 24202 6169
rect 24254 6135 24304 6169
rect 24338 6135 24345 6169
rect 24430 6135 24459 6169
rect 10753 6120 11261 6132
rect 10753 5974 10955 6120
rect 11105 5986 11261 6120
rect 11411 5986 11429 6132
rect 23020 6121 23052 6122
rect 23020 6117 23101 6121
rect 23020 6065 23026 6117
rect 23078 6107 23101 6117
rect 23381 6107 23440 6113
rect 23078 6073 23394 6107
rect 23428 6073 23440 6107
rect 23078 6072 23440 6073
rect 23078 6065 23101 6072
rect 23381 6066 23440 6072
rect 11607 6051 11665 6057
rect 11607 6017 11619 6051
rect 11653 6048 11665 6051
rect 11975 6051 12033 6057
rect 11975 6048 11987 6051
rect 11653 6020 11987 6048
rect 11653 6017 11665 6020
rect 11607 6011 11665 6017
rect 11975 6017 11987 6020
rect 12021 6048 12033 6051
rect 12711 6051 12769 6057
rect 12711 6048 12723 6051
rect 12021 6020 12723 6048
rect 12021 6017 12033 6020
rect 11975 6011 12033 6017
rect 12711 6017 12723 6020
rect 12757 6017 12769 6051
rect 12711 6011 12769 6017
rect 13999 6051 14057 6057
rect 13999 6017 14011 6051
rect 14045 6048 14057 6051
rect 14367 6051 14425 6057
rect 14367 6048 14379 6051
rect 14045 6020 14379 6048
rect 14045 6017 14057 6020
rect 13999 6011 14057 6017
rect 14367 6017 14379 6020
rect 14413 6048 14425 6051
rect 15103 6051 15161 6057
rect 15103 6048 15115 6051
rect 14413 6020 15115 6048
rect 14413 6017 14425 6020
rect 14367 6011 14425 6017
rect 15103 6017 15115 6020
rect 15149 6017 15161 6051
rect 15103 6011 15161 6017
rect 16391 6051 16449 6057
rect 16391 6017 16403 6051
rect 16437 6048 16449 6051
rect 16759 6051 16817 6057
rect 16759 6048 16771 6051
rect 16437 6020 16771 6048
rect 16437 6017 16449 6020
rect 16391 6011 16449 6017
rect 16759 6017 16771 6020
rect 16805 6048 16817 6051
rect 17495 6051 17553 6057
rect 17495 6048 17507 6051
rect 16805 6020 17507 6048
rect 16805 6017 16817 6020
rect 16759 6011 16817 6017
rect 17495 6017 17507 6020
rect 17541 6017 17553 6051
rect 17495 6011 17553 6017
rect 18783 6051 18841 6057
rect 18783 6017 18795 6051
rect 18829 6048 18841 6051
rect 19151 6051 19209 6057
rect 19151 6048 19163 6051
rect 18829 6020 19163 6048
rect 18829 6017 18841 6020
rect 18783 6011 18841 6017
rect 19151 6017 19163 6020
rect 19197 6048 19209 6051
rect 19887 6051 19945 6057
rect 19887 6048 19899 6051
rect 19197 6020 19899 6048
rect 19197 6017 19209 6020
rect 19151 6011 19209 6017
rect 19887 6017 19899 6020
rect 19933 6017 19945 6051
rect 19887 6011 19945 6017
rect 21175 6051 21233 6057
rect 21175 6017 21187 6051
rect 21221 6048 21233 6051
rect 21543 6051 21601 6057
rect 21543 6048 21555 6051
rect 21221 6020 21555 6048
rect 21221 6017 21233 6020
rect 21175 6011 21233 6017
rect 21543 6017 21555 6020
rect 21589 6048 21601 6051
rect 22279 6051 22337 6057
rect 23020 6056 23101 6065
rect 23020 6055 23052 6056
rect 22279 6048 22291 6051
rect 21589 6020 22291 6048
rect 21589 6017 21601 6020
rect 21543 6011 21601 6017
rect 22279 6017 22291 6020
rect 22325 6017 22337 6051
rect 22279 6011 22337 6017
rect 23531 6040 23795 6132
rect 23999 6126 24082 6135
rect 24134 6126 24202 6135
rect 24254 6126 24345 6135
rect 24397 6126 24459 6135
rect 23999 6104 24459 6126
rect 11105 5974 11429 5986
rect 10753 5864 11429 5974
rect 11874 5980 11937 5987
rect 12478 5980 12485 5992
rect 11874 5946 11891 5980
rect 11925 5952 12485 5980
rect 11925 5946 11937 5952
rect 11874 5940 11937 5946
rect 12478 5940 12485 5952
rect 12537 5940 12544 5992
rect 12619 5983 12677 5989
rect 12619 5949 12631 5983
rect 12665 5980 12677 5983
rect 13263 5983 13321 5989
rect 13263 5980 13275 5983
rect 12665 5952 13275 5980
rect 12665 5949 12677 5952
rect 12619 5943 12677 5949
rect 13263 5949 13275 5952
rect 13309 5949 13321 5983
rect 13263 5943 13321 5949
rect 13819 5987 13878 5993
rect 13819 5953 13831 5987
rect 13865 5983 13878 5987
rect 14230 5983 14289 5989
rect 13865 5955 14242 5983
rect 13865 5953 13878 5955
rect 13819 5946 13878 5953
rect 14230 5949 14242 5955
rect 14276 5949 14289 5983
rect 14230 5942 14289 5949
rect 15011 5983 15069 5989
rect 15011 5949 15023 5983
rect 15057 5980 15069 5983
rect 15655 5983 15713 5989
rect 15655 5980 15667 5983
rect 15057 5952 15667 5980
rect 15057 5949 15069 5952
rect 15011 5943 15069 5949
rect 15655 5949 15667 5952
rect 15701 5949 15713 5983
rect 15655 5943 15713 5949
rect 16208 5986 16267 5992
rect 16208 5952 16220 5986
rect 16254 5982 16267 5986
rect 16619 5982 16678 5988
rect 16254 5954 16631 5982
rect 16254 5952 16267 5954
rect 16208 5945 16267 5952
rect 16619 5948 16631 5954
rect 16665 5948 16678 5982
rect 16619 5941 16678 5948
rect 17403 5983 17461 5989
rect 17403 5949 17415 5983
rect 17449 5980 17461 5983
rect 18047 5983 18105 5989
rect 18047 5980 18059 5983
rect 17449 5952 18059 5980
rect 17449 5949 17461 5952
rect 17403 5943 17461 5949
rect 18047 5949 18059 5952
rect 18093 5949 18105 5983
rect 18047 5943 18105 5949
rect 18603 5984 18662 5990
rect 18603 5950 18615 5984
rect 18649 5980 18662 5984
rect 19014 5980 19073 5986
rect 18649 5952 19026 5980
rect 18649 5950 18662 5952
rect 18603 5943 18662 5950
rect 19014 5946 19026 5952
rect 19060 5946 19073 5980
rect 19014 5939 19073 5946
rect 19795 5983 19853 5989
rect 19795 5949 19807 5983
rect 19841 5980 19853 5983
rect 20439 5983 20497 5989
rect 20439 5980 20451 5983
rect 19841 5952 20451 5980
rect 19841 5949 19853 5952
rect 19795 5943 19853 5949
rect 20439 5949 20451 5952
rect 20485 5949 20497 5983
rect 20439 5943 20497 5949
rect 20994 5983 21053 5989
rect 20994 5949 21006 5983
rect 21040 5979 21053 5983
rect 21405 5979 21464 5985
rect 21040 5951 21417 5979
rect 21040 5949 21053 5951
rect 20994 5942 21053 5949
rect 21405 5945 21417 5951
rect 21451 5945 21464 5979
rect 21405 5938 21464 5945
rect 22187 5983 22245 5989
rect 22187 5949 22199 5983
rect 22233 5980 22245 5983
rect 22831 5983 22889 5989
rect 22831 5980 22843 5983
rect 22233 5952 22843 5980
rect 22233 5949 22245 5952
rect 22187 5943 22245 5949
rect 22831 5949 22843 5952
rect 22877 5949 22889 5983
rect 22831 5943 22889 5949
rect 12711 5915 12769 5921
rect 12711 5912 12723 5915
rect 11515 5909 11581 5910
rect 11515 5857 11522 5909
rect 11574 5857 11581 5909
rect 12082 5884 12723 5912
rect 12082 5853 12121 5884
rect 12711 5881 12723 5884
rect 12757 5881 12769 5915
rect 15103 5915 15161 5921
rect 15103 5912 15115 5915
rect 12711 5875 12769 5881
rect 13905 5909 13971 5910
rect 13905 5857 13912 5909
rect 13964 5857 13971 5909
rect 14474 5884 15115 5912
rect 12983 5854 13049 5855
rect 11699 5847 11757 5853
rect 11699 5813 11711 5847
rect 11745 5844 11757 5847
rect 12063 5847 12121 5853
rect 12063 5844 12075 5847
rect 11745 5816 12075 5844
rect 11745 5813 11757 5816
rect 11699 5807 11757 5813
rect 12063 5813 12075 5816
rect 12109 5813 12121 5847
rect 12063 5807 12121 5813
rect 12251 5847 12309 5853
rect 12251 5813 12263 5847
rect 12297 5844 12309 5847
rect 12983 5844 12990 5854
rect 12297 5816 12990 5844
rect 12297 5813 12309 5816
rect 12251 5807 12309 5813
rect 12983 5802 12990 5816
rect 13042 5802 13049 5854
rect 14474 5853 14513 5884
rect 15103 5881 15115 5884
rect 15149 5881 15161 5915
rect 15103 5875 15161 5881
rect 15749 5876 15756 5928
rect 15808 5876 15814 5928
rect 18149 5927 18202 5934
rect 17495 5915 17553 5921
rect 17495 5912 17507 5915
rect 16298 5910 16364 5911
rect 16298 5858 16305 5910
rect 16357 5858 16364 5910
rect 16866 5884 17507 5912
rect 16866 5853 16905 5884
rect 17495 5881 17507 5884
rect 17541 5881 17553 5915
rect 17495 5875 17553 5881
rect 18201 5875 18202 5927
rect 20540 5929 20593 5936
rect 19887 5915 19945 5921
rect 19887 5912 19899 5915
rect 18149 5868 18202 5875
rect 18690 5909 18756 5910
rect 18690 5857 18697 5909
rect 18749 5857 18756 5909
rect 19258 5884 19899 5912
rect 19258 5853 19297 5884
rect 19887 5881 19899 5884
rect 19933 5881 19945 5915
rect 19887 5875 19945 5881
rect 20592 5877 20593 5929
rect 22931 5927 22984 5934
rect 22279 5915 22337 5921
rect 22279 5912 22291 5915
rect 20540 5870 20593 5877
rect 21085 5911 21151 5912
rect 21085 5859 21092 5911
rect 21144 5859 21151 5911
rect 21650 5884 22291 5912
rect 21650 5853 21689 5884
rect 22279 5881 22291 5884
rect 22325 5881 22337 5915
rect 22279 5875 22337 5881
rect 22983 5875 22984 5927
rect 22931 5868 22984 5875
rect 23531 5894 23609 6040
rect 23759 5894 23795 6040
rect 23914 5985 23921 6037
rect 23973 6035 23979 6037
rect 24594 6035 24642 6435
rect 23973 5988 24642 6035
rect 23973 5985 23979 5988
rect 23914 5984 23979 5985
rect 14091 5847 14149 5853
rect 14091 5813 14103 5847
rect 14137 5844 14149 5847
rect 14455 5847 14513 5853
rect 14455 5844 14467 5847
rect 14137 5816 14467 5844
rect 14137 5813 14149 5816
rect 14091 5807 14149 5813
rect 14455 5813 14467 5816
rect 14501 5813 14513 5847
rect 14455 5807 14513 5813
rect 14643 5847 14701 5853
rect 14643 5813 14655 5847
rect 14689 5844 14701 5847
rect 15379 5847 15437 5853
rect 15379 5844 15391 5847
rect 14689 5816 15391 5844
rect 14689 5813 14701 5816
rect 14643 5807 14701 5813
rect 15379 5813 15391 5816
rect 15425 5813 15437 5847
rect 16483 5847 16541 5853
rect 16039 5821 16092 5828
rect 15379 5807 15437 5813
rect 15923 5810 15987 5816
rect 13533 5796 13599 5797
rect 13533 5744 13540 5796
rect 13592 5744 13599 5796
rect 15923 5758 15930 5810
rect 15982 5758 15987 5810
rect 16039 5769 16040 5821
rect 16200 5817 16261 5821
rect 16199 5812 16261 5817
rect 16092 5778 16211 5812
rect 16245 5778 16261 5812
rect 16483 5813 16495 5847
rect 16529 5844 16541 5847
rect 16847 5847 16905 5853
rect 16847 5844 16859 5847
rect 16529 5816 16859 5844
rect 16529 5813 16541 5816
rect 16483 5807 16541 5813
rect 16847 5813 16859 5816
rect 16893 5813 16905 5847
rect 16847 5807 16905 5813
rect 17035 5847 17093 5853
rect 17035 5813 17047 5847
rect 17081 5844 17093 5847
rect 17771 5847 17829 5853
rect 17771 5844 17783 5847
rect 17081 5816 17783 5844
rect 17081 5813 17093 5816
rect 17035 5807 17093 5813
rect 17771 5813 17783 5816
rect 17817 5813 17829 5847
rect 18875 5847 18933 5853
rect 17771 5807 17829 5813
rect 16199 5773 16261 5778
rect 16200 5770 16261 5773
rect 16039 5762 16092 5769
rect 18313 5766 18319 5818
rect 18371 5766 18377 5818
rect 18313 5758 18377 5766
rect 18435 5810 18488 5817
rect 18875 5813 18887 5847
rect 18921 5844 18933 5847
rect 19239 5847 19297 5853
rect 19239 5844 19251 5847
rect 18921 5816 19251 5844
rect 18921 5813 18933 5816
rect 18435 5758 18436 5810
rect 18598 5806 18659 5811
rect 18875 5807 18933 5813
rect 19239 5813 19251 5816
rect 19285 5813 19297 5847
rect 19239 5807 19297 5813
rect 19427 5847 19485 5853
rect 19427 5813 19439 5847
rect 19473 5844 19485 5847
rect 20163 5847 20221 5853
rect 20163 5844 20175 5847
rect 19473 5816 20175 5844
rect 19473 5813 19485 5816
rect 19427 5807 19485 5813
rect 20163 5813 20175 5816
rect 20209 5813 20221 5847
rect 21267 5847 21325 5853
rect 20163 5807 20221 5813
rect 20835 5826 20888 5833
rect 18595 5801 18659 5806
rect 18488 5767 18607 5801
rect 18641 5767 18659 5801
rect 18595 5762 18659 5767
rect 18598 5760 18659 5762
rect 20715 5795 20768 5802
rect 15923 5757 15987 5758
rect 15923 5752 15986 5757
rect 18435 5751 18488 5758
rect 20767 5743 20768 5795
rect 20835 5774 20836 5826
rect 20995 5817 21056 5826
rect 20888 5783 21007 5817
rect 21041 5783 21056 5817
rect 21267 5813 21279 5847
rect 21313 5844 21325 5847
rect 21631 5847 21689 5853
rect 21631 5844 21643 5847
rect 21313 5816 21643 5844
rect 21313 5813 21325 5816
rect 21267 5807 21325 5813
rect 21631 5813 21643 5816
rect 21677 5813 21689 5847
rect 21631 5807 21689 5813
rect 21819 5847 21877 5853
rect 21819 5813 21831 5847
rect 21865 5844 21877 5847
rect 22555 5847 22613 5853
rect 22555 5844 22567 5847
rect 21865 5816 22567 5844
rect 21865 5813 21877 5816
rect 21819 5807 21877 5813
rect 22555 5813 22567 5816
rect 22601 5813 22613 5847
rect 22555 5807 22613 5813
rect 23230 5826 23283 5833
rect 20995 5775 21056 5783
rect 23106 5796 23159 5803
rect 20835 5767 20888 5774
rect 20715 5736 20768 5743
rect 23158 5744 23159 5796
rect 23230 5774 23231 5826
rect 23389 5817 23450 5826
rect 23283 5783 23402 5817
rect 23436 5783 23450 5817
rect 23389 5775 23450 5783
rect 23531 5814 23795 5894
rect 24594 5847 24642 5988
rect 24584 5841 24642 5847
rect 24343 5835 24408 5836
rect 24343 5834 24349 5835
rect 23230 5767 23283 5774
rect 23106 5737 23159 5744
rect 10871 5701 23490 5708
rect 23531 5701 23609 5814
rect 10871 5677 23609 5701
rect 10871 5643 11526 5677
rect 11560 5643 11618 5677
rect 11652 5643 11710 5677
rect 11744 5643 11802 5677
rect 11836 5643 11894 5677
rect 11928 5643 11986 5677
rect 12020 5643 12078 5677
rect 12112 5643 12170 5677
rect 12204 5643 12262 5677
rect 12296 5643 12354 5677
rect 12388 5643 12446 5677
rect 12480 5643 12538 5677
rect 12572 5643 12630 5677
rect 12664 5643 12722 5677
rect 12756 5643 12814 5677
rect 12848 5643 12906 5677
rect 12940 5643 12998 5677
rect 13032 5643 13090 5677
rect 13124 5643 13182 5677
rect 13216 5643 13274 5677
rect 13308 5643 13366 5677
rect 13400 5643 13458 5677
rect 13492 5643 13550 5677
rect 13584 5643 13642 5677
rect 13676 5643 13734 5677
rect 13768 5643 13826 5677
rect 13860 5643 13918 5677
rect 13952 5643 14010 5677
rect 14044 5643 14102 5677
rect 14136 5643 14194 5677
rect 14228 5643 14286 5677
rect 14320 5643 14378 5677
rect 14412 5643 14470 5677
rect 14504 5643 14562 5677
rect 14596 5643 14654 5677
rect 14688 5643 14746 5677
rect 14780 5643 14838 5677
rect 14872 5643 14930 5677
rect 14964 5643 15022 5677
rect 15056 5643 15114 5677
rect 15148 5643 15206 5677
rect 15240 5643 15298 5677
rect 15332 5643 15390 5677
rect 15424 5643 15482 5677
rect 15516 5643 15574 5677
rect 15608 5643 15666 5677
rect 15700 5643 15758 5677
rect 15792 5643 15850 5677
rect 15884 5643 15942 5677
rect 15976 5643 16034 5677
rect 16068 5643 16126 5677
rect 16160 5643 16218 5677
rect 16252 5643 16310 5677
rect 16344 5643 16402 5677
rect 16436 5643 16494 5677
rect 16528 5643 16586 5677
rect 16620 5643 16678 5677
rect 16712 5643 16770 5677
rect 16804 5643 16862 5677
rect 16896 5643 16954 5677
rect 16988 5643 17046 5677
rect 17080 5643 17138 5677
rect 17172 5643 17230 5677
rect 17264 5643 17322 5677
rect 17356 5643 17414 5677
rect 17448 5643 17506 5677
rect 17540 5643 17598 5677
rect 17632 5643 17690 5677
rect 17724 5643 17782 5677
rect 17816 5643 17874 5677
rect 17908 5643 17966 5677
rect 18000 5643 18058 5677
rect 18092 5643 18150 5677
rect 18184 5643 18242 5677
rect 18276 5643 18334 5677
rect 18368 5643 18426 5677
rect 18460 5643 18518 5677
rect 18552 5643 18610 5677
rect 18644 5643 18702 5677
rect 18736 5643 18794 5677
rect 18828 5643 18886 5677
rect 18920 5643 18978 5677
rect 19012 5643 19070 5677
rect 19104 5643 19162 5677
rect 19196 5643 19254 5677
rect 19288 5643 19346 5677
rect 19380 5643 19438 5677
rect 19472 5643 19530 5677
rect 19564 5643 19622 5677
rect 19656 5643 19714 5677
rect 19748 5643 19806 5677
rect 19840 5643 19898 5677
rect 19932 5643 19990 5677
rect 20024 5643 20082 5677
rect 20116 5643 20174 5677
rect 20208 5643 20266 5677
rect 20300 5643 20358 5677
rect 20392 5643 20450 5677
rect 20484 5643 20542 5677
rect 20576 5643 20634 5677
rect 20668 5643 20726 5677
rect 20760 5643 20818 5677
rect 20852 5643 20910 5677
rect 20944 5643 21002 5677
rect 21036 5643 21094 5677
rect 21128 5643 21186 5677
rect 21220 5643 21278 5677
rect 21312 5643 21370 5677
rect 21404 5643 21462 5677
rect 21496 5643 21554 5677
rect 21588 5643 21646 5677
rect 21680 5643 21738 5677
rect 21772 5643 21830 5677
rect 21864 5643 21922 5677
rect 21956 5643 22014 5677
rect 22048 5643 22106 5677
rect 22140 5643 22198 5677
rect 22232 5643 22290 5677
rect 22324 5643 22382 5677
rect 22416 5643 22474 5677
rect 22508 5643 22566 5677
rect 22600 5643 22658 5677
rect 22692 5643 22750 5677
rect 22784 5643 22842 5677
rect 22876 5643 22934 5677
rect 22968 5643 23026 5677
rect 23060 5643 23118 5677
rect 23152 5643 23210 5677
rect 23244 5643 23302 5677
rect 23336 5643 23394 5677
rect 23428 5668 23609 5677
rect 23759 5668 23795 5814
rect 24237 5786 24349 5834
rect 24343 5783 24349 5786
rect 24401 5783 24408 5835
rect 24584 5807 24596 5841
rect 24630 5807 24642 5841
rect 24584 5801 24642 5807
rect 24680 6032 24726 6522
rect 30394 6402 30484 6418
rect 30394 6391 30413 6402
rect 30319 6350 30413 6391
rect 30465 6350 30484 6402
rect 30771 6410 30861 6426
rect 30771 6399 30790 6410
rect 30752 6367 30790 6399
rect 24776 6335 24825 6342
rect 24776 6330 25395 6335
rect 24776 6296 24785 6330
rect 24819 6296 25395 6330
rect 24776 6288 25395 6296
rect 24776 6283 24825 6288
rect 24777 6241 24826 6249
rect 25346 6241 25395 6288
rect 30319 6332 30484 6350
rect 30679 6358 30790 6367
rect 30842 6367 30861 6410
rect 30971 6410 31061 6426
rect 30971 6399 30990 6410
rect 30952 6367 30990 6399
rect 30842 6358 30990 6367
rect 31042 6358 31061 6410
rect 30679 6340 31061 6358
rect 30679 6336 31047 6340
rect 30319 6286 30366 6332
rect 30679 6302 30708 6336
rect 30742 6302 30800 6336
rect 30834 6302 30892 6336
rect 30926 6302 30984 6336
rect 31018 6302 31047 6336
rect 30320 6283 30366 6286
rect 24777 6237 25278 6241
rect 24777 6203 24786 6237
rect 24820 6232 25278 6237
rect 24820 6203 25227 6232
rect 24777 6198 25227 6203
rect 25261 6198 25278 6232
rect 24777 6195 25278 6198
rect 25346 6235 29767 6241
rect 25346 6201 25959 6235
rect 25993 6201 26085 6235
rect 26119 6201 27171 6235
rect 27205 6201 27297 6235
rect 27331 6201 28383 6235
rect 28417 6201 28509 6235
rect 28543 6201 29595 6235
rect 29629 6201 29721 6235
rect 29755 6201 29767 6235
rect 30320 6223 30326 6283
rect 30360 6223 30366 6283
rect 30320 6211 30366 6223
rect 30408 6283 30454 6295
rect 30408 6223 30414 6283
rect 30448 6223 30454 6283
rect 30679 6271 31047 6302
rect 30408 6214 30454 6223
rect 25346 6195 29767 6201
rect 24777 6194 25273 6195
rect 25346 6194 25792 6195
rect 24777 6190 24826 6194
rect 25215 6192 25273 6194
rect 30408 6185 30646 6214
rect 25177 6143 25223 6151
rect 25154 6142 25233 6143
rect 25154 6078 25161 6142
rect 25225 6078 25233 6142
rect 25265 6142 25311 6154
rect 25909 6146 25955 6154
rect 25265 6082 25271 6142
rect 25305 6082 25311 6142
rect 25177 6067 25223 6078
rect 25265 6032 25311 6082
rect 25886 6145 25965 6146
rect 25886 6081 25893 6145
rect 25957 6081 25965 6145
rect 26014 6142 26060 6154
rect 26123 6146 26169 6154
rect 27121 6146 27167 6154
rect 26014 6082 26020 6142
rect 26054 6082 26060 6142
rect 25909 6070 25955 6081
rect 26014 6032 26060 6082
rect 26113 6145 26192 6146
rect 26113 6081 26121 6145
rect 26185 6081 26192 6145
rect 27098 6145 27177 6146
rect 27098 6081 27105 6145
rect 27169 6081 27177 6145
rect 27225 6142 27271 6154
rect 27335 6146 27381 6154
rect 28333 6146 28379 6154
rect 27225 6082 27231 6142
rect 27265 6082 27271 6142
rect 26123 6070 26169 6081
rect 27121 6070 27167 6081
rect 27225 6032 27271 6082
rect 27325 6145 27404 6146
rect 27325 6081 27333 6145
rect 27397 6081 27404 6145
rect 28310 6145 28389 6146
rect 28310 6081 28317 6145
rect 28381 6081 28389 6145
rect 28438 6142 28484 6154
rect 28547 6146 28593 6154
rect 29545 6146 29591 6154
rect 28438 6082 28444 6142
rect 28478 6082 28484 6142
rect 27335 6070 27381 6081
rect 28333 6070 28379 6081
rect 28438 6032 28484 6082
rect 28537 6145 28616 6146
rect 28537 6081 28545 6145
rect 28609 6081 28616 6145
rect 29522 6145 29601 6146
rect 29522 6081 29529 6145
rect 29593 6081 29601 6145
rect 29652 6142 29698 6154
rect 29759 6146 29805 6154
rect 29652 6082 29658 6142
rect 29692 6082 29698 6142
rect 28547 6070 28593 6081
rect 29545 6070 29591 6081
rect 29652 6032 29698 6082
rect 29749 6145 29828 6146
rect 29749 6081 29757 6145
rect 29821 6081 29828 6145
rect 30320 6145 30366 6157
rect 30320 6085 30326 6145
rect 30360 6085 30366 6145
rect 29759 6070 29805 6081
rect 30320 6073 30366 6085
rect 30408 6145 30454 6185
rect 30408 6085 30414 6145
rect 30448 6085 30454 6145
rect 30408 6073 30454 6085
rect 30482 6145 30572 6157
rect 30482 6141 30510 6145
rect 30544 6141 30572 6145
rect 30482 6089 30501 6141
rect 30553 6089 30572 6141
rect 30482 6085 30510 6089
rect 30544 6085 30572 6089
rect 30482 6073 30572 6085
rect 30600 6145 30646 6185
rect 30600 6085 30606 6145
rect 30640 6085 30646 6145
rect 30600 6073 30646 6085
rect 30239 6032 30305 6034
rect 24680 6028 30305 6032
rect 24680 5994 30255 6028
rect 30289 5994 30305 6028
rect 24680 5990 30305 5994
rect 24680 5769 24726 5990
rect 25530 5943 25576 5953
rect 25508 5879 25517 5943
rect 25581 5879 25590 5943
rect 25508 5878 25590 5879
rect 25620 5941 25666 5990
rect 26262 5943 26308 5953
rect 25620 5881 25626 5941
rect 25660 5881 25666 5941
rect 25530 5869 25576 5878
rect 25620 5869 25666 5881
rect 26240 5879 26249 5943
rect 26313 5879 26322 5943
rect 26240 5878 26322 5879
rect 26369 5941 26415 5990
rect 26472 5943 26518 5953
rect 27474 5943 27520 5953
rect 26369 5881 26375 5941
rect 26409 5881 26415 5941
rect 26262 5869 26308 5878
rect 26369 5869 26415 5881
rect 26458 5879 26467 5943
rect 26531 5879 26540 5943
rect 26458 5878 26540 5879
rect 27452 5879 27461 5943
rect 27525 5879 27534 5943
rect 27452 5878 27534 5879
rect 27580 5941 27626 5990
rect 27684 5943 27730 5953
rect 28812 5943 28858 5953
rect 27580 5881 27586 5941
rect 27620 5881 27626 5941
rect 26472 5869 26518 5878
rect 27474 5869 27520 5878
rect 27580 5869 27626 5881
rect 27670 5879 27679 5943
rect 27743 5879 27752 5943
rect 27670 5878 27752 5879
rect 28790 5879 28799 5943
rect 28863 5879 28872 5943
rect 28790 5878 28872 5879
rect 28920 5941 28966 5990
rect 29022 5943 29068 5953
rect 28920 5881 28926 5941
rect 28960 5881 28966 5941
rect 27684 5869 27730 5878
rect 28812 5869 28858 5878
rect 28920 5869 28966 5881
rect 29008 5879 29017 5943
rect 29081 5879 29090 5943
rect 29008 5878 29090 5879
rect 29667 5941 29713 5990
rect 30243 5988 30305 5990
rect 30338 6025 30366 6073
rect 30450 6026 30749 6032
rect 30450 6025 30462 6026
rect 30338 5996 30462 6025
rect 30338 5954 30366 5996
rect 30450 5992 30462 5996
rect 30496 5992 30702 6026
rect 30736 5992 30749 6026
rect 30450 5986 30749 5992
rect 30897 6026 30955 6032
rect 30897 5992 30909 6026
rect 30943 6023 30955 6026
rect 30943 5995 31104 6023
rect 30943 5992 30955 5995
rect 30897 5986 30955 5992
rect 29756 5943 29802 5953
rect 29667 5881 29673 5941
rect 29707 5881 29713 5941
rect 29022 5869 29068 5878
rect 29667 5869 29713 5881
rect 29742 5879 29751 5943
rect 29815 5879 29824 5943
rect 29742 5878 29824 5879
rect 30320 5942 30366 5954
rect 30320 5882 30326 5942
rect 30360 5882 30366 5942
rect 29756 5869 29802 5878
rect 30320 5870 30366 5882
rect 30408 5942 30454 5954
rect 30408 5882 30414 5942
rect 30448 5882 30454 5942
rect 30408 5842 30454 5882
rect 30482 5942 30572 5954
rect 30482 5938 30510 5942
rect 30544 5938 30572 5942
rect 30482 5886 30501 5938
rect 30553 5886 30572 5938
rect 30482 5882 30510 5886
rect 30544 5882 30572 5886
rect 30482 5870 30572 5882
rect 30600 5942 30646 5954
rect 30600 5882 30606 5942
rect 30640 5882 30646 5942
rect 30600 5842 30646 5882
rect 29708 5837 29767 5840
rect 24830 5783 24837 5835
rect 24889 5833 24895 5835
rect 25568 5833 25626 5837
rect 24889 5831 25626 5833
rect 24889 5797 25580 5831
rect 25614 5816 25626 5831
rect 26300 5831 27696 5837
rect 25614 5797 25628 5816
rect 24889 5786 25628 5797
rect 26300 5797 26312 5831
rect 26346 5797 26434 5831
rect 26468 5797 27524 5831
rect 27558 5797 27646 5831
rect 27680 5797 27696 5831
rect 26300 5791 27696 5797
rect 28850 5831 29034 5837
rect 28850 5797 28862 5831
rect 28896 5797 28984 5831
rect 29018 5797 29034 5831
rect 28850 5791 29034 5797
rect 29706 5831 29767 5837
rect 29706 5797 29718 5831
rect 29752 5797 29767 5831
rect 29706 5791 29767 5797
rect 24889 5783 24895 5786
rect 24830 5782 24895 5783
rect 25570 5781 25628 5786
rect 23428 5643 23795 5668
rect 10871 5625 23795 5643
rect 24510 5757 24556 5769
rect 24510 5697 24516 5757
rect 24550 5697 24556 5757
rect 10871 5612 23490 5625
rect 24510 5619 24556 5697
rect 24670 5757 24726 5769
rect 24670 5697 24676 5757
rect 24710 5697 24726 5757
rect 24670 5685 24726 5697
rect 10871 5556 23490 5563
rect 10753 5532 23490 5556
rect 24510 5559 24516 5619
rect 24550 5559 24556 5619
rect 24510 5547 24556 5559
rect 24670 5619 24716 5631
rect 24670 5559 24676 5619
rect 24710 5559 24716 5619
rect 10753 5498 11086 5532
rect 11120 5498 11178 5532
rect 11212 5498 11270 5532
rect 11304 5498 11362 5532
rect 11396 5498 11454 5532
rect 11488 5498 11546 5532
rect 11580 5498 11638 5532
rect 11672 5498 11730 5532
rect 11764 5498 11822 5532
rect 11856 5498 11894 5532
rect 11928 5498 11986 5532
rect 12020 5498 12078 5532
rect 12112 5498 12170 5532
rect 12204 5498 12262 5532
rect 12296 5498 12354 5532
rect 12388 5498 12446 5532
rect 12480 5498 12538 5532
rect 12572 5498 12630 5532
rect 12664 5498 12722 5532
rect 12756 5498 12814 5532
rect 12848 5498 12906 5532
rect 12940 5498 12998 5532
rect 13032 5498 13090 5532
rect 13124 5498 13182 5532
rect 13216 5498 13274 5532
rect 13308 5498 13366 5532
rect 13400 5498 13458 5532
rect 13492 5498 13550 5532
rect 13584 5498 13642 5532
rect 13676 5498 13734 5532
rect 13768 5498 13826 5532
rect 13860 5498 13918 5532
rect 13952 5498 14010 5532
rect 14044 5498 14102 5532
rect 14136 5498 14194 5532
rect 14228 5498 14286 5532
rect 14320 5498 14378 5532
rect 14412 5498 14470 5532
rect 14504 5498 14562 5532
rect 14596 5498 14654 5532
rect 14688 5498 14746 5532
rect 14780 5498 14838 5532
rect 14872 5498 14930 5532
rect 14964 5498 15022 5532
rect 15056 5498 15114 5532
rect 15148 5498 15206 5532
rect 15240 5498 15298 5532
rect 15332 5498 15390 5532
rect 15424 5498 15482 5532
rect 15516 5498 15574 5532
rect 15608 5498 15666 5532
rect 15700 5498 15758 5532
rect 15792 5498 15850 5532
rect 15884 5498 15942 5532
rect 15976 5498 16034 5532
rect 16068 5498 16126 5532
rect 16160 5498 16218 5532
rect 16252 5498 16310 5532
rect 16344 5498 16402 5532
rect 16436 5498 16494 5532
rect 16528 5498 16586 5532
rect 16620 5498 16678 5532
rect 16712 5498 16770 5532
rect 16804 5498 16862 5532
rect 16896 5498 16954 5532
rect 16988 5498 17046 5532
rect 17080 5498 17138 5532
rect 17172 5498 17230 5532
rect 17264 5498 17322 5532
rect 17356 5498 17414 5532
rect 17448 5498 17506 5532
rect 17540 5498 17598 5532
rect 17632 5498 17690 5532
rect 17724 5498 17782 5532
rect 17816 5498 17874 5532
rect 17908 5498 17966 5532
rect 18000 5498 18058 5532
rect 18092 5498 18150 5532
rect 18184 5498 18242 5532
rect 18276 5498 18334 5532
rect 18368 5498 18426 5532
rect 18460 5498 18518 5532
rect 18552 5498 18610 5532
rect 18644 5498 18702 5532
rect 18736 5498 18794 5532
rect 18828 5498 18886 5532
rect 18920 5498 18978 5532
rect 19012 5498 19070 5532
rect 19104 5498 19162 5532
rect 19196 5498 19254 5532
rect 19288 5498 19346 5532
rect 19380 5498 19438 5532
rect 19472 5498 19530 5532
rect 19564 5498 19622 5532
rect 19656 5498 19714 5532
rect 19748 5498 19806 5532
rect 19840 5498 19898 5532
rect 19932 5498 19990 5532
rect 20024 5498 20082 5532
rect 20116 5498 20174 5532
rect 20208 5498 20266 5532
rect 20300 5498 20358 5532
rect 20392 5498 20450 5532
rect 20484 5498 20542 5532
rect 20576 5498 20634 5532
rect 20668 5498 20726 5532
rect 20760 5498 20818 5532
rect 20852 5498 20910 5532
rect 20944 5498 21002 5532
rect 21036 5498 21094 5532
rect 21128 5498 21186 5532
rect 21220 5498 21278 5532
rect 21312 5498 21370 5532
rect 21404 5498 21462 5532
rect 21496 5498 21554 5532
rect 21588 5498 21646 5532
rect 21680 5498 21738 5532
rect 21772 5498 21830 5532
rect 21864 5498 21922 5532
rect 21956 5498 22014 5532
rect 22048 5498 22106 5532
rect 22140 5498 22198 5532
rect 22232 5498 22290 5532
rect 22324 5498 22382 5532
rect 22416 5498 22474 5532
rect 22508 5498 22566 5532
rect 22600 5498 22658 5532
rect 22692 5498 22750 5532
rect 22784 5498 22842 5532
rect 22876 5498 22934 5532
rect 22968 5498 23026 5532
rect 23060 5498 23118 5532
rect 23152 5498 23210 5532
rect 23244 5498 23302 5532
rect 23336 5498 23394 5532
rect 23428 5498 23490 5532
rect 10753 5492 23490 5498
rect 10753 5346 10787 5492
rect 10937 5467 23490 5492
rect 24510 5481 24556 5493
rect 10937 5346 10983 5467
rect 10753 5284 10983 5346
rect 12990 5404 13043 5411
rect 12990 5352 12991 5404
rect 13899 5386 13905 5438
rect 13957 5386 13963 5438
rect 24510 5421 24516 5481
rect 24550 5421 24556 5481
rect 16296 5420 16362 5421
rect 16296 5368 16303 5420
rect 16355 5405 16362 5420
rect 18687 5420 18753 5421
rect 16355 5368 16415 5405
rect 18687 5368 18694 5420
rect 18746 5405 18753 5420
rect 21081 5411 21134 5417
rect 18746 5368 18807 5405
rect 12990 5345 13043 5352
rect 15009 5362 15067 5368
rect 15009 5328 15021 5362
rect 15055 5359 15067 5362
rect 15745 5362 15803 5368
rect 15745 5359 15757 5362
rect 15055 5331 15757 5359
rect 15055 5328 15067 5331
rect 15009 5322 15067 5328
rect 15745 5328 15757 5331
rect 15791 5359 15803 5362
rect 16113 5362 16171 5368
rect 16113 5359 16125 5362
rect 15791 5331 16125 5359
rect 15791 5328 15803 5331
rect 15745 5322 15803 5328
rect 16113 5328 16125 5331
rect 16159 5328 16171 5362
rect 16113 5322 16171 5328
rect 16296 5303 16349 5310
rect 16296 5302 16297 5303
rect 14457 5294 14515 5300
rect 14457 5260 14469 5294
rect 14503 5291 14515 5294
rect 15101 5294 15159 5300
rect 15101 5291 15113 5294
rect 14503 5263 15113 5291
rect 14503 5260 14515 5263
rect 14457 5254 14515 5260
rect 15101 5260 15113 5263
rect 15147 5260 15159 5294
rect 15101 5254 15159 5260
rect 15880 5292 15939 5298
rect 16291 5292 16297 5302
rect 15880 5258 15893 5292
rect 15927 5264 16297 5292
rect 15927 5258 15939 5264
rect 15880 5251 15939 5258
rect 16291 5255 16297 5264
rect 16296 5251 16297 5255
rect 16349 5255 16350 5302
rect 10311 5240 10363 5246
rect 14351 5238 14404 5245
rect 16296 5244 16349 5251
rect 11080 5234 11145 5235
rect 10363 5228 10949 5231
rect 10363 5225 10967 5228
rect 11074 5225 11145 5234
rect 10363 5224 11145 5225
rect 10363 5197 11088 5224
rect 10933 5194 10967 5197
rect 10311 5182 10363 5188
rect 11074 5190 11088 5197
rect 11122 5190 11145 5224
rect 11074 5184 11145 5190
rect 11080 5183 11145 5184
rect 14403 5186 14404 5238
rect 15009 5226 15067 5232
rect 15009 5192 15021 5226
rect 15055 5223 15067 5226
rect 15055 5195 15696 5223
rect 15055 5192 15067 5195
rect 15009 5186 15067 5192
rect 14351 5179 14404 5186
rect 15657 5164 15696 5195
rect 16199 5213 16249 5214
rect 16199 5211 16259 5213
rect 16378 5211 16415 5368
rect 17401 5362 17459 5368
rect 17401 5328 17413 5362
rect 17447 5359 17459 5362
rect 18137 5362 18195 5368
rect 18137 5359 18149 5362
rect 17447 5331 18149 5359
rect 17447 5328 17459 5331
rect 17401 5322 17459 5328
rect 18137 5328 18149 5331
rect 18183 5359 18195 5362
rect 18505 5362 18563 5368
rect 18505 5359 18517 5362
rect 18183 5331 18517 5359
rect 18183 5328 18195 5331
rect 18137 5322 18195 5328
rect 18505 5328 18517 5331
rect 18551 5328 18563 5362
rect 18505 5322 18563 5328
rect 18684 5302 18737 5308
rect 18683 5301 18742 5302
rect 16849 5294 16907 5300
rect 16849 5260 16861 5294
rect 16895 5291 16907 5294
rect 17493 5294 17551 5300
rect 17493 5291 17505 5294
rect 16895 5263 17505 5291
rect 16895 5260 16907 5263
rect 16849 5254 16907 5260
rect 17493 5260 17505 5263
rect 17539 5260 17551 5294
rect 17493 5254 17551 5260
rect 18272 5292 18331 5298
rect 18683 5292 18685 5301
rect 18272 5258 18285 5292
rect 18319 5264 18685 5292
rect 18319 5258 18331 5264
rect 18272 5251 18331 5258
rect 18683 5255 18685 5264
rect 18684 5249 18685 5255
rect 18737 5255 18742 5301
rect 16199 5207 16415 5211
rect 16199 5173 16213 5207
rect 16247 5174 16415 5207
rect 16746 5239 16799 5246
rect 18684 5242 18737 5249
rect 16798 5187 16799 5239
rect 16746 5180 16799 5187
rect 17401 5226 17459 5232
rect 17401 5192 17413 5226
rect 17447 5223 17459 5226
rect 17447 5195 18088 5223
rect 17447 5192 17459 5195
rect 17401 5186 17459 5192
rect 16247 5173 16259 5174
rect 16199 5166 16259 5173
rect 18049 5164 18088 5195
rect 18596 5211 18653 5214
rect 18770 5211 18807 5368
rect 19793 5362 19851 5368
rect 19793 5328 19805 5362
rect 19839 5359 19851 5362
rect 20529 5362 20587 5368
rect 20529 5359 20541 5362
rect 19839 5331 20541 5359
rect 19839 5328 19851 5331
rect 19793 5322 19851 5328
rect 20529 5328 20541 5331
rect 20575 5359 20587 5362
rect 20897 5362 20955 5368
rect 20897 5359 20909 5362
rect 20575 5331 20909 5359
rect 20575 5328 20587 5331
rect 20529 5322 20587 5328
rect 20897 5328 20909 5331
rect 20943 5328 20955 5362
rect 21081 5359 21082 5411
rect 21134 5368 21199 5405
rect 21081 5351 21134 5359
rect 20897 5322 20955 5328
rect 21076 5303 21129 5309
rect 21075 5302 21134 5303
rect 19241 5294 19299 5300
rect 19241 5260 19253 5294
rect 19287 5291 19299 5294
rect 19885 5294 19943 5300
rect 19885 5291 19897 5294
rect 19287 5263 19897 5291
rect 19287 5260 19299 5263
rect 19241 5254 19299 5260
rect 19885 5260 19897 5263
rect 19931 5260 19943 5294
rect 19885 5254 19943 5260
rect 20664 5293 20723 5299
rect 21075 5293 21077 5302
rect 20664 5259 20677 5293
rect 20711 5265 21077 5293
rect 20711 5259 20723 5265
rect 20664 5252 20723 5259
rect 21075 5256 21077 5265
rect 21076 5250 21077 5256
rect 21129 5256 21134 5302
rect 18596 5208 18807 5211
rect 18596 5174 18610 5208
rect 18644 5174 18807 5208
rect 19136 5240 19189 5247
rect 21076 5243 21129 5250
rect 19188 5188 19189 5240
rect 19136 5181 19189 5188
rect 19793 5226 19851 5232
rect 19793 5192 19805 5226
rect 19839 5223 19851 5226
rect 19839 5195 20480 5223
rect 19839 5192 19851 5195
rect 19793 5186 19851 5192
rect 14733 5158 14791 5164
rect 14733 5124 14745 5158
rect 14779 5155 14791 5158
rect 15469 5158 15527 5164
rect 15469 5155 15481 5158
rect 14779 5127 15481 5155
rect 14779 5124 14791 5127
rect 14733 5118 14791 5124
rect 15469 5124 15481 5127
rect 15515 5124 15527 5158
rect 15469 5118 15527 5124
rect 15657 5158 15715 5164
rect 15657 5124 15669 5158
rect 15703 5155 15715 5158
rect 16021 5158 16079 5164
rect 16021 5155 16033 5158
rect 15703 5127 16033 5155
rect 15703 5124 15715 5127
rect 15657 5118 15715 5124
rect 16021 5124 16033 5127
rect 16067 5124 16079 5158
rect 17125 5158 17183 5164
rect 16439 5135 16492 5142
rect 16021 5118 16079 5124
rect 16294 5128 16356 5134
rect 13812 5100 13878 5101
rect 13812 5048 13819 5100
rect 13871 5048 13878 5100
rect 16294 5094 16308 5128
rect 16342 5127 16356 5128
rect 16342 5094 16439 5127
rect 16294 5093 16439 5094
rect 16294 5088 16356 5093
rect 16491 5083 16492 5135
rect 17125 5124 17137 5158
rect 17171 5155 17183 5158
rect 17861 5158 17919 5164
rect 17861 5155 17873 5158
rect 17171 5127 17873 5155
rect 17171 5124 17183 5127
rect 17125 5118 17183 5124
rect 17861 5124 17873 5127
rect 17907 5124 17919 5158
rect 17861 5118 17919 5124
rect 18049 5158 18107 5164
rect 18049 5124 18061 5158
rect 18095 5155 18107 5158
rect 18413 5158 18471 5164
rect 18596 5161 18653 5174
rect 20441 5164 20480 5195
rect 20988 5211 21042 5215
rect 21162 5211 21199 5368
rect 22185 5362 22243 5368
rect 22185 5328 22197 5362
rect 22231 5359 22243 5362
rect 22921 5362 22979 5368
rect 22921 5359 22933 5362
rect 22231 5331 22933 5359
rect 22231 5328 22243 5331
rect 22185 5322 22243 5328
rect 22921 5328 22933 5331
rect 22967 5359 22979 5362
rect 23289 5362 23347 5368
rect 23289 5359 23301 5362
rect 22967 5331 23301 5359
rect 22967 5328 22979 5331
rect 22921 5322 22979 5328
rect 23289 5328 23301 5331
rect 23335 5328 23347 5362
rect 23289 5322 23347 5328
rect 24510 5343 24556 5421
rect 24670 5481 24716 5559
rect 24670 5421 24676 5481
rect 24710 5421 24716 5481
rect 24670 5409 24716 5421
rect 21633 5294 21691 5300
rect 21633 5260 21645 5294
rect 21679 5291 21691 5294
rect 22277 5294 22335 5300
rect 22277 5291 22289 5294
rect 21679 5263 22289 5291
rect 21679 5260 21691 5263
rect 21633 5254 21691 5260
rect 22277 5260 22289 5263
rect 22323 5260 22335 5294
rect 22277 5254 22335 5260
rect 23021 5294 23092 5302
rect 20988 5208 21199 5211
rect 20988 5174 21001 5208
rect 21035 5174 21199 5208
rect 21530 5237 21583 5244
rect 23021 5242 23029 5294
rect 23081 5242 23092 5294
rect 21582 5185 21583 5237
rect 23377 5237 23383 5289
rect 23435 5237 23441 5289
rect 24510 5283 24516 5343
rect 24550 5283 24556 5343
rect 24510 5271 24556 5283
rect 24670 5343 24716 5355
rect 24670 5283 24676 5343
rect 24710 5283 24716 5343
rect 23377 5236 23441 5237
rect 22185 5226 22243 5232
rect 22185 5192 22197 5226
rect 22231 5223 22243 5226
rect 22231 5195 22872 5223
rect 22231 5192 22243 5195
rect 22185 5186 22243 5192
rect 21530 5178 21583 5185
rect 18413 5155 18425 5158
rect 18095 5127 18425 5155
rect 18095 5124 18107 5127
rect 18049 5118 18107 5124
rect 18413 5124 18425 5127
rect 18459 5124 18471 5158
rect 19517 5158 19575 5164
rect 18413 5118 18471 5124
rect 18690 5115 18757 5125
rect 18861 5124 18914 5131
rect 16439 5076 16492 5083
rect 16581 5089 16634 5101
rect 16581 5055 16594 5089
rect 16628 5080 16634 5089
rect 17030 5099 17096 5100
rect 17030 5080 17037 5099
rect 16628 5055 17037 5080
rect 16581 5052 17037 5055
rect 16581 5049 16634 5052
rect 17030 5047 17037 5052
rect 17089 5080 17096 5099
rect 18690 5081 18708 5115
rect 18742 5081 18861 5115
rect 17089 5052 17295 5080
rect 18690 5071 18757 5081
rect 18913 5072 18914 5124
rect 19517 5124 19529 5158
rect 19563 5155 19575 5158
rect 20253 5158 20311 5164
rect 20253 5155 20265 5158
rect 19563 5127 20265 5155
rect 19563 5124 19575 5127
rect 19517 5118 19575 5124
rect 20253 5124 20265 5127
rect 20299 5124 20311 5158
rect 20253 5118 20311 5124
rect 20441 5158 20499 5164
rect 20441 5124 20453 5158
rect 20487 5155 20499 5158
rect 20805 5158 20863 5164
rect 20988 5163 21042 5174
rect 22833 5164 22872 5195
rect 24510 5205 24556 5217
rect 20805 5155 20817 5158
rect 20487 5127 20817 5155
rect 20487 5124 20499 5127
rect 20441 5118 20499 5124
rect 20805 5124 20817 5127
rect 20851 5124 20863 5158
rect 21909 5158 21967 5164
rect 20805 5118 20863 5124
rect 21078 5123 21145 5133
rect 21249 5132 21302 5139
rect 19422 5100 19488 5101
rect 18861 5065 18914 5072
rect 18970 5088 19028 5095
rect 18970 5054 18982 5088
rect 19016 5079 19028 5088
rect 19422 5079 19429 5100
rect 19016 5054 19429 5079
rect 17089 5047 17096 5052
rect 18970 5051 19429 5054
rect 18970 5048 19028 5051
rect 19422 5048 19429 5051
rect 19481 5079 19488 5100
rect 21078 5089 21096 5123
rect 21130 5089 21249 5123
rect 21078 5079 21145 5089
rect 21301 5080 21302 5132
rect 21909 5124 21921 5158
rect 21955 5155 21967 5158
rect 22645 5158 22703 5164
rect 22645 5155 22657 5158
rect 21955 5127 22657 5155
rect 21955 5124 21967 5127
rect 21909 5118 21967 5124
rect 22645 5124 22657 5127
rect 22691 5124 22703 5158
rect 22645 5118 22703 5124
rect 22833 5158 22891 5164
rect 22833 5124 22845 5158
rect 22879 5155 22891 5158
rect 23197 5158 23255 5164
rect 23197 5155 23209 5158
rect 22879 5127 23209 5155
rect 22879 5124 22891 5127
rect 22833 5118 22891 5124
rect 23197 5124 23209 5127
rect 23243 5124 23255 5158
rect 23197 5118 23255 5124
rect 21811 5101 21877 5102
rect 19481 5051 19688 5079
rect 21249 5073 21302 5080
rect 21361 5094 21422 5100
rect 21361 5060 21376 5094
rect 21410 5080 21422 5094
rect 21811 5080 21818 5101
rect 21410 5060 21818 5080
rect 21361 5052 21818 5060
rect 19481 5048 19488 5051
rect 21361 5048 21422 5052
rect 21811 5049 21818 5052
rect 21870 5080 21877 5101
rect 23543 5080 23795 5162
rect 21870 5052 22080 5080
rect 21870 5049 21877 5052
rect 23543 5019 23625 5080
rect 10932 4988 23625 5019
rect 10932 4954 11086 4988
rect 11120 4954 11178 4988
rect 11212 4954 11270 4988
rect 11304 4954 11362 4988
rect 11396 4954 11454 4988
rect 11488 4954 11546 4988
rect 11580 4954 11638 4988
rect 11672 4954 11730 4988
rect 11764 4954 11822 4988
rect 11856 4954 11894 4988
rect 11928 4954 11986 4988
rect 12020 4954 12078 4988
rect 12112 4954 12170 4988
rect 12204 4954 12262 4988
rect 12296 4954 12354 4988
rect 12388 4954 12446 4988
rect 12480 4954 12538 4988
rect 12572 4954 12630 4988
rect 12664 4954 12722 4988
rect 12756 4954 12814 4988
rect 12848 4954 12906 4988
rect 12940 4954 12998 4988
rect 13032 4954 13090 4988
rect 13124 4954 13182 4988
rect 13216 4954 13274 4988
rect 13308 4954 13366 4988
rect 13400 4954 13458 4988
rect 13492 4954 13550 4988
rect 13584 4954 13642 4988
rect 13676 4954 13734 4988
rect 13768 4954 13826 4988
rect 13860 4954 13918 4988
rect 13952 4954 14010 4988
rect 14044 4954 14102 4988
rect 14136 4954 14194 4988
rect 14228 4954 14286 4988
rect 14320 4954 14378 4988
rect 14412 4954 14470 4988
rect 14504 4954 14562 4988
rect 14596 4954 14654 4988
rect 14688 4954 14746 4988
rect 14780 4954 14838 4988
rect 14872 4954 14930 4988
rect 14964 4954 15022 4988
rect 15056 4954 15114 4988
rect 15148 4954 15206 4988
rect 15240 4954 15298 4988
rect 15332 4954 15390 4988
rect 15424 4954 15482 4988
rect 15516 4954 15574 4988
rect 15608 4954 15666 4988
rect 15700 4954 15758 4988
rect 15792 4954 15850 4988
rect 15884 4954 15942 4988
rect 15976 4954 16034 4988
rect 16068 4954 16126 4988
rect 16160 4954 16218 4988
rect 16252 4954 16310 4988
rect 16344 4954 16402 4988
rect 16436 4954 16494 4988
rect 16528 4954 16586 4988
rect 16620 4954 16678 4988
rect 16712 4954 16770 4988
rect 16804 4954 16862 4988
rect 16896 4954 16954 4988
rect 16988 4954 17046 4988
rect 17080 4954 17138 4988
rect 17172 4954 17230 4988
rect 17264 4954 17322 4988
rect 17356 4954 17414 4988
rect 17448 4954 17506 4988
rect 17540 4954 17598 4988
rect 17632 4954 17690 4988
rect 17724 4954 17782 4988
rect 17816 4954 17874 4988
rect 17908 4954 17966 4988
rect 18000 4954 18058 4988
rect 18092 4954 18150 4988
rect 18184 4954 18242 4988
rect 18276 4954 18334 4988
rect 18368 4954 18426 4988
rect 18460 4954 18518 4988
rect 18552 4954 18610 4988
rect 18644 4954 18702 4988
rect 18736 4954 18794 4988
rect 18828 4954 18886 4988
rect 18920 4954 18978 4988
rect 19012 4954 19070 4988
rect 19104 4954 19162 4988
rect 19196 4954 19254 4988
rect 19288 4954 19346 4988
rect 19380 4954 19438 4988
rect 19472 4954 19530 4988
rect 19564 4954 19622 4988
rect 19656 4954 19714 4988
rect 19748 4954 19806 4988
rect 19840 4954 19898 4988
rect 19932 4954 19990 4988
rect 20024 4954 20082 4988
rect 20116 4954 20174 4988
rect 20208 4954 20266 4988
rect 20300 4954 20358 4988
rect 20392 4954 20450 4988
rect 20484 4954 20542 4988
rect 20576 4954 20634 4988
rect 20668 4954 20726 4988
rect 20760 4954 20818 4988
rect 20852 4954 20910 4988
rect 20944 4954 21002 4988
rect 21036 4954 21094 4988
rect 21128 4954 21186 4988
rect 21220 4954 21278 4988
rect 21312 4954 21370 4988
rect 21404 4954 21462 4988
rect 21496 4954 21554 4988
rect 21588 4954 21646 4988
rect 21680 4954 21738 4988
rect 21772 4954 21830 4988
rect 21864 4954 21922 4988
rect 21956 4954 22014 4988
rect 22048 4954 22106 4988
rect 22140 4954 22198 4988
rect 22232 4954 22290 4988
rect 22324 4954 22382 4988
rect 22416 4954 22474 4988
rect 22508 4954 22566 4988
rect 22600 4954 22658 4988
rect 22692 4954 22750 4988
rect 22784 4954 22842 4988
rect 22876 4954 22934 4988
rect 22968 4954 23026 4988
rect 23060 4954 23118 4988
rect 23152 4954 23210 4988
rect 23244 4954 23302 4988
rect 23336 4954 23394 4988
rect 23428 4954 23625 4988
rect 10932 4934 23625 4954
rect 23775 4934 23795 5080
rect 24510 5145 24516 5205
rect 24550 5145 24556 5205
rect 24510 5067 24556 5145
rect 24670 5205 24716 5283
rect 24670 5145 24676 5205
rect 24710 5145 24716 5205
rect 24670 5133 24716 5145
rect 24510 5007 24516 5067
rect 24550 5007 24556 5067
rect 24510 4995 24556 5007
rect 24670 5067 24716 5079
rect 24670 5007 24676 5067
rect 24710 5007 24716 5067
rect 10932 4923 23795 4934
rect 13812 4858 13878 4859
rect 11952 4847 11959 4858
rect 11947 4818 11959 4847
rect 11952 4806 11959 4818
rect 12011 4847 12018 4858
rect 13812 4847 13819 4858
rect 12011 4818 13819 4847
rect 12011 4806 12018 4818
rect 13812 4806 13819 4818
rect 13871 4847 13878 4858
rect 14344 4858 14410 4859
rect 14344 4847 14351 4858
rect 13871 4818 14351 4847
rect 13871 4806 13878 4818
rect 14344 4806 14351 4818
rect 14403 4847 14410 4858
rect 15748 4858 15814 4859
rect 15748 4847 15755 4858
rect 14403 4819 15755 4847
rect 14403 4806 14410 4819
rect 15748 4806 15755 4819
rect 15807 4847 15814 4858
rect 16733 4858 16799 4859
rect 16733 4847 16740 4858
rect 15807 4819 16740 4847
rect 15807 4806 15814 4819
rect 16733 4806 16740 4819
rect 16792 4847 16799 4858
rect 18140 4858 18206 4859
rect 18140 4847 18147 4858
rect 16792 4819 18147 4847
rect 16792 4806 16799 4819
rect 18140 4806 18147 4819
rect 18199 4847 18206 4858
rect 19123 4858 19189 4859
rect 19123 4847 19130 4858
rect 18199 4819 19130 4847
rect 18199 4806 18206 4819
rect 19123 4806 19130 4819
rect 19182 4847 19189 4858
rect 20537 4858 20603 4859
rect 20537 4847 20544 4858
rect 19182 4819 20544 4847
rect 19182 4806 19189 4819
rect 20537 4806 20544 4819
rect 20596 4847 20603 4858
rect 21513 4858 21579 4859
rect 21513 4847 21520 4858
rect 20596 4819 21520 4847
rect 20596 4806 20603 4819
rect 21513 4806 21520 4819
rect 21572 4847 21579 4858
rect 22925 4858 22991 4859
rect 22925 4847 22932 4858
rect 21572 4819 22932 4847
rect 21572 4806 21579 4819
rect 22925 4806 22932 4819
rect 22984 4847 22991 4858
rect 22984 4819 23404 4847
rect 22984 4806 22991 4819
rect 23537 4746 23795 4923
rect 10952 4718 23795 4746
rect 24510 4929 24556 4941
rect 24510 4869 24516 4929
rect 24550 4869 24556 4929
rect 24510 4791 24556 4869
rect 24670 4929 24716 5007
rect 24670 4869 24676 4929
rect 24710 4869 24716 4929
rect 24670 4857 24716 4869
rect 24510 4731 24516 4791
rect 24550 4731 24556 4791
rect 24670 4791 24716 4803
rect 24670 4767 24676 4791
rect 24510 4719 24556 4731
rect 24631 4751 24676 4767
rect 24710 4767 24716 4791
rect 24710 4751 24738 4767
rect 24631 4699 24667 4751
rect 24719 4699 24738 4751
rect 10949 4685 23568 4690
rect 10753 4659 23568 4685
rect 24631 4683 24738 4699
rect 25191 4754 25523 4760
rect 25191 4702 25209 4754
rect 25261 4702 25289 4754
rect 25341 4702 25369 4754
rect 25421 4702 25449 4754
rect 25501 4702 25523 4754
rect 25191 4692 25523 4702
rect 25923 4754 26255 4760
rect 25923 4702 25941 4754
rect 25993 4702 26021 4754
rect 26073 4702 26101 4754
rect 26153 4702 26181 4754
rect 26233 4702 26255 4754
rect 25923 4692 26255 4702
rect 26426 4663 26484 5791
rect 26525 4754 26857 4760
rect 26525 4702 26547 4754
rect 26599 4702 26627 4754
rect 26679 4702 26707 4754
rect 26759 4702 26787 4754
rect 26839 4702 26857 4754
rect 26525 4692 26857 4702
rect 27135 4754 27467 4760
rect 27135 4702 27153 4754
rect 27205 4702 27233 4754
rect 27285 4702 27313 4754
rect 27365 4702 27393 4754
rect 27445 4702 27467 4754
rect 27135 4692 27467 4702
rect 27737 4754 28069 4760
rect 27737 4702 27759 4754
rect 27811 4702 27839 4754
rect 27891 4702 27919 4754
rect 27971 4702 27999 4754
rect 28051 4702 28069 4754
rect 27737 4692 28069 4702
rect 28473 4754 28805 4760
rect 28473 4702 28491 4754
rect 28543 4702 28571 4754
rect 28623 4702 28651 4754
rect 28703 4702 28731 4754
rect 28783 4702 28805 4754
rect 28473 4692 28805 4702
rect 10753 4658 13660 4659
rect 10753 4646 11118 4658
rect 10753 4500 10823 4646
rect 10973 4624 11118 4646
rect 11152 4650 11210 4658
rect 11244 4650 11302 4658
rect 11152 4624 11175 4650
rect 11336 4624 11394 4658
rect 11428 4624 11486 4658
rect 11520 4624 11578 4658
rect 11612 4650 11670 4658
rect 11704 4650 11762 4658
rect 11612 4624 11621 4650
rect 11796 4624 11854 4658
rect 11888 4654 13660 4658
rect 11888 4624 12187 4654
rect 10973 4504 11175 4624
rect 11325 4504 11621 4624
rect 11771 4508 12187 4624
rect 12337 4508 12853 4654
rect 13003 4638 13660 4654
rect 13003 4508 13235 4638
rect 11771 4504 13235 4508
rect 10973 4500 13235 4504
rect 10753 4492 13235 4500
rect 13385 4625 13660 4638
rect 13694 4625 13752 4659
rect 13786 4625 13844 4659
rect 13878 4625 13917 4659
rect 13951 4625 14009 4659
rect 14043 4625 14101 4659
rect 14135 4625 14193 4659
rect 14227 4625 14285 4659
rect 14319 4625 14377 4659
rect 14411 4625 14469 4659
rect 14503 4625 14561 4659
rect 14595 4625 14653 4659
rect 14687 4625 14745 4659
rect 14779 4625 14837 4659
rect 14871 4625 14929 4659
rect 14963 4625 15021 4659
rect 15055 4625 15113 4659
rect 15147 4625 15205 4659
rect 15239 4625 15297 4659
rect 15331 4625 15389 4659
rect 15423 4625 15481 4659
rect 15515 4625 15573 4659
rect 15607 4625 15665 4659
rect 15699 4625 15757 4659
rect 15791 4625 15849 4659
rect 15883 4625 15941 4659
rect 15975 4625 16033 4659
rect 16067 4625 16125 4659
rect 16159 4625 16217 4659
rect 16251 4625 16309 4659
rect 16343 4625 16401 4659
rect 16435 4625 16493 4659
rect 16527 4625 16585 4659
rect 16619 4625 16677 4659
rect 16711 4625 16769 4659
rect 16803 4625 16861 4659
rect 16895 4625 16953 4659
rect 16987 4625 17045 4659
rect 17079 4625 17137 4659
rect 17171 4625 17229 4659
rect 17263 4625 17321 4659
rect 17355 4625 17413 4659
rect 17447 4625 17505 4659
rect 17539 4625 17597 4659
rect 17631 4625 17689 4659
rect 17723 4625 17781 4659
rect 17815 4625 17873 4659
rect 17907 4625 17965 4659
rect 17999 4625 18057 4659
rect 18091 4625 18149 4659
rect 18183 4625 18241 4659
rect 18275 4625 18333 4659
rect 18367 4625 18425 4659
rect 18459 4625 18517 4659
rect 18551 4625 18609 4659
rect 18643 4625 18701 4659
rect 18735 4625 18793 4659
rect 18827 4625 18885 4659
rect 18919 4625 18977 4659
rect 19011 4625 19069 4659
rect 19103 4625 19161 4659
rect 19195 4625 19253 4659
rect 19287 4625 19345 4659
rect 19379 4625 19437 4659
rect 19471 4625 19529 4659
rect 19563 4625 19621 4659
rect 19655 4625 19713 4659
rect 19747 4625 19805 4659
rect 19839 4625 19897 4659
rect 19931 4625 19989 4659
rect 20023 4625 20081 4659
rect 20115 4625 20173 4659
rect 20207 4625 20265 4659
rect 20299 4625 20357 4659
rect 20391 4625 20449 4659
rect 20483 4625 20541 4659
rect 20575 4625 20633 4659
rect 20667 4625 20725 4659
rect 20759 4625 20817 4659
rect 20851 4625 20909 4659
rect 20943 4625 21001 4659
rect 21035 4625 21093 4659
rect 21127 4625 21185 4659
rect 21219 4625 21277 4659
rect 21311 4625 21369 4659
rect 21403 4625 21461 4659
rect 21495 4625 21553 4659
rect 21587 4625 21645 4659
rect 21679 4625 21737 4659
rect 21771 4625 21829 4659
rect 21863 4625 21921 4659
rect 21955 4625 22013 4659
rect 22047 4625 22105 4659
rect 22139 4625 22197 4659
rect 22231 4625 22289 4659
rect 22323 4625 22381 4659
rect 22415 4625 22473 4659
rect 22507 4625 22565 4659
rect 22599 4625 22657 4659
rect 22691 4625 22749 4659
rect 22783 4625 22841 4659
rect 22875 4625 22933 4659
rect 22967 4625 23025 4659
rect 23059 4625 23117 4659
rect 23151 4625 23209 4659
rect 23243 4625 23301 4659
rect 23335 4625 23393 4659
rect 23427 4625 23568 4659
rect 25545 4635 26484 4663
rect 13385 4594 23568 4625
rect 28852 4607 28910 5791
rect 29075 4754 29407 4760
rect 29075 4702 29097 4754
rect 29149 4702 29177 4754
rect 29229 4702 29257 4754
rect 29309 4702 29337 4754
rect 29389 4702 29407 4754
rect 29075 4692 29407 4702
rect 13385 4492 13489 4594
rect 25545 4579 28910 4607
rect 29708 4551 29767 5791
rect 30320 5804 30366 5816
rect 30320 5744 30326 5804
rect 30360 5744 30366 5804
rect 30320 5692 30366 5744
rect 30408 5813 30646 5842
rect 30408 5804 30454 5813
rect 30408 5744 30414 5804
rect 30448 5744 30454 5804
rect 30679 5792 31047 5823
rect 30679 5784 30708 5792
rect 30408 5732 30454 5744
rect 30565 5768 30708 5784
rect 30565 5716 30601 5768
rect 30653 5758 30708 5768
rect 30742 5758 30800 5792
rect 30834 5758 30892 5792
rect 30926 5758 30984 5792
rect 31018 5784 31047 5792
rect 31018 5758 31048 5784
rect 30653 5716 31048 5758
rect 30565 5700 31048 5716
rect 30320 5676 30481 5692
rect 30320 5624 30410 5676
rect 30462 5624 30481 5676
rect 30320 5608 30481 5624
rect 25545 4523 29767 4551
rect 29809 4754 30141 4760
rect 29809 4702 29831 4754
rect 29883 4702 29911 4754
rect 29963 4702 29991 4754
rect 30043 4702 30071 4754
rect 30123 4702 30141 4754
rect 29809 4495 30141 4702
rect 10753 4460 13489 4492
rect 13998 4489 14056 4495
rect 13998 4455 14010 4489
rect 14044 4486 14056 4489
rect 14366 4489 14424 4495
rect 14366 4486 14378 4489
rect 14044 4458 14378 4486
rect 14044 4455 14056 4458
rect 13998 4449 14056 4455
rect 14366 4455 14378 4458
rect 14412 4486 14424 4489
rect 15102 4489 15160 4495
rect 15102 4486 15114 4489
rect 14412 4458 15114 4486
rect 14412 4455 14424 4458
rect 14366 4449 14424 4455
rect 15102 4455 15114 4458
rect 15148 4455 15160 4489
rect 15102 4449 15160 4455
rect 16390 4489 16448 4495
rect 16390 4455 16402 4489
rect 16436 4486 16448 4489
rect 16758 4489 16816 4495
rect 16758 4486 16770 4489
rect 16436 4458 16770 4486
rect 16436 4455 16448 4458
rect 16390 4449 16448 4455
rect 16758 4455 16770 4458
rect 16804 4486 16816 4489
rect 17494 4489 17552 4495
rect 17494 4486 17506 4489
rect 16804 4458 17506 4486
rect 16804 4455 16816 4458
rect 16758 4449 16816 4455
rect 17494 4455 17506 4458
rect 17540 4455 17552 4489
rect 17494 4449 17552 4455
rect 18782 4489 18840 4495
rect 18782 4455 18794 4489
rect 18828 4486 18840 4489
rect 19150 4489 19208 4495
rect 19150 4486 19162 4489
rect 18828 4458 19162 4486
rect 18828 4455 18840 4458
rect 18782 4449 18840 4455
rect 19150 4455 19162 4458
rect 19196 4486 19208 4489
rect 19886 4489 19944 4495
rect 19886 4486 19898 4489
rect 19196 4458 19898 4486
rect 19196 4455 19208 4458
rect 19150 4449 19208 4455
rect 19886 4455 19898 4458
rect 19932 4455 19944 4489
rect 19886 4449 19944 4455
rect 21174 4489 21232 4495
rect 21174 4455 21186 4489
rect 21220 4486 21232 4489
rect 21542 4489 21600 4495
rect 21542 4486 21554 4489
rect 21220 4458 21554 4486
rect 21220 4455 21232 4458
rect 21174 4449 21232 4455
rect 21542 4455 21554 4458
rect 21588 4486 21600 4489
rect 22278 4489 22336 4495
rect 22278 4486 22290 4489
rect 21588 4458 22290 4486
rect 21588 4455 21600 4458
rect 21542 4449 21600 4455
rect 22278 4455 22290 4458
rect 22324 4455 22336 4489
rect 22278 4449 22336 4455
rect 25492 4467 30141 4495
rect 13077 4430 13144 4431
rect 10931 4389 12095 4417
rect 10623 4311 10630 4363
rect 10682 4354 10688 4363
rect 10931 4354 10965 4389
rect 10682 4320 10965 4354
rect 10682 4311 10688 4320
rect 11113 4303 11119 4355
rect 11171 4303 11177 4355
rect 11720 4303 11726 4355
rect 11778 4303 11784 4355
rect 12061 4349 12095 4389
rect 13077 4378 13085 4430
rect 13137 4405 13144 4430
rect 13523 4429 13589 4430
rect 13523 4405 13530 4429
rect 13137 4378 13530 4405
rect 13085 4377 13530 4378
rect 13582 4377 13589 4429
rect 13796 4426 13857 4433
rect 13796 4392 13810 4426
rect 13844 4421 13857 4426
rect 14644 4421 14652 4430
rect 13844 4393 14652 4421
rect 13844 4392 13857 4393
rect 13796 4386 13857 4392
rect 14644 4378 14652 4393
rect 14704 4378 14711 4430
rect 15010 4421 15068 4427
rect 15010 4387 15022 4421
rect 15056 4418 15068 4421
rect 15654 4421 15712 4427
rect 15654 4418 15666 4421
rect 15056 4390 15666 4418
rect 15056 4387 15068 4390
rect 15010 4381 15068 4387
rect 15654 4387 15666 4390
rect 15700 4387 15712 4421
rect 15654 4381 15712 4387
rect 17402 4421 17460 4427
rect 17402 4387 17414 4421
rect 17448 4418 17460 4421
rect 18046 4421 18104 4427
rect 18046 4418 18058 4421
rect 17448 4390 18058 4418
rect 17448 4387 17460 4390
rect 17402 4381 17460 4387
rect 18046 4387 18058 4390
rect 18092 4387 18104 4421
rect 18046 4381 18104 4387
rect 19794 4421 19852 4427
rect 19794 4387 19806 4421
rect 19840 4418 19852 4421
rect 20438 4421 20496 4427
rect 20438 4418 20450 4421
rect 19840 4390 20450 4418
rect 19840 4387 19852 4390
rect 19794 4381 19852 4387
rect 20438 4387 20450 4390
rect 20484 4387 20496 4421
rect 20438 4381 20496 4387
rect 22186 4421 22244 4427
rect 22186 4387 22198 4421
rect 22232 4418 22244 4421
rect 22830 4421 22888 4427
rect 22830 4418 22842 4421
rect 22232 4390 22842 4418
rect 22232 4387 22244 4390
rect 22186 4381 22244 4387
rect 22830 4387 22842 4390
rect 22876 4387 22888 4421
rect 22830 4381 22888 4387
rect 18147 4369 18200 4376
rect 12475 4357 12541 4358
rect 12475 4349 12482 4357
rect 12061 4321 12482 4349
rect 12475 4305 12482 4321
rect 12534 4349 12541 4357
rect 13619 4352 13665 4364
rect 13619 4349 13625 4352
rect 12534 4321 13625 4349
rect 12534 4305 12541 4321
rect 13619 4318 13625 4321
rect 13659 4318 13665 4352
rect 13619 4306 13665 4318
rect 13909 4351 13958 4364
rect 13909 4317 13918 4351
rect 13952 4317 13958 4351
rect 13909 4310 13958 4317
rect 14004 4359 14300 4365
rect 15756 4359 15809 4366
rect 14004 4326 14247 4359
rect 13916 4146 13955 4310
rect 14004 4146 14043 4326
rect 14239 4325 14247 4326
rect 14281 4325 14300 4359
rect 15102 4353 15160 4359
rect 15102 4350 15114 4353
rect 14239 4313 14300 4325
rect 14473 4322 15114 4350
rect 14473 4291 14512 4322
rect 15102 4319 15114 4322
rect 15148 4319 15160 4353
rect 15102 4313 15160 4319
rect 15808 4307 15809 4359
rect 16647 4311 16654 4363
rect 16706 4311 16713 4363
rect 17494 4353 17552 4359
rect 17494 4350 17506 4353
rect 16865 4322 17506 4350
rect 15756 4300 15809 4307
rect 14090 4285 14148 4291
rect 14090 4251 14102 4285
rect 14136 4282 14148 4285
rect 14454 4285 14512 4291
rect 14454 4282 14466 4285
rect 14136 4254 14466 4282
rect 14136 4251 14148 4254
rect 14090 4245 14148 4251
rect 14454 4251 14466 4254
rect 14500 4251 14512 4285
rect 14454 4245 14512 4251
rect 14638 4293 14702 4294
rect 14638 4241 14644 4293
rect 14696 4282 14702 4293
rect 16865 4291 16904 4322
rect 17494 4319 17506 4322
rect 17540 4319 17552 4353
rect 17494 4313 17552 4319
rect 18199 4317 18200 4369
rect 20538 4365 20591 4372
rect 18147 4310 18200 4317
rect 19034 4311 19041 4363
rect 19093 4311 19100 4363
rect 19886 4353 19944 4359
rect 19886 4350 19898 4353
rect 19257 4322 19898 4350
rect 15378 4285 15436 4291
rect 15378 4282 15390 4285
rect 14696 4254 15390 4282
rect 14696 4241 14702 4254
rect 15378 4251 15390 4254
rect 15424 4251 15436 4285
rect 15378 4245 15436 4251
rect 16482 4285 16540 4291
rect 16482 4251 16494 4285
rect 16528 4282 16540 4285
rect 16846 4285 16904 4291
rect 16846 4282 16858 4285
rect 16528 4254 16858 4282
rect 16528 4251 16540 4254
rect 16482 4245 16540 4251
rect 16846 4251 16858 4254
rect 16892 4251 16904 4285
rect 16846 4245 16904 4251
rect 17031 4292 17097 4293
rect 17031 4240 17038 4292
rect 17090 4282 17097 4292
rect 19257 4291 19296 4322
rect 19886 4319 19898 4322
rect 19932 4319 19944 4353
rect 19886 4313 19944 4319
rect 20590 4313 20591 4365
rect 22930 4364 22983 4371
rect 20538 4306 20591 4313
rect 21437 4310 21444 4362
rect 21496 4310 21503 4362
rect 22278 4353 22336 4359
rect 22278 4350 22290 4353
rect 21649 4322 22290 4350
rect 17770 4285 17828 4291
rect 17770 4282 17782 4285
rect 17090 4254 17782 4282
rect 17090 4240 17097 4254
rect 17770 4251 17782 4254
rect 17816 4251 17828 4285
rect 18874 4285 18932 4291
rect 17770 4245 17828 4251
rect 18604 4261 18657 4268
rect 18656 4209 18657 4261
rect 18874 4251 18886 4285
rect 18920 4282 18932 4285
rect 19238 4285 19296 4291
rect 19238 4282 19250 4285
rect 18920 4254 19250 4282
rect 18920 4251 18932 4254
rect 18874 4245 18932 4251
rect 19238 4251 19250 4254
rect 19284 4251 19296 4285
rect 19238 4245 19296 4251
rect 19425 4291 19491 4292
rect 21649 4291 21688 4322
rect 22278 4319 22290 4322
rect 22324 4319 22336 4353
rect 22278 4313 22336 4319
rect 22982 4312 22983 4364
rect 22930 4305 22983 4312
rect 25492 4329 25546 4467
rect 25616 4372 25622 4424
rect 25674 4412 25680 4424
rect 28010 4412 28016 4424
rect 25674 4384 28016 4412
rect 25674 4372 25680 4384
rect 28010 4372 28016 4384
rect 28068 4412 28074 4424
rect 31076 4412 31104 5995
rect 28068 4384 31104 4412
rect 28068 4372 28074 4384
rect 25698 4329 25732 4332
rect 25790 4329 25824 4332
rect 25882 4329 25916 4332
rect 25974 4329 26008 4332
rect 26066 4329 26100 4332
rect 26158 4329 26192 4332
rect 26250 4329 26284 4332
rect 26342 4329 26376 4332
rect 26433 4329 26467 4332
rect 26526 4329 26560 4332
rect 26618 4329 26652 4332
rect 26710 4329 26744 4332
rect 26802 4329 26836 4332
rect 26894 4329 26928 4332
rect 26986 4329 27020 4332
rect 27078 4329 27112 4332
rect 27170 4329 27204 4332
rect 27262 4329 27296 4332
rect 27354 4329 27388 4332
rect 27446 4329 27480 4332
rect 27538 4329 27572 4332
rect 27630 4329 27664 4332
rect 27722 4329 27756 4332
rect 27814 4329 27848 4332
rect 27906 4329 27940 4332
rect 27998 4329 28032 4332
rect 28090 4329 28124 4332
rect 28182 4329 28216 4332
rect 28274 4329 28308 4332
rect 28366 4329 28400 4332
rect 28458 4329 28492 4332
rect 28550 4329 28584 4332
rect 28642 4329 28676 4332
rect 28734 4329 28768 4332
rect 28826 4329 28860 4332
rect 28918 4329 28952 4332
rect 29010 4329 29044 4332
rect 29102 4329 29136 4332
rect 29194 4329 29228 4332
rect 29286 4329 29320 4332
rect 29378 4329 29412 4332
rect 29470 4329 29504 4332
rect 29562 4329 29596 4332
rect 29654 4329 29688 4332
rect 29746 4329 29780 4332
rect 29838 4329 29872 4332
rect 29930 4329 29964 4332
rect 30022 4329 30056 4332
rect 30114 4329 30148 4332
rect 30206 4329 30240 4332
rect 30298 4329 30332 4332
rect 25492 4313 30361 4329
rect 25492 4312 29110 4313
rect 25492 4309 26746 4312
rect 25492 4307 26314 4309
rect 25492 4306 26113 4307
rect 25492 4298 25714 4306
rect 25766 4305 26113 4306
rect 25766 4298 25888 4305
rect 25940 4298 26113 4305
rect 26165 4298 26314 4307
rect 26366 4307 26746 4309
rect 26366 4298 26537 4307
rect 26589 4298 26746 4307
rect 19425 4239 19432 4291
rect 19484 4282 19491 4291
rect 20162 4285 20220 4291
rect 20162 4282 20174 4285
rect 19484 4254 20174 4282
rect 19484 4239 19491 4254
rect 20162 4251 20174 4254
rect 20208 4251 20220 4285
rect 21266 4285 21324 4291
rect 20162 4245 20220 4251
rect 20996 4262 21049 4269
rect 18604 4202 18657 4209
rect 21048 4210 21049 4262
rect 21266 4251 21278 4285
rect 21312 4282 21324 4285
rect 21630 4285 21688 4291
rect 21630 4282 21642 4285
rect 21312 4254 21642 4282
rect 21312 4251 21324 4254
rect 21266 4245 21324 4251
rect 21630 4251 21642 4254
rect 21676 4251 21688 4285
rect 21630 4245 21688 4251
rect 21811 4292 21877 4293
rect 21811 4240 21818 4292
rect 21870 4282 21877 4292
rect 22554 4285 22612 4291
rect 22554 4282 22566 4285
rect 21870 4254 22566 4282
rect 21870 4240 21877 4254
rect 22554 4251 22566 4254
rect 22600 4251 22612 4285
rect 22554 4245 22612 4251
rect 23386 4265 23439 4272
rect 20996 4203 21049 4210
rect 23438 4213 23439 4265
rect 25492 4264 25606 4298
rect 25640 4264 25698 4298
rect 25766 4264 25790 4298
rect 25824 4264 25882 4298
rect 25940 4264 25974 4298
rect 26008 4264 26066 4298
rect 26100 4264 26113 4298
rect 26192 4264 26250 4298
rect 26284 4264 26314 4298
rect 26376 4264 26434 4298
rect 26468 4264 26526 4298
rect 26589 4264 26618 4298
rect 26652 4264 26710 4298
rect 26744 4264 26746 4298
rect 25492 4254 25714 4264
rect 25766 4254 25888 4264
rect 25492 4253 25888 4254
rect 25940 4255 26113 4264
rect 26165 4257 26314 4264
rect 26366 4257 26537 4264
rect 26165 4255 26537 4257
rect 26589 4260 26746 4264
rect 26798 4309 27369 4312
rect 26798 4305 27164 4309
rect 26798 4298 26974 4305
rect 27026 4298 27164 4305
rect 27216 4298 27369 4309
rect 27421 4298 27568 4312
rect 27620 4307 28172 4312
rect 27620 4298 27784 4307
rect 27836 4298 28172 4307
rect 28224 4310 29110 4312
rect 28224 4309 28881 4310
rect 28224 4307 28649 4309
rect 28224 4298 28407 4307
rect 28459 4298 28649 4307
rect 28701 4298 28881 4309
rect 28933 4298 29110 4310
rect 29162 4312 30361 4313
rect 29162 4309 30243 4312
rect 29162 4305 29577 4309
rect 29162 4298 29359 4305
rect 29411 4298 29577 4305
rect 29629 4307 30243 4309
rect 29629 4305 30027 4307
rect 29629 4298 29806 4305
rect 29858 4298 30027 4305
rect 30079 4298 30243 4307
rect 26798 4264 26802 4298
rect 26836 4264 26894 4298
rect 26928 4264 26974 4298
rect 27026 4264 27078 4298
rect 27112 4264 27164 4298
rect 27216 4264 27262 4298
rect 27296 4264 27354 4298
rect 27421 4264 27446 4298
rect 27480 4264 27538 4298
rect 27620 4264 27630 4298
rect 27664 4264 27722 4298
rect 27756 4264 27784 4298
rect 27848 4264 27906 4298
rect 27940 4264 27998 4298
rect 28032 4264 28090 4298
rect 28124 4264 28172 4298
rect 28224 4264 28274 4298
rect 28308 4264 28366 4298
rect 28400 4264 28407 4298
rect 28492 4264 28550 4298
rect 28584 4264 28642 4298
rect 28701 4264 28734 4298
rect 28768 4264 28826 4298
rect 28860 4264 28881 4298
rect 28952 4264 29010 4298
rect 29044 4264 29102 4298
rect 29162 4264 29194 4298
rect 29228 4264 29286 4298
rect 29320 4264 29359 4298
rect 29412 4264 29470 4298
rect 29504 4264 29562 4298
rect 29629 4264 29654 4298
rect 29688 4264 29746 4298
rect 29780 4264 29806 4298
rect 29872 4264 29930 4298
rect 29964 4264 30022 4298
rect 30079 4264 30114 4298
rect 30148 4264 30206 4298
rect 30240 4264 30243 4298
rect 26798 4260 26974 4264
rect 26589 4255 26974 4260
rect 25940 4253 26974 4255
rect 27026 4257 27164 4264
rect 27216 4260 27369 4264
rect 27421 4260 27568 4264
rect 27620 4260 27784 4264
rect 27216 4257 27784 4260
rect 27026 4255 27784 4257
rect 27836 4260 28172 4264
rect 28224 4260 28407 4264
rect 27836 4255 28407 4260
rect 28459 4257 28649 4264
rect 28701 4258 28881 4264
rect 28933 4261 29110 4264
rect 29162 4261 29359 4264
rect 28933 4258 29359 4261
rect 28701 4257 29359 4258
rect 28459 4255 29359 4257
rect 27026 4253 29359 4255
rect 29411 4257 29577 4264
rect 29629 4257 29806 4264
rect 29411 4253 29806 4257
rect 29858 4255 30027 4264
rect 30079 4260 30243 4264
rect 30295 4298 30361 4312
rect 30295 4264 30298 4298
rect 30332 4264 30361 4298
rect 30295 4260 30361 4264
rect 30079 4255 30361 4260
rect 29858 4253 30361 4255
rect 25492 4233 30361 4253
rect 23386 4206 23439 4213
rect 23529 4146 23795 4216
rect 10928 4115 23795 4146
rect 10928 4114 13660 4115
rect 10928 4080 11118 4114
rect 11152 4080 11210 4114
rect 11244 4080 11302 4114
rect 11336 4080 11394 4114
rect 11428 4080 11486 4114
rect 11520 4080 11578 4114
rect 11612 4080 11670 4114
rect 11704 4080 11762 4114
rect 11796 4080 11854 4114
rect 11888 4081 13660 4114
rect 13694 4081 13752 4115
rect 13786 4081 13844 4115
rect 13878 4081 13917 4115
rect 13951 4081 14009 4115
rect 14043 4081 14101 4115
rect 14135 4081 14193 4115
rect 14227 4081 14285 4115
rect 14319 4081 14377 4115
rect 14411 4081 14469 4115
rect 14503 4081 14561 4115
rect 14595 4081 14653 4115
rect 14687 4081 14745 4115
rect 14779 4081 14837 4115
rect 14871 4081 14929 4115
rect 14963 4081 15021 4115
rect 15055 4081 15113 4115
rect 15147 4081 15205 4115
rect 15239 4081 15297 4115
rect 15331 4081 15389 4115
rect 15423 4081 15481 4115
rect 15515 4081 15573 4115
rect 15607 4081 15665 4115
rect 15699 4081 15757 4115
rect 15791 4081 15849 4115
rect 15883 4081 15941 4115
rect 15975 4081 16033 4115
rect 16067 4081 16125 4115
rect 16159 4081 16217 4115
rect 16251 4081 16309 4115
rect 16343 4081 16401 4115
rect 16435 4081 16493 4115
rect 16527 4081 16585 4115
rect 16619 4081 16677 4115
rect 16711 4081 16769 4115
rect 16803 4081 16861 4115
rect 16895 4081 16953 4115
rect 16987 4081 17045 4115
rect 17079 4081 17137 4115
rect 17171 4081 17229 4115
rect 17263 4081 17321 4115
rect 17355 4081 17413 4115
rect 17447 4081 17505 4115
rect 17539 4081 17597 4115
rect 17631 4081 17689 4115
rect 17723 4081 17781 4115
rect 17815 4081 17873 4115
rect 17907 4081 17965 4115
rect 17999 4081 18057 4115
rect 18091 4081 18149 4115
rect 18183 4081 18241 4115
rect 18275 4081 18333 4115
rect 18367 4081 18425 4115
rect 18459 4081 18517 4115
rect 18551 4081 18609 4115
rect 18643 4081 18701 4115
rect 18735 4081 18793 4115
rect 18827 4081 18885 4115
rect 18919 4081 18977 4115
rect 19011 4081 19069 4115
rect 19103 4081 19161 4115
rect 19195 4081 19253 4115
rect 19287 4081 19345 4115
rect 19379 4081 19437 4115
rect 19471 4081 19529 4115
rect 19563 4081 19621 4115
rect 19655 4081 19713 4115
rect 19747 4081 19805 4115
rect 19839 4081 19897 4115
rect 19931 4081 19989 4115
rect 20023 4081 20081 4115
rect 20115 4081 20173 4115
rect 20207 4081 20265 4115
rect 20299 4081 20357 4115
rect 20391 4081 20449 4115
rect 20483 4081 20541 4115
rect 20575 4081 20633 4115
rect 20667 4081 20725 4115
rect 20759 4081 20817 4115
rect 20851 4081 20909 4115
rect 20943 4081 21001 4115
rect 21035 4081 21093 4115
rect 21127 4081 21185 4115
rect 21219 4081 21277 4115
rect 21311 4081 21369 4115
rect 21403 4081 21461 4115
rect 21495 4081 21553 4115
rect 21587 4081 21645 4115
rect 21679 4081 21737 4115
rect 21771 4081 21829 4115
rect 21863 4081 21921 4115
rect 21955 4081 22013 4115
rect 22047 4081 22105 4115
rect 22139 4081 22197 4115
rect 22231 4081 22289 4115
rect 22323 4081 22381 4115
rect 22415 4081 22473 4115
rect 22507 4081 22565 4115
rect 22599 4081 22657 4115
rect 22691 4081 22749 4115
rect 22783 4081 22841 4115
rect 22875 4081 22933 4115
rect 22967 4081 23025 4115
rect 23059 4081 23117 4115
rect 23151 4081 23209 4115
rect 23243 4081 23301 4115
rect 23335 4081 23393 4115
rect 23427 4088 23795 4115
rect 23427 4081 23605 4088
rect 11888 4080 23605 4081
rect 10928 4050 23605 4080
rect 11089 4049 11917 4050
rect 10933 3972 10967 3977
rect 11103 3972 11109 3988
rect 10931 3944 11109 3972
rect 10933 3942 10967 3944
rect 11103 3936 11109 3944
rect 11161 3936 11167 3988
rect 11723 3933 11729 3985
rect 11781 3972 11787 3985
rect 13463 3972 13470 3983
rect 11781 3944 13470 3972
rect 11781 3933 11787 3944
rect 13463 3931 13470 3944
rect 13522 3972 13529 3983
rect 15843 3972 15850 3984
rect 13522 3944 15850 3972
rect 13522 3931 13529 3944
rect 15843 3932 15850 3944
rect 15902 3972 15909 3984
rect 16642 3972 16649 3983
rect 15902 3944 16649 3972
rect 15902 3932 15909 3944
rect 16642 3931 16649 3944
rect 16701 3972 16708 3983
rect 18236 3972 18243 3983
rect 16701 3944 18243 3972
rect 16701 3931 16708 3944
rect 18236 3931 18243 3944
rect 18295 3972 18302 3983
rect 19031 3972 19038 3984
rect 18295 3944 19038 3972
rect 18295 3931 18302 3944
rect 19031 3932 19038 3944
rect 19090 3972 19097 3984
rect 20623 3972 20630 3983
rect 19090 3944 20630 3972
rect 19090 3932 19097 3944
rect 20623 3931 20630 3944
rect 20682 3972 20689 3983
rect 21440 3972 21447 3984
rect 20682 3944 21447 3972
rect 20682 3931 20689 3944
rect 21440 3932 21447 3944
rect 21499 3972 21506 3984
rect 23018 3972 23025 3984
rect 21499 3944 23025 3972
rect 21499 3932 21506 3944
rect 23018 3932 23025 3944
rect 23077 3972 23084 3984
rect 23077 3944 23461 3972
rect 23077 3932 23084 3944
rect 23525 3942 23605 4050
rect 23755 3942 23795 4088
rect 23525 3874 23795 3942
rect 11018 3846 23795 3874
rect 25226 4193 25541 4203
rect 25226 4165 28114 4193
rect 30414 4183 30754 4193
rect 30285 4177 30754 4183
rect 25226 4155 25541 4165
rect 11018 3845 23521 3846
rect 10826 3813 23675 3817
rect 10753 3800 23675 3813
rect 10753 3792 11255 3800
rect 10753 3646 10905 3792
rect 11055 3654 11255 3792
rect 11405 3786 23675 3800
rect 11405 3752 11525 3786
rect 11559 3752 11617 3786
rect 11651 3752 11709 3786
rect 11743 3752 11801 3786
rect 11835 3752 11893 3786
rect 11927 3752 11985 3786
rect 12019 3752 12077 3786
rect 12111 3752 12169 3786
rect 12203 3752 12261 3786
rect 12295 3752 12353 3786
rect 12387 3752 12445 3786
rect 12479 3752 12537 3786
rect 12571 3752 12629 3786
rect 12663 3752 12721 3786
rect 12755 3752 12813 3786
rect 12847 3752 12905 3786
rect 12939 3752 12997 3786
rect 13031 3752 13089 3786
rect 13123 3752 13181 3786
rect 13215 3752 13273 3786
rect 13307 3752 13365 3786
rect 13399 3752 13457 3786
rect 13491 3752 13549 3786
rect 13583 3752 13641 3786
rect 13675 3752 13733 3786
rect 13767 3752 13825 3786
rect 13859 3752 13917 3786
rect 13951 3752 14009 3786
rect 14043 3752 14101 3786
rect 14135 3752 14193 3786
rect 14227 3752 14285 3786
rect 14319 3752 14377 3786
rect 14411 3752 14469 3786
rect 14503 3752 14561 3786
rect 14595 3752 14653 3786
rect 14687 3752 14745 3786
rect 14779 3752 14837 3786
rect 14871 3752 14929 3786
rect 14963 3752 15021 3786
rect 15055 3752 15113 3786
rect 15147 3752 15205 3786
rect 15239 3752 15297 3786
rect 15331 3752 15389 3786
rect 15423 3752 15481 3786
rect 15515 3752 15573 3786
rect 15607 3752 15665 3786
rect 15699 3752 15757 3786
rect 15791 3752 15849 3786
rect 15883 3752 15941 3786
rect 15975 3752 16033 3786
rect 16067 3752 16125 3786
rect 16159 3752 16217 3786
rect 16251 3752 16309 3786
rect 16343 3752 16401 3786
rect 16435 3752 16493 3786
rect 16527 3752 16585 3786
rect 16619 3752 16677 3786
rect 16711 3752 16769 3786
rect 16803 3752 16861 3786
rect 16895 3752 16953 3786
rect 16987 3752 17045 3786
rect 17079 3752 17137 3786
rect 17171 3752 17229 3786
rect 17263 3752 17321 3786
rect 17355 3752 17413 3786
rect 17447 3752 17505 3786
rect 17539 3752 17597 3786
rect 17631 3752 17689 3786
rect 17723 3752 17781 3786
rect 17815 3752 17873 3786
rect 17907 3752 17965 3786
rect 17999 3752 18057 3786
rect 18091 3752 18149 3786
rect 18183 3752 18241 3786
rect 18275 3752 18333 3786
rect 18367 3752 18425 3786
rect 18459 3752 18517 3786
rect 18551 3752 18609 3786
rect 18643 3752 18701 3786
rect 18735 3752 18793 3786
rect 18827 3752 18885 3786
rect 18919 3752 18977 3786
rect 19011 3752 19069 3786
rect 19103 3752 19161 3786
rect 19195 3752 19253 3786
rect 19287 3752 19345 3786
rect 19379 3752 19437 3786
rect 19471 3752 19529 3786
rect 19563 3752 19621 3786
rect 19655 3752 19713 3786
rect 19747 3752 19805 3786
rect 19839 3752 19897 3786
rect 19931 3752 19989 3786
rect 20023 3752 20081 3786
rect 20115 3752 20173 3786
rect 20207 3752 20265 3786
rect 20299 3752 20357 3786
rect 20391 3752 20449 3786
rect 20483 3752 20541 3786
rect 20575 3752 20633 3786
rect 20667 3752 20725 3786
rect 20759 3752 20817 3786
rect 20851 3752 20909 3786
rect 20943 3752 21001 3786
rect 21035 3752 21093 3786
rect 21127 3752 21185 3786
rect 21219 3752 21277 3786
rect 21311 3752 21369 3786
rect 21403 3752 21461 3786
rect 21495 3752 21553 3786
rect 21587 3752 21645 3786
rect 21679 3752 21737 3786
rect 21771 3752 21829 3786
rect 21863 3752 21921 3786
rect 21955 3752 22013 3786
rect 22047 3752 22105 3786
rect 22139 3752 22197 3786
rect 22231 3752 22289 3786
rect 22323 3752 22381 3786
rect 22415 3752 22473 3786
rect 22507 3752 22565 3786
rect 22599 3752 22657 3786
rect 22691 3752 22749 3786
rect 22783 3752 22841 3786
rect 22875 3752 22933 3786
rect 22967 3752 23025 3786
rect 23059 3752 23117 3786
rect 23151 3752 23209 3786
rect 23243 3752 23301 3786
rect 23335 3752 23393 3786
rect 23427 3752 23675 3786
rect 11405 3721 23675 3752
rect 11405 3654 11437 3721
rect 11055 3646 11437 3654
rect 10753 3372 11437 3646
rect 12616 3616 12674 3622
rect 12616 3582 12628 3616
rect 12662 3613 12674 3616
rect 13352 3616 13410 3622
rect 13352 3613 13364 3616
rect 12662 3585 13364 3613
rect 12662 3582 12674 3585
rect 12616 3576 12674 3582
rect 13352 3582 13364 3585
rect 13398 3613 13410 3616
rect 13720 3616 13778 3622
rect 13720 3613 13732 3616
rect 13398 3585 13732 3613
rect 13398 3582 13410 3585
rect 13352 3576 13410 3582
rect 13720 3582 13732 3585
rect 13766 3582 13778 3616
rect 13720 3576 13778 3582
rect 15008 3616 15066 3622
rect 15008 3582 15020 3616
rect 15054 3613 15066 3616
rect 15744 3616 15802 3622
rect 15744 3613 15756 3616
rect 15054 3585 15756 3613
rect 15054 3582 15066 3585
rect 15008 3576 15066 3582
rect 15744 3582 15756 3585
rect 15790 3613 15802 3616
rect 16112 3616 16170 3622
rect 16112 3613 16124 3616
rect 15790 3585 16124 3613
rect 15790 3582 15802 3585
rect 15744 3576 15802 3582
rect 16112 3582 16124 3585
rect 16158 3582 16170 3616
rect 16112 3576 16170 3582
rect 17400 3616 17458 3622
rect 17400 3582 17412 3616
rect 17446 3613 17458 3616
rect 18136 3616 18194 3622
rect 18136 3613 18148 3616
rect 17446 3585 18148 3613
rect 17446 3582 17458 3585
rect 17400 3576 17458 3582
rect 18136 3582 18148 3585
rect 18182 3613 18194 3616
rect 18504 3616 18562 3622
rect 18504 3613 18516 3616
rect 18182 3585 18516 3613
rect 18182 3582 18194 3585
rect 18136 3576 18194 3582
rect 18504 3582 18516 3585
rect 18550 3582 18562 3616
rect 18504 3576 18562 3582
rect 19792 3616 19850 3622
rect 19792 3582 19804 3616
rect 19838 3613 19850 3616
rect 20528 3616 20586 3622
rect 20528 3613 20540 3616
rect 19838 3585 20540 3613
rect 19838 3582 19850 3585
rect 19792 3576 19850 3582
rect 20528 3582 20540 3585
rect 20574 3613 20586 3616
rect 20896 3616 20954 3622
rect 20896 3613 20908 3616
rect 20574 3585 20908 3613
rect 20574 3582 20586 3585
rect 20528 3576 20586 3582
rect 20896 3582 20908 3585
rect 20942 3582 20954 3616
rect 20896 3576 20954 3582
rect 22184 3616 22242 3622
rect 22184 3582 22196 3616
rect 22230 3613 22242 3616
rect 22920 3616 22978 3622
rect 22920 3613 22932 3616
rect 22230 3585 22932 3613
rect 22230 3582 22242 3585
rect 22184 3576 22242 3582
rect 22920 3582 22932 3585
rect 22966 3613 22978 3616
rect 23288 3616 23346 3622
rect 23288 3613 23300 3616
rect 22966 3585 23300 3613
rect 22966 3582 22978 3585
rect 22920 3576 22978 3582
rect 23288 3582 23300 3585
rect 23334 3582 23346 3616
rect 23288 3576 23346 3582
rect 12064 3548 12122 3554
rect 12064 3514 12076 3548
rect 12110 3545 12122 3548
rect 12708 3548 12766 3554
rect 12708 3545 12720 3548
rect 12110 3517 12720 3545
rect 12110 3514 12122 3517
rect 12064 3508 12122 3514
rect 12708 3514 12720 3517
rect 12754 3514 12766 3548
rect 14456 3548 14514 3554
rect 12708 3508 12766 3514
rect 13462 3494 13469 3546
rect 13521 3494 13528 3546
rect 14456 3514 14468 3548
rect 14502 3545 14514 3548
rect 15100 3548 15158 3554
rect 15100 3545 15112 3548
rect 14502 3517 15112 3545
rect 14502 3514 14514 3517
rect 14456 3508 14514 3514
rect 15100 3514 15112 3517
rect 15146 3514 15158 3548
rect 16848 3548 16906 3554
rect 15100 3508 15158 3514
rect 14350 3494 14403 3501
rect 11951 3436 11961 3488
rect 12013 3436 12025 3488
rect 12616 3480 12674 3486
rect 12616 3446 12628 3480
rect 12662 3477 12674 3480
rect 12662 3449 13303 3477
rect 12662 3446 12674 3449
rect 12616 3440 12674 3446
rect 11951 3434 12025 3436
rect 13075 3420 13141 3421
rect 12340 3412 12398 3418
rect 12340 3378 12352 3412
rect 12386 3409 12398 3412
rect 13075 3409 13082 3420
rect 12386 3381 13082 3409
rect 12386 3378 12398 3381
rect 12340 3372 12398 3378
rect 13075 3368 13082 3381
rect 13134 3368 13141 3420
rect 13264 3418 13303 3449
rect 14350 3442 14351 3494
rect 15843 3491 15850 3543
rect 15902 3491 15909 3543
rect 16848 3514 16860 3548
rect 16894 3545 16906 3548
rect 17492 3548 17550 3554
rect 17492 3545 17504 3548
rect 16894 3517 17504 3545
rect 16894 3514 16906 3517
rect 16848 3508 16906 3514
rect 17492 3514 17504 3517
rect 17538 3514 17550 3548
rect 19240 3548 19298 3554
rect 17492 3508 17550 3514
rect 16744 3492 16797 3499
rect 18234 3495 18241 3547
rect 18293 3495 18300 3547
rect 19240 3514 19252 3548
rect 19286 3545 19298 3548
rect 19884 3548 19942 3554
rect 21632 3548 21690 3554
rect 19884 3545 19896 3548
rect 19286 3517 19896 3545
rect 19286 3514 19298 3517
rect 19240 3508 19298 3514
rect 19884 3514 19896 3517
rect 19930 3514 19942 3548
rect 19884 3508 19942 3514
rect 14350 3435 14403 3442
rect 15008 3480 15066 3486
rect 15008 3446 15020 3480
rect 15054 3477 15066 3480
rect 15054 3449 15695 3477
rect 15054 3446 15066 3449
rect 15008 3440 15066 3446
rect 15656 3418 15695 3449
rect 16796 3440 16797 3492
rect 19136 3493 19189 3500
rect 20623 3496 20630 3548
rect 20682 3496 20689 3548
rect 21632 3514 21644 3548
rect 21678 3545 21690 3548
rect 22276 3548 22334 3554
rect 22276 3545 22288 3548
rect 21678 3517 22288 3545
rect 21678 3514 21690 3517
rect 21632 3508 21690 3514
rect 22276 3514 22288 3517
rect 22322 3514 22334 3548
rect 22276 3508 22334 3514
rect 17400 3480 17458 3486
rect 17400 3446 17412 3480
rect 17446 3477 17458 3480
rect 17446 3449 18087 3477
rect 17446 3446 17458 3449
rect 17400 3440 17458 3446
rect 16744 3433 16797 3440
rect 18048 3418 18087 3449
rect 19188 3441 19189 3493
rect 21529 3494 21582 3501
rect 23017 3496 23024 3548
rect 23076 3496 23083 3548
rect 23382 3501 23434 3503
rect 23379 3497 23436 3501
rect 19136 3434 19189 3441
rect 19792 3480 19850 3486
rect 19792 3446 19804 3480
rect 19838 3477 19850 3480
rect 19838 3449 20479 3477
rect 19838 3446 19850 3449
rect 19792 3440 19850 3446
rect 20440 3418 20479 3449
rect 21581 3442 21582 3494
rect 21529 3435 21582 3442
rect 22184 3480 22242 3486
rect 22184 3446 22196 3480
rect 22230 3477 22242 3480
rect 22230 3449 22871 3477
rect 22230 3446 22242 3449
rect 22184 3440 22242 3446
rect 22832 3418 22871 3449
rect 23379 3445 23382 3497
rect 23434 3445 23436 3497
rect 23379 3442 23436 3445
rect 23382 3439 23434 3442
rect 13264 3412 13322 3418
rect 13264 3378 13276 3412
rect 13310 3409 13322 3412
rect 13628 3412 13686 3418
rect 13628 3409 13640 3412
rect 13310 3381 13640 3409
rect 13310 3378 13322 3381
rect 13264 3372 13322 3378
rect 13628 3378 13640 3381
rect 13674 3378 13686 3412
rect 14732 3412 14790 3418
rect 13628 3372 13686 3378
rect 13905 3384 13958 3391
rect 11514 3361 11567 3368
rect 11566 3309 11567 3361
rect 13957 3332 13958 3384
rect 14732 3378 14744 3412
rect 14778 3409 14790 3412
rect 15468 3412 15526 3418
rect 15468 3409 15480 3412
rect 14778 3381 15480 3409
rect 14778 3378 14790 3381
rect 14732 3372 14790 3378
rect 15468 3378 15480 3381
rect 15514 3378 15526 3412
rect 15468 3372 15526 3378
rect 15656 3412 15714 3418
rect 15656 3378 15668 3412
rect 15702 3409 15714 3412
rect 16020 3412 16078 3418
rect 16020 3409 16032 3412
rect 15702 3381 16032 3409
rect 15702 3378 15714 3381
rect 15656 3372 15714 3378
rect 16020 3378 16032 3381
rect 16066 3378 16078 3412
rect 17124 3412 17182 3418
rect 16020 3372 16078 3378
rect 16296 3383 16349 3390
rect 13905 3325 13958 3332
rect 15480 3344 15514 3372
rect 15923 3344 15929 3353
rect 15480 3316 15929 3344
rect 11514 3302 11567 3309
rect 15923 3301 15929 3316
rect 15981 3301 15987 3353
rect 16348 3331 16349 3383
rect 17124 3378 17136 3412
rect 17170 3409 17182 3412
rect 17860 3412 17918 3418
rect 17860 3409 17872 3412
rect 17170 3381 17872 3409
rect 17170 3378 17182 3381
rect 17124 3372 17182 3378
rect 17860 3378 17872 3381
rect 17906 3378 17918 3412
rect 17860 3372 17918 3378
rect 18048 3412 18106 3418
rect 18048 3378 18060 3412
rect 18094 3409 18106 3412
rect 18412 3412 18470 3418
rect 18412 3409 18424 3412
rect 18094 3381 18424 3409
rect 18094 3378 18106 3381
rect 18048 3372 18106 3378
rect 18412 3378 18424 3381
rect 18458 3378 18470 3412
rect 19516 3412 19574 3418
rect 18412 3372 18470 3378
rect 18691 3386 18744 3393
rect 16296 3324 16349 3331
rect 17872 3344 17906 3372
rect 18315 3344 18321 3353
rect 17872 3316 18321 3344
rect 18315 3301 18321 3316
rect 18373 3301 18379 3353
rect 18743 3334 18744 3386
rect 19516 3378 19528 3412
rect 19562 3409 19574 3412
rect 20252 3412 20310 3418
rect 20252 3409 20264 3412
rect 19562 3381 20264 3409
rect 19562 3378 19574 3381
rect 19516 3372 19574 3378
rect 20252 3378 20264 3381
rect 20298 3378 20310 3412
rect 20252 3372 20310 3378
rect 20440 3412 20498 3418
rect 20440 3378 20452 3412
rect 20486 3409 20498 3412
rect 20804 3412 20862 3418
rect 20804 3409 20816 3412
rect 20486 3381 20816 3409
rect 20486 3378 20498 3381
rect 20440 3372 20498 3378
rect 20804 3378 20816 3381
rect 20850 3378 20862 3412
rect 21908 3412 21966 3418
rect 20804 3372 20862 3378
rect 21080 3384 21133 3391
rect 18691 3327 18744 3334
rect 20264 3344 20298 3372
rect 20707 3344 20713 3353
rect 20264 3316 20713 3344
rect 20707 3301 20713 3316
rect 20765 3301 20771 3353
rect 21132 3332 21133 3384
rect 21908 3378 21920 3412
rect 21954 3409 21966 3412
rect 22644 3412 22702 3418
rect 22644 3409 22656 3412
rect 21954 3381 22656 3409
rect 21954 3378 21966 3381
rect 21908 3372 21966 3378
rect 22644 3378 22656 3381
rect 22690 3378 22702 3412
rect 22644 3372 22702 3378
rect 22832 3412 22890 3418
rect 22832 3378 22844 3412
rect 22878 3409 22890 3412
rect 23196 3412 23254 3418
rect 23196 3409 23208 3412
rect 22878 3381 23208 3409
rect 22878 3378 22890 3381
rect 22832 3372 22890 3378
rect 23196 3378 23208 3381
rect 23242 3378 23254 3412
rect 23196 3372 23254 3378
rect 23535 3410 23795 3572
rect 21080 3325 21133 3332
rect 22656 3344 22690 3372
rect 23098 3344 23104 3353
rect 22656 3316 23104 3344
rect 23098 3301 23104 3316
rect 23156 3301 23162 3353
rect 23535 3273 23611 3410
rect 10853 3264 23611 3273
rect 23761 3264 23795 3410
rect 10853 3242 23795 3264
rect 10853 3208 11525 3242
rect 11559 3208 11617 3242
rect 11651 3208 11709 3242
rect 11743 3208 11801 3242
rect 11835 3208 11893 3242
rect 11927 3208 11985 3242
rect 12019 3208 12077 3242
rect 12111 3208 12169 3242
rect 12203 3208 12261 3242
rect 12295 3208 12353 3242
rect 12387 3208 12445 3242
rect 12479 3208 12537 3242
rect 12571 3208 12629 3242
rect 12663 3208 12721 3242
rect 12755 3208 12813 3242
rect 12847 3208 12905 3242
rect 12939 3208 12997 3242
rect 13031 3208 13089 3242
rect 13123 3208 13181 3242
rect 13215 3208 13273 3242
rect 13307 3208 13365 3242
rect 13399 3208 13457 3242
rect 13491 3208 13549 3242
rect 13583 3208 13641 3242
rect 13675 3208 13733 3242
rect 13767 3208 13825 3242
rect 13859 3208 13917 3242
rect 13951 3208 14009 3242
rect 14043 3208 14101 3242
rect 14135 3208 14193 3242
rect 14227 3208 14285 3242
rect 14319 3208 14377 3242
rect 14411 3208 14469 3242
rect 14503 3208 14561 3242
rect 14595 3208 14653 3242
rect 14687 3208 14745 3242
rect 14779 3208 14837 3242
rect 14871 3208 14929 3242
rect 14963 3208 15021 3242
rect 15055 3208 15113 3242
rect 15147 3208 15205 3242
rect 15239 3208 15297 3242
rect 15331 3208 15389 3242
rect 15423 3208 15481 3242
rect 15515 3208 15573 3242
rect 15607 3208 15665 3242
rect 15699 3208 15757 3242
rect 15791 3208 15849 3242
rect 15883 3208 15941 3242
rect 15975 3208 16033 3242
rect 16067 3208 16125 3242
rect 16159 3208 16217 3242
rect 16251 3208 16309 3242
rect 16343 3208 16401 3242
rect 16435 3208 16493 3242
rect 16527 3208 16585 3242
rect 16619 3208 16677 3242
rect 16711 3208 16769 3242
rect 16803 3208 16861 3242
rect 16895 3208 16953 3242
rect 16987 3208 17045 3242
rect 17079 3208 17137 3242
rect 17171 3208 17229 3242
rect 17263 3208 17321 3242
rect 17355 3208 17413 3242
rect 17447 3208 17505 3242
rect 17539 3208 17597 3242
rect 17631 3208 17689 3242
rect 17723 3208 17781 3242
rect 17815 3208 17873 3242
rect 17907 3208 17965 3242
rect 17999 3208 18057 3242
rect 18091 3208 18149 3242
rect 18183 3208 18241 3242
rect 18275 3208 18333 3242
rect 18367 3208 18425 3242
rect 18459 3208 18517 3242
rect 18551 3208 18609 3242
rect 18643 3208 18701 3242
rect 18735 3208 18793 3242
rect 18827 3208 18885 3242
rect 18919 3208 18977 3242
rect 19011 3208 19069 3242
rect 19103 3208 19161 3242
rect 19195 3208 19253 3242
rect 19287 3208 19345 3242
rect 19379 3208 19437 3242
rect 19471 3208 19529 3242
rect 19563 3208 19621 3242
rect 19655 3208 19713 3242
rect 19747 3208 19805 3242
rect 19839 3208 19897 3242
rect 19931 3208 19989 3242
rect 20023 3208 20081 3242
rect 20115 3208 20173 3242
rect 20207 3208 20265 3242
rect 20299 3208 20357 3242
rect 20391 3208 20449 3242
rect 20483 3208 20541 3242
rect 20575 3208 20633 3242
rect 20667 3208 20725 3242
rect 20759 3208 20817 3242
rect 20851 3208 20909 3242
rect 20943 3208 21001 3242
rect 21035 3208 21093 3242
rect 21127 3208 21185 3242
rect 21219 3208 21277 3242
rect 21311 3208 21369 3242
rect 21403 3208 21461 3242
rect 21495 3208 21553 3242
rect 21587 3208 21645 3242
rect 21679 3208 21737 3242
rect 21771 3208 21829 3242
rect 21863 3208 21921 3242
rect 21955 3208 22013 3242
rect 22047 3208 22105 3242
rect 22139 3208 22197 3242
rect 22231 3208 22289 3242
rect 22323 3208 22381 3242
rect 22415 3208 22473 3242
rect 22507 3208 22565 3242
rect 22599 3208 22657 3242
rect 22691 3208 22749 3242
rect 22783 3208 22841 3242
rect 22875 3208 22933 3242
rect 22967 3208 23025 3242
rect 23059 3208 23117 3242
rect 23151 3208 23209 3242
rect 23243 3208 23301 3242
rect 23335 3208 23393 3242
rect 23427 3208 23795 3242
rect 10853 3177 23795 3208
rect 23535 3176 23795 3177
rect 14907 3096 14914 3148
rect 14966 3143 14972 3148
rect 20834 3143 20840 3149
rect 14966 3115 20840 3143
rect 14966 3096 14972 3115
rect 20834 3097 20840 3115
rect 20892 3097 20898 3149
rect 20996 3097 21002 3149
rect 21054 3142 21060 3149
rect 24881 3142 24887 3155
rect 21054 3114 24887 3142
rect 21054 3097 21060 3114
rect 24881 3103 24887 3114
rect 24940 3142 24946 3155
rect 25226 3142 25254 4155
rect 25779 4128 25837 4134
rect 25779 4094 25791 4128
rect 25825 4125 25837 4128
rect 26143 4128 26201 4134
rect 26143 4125 26155 4128
rect 25825 4097 26155 4125
rect 25825 4094 25837 4097
rect 25779 4088 25837 4094
rect 26143 4094 26155 4097
rect 26189 4094 26201 4128
rect 26143 4088 26201 4094
rect 26331 4128 26389 4134
rect 26331 4094 26343 4128
rect 26377 4125 26389 4128
rect 27067 4128 27125 4134
rect 27067 4125 27079 4128
rect 26377 4119 27079 4125
rect 27113 4119 27125 4128
rect 26377 4097 27072 4119
rect 26377 4094 26389 4097
rect 26331 4088 26389 4094
rect 25613 4081 25665 4087
rect 26162 4057 26201 4088
rect 27065 4067 27072 4097
rect 27124 4067 27131 4119
rect 26791 4060 26849 4066
rect 26791 4057 26803 4060
rect 26162 4029 26803 4057
rect 25613 4023 25665 4029
rect 26791 4026 26803 4029
rect 26837 4026 26849 4060
rect 26791 4020 26849 4026
rect 27450 4016 27457 4068
rect 27509 4016 27516 4068
rect 28085 4059 28113 4165
rect 30285 4143 30298 4177
rect 30332 4154 30754 4177
rect 30332 4143 30344 4154
rect 30414 4145 30754 4154
rect 30285 4137 30344 4143
rect 28171 4128 28229 4134
rect 28171 4094 28183 4128
rect 28217 4125 28229 4128
rect 28535 4128 28593 4134
rect 28535 4125 28547 4128
rect 28217 4097 28547 4125
rect 28217 4094 28229 4097
rect 28171 4088 28229 4094
rect 28535 4094 28547 4097
rect 28581 4094 28593 4128
rect 28535 4088 28593 4094
rect 28723 4128 28781 4134
rect 28723 4094 28735 4128
rect 28769 4125 28781 4128
rect 29459 4128 29517 4134
rect 29459 4125 29471 4128
rect 28769 4118 29471 4125
rect 29505 4118 29517 4128
rect 28769 4097 29467 4118
rect 28769 4094 28781 4097
rect 28723 4088 28781 4094
rect 29459 4088 29467 4097
rect 28327 4060 28394 4069
rect 28327 4059 28345 4060
rect 28005 4039 28057 4045
rect 28085 4031 28345 4059
rect 24940 3114 25254 3142
rect 25282 3997 25525 3999
rect 25928 3998 25989 4004
rect 25282 3986 25549 3997
rect 25928 3986 25943 3998
rect 25282 3964 25943 3986
rect 25977 3964 25989 3998
rect 25282 3958 25989 3964
rect 26699 3992 26757 3998
rect 26699 3958 26711 3992
rect 26745 3989 26757 3992
rect 27343 3992 27401 3998
rect 27343 3989 27355 3992
rect 26745 3961 27355 3989
rect 26745 3958 26757 3961
rect 25282 3951 25549 3958
rect 26699 3952 26757 3958
rect 27343 3958 27355 3961
rect 27389 3958 27401 3992
rect 28327 4026 28345 4031
rect 28379 4026 28394 4060
rect 28554 4057 28593 4088
rect 29460 4066 29467 4088
rect 29519 4066 29526 4118
rect 29183 4060 29241 4066
rect 29183 4057 29195 4060
rect 28554 4029 29195 4057
rect 28327 4018 28394 4026
rect 29183 4026 29195 4029
rect 29229 4026 29241 4060
rect 29183 4020 29241 4026
rect 29845 4017 29852 4069
rect 29904 4017 29911 4069
rect 28005 3981 28057 3987
rect 29091 3992 29149 3998
rect 27343 3952 27401 3958
rect 29091 3958 29103 3992
rect 29137 3989 29149 3992
rect 29735 3992 29793 3998
rect 29735 3989 29747 3992
rect 29137 3961 29747 3989
rect 29137 3958 29149 3961
rect 29091 3952 29149 3958
rect 29735 3958 29747 3961
rect 29781 3958 29793 3992
rect 29735 3952 29793 3958
rect 24940 3103 24946 3114
rect 18599 3018 18605 3086
rect 18657 3069 18663 3086
rect 25282 3069 25310 3951
rect 25504 3949 25549 3951
rect 25687 3924 25745 3930
rect 25687 3890 25699 3924
rect 25733 3921 25745 3924
rect 26055 3924 26113 3930
rect 26055 3921 26067 3924
rect 25733 3893 26067 3921
rect 25733 3890 25745 3893
rect 25687 3884 25745 3890
rect 26055 3890 26067 3893
rect 26101 3921 26113 3924
rect 26791 3924 26849 3930
rect 26791 3921 26803 3924
rect 26101 3893 26803 3921
rect 26101 3890 26113 3893
rect 26055 3884 26113 3890
rect 26791 3890 26803 3893
rect 26837 3890 26849 3924
rect 26791 3884 26849 3890
rect 28079 3924 28137 3930
rect 28079 3890 28091 3924
rect 28125 3921 28137 3924
rect 28447 3924 28505 3930
rect 28447 3921 28459 3924
rect 28125 3893 28459 3921
rect 28125 3890 28137 3893
rect 28079 3884 28137 3890
rect 28447 3890 28459 3893
rect 28493 3921 28505 3924
rect 29183 3924 29241 3930
rect 29183 3921 29195 3924
rect 28493 3893 29195 3921
rect 28493 3890 28505 3893
rect 28447 3884 28505 3890
rect 29183 3890 29195 3893
rect 29229 3890 29241 3924
rect 29183 3884 29241 3890
rect 27898 3860 27956 3867
rect 27898 3826 27910 3860
rect 27944 3853 27956 3860
rect 30414 3853 30764 3863
rect 27944 3826 30764 3853
rect 27898 3825 30764 3826
rect 27898 3819 27956 3825
rect 30414 3815 30764 3825
rect 25577 3754 30361 3785
rect 25577 3720 25606 3754
rect 25640 3720 25698 3754
rect 25732 3723 25790 3754
rect 25768 3720 25790 3723
rect 25824 3720 25882 3754
rect 25916 3721 25974 3754
rect 25943 3720 25974 3721
rect 26008 3720 26066 3754
rect 26100 3723 26158 3754
rect 26140 3720 26158 3723
rect 26192 3720 26250 3754
rect 26284 3726 26342 3754
rect 26284 3720 26307 3726
rect 26376 3720 26434 3754
rect 26468 3720 26526 3754
rect 26560 3722 26618 3754
rect 26591 3720 26618 3722
rect 26652 3720 26710 3754
rect 26744 3729 26802 3754
rect 26744 3720 26763 3729
rect 26836 3720 26894 3754
rect 26928 3720 26986 3754
rect 27020 3720 27078 3754
rect 27112 3720 27170 3754
rect 27204 3720 27262 3754
rect 27296 3720 27354 3754
rect 27388 3720 27446 3754
rect 27480 3720 27538 3754
rect 27572 3720 27630 3754
rect 27664 3720 27722 3754
rect 27756 3720 27814 3754
rect 27848 3720 27906 3754
rect 27940 3720 27998 3754
rect 28032 3720 28090 3754
rect 28124 3720 28182 3754
rect 28216 3720 28274 3754
rect 28308 3720 28366 3754
rect 28400 3720 28458 3754
rect 28492 3720 28550 3754
rect 28584 3720 28642 3754
rect 28676 3720 28734 3754
rect 28768 3720 28826 3754
rect 28860 3720 28918 3754
rect 28952 3720 29010 3754
rect 29044 3720 29102 3754
rect 29136 3720 29194 3754
rect 29228 3720 29286 3754
rect 29320 3720 29378 3754
rect 29412 3720 29470 3754
rect 29504 3720 29562 3754
rect 29596 3720 29654 3754
rect 29688 3720 29746 3754
rect 29780 3720 29838 3754
rect 29872 3720 29930 3754
rect 29964 3720 30022 3754
rect 30056 3720 30114 3754
rect 30148 3720 30206 3754
rect 30240 3720 30298 3754
rect 30332 3720 30361 3754
rect 25577 3671 25716 3720
rect 25768 3671 25891 3720
rect 25577 3669 25891 3671
rect 25943 3671 26088 3720
rect 26140 3674 26307 3720
rect 26359 3674 26539 3720
rect 26140 3671 26539 3674
rect 25943 3670 26539 3671
rect 26591 3677 26763 3720
rect 26815 3719 30192 3720
rect 26815 3717 29970 3719
rect 26815 3677 26975 3717
rect 26591 3670 26975 3677
rect 25943 3669 26975 3670
rect 25577 3665 26975 3669
rect 27027 3713 29970 3717
rect 27027 3665 27197 3713
rect 25577 3661 27197 3665
rect 27249 3712 29970 3713
rect 27249 3710 28934 3712
rect 27249 3661 27420 3710
rect 25577 3658 27420 3661
rect 27472 3658 27630 3710
rect 27682 3658 27843 3710
rect 27895 3708 28934 3710
rect 27895 3707 28742 3708
rect 27895 3706 28563 3707
rect 27895 3703 28362 3706
rect 27895 3658 28160 3703
rect 28212 3658 28362 3703
rect 28414 3658 28563 3706
rect 28615 3658 28742 3707
rect 28794 3660 28934 3708
rect 28986 3710 29762 3712
rect 28986 3709 29556 3710
rect 28986 3660 29119 3709
rect 28794 3658 29119 3660
rect 29171 3708 29556 3709
rect 29171 3658 29351 3708
rect 29403 3658 29556 3708
rect 29608 3660 29762 3710
rect 29814 3709 29970 3712
rect 29814 3660 29862 3709
rect 29608 3658 29862 3660
rect 29914 3667 29970 3709
rect 30022 3668 30192 3719
rect 30244 3668 30361 3720
rect 30022 3667 30361 3668
rect 29914 3658 30361 3667
rect 25577 3624 25606 3658
rect 25640 3624 25698 3658
rect 25732 3624 25790 3658
rect 25824 3624 25882 3658
rect 25916 3624 25974 3658
rect 26008 3624 26066 3658
rect 26100 3624 26158 3658
rect 26192 3624 26250 3658
rect 26284 3624 26342 3658
rect 26376 3624 26434 3658
rect 26468 3624 26526 3658
rect 26560 3624 26618 3658
rect 26652 3624 26710 3658
rect 26744 3624 26802 3658
rect 26836 3624 26894 3658
rect 26928 3624 26986 3658
rect 27020 3624 27078 3658
rect 27112 3624 27170 3658
rect 27204 3624 27262 3658
rect 27296 3624 27354 3658
rect 27388 3624 27446 3658
rect 27480 3624 27538 3658
rect 27572 3624 27630 3658
rect 27664 3624 27722 3658
rect 27756 3624 27814 3658
rect 27848 3624 27906 3658
rect 27940 3624 27998 3658
rect 28032 3624 28090 3658
rect 28124 3651 28160 3658
rect 28124 3624 28182 3651
rect 28216 3624 28274 3658
rect 28308 3654 28362 3658
rect 28414 3654 28458 3658
rect 28308 3624 28366 3654
rect 28400 3624 28458 3654
rect 28492 3624 28550 3658
rect 28615 3655 28642 3658
rect 28584 3624 28642 3655
rect 28676 3624 28734 3658
rect 28794 3656 28826 3658
rect 28768 3624 28826 3656
rect 28860 3624 28918 3658
rect 28952 3624 29010 3658
rect 29044 3624 29102 3658
rect 29171 3657 29194 3658
rect 29136 3624 29194 3657
rect 29228 3624 29286 3658
rect 29320 3656 29351 3658
rect 29320 3624 29378 3656
rect 29412 3624 29470 3658
rect 29504 3624 29562 3658
rect 29596 3624 29654 3658
rect 29688 3624 29746 3658
rect 29780 3624 29838 3658
rect 29914 3657 29930 3658
rect 29872 3624 29930 3657
rect 29964 3624 30022 3658
rect 30056 3624 30114 3658
rect 30148 3624 30206 3658
rect 30240 3624 30298 3658
rect 30332 3624 30361 3658
rect 25577 3593 30361 3624
rect 30414 3554 30756 3564
rect 27896 3548 30756 3554
rect 27896 3514 27909 3548
rect 27943 3526 30756 3548
rect 27943 3514 27957 3526
rect 30414 3516 30756 3526
rect 27896 3507 27957 3514
rect 25687 3488 25745 3494
rect 25687 3454 25699 3488
rect 25733 3485 25745 3488
rect 26055 3488 26113 3494
rect 26055 3485 26067 3488
rect 25733 3457 26067 3485
rect 25733 3454 25745 3457
rect 25687 3448 25745 3454
rect 26055 3454 26067 3457
rect 26101 3485 26113 3488
rect 26791 3488 26849 3494
rect 26791 3485 26803 3488
rect 26101 3457 26803 3485
rect 26101 3454 26113 3457
rect 26055 3448 26113 3454
rect 26791 3454 26803 3457
rect 26837 3454 26849 3488
rect 26791 3448 26849 3454
rect 28079 3488 28137 3494
rect 28079 3454 28091 3488
rect 28125 3485 28137 3488
rect 28447 3488 28505 3494
rect 28447 3485 28459 3488
rect 28125 3457 28459 3485
rect 28125 3454 28137 3457
rect 28079 3448 28137 3454
rect 28447 3454 28459 3457
rect 28493 3485 28505 3488
rect 29183 3488 29241 3494
rect 29183 3485 29195 3488
rect 28493 3457 29195 3485
rect 28493 3454 28505 3457
rect 28447 3448 28505 3454
rect 29183 3454 29195 3457
rect 29229 3454 29241 3488
rect 29183 3448 29241 3454
rect 25608 3432 25660 3438
rect 26699 3420 26757 3426
rect 26699 3386 26711 3420
rect 26745 3417 26757 3420
rect 27343 3420 27401 3426
rect 27343 3417 27355 3420
rect 26745 3389 27355 3417
rect 26745 3386 26757 3389
rect 26699 3380 26757 3386
rect 27343 3386 27355 3389
rect 27389 3386 27401 3420
rect 29091 3420 29149 3426
rect 27343 3380 27401 3386
rect 28004 3390 28056 3396
rect 25608 3374 25660 3380
rect 29091 3386 29103 3420
rect 29137 3417 29149 3420
rect 29735 3420 29793 3426
rect 29735 3417 29747 3420
rect 29137 3389 29747 3417
rect 29137 3386 29149 3389
rect 29091 3380 29149 3386
rect 29735 3386 29747 3389
rect 29781 3386 29793 3420
rect 29735 3380 29793 3386
rect 18657 3041 25310 3069
rect 25338 3346 25559 3356
rect 25930 3352 25997 3361
rect 25930 3346 25948 3352
rect 25338 3318 25948 3346
rect 25982 3318 25997 3352
rect 26791 3352 26849 3358
rect 26791 3349 26803 3352
rect 25338 3308 25559 3318
rect 25930 3310 25997 3318
rect 26162 3321 26803 3349
rect 18657 3018 18663 3041
rect 9983 2924 9989 2976
rect 10041 2965 10047 2976
rect 11905 2965 11911 2978
rect 10041 2937 11911 2965
rect 10041 2924 10047 2937
rect 11905 2926 11911 2937
rect 11963 2926 11969 2978
rect 19695 2961 19701 3013
rect 19753 3003 19759 3013
rect 21245 3003 21251 3013
rect 19753 2975 21251 3003
rect 19753 2961 19759 2975
rect 21245 2961 21251 2975
rect 21303 2961 21309 3013
rect 22486 2961 22493 3013
rect 22545 3003 22551 3013
rect 23380 3003 23386 3013
rect 22545 2975 23386 3003
rect 22545 2961 22551 2975
rect 23380 2961 23386 2975
rect 23438 3003 23444 3013
rect 25338 3003 25366 3308
rect 26162 3290 26201 3321
rect 26791 3318 26803 3321
rect 26837 3318 26849 3352
rect 26791 3312 26849 3318
rect 27449 3305 27455 3357
rect 27507 3305 27513 3357
rect 28328 3351 28395 3360
rect 28328 3346 28346 3351
rect 28004 3332 28056 3338
rect 28092 3318 28346 3346
rect 25779 3284 25837 3290
rect 25779 3250 25791 3284
rect 25825 3281 25837 3284
rect 26143 3284 26201 3290
rect 26143 3281 26155 3284
rect 25825 3253 26155 3281
rect 25825 3250 25837 3253
rect 25779 3244 25837 3250
rect 26143 3250 26155 3253
rect 26189 3250 26201 3284
rect 26143 3244 26201 3250
rect 26331 3284 26389 3290
rect 26331 3250 26343 3284
rect 26377 3281 26389 3284
rect 26691 3281 26697 3293
rect 26377 3253 26697 3281
rect 26377 3250 26389 3253
rect 26331 3244 26389 3250
rect 26691 3241 26697 3253
rect 26749 3281 26755 3293
rect 27067 3284 27125 3290
rect 27067 3281 27079 3284
rect 26749 3253 27079 3281
rect 26749 3241 26755 3253
rect 27067 3250 27079 3253
rect 27113 3250 27125 3284
rect 27067 3244 27125 3250
rect 26691 3240 26755 3241
rect 23438 2975 25366 3003
rect 25394 3212 25562 3222
rect 28092 3212 28120 3318
rect 28328 3317 28346 3318
rect 28380 3317 28395 3351
rect 29183 3352 29241 3358
rect 29183 3349 29195 3352
rect 28328 3309 28395 3317
rect 28554 3321 29195 3349
rect 28554 3290 28593 3321
rect 29183 3318 29195 3321
rect 29229 3318 29241 3352
rect 29183 3312 29241 3318
rect 29842 3306 29848 3358
rect 29900 3306 29906 3358
rect 28171 3284 28229 3290
rect 28171 3250 28183 3284
rect 28217 3281 28229 3284
rect 28535 3284 28593 3290
rect 28535 3281 28547 3284
rect 28217 3253 28547 3281
rect 28217 3250 28229 3253
rect 28171 3244 28229 3250
rect 28535 3250 28547 3253
rect 28581 3250 28593 3284
rect 28535 3244 28593 3250
rect 28723 3284 28781 3290
rect 28723 3250 28735 3284
rect 28769 3281 28781 3284
rect 29086 3281 29092 3293
rect 28769 3253 29092 3281
rect 28769 3250 28781 3253
rect 28723 3244 28781 3250
rect 29086 3241 29092 3253
rect 29144 3281 29150 3293
rect 29459 3284 29517 3290
rect 29459 3281 29471 3284
rect 29144 3253 29471 3281
rect 29144 3241 29150 3253
rect 29459 3250 29471 3253
rect 29505 3250 29517 3284
rect 29459 3244 29517 3250
rect 30287 3219 30344 3231
rect 25394 3184 28121 3212
rect 30287 3185 30299 3219
rect 30333 3216 30344 3219
rect 30419 3216 30770 3222
rect 30333 3185 30770 3216
rect 25394 3174 25562 3184
rect 30287 3182 30770 3185
rect 30287 3179 30344 3182
rect 30419 3174 30770 3182
rect 23438 2961 23444 2975
rect 12518 2904 12524 2956
rect 12576 2949 12583 2956
rect 18429 2949 18435 2954
rect 12576 2907 18435 2949
rect 12576 2904 12583 2907
rect 18429 2902 18435 2907
rect 18487 2902 18494 2954
rect 20092 2892 20099 2944
rect 20151 2933 20157 2944
rect 21076 2933 21082 2944
rect 20151 2905 21082 2933
rect 20151 2892 20157 2905
rect 21076 2892 21082 2905
rect 21134 2933 21140 2944
rect 25394 2933 25422 3174
rect 25577 3114 30361 3145
rect 25577 3080 25606 3114
rect 25640 3080 25698 3114
rect 25732 3080 25790 3114
rect 25824 3080 25882 3114
rect 25916 3080 25974 3114
rect 26008 3080 26066 3114
rect 26100 3080 26158 3114
rect 26192 3080 26250 3114
rect 26284 3080 26342 3114
rect 26376 3080 26434 3114
rect 26468 3080 26526 3114
rect 26560 3080 26618 3114
rect 26652 3080 26710 3114
rect 26744 3080 26802 3114
rect 26836 3080 26894 3114
rect 26928 3080 26986 3114
rect 27020 3080 27078 3114
rect 27112 3080 27170 3114
rect 27204 3080 27262 3114
rect 27296 3080 27354 3114
rect 27388 3080 27446 3114
rect 27480 3080 27538 3114
rect 27572 3080 27630 3114
rect 27664 3080 27722 3114
rect 27756 3080 27814 3114
rect 27848 3080 27906 3114
rect 27940 3080 27998 3114
rect 28032 3080 28090 3114
rect 28124 3080 28182 3114
rect 28216 3080 28274 3114
rect 28308 3080 28366 3114
rect 28400 3080 28458 3114
rect 28492 3080 28550 3114
rect 28584 3080 28642 3114
rect 28676 3080 28734 3114
rect 28768 3080 28826 3114
rect 28860 3080 28918 3114
rect 28952 3080 29010 3114
rect 29044 3083 29102 3114
rect 29136 3083 29194 3114
rect 29044 3080 29086 3083
rect 29138 3080 29194 3083
rect 29228 3080 29286 3114
rect 29320 3080 29378 3114
rect 29412 3080 29470 3114
rect 29504 3080 29562 3114
rect 29596 3080 29654 3114
rect 29688 3080 29746 3114
rect 29780 3080 29838 3114
rect 29872 3080 29930 3114
rect 29964 3080 30022 3114
rect 30056 3080 30114 3114
rect 30148 3080 30206 3114
rect 30240 3080 30298 3114
rect 30332 3080 30361 3114
rect 25577 3079 26165 3080
rect 25577 3074 25959 3079
rect 25577 3022 25743 3074
rect 25795 3027 25959 3074
rect 26011 3028 26165 3079
rect 26217 3077 28863 3080
rect 26217 3076 28418 3077
rect 26217 3074 26788 3076
rect 26217 3072 26563 3074
rect 26217 3028 26367 3072
rect 26011 3027 26367 3028
rect 25795 3022 26367 3027
rect 25577 3020 26367 3022
rect 26419 3022 26563 3072
rect 26615 3024 26788 3074
rect 26840 3075 27886 3076
rect 26840 3072 27446 3075
rect 26840 3024 27003 3072
rect 26615 3022 27003 3024
rect 26419 3020 27003 3022
rect 27055 3020 27238 3072
rect 27290 3023 27446 3072
rect 27498 3023 27688 3075
rect 27740 3024 27886 3075
rect 27938 3024 28193 3076
rect 28245 3025 28418 3076
rect 28470 3076 28863 3077
rect 28470 3025 28647 3076
rect 28245 3024 28647 3025
rect 28699 3028 28863 3076
rect 28915 3031 29086 3080
rect 29138 3079 30361 3080
rect 29138 3031 29310 3079
rect 28915 3028 29310 3031
rect 28699 3027 29310 3028
rect 29362 3072 30361 3079
rect 29362 3071 30188 3072
rect 29362 3068 29961 3071
rect 29362 3027 29537 3068
rect 28699 3024 29537 3027
rect 27740 3023 29537 3024
rect 27290 3020 29537 3023
rect 25577 3018 29537 3020
rect 29589 3067 29961 3068
rect 29589 3018 29750 3067
rect 29802 3019 29961 3067
rect 30013 3020 30188 3071
rect 30240 3020 30361 3072
rect 30013 3019 30361 3020
rect 29802 3018 30361 3019
rect 25577 2984 25606 3018
rect 25640 2984 25698 3018
rect 25732 2984 25790 3018
rect 25824 2984 25882 3018
rect 25916 2984 25974 3018
rect 26008 2984 26066 3018
rect 26100 2984 26158 3018
rect 26192 2984 26250 3018
rect 26284 2984 26342 3018
rect 26376 2984 26434 3018
rect 26468 2984 26526 3018
rect 26560 2984 26618 3018
rect 26652 2984 26710 3018
rect 26744 2984 26802 3018
rect 26836 2984 26894 3018
rect 26928 2984 26986 3018
rect 27020 2984 27078 3018
rect 27112 2984 27170 3018
rect 27204 2984 27262 3018
rect 27296 2984 27354 3018
rect 27388 2984 27446 3018
rect 27480 2984 27538 3018
rect 27572 2984 27630 3018
rect 27664 2984 27722 3018
rect 27756 2984 27814 3018
rect 27848 2984 27906 3018
rect 27940 2984 27998 3018
rect 28032 2984 28090 3018
rect 28124 2984 28182 3018
rect 28216 2984 28274 3018
rect 28308 2984 28366 3018
rect 28400 2984 28458 3018
rect 28492 2984 28550 3018
rect 28584 2984 28642 3018
rect 28676 2984 28734 3018
rect 28768 2984 28826 3018
rect 28860 2984 28918 3018
rect 28952 2984 29010 3018
rect 29044 2984 29102 3018
rect 29136 2984 29194 3018
rect 29228 2984 29286 3018
rect 29320 2984 29378 3018
rect 29412 2984 29470 3018
rect 29504 3016 29537 3018
rect 29504 2984 29562 3016
rect 29596 2984 29654 3018
rect 29688 2984 29746 3018
rect 29802 3015 29838 3018
rect 29780 2984 29838 3015
rect 29872 2984 29930 3018
rect 29964 2984 30022 3018
rect 30056 2984 30114 3018
rect 30148 2984 30206 3018
rect 30240 2984 30298 3018
rect 30332 2984 30361 3018
rect 25577 2953 30361 2984
rect 21134 2905 25422 2933
rect 25504 2913 25549 2922
rect 21134 2892 21140 2905
rect 25504 2885 28135 2913
rect 30410 2906 30759 2912
rect 30277 2896 30759 2906
rect 15309 2824 15316 2876
rect 15368 2864 15374 2876
rect 16296 2864 16302 2877
rect 15368 2836 16302 2864
rect 15368 2824 15374 2836
rect 16296 2825 16302 2836
rect 16354 2864 16360 2877
rect 25504 2864 25549 2885
rect 16354 2836 25549 2864
rect 25779 2848 25837 2854
rect 16354 2825 16360 2836
rect 25616 2817 25668 2823
rect 8498 2735 8505 2787
rect 8557 2773 8563 2787
rect 10303 2773 10310 2783
rect 8557 2745 10310 2773
rect 8557 2735 8563 2745
rect 8498 2734 8563 2735
rect 10303 2731 10310 2745
rect 10362 2731 10368 2783
rect 17701 2756 17708 2808
rect 17760 2797 17766 2808
rect 18685 2797 18691 2808
rect 17760 2769 18691 2797
rect 17760 2756 17766 2769
rect 18685 2756 18691 2769
rect 18743 2797 18750 2808
rect 25779 2814 25791 2848
rect 25825 2845 25837 2848
rect 26143 2848 26201 2854
rect 26143 2845 26155 2848
rect 25825 2817 26155 2845
rect 25825 2814 25837 2817
rect 25779 2808 25837 2814
rect 26143 2814 26155 2817
rect 26189 2814 26201 2848
rect 26143 2808 26201 2814
rect 26331 2848 26389 2854
rect 26331 2814 26343 2848
rect 26377 2845 26389 2848
rect 27067 2848 27125 2854
rect 27067 2845 27079 2848
rect 27113 2845 27125 2848
rect 26377 2817 27077 2845
rect 26377 2814 26389 2817
rect 26331 2808 26389 2814
rect 27067 2808 27077 2817
rect 18743 2769 25550 2797
rect 18743 2756 18750 2769
rect 10303 2730 10368 2731
rect 12922 2700 12928 2752
rect 12980 2728 12987 2752
rect 13898 2728 13904 2752
rect 12980 2700 13904 2728
rect 13956 2728 13963 2752
rect 13956 2700 25477 2728
rect 10529 2637 10535 2689
rect 10587 2672 10594 2689
rect 11509 2672 11515 2686
rect 10587 2644 11515 2672
rect 10587 2637 10594 2644
rect 11509 2634 11515 2644
rect 11567 2672 11574 2686
rect 11567 2644 25420 2672
rect 11567 2634 11574 2644
rect 10126 2568 10132 2620
rect 10184 2605 10191 2620
rect 16033 2605 16039 2614
rect 10184 2577 16039 2605
rect 10184 2568 10191 2577
rect 16033 2562 16039 2577
rect 16091 2562 16097 2614
rect 16434 2561 16440 2613
rect 16492 2605 16498 2613
rect 24475 2605 24482 2616
rect 16492 2577 24482 2605
rect 16492 2561 16498 2577
rect 24475 2564 24482 2577
rect 24534 2564 24540 2616
rect 17301 2496 17307 2548
rect 17359 2537 17366 2548
rect 23224 2537 23230 2549
rect 17359 2509 23230 2537
rect 17359 2496 17366 2509
rect 23224 2497 23230 2509
rect 23282 2497 23288 2549
rect 18857 2429 18863 2481
rect 18915 2469 18922 2481
rect 22083 2469 22089 2481
rect 18915 2441 22089 2469
rect 18915 2429 18922 2441
rect 22083 2429 22089 2441
rect 22141 2429 22147 2481
rect 9823 2360 9829 2412
rect 9881 2401 9887 2412
rect 25247 2401 25253 2413
rect 9881 2371 25253 2401
rect 9881 2360 9887 2371
rect 25247 2361 25253 2371
rect 25305 2361 25312 2413
rect 9736 2291 9742 2343
rect 9794 2332 9800 2343
rect 22853 2332 22859 2342
rect 9794 2302 22859 2332
rect 9794 2291 9800 2302
rect 22853 2290 22859 2302
rect 22911 2290 22918 2342
rect 9649 2222 9655 2274
rect 9707 2262 9713 2274
rect 20462 2262 20468 2271
rect 9707 2232 20468 2262
rect 9707 2222 9713 2232
rect 20462 2219 20468 2232
rect 20520 2219 20527 2271
rect 9563 2152 9569 2204
rect 9621 2192 9627 2204
rect 18070 2192 18076 2203
rect 9621 2162 18076 2192
rect 9621 2152 9627 2162
rect 18070 2151 18076 2162
rect 18128 2151 18135 2203
rect 9477 2082 9483 2134
rect 9535 2123 9541 2134
rect 15679 2123 15685 2133
rect 9535 2093 15685 2123
rect 9535 2082 9541 2093
rect 15679 2081 15685 2093
rect 15737 2081 15744 2133
rect 9390 2013 9396 2065
rect 9448 2053 9454 2065
rect 13285 2053 13291 2064
rect 9448 2023 13291 2053
rect 9448 2013 9454 2023
rect 13285 2012 13291 2023
rect 13343 2012 13350 2064
rect 9304 1943 9310 1995
rect 9362 1983 9368 1995
rect 10893 1983 10899 1994
rect 9362 1953 10899 1983
rect 9362 1943 9368 1953
rect 10893 1942 10899 1953
rect 10951 1942 10958 1994
rect 25391 1942 25420 2644
rect 25448 2141 25477 2700
rect 25505 2707 25550 2769
rect 25616 2759 25668 2765
rect 26162 2777 26201 2808
rect 27070 2793 27077 2808
rect 27129 2793 27136 2845
rect 26791 2780 26849 2786
rect 26791 2777 26803 2780
rect 26162 2749 26803 2777
rect 26791 2746 26803 2749
rect 26837 2746 26849 2780
rect 26791 2740 26849 2746
rect 27453 2734 27460 2786
rect 27512 2734 27519 2786
rect 28003 2774 28055 2780
rect 25935 2722 26002 2731
rect 25935 2707 25953 2722
rect 25505 2688 25953 2707
rect 25987 2688 26002 2722
rect 28106 2779 28134 2885
rect 30277 2862 30293 2896
rect 30327 2872 30759 2896
rect 30327 2862 30344 2872
rect 30410 2864 30759 2872
rect 28171 2848 28229 2854
rect 28171 2814 28183 2848
rect 28217 2845 28229 2848
rect 28535 2848 28593 2854
rect 28535 2845 28547 2848
rect 28217 2817 28547 2845
rect 28217 2814 28229 2817
rect 28171 2808 28229 2814
rect 28535 2814 28547 2817
rect 28581 2814 28593 2848
rect 28535 2808 28593 2814
rect 28723 2848 28781 2854
rect 28723 2814 28735 2848
rect 28769 2845 28781 2848
rect 29459 2848 29517 2854
rect 30277 2852 30344 2862
rect 29459 2847 29471 2848
rect 29505 2847 29517 2848
rect 29459 2845 29469 2847
rect 28769 2817 29469 2845
rect 28769 2814 28781 2817
rect 28723 2808 28781 2814
rect 29459 2808 29469 2817
rect 28329 2779 28396 2788
rect 28106 2751 28347 2779
rect 28329 2745 28347 2751
rect 28381 2745 28396 2779
rect 28554 2777 28593 2808
rect 29462 2795 29469 2808
rect 29521 2795 29528 2847
rect 29183 2780 29241 2786
rect 29183 2777 29195 2780
rect 28554 2749 29195 2777
rect 28329 2737 28396 2745
rect 29183 2746 29195 2749
rect 29229 2746 29241 2780
rect 29183 2740 29241 2746
rect 29839 2741 29846 2793
rect 29898 2741 29905 2793
rect 25505 2680 26002 2688
rect 26699 2712 26757 2718
rect 25505 2679 25951 2680
rect 25505 2671 25550 2679
rect 26699 2678 26711 2712
rect 26745 2709 26757 2712
rect 27343 2712 27401 2718
rect 28003 2716 28055 2722
rect 27343 2709 27355 2712
rect 26745 2681 27355 2709
rect 26745 2678 26757 2681
rect 26699 2672 26757 2678
rect 27343 2678 27355 2681
rect 27389 2678 27401 2712
rect 27343 2672 27401 2678
rect 29091 2712 29149 2718
rect 29091 2678 29103 2712
rect 29137 2709 29149 2712
rect 29735 2712 29793 2718
rect 29735 2709 29747 2712
rect 29137 2681 29747 2709
rect 29137 2678 29149 2681
rect 29091 2672 29149 2678
rect 29735 2678 29747 2681
rect 29781 2678 29793 2712
rect 29735 2672 29793 2678
rect 25687 2644 25745 2650
rect 25687 2610 25699 2644
rect 25733 2641 25745 2644
rect 26055 2644 26113 2650
rect 26055 2641 26067 2644
rect 25733 2613 26067 2641
rect 25733 2610 25745 2613
rect 25687 2604 25745 2610
rect 26055 2610 26067 2613
rect 26101 2641 26113 2644
rect 26791 2644 26849 2650
rect 26791 2641 26803 2644
rect 26101 2613 26803 2641
rect 26101 2610 26113 2613
rect 26055 2604 26113 2610
rect 26791 2610 26803 2613
rect 26837 2610 26849 2644
rect 26791 2604 26849 2610
rect 28079 2644 28137 2650
rect 28079 2610 28091 2644
rect 28125 2641 28137 2644
rect 28447 2644 28505 2650
rect 28447 2641 28459 2644
rect 28125 2613 28459 2641
rect 28125 2610 28137 2613
rect 28079 2604 28137 2610
rect 28447 2610 28459 2613
rect 28493 2641 28505 2644
rect 29183 2644 29241 2650
rect 29183 2641 29195 2644
rect 28493 2613 29195 2641
rect 28493 2610 28505 2613
rect 28447 2604 28505 2610
rect 29183 2610 29195 2613
rect 29229 2610 29241 2644
rect 29183 2604 29241 2610
rect 27891 2585 27954 2591
rect 27891 2551 27906 2585
rect 27940 2572 27954 2585
rect 30413 2572 30765 2581
rect 27940 2551 30765 2572
rect 27891 2544 30765 2551
rect 30413 2533 30765 2544
rect 25577 2474 30361 2505
rect 25577 2440 25606 2474
rect 25640 2440 25698 2474
rect 25732 2440 25790 2474
rect 25824 2440 25882 2474
rect 25916 2440 25974 2474
rect 26008 2440 26066 2474
rect 26100 2440 26158 2474
rect 26192 2440 26250 2474
rect 26284 2440 26342 2474
rect 26376 2440 26434 2474
rect 26468 2440 26526 2474
rect 26560 2440 26618 2474
rect 26652 2440 26710 2474
rect 26744 2440 26802 2474
rect 26836 2440 26894 2474
rect 26928 2440 26986 2474
rect 27020 2440 27078 2474
rect 27112 2440 27170 2474
rect 27204 2440 27262 2474
rect 27296 2440 27354 2474
rect 27388 2443 27446 2474
rect 27388 2440 27395 2443
rect 27480 2440 27538 2474
rect 27572 2440 27630 2474
rect 27664 2445 27722 2474
rect 27685 2440 27722 2445
rect 27756 2440 27814 2474
rect 27848 2447 27906 2474
rect 27898 2440 27906 2447
rect 27940 2440 27998 2474
rect 28032 2440 28090 2474
rect 28124 2440 28182 2474
rect 28216 2440 28274 2474
rect 28308 2440 28366 2474
rect 28400 2440 28458 2474
rect 28492 2440 28550 2474
rect 28584 2440 28642 2474
rect 28676 2440 28734 2474
rect 28768 2440 28826 2474
rect 28860 2440 28918 2474
rect 28952 2440 29010 2474
rect 29044 2440 29102 2474
rect 29136 2440 29194 2474
rect 29228 2440 29286 2474
rect 29320 2440 29378 2474
rect 29412 2440 29470 2474
rect 29504 2440 29562 2474
rect 29596 2440 29654 2474
rect 29688 2440 29746 2474
rect 29780 2440 29838 2474
rect 29872 2440 29930 2474
rect 29964 2440 30022 2474
rect 30056 2440 30114 2474
rect 30148 2440 30206 2474
rect 30240 2440 30298 2474
rect 30332 2440 30361 2474
rect 25577 2439 27395 2440
rect 25577 2438 26963 2439
rect 25577 2429 25994 2438
rect 25577 2378 25769 2429
rect 25821 2386 25994 2429
rect 26046 2435 26492 2438
rect 26046 2386 26271 2435
rect 25821 2383 26271 2386
rect 26323 2386 26492 2435
rect 26544 2435 26963 2438
rect 26544 2386 26737 2435
rect 26323 2383 26737 2386
rect 26789 2387 26963 2435
rect 27015 2437 27395 2439
rect 27015 2387 27175 2437
rect 26789 2385 27175 2387
rect 27227 2391 27395 2437
rect 27447 2393 27633 2440
rect 27685 2395 27846 2440
rect 27898 2438 30361 2440
rect 27898 2437 28580 2438
rect 27898 2395 28233 2437
rect 27685 2393 28233 2395
rect 27447 2391 28233 2393
rect 27227 2385 28233 2391
rect 28285 2386 28580 2437
rect 28632 2435 30361 2438
rect 28632 2433 29239 2435
rect 28632 2386 28816 2433
rect 28285 2385 28816 2386
rect 26789 2383 28816 2385
rect 25821 2381 28816 2383
rect 28868 2381 29000 2433
rect 29052 2383 29239 2433
rect 29291 2434 30361 2435
rect 29291 2431 30009 2434
rect 29291 2383 29442 2431
rect 29052 2381 29442 2383
rect 25821 2379 29442 2381
rect 29494 2430 30009 2431
rect 29494 2428 29818 2430
rect 29494 2379 29627 2428
rect 25821 2378 29627 2379
rect 29679 2378 29818 2428
rect 29870 2382 30009 2430
rect 30061 2430 30361 2434
rect 30061 2382 30195 2430
rect 29870 2378 30195 2382
rect 30247 2378 30361 2430
rect 25577 2344 25606 2378
rect 25640 2344 25698 2378
rect 25732 2377 25769 2378
rect 25732 2344 25790 2377
rect 25824 2344 25882 2378
rect 25916 2344 25974 2378
rect 26008 2344 26066 2378
rect 26100 2344 26158 2378
rect 26192 2344 26250 2378
rect 26284 2344 26342 2378
rect 26376 2344 26434 2378
rect 26468 2344 26526 2378
rect 26560 2344 26618 2378
rect 26652 2344 26710 2378
rect 26744 2344 26802 2378
rect 26836 2344 26894 2378
rect 26928 2344 26986 2378
rect 27020 2344 27078 2378
rect 27112 2344 27170 2378
rect 27204 2344 27262 2378
rect 27296 2344 27354 2378
rect 27388 2344 27446 2378
rect 27480 2344 27538 2378
rect 27572 2344 27630 2378
rect 27664 2344 27722 2378
rect 27756 2344 27814 2378
rect 27848 2344 27906 2378
rect 27940 2344 27998 2378
rect 28032 2344 28090 2378
rect 28124 2344 28182 2378
rect 28216 2344 28274 2378
rect 28308 2344 28366 2378
rect 28400 2344 28458 2378
rect 28492 2344 28550 2378
rect 28584 2344 28642 2378
rect 28676 2344 28734 2378
rect 28768 2344 28826 2378
rect 28860 2344 28918 2378
rect 28952 2344 29010 2378
rect 29044 2344 29102 2378
rect 29136 2344 29194 2378
rect 29228 2344 29286 2378
rect 29320 2344 29378 2378
rect 29412 2344 29470 2378
rect 29504 2344 29562 2378
rect 29596 2376 29627 2378
rect 29596 2344 29654 2376
rect 29688 2344 29746 2378
rect 29780 2344 29838 2378
rect 29872 2344 29930 2378
rect 29964 2344 30022 2378
rect 30056 2344 30114 2378
rect 30148 2344 30206 2378
rect 30240 2344 30298 2378
rect 30332 2344 30361 2378
rect 25577 2313 30361 2344
rect 30416 2277 30762 2285
rect 27894 2270 30762 2277
rect 27894 2236 27906 2270
rect 27940 2249 30762 2270
rect 27940 2236 27952 2249
rect 30416 2237 30762 2249
rect 27894 2229 27952 2236
rect 25687 2208 25745 2214
rect 25687 2174 25699 2208
rect 25733 2205 25745 2208
rect 26055 2208 26113 2214
rect 26055 2205 26067 2208
rect 25733 2177 26067 2205
rect 25733 2174 25745 2177
rect 25687 2168 25745 2174
rect 26055 2174 26067 2177
rect 26101 2205 26113 2208
rect 26791 2208 26849 2214
rect 26791 2205 26803 2208
rect 26101 2177 26803 2205
rect 26101 2174 26113 2177
rect 26055 2168 26113 2174
rect 26791 2174 26803 2177
rect 26837 2174 26849 2208
rect 26791 2168 26849 2174
rect 28079 2208 28137 2214
rect 28079 2174 28091 2208
rect 28125 2205 28137 2208
rect 28447 2208 28505 2214
rect 28447 2205 28459 2208
rect 28125 2177 28459 2205
rect 28125 2174 28137 2177
rect 28079 2168 28137 2174
rect 28447 2174 28459 2177
rect 28493 2205 28505 2208
rect 29183 2208 29241 2214
rect 29183 2205 29195 2208
rect 28493 2177 29195 2205
rect 28493 2174 28505 2177
rect 28447 2168 28505 2174
rect 29183 2174 29195 2177
rect 29229 2174 29241 2208
rect 29183 2168 29241 2174
rect 25448 2129 25551 2141
rect 26699 2140 26757 2146
rect 25932 2130 25999 2139
rect 25932 2129 25950 2130
rect 25448 2101 25950 2129
rect 25448 2093 25551 2101
rect 25932 2096 25950 2101
rect 25984 2096 25999 2130
rect 26699 2106 26711 2140
rect 26745 2137 26757 2140
rect 27343 2140 27401 2146
rect 27343 2137 27355 2140
rect 26745 2109 27355 2137
rect 26745 2106 26757 2109
rect 26699 2100 26757 2106
rect 27343 2106 27355 2109
rect 27389 2106 27401 2140
rect 27343 2100 27401 2106
rect 29091 2140 29149 2146
rect 29091 2106 29103 2140
rect 29137 2137 29149 2140
rect 29735 2140 29793 2146
rect 29735 2137 29747 2140
rect 29137 2109 29747 2137
rect 29137 2106 29149 2109
rect 29091 2100 29149 2106
rect 29735 2106 29747 2109
rect 29781 2106 29793 2140
rect 29735 2100 29793 2106
rect 25932 2088 25999 2096
rect 28004 2087 28056 2093
rect 27449 2078 27514 2079
rect 26791 2072 26849 2078
rect 26791 2069 26803 2072
rect 25611 2057 25663 2063
rect 26162 2041 26803 2069
rect 26162 2010 26201 2041
rect 26791 2038 26803 2041
rect 26837 2038 26849 2072
rect 26791 2032 26849 2038
rect 27449 2026 27455 2078
rect 27507 2026 27514 2078
rect 28330 2071 28397 2080
rect 29841 2079 29905 2080
rect 28330 2066 28348 2071
rect 28004 2029 28056 2035
rect 28093 2038 28348 2066
rect 25611 1999 25663 2005
rect 25779 2004 25837 2010
rect 25779 1970 25791 2004
rect 25825 2001 25837 2004
rect 26143 2004 26201 2010
rect 26143 2001 26155 2004
rect 25825 1973 26155 2001
rect 25825 1970 25837 1973
rect 25779 1964 25837 1970
rect 26143 1970 26155 1973
rect 26189 1970 26201 2004
rect 26143 1964 26201 1970
rect 26331 2004 26389 2010
rect 26331 1970 26343 2004
rect 26377 2001 26389 2004
rect 26698 2001 26706 2013
rect 26377 1973 26706 2001
rect 26377 1970 26389 1973
rect 26331 1964 26389 1970
rect 26698 1961 26706 1973
rect 26758 2001 26764 2013
rect 27067 2004 27125 2010
rect 27067 2001 27079 2004
rect 26758 1973 27079 2001
rect 26758 1961 26764 1973
rect 27067 1970 27079 1973
rect 27113 1970 27125 2004
rect 27067 1964 27125 1970
rect 25391 1932 25534 1942
rect 28093 1932 28121 2038
rect 28330 2037 28348 2038
rect 28382 2037 28397 2071
rect 29183 2072 29241 2078
rect 29183 2069 29195 2072
rect 28330 2029 28397 2037
rect 28554 2041 29195 2069
rect 28554 2010 28593 2041
rect 29183 2038 29195 2041
rect 29229 2038 29241 2072
rect 29183 2032 29241 2038
rect 29841 2027 29847 2079
rect 29899 2027 29905 2079
rect 28171 2004 28229 2010
rect 28171 1970 28183 2004
rect 28217 2001 28229 2004
rect 28535 2004 28593 2010
rect 28535 2001 28547 2004
rect 28217 1973 28547 2001
rect 28217 1970 28229 1973
rect 28171 1964 28229 1970
rect 28535 1970 28547 1973
rect 28581 1970 28593 2004
rect 28535 1964 28593 1970
rect 28723 2004 28781 2010
rect 28723 1970 28735 2004
rect 28769 2001 28781 2004
rect 29089 2001 29096 2013
rect 28769 1973 29096 2001
rect 28769 1970 28781 1973
rect 28723 1964 28781 1970
rect 29089 1961 29096 1973
rect 29149 2001 29156 2013
rect 29459 2004 29517 2010
rect 29459 2001 29471 2004
rect 29149 1973 29471 2001
rect 29149 1961 29156 1973
rect 29459 1970 29471 1973
rect 29505 1970 29517 2004
rect 29459 1964 29517 1970
rect 30282 1937 30340 1944
rect 9218 1873 9224 1925
rect 9276 1913 9282 1925
rect 23055 1913 23061 1924
rect 9276 1883 23061 1913
rect 9276 1873 9282 1883
rect 23055 1872 23061 1883
rect 23113 1872 23120 1924
rect 25391 1904 28122 1932
rect 25391 1894 25534 1904
rect 30282 1903 30294 1937
rect 30328 1935 30340 1937
rect 30412 1935 30760 1941
rect 30328 1903 30760 1935
rect 30282 1901 30760 1903
rect 30282 1897 30340 1901
rect 30412 1893 30760 1901
rect 9132 1803 9138 1855
rect 9190 1844 9196 1855
rect 20666 1844 20672 1854
rect 9190 1814 20672 1844
rect 9190 1803 9196 1814
rect 20666 1802 20672 1814
rect 20724 1802 20731 1854
rect 25577 1849 30361 1865
rect 25577 1848 28357 1849
rect 25577 1847 26033 1848
rect 25577 1834 25642 1847
rect 25577 1800 25606 1834
rect 25640 1800 25642 1834
rect 25577 1795 25642 1800
rect 25694 1843 26033 1847
rect 25694 1834 25847 1843
rect 25899 1834 26033 1843
rect 26085 1846 28357 1848
rect 26085 1841 26446 1846
rect 26085 1834 26227 1841
rect 26279 1834 26446 1841
rect 26498 1834 26656 1846
rect 25694 1800 25698 1834
rect 25732 1800 25790 1834
rect 25824 1800 25847 1834
rect 25916 1800 25974 1834
rect 26008 1800 26033 1834
rect 26100 1800 26158 1834
rect 26192 1800 26227 1834
rect 26284 1800 26342 1834
rect 26376 1800 26434 1834
rect 26498 1800 26526 1834
rect 26560 1800 26618 1834
rect 26652 1800 26656 1834
rect 25694 1795 25847 1800
rect 25577 1791 25847 1795
rect 25899 1796 26033 1800
rect 26085 1796 26227 1800
rect 25899 1791 26227 1796
rect 25577 1789 26227 1791
rect 26279 1794 26446 1800
rect 26498 1794 26656 1800
rect 26708 1843 28139 1846
rect 26708 1834 26885 1843
rect 26937 1834 27131 1843
rect 27183 1834 27405 1843
rect 27457 1834 27680 1843
rect 27732 1834 27916 1843
rect 27968 1834 28139 1843
rect 28191 1834 28357 1846
rect 28409 1847 30361 1849
rect 28409 1843 29802 1847
rect 28409 1842 29382 1843
rect 28409 1840 28774 1842
rect 28409 1834 28535 1840
rect 28587 1834 28774 1840
rect 26708 1800 26710 1834
rect 26744 1800 26802 1834
rect 26836 1800 26885 1834
rect 26937 1800 26986 1834
rect 27020 1800 27078 1834
rect 27112 1800 27131 1834
rect 27204 1800 27262 1834
rect 27296 1800 27354 1834
rect 27388 1800 27405 1834
rect 27480 1800 27538 1834
rect 27572 1800 27630 1834
rect 27664 1800 27680 1834
rect 27756 1800 27814 1834
rect 27848 1800 27906 1834
rect 27968 1800 27998 1834
rect 28032 1800 28090 1834
rect 28124 1800 28139 1834
rect 28216 1800 28274 1834
rect 28308 1800 28357 1834
rect 28409 1800 28458 1834
rect 28492 1800 28535 1834
rect 28587 1800 28642 1834
rect 28676 1800 28734 1834
rect 28768 1800 28774 1834
rect 26708 1794 26885 1800
rect 26279 1791 26885 1794
rect 26937 1791 27131 1800
rect 27183 1791 27405 1800
rect 27457 1791 27680 1800
rect 27732 1791 27916 1800
rect 27968 1794 28139 1800
rect 28191 1797 28357 1800
rect 28409 1797 28535 1800
rect 28191 1794 28535 1797
rect 27968 1791 28535 1794
rect 26279 1789 28535 1791
rect 25577 1788 28535 1789
rect 28587 1790 28774 1800
rect 28826 1834 28971 1842
rect 29023 1834 29169 1842
rect 29221 1834 29382 1842
rect 29434 1842 29802 1843
rect 29434 1834 29605 1842
rect 29657 1834 29802 1842
rect 29854 1845 30361 1847
rect 29854 1834 30018 1845
rect 30070 1834 30227 1845
rect 30279 1834 30361 1845
rect 28860 1800 28918 1834
rect 28952 1800 28971 1834
rect 29044 1800 29102 1834
rect 29136 1800 29169 1834
rect 29228 1800 29286 1834
rect 29320 1800 29378 1834
rect 29434 1800 29470 1834
rect 29504 1800 29562 1834
rect 29596 1800 29605 1834
rect 29688 1800 29746 1834
rect 29780 1800 29802 1834
rect 29872 1800 29930 1834
rect 29964 1800 30018 1834
rect 30070 1800 30114 1834
rect 30148 1800 30206 1834
rect 30279 1800 30298 1834
rect 30332 1800 30361 1834
rect 28826 1790 28971 1800
rect 29023 1790 29169 1800
rect 29221 1791 29382 1800
rect 29434 1791 29605 1800
rect 29221 1790 29605 1791
rect 29657 1795 29802 1800
rect 29854 1795 30018 1800
rect 29657 1793 30018 1795
rect 30070 1793 30227 1800
rect 30279 1793 30361 1800
rect 29657 1790 30361 1793
rect 28587 1788 30361 1790
rect 9045 1734 9051 1786
rect 9103 1774 9109 1786
rect 18273 1774 18279 1785
rect 9103 1744 18279 1774
rect 9103 1734 9109 1744
rect 18273 1733 18279 1744
rect 18331 1733 18338 1785
rect 25577 1769 30361 1788
rect 25606 1766 25640 1769
rect 25698 1766 25732 1769
rect 25790 1766 25824 1769
rect 25882 1766 25916 1769
rect 25974 1766 26008 1769
rect 26066 1766 26100 1769
rect 26158 1766 26192 1769
rect 26250 1766 26284 1769
rect 26342 1766 26376 1769
rect 26434 1766 26468 1769
rect 26526 1766 26560 1769
rect 26618 1766 26652 1769
rect 26710 1766 26744 1769
rect 26802 1766 26836 1769
rect 26894 1766 26928 1769
rect 26986 1766 27020 1769
rect 27078 1766 27112 1769
rect 27170 1766 27204 1769
rect 27262 1766 27296 1769
rect 27354 1766 27388 1769
rect 27446 1766 27480 1769
rect 27538 1766 27572 1769
rect 27630 1766 27664 1769
rect 27722 1766 27756 1769
rect 27814 1766 27848 1769
rect 27906 1766 27940 1769
rect 27998 1766 28032 1769
rect 28090 1766 28124 1769
rect 28182 1766 28216 1769
rect 28274 1766 28308 1769
rect 28366 1766 28400 1769
rect 28458 1766 28492 1769
rect 28550 1766 28584 1769
rect 28642 1766 28676 1769
rect 28734 1766 28768 1769
rect 28826 1766 28860 1769
rect 28918 1766 28952 1769
rect 29010 1766 29044 1769
rect 29102 1766 29136 1769
rect 29194 1766 29228 1769
rect 29286 1766 29320 1769
rect 29378 1766 29412 1769
rect 29470 1766 29504 1769
rect 29562 1766 29596 1769
rect 29654 1766 29688 1769
rect 29746 1766 29780 1769
rect 29838 1766 29872 1769
rect 29930 1766 29964 1769
rect 30022 1766 30056 1769
rect 30114 1766 30148 1769
rect 30206 1766 30240 1769
rect 30298 1766 30332 1769
rect 8959 1664 8965 1716
rect 9017 1705 9023 1716
rect 15880 1705 15886 1715
rect 9017 1675 15886 1705
rect 9017 1664 9023 1675
rect 15880 1663 15886 1675
rect 15938 1663 15945 1715
rect 8872 1595 8878 1647
rect 8930 1635 8936 1647
rect 13488 1635 13494 1646
rect 8930 1605 13494 1635
rect 8930 1595 8936 1605
rect 13488 1594 13494 1605
rect 13546 1594 13553 1646
rect 8786 1525 8792 1577
rect 8844 1565 8850 1577
rect 11098 1565 11104 1575
rect 8844 1535 11104 1565
rect 8844 1525 8850 1535
rect 11098 1523 11104 1535
rect 11156 1523 11163 1575
rect 8449 1415 24265 1437
rect 8449 1413 9840 1415
rect 8449 1411 8830 1413
rect 8449 1406 8628 1411
rect 8680 1406 8830 1411
rect 8449 1372 8606 1406
rect 8680 1372 8698 1406
rect 8732 1372 8790 1406
rect 8824 1372 8830 1406
rect 8449 1359 8628 1372
rect 8680 1361 8830 1372
rect 8882 1411 9439 1413
rect 8882 1406 9041 1411
rect 9093 1406 9231 1411
rect 9283 1406 9439 1411
rect 9491 1406 9641 1413
rect 9693 1406 9840 1413
rect 8916 1372 8974 1406
rect 9008 1372 9041 1406
rect 9100 1372 9158 1406
rect 9192 1372 9231 1406
rect 9284 1372 9342 1406
rect 9376 1372 9434 1406
rect 9491 1372 9526 1406
rect 9560 1372 9618 1406
rect 9693 1372 9710 1406
rect 9744 1372 9802 1406
rect 9836 1372 9840 1406
rect 8882 1361 9041 1372
rect 8680 1359 9041 1361
rect 9093 1359 9231 1372
rect 9283 1361 9439 1372
rect 9491 1361 9641 1372
rect 9693 1363 9840 1372
rect 9892 1414 10727 1415
rect 9892 1412 10236 1414
rect 9892 1406 10035 1412
rect 10087 1406 10236 1412
rect 10288 1412 10727 1414
rect 10288 1406 10453 1412
rect 10505 1406 10727 1412
rect 10779 1411 24265 1415
rect 10779 1408 11227 1411
rect 10779 1406 11004 1408
rect 11056 1406 11227 1408
rect 11279 1410 24265 1411
rect 11279 1406 11459 1410
rect 9892 1372 9894 1406
rect 9928 1372 9986 1406
rect 10020 1372 10035 1406
rect 10112 1372 10170 1406
rect 10204 1372 10236 1406
rect 10296 1372 10354 1406
rect 10388 1372 10446 1406
rect 10505 1372 10538 1406
rect 10572 1372 10630 1406
rect 10664 1372 10722 1406
rect 10779 1372 10814 1406
rect 10848 1372 10906 1406
rect 10940 1372 10998 1406
rect 11056 1372 11090 1406
rect 11124 1372 11182 1406
rect 11216 1372 11227 1406
rect 11308 1372 11366 1406
rect 11400 1372 11459 1406
rect 9892 1363 10035 1372
rect 9693 1361 10035 1363
rect 9283 1360 10035 1361
rect 10087 1362 10236 1372
rect 10288 1362 10453 1372
rect 10087 1360 10453 1362
rect 10505 1363 10727 1372
rect 10779 1363 11004 1372
rect 10505 1360 11004 1363
rect 9283 1359 11004 1360
rect 8449 1356 11004 1359
rect 11056 1359 11227 1372
rect 11279 1359 11459 1372
rect 11056 1358 11459 1359
rect 11511 1409 14478 1410
rect 11511 1408 13603 1409
rect 11511 1407 13403 1408
rect 11511 1406 13095 1407
rect 13147 1406 13403 1407
rect 13455 1406 13603 1408
rect 13655 1408 14276 1409
rect 13655 1406 13822 1408
rect 13874 1407 14276 1408
rect 13874 1406 14068 1407
rect 14120 1406 14276 1407
rect 14328 1406 14478 1409
rect 14530 1409 24265 1410
rect 14530 1406 14671 1409
rect 14723 1408 24265 1409
rect 14723 1406 15043 1408
rect 15095 1406 15795 1408
rect 11511 1372 12990 1406
rect 13024 1372 13082 1406
rect 13147 1372 13174 1406
rect 13208 1372 13266 1406
rect 13300 1372 13358 1406
rect 13392 1372 13403 1406
rect 13484 1372 13542 1406
rect 13576 1372 13603 1406
rect 13668 1372 13726 1406
rect 13760 1372 13818 1406
rect 13874 1372 13910 1406
rect 13944 1372 14002 1406
rect 14036 1372 14068 1406
rect 14128 1372 14186 1406
rect 14220 1372 14276 1406
rect 14328 1372 14370 1406
rect 14404 1372 14462 1406
rect 14530 1372 14554 1406
rect 14588 1372 14646 1406
rect 14723 1372 14738 1406
rect 14772 1372 14830 1406
rect 14864 1372 14922 1406
rect 14956 1372 15014 1406
rect 15095 1372 15106 1406
rect 15140 1372 15198 1406
rect 11511 1358 13095 1372
rect 11056 1356 13095 1358
rect 8449 1355 13095 1356
rect 13147 1356 13403 1372
rect 13455 1357 13603 1372
rect 13655 1357 13822 1372
rect 13455 1356 13822 1357
rect 13874 1356 14068 1372
rect 13147 1355 14068 1356
rect 14120 1357 14276 1372
rect 14328 1358 14478 1372
rect 14530 1358 14671 1372
rect 14328 1357 14671 1358
rect 14723 1357 15043 1372
rect 14120 1356 15043 1357
rect 15095 1356 15232 1372
rect 14120 1355 15232 1356
rect 8449 1354 15232 1355
rect 15284 1372 15290 1406
rect 15324 1372 15382 1406
rect 15416 1372 15474 1406
rect 15508 1372 15522 1406
rect 15600 1372 15658 1406
rect 15692 1372 15750 1406
rect 15784 1372 15795 1406
rect 15284 1354 15522 1372
rect 15574 1356 15795 1372
rect 15847 1356 24265 1408
rect 15574 1354 24265 1356
rect 8449 1341 24265 1354
rect 8489 1191 8497 1216
rect 8449 1164 8497 1191
rect 8549 1164 8555 1216
rect 8449 1157 8541 1164
rect 8507 1116 8541 1157
rect 8602 1116 8660 1122
rect 8507 1110 8660 1116
rect 8507 1082 8614 1110
rect 8601 1076 8614 1082
rect 8648 1076 8660 1110
rect 8601 1066 8660 1076
rect 11435 1057 11441 1109
rect 11493 1057 11499 1109
rect 15739 1103 15791 1109
rect 15996 1103 16002 1109
rect 15739 1101 16002 1103
rect 12986 1093 13044 1099
rect 12986 1091 12998 1093
rect 12845 1059 12998 1091
rect 13032 1059 13044 1093
rect 11910 995 11916 1019
rect 8449 967 11916 995
rect 11968 995 11974 1019
rect 12845 995 12877 1059
rect 12986 1053 13044 1059
rect 15739 1067 15751 1101
rect 15785 1067 16002 1101
rect 15739 1061 16002 1067
rect 15739 1055 15791 1061
rect 15996 1057 16002 1061
rect 16054 1057 16060 1109
rect 11968 967 12877 995
rect 8449 961 12877 967
rect 8449 883 25436 893
rect 8449 876 25451 883
rect 8449 872 9965 876
rect 8449 862 9746 872
rect 8449 828 8606 862
rect 8640 828 8698 862
rect 8732 828 8790 862
rect 8824 828 8882 862
rect 8916 828 8974 862
rect 9008 828 9066 862
rect 9100 828 9158 862
rect 9192 828 9250 862
rect 9284 828 9342 862
rect 9376 828 9434 862
rect 9468 828 9526 862
rect 9560 828 9618 862
rect 9652 828 9710 862
rect 9744 828 9746 862
rect 8449 820 9746 828
rect 9798 862 9965 872
rect 10017 862 10248 876
rect 10300 862 10457 876
rect 10509 875 25451 876
rect 10509 874 13052 875
rect 10509 862 10728 874
rect 10780 872 13052 874
rect 10780 862 12803 872
rect 9798 828 9802 862
rect 9836 828 9894 862
rect 9928 828 9965 862
rect 10020 828 10078 862
rect 10112 828 10170 862
rect 10204 828 10248 862
rect 10300 828 10354 862
rect 10388 828 10446 862
rect 10509 828 10538 862
rect 10572 828 10630 862
rect 10664 828 10722 862
rect 10780 828 10814 862
rect 10848 828 10906 862
rect 10940 828 10998 862
rect 11032 828 11090 862
rect 11124 828 11182 862
rect 11216 828 11274 862
rect 11308 828 11366 862
rect 11400 828 12803 862
rect 9798 824 9965 828
rect 10017 824 10248 828
rect 10300 824 10457 828
rect 10509 824 10728 828
rect 9798 822 10728 824
rect 10780 822 12803 828
rect 9798 820 12803 822
rect 12855 862 13052 872
rect 13104 874 25451 875
rect 13104 872 15801 874
rect 13104 867 15597 872
rect 13104 862 13650 867
rect 13702 862 13879 867
rect 13931 862 15597 867
rect 15649 862 15801 872
rect 12855 828 12990 862
rect 13024 828 13052 862
rect 13116 828 13174 862
rect 13208 828 13266 862
rect 13300 828 13358 862
rect 13392 861 13450 862
rect 13392 828 13396 861
rect 12855 823 13052 828
rect 13104 823 13396 828
rect 12855 820 13396 823
rect 8449 809 13396 820
rect 13448 828 13450 861
rect 13484 828 13542 862
rect 13576 828 13634 862
rect 13702 828 13726 862
rect 13760 828 13818 862
rect 13852 828 13879 862
rect 13944 828 14002 862
rect 14036 828 14094 862
rect 14128 828 14186 862
rect 14220 828 14278 862
rect 14312 828 14370 862
rect 14404 828 14462 862
rect 14496 828 14554 862
rect 14588 828 14646 862
rect 14680 828 14738 862
rect 14772 828 14830 862
rect 14864 828 14922 862
rect 14956 828 15014 862
rect 15048 828 15106 862
rect 15140 828 15198 862
rect 15232 828 15290 862
rect 15324 828 15382 862
rect 15416 828 15474 862
rect 15508 828 15566 862
rect 15649 828 15658 862
rect 15692 828 15750 862
rect 15784 828 15801 862
rect 13448 815 13650 828
rect 13702 815 13879 828
rect 13931 820 15597 828
rect 15649 822 15801 828
rect 15853 872 25451 874
rect 15853 822 16124 872
rect 15649 820 16124 822
rect 16176 820 25451 872
rect 13931 815 25451 820
rect 13448 809 25451 815
rect 8449 797 25451 809
rect 9593 729 9599 738
rect 8670 695 9599 729
rect 9593 685 9599 695
rect 9652 729 9658 738
rect 11435 729 11441 737
rect 9652 695 11441 729
rect 9652 685 9658 695
rect 11435 685 11441 695
rect 11493 729 11499 737
rect 11987 729 11993 744
rect 11493 695 11993 729
rect 11493 685 11499 695
rect 11987 691 11993 695
rect 12046 729 12052 744
rect 14378 729 14384 744
rect 12046 695 14384 729
rect 12046 691 12052 695
rect 11987 690 12052 691
rect 14378 691 14384 695
rect 14437 729 14443 744
rect 16769 729 16775 744
rect 14437 695 16775 729
rect 14437 691 14443 695
rect 15991 694 16108 695
rect 14378 690 14443 691
rect 16769 691 16775 695
rect 16828 729 16834 744
rect 19161 729 19167 744
rect 16828 695 19167 729
rect 16828 691 16834 695
rect 16769 690 16834 691
rect 19161 691 19167 695
rect 19220 729 19226 744
rect 21552 729 21558 744
rect 19220 695 21558 729
rect 19220 691 19226 695
rect 19161 690 19226 691
rect 21552 691 21558 695
rect 21611 729 21617 744
rect 23945 729 23951 744
rect 21611 695 23951 729
rect 21611 691 21617 695
rect 21552 690 21617 691
rect 23945 691 23951 695
rect 24004 729 24010 744
rect 24004 695 25436 729
rect 24004 691 24010 695
rect 23945 690 24010 691
rect 9593 684 9658 685
rect 8670 621 25436 623
rect 8670 589 25451 621
rect 15994 588 16103 589
rect 9042 517 9049 526
rect 8670 483 9049 517
rect 9042 474 9049 483
rect 9101 517 9108 526
rect 10304 517 10311 526
rect 9101 483 10311 517
rect 9101 474 9108 483
rect 10304 474 10311 483
rect 10363 517 10370 526
rect 11435 517 11442 525
rect 10363 483 11442 517
rect 10363 474 10370 483
rect 11435 473 11442 483
rect 11494 517 11501 525
rect 12696 517 12703 526
rect 11494 483 12703 517
rect 11494 473 11501 483
rect 12696 474 12703 483
rect 12755 517 12762 526
rect 13827 517 13834 525
rect 12755 483 13834 517
rect 12755 474 12762 483
rect 13827 473 13834 483
rect 13886 517 13893 525
rect 15087 517 15094 527
rect 13886 483 15094 517
rect 13886 473 13893 483
rect 15087 475 15094 483
rect 15146 517 15153 527
rect 15996 517 16002 525
rect 15146 483 16002 517
rect 15146 475 15153 483
rect 15996 473 16002 483
rect 16054 517 16060 525
rect 16219 517 16226 526
rect 16054 483 16226 517
rect 16054 473 16060 483
rect 16219 474 16226 483
rect 16278 517 16285 526
rect 17480 517 17487 527
rect 16278 483 17487 517
rect 16278 474 16285 483
rect 17480 475 17487 483
rect 17539 517 17546 527
rect 18610 517 18617 525
rect 17539 483 18617 517
rect 17539 475 17546 483
rect 18610 473 18617 483
rect 18669 517 18676 525
rect 19873 517 19880 527
rect 18669 483 19880 517
rect 18669 473 18676 483
rect 19873 475 19880 483
rect 19932 517 19939 527
rect 21002 517 21009 524
rect 19932 483 21009 517
rect 19932 475 19939 483
rect 21002 472 21009 483
rect 21061 517 21068 524
rect 22262 517 22269 527
rect 21061 483 22269 517
rect 21061 472 21068 483
rect 22262 475 22269 483
rect 22321 517 22328 527
rect 23394 517 23401 525
rect 22321 483 23401 517
rect 22321 475 22328 483
rect 23394 473 23401 483
rect 23453 517 23460 525
rect 24657 517 24664 527
rect 23453 483 24664 517
rect 23453 473 23460 483
rect 24657 475 24664 483
rect 24716 517 24723 527
rect 24716 483 25436 517
rect 24716 475 24723 483
rect 8670 379 25451 411
rect 8670 377 25436 379
rect 8449 291 25436 295
rect 8431 275 25436 291
rect 8431 272 14537 275
rect 8431 271 14171 272
rect 8431 269 11603 271
rect 8431 267 11278 269
rect 8431 215 8594 267
rect 8646 265 11278 267
rect 8646 264 8834 265
rect 8886 264 9374 265
rect 8646 230 8696 264
rect 8730 230 8788 264
rect 8822 230 8834 264
rect 8914 230 8972 264
rect 9006 230 9064 264
rect 9098 230 9156 264
rect 9208 230 9248 264
rect 9282 230 9340 264
rect 8646 215 8834 230
rect 8431 213 8834 215
rect 8886 213 9156 230
rect 8431 212 9156 213
rect 9208 213 9374 230
rect 9426 264 11278 265
rect 11330 264 11603 269
rect 11655 264 11871 271
rect 9426 230 10038 264
rect 10072 230 10130 264
rect 10164 230 10222 264
rect 10256 230 10314 264
rect 10348 230 10406 264
rect 10440 230 10498 264
rect 10532 230 10590 264
rect 10624 230 10682 264
rect 10716 230 10774 264
rect 10808 230 10996 264
rect 11030 230 11088 264
rect 11122 230 11180 264
rect 11214 230 11272 264
rect 11330 230 11364 264
rect 11398 230 11456 264
rect 11490 230 11548 264
rect 11582 230 11603 264
rect 11674 230 11732 264
rect 11766 230 11871 264
rect 9426 217 11278 230
rect 11330 219 11603 230
rect 11655 219 11871 230
rect 11923 219 12137 271
rect 12189 269 14171 271
rect 12189 219 12377 269
rect 11330 217 12377 219
rect 12429 264 14171 269
rect 12429 230 12430 264
rect 12464 230 12522 264
rect 12556 230 12614 264
rect 12648 230 12706 264
rect 12740 230 12798 264
rect 12832 230 12890 264
rect 12924 230 12982 264
rect 13016 230 13074 264
rect 13108 230 13166 264
rect 13200 230 13388 264
rect 13422 230 13480 264
rect 13514 230 13572 264
rect 13606 230 13664 264
rect 13698 230 13756 264
rect 13790 230 13848 264
rect 13882 230 13940 264
rect 13974 230 14032 264
rect 14066 230 14124 264
rect 14158 230 14171 264
rect 12429 220 14171 230
rect 14223 223 14537 272
rect 14589 223 14781 275
rect 14833 273 25436 275
rect 14833 268 17605 273
rect 14833 266 17147 268
rect 14833 264 15204 266
rect 15256 264 17147 266
rect 14854 230 14912 264
rect 14946 230 15004 264
rect 15038 230 15096 264
rect 15130 230 15188 264
rect 15256 230 15280 264
rect 15314 230 15372 264
rect 15406 230 15464 264
rect 15498 230 15556 264
rect 15590 230 15780 264
rect 15814 230 15872 264
rect 15906 230 15964 264
rect 15998 230 16056 264
rect 16090 230 16148 264
rect 16182 230 16240 264
rect 16274 230 16332 264
rect 16366 230 16424 264
rect 16458 230 16516 264
rect 16550 230 17147 264
rect 14833 223 15204 230
rect 14223 220 15204 223
rect 12429 217 15204 220
rect 9426 214 15204 217
rect 15256 216 17147 230
rect 17199 265 17605 268
rect 17199 264 17399 265
rect 17451 264 17605 265
rect 17657 271 25436 273
rect 17657 269 20228 271
rect 17657 268 20018 269
rect 17657 267 18186 268
rect 17657 264 17888 267
rect 17940 264 18186 267
rect 18238 264 20018 268
rect 20070 264 20228 269
rect 20280 269 25436 271
rect 20280 264 20579 269
rect 20631 264 20859 269
rect 20911 268 24122 269
rect 20911 264 21176 268
rect 21228 266 24122 268
rect 21228 264 22966 266
rect 23018 264 23261 266
rect 23313 264 23548 266
rect 17199 230 17214 264
rect 17248 230 17306 264
rect 17340 230 17398 264
rect 17451 230 17490 264
rect 17524 230 17582 264
rect 17657 230 17674 264
rect 17708 230 17766 264
rect 17800 230 17858 264
rect 17940 230 17950 264
rect 17984 230 18172 264
rect 18238 230 18264 264
rect 18298 230 18356 264
rect 18390 230 18448 264
rect 18482 230 18540 264
rect 18574 230 18632 264
rect 18666 230 18724 264
rect 18758 230 18816 264
rect 18850 230 18908 264
rect 18942 230 19606 264
rect 19640 230 19698 264
rect 19732 230 19790 264
rect 19824 230 19882 264
rect 19916 230 19974 264
rect 20008 230 20018 264
rect 20100 230 20158 264
rect 20192 230 20228 264
rect 20284 230 20342 264
rect 20376 230 20564 264
rect 20631 230 20656 264
rect 20690 230 20748 264
rect 20782 230 20840 264
rect 20911 230 20932 264
rect 20966 230 21024 264
rect 21058 230 21116 264
rect 21150 230 21176 264
rect 21242 230 21300 264
rect 21334 230 21996 264
rect 22030 230 22088 264
rect 22122 230 22180 264
rect 22214 230 22272 264
rect 22306 230 22364 264
rect 22398 230 22456 264
rect 22490 230 22548 264
rect 22582 230 22640 264
rect 22674 230 22732 264
rect 22766 230 22956 264
rect 23018 230 23048 264
rect 23082 230 23140 264
rect 23174 230 23232 264
rect 23313 230 23324 264
rect 23358 230 23416 264
rect 23450 230 23508 264
rect 23542 230 23548 264
rect 17199 216 17399 230
rect 15256 214 17399 216
rect 9426 213 17399 214
rect 17451 221 17605 230
rect 17657 221 17888 230
rect 17451 215 17888 221
rect 17940 216 18186 230
rect 18238 217 20018 230
rect 20070 219 20228 230
rect 20280 219 20579 230
rect 20070 217 20579 219
rect 20631 217 20859 230
rect 20911 217 21176 230
rect 18238 216 21176 217
rect 21228 216 22966 230
rect 17940 215 22966 216
rect 17451 214 22966 215
rect 23018 214 23261 230
rect 23313 214 23548 230
rect 23600 264 23838 266
rect 23634 230 23692 264
rect 23726 230 23838 264
rect 23600 214 23838 230
rect 23890 217 24122 266
rect 24174 264 25436 269
rect 24174 230 24390 264
rect 24424 230 24482 264
rect 24516 230 24574 264
rect 24608 230 24666 264
rect 24700 230 24758 264
rect 24792 230 24850 264
rect 24884 230 24942 264
rect 24976 230 25034 264
rect 25068 230 25126 264
rect 25160 230 25436 264
rect 24174 217 25436 230
rect 23890 214 25436 217
rect 17451 213 25436 214
rect 9208 212 25436 213
rect 8431 205 25436 212
rect 8449 199 25436 205
rect 9043 0 9050 52
rect 9102 0 9109 52
rect 9216 26 9285 43
rect 10126 26 10132 38
rect 9216 -8 9231 26
rect 9265 -8 10132 26
rect 9216 -23 9285 -8
rect 10126 -15 10132 -8
rect 10184 -15 10191 38
rect 10305 0 10312 52
rect 10364 0 10371 52
rect 11436 -1 11443 51
rect 11495 -1 11502 51
rect 11608 25 11678 46
rect 12518 25 12524 37
rect 10126 -16 10191 -15
rect 11608 -9 11623 25
rect 11657 -9 12524 25
rect 11608 -24 11678 -9
rect 12518 -16 12524 -9
rect 12576 -16 12583 37
rect 12697 0 12704 52
rect 12756 0 12763 52
rect 13828 -1 13835 51
rect 13887 -1 13894 51
rect 13999 37 14063 40
rect 13999 26 14064 37
rect 12518 -17 12583 -16
rect 13999 -8 14014 26
rect 14048 25 14064 26
rect 14908 25 14914 37
rect 14048 -6 14914 25
rect 14048 -8 14064 -6
rect 13999 -17 14064 -8
rect 14908 -16 14914 -6
rect 14966 -16 14973 37
rect 15088 1 15095 53
rect 15147 1 15154 53
rect 16220 0 16227 52
rect 16279 0 16286 52
rect 16392 26 16459 39
rect 17302 26 17308 38
rect 14908 -17 14973 -16
rect 16392 -8 16407 26
rect 16441 -7 17308 26
rect 16441 -8 16459 -7
rect 13999 -19 14063 -17
rect 16392 -22 16459 -8
rect 17302 -15 17308 -7
rect 17360 -15 17367 38
rect 17481 1 17488 53
rect 17540 1 17547 53
rect 18611 -1 18618 51
rect 18670 -1 18677 51
rect 18783 27 18845 42
rect 17302 -16 17367 -15
rect 18783 -7 18798 27
rect 18832 26 18845 27
rect 19694 26 19700 37
rect 18832 -6 19700 26
rect 18832 -7 18845 -6
rect 18783 -21 18845 -7
rect 19694 -16 19700 -6
rect 19752 -16 19759 37
rect 19874 1 19881 53
rect 19933 1 19940 53
rect 21003 -2 21010 50
rect 21062 -2 21069 50
rect 21175 28 21233 39
rect 22083 28 22089 37
rect 21175 27 22089 28
rect 19694 -17 19759 -16
rect 21175 -7 21190 27
rect 21224 -6 22089 27
rect 21224 -7 21233 -6
rect 21175 -19 21233 -7
rect 22083 -16 22089 -6
rect 22141 -16 22148 37
rect 22263 1 22270 53
rect 22322 1 22329 53
rect 23395 -1 23402 51
rect 23454 -1 23461 51
rect 23571 27 23623 33
rect 24478 27 24484 38
rect 23571 -7 23583 27
rect 23617 -7 24484 27
rect 23571 -13 23623 -7
rect 24478 -15 24484 -7
rect 24536 -15 24543 38
rect 24658 1 24665 53
rect 24717 1 24724 53
rect 24478 -16 24543 -15
rect 22083 -17 22148 -16
rect 8592 -151 8646 -145
rect 8592 -203 8593 -151
rect 8645 -203 8646 -151
rect 8924 -165 8931 -113
rect 8983 -117 8989 -113
rect 10525 -117 10532 -112
rect 8983 -159 10532 -117
rect 8983 -165 8989 -159
rect 10525 -164 10532 -159
rect 10584 -164 10590 -112
rect 10984 -151 11038 -145
rect 10763 -203 10769 -151
rect 10821 -203 10829 -151
rect 10984 -203 10985 -151
rect 11037 -203 11038 -151
rect 11316 -165 11323 -113
rect 11375 -117 11381 -113
rect 12917 -117 12924 -112
rect 11375 -159 12924 -117
rect 11375 -165 11381 -159
rect 12917 -164 12924 -159
rect 12976 -164 12982 -112
rect 13376 -151 13430 -145
rect 13157 -203 13163 -151
rect 13215 -203 13223 -151
rect 13376 -203 13377 -151
rect 13429 -203 13430 -151
rect 13707 -164 13714 -112
rect 13766 -116 13772 -112
rect 15308 -116 15315 -111
rect 13766 -158 15315 -116
rect 13766 -164 13772 -158
rect 15308 -163 15315 -158
rect 15367 -163 15373 -111
rect 15547 -201 15553 -149
rect 15605 -201 15613 -149
rect 15768 -151 15822 -145
rect 8592 -209 8646 -203
rect 10984 -209 11038 -203
rect 13376 -209 13430 -203
rect 15768 -203 15769 -151
rect 15821 -203 15822 -151
rect 16100 -165 16107 -113
rect 16159 -117 16165 -113
rect 17701 -117 17708 -112
rect 16159 -159 17708 -117
rect 16159 -165 16165 -159
rect 17701 -164 17708 -159
rect 17760 -164 17766 -112
rect 18159 -150 18213 -144
rect 17939 -203 17945 -151
rect 17997 -203 18005 -151
rect 18159 -202 18160 -150
rect 18212 -202 18213 -150
rect 18492 -164 18499 -112
rect 18551 -116 18557 -112
rect 20093 -116 20100 -111
rect 18551 -158 20100 -116
rect 18551 -164 18557 -158
rect 20093 -163 20100 -158
rect 20152 -163 20158 -111
rect 20331 -201 20337 -149
rect 20389 -201 20397 -149
rect 20551 -151 20605 -145
rect 15768 -209 15822 -203
rect 18159 -208 18213 -202
rect 20551 -203 20552 -151
rect 20604 -203 20605 -151
rect 20884 -164 20891 -112
rect 20943 -116 20949 -112
rect 22485 -116 22492 -111
rect 20943 -158 22492 -116
rect 20943 -164 20949 -158
rect 22485 -163 22492 -158
rect 22544 -163 22550 -111
rect 22944 -150 22998 -144
rect 22723 -203 22729 -151
rect 22781 -203 22789 -151
rect 22944 -202 22945 -150
rect 22997 -202 22998 -150
rect 23279 -164 23286 -112
rect 23338 -116 23344 -112
rect 24880 -116 24887 -111
rect 23338 -158 24887 -116
rect 23338 -164 23344 -158
rect 24880 -163 24887 -158
rect 24939 -163 24945 -111
rect 25115 -201 25121 -149
rect 25173 -201 25181 -149
rect 20551 -209 20605 -203
rect 22944 -208 22998 -202
rect 24750 -249 24780 -203
rect 8449 -251 25436 -249
rect 8449 -264 25451 -251
rect 8449 -266 19085 -264
rect 8449 -268 16433 -266
rect 8449 -271 16243 -268
rect 8449 -280 9785 -271
rect 8449 -314 8604 -280
rect 8638 -314 8696 -280
rect 8730 -314 8788 -280
rect 8822 -314 8880 -280
rect 8914 -314 8972 -280
rect 9006 -314 9064 -280
rect 9098 -314 9156 -280
rect 9190 -314 9248 -280
rect 9282 -314 9340 -280
rect 9374 -314 9785 -280
rect 8449 -323 9785 -314
rect 9837 -323 10002 -271
rect 10054 -280 10221 -271
rect 10273 -275 13619 -271
rect 10273 -280 10434 -275
rect 10486 -280 10645 -275
rect 10697 -280 12769 -275
rect 12821 -276 13619 -275
rect 12821 -280 13047 -276
rect 13099 -280 13619 -276
rect 13671 -280 13858 -271
rect 13910 -273 16243 -271
rect 13910 -280 16016 -273
rect 16068 -280 16243 -273
rect 16295 -280 16433 -268
rect 16485 -269 19085 -266
rect 16485 -272 18859 -269
rect 16485 -275 18630 -272
rect 16485 -280 16649 -275
rect 10072 -314 10130 -280
rect 10164 -314 10221 -280
rect 10273 -314 10314 -280
rect 10348 -314 10406 -280
rect 10486 -314 10498 -280
rect 10532 -314 10590 -280
rect 10624 -314 10645 -280
rect 10716 -314 10774 -280
rect 10808 -314 10996 -280
rect 11030 -314 11088 -280
rect 11122 -314 11180 -280
rect 11214 -314 11272 -280
rect 11306 -314 11364 -280
rect 11398 -314 11456 -280
rect 11490 -314 11548 -280
rect 11582 -314 11640 -280
rect 11674 -314 11732 -280
rect 11766 -314 12430 -280
rect 12464 -314 12522 -280
rect 12556 -314 12614 -280
rect 12648 -314 12706 -280
rect 12740 -314 12769 -280
rect 12832 -314 12890 -280
rect 12924 -314 12982 -280
rect 13016 -314 13047 -280
rect 13108 -314 13166 -280
rect 13200 -314 13388 -280
rect 13422 -314 13480 -280
rect 13514 -314 13572 -280
rect 13606 -314 13619 -280
rect 13698 -314 13756 -280
rect 13790 -314 13848 -280
rect 13910 -314 13940 -280
rect 13974 -314 14032 -280
rect 14066 -314 14124 -280
rect 14158 -314 14820 -280
rect 14854 -314 14912 -280
rect 14946 -314 15004 -280
rect 15038 -314 15096 -280
rect 15130 -314 15188 -280
rect 15222 -314 15280 -280
rect 15314 -314 15372 -280
rect 15406 -314 15464 -280
rect 15498 -314 15556 -280
rect 15590 -314 15780 -280
rect 15814 -314 15872 -280
rect 15906 -314 15964 -280
rect 15998 -314 16016 -280
rect 16090 -314 16148 -280
rect 16182 -314 16240 -280
rect 16295 -314 16332 -280
rect 16366 -314 16424 -280
rect 16485 -314 16516 -280
rect 16550 -314 16649 -280
rect 10054 -323 10221 -314
rect 10273 -323 10434 -314
rect 8449 -327 10434 -323
rect 10486 -327 10645 -314
rect 10697 -327 12769 -314
rect 12821 -327 13047 -314
rect 8449 -328 13047 -327
rect 13099 -323 13619 -314
rect 13671 -323 13858 -314
rect 13910 -323 16016 -314
rect 13099 -325 16016 -323
rect 16068 -320 16243 -314
rect 16295 -318 16433 -314
rect 16485 -318 16649 -314
rect 16295 -320 16649 -318
rect 16068 -325 16649 -320
rect 13099 -327 16649 -325
rect 16701 -280 18630 -275
rect 18682 -280 18859 -272
rect 18911 -280 19085 -269
rect 16701 -314 17214 -280
rect 17248 -314 17306 -280
rect 17340 -314 17398 -280
rect 17432 -314 17490 -280
rect 17524 -314 17582 -280
rect 17616 -314 17674 -280
rect 17708 -314 17766 -280
rect 17800 -314 17858 -280
rect 17892 -314 17950 -280
rect 17984 -314 18172 -280
rect 18206 -314 18264 -280
rect 18298 -314 18356 -280
rect 18390 -314 18448 -280
rect 18482 -314 18540 -280
rect 18574 -314 18630 -280
rect 18682 -314 18724 -280
rect 18758 -314 18816 -280
rect 18850 -314 18859 -280
rect 18942 -314 19085 -280
rect 16701 -324 18630 -314
rect 18682 -321 18859 -314
rect 18911 -316 19085 -314
rect 19137 -266 25451 -264
rect 19137 -272 19549 -266
rect 19137 -316 19313 -272
rect 18911 -321 19313 -316
rect 18682 -324 19313 -321
rect 19365 -318 19549 -272
rect 19601 -267 25451 -266
rect 19601 -270 24597 -267
rect 19601 -275 21680 -270
rect 19601 -280 19741 -275
rect 19793 -280 21476 -275
rect 19601 -314 19606 -280
rect 19640 -314 19698 -280
rect 19732 -314 19741 -280
rect 19824 -314 19882 -280
rect 19916 -314 19974 -280
rect 20008 -314 20066 -280
rect 20100 -314 20158 -280
rect 20192 -314 20250 -280
rect 20284 -314 20342 -280
rect 20376 -314 20564 -280
rect 20598 -314 20656 -280
rect 20690 -314 20748 -280
rect 20782 -314 20840 -280
rect 20874 -314 20932 -280
rect 20966 -314 21024 -280
rect 21058 -314 21116 -280
rect 21150 -314 21208 -280
rect 21242 -314 21300 -280
rect 21334 -314 21476 -280
rect 19601 -318 19741 -314
rect 19365 -324 19741 -318
rect 16701 -327 19741 -324
rect 19793 -327 21476 -314
rect 21528 -322 21680 -275
rect 21732 -271 24597 -270
rect 21732 -275 24403 -271
rect 21732 -322 21871 -275
rect 21528 -327 21871 -322
rect 21923 -276 22363 -275
rect 21923 -280 22073 -276
rect 22125 -280 22363 -276
rect 22415 -276 24403 -275
rect 22415 -280 22648 -276
rect 22700 -280 24403 -276
rect 24455 -280 24597 -271
rect 24649 -268 25451 -267
rect 24649 -270 25009 -268
rect 24649 -280 24786 -270
rect 24838 -280 25009 -270
rect 25061 -280 25451 -268
rect 21923 -314 21996 -280
rect 22030 -314 22073 -280
rect 22125 -314 22180 -280
rect 22214 -314 22272 -280
rect 22306 -314 22363 -280
rect 22415 -314 22456 -280
rect 22490 -314 22548 -280
rect 22582 -314 22640 -280
rect 22700 -314 22732 -280
rect 22766 -314 22956 -280
rect 22990 -314 23048 -280
rect 23082 -314 23140 -280
rect 23174 -314 23232 -280
rect 23266 -314 23324 -280
rect 23358 -314 23416 -280
rect 23450 -314 23508 -280
rect 23542 -314 23600 -280
rect 23634 -314 23692 -280
rect 23726 -314 24390 -280
rect 24455 -314 24482 -280
rect 24516 -314 24574 -280
rect 24649 -314 24666 -280
rect 24700 -314 24758 -280
rect 24838 -314 24850 -280
rect 24884 -314 24942 -280
rect 24976 -314 25009 -280
rect 25068 -314 25126 -280
rect 25160 -314 25451 -280
rect 21923 -327 22073 -314
rect 13099 -328 22073 -327
rect 22125 -327 22363 -314
rect 22415 -327 22648 -314
rect 22125 -328 22648 -327
rect 22700 -323 24403 -314
rect 24455 -319 24597 -314
rect 24649 -319 24786 -314
rect 24455 -322 24786 -319
rect 24838 -320 25009 -314
rect 25061 -320 25451 -314
rect 24838 -322 25451 -320
rect 24455 -323 25451 -322
rect 22700 -328 25451 -323
rect 8449 -337 25451 -328
rect 8449 -345 25436 -337
rect 24812 -393 24878 -392
rect 8449 -401 25357 -393
rect 8431 -414 25357 -401
rect 8431 -415 17328 -414
rect 8431 -416 11837 -415
rect 8431 -424 8840 -416
rect 8892 -419 11837 -416
rect 8892 -420 11229 -419
rect 8892 -424 9042 -420
rect 9094 -422 11229 -420
rect 9094 -423 9460 -422
rect 9094 -424 9231 -423
rect 9283 -424 9460 -423
rect 9512 -424 11229 -422
rect 11281 -422 11837 -419
rect 11281 -424 11444 -422
rect 11496 -424 11837 -422
rect 11889 -416 17328 -415
rect 11889 -417 17138 -416
rect 11889 -424 12117 -417
rect 12169 -418 17138 -417
rect 12169 -419 15093 -418
rect 12169 -424 12336 -419
rect 12388 -420 15093 -419
rect 12388 -422 14902 -420
rect 12388 -424 14157 -422
rect 14209 -424 14902 -422
rect 14954 -424 15093 -420
rect 15145 -424 17138 -418
rect 17190 -424 17328 -416
rect 17380 -415 25357 -414
rect 17380 -416 23188 -415
rect 17380 -424 17522 -416
rect 17574 -420 23188 -416
rect 17574 -424 17833 -420
rect 17885 -421 23188 -420
rect 17885 -424 20016 -421
rect 20068 -424 20220 -421
rect 20272 -423 23188 -421
rect 20272 -424 21024 -423
rect 21076 -424 21228 -423
rect 21280 -424 23188 -423
rect 23240 -417 24117 -415
rect 23240 -424 23421 -417
rect 23473 -419 23837 -417
rect 23473 -424 23628 -419
rect 23680 -424 23837 -419
rect 23889 -424 24117 -417
rect 24169 -424 25357 -415
rect 8431 -458 8604 -424
rect 8638 -458 8696 -424
rect 8730 -458 8788 -424
rect 8822 -458 8840 -424
rect 8914 -458 8972 -424
rect 9006 -458 9042 -424
rect 9098 -458 9156 -424
rect 9190 -458 9231 -424
rect 9283 -458 9340 -424
rect 9374 -458 9432 -424
rect 9512 -458 9524 -424
rect 9558 -458 9616 -424
rect 9650 -458 9708 -424
rect 9742 -458 9800 -424
rect 9834 -458 9892 -424
rect 9926 -458 9984 -424
rect 10018 -458 10076 -424
rect 10110 -458 10168 -424
rect 10202 -458 10260 -424
rect 10294 -458 10352 -424
rect 10386 -458 10444 -424
rect 10478 -458 10536 -424
rect 10570 -458 10628 -424
rect 10662 -458 10720 -424
rect 10754 -458 10812 -424
rect 10846 -458 10904 -424
rect 10938 -458 10996 -424
rect 11030 -458 11088 -424
rect 11122 -458 11180 -424
rect 11214 -458 11229 -424
rect 11306 -458 11364 -424
rect 11398 -458 11444 -424
rect 11496 -458 11548 -424
rect 11582 -458 11640 -424
rect 11674 -425 11732 -424
rect 11694 -458 11732 -425
rect 11766 -458 11824 -424
rect 11889 -458 11916 -424
rect 11950 -458 12008 -424
rect 12042 -458 12100 -424
rect 12169 -458 12192 -424
rect 12226 -458 12284 -424
rect 12318 -458 12336 -424
rect 12410 -458 12468 -424
rect 12502 -458 12560 -424
rect 12594 -458 12652 -424
rect 12686 -458 12744 -424
rect 12778 -458 12836 -424
rect 12870 -458 12928 -424
rect 12962 -458 13020 -424
rect 13054 -458 13112 -424
rect 13146 -458 13204 -424
rect 13238 -458 13296 -424
rect 13330 -458 13388 -424
rect 13422 -458 13480 -424
rect 13514 -458 13572 -424
rect 13606 -458 13664 -424
rect 13698 -458 13756 -424
rect 13790 -458 13848 -424
rect 13882 -458 13940 -424
rect 13974 -458 14032 -424
rect 14066 -458 14124 -424
rect 14209 -458 14216 -424
rect 14250 -458 14308 -424
rect 14342 -458 14400 -424
rect 14434 -458 14492 -424
rect 14526 -425 14584 -424
rect 14560 -458 14584 -425
rect 14618 -458 14676 -424
rect 14710 -427 14768 -424
rect 14749 -458 14768 -427
rect 14802 -458 14860 -424
rect 14894 -458 14902 -424
rect 14986 -458 15044 -424
rect 15078 -458 15093 -424
rect 15170 -458 15228 -424
rect 15262 -458 15320 -424
rect 15354 -458 15412 -424
rect 15446 -458 15504 -424
rect 15538 -458 15596 -424
rect 15630 -458 15688 -424
rect 15722 -458 15780 -424
rect 15814 -458 15872 -424
rect 15906 -458 15964 -424
rect 15998 -458 16056 -424
rect 16090 -458 16148 -424
rect 16182 -458 16240 -424
rect 16274 -458 16332 -424
rect 16366 -458 16424 -424
rect 16458 -458 16516 -424
rect 16550 -458 16608 -424
rect 16642 -458 16700 -424
rect 16734 -458 16792 -424
rect 16826 -458 16884 -424
rect 16918 -458 16976 -424
rect 17010 -458 17068 -424
rect 17102 -458 17138 -424
rect 17194 -458 17252 -424
rect 17286 -458 17328 -424
rect 17380 -458 17436 -424
rect 17470 -458 17522 -424
rect 17574 -458 17620 -424
rect 17654 -458 17712 -424
rect 17746 -458 17804 -424
rect 17885 -458 17896 -424
rect 17930 -458 17988 -424
rect 18022 -458 18080 -424
rect 18114 -458 18172 -424
rect 18206 -458 18264 -424
rect 18298 -458 18356 -424
rect 18390 -458 18448 -424
rect 18482 -458 18540 -424
rect 18574 -458 18632 -424
rect 18666 -458 18724 -424
rect 18758 -458 18816 -424
rect 18850 -458 18908 -424
rect 18942 -458 19000 -424
rect 19034 -458 19092 -424
rect 19126 -458 19184 -424
rect 19218 -458 19276 -424
rect 19310 -458 19368 -424
rect 19402 -458 19460 -424
rect 19494 -458 19552 -424
rect 19586 -458 19644 -424
rect 19678 -458 19736 -424
rect 19770 -458 19828 -424
rect 19862 -458 19920 -424
rect 19954 -458 20012 -424
rect 20068 -458 20104 -424
rect 20138 -458 20196 -424
rect 20272 -458 20288 -424
rect 20322 -458 20380 -424
rect 20414 -458 20472 -424
rect 20506 -458 20564 -424
rect 20598 -458 20656 -424
rect 20690 -458 20748 -424
rect 20782 -425 20840 -424
rect 20782 -458 20785 -425
rect 8431 -468 8840 -458
rect 8892 -468 9042 -458
rect 8431 -472 9042 -468
rect 9094 -472 9231 -458
rect 8431 -475 9231 -472
rect 9283 -474 9460 -458
rect 9512 -471 11229 -458
rect 11281 -471 11444 -458
rect 9512 -474 11444 -471
rect 11496 -474 11642 -458
rect 9283 -475 11642 -474
rect 8431 -477 11642 -475
rect 11694 -467 11837 -458
rect 11889 -467 12117 -458
rect 11694 -469 12117 -467
rect 12169 -469 12336 -458
rect 11694 -471 12336 -469
rect 12388 -471 14157 -458
rect 11694 -474 14157 -471
rect 14209 -474 14508 -458
rect 11694 -477 14508 -474
rect 14560 -477 14697 -458
rect 8431 -479 14697 -477
rect 14749 -472 14902 -458
rect 14954 -470 15093 -458
rect 15145 -468 17138 -458
rect 17190 -466 17328 -458
rect 17380 -466 17522 -458
rect 17190 -468 17522 -466
rect 17574 -468 17833 -458
rect 15145 -470 17833 -468
rect 14954 -472 17833 -470
rect 17885 -472 20016 -458
rect 14749 -473 20016 -472
rect 20068 -473 20220 -458
rect 20272 -473 20785 -458
rect 14749 -477 20785 -473
rect 20837 -458 20840 -425
rect 20874 -458 20932 -424
rect 20966 -458 21024 -424
rect 21076 -458 21116 -424
rect 21150 -458 21208 -424
rect 21280 -458 21300 -424
rect 21334 -458 21392 -424
rect 21426 -458 21484 -424
rect 21518 -458 21576 -424
rect 21610 -458 21668 -424
rect 21702 -458 21760 -424
rect 21794 -458 21852 -424
rect 21886 -458 21944 -424
rect 21978 -458 22036 -424
rect 22070 -458 22128 -424
rect 22162 -458 22220 -424
rect 22254 -458 22312 -424
rect 22346 -458 22404 -424
rect 22438 -458 22496 -424
rect 22530 -458 22588 -424
rect 22622 -458 22680 -424
rect 22714 -458 22772 -424
rect 22806 -458 22864 -424
rect 22898 -458 22956 -424
rect 22990 -458 23048 -424
rect 23082 -458 23140 -424
rect 23174 -458 23188 -424
rect 23266 -458 23324 -424
rect 23358 -458 23416 -424
rect 23473 -458 23508 -424
rect 23542 -458 23600 -424
rect 23680 -458 23692 -424
rect 23726 -458 23784 -424
rect 23818 -458 23837 -424
rect 23910 -458 23968 -424
rect 24002 -458 24060 -424
rect 24094 -458 24117 -424
rect 24186 -458 24244 -424
rect 24278 -458 24336 -424
rect 24370 -458 24428 -424
rect 24462 -458 24520 -424
rect 24554 -458 24612 -424
rect 24646 -458 24704 -424
rect 24738 -458 24796 -424
rect 24830 -458 24888 -424
rect 24922 -458 24980 -424
rect 25014 -458 25072 -424
rect 25106 -458 25164 -424
rect 25198 -458 25256 -424
rect 25290 -458 25357 -424
rect 20837 -475 21024 -458
rect 21076 -475 21228 -458
rect 21280 -467 23188 -458
rect 23240 -467 23421 -458
rect 21280 -469 23421 -467
rect 23473 -469 23628 -458
rect 21280 -471 23628 -469
rect 23680 -469 23837 -458
rect 23889 -467 24117 -458
rect 24169 -467 25357 -458
rect 23889 -469 25357 -467
rect 23680 -471 25357 -469
rect 21280 -475 25357 -471
rect 20837 -477 25357 -475
rect 14749 -479 25357 -477
rect 8431 -487 25357 -479
rect 8449 -489 25357 -487
rect 10899 -523 10951 -517
rect 10899 -581 10951 -575
rect 13291 -523 13343 -517
rect 13291 -581 13343 -575
rect 15683 -523 15735 -517
rect 15683 -581 15735 -575
rect 18075 -523 18127 -517
rect 18075 -581 18127 -575
rect 20467 -523 20519 -517
rect 20467 -581 20519 -575
rect 22859 -523 22911 -517
rect 22859 -581 22911 -575
rect 25251 -523 25303 -517
rect 25251 -581 25303 -575
rect 8776 -594 8834 -588
rect 8776 -628 8788 -594
rect 8822 -597 8834 -594
rect 9052 -594 9110 -588
rect 9052 -597 9064 -594
rect 8822 -625 9064 -597
rect 8822 -628 8834 -625
rect 8776 -634 8834 -628
rect 9052 -628 9064 -625
rect 9098 -597 9110 -594
rect 9788 -594 9846 -588
rect 11168 -594 11226 -588
rect 9788 -597 9800 -594
rect 9098 -625 9800 -597
rect 9098 -628 9110 -625
rect 9052 -634 9110 -628
rect 9788 -628 9800 -625
rect 9834 -628 9846 -594
rect 9788 -634 9846 -628
rect 10617 -600 10669 -594
rect 11168 -628 11180 -594
rect 11214 -597 11226 -594
rect 11444 -594 11502 -588
rect 11444 -597 11456 -594
rect 11214 -625 11456 -597
rect 11214 -628 11226 -625
rect 11168 -634 11226 -628
rect 11444 -628 11456 -625
rect 11490 -597 11502 -594
rect 12180 -594 12238 -588
rect 12180 -597 12192 -594
rect 11490 -625 12192 -597
rect 11490 -628 11502 -625
rect 11444 -634 11502 -628
rect 12180 -628 12192 -625
rect 12226 -628 12238 -594
rect 12180 -634 12238 -628
rect 13009 -599 13061 -593
rect 9696 -662 9754 -656
rect 8592 -696 8646 -690
rect 8592 -748 8593 -696
rect 8645 -748 8646 -696
rect 8926 -724 8932 -671
rect 8984 -724 8991 -671
rect 9696 -696 9708 -662
rect 9742 -665 9754 -662
rect 10334 -662 10392 -656
rect 10617 -658 10669 -652
rect 13560 -594 13618 -588
rect 13560 -628 13572 -594
rect 13606 -597 13618 -594
rect 13836 -594 13894 -588
rect 13836 -597 13848 -594
rect 13606 -625 13848 -597
rect 13606 -628 13618 -625
rect 13560 -634 13618 -628
rect 13836 -628 13848 -625
rect 13882 -597 13894 -594
rect 14572 -594 14630 -588
rect 14572 -597 14584 -594
rect 13882 -625 14584 -597
rect 13882 -628 13894 -625
rect 13836 -634 13894 -628
rect 14572 -628 14584 -625
rect 14618 -628 14630 -594
rect 14572 -634 14630 -628
rect 15400 -599 15452 -593
rect 10334 -665 10346 -662
rect 9742 -693 10346 -665
rect 9742 -696 9754 -693
rect 9696 -702 9754 -696
rect 10334 -696 10346 -693
rect 10380 -696 10392 -662
rect 12088 -662 12146 -656
rect 10334 -702 10392 -696
rect 10984 -696 11038 -690
rect 8926 -725 8991 -724
rect 9788 -730 9846 -724
rect 9788 -733 9800 -730
rect 8592 -754 8646 -748
rect 9159 -761 9800 -733
rect 9159 -792 9202 -761
rect 9788 -764 9800 -761
rect 9834 -764 9846 -730
rect 10984 -748 10985 -696
rect 11037 -748 11038 -696
rect 11318 -724 11324 -671
rect 11376 -724 11383 -671
rect 12088 -696 12100 -662
rect 12134 -665 12146 -662
rect 12726 -662 12784 -656
rect 13009 -657 13061 -651
rect 15952 -594 16010 -588
rect 15952 -628 15964 -594
rect 15998 -597 16010 -594
rect 16228 -594 16286 -588
rect 16228 -597 16240 -594
rect 15998 -625 16240 -597
rect 15998 -628 16010 -625
rect 15952 -634 16010 -628
rect 16228 -628 16240 -625
rect 16274 -597 16286 -594
rect 16964 -594 17022 -588
rect 16964 -597 16976 -594
rect 16274 -625 16976 -597
rect 16274 -628 16286 -625
rect 16228 -634 16286 -628
rect 16964 -628 16976 -625
rect 17010 -628 17022 -594
rect 16964 -634 17022 -628
rect 17793 -598 17845 -592
rect 12726 -665 12738 -662
rect 12134 -693 12738 -665
rect 12134 -696 12146 -693
rect 12088 -702 12146 -696
rect 12726 -696 12738 -693
rect 12772 -696 12784 -662
rect 14480 -662 14538 -656
rect 12726 -702 12784 -696
rect 13376 -696 13430 -690
rect 11318 -725 11383 -724
rect 12180 -730 12238 -724
rect 12180 -733 12192 -730
rect 10984 -754 11038 -748
rect 9788 -770 9846 -764
rect 11551 -761 12192 -733
rect 8685 -798 8743 -792
rect 8685 -832 8697 -798
rect 8731 -801 8743 -798
rect 9144 -798 9202 -792
rect 9144 -801 9156 -798
rect 8731 -829 9156 -801
rect 8731 -832 8743 -829
rect 8685 -838 8743 -832
rect 9144 -832 9156 -829
rect 9190 -832 9202 -798
rect 9144 -838 9202 -832
rect 9328 -798 9386 -792
rect 9328 -832 9340 -798
rect 9374 -801 9386 -798
rect 9599 -795 9653 -789
rect 11551 -792 11594 -761
rect 12180 -764 12192 -761
rect 12226 -764 12238 -730
rect 13376 -748 13377 -696
rect 13429 -748 13430 -696
rect 13710 -723 13716 -670
rect 13768 -723 13775 -670
rect 14480 -696 14492 -662
rect 14526 -665 14538 -662
rect 15118 -662 15176 -656
rect 15400 -657 15452 -651
rect 18344 -594 18402 -588
rect 18344 -628 18356 -594
rect 18390 -597 18402 -594
rect 18620 -594 18678 -588
rect 18620 -597 18632 -594
rect 18390 -625 18632 -597
rect 18390 -628 18402 -625
rect 18344 -634 18402 -628
rect 18620 -628 18632 -625
rect 18666 -597 18678 -594
rect 19356 -594 19414 -588
rect 19356 -597 19368 -594
rect 18666 -625 19368 -597
rect 18666 -628 18678 -625
rect 18620 -634 18678 -628
rect 19356 -628 19368 -625
rect 19402 -628 19414 -594
rect 19356 -634 19414 -628
rect 20184 -599 20236 -593
rect 17793 -656 17845 -650
rect 20736 -594 20794 -588
rect 20736 -628 20748 -594
rect 20782 -597 20794 -594
rect 21012 -594 21070 -588
rect 21012 -597 21024 -594
rect 20782 -625 21024 -597
rect 20782 -628 20794 -625
rect 20736 -634 20794 -628
rect 21012 -628 21024 -625
rect 21058 -597 21070 -594
rect 21748 -594 21806 -588
rect 23128 -594 23186 -588
rect 21748 -597 21760 -594
rect 21058 -625 21760 -597
rect 21058 -628 21070 -625
rect 21012 -634 21070 -628
rect 21748 -628 21760 -625
rect 21794 -628 21806 -594
rect 21748 -634 21806 -628
rect 22577 -600 22629 -594
rect 15118 -665 15130 -662
rect 14526 -693 15130 -665
rect 14526 -696 14538 -693
rect 14480 -702 14538 -696
rect 15118 -696 15130 -693
rect 15164 -696 15176 -662
rect 16872 -662 16930 -656
rect 15118 -702 15176 -696
rect 15768 -696 15822 -690
rect 13710 -724 13775 -723
rect 14572 -730 14630 -724
rect 14572 -733 14584 -730
rect 13376 -754 13430 -748
rect 12180 -770 12238 -764
rect 13943 -761 14584 -733
rect 9599 -801 9600 -795
rect 9374 -829 9600 -801
rect 9374 -832 9386 -829
rect 9328 -838 9386 -832
rect 9599 -847 9600 -829
rect 9652 -801 9653 -795
rect 10078 -798 10136 -792
rect 10078 -801 10090 -798
rect 9652 -829 10090 -801
rect 9652 -847 9653 -829
rect 10078 -832 10090 -829
rect 10124 -832 10136 -798
rect 10078 -838 10136 -832
rect 11077 -798 11135 -792
rect 11077 -832 11089 -798
rect 11123 -801 11135 -798
rect 11536 -798 11594 -792
rect 11536 -801 11548 -798
rect 11123 -829 11548 -801
rect 11123 -832 11135 -829
rect 11077 -838 11135 -832
rect 11536 -832 11548 -829
rect 11582 -832 11594 -798
rect 11536 -838 11594 -832
rect 11720 -798 11778 -792
rect 11720 -832 11732 -798
rect 11766 -801 11778 -798
rect 11992 -795 12046 -789
rect 13943 -792 13986 -761
rect 14572 -764 14584 -761
rect 14618 -764 14630 -730
rect 15768 -748 15769 -696
rect 15821 -748 15822 -696
rect 16102 -723 16108 -670
rect 16160 -723 16167 -670
rect 16872 -696 16884 -662
rect 16918 -665 16930 -662
rect 17510 -662 17568 -656
rect 17510 -665 17522 -662
rect 16918 -693 17522 -665
rect 16918 -696 16930 -693
rect 16872 -702 16930 -696
rect 17510 -696 17522 -693
rect 17556 -696 17568 -662
rect 19264 -662 19322 -656
rect 17510 -702 17568 -696
rect 18159 -695 18213 -689
rect 16102 -724 16167 -723
rect 16964 -730 17022 -724
rect 16964 -733 16976 -730
rect 15768 -754 15822 -748
rect 14572 -770 14630 -764
rect 16335 -761 16976 -733
rect 11992 -801 11993 -795
rect 11766 -829 11993 -801
rect 11766 -832 11778 -829
rect 11720 -838 11778 -832
rect 9599 -853 9653 -847
rect 11992 -847 11993 -829
rect 12045 -801 12046 -795
rect 12470 -798 12528 -792
rect 12470 -801 12482 -798
rect 12045 -829 12482 -801
rect 12045 -847 12046 -829
rect 12470 -832 12482 -829
rect 12516 -832 12528 -798
rect 12470 -838 12528 -832
rect 13469 -798 13527 -792
rect 13469 -832 13481 -798
rect 13515 -801 13527 -798
rect 13928 -798 13986 -792
rect 13928 -801 13940 -798
rect 13515 -829 13940 -801
rect 13515 -832 13527 -829
rect 13469 -838 13527 -832
rect 13928 -832 13940 -829
rect 13974 -832 13986 -798
rect 13928 -838 13986 -832
rect 14112 -798 14170 -792
rect 14112 -832 14124 -798
rect 14158 -801 14170 -798
rect 14384 -795 14438 -789
rect 16335 -792 16378 -761
rect 16964 -764 16976 -761
rect 17010 -764 17022 -730
rect 18159 -747 18160 -695
rect 18212 -747 18213 -695
rect 18494 -724 18500 -671
rect 18552 -724 18559 -671
rect 19264 -696 19276 -662
rect 19310 -665 19322 -662
rect 19902 -662 19960 -656
rect 20184 -657 20236 -651
rect 23128 -628 23140 -594
rect 23174 -597 23186 -594
rect 23404 -594 23462 -588
rect 23404 -597 23416 -594
rect 23174 -625 23416 -597
rect 23174 -628 23186 -625
rect 23128 -634 23186 -628
rect 23404 -628 23416 -625
rect 23450 -597 23462 -594
rect 24140 -594 24198 -588
rect 24140 -597 24152 -594
rect 23450 -625 24152 -597
rect 23450 -628 23462 -625
rect 23404 -634 23462 -628
rect 24140 -628 24152 -625
rect 24186 -628 24198 -594
rect 24140 -634 24198 -628
rect 24970 -598 25022 -592
rect 19902 -665 19914 -662
rect 19310 -693 19914 -665
rect 19310 -696 19322 -693
rect 19264 -702 19322 -696
rect 19902 -696 19914 -693
rect 19948 -696 19960 -662
rect 21656 -662 21714 -656
rect 19902 -702 19960 -696
rect 20551 -696 20605 -690
rect 18494 -725 18559 -724
rect 19356 -730 19414 -724
rect 19356 -733 19368 -730
rect 18159 -753 18213 -747
rect 16964 -770 17022 -764
rect 18727 -761 19368 -733
rect 14384 -801 14385 -795
rect 14158 -829 14385 -801
rect 14158 -832 14170 -829
rect 14112 -838 14170 -832
rect 11992 -853 12046 -847
rect 14384 -847 14385 -829
rect 14437 -801 14438 -795
rect 14862 -798 14920 -792
rect 14862 -801 14874 -798
rect 14437 -829 14874 -801
rect 14437 -847 14438 -829
rect 14862 -832 14874 -829
rect 14908 -832 14920 -798
rect 14862 -838 14920 -832
rect 15861 -798 15919 -792
rect 15861 -832 15873 -798
rect 15907 -801 15919 -798
rect 16320 -798 16378 -792
rect 16320 -801 16332 -798
rect 15907 -829 16332 -801
rect 15907 -832 15919 -829
rect 15861 -838 15919 -832
rect 16320 -832 16332 -829
rect 16366 -832 16378 -798
rect 16320 -838 16378 -832
rect 16504 -798 16562 -792
rect 16504 -832 16516 -798
rect 16550 -801 16562 -798
rect 16776 -795 16830 -789
rect 18727 -792 18770 -761
rect 19356 -764 19368 -761
rect 19402 -764 19414 -730
rect 20551 -748 20552 -696
rect 20604 -748 20605 -696
rect 20886 -723 20892 -670
rect 20944 -723 20951 -670
rect 21656 -696 21668 -662
rect 21702 -665 21714 -662
rect 22294 -662 22352 -656
rect 22577 -658 22629 -652
rect 24970 -656 25022 -650
rect 22294 -665 22306 -662
rect 21702 -693 22306 -665
rect 21702 -696 21714 -693
rect 21656 -702 21714 -696
rect 22294 -696 22306 -693
rect 22340 -696 22352 -662
rect 24048 -662 24106 -656
rect 22294 -702 22352 -696
rect 22944 -695 22998 -689
rect 20886 -724 20951 -723
rect 21748 -730 21806 -724
rect 21748 -733 21760 -730
rect 20551 -754 20605 -748
rect 19356 -770 19414 -764
rect 21119 -761 21760 -733
rect 16776 -801 16777 -795
rect 16550 -829 16777 -801
rect 16550 -832 16562 -829
rect 16504 -838 16562 -832
rect 14384 -853 14438 -847
rect 16776 -847 16777 -829
rect 16829 -801 16830 -795
rect 17254 -798 17312 -792
rect 17254 -801 17266 -798
rect 16829 -829 17266 -801
rect 16829 -847 16830 -829
rect 17254 -832 17266 -829
rect 17300 -832 17312 -798
rect 17254 -838 17312 -832
rect 18253 -798 18311 -792
rect 18253 -832 18265 -798
rect 18299 -801 18311 -798
rect 18712 -798 18770 -792
rect 18712 -801 18724 -798
rect 18299 -829 18724 -801
rect 18299 -832 18311 -829
rect 18253 -838 18311 -832
rect 18712 -832 18724 -829
rect 18758 -832 18770 -798
rect 18712 -838 18770 -832
rect 18896 -798 18954 -792
rect 18896 -832 18908 -798
rect 18942 -801 18954 -798
rect 19167 -795 19221 -789
rect 21119 -792 21162 -761
rect 21748 -764 21760 -761
rect 21794 -764 21806 -730
rect 22944 -747 22945 -695
rect 22997 -747 22998 -695
rect 23279 -724 23285 -671
rect 23337 -724 23344 -671
rect 24048 -696 24060 -662
rect 24094 -665 24106 -662
rect 24686 -662 24744 -656
rect 24686 -665 24698 -662
rect 24094 -693 24698 -665
rect 24094 -696 24106 -693
rect 24048 -702 24106 -696
rect 24686 -696 24698 -693
rect 24732 -696 24744 -662
rect 24686 -702 24744 -696
rect 23279 -725 23344 -724
rect 24140 -730 24198 -724
rect 24140 -733 24152 -730
rect 22944 -753 22998 -747
rect 21748 -770 21806 -764
rect 23511 -761 24152 -733
rect 19167 -801 19168 -795
rect 18942 -829 19168 -801
rect 18942 -832 18954 -829
rect 18896 -838 18954 -832
rect 16776 -853 16830 -847
rect 19167 -847 19168 -829
rect 19220 -801 19221 -795
rect 19646 -798 19704 -792
rect 19646 -801 19658 -798
rect 19220 -829 19658 -801
rect 19220 -847 19221 -829
rect 19646 -832 19658 -829
rect 19692 -832 19704 -798
rect 19646 -838 19704 -832
rect 20645 -798 20703 -792
rect 20645 -832 20657 -798
rect 20691 -801 20703 -798
rect 21104 -798 21162 -792
rect 21104 -801 21116 -798
rect 20691 -829 21116 -801
rect 20691 -832 20703 -829
rect 20645 -838 20703 -832
rect 21104 -832 21116 -829
rect 21150 -832 21162 -798
rect 21104 -838 21162 -832
rect 21288 -798 21346 -792
rect 21288 -832 21300 -798
rect 21334 -801 21346 -798
rect 21559 -795 21613 -789
rect 23511 -792 23554 -761
rect 24140 -764 24152 -761
rect 24186 -764 24198 -730
rect 24140 -770 24198 -764
rect 21559 -801 21560 -795
rect 21334 -829 21560 -801
rect 21334 -832 21346 -829
rect 21288 -838 21346 -832
rect 19167 -855 19221 -847
rect 21559 -847 21560 -829
rect 21612 -801 21613 -795
rect 22038 -798 22096 -792
rect 22038 -801 22050 -798
rect 21612 -829 22050 -801
rect 21612 -847 21613 -829
rect 22038 -832 22050 -829
rect 22084 -832 22096 -798
rect 22038 -838 22096 -832
rect 23037 -798 23095 -792
rect 23037 -832 23049 -798
rect 23083 -801 23095 -798
rect 23496 -798 23554 -792
rect 23496 -801 23508 -798
rect 23083 -829 23508 -801
rect 23083 -832 23095 -829
rect 23037 -838 23095 -832
rect 23496 -832 23508 -829
rect 23542 -832 23554 -798
rect 23496 -838 23554 -832
rect 23680 -798 23738 -792
rect 23680 -832 23692 -798
rect 23726 -801 23738 -798
rect 23951 -795 24005 -789
rect 23951 -801 23952 -795
rect 23726 -829 23952 -801
rect 23726 -832 23738 -829
rect 23680 -838 23738 -832
rect 21559 -853 21613 -847
rect 23951 -847 23952 -829
rect 24004 -801 24005 -795
rect 24430 -798 24488 -792
rect 24430 -801 24442 -798
rect 24004 -829 24442 -801
rect 24004 -847 24005 -829
rect 24430 -832 24442 -829
rect 24476 -832 24488 -798
rect 24430 -838 24488 -832
rect 23951 -853 24005 -847
rect 25391 -937 25436 -933
rect 8449 -953 25451 -937
rect 8449 -965 9996 -953
rect 8449 -968 9767 -965
rect 9819 -968 9996 -965
rect 10048 -954 25451 -953
rect 10048 -956 13613 -954
rect 10048 -959 13283 -956
rect 10048 -963 10407 -959
rect 10048 -968 10215 -963
rect 10267 -968 10407 -963
rect 10459 -961 13283 -959
rect 10459 -968 10901 -961
rect 10953 -962 13283 -961
rect 10953 -968 12693 -962
rect 12745 -964 13283 -962
rect 12745 -968 13086 -964
rect 13138 -968 13283 -964
rect 13335 -968 13613 -956
rect 13665 -968 13809 -954
rect 13861 -956 16644 -954
rect 13861 -957 16223 -956
rect 13861 -961 16017 -957
rect 13861 -968 15716 -961
rect 15768 -968 16017 -961
rect 16069 -968 16223 -957
rect 16275 -960 16644 -956
rect 16275 -968 16433 -960
rect 16485 -968 16644 -960
rect 8449 -1002 8604 -968
rect 8638 -1002 8696 -968
rect 8730 -1002 8788 -968
rect 8822 -1002 8880 -968
rect 8914 -1002 8972 -968
rect 9006 -1002 9064 -968
rect 9098 -1002 9156 -968
rect 9190 -1002 9248 -968
rect 9282 -1002 9340 -968
rect 9374 -1002 9432 -968
rect 9466 -1002 9524 -968
rect 9558 -1002 9616 -968
rect 9650 -1002 9708 -968
rect 9742 -1002 9767 -968
rect 9834 -1002 9892 -968
rect 9926 -1002 9984 -968
rect 10048 -1002 10076 -968
rect 10110 -1002 10168 -968
rect 10202 -1002 10215 -968
rect 10294 -1002 10352 -968
rect 10386 -1002 10407 -968
rect 10478 -1002 10536 -968
rect 10570 -1002 10628 -968
rect 10662 -1002 10720 -968
rect 10754 -1002 10812 -968
rect 10846 -1002 10901 -968
rect 10953 -1002 10996 -968
rect 11030 -1002 11088 -968
rect 11122 -1002 11180 -968
rect 11214 -1002 11272 -968
rect 11306 -1002 11364 -968
rect 11398 -1002 11456 -968
rect 11490 -1002 11548 -968
rect 11582 -1002 11640 -968
rect 11674 -1002 11732 -968
rect 11766 -1002 11824 -968
rect 11858 -1002 11916 -968
rect 11950 -1002 12008 -968
rect 12042 -1002 12100 -968
rect 12134 -1002 12192 -968
rect 12226 -1002 12284 -968
rect 12318 -1002 12376 -968
rect 12410 -1002 12468 -968
rect 12502 -1002 12560 -968
rect 12594 -1002 12652 -968
rect 12686 -1002 12693 -968
rect 12778 -1002 12836 -968
rect 12870 -1002 12928 -968
rect 12962 -1002 13020 -968
rect 13054 -1002 13086 -968
rect 13146 -1002 13204 -968
rect 13238 -1002 13283 -968
rect 13335 -1002 13388 -968
rect 13422 -1002 13480 -968
rect 13514 -1002 13572 -968
rect 13606 -1002 13613 -968
rect 13698 -1002 13756 -968
rect 13790 -1002 13809 -968
rect 13882 -1002 13940 -968
rect 13974 -1002 14032 -968
rect 14066 -1002 14124 -968
rect 14158 -1002 14216 -968
rect 14250 -1002 14308 -968
rect 14342 -1002 14400 -968
rect 14434 -1002 14492 -968
rect 14526 -1002 14584 -968
rect 14618 -1002 14676 -968
rect 14710 -1002 14768 -968
rect 14802 -1002 14860 -968
rect 14894 -1002 14952 -968
rect 14986 -1002 15044 -968
rect 15078 -1002 15136 -968
rect 15170 -1002 15228 -968
rect 15262 -1002 15320 -968
rect 15354 -1002 15412 -968
rect 15446 -1002 15504 -968
rect 15538 -1002 15596 -968
rect 15630 -1002 15688 -968
rect 15768 -1002 15780 -968
rect 15814 -1002 15872 -968
rect 15906 -1002 15964 -968
rect 15998 -1002 16017 -968
rect 16090 -1002 16148 -968
rect 16182 -1002 16223 -968
rect 16275 -1002 16332 -968
rect 16366 -1002 16424 -968
rect 16485 -1002 16516 -968
rect 16550 -1002 16608 -968
rect 16642 -1002 16644 -968
rect 8449 -1017 9767 -1002
rect 9819 -1005 9996 -1002
rect 10048 -1005 10215 -1002
rect 9819 -1015 10215 -1005
rect 10267 -1011 10407 -1002
rect 10459 -1011 10901 -1002
rect 10267 -1013 10901 -1011
rect 10953 -1013 12693 -1002
rect 10267 -1014 12693 -1013
rect 12745 -1014 13086 -1002
rect 10267 -1015 13086 -1014
rect 9819 -1016 13086 -1015
rect 13138 -1008 13283 -1002
rect 13335 -1006 13613 -1002
rect 13665 -1006 13809 -1002
rect 13861 -1006 15716 -1002
rect 13335 -1008 15716 -1006
rect 13138 -1013 15716 -1008
rect 15768 -1009 16017 -1002
rect 16069 -1008 16223 -1002
rect 16275 -1008 16433 -1002
rect 16069 -1009 16433 -1008
rect 15768 -1012 16433 -1009
rect 16485 -1006 16644 -1002
rect 16696 -957 19543 -954
rect 16696 -958 19302 -957
rect 16696 -965 18781 -958
rect 16696 -968 18524 -965
rect 18576 -968 18781 -965
rect 18833 -962 19302 -958
rect 18833 -968 19031 -962
rect 19083 -968 19302 -962
rect 19354 -968 19543 -957
rect 19595 -955 25451 -954
rect 19595 -957 24791 -955
rect 19595 -958 24596 -957
rect 19595 -968 19768 -958
rect 19820 -959 24596 -958
rect 19820 -960 21676 -959
rect 19820 -968 21475 -960
rect 21527 -968 21676 -960
rect 21728 -963 22101 -959
rect 21728 -968 21894 -963
rect 21946 -968 22101 -963
rect 22153 -960 24596 -959
rect 22153 -968 22306 -960
rect 22358 -964 24405 -960
rect 22358 -968 22653 -964
rect 22705 -968 24405 -964
rect 24457 -968 24596 -960
rect 24648 -968 24791 -957
rect 24843 -960 25451 -955
rect 24843 -968 25238 -960
rect 16696 -1002 16700 -968
rect 16734 -1002 16792 -968
rect 16826 -1002 16884 -968
rect 16918 -1002 16976 -968
rect 17010 -1002 17068 -968
rect 17102 -1002 17160 -968
rect 17194 -1002 17252 -968
rect 17286 -1002 17344 -968
rect 17378 -1002 17436 -968
rect 17470 -1002 17528 -968
rect 17562 -1002 17620 -968
rect 17654 -1002 17712 -968
rect 17746 -1002 17804 -968
rect 17838 -1002 17896 -968
rect 17930 -1002 17988 -968
rect 18022 -1002 18080 -968
rect 18114 -1002 18172 -968
rect 18206 -1002 18264 -968
rect 18298 -1002 18356 -968
rect 18390 -1002 18448 -968
rect 18482 -1002 18524 -968
rect 18576 -1002 18632 -968
rect 18666 -1002 18724 -968
rect 18758 -1002 18781 -968
rect 18850 -1002 18908 -968
rect 18942 -1002 19000 -968
rect 19083 -1002 19092 -968
rect 19126 -1002 19184 -968
rect 19218 -1002 19276 -968
rect 19354 -1002 19368 -968
rect 19402 -1002 19460 -968
rect 19494 -1002 19543 -968
rect 19595 -1002 19644 -968
rect 19678 -1002 19736 -968
rect 19820 -1002 19828 -968
rect 19862 -1002 19920 -968
rect 19954 -1002 20012 -968
rect 20046 -1002 20104 -968
rect 20138 -1002 20196 -968
rect 20230 -1002 20288 -968
rect 20322 -1002 20380 -968
rect 20414 -1002 20472 -968
rect 20506 -1002 20564 -968
rect 20598 -1002 20656 -968
rect 20690 -1002 20748 -968
rect 20782 -1002 20840 -968
rect 20874 -1002 20932 -968
rect 20966 -1002 21024 -968
rect 21058 -1002 21116 -968
rect 21150 -1002 21208 -968
rect 21242 -1002 21300 -968
rect 21334 -1002 21392 -968
rect 21426 -1002 21475 -968
rect 21527 -1002 21576 -968
rect 21610 -1002 21668 -968
rect 21728 -1002 21760 -968
rect 21794 -1002 21852 -968
rect 21886 -1002 21894 -968
rect 21978 -1002 22036 -968
rect 22070 -1002 22101 -968
rect 22162 -1002 22220 -968
rect 22254 -1002 22306 -968
rect 22358 -1002 22404 -968
rect 22438 -1002 22496 -968
rect 22530 -1002 22588 -968
rect 22622 -1002 22653 -968
rect 22714 -1002 22772 -968
rect 22806 -1002 22864 -968
rect 22898 -1002 22956 -968
rect 22990 -1002 23048 -968
rect 23082 -1002 23140 -968
rect 23174 -1002 23232 -968
rect 23266 -1002 23324 -968
rect 23358 -1002 23416 -968
rect 23450 -1002 23508 -968
rect 23542 -1002 23600 -968
rect 23634 -1002 23692 -968
rect 23726 -1002 23784 -968
rect 23818 -1002 23876 -968
rect 23910 -1002 23968 -968
rect 24002 -1002 24060 -968
rect 24094 -1002 24152 -968
rect 24186 -1002 24244 -968
rect 24278 -1002 24336 -968
rect 24370 -1002 24405 -968
rect 24462 -1002 24520 -968
rect 24554 -1002 24596 -968
rect 24648 -1002 24704 -968
rect 24738 -1002 24791 -968
rect 24843 -1002 24888 -968
rect 24922 -1002 24980 -968
rect 25014 -1002 25072 -968
rect 25106 -1002 25164 -968
rect 25198 -1002 25238 -968
rect 16696 -1006 18524 -1002
rect 16485 -1012 18524 -1006
rect 15768 -1013 18524 -1012
rect 13138 -1016 18524 -1013
rect 9819 -1017 18524 -1016
rect 18576 -1010 18781 -1002
rect 18833 -1010 19031 -1002
rect 18576 -1014 19031 -1010
rect 19083 -1009 19302 -1002
rect 19354 -1006 19543 -1002
rect 19595 -1006 19768 -1002
rect 19354 -1009 19768 -1006
rect 19083 -1010 19768 -1009
rect 19820 -1010 21475 -1002
rect 19083 -1012 21475 -1010
rect 21527 -1011 21676 -1002
rect 21728 -1011 21894 -1002
rect 21527 -1012 21894 -1011
rect 19083 -1014 21894 -1012
rect 18576 -1015 21894 -1014
rect 21946 -1011 22101 -1002
rect 22153 -1011 22306 -1002
rect 21946 -1012 22306 -1011
rect 22358 -1012 22653 -1002
rect 21946 -1015 22653 -1012
rect 18576 -1016 22653 -1015
rect 22705 -1012 24405 -1002
rect 24457 -1009 24596 -1002
rect 24648 -1007 24791 -1002
rect 24843 -1007 25238 -1002
rect 24648 -1009 25238 -1007
rect 24457 -1012 25238 -1009
rect 25290 -1012 25451 -960
rect 22705 -1016 25451 -1012
rect 18576 -1017 25451 -1016
rect 8449 -1023 25451 -1017
rect 8449 -1029 25436 -1023
rect 8449 -1033 25391 -1029
rect 10166 -1082 10232 -1078
rect 12558 -1082 12624 -1078
rect 14950 -1082 15016 -1078
rect 17342 -1082 17408 -1078
rect 19734 -1082 19800 -1078
rect 22126 -1082 22192 -1078
rect 24518 -1082 24584 -1080
rect 25391 -1082 25436 -1078
rect 8449 -1089 25436 -1082
rect 8431 -1101 25436 -1089
rect 8431 -1104 23597 -1101
rect 8431 -1106 12361 -1104
rect 8431 -1109 9070 -1106
rect 8431 -1113 8622 -1109
rect 8674 -1113 9070 -1109
rect 9122 -1108 12361 -1106
rect 9122 -1109 9504 -1108
rect 9122 -1113 9288 -1109
rect 8431 -1147 8604 -1113
rect 8674 -1147 8696 -1113
rect 8730 -1147 8788 -1113
rect 8822 -1147 8855 -1113
rect 8914 -1147 8972 -1113
rect 9006 -1147 9064 -1113
rect 9122 -1147 9156 -1113
rect 9190 -1147 9248 -1113
rect 9282 -1147 9288 -1113
rect 8431 -1161 8622 -1147
rect 8674 -1161 8855 -1147
rect 8431 -1165 8855 -1161
rect 8907 -1158 9070 -1147
rect 9122 -1158 9288 -1147
rect 8907 -1161 9288 -1158
rect 9340 -1113 9504 -1109
rect 9556 -1109 12361 -1108
rect 9556 -1112 11625 -1109
rect 9556 -1113 11225 -1112
rect 11277 -1113 11415 -1112
rect 11467 -1113 11625 -1112
rect 11677 -1112 12137 -1109
rect 11677 -1113 11842 -1112
rect 11894 -1113 12137 -1112
rect 9374 -1147 9432 -1113
rect 9466 -1147 9504 -1113
rect 9558 -1147 9616 -1113
rect 9650 -1147 9708 -1113
rect 9742 -1147 9800 -1113
rect 9834 -1147 9892 -1113
rect 9926 -1147 9984 -1113
rect 10018 -1147 10076 -1113
rect 10110 -1147 10168 -1113
rect 10202 -1147 10260 -1113
rect 10294 -1147 10352 -1113
rect 10386 -1147 10444 -1113
rect 10478 -1147 10536 -1113
rect 10570 -1147 10628 -1113
rect 10662 -1147 10720 -1113
rect 10754 -1147 10812 -1113
rect 10846 -1147 10904 -1113
rect 10938 -1147 10996 -1113
rect 11030 -1147 11088 -1113
rect 11122 -1147 11180 -1113
rect 11214 -1147 11225 -1113
rect 11306 -1147 11364 -1113
rect 11398 -1147 11415 -1113
rect 11490 -1147 11548 -1113
rect 11582 -1147 11625 -1113
rect 11677 -1147 11732 -1113
rect 11766 -1147 11824 -1113
rect 11894 -1147 11916 -1113
rect 11950 -1147 12008 -1113
rect 12042 -1147 12100 -1113
rect 12134 -1147 12137 -1113
rect 9340 -1160 9504 -1147
rect 9556 -1160 11225 -1147
rect 9340 -1161 11225 -1160
rect 8907 -1164 11225 -1161
rect 11277 -1164 11415 -1147
rect 11467 -1161 11625 -1147
rect 11677 -1161 11842 -1147
rect 11467 -1164 11842 -1161
rect 11894 -1161 12137 -1147
rect 12189 -1113 12361 -1109
rect 12413 -1109 15008 -1104
rect 12413 -1111 14791 -1109
rect 12413 -1113 14239 -1111
rect 14291 -1113 14791 -1111
rect 14843 -1113 15008 -1109
rect 15060 -1107 22965 -1104
rect 15060 -1113 15209 -1107
rect 15261 -1108 22965 -1107
rect 15261 -1113 18104 -1108
rect 18156 -1110 22965 -1108
rect 18156 -1112 20785 -1110
rect 18156 -1113 20005 -1112
rect 20057 -1113 20261 -1112
rect 20313 -1113 20496 -1112
rect 20548 -1113 20785 -1112
rect 12189 -1147 12192 -1113
rect 12226 -1147 12284 -1113
rect 12318 -1147 12361 -1113
rect 12413 -1147 12468 -1113
rect 12502 -1147 12560 -1113
rect 12594 -1147 12652 -1113
rect 12686 -1147 12744 -1113
rect 12778 -1147 12836 -1113
rect 12870 -1147 12928 -1113
rect 12962 -1147 13020 -1113
rect 13054 -1147 13112 -1113
rect 13146 -1147 13204 -1113
rect 13238 -1147 13296 -1113
rect 13330 -1147 13388 -1113
rect 13422 -1147 13480 -1113
rect 13514 -1147 13572 -1113
rect 13606 -1147 13664 -1113
rect 13698 -1147 13756 -1113
rect 13790 -1147 13848 -1113
rect 13882 -1147 13940 -1113
rect 13974 -1147 14032 -1113
rect 14066 -1147 14124 -1113
rect 14158 -1147 14216 -1113
rect 14291 -1147 14308 -1113
rect 14342 -1147 14400 -1113
rect 14434 -1147 14492 -1113
rect 14526 -1147 14539 -1113
rect 14618 -1147 14676 -1113
rect 14710 -1147 14768 -1113
rect 14843 -1147 14860 -1113
rect 14894 -1147 14952 -1113
rect 14986 -1147 15008 -1113
rect 15078 -1147 15136 -1113
rect 15170 -1147 15209 -1113
rect 15262 -1147 15320 -1113
rect 15354 -1147 15412 -1113
rect 15446 -1147 15504 -1113
rect 15538 -1147 15596 -1113
rect 15630 -1147 15688 -1113
rect 15722 -1147 15780 -1113
rect 15814 -1147 15872 -1113
rect 15906 -1147 15964 -1113
rect 15998 -1147 16056 -1113
rect 16090 -1147 16148 -1113
rect 16182 -1147 16240 -1113
rect 16274 -1147 16332 -1113
rect 16366 -1147 16424 -1113
rect 16458 -1147 16516 -1113
rect 16550 -1147 16608 -1113
rect 16642 -1147 16700 -1113
rect 16734 -1147 16792 -1113
rect 16826 -1147 16884 -1113
rect 16918 -1147 16976 -1113
rect 17010 -1147 17068 -1113
rect 17102 -1116 17160 -1113
rect 17146 -1147 17160 -1116
rect 17194 -1147 17252 -1113
rect 17286 -1116 17344 -1113
rect 12189 -1156 12361 -1147
rect 12413 -1156 14239 -1147
rect 12189 -1161 14239 -1156
rect 11894 -1163 14239 -1161
rect 14291 -1163 14539 -1147
rect 11894 -1164 14539 -1163
rect 8907 -1165 14539 -1164
rect 14591 -1161 14791 -1147
rect 14843 -1156 15008 -1147
rect 15060 -1156 15209 -1147
rect 14843 -1159 15209 -1156
rect 15261 -1159 17094 -1147
rect 14843 -1161 17094 -1159
rect 14591 -1165 17094 -1161
rect 8431 -1168 17094 -1165
rect 17146 -1168 17286 -1147
rect 17338 -1147 17344 -1116
rect 17378 -1147 17436 -1113
rect 17470 -1116 17528 -1113
rect 17470 -1147 17486 -1116
rect 17562 -1147 17620 -1113
rect 17654 -1147 17712 -1113
rect 17746 -1147 17804 -1113
rect 17838 -1147 17896 -1113
rect 17930 -1147 17988 -1113
rect 18022 -1147 18080 -1113
rect 18156 -1147 18172 -1113
rect 18206 -1147 18264 -1113
rect 18298 -1147 18356 -1113
rect 18390 -1147 18448 -1113
rect 18482 -1147 18540 -1113
rect 18574 -1147 18632 -1113
rect 18666 -1147 18724 -1113
rect 18758 -1147 18816 -1113
rect 18850 -1147 18908 -1113
rect 18942 -1147 19000 -1113
rect 19034 -1147 19092 -1113
rect 19126 -1147 19184 -1113
rect 19218 -1147 19276 -1113
rect 19310 -1147 19368 -1113
rect 19402 -1147 19460 -1113
rect 19494 -1147 19552 -1113
rect 19586 -1147 19644 -1113
rect 19678 -1147 19736 -1113
rect 19770 -1147 19828 -1113
rect 19862 -1147 19920 -1113
rect 19954 -1147 20005 -1113
rect 20057 -1147 20104 -1113
rect 20138 -1147 20196 -1113
rect 20230 -1147 20261 -1113
rect 20322 -1147 20380 -1113
rect 20414 -1147 20472 -1113
rect 20548 -1147 20564 -1113
rect 20598 -1147 20656 -1113
rect 20690 -1147 20748 -1113
rect 20782 -1147 20785 -1113
rect 17338 -1168 17486 -1147
rect 17538 -1160 18104 -1147
rect 18156 -1160 20005 -1147
rect 17538 -1164 20005 -1160
rect 20057 -1164 20261 -1147
rect 20313 -1164 20496 -1147
rect 20548 -1162 20785 -1147
rect 20837 -1112 21179 -1110
rect 20837 -1113 20975 -1112
rect 21027 -1113 21179 -1112
rect 21231 -1113 22965 -1110
rect 23017 -1108 23597 -1104
rect 23017 -1113 23207 -1108
rect 23259 -1109 23597 -1108
rect 23259 -1113 23407 -1109
rect 23459 -1113 23597 -1109
rect 23649 -1103 25436 -1101
rect 23649 -1113 23818 -1103
rect 20837 -1147 20840 -1113
rect 20874 -1147 20932 -1113
rect 20966 -1147 20975 -1113
rect 21058 -1147 21116 -1113
rect 21150 -1147 21179 -1113
rect 21242 -1147 21300 -1113
rect 21334 -1147 21392 -1113
rect 21426 -1147 21484 -1113
rect 21518 -1147 21576 -1113
rect 21610 -1147 21668 -1113
rect 21702 -1147 21760 -1113
rect 21794 -1147 21852 -1113
rect 21886 -1147 21944 -1113
rect 21978 -1147 22036 -1113
rect 22070 -1147 22128 -1113
rect 22162 -1147 22220 -1113
rect 22254 -1147 22312 -1113
rect 22346 -1147 22404 -1113
rect 22438 -1147 22496 -1113
rect 22530 -1147 22588 -1113
rect 22622 -1147 22680 -1113
rect 22714 -1147 22772 -1113
rect 22806 -1147 22864 -1113
rect 22898 -1147 22956 -1113
rect 23017 -1147 23048 -1113
rect 23082 -1147 23140 -1113
rect 23174 -1147 23207 -1113
rect 23266 -1147 23324 -1113
rect 23358 -1147 23407 -1113
rect 23459 -1147 23508 -1113
rect 23542 -1147 23597 -1113
rect 23649 -1147 23692 -1113
rect 23726 -1147 23784 -1113
rect 20837 -1162 20975 -1147
rect 20548 -1164 20975 -1162
rect 21027 -1162 21179 -1147
rect 21231 -1156 22965 -1147
rect 23017 -1156 23207 -1147
rect 21231 -1160 23207 -1156
rect 23259 -1160 23407 -1147
rect 21231 -1161 23407 -1160
rect 23459 -1153 23597 -1147
rect 23649 -1153 23818 -1147
rect 23459 -1155 23818 -1153
rect 23870 -1108 25436 -1103
rect 23870 -1113 24114 -1108
rect 24166 -1113 25436 -1108
rect 23870 -1147 23876 -1113
rect 23910 -1147 23968 -1113
rect 24002 -1147 24060 -1113
rect 24094 -1147 24114 -1113
rect 24186 -1147 24244 -1113
rect 24278 -1147 24336 -1113
rect 24370 -1147 24428 -1113
rect 24462 -1147 24520 -1113
rect 24554 -1147 24612 -1113
rect 24646 -1147 24704 -1113
rect 24738 -1147 24796 -1113
rect 24830 -1147 24888 -1113
rect 24922 -1147 24980 -1113
rect 25014 -1147 25072 -1113
rect 25106 -1147 25164 -1113
rect 25198 -1147 25256 -1113
rect 25290 -1147 25436 -1113
rect 23870 -1155 24114 -1147
rect 23459 -1160 24114 -1155
rect 24166 -1160 25436 -1147
rect 23459 -1161 25436 -1160
rect 21231 -1162 25436 -1161
rect 21027 -1164 25436 -1162
rect 17538 -1168 25436 -1164
rect 8431 -1174 25436 -1168
rect 8431 -1175 25391 -1174
rect 8449 -1178 25391 -1175
rect 20959 -1179 21056 -1178
rect 8592 -1215 8644 -1209
rect 10984 -1215 11036 -1209
rect 9594 -1263 9600 -1251
rect 8592 -1273 8644 -1267
rect 8872 -1279 8924 -1273
rect 8872 -1337 8924 -1331
rect 9083 -1294 9600 -1263
rect 9083 -1411 9112 -1294
rect 9594 -1303 9600 -1294
rect 9652 -1303 9658 -1251
rect 13377 -1215 13429 -1209
rect 11986 -1262 11992 -1250
rect 10984 -1273 11036 -1267
rect 9696 -1283 9754 -1277
rect 9696 -1317 9708 -1283
rect 9742 -1286 9754 -1283
rect 10432 -1283 10490 -1277
rect 10432 -1286 10444 -1283
rect 9742 -1314 10444 -1286
rect 9742 -1317 9754 -1314
rect 9696 -1323 9754 -1317
rect 10432 -1317 10444 -1314
rect 10478 -1286 10490 -1283
rect 10708 -1283 10766 -1277
rect 10708 -1286 10720 -1283
rect 10478 -1314 10720 -1286
rect 10478 -1317 10490 -1314
rect 10432 -1323 10490 -1317
rect 10708 -1317 10720 -1314
rect 10754 -1317 10766 -1283
rect 10708 -1323 10766 -1317
rect 11264 -1279 11316 -1273
rect 11264 -1337 11316 -1331
rect 11475 -1293 11992 -1262
rect 9150 -1351 9208 -1345
rect 9150 -1385 9162 -1351
rect 9196 -1354 9208 -1351
rect 9788 -1351 9846 -1345
rect 9788 -1354 9800 -1351
rect 9196 -1382 9800 -1354
rect 9196 -1385 9208 -1382
rect 9150 -1391 9208 -1385
rect 9788 -1385 9800 -1382
rect 9834 -1385 9846 -1351
rect 9788 -1391 9846 -1385
rect 10873 -1402 10879 -1350
rect 10933 -1402 10939 -1350
rect 9065 -1417 9123 -1411
rect 9065 -1451 9077 -1417
rect 9111 -1451 9123 -1417
rect 9065 -1457 9123 -1451
rect 9696 -1419 9754 -1413
rect 9696 -1453 9708 -1419
rect 9742 -1422 9754 -1419
rect 9742 -1450 10383 -1422
rect 9742 -1453 9754 -1450
rect 9083 -1458 9112 -1457
rect 9696 -1459 9754 -1453
rect 10340 -1481 10383 -1450
rect 10528 -1458 10534 -1405
rect 10586 -1458 10593 -1405
rect 11475 -1409 11504 -1293
rect 11986 -1302 11992 -1293
rect 12044 -1302 12050 -1250
rect 15768 -1215 15820 -1209
rect 14378 -1263 14384 -1251
rect 13377 -1273 13429 -1267
rect 12088 -1283 12146 -1277
rect 12088 -1317 12100 -1283
rect 12134 -1286 12146 -1283
rect 12824 -1283 12882 -1277
rect 12824 -1286 12836 -1283
rect 12134 -1314 12836 -1286
rect 12134 -1317 12146 -1314
rect 12088 -1323 12146 -1317
rect 12824 -1317 12836 -1314
rect 12870 -1286 12882 -1283
rect 13100 -1283 13158 -1277
rect 13100 -1286 13112 -1283
rect 12870 -1314 13112 -1286
rect 12870 -1317 12882 -1314
rect 12824 -1323 12882 -1317
rect 13100 -1317 13112 -1314
rect 13146 -1317 13158 -1283
rect 13100 -1323 13158 -1317
rect 13655 -1279 13707 -1273
rect 13655 -1337 13707 -1331
rect 13867 -1294 14384 -1263
rect 11542 -1351 11600 -1345
rect 11542 -1385 11554 -1351
rect 11588 -1354 11600 -1351
rect 12180 -1351 12238 -1345
rect 12180 -1354 12192 -1351
rect 11588 -1382 12192 -1354
rect 11588 -1385 11600 -1382
rect 11542 -1391 11600 -1385
rect 12180 -1385 12192 -1382
rect 12226 -1385 12238 -1351
rect 12180 -1391 12238 -1385
rect 13267 -1402 13273 -1350
rect 13327 -1402 13333 -1350
rect 11454 -1415 11512 -1409
rect 11454 -1449 11466 -1415
rect 11500 -1449 11512 -1415
rect 11454 -1455 11512 -1449
rect 12088 -1419 12146 -1413
rect 12088 -1453 12100 -1419
rect 12134 -1422 12146 -1419
rect 12134 -1450 12775 -1422
rect 12134 -1453 12146 -1450
rect 11475 -1457 11504 -1455
rect 10528 -1459 10593 -1458
rect 12088 -1459 12146 -1453
rect 12732 -1481 12775 -1450
rect 12920 -1458 12926 -1405
rect 12978 -1458 12985 -1405
rect 13867 -1409 13896 -1294
rect 14378 -1303 14384 -1294
rect 14436 -1303 14442 -1251
rect 18160 -1216 18212 -1210
rect 16770 -1263 16776 -1251
rect 15768 -1273 15820 -1267
rect 14480 -1283 14538 -1277
rect 14480 -1317 14492 -1283
rect 14526 -1286 14538 -1283
rect 15216 -1283 15274 -1277
rect 15216 -1286 15228 -1283
rect 14526 -1314 15228 -1286
rect 14526 -1317 14538 -1314
rect 14480 -1323 14538 -1317
rect 15216 -1317 15228 -1314
rect 15262 -1286 15274 -1283
rect 15492 -1283 15550 -1277
rect 15492 -1286 15504 -1283
rect 15262 -1314 15504 -1286
rect 15262 -1317 15274 -1314
rect 15216 -1323 15274 -1317
rect 15492 -1317 15504 -1314
rect 15538 -1317 15550 -1283
rect 15492 -1323 15550 -1317
rect 16048 -1279 16100 -1273
rect 16048 -1337 16100 -1331
rect 16259 -1294 16776 -1263
rect 13934 -1351 13992 -1345
rect 13934 -1385 13946 -1351
rect 13980 -1354 13992 -1351
rect 14572 -1351 14630 -1345
rect 14572 -1354 14584 -1351
rect 13980 -1382 14584 -1354
rect 13980 -1385 13992 -1382
rect 13934 -1391 13992 -1385
rect 14572 -1385 14584 -1382
rect 14618 -1385 14630 -1351
rect 14572 -1391 14630 -1385
rect 15657 -1400 15663 -1348
rect 15717 -1400 15723 -1348
rect 15311 -1405 15376 -1404
rect 13847 -1415 13905 -1409
rect 13847 -1449 13859 -1415
rect 13893 -1449 13905 -1415
rect 13847 -1455 13905 -1449
rect 14480 -1419 14538 -1413
rect 14480 -1453 14492 -1419
rect 14526 -1422 14538 -1419
rect 14526 -1450 15167 -1422
rect 14526 -1453 14538 -1450
rect 13867 -1458 13896 -1455
rect 12920 -1459 12985 -1458
rect 14480 -1459 14538 -1453
rect 15124 -1481 15167 -1450
rect 15311 -1457 15317 -1405
rect 15369 -1457 15376 -1405
rect 16259 -1409 16288 -1294
rect 16770 -1303 16776 -1294
rect 16828 -1303 16834 -1251
rect 20553 -1214 20605 -1208
rect 19162 -1263 19168 -1251
rect 18160 -1274 18212 -1268
rect 16872 -1283 16930 -1277
rect 16872 -1317 16884 -1283
rect 16918 -1286 16930 -1283
rect 17608 -1283 17666 -1277
rect 17608 -1286 17620 -1283
rect 16918 -1314 17620 -1286
rect 16918 -1317 16930 -1314
rect 16872 -1323 16930 -1317
rect 17608 -1317 17620 -1314
rect 17654 -1286 17666 -1283
rect 17884 -1283 17942 -1277
rect 17884 -1286 17896 -1283
rect 17654 -1314 17896 -1286
rect 17654 -1317 17666 -1314
rect 17608 -1323 17666 -1317
rect 17884 -1317 17896 -1314
rect 17930 -1317 17942 -1283
rect 17884 -1323 17942 -1317
rect 18440 -1279 18492 -1273
rect 18440 -1337 18492 -1331
rect 18651 -1294 19168 -1263
rect 16326 -1351 16384 -1345
rect 16326 -1385 16338 -1351
rect 16372 -1354 16384 -1351
rect 16964 -1351 17022 -1345
rect 16964 -1354 16976 -1351
rect 16372 -1382 16976 -1354
rect 16372 -1385 16384 -1382
rect 16326 -1391 16384 -1385
rect 16964 -1385 16976 -1382
rect 17010 -1385 17022 -1351
rect 16964 -1391 17022 -1385
rect 18049 -1402 18055 -1350
rect 18109 -1402 18115 -1350
rect 16240 -1415 16298 -1409
rect 16240 -1449 16252 -1415
rect 16286 -1449 16298 -1415
rect 16240 -1455 16298 -1449
rect 16872 -1419 16930 -1413
rect 16872 -1453 16884 -1419
rect 16918 -1422 16930 -1419
rect 16918 -1450 17559 -1422
rect 16918 -1453 16930 -1450
rect 15311 -1458 15376 -1457
rect 16259 -1458 16288 -1455
rect 16872 -1459 16930 -1453
rect 17516 -1481 17559 -1450
rect 17704 -1458 17710 -1405
rect 17762 -1458 17769 -1405
rect 18651 -1409 18680 -1294
rect 19162 -1303 19168 -1294
rect 19220 -1303 19226 -1251
rect 22944 -1214 22996 -1208
rect 21554 -1262 21560 -1250
rect 20553 -1272 20605 -1266
rect 19264 -1283 19322 -1277
rect 19264 -1317 19276 -1283
rect 19310 -1286 19322 -1283
rect 20000 -1283 20058 -1277
rect 20000 -1286 20012 -1283
rect 19310 -1314 20012 -1286
rect 19310 -1317 19322 -1314
rect 19264 -1323 19322 -1317
rect 20000 -1317 20012 -1314
rect 20046 -1286 20058 -1283
rect 20276 -1283 20334 -1277
rect 20276 -1286 20288 -1283
rect 20046 -1314 20288 -1286
rect 20046 -1317 20058 -1314
rect 20000 -1323 20058 -1317
rect 20276 -1317 20288 -1314
rect 20322 -1317 20334 -1283
rect 20276 -1323 20334 -1317
rect 20831 -1278 20883 -1272
rect 20831 -1336 20883 -1330
rect 21043 -1293 21560 -1262
rect 18718 -1351 18776 -1345
rect 18718 -1385 18730 -1351
rect 18764 -1354 18776 -1351
rect 19356 -1351 19414 -1345
rect 19356 -1354 19368 -1351
rect 18764 -1382 19368 -1354
rect 18764 -1385 18776 -1382
rect 18718 -1391 18776 -1385
rect 19356 -1385 19368 -1382
rect 19402 -1385 19414 -1351
rect 19356 -1391 19414 -1385
rect 20441 -1400 20447 -1348
rect 20501 -1400 20507 -1348
rect 18631 -1415 18689 -1409
rect 18631 -1449 18643 -1415
rect 18677 -1449 18689 -1415
rect 18631 -1455 18689 -1449
rect 19264 -1419 19322 -1413
rect 19264 -1453 19276 -1419
rect 19310 -1422 19322 -1419
rect 19310 -1450 19951 -1422
rect 19310 -1453 19322 -1450
rect 18651 -1458 18680 -1455
rect 17704 -1459 17769 -1458
rect 19264 -1459 19322 -1453
rect 19908 -1481 19951 -1450
rect 20095 -1458 20101 -1405
rect 20153 -1458 20160 -1405
rect 21043 -1409 21072 -1293
rect 21554 -1302 21560 -1293
rect 21612 -1302 21618 -1250
rect 23946 -1262 23952 -1250
rect 22944 -1272 22996 -1266
rect 21656 -1283 21714 -1277
rect 21656 -1317 21668 -1283
rect 21702 -1286 21714 -1283
rect 22392 -1283 22450 -1277
rect 22392 -1286 22404 -1283
rect 21702 -1314 22404 -1286
rect 21702 -1317 21714 -1314
rect 21656 -1323 21714 -1317
rect 22392 -1317 22404 -1314
rect 22438 -1286 22450 -1283
rect 22668 -1283 22726 -1277
rect 22668 -1286 22680 -1283
rect 22438 -1314 22680 -1286
rect 22438 -1317 22450 -1314
rect 22392 -1323 22450 -1317
rect 22668 -1317 22680 -1314
rect 22714 -1317 22726 -1283
rect 22668 -1323 22726 -1317
rect 23224 -1279 23276 -1273
rect 23224 -1337 23276 -1331
rect 23435 -1293 23952 -1262
rect 21110 -1351 21168 -1345
rect 21110 -1385 21122 -1351
rect 21156 -1354 21168 -1351
rect 21748 -1351 21806 -1345
rect 21748 -1354 21760 -1351
rect 21156 -1382 21760 -1354
rect 21156 -1385 21168 -1382
rect 21110 -1391 21168 -1385
rect 21748 -1385 21760 -1382
rect 21794 -1385 21806 -1351
rect 21748 -1391 21806 -1385
rect 22833 -1402 22839 -1350
rect 22893 -1402 22899 -1350
rect 21024 -1415 21082 -1409
rect 21024 -1449 21036 -1415
rect 21070 -1449 21082 -1415
rect 21024 -1455 21082 -1449
rect 21656 -1419 21714 -1413
rect 21656 -1453 21668 -1419
rect 21702 -1422 21714 -1419
rect 21702 -1450 22343 -1422
rect 21702 -1453 21714 -1450
rect 21043 -1457 21072 -1455
rect 20095 -1459 20160 -1458
rect 21656 -1459 21714 -1453
rect 22300 -1481 22343 -1450
rect 22488 -1458 22494 -1405
rect 22546 -1458 22553 -1405
rect 23435 -1409 23464 -1293
rect 23946 -1302 23952 -1293
rect 24004 -1302 24010 -1250
rect 24048 -1283 24106 -1277
rect 24048 -1317 24060 -1283
rect 24094 -1286 24106 -1283
rect 24784 -1283 24842 -1277
rect 24784 -1286 24796 -1283
rect 24094 -1314 24796 -1286
rect 24094 -1317 24106 -1314
rect 24048 -1323 24106 -1317
rect 24784 -1317 24796 -1314
rect 24830 -1286 24842 -1283
rect 25060 -1283 25118 -1277
rect 25060 -1286 25072 -1283
rect 24830 -1314 25072 -1286
rect 24830 -1317 24842 -1314
rect 24784 -1323 24842 -1317
rect 25060 -1317 25072 -1314
rect 25106 -1317 25118 -1283
rect 25060 -1323 25118 -1317
rect 23502 -1351 23560 -1345
rect 23502 -1385 23514 -1351
rect 23548 -1354 23560 -1351
rect 24140 -1351 24198 -1345
rect 24140 -1354 24152 -1351
rect 23548 -1382 24152 -1354
rect 23548 -1385 23560 -1382
rect 23502 -1391 23560 -1385
rect 24140 -1385 24152 -1382
rect 24186 -1385 24198 -1351
rect 24140 -1391 24198 -1385
rect 25225 -1400 25231 -1348
rect 25285 -1400 25291 -1348
rect 23415 -1415 23473 -1409
rect 23415 -1449 23427 -1415
rect 23461 -1449 23473 -1415
rect 23415 -1455 23473 -1449
rect 24048 -1419 24106 -1413
rect 24048 -1453 24060 -1419
rect 24094 -1422 24106 -1419
rect 24094 -1450 24735 -1422
rect 24094 -1453 24106 -1450
rect 23435 -1457 23464 -1455
rect 22488 -1459 22553 -1458
rect 24048 -1459 24106 -1453
rect 24692 -1481 24735 -1450
rect 24881 -1458 24887 -1405
rect 24939 -1458 24946 -1405
rect 24881 -1459 24946 -1458
rect 9406 -1487 9464 -1481
rect 9406 -1521 9418 -1487
rect 9452 -1490 9464 -1487
rect 10156 -1487 10214 -1481
rect 10156 -1490 10168 -1487
rect 9452 -1518 10168 -1490
rect 9452 -1521 9464 -1518
rect 9406 -1527 9464 -1521
rect 10156 -1521 10168 -1518
rect 10202 -1521 10214 -1487
rect 10156 -1527 10214 -1521
rect 10340 -1487 10398 -1481
rect 10340 -1521 10352 -1487
rect 10386 -1490 10398 -1487
rect 10799 -1487 10857 -1481
rect 10799 -1490 10811 -1487
rect 10386 -1518 10811 -1490
rect 10386 -1521 10398 -1518
rect 10340 -1527 10398 -1521
rect 10799 -1521 10811 -1518
rect 10845 -1521 10857 -1487
rect 10799 -1527 10857 -1521
rect 11798 -1487 11856 -1481
rect 11798 -1521 11810 -1487
rect 11844 -1490 11856 -1487
rect 12548 -1487 12606 -1481
rect 12548 -1490 12560 -1487
rect 11844 -1518 12560 -1490
rect 11844 -1521 11856 -1518
rect 11798 -1527 11856 -1521
rect 12548 -1521 12560 -1518
rect 12594 -1521 12606 -1487
rect 12548 -1527 12606 -1521
rect 12732 -1487 12790 -1481
rect 12732 -1521 12744 -1487
rect 12778 -1490 12790 -1487
rect 13191 -1487 13249 -1481
rect 13191 -1490 13203 -1487
rect 12778 -1518 13203 -1490
rect 12778 -1521 12790 -1518
rect 12732 -1527 12790 -1521
rect 13191 -1521 13203 -1518
rect 13237 -1521 13249 -1487
rect 13191 -1527 13249 -1521
rect 14190 -1487 14248 -1481
rect 14190 -1521 14202 -1487
rect 14236 -1490 14248 -1487
rect 14940 -1487 14998 -1481
rect 14940 -1490 14952 -1487
rect 14236 -1518 14952 -1490
rect 14236 -1521 14248 -1518
rect 14190 -1527 14248 -1521
rect 14940 -1521 14952 -1518
rect 14986 -1521 14998 -1487
rect 14940 -1527 14998 -1521
rect 15124 -1487 15182 -1481
rect 15124 -1521 15136 -1487
rect 15170 -1490 15182 -1487
rect 15583 -1487 15641 -1481
rect 15583 -1490 15595 -1487
rect 15170 -1518 15595 -1490
rect 15170 -1521 15182 -1518
rect 15124 -1527 15182 -1521
rect 15583 -1521 15595 -1518
rect 15629 -1521 15641 -1487
rect 15583 -1527 15641 -1521
rect 16582 -1487 16640 -1481
rect 16582 -1521 16594 -1487
rect 16628 -1490 16640 -1487
rect 17332 -1487 17390 -1481
rect 17332 -1490 17344 -1487
rect 16628 -1518 17344 -1490
rect 16628 -1521 16640 -1518
rect 16582 -1527 16640 -1521
rect 17332 -1521 17344 -1518
rect 17378 -1521 17390 -1487
rect 17332 -1527 17390 -1521
rect 17516 -1487 17574 -1481
rect 17516 -1521 17528 -1487
rect 17562 -1490 17574 -1487
rect 17975 -1487 18033 -1481
rect 17975 -1490 17987 -1487
rect 17562 -1518 17987 -1490
rect 17562 -1521 17574 -1518
rect 17516 -1527 17574 -1521
rect 17975 -1521 17987 -1518
rect 18021 -1521 18033 -1487
rect 17975 -1527 18033 -1521
rect 18974 -1487 19032 -1481
rect 18974 -1521 18986 -1487
rect 19020 -1490 19032 -1487
rect 19724 -1487 19782 -1481
rect 19724 -1490 19736 -1487
rect 19020 -1518 19736 -1490
rect 19020 -1521 19032 -1518
rect 18974 -1527 19032 -1521
rect 19724 -1521 19736 -1518
rect 19770 -1521 19782 -1487
rect 19724 -1527 19782 -1521
rect 19908 -1487 19966 -1481
rect 19908 -1521 19920 -1487
rect 19954 -1490 19966 -1487
rect 20367 -1487 20425 -1481
rect 20367 -1490 20379 -1487
rect 19954 -1518 20379 -1490
rect 19954 -1521 19966 -1518
rect 19908 -1527 19966 -1521
rect 20367 -1521 20379 -1518
rect 20413 -1521 20425 -1487
rect 20367 -1527 20425 -1521
rect 21366 -1487 21424 -1481
rect 21366 -1521 21378 -1487
rect 21412 -1490 21424 -1487
rect 22116 -1487 22174 -1481
rect 22116 -1490 22128 -1487
rect 21412 -1518 22128 -1490
rect 21412 -1521 21424 -1518
rect 21366 -1527 21424 -1521
rect 22116 -1521 22128 -1518
rect 22162 -1521 22174 -1487
rect 22116 -1527 22174 -1521
rect 22300 -1487 22358 -1481
rect 22300 -1521 22312 -1487
rect 22346 -1490 22358 -1487
rect 22759 -1487 22817 -1481
rect 22759 -1490 22771 -1487
rect 22346 -1518 22771 -1490
rect 22346 -1521 22358 -1518
rect 22300 -1527 22358 -1521
rect 22759 -1521 22771 -1518
rect 22805 -1521 22817 -1487
rect 22759 -1527 22817 -1521
rect 23758 -1487 23816 -1481
rect 23758 -1521 23770 -1487
rect 23804 -1490 23816 -1487
rect 24508 -1487 24566 -1481
rect 24508 -1490 24520 -1487
rect 23804 -1518 24520 -1490
rect 23804 -1521 23816 -1518
rect 23758 -1527 23816 -1521
rect 24508 -1521 24520 -1518
rect 24554 -1521 24566 -1487
rect 24508 -1527 24566 -1521
rect 24692 -1487 24750 -1481
rect 24692 -1521 24704 -1487
rect 24738 -1490 24750 -1487
rect 25151 -1487 25209 -1481
rect 25151 -1490 25163 -1487
rect 24738 -1518 25163 -1490
rect 24738 -1521 24750 -1518
rect 24692 -1527 24750 -1521
rect 25151 -1521 25163 -1518
rect 25197 -1521 25209 -1487
rect 25151 -1527 25209 -1521
rect 25391 -1626 25436 -1622
rect 8449 -1629 25436 -1626
rect 8449 -1639 25451 -1629
rect 8449 -1641 10738 -1639
rect 8449 -1657 8996 -1641
rect 9048 -1644 10738 -1641
rect 9048 -1657 9195 -1644
rect 8449 -1691 8604 -1657
rect 8638 -1691 8696 -1657
rect 8730 -1691 8788 -1657
rect 8822 -1691 8880 -1657
rect 8914 -1691 8972 -1657
rect 9048 -1691 9064 -1657
rect 9098 -1691 9156 -1657
rect 9190 -1691 9195 -1657
rect 8449 -1693 8996 -1691
rect 9048 -1693 9195 -1691
rect 8449 -1696 9195 -1693
rect 9247 -1657 9406 -1644
rect 9458 -1657 9612 -1644
rect 9664 -1646 10314 -1644
rect 9664 -1657 9840 -1646
rect 9247 -1691 9248 -1657
rect 9282 -1691 9340 -1657
rect 9374 -1691 9406 -1657
rect 9466 -1691 9524 -1657
rect 9558 -1691 9612 -1657
rect 9664 -1691 9708 -1657
rect 9742 -1691 9800 -1657
rect 9834 -1691 9840 -1657
rect 9247 -1696 9406 -1691
rect 9458 -1696 9612 -1691
rect 9664 -1696 9840 -1691
rect 8449 -1698 9840 -1696
rect 9892 -1657 10084 -1646
rect 10136 -1657 10314 -1646
rect 10366 -1657 10520 -1644
rect 10572 -1657 10738 -1644
rect 10790 -1642 25451 -1639
rect 10790 -1645 11149 -1642
rect 10790 -1657 10941 -1645
rect 9926 -1691 9984 -1657
rect 10018 -1691 10076 -1657
rect 10136 -1691 10168 -1657
rect 10202 -1691 10260 -1657
rect 10294 -1691 10314 -1657
rect 10386 -1691 10444 -1657
rect 10478 -1691 10520 -1657
rect 10572 -1691 10628 -1657
rect 10662 -1691 10720 -1657
rect 10790 -1691 10812 -1657
rect 10846 -1691 10904 -1657
rect 10938 -1691 10941 -1657
rect 9892 -1698 10084 -1691
rect 10136 -1696 10314 -1691
rect 10366 -1696 10520 -1691
rect 10572 -1696 10941 -1691
rect 10136 -1697 10941 -1696
rect 10993 -1657 11149 -1645
rect 11201 -1645 12030 -1642
rect 11201 -1646 11620 -1645
rect 11201 -1657 11412 -1646
rect 11464 -1657 11620 -1646
rect 11672 -1648 12030 -1645
rect 11672 -1657 11830 -1648
rect 11882 -1657 12030 -1648
rect 12082 -1643 15910 -1642
rect 12082 -1644 12860 -1643
rect 12082 -1645 12644 -1644
rect 12082 -1657 12233 -1645
rect 12285 -1657 12443 -1645
rect 12495 -1657 12644 -1645
rect 12696 -1657 12860 -1644
rect 12912 -1645 13787 -1643
rect 12912 -1657 13141 -1645
rect 13193 -1649 13787 -1645
rect 13193 -1650 13566 -1649
rect 13193 -1657 13361 -1650
rect 13413 -1657 13566 -1650
rect 13618 -1657 13787 -1649
rect 13839 -1644 15910 -1643
rect 13839 -1649 14632 -1644
rect 13839 -1650 14201 -1649
rect 13839 -1657 13992 -1650
rect 14044 -1657 14201 -1650
rect 14253 -1657 14418 -1649
rect 14470 -1657 14632 -1649
rect 14684 -1645 15707 -1644
rect 14684 -1646 15508 -1645
rect 14684 -1657 14827 -1646
rect 14879 -1649 15224 -1646
rect 14879 -1657 15022 -1649
rect 15074 -1657 15224 -1649
rect 15276 -1657 15508 -1646
rect 15560 -1657 15707 -1645
rect 15759 -1657 15910 -1644
rect 10993 -1691 10996 -1657
rect 11030 -1691 11088 -1657
rect 11122 -1691 11149 -1657
rect 11214 -1691 11272 -1657
rect 11306 -1691 11364 -1657
rect 11398 -1691 11412 -1657
rect 11490 -1691 11548 -1657
rect 11582 -1691 11620 -1657
rect 11674 -1691 11732 -1657
rect 11766 -1691 11824 -1657
rect 11882 -1691 11916 -1657
rect 11950 -1691 12008 -1657
rect 12082 -1691 12100 -1657
rect 12134 -1691 12192 -1657
rect 12226 -1691 12233 -1657
rect 12318 -1691 12376 -1657
rect 12410 -1691 12443 -1657
rect 12502 -1691 12560 -1657
rect 12594 -1691 12644 -1657
rect 12696 -1691 12744 -1657
rect 12778 -1691 12836 -1657
rect 12912 -1691 12928 -1657
rect 12962 -1691 13020 -1657
rect 13054 -1691 13112 -1657
rect 13193 -1691 13204 -1657
rect 13238 -1691 13296 -1657
rect 13330 -1691 13361 -1657
rect 13422 -1691 13480 -1657
rect 13514 -1691 13566 -1657
rect 13618 -1691 13664 -1657
rect 13698 -1691 13756 -1657
rect 13839 -1691 13848 -1657
rect 13882 -1691 13940 -1657
rect 13974 -1691 13992 -1657
rect 14066 -1691 14124 -1657
rect 14158 -1691 14201 -1657
rect 14253 -1691 14308 -1657
rect 14342 -1691 14400 -1657
rect 14470 -1691 14492 -1657
rect 14526 -1691 14584 -1657
rect 14618 -1691 14632 -1657
rect 14710 -1691 14768 -1657
rect 14802 -1691 14827 -1657
rect 14894 -1691 14952 -1657
rect 14986 -1691 15022 -1657
rect 15078 -1691 15136 -1657
rect 15170 -1691 15224 -1657
rect 15276 -1691 15320 -1657
rect 15354 -1691 15412 -1657
rect 15446 -1691 15504 -1657
rect 15560 -1691 15596 -1657
rect 15630 -1691 15688 -1657
rect 15759 -1691 15780 -1657
rect 15814 -1691 15872 -1657
rect 15906 -1691 15910 -1657
rect 10993 -1694 11149 -1691
rect 11201 -1694 11412 -1691
rect 10993 -1697 11412 -1694
rect 10136 -1698 11412 -1697
rect 11464 -1697 11620 -1691
rect 11672 -1697 11830 -1691
rect 11464 -1698 11830 -1697
rect 8449 -1700 11830 -1698
rect 11882 -1694 12030 -1691
rect 12082 -1694 12233 -1691
rect 11882 -1697 12233 -1694
rect 12285 -1697 12443 -1691
rect 12495 -1696 12644 -1691
rect 12696 -1695 12860 -1691
rect 12912 -1695 13141 -1691
rect 12696 -1696 13141 -1695
rect 12495 -1697 13141 -1696
rect 13193 -1697 13361 -1691
rect 11882 -1700 13361 -1697
rect 8449 -1702 13361 -1700
rect 13413 -1701 13566 -1691
rect 13618 -1695 13787 -1691
rect 13839 -1695 13992 -1691
rect 13618 -1701 13992 -1695
rect 13413 -1702 13992 -1701
rect 14044 -1701 14201 -1691
rect 14253 -1701 14418 -1691
rect 14470 -1696 14632 -1691
rect 14684 -1696 14827 -1691
rect 14470 -1698 14827 -1696
rect 14879 -1698 15022 -1691
rect 14470 -1701 15022 -1698
rect 15074 -1698 15224 -1691
rect 15276 -1697 15508 -1691
rect 15560 -1696 15707 -1691
rect 15759 -1694 15910 -1691
rect 15962 -1643 19392 -1642
rect 15962 -1644 17609 -1643
rect 15962 -1645 16562 -1644
rect 15962 -1657 16175 -1645
rect 16227 -1646 16562 -1645
rect 16227 -1657 16373 -1646
rect 16425 -1657 16562 -1646
rect 16614 -1657 16774 -1644
rect 16826 -1657 16991 -1644
rect 17043 -1648 17609 -1644
rect 17043 -1657 17196 -1648
rect 15962 -1691 15964 -1657
rect 15998 -1691 16056 -1657
rect 16090 -1691 16148 -1657
rect 16227 -1691 16240 -1657
rect 16274 -1691 16332 -1657
rect 16366 -1691 16373 -1657
rect 16458 -1691 16516 -1657
rect 16550 -1691 16562 -1657
rect 16642 -1691 16700 -1657
rect 16734 -1691 16774 -1657
rect 16826 -1691 16884 -1657
rect 16918 -1691 16976 -1657
rect 17043 -1691 17068 -1657
rect 17102 -1691 17160 -1657
rect 17194 -1691 17196 -1657
rect 15962 -1694 16175 -1691
rect 15759 -1696 16175 -1694
rect 15560 -1697 16175 -1696
rect 16227 -1697 16373 -1691
rect 15276 -1698 16373 -1697
rect 16425 -1696 16562 -1691
rect 16614 -1696 16774 -1691
rect 16826 -1696 16991 -1691
rect 17043 -1696 17196 -1691
rect 16425 -1698 17196 -1696
rect 15074 -1700 17196 -1698
rect 17248 -1657 17401 -1648
rect 17453 -1657 17609 -1648
rect 17661 -1644 19392 -1643
rect 17661 -1657 17892 -1644
rect 17944 -1646 18770 -1644
rect 17944 -1657 18085 -1646
rect 18137 -1648 18770 -1646
rect 18137 -1657 18311 -1648
rect 18363 -1657 18576 -1648
rect 17248 -1691 17252 -1657
rect 17286 -1691 17344 -1657
rect 17378 -1691 17401 -1657
rect 17470 -1691 17528 -1657
rect 17562 -1691 17609 -1657
rect 17661 -1691 17712 -1657
rect 17746 -1691 17804 -1657
rect 17838 -1691 17892 -1657
rect 17944 -1691 17988 -1657
rect 18022 -1691 18080 -1657
rect 18137 -1691 18172 -1657
rect 18206 -1691 18264 -1657
rect 18298 -1691 18311 -1657
rect 18390 -1691 18448 -1657
rect 18482 -1691 18540 -1657
rect 18574 -1691 18576 -1657
rect 17248 -1700 17401 -1691
rect 17453 -1695 17609 -1691
rect 17661 -1695 17892 -1691
rect 17453 -1696 17892 -1695
rect 17944 -1696 18085 -1691
rect 17453 -1698 18085 -1696
rect 18137 -1698 18311 -1691
rect 17453 -1700 18311 -1698
rect 18363 -1700 18576 -1691
rect 18628 -1657 18770 -1648
rect 18822 -1645 19392 -1644
rect 18822 -1653 19172 -1645
rect 18822 -1657 18968 -1653
rect 19020 -1657 19172 -1653
rect 19224 -1657 19392 -1645
rect 19444 -1643 25451 -1642
rect 19444 -1646 19835 -1643
rect 19444 -1657 19607 -1646
rect 19659 -1657 19835 -1646
rect 19887 -1644 20470 -1643
rect 19887 -1646 20277 -1644
rect 19887 -1657 20039 -1646
rect 20091 -1657 20277 -1646
rect 20329 -1657 20470 -1644
rect 20522 -1645 25451 -1643
rect 20522 -1648 20923 -1645
rect 20522 -1657 20667 -1648
rect 20719 -1657 20923 -1648
rect 20975 -1646 25451 -1645
rect 20975 -1648 22035 -1646
rect 20975 -1649 21616 -1648
rect 20975 -1657 21162 -1649
rect 21214 -1653 21616 -1649
rect 21214 -1657 21395 -1653
rect 21447 -1657 21616 -1653
rect 18628 -1691 18632 -1657
rect 18666 -1691 18724 -1657
rect 18758 -1691 18770 -1657
rect 18850 -1691 18908 -1657
rect 18942 -1691 18968 -1657
rect 19034 -1691 19092 -1657
rect 19126 -1691 19172 -1657
rect 19224 -1691 19276 -1657
rect 19310 -1691 19368 -1657
rect 19444 -1691 19460 -1657
rect 19494 -1691 19552 -1657
rect 19586 -1691 19607 -1657
rect 19678 -1691 19736 -1657
rect 19770 -1691 19828 -1657
rect 19887 -1691 19920 -1657
rect 19954 -1691 20012 -1657
rect 20091 -1691 20104 -1657
rect 20138 -1691 20196 -1657
rect 20230 -1691 20277 -1657
rect 20329 -1691 20380 -1657
rect 20414 -1691 20470 -1657
rect 20522 -1691 20564 -1657
rect 20598 -1691 20656 -1657
rect 20719 -1691 20748 -1657
rect 20782 -1691 20840 -1657
rect 20874 -1691 20923 -1657
rect 20975 -1691 21024 -1657
rect 21058 -1691 21116 -1657
rect 21150 -1691 21162 -1657
rect 21242 -1691 21300 -1657
rect 21334 -1691 21392 -1657
rect 21447 -1691 21484 -1657
rect 21518 -1691 21576 -1657
rect 21610 -1691 21616 -1657
rect 18628 -1696 18770 -1691
rect 18822 -1696 18968 -1691
rect 18628 -1700 18968 -1696
rect 15074 -1701 18968 -1700
rect 14044 -1702 18968 -1701
rect 8449 -1705 18968 -1702
rect 19020 -1697 19172 -1691
rect 19224 -1694 19392 -1691
rect 19444 -1694 19607 -1691
rect 19224 -1697 19607 -1694
rect 19020 -1698 19607 -1697
rect 19659 -1695 19835 -1691
rect 19887 -1695 20039 -1691
rect 19659 -1698 20039 -1695
rect 20091 -1696 20277 -1691
rect 20329 -1695 20470 -1691
rect 20522 -1695 20667 -1691
rect 20329 -1696 20667 -1695
rect 20091 -1698 20667 -1696
rect 19020 -1700 20667 -1698
rect 20719 -1697 20923 -1691
rect 20975 -1697 21162 -1691
rect 20719 -1700 21162 -1697
rect 19020 -1701 21162 -1700
rect 21214 -1701 21395 -1691
rect 19020 -1705 21395 -1701
rect 21447 -1700 21616 -1691
rect 21668 -1657 21807 -1648
rect 21859 -1657 22035 -1648
rect 22087 -1647 23086 -1646
rect 22087 -1648 22860 -1647
rect 22087 -1651 22671 -1648
rect 22087 -1657 22232 -1651
rect 22284 -1657 22444 -1651
rect 21702 -1691 21760 -1657
rect 21794 -1691 21807 -1657
rect 21886 -1691 21944 -1657
rect 21978 -1691 22035 -1657
rect 22087 -1691 22128 -1657
rect 22162 -1691 22220 -1657
rect 22284 -1691 22312 -1657
rect 22346 -1691 22404 -1657
rect 22438 -1691 22444 -1657
rect 21668 -1700 21807 -1691
rect 21859 -1698 22035 -1691
rect 22087 -1698 22232 -1691
rect 21859 -1700 22232 -1698
rect 21447 -1703 22232 -1700
rect 22284 -1703 22444 -1691
rect 22496 -1657 22671 -1651
rect 22723 -1657 22860 -1648
rect 22912 -1657 23086 -1647
rect 22530 -1691 22588 -1657
rect 22622 -1691 22671 -1657
rect 22723 -1691 22772 -1657
rect 22806 -1691 22860 -1657
rect 22912 -1691 22956 -1657
rect 22990 -1691 23048 -1657
rect 23082 -1691 23086 -1657
rect 22496 -1700 22671 -1691
rect 22723 -1699 22860 -1691
rect 22912 -1698 23086 -1691
rect 23138 -1657 23340 -1646
rect 23392 -1647 25072 -1646
rect 23392 -1649 24072 -1647
rect 23392 -1657 23584 -1649
rect 23636 -1650 24072 -1649
rect 23636 -1657 23814 -1650
rect 23866 -1657 24072 -1650
rect 24124 -1657 24282 -1647
rect 23138 -1691 23140 -1657
rect 23174 -1691 23232 -1657
rect 23266 -1691 23324 -1657
rect 23392 -1691 23416 -1657
rect 23450 -1691 23508 -1657
rect 23542 -1691 23584 -1657
rect 23636 -1691 23692 -1657
rect 23726 -1691 23784 -1657
rect 23866 -1691 23876 -1657
rect 23910 -1691 23968 -1657
rect 24002 -1691 24060 -1657
rect 24124 -1691 24152 -1657
rect 24186 -1691 24244 -1657
rect 24278 -1691 24282 -1657
rect 23138 -1698 23340 -1691
rect 23392 -1698 23584 -1691
rect 22912 -1699 23584 -1698
rect 22723 -1700 23584 -1699
rect 22496 -1701 23584 -1700
rect 23636 -1701 23814 -1691
rect 22496 -1702 23814 -1701
rect 23866 -1699 24072 -1691
rect 24124 -1699 24282 -1691
rect 24334 -1657 24507 -1647
rect 24559 -1650 25072 -1647
rect 24559 -1657 24726 -1650
rect 24778 -1657 25072 -1650
rect 25124 -1649 25451 -1646
rect 25124 -1657 25271 -1649
rect 24334 -1691 24336 -1657
rect 24370 -1691 24428 -1657
rect 24462 -1691 24507 -1657
rect 24559 -1691 24612 -1657
rect 24646 -1691 24704 -1657
rect 24778 -1691 24796 -1657
rect 24830 -1691 24888 -1657
rect 24922 -1691 24980 -1657
rect 25014 -1691 25072 -1657
rect 25124 -1691 25164 -1657
rect 25198 -1691 25256 -1657
rect 24334 -1699 24507 -1691
rect 24559 -1699 24726 -1691
rect 23866 -1702 24726 -1699
rect 24778 -1698 25072 -1691
rect 25124 -1698 25271 -1691
rect 24778 -1701 25271 -1698
rect 25323 -1701 25451 -1649
rect 24778 -1702 25451 -1701
rect 22496 -1703 25451 -1702
rect 21447 -1705 25451 -1703
rect 8449 -1715 25451 -1705
rect 8449 -1718 25436 -1715
rect 8449 -1722 25391 -1718
<< via1 >>
rect 13956 13574 14008 13626
rect 14054 13605 14106 13617
rect 14054 13571 14064 13605
rect 14064 13571 14098 13605
rect 14098 13571 14106 13605
rect 14054 13565 14106 13571
rect 14134 13605 14186 13617
rect 14134 13571 14144 13605
rect 14144 13571 14178 13605
rect 14178 13571 14186 13605
rect 14134 13565 14186 13571
rect 14214 13605 14266 13617
rect 14214 13571 14224 13605
rect 14224 13571 14258 13605
rect 14258 13571 14266 13605
rect 14214 13565 14266 13571
rect 14294 13605 14346 13617
rect 14294 13571 14304 13605
rect 14304 13571 14338 13605
rect 14338 13571 14346 13605
rect 14294 13565 14346 13571
rect 14374 13605 14426 13617
rect 14374 13571 14384 13605
rect 14384 13571 14418 13605
rect 14418 13571 14426 13605
rect 14374 13565 14426 13571
rect 14454 13605 14506 13617
rect 14454 13571 14464 13605
rect 14464 13571 14498 13605
rect 14498 13571 14506 13605
rect 14454 13565 14506 13571
rect 14786 13608 14838 13620
rect 14786 13574 14796 13608
rect 14796 13574 14830 13608
rect 14830 13574 14838 13608
rect 14786 13568 14838 13574
rect 14866 13608 14918 13620
rect 14866 13574 14876 13608
rect 14876 13574 14910 13608
rect 14910 13574 14918 13608
rect 14866 13568 14918 13574
rect 14946 13608 14998 13620
rect 14946 13574 14956 13608
rect 14956 13574 14990 13608
rect 14990 13574 14998 13608
rect 14946 13568 14998 13574
rect 15026 13608 15078 13620
rect 15026 13574 15036 13608
rect 15036 13574 15070 13608
rect 15070 13574 15078 13608
rect 15026 13568 15078 13574
rect 15106 13608 15158 13620
rect 15106 13574 15116 13608
rect 15116 13574 15150 13608
rect 15150 13574 15158 13608
rect 15106 13568 15158 13574
rect 15186 13608 15238 13620
rect 15186 13574 15196 13608
rect 15196 13574 15230 13608
rect 15230 13574 15238 13608
rect 15186 13568 15238 13574
rect 15390 13608 15442 13620
rect 15390 13574 15398 13608
rect 15398 13574 15432 13608
rect 15432 13574 15442 13608
rect 15390 13568 15442 13574
rect 15470 13608 15522 13620
rect 15470 13574 15478 13608
rect 15478 13574 15512 13608
rect 15512 13574 15522 13608
rect 15470 13568 15522 13574
rect 15550 13608 15602 13620
rect 15550 13574 15558 13608
rect 15558 13574 15592 13608
rect 15592 13574 15602 13608
rect 15550 13568 15602 13574
rect 15630 13608 15682 13620
rect 15630 13574 15638 13608
rect 15638 13574 15672 13608
rect 15672 13574 15682 13608
rect 15630 13568 15682 13574
rect 15710 13608 15762 13620
rect 15710 13574 15718 13608
rect 15718 13574 15752 13608
rect 15752 13574 15762 13608
rect 15710 13568 15762 13574
rect 15790 13608 15842 13620
rect 15790 13574 15798 13608
rect 15798 13574 15832 13608
rect 15832 13574 15842 13608
rect 15790 13568 15842 13574
rect 15998 13608 16050 13620
rect 15998 13574 16008 13608
rect 16008 13574 16042 13608
rect 16042 13574 16050 13608
rect 15998 13568 16050 13574
rect 16078 13608 16130 13620
rect 16078 13574 16088 13608
rect 16088 13574 16122 13608
rect 16122 13574 16130 13608
rect 16078 13568 16130 13574
rect 16158 13608 16210 13620
rect 16158 13574 16168 13608
rect 16168 13574 16202 13608
rect 16202 13574 16210 13608
rect 16158 13568 16210 13574
rect 16238 13608 16290 13620
rect 16238 13574 16248 13608
rect 16248 13574 16282 13608
rect 16282 13574 16290 13608
rect 16238 13568 16290 13574
rect 16318 13608 16370 13620
rect 16318 13574 16328 13608
rect 16328 13574 16362 13608
rect 16362 13574 16370 13608
rect 16318 13568 16370 13574
rect 16398 13608 16450 13620
rect 16398 13574 16408 13608
rect 16408 13574 16442 13608
rect 16442 13574 16450 13608
rect 16398 13568 16450 13574
rect 16602 13608 16654 13620
rect 16602 13574 16610 13608
rect 16610 13574 16644 13608
rect 16644 13574 16654 13608
rect 16602 13568 16654 13574
rect 16682 13608 16734 13620
rect 16682 13574 16690 13608
rect 16690 13574 16724 13608
rect 16724 13574 16734 13608
rect 16682 13568 16734 13574
rect 16762 13608 16814 13620
rect 16762 13574 16770 13608
rect 16770 13574 16804 13608
rect 16804 13574 16814 13608
rect 16762 13568 16814 13574
rect 16842 13608 16894 13620
rect 16842 13574 16850 13608
rect 16850 13574 16884 13608
rect 16884 13574 16894 13608
rect 16842 13568 16894 13574
rect 16922 13608 16974 13620
rect 16922 13574 16930 13608
rect 16930 13574 16964 13608
rect 16964 13574 16974 13608
rect 16922 13568 16974 13574
rect 17002 13608 17054 13620
rect 17002 13574 17010 13608
rect 17010 13574 17044 13608
rect 17044 13574 17054 13608
rect 17002 13568 17054 13574
rect 17210 13608 17262 13620
rect 17210 13574 17220 13608
rect 17220 13574 17254 13608
rect 17254 13574 17262 13608
rect 17210 13568 17262 13574
rect 17290 13608 17342 13620
rect 17290 13574 17300 13608
rect 17300 13574 17334 13608
rect 17334 13574 17342 13608
rect 17290 13568 17342 13574
rect 17370 13608 17422 13620
rect 17370 13574 17380 13608
rect 17380 13574 17414 13608
rect 17414 13574 17422 13608
rect 17370 13568 17422 13574
rect 17450 13608 17502 13620
rect 17450 13574 17460 13608
rect 17460 13574 17494 13608
rect 17494 13574 17502 13608
rect 17450 13568 17502 13574
rect 17530 13608 17582 13620
rect 17530 13574 17540 13608
rect 17540 13574 17574 13608
rect 17574 13574 17582 13608
rect 17530 13568 17582 13574
rect 17610 13608 17662 13620
rect 17610 13574 17620 13608
rect 17620 13574 17654 13608
rect 17654 13574 17662 13608
rect 17610 13568 17662 13574
rect 17814 13608 17866 13620
rect 17814 13574 17822 13608
rect 17822 13574 17856 13608
rect 17856 13574 17866 13608
rect 17814 13568 17866 13574
rect 17894 13608 17946 13620
rect 17894 13574 17902 13608
rect 17902 13574 17936 13608
rect 17936 13574 17946 13608
rect 17894 13568 17946 13574
rect 17974 13608 18026 13620
rect 17974 13574 17982 13608
rect 17982 13574 18016 13608
rect 18016 13574 18026 13608
rect 17974 13568 18026 13574
rect 18054 13608 18106 13620
rect 18054 13574 18062 13608
rect 18062 13574 18096 13608
rect 18096 13574 18106 13608
rect 18054 13568 18106 13574
rect 18134 13608 18186 13620
rect 18134 13574 18142 13608
rect 18142 13574 18176 13608
rect 18176 13574 18186 13608
rect 18134 13568 18186 13574
rect 18214 13608 18266 13620
rect 18214 13574 18222 13608
rect 18222 13574 18256 13608
rect 18256 13574 18266 13608
rect 18214 13568 18266 13574
rect 18422 13608 18474 13620
rect 18422 13574 18432 13608
rect 18432 13574 18466 13608
rect 18466 13574 18474 13608
rect 18422 13568 18474 13574
rect 18502 13608 18554 13620
rect 18502 13574 18512 13608
rect 18512 13574 18546 13608
rect 18546 13574 18554 13608
rect 18502 13568 18554 13574
rect 18582 13608 18634 13620
rect 18582 13574 18592 13608
rect 18592 13574 18626 13608
rect 18626 13574 18634 13608
rect 18582 13568 18634 13574
rect 18662 13608 18714 13620
rect 18662 13574 18672 13608
rect 18672 13574 18706 13608
rect 18706 13574 18714 13608
rect 18662 13568 18714 13574
rect 18742 13608 18794 13620
rect 18742 13574 18752 13608
rect 18752 13574 18786 13608
rect 18786 13574 18794 13608
rect 18742 13568 18794 13574
rect 18822 13608 18874 13620
rect 18822 13574 18832 13608
rect 18832 13574 18866 13608
rect 18866 13574 18874 13608
rect 18822 13568 18874 13574
rect 19026 13608 19078 13620
rect 19026 13574 19034 13608
rect 19034 13574 19068 13608
rect 19068 13574 19078 13608
rect 19026 13568 19078 13574
rect 19106 13608 19158 13620
rect 19106 13574 19114 13608
rect 19114 13574 19148 13608
rect 19148 13574 19158 13608
rect 19106 13568 19158 13574
rect 19186 13608 19238 13620
rect 19186 13574 19194 13608
rect 19194 13574 19228 13608
rect 19228 13574 19238 13608
rect 19186 13568 19238 13574
rect 19266 13608 19318 13620
rect 19266 13574 19274 13608
rect 19274 13574 19308 13608
rect 19308 13574 19318 13608
rect 19266 13568 19318 13574
rect 19346 13608 19398 13620
rect 19346 13574 19354 13608
rect 19354 13574 19388 13608
rect 19388 13574 19398 13608
rect 19346 13568 19398 13574
rect 19426 13608 19478 13620
rect 19426 13574 19434 13608
rect 19434 13574 19468 13608
rect 19468 13574 19478 13608
rect 19426 13568 19478 13574
rect 19765 13557 19817 13564
rect 19765 13523 19776 13557
rect 19776 13523 19810 13557
rect 19810 13523 19817 13557
rect 19765 13512 19817 13523
rect 20242 13560 20294 13567
rect 20242 13526 20253 13560
rect 20253 13526 20287 13560
rect 20287 13526 20294 13560
rect 20242 13515 20294 13526
rect 20665 13574 20717 13626
rect 20763 13605 20815 13617
rect 20763 13571 20773 13605
rect 20773 13571 20807 13605
rect 20807 13571 20815 13605
rect 20763 13565 20815 13571
rect 20843 13605 20895 13617
rect 20843 13571 20853 13605
rect 20853 13571 20887 13605
rect 20887 13571 20895 13605
rect 20843 13565 20895 13571
rect 20923 13605 20975 13617
rect 20923 13571 20933 13605
rect 20933 13571 20967 13605
rect 20967 13571 20975 13605
rect 20923 13565 20975 13571
rect 21003 13605 21055 13617
rect 21003 13571 21013 13605
rect 21013 13571 21047 13605
rect 21047 13571 21055 13605
rect 21003 13565 21055 13571
rect 21083 13605 21135 13617
rect 21083 13571 21093 13605
rect 21093 13571 21127 13605
rect 21127 13571 21135 13605
rect 21083 13565 21135 13571
rect 21163 13605 21215 13617
rect 21163 13571 21173 13605
rect 21173 13571 21207 13605
rect 21207 13571 21215 13605
rect 21163 13565 21215 13571
rect 21495 13608 21547 13620
rect 21495 13574 21505 13608
rect 21505 13574 21539 13608
rect 21539 13574 21547 13608
rect 21495 13568 21547 13574
rect 21575 13608 21627 13620
rect 21575 13574 21585 13608
rect 21585 13574 21619 13608
rect 21619 13574 21627 13608
rect 21575 13568 21627 13574
rect 21655 13608 21707 13620
rect 21655 13574 21665 13608
rect 21665 13574 21699 13608
rect 21699 13574 21707 13608
rect 21655 13568 21707 13574
rect 21735 13608 21787 13620
rect 21735 13574 21745 13608
rect 21745 13574 21779 13608
rect 21779 13574 21787 13608
rect 21735 13568 21787 13574
rect 21815 13608 21867 13620
rect 21815 13574 21825 13608
rect 21825 13574 21859 13608
rect 21859 13574 21867 13608
rect 21815 13568 21867 13574
rect 21895 13608 21947 13620
rect 21895 13574 21905 13608
rect 21905 13574 21939 13608
rect 21939 13574 21947 13608
rect 21895 13568 21947 13574
rect 22099 13608 22151 13620
rect 22099 13574 22107 13608
rect 22107 13574 22141 13608
rect 22141 13574 22151 13608
rect 22099 13568 22151 13574
rect 22179 13608 22231 13620
rect 22179 13574 22187 13608
rect 22187 13574 22221 13608
rect 22221 13574 22231 13608
rect 22179 13568 22231 13574
rect 22259 13608 22311 13620
rect 22259 13574 22267 13608
rect 22267 13574 22301 13608
rect 22301 13574 22311 13608
rect 22259 13568 22311 13574
rect 22339 13608 22391 13620
rect 22339 13574 22347 13608
rect 22347 13574 22381 13608
rect 22381 13574 22391 13608
rect 22339 13568 22391 13574
rect 22419 13608 22471 13620
rect 22419 13574 22427 13608
rect 22427 13574 22461 13608
rect 22461 13574 22471 13608
rect 22419 13568 22471 13574
rect 22499 13608 22551 13620
rect 22499 13574 22507 13608
rect 22507 13574 22541 13608
rect 22541 13574 22551 13608
rect 22499 13568 22551 13574
rect 22707 13608 22759 13620
rect 22707 13574 22717 13608
rect 22717 13574 22751 13608
rect 22751 13574 22759 13608
rect 22707 13568 22759 13574
rect 22787 13608 22839 13620
rect 22787 13574 22797 13608
rect 22797 13574 22831 13608
rect 22831 13574 22839 13608
rect 22787 13568 22839 13574
rect 22867 13608 22919 13620
rect 22867 13574 22877 13608
rect 22877 13574 22911 13608
rect 22911 13574 22919 13608
rect 22867 13568 22919 13574
rect 22947 13608 22999 13620
rect 22947 13574 22957 13608
rect 22957 13574 22991 13608
rect 22991 13574 22999 13608
rect 22947 13568 22999 13574
rect 23027 13608 23079 13620
rect 23027 13574 23037 13608
rect 23037 13574 23071 13608
rect 23071 13574 23079 13608
rect 23027 13568 23079 13574
rect 23107 13608 23159 13620
rect 23107 13574 23117 13608
rect 23117 13574 23151 13608
rect 23151 13574 23159 13608
rect 23107 13568 23159 13574
rect 23311 13608 23363 13620
rect 23311 13574 23319 13608
rect 23319 13574 23353 13608
rect 23353 13574 23363 13608
rect 23311 13568 23363 13574
rect 23391 13608 23443 13620
rect 23391 13574 23399 13608
rect 23399 13574 23433 13608
rect 23433 13574 23443 13608
rect 23391 13568 23443 13574
rect 23471 13608 23523 13620
rect 23471 13574 23479 13608
rect 23479 13574 23513 13608
rect 23513 13574 23523 13608
rect 23471 13568 23523 13574
rect 23551 13608 23603 13620
rect 23551 13574 23559 13608
rect 23559 13574 23593 13608
rect 23593 13574 23603 13608
rect 23551 13568 23603 13574
rect 23631 13608 23683 13620
rect 23631 13574 23639 13608
rect 23639 13574 23673 13608
rect 23673 13574 23683 13608
rect 23631 13568 23683 13574
rect 23711 13608 23763 13620
rect 23711 13574 23719 13608
rect 23719 13574 23753 13608
rect 23753 13574 23763 13608
rect 23711 13568 23763 13574
rect 23919 13608 23971 13620
rect 23919 13574 23929 13608
rect 23929 13574 23963 13608
rect 23963 13574 23971 13608
rect 23919 13568 23971 13574
rect 23999 13608 24051 13620
rect 23999 13574 24009 13608
rect 24009 13574 24043 13608
rect 24043 13574 24051 13608
rect 23999 13568 24051 13574
rect 24079 13608 24131 13620
rect 24079 13574 24089 13608
rect 24089 13574 24123 13608
rect 24123 13574 24131 13608
rect 24079 13568 24131 13574
rect 24159 13608 24211 13620
rect 24159 13574 24169 13608
rect 24169 13574 24203 13608
rect 24203 13574 24211 13608
rect 24159 13568 24211 13574
rect 24239 13608 24291 13620
rect 24239 13574 24249 13608
rect 24249 13574 24283 13608
rect 24283 13574 24291 13608
rect 24239 13568 24291 13574
rect 24319 13608 24371 13620
rect 24319 13574 24329 13608
rect 24329 13574 24363 13608
rect 24363 13574 24371 13608
rect 24319 13568 24371 13574
rect 24523 13608 24575 13620
rect 24523 13574 24531 13608
rect 24531 13574 24565 13608
rect 24565 13574 24575 13608
rect 24523 13568 24575 13574
rect 24603 13608 24655 13620
rect 24603 13574 24611 13608
rect 24611 13574 24645 13608
rect 24645 13574 24655 13608
rect 24603 13568 24655 13574
rect 24683 13608 24735 13620
rect 24683 13574 24691 13608
rect 24691 13574 24725 13608
rect 24725 13574 24735 13608
rect 24683 13568 24735 13574
rect 24763 13608 24815 13620
rect 24763 13574 24771 13608
rect 24771 13574 24805 13608
rect 24805 13574 24815 13608
rect 24763 13568 24815 13574
rect 24843 13608 24895 13620
rect 24843 13574 24851 13608
rect 24851 13574 24885 13608
rect 24885 13574 24895 13608
rect 24843 13568 24895 13574
rect 24923 13608 24975 13620
rect 24923 13574 24931 13608
rect 24931 13574 24965 13608
rect 24965 13574 24975 13608
rect 24923 13568 24975 13574
rect 25131 13608 25183 13620
rect 25131 13574 25141 13608
rect 25141 13574 25175 13608
rect 25175 13574 25183 13608
rect 25131 13568 25183 13574
rect 25211 13608 25263 13620
rect 25211 13574 25221 13608
rect 25221 13574 25255 13608
rect 25255 13574 25263 13608
rect 25211 13568 25263 13574
rect 25291 13608 25343 13620
rect 25291 13574 25301 13608
rect 25301 13574 25335 13608
rect 25335 13574 25343 13608
rect 25291 13568 25343 13574
rect 25371 13608 25423 13620
rect 25371 13574 25381 13608
rect 25381 13574 25415 13608
rect 25415 13574 25423 13608
rect 25371 13568 25423 13574
rect 25451 13608 25503 13620
rect 25451 13574 25461 13608
rect 25461 13574 25495 13608
rect 25495 13574 25503 13608
rect 25451 13568 25503 13574
rect 25531 13608 25583 13620
rect 25531 13574 25541 13608
rect 25541 13574 25575 13608
rect 25575 13574 25583 13608
rect 25531 13568 25583 13574
rect 25735 13608 25787 13620
rect 25735 13574 25743 13608
rect 25743 13574 25777 13608
rect 25777 13574 25787 13608
rect 25735 13568 25787 13574
rect 25815 13608 25867 13620
rect 25815 13574 25823 13608
rect 25823 13574 25857 13608
rect 25857 13574 25867 13608
rect 25815 13568 25867 13574
rect 25895 13608 25947 13620
rect 25895 13574 25903 13608
rect 25903 13574 25937 13608
rect 25937 13574 25947 13608
rect 25895 13568 25947 13574
rect 25975 13608 26027 13620
rect 25975 13574 25983 13608
rect 25983 13574 26017 13608
rect 26017 13574 26027 13608
rect 25975 13568 26027 13574
rect 26055 13608 26107 13620
rect 26055 13574 26063 13608
rect 26063 13574 26097 13608
rect 26097 13574 26107 13608
rect 26055 13568 26107 13574
rect 26135 13608 26187 13620
rect 26135 13574 26143 13608
rect 26143 13574 26177 13608
rect 26177 13574 26187 13608
rect 26135 13568 26187 13574
rect 26474 13557 26526 13564
rect 26474 13523 26485 13557
rect 26485 13523 26519 13557
rect 26519 13523 26526 13557
rect 26474 13512 26526 13523
rect 19770 13413 19822 13420
rect 19770 13379 19781 13413
rect 19781 13379 19815 13413
rect 19815 13379 19822 13413
rect 19770 13368 19822 13379
rect 20231 13388 20283 13395
rect 20231 13354 20242 13388
rect 20242 13354 20276 13388
rect 20276 13354 20283 13388
rect 20231 13343 20283 13354
rect 19771 13261 19823 13268
rect 19771 13227 19782 13261
rect 19782 13227 19816 13261
rect 19816 13227 19823 13261
rect 19771 13216 19823 13227
rect 3068 13099 3120 13151
rect 3166 13130 3218 13142
rect 3166 13096 3176 13130
rect 3176 13096 3210 13130
rect 3210 13096 3218 13130
rect 3166 13090 3218 13096
rect 3246 13130 3298 13142
rect 3246 13096 3256 13130
rect 3256 13096 3290 13130
rect 3290 13096 3298 13130
rect 3246 13090 3298 13096
rect 3326 13130 3378 13142
rect 3326 13096 3336 13130
rect 3336 13096 3370 13130
rect 3370 13096 3378 13130
rect 3326 13090 3378 13096
rect 3406 13130 3458 13142
rect 3406 13096 3416 13130
rect 3416 13096 3450 13130
rect 3450 13096 3458 13130
rect 3406 13090 3458 13096
rect 3486 13130 3538 13142
rect 3486 13096 3496 13130
rect 3496 13096 3530 13130
rect 3530 13096 3538 13130
rect 3486 13090 3538 13096
rect 3566 13130 3618 13142
rect 3566 13096 3576 13130
rect 3576 13096 3610 13130
rect 3610 13096 3618 13130
rect 3566 13090 3618 13096
rect 3898 13133 3950 13145
rect 3898 13099 3908 13133
rect 3908 13099 3942 13133
rect 3942 13099 3950 13133
rect 3898 13093 3950 13099
rect 3978 13133 4030 13145
rect 3978 13099 3988 13133
rect 3988 13099 4022 13133
rect 4022 13099 4030 13133
rect 3978 13093 4030 13099
rect 4058 13133 4110 13145
rect 4058 13099 4068 13133
rect 4068 13099 4102 13133
rect 4102 13099 4110 13133
rect 4058 13093 4110 13099
rect 4138 13133 4190 13145
rect 4138 13099 4148 13133
rect 4148 13099 4182 13133
rect 4182 13099 4190 13133
rect 4138 13093 4190 13099
rect 4218 13133 4270 13145
rect 4218 13099 4228 13133
rect 4228 13099 4262 13133
rect 4262 13099 4270 13133
rect 4218 13093 4270 13099
rect 4298 13133 4350 13145
rect 4298 13099 4308 13133
rect 4308 13099 4342 13133
rect 4342 13099 4350 13133
rect 4298 13093 4350 13099
rect 4502 13133 4554 13145
rect 4502 13099 4510 13133
rect 4510 13099 4544 13133
rect 4544 13099 4554 13133
rect 4502 13093 4554 13099
rect 4582 13133 4634 13145
rect 4582 13099 4590 13133
rect 4590 13099 4624 13133
rect 4624 13099 4634 13133
rect 4582 13093 4634 13099
rect 4662 13133 4714 13145
rect 4662 13099 4670 13133
rect 4670 13099 4704 13133
rect 4704 13099 4714 13133
rect 4662 13093 4714 13099
rect 4742 13133 4794 13145
rect 4742 13099 4750 13133
rect 4750 13099 4784 13133
rect 4784 13099 4794 13133
rect 4742 13093 4794 13099
rect 4822 13133 4874 13145
rect 4822 13099 4830 13133
rect 4830 13099 4864 13133
rect 4864 13099 4874 13133
rect 4822 13093 4874 13099
rect 4902 13133 4954 13145
rect 4902 13099 4910 13133
rect 4910 13099 4944 13133
rect 4944 13099 4954 13133
rect 4902 13093 4954 13099
rect 5110 13133 5162 13145
rect 5110 13099 5120 13133
rect 5120 13099 5154 13133
rect 5154 13099 5162 13133
rect 5110 13093 5162 13099
rect 5190 13133 5242 13145
rect 5190 13099 5200 13133
rect 5200 13099 5234 13133
rect 5234 13099 5242 13133
rect 5190 13093 5242 13099
rect 5270 13133 5322 13145
rect 5270 13099 5280 13133
rect 5280 13099 5314 13133
rect 5314 13099 5322 13133
rect 5270 13093 5322 13099
rect 5350 13133 5402 13145
rect 5350 13099 5360 13133
rect 5360 13099 5394 13133
rect 5394 13099 5402 13133
rect 5350 13093 5402 13099
rect 5430 13133 5482 13145
rect 5430 13099 5440 13133
rect 5440 13099 5474 13133
rect 5474 13099 5482 13133
rect 5430 13093 5482 13099
rect 5510 13133 5562 13145
rect 5510 13099 5520 13133
rect 5520 13099 5554 13133
rect 5554 13099 5562 13133
rect 5510 13093 5562 13099
rect 5714 13133 5766 13145
rect 5714 13099 5722 13133
rect 5722 13099 5756 13133
rect 5756 13099 5766 13133
rect 5714 13093 5766 13099
rect 5794 13133 5846 13145
rect 5794 13099 5802 13133
rect 5802 13099 5836 13133
rect 5836 13099 5846 13133
rect 5794 13093 5846 13099
rect 5874 13133 5926 13145
rect 5874 13099 5882 13133
rect 5882 13099 5916 13133
rect 5916 13099 5926 13133
rect 5874 13093 5926 13099
rect 5954 13133 6006 13145
rect 5954 13099 5962 13133
rect 5962 13099 5996 13133
rect 5996 13099 6006 13133
rect 5954 13093 6006 13099
rect 6034 13133 6086 13145
rect 6034 13099 6042 13133
rect 6042 13099 6076 13133
rect 6076 13099 6086 13133
rect 6034 13093 6086 13099
rect 6114 13133 6166 13145
rect 6114 13099 6122 13133
rect 6122 13099 6156 13133
rect 6156 13099 6166 13133
rect 6114 13093 6166 13099
rect 6322 13133 6374 13145
rect 6322 13099 6332 13133
rect 6332 13099 6366 13133
rect 6366 13099 6374 13133
rect 6322 13093 6374 13099
rect 6402 13133 6454 13145
rect 6402 13099 6412 13133
rect 6412 13099 6446 13133
rect 6446 13099 6454 13133
rect 6402 13093 6454 13099
rect 6482 13133 6534 13145
rect 6482 13099 6492 13133
rect 6492 13099 6526 13133
rect 6526 13099 6534 13133
rect 6482 13093 6534 13099
rect 6562 13133 6614 13145
rect 6562 13099 6572 13133
rect 6572 13099 6606 13133
rect 6606 13099 6614 13133
rect 6562 13093 6614 13099
rect 6642 13133 6694 13145
rect 6642 13099 6652 13133
rect 6652 13099 6686 13133
rect 6686 13099 6694 13133
rect 6642 13093 6694 13099
rect 6722 13133 6774 13145
rect 6722 13099 6732 13133
rect 6732 13099 6766 13133
rect 6766 13099 6774 13133
rect 6722 13093 6774 13099
rect 6926 13133 6978 13145
rect 6926 13099 6934 13133
rect 6934 13099 6968 13133
rect 6968 13099 6978 13133
rect 6926 13093 6978 13099
rect 7006 13133 7058 13145
rect 7006 13099 7014 13133
rect 7014 13099 7048 13133
rect 7048 13099 7058 13133
rect 7006 13093 7058 13099
rect 7086 13133 7138 13145
rect 7086 13099 7094 13133
rect 7094 13099 7128 13133
rect 7128 13099 7138 13133
rect 7086 13093 7138 13099
rect 7166 13133 7218 13145
rect 7166 13099 7174 13133
rect 7174 13099 7208 13133
rect 7208 13099 7218 13133
rect 7166 13093 7218 13099
rect 7246 13133 7298 13145
rect 7246 13099 7254 13133
rect 7254 13099 7288 13133
rect 7288 13099 7298 13133
rect 7246 13093 7298 13099
rect 7326 13133 7378 13145
rect 7326 13099 7334 13133
rect 7334 13099 7368 13133
rect 7368 13099 7378 13133
rect 7326 13093 7378 13099
rect 7534 13133 7586 13145
rect 7534 13099 7544 13133
rect 7544 13099 7578 13133
rect 7578 13099 7586 13133
rect 7534 13093 7586 13099
rect 7614 13133 7666 13145
rect 7614 13099 7624 13133
rect 7624 13099 7658 13133
rect 7658 13099 7666 13133
rect 7614 13093 7666 13099
rect 7694 13133 7746 13145
rect 7694 13099 7704 13133
rect 7704 13099 7738 13133
rect 7738 13099 7746 13133
rect 7694 13093 7746 13099
rect 7774 13133 7826 13145
rect 7774 13099 7784 13133
rect 7784 13099 7818 13133
rect 7818 13099 7826 13133
rect 7774 13093 7826 13099
rect 7854 13133 7906 13145
rect 7854 13099 7864 13133
rect 7864 13099 7898 13133
rect 7898 13099 7906 13133
rect 7854 13093 7906 13099
rect 7934 13133 7986 13145
rect 7934 13099 7944 13133
rect 7944 13099 7978 13133
rect 7978 13099 7986 13133
rect 7934 13093 7986 13099
rect 8138 13133 8190 13145
rect 8138 13099 8146 13133
rect 8146 13099 8180 13133
rect 8180 13099 8190 13133
rect 8138 13093 8190 13099
rect 8218 13133 8270 13145
rect 8218 13099 8226 13133
rect 8226 13099 8260 13133
rect 8260 13099 8270 13133
rect 8218 13093 8270 13099
rect 8298 13133 8350 13145
rect 8298 13099 8306 13133
rect 8306 13099 8340 13133
rect 8340 13099 8350 13133
rect 8298 13093 8350 13099
rect 8378 13133 8430 13145
rect 8378 13099 8386 13133
rect 8386 13099 8420 13133
rect 8420 13099 8430 13133
rect 8378 13093 8430 13099
rect 8458 13133 8510 13145
rect 8458 13099 8466 13133
rect 8466 13099 8500 13133
rect 8500 13099 8510 13133
rect 8458 13093 8510 13099
rect 8538 13133 8590 13145
rect 8538 13099 8546 13133
rect 8546 13099 8580 13133
rect 8580 13099 8590 13133
rect 8538 13093 8590 13099
rect 20231 13196 20283 13203
rect 20231 13162 20242 13196
rect 20242 13162 20276 13196
rect 20276 13162 20283 13196
rect 20231 13151 20283 13162
rect 26479 13413 26531 13420
rect 26479 13379 26490 13413
rect 26490 13379 26524 13413
rect 26524 13379 26531 13413
rect 26479 13368 26531 13379
rect 26480 13261 26532 13268
rect 26480 13227 26491 13261
rect 26491 13227 26525 13261
rect 26525 13227 26532 13261
rect 26480 13216 26532 13227
rect 8877 13082 8929 13089
rect 8877 13048 8888 13082
rect 8888 13048 8922 13082
rect 8922 13048 8929 13082
rect 8877 13037 8929 13048
rect 13339 12969 13391 13021
rect 13470 13010 13522 13020
rect 13470 12976 13487 13010
rect 13487 12976 13521 13010
rect 13521 12976 13522 13010
rect 13470 12968 13522 12976
rect 13614 12969 13666 13021
rect 8882 12938 8934 12945
rect 8882 12904 8893 12938
rect 8893 12904 8927 12938
rect 8927 12904 8934 12938
rect 8882 12893 8934 12904
rect 19771 13091 19823 13098
rect 19771 13057 19782 13091
rect 19782 13057 19816 13091
rect 19816 13057 19823 13091
rect 19771 13046 19823 13057
rect 20048 12969 20100 13021
rect 20179 13010 20231 13020
rect 20179 12976 20196 13010
rect 20196 12976 20230 13010
rect 20230 12976 20231 13010
rect 20179 12968 20231 12976
rect 20323 12969 20375 13021
rect 8883 12786 8935 12793
rect 8883 12752 8894 12786
rect 8894 12752 8928 12786
rect 8928 12752 8935 12786
rect 8883 12741 8935 12752
rect 13612 12701 13664 12710
rect 13612 12667 13624 12701
rect 13624 12667 13658 12701
rect 13658 12667 13664 12701
rect 13612 12658 13664 12667
rect 2451 12494 2503 12546
rect 2582 12535 2634 12545
rect 2582 12501 2599 12535
rect 2599 12501 2633 12535
rect 2633 12501 2634 12535
rect 2582 12493 2634 12501
rect 2726 12494 2778 12546
rect 8883 12616 8935 12623
rect 8883 12582 8894 12616
rect 8894 12582 8928 12616
rect 8928 12582 8935 12616
rect 8883 12571 8935 12582
rect 19770 12934 19822 12941
rect 19770 12900 19781 12934
rect 19781 12900 19815 12934
rect 19815 12900 19822 12934
rect 19770 12889 19822 12900
rect 26480 13091 26532 13098
rect 26480 13057 26491 13091
rect 26491 13057 26525 13091
rect 26525 13057 26532 13091
rect 26480 13046 26532 13057
rect 10987 12502 11039 12554
rect 11174 12504 11226 12556
rect 11359 12506 11411 12558
rect 11544 12507 11596 12559
rect 11747 12509 11799 12561
rect 11932 12511 11984 12563
rect 12131 12513 12183 12565
rect 12333 12512 12385 12564
rect 12543 12515 12595 12567
rect 12767 12515 12819 12567
rect 12973 12514 13025 12566
rect 13194 12513 13246 12565
rect 2724 12226 2776 12235
rect 2724 12192 2736 12226
rect 2736 12192 2770 12226
rect 2770 12192 2776 12226
rect 2724 12183 2776 12192
rect 8882 12459 8934 12466
rect 8882 12425 8893 12459
rect 8893 12425 8927 12459
rect 8927 12425 8934 12459
rect 8882 12414 8934 12425
rect 13357 12466 13409 12475
rect 13477 12466 13529 12475
rect 13620 12466 13672 12475
rect 13357 12432 13395 12466
rect 13395 12432 13409 12466
rect 13477 12432 13487 12466
rect 13487 12432 13521 12466
rect 13521 12432 13529 12466
rect 13620 12432 13671 12466
rect 13671 12432 13672 12466
rect 13357 12423 13409 12432
rect 13477 12423 13529 12432
rect 13620 12423 13672 12432
rect 2469 11991 2521 12000
rect 2589 11991 2641 12000
rect 2732 11991 2784 12000
rect 2469 11957 2507 11991
rect 2507 11957 2521 11991
rect 2589 11957 2599 11991
rect 2599 11957 2633 11991
rect 2633 11957 2641 11991
rect 2732 11957 2783 11991
rect 2783 11957 2784 11991
rect 2469 11948 2521 11957
rect 2589 11948 2641 11957
rect 2732 11948 2784 11957
rect 2736 11605 2788 11657
rect 8800 12172 8852 12224
rect 9177 12224 9229 12276
rect 11638 12296 11690 12311
rect 11638 12262 11648 12296
rect 11648 12262 11682 12296
rect 11682 12262 11690 12296
rect 11638 12259 11690 12262
rect 11256 12189 11308 12197
rect 11256 12155 11263 12189
rect 11263 12155 11297 12189
rect 11297 12155 11308 12189
rect 11256 12145 11308 12155
rect 12759 12225 12811 12239
rect 12759 12191 12768 12225
rect 12768 12191 12802 12225
rect 12802 12191 12811 12225
rect 12759 12186 12811 12191
rect 13624 12080 13676 12132
rect 19688 12647 19740 12699
rect 20321 12701 20373 12710
rect 20321 12667 20333 12701
rect 20333 12667 20367 12701
rect 20367 12667 20373 12701
rect 20321 12658 20373 12667
rect 26479 12934 26531 12941
rect 26479 12900 26490 12934
rect 26490 12900 26524 12934
rect 26524 12900 26531 12934
rect 26479 12889 26531 12900
rect 14436 12436 14500 12439
rect 14436 12376 14458 12436
rect 14458 12376 14492 12436
rect 14492 12376 14500 12436
rect 14436 12375 14500 12376
rect 15168 12439 15232 12442
rect 15168 12379 15190 12439
rect 15190 12379 15224 12439
rect 15224 12379 15232 12439
rect 15168 12378 15232 12379
rect 15396 12439 15460 12442
rect 15396 12379 15404 12439
rect 15404 12379 15438 12439
rect 15438 12379 15460 12439
rect 15396 12378 15460 12379
rect 16380 12439 16444 12442
rect 16380 12379 16402 12439
rect 16402 12379 16436 12439
rect 16436 12379 16444 12439
rect 16380 12378 16444 12379
rect 16608 12439 16672 12442
rect 16608 12379 16616 12439
rect 16616 12379 16650 12439
rect 16650 12379 16672 12439
rect 16608 12378 16672 12379
rect 17592 12439 17656 12442
rect 17592 12379 17614 12439
rect 17614 12379 17648 12439
rect 17648 12379 17656 12439
rect 17592 12378 17656 12379
rect 17820 12439 17884 12442
rect 17820 12379 17828 12439
rect 17828 12379 17862 12439
rect 17862 12379 17884 12439
rect 17820 12378 17884 12379
rect 18804 12439 18868 12442
rect 18804 12379 18826 12439
rect 18826 12379 18860 12439
rect 18860 12379 18868 12439
rect 18804 12378 18868 12379
rect 19032 12439 19096 12442
rect 19032 12379 19040 12439
rect 19040 12379 19074 12439
rect 19074 12379 19096 12439
rect 19032 12378 19096 12379
rect 19776 12386 19785 12438
rect 19785 12386 19819 12438
rect 19819 12386 19828 12438
rect 20066 12466 20118 12475
rect 20186 12466 20238 12475
rect 20329 12466 20381 12475
rect 20066 12432 20104 12466
rect 20104 12432 20118 12466
rect 20186 12432 20196 12466
rect 20196 12432 20230 12466
rect 20230 12432 20238 12466
rect 20329 12432 20380 12466
rect 20380 12432 20381 12466
rect 20066 12423 20118 12432
rect 20186 12423 20238 12432
rect 20329 12423 20381 12432
rect 14792 12238 14856 12240
rect 14792 12178 14811 12238
rect 14811 12178 14845 12238
rect 14845 12178 14856 12238
rect 14792 12176 14856 12178
rect 15524 12238 15588 12240
rect 15524 12178 15543 12238
rect 15543 12178 15577 12238
rect 15577 12178 15588 12238
rect 15524 12176 15588 12178
rect 15742 12238 15806 12240
rect 15742 12178 15753 12238
rect 15753 12178 15787 12238
rect 15787 12178 15806 12238
rect 15742 12176 15806 12178
rect 16736 12238 16800 12240
rect 16736 12178 16755 12238
rect 16755 12178 16789 12238
rect 16789 12178 16800 12238
rect 16736 12176 16800 12178
rect 16954 12238 17018 12240
rect 16954 12178 16965 12238
rect 16965 12178 16999 12238
rect 16999 12178 17018 12238
rect 16954 12176 17018 12178
rect 18074 12238 18138 12240
rect 18074 12178 18093 12238
rect 18093 12178 18127 12238
rect 18127 12178 18138 12238
rect 18074 12176 18138 12178
rect 18292 12238 18356 12240
rect 18292 12178 18303 12238
rect 18303 12178 18337 12238
rect 18337 12178 18356 12238
rect 18292 12176 18356 12178
rect 19026 12238 19090 12240
rect 19026 12178 19037 12238
rect 19037 12178 19071 12238
rect 19071 12178 19090 12238
rect 19026 12176 19090 12178
rect 19776 12183 19785 12235
rect 19785 12183 19819 12235
rect 19819 12183 19828 12235
rect 14112 12080 14164 12132
rect 3548 11961 3612 11964
rect 3548 11901 3570 11961
rect 3570 11901 3604 11961
rect 3604 11901 3612 11961
rect 3548 11900 3612 11901
rect 4280 11964 4344 11967
rect 4280 11904 4302 11964
rect 4302 11904 4336 11964
rect 4336 11904 4344 11964
rect 4280 11903 4344 11904
rect 4508 11964 4572 11967
rect 4508 11904 4516 11964
rect 4516 11904 4550 11964
rect 4550 11904 4572 11964
rect 4508 11903 4572 11904
rect 5492 11964 5556 11967
rect 5492 11904 5514 11964
rect 5514 11904 5548 11964
rect 5548 11904 5556 11964
rect 5492 11903 5556 11904
rect 5720 11964 5784 11967
rect 5720 11904 5728 11964
rect 5728 11904 5762 11964
rect 5762 11904 5784 11964
rect 5720 11903 5784 11904
rect 6704 11964 6768 11967
rect 6704 11904 6726 11964
rect 6726 11904 6760 11964
rect 6760 11904 6768 11964
rect 6704 11903 6768 11904
rect 6932 11964 6996 11967
rect 6932 11904 6940 11964
rect 6940 11904 6974 11964
rect 6974 11904 6996 11964
rect 6932 11903 6996 11904
rect 7916 11964 7980 11967
rect 7916 11904 7938 11964
rect 7938 11904 7972 11964
rect 7972 11904 7980 11964
rect 7916 11903 7980 11904
rect 8144 11964 8208 11967
rect 8144 11904 8152 11964
rect 8152 11904 8186 11964
rect 8186 11904 8208 11964
rect 8144 11903 8208 11904
rect 8888 11911 8897 11963
rect 8897 11911 8931 11963
rect 8931 11911 8940 11963
rect 11264 11981 11317 12033
rect 13205 12044 13257 12054
rect 13205 12010 13215 12044
rect 13215 12010 13249 12044
rect 13249 12010 13257 12044
rect 13205 12002 13257 12010
rect 3904 11763 3968 11765
rect 3904 11703 3923 11763
rect 3923 11703 3957 11763
rect 3957 11703 3968 11763
rect 3904 11701 3968 11703
rect 4636 11763 4700 11765
rect 4636 11703 4655 11763
rect 4655 11703 4689 11763
rect 4689 11703 4700 11763
rect 4636 11701 4700 11703
rect 4854 11763 4918 11765
rect 4854 11703 4865 11763
rect 4865 11703 4899 11763
rect 4899 11703 4918 11763
rect 4854 11701 4918 11703
rect 5848 11763 5912 11765
rect 5848 11703 5867 11763
rect 5867 11703 5901 11763
rect 5901 11703 5912 11763
rect 5848 11701 5912 11703
rect 6066 11763 6130 11765
rect 6066 11703 6077 11763
rect 6077 11703 6111 11763
rect 6111 11703 6130 11763
rect 6066 11701 6130 11703
rect 7186 11763 7250 11765
rect 7186 11703 7205 11763
rect 7205 11703 7239 11763
rect 7239 11703 7250 11763
rect 7186 11701 7250 11703
rect 7404 11763 7468 11765
rect 7404 11703 7415 11763
rect 7415 11703 7449 11763
rect 7449 11703 7468 11763
rect 7404 11701 7468 11703
rect 10298 11808 10352 11862
rect 10917 11829 10970 11882
rect 11117 11832 11170 11885
rect 11353 11830 11406 11883
rect 11786 11824 11839 11877
rect 11987 11825 12040 11878
rect 12173 11823 12226 11876
rect 12364 11826 12417 11879
rect 12577 11825 12630 11878
rect 8138 11763 8202 11765
rect 8138 11703 8149 11763
rect 8149 11703 8183 11763
rect 8183 11703 8202 11763
rect 8138 11701 8202 11703
rect 8888 11708 8897 11760
rect 8897 11708 8931 11760
rect 8931 11708 8940 11760
rect 12761 11693 12813 11745
rect 3224 11605 3276 11657
rect 3054 10553 3063 10573
rect 3063 10553 3097 10573
rect 3097 10553 3106 10573
rect 3054 10521 3106 10553
rect 3596 10566 3648 10576
rect 3596 10532 3604 10566
rect 3604 10532 3638 10566
rect 3638 10532 3648 10566
rect 3596 10524 3648 10532
rect 3676 10566 3728 10576
rect 3676 10532 3684 10566
rect 3684 10532 3718 10566
rect 3718 10532 3728 10566
rect 3676 10524 3728 10532
rect 3756 10566 3808 10576
rect 3756 10532 3764 10566
rect 3764 10532 3798 10566
rect 3798 10532 3808 10566
rect 3756 10524 3808 10532
rect 3836 10566 3888 10576
rect 3836 10532 3844 10566
rect 3844 10532 3878 10566
rect 3878 10532 3888 10566
rect 3836 10524 3888 10532
rect 4328 10566 4380 10576
rect 4328 10532 4336 10566
rect 4336 10532 4370 10566
rect 4370 10532 4380 10566
rect 4328 10524 4380 10532
rect 4408 10566 4460 10576
rect 4408 10532 4416 10566
rect 4416 10532 4450 10566
rect 4450 10532 4460 10566
rect 4408 10524 4460 10532
rect 4488 10566 4540 10576
rect 4488 10532 4496 10566
rect 4496 10532 4530 10566
rect 4530 10532 4540 10566
rect 4488 10524 4540 10532
rect 4568 10566 4620 10576
rect 4568 10532 4576 10566
rect 4576 10532 4610 10566
rect 4610 10532 4620 10566
rect 4568 10524 4620 10532
rect 4934 10566 4986 10576
rect 4934 10532 4944 10566
rect 4944 10532 4978 10566
rect 4978 10532 4986 10566
rect 4934 10524 4986 10532
rect 5014 10566 5066 10576
rect 5014 10532 5024 10566
rect 5024 10532 5058 10566
rect 5058 10532 5066 10566
rect 5014 10524 5066 10532
rect 5094 10566 5146 10576
rect 5094 10532 5104 10566
rect 5104 10532 5138 10566
rect 5138 10532 5146 10566
rect 5094 10524 5146 10532
rect 5174 10566 5226 10576
rect 5174 10532 5184 10566
rect 5184 10532 5218 10566
rect 5218 10532 5226 10566
rect 5174 10524 5226 10532
rect 5540 10566 5592 10576
rect 5540 10532 5548 10566
rect 5548 10532 5582 10566
rect 5582 10532 5592 10566
rect 5540 10524 5592 10532
rect 5620 10566 5672 10576
rect 5620 10532 5628 10566
rect 5628 10532 5662 10566
rect 5662 10532 5672 10566
rect 5620 10524 5672 10532
rect 5700 10566 5752 10576
rect 5700 10532 5708 10566
rect 5708 10532 5742 10566
rect 5742 10532 5752 10566
rect 5700 10524 5752 10532
rect 5780 10566 5832 10576
rect 5780 10532 5788 10566
rect 5788 10532 5822 10566
rect 5822 10532 5832 10566
rect 5780 10524 5832 10532
rect 6146 10566 6198 10576
rect 6146 10532 6156 10566
rect 6156 10532 6190 10566
rect 6190 10532 6198 10566
rect 6146 10524 6198 10532
rect 6226 10566 6278 10576
rect 6226 10532 6236 10566
rect 6236 10532 6270 10566
rect 6270 10532 6278 10566
rect 6226 10524 6278 10532
rect 6306 10566 6358 10576
rect 6306 10532 6316 10566
rect 6316 10532 6350 10566
rect 6350 10532 6358 10566
rect 6306 10524 6358 10532
rect 6386 10566 6438 10576
rect 6386 10532 6396 10566
rect 6396 10532 6430 10566
rect 6430 10532 6438 10566
rect 6386 10524 6438 10532
rect 6878 10566 6930 10576
rect 6878 10532 6886 10566
rect 6886 10532 6920 10566
rect 6920 10532 6930 10566
rect 6878 10524 6930 10532
rect 6958 10566 7010 10576
rect 6958 10532 6966 10566
rect 6966 10532 7000 10566
rect 7000 10532 7010 10566
rect 6958 10524 7010 10532
rect 7038 10566 7090 10576
rect 7038 10532 7046 10566
rect 7046 10532 7080 10566
rect 7080 10532 7090 10566
rect 7038 10524 7090 10532
rect 7118 10566 7170 10576
rect 7118 10532 7126 10566
rect 7126 10532 7160 10566
rect 7160 10532 7170 10566
rect 7118 10524 7170 10532
rect 7484 10566 7536 10576
rect 7484 10532 7494 10566
rect 7494 10532 7528 10566
rect 7528 10532 7536 10566
rect 7484 10524 7536 10532
rect 7564 10566 7616 10576
rect 7564 10532 7574 10566
rect 7574 10532 7608 10566
rect 7608 10532 7616 10566
rect 7564 10524 7616 10532
rect 7644 10566 7696 10576
rect 7644 10532 7654 10566
rect 7654 10532 7688 10566
rect 7688 10532 7696 10566
rect 7644 10524 7696 10532
rect 7724 10566 7776 10576
rect 7724 10532 7734 10566
rect 7734 10532 7768 10566
rect 7768 10532 7776 10566
rect 7724 10524 7776 10532
rect 11634 11620 11686 11672
rect 13317 11543 13375 11594
rect 13375 11543 13377 11594
rect 13317 11538 13377 11543
rect 8797 11446 8849 11498
rect 9200 11467 9252 11519
rect 10935 11248 10945 11257
rect 10945 11248 10987 11257
rect 11123 11248 11129 11254
rect 11129 11248 11175 11254
rect 11320 11248 11371 11252
rect 11371 11248 11372 11252
rect 10935 11205 10987 11248
rect 11123 11202 11175 11248
rect 11320 11200 11372 11248
rect 13942 11028 13951 11048
rect 13951 11028 13985 11048
rect 13985 11028 13994 11048
rect 13942 10996 13994 11028
rect 14484 11041 14536 11051
rect 14484 11007 14492 11041
rect 14492 11007 14526 11041
rect 14526 11007 14536 11041
rect 14484 10999 14536 11007
rect 14564 11041 14616 11051
rect 14564 11007 14572 11041
rect 14572 11007 14606 11041
rect 14606 11007 14616 11041
rect 14564 10999 14616 11007
rect 14644 11041 14696 11051
rect 14644 11007 14652 11041
rect 14652 11007 14686 11041
rect 14686 11007 14696 11041
rect 14644 10999 14696 11007
rect 14724 11041 14776 11051
rect 14724 11007 14732 11041
rect 14732 11007 14766 11041
rect 14766 11007 14776 11041
rect 14724 10999 14776 11007
rect 15216 11041 15268 11051
rect 15216 11007 15224 11041
rect 15224 11007 15258 11041
rect 15258 11007 15268 11041
rect 15216 10999 15268 11007
rect 15296 11041 15348 11051
rect 15296 11007 15304 11041
rect 15304 11007 15338 11041
rect 15338 11007 15348 11041
rect 15296 10999 15348 11007
rect 15376 11041 15428 11051
rect 15376 11007 15384 11041
rect 15384 11007 15418 11041
rect 15418 11007 15428 11041
rect 15376 10999 15428 11007
rect 15456 11041 15508 11051
rect 15456 11007 15464 11041
rect 15464 11007 15498 11041
rect 15498 11007 15508 11041
rect 15456 10999 15508 11007
rect 15822 11041 15874 11051
rect 15822 11007 15832 11041
rect 15832 11007 15866 11041
rect 15866 11007 15874 11041
rect 15822 10999 15874 11007
rect 15902 11041 15954 11051
rect 15902 11007 15912 11041
rect 15912 11007 15946 11041
rect 15946 11007 15954 11041
rect 15902 10999 15954 11007
rect 15982 11041 16034 11051
rect 15982 11007 15992 11041
rect 15992 11007 16026 11041
rect 16026 11007 16034 11041
rect 15982 10999 16034 11007
rect 16062 11041 16114 11051
rect 16062 11007 16072 11041
rect 16072 11007 16106 11041
rect 16106 11007 16114 11041
rect 16062 10999 16114 11007
rect 16428 11041 16480 11051
rect 16428 11007 16436 11041
rect 16436 11007 16470 11041
rect 16470 11007 16480 11041
rect 16428 10999 16480 11007
rect 16508 11041 16560 11051
rect 16508 11007 16516 11041
rect 16516 11007 16550 11041
rect 16550 11007 16560 11041
rect 16508 10999 16560 11007
rect 16588 11041 16640 11051
rect 16588 11007 16596 11041
rect 16596 11007 16630 11041
rect 16630 11007 16640 11041
rect 16588 10999 16640 11007
rect 16668 11041 16720 11051
rect 16668 11007 16676 11041
rect 16676 11007 16710 11041
rect 16710 11007 16720 11041
rect 16668 10999 16720 11007
rect 17034 11041 17086 11051
rect 17034 11007 17044 11041
rect 17044 11007 17078 11041
rect 17078 11007 17086 11041
rect 17034 10999 17086 11007
rect 17114 11041 17166 11051
rect 17114 11007 17124 11041
rect 17124 11007 17158 11041
rect 17158 11007 17166 11041
rect 17114 10999 17166 11007
rect 17194 11041 17246 11051
rect 17194 11007 17204 11041
rect 17204 11007 17238 11041
rect 17238 11007 17246 11041
rect 17194 10999 17246 11007
rect 17274 11041 17326 11051
rect 17274 11007 17284 11041
rect 17284 11007 17318 11041
rect 17318 11007 17326 11041
rect 17274 10999 17326 11007
rect 17766 11041 17818 11051
rect 17766 11007 17774 11041
rect 17774 11007 17808 11041
rect 17808 11007 17818 11041
rect 17766 10999 17818 11007
rect 17846 11041 17898 11051
rect 17846 11007 17854 11041
rect 17854 11007 17888 11041
rect 17888 11007 17898 11041
rect 17846 10999 17898 11007
rect 17926 11041 17978 11051
rect 17926 11007 17934 11041
rect 17934 11007 17968 11041
rect 17968 11007 17978 11041
rect 17926 10999 17978 11007
rect 18006 11041 18058 11051
rect 18006 11007 18014 11041
rect 18014 11007 18048 11041
rect 18048 11007 18058 11041
rect 18006 10999 18058 11007
rect 18372 11041 18424 11051
rect 18372 11007 18382 11041
rect 18382 11007 18416 11041
rect 18416 11007 18424 11041
rect 18372 10999 18424 11007
rect 18452 11041 18504 11051
rect 18452 11007 18462 11041
rect 18462 11007 18496 11041
rect 18496 11007 18504 11041
rect 18452 10999 18504 11007
rect 18532 11041 18584 11051
rect 18532 11007 18542 11041
rect 18542 11007 18576 11041
rect 18576 11007 18584 11041
rect 18532 10999 18584 11007
rect 18612 11041 18664 11051
rect 18612 11007 18622 11041
rect 18622 11007 18656 11041
rect 18656 11007 18664 11041
rect 18612 10999 18664 11007
rect 20333 12080 20385 12132
rect 26397 12647 26449 12699
rect 21145 12436 21209 12439
rect 21145 12376 21167 12436
rect 21167 12376 21201 12436
rect 21201 12376 21209 12436
rect 21145 12375 21209 12376
rect 21877 12439 21941 12442
rect 21877 12379 21899 12439
rect 21899 12379 21933 12439
rect 21933 12379 21941 12439
rect 21877 12378 21941 12379
rect 22105 12439 22169 12442
rect 22105 12379 22113 12439
rect 22113 12379 22147 12439
rect 22147 12379 22169 12439
rect 22105 12378 22169 12379
rect 23089 12439 23153 12442
rect 23089 12379 23111 12439
rect 23111 12379 23145 12439
rect 23145 12379 23153 12439
rect 23089 12378 23153 12379
rect 23317 12439 23381 12442
rect 23317 12379 23325 12439
rect 23325 12379 23359 12439
rect 23359 12379 23381 12439
rect 23317 12378 23381 12379
rect 24301 12439 24365 12442
rect 24301 12379 24323 12439
rect 24323 12379 24357 12439
rect 24357 12379 24365 12439
rect 24301 12378 24365 12379
rect 24529 12439 24593 12442
rect 24529 12379 24537 12439
rect 24537 12379 24571 12439
rect 24571 12379 24593 12439
rect 24529 12378 24593 12379
rect 25513 12439 25577 12442
rect 25513 12379 25535 12439
rect 25535 12379 25569 12439
rect 25569 12379 25577 12439
rect 25513 12378 25577 12379
rect 25741 12439 25805 12442
rect 25741 12379 25749 12439
rect 25749 12379 25783 12439
rect 25783 12379 25805 12439
rect 25741 12378 25805 12379
rect 26485 12386 26494 12438
rect 26494 12386 26528 12438
rect 26528 12386 26537 12438
rect 21501 12238 21565 12240
rect 21501 12178 21520 12238
rect 21520 12178 21554 12238
rect 21554 12178 21565 12238
rect 21501 12176 21565 12178
rect 22233 12238 22297 12240
rect 22233 12178 22252 12238
rect 22252 12178 22286 12238
rect 22286 12178 22297 12238
rect 22233 12176 22297 12178
rect 22451 12238 22515 12240
rect 22451 12178 22462 12238
rect 22462 12178 22496 12238
rect 22496 12178 22515 12238
rect 22451 12176 22515 12178
rect 23445 12238 23509 12240
rect 23445 12178 23464 12238
rect 23464 12178 23498 12238
rect 23498 12178 23509 12238
rect 23445 12176 23509 12178
rect 23663 12238 23727 12240
rect 23663 12178 23674 12238
rect 23674 12178 23708 12238
rect 23708 12178 23727 12238
rect 23663 12176 23727 12178
rect 24783 12238 24847 12240
rect 24783 12178 24802 12238
rect 24802 12178 24836 12238
rect 24836 12178 24847 12238
rect 24783 12176 24847 12178
rect 25001 12238 25065 12240
rect 25001 12178 25012 12238
rect 25012 12178 25046 12238
rect 25046 12178 25065 12238
rect 25001 12176 25065 12178
rect 25735 12238 25799 12240
rect 25735 12178 25746 12238
rect 25746 12178 25780 12238
rect 25780 12178 25799 12238
rect 25735 12176 25799 12178
rect 26485 12183 26494 12235
rect 26494 12183 26528 12235
rect 26528 12183 26537 12235
rect 20821 12080 20873 12132
rect 19685 11921 19737 11973
rect 19106 11041 19158 11051
rect 19106 11007 19116 11041
rect 19116 11007 19150 11041
rect 19150 11007 19158 11041
rect 19106 10999 19158 11007
rect 19186 11041 19238 11051
rect 19186 11007 19196 11041
rect 19196 11007 19230 11041
rect 19230 11007 19238 11041
rect 19186 10999 19238 11007
rect 19266 11041 19318 11051
rect 19266 11007 19276 11041
rect 19276 11007 19310 11041
rect 19310 11007 19318 11041
rect 19266 10999 19318 11007
rect 19346 11041 19398 11051
rect 19346 11007 19356 11041
rect 19356 11007 19390 11041
rect 19390 11007 19398 11041
rect 19346 10999 19398 11007
rect 20651 11028 20660 11048
rect 20660 11028 20694 11048
rect 20694 11028 20703 11048
rect 20651 10996 20703 11028
rect 21193 11041 21245 11051
rect 21193 11007 21201 11041
rect 21201 11007 21235 11041
rect 21235 11007 21245 11041
rect 21193 10999 21245 11007
rect 21273 11041 21325 11051
rect 21273 11007 21281 11041
rect 21281 11007 21315 11041
rect 21315 11007 21325 11041
rect 21273 10999 21325 11007
rect 21353 11041 21405 11051
rect 21353 11007 21361 11041
rect 21361 11007 21395 11041
rect 21395 11007 21405 11041
rect 21353 10999 21405 11007
rect 21433 11041 21485 11051
rect 21433 11007 21441 11041
rect 21441 11007 21475 11041
rect 21475 11007 21485 11041
rect 21433 10999 21485 11007
rect 21925 11041 21977 11051
rect 21925 11007 21933 11041
rect 21933 11007 21967 11041
rect 21967 11007 21977 11041
rect 21925 10999 21977 11007
rect 22005 11041 22057 11051
rect 22005 11007 22013 11041
rect 22013 11007 22047 11041
rect 22047 11007 22057 11041
rect 22005 10999 22057 11007
rect 22085 11041 22137 11051
rect 22085 11007 22093 11041
rect 22093 11007 22127 11041
rect 22127 11007 22137 11041
rect 22085 10999 22137 11007
rect 22165 11041 22217 11051
rect 22165 11007 22173 11041
rect 22173 11007 22207 11041
rect 22207 11007 22217 11041
rect 22165 10999 22217 11007
rect 22531 11041 22583 11051
rect 22531 11007 22541 11041
rect 22541 11007 22575 11041
rect 22575 11007 22583 11041
rect 22531 10999 22583 11007
rect 22611 11041 22663 11051
rect 22611 11007 22621 11041
rect 22621 11007 22655 11041
rect 22655 11007 22663 11041
rect 22611 10999 22663 11007
rect 22691 11041 22743 11051
rect 22691 11007 22701 11041
rect 22701 11007 22735 11041
rect 22735 11007 22743 11041
rect 22691 10999 22743 11007
rect 22771 11041 22823 11051
rect 22771 11007 22781 11041
rect 22781 11007 22815 11041
rect 22815 11007 22823 11041
rect 22771 10999 22823 11007
rect 23137 11041 23189 11051
rect 23137 11007 23145 11041
rect 23145 11007 23179 11041
rect 23179 11007 23189 11041
rect 23137 10999 23189 11007
rect 23217 11041 23269 11051
rect 23217 11007 23225 11041
rect 23225 11007 23259 11041
rect 23259 11007 23269 11041
rect 23217 10999 23269 11007
rect 23297 11041 23349 11051
rect 23297 11007 23305 11041
rect 23305 11007 23339 11041
rect 23339 11007 23349 11041
rect 23297 10999 23349 11007
rect 23377 11041 23429 11051
rect 23377 11007 23385 11041
rect 23385 11007 23419 11041
rect 23419 11007 23429 11041
rect 23377 10999 23429 11007
rect 23743 11041 23795 11051
rect 23743 11007 23753 11041
rect 23753 11007 23787 11041
rect 23787 11007 23795 11041
rect 23743 10999 23795 11007
rect 23823 11041 23875 11051
rect 23823 11007 23833 11041
rect 23833 11007 23867 11041
rect 23867 11007 23875 11041
rect 23823 10999 23875 11007
rect 23903 11041 23955 11051
rect 23903 11007 23913 11041
rect 23913 11007 23947 11041
rect 23947 11007 23955 11041
rect 23903 10999 23955 11007
rect 23983 11041 24035 11051
rect 23983 11007 23993 11041
rect 23993 11007 24027 11041
rect 24027 11007 24035 11041
rect 23983 10999 24035 11007
rect 24475 11041 24527 11051
rect 24475 11007 24483 11041
rect 24483 11007 24517 11041
rect 24517 11007 24527 11041
rect 24475 10999 24527 11007
rect 24555 11041 24607 11051
rect 24555 11007 24563 11041
rect 24563 11007 24597 11041
rect 24597 11007 24607 11041
rect 24555 10999 24607 11007
rect 24635 11041 24687 11051
rect 24635 11007 24643 11041
rect 24643 11007 24677 11041
rect 24677 11007 24687 11041
rect 24635 10999 24687 11007
rect 24715 11041 24767 11051
rect 24715 11007 24723 11041
rect 24723 11007 24757 11041
rect 24757 11007 24767 11041
rect 24715 10999 24767 11007
rect 25081 11041 25133 11051
rect 25081 11007 25091 11041
rect 25091 11007 25125 11041
rect 25125 11007 25133 11041
rect 25081 10999 25133 11007
rect 25161 11041 25213 11051
rect 25161 11007 25171 11041
rect 25171 11007 25205 11041
rect 25205 11007 25213 11041
rect 25161 10999 25213 11007
rect 25241 11041 25293 11051
rect 25241 11007 25251 11041
rect 25251 11007 25285 11041
rect 25285 11007 25293 11041
rect 25241 10999 25293 11007
rect 25321 11041 25373 11051
rect 25321 11007 25331 11041
rect 25331 11007 25365 11041
rect 25365 11007 25373 11041
rect 25321 10999 25373 11007
rect 26394 11921 26446 11973
rect 25815 11041 25867 11051
rect 25815 11007 25825 11041
rect 25825 11007 25859 11041
rect 25859 11007 25867 11041
rect 25815 10999 25867 11007
rect 25895 11041 25947 11051
rect 25895 11007 25905 11041
rect 25905 11007 25939 11041
rect 25939 11007 25947 11041
rect 25895 10999 25947 11007
rect 25975 11041 26027 11051
rect 25975 11007 25985 11041
rect 25985 11007 26019 11041
rect 26019 11007 26027 11041
rect 25975 10999 26027 11007
rect 26055 11041 26107 11051
rect 26055 11007 26065 11041
rect 26065 11007 26099 11041
rect 26099 11007 26107 11041
rect 26055 10999 26107 11007
rect 8218 10566 8270 10576
rect 8218 10532 8228 10566
rect 8228 10532 8262 10566
rect 8262 10532 8270 10566
rect 8218 10524 8270 10532
rect 8298 10566 8350 10576
rect 8298 10532 8308 10566
rect 8308 10532 8342 10566
rect 8342 10532 8350 10566
rect 8298 10524 8350 10532
rect 8378 10566 8430 10576
rect 8378 10532 8388 10566
rect 8388 10532 8422 10566
rect 8422 10532 8430 10566
rect 8378 10524 8430 10532
rect 8458 10566 8510 10576
rect 8458 10532 8468 10566
rect 8468 10532 8502 10566
rect 8502 10532 8510 10566
rect 8458 10524 8510 10532
rect 14112 10526 14164 10578
rect 19012 10516 19065 10568
rect 20821 10518 20873 10571
rect 25716 10515 25780 10579
rect 3054 10093 3106 10125
rect 3054 10073 3063 10093
rect 3063 10073 3097 10093
rect 3097 10073 3106 10093
rect 3596 10114 3648 10122
rect 3596 10080 3604 10114
rect 3604 10080 3638 10114
rect 3638 10080 3648 10114
rect 3596 10070 3648 10080
rect 3676 10114 3728 10122
rect 3676 10080 3684 10114
rect 3684 10080 3718 10114
rect 3718 10080 3728 10114
rect 3676 10070 3728 10080
rect 3756 10114 3808 10122
rect 3756 10080 3764 10114
rect 3764 10080 3798 10114
rect 3798 10080 3808 10114
rect 3756 10070 3808 10080
rect 3836 10114 3888 10122
rect 3836 10080 3844 10114
rect 3844 10080 3878 10114
rect 3878 10080 3888 10114
rect 3836 10070 3888 10080
rect 4328 10114 4380 10122
rect 4328 10080 4336 10114
rect 4336 10080 4370 10114
rect 4370 10080 4380 10114
rect 4328 10070 4380 10080
rect 4408 10114 4460 10122
rect 4408 10080 4416 10114
rect 4416 10080 4450 10114
rect 4450 10080 4460 10114
rect 4408 10070 4460 10080
rect 4488 10114 4540 10122
rect 4488 10080 4496 10114
rect 4496 10080 4530 10114
rect 4530 10080 4540 10114
rect 4488 10070 4540 10080
rect 4568 10114 4620 10122
rect 4568 10080 4576 10114
rect 4576 10080 4610 10114
rect 4610 10080 4620 10114
rect 4568 10070 4620 10080
rect 2736 8989 2788 9041
rect 2469 8689 2521 8698
rect 2589 8689 2641 8698
rect 2732 8689 2784 8698
rect 2469 8655 2507 8689
rect 2507 8655 2521 8689
rect 2589 8655 2599 8689
rect 2599 8655 2633 8689
rect 2633 8655 2641 8689
rect 2732 8655 2783 8689
rect 2783 8655 2784 8689
rect 2469 8646 2521 8655
rect 2589 8646 2641 8655
rect 2732 8646 2784 8655
rect 2724 8454 2776 8463
rect 2724 8420 2736 8454
rect 2736 8420 2770 8454
rect 2770 8420 2776 8454
rect 2724 8411 2776 8420
rect 3224 8989 3276 9041
rect 4934 10114 4986 10122
rect 4934 10080 4944 10114
rect 4944 10080 4978 10114
rect 4978 10080 4986 10114
rect 4934 10070 4986 10080
rect 5014 10114 5066 10122
rect 5014 10080 5024 10114
rect 5024 10080 5058 10114
rect 5058 10080 5066 10114
rect 5014 10070 5066 10080
rect 5094 10114 5146 10122
rect 5094 10080 5104 10114
rect 5104 10080 5138 10114
rect 5138 10080 5146 10114
rect 5094 10070 5146 10080
rect 5174 10114 5226 10122
rect 5174 10080 5184 10114
rect 5184 10080 5218 10114
rect 5218 10080 5226 10114
rect 5174 10070 5226 10080
rect 5540 10114 5592 10122
rect 5540 10080 5548 10114
rect 5548 10080 5582 10114
rect 5582 10080 5592 10114
rect 5540 10070 5592 10080
rect 5620 10114 5672 10122
rect 5620 10080 5628 10114
rect 5628 10080 5662 10114
rect 5662 10080 5672 10114
rect 5620 10070 5672 10080
rect 5700 10114 5752 10122
rect 5700 10080 5708 10114
rect 5708 10080 5742 10114
rect 5742 10080 5752 10114
rect 5700 10070 5752 10080
rect 5780 10114 5832 10122
rect 5780 10080 5788 10114
rect 5788 10080 5822 10114
rect 5822 10080 5832 10114
rect 5780 10070 5832 10080
rect 6146 10114 6198 10122
rect 6146 10080 6156 10114
rect 6156 10080 6190 10114
rect 6190 10080 6198 10114
rect 6146 10070 6198 10080
rect 6226 10114 6278 10122
rect 6226 10080 6236 10114
rect 6236 10080 6270 10114
rect 6270 10080 6278 10114
rect 6226 10070 6278 10080
rect 6306 10114 6358 10122
rect 6306 10080 6316 10114
rect 6316 10080 6350 10114
rect 6350 10080 6358 10114
rect 6306 10070 6358 10080
rect 6386 10114 6438 10122
rect 6386 10080 6396 10114
rect 6396 10080 6430 10114
rect 6430 10080 6438 10114
rect 6386 10070 6438 10080
rect 6878 10114 6930 10122
rect 6878 10080 6886 10114
rect 6886 10080 6920 10114
rect 6920 10080 6930 10114
rect 6878 10070 6930 10080
rect 6958 10114 7010 10122
rect 6958 10080 6966 10114
rect 6966 10080 7000 10114
rect 7000 10080 7010 10114
rect 6958 10070 7010 10080
rect 7038 10114 7090 10122
rect 7038 10080 7046 10114
rect 7046 10080 7080 10114
rect 7080 10080 7090 10114
rect 7038 10070 7090 10080
rect 7118 10114 7170 10122
rect 7118 10080 7126 10114
rect 7126 10080 7160 10114
rect 7160 10080 7170 10114
rect 7118 10070 7170 10080
rect 7484 10114 7536 10122
rect 7484 10080 7494 10114
rect 7494 10080 7528 10114
rect 7528 10080 7536 10114
rect 7484 10070 7536 10080
rect 7564 10114 7616 10122
rect 7564 10080 7574 10114
rect 7574 10080 7608 10114
rect 7608 10080 7616 10114
rect 7564 10070 7616 10080
rect 7644 10114 7696 10122
rect 7644 10080 7654 10114
rect 7654 10080 7688 10114
rect 7688 10080 7696 10114
rect 7644 10070 7696 10080
rect 7724 10114 7776 10122
rect 7724 10080 7734 10114
rect 7734 10080 7768 10114
rect 7768 10080 7776 10114
rect 7724 10070 7776 10080
rect 8218 10114 8270 10122
rect 8218 10080 8228 10114
rect 8228 10080 8262 10114
rect 8262 10080 8270 10114
rect 8218 10070 8270 10080
rect 8298 10114 8350 10122
rect 8298 10080 8308 10114
rect 8308 10080 8342 10114
rect 8342 10080 8350 10114
rect 8298 10070 8350 10080
rect 8378 10114 8430 10122
rect 8378 10080 8388 10114
rect 8388 10080 8422 10114
rect 8422 10080 8430 10114
rect 8378 10070 8430 10080
rect 8458 10114 8510 10122
rect 8458 10080 8468 10114
rect 8468 10080 8502 10114
rect 8502 10080 8510 10114
rect 8458 10070 8510 10080
rect 13781 10102 13833 10110
rect 13781 10068 13789 10102
rect 13789 10068 13823 10102
rect 13823 10068 13833 10102
rect 13781 10058 13833 10068
rect 13861 10102 13913 10110
rect 13861 10068 13869 10102
rect 13869 10068 13903 10102
rect 13903 10068 13913 10102
rect 13861 10058 13913 10068
rect 13941 10102 13993 10110
rect 13941 10068 13949 10102
rect 13949 10068 13983 10102
rect 13983 10068 13993 10102
rect 13941 10058 13993 10068
rect 14021 10102 14073 10110
rect 14021 10068 14029 10102
rect 14029 10068 14063 10102
rect 14063 10068 14073 10102
rect 14021 10058 14073 10068
rect 12677 9976 12729 10028
rect 13205 9978 13257 10030
rect 8797 9148 8849 9200
rect 9225 9107 9277 9159
rect 9702 9107 9754 9159
rect 10122 9096 10174 9148
rect 10498 9104 10550 9156
rect 10846 9104 10898 9156
rect 11104 9110 11156 9162
rect 11330 9110 11382 9162
rect 11589 9113 11641 9165
rect 12196 9075 12248 9127
rect 12428 9076 12480 9128
rect 12864 9082 12916 9134
rect 13099 9084 13151 9136
rect 13442 9136 13494 9188
rect 3904 8943 3968 8945
rect 3904 8883 3923 8943
rect 3923 8883 3957 8943
rect 3957 8883 3968 8943
rect 3904 8881 3968 8883
rect 4636 8943 4700 8945
rect 4636 8883 4655 8943
rect 4655 8883 4689 8943
rect 4689 8883 4700 8943
rect 4636 8881 4700 8883
rect 4854 8943 4918 8945
rect 4854 8883 4865 8943
rect 4865 8883 4899 8943
rect 4899 8883 4918 8943
rect 4854 8881 4918 8883
rect 5848 8943 5912 8945
rect 5848 8883 5867 8943
rect 5867 8883 5901 8943
rect 5901 8883 5912 8943
rect 5848 8881 5912 8883
rect 6066 8943 6130 8945
rect 6066 8883 6077 8943
rect 6077 8883 6111 8943
rect 6111 8883 6130 8943
rect 6066 8881 6130 8883
rect 7186 8943 7250 8945
rect 7186 8883 7205 8943
rect 7205 8883 7239 8943
rect 7239 8883 7250 8943
rect 7186 8881 7250 8883
rect 7404 8943 7468 8945
rect 7404 8883 7415 8943
rect 7415 8883 7449 8943
rect 7449 8883 7468 8943
rect 7404 8881 7468 8883
rect 8138 8943 8202 8945
rect 8138 8883 8149 8943
rect 8149 8883 8183 8943
rect 8183 8883 8202 8943
rect 8138 8881 8202 8883
rect 8888 8886 8897 8938
rect 8897 8886 8931 8938
rect 8931 8886 8940 8938
rect 2984 8383 3036 8392
rect 2984 8349 3006 8383
rect 3006 8349 3036 8383
rect 2984 8340 3036 8349
rect 3548 8745 3612 8746
rect 3548 8685 3570 8745
rect 3570 8685 3604 8745
rect 3604 8685 3612 8745
rect 3548 8682 3612 8685
rect 4280 8742 4344 8743
rect 4280 8682 4302 8742
rect 4302 8682 4336 8742
rect 4336 8682 4344 8742
rect 4280 8679 4344 8682
rect 4508 8742 4572 8743
rect 4508 8682 4516 8742
rect 4516 8682 4550 8742
rect 4550 8682 4572 8742
rect 4508 8679 4572 8682
rect 5492 8742 5556 8743
rect 5492 8682 5514 8742
rect 5514 8682 5548 8742
rect 5548 8682 5556 8742
rect 5492 8679 5556 8682
rect 5720 8742 5784 8743
rect 5720 8682 5728 8742
rect 5728 8682 5762 8742
rect 5762 8682 5784 8742
rect 5720 8679 5784 8682
rect 6704 8742 6768 8743
rect 6704 8682 6726 8742
rect 6726 8682 6760 8742
rect 6760 8682 6768 8742
rect 6704 8679 6768 8682
rect 6932 8742 6996 8743
rect 6932 8682 6940 8742
rect 6940 8682 6974 8742
rect 6974 8682 6996 8742
rect 6932 8679 6996 8682
rect 7916 8742 7980 8743
rect 7916 8682 7938 8742
rect 7938 8682 7972 8742
rect 7972 8682 7980 8742
rect 7916 8679 7980 8682
rect 10303 8859 10357 8913
rect 8144 8742 8208 8743
rect 8144 8682 8152 8742
rect 8152 8682 8186 8742
rect 8186 8682 8208 8742
rect 8144 8679 8208 8682
rect 8888 8683 8897 8735
rect 8897 8683 8931 8735
rect 8931 8683 8940 8735
rect 11544 8728 11596 8780
rect 14515 10102 14567 10110
rect 14515 10068 14523 10102
rect 14523 10068 14557 10102
rect 14557 10068 14567 10102
rect 14515 10058 14567 10068
rect 14595 10102 14647 10110
rect 14595 10068 14603 10102
rect 14603 10068 14637 10102
rect 14637 10068 14647 10102
rect 14595 10058 14647 10068
rect 14675 10102 14727 10110
rect 14675 10068 14683 10102
rect 14683 10068 14717 10102
rect 14717 10068 14727 10102
rect 14675 10058 14727 10068
rect 14755 10102 14807 10110
rect 14755 10068 14763 10102
rect 14763 10068 14797 10102
rect 14797 10068 14807 10102
rect 14755 10058 14807 10068
rect 15121 10102 15173 10110
rect 15121 10068 15131 10102
rect 15131 10068 15165 10102
rect 15165 10068 15173 10102
rect 15121 10058 15173 10068
rect 15201 10102 15253 10110
rect 15201 10068 15211 10102
rect 15211 10068 15245 10102
rect 15245 10068 15253 10102
rect 15201 10058 15253 10068
rect 15281 10102 15333 10110
rect 15281 10068 15291 10102
rect 15291 10068 15325 10102
rect 15325 10068 15333 10102
rect 15281 10058 15333 10068
rect 15361 10102 15413 10110
rect 15361 10068 15371 10102
rect 15371 10068 15405 10102
rect 15405 10068 15413 10102
rect 15361 10058 15413 10068
rect 15853 10102 15905 10110
rect 15853 10068 15861 10102
rect 15861 10068 15895 10102
rect 15895 10068 15905 10102
rect 15853 10058 15905 10068
rect 15933 10102 15985 10110
rect 15933 10068 15941 10102
rect 15941 10068 15975 10102
rect 15975 10068 15985 10102
rect 15933 10058 15985 10068
rect 16013 10102 16065 10110
rect 16013 10068 16021 10102
rect 16021 10068 16055 10102
rect 16055 10068 16065 10102
rect 16013 10058 16065 10068
rect 16093 10102 16145 10110
rect 16093 10068 16101 10102
rect 16101 10068 16135 10102
rect 16135 10068 16145 10102
rect 16093 10058 16145 10068
rect 16459 10102 16511 10110
rect 16459 10068 16469 10102
rect 16469 10068 16503 10102
rect 16503 10068 16511 10102
rect 16459 10058 16511 10068
rect 16539 10102 16591 10110
rect 16539 10068 16549 10102
rect 16549 10068 16583 10102
rect 16583 10068 16591 10102
rect 16539 10058 16591 10068
rect 16619 10102 16671 10110
rect 16619 10068 16629 10102
rect 16629 10068 16663 10102
rect 16663 10068 16671 10102
rect 16619 10058 16671 10068
rect 16699 10102 16751 10110
rect 16699 10068 16709 10102
rect 16709 10068 16743 10102
rect 16743 10068 16751 10102
rect 16699 10058 16751 10068
rect 17065 10102 17117 10110
rect 17065 10068 17073 10102
rect 17073 10068 17107 10102
rect 17107 10068 17117 10102
rect 17065 10058 17117 10068
rect 17145 10102 17197 10110
rect 17145 10068 17153 10102
rect 17153 10068 17187 10102
rect 17187 10068 17197 10102
rect 17145 10058 17197 10068
rect 17225 10102 17277 10110
rect 17225 10068 17233 10102
rect 17233 10068 17267 10102
rect 17267 10068 17277 10102
rect 17225 10058 17277 10068
rect 17305 10102 17357 10110
rect 17305 10068 17313 10102
rect 17313 10068 17347 10102
rect 17347 10068 17357 10102
rect 17305 10058 17357 10068
rect 17671 10102 17723 10110
rect 17671 10068 17681 10102
rect 17681 10068 17715 10102
rect 17715 10068 17723 10102
rect 17671 10058 17723 10068
rect 17751 10102 17803 10110
rect 17751 10068 17761 10102
rect 17761 10068 17795 10102
rect 17795 10068 17803 10102
rect 17751 10058 17803 10068
rect 17831 10102 17883 10110
rect 17831 10068 17841 10102
rect 17841 10068 17875 10102
rect 17875 10068 17883 10102
rect 17831 10058 17883 10068
rect 17911 10102 17963 10110
rect 17911 10068 17921 10102
rect 17921 10068 17955 10102
rect 17955 10068 17963 10102
rect 17911 10058 17963 10068
rect 18403 10102 18455 10110
rect 18403 10068 18413 10102
rect 18413 10068 18447 10102
rect 18447 10068 18455 10102
rect 18403 10058 18455 10068
rect 18483 10102 18535 10110
rect 18483 10068 18493 10102
rect 18493 10068 18527 10102
rect 18527 10068 18535 10102
rect 18483 10058 18535 10068
rect 18563 10102 18615 10110
rect 18563 10068 18573 10102
rect 18573 10068 18607 10102
rect 18607 10068 18615 10102
rect 18563 10058 18615 10068
rect 18643 10102 18695 10110
rect 18643 10068 18653 10102
rect 18653 10068 18687 10102
rect 18687 10068 18695 10102
rect 18643 10058 18695 10068
rect 19185 10081 19237 10113
rect 19185 10061 19194 10081
rect 19194 10061 19228 10081
rect 19228 10061 19237 10081
rect 20490 10102 20542 10110
rect 20490 10068 20498 10102
rect 20498 10068 20532 10102
rect 20532 10068 20542 10102
rect 20490 10058 20542 10068
rect 20570 10102 20622 10110
rect 20570 10068 20578 10102
rect 20578 10068 20612 10102
rect 20612 10068 20622 10102
rect 20570 10058 20622 10068
rect 20650 10102 20702 10110
rect 20650 10068 20658 10102
rect 20658 10068 20692 10102
rect 20692 10068 20702 10102
rect 20650 10058 20702 10068
rect 20730 10102 20782 10110
rect 20730 10068 20738 10102
rect 20738 10068 20772 10102
rect 20772 10068 20782 10102
rect 20730 10058 20782 10068
rect 20151 9136 20203 9188
rect 19015 8977 19067 9029
rect 13351 8874 13360 8926
rect 13360 8874 13394 8926
rect 13394 8874 13403 8926
rect 14089 8931 14153 8933
rect 14089 8871 14108 8931
rect 14108 8871 14142 8931
rect 14142 8871 14153 8931
rect 14089 8869 14153 8871
rect 9333 8635 9385 8654
rect 9333 8601 9343 8635
rect 9343 8601 9377 8635
rect 9377 8601 9385 8635
rect 8800 8422 8852 8474
rect 12585 8781 12637 8834
rect 12677 8816 12729 8824
rect 12677 8782 12687 8816
rect 12687 8782 12721 8816
rect 12721 8782 12729 8816
rect 12677 8772 12729 8782
rect 14823 8931 14887 8933
rect 14823 8871 14842 8931
rect 14842 8871 14876 8931
rect 14876 8871 14887 8931
rect 14823 8869 14887 8871
rect 15041 8931 15105 8933
rect 15041 8871 15052 8931
rect 15052 8871 15086 8931
rect 15086 8871 15105 8931
rect 15041 8869 15105 8871
rect 16161 8931 16225 8933
rect 16161 8871 16180 8931
rect 16180 8871 16214 8931
rect 16214 8871 16225 8931
rect 16161 8869 16225 8871
rect 16379 8931 16443 8933
rect 16379 8871 16390 8931
rect 16390 8871 16424 8931
rect 16424 8871 16443 8931
rect 16379 8869 16443 8871
rect 17373 8931 17437 8933
rect 17373 8871 17392 8931
rect 17392 8871 17426 8931
rect 17426 8871 17437 8931
rect 17373 8869 17437 8871
rect 17591 8931 17655 8933
rect 17591 8871 17602 8931
rect 17602 8871 17636 8931
rect 17636 8871 17655 8931
rect 17591 8869 17655 8871
rect 18323 8931 18387 8933
rect 18323 8871 18334 8931
rect 18334 8871 18368 8931
rect 18368 8871 18387 8931
rect 18323 8869 18387 8871
rect 12594 8590 12646 8642
rect 12923 8587 12975 8639
rect 13351 8671 13360 8723
rect 13360 8671 13394 8723
rect 13394 8671 13403 8723
rect 14083 8730 14147 8731
rect 14083 8670 14105 8730
rect 14105 8670 14139 8730
rect 14139 8670 14147 8730
rect 14083 8667 14147 8670
rect 14311 8730 14375 8731
rect 14311 8670 14319 8730
rect 14319 8670 14353 8730
rect 14353 8670 14375 8730
rect 14311 8667 14375 8670
rect 15295 8730 15359 8731
rect 15295 8670 15317 8730
rect 15317 8670 15351 8730
rect 15351 8670 15359 8730
rect 15295 8667 15359 8670
rect 15523 8730 15587 8731
rect 15523 8670 15531 8730
rect 15531 8670 15565 8730
rect 15565 8670 15587 8730
rect 15523 8667 15587 8670
rect 16507 8730 16571 8731
rect 16507 8670 16529 8730
rect 16529 8670 16563 8730
rect 16563 8670 16571 8730
rect 16507 8667 16571 8670
rect 16735 8730 16799 8731
rect 16735 8670 16743 8730
rect 16743 8670 16777 8730
rect 16777 8670 16799 8730
rect 16735 8667 16799 8670
rect 17719 8730 17783 8731
rect 17719 8670 17741 8730
rect 17741 8670 17775 8730
rect 17775 8670 17783 8730
rect 17719 8667 17783 8670
rect 17947 8730 18011 8731
rect 17947 8670 17955 8730
rect 17955 8670 17989 8730
rect 17989 8670 18011 8730
rect 17947 8667 18011 8670
rect 18679 8733 18743 8734
rect 18679 8673 18687 8733
rect 18687 8673 18721 8733
rect 18721 8673 18743 8733
rect 18679 8670 18743 8673
rect 12723 8477 12770 8509
rect 12770 8477 12776 8509
rect 13097 8477 13138 8509
rect 13138 8477 13150 8509
rect 9210 8396 9262 8448
rect 9472 8397 9524 8449
rect 9744 8397 9796 8449
rect 10071 8397 10123 8449
rect 10452 8397 10504 8449
rect 10829 8397 10881 8449
rect 12723 8456 12776 8477
rect 13097 8456 13150 8477
rect 12228 8427 12281 8439
rect 2451 8100 2503 8152
rect 2582 8145 2634 8153
rect 2582 8111 2599 8145
rect 2599 8111 2633 8145
rect 2633 8111 2634 8145
rect 2582 8101 2634 8111
rect 2726 8100 2778 8152
rect 8882 8221 8934 8232
rect 8882 8187 8893 8221
rect 8893 8187 8927 8221
rect 8927 8187 8934 8221
rect 8882 8180 8934 8187
rect 8883 8064 8935 8075
rect 8883 8030 8894 8064
rect 8894 8030 8928 8064
rect 8928 8030 8935 8064
rect 8883 8023 8935 8030
rect 10706 8112 10758 8121
rect 10706 8078 10715 8112
rect 10715 8078 10749 8112
rect 10749 8078 10758 8112
rect 10706 8069 10758 8078
rect 11524 8112 11576 8122
rect 11524 8078 11538 8112
rect 11538 8078 11572 8112
rect 11572 8078 11576 8112
rect 11524 8070 11576 8078
rect 12228 8393 12234 8427
rect 12234 8393 12274 8427
rect 12274 8393 12281 8427
rect 12228 8386 12281 8393
rect 13439 8410 13491 8462
rect 9340 7996 9392 8049
rect 12585 8313 12638 8366
rect 12769 8310 12822 8363
rect 13071 8304 13124 8357
rect 19503 8977 19555 9029
rect 21224 10102 21276 10110
rect 21224 10068 21232 10102
rect 21232 10068 21266 10102
rect 21266 10068 21276 10102
rect 21224 10058 21276 10068
rect 21304 10102 21356 10110
rect 21304 10068 21312 10102
rect 21312 10068 21346 10102
rect 21346 10068 21356 10102
rect 21304 10058 21356 10068
rect 21384 10102 21436 10110
rect 21384 10068 21392 10102
rect 21392 10068 21426 10102
rect 21426 10068 21436 10102
rect 21384 10058 21436 10068
rect 21464 10102 21516 10110
rect 21464 10068 21472 10102
rect 21472 10068 21506 10102
rect 21506 10068 21516 10102
rect 21464 10058 21516 10068
rect 21830 10102 21882 10110
rect 21830 10068 21840 10102
rect 21840 10068 21874 10102
rect 21874 10068 21882 10102
rect 21830 10058 21882 10068
rect 21910 10102 21962 10110
rect 21910 10068 21920 10102
rect 21920 10068 21954 10102
rect 21954 10068 21962 10102
rect 21910 10058 21962 10068
rect 21990 10102 22042 10110
rect 21990 10068 22000 10102
rect 22000 10068 22034 10102
rect 22034 10068 22042 10102
rect 21990 10058 22042 10068
rect 22070 10102 22122 10110
rect 22070 10068 22080 10102
rect 22080 10068 22114 10102
rect 22114 10068 22122 10102
rect 22070 10058 22122 10068
rect 22562 10102 22614 10110
rect 22562 10068 22570 10102
rect 22570 10068 22604 10102
rect 22604 10068 22614 10102
rect 22562 10058 22614 10068
rect 22642 10102 22694 10110
rect 22642 10068 22650 10102
rect 22650 10068 22684 10102
rect 22684 10068 22694 10102
rect 22642 10058 22694 10068
rect 22722 10102 22774 10110
rect 22722 10068 22730 10102
rect 22730 10068 22764 10102
rect 22764 10068 22774 10102
rect 22722 10058 22774 10068
rect 22802 10102 22854 10110
rect 22802 10068 22810 10102
rect 22810 10068 22844 10102
rect 22844 10068 22854 10102
rect 22802 10058 22854 10068
rect 23168 10102 23220 10110
rect 23168 10068 23178 10102
rect 23178 10068 23212 10102
rect 23212 10068 23220 10102
rect 23168 10058 23220 10068
rect 23248 10102 23300 10110
rect 23248 10068 23258 10102
rect 23258 10068 23292 10102
rect 23292 10068 23300 10102
rect 23248 10058 23300 10068
rect 23328 10102 23380 10110
rect 23328 10068 23338 10102
rect 23338 10068 23372 10102
rect 23372 10068 23380 10102
rect 23328 10058 23380 10068
rect 23408 10102 23460 10110
rect 23408 10068 23418 10102
rect 23418 10068 23452 10102
rect 23452 10068 23460 10102
rect 23408 10058 23460 10068
rect 23774 10102 23826 10110
rect 23774 10068 23782 10102
rect 23782 10068 23816 10102
rect 23816 10068 23826 10102
rect 23774 10058 23826 10068
rect 23854 10102 23906 10110
rect 23854 10068 23862 10102
rect 23862 10068 23896 10102
rect 23896 10068 23906 10102
rect 23854 10058 23906 10068
rect 23934 10102 23986 10110
rect 23934 10068 23942 10102
rect 23942 10068 23976 10102
rect 23976 10068 23986 10102
rect 23934 10058 23986 10068
rect 24014 10102 24066 10110
rect 24014 10068 24022 10102
rect 24022 10068 24056 10102
rect 24056 10068 24066 10102
rect 24014 10058 24066 10068
rect 24380 10102 24432 10110
rect 24380 10068 24390 10102
rect 24390 10068 24424 10102
rect 24424 10068 24432 10102
rect 24380 10058 24432 10068
rect 24460 10102 24512 10110
rect 24460 10068 24470 10102
rect 24470 10068 24504 10102
rect 24504 10068 24512 10102
rect 24460 10058 24512 10068
rect 24540 10102 24592 10110
rect 24540 10068 24550 10102
rect 24550 10068 24584 10102
rect 24584 10068 24592 10102
rect 24540 10058 24592 10068
rect 24620 10102 24672 10110
rect 24620 10068 24630 10102
rect 24630 10068 24664 10102
rect 24664 10068 24672 10102
rect 24620 10058 24672 10068
rect 25112 10102 25164 10110
rect 25112 10068 25122 10102
rect 25122 10068 25156 10102
rect 25156 10068 25164 10102
rect 25112 10058 25164 10068
rect 25192 10102 25244 10110
rect 25192 10068 25202 10102
rect 25202 10068 25236 10102
rect 25236 10068 25244 10102
rect 25192 10058 25244 10068
rect 25272 10102 25324 10110
rect 25272 10068 25282 10102
rect 25282 10068 25316 10102
rect 25316 10068 25324 10102
rect 25272 10058 25324 10068
rect 25352 10102 25404 10110
rect 25352 10068 25362 10102
rect 25362 10068 25396 10102
rect 25396 10068 25404 10102
rect 25352 10058 25404 10068
rect 25894 10081 25946 10113
rect 25894 10061 25903 10081
rect 25903 10061 25937 10081
rect 25937 10061 25946 10081
rect 25724 8977 25776 9029
rect 20060 8874 20069 8926
rect 20069 8874 20103 8926
rect 20103 8874 20112 8926
rect 20798 8931 20862 8933
rect 20798 8871 20817 8931
rect 20817 8871 20851 8931
rect 20851 8871 20862 8931
rect 20798 8869 20862 8871
rect 21532 8931 21596 8933
rect 21532 8871 21551 8931
rect 21551 8871 21585 8931
rect 21585 8871 21596 8931
rect 21532 8869 21596 8871
rect 21750 8931 21814 8933
rect 21750 8871 21761 8931
rect 21761 8871 21795 8931
rect 21795 8871 21814 8931
rect 21750 8869 21814 8871
rect 22870 8931 22934 8933
rect 22870 8871 22889 8931
rect 22889 8871 22923 8931
rect 22923 8871 22934 8931
rect 22870 8869 22934 8871
rect 23088 8931 23152 8933
rect 23088 8871 23099 8931
rect 23099 8871 23133 8931
rect 23133 8871 23152 8931
rect 23088 8869 23152 8871
rect 24082 8931 24146 8933
rect 24082 8871 24101 8931
rect 24101 8871 24135 8931
rect 24135 8871 24146 8931
rect 24082 8869 24146 8871
rect 24300 8931 24364 8933
rect 24300 8871 24311 8931
rect 24311 8871 24345 8931
rect 24345 8871 24364 8931
rect 24300 8869 24364 8871
rect 25032 8931 25096 8933
rect 25032 8871 25043 8931
rect 25043 8871 25077 8931
rect 25077 8871 25096 8931
rect 25032 8869 25096 8871
rect 19507 8677 19559 8686
rect 19650 8677 19702 8686
rect 19770 8677 19822 8686
rect 19507 8643 19508 8677
rect 19508 8643 19559 8677
rect 19650 8643 19658 8677
rect 19658 8643 19692 8677
rect 19692 8643 19702 8677
rect 19770 8643 19784 8677
rect 19784 8643 19822 8677
rect 19507 8634 19559 8643
rect 19650 8634 19702 8643
rect 19770 8634 19822 8643
rect 20060 8671 20069 8723
rect 20069 8671 20103 8723
rect 20103 8671 20112 8723
rect 20792 8730 20856 8731
rect 20792 8670 20814 8730
rect 20814 8670 20848 8730
rect 20848 8670 20856 8730
rect 20792 8667 20856 8670
rect 21020 8730 21084 8731
rect 21020 8670 21028 8730
rect 21028 8670 21062 8730
rect 21062 8670 21084 8730
rect 21020 8667 21084 8670
rect 22004 8730 22068 8731
rect 22004 8670 22026 8730
rect 22026 8670 22060 8730
rect 22060 8670 22068 8730
rect 22004 8667 22068 8670
rect 22232 8730 22296 8731
rect 22232 8670 22240 8730
rect 22240 8670 22274 8730
rect 22274 8670 22296 8730
rect 22232 8667 22296 8670
rect 23216 8730 23280 8731
rect 23216 8670 23238 8730
rect 23238 8670 23272 8730
rect 23272 8670 23280 8730
rect 23216 8667 23280 8670
rect 23444 8730 23508 8731
rect 23444 8670 23452 8730
rect 23452 8670 23486 8730
rect 23486 8670 23508 8730
rect 23444 8667 23508 8670
rect 24428 8730 24492 8731
rect 24428 8670 24450 8730
rect 24450 8670 24484 8730
rect 24484 8670 24492 8730
rect 24428 8667 24492 8670
rect 24656 8730 24720 8731
rect 24656 8670 24664 8730
rect 24664 8670 24698 8730
rect 24698 8670 24720 8730
rect 24656 8667 24720 8670
rect 25388 8733 25452 8734
rect 25388 8673 25396 8733
rect 25396 8673 25430 8733
rect 25430 8673 25452 8733
rect 25388 8670 25452 8673
rect 13357 8209 13409 8220
rect 13357 8175 13364 8209
rect 13364 8175 13398 8209
rect 13398 8175 13409 8209
rect 13357 8168 13409 8175
rect 19515 8442 19567 8451
rect 19515 8408 19521 8442
rect 19521 8408 19555 8442
rect 19555 8408 19567 8442
rect 19515 8399 19567 8408
rect 20148 8410 20200 8462
rect 26212 8977 26264 9029
rect 26216 8677 26268 8686
rect 26359 8677 26411 8686
rect 26479 8677 26531 8686
rect 26216 8643 26217 8677
rect 26217 8643 26268 8677
rect 26359 8643 26367 8677
rect 26367 8643 26401 8677
rect 26401 8643 26411 8677
rect 26479 8643 26493 8677
rect 26493 8643 26531 8677
rect 26216 8634 26268 8643
rect 26359 8634 26411 8643
rect 26479 8634 26531 8643
rect 8883 7894 8935 7905
rect 8883 7860 8894 7894
rect 8894 7860 8928 7894
rect 8928 7860 8935 7894
rect 8883 7853 8935 7860
rect 8882 7742 8934 7753
rect 8882 7708 8893 7742
rect 8893 7708 8927 7742
rect 8927 7708 8934 7742
rect 8882 7701 8934 7708
rect 3166 7550 3218 7556
rect 3068 7495 3120 7547
rect 3166 7516 3176 7550
rect 3176 7516 3210 7550
rect 3210 7516 3218 7550
rect 3166 7504 3218 7516
rect 3246 7550 3298 7556
rect 3246 7516 3256 7550
rect 3256 7516 3290 7550
rect 3290 7516 3298 7550
rect 3246 7504 3298 7516
rect 3326 7550 3378 7556
rect 3326 7516 3336 7550
rect 3336 7516 3370 7550
rect 3370 7516 3378 7550
rect 3326 7504 3378 7516
rect 3406 7550 3458 7556
rect 3406 7516 3416 7550
rect 3416 7516 3450 7550
rect 3450 7516 3458 7550
rect 3406 7504 3458 7516
rect 3486 7550 3538 7556
rect 3486 7516 3496 7550
rect 3496 7516 3530 7550
rect 3530 7516 3538 7550
rect 3486 7504 3538 7516
rect 3566 7550 3618 7556
rect 3566 7516 3576 7550
rect 3576 7516 3610 7550
rect 3610 7516 3618 7550
rect 3566 7504 3618 7516
rect 3898 7547 3950 7553
rect 3898 7513 3908 7547
rect 3908 7513 3942 7547
rect 3942 7513 3950 7547
rect 3898 7501 3950 7513
rect 3978 7547 4030 7553
rect 3978 7513 3988 7547
rect 3988 7513 4022 7547
rect 4022 7513 4030 7547
rect 3978 7501 4030 7513
rect 4058 7547 4110 7553
rect 4058 7513 4068 7547
rect 4068 7513 4102 7547
rect 4102 7513 4110 7547
rect 4058 7501 4110 7513
rect 4138 7547 4190 7553
rect 4138 7513 4148 7547
rect 4148 7513 4182 7547
rect 4182 7513 4190 7547
rect 4138 7501 4190 7513
rect 4218 7547 4270 7553
rect 4218 7513 4228 7547
rect 4228 7513 4262 7547
rect 4262 7513 4270 7547
rect 4218 7501 4270 7513
rect 4298 7547 4350 7553
rect 4298 7513 4308 7547
rect 4308 7513 4342 7547
rect 4342 7513 4350 7547
rect 4298 7501 4350 7513
rect 4502 7547 4554 7553
rect 4502 7513 4510 7547
rect 4510 7513 4544 7547
rect 4544 7513 4554 7547
rect 4502 7501 4554 7513
rect 4582 7547 4634 7553
rect 4582 7513 4590 7547
rect 4590 7513 4624 7547
rect 4624 7513 4634 7547
rect 4582 7501 4634 7513
rect 4662 7547 4714 7553
rect 4662 7513 4670 7547
rect 4670 7513 4704 7547
rect 4704 7513 4714 7547
rect 4662 7501 4714 7513
rect 4742 7547 4794 7553
rect 4742 7513 4750 7547
rect 4750 7513 4784 7547
rect 4784 7513 4794 7547
rect 4742 7501 4794 7513
rect 4822 7547 4874 7553
rect 4822 7513 4830 7547
rect 4830 7513 4864 7547
rect 4864 7513 4874 7547
rect 4822 7501 4874 7513
rect 4902 7547 4954 7553
rect 4902 7513 4910 7547
rect 4910 7513 4944 7547
rect 4944 7513 4954 7547
rect 4902 7501 4954 7513
rect 5110 7547 5162 7553
rect 5110 7513 5120 7547
rect 5120 7513 5154 7547
rect 5154 7513 5162 7547
rect 5110 7501 5162 7513
rect 5190 7547 5242 7553
rect 5190 7513 5200 7547
rect 5200 7513 5234 7547
rect 5234 7513 5242 7547
rect 5190 7501 5242 7513
rect 5270 7547 5322 7553
rect 5270 7513 5280 7547
rect 5280 7513 5314 7547
rect 5314 7513 5322 7547
rect 5270 7501 5322 7513
rect 5350 7547 5402 7553
rect 5350 7513 5360 7547
rect 5360 7513 5394 7547
rect 5394 7513 5402 7547
rect 5350 7501 5402 7513
rect 5430 7547 5482 7553
rect 5430 7513 5440 7547
rect 5440 7513 5474 7547
rect 5474 7513 5482 7547
rect 5430 7501 5482 7513
rect 5510 7547 5562 7553
rect 5510 7513 5520 7547
rect 5520 7513 5554 7547
rect 5554 7513 5562 7547
rect 5510 7501 5562 7513
rect 5714 7547 5766 7553
rect 5714 7513 5722 7547
rect 5722 7513 5756 7547
rect 5756 7513 5766 7547
rect 5714 7501 5766 7513
rect 5794 7547 5846 7553
rect 5794 7513 5802 7547
rect 5802 7513 5836 7547
rect 5836 7513 5846 7547
rect 5794 7501 5846 7513
rect 5874 7547 5926 7553
rect 5874 7513 5882 7547
rect 5882 7513 5916 7547
rect 5916 7513 5926 7547
rect 5874 7501 5926 7513
rect 5954 7547 6006 7553
rect 5954 7513 5962 7547
rect 5962 7513 5996 7547
rect 5996 7513 6006 7547
rect 5954 7501 6006 7513
rect 6034 7547 6086 7553
rect 6034 7513 6042 7547
rect 6042 7513 6076 7547
rect 6076 7513 6086 7547
rect 6034 7501 6086 7513
rect 6114 7547 6166 7553
rect 6114 7513 6122 7547
rect 6122 7513 6156 7547
rect 6156 7513 6166 7547
rect 6114 7501 6166 7513
rect 6322 7547 6374 7553
rect 6322 7513 6332 7547
rect 6332 7513 6366 7547
rect 6366 7513 6374 7547
rect 6322 7501 6374 7513
rect 6402 7547 6454 7553
rect 6402 7513 6412 7547
rect 6412 7513 6446 7547
rect 6446 7513 6454 7547
rect 6402 7501 6454 7513
rect 6482 7547 6534 7553
rect 6482 7513 6492 7547
rect 6492 7513 6526 7547
rect 6526 7513 6534 7547
rect 6482 7501 6534 7513
rect 6562 7547 6614 7553
rect 6562 7513 6572 7547
rect 6572 7513 6606 7547
rect 6606 7513 6614 7547
rect 6562 7501 6614 7513
rect 6642 7547 6694 7553
rect 6642 7513 6652 7547
rect 6652 7513 6686 7547
rect 6686 7513 6694 7547
rect 6642 7501 6694 7513
rect 6722 7547 6774 7553
rect 6722 7513 6732 7547
rect 6732 7513 6766 7547
rect 6766 7513 6774 7547
rect 6722 7501 6774 7513
rect 6926 7547 6978 7553
rect 6926 7513 6934 7547
rect 6934 7513 6968 7547
rect 6968 7513 6978 7547
rect 6926 7501 6978 7513
rect 7006 7547 7058 7553
rect 7006 7513 7014 7547
rect 7014 7513 7048 7547
rect 7048 7513 7058 7547
rect 7006 7501 7058 7513
rect 7086 7547 7138 7553
rect 7086 7513 7094 7547
rect 7094 7513 7128 7547
rect 7128 7513 7138 7547
rect 7086 7501 7138 7513
rect 7166 7547 7218 7553
rect 7166 7513 7174 7547
rect 7174 7513 7208 7547
rect 7208 7513 7218 7547
rect 7166 7501 7218 7513
rect 7246 7547 7298 7553
rect 7246 7513 7254 7547
rect 7254 7513 7288 7547
rect 7288 7513 7298 7547
rect 7246 7501 7298 7513
rect 7326 7547 7378 7553
rect 7326 7513 7334 7547
rect 7334 7513 7368 7547
rect 7368 7513 7378 7547
rect 7326 7501 7378 7513
rect 7534 7547 7586 7553
rect 7534 7513 7544 7547
rect 7544 7513 7578 7547
rect 7578 7513 7586 7547
rect 7534 7501 7586 7513
rect 7614 7547 7666 7553
rect 7614 7513 7624 7547
rect 7624 7513 7658 7547
rect 7658 7513 7666 7547
rect 7614 7501 7666 7513
rect 7694 7547 7746 7553
rect 7694 7513 7704 7547
rect 7704 7513 7738 7547
rect 7738 7513 7746 7547
rect 7694 7501 7746 7513
rect 7774 7547 7826 7553
rect 7774 7513 7784 7547
rect 7784 7513 7818 7547
rect 7818 7513 7826 7547
rect 7774 7501 7826 7513
rect 7854 7547 7906 7553
rect 7854 7513 7864 7547
rect 7864 7513 7898 7547
rect 7898 7513 7906 7547
rect 7854 7501 7906 7513
rect 7934 7547 7986 7553
rect 7934 7513 7944 7547
rect 7944 7513 7978 7547
rect 7978 7513 7986 7547
rect 7934 7501 7986 7513
rect 8138 7547 8190 7553
rect 8138 7513 8146 7547
rect 8146 7513 8180 7547
rect 8180 7513 8190 7547
rect 8138 7501 8190 7513
rect 8218 7547 8270 7553
rect 8218 7513 8226 7547
rect 8226 7513 8260 7547
rect 8260 7513 8270 7547
rect 8218 7501 8270 7513
rect 8298 7547 8350 7553
rect 8298 7513 8306 7547
rect 8306 7513 8340 7547
rect 8340 7513 8350 7547
rect 8298 7501 8350 7513
rect 8378 7547 8430 7553
rect 8378 7513 8386 7547
rect 8386 7513 8420 7547
rect 8420 7513 8430 7547
rect 8378 7501 8430 7513
rect 8458 7547 8510 7553
rect 8458 7513 8466 7547
rect 8466 7513 8500 7547
rect 8500 7513 8510 7547
rect 8458 7501 8510 7513
rect 8538 7547 8590 7553
rect 8538 7513 8546 7547
rect 8546 7513 8580 7547
rect 8580 7513 8590 7547
rect 8538 7501 8590 7513
rect 8877 7598 8929 7609
rect 8877 7564 8888 7598
rect 8888 7564 8922 7598
rect 8922 7564 8929 7598
rect 8877 7557 8929 7564
rect 11750 7797 11802 7849
rect 10146 7671 10198 7723
rect 10394 7671 10446 7723
rect 10691 7671 10743 7723
rect 11035 7673 11087 7725
rect 11354 7673 11406 7725
rect 11966 7728 11976 7734
rect 11976 7728 12014 7734
rect 12014 7728 12018 7734
rect 11966 7690 12018 7728
rect 12220 7727 12232 7738
rect 12232 7727 12266 7738
rect 12266 7727 12272 7738
rect 11966 7682 11975 7690
rect 11975 7682 12013 7690
rect 12013 7682 12018 7690
rect 12220 7689 12272 7727
rect 12220 7686 12231 7689
rect 12231 7686 12265 7689
rect 12265 7686 12272 7689
rect 11976 7584 12013 7589
rect 12013 7584 12028 7589
rect 11976 7546 12028 7584
rect 12228 7583 12231 7592
rect 12231 7583 12265 7592
rect 12265 7583 12280 7592
rect 12919 7987 12971 8040
rect 13356 8052 13408 8063
rect 13356 8018 13363 8052
rect 13363 8018 13397 8052
rect 13397 8018 13408 8052
rect 13356 8011 13408 8018
rect 20066 8209 20118 8220
rect 20066 8175 20073 8209
rect 20073 8175 20107 8209
rect 20107 8175 20118 8209
rect 20066 8168 20118 8175
rect 26224 8442 26276 8451
rect 26224 8408 26230 8442
rect 26230 8408 26264 8442
rect 26264 8408 26276 8442
rect 26224 8399 26276 8408
rect 19513 8088 19565 8140
rect 19657 8133 19709 8141
rect 19657 8099 19658 8133
rect 19658 8099 19692 8133
rect 19692 8099 19709 8133
rect 19657 8089 19709 8099
rect 19788 8088 19840 8140
rect 20065 8052 20117 8063
rect 20065 8018 20072 8052
rect 20072 8018 20106 8052
rect 20106 8018 20117 8052
rect 20065 8011 20117 8018
rect 12940 7918 12992 7929
rect 12940 7884 12947 7918
rect 12947 7884 12981 7918
rect 12981 7884 12992 7918
rect 12940 7877 12992 7884
rect 13356 7882 13408 7893
rect 13356 7848 13363 7882
rect 13363 7848 13397 7882
rect 13397 7848 13408 7882
rect 13356 7841 13408 7848
rect 12932 7698 12984 7709
rect 12932 7664 12939 7698
rect 12939 7664 12973 7698
rect 12973 7664 12984 7698
rect 12932 7657 12984 7664
rect 13357 7730 13409 7741
rect 13357 7696 13364 7730
rect 13364 7696 13398 7730
rect 13398 7696 13409 7730
rect 13357 7689 13409 7696
rect 26222 8088 26274 8140
rect 26366 8133 26418 8141
rect 26366 8099 26367 8133
rect 26367 8099 26401 8133
rect 26401 8099 26418 8133
rect 26366 8089 26418 8099
rect 26497 8088 26549 8140
rect 19643 7980 19695 7991
rect 19643 7946 19650 7980
rect 19650 7946 19684 7980
rect 19684 7946 19695 7980
rect 19643 7939 19695 7946
rect 20065 7882 20117 7893
rect 20065 7848 20072 7882
rect 20072 7848 20106 7882
rect 20106 7848 20117 7882
rect 20065 7841 20117 7848
rect 19643 7784 19695 7795
rect 19643 7750 19650 7784
rect 19650 7750 19684 7784
rect 19684 7750 19695 7784
rect 19643 7743 19695 7750
rect 20066 7730 20118 7741
rect 20066 7696 20073 7730
rect 20073 7696 20107 7730
rect 20107 7696 20118 7730
rect 20066 7689 20118 7696
rect 10311 7481 10363 7533
rect 11749 7480 11801 7532
rect 11976 7537 12012 7546
rect 12012 7537 12028 7546
rect 12228 7545 12280 7583
rect 12228 7540 12230 7545
rect 12230 7540 12264 7545
rect 12264 7540 12280 7545
rect 13362 7586 13414 7597
rect 13362 7552 13369 7586
rect 13369 7552 13403 7586
rect 13403 7552 13414 7586
rect 13362 7545 13414 7552
rect 13701 7535 13753 7541
rect 13701 7501 13711 7535
rect 13711 7501 13745 7535
rect 13745 7501 13753 7535
rect 13701 7489 13753 7501
rect 13781 7535 13833 7541
rect 13781 7501 13791 7535
rect 13791 7501 13825 7535
rect 13825 7501 13833 7535
rect 13781 7489 13833 7501
rect 13861 7535 13913 7541
rect 13861 7501 13871 7535
rect 13871 7501 13905 7535
rect 13905 7501 13913 7535
rect 13861 7489 13913 7501
rect 13941 7535 13993 7541
rect 13941 7501 13951 7535
rect 13951 7501 13985 7535
rect 13985 7501 13993 7535
rect 13941 7489 13993 7501
rect 14021 7535 14073 7541
rect 14021 7501 14031 7535
rect 14031 7501 14065 7535
rect 14065 7501 14073 7535
rect 14021 7489 14073 7501
rect 14101 7535 14153 7541
rect 14101 7501 14111 7535
rect 14111 7501 14145 7535
rect 14145 7501 14153 7535
rect 14101 7489 14153 7501
rect 14305 7535 14357 7541
rect 14305 7501 14313 7535
rect 14313 7501 14347 7535
rect 14347 7501 14357 7535
rect 14305 7489 14357 7501
rect 14385 7535 14437 7541
rect 14385 7501 14393 7535
rect 14393 7501 14427 7535
rect 14427 7501 14437 7535
rect 14385 7489 14437 7501
rect 14465 7535 14517 7541
rect 14465 7501 14473 7535
rect 14473 7501 14507 7535
rect 14507 7501 14517 7535
rect 14465 7489 14517 7501
rect 14545 7535 14597 7541
rect 14545 7501 14553 7535
rect 14553 7501 14587 7535
rect 14587 7501 14597 7535
rect 14545 7489 14597 7501
rect 14625 7535 14677 7541
rect 14625 7501 14633 7535
rect 14633 7501 14667 7535
rect 14667 7501 14677 7535
rect 14625 7489 14677 7501
rect 14705 7535 14757 7541
rect 14705 7501 14713 7535
rect 14713 7501 14747 7535
rect 14747 7501 14757 7535
rect 14705 7489 14757 7501
rect 14913 7535 14965 7541
rect 14913 7501 14923 7535
rect 14923 7501 14957 7535
rect 14957 7501 14965 7535
rect 14913 7489 14965 7501
rect 14993 7535 15045 7541
rect 14993 7501 15003 7535
rect 15003 7501 15037 7535
rect 15037 7501 15045 7535
rect 14993 7489 15045 7501
rect 15073 7535 15125 7541
rect 15073 7501 15083 7535
rect 15083 7501 15117 7535
rect 15117 7501 15125 7535
rect 15073 7489 15125 7501
rect 15153 7535 15205 7541
rect 15153 7501 15163 7535
rect 15163 7501 15197 7535
rect 15197 7501 15205 7535
rect 15153 7489 15205 7501
rect 15233 7535 15285 7541
rect 15233 7501 15243 7535
rect 15243 7501 15277 7535
rect 15277 7501 15285 7535
rect 15233 7489 15285 7501
rect 15313 7535 15365 7541
rect 15313 7501 15323 7535
rect 15323 7501 15357 7535
rect 15357 7501 15365 7535
rect 15313 7489 15365 7501
rect 15517 7535 15569 7541
rect 15517 7501 15525 7535
rect 15525 7501 15559 7535
rect 15559 7501 15569 7535
rect 15517 7489 15569 7501
rect 15597 7535 15649 7541
rect 15597 7501 15605 7535
rect 15605 7501 15639 7535
rect 15639 7501 15649 7535
rect 15597 7489 15649 7501
rect 15677 7535 15729 7541
rect 15677 7501 15685 7535
rect 15685 7501 15719 7535
rect 15719 7501 15729 7535
rect 15677 7489 15729 7501
rect 15757 7535 15809 7541
rect 15757 7501 15765 7535
rect 15765 7501 15799 7535
rect 15799 7501 15809 7535
rect 15757 7489 15809 7501
rect 15837 7535 15889 7541
rect 15837 7501 15845 7535
rect 15845 7501 15879 7535
rect 15879 7501 15889 7535
rect 15837 7489 15889 7501
rect 15917 7535 15969 7541
rect 15917 7501 15925 7535
rect 15925 7501 15959 7535
rect 15959 7501 15969 7535
rect 15917 7489 15969 7501
rect 16125 7535 16177 7541
rect 16125 7501 16135 7535
rect 16135 7501 16169 7535
rect 16169 7501 16177 7535
rect 16125 7489 16177 7501
rect 16205 7535 16257 7541
rect 16205 7501 16215 7535
rect 16215 7501 16249 7535
rect 16249 7501 16257 7535
rect 16205 7489 16257 7501
rect 16285 7535 16337 7541
rect 16285 7501 16295 7535
rect 16295 7501 16329 7535
rect 16329 7501 16337 7535
rect 16285 7489 16337 7501
rect 16365 7535 16417 7541
rect 16365 7501 16375 7535
rect 16375 7501 16409 7535
rect 16409 7501 16417 7535
rect 16365 7489 16417 7501
rect 16445 7535 16497 7541
rect 16445 7501 16455 7535
rect 16455 7501 16489 7535
rect 16489 7501 16497 7535
rect 16445 7489 16497 7501
rect 16525 7535 16577 7541
rect 16525 7501 16535 7535
rect 16535 7501 16569 7535
rect 16569 7501 16577 7535
rect 16525 7489 16577 7501
rect 16729 7535 16781 7541
rect 16729 7501 16737 7535
rect 16737 7501 16771 7535
rect 16771 7501 16781 7535
rect 16729 7489 16781 7501
rect 16809 7535 16861 7541
rect 16809 7501 16817 7535
rect 16817 7501 16851 7535
rect 16851 7501 16861 7535
rect 16809 7489 16861 7501
rect 16889 7535 16941 7541
rect 16889 7501 16897 7535
rect 16897 7501 16931 7535
rect 16931 7501 16941 7535
rect 16889 7489 16941 7501
rect 16969 7535 17021 7541
rect 16969 7501 16977 7535
rect 16977 7501 17011 7535
rect 17011 7501 17021 7535
rect 16969 7489 17021 7501
rect 17049 7535 17101 7541
rect 17049 7501 17057 7535
rect 17057 7501 17091 7535
rect 17091 7501 17101 7535
rect 17049 7489 17101 7501
rect 17129 7535 17181 7541
rect 17129 7501 17137 7535
rect 17137 7501 17171 7535
rect 17171 7501 17181 7535
rect 17129 7489 17181 7501
rect 17337 7535 17389 7541
rect 17337 7501 17347 7535
rect 17347 7501 17381 7535
rect 17381 7501 17389 7535
rect 17337 7489 17389 7501
rect 17417 7535 17469 7541
rect 17417 7501 17427 7535
rect 17427 7501 17461 7535
rect 17461 7501 17469 7535
rect 17417 7489 17469 7501
rect 17497 7535 17549 7541
rect 17497 7501 17507 7535
rect 17507 7501 17541 7535
rect 17541 7501 17549 7535
rect 17497 7489 17549 7501
rect 17577 7535 17629 7541
rect 17577 7501 17587 7535
rect 17587 7501 17621 7535
rect 17621 7501 17629 7535
rect 17577 7489 17629 7501
rect 17657 7535 17709 7541
rect 17657 7501 17667 7535
rect 17667 7501 17701 7535
rect 17701 7501 17709 7535
rect 17657 7489 17709 7501
rect 17737 7535 17789 7541
rect 17737 7501 17747 7535
rect 17747 7501 17781 7535
rect 17781 7501 17789 7535
rect 17737 7489 17789 7501
rect 17941 7535 17993 7541
rect 17941 7501 17949 7535
rect 17949 7501 17983 7535
rect 17983 7501 17993 7535
rect 17941 7489 17993 7501
rect 18021 7535 18073 7541
rect 18021 7501 18029 7535
rect 18029 7501 18063 7535
rect 18063 7501 18073 7535
rect 18021 7489 18073 7501
rect 18101 7535 18153 7541
rect 18101 7501 18109 7535
rect 18109 7501 18143 7535
rect 18143 7501 18153 7535
rect 18101 7489 18153 7501
rect 18181 7535 18233 7541
rect 18181 7501 18189 7535
rect 18189 7501 18223 7535
rect 18223 7501 18233 7535
rect 18181 7489 18233 7501
rect 18261 7535 18313 7541
rect 18261 7501 18269 7535
rect 18269 7501 18303 7535
rect 18303 7501 18313 7535
rect 18261 7489 18313 7501
rect 18341 7535 18393 7541
rect 18341 7501 18349 7535
rect 18349 7501 18383 7535
rect 18383 7501 18393 7535
rect 18341 7489 18393 7501
rect 18673 7538 18725 7544
rect 18673 7504 18681 7538
rect 18681 7504 18715 7538
rect 18715 7504 18725 7538
rect 18673 7492 18725 7504
rect 18753 7538 18805 7544
rect 18753 7504 18761 7538
rect 18761 7504 18795 7538
rect 18795 7504 18805 7538
rect 18753 7492 18805 7504
rect 18833 7538 18885 7544
rect 18833 7504 18841 7538
rect 18841 7504 18875 7538
rect 18875 7504 18885 7538
rect 18833 7492 18885 7504
rect 18913 7538 18965 7544
rect 18913 7504 18921 7538
rect 18921 7504 18955 7538
rect 18955 7504 18965 7538
rect 18913 7492 18965 7504
rect 18993 7538 19045 7544
rect 18993 7504 19001 7538
rect 19001 7504 19035 7538
rect 19035 7504 19045 7538
rect 18993 7492 19045 7504
rect 19073 7538 19125 7544
rect 19073 7504 19081 7538
rect 19081 7504 19115 7538
rect 19115 7504 19125 7538
rect 19073 7492 19125 7504
rect 19171 7483 19223 7535
rect 19643 7609 19695 7620
rect 19643 7575 19650 7609
rect 19650 7575 19684 7609
rect 19684 7575 19695 7609
rect 19643 7568 19695 7575
rect 20071 7586 20123 7597
rect 20071 7552 20078 7586
rect 20078 7552 20112 7586
rect 20112 7552 20123 7586
rect 20071 7545 20123 7552
rect 20410 7535 20462 7541
rect 20410 7501 20420 7535
rect 20420 7501 20454 7535
rect 20454 7501 20462 7535
rect 20410 7489 20462 7501
rect 20490 7535 20542 7541
rect 20490 7501 20500 7535
rect 20500 7501 20534 7535
rect 20534 7501 20542 7535
rect 20490 7489 20542 7501
rect 20570 7535 20622 7541
rect 20570 7501 20580 7535
rect 20580 7501 20614 7535
rect 20614 7501 20622 7535
rect 20570 7489 20622 7501
rect 20650 7535 20702 7541
rect 20650 7501 20660 7535
rect 20660 7501 20694 7535
rect 20694 7501 20702 7535
rect 20650 7489 20702 7501
rect 20730 7535 20782 7541
rect 20730 7501 20740 7535
rect 20740 7501 20774 7535
rect 20774 7501 20782 7535
rect 20730 7489 20782 7501
rect 20810 7535 20862 7541
rect 20810 7501 20820 7535
rect 20820 7501 20854 7535
rect 20854 7501 20862 7535
rect 20810 7489 20862 7501
rect 21014 7535 21066 7541
rect 21014 7501 21022 7535
rect 21022 7501 21056 7535
rect 21056 7501 21066 7535
rect 21014 7489 21066 7501
rect 21094 7535 21146 7541
rect 21094 7501 21102 7535
rect 21102 7501 21136 7535
rect 21136 7501 21146 7535
rect 21094 7489 21146 7501
rect 21174 7535 21226 7541
rect 21174 7501 21182 7535
rect 21182 7501 21216 7535
rect 21216 7501 21226 7535
rect 21174 7489 21226 7501
rect 21254 7535 21306 7541
rect 21254 7501 21262 7535
rect 21262 7501 21296 7535
rect 21296 7501 21306 7535
rect 21254 7489 21306 7501
rect 21334 7535 21386 7541
rect 21334 7501 21342 7535
rect 21342 7501 21376 7535
rect 21376 7501 21386 7535
rect 21334 7489 21386 7501
rect 21414 7535 21466 7541
rect 21414 7501 21422 7535
rect 21422 7501 21456 7535
rect 21456 7501 21466 7535
rect 21414 7489 21466 7501
rect 21622 7535 21674 7541
rect 21622 7501 21632 7535
rect 21632 7501 21666 7535
rect 21666 7501 21674 7535
rect 21622 7489 21674 7501
rect 21702 7535 21754 7541
rect 21702 7501 21712 7535
rect 21712 7501 21746 7535
rect 21746 7501 21754 7535
rect 21702 7489 21754 7501
rect 21782 7535 21834 7541
rect 21782 7501 21792 7535
rect 21792 7501 21826 7535
rect 21826 7501 21834 7535
rect 21782 7489 21834 7501
rect 21862 7535 21914 7541
rect 21862 7501 21872 7535
rect 21872 7501 21906 7535
rect 21906 7501 21914 7535
rect 21862 7489 21914 7501
rect 21942 7535 21994 7541
rect 21942 7501 21952 7535
rect 21952 7501 21986 7535
rect 21986 7501 21994 7535
rect 21942 7489 21994 7501
rect 22022 7535 22074 7541
rect 22022 7501 22032 7535
rect 22032 7501 22066 7535
rect 22066 7501 22074 7535
rect 22022 7489 22074 7501
rect 22226 7535 22278 7541
rect 22226 7501 22234 7535
rect 22234 7501 22268 7535
rect 22268 7501 22278 7535
rect 22226 7489 22278 7501
rect 22306 7535 22358 7541
rect 22306 7501 22314 7535
rect 22314 7501 22348 7535
rect 22348 7501 22358 7535
rect 22306 7489 22358 7501
rect 22386 7535 22438 7541
rect 22386 7501 22394 7535
rect 22394 7501 22428 7535
rect 22428 7501 22438 7535
rect 22386 7489 22438 7501
rect 22466 7535 22518 7541
rect 22466 7501 22474 7535
rect 22474 7501 22508 7535
rect 22508 7501 22518 7535
rect 22466 7489 22518 7501
rect 22546 7535 22598 7541
rect 22546 7501 22554 7535
rect 22554 7501 22588 7535
rect 22588 7501 22598 7535
rect 22546 7489 22598 7501
rect 22626 7535 22678 7541
rect 22626 7501 22634 7535
rect 22634 7501 22668 7535
rect 22668 7501 22678 7535
rect 22626 7489 22678 7501
rect 22834 7535 22886 7541
rect 22834 7501 22844 7535
rect 22844 7501 22878 7535
rect 22878 7501 22886 7535
rect 22834 7489 22886 7501
rect 22914 7535 22966 7541
rect 22914 7501 22924 7535
rect 22924 7501 22958 7535
rect 22958 7501 22966 7535
rect 22914 7489 22966 7501
rect 22994 7535 23046 7541
rect 22994 7501 23004 7535
rect 23004 7501 23038 7535
rect 23038 7501 23046 7535
rect 22994 7489 23046 7501
rect 23074 7535 23126 7541
rect 23074 7501 23084 7535
rect 23084 7501 23118 7535
rect 23118 7501 23126 7535
rect 23074 7489 23126 7501
rect 23154 7535 23206 7541
rect 23154 7501 23164 7535
rect 23164 7501 23198 7535
rect 23198 7501 23206 7535
rect 23154 7489 23206 7501
rect 23234 7535 23286 7541
rect 23234 7501 23244 7535
rect 23244 7501 23278 7535
rect 23278 7501 23286 7535
rect 23234 7489 23286 7501
rect 23438 7535 23490 7541
rect 23438 7501 23446 7535
rect 23446 7501 23480 7535
rect 23480 7501 23490 7535
rect 23438 7489 23490 7501
rect 23518 7535 23570 7541
rect 23518 7501 23526 7535
rect 23526 7501 23560 7535
rect 23560 7501 23570 7535
rect 23518 7489 23570 7501
rect 23598 7535 23650 7541
rect 23598 7501 23606 7535
rect 23606 7501 23640 7535
rect 23640 7501 23650 7535
rect 23598 7489 23650 7501
rect 23678 7535 23730 7541
rect 23678 7501 23686 7535
rect 23686 7501 23720 7535
rect 23720 7501 23730 7535
rect 23678 7489 23730 7501
rect 23758 7535 23810 7541
rect 23758 7501 23766 7535
rect 23766 7501 23800 7535
rect 23800 7501 23810 7535
rect 23758 7489 23810 7501
rect 23838 7535 23890 7541
rect 23838 7501 23846 7535
rect 23846 7501 23880 7535
rect 23880 7501 23890 7535
rect 23838 7489 23890 7501
rect 24046 7535 24098 7541
rect 24046 7501 24056 7535
rect 24056 7501 24090 7535
rect 24090 7501 24098 7535
rect 24046 7489 24098 7501
rect 24126 7535 24178 7541
rect 24126 7501 24136 7535
rect 24136 7501 24170 7535
rect 24170 7501 24178 7535
rect 24126 7489 24178 7501
rect 24206 7535 24258 7541
rect 24206 7501 24216 7535
rect 24216 7501 24250 7535
rect 24250 7501 24258 7535
rect 24206 7489 24258 7501
rect 24286 7535 24338 7541
rect 24286 7501 24296 7535
rect 24296 7501 24330 7535
rect 24330 7501 24338 7535
rect 24286 7489 24338 7501
rect 24366 7535 24418 7541
rect 24366 7501 24376 7535
rect 24376 7501 24410 7535
rect 24410 7501 24418 7535
rect 24366 7489 24418 7501
rect 24446 7535 24498 7541
rect 24446 7501 24456 7535
rect 24456 7501 24490 7535
rect 24490 7501 24498 7535
rect 24446 7489 24498 7501
rect 24650 7535 24702 7541
rect 24650 7501 24658 7535
rect 24658 7501 24692 7535
rect 24692 7501 24702 7535
rect 24650 7489 24702 7501
rect 24730 7535 24782 7541
rect 24730 7501 24738 7535
rect 24738 7501 24772 7535
rect 24772 7501 24782 7535
rect 24730 7489 24782 7501
rect 24810 7535 24862 7541
rect 24810 7501 24818 7535
rect 24818 7501 24852 7535
rect 24852 7501 24862 7535
rect 24810 7489 24862 7501
rect 24890 7535 24942 7541
rect 24890 7501 24898 7535
rect 24898 7501 24932 7535
rect 24932 7501 24942 7535
rect 24890 7489 24942 7501
rect 24970 7535 25022 7541
rect 24970 7501 24978 7535
rect 24978 7501 25012 7535
rect 25012 7501 25022 7535
rect 24970 7489 25022 7501
rect 25050 7535 25102 7541
rect 25050 7501 25058 7535
rect 25058 7501 25092 7535
rect 25092 7501 25102 7535
rect 25050 7489 25102 7501
rect 25382 7538 25434 7544
rect 25382 7504 25390 7538
rect 25390 7504 25424 7538
rect 25424 7504 25434 7538
rect 25382 7492 25434 7504
rect 25462 7538 25514 7544
rect 25462 7504 25470 7538
rect 25470 7504 25504 7538
rect 25504 7504 25514 7538
rect 25462 7492 25514 7504
rect 25542 7538 25594 7544
rect 25542 7504 25550 7538
rect 25550 7504 25584 7538
rect 25584 7504 25594 7538
rect 25542 7492 25594 7504
rect 25622 7538 25674 7544
rect 25622 7504 25630 7538
rect 25630 7504 25664 7538
rect 25664 7504 25674 7538
rect 25622 7492 25674 7504
rect 25702 7538 25754 7544
rect 25702 7504 25710 7538
rect 25710 7504 25744 7538
rect 25744 7504 25754 7538
rect 25702 7492 25754 7504
rect 25782 7538 25834 7544
rect 25782 7504 25790 7538
rect 25790 7504 25824 7538
rect 25824 7504 25834 7538
rect 25782 7492 25834 7504
rect 25880 7483 25932 7535
rect 2985 7358 3038 7410
rect 9951 7358 10003 7410
rect 10629 7282 10681 7334
rect 23921 7281 23973 7333
rect 24681 7277 24733 7329
rect 24779 7308 24831 7320
rect 24779 7274 24789 7308
rect 24789 7274 24823 7308
rect 24823 7274 24831 7308
rect 24779 7268 24831 7274
rect 24859 7308 24911 7320
rect 24859 7274 24869 7308
rect 24869 7274 24903 7308
rect 24903 7274 24911 7308
rect 24859 7268 24911 7274
rect 24939 7308 24991 7320
rect 24939 7274 24949 7308
rect 24949 7274 24983 7308
rect 24983 7274 24991 7308
rect 24939 7268 24991 7274
rect 25019 7308 25071 7320
rect 25019 7274 25029 7308
rect 25029 7274 25063 7308
rect 25063 7274 25071 7308
rect 25019 7268 25071 7274
rect 25099 7308 25151 7320
rect 25099 7274 25109 7308
rect 25109 7274 25143 7308
rect 25143 7274 25151 7308
rect 25099 7268 25151 7274
rect 25179 7308 25231 7320
rect 25179 7274 25189 7308
rect 25189 7274 25223 7308
rect 25223 7274 25231 7308
rect 25179 7268 25231 7274
rect 25511 7311 25563 7323
rect 25511 7277 25521 7311
rect 25521 7277 25555 7311
rect 25555 7277 25563 7311
rect 25511 7271 25563 7277
rect 25591 7311 25643 7323
rect 25591 7277 25601 7311
rect 25601 7277 25635 7311
rect 25635 7277 25643 7311
rect 25591 7271 25643 7277
rect 25671 7311 25723 7323
rect 25671 7277 25681 7311
rect 25681 7277 25715 7311
rect 25715 7277 25723 7311
rect 25671 7271 25723 7277
rect 25751 7311 25803 7323
rect 25751 7277 25761 7311
rect 25761 7277 25795 7311
rect 25795 7277 25803 7311
rect 25751 7271 25803 7277
rect 25831 7311 25883 7323
rect 25831 7277 25841 7311
rect 25841 7277 25875 7311
rect 25875 7277 25883 7311
rect 25831 7271 25883 7277
rect 25911 7311 25963 7323
rect 25911 7277 25921 7311
rect 25921 7277 25955 7311
rect 25955 7277 25963 7311
rect 25911 7271 25963 7277
rect 26115 7311 26167 7323
rect 26115 7277 26123 7311
rect 26123 7277 26157 7311
rect 26157 7277 26167 7311
rect 26115 7271 26167 7277
rect 26195 7311 26247 7323
rect 26195 7277 26203 7311
rect 26203 7277 26237 7311
rect 26237 7277 26247 7311
rect 26195 7271 26247 7277
rect 26275 7311 26327 7323
rect 26275 7277 26283 7311
rect 26283 7277 26317 7311
rect 26317 7277 26327 7311
rect 26275 7271 26327 7277
rect 26355 7311 26407 7323
rect 26355 7277 26363 7311
rect 26363 7277 26397 7311
rect 26397 7277 26407 7311
rect 26355 7271 26407 7277
rect 26435 7311 26487 7323
rect 26435 7277 26443 7311
rect 26443 7277 26477 7311
rect 26477 7277 26487 7311
rect 26435 7271 26487 7277
rect 26515 7311 26567 7323
rect 26515 7277 26523 7311
rect 26523 7277 26557 7311
rect 26557 7277 26567 7311
rect 26515 7271 26567 7277
rect 26723 7311 26775 7323
rect 26723 7277 26733 7311
rect 26733 7277 26767 7311
rect 26767 7277 26775 7311
rect 26723 7271 26775 7277
rect 26803 7311 26855 7323
rect 26803 7277 26813 7311
rect 26813 7277 26847 7311
rect 26847 7277 26855 7311
rect 26803 7271 26855 7277
rect 26883 7311 26935 7323
rect 26883 7277 26893 7311
rect 26893 7277 26927 7311
rect 26927 7277 26935 7311
rect 26883 7271 26935 7277
rect 26963 7311 27015 7323
rect 26963 7277 26973 7311
rect 26973 7277 27007 7311
rect 27007 7277 27015 7311
rect 26963 7271 27015 7277
rect 27043 7311 27095 7323
rect 27043 7277 27053 7311
rect 27053 7277 27087 7311
rect 27087 7277 27095 7311
rect 27043 7271 27095 7277
rect 27123 7311 27175 7323
rect 27123 7277 27133 7311
rect 27133 7277 27167 7311
rect 27167 7277 27175 7311
rect 27123 7271 27175 7277
rect 27327 7311 27379 7323
rect 27327 7277 27335 7311
rect 27335 7277 27369 7311
rect 27369 7277 27379 7311
rect 27327 7271 27379 7277
rect 27407 7311 27459 7323
rect 27407 7277 27415 7311
rect 27415 7277 27449 7311
rect 27449 7277 27459 7311
rect 27407 7271 27459 7277
rect 27487 7311 27539 7323
rect 27487 7277 27495 7311
rect 27495 7277 27529 7311
rect 27529 7277 27539 7311
rect 27487 7271 27539 7277
rect 27567 7311 27619 7323
rect 27567 7277 27575 7311
rect 27575 7277 27609 7311
rect 27609 7277 27619 7311
rect 27567 7271 27619 7277
rect 27647 7311 27699 7323
rect 27647 7277 27655 7311
rect 27655 7277 27689 7311
rect 27689 7277 27699 7311
rect 27647 7271 27699 7277
rect 27727 7311 27779 7323
rect 27727 7277 27735 7311
rect 27735 7277 27769 7311
rect 27769 7277 27779 7311
rect 27727 7271 27779 7277
rect 27935 7311 27987 7323
rect 27935 7277 27945 7311
rect 27945 7277 27979 7311
rect 27979 7277 27987 7311
rect 27935 7271 27987 7277
rect 28015 7311 28067 7323
rect 28015 7277 28025 7311
rect 28025 7277 28059 7311
rect 28059 7277 28067 7311
rect 28015 7271 28067 7277
rect 28095 7311 28147 7323
rect 28095 7277 28105 7311
rect 28105 7277 28139 7311
rect 28139 7277 28147 7311
rect 28095 7271 28147 7277
rect 28175 7311 28227 7323
rect 28175 7277 28185 7311
rect 28185 7277 28219 7311
rect 28219 7277 28227 7311
rect 28175 7271 28227 7277
rect 28255 7311 28307 7323
rect 28255 7277 28265 7311
rect 28265 7277 28299 7311
rect 28299 7277 28307 7311
rect 28255 7271 28307 7277
rect 28335 7311 28387 7323
rect 28335 7277 28345 7311
rect 28345 7277 28379 7311
rect 28379 7277 28387 7311
rect 28335 7271 28387 7277
rect 28539 7311 28591 7323
rect 28539 7277 28547 7311
rect 28547 7277 28581 7311
rect 28581 7277 28591 7311
rect 28539 7271 28591 7277
rect 28619 7311 28671 7323
rect 28619 7277 28627 7311
rect 28627 7277 28661 7311
rect 28661 7277 28671 7311
rect 28619 7271 28671 7277
rect 28699 7311 28751 7323
rect 28699 7277 28707 7311
rect 28707 7277 28741 7311
rect 28741 7277 28751 7311
rect 28699 7271 28751 7277
rect 28779 7311 28831 7323
rect 28779 7277 28787 7311
rect 28787 7277 28821 7311
rect 28821 7277 28831 7311
rect 28779 7271 28831 7277
rect 28859 7311 28911 7323
rect 28859 7277 28867 7311
rect 28867 7277 28901 7311
rect 28901 7277 28911 7311
rect 28859 7271 28911 7277
rect 28939 7311 28991 7323
rect 28939 7277 28947 7311
rect 28947 7277 28981 7311
rect 28981 7277 28991 7311
rect 28939 7271 28991 7277
rect 29147 7311 29199 7323
rect 29147 7277 29157 7311
rect 29157 7277 29191 7311
rect 29191 7277 29199 7311
rect 29147 7271 29199 7277
rect 29227 7311 29279 7323
rect 29227 7277 29237 7311
rect 29237 7277 29271 7311
rect 29271 7277 29279 7311
rect 29227 7271 29279 7277
rect 29307 7311 29359 7323
rect 29307 7277 29317 7311
rect 29317 7277 29351 7311
rect 29351 7277 29359 7311
rect 29307 7271 29359 7277
rect 29387 7311 29439 7323
rect 29387 7277 29397 7311
rect 29397 7277 29431 7311
rect 29431 7277 29439 7311
rect 29387 7271 29439 7277
rect 29467 7311 29519 7323
rect 29467 7277 29477 7311
rect 29477 7277 29511 7311
rect 29511 7277 29519 7311
rect 29467 7271 29519 7277
rect 29547 7311 29599 7323
rect 29547 7277 29557 7311
rect 29557 7277 29591 7311
rect 29591 7277 29599 7311
rect 29547 7271 29599 7277
rect 29751 7311 29803 7323
rect 29751 7277 29759 7311
rect 29759 7277 29793 7311
rect 29793 7277 29803 7311
rect 29751 7271 29803 7277
rect 29831 7311 29883 7323
rect 29831 7277 29839 7311
rect 29839 7277 29873 7311
rect 29873 7277 29883 7311
rect 29831 7271 29883 7277
rect 29911 7311 29963 7323
rect 29911 7277 29919 7311
rect 29919 7277 29953 7311
rect 29953 7277 29963 7311
rect 29911 7271 29963 7277
rect 29991 7311 30043 7323
rect 29991 7277 29999 7311
rect 29999 7277 30033 7311
rect 30033 7277 30043 7311
rect 29991 7271 30043 7277
rect 30071 7311 30123 7323
rect 30071 7277 30079 7311
rect 30079 7277 30113 7311
rect 30113 7277 30123 7311
rect 30071 7271 30123 7277
rect 30151 7311 30203 7323
rect 30151 7277 30159 7311
rect 30159 7277 30193 7311
rect 30193 7277 30203 7311
rect 30151 7271 30203 7277
rect 30490 7260 30542 7267
rect 30490 7226 30501 7260
rect 30501 7226 30535 7260
rect 30535 7226 30542 7260
rect 30490 7215 30542 7226
rect 10891 6934 11041 7080
rect 11203 6918 11353 7064
rect 30495 7116 30547 7123
rect 30495 7082 30506 7116
rect 30506 7082 30540 7116
rect 30540 7082 30547 7116
rect 30495 7071 30547 7082
rect 30496 6964 30548 6971
rect 30496 6930 30507 6964
rect 30507 6930 30541 6964
rect 30541 6930 30548 6964
rect 30496 6919 30548 6930
rect 9988 6744 10040 6796
rect 12160 6789 12212 6797
rect 12160 6755 12175 6789
rect 12175 6755 12209 6789
rect 12209 6755 12212 6789
rect 12160 6745 12212 6755
rect 12483 6744 12535 6796
rect 18583 6757 18635 6809
rect 14065 6719 14117 6727
rect 14065 6685 14076 6719
rect 14076 6685 14110 6719
rect 14110 6685 14117 6719
rect 14065 6675 14117 6685
rect 20991 6681 21043 6733
rect 24064 6672 24116 6724
rect 24195 6713 24247 6723
rect 24195 6679 24212 6713
rect 24212 6679 24246 6713
rect 24246 6679 24247 6713
rect 24195 6671 24247 6679
rect 24339 6672 24391 6724
rect 14345 6658 14397 6665
rect 14345 6624 14354 6658
rect 14354 6624 14388 6658
rect 14388 6624 14397 6658
rect 14345 6613 14397 6624
rect 16194 6613 16246 6665
rect 30496 6794 30548 6801
rect 30496 6760 30507 6794
rect 30507 6760 30541 6794
rect 30541 6760 30548 6794
rect 30496 6749 30548 6760
rect 11523 6370 11575 6422
rect 12184 6370 12236 6422
rect 13914 6370 13966 6422
rect 16297 6370 16349 6422
rect 18692 6370 18744 6422
rect 21087 6370 21139 6422
rect 23383 6370 23435 6422
rect 23609 6320 23759 6466
rect 24337 6404 24389 6413
rect 24337 6370 24349 6404
rect 24349 6370 24383 6404
rect 24383 6370 24389 6404
rect 24337 6361 24389 6370
rect 30495 6637 30547 6644
rect 30495 6603 30506 6637
rect 30506 6603 30540 6637
rect 30540 6603 30547 6637
rect 30495 6592 30547 6603
rect 24082 6169 24134 6178
rect 24202 6169 24254 6178
rect 24345 6169 24397 6178
rect 24082 6135 24120 6169
rect 24120 6135 24134 6169
rect 24202 6135 24212 6169
rect 24212 6135 24246 6169
rect 24246 6135 24254 6169
rect 24345 6135 24396 6169
rect 24396 6135 24397 6169
rect 10955 5974 11105 6120
rect 11261 5986 11411 6132
rect 23026 6065 23078 6117
rect 24082 6126 24134 6135
rect 24202 6126 24254 6135
rect 24345 6126 24397 6135
rect 12485 5940 12537 5992
rect 11522 5900 11574 5909
rect 11522 5866 11530 5900
rect 11530 5866 11564 5900
rect 11564 5866 11574 5900
rect 11522 5857 11574 5866
rect 13912 5900 13964 5909
rect 13912 5866 13920 5900
rect 13920 5866 13954 5900
rect 13954 5866 13964 5900
rect 13912 5857 13964 5866
rect 12990 5847 13042 5854
rect 12990 5813 12999 5847
rect 12999 5813 13033 5847
rect 13033 5813 13042 5847
rect 12990 5802 13042 5813
rect 15756 5917 15808 5928
rect 15756 5883 15768 5917
rect 15768 5883 15802 5917
rect 15802 5883 15808 5917
rect 15756 5876 15808 5883
rect 16305 5901 16357 5910
rect 16305 5867 16313 5901
rect 16313 5867 16347 5901
rect 16347 5867 16357 5901
rect 16305 5858 16357 5867
rect 18149 5918 18201 5927
rect 18149 5884 18158 5918
rect 18158 5884 18192 5918
rect 18192 5884 18201 5918
rect 18149 5875 18201 5884
rect 18697 5900 18749 5909
rect 18697 5866 18705 5900
rect 18705 5866 18739 5900
rect 18739 5866 18749 5900
rect 18697 5857 18749 5866
rect 20540 5920 20592 5929
rect 20540 5886 20549 5920
rect 20549 5886 20583 5920
rect 20583 5886 20592 5920
rect 20540 5877 20592 5886
rect 21092 5902 21144 5911
rect 21092 5868 21100 5902
rect 21100 5868 21134 5902
rect 21134 5868 21144 5902
rect 21092 5859 21144 5868
rect 22931 5918 22983 5927
rect 22931 5884 22940 5918
rect 22940 5884 22974 5918
rect 22974 5884 22983 5918
rect 22931 5875 22983 5884
rect 23609 5894 23759 6040
rect 23921 5985 23973 6037
rect 13540 5789 13592 5796
rect 13540 5755 13550 5789
rect 13550 5755 13584 5789
rect 13584 5755 13592 5789
rect 13540 5744 13592 5755
rect 15930 5800 15982 5810
rect 15930 5766 15939 5800
rect 15939 5766 15973 5800
rect 15973 5766 15982 5800
rect 15930 5758 15982 5766
rect 16040 5769 16092 5821
rect 18319 5803 18371 5818
rect 18319 5769 18327 5803
rect 18327 5769 18361 5803
rect 18361 5769 18371 5803
rect 18319 5766 18371 5769
rect 18436 5758 18488 5810
rect 20715 5786 20767 5795
rect 20715 5752 20724 5786
rect 20724 5752 20758 5786
rect 20758 5752 20767 5786
rect 20715 5743 20767 5752
rect 20836 5774 20888 5826
rect 23106 5787 23158 5796
rect 23106 5753 23115 5787
rect 23115 5753 23149 5787
rect 23149 5753 23158 5787
rect 23106 5744 23158 5753
rect 23231 5774 23283 5826
rect 23609 5668 23759 5814
rect 24349 5783 24401 5835
rect 30413 6350 30465 6402
rect 30790 6358 30842 6410
rect 30990 6358 31042 6410
rect 25161 6139 25225 6142
rect 25161 6079 25183 6139
rect 25183 6079 25217 6139
rect 25217 6079 25225 6139
rect 25161 6078 25225 6079
rect 25893 6142 25957 6145
rect 25893 6082 25915 6142
rect 25915 6082 25949 6142
rect 25949 6082 25957 6142
rect 25893 6081 25957 6082
rect 26121 6142 26185 6145
rect 26121 6082 26129 6142
rect 26129 6082 26163 6142
rect 26163 6082 26185 6142
rect 26121 6081 26185 6082
rect 27105 6142 27169 6145
rect 27105 6082 27127 6142
rect 27127 6082 27161 6142
rect 27161 6082 27169 6142
rect 27105 6081 27169 6082
rect 27333 6142 27397 6145
rect 27333 6082 27341 6142
rect 27341 6082 27375 6142
rect 27375 6082 27397 6142
rect 27333 6081 27397 6082
rect 28317 6142 28381 6145
rect 28317 6082 28339 6142
rect 28339 6082 28373 6142
rect 28373 6082 28381 6142
rect 28317 6081 28381 6082
rect 28545 6142 28609 6145
rect 28545 6082 28553 6142
rect 28553 6082 28587 6142
rect 28587 6082 28609 6142
rect 28545 6081 28609 6082
rect 29529 6142 29593 6145
rect 29529 6082 29551 6142
rect 29551 6082 29585 6142
rect 29585 6082 29593 6142
rect 29529 6081 29593 6082
rect 29757 6142 29821 6145
rect 29757 6082 29765 6142
rect 29765 6082 29799 6142
rect 29799 6082 29821 6142
rect 29757 6081 29821 6082
rect 30501 6089 30510 6141
rect 30510 6089 30544 6141
rect 30544 6089 30553 6141
rect 25517 5941 25581 5943
rect 25517 5881 25536 5941
rect 25536 5881 25570 5941
rect 25570 5881 25581 5941
rect 25517 5879 25581 5881
rect 26249 5941 26313 5943
rect 26249 5881 26268 5941
rect 26268 5881 26302 5941
rect 26302 5881 26313 5941
rect 26249 5879 26313 5881
rect 26467 5941 26531 5943
rect 26467 5881 26478 5941
rect 26478 5881 26512 5941
rect 26512 5881 26531 5941
rect 26467 5879 26531 5881
rect 27461 5941 27525 5943
rect 27461 5881 27480 5941
rect 27480 5881 27514 5941
rect 27514 5881 27525 5941
rect 27461 5879 27525 5881
rect 27679 5941 27743 5943
rect 27679 5881 27690 5941
rect 27690 5881 27724 5941
rect 27724 5881 27743 5941
rect 27679 5879 27743 5881
rect 28799 5941 28863 5943
rect 28799 5881 28818 5941
rect 28818 5881 28852 5941
rect 28852 5881 28863 5941
rect 28799 5879 28863 5881
rect 29017 5941 29081 5943
rect 29017 5881 29028 5941
rect 29028 5881 29062 5941
rect 29062 5881 29081 5941
rect 29017 5879 29081 5881
rect 29751 5941 29815 5943
rect 29751 5881 29762 5941
rect 29762 5881 29796 5941
rect 29796 5881 29815 5941
rect 29751 5879 29815 5881
rect 30501 5886 30510 5938
rect 30510 5886 30544 5938
rect 30544 5886 30553 5938
rect 24837 5783 24889 5835
rect 10787 5346 10937 5492
rect 12991 5394 13043 5404
rect 12991 5360 13001 5394
rect 13001 5360 13035 5394
rect 13035 5360 13043 5394
rect 13905 5430 13957 5438
rect 13905 5396 13915 5430
rect 13915 5396 13949 5430
rect 13949 5396 13957 5430
rect 13905 5386 13957 5396
rect 16303 5368 16355 5420
rect 18694 5368 18746 5420
rect 12991 5352 13043 5360
rect 16297 5296 16349 5303
rect 16297 5262 16304 5296
rect 16304 5262 16338 5296
rect 16338 5262 16349 5296
rect 16297 5251 16349 5262
rect 10311 5188 10363 5240
rect 14351 5228 14403 5238
rect 14351 5194 14361 5228
rect 14361 5194 14395 5228
rect 14395 5194 14403 5228
rect 14351 5186 14403 5194
rect 18685 5296 18737 5301
rect 18685 5262 18696 5296
rect 18696 5262 18730 5296
rect 18730 5262 18737 5296
rect 18685 5249 18737 5262
rect 16746 5230 16798 5239
rect 16746 5196 16755 5230
rect 16755 5196 16789 5230
rect 16789 5196 16798 5230
rect 16746 5187 16798 5196
rect 21082 5359 21134 5411
rect 21077 5297 21129 5302
rect 21077 5263 21088 5297
rect 21088 5263 21122 5297
rect 21122 5263 21129 5297
rect 21077 5250 21129 5263
rect 19136 5231 19188 5240
rect 19136 5197 19145 5231
rect 19145 5197 19179 5231
rect 19179 5197 19188 5231
rect 19136 5188 19188 5197
rect 13819 5093 13871 5100
rect 13819 5059 13829 5093
rect 13829 5059 13863 5093
rect 13863 5059 13871 5093
rect 13819 5048 13871 5059
rect 16439 5083 16491 5135
rect 23029 5289 23081 5294
rect 23029 5255 23038 5289
rect 23038 5255 23072 5289
rect 23072 5255 23081 5289
rect 23029 5242 23081 5255
rect 21530 5228 21582 5237
rect 21530 5194 21539 5228
rect 21539 5194 21573 5228
rect 21573 5194 21582 5228
rect 21530 5185 21582 5194
rect 23383 5281 23435 5289
rect 23383 5247 23393 5281
rect 23393 5247 23427 5281
rect 23427 5247 23435 5281
rect 23383 5237 23435 5247
rect 17037 5047 17089 5099
rect 18861 5072 18913 5124
rect 19429 5048 19481 5100
rect 21249 5080 21301 5132
rect 21818 5049 21870 5101
rect 23625 4934 23775 5080
rect 11959 4806 12011 4858
rect 13819 4806 13871 4858
rect 14351 4806 14403 4858
rect 15755 4806 15807 4858
rect 16740 4806 16792 4858
rect 18147 4806 18199 4858
rect 19130 4806 19182 4858
rect 20544 4806 20596 4858
rect 21520 4806 21572 4858
rect 22932 4806 22984 4858
rect 24667 4731 24676 4751
rect 24676 4731 24710 4751
rect 24710 4731 24719 4751
rect 24667 4699 24719 4731
rect 25209 4744 25261 4754
rect 25209 4710 25217 4744
rect 25217 4710 25251 4744
rect 25251 4710 25261 4744
rect 25209 4702 25261 4710
rect 25289 4744 25341 4754
rect 25289 4710 25297 4744
rect 25297 4710 25331 4744
rect 25331 4710 25341 4744
rect 25289 4702 25341 4710
rect 25369 4744 25421 4754
rect 25369 4710 25377 4744
rect 25377 4710 25411 4744
rect 25411 4710 25421 4744
rect 25369 4702 25421 4710
rect 25449 4744 25501 4754
rect 25449 4710 25457 4744
rect 25457 4710 25491 4744
rect 25491 4710 25501 4744
rect 25449 4702 25501 4710
rect 25941 4744 25993 4754
rect 25941 4710 25949 4744
rect 25949 4710 25983 4744
rect 25983 4710 25993 4744
rect 25941 4702 25993 4710
rect 26021 4744 26073 4754
rect 26021 4710 26029 4744
rect 26029 4710 26063 4744
rect 26063 4710 26073 4744
rect 26021 4702 26073 4710
rect 26101 4744 26153 4754
rect 26101 4710 26109 4744
rect 26109 4710 26143 4744
rect 26143 4710 26153 4744
rect 26101 4702 26153 4710
rect 26181 4744 26233 4754
rect 26181 4710 26189 4744
rect 26189 4710 26223 4744
rect 26223 4710 26233 4744
rect 26181 4702 26233 4710
rect 26547 4744 26599 4754
rect 26547 4710 26557 4744
rect 26557 4710 26591 4744
rect 26591 4710 26599 4744
rect 26547 4702 26599 4710
rect 26627 4744 26679 4754
rect 26627 4710 26637 4744
rect 26637 4710 26671 4744
rect 26671 4710 26679 4744
rect 26627 4702 26679 4710
rect 26707 4744 26759 4754
rect 26707 4710 26717 4744
rect 26717 4710 26751 4744
rect 26751 4710 26759 4744
rect 26707 4702 26759 4710
rect 26787 4744 26839 4754
rect 26787 4710 26797 4744
rect 26797 4710 26831 4744
rect 26831 4710 26839 4744
rect 26787 4702 26839 4710
rect 27153 4744 27205 4754
rect 27153 4710 27161 4744
rect 27161 4710 27195 4744
rect 27195 4710 27205 4744
rect 27153 4702 27205 4710
rect 27233 4744 27285 4754
rect 27233 4710 27241 4744
rect 27241 4710 27275 4744
rect 27275 4710 27285 4744
rect 27233 4702 27285 4710
rect 27313 4744 27365 4754
rect 27313 4710 27321 4744
rect 27321 4710 27355 4744
rect 27355 4710 27365 4744
rect 27313 4702 27365 4710
rect 27393 4744 27445 4754
rect 27393 4710 27401 4744
rect 27401 4710 27435 4744
rect 27435 4710 27445 4744
rect 27393 4702 27445 4710
rect 27759 4744 27811 4754
rect 27759 4710 27769 4744
rect 27769 4710 27803 4744
rect 27803 4710 27811 4744
rect 27759 4702 27811 4710
rect 27839 4744 27891 4754
rect 27839 4710 27849 4744
rect 27849 4710 27883 4744
rect 27883 4710 27891 4744
rect 27839 4702 27891 4710
rect 27919 4744 27971 4754
rect 27919 4710 27929 4744
rect 27929 4710 27963 4744
rect 27963 4710 27971 4744
rect 27919 4702 27971 4710
rect 27999 4744 28051 4754
rect 27999 4710 28009 4744
rect 28009 4710 28043 4744
rect 28043 4710 28051 4744
rect 27999 4702 28051 4710
rect 28491 4744 28543 4754
rect 28491 4710 28499 4744
rect 28499 4710 28533 4744
rect 28533 4710 28543 4744
rect 28491 4702 28543 4710
rect 28571 4744 28623 4754
rect 28571 4710 28579 4744
rect 28579 4710 28613 4744
rect 28613 4710 28623 4744
rect 28571 4702 28623 4710
rect 28651 4744 28703 4754
rect 28651 4710 28659 4744
rect 28659 4710 28693 4744
rect 28693 4710 28703 4744
rect 28651 4702 28703 4710
rect 28731 4744 28783 4754
rect 28731 4710 28739 4744
rect 28739 4710 28773 4744
rect 28773 4710 28783 4744
rect 28731 4702 28783 4710
rect 10823 4500 10973 4646
rect 11175 4624 11210 4650
rect 11210 4624 11244 4650
rect 11244 4624 11302 4650
rect 11302 4624 11325 4650
rect 11621 4624 11670 4650
rect 11670 4624 11704 4650
rect 11704 4624 11762 4650
rect 11762 4624 11771 4650
rect 11175 4504 11325 4624
rect 11621 4504 11771 4624
rect 12187 4508 12337 4654
rect 12853 4508 13003 4654
rect 13235 4492 13385 4638
rect 29097 4744 29149 4754
rect 29097 4710 29107 4744
rect 29107 4710 29141 4744
rect 29141 4710 29149 4744
rect 29097 4702 29149 4710
rect 29177 4744 29229 4754
rect 29177 4710 29187 4744
rect 29187 4710 29221 4744
rect 29221 4710 29229 4744
rect 29177 4702 29229 4710
rect 29257 4744 29309 4754
rect 29257 4710 29267 4744
rect 29267 4710 29301 4744
rect 29301 4710 29309 4744
rect 29257 4702 29309 4710
rect 29337 4744 29389 4754
rect 29337 4710 29347 4744
rect 29347 4710 29381 4744
rect 29381 4710 29389 4744
rect 29337 4702 29389 4710
rect 30601 5716 30653 5768
rect 30410 5624 30462 5676
rect 29831 4744 29883 4754
rect 29831 4710 29841 4744
rect 29841 4710 29875 4744
rect 29875 4710 29883 4744
rect 29831 4702 29883 4710
rect 29911 4744 29963 4754
rect 29911 4710 29921 4744
rect 29921 4710 29955 4744
rect 29955 4710 29963 4744
rect 29911 4702 29963 4710
rect 29991 4744 30043 4754
rect 29991 4710 30001 4744
rect 30001 4710 30035 4744
rect 30035 4710 30043 4744
rect 29991 4702 30043 4710
rect 30071 4744 30123 4754
rect 30071 4710 30081 4744
rect 30081 4710 30115 4744
rect 30115 4710 30123 4744
rect 30071 4702 30123 4710
rect 10630 4311 10682 4363
rect 11119 4345 11171 4355
rect 11119 4311 11128 4345
rect 11128 4311 11162 4345
rect 11162 4311 11171 4345
rect 11119 4303 11171 4311
rect 11726 4346 11778 4355
rect 11726 4312 11733 4346
rect 11733 4312 11767 4346
rect 11767 4312 11778 4346
rect 11726 4303 11778 4312
rect 13085 4378 13137 4430
rect 13530 4377 13582 4429
rect 14652 4378 14704 4430
rect 12482 4305 12534 4357
rect 15756 4352 15808 4359
rect 15756 4318 15766 4352
rect 15766 4318 15800 4352
rect 15800 4318 15808 4352
rect 15756 4307 15808 4318
rect 16654 4355 16706 4363
rect 16654 4321 16663 4355
rect 16663 4321 16697 4355
rect 16697 4321 16706 4355
rect 16654 4311 16706 4321
rect 18147 4360 18199 4369
rect 14644 4285 14696 4293
rect 14644 4251 14654 4285
rect 14654 4251 14688 4285
rect 14688 4251 14696 4285
rect 18147 4326 18156 4360
rect 18156 4326 18190 4360
rect 18190 4326 18199 4360
rect 18147 4317 18199 4326
rect 19041 4355 19093 4363
rect 19041 4321 19050 4355
rect 19050 4321 19084 4355
rect 19084 4321 19093 4355
rect 19041 4311 19093 4321
rect 14644 4241 14696 4251
rect 17038 4285 17090 4292
rect 17038 4251 17046 4285
rect 17046 4251 17080 4285
rect 17080 4251 17090 4285
rect 20538 4356 20590 4365
rect 20538 4322 20547 4356
rect 20547 4322 20581 4356
rect 20581 4322 20590 4356
rect 20538 4313 20590 4322
rect 21444 4354 21496 4362
rect 21444 4320 21453 4354
rect 21453 4320 21487 4354
rect 21487 4320 21496 4354
rect 21444 4310 21496 4320
rect 17038 4240 17090 4251
rect 18604 4253 18656 4261
rect 18604 4219 18612 4253
rect 18612 4219 18646 4253
rect 18646 4219 18656 4253
rect 18604 4209 18656 4219
rect 22930 4355 22982 4364
rect 22930 4321 22939 4355
rect 22939 4321 22973 4355
rect 22973 4321 22982 4355
rect 22930 4312 22982 4321
rect 25622 4372 25674 4424
rect 28016 4372 28068 4424
rect 25714 4298 25766 4306
rect 25888 4298 25940 4305
rect 26113 4298 26165 4307
rect 26314 4298 26366 4309
rect 26537 4298 26589 4307
rect 19432 4285 19484 4291
rect 19432 4251 19438 4285
rect 19438 4251 19472 4285
rect 19472 4251 19484 4285
rect 19432 4239 19484 4251
rect 20996 4254 21048 4262
rect 20996 4220 21004 4254
rect 21004 4220 21038 4254
rect 21038 4220 21048 4254
rect 20996 4210 21048 4220
rect 21818 4285 21870 4292
rect 21818 4251 21830 4285
rect 21830 4251 21864 4285
rect 21864 4251 21870 4285
rect 21818 4240 21870 4251
rect 23386 4257 23438 4265
rect 23386 4223 23394 4257
rect 23394 4223 23428 4257
rect 23428 4223 23438 4257
rect 23386 4213 23438 4223
rect 25714 4264 25732 4298
rect 25732 4264 25766 4298
rect 25888 4264 25916 4298
rect 25916 4264 25940 4298
rect 26113 4264 26158 4298
rect 26158 4264 26165 4298
rect 26314 4264 26342 4298
rect 26342 4264 26366 4298
rect 26537 4264 26560 4298
rect 26560 4264 26589 4298
rect 25714 4254 25766 4264
rect 25888 4253 25940 4264
rect 26113 4255 26165 4264
rect 26314 4257 26366 4264
rect 26537 4255 26589 4264
rect 26746 4260 26798 4312
rect 26974 4298 27026 4305
rect 27164 4298 27216 4309
rect 27369 4298 27421 4312
rect 27568 4298 27620 4312
rect 27784 4298 27836 4307
rect 28172 4298 28224 4312
rect 28407 4298 28459 4307
rect 28649 4298 28701 4309
rect 28881 4298 28933 4310
rect 29110 4298 29162 4313
rect 29359 4298 29411 4305
rect 29577 4298 29629 4309
rect 29806 4298 29858 4305
rect 30027 4298 30079 4307
rect 26974 4264 26986 4298
rect 26986 4264 27020 4298
rect 27020 4264 27026 4298
rect 27164 4264 27170 4298
rect 27170 4264 27204 4298
rect 27204 4264 27216 4298
rect 27369 4264 27388 4298
rect 27388 4264 27421 4298
rect 27568 4264 27572 4298
rect 27572 4264 27620 4298
rect 27784 4264 27814 4298
rect 27814 4264 27836 4298
rect 28172 4264 28182 4298
rect 28182 4264 28216 4298
rect 28216 4264 28224 4298
rect 28407 4264 28458 4298
rect 28458 4264 28459 4298
rect 28649 4264 28676 4298
rect 28676 4264 28701 4298
rect 28881 4264 28918 4298
rect 28918 4264 28933 4298
rect 29110 4264 29136 4298
rect 29136 4264 29162 4298
rect 29359 4264 29378 4298
rect 29378 4264 29411 4298
rect 29577 4264 29596 4298
rect 29596 4264 29629 4298
rect 29806 4264 29838 4298
rect 29838 4264 29858 4298
rect 30027 4264 30056 4298
rect 30056 4264 30079 4298
rect 26974 4253 27026 4264
rect 27164 4257 27216 4264
rect 27369 4260 27421 4264
rect 27568 4260 27620 4264
rect 27784 4255 27836 4264
rect 28172 4260 28224 4264
rect 28407 4255 28459 4264
rect 28649 4257 28701 4264
rect 28881 4258 28933 4264
rect 29110 4261 29162 4264
rect 29359 4253 29411 4264
rect 29577 4257 29629 4264
rect 29806 4253 29858 4264
rect 30027 4255 30079 4264
rect 30243 4260 30295 4312
rect 11109 3936 11161 3988
rect 11729 3933 11781 3985
rect 13470 3931 13522 3983
rect 15850 3932 15902 3984
rect 16649 3931 16701 3983
rect 18243 3931 18295 3983
rect 19038 3932 19090 3984
rect 20630 3931 20682 3983
rect 21447 3932 21499 3984
rect 23025 3932 23077 3984
rect 23605 3942 23755 4088
rect 10905 3646 11055 3792
rect 11255 3654 11405 3800
rect 13469 3538 13521 3546
rect 13469 3504 13478 3538
rect 13478 3504 13512 3538
rect 13512 3504 13521 3538
rect 13469 3494 13521 3504
rect 11961 3478 12013 3488
rect 11961 3444 11966 3478
rect 11966 3444 12000 3478
rect 12000 3444 12013 3478
rect 11961 3436 12013 3444
rect 13082 3412 13134 3420
rect 13082 3378 13088 3412
rect 13088 3378 13122 3412
rect 13122 3378 13134 3412
rect 13082 3368 13134 3378
rect 14351 3483 14403 3494
rect 15850 3535 15902 3543
rect 15850 3501 15859 3535
rect 15859 3501 15893 3535
rect 15893 3501 15902 3535
rect 15850 3491 15902 3501
rect 18241 3539 18293 3547
rect 18241 3505 18250 3539
rect 18250 3505 18284 3539
rect 18284 3505 18293 3539
rect 18241 3495 18293 3505
rect 14351 3449 14359 3483
rect 14359 3449 14393 3483
rect 14393 3449 14403 3483
rect 14351 3442 14403 3449
rect 16744 3483 16796 3492
rect 16744 3449 16753 3483
rect 16753 3449 16787 3483
rect 16787 3449 16796 3483
rect 16744 3440 16796 3449
rect 20630 3540 20682 3548
rect 20630 3506 20639 3540
rect 20639 3506 20673 3540
rect 20673 3506 20682 3540
rect 20630 3496 20682 3506
rect 19136 3484 19188 3493
rect 19136 3450 19145 3484
rect 19145 3450 19179 3484
rect 19179 3450 19188 3484
rect 19136 3441 19188 3450
rect 23024 3540 23076 3548
rect 23024 3506 23033 3540
rect 23033 3506 23067 3540
rect 23067 3506 23076 3540
rect 23024 3496 23076 3506
rect 21529 3485 21581 3494
rect 21529 3451 21538 3485
rect 21538 3451 21572 3485
rect 21572 3451 21581 3485
rect 21529 3442 21581 3451
rect 23382 3489 23434 3497
rect 23382 3455 23390 3489
rect 23390 3455 23424 3489
rect 23424 3455 23434 3489
rect 23382 3445 23434 3455
rect 13905 3376 13957 3384
rect 11514 3353 11566 3361
rect 11514 3319 11522 3353
rect 11522 3319 11556 3353
rect 11556 3319 11566 3353
rect 11514 3309 11566 3319
rect 13905 3342 13913 3376
rect 13913 3342 13947 3376
rect 13947 3342 13957 3376
rect 13905 3332 13957 3342
rect 16296 3375 16348 3383
rect 15929 3301 15981 3353
rect 16296 3341 16304 3375
rect 16304 3341 16338 3375
rect 16338 3341 16348 3375
rect 16296 3331 16348 3341
rect 18691 3378 18743 3386
rect 18321 3301 18373 3353
rect 18691 3344 18699 3378
rect 18699 3344 18733 3378
rect 18733 3344 18743 3378
rect 18691 3334 18743 3344
rect 21080 3376 21132 3384
rect 20713 3301 20765 3353
rect 21080 3342 21088 3376
rect 21088 3342 21122 3376
rect 21122 3342 21132 3376
rect 21080 3332 21132 3342
rect 23104 3301 23156 3353
rect 23611 3264 23761 3410
rect 14914 3096 14966 3148
rect 20840 3097 20892 3149
rect 21002 3097 21054 3149
rect 24887 3103 24940 3155
rect 25613 4072 25665 4081
rect 25613 4038 25623 4072
rect 25623 4038 25657 4072
rect 25657 4038 25665 4072
rect 25613 4029 25665 4038
rect 27072 4094 27079 4119
rect 27079 4094 27113 4119
rect 27113 4094 27124 4119
rect 27072 4067 27124 4094
rect 27457 4057 27509 4068
rect 27457 4023 27462 4057
rect 27462 4023 27496 4057
rect 27496 4023 27509 4057
rect 27457 4016 27509 4023
rect 29467 4094 29471 4118
rect 29471 4094 29505 4118
rect 29505 4094 29519 4118
rect 28005 4027 28057 4039
rect 28005 3993 28012 4027
rect 28012 3993 28046 4027
rect 28046 3993 28057 4027
rect 29467 4066 29519 4094
rect 29852 4061 29904 4069
rect 29852 4027 29861 4061
rect 29861 4027 29895 4061
rect 29895 4027 29904 4061
rect 29852 4017 29904 4027
rect 28005 3987 28057 3993
rect 18605 3018 18657 3086
rect 25716 3720 25732 3723
rect 25732 3720 25768 3723
rect 25891 3720 25916 3721
rect 25916 3720 25943 3721
rect 26088 3720 26100 3723
rect 26100 3720 26140 3723
rect 26307 3720 26342 3726
rect 26342 3720 26359 3726
rect 26539 3720 26560 3722
rect 26560 3720 26591 3722
rect 26763 3720 26802 3729
rect 26802 3720 26815 3729
rect 25716 3671 25768 3720
rect 25891 3669 25943 3720
rect 26088 3671 26140 3720
rect 26307 3674 26359 3720
rect 26539 3670 26591 3720
rect 26763 3677 26815 3720
rect 26975 3665 27027 3717
rect 27197 3661 27249 3713
rect 27420 3658 27472 3710
rect 27630 3658 27682 3710
rect 27843 3658 27895 3710
rect 28160 3658 28212 3703
rect 28362 3658 28414 3706
rect 28563 3658 28615 3707
rect 28742 3658 28794 3708
rect 28934 3660 28986 3712
rect 29119 3658 29171 3709
rect 29351 3658 29403 3708
rect 29556 3658 29608 3710
rect 29762 3660 29814 3712
rect 29862 3658 29914 3709
rect 29970 3667 30022 3719
rect 30192 3668 30244 3720
rect 28160 3651 28182 3658
rect 28182 3651 28212 3658
rect 28362 3654 28366 3658
rect 28366 3654 28400 3658
rect 28400 3654 28414 3658
rect 28563 3655 28584 3658
rect 28584 3655 28615 3658
rect 28742 3656 28768 3658
rect 28768 3656 28794 3658
rect 29119 3657 29136 3658
rect 29136 3657 29171 3658
rect 29351 3656 29378 3658
rect 29378 3656 29403 3658
rect 29862 3657 29872 3658
rect 29872 3657 29914 3658
rect 25608 3422 25660 3432
rect 25608 3388 25618 3422
rect 25618 3388 25652 3422
rect 25652 3388 25660 3422
rect 25608 3380 25660 3388
rect 28004 3379 28056 3390
rect 9989 2924 10041 2976
rect 11911 2926 11963 2978
rect 19701 2961 19753 3013
rect 21251 2961 21303 3013
rect 22493 2961 22545 3013
rect 23386 2961 23438 3013
rect 27455 3350 27507 3357
rect 27455 3316 27463 3350
rect 27463 3316 27497 3350
rect 27497 3316 27507 3350
rect 27455 3305 27507 3316
rect 28004 3345 28013 3379
rect 28013 3345 28047 3379
rect 28047 3345 28056 3379
rect 28004 3338 28056 3345
rect 26697 3241 26749 3293
rect 29848 3351 29900 3358
rect 29848 3317 29856 3351
rect 29856 3317 29890 3351
rect 29890 3317 29900 3351
rect 29848 3306 29900 3317
rect 29092 3241 29144 3293
rect 12524 2904 12576 2956
rect 18435 2902 18487 2954
rect 20099 2892 20151 2944
rect 21082 2892 21134 2944
rect 29086 3080 29102 3083
rect 29102 3080 29136 3083
rect 29136 3080 29138 3083
rect 25743 3022 25795 3074
rect 25959 3027 26011 3079
rect 26165 3028 26217 3080
rect 26367 3020 26419 3072
rect 26563 3022 26615 3074
rect 26788 3024 26840 3076
rect 27003 3020 27055 3072
rect 27238 3020 27290 3072
rect 27446 3023 27498 3075
rect 27688 3023 27740 3075
rect 27886 3024 27938 3076
rect 28193 3024 28245 3076
rect 28418 3025 28470 3077
rect 28647 3024 28699 3076
rect 28863 3028 28915 3080
rect 29086 3031 29138 3080
rect 29310 3027 29362 3079
rect 29537 3018 29589 3068
rect 29750 3018 29802 3067
rect 29961 3019 30013 3071
rect 30188 3020 30240 3072
rect 29537 3016 29562 3018
rect 29562 3016 29589 3018
rect 29750 3015 29780 3018
rect 29780 3015 29802 3018
rect 15316 2824 15368 2876
rect 16302 2825 16354 2877
rect 8505 2735 8557 2787
rect 10310 2731 10362 2783
rect 17708 2756 17760 2808
rect 18691 2756 18743 2808
rect 25616 2806 25668 2817
rect 27077 2814 27079 2845
rect 27079 2814 27113 2845
rect 27113 2814 27129 2845
rect 12928 2700 12980 2752
rect 13904 2700 13956 2752
rect 10535 2637 10587 2689
rect 11515 2634 11567 2686
rect 10132 2568 10184 2620
rect 16039 2562 16091 2614
rect 16440 2561 16492 2613
rect 24482 2564 24534 2616
rect 17307 2496 17359 2548
rect 23230 2497 23282 2549
rect 18863 2429 18915 2481
rect 22089 2429 22141 2481
rect 9829 2360 9881 2412
rect 25253 2361 25305 2413
rect 9742 2291 9794 2343
rect 22859 2290 22911 2342
rect 9655 2222 9707 2274
rect 20468 2219 20520 2271
rect 9569 2152 9621 2204
rect 18076 2151 18128 2203
rect 9483 2082 9535 2134
rect 15685 2081 15737 2133
rect 9396 2013 9448 2065
rect 13291 2012 13343 2064
rect 9310 1943 9362 1995
rect 10899 1942 10951 1994
rect 25616 2772 25626 2806
rect 25626 2772 25660 2806
rect 25660 2772 25668 2806
rect 25616 2765 25668 2772
rect 27077 2793 27129 2814
rect 27460 2780 27512 2786
rect 27460 2746 27472 2780
rect 27472 2746 27506 2780
rect 27506 2746 27512 2780
rect 27460 2734 27512 2746
rect 28003 2762 28055 2774
rect 28003 2728 28010 2762
rect 28010 2728 28044 2762
rect 28044 2728 28055 2762
rect 29469 2814 29471 2847
rect 29471 2814 29505 2847
rect 29505 2814 29521 2847
rect 29469 2795 29521 2814
rect 29846 2782 29898 2793
rect 29846 2748 29856 2782
rect 29856 2748 29890 2782
rect 29890 2748 29898 2782
rect 29846 2741 29898 2748
rect 28003 2722 28055 2728
rect 27395 2440 27446 2443
rect 27446 2440 27447 2443
rect 27633 2440 27664 2445
rect 27664 2440 27685 2445
rect 27846 2440 27848 2447
rect 27848 2440 27898 2447
rect 25769 2378 25821 2429
rect 25994 2386 26046 2438
rect 26271 2383 26323 2435
rect 26492 2386 26544 2438
rect 26737 2383 26789 2435
rect 26963 2387 27015 2439
rect 27175 2385 27227 2437
rect 27395 2391 27447 2440
rect 27633 2393 27685 2440
rect 27846 2395 27898 2440
rect 28233 2385 28285 2437
rect 28580 2386 28632 2438
rect 28816 2381 28868 2433
rect 29000 2381 29052 2433
rect 29239 2383 29291 2435
rect 29442 2379 29494 2431
rect 29627 2378 29679 2428
rect 29818 2378 29870 2430
rect 30009 2382 30061 2434
rect 30195 2378 30247 2430
rect 25769 2377 25790 2378
rect 25790 2377 25821 2378
rect 29627 2376 29654 2378
rect 29654 2376 29679 2378
rect 25611 2046 25663 2057
rect 25611 2012 25622 2046
rect 25622 2012 25656 2046
rect 25656 2012 25663 2046
rect 25611 2005 25663 2012
rect 27455 2070 27507 2078
rect 27455 2036 27464 2070
rect 27464 2036 27498 2070
rect 27498 2036 27507 2070
rect 27455 2026 27507 2036
rect 28004 2076 28056 2087
rect 28004 2042 28011 2076
rect 28011 2042 28045 2076
rect 28045 2042 28056 2076
rect 28004 2035 28056 2042
rect 26706 1961 26758 2013
rect 29847 2071 29899 2079
rect 29847 2037 29856 2071
rect 29856 2037 29890 2071
rect 29890 2037 29899 2071
rect 29847 2027 29899 2037
rect 29096 1961 29149 2013
rect 9224 1873 9276 1925
rect 23061 1872 23113 1924
rect 9138 1803 9190 1855
rect 20672 1802 20724 1854
rect 25642 1795 25694 1847
rect 25847 1834 25899 1843
rect 26033 1834 26085 1848
rect 26227 1834 26279 1841
rect 26446 1834 26498 1846
rect 25847 1800 25882 1834
rect 25882 1800 25899 1834
rect 26033 1800 26066 1834
rect 26066 1800 26085 1834
rect 26227 1800 26250 1834
rect 26250 1800 26279 1834
rect 26446 1800 26468 1834
rect 26468 1800 26498 1834
rect 25847 1791 25899 1800
rect 26033 1796 26085 1800
rect 26227 1789 26279 1800
rect 26446 1794 26498 1800
rect 26656 1794 26708 1846
rect 26885 1834 26937 1843
rect 27131 1834 27183 1843
rect 27405 1834 27457 1843
rect 27680 1834 27732 1843
rect 27916 1834 27968 1843
rect 28139 1834 28191 1846
rect 28357 1834 28409 1849
rect 28535 1834 28587 1840
rect 26885 1800 26894 1834
rect 26894 1800 26928 1834
rect 26928 1800 26937 1834
rect 27131 1800 27170 1834
rect 27170 1800 27183 1834
rect 27405 1800 27446 1834
rect 27446 1800 27457 1834
rect 27680 1800 27722 1834
rect 27722 1800 27732 1834
rect 27916 1800 27940 1834
rect 27940 1800 27968 1834
rect 28139 1800 28182 1834
rect 28182 1800 28191 1834
rect 28357 1800 28366 1834
rect 28366 1800 28400 1834
rect 28400 1800 28409 1834
rect 28535 1800 28550 1834
rect 28550 1800 28584 1834
rect 28584 1800 28587 1834
rect 26885 1791 26937 1800
rect 27131 1791 27183 1800
rect 27405 1791 27457 1800
rect 27680 1791 27732 1800
rect 27916 1791 27968 1800
rect 28139 1794 28191 1800
rect 28357 1797 28409 1800
rect 28535 1788 28587 1800
rect 28774 1790 28826 1842
rect 28971 1834 29023 1842
rect 29169 1834 29221 1842
rect 29382 1834 29434 1843
rect 29605 1834 29657 1842
rect 29802 1834 29854 1847
rect 30018 1834 30070 1845
rect 30227 1834 30279 1845
rect 28971 1800 29010 1834
rect 29010 1800 29023 1834
rect 29169 1800 29194 1834
rect 29194 1800 29221 1834
rect 29382 1800 29412 1834
rect 29412 1800 29434 1834
rect 29605 1800 29654 1834
rect 29654 1800 29657 1834
rect 29802 1800 29838 1834
rect 29838 1800 29854 1834
rect 30018 1800 30022 1834
rect 30022 1800 30056 1834
rect 30056 1800 30070 1834
rect 30227 1800 30240 1834
rect 30240 1800 30279 1834
rect 28971 1790 29023 1800
rect 29169 1790 29221 1800
rect 29382 1791 29434 1800
rect 29605 1790 29657 1800
rect 29802 1795 29854 1800
rect 30018 1793 30070 1800
rect 30227 1793 30279 1800
rect 9051 1734 9103 1786
rect 18279 1733 18331 1785
rect 8965 1664 9017 1716
rect 15886 1663 15938 1715
rect 8878 1595 8930 1647
rect 13494 1594 13546 1646
rect 8792 1525 8844 1577
rect 11104 1523 11156 1575
rect 8628 1406 8680 1411
rect 8628 1372 8640 1406
rect 8640 1372 8680 1406
rect 8628 1359 8680 1372
rect 8830 1361 8882 1413
rect 9041 1406 9093 1411
rect 9231 1406 9283 1411
rect 9439 1406 9491 1413
rect 9641 1406 9693 1413
rect 9041 1372 9066 1406
rect 9066 1372 9093 1406
rect 9231 1372 9250 1406
rect 9250 1372 9283 1406
rect 9439 1372 9468 1406
rect 9468 1372 9491 1406
rect 9641 1372 9652 1406
rect 9652 1372 9693 1406
rect 9041 1359 9093 1372
rect 9231 1359 9283 1372
rect 9439 1361 9491 1372
rect 9641 1361 9693 1372
rect 9840 1363 9892 1415
rect 10035 1406 10087 1412
rect 10236 1406 10288 1414
rect 10453 1406 10505 1412
rect 10727 1406 10779 1415
rect 11004 1406 11056 1408
rect 11227 1406 11279 1411
rect 10035 1372 10078 1406
rect 10078 1372 10087 1406
rect 10236 1372 10262 1406
rect 10262 1372 10288 1406
rect 10453 1372 10480 1406
rect 10480 1372 10505 1406
rect 10727 1372 10756 1406
rect 10756 1372 10779 1406
rect 11004 1372 11032 1406
rect 11032 1372 11056 1406
rect 11227 1372 11274 1406
rect 11274 1372 11279 1406
rect 10035 1360 10087 1372
rect 10236 1362 10288 1372
rect 10453 1360 10505 1372
rect 10727 1363 10779 1372
rect 11004 1356 11056 1372
rect 11227 1359 11279 1372
rect 11459 1358 11511 1410
rect 13095 1406 13147 1407
rect 13403 1406 13455 1408
rect 13603 1406 13655 1409
rect 13822 1406 13874 1408
rect 14068 1406 14120 1407
rect 14276 1406 14328 1409
rect 14478 1406 14530 1410
rect 14671 1406 14723 1409
rect 15043 1406 15095 1408
rect 13095 1372 13116 1406
rect 13116 1372 13147 1406
rect 13403 1372 13450 1406
rect 13450 1372 13455 1406
rect 13603 1372 13634 1406
rect 13634 1372 13655 1406
rect 13822 1372 13852 1406
rect 13852 1372 13874 1406
rect 14068 1372 14094 1406
rect 14094 1372 14120 1406
rect 14276 1372 14278 1406
rect 14278 1372 14312 1406
rect 14312 1372 14328 1406
rect 14478 1372 14496 1406
rect 14496 1372 14530 1406
rect 14671 1372 14680 1406
rect 14680 1372 14723 1406
rect 15043 1372 15048 1406
rect 15048 1372 15095 1406
rect 13095 1355 13147 1372
rect 13403 1356 13455 1372
rect 13603 1357 13655 1372
rect 13822 1356 13874 1372
rect 14068 1355 14120 1372
rect 14276 1357 14328 1372
rect 14478 1358 14530 1372
rect 14671 1357 14723 1372
rect 15043 1356 15095 1372
rect 15232 1354 15284 1406
rect 15522 1372 15566 1406
rect 15566 1372 15574 1406
rect 15522 1354 15574 1372
rect 15795 1356 15847 1408
rect 8497 1164 8549 1216
rect 11441 1099 11493 1109
rect 11441 1065 11451 1099
rect 11451 1065 11485 1099
rect 11485 1065 11493 1099
rect 11441 1057 11493 1065
rect 11916 967 11968 1019
rect 16002 1057 16054 1109
rect 9746 820 9798 872
rect 9965 862 10017 876
rect 10248 862 10300 876
rect 10457 862 10509 876
rect 10728 862 10780 874
rect 9965 828 9986 862
rect 9986 828 10017 862
rect 10248 828 10262 862
rect 10262 828 10296 862
rect 10296 828 10300 862
rect 10457 828 10480 862
rect 10480 828 10509 862
rect 10728 828 10756 862
rect 10756 828 10780 862
rect 9965 824 10017 828
rect 10248 824 10300 828
rect 10457 824 10509 828
rect 10728 822 10780 828
rect 12803 820 12855 872
rect 13052 862 13104 875
rect 13650 862 13702 867
rect 13879 862 13931 867
rect 15597 862 15649 872
rect 13052 828 13082 862
rect 13082 828 13104 862
rect 13052 823 13104 828
rect 13396 809 13448 861
rect 13650 828 13668 862
rect 13668 828 13702 862
rect 13879 828 13910 862
rect 13910 828 13931 862
rect 15597 828 15600 862
rect 15600 828 15649 862
rect 13650 815 13702 828
rect 13879 815 13931 828
rect 15597 820 15649 828
rect 15801 822 15853 874
rect 16124 820 16176 872
rect 9599 685 9652 738
rect 11441 685 11493 737
rect 11993 691 12046 744
rect 14384 691 14437 744
rect 16775 691 16828 744
rect 19167 691 19220 744
rect 21558 691 21611 744
rect 23951 691 24004 744
rect 9049 474 9101 526
rect 10311 474 10363 526
rect 11442 473 11494 525
rect 12703 474 12755 526
rect 13834 473 13886 525
rect 15094 475 15146 527
rect 16002 473 16054 525
rect 16226 474 16278 526
rect 17487 475 17539 527
rect 18617 473 18669 525
rect 19880 475 19932 527
rect 21009 472 21061 524
rect 22269 475 22321 527
rect 23401 473 23453 525
rect 24664 475 24716 527
rect 8594 264 8646 267
rect 8834 264 8886 265
rect 8594 230 8604 264
rect 8604 230 8638 264
rect 8638 230 8646 264
rect 8834 230 8880 264
rect 8880 230 8886 264
rect 9156 230 9190 264
rect 9190 230 9208 264
rect 8594 215 8646 230
rect 8834 213 8886 230
rect 9156 212 9208 230
rect 9374 213 9426 265
rect 11278 264 11330 269
rect 11603 264 11655 271
rect 11278 230 11306 264
rect 11306 230 11330 264
rect 11603 230 11640 264
rect 11640 230 11655 264
rect 11278 217 11330 230
rect 11603 219 11655 230
rect 11871 219 11923 271
rect 12137 219 12189 271
rect 12377 217 12429 269
rect 14171 220 14223 272
rect 14537 223 14589 275
rect 14781 264 14833 275
rect 15204 264 15256 266
rect 14781 230 14820 264
rect 14820 230 14833 264
rect 15204 230 15222 264
rect 15222 230 15256 264
rect 14781 223 14833 230
rect 15204 214 15256 230
rect 17147 216 17199 268
rect 17399 264 17451 265
rect 17605 264 17657 273
rect 17888 264 17940 267
rect 18186 264 18238 268
rect 20018 264 20070 269
rect 20228 264 20280 271
rect 20579 264 20631 269
rect 20859 264 20911 269
rect 21176 264 21228 268
rect 22966 264 23018 266
rect 23261 264 23313 266
rect 17399 230 17432 264
rect 17432 230 17451 264
rect 17605 230 17616 264
rect 17616 230 17657 264
rect 17888 230 17892 264
rect 17892 230 17940 264
rect 18186 230 18206 264
rect 18206 230 18238 264
rect 20018 230 20066 264
rect 20066 230 20070 264
rect 20228 230 20250 264
rect 20250 230 20280 264
rect 20579 230 20598 264
rect 20598 230 20631 264
rect 20859 230 20874 264
rect 20874 230 20911 264
rect 21176 230 21208 264
rect 21208 230 21228 264
rect 22966 230 22990 264
rect 22990 230 23018 264
rect 23261 230 23266 264
rect 23266 230 23313 264
rect 17399 213 17451 230
rect 17605 221 17657 230
rect 17888 215 17940 230
rect 18186 216 18238 230
rect 20018 217 20070 230
rect 20228 219 20280 230
rect 20579 217 20631 230
rect 20859 217 20911 230
rect 21176 216 21228 230
rect 22966 214 23018 230
rect 23261 214 23313 230
rect 23548 214 23600 266
rect 23838 214 23890 266
rect 24122 217 24174 269
rect 9050 42 9102 52
rect 9050 8 9059 42
rect 9059 8 9093 42
rect 9093 8 9102 42
rect 9050 0 9102 8
rect 10132 27 10184 38
rect 10132 -7 10141 27
rect 10141 -7 10175 27
rect 10175 -7 10184 27
rect 10132 -15 10184 -7
rect 10312 42 10364 52
rect 10312 8 10321 42
rect 10321 8 10355 42
rect 10355 8 10364 42
rect 10312 0 10364 8
rect 11443 41 11495 51
rect 11443 7 11452 41
rect 11452 7 11486 41
rect 11486 7 11495 41
rect 11443 -1 11495 7
rect 12524 26 12576 37
rect 12524 -8 12533 26
rect 12533 -8 12567 26
rect 12567 -8 12576 26
rect 12524 -16 12576 -8
rect 12704 42 12756 52
rect 12704 8 12713 42
rect 12713 8 12747 42
rect 12747 8 12756 42
rect 12704 0 12756 8
rect 13835 41 13887 51
rect 13835 7 13844 41
rect 13844 7 13878 41
rect 13878 7 13887 41
rect 13835 -1 13887 7
rect 14914 26 14966 37
rect 14914 -8 14923 26
rect 14923 -8 14957 26
rect 14957 -8 14966 26
rect 14914 -16 14966 -8
rect 15095 43 15147 53
rect 15095 9 15104 43
rect 15104 9 15138 43
rect 15138 9 15147 43
rect 15095 1 15147 9
rect 16227 42 16279 52
rect 16227 8 16236 42
rect 16236 8 16270 42
rect 16270 8 16279 42
rect 16227 0 16279 8
rect 17308 27 17360 38
rect 17308 -7 17317 27
rect 17317 -7 17351 27
rect 17351 -7 17360 27
rect 17308 -15 17360 -7
rect 17488 43 17540 53
rect 17488 9 17497 43
rect 17497 9 17531 43
rect 17531 9 17540 43
rect 17488 1 17540 9
rect 18618 41 18670 51
rect 18618 7 18627 41
rect 18627 7 18661 41
rect 18661 7 18670 41
rect 18618 -1 18670 7
rect 19700 26 19752 37
rect 19700 -8 19709 26
rect 19709 -8 19743 26
rect 19743 -8 19752 26
rect 19700 -16 19752 -8
rect 19881 43 19933 53
rect 19881 9 19890 43
rect 19890 9 19924 43
rect 19924 9 19933 43
rect 19881 1 19933 9
rect 21010 40 21062 50
rect 21010 6 21019 40
rect 21019 6 21053 40
rect 21053 6 21062 40
rect 21010 -2 21062 6
rect 22089 26 22141 37
rect 22089 -8 22098 26
rect 22098 -8 22132 26
rect 22132 -8 22141 26
rect 22089 -16 22141 -8
rect 22270 43 22322 53
rect 22270 9 22279 43
rect 22279 9 22313 43
rect 22313 9 22322 43
rect 22270 1 22322 9
rect 23402 41 23454 51
rect 23402 7 23411 41
rect 23411 7 23445 41
rect 23445 7 23454 41
rect 23402 -1 23454 7
rect 24484 27 24536 38
rect 24484 -7 24493 27
rect 24493 -7 24527 27
rect 24527 -7 24536 27
rect 24484 -15 24536 -7
rect 24665 43 24717 53
rect 24665 9 24674 43
rect 24674 9 24708 43
rect 24708 9 24717 43
rect 24665 1 24717 9
rect 8593 -159 8645 -151
rect 8593 -193 8603 -159
rect 8603 -193 8637 -159
rect 8637 -193 8645 -159
rect 8593 -203 8645 -193
rect 8931 -165 8983 -113
rect 10532 -164 10584 -112
rect 10769 -161 10821 -151
rect 10769 -195 10779 -161
rect 10779 -195 10813 -161
rect 10813 -195 10821 -161
rect 10769 -203 10821 -195
rect 10985 -159 11037 -151
rect 10985 -193 10995 -159
rect 10995 -193 11029 -159
rect 11029 -193 11037 -159
rect 10985 -203 11037 -193
rect 11323 -165 11375 -113
rect 12924 -164 12976 -112
rect 13163 -161 13215 -151
rect 13163 -195 13173 -161
rect 13173 -195 13207 -161
rect 13207 -195 13215 -161
rect 13163 -203 13215 -195
rect 13377 -159 13429 -151
rect 13377 -193 13387 -159
rect 13387 -193 13421 -159
rect 13421 -193 13429 -159
rect 13377 -203 13429 -193
rect 13714 -164 13766 -112
rect 15315 -163 15367 -111
rect 15553 -159 15605 -149
rect 15553 -193 15563 -159
rect 15563 -193 15597 -159
rect 15597 -193 15605 -159
rect 15553 -201 15605 -193
rect 15769 -159 15821 -151
rect 15769 -193 15779 -159
rect 15779 -193 15813 -159
rect 15813 -193 15821 -159
rect 15769 -203 15821 -193
rect 16107 -165 16159 -113
rect 17708 -164 17760 -112
rect 17945 -161 17997 -151
rect 17945 -195 17955 -161
rect 17955 -195 17989 -161
rect 17989 -195 17997 -161
rect 17945 -203 17997 -195
rect 18160 -158 18212 -150
rect 18160 -192 18170 -158
rect 18170 -192 18204 -158
rect 18204 -192 18212 -158
rect 18160 -202 18212 -192
rect 18499 -164 18551 -112
rect 20100 -163 20152 -111
rect 20337 -159 20389 -149
rect 20337 -193 20347 -159
rect 20347 -193 20381 -159
rect 20381 -193 20389 -159
rect 20337 -201 20389 -193
rect 20552 -159 20604 -151
rect 20552 -193 20562 -159
rect 20562 -193 20596 -159
rect 20596 -193 20604 -159
rect 20552 -203 20604 -193
rect 20891 -164 20943 -112
rect 22492 -163 22544 -111
rect 22729 -161 22781 -151
rect 22729 -195 22739 -161
rect 22739 -195 22773 -161
rect 22773 -195 22781 -161
rect 22729 -203 22781 -195
rect 22945 -158 22997 -150
rect 22945 -192 22955 -158
rect 22955 -192 22989 -158
rect 22989 -192 22997 -158
rect 22945 -202 22997 -192
rect 23286 -164 23338 -112
rect 24887 -163 24939 -111
rect 25121 -159 25173 -149
rect 25121 -193 25131 -159
rect 25131 -193 25165 -159
rect 25165 -193 25173 -159
rect 25121 -201 25173 -193
rect 9785 -323 9837 -271
rect 10002 -280 10054 -271
rect 10221 -280 10273 -271
rect 10434 -280 10486 -275
rect 10645 -280 10697 -275
rect 12769 -280 12821 -275
rect 13047 -280 13099 -276
rect 13619 -280 13671 -271
rect 13858 -280 13910 -271
rect 16016 -280 16068 -273
rect 16243 -280 16295 -268
rect 16433 -280 16485 -266
rect 10002 -314 10038 -280
rect 10038 -314 10054 -280
rect 10221 -314 10222 -280
rect 10222 -314 10256 -280
rect 10256 -314 10273 -280
rect 10434 -314 10440 -280
rect 10440 -314 10486 -280
rect 10645 -314 10682 -280
rect 10682 -314 10697 -280
rect 12769 -314 12798 -280
rect 12798 -314 12821 -280
rect 13047 -314 13074 -280
rect 13074 -314 13099 -280
rect 13619 -314 13664 -280
rect 13664 -314 13671 -280
rect 13858 -314 13882 -280
rect 13882 -314 13910 -280
rect 16016 -314 16056 -280
rect 16056 -314 16068 -280
rect 16243 -314 16274 -280
rect 16274 -314 16295 -280
rect 16433 -314 16458 -280
rect 16458 -314 16485 -280
rect 10002 -323 10054 -314
rect 10221 -323 10273 -314
rect 10434 -327 10486 -314
rect 10645 -327 10697 -314
rect 12769 -327 12821 -314
rect 13047 -328 13099 -314
rect 13619 -323 13671 -314
rect 13858 -323 13910 -314
rect 16016 -325 16068 -314
rect 16243 -320 16295 -314
rect 16433 -318 16485 -314
rect 16649 -327 16701 -275
rect 18630 -280 18682 -272
rect 18859 -280 18911 -269
rect 18630 -314 18632 -280
rect 18632 -314 18666 -280
rect 18666 -314 18682 -280
rect 18859 -314 18908 -280
rect 18908 -314 18911 -280
rect 18630 -324 18682 -314
rect 18859 -321 18911 -314
rect 19085 -316 19137 -264
rect 19313 -324 19365 -272
rect 19549 -318 19601 -266
rect 19741 -280 19793 -275
rect 19741 -314 19790 -280
rect 19790 -314 19793 -280
rect 19741 -327 19793 -314
rect 21476 -327 21528 -275
rect 21680 -322 21732 -270
rect 21871 -327 21923 -275
rect 22073 -280 22125 -276
rect 22363 -280 22415 -275
rect 22648 -280 22700 -276
rect 24403 -280 24455 -271
rect 24597 -280 24649 -267
rect 24786 -280 24838 -270
rect 25009 -280 25061 -268
rect 22073 -314 22088 -280
rect 22088 -314 22122 -280
rect 22122 -314 22125 -280
rect 22363 -314 22364 -280
rect 22364 -314 22398 -280
rect 22398 -314 22415 -280
rect 22648 -314 22674 -280
rect 22674 -314 22700 -280
rect 24403 -314 24424 -280
rect 24424 -314 24455 -280
rect 24597 -314 24608 -280
rect 24608 -314 24649 -280
rect 24786 -314 24792 -280
rect 24792 -314 24838 -280
rect 25009 -314 25034 -280
rect 25034 -314 25061 -280
rect 22073 -328 22125 -314
rect 22363 -327 22415 -314
rect 22648 -328 22700 -314
rect 24403 -323 24455 -314
rect 24597 -319 24649 -314
rect 24786 -322 24838 -314
rect 25009 -320 25061 -314
rect 8840 -424 8892 -416
rect 9042 -424 9094 -420
rect 9231 -424 9283 -423
rect 9460 -424 9512 -422
rect 11229 -424 11281 -419
rect 11444 -424 11496 -422
rect 11837 -424 11889 -415
rect 12117 -424 12169 -417
rect 12336 -424 12388 -419
rect 14157 -424 14209 -422
rect 14902 -424 14954 -420
rect 15093 -424 15145 -418
rect 17138 -424 17190 -416
rect 17328 -424 17380 -414
rect 17522 -424 17574 -416
rect 17833 -424 17885 -420
rect 20016 -424 20068 -421
rect 20220 -424 20272 -421
rect 21024 -424 21076 -423
rect 21228 -424 21280 -423
rect 23188 -424 23240 -415
rect 23421 -424 23473 -417
rect 23628 -424 23680 -419
rect 23837 -424 23889 -417
rect 24117 -424 24169 -415
rect 8840 -458 8880 -424
rect 8880 -458 8892 -424
rect 9042 -458 9064 -424
rect 9064 -458 9094 -424
rect 9231 -458 9248 -424
rect 9248 -458 9282 -424
rect 9282 -458 9283 -424
rect 9460 -458 9466 -424
rect 9466 -458 9512 -424
rect 11229 -458 11272 -424
rect 11272 -458 11281 -424
rect 11444 -458 11456 -424
rect 11456 -458 11490 -424
rect 11490 -458 11496 -424
rect 11642 -458 11674 -425
rect 11674 -458 11694 -425
rect 11837 -458 11858 -424
rect 11858 -458 11889 -424
rect 12117 -458 12134 -424
rect 12134 -458 12169 -424
rect 12336 -458 12376 -424
rect 12376 -458 12388 -424
rect 14157 -458 14158 -424
rect 14158 -458 14209 -424
rect 14508 -458 14526 -425
rect 14526 -458 14560 -425
rect 14697 -458 14710 -427
rect 14710 -458 14749 -427
rect 14902 -458 14952 -424
rect 14952 -458 14954 -424
rect 15093 -458 15136 -424
rect 15136 -458 15145 -424
rect 17138 -458 17160 -424
rect 17160 -458 17190 -424
rect 17328 -458 17344 -424
rect 17344 -458 17378 -424
rect 17378 -458 17380 -424
rect 17522 -458 17528 -424
rect 17528 -458 17562 -424
rect 17562 -458 17574 -424
rect 17833 -458 17838 -424
rect 17838 -458 17885 -424
rect 20016 -458 20046 -424
rect 20046 -458 20068 -424
rect 20220 -458 20230 -424
rect 20230 -458 20272 -424
rect 8840 -468 8892 -458
rect 9042 -472 9094 -458
rect 9231 -475 9283 -458
rect 9460 -474 9512 -458
rect 11229 -471 11281 -458
rect 11444 -474 11496 -458
rect 11642 -477 11694 -458
rect 11837 -467 11889 -458
rect 12117 -469 12169 -458
rect 12336 -471 12388 -458
rect 14157 -474 14209 -458
rect 14508 -477 14560 -458
rect 14697 -479 14749 -458
rect 14902 -472 14954 -458
rect 15093 -470 15145 -458
rect 17138 -468 17190 -458
rect 17328 -466 17380 -458
rect 17522 -468 17574 -458
rect 17833 -472 17885 -458
rect 20016 -473 20068 -458
rect 20220 -473 20272 -458
rect 20785 -477 20837 -425
rect 21024 -458 21058 -424
rect 21058 -458 21076 -424
rect 21228 -458 21242 -424
rect 21242 -458 21280 -424
rect 23188 -458 23232 -424
rect 23232 -458 23240 -424
rect 23421 -458 23450 -424
rect 23450 -458 23473 -424
rect 23628 -458 23634 -424
rect 23634 -458 23680 -424
rect 23837 -458 23876 -424
rect 23876 -458 23889 -424
rect 24117 -458 24152 -424
rect 24152 -458 24169 -424
rect 21024 -475 21076 -458
rect 21228 -475 21280 -458
rect 23188 -467 23240 -458
rect 23421 -469 23473 -458
rect 23628 -471 23680 -458
rect 23837 -469 23889 -458
rect 24117 -467 24169 -458
rect 10899 -531 10951 -523
rect 10899 -565 10909 -531
rect 10909 -565 10943 -531
rect 10943 -565 10951 -531
rect 10899 -575 10951 -565
rect 13291 -531 13343 -523
rect 13291 -565 13301 -531
rect 13301 -565 13335 -531
rect 13335 -565 13343 -531
rect 13291 -575 13343 -565
rect 15683 -531 15735 -523
rect 15683 -565 15693 -531
rect 15693 -565 15727 -531
rect 15727 -565 15735 -531
rect 15683 -575 15735 -565
rect 18075 -531 18127 -523
rect 18075 -565 18085 -531
rect 18085 -565 18119 -531
rect 18119 -565 18127 -531
rect 18075 -575 18127 -565
rect 20467 -531 20519 -523
rect 20467 -565 20477 -531
rect 20477 -565 20511 -531
rect 20511 -565 20519 -531
rect 20467 -575 20519 -565
rect 22859 -531 22911 -523
rect 22859 -565 22869 -531
rect 22869 -565 22903 -531
rect 22903 -565 22911 -531
rect 22859 -575 22911 -565
rect 25251 -531 25303 -523
rect 25251 -565 25261 -531
rect 25261 -565 25295 -531
rect 25295 -565 25303 -531
rect 25251 -575 25303 -565
rect 10617 -610 10669 -600
rect 10617 -644 10626 -610
rect 10626 -644 10660 -610
rect 10660 -644 10669 -610
rect 13009 -609 13061 -599
rect 10617 -652 10669 -644
rect 8593 -706 8645 -696
rect 8593 -740 8601 -706
rect 8601 -740 8635 -706
rect 8635 -740 8645 -706
rect 8593 -748 8645 -740
rect 8932 -682 8984 -671
rect 8932 -716 8941 -682
rect 8941 -716 8975 -682
rect 8975 -716 8984 -682
rect 8932 -724 8984 -716
rect 13009 -643 13018 -609
rect 13018 -643 13052 -609
rect 13052 -643 13061 -609
rect 15400 -609 15452 -599
rect 13009 -651 13061 -643
rect 10985 -706 11037 -696
rect 10985 -740 10993 -706
rect 10993 -740 11027 -706
rect 11027 -740 11037 -706
rect 10985 -748 11037 -740
rect 11324 -682 11376 -671
rect 11324 -716 11333 -682
rect 11333 -716 11367 -682
rect 11367 -716 11376 -682
rect 11324 -724 11376 -716
rect 15400 -643 15409 -609
rect 15409 -643 15443 -609
rect 15443 -643 15452 -609
rect 17793 -608 17845 -598
rect 15400 -651 15452 -643
rect 13377 -706 13429 -696
rect 13377 -740 13385 -706
rect 13385 -740 13419 -706
rect 13419 -740 13429 -706
rect 13377 -748 13429 -740
rect 13716 -681 13768 -670
rect 13716 -715 13725 -681
rect 13725 -715 13759 -681
rect 13759 -715 13768 -681
rect 13716 -723 13768 -715
rect 17793 -642 17802 -608
rect 17802 -642 17836 -608
rect 17836 -642 17845 -608
rect 20184 -609 20236 -599
rect 17793 -650 17845 -642
rect 20184 -643 20193 -609
rect 20193 -643 20227 -609
rect 20227 -643 20236 -609
rect 22577 -610 22629 -600
rect 20184 -651 20236 -643
rect 9600 -847 9652 -795
rect 15769 -706 15821 -696
rect 15769 -740 15777 -706
rect 15777 -740 15811 -706
rect 15811 -740 15821 -706
rect 15769 -748 15821 -740
rect 16108 -681 16160 -670
rect 16108 -715 16117 -681
rect 16117 -715 16151 -681
rect 16151 -715 16160 -681
rect 16108 -723 16160 -715
rect 11993 -847 12045 -795
rect 18160 -705 18212 -695
rect 18160 -739 18168 -705
rect 18168 -739 18202 -705
rect 18202 -739 18212 -705
rect 18160 -747 18212 -739
rect 18500 -682 18552 -671
rect 18500 -716 18509 -682
rect 18509 -716 18543 -682
rect 18543 -716 18552 -682
rect 18500 -724 18552 -716
rect 22577 -644 22586 -610
rect 22586 -644 22620 -610
rect 22620 -644 22629 -610
rect 24970 -608 25022 -598
rect 22577 -652 22629 -644
rect 14385 -847 14437 -795
rect 20552 -706 20604 -696
rect 20552 -740 20560 -706
rect 20560 -740 20594 -706
rect 20594 -740 20604 -706
rect 20552 -748 20604 -740
rect 20892 -681 20944 -670
rect 20892 -715 20901 -681
rect 20901 -715 20935 -681
rect 20935 -715 20944 -681
rect 20892 -723 20944 -715
rect 24970 -642 24979 -608
rect 24979 -642 25013 -608
rect 25013 -642 25022 -608
rect 24970 -650 25022 -642
rect 16777 -847 16829 -795
rect 22945 -705 22997 -695
rect 22945 -739 22953 -705
rect 22953 -739 22987 -705
rect 22987 -739 22997 -705
rect 22945 -747 22997 -739
rect 23285 -682 23337 -671
rect 23285 -716 23294 -682
rect 23294 -716 23328 -682
rect 23328 -716 23337 -682
rect 23285 -724 23337 -716
rect 19168 -847 19220 -795
rect 21560 -847 21612 -795
rect 23952 -847 24004 -795
rect 9767 -968 9819 -965
rect 9996 -968 10048 -953
rect 10215 -968 10267 -963
rect 10407 -968 10459 -959
rect 10901 -968 10953 -961
rect 12693 -968 12745 -962
rect 13086 -968 13138 -964
rect 13283 -968 13335 -956
rect 13613 -968 13665 -954
rect 13809 -968 13861 -954
rect 15716 -968 15768 -961
rect 16017 -968 16069 -957
rect 16223 -968 16275 -956
rect 16433 -968 16485 -960
rect 9767 -1002 9800 -968
rect 9800 -1002 9819 -968
rect 9996 -1002 10018 -968
rect 10018 -1002 10048 -968
rect 10215 -1002 10260 -968
rect 10260 -1002 10267 -968
rect 10407 -1002 10444 -968
rect 10444 -1002 10459 -968
rect 10901 -1002 10904 -968
rect 10904 -1002 10938 -968
rect 10938 -1002 10953 -968
rect 12693 -1002 12744 -968
rect 12744 -1002 12745 -968
rect 13086 -1002 13112 -968
rect 13112 -1002 13138 -968
rect 13283 -1002 13296 -968
rect 13296 -1002 13330 -968
rect 13330 -1002 13335 -968
rect 13613 -1002 13664 -968
rect 13664 -1002 13665 -968
rect 13809 -1002 13848 -968
rect 13848 -1002 13861 -968
rect 15716 -1002 15722 -968
rect 15722 -1002 15768 -968
rect 16017 -1002 16056 -968
rect 16056 -1002 16069 -968
rect 16223 -1002 16240 -968
rect 16240 -1002 16274 -968
rect 16274 -1002 16275 -968
rect 16433 -1002 16458 -968
rect 16458 -1002 16485 -968
rect 9767 -1017 9819 -1002
rect 9996 -1005 10048 -1002
rect 10215 -1015 10267 -1002
rect 10407 -1011 10459 -1002
rect 10901 -1013 10953 -1002
rect 12693 -1014 12745 -1002
rect 13086 -1016 13138 -1002
rect 13283 -1008 13335 -1002
rect 13613 -1006 13665 -1002
rect 13809 -1006 13861 -1002
rect 15716 -1013 15768 -1002
rect 16017 -1009 16069 -1002
rect 16223 -1008 16275 -1002
rect 16433 -1012 16485 -1002
rect 16644 -1006 16696 -954
rect 18524 -968 18576 -965
rect 18781 -968 18833 -958
rect 19031 -968 19083 -962
rect 19302 -968 19354 -957
rect 19543 -968 19595 -954
rect 19768 -968 19820 -958
rect 21475 -968 21527 -960
rect 21676 -968 21728 -959
rect 21894 -968 21946 -963
rect 22101 -968 22153 -959
rect 22306 -968 22358 -960
rect 22653 -968 22705 -964
rect 24405 -968 24457 -960
rect 24596 -968 24648 -957
rect 24791 -968 24843 -955
rect 25238 -968 25290 -960
rect 18524 -1002 18540 -968
rect 18540 -1002 18574 -968
rect 18574 -1002 18576 -968
rect 18781 -1002 18816 -968
rect 18816 -1002 18833 -968
rect 19031 -1002 19034 -968
rect 19034 -1002 19083 -968
rect 19302 -1002 19310 -968
rect 19310 -1002 19354 -968
rect 19543 -1002 19552 -968
rect 19552 -1002 19586 -968
rect 19586 -1002 19595 -968
rect 19768 -1002 19770 -968
rect 19770 -1002 19820 -968
rect 21475 -1002 21484 -968
rect 21484 -1002 21518 -968
rect 21518 -1002 21527 -968
rect 21676 -1002 21702 -968
rect 21702 -1002 21728 -968
rect 21894 -1002 21944 -968
rect 21944 -1002 21946 -968
rect 22101 -1002 22128 -968
rect 22128 -1002 22153 -968
rect 22306 -1002 22312 -968
rect 22312 -1002 22346 -968
rect 22346 -1002 22358 -968
rect 22653 -1002 22680 -968
rect 22680 -1002 22705 -968
rect 24405 -1002 24428 -968
rect 24428 -1002 24457 -968
rect 24596 -1002 24612 -968
rect 24612 -1002 24646 -968
rect 24646 -1002 24648 -968
rect 24791 -1002 24796 -968
rect 24796 -1002 24830 -968
rect 24830 -1002 24843 -968
rect 25238 -1002 25256 -968
rect 25256 -1002 25290 -968
rect 18524 -1017 18576 -1002
rect 18781 -1010 18833 -1002
rect 19031 -1014 19083 -1002
rect 19302 -1009 19354 -1002
rect 19543 -1006 19595 -1002
rect 19768 -1010 19820 -1002
rect 21475 -1012 21527 -1002
rect 21676 -1011 21728 -1002
rect 21894 -1015 21946 -1002
rect 22101 -1011 22153 -1002
rect 22306 -1012 22358 -1002
rect 22653 -1016 22705 -1002
rect 24405 -1012 24457 -1002
rect 24596 -1009 24648 -1002
rect 24791 -1007 24843 -1002
rect 25238 -1012 25290 -1002
rect 8622 -1113 8674 -1109
rect 9070 -1113 9122 -1106
rect 8622 -1147 8638 -1113
rect 8638 -1147 8674 -1113
rect 8855 -1147 8880 -1113
rect 8880 -1147 8907 -1113
rect 9070 -1147 9098 -1113
rect 9098 -1147 9122 -1113
rect 8622 -1161 8674 -1147
rect 8855 -1165 8907 -1147
rect 9070 -1158 9122 -1147
rect 9288 -1161 9340 -1109
rect 9504 -1113 9556 -1108
rect 11225 -1113 11277 -1112
rect 11415 -1113 11467 -1112
rect 11625 -1113 11677 -1109
rect 11842 -1113 11894 -1112
rect 9504 -1147 9524 -1113
rect 9524 -1147 9556 -1113
rect 11225 -1147 11272 -1113
rect 11272 -1147 11277 -1113
rect 11415 -1147 11456 -1113
rect 11456 -1147 11467 -1113
rect 11625 -1147 11640 -1113
rect 11640 -1147 11674 -1113
rect 11674 -1147 11677 -1113
rect 11842 -1147 11858 -1113
rect 11858 -1147 11894 -1113
rect 9504 -1160 9556 -1147
rect 11225 -1164 11277 -1147
rect 11415 -1164 11467 -1147
rect 11625 -1161 11677 -1147
rect 11842 -1164 11894 -1147
rect 12137 -1161 12189 -1109
rect 12361 -1113 12413 -1104
rect 14239 -1113 14291 -1111
rect 14791 -1113 14843 -1109
rect 15008 -1113 15060 -1104
rect 15209 -1113 15261 -1107
rect 18104 -1113 18156 -1108
rect 20005 -1113 20057 -1112
rect 20261 -1113 20313 -1112
rect 20496 -1113 20548 -1112
rect 12361 -1147 12376 -1113
rect 12376 -1147 12410 -1113
rect 12410 -1147 12413 -1113
rect 14239 -1147 14250 -1113
rect 14250 -1147 14291 -1113
rect 14539 -1147 14584 -1113
rect 14584 -1147 14591 -1113
rect 14791 -1147 14802 -1113
rect 14802 -1147 14843 -1113
rect 15008 -1147 15044 -1113
rect 15044 -1147 15060 -1113
rect 15209 -1147 15228 -1113
rect 15228 -1147 15261 -1113
rect 17094 -1147 17102 -1116
rect 17102 -1147 17146 -1116
rect 12361 -1156 12413 -1147
rect 14239 -1163 14291 -1147
rect 14539 -1165 14591 -1147
rect 14791 -1161 14843 -1147
rect 15008 -1156 15060 -1147
rect 15209 -1159 15261 -1147
rect 17094 -1168 17146 -1147
rect 17286 -1168 17338 -1116
rect 17486 -1147 17528 -1116
rect 17528 -1147 17538 -1116
rect 18104 -1147 18114 -1113
rect 18114 -1147 18156 -1113
rect 20005 -1147 20012 -1113
rect 20012 -1147 20046 -1113
rect 20046 -1147 20057 -1113
rect 20261 -1147 20288 -1113
rect 20288 -1147 20313 -1113
rect 20496 -1147 20506 -1113
rect 20506 -1147 20548 -1113
rect 17486 -1168 17538 -1147
rect 18104 -1160 18156 -1147
rect 20005 -1164 20057 -1147
rect 20261 -1164 20313 -1147
rect 20496 -1164 20548 -1147
rect 20785 -1162 20837 -1110
rect 20975 -1113 21027 -1112
rect 21179 -1113 21231 -1110
rect 22965 -1113 23017 -1104
rect 23207 -1113 23259 -1108
rect 23407 -1113 23459 -1109
rect 23597 -1113 23649 -1101
rect 20975 -1147 21024 -1113
rect 21024 -1147 21027 -1113
rect 21179 -1147 21208 -1113
rect 21208 -1147 21231 -1113
rect 22965 -1147 22990 -1113
rect 22990 -1147 23017 -1113
rect 23207 -1147 23232 -1113
rect 23232 -1147 23259 -1113
rect 23407 -1147 23416 -1113
rect 23416 -1147 23450 -1113
rect 23450 -1147 23459 -1113
rect 23597 -1147 23600 -1113
rect 23600 -1147 23634 -1113
rect 23634 -1147 23649 -1113
rect 20975 -1164 21027 -1147
rect 21179 -1162 21231 -1147
rect 22965 -1156 23017 -1147
rect 23207 -1160 23259 -1147
rect 23407 -1161 23459 -1147
rect 23597 -1153 23649 -1147
rect 23818 -1155 23870 -1103
rect 24114 -1113 24166 -1108
rect 24114 -1147 24152 -1113
rect 24152 -1147 24166 -1113
rect 24114 -1160 24166 -1147
rect 8592 -1223 8644 -1215
rect 8592 -1257 8601 -1223
rect 8601 -1257 8635 -1223
rect 8635 -1257 8644 -1223
rect 10984 -1223 11036 -1215
rect 8592 -1267 8644 -1257
rect 8872 -1289 8924 -1279
rect 8872 -1323 8881 -1289
rect 8881 -1323 8915 -1289
rect 8915 -1323 8924 -1289
rect 8872 -1331 8924 -1323
rect 9600 -1303 9652 -1251
rect 10984 -1257 10993 -1223
rect 10993 -1257 11027 -1223
rect 11027 -1257 11036 -1223
rect 13377 -1223 13429 -1215
rect 10984 -1267 11036 -1257
rect 11264 -1289 11316 -1279
rect 11264 -1323 11273 -1289
rect 11273 -1323 11307 -1289
rect 11307 -1323 11316 -1289
rect 11264 -1331 11316 -1323
rect 10879 -1360 10933 -1350
rect 10879 -1394 10889 -1360
rect 10889 -1394 10923 -1360
rect 10923 -1394 10933 -1360
rect 10879 -1402 10933 -1394
rect 10534 -1416 10586 -1405
rect 10534 -1450 10543 -1416
rect 10543 -1450 10577 -1416
rect 10577 -1450 10586 -1416
rect 10534 -1458 10586 -1450
rect 11992 -1302 12044 -1250
rect 13377 -1257 13386 -1223
rect 13386 -1257 13420 -1223
rect 13420 -1257 13429 -1223
rect 15768 -1223 15820 -1215
rect 13377 -1267 13429 -1257
rect 13655 -1289 13707 -1279
rect 13655 -1323 13664 -1289
rect 13664 -1323 13698 -1289
rect 13698 -1323 13707 -1289
rect 13655 -1331 13707 -1323
rect 13273 -1360 13327 -1350
rect 13273 -1394 13283 -1360
rect 13283 -1394 13317 -1360
rect 13317 -1394 13327 -1360
rect 13273 -1402 13327 -1394
rect 12926 -1416 12978 -1405
rect 12926 -1450 12935 -1416
rect 12935 -1450 12969 -1416
rect 12969 -1450 12978 -1416
rect 12926 -1458 12978 -1450
rect 14384 -1303 14436 -1251
rect 15768 -1257 15777 -1223
rect 15777 -1257 15811 -1223
rect 15811 -1257 15820 -1223
rect 18160 -1224 18212 -1216
rect 15768 -1267 15820 -1257
rect 16048 -1289 16100 -1279
rect 16048 -1323 16057 -1289
rect 16057 -1323 16091 -1289
rect 16091 -1323 16100 -1289
rect 16048 -1331 16100 -1323
rect 15663 -1358 15717 -1348
rect 15663 -1392 15673 -1358
rect 15673 -1392 15707 -1358
rect 15707 -1392 15717 -1358
rect 15663 -1400 15717 -1392
rect 15317 -1415 15369 -1405
rect 15317 -1449 15326 -1415
rect 15326 -1449 15360 -1415
rect 15360 -1449 15369 -1415
rect 15317 -1457 15369 -1449
rect 16776 -1303 16828 -1251
rect 18160 -1258 18169 -1224
rect 18169 -1258 18203 -1224
rect 18203 -1258 18212 -1224
rect 20553 -1222 20605 -1214
rect 18160 -1268 18212 -1258
rect 18440 -1289 18492 -1279
rect 18440 -1323 18449 -1289
rect 18449 -1323 18483 -1289
rect 18483 -1323 18492 -1289
rect 18440 -1331 18492 -1323
rect 18055 -1360 18109 -1350
rect 18055 -1394 18065 -1360
rect 18065 -1394 18099 -1360
rect 18099 -1394 18109 -1360
rect 18055 -1402 18109 -1394
rect 17710 -1416 17762 -1405
rect 17710 -1450 17719 -1416
rect 17719 -1450 17753 -1416
rect 17753 -1450 17762 -1416
rect 17710 -1458 17762 -1450
rect 19168 -1303 19220 -1251
rect 20553 -1256 20562 -1222
rect 20562 -1256 20596 -1222
rect 20596 -1256 20605 -1222
rect 22944 -1222 22996 -1214
rect 20553 -1266 20605 -1256
rect 20831 -1288 20883 -1278
rect 20831 -1322 20840 -1288
rect 20840 -1322 20874 -1288
rect 20874 -1322 20883 -1288
rect 20831 -1330 20883 -1322
rect 20447 -1358 20501 -1348
rect 20447 -1392 20457 -1358
rect 20457 -1392 20491 -1358
rect 20491 -1392 20501 -1358
rect 20447 -1400 20501 -1392
rect 20101 -1416 20153 -1405
rect 20101 -1450 20110 -1416
rect 20110 -1450 20144 -1416
rect 20144 -1450 20153 -1416
rect 20101 -1458 20153 -1450
rect 21560 -1302 21612 -1250
rect 22944 -1256 22953 -1222
rect 22953 -1256 22987 -1222
rect 22987 -1256 22996 -1222
rect 22944 -1266 22996 -1256
rect 23224 -1289 23276 -1279
rect 23224 -1323 23233 -1289
rect 23233 -1323 23267 -1289
rect 23267 -1323 23276 -1289
rect 23224 -1331 23276 -1323
rect 22839 -1360 22893 -1350
rect 22839 -1394 22849 -1360
rect 22849 -1394 22883 -1360
rect 22883 -1394 22893 -1360
rect 22839 -1402 22893 -1394
rect 22494 -1416 22546 -1405
rect 22494 -1450 22503 -1416
rect 22503 -1450 22537 -1416
rect 22537 -1450 22546 -1416
rect 22494 -1458 22546 -1450
rect 23952 -1302 24004 -1250
rect 25231 -1358 25285 -1348
rect 25231 -1392 25241 -1358
rect 25241 -1392 25275 -1358
rect 25275 -1392 25285 -1358
rect 25231 -1400 25285 -1392
rect 24887 -1416 24939 -1405
rect 24887 -1450 24896 -1416
rect 24896 -1450 24930 -1416
rect 24930 -1450 24939 -1416
rect 24887 -1458 24939 -1450
rect 8996 -1657 9048 -1641
rect 8996 -1691 9006 -1657
rect 9006 -1691 9048 -1657
rect 8996 -1693 9048 -1691
rect 9195 -1696 9247 -1644
rect 9406 -1657 9458 -1644
rect 9612 -1657 9664 -1644
rect 9406 -1691 9432 -1657
rect 9432 -1691 9458 -1657
rect 9612 -1691 9616 -1657
rect 9616 -1691 9650 -1657
rect 9650 -1691 9664 -1657
rect 9406 -1696 9458 -1691
rect 9612 -1696 9664 -1691
rect 9840 -1698 9892 -1646
rect 10084 -1657 10136 -1646
rect 10314 -1657 10366 -1644
rect 10520 -1657 10572 -1644
rect 10738 -1657 10790 -1639
rect 10084 -1691 10110 -1657
rect 10110 -1691 10136 -1657
rect 10314 -1691 10352 -1657
rect 10352 -1691 10366 -1657
rect 10520 -1691 10536 -1657
rect 10536 -1691 10570 -1657
rect 10570 -1691 10572 -1657
rect 10738 -1691 10754 -1657
rect 10754 -1691 10790 -1657
rect 10084 -1698 10136 -1691
rect 10314 -1696 10366 -1691
rect 10520 -1696 10572 -1691
rect 10941 -1697 10993 -1645
rect 11149 -1657 11201 -1642
rect 11412 -1657 11464 -1646
rect 11620 -1657 11672 -1645
rect 11830 -1657 11882 -1648
rect 12030 -1657 12082 -1642
rect 12233 -1657 12285 -1645
rect 12443 -1657 12495 -1645
rect 12644 -1657 12696 -1644
rect 12860 -1657 12912 -1643
rect 13141 -1657 13193 -1645
rect 13361 -1657 13413 -1650
rect 13566 -1657 13618 -1649
rect 13787 -1657 13839 -1643
rect 13992 -1657 14044 -1650
rect 14201 -1657 14253 -1649
rect 14418 -1657 14470 -1649
rect 14632 -1657 14684 -1644
rect 14827 -1657 14879 -1646
rect 15022 -1657 15074 -1649
rect 15224 -1657 15276 -1646
rect 15508 -1657 15560 -1645
rect 15707 -1657 15759 -1644
rect 11149 -1691 11180 -1657
rect 11180 -1691 11201 -1657
rect 11412 -1691 11456 -1657
rect 11456 -1691 11464 -1657
rect 11620 -1691 11640 -1657
rect 11640 -1691 11672 -1657
rect 11830 -1691 11858 -1657
rect 11858 -1691 11882 -1657
rect 12030 -1691 12042 -1657
rect 12042 -1691 12082 -1657
rect 12233 -1691 12284 -1657
rect 12284 -1691 12285 -1657
rect 12443 -1691 12468 -1657
rect 12468 -1691 12495 -1657
rect 12644 -1691 12652 -1657
rect 12652 -1691 12686 -1657
rect 12686 -1691 12696 -1657
rect 12860 -1691 12870 -1657
rect 12870 -1691 12912 -1657
rect 13141 -1691 13146 -1657
rect 13146 -1691 13193 -1657
rect 13361 -1691 13388 -1657
rect 13388 -1691 13413 -1657
rect 13566 -1691 13572 -1657
rect 13572 -1691 13606 -1657
rect 13606 -1691 13618 -1657
rect 13787 -1691 13790 -1657
rect 13790 -1691 13839 -1657
rect 13992 -1691 14032 -1657
rect 14032 -1691 14044 -1657
rect 14201 -1691 14216 -1657
rect 14216 -1691 14250 -1657
rect 14250 -1691 14253 -1657
rect 14418 -1691 14434 -1657
rect 14434 -1691 14470 -1657
rect 14632 -1691 14676 -1657
rect 14676 -1691 14684 -1657
rect 14827 -1691 14860 -1657
rect 14860 -1691 14879 -1657
rect 15022 -1691 15044 -1657
rect 15044 -1691 15074 -1657
rect 15224 -1691 15228 -1657
rect 15228 -1691 15262 -1657
rect 15262 -1691 15276 -1657
rect 15508 -1691 15538 -1657
rect 15538 -1691 15560 -1657
rect 15707 -1691 15722 -1657
rect 15722 -1691 15759 -1657
rect 11149 -1694 11201 -1691
rect 11412 -1698 11464 -1691
rect 11620 -1697 11672 -1691
rect 11830 -1700 11882 -1691
rect 12030 -1694 12082 -1691
rect 12233 -1697 12285 -1691
rect 12443 -1697 12495 -1691
rect 12644 -1696 12696 -1691
rect 12860 -1695 12912 -1691
rect 13141 -1697 13193 -1691
rect 13361 -1702 13413 -1691
rect 13566 -1701 13618 -1691
rect 13787 -1695 13839 -1691
rect 13992 -1702 14044 -1691
rect 14201 -1701 14253 -1691
rect 14418 -1701 14470 -1691
rect 14632 -1696 14684 -1691
rect 14827 -1698 14879 -1691
rect 15022 -1701 15074 -1691
rect 15224 -1698 15276 -1691
rect 15508 -1697 15560 -1691
rect 15707 -1696 15759 -1691
rect 15910 -1694 15962 -1642
rect 16175 -1657 16227 -1645
rect 16373 -1657 16425 -1646
rect 16562 -1657 16614 -1644
rect 16774 -1657 16826 -1644
rect 16991 -1657 17043 -1644
rect 16175 -1691 16182 -1657
rect 16182 -1691 16227 -1657
rect 16373 -1691 16424 -1657
rect 16424 -1691 16425 -1657
rect 16562 -1691 16608 -1657
rect 16608 -1691 16614 -1657
rect 16774 -1691 16792 -1657
rect 16792 -1691 16826 -1657
rect 16991 -1691 17010 -1657
rect 17010 -1691 17043 -1657
rect 16175 -1697 16227 -1691
rect 16373 -1698 16425 -1691
rect 16562 -1696 16614 -1691
rect 16774 -1696 16826 -1691
rect 16991 -1696 17043 -1691
rect 17196 -1700 17248 -1648
rect 17401 -1657 17453 -1648
rect 17609 -1657 17661 -1643
rect 17892 -1657 17944 -1644
rect 18085 -1657 18137 -1646
rect 18311 -1657 18363 -1648
rect 17401 -1691 17436 -1657
rect 17436 -1691 17453 -1657
rect 17609 -1691 17620 -1657
rect 17620 -1691 17654 -1657
rect 17654 -1691 17661 -1657
rect 17892 -1691 17896 -1657
rect 17896 -1691 17930 -1657
rect 17930 -1691 17944 -1657
rect 18085 -1691 18114 -1657
rect 18114 -1691 18137 -1657
rect 18311 -1691 18356 -1657
rect 18356 -1691 18363 -1657
rect 17401 -1700 17453 -1691
rect 17609 -1695 17661 -1691
rect 17892 -1696 17944 -1691
rect 18085 -1698 18137 -1691
rect 18311 -1700 18363 -1691
rect 18576 -1700 18628 -1648
rect 18770 -1657 18822 -1644
rect 18968 -1657 19020 -1653
rect 19172 -1657 19224 -1645
rect 19392 -1657 19444 -1642
rect 19607 -1657 19659 -1646
rect 19835 -1657 19887 -1643
rect 20039 -1657 20091 -1646
rect 20277 -1657 20329 -1644
rect 20470 -1657 20522 -1643
rect 20667 -1657 20719 -1648
rect 20923 -1657 20975 -1645
rect 21162 -1657 21214 -1649
rect 21395 -1657 21447 -1653
rect 18770 -1691 18816 -1657
rect 18816 -1691 18822 -1657
rect 18968 -1691 19000 -1657
rect 19000 -1691 19020 -1657
rect 19172 -1691 19184 -1657
rect 19184 -1691 19218 -1657
rect 19218 -1691 19224 -1657
rect 19392 -1691 19402 -1657
rect 19402 -1691 19444 -1657
rect 19607 -1691 19644 -1657
rect 19644 -1691 19659 -1657
rect 19835 -1691 19862 -1657
rect 19862 -1691 19887 -1657
rect 20039 -1691 20046 -1657
rect 20046 -1691 20091 -1657
rect 20277 -1691 20288 -1657
rect 20288 -1691 20322 -1657
rect 20322 -1691 20329 -1657
rect 20470 -1691 20472 -1657
rect 20472 -1691 20506 -1657
rect 20506 -1691 20522 -1657
rect 20667 -1691 20690 -1657
rect 20690 -1691 20719 -1657
rect 20923 -1691 20932 -1657
rect 20932 -1691 20966 -1657
rect 20966 -1691 20975 -1657
rect 21162 -1691 21208 -1657
rect 21208 -1691 21214 -1657
rect 21395 -1691 21426 -1657
rect 21426 -1691 21447 -1657
rect 18770 -1696 18822 -1691
rect 18968 -1705 19020 -1691
rect 19172 -1697 19224 -1691
rect 19392 -1694 19444 -1691
rect 19607 -1698 19659 -1691
rect 19835 -1695 19887 -1691
rect 20039 -1698 20091 -1691
rect 20277 -1696 20329 -1691
rect 20470 -1695 20522 -1691
rect 20667 -1700 20719 -1691
rect 20923 -1697 20975 -1691
rect 21162 -1701 21214 -1691
rect 21395 -1705 21447 -1691
rect 21616 -1700 21668 -1648
rect 21807 -1657 21859 -1648
rect 22035 -1657 22087 -1646
rect 22232 -1657 22284 -1651
rect 21807 -1691 21852 -1657
rect 21852 -1691 21859 -1657
rect 22035 -1691 22036 -1657
rect 22036 -1691 22070 -1657
rect 22070 -1691 22087 -1657
rect 22232 -1691 22254 -1657
rect 22254 -1691 22284 -1657
rect 21807 -1700 21859 -1691
rect 22035 -1698 22087 -1691
rect 22232 -1703 22284 -1691
rect 22444 -1703 22496 -1651
rect 22671 -1657 22723 -1648
rect 22860 -1657 22912 -1647
rect 22671 -1691 22680 -1657
rect 22680 -1691 22714 -1657
rect 22714 -1691 22723 -1657
rect 22860 -1691 22864 -1657
rect 22864 -1691 22898 -1657
rect 22898 -1691 22912 -1657
rect 22671 -1700 22723 -1691
rect 22860 -1699 22912 -1691
rect 23086 -1698 23138 -1646
rect 23340 -1657 23392 -1646
rect 23584 -1657 23636 -1649
rect 23814 -1657 23866 -1650
rect 24072 -1657 24124 -1647
rect 23340 -1691 23358 -1657
rect 23358 -1691 23392 -1657
rect 23584 -1691 23600 -1657
rect 23600 -1691 23634 -1657
rect 23634 -1691 23636 -1657
rect 23814 -1691 23818 -1657
rect 23818 -1691 23866 -1657
rect 24072 -1691 24094 -1657
rect 24094 -1691 24124 -1657
rect 23340 -1698 23392 -1691
rect 23584 -1701 23636 -1691
rect 23814 -1702 23866 -1691
rect 24072 -1699 24124 -1691
rect 24282 -1699 24334 -1647
rect 24507 -1657 24559 -1647
rect 24726 -1657 24778 -1650
rect 25072 -1657 25124 -1646
rect 25271 -1657 25323 -1649
rect 24507 -1691 24520 -1657
rect 24520 -1691 24554 -1657
rect 24554 -1691 24559 -1657
rect 24726 -1691 24738 -1657
rect 24738 -1691 24778 -1657
rect 25072 -1691 25106 -1657
rect 25106 -1691 25124 -1657
rect 25271 -1691 25290 -1657
rect 25290 -1691 25323 -1657
rect 24507 -1699 24559 -1691
rect 24726 -1702 24778 -1691
rect 25072 -1698 25124 -1691
rect 25271 -1701 25323 -1691
<< metal2 >>
rect 13945 13628 14019 13632
rect 13945 13572 13954 13628
rect 14010 13623 14019 13628
rect 20654 13628 20728 13632
rect 14010 13619 14616 13623
rect 14010 13572 14050 13619
rect 13945 13568 14050 13572
rect 13946 13563 14050 13568
rect 14106 13563 14130 13619
rect 14186 13563 14210 13619
rect 14266 13563 14290 13619
rect 14346 13563 14370 13619
rect 14426 13563 14450 13619
rect 14506 13563 14616 13619
rect 13946 13557 14616 13563
rect 14678 13622 19586 13626
rect 14678 13566 14782 13622
rect 14838 13566 14862 13622
rect 14918 13566 14942 13622
rect 14998 13566 15022 13622
rect 15078 13566 15102 13622
rect 15158 13566 15182 13622
rect 15238 13566 15390 13622
rect 15446 13566 15470 13622
rect 15526 13566 15550 13622
rect 15606 13566 15630 13622
rect 15686 13566 15710 13622
rect 15766 13566 15790 13622
rect 15846 13566 15994 13622
rect 16050 13566 16074 13622
rect 16130 13566 16154 13622
rect 16210 13566 16234 13622
rect 16290 13566 16314 13622
rect 16370 13566 16394 13622
rect 16450 13566 16602 13622
rect 16658 13566 16682 13622
rect 16738 13566 16762 13622
rect 16818 13566 16842 13622
rect 16898 13566 16922 13622
rect 16978 13566 17002 13622
rect 17058 13566 17206 13622
rect 17262 13566 17286 13622
rect 17342 13566 17366 13622
rect 17422 13566 17446 13622
rect 17502 13566 17526 13622
rect 17582 13566 17606 13622
rect 17662 13566 17814 13622
rect 17870 13566 17894 13622
rect 17950 13566 17974 13622
rect 18030 13566 18054 13622
rect 18110 13566 18134 13622
rect 18190 13566 18214 13622
rect 18270 13566 18418 13622
rect 18474 13566 18498 13622
rect 18554 13566 18578 13622
rect 18634 13566 18658 13622
rect 18714 13566 18738 13622
rect 18794 13566 18818 13622
rect 18874 13566 19026 13622
rect 19082 13566 19106 13622
rect 19162 13566 19186 13622
rect 19242 13566 19266 13622
rect 19322 13566 19346 13622
rect 19402 13566 19426 13622
rect 19482 13566 19586 13622
rect 14678 13560 19586 13566
rect 19754 13566 19828 13570
rect 19754 13510 19763 13566
rect 19819 13510 19828 13566
rect 19754 13506 19828 13510
rect 20231 13569 20305 13573
rect 20231 13513 20240 13569
rect 20296 13513 20305 13569
rect 20654 13572 20663 13628
rect 20719 13623 20728 13628
rect 20719 13619 21325 13623
rect 20719 13572 20759 13619
rect 20654 13568 20759 13572
rect 20655 13563 20759 13568
rect 20815 13563 20839 13619
rect 20895 13563 20919 13619
rect 20975 13563 20999 13619
rect 21055 13563 21079 13619
rect 21135 13563 21159 13619
rect 21215 13563 21325 13619
rect 20655 13557 21325 13563
rect 21387 13622 26295 13626
rect 21387 13566 21491 13622
rect 21547 13566 21571 13622
rect 21627 13566 21651 13622
rect 21707 13566 21731 13622
rect 21787 13566 21811 13622
rect 21867 13566 21891 13622
rect 21947 13566 22099 13622
rect 22155 13566 22179 13622
rect 22235 13566 22259 13622
rect 22315 13566 22339 13622
rect 22395 13566 22419 13622
rect 22475 13566 22499 13622
rect 22555 13566 22703 13622
rect 22759 13566 22783 13622
rect 22839 13566 22863 13622
rect 22919 13566 22943 13622
rect 22999 13566 23023 13622
rect 23079 13566 23103 13622
rect 23159 13566 23311 13622
rect 23367 13566 23391 13622
rect 23447 13566 23471 13622
rect 23527 13566 23551 13622
rect 23607 13566 23631 13622
rect 23687 13566 23711 13622
rect 23767 13566 23915 13622
rect 23971 13566 23995 13622
rect 24051 13566 24075 13622
rect 24131 13566 24155 13622
rect 24211 13566 24235 13622
rect 24291 13566 24315 13622
rect 24371 13566 24523 13622
rect 24579 13566 24603 13622
rect 24659 13566 24683 13622
rect 24739 13566 24763 13622
rect 24819 13566 24843 13622
rect 24899 13566 24923 13622
rect 24979 13566 25127 13622
rect 25183 13566 25207 13622
rect 25263 13566 25287 13622
rect 25343 13566 25367 13622
rect 25423 13566 25447 13622
rect 25503 13566 25527 13622
rect 25583 13566 25735 13622
rect 25791 13566 25815 13622
rect 25871 13566 25895 13622
rect 25951 13566 25975 13622
rect 26031 13566 26055 13622
rect 26111 13566 26135 13622
rect 26191 13566 26295 13622
rect 21387 13560 26295 13566
rect 26463 13566 26537 13570
rect 20231 13509 20305 13513
rect 26463 13510 26472 13566
rect 26528 13510 26537 13566
rect 26463 13506 26537 13510
rect 19759 13422 19833 13426
rect 19759 13366 19768 13422
rect 19824 13366 19833 13422
rect 26468 13422 26542 13426
rect 19759 13362 19833 13366
rect 20220 13397 20294 13401
rect 3057 13153 3131 13157
rect 3057 13097 3066 13153
rect 3122 13148 3131 13153
rect 3356 13148 3390 13362
rect 20220 13341 20229 13397
rect 20285 13341 20294 13397
rect 26468 13366 26477 13422
rect 26533 13366 26542 13422
rect 26468 13362 26542 13366
rect 20220 13337 20294 13341
rect 19760 13270 19834 13274
rect 19760 13214 19769 13270
rect 19825 13214 19834 13270
rect 19760 13210 19834 13214
rect 26469 13270 26543 13274
rect 26469 13214 26478 13270
rect 26534 13214 26543 13270
rect 26469 13210 26543 13214
rect 20220 13205 20294 13209
rect 3122 13144 3728 13148
rect 3122 13097 3162 13144
rect 3057 13093 3162 13097
rect 3058 13088 3162 13093
rect 3218 13088 3242 13144
rect 3298 13088 3322 13144
rect 3378 13088 3402 13144
rect 3458 13088 3482 13144
rect 3538 13088 3562 13144
rect 3618 13088 3728 13144
rect 3058 13082 3728 13088
rect 3790 13147 8698 13151
rect 3790 13091 3894 13147
rect 3950 13091 3974 13147
rect 4030 13091 4054 13147
rect 4110 13091 4134 13147
rect 4190 13091 4214 13147
rect 4270 13091 4294 13147
rect 4350 13091 4502 13147
rect 4558 13091 4582 13147
rect 4638 13091 4662 13147
rect 4718 13091 4742 13147
rect 4798 13091 4822 13147
rect 4878 13091 4902 13147
rect 4958 13091 5106 13147
rect 5162 13091 5186 13147
rect 5242 13091 5266 13147
rect 5322 13091 5346 13147
rect 5402 13091 5426 13147
rect 5482 13091 5506 13147
rect 5562 13091 5714 13147
rect 5770 13091 5794 13147
rect 5850 13091 5874 13147
rect 5930 13091 5954 13147
rect 6010 13091 6034 13147
rect 6090 13091 6114 13147
rect 6170 13091 6318 13147
rect 6374 13091 6398 13147
rect 6454 13091 6478 13147
rect 6534 13091 6558 13147
rect 6614 13091 6638 13147
rect 6694 13091 6718 13147
rect 6774 13091 6926 13147
rect 6982 13091 7006 13147
rect 7062 13091 7086 13147
rect 7142 13091 7166 13147
rect 7222 13091 7246 13147
rect 7302 13091 7326 13147
rect 7382 13091 7530 13147
rect 7586 13091 7610 13147
rect 7666 13091 7690 13147
rect 7746 13091 7770 13147
rect 7826 13091 7850 13147
rect 7906 13091 7930 13147
rect 7986 13091 8138 13147
rect 8194 13091 8218 13147
rect 8274 13091 8298 13147
rect 8354 13091 8378 13147
rect 8434 13091 8458 13147
rect 8514 13091 8538 13147
rect 8594 13091 8698 13147
rect 20220 13149 20229 13205
rect 20285 13149 20294 13205
rect 20220 13145 20294 13149
rect 19760 13100 19834 13104
rect 3790 13085 8698 13091
rect 8866 13091 8940 13095
rect 2449 12548 2505 12557
rect 2449 12483 2505 12492
rect 2580 12547 2636 12556
rect 2580 12482 2636 12491
rect 2724 12548 2780 12557
rect 2724 12483 2780 12492
rect 3356 12297 3390 13082
rect 8866 13035 8875 13091
rect 8931 13035 8940 13091
rect 19760 13044 19769 13100
rect 19825 13044 19834 13100
rect 19760 13040 19834 13044
rect 26469 13100 26543 13104
rect 26469 13044 26478 13100
rect 26534 13044 26543 13100
rect 26469 13040 26543 13044
rect 8866 13031 8940 13035
rect 13337 13023 13393 13032
rect 13337 12958 13393 12967
rect 13468 13022 13524 13031
rect 13468 12957 13524 12966
rect 13612 13023 13668 13032
rect 13612 12958 13668 12967
rect 20046 13023 20102 13032
rect 20046 12958 20102 12967
rect 20177 13022 20233 13031
rect 20177 12957 20233 12966
rect 20321 13023 20377 13032
rect 20321 12958 20377 12967
rect 8871 12947 8945 12951
rect 8871 12891 8880 12947
rect 8936 12891 8945 12947
rect 8871 12887 8945 12891
rect 19759 12943 19833 12947
rect 19759 12887 19768 12943
rect 19824 12887 19833 12943
rect 19759 12883 19833 12887
rect 26468 12943 26542 12947
rect 26468 12887 26477 12943
rect 26533 12887 26542 12943
rect 26468 12883 26542 12887
rect 8872 12795 8946 12799
rect 8872 12739 8881 12795
rect 8937 12739 8946 12795
rect 8872 12735 8946 12739
rect 13604 12658 13612 12710
rect 13664 12658 13670 12710
rect 13604 12657 13670 12658
rect 19677 12701 19751 12705
rect 8872 12625 8946 12629
rect 8872 12569 8881 12625
rect 8937 12569 8946 12625
rect 13622 12581 13668 12657
rect 19677 12645 19686 12701
rect 19742 12645 19751 12701
rect 20313 12658 20321 12710
rect 20373 12658 20379 12710
rect 20313 12657 20379 12658
rect 26386 12701 26460 12705
rect 19677 12641 19751 12645
rect 20331 12581 20377 12657
rect 26386 12645 26395 12701
rect 26451 12645 26460 12701
rect 26386 12641 26460 12645
rect 8872 12565 8946 12569
rect 10976 12556 11050 12560
rect 10976 12500 10985 12556
rect 11041 12500 11050 12556
rect 10976 12496 11050 12500
rect 11163 12558 11237 12562
rect 11163 12502 11172 12558
rect 11228 12502 11237 12558
rect 11163 12498 11237 12502
rect 11348 12560 11422 12564
rect 11348 12504 11357 12560
rect 11413 12504 11422 12560
rect 11348 12500 11422 12504
rect 11533 12561 11607 12565
rect 11533 12505 11542 12561
rect 11598 12505 11607 12561
rect 11533 12501 11607 12505
rect 11736 12563 11810 12567
rect 11736 12507 11745 12563
rect 11801 12507 11810 12563
rect 11736 12503 11810 12507
rect 11921 12565 11995 12569
rect 11921 12509 11930 12565
rect 11986 12509 11995 12565
rect 11921 12505 11995 12509
rect 12120 12567 12194 12571
rect 12120 12511 12129 12567
rect 12185 12511 12194 12567
rect 12120 12507 12194 12511
rect 12322 12566 12396 12570
rect 12322 12510 12331 12566
rect 12387 12510 12396 12566
rect 12322 12506 12396 12510
rect 12532 12569 12606 12573
rect 12532 12513 12541 12569
rect 12597 12513 12606 12569
rect 12532 12509 12606 12513
rect 12756 12569 12830 12573
rect 12756 12513 12765 12569
rect 12821 12513 12830 12569
rect 12756 12509 12830 12513
rect 12962 12568 13036 12572
rect 12962 12512 12971 12568
rect 13027 12512 13036 12568
rect 12962 12508 13036 12512
rect 13183 12567 13257 12571
rect 13183 12511 13192 12567
rect 13248 12511 13257 12567
rect 13622 12535 13861 12581
rect 20331 12535 20570 12581
rect 13183 12507 13257 12511
rect 13355 12477 13411 12486
rect 8871 12468 8945 12472
rect 8871 12412 8880 12468
rect 8936 12412 8945 12468
rect 13355 12412 13411 12421
rect 13475 12477 13531 12486
rect 13475 12412 13531 12421
rect 13618 12477 13674 12486
rect 13618 12412 13674 12421
rect 8871 12408 8945 12412
rect 11632 12311 11696 12312
rect 9166 12278 9240 12282
rect 2716 12183 2724 12235
rect 2776 12183 2782 12235
rect 2716 12182 2782 12183
rect 8789 12226 8863 12230
rect 2734 12106 2780 12182
rect 8789 12170 8798 12226
rect 8854 12170 8863 12226
rect 9166 12222 9175 12278
rect 9231 12222 9240 12278
rect 11632 12259 11638 12311
rect 11690 12259 11696 12311
rect 9166 12218 9240 12222
rect 8789 12166 8863 12170
rect 11248 12145 11256 12197
rect 11308 12145 11314 12197
rect 2734 12060 2973 12106
rect 2467 12002 2523 12011
rect 2467 11937 2523 11946
rect 2587 12002 2643 12011
rect 2587 11937 2643 11946
rect 2730 12002 2786 12011
rect 2730 11937 2786 11946
rect 2730 11657 2795 11658
rect 2730 11605 2736 11657
rect 2788 11654 2795 11657
rect 2927 11654 2973 12060
rect 11274 12033 11305 12145
rect 11258 11981 11264 12033
rect 11317 11981 11324 12033
rect 4273 11967 4352 11968
rect 4500 11967 4579 11968
rect 5485 11967 5564 11968
rect 5712 11967 5791 11968
rect 6697 11967 6776 11968
rect 6924 11967 7003 11968
rect 7909 11967 7988 11968
rect 8136 11967 8215 11968
rect 3541 11964 3620 11965
rect 3538 11900 3548 11964
rect 3612 11900 3621 11964
rect 4270 11903 4280 11967
rect 4344 11903 4353 11967
rect 4499 11903 4508 11967
rect 4572 11903 4582 11967
rect 5482 11903 5492 11967
rect 5556 11903 5565 11967
rect 5711 11903 5720 11967
rect 5784 11903 5794 11967
rect 6694 11903 6704 11967
rect 6768 11903 6777 11967
rect 6923 11903 6932 11967
rect 6996 11903 7006 11967
rect 7906 11903 7916 11967
rect 7980 11903 7989 11967
rect 8135 11903 8144 11967
rect 8208 11903 8218 11967
rect 8877 11965 8951 11969
rect 8877 11909 8886 11965
rect 8942 11909 8951 11965
rect 8877 11905 8951 11909
rect 10906 11883 10981 11887
rect 10291 11808 10298 11862
rect 10352 11808 10359 11862
rect 10906 11827 10916 11883
rect 10972 11827 10981 11883
rect 11106 11886 11181 11890
rect 11106 11830 11116 11886
rect 11172 11830 11181 11886
rect 11106 11829 11181 11830
rect 11342 11884 11417 11888
rect 11342 11828 11352 11884
rect 11408 11828 11417 11884
rect 11342 11827 11417 11828
rect 10906 11826 10981 11827
rect 3895 11701 3904 11765
rect 3968 11701 3977 11765
rect 3895 11700 3977 11701
rect 4627 11701 4636 11765
rect 4700 11701 4709 11765
rect 4627 11700 4709 11701
rect 4845 11701 4854 11765
rect 4918 11701 4927 11765
rect 4845 11700 4927 11701
rect 5839 11701 5848 11765
rect 5912 11701 5921 11765
rect 5839 11700 5921 11701
rect 6057 11701 6066 11765
rect 6130 11701 6139 11765
rect 6057 11700 6139 11701
rect 7177 11701 7186 11765
rect 7250 11701 7259 11765
rect 7177 11700 7259 11701
rect 7395 11701 7404 11765
rect 7468 11701 7477 11765
rect 7395 11700 7477 11701
rect 8129 11701 8138 11765
rect 8202 11701 8211 11765
rect 8877 11762 8951 11766
rect 8877 11706 8886 11762
rect 8942 11706 8951 11762
rect 8877 11702 8951 11706
rect 8129 11700 8211 11701
rect 3217 11654 3224 11657
rect 2788 11608 3224 11654
rect 2788 11605 2795 11608
rect 3217 11605 3224 11608
rect 3276 11605 3282 11657
rect 2737 9041 2790 11605
rect 3217 11604 3282 11605
rect 9189 11521 9263 11525
rect 8786 11500 8860 11504
rect 8786 11444 8795 11500
rect 8851 11444 8860 11500
rect 9189 11465 9198 11521
rect 9254 11465 9263 11521
rect 9189 11461 9263 11465
rect 8786 11440 8860 11444
rect 3043 10575 3117 10579
rect 3043 10519 3052 10575
rect 3108 10519 3117 10575
rect 3043 10515 3117 10519
rect 3578 10578 3910 10582
rect 3578 10522 3594 10578
rect 3650 10522 3674 10578
rect 3730 10522 3754 10578
rect 3810 10522 3834 10578
rect 3890 10522 3910 10578
rect 3578 10514 3910 10522
rect 4310 10578 4642 10582
rect 4310 10522 4326 10578
rect 4382 10522 4406 10578
rect 4462 10522 4486 10578
rect 4542 10522 4566 10578
rect 4622 10522 4642 10578
rect 4310 10514 4642 10522
rect 4912 10578 5244 10582
rect 4912 10522 4932 10578
rect 4988 10522 5012 10578
rect 5068 10522 5092 10578
rect 5148 10522 5172 10578
rect 5228 10522 5244 10578
rect 4912 10514 5244 10522
rect 5522 10578 5854 10582
rect 5522 10522 5538 10578
rect 5594 10522 5618 10578
rect 5674 10522 5698 10578
rect 5754 10522 5778 10578
rect 5834 10522 5854 10578
rect 5522 10514 5854 10522
rect 6124 10578 6456 10582
rect 6124 10522 6144 10578
rect 6200 10522 6224 10578
rect 6280 10522 6304 10578
rect 6360 10522 6384 10578
rect 6440 10522 6456 10578
rect 6124 10514 6456 10522
rect 6860 10578 7192 10582
rect 6860 10522 6876 10578
rect 6932 10522 6956 10578
rect 7012 10522 7036 10578
rect 7092 10522 7116 10578
rect 7172 10522 7192 10578
rect 6860 10514 7192 10522
rect 7462 10578 7794 10582
rect 7462 10522 7482 10578
rect 7538 10522 7562 10578
rect 7618 10522 7642 10578
rect 7698 10522 7722 10578
rect 7778 10522 7794 10578
rect 7462 10514 7794 10522
rect 8196 10578 8528 10582
rect 8196 10522 8216 10578
rect 8272 10522 8296 10578
rect 8352 10522 8376 10578
rect 8432 10522 8456 10578
rect 8512 10522 8528 10578
rect 8196 10514 8528 10522
rect 3043 10127 3117 10131
rect 3043 10071 3052 10127
rect 3108 10071 3117 10127
rect 3043 10067 3117 10071
rect 3578 10124 3910 10132
rect 3578 10068 3594 10124
rect 3650 10068 3674 10124
rect 3730 10068 3754 10124
rect 3810 10068 3834 10124
rect 3890 10068 3910 10124
rect 3578 10064 3910 10068
rect 4310 10124 4642 10132
rect 4310 10068 4326 10124
rect 4382 10068 4406 10124
rect 4462 10068 4486 10124
rect 4542 10068 4566 10124
rect 4622 10068 4642 10124
rect 4310 10064 4642 10068
rect 4912 10124 5244 10132
rect 4912 10068 4932 10124
rect 4988 10068 5012 10124
rect 5068 10068 5092 10124
rect 5148 10068 5172 10124
rect 5228 10068 5244 10124
rect 4912 10064 5244 10068
rect 5522 10124 5854 10132
rect 5522 10068 5538 10124
rect 5594 10068 5618 10124
rect 5674 10068 5698 10124
rect 5754 10068 5778 10124
rect 5834 10068 5854 10124
rect 5522 10064 5854 10068
rect 6124 10124 6456 10132
rect 6124 10068 6144 10124
rect 6200 10068 6224 10124
rect 6280 10068 6304 10124
rect 6360 10068 6384 10124
rect 6440 10068 6456 10124
rect 6124 10064 6456 10068
rect 6860 10124 7192 10132
rect 6860 10068 6876 10124
rect 6932 10068 6956 10124
rect 7012 10068 7036 10124
rect 7092 10068 7116 10124
rect 7172 10068 7192 10124
rect 6860 10064 7192 10068
rect 7462 10124 7794 10132
rect 7462 10068 7482 10124
rect 7538 10068 7562 10124
rect 7618 10068 7642 10124
rect 7698 10068 7722 10124
rect 7778 10068 7794 10124
rect 7462 10064 7794 10068
rect 8196 10124 8528 10132
rect 8196 10068 8216 10124
rect 8272 10068 8296 10124
rect 8352 10068 8376 10124
rect 8432 10068 8456 10124
rect 8512 10068 8528 10124
rect 8196 10064 8528 10068
rect 8786 9202 8860 9206
rect 8786 9146 8795 9202
rect 8851 9146 8860 9202
rect 8786 9142 8860 9146
rect 9214 9161 9288 9165
rect 9214 9105 9223 9161
rect 9279 9105 9288 9161
rect 9214 9101 9288 9105
rect 9691 9161 9765 9165
rect 9691 9105 9700 9161
rect 9756 9105 9765 9161
rect 9691 9101 9765 9105
rect 10111 9150 10185 9154
rect 10111 9094 10120 9150
rect 10176 9094 10185 9150
rect 10111 9090 10185 9094
rect 3217 9041 3282 9042
rect 2730 8989 2736 9041
rect 2788 9038 2795 9041
rect 3217 9038 3224 9041
rect 2788 8992 3224 9038
rect 2788 8989 2795 8992
rect 2730 8988 2795 8989
rect 2467 8700 2523 8709
rect 2467 8635 2523 8644
rect 2587 8700 2643 8709
rect 2587 8635 2643 8644
rect 2730 8700 2786 8709
rect 2730 8635 2786 8644
rect 2927 8586 2973 8992
rect 3217 8989 3224 8992
rect 3276 8989 3282 9041
rect 3895 8945 3977 8946
rect 3895 8881 3904 8945
rect 3968 8881 3977 8945
rect 4627 8945 4709 8946
rect 4627 8881 4636 8945
rect 4700 8881 4709 8945
rect 4845 8945 4927 8946
rect 4845 8881 4854 8945
rect 4918 8881 4927 8945
rect 5839 8945 5921 8946
rect 5839 8881 5848 8945
rect 5912 8881 5921 8945
rect 6057 8945 6139 8946
rect 6057 8881 6066 8945
rect 6130 8881 6139 8945
rect 7177 8945 7259 8946
rect 7177 8881 7186 8945
rect 7250 8881 7259 8945
rect 7395 8945 7477 8946
rect 7395 8881 7404 8945
rect 7468 8881 7477 8945
rect 8129 8945 8211 8946
rect 8129 8881 8138 8945
rect 8202 8881 8211 8945
rect 8877 8940 8951 8944
rect 8877 8884 8886 8940
rect 8942 8884 8951 8940
rect 10314 8923 10342 11808
rect 11646 11672 11674 12259
rect 12753 12186 12759 12239
rect 12811 12186 12817 12239
rect 12753 12185 12817 12186
rect 11775 11878 11850 11882
rect 11775 11822 11785 11878
rect 11841 11822 11850 11878
rect 11976 11879 12051 11883
rect 11976 11823 11986 11879
rect 12042 11823 12051 11879
rect 11976 11822 12051 11823
rect 12162 11877 12237 11881
rect 11775 11821 11850 11822
rect 12162 11821 12172 11877
rect 12228 11821 12237 11877
rect 12353 11880 12428 11884
rect 12353 11824 12363 11880
rect 12419 11824 12428 11880
rect 12353 11823 12428 11824
rect 12566 11879 12641 11883
rect 12566 11823 12576 11879
rect 12632 11823 12641 11879
rect 12566 11822 12641 11823
rect 12162 11820 12237 11821
rect 12774 11745 12802 12185
rect 13618 12132 13683 12133
rect 13618 12080 13624 12132
rect 13676 12129 13683 12132
rect 13815 12129 13861 12535
rect 20064 12477 20120 12486
rect 15161 12442 15240 12443
rect 15388 12442 15467 12443
rect 16373 12442 16452 12443
rect 16600 12442 16679 12443
rect 17585 12442 17664 12443
rect 17812 12442 17891 12443
rect 18797 12442 18876 12443
rect 19024 12442 19103 12443
rect 14429 12439 14508 12440
rect 14426 12375 14436 12439
rect 14500 12375 14509 12439
rect 15158 12378 15168 12442
rect 15232 12378 15241 12442
rect 15387 12378 15396 12442
rect 15460 12378 15470 12442
rect 16370 12378 16380 12442
rect 16444 12378 16453 12442
rect 16599 12378 16608 12442
rect 16672 12378 16682 12442
rect 17582 12378 17592 12442
rect 17656 12378 17665 12442
rect 17811 12378 17820 12442
rect 17884 12378 17894 12442
rect 18794 12378 18804 12442
rect 18868 12378 18877 12442
rect 19023 12378 19032 12442
rect 19096 12378 19106 12442
rect 19765 12440 19839 12444
rect 19765 12384 19774 12440
rect 19830 12384 19839 12440
rect 20064 12412 20120 12421
rect 20184 12477 20240 12486
rect 20184 12412 20240 12421
rect 20327 12477 20383 12486
rect 20327 12412 20383 12421
rect 19765 12380 19839 12384
rect 14783 12176 14792 12240
rect 14856 12176 14865 12240
rect 14783 12175 14865 12176
rect 15515 12176 15524 12240
rect 15588 12176 15597 12240
rect 15515 12175 15597 12176
rect 15733 12176 15742 12240
rect 15806 12176 15815 12240
rect 15733 12175 15815 12176
rect 16727 12176 16736 12240
rect 16800 12176 16809 12240
rect 16727 12175 16809 12176
rect 16945 12176 16954 12240
rect 17018 12176 17027 12240
rect 16945 12175 17027 12176
rect 18065 12176 18074 12240
rect 18138 12176 18147 12240
rect 18065 12175 18147 12176
rect 18283 12176 18292 12240
rect 18356 12176 18365 12240
rect 18283 12175 18365 12176
rect 19017 12176 19026 12240
rect 19090 12176 19099 12240
rect 19765 12237 19839 12241
rect 19765 12181 19774 12237
rect 19830 12181 19839 12237
rect 19765 12177 19839 12181
rect 19017 12175 19099 12176
rect 20327 12132 20392 12133
rect 14105 12129 14112 12132
rect 13676 12083 14112 12129
rect 13676 12080 13683 12083
rect 14105 12080 14112 12083
rect 14164 12080 14170 12132
rect 20327 12080 20333 12132
rect 20385 12129 20392 12132
rect 20524 12129 20570 12535
rect 21870 12442 21949 12443
rect 22097 12442 22176 12443
rect 23082 12442 23161 12443
rect 23309 12442 23388 12443
rect 24294 12442 24373 12443
rect 24521 12442 24600 12443
rect 25506 12442 25585 12443
rect 25733 12442 25812 12443
rect 21138 12439 21217 12440
rect 21135 12375 21145 12439
rect 21209 12375 21218 12439
rect 21867 12378 21877 12442
rect 21941 12378 21950 12442
rect 22096 12378 22105 12442
rect 22169 12378 22179 12442
rect 23079 12378 23089 12442
rect 23153 12378 23162 12442
rect 23308 12378 23317 12442
rect 23381 12378 23391 12442
rect 24291 12378 24301 12442
rect 24365 12378 24374 12442
rect 24520 12378 24529 12442
rect 24593 12378 24603 12442
rect 25503 12378 25513 12442
rect 25577 12378 25586 12442
rect 25732 12378 25741 12442
rect 25805 12378 25815 12442
rect 26474 12440 26548 12444
rect 26474 12384 26483 12440
rect 26539 12384 26548 12440
rect 26474 12380 26548 12384
rect 21492 12176 21501 12240
rect 21565 12176 21574 12240
rect 21492 12175 21574 12176
rect 22224 12176 22233 12240
rect 22297 12176 22306 12240
rect 22224 12175 22306 12176
rect 22442 12176 22451 12240
rect 22515 12176 22524 12240
rect 22442 12175 22524 12176
rect 23436 12176 23445 12240
rect 23509 12176 23518 12240
rect 23436 12175 23518 12176
rect 23654 12176 23663 12240
rect 23727 12176 23736 12240
rect 23654 12175 23736 12176
rect 24774 12176 24783 12240
rect 24847 12176 24856 12240
rect 24774 12175 24856 12176
rect 24992 12176 25001 12240
rect 25065 12176 25074 12240
rect 24992 12175 25074 12176
rect 25726 12176 25735 12240
rect 25799 12176 25808 12240
rect 26474 12237 26548 12241
rect 26474 12181 26483 12237
rect 26539 12181 26548 12237
rect 26474 12177 26548 12181
rect 25726 12175 25808 12176
rect 20814 12129 20821 12132
rect 20385 12083 20821 12129
rect 20385 12080 20392 12083
rect 20814 12080 20821 12083
rect 20873 12080 20879 12132
rect 14105 12079 14170 12080
rect 20814 12079 20879 12080
rect 13199 12002 13205 12054
rect 13257 12002 13263 12054
rect 12755 11693 12761 11745
rect 12813 11693 12819 11745
rect 11628 11620 11634 11672
rect 11686 11620 11692 11672
rect 10924 11259 10998 11263
rect 10924 11203 10933 11259
rect 10989 11203 10998 11259
rect 10924 11199 10998 11203
rect 11112 11256 11186 11260
rect 11112 11200 11121 11256
rect 11177 11200 11186 11256
rect 11112 11196 11186 11200
rect 11309 11254 11383 11258
rect 11309 11198 11318 11254
rect 11374 11198 11383 11254
rect 11309 11194 11383 11198
rect 13209 10030 13253 12002
rect 13284 11595 13411 11610
rect 13284 11537 13314 11595
rect 13381 11537 13411 11595
rect 13284 11519 13411 11537
rect 13931 11050 14005 11054
rect 13931 10994 13940 11050
rect 13996 10994 14005 11050
rect 13931 10990 14005 10994
rect 14112 10581 14164 12079
rect 19674 11975 19748 11979
rect 19674 11919 19683 11975
rect 19739 11919 19748 11975
rect 19674 11915 19748 11919
rect 14466 11053 14798 11057
rect 14466 10997 14482 11053
rect 14538 10997 14562 11053
rect 14618 10997 14642 11053
rect 14698 10997 14722 11053
rect 14778 10997 14798 11053
rect 14466 10989 14798 10997
rect 15198 11053 15530 11057
rect 15198 10997 15214 11053
rect 15270 10997 15294 11053
rect 15350 10997 15374 11053
rect 15430 10997 15454 11053
rect 15510 10997 15530 11053
rect 15198 10989 15530 10997
rect 15800 11053 16132 11057
rect 15800 10997 15820 11053
rect 15876 10997 15900 11053
rect 15956 10997 15980 11053
rect 16036 10997 16060 11053
rect 16116 10997 16132 11053
rect 15800 10989 16132 10997
rect 16410 11053 16742 11057
rect 16410 10997 16426 11053
rect 16482 10997 16506 11053
rect 16562 10997 16586 11053
rect 16642 10997 16666 11053
rect 16722 10997 16742 11053
rect 16410 10989 16742 10997
rect 17012 11053 17344 11057
rect 17012 10997 17032 11053
rect 17088 10997 17112 11053
rect 17168 10997 17192 11053
rect 17248 10997 17272 11053
rect 17328 10997 17344 11053
rect 17012 10989 17344 10997
rect 17748 11053 18080 11057
rect 17748 10997 17764 11053
rect 17820 10997 17844 11053
rect 17900 10997 17924 11053
rect 17980 10997 18004 11053
rect 18060 10997 18080 11053
rect 17748 10989 18080 10997
rect 18350 11053 18682 11057
rect 18350 10997 18370 11053
rect 18426 10997 18450 11053
rect 18506 10997 18530 11053
rect 18586 10997 18610 11053
rect 18666 10997 18682 11053
rect 18350 10989 18682 10997
rect 19084 11053 19416 11057
rect 19084 10997 19104 11053
rect 19160 10997 19184 11053
rect 19240 10997 19264 11053
rect 19320 10997 19344 11053
rect 19400 10997 19416 11053
rect 19084 10989 19416 10997
rect 20640 11050 20714 11054
rect 20640 10994 20649 11050
rect 20705 10994 20714 11050
rect 20640 10990 20714 10994
rect 14103 10578 14173 10581
rect 14103 10526 14112 10578
rect 14164 10526 14173 10578
rect 20821 10575 20873 12079
rect 26383 11975 26457 11979
rect 26383 11919 26392 11975
rect 26448 11919 26457 11975
rect 26383 11915 26457 11919
rect 21175 11053 21507 11057
rect 21175 10997 21191 11053
rect 21247 10997 21271 11053
rect 21327 10997 21351 11053
rect 21407 10997 21431 11053
rect 21487 10997 21507 11053
rect 21175 10989 21507 10997
rect 21907 11053 22239 11057
rect 21907 10997 21923 11053
rect 21979 10997 22003 11053
rect 22059 10997 22083 11053
rect 22139 10997 22163 11053
rect 22219 10997 22239 11053
rect 21907 10989 22239 10997
rect 22509 11053 22841 11057
rect 22509 10997 22529 11053
rect 22585 10997 22609 11053
rect 22665 10997 22689 11053
rect 22745 10997 22769 11053
rect 22825 10997 22841 11053
rect 22509 10989 22841 10997
rect 23119 11053 23451 11057
rect 23119 10997 23135 11053
rect 23191 10997 23215 11053
rect 23271 10997 23295 11053
rect 23351 10997 23375 11053
rect 23431 10997 23451 11053
rect 23119 10989 23451 10997
rect 23721 11053 24053 11057
rect 23721 10997 23741 11053
rect 23797 10997 23821 11053
rect 23877 10997 23901 11053
rect 23957 10997 23981 11053
rect 24037 10997 24053 11053
rect 23721 10989 24053 10997
rect 24457 11053 24789 11057
rect 24457 10997 24473 11053
rect 24529 10997 24553 11053
rect 24609 10997 24633 11053
rect 24689 10997 24713 11053
rect 24769 10997 24789 11053
rect 24457 10989 24789 10997
rect 25059 11053 25391 11057
rect 25059 10997 25079 11053
rect 25135 10997 25159 11053
rect 25215 10997 25239 11053
rect 25295 10997 25319 11053
rect 25375 10997 25391 11053
rect 25059 10989 25391 10997
rect 25793 11053 26125 11057
rect 25793 10997 25813 11053
rect 25869 10997 25893 11053
rect 25949 10997 25973 11053
rect 26029 10997 26053 11053
rect 26109 10997 26125 11053
rect 25793 10989 26125 10997
rect 25710 10579 25786 10580
rect 14103 10518 14173 10526
rect 19003 10568 19073 10575
rect 19003 10516 19012 10568
rect 19065 10516 19073 10568
rect 20814 10571 20882 10575
rect 20814 10518 20821 10571
rect 20873 10518 20882 10571
rect 19003 10508 19073 10516
rect 25710 10515 25716 10579
rect 25780 10515 25786 10579
rect 13763 10112 14095 10120
rect 13763 10056 13779 10112
rect 13835 10056 13859 10112
rect 13915 10056 13939 10112
rect 13995 10056 14019 10112
rect 14075 10056 14095 10112
rect 13763 10052 14095 10056
rect 14497 10112 14829 10120
rect 14497 10056 14513 10112
rect 14569 10056 14593 10112
rect 14649 10056 14673 10112
rect 14729 10056 14753 10112
rect 14809 10056 14829 10112
rect 14497 10052 14829 10056
rect 15099 10112 15431 10120
rect 15099 10056 15119 10112
rect 15175 10056 15199 10112
rect 15255 10056 15279 10112
rect 15335 10056 15359 10112
rect 15415 10056 15431 10112
rect 15099 10052 15431 10056
rect 15835 10112 16167 10120
rect 15835 10056 15851 10112
rect 15907 10056 15931 10112
rect 15987 10056 16011 10112
rect 16067 10056 16091 10112
rect 16147 10056 16167 10112
rect 15835 10052 16167 10056
rect 16437 10112 16769 10120
rect 16437 10056 16457 10112
rect 16513 10056 16537 10112
rect 16593 10056 16617 10112
rect 16673 10056 16697 10112
rect 16753 10056 16769 10112
rect 16437 10052 16769 10056
rect 17047 10112 17379 10120
rect 17047 10056 17063 10112
rect 17119 10056 17143 10112
rect 17199 10056 17223 10112
rect 17279 10056 17303 10112
rect 17359 10056 17379 10112
rect 17047 10052 17379 10056
rect 17649 10112 17981 10120
rect 17649 10056 17669 10112
rect 17725 10056 17749 10112
rect 17805 10056 17829 10112
rect 17885 10056 17909 10112
rect 17965 10056 17981 10112
rect 17649 10052 17981 10056
rect 18381 10112 18713 10120
rect 18381 10056 18401 10112
rect 18457 10056 18481 10112
rect 18537 10056 18561 10112
rect 18617 10056 18641 10112
rect 18697 10056 18713 10112
rect 18381 10052 18713 10056
rect 12671 9976 12677 10028
rect 12729 9976 12735 10028
rect 13199 9978 13205 10030
rect 13257 9978 13263 10030
rect 10487 9158 10561 9162
rect 10487 9102 10496 9158
rect 10552 9102 10561 9158
rect 10487 9098 10561 9102
rect 8877 8880 8951 8884
rect 10302 8913 10357 8923
rect 10302 8859 10303 8913
rect 10302 8852 10357 8859
rect 3538 8682 3548 8746
rect 3612 8682 3621 8746
rect 3541 8681 3620 8682
rect 4270 8679 4280 8743
rect 4344 8679 4353 8743
rect 4499 8679 4508 8743
rect 4572 8679 4582 8743
rect 5482 8679 5492 8743
rect 5556 8679 5565 8743
rect 5711 8679 5720 8743
rect 5784 8679 5794 8743
rect 6694 8679 6704 8743
rect 6768 8679 6777 8743
rect 6923 8679 6932 8743
rect 6996 8679 7006 8743
rect 7906 8679 7916 8743
rect 7980 8679 7989 8743
rect 8135 8679 8144 8743
rect 8208 8679 8218 8743
rect 8877 8737 8951 8741
rect 8877 8681 8886 8737
rect 8942 8681 8951 8737
rect 4273 8678 4352 8679
rect 4500 8678 4579 8679
rect 5485 8678 5564 8679
rect 5712 8678 5791 8679
rect 6697 8678 6776 8679
rect 6924 8678 7003 8679
rect 7909 8678 7988 8679
rect 8136 8678 8215 8679
rect 8877 8677 8951 8681
rect 9333 8654 9386 8666
rect 9385 8601 9386 8654
rect 9333 8589 9386 8601
rect 2734 8540 2973 8586
rect 2734 8464 2780 8540
rect 8789 8476 8863 8480
rect 2716 8463 2782 8464
rect 2716 8411 2724 8463
rect 2776 8411 2782 8463
rect 8789 8420 8798 8476
rect 8854 8420 8863 8476
rect 8789 8416 8863 8420
rect 9199 8450 9273 8454
rect 2984 8392 3036 8399
rect 9199 8394 9208 8450
rect 9264 8394 9273 8450
rect 9199 8390 9273 8394
rect 2984 8334 3036 8340
rect 2449 8154 2505 8163
rect 2449 8089 2505 8098
rect 2580 8155 2636 8164
rect 2580 8090 2636 8099
rect 2724 8154 2780 8163
rect 2724 8089 2780 8098
rect 2993 7410 3027 8334
rect 8871 8234 8945 8238
rect 8871 8178 8880 8234
rect 8936 8178 8945 8234
rect 8871 8174 8945 8178
rect 8872 8077 8946 8081
rect 8872 8021 8881 8077
rect 8937 8021 8946 8077
rect 9351 8050 9379 8589
rect 9461 8451 9535 8455
rect 9461 8395 9470 8451
rect 9526 8395 9535 8451
rect 9461 8391 9535 8395
rect 9733 8451 9807 8455
rect 9733 8395 9742 8451
rect 9798 8395 9807 8451
rect 9733 8391 9807 8395
rect 10060 8451 10134 8455
rect 10060 8395 10069 8451
rect 10125 8395 10134 8451
rect 10060 8391 10134 8395
rect 10441 8451 10515 8455
rect 10441 8395 10450 8451
rect 10506 8395 10515 8451
rect 10441 8391 10515 8395
rect 10746 8124 10780 9459
rect 11093 9164 11167 9168
rect 10835 9158 10909 9162
rect 10835 9102 10844 9158
rect 10900 9102 10909 9158
rect 11093 9108 11102 9164
rect 11158 9108 11167 9164
rect 11093 9104 11167 9108
rect 11319 9164 11393 9168
rect 11319 9108 11328 9164
rect 11384 9108 11393 9164
rect 11319 9104 11393 9108
rect 11578 9167 11652 9171
rect 11578 9111 11587 9167
rect 11643 9111 11652 9167
rect 11578 9107 11652 9111
rect 12185 9129 12259 9133
rect 10835 9098 10909 9102
rect 12185 9073 12194 9129
rect 12250 9073 12259 9129
rect 12185 9069 12259 9073
rect 12417 9130 12491 9134
rect 12417 9074 12426 9130
rect 12482 9074 12491 9130
rect 12417 9070 12491 9074
rect 12579 8834 12643 8835
rect 12579 8781 12585 8834
rect 12637 8781 12643 8834
rect 12681 8824 12725 9976
rect 13431 9190 13505 9194
rect 12853 9136 12927 9140
rect 12853 9080 12862 9136
rect 12918 9080 12927 9136
rect 12853 9076 12927 9080
rect 13088 9138 13162 9142
rect 13088 9082 13097 9138
rect 13153 9082 13162 9138
rect 13431 9134 13440 9190
rect 13496 9134 13505 9190
rect 13431 9130 13505 9134
rect 13088 9078 13162 9082
rect 19011 9030 19063 10508
rect 19174 10115 19248 10119
rect 19174 10059 19183 10115
rect 19239 10059 19248 10115
rect 19174 10055 19248 10059
rect 20472 10112 20804 10120
rect 20472 10056 20488 10112
rect 20544 10056 20568 10112
rect 20624 10056 20648 10112
rect 20704 10056 20728 10112
rect 20784 10056 20804 10112
rect 20472 10052 20804 10056
rect 21206 10112 21538 10120
rect 21206 10056 21222 10112
rect 21278 10056 21302 10112
rect 21358 10056 21382 10112
rect 21438 10056 21462 10112
rect 21518 10056 21538 10112
rect 21206 10052 21538 10056
rect 21808 10112 22140 10120
rect 21808 10056 21828 10112
rect 21884 10056 21908 10112
rect 21964 10056 21988 10112
rect 22044 10056 22068 10112
rect 22124 10056 22140 10112
rect 21808 10052 22140 10056
rect 22544 10112 22876 10120
rect 22544 10056 22560 10112
rect 22616 10056 22640 10112
rect 22696 10056 22720 10112
rect 22776 10056 22800 10112
rect 22856 10056 22876 10112
rect 22544 10052 22876 10056
rect 23146 10112 23478 10120
rect 23146 10056 23166 10112
rect 23222 10056 23246 10112
rect 23302 10056 23326 10112
rect 23382 10056 23406 10112
rect 23462 10056 23478 10112
rect 23146 10052 23478 10056
rect 23756 10112 24088 10120
rect 23756 10056 23772 10112
rect 23828 10056 23852 10112
rect 23908 10056 23932 10112
rect 23988 10056 24012 10112
rect 24068 10056 24088 10112
rect 23756 10052 24088 10056
rect 24358 10112 24690 10120
rect 24358 10056 24378 10112
rect 24434 10056 24458 10112
rect 24514 10056 24538 10112
rect 24594 10056 24618 10112
rect 24674 10056 24690 10112
rect 24358 10052 24690 10056
rect 25090 10112 25422 10120
rect 25090 10056 25110 10112
rect 25166 10056 25190 10112
rect 25246 10056 25270 10112
rect 25326 10056 25350 10112
rect 25406 10056 25422 10112
rect 25090 10052 25422 10056
rect 20140 9190 20214 9194
rect 20140 9134 20149 9190
rect 20205 9134 20214 9190
rect 20140 9130 20214 9134
rect 25723 9030 25775 10515
rect 25883 10115 25957 10119
rect 25883 10059 25892 10115
rect 25948 10059 25957 10115
rect 25883 10055 25957 10059
rect 19009 9029 19074 9030
rect 25718 9029 25783 9030
rect 19009 8977 19015 9029
rect 19067 9026 19074 9029
rect 19496 9026 19503 9029
rect 19067 8980 19503 9026
rect 19067 8977 19074 8980
rect 14080 8933 14162 8934
rect 13340 8928 13414 8932
rect 13340 8872 13349 8928
rect 13405 8872 13414 8928
rect 13340 8868 13414 8872
rect 14080 8869 14089 8933
rect 14153 8869 14162 8933
rect 14814 8933 14896 8934
rect 14814 8869 14823 8933
rect 14887 8869 14896 8933
rect 15032 8933 15114 8934
rect 15032 8869 15041 8933
rect 15105 8869 15114 8933
rect 16152 8933 16234 8934
rect 16152 8869 16161 8933
rect 16225 8869 16234 8933
rect 16370 8933 16452 8934
rect 16370 8869 16379 8933
rect 16443 8869 16452 8933
rect 17364 8933 17446 8934
rect 17364 8869 17373 8933
rect 17437 8869 17446 8933
rect 17582 8933 17664 8934
rect 17582 8869 17591 8933
rect 17655 8869 17664 8933
rect 18314 8933 18396 8934
rect 18314 8869 18323 8933
rect 18387 8869 18396 8933
rect 11538 8728 11544 8780
rect 11596 8728 11602 8780
rect 10817 8451 10892 8455
rect 10817 8395 10827 8451
rect 10883 8395 10892 8451
rect 10817 8391 10892 8395
rect 11556 8130 11590 8728
rect 12590 8648 12633 8781
rect 12671 8772 12677 8824
rect 12729 8772 12735 8824
rect 13340 8725 13414 8729
rect 13340 8669 13349 8725
rect 13405 8669 13414 8725
rect 13340 8665 13414 8669
rect 14073 8667 14083 8731
rect 14147 8667 14156 8731
rect 14302 8667 14311 8731
rect 14375 8667 14385 8731
rect 15285 8667 15295 8731
rect 15359 8667 15368 8731
rect 15514 8667 15523 8731
rect 15587 8667 15597 8731
rect 16497 8667 16507 8731
rect 16571 8667 16580 8731
rect 16726 8667 16735 8731
rect 16799 8667 16809 8731
rect 17709 8667 17719 8731
rect 17783 8667 17792 8731
rect 17938 8667 17947 8731
rect 18011 8667 18021 8731
rect 18670 8670 18679 8734
rect 18743 8670 18753 8734
rect 18671 8669 18750 8670
rect 14076 8666 14155 8667
rect 14303 8666 14382 8667
rect 15288 8666 15367 8667
rect 15515 8666 15594 8667
rect 16500 8666 16579 8667
rect 16727 8666 16806 8667
rect 17712 8666 17791 8667
rect 17939 8666 18018 8667
rect 12590 8642 12646 8648
rect 12926 8645 12967 8646
rect 12590 8590 12594 8642
rect 12590 8587 12646 8590
rect 12594 8584 12646 8587
rect 12922 8639 12975 8645
rect 12922 8587 12923 8639
rect 12922 8584 12975 8587
rect 12923 8581 12975 8584
rect 12712 8510 12787 8514
rect 12712 8454 12722 8510
rect 12778 8454 12787 8510
rect 12712 8453 12787 8454
rect 12217 8440 12292 8444
rect 12217 8384 12227 8440
rect 12283 8384 12292 8440
rect 12217 8383 12292 8384
rect 12574 8367 12649 8371
rect 12574 8311 12584 8367
rect 12640 8311 12649 8367
rect 12574 8310 12649 8311
rect 12758 8364 12833 8368
rect 12758 8308 12768 8364
rect 12824 8308 12833 8364
rect 12758 8307 12833 8308
rect 10624 8121 10780 8124
rect 10624 8069 10706 8121
rect 10758 8069 10780 8121
rect 10624 8067 10780 8069
rect 8872 8017 8946 8021
rect 9333 8049 9398 8050
rect 9333 7996 9340 8049
rect 9392 7996 9398 8049
rect 8872 7907 8946 7911
rect 8872 7851 8881 7907
rect 8937 7851 8946 7907
rect 8872 7847 8946 7851
rect 8871 7755 8945 7759
rect 8871 7699 8880 7755
rect 8936 7699 8945 7755
rect 8871 7695 8945 7699
rect 10135 7725 10209 7729
rect 10135 7669 10144 7725
rect 10200 7669 10209 7725
rect 10135 7665 10209 7669
rect 10383 7725 10457 7729
rect 10383 7669 10392 7725
rect 10448 7669 10457 7725
rect 10383 7665 10457 7669
rect 8866 7611 8940 7615
rect 3058 7558 3728 7564
rect 3058 7553 3162 7558
rect 3057 7549 3162 7553
rect 3057 7493 3066 7549
rect 3122 7502 3162 7549
rect 3218 7502 3242 7558
rect 3298 7502 3322 7558
rect 3378 7502 3402 7558
rect 3458 7502 3482 7558
rect 3538 7502 3562 7558
rect 3618 7502 3728 7558
rect 3122 7498 3728 7502
rect 3790 7555 8698 7561
rect 3790 7499 3894 7555
rect 3950 7499 3974 7555
rect 4030 7499 4054 7555
rect 4110 7499 4134 7555
rect 4190 7499 4214 7555
rect 4270 7499 4294 7555
rect 4350 7499 4502 7555
rect 4558 7499 4582 7555
rect 4638 7499 4662 7555
rect 4718 7499 4742 7555
rect 4798 7499 4822 7555
rect 4878 7499 4902 7555
rect 4958 7499 5106 7555
rect 5162 7499 5186 7555
rect 5242 7499 5266 7555
rect 5322 7499 5346 7555
rect 5402 7499 5426 7555
rect 5482 7499 5506 7555
rect 5562 7499 5714 7555
rect 5770 7499 5794 7555
rect 5850 7499 5874 7555
rect 5930 7499 5954 7555
rect 6010 7499 6034 7555
rect 6090 7499 6114 7555
rect 6170 7499 6318 7555
rect 6374 7499 6398 7555
rect 6454 7499 6478 7555
rect 6534 7499 6558 7555
rect 6614 7499 6638 7555
rect 6694 7499 6718 7555
rect 6774 7499 6926 7555
rect 6982 7499 7006 7555
rect 7062 7499 7086 7555
rect 7142 7499 7166 7555
rect 7222 7499 7246 7555
rect 7302 7499 7326 7555
rect 7382 7499 7530 7555
rect 7586 7499 7610 7555
rect 7666 7499 7690 7555
rect 7746 7499 7770 7555
rect 7826 7499 7850 7555
rect 7906 7499 7930 7555
rect 7986 7499 8138 7555
rect 8194 7499 8218 7555
rect 8274 7499 8298 7555
rect 8354 7499 8378 7555
rect 8434 7499 8458 7555
rect 8514 7499 8538 7555
rect 8594 7499 8698 7555
rect 8866 7555 8875 7611
rect 8931 7555 8940 7611
rect 8866 7551 8940 7555
rect 3122 7493 3131 7498
rect 3790 7495 8698 7499
rect 3057 7489 3131 7493
rect 10305 7481 10311 7533
rect 10363 7481 10369 7533
rect 2978 7358 2985 7410
rect 3038 7358 3044 7410
rect 9945 7358 9951 7410
rect 10003 7358 10029 7410
rect 10001 6796 10029 7358
rect 9982 6744 9988 6796
rect 10040 6744 10046 6796
rect 10001 2976 10029 6744
rect 10323 5246 10351 7481
rect 10624 7334 10652 8067
rect 10746 8063 10780 8067
rect 11518 8122 11590 8130
rect 11518 8070 11524 8122
rect 11576 8070 11590 8122
rect 11518 8064 11590 8070
rect 10680 7725 10754 7729
rect 10680 7669 10689 7725
rect 10745 7669 10754 7725
rect 10680 7665 10754 7669
rect 11024 7727 11098 7731
rect 11024 7671 11033 7727
rect 11089 7671 11098 7727
rect 11024 7667 11098 7671
rect 11343 7727 11417 7731
rect 11343 7671 11352 7727
rect 11408 7671 11417 7727
rect 11343 7667 11417 7671
rect 11556 7587 11590 8064
rect 12926 8040 12967 8581
rect 19318 8574 19364 8980
rect 19496 8977 19503 8980
rect 19555 8977 19561 9029
rect 25718 8977 25724 9029
rect 25776 9026 25783 9029
rect 26205 9026 26212 9029
rect 25776 8980 26212 9026
rect 25776 8977 25783 8980
rect 19496 8976 19561 8977
rect 20789 8933 20871 8934
rect 20049 8928 20123 8932
rect 20049 8872 20058 8928
rect 20114 8872 20123 8928
rect 20049 8868 20123 8872
rect 20789 8869 20798 8933
rect 20862 8869 20871 8933
rect 21523 8933 21605 8934
rect 21523 8869 21532 8933
rect 21596 8869 21605 8933
rect 21741 8933 21823 8934
rect 21741 8869 21750 8933
rect 21814 8869 21823 8933
rect 22861 8933 22943 8934
rect 22861 8869 22870 8933
rect 22934 8869 22943 8933
rect 23079 8933 23161 8934
rect 23079 8869 23088 8933
rect 23152 8869 23161 8933
rect 24073 8933 24155 8934
rect 24073 8869 24082 8933
rect 24146 8869 24155 8933
rect 24291 8933 24373 8934
rect 24291 8869 24300 8933
rect 24364 8869 24373 8933
rect 25023 8933 25105 8934
rect 25023 8869 25032 8933
rect 25096 8869 25105 8933
rect 20049 8725 20123 8729
rect 19505 8688 19561 8697
rect 19505 8623 19561 8632
rect 19648 8688 19704 8697
rect 19648 8623 19704 8632
rect 19768 8688 19824 8697
rect 20049 8669 20058 8725
rect 20114 8669 20123 8725
rect 20049 8665 20123 8669
rect 20782 8667 20792 8731
rect 20856 8667 20865 8731
rect 21011 8667 21020 8731
rect 21084 8667 21094 8731
rect 21994 8667 22004 8731
rect 22068 8667 22077 8731
rect 22223 8667 22232 8731
rect 22296 8667 22306 8731
rect 23206 8667 23216 8731
rect 23280 8667 23289 8731
rect 23435 8667 23444 8731
rect 23508 8667 23518 8731
rect 24418 8667 24428 8731
rect 24492 8667 24501 8731
rect 24647 8667 24656 8731
rect 24720 8667 24730 8731
rect 25379 8670 25388 8734
rect 25452 8670 25462 8734
rect 25380 8669 25459 8670
rect 20785 8666 20864 8667
rect 21012 8666 21091 8667
rect 21997 8666 22076 8667
rect 22224 8666 22303 8667
rect 23209 8666 23288 8667
rect 23436 8666 23515 8667
rect 24421 8666 24500 8667
rect 24648 8666 24727 8667
rect 19768 8623 19824 8632
rect 26027 8574 26073 8980
rect 26205 8977 26212 8980
rect 26264 8977 26270 9029
rect 26205 8976 26270 8977
rect 26214 8688 26270 8697
rect 26214 8623 26270 8632
rect 26357 8688 26413 8697
rect 26357 8623 26413 8632
rect 26477 8688 26533 8697
rect 26477 8623 26533 8632
rect 19318 8528 19557 8574
rect 26027 8528 26266 8574
rect 13086 8510 13161 8514
rect 13086 8454 13096 8510
rect 13152 8454 13161 8510
rect 13086 8453 13161 8454
rect 13428 8464 13502 8468
rect 13428 8408 13437 8464
rect 13493 8408 13502 8464
rect 19511 8452 19557 8528
rect 20137 8464 20211 8468
rect 13428 8404 13502 8408
rect 19509 8451 19575 8452
rect 19509 8399 19515 8451
rect 19567 8399 19575 8451
rect 20137 8408 20146 8464
rect 20202 8408 20211 8464
rect 26220 8452 26266 8528
rect 20137 8404 20211 8408
rect 26218 8451 26284 8452
rect 26218 8399 26224 8451
rect 26276 8399 26284 8451
rect 13060 8358 13135 8362
rect 13060 8302 13070 8358
rect 13126 8302 13135 8358
rect 13060 8301 13135 8302
rect 13346 8222 13420 8226
rect 13346 8166 13355 8222
rect 13411 8166 13420 8222
rect 13346 8162 13420 8166
rect 20055 8222 20129 8226
rect 20055 8166 20064 8222
rect 20120 8166 20129 8222
rect 20055 8162 20129 8166
rect 19511 8142 19567 8151
rect 19511 8077 19567 8086
rect 19655 8143 19711 8152
rect 19655 8078 19711 8087
rect 19786 8142 19842 8151
rect 19786 8077 19842 8086
rect 26220 8142 26276 8151
rect 26220 8077 26276 8086
rect 26364 8143 26420 8152
rect 26364 8078 26420 8087
rect 26495 8142 26551 8151
rect 26495 8077 26551 8086
rect 13345 8065 13419 8069
rect 12911 7987 12919 8040
rect 12971 7987 12977 8040
rect 13345 8009 13354 8065
rect 13410 8009 13419 8065
rect 13345 8005 13419 8009
rect 20054 8065 20128 8069
rect 20054 8009 20063 8065
rect 20119 8009 20128 8065
rect 20054 8005 20128 8009
rect 12911 7986 12977 7987
rect 19632 7993 19706 7997
rect 19632 7937 19641 7993
rect 19697 7937 19706 7993
rect 12929 7931 13003 7935
rect 19632 7933 19706 7937
rect 12929 7875 12938 7931
rect 12994 7875 13003 7931
rect 12929 7871 13003 7875
rect 13345 7895 13419 7899
rect 11750 7849 11802 7855
rect 13345 7839 13354 7895
rect 13410 7839 13419 7895
rect 13345 7835 13419 7839
rect 20054 7895 20128 7899
rect 20054 7839 20063 7895
rect 20119 7839 20128 7895
rect 20054 7835 20128 7839
rect 11750 7790 11802 7797
rect 19632 7797 19706 7801
rect 11762 7532 11790 7790
rect 12209 7740 12283 7744
rect 11955 7736 12029 7740
rect 11955 7680 11964 7736
rect 12020 7680 12029 7736
rect 12209 7684 12218 7740
rect 12274 7684 12283 7740
rect 13346 7743 13420 7747
rect 12209 7680 12283 7684
rect 12921 7711 12995 7715
rect 11955 7676 12029 7680
rect 12921 7655 12930 7711
rect 12986 7655 12995 7711
rect 13346 7687 13355 7743
rect 13411 7687 13420 7743
rect 19632 7741 19641 7797
rect 19697 7741 19706 7797
rect 19632 7737 19706 7741
rect 20055 7743 20129 7747
rect 13346 7683 13420 7687
rect 20055 7687 20064 7743
rect 20120 7687 20129 7743
rect 20055 7683 20129 7687
rect 12921 7651 12995 7655
rect 19632 7622 19706 7626
rect 13351 7599 13425 7603
rect 11965 7591 12039 7595
rect 11965 7535 11974 7591
rect 12030 7535 12039 7591
rect 11743 7480 11749 7532
rect 11801 7480 11807 7532
rect 11965 7531 12039 7535
rect 12217 7594 12291 7598
rect 12217 7538 12226 7594
rect 12282 7538 12291 7594
rect 13351 7543 13360 7599
rect 13416 7543 13425 7599
rect 19632 7566 19641 7622
rect 19697 7566 19706 7622
rect 19632 7562 19706 7566
rect 20060 7599 20134 7603
rect 13351 7539 13425 7543
rect 13593 7543 18501 7549
rect 12217 7534 12291 7538
rect 13593 7487 13697 7543
rect 13753 7487 13777 7543
rect 13833 7487 13857 7543
rect 13913 7487 13937 7543
rect 13993 7487 14017 7543
rect 14073 7487 14097 7543
rect 14153 7487 14305 7543
rect 14361 7487 14385 7543
rect 14441 7487 14465 7543
rect 14521 7487 14545 7543
rect 14601 7487 14625 7543
rect 14681 7487 14705 7543
rect 14761 7487 14909 7543
rect 14965 7487 14989 7543
rect 15045 7487 15069 7543
rect 15125 7487 15149 7543
rect 15205 7487 15229 7543
rect 15285 7487 15309 7543
rect 15365 7487 15517 7543
rect 15573 7487 15597 7543
rect 15653 7487 15677 7543
rect 15733 7487 15757 7543
rect 15813 7487 15837 7543
rect 15893 7487 15917 7543
rect 15973 7487 16121 7543
rect 16177 7487 16201 7543
rect 16257 7487 16281 7543
rect 16337 7487 16361 7543
rect 16417 7487 16441 7543
rect 16497 7487 16521 7543
rect 16577 7487 16729 7543
rect 16785 7487 16809 7543
rect 16865 7487 16889 7543
rect 16945 7487 16969 7543
rect 17025 7487 17049 7543
rect 17105 7487 17129 7543
rect 17185 7487 17333 7543
rect 17389 7487 17413 7543
rect 17469 7487 17493 7543
rect 17549 7487 17573 7543
rect 17629 7487 17653 7543
rect 17709 7487 17733 7543
rect 17789 7487 17941 7543
rect 17997 7487 18021 7543
rect 18077 7487 18101 7543
rect 18157 7487 18181 7543
rect 18237 7487 18261 7543
rect 18317 7487 18341 7543
rect 18397 7487 18501 7543
rect 13593 7483 18501 7487
rect 18563 7546 19233 7552
rect 18563 7490 18673 7546
rect 18729 7490 18753 7546
rect 18809 7490 18833 7546
rect 18889 7490 18913 7546
rect 18969 7490 18993 7546
rect 19049 7490 19073 7546
rect 19129 7541 19233 7546
rect 20060 7543 20069 7599
rect 20125 7543 20134 7599
rect 19129 7537 19234 7541
rect 20060 7539 20134 7543
rect 20302 7543 25210 7549
rect 19129 7490 19169 7537
rect 18563 7486 19169 7490
rect 19160 7481 19169 7486
rect 19225 7481 19234 7537
rect 20302 7487 20406 7543
rect 20462 7487 20486 7543
rect 20542 7487 20566 7543
rect 20622 7487 20646 7543
rect 20702 7487 20726 7543
rect 20782 7487 20806 7543
rect 20862 7487 21014 7543
rect 21070 7487 21094 7543
rect 21150 7487 21174 7543
rect 21230 7487 21254 7543
rect 21310 7487 21334 7543
rect 21390 7487 21414 7543
rect 21470 7487 21618 7543
rect 21674 7487 21698 7543
rect 21754 7487 21778 7543
rect 21834 7487 21858 7543
rect 21914 7487 21938 7543
rect 21994 7487 22018 7543
rect 22074 7487 22226 7543
rect 22282 7487 22306 7543
rect 22362 7487 22386 7543
rect 22442 7487 22466 7543
rect 22522 7487 22546 7543
rect 22602 7487 22626 7543
rect 22682 7487 22830 7543
rect 22886 7487 22910 7543
rect 22966 7487 22990 7543
rect 23046 7487 23070 7543
rect 23126 7487 23150 7543
rect 23206 7487 23230 7543
rect 23286 7487 23438 7543
rect 23494 7487 23518 7543
rect 23574 7487 23598 7543
rect 23654 7487 23678 7543
rect 23734 7487 23758 7543
rect 23814 7487 23838 7543
rect 23894 7487 24042 7543
rect 24098 7487 24122 7543
rect 24178 7487 24202 7543
rect 24258 7487 24282 7543
rect 24338 7487 24362 7543
rect 24418 7487 24442 7543
rect 24498 7487 24650 7543
rect 24706 7487 24730 7543
rect 24786 7487 24810 7543
rect 24866 7487 24890 7543
rect 24946 7487 24970 7543
rect 25026 7487 25050 7543
rect 25106 7487 25210 7543
rect 20302 7483 25210 7487
rect 25272 7546 25942 7552
rect 25272 7490 25382 7546
rect 25438 7490 25462 7546
rect 25518 7490 25542 7546
rect 25598 7490 25622 7546
rect 25678 7490 25702 7546
rect 25758 7490 25782 7546
rect 25838 7541 25942 7546
rect 25838 7537 25943 7541
rect 25838 7490 25878 7537
rect 25272 7486 25878 7490
rect 19160 7477 19234 7481
rect 25869 7481 25878 7486
rect 25934 7481 25943 7537
rect 25869 7477 25943 7481
rect 10623 7282 10629 7334
rect 10681 7282 10687 7334
rect 10623 7281 10687 7282
rect 23915 7281 23921 7333
rect 23973 7281 23979 7333
rect 10311 5240 10363 5246
rect 10311 5182 10363 5188
rect 8498 2735 8505 2787
rect 8557 2735 8563 2787
rect 8498 2734 8563 2735
rect 8506 1216 8543 2734
rect 8626 1413 8682 1422
rect 8626 1348 8682 1357
rect 8489 1164 8497 1216
rect 8549 1164 8555 1216
rect 8592 269 8648 278
rect 8592 204 8648 213
rect 8592 -151 8646 -145
rect 8592 -203 8593 -151
rect 8645 -203 8646 -151
rect 8592 -209 8646 -203
rect 8598 -690 8640 -209
rect 8592 -696 8646 -690
rect 8592 -748 8593 -696
rect 8645 -748 8646 -696
rect 8592 -754 8646 -748
rect 8620 -1107 8676 -1098
rect 8620 -1172 8676 -1163
rect 8592 -1215 8644 -1209
rect 8716 -1219 8758 2925
rect 8798 1577 8840 2925
rect 8882 1647 8924 2925
rect 8970 1716 9012 2925
rect 9057 1786 9099 2925
rect 9143 1855 9185 2925
rect 9229 1925 9271 2925
rect 9316 1995 9358 2925
rect 9402 2065 9444 2925
rect 9488 2134 9530 2925
rect 9575 2204 9617 2925
rect 9660 2274 9702 2925
rect 9747 2343 9789 2925
rect 9834 2412 9876 2925
rect 9983 2924 9989 2976
rect 10041 2924 10047 2976
rect 10323 2783 10351 5182
rect 10642 4363 10670 7281
rect 23915 7280 23979 7281
rect 24670 7331 24744 7335
rect 10881 7080 11053 7090
rect 10881 6934 10891 7080
rect 11041 6934 11053 7080
rect 10881 6924 11053 6934
rect 11193 7064 11365 7074
rect 11193 6918 11203 7064
rect 11353 6918 11365 7064
rect 11193 6908 11365 6918
rect 18583 6809 18636 6816
rect 12153 6745 12160 6797
rect 12212 6745 12221 6797
rect 12193 6423 12221 6745
rect 12476 6796 12542 6797
rect 12476 6744 12483 6796
rect 12535 6744 12542 6796
rect 18635 6757 18636 6809
rect 18583 6750 18636 6757
rect 11516 6422 11582 6423
rect 11516 6370 11523 6422
rect 11575 6370 11582 6422
rect 12177 6422 12243 6423
rect 12177 6370 12184 6422
rect 12236 6370 12243 6422
rect 11251 6132 11423 6142
rect 10945 6120 11117 6130
rect 10945 5974 10955 6120
rect 11105 5974 11117 6120
rect 11251 5986 11261 6132
rect 11411 5986 11423 6132
rect 11251 5976 11423 5986
rect 10945 5964 11117 5974
rect 11534 5935 11562 6370
rect 12495 5992 12523 6744
rect 14059 6675 14065 6727
rect 14117 6675 14123 6727
rect 13907 6422 13973 6423
rect 13907 6370 13914 6422
rect 13966 6370 13973 6422
rect 12478 5940 12485 5992
rect 12537 5940 12544 5992
rect 11533 5910 11562 5935
rect 11515 5909 11581 5910
rect 11515 5857 11522 5909
rect 11574 5857 11581 5909
rect 10777 5492 10949 5502
rect 10777 5346 10787 5492
rect 10937 5346 10949 5492
rect 10777 5336 10949 5346
rect 11952 4806 11959 4858
rect 12011 4806 12018 4858
rect 10813 4646 10985 4656
rect 10813 4500 10823 4646
rect 10973 4500 10985 4646
rect 10813 4490 10985 4500
rect 11165 4650 11337 4660
rect 11165 4504 11175 4650
rect 11325 4504 11337 4650
rect 11165 4494 11337 4504
rect 11611 4650 11783 4660
rect 11611 4504 11621 4650
rect 11771 4504 11783 4650
rect 11611 4494 11783 4504
rect 10623 4311 10630 4363
rect 10682 4311 10688 4363
rect 11113 4303 11119 4355
rect 11171 4303 11177 4355
rect 11720 4303 11726 4355
rect 11778 4303 11784 4355
rect 11117 3988 11153 4303
rect 11103 3936 11109 3988
rect 11161 3936 11167 3988
rect 11734 3985 11770 4303
rect 11723 3933 11729 3985
rect 11781 3933 11787 3985
rect 10895 3792 11067 3802
rect 10895 3646 10905 3792
rect 11055 3646 11067 3792
rect 10895 3636 11067 3646
rect 11245 3800 11417 3810
rect 11245 3654 11255 3800
rect 11405 3654 11417 3800
rect 11245 3644 11417 3654
rect 11971 3488 11999 4806
rect 12177 4654 12349 4664
rect 12177 4508 12187 4654
rect 12337 4508 12349 4654
rect 12177 4498 12349 4508
rect 12495 4358 12523 5940
rect 13927 5910 13955 6370
rect 13905 5909 13971 5910
rect 13905 5857 13912 5909
rect 13964 5857 13971 5909
rect 12983 5854 13049 5855
rect 12983 5802 12990 5854
rect 13042 5802 13049 5854
rect 12998 5411 13031 5802
rect 13533 5796 13599 5797
rect 13533 5744 13540 5796
rect 13592 5744 13599 5796
rect 12990 5404 13043 5411
rect 12990 5352 12991 5404
rect 12990 5345 13043 5352
rect 12843 4654 13015 4664
rect 12843 4508 12853 4654
rect 13003 4508 13015 4654
rect 12843 4498 13015 4508
rect 13225 4638 13397 4648
rect 13225 4492 13235 4638
rect 13385 4492 13397 4638
rect 13225 4482 13397 4492
rect 13079 4431 13144 4432
rect 13078 4430 13144 4431
rect 13557 4430 13585 5744
rect 13899 5386 13905 5438
rect 13957 5431 13963 5438
rect 14071 5431 14104 6675
rect 14338 6613 14345 6665
rect 14397 6613 14404 6665
rect 16187 6613 16194 6665
rect 16246 6613 16253 6665
rect 14338 6612 14404 6613
rect 15749 5876 15756 5928
rect 15808 5876 15814 5928
rect 13957 5396 14104 5431
rect 13957 5386 13963 5396
rect 14351 5238 14404 5245
rect 14403 5186 14404 5238
rect 14351 5179 14404 5186
rect 13812 5100 13878 5101
rect 13812 5048 13819 5100
rect 13871 5048 13878 5100
rect 13832 4859 13860 5048
rect 14363 4859 14391 5179
rect 15768 4859 15796 5876
rect 16039 5821 16092 5828
rect 15923 5810 15987 5816
rect 15923 5758 15930 5810
rect 15982 5758 15987 5810
rect 16039 5769 16040 5821
rect 16039 5762 16092 5769
rect 15923 5757 15987 5758
rect 15923 5752 15986 5757
rect 13812 4858 13878 4859
rect 13812 4806 13819 4858
rect 13871 4806 13878 4858
rect 14344 4858 14410 4859
rect 14344 4806 14351 4858
rect 14403 4806 14410 4858
rect 15748 4858 15814 4859
rect 15748 4806 15755 4858
rect 15807 4806 15814 4858
rect 13078 4378 13085 4430
rect 13137 4378 13144 4430
rect 13523 4429 13589 4430
rect 12475 4357 12541 4358
rect 12475 4305 12482 4357
rect 12534 4305 12541 4357
rect 11951 3436 11961 3488
rect 12013 3436 12025 3488
rect 11951 3434 12025 3436
rect 13092 3421 13120 4378
rect 13523 4377 13530 4429
rect 13582 4377 13589 4429
rect 13463 3931 13470 3983
rect 13522 3931 13529 3983
rect 13483 3546 13511 3931
rect 13462 3494 13469 3546
rect 13521 3494 13528 3546
rect 14363 3501 14391 4806
rect 14644 4378 14652 4430
rect 14704 4378 14711 4430
rect 14657 4294 14685 4378
rect 15768 4366 15796 4806
rect 15756 4359 15809 4366
rect 15808 4307 15809 4359
rect 15756 4300 15809 4307
rect 14638 4293 14702 4294
rect 14638 4241 14644 4293
rect 14696 4241 14702 4293
rect 15843 3932 15850 3984
rect 15902 3932 15909 3984
rect 15863 3543 15891 3932
rect 14350 3494 14403 3501
rect 14350 3442 14351 3494
rect 15843 3491 15850 3543
rect 15902 3491 15909 3543
rect 14350 3435 14403 3442
rect 13075 3420 13141 3421
rect 13075 3368 13082 3420
rect 13134 3368 13141 3420
rect 13905 3384 13958 3391
rect 11514 3361 11567 3368
rect 11566 3309 11567 3361
rect 13957 3332 13958 3384
rect 15939 3353 15972 5752
rect 13905 3325 13958 3332
rect 11514 3302 11567 3309
rect 10303 2731 10310 2783
rect 10362 2731 10368 2783
rect 10303 2730 10368 2731
rect 11526 2690 11554 3302
rect 11905 2926 11911 2978
rect 11963 2926 11969 2978
rect 10529 2637 10535 2689
rect 10587 2637 10594 2689
rect 11521 2686 11555 2690
rect 10126 2568 10132 2620
rect 10184 2568 10191 2620
rect 9823 2360 9829 2412
rect 9881 2360 9887 2412
rect 9736 2291 9742 2343
rect 9794 2291 9800 2343
rect 9649 2222 9655 2274
rect 9707 2222 9713 2274
rect 9563 2152 9569 2204
rect 9621 2152 9627 2204
rect 9477 2082 9483 2134
rect 9535 2082 9541 2134
rect 9390 2013 9396 2065
rect 9448 2013 9454 2065
rect 9304 1943 9310 1995
rect 9362 1943 9368 1995
rect 9218 1873 9224 1925
rect 9276 1873 9282 1925
rect 9132 1803 9138 1855
rect 9190 1803 9196 1855
rect 9045 1734 9051 1786
rect 9103 1734 9109 1786
rect 8959 1664 8965 1716
rect 9017 1664 9023 1716
rect 8872 1595 8878 1647
rect 8930 1595 8936 1647
rect 8786 1525 8792 1577
rect 8844 1525 8850 1577
rect 8828 1415 8884 1424
rect 8828 1350 8884 1359
rect 9039 1413 9095 1422
rect 9039 1348 9095 1357
rect 9229 1413 9285 1422
rect 9229 1348 9285 1357
rect 9437 1415 9493 1424
rect 9437 1350 9493 1359
rect 9639 1415 9695 1424
rect 9639 1350 9695 1359
rect 9838 1417 9894 1426
rect 9838 1352 9894 1361
rect 10033 1414 10089 1423
rect 10033 1349 10089 1358
rect 9744 874 9800 883
rect 9744 809 9800 818
rect 9963 878 10019 887
rect 9963 813 10019 822
rect 9593 685 9599 738
rect 9652 685 9658 738
rect 9593 684 9658 685
rect 9042 474 9049 526
rect 9101 474 9108 526
rect 8832 267 8888 276
rect 8832 202 8888 211
rect 9057 52 9094 474
rect 9154 266 9210 275
rect 9154 201 9210 210
rect 9372 267 9428 276
rect 9372 202 9428 211
rect 9043 0 9050 52
rect 9102 0 9109 52
rect 8924 -165 8931 -113
rect 8983 -165 8989 -113
rect 8838 -414 8894 -405
rect 8838 -479 8894 -470
rect 8937 -671 8979 -165
rect 9040 -418 9096 -409
rect 9040 -483 9096 -474
rect 9229 -421 9285 -412
rect 9229 -486 9285 -477
rect 9458 -420 9514 -411
rect 9458 -485 9514 -476
rect 8926 -724 8932 -671
rect 8984 -724 8991 -671
rect 8926 -725 8991 -724
rect 9605 -789 9647 684
rect 10137 38 10179 2568
rect 10234 1416 10290 1425
rect 10234 1351 10290 1360
rect 10451 1414 10507 1423
rect 10451 1349 10507 1358
rect 10246 878 10302 887
rect 10246 813 10302 822
rect 10455 878 10511 887
rect 10455 813 10511 822
rect 10304 474 10311 526
rect 10363 474 10370 526
rect 10319 52 10356 474
rect 10126 -15 10132 38
rect 10184 -15 10191 38
rect 10305 0 10312 52
rect 10364 0 10371 52
rect 10126 -16 10191 -15
rect 10539 -112 10581 2637
rect 11509 2634 11515 2686
rect 11567 2634 11574 2686
rect 10893 1942 10899 1994
rect 10951 1942 10958 1994
rect 10725 1417 10781 1426
rect 10725 1352 10781 1361
rect 10726 876 10782 885
rect 10726 811 10782 820
rect 10525 -164 10532 -112
rect 10584 -164 10590 -112
rect 9783 -269 9839 -260
rect 9783 -334 9839 -325
rect 10000 -269 10056 -260
rect 10000 -334 10056 -325
rect 10219 -269 10275 -260
rect 10219 -334 10275 -325
rect 10432 -273 10488 -264
rect 10432 -338 10488 -329
rect 9599 -795 9653 -789
rect 9599 -847 9600 -795
rect 9652 -847 9653 -795
rect 9599 -853 9653 -847
rect 8853 -1111 8909 -1102
rect 8853 -1176 8909 -1167
rect 9068 -1104 9124 -1095
rect 9068 -1169 9124 -1160
rect 9286 -1107 9342 -1098
rect 9286 -1172 9342 -1163
rect 9502 -1106 9558 -1097
rect 9502 -1171 9558 -1162
rect 8644 -1261 8758 -1219
rect 9605 -1251 9647 -853
rect 9994 -951 10050 -942
rect 9765 -963 9821 -954
rect 9994 -1016 10050 -1007
rect 10213 -961 10269 -952
rect 9765 -1028 9821 -1019
rect 10213 -1026 10269 -1017
rect 10405 -957 10461 -948
rect 10405 -1022 10461 -1013
rect 8592 -1273 8644 -1267
rect 8872 -1279 8924 -1273
rect 9594 -1303 9600 -1251
rect 9652 -1303 9658 -1251
rect 8872 -1337 8924 -1331
rect 8876 -1908 8918 -1337
rect 10539 -1405 10581 -164
rect 10763 -203 10769 -151
rect 10821 -203 10829 -151
rect 10643 -273 10699 -264
rect 10643 -338 10699 -329
rect 10617 -600 10669 -594
rect 10617 -658 10669 -652
rect 10528 -1458 10534 -1405
rect 10586 -1458 10593 -1405
rect 10528 -1459 10593 -1458
rect 8994 -1639 9050 -1630
rect 8994 -1704 9050 -1695
rect 9193 -1642 9249 -1633
rect 9193 -1707 9249 -1698
rect 9404 -1642 9460 -1633
rect 9404 -1707 9460 -1698
rect 9610 -1642 9666 -1633
rect 9610 -1707 9666 -1698
rect 9838 -1644 9894 -1635
rect 9838 -1709 9894 -1700
rect 10082 -1644 10138 -1635
rect 10082 -1709 10138 -1700
rect 10312 -1642 10368 -1633
rect 10312 -1707 10368 -1698
rect 10518 -1642 10574 -1633
rect 10518 -1707 10574 -1698
rect 10621 -1908 10663 -658
rect 10775 -1350 10817 -203
rect 10905 -517 10947 1942
rect 11108 1575 11150 1735
rect 11098 1523 11104 1575
rect 11156 1523 11163 1575
rect 11002 1410 11058 1419
rect 11002 1345 11058 1354
rect 10984 -151 11038 -145
rect 10984 -203 10985 -151
rect 11037 -203 11038 -151
rect 10984 -209 11038 -203
rect 10899 -523 10951 -517
rect 10899 -581 10951 -575
rect 10990 -690 11032 -209
rect 10984 -696 11038 -690
rect 10984 -748 10985 -696
rect 11037 -748 11038 -696
rect 10984 -754 11038 -748
rect 10899 -959 10955 -950
rect 10899 -1024 10955 -1015
rect 10984 -1215 11036 -1209
rect 11108 -1219 11150 1523
rect 11225 1413 11281 1422
rect 11225 1348 11281 1357
rect 11457 1412 11513 1421
rect 11457 1347 11513 1356
rect 11435 1057 11441 1109
rect 11493 1057 11499 1109
rect 11441 737 11493 1057
rect 11922 1019 11950 2926
rect 12518 2904 12524 2956
rect 12576 2904 12583 2956
rect 12529 2703 12571 2904
rect 13917 2752 13945 3325
rect 15923 3301 15929 3353
rect 15981 3301 15987 3353
rect 15939 3298 15972 3301
rect 14907 3096 14914 3148
rect 14966 3096 14972 3148
rect 12528 1703 12571 2703
rect 12922 2700 12928 2752
rect 12980 2700 12987 2752
rect 13898 2700 13904 2752
rect 13956 2700 13963 2752
rect 11910 967 11916 1019
rect 11968 967 11974 1019
rect 11435 685 11441 737
rect 11493 685 11499 737
rect 11987 691 11993 744
rect 12046 691 12052 744
rect 11987 690 12052 691
rect 11435 473 11442 525
rect 11494 473 11501 525
rect 11276 271 11332 280
rect 11276 206 11332 215
rect 11450 51 11487 473
rect 11601 273 11657 282
rect 11601 208 11657 217
rect 11869 273 11925 282
rect 11869 208 11925 217
rect 11436 -1 11443 51
rect 11495 -1 11502 51
rect 11316 -165 11323 -113
rect 11375 -165 11381 -113
rect 11227 -417 11283 -408
rect 11227 -482 11283 -473
rect 11329 -671 11371 -165
rect 11442 -420 11498 -411
rect 11835 -413 11891 -404
rect 11442 -485 11498 -476
rect 11640 -423 11696 -414
rect 11835 -478 11891 -469
rect 11640 -488 11696 -479
rect 11318 -724 11324 -671
rect 11376 -724 11383 -671
rect 11318 -725 11383 -724
rect 11999 -789 12041 690
rect 12135 273 12191 282
rect 12135 208 12191 217
rect 12375 271 12431 280
rect 12375 206 12431 215
rect 12529 37 12571 1703
rect 12801 874 12857 883
rect 12801 809 12857 818
rect 12696 474 12703 526
rect 12755 474 12762 526
rect 12711 52 12748 474
rect 12518 -16 12524 37
rect 12576 -16 12583 37
rect 12697 0 12704 52
rect 12756 0 12763 52
rect 12518 -17 12583 -16
rect 12931 -112 12973 2700
rect 13913 2656 13947 2700
rect 13917 2654 13945 2656
rect 13285 2012 13291 2064
rect 13343 2012 13350 2064
rect 13093 1409 13149 1418
rect 13093 1344 13149 1353
rect 13050 877 13106 886
rect 13050 812 13106 821
rect 12917 -164 12924 -112
rect 12976 -164 12982 -112
rect 12767 -273 12823 -264
rect 12767 -338 12823 -329
rect 12115 -415 12171 -406
rect 12115 -480 12171 -471
rect 12334 -417 12390 -408
rect 12334 -482 12390 -473
rect 11992 -795 12046 -789
rect 11992 -847 11993 -795
rect 12045 -847 12046 -795
rect 11992 -853 12046 -847
rect 11223 -1110 11279 -1101
rect 11223 -1175 11279 -1166
rect 11413 -1110 11469 -1101
rect 11413 -1175 11469 -1166
rect 11623 -1107 11679 -1098
rect 11623 -1172 11679 -1163
rect 11840 -1110 11896 -1101
rect 11840 -1175 11896 -1166
rect 11036 -1261 11150 -1219
rect 11997 -1250 12039 -853
rect 12691 -960 12747 -951
rect 12691 -1025 12747 -1016
rect 12135 -1107 12191 -1098
rect 12135 -1172 12191 -1163
rect 12359 -1102 12415 -1093
rect 12359 -1167 12415 -1158
rect 10984 -1273 11036 -1267
rect 11264 -1279 11316 -1273
rect 11986 -1302 11992 -1250
rect 12044 -1302 12050 -1250
rect 11264 -1337 11316 -1331
rect 10775 -1390 10879 -1350
rect 10873 -1402 10879 -1390
rect 10933 -1402 10939 -1350
rect 10736 -1637 10792 -1628
rect 10736 -1702 10792 -1693
rect 10939 -1643 10995 -1634
rect 10939 -1708 10995 -1699
rect 11147 -1640 11203 -1631
rect 11147 -1705 11203 -1696
rect 11268 -1908 11310 -1337
rect 12931 -1405 12973 -164
rect 13157 -203 13163 -151
rect 13215 -203 13223 -151
rect 13045 -274 13101 -265
rect 13045 -339 13101 -330
rect 13009 -599 13061 -593
rect 13009 -657 13061 -651
rect 12920 -1458 12926 -1405
rect 12978 -1458 12985 -1405
rect 12920 -1459 12985 -1458
rect 11410 -1644 11466 -1635
rect 11410 -1709 11466 -1700
rect 11618 -1643 11674 -1634
rect 11618 -1708 11674 -1699
rect 11828 -1646 11884 -1637
rect 11828 -1711 11884 -1702
rect 12028 -1640 12084 -1631
rect 12028 -1705 12084 -1696
rect 12231 -1643 12287 -1634
rect 12231 -1708 12287 -1699
rect 12441 -1643 12497 -1634
rect 12441 -1708 12497 -1699
rect 12642 -1642 12698 -1633
rect 12642 -1707 12698 -1698
rect 12858 -1641 12914 -1632
rect 12858 -1706 12914 -1697
rect 13013 -1908 13055 -657
rect 13084 -962 13140 -953
rect 13084 -1027 13140 -1018
rect 13169 -1350 13211 -203
rect 13297 -517 13339 2012
rect 13501 1646 13543 1735
rect 13488 1594 13494 1646
rect 13546 1594 13553 1646
rect 13401 1410 13457 1419
rect 13401 1345 13457 1354
rect 13394 863 13450 872
rect 13394 798 13450 807
rect 13376 -151 13430 -145
rect 13376 -203 13377 -151
rect 13429 -203 13430 -151
rect 13376 -209 13430 -203
rect 13291 -523 13343 -517
rect 13291 -581 13343 -575
rect 13382 -690 13424 -209
rect 13376 -696 13430 -690
rect 13376 -748 13377 -696
rect 13429 -748 13430 -696
rect 13376 -754 13430 -748
rect 13281 -954 13337 -945
rect 13281 -1019 13337 -1010
rect 13377 -1215 13429 -1209
rect 13501 -1219 13543 1594
rect 13601 1411 13657 1420
rect 13601 1346 13657 1355
rect 13820 1410 13876 1419
rect 13820 1345 13876 1354
rect 14066 1409 14122 1418
rect 14066 1344 14122 1353
rect 14274 1411 14330 1420
rect 14274 1346 14330 1355
rect 14476 1412 14532 1421
rect 14476 1347 14532 1356
rect 14669 1411 14725 1420
rect 14669 1346 14725 1355
rect 13648 869 13704 878
rect 13648 804 13704 813
rect 13877 869 13933 878
rect 13877 804 13933 813
rect 14378 691 14384 744
rect 14437 691 14443 744
rect 14378 690 14443 691
rect 13827 473 13834 525
rect 13886 473 13893 525
rect 13842 51 13879 473
rect 14169 274 14225 283
rect 14169 209 14225 218
rect 13828 -1 13835 51
rect 13887 -1 13894 51
rect 13707 -164 13714 -112
rect 13766 -164 13772 -112
rect 13617 -269 13673 -260
rect 13617 -334 13673 -325
rect 13721 -670 13763 -164
rect 13856 -269 13912 -260
rect 13856 -334 13912 -325
rect 14155 -420 14211 -411
rect 14155 -485 14211 -476
rect 13710 -723 13716 -670
rect 13768 -723 13775 -670
rect 13710 -724 13775 -723
rect 14390 -789 14432 690
rect 14535 277 14591 286
rect 14535 212 14591 221
rect 14779 277 14835 286
rect 14779 212 14835 221
rect 14919 37 14961 3096
rect 15309 2824 15316 2876
rect 15368 2824 15374 2876
rect 15041 1410 15097 1419
rect 15041 1345 15097 1354
rect 15230 1408 15286 1417
rect 15230 1343 15286 1352
rect 15087 475 15094 527
rect 15146 475 15153 527
rect 15102 288 15139 475
rect 15096 254 15139 288
rect 15102 53 15139 254
rect 15202 268 15258 277
rect 15202 203 15258 212
rect 14908 -16 14914 37
rect 14966 -16 14973 37
rect 15088 1 15095 53
rect 15147 1 15154 53
rect 14908 -17 14973 -16
rect 15322 -111 15364 2824
rect 16052 2688 16080 5762
rect 16202 5296 16235 6613
rect 16290 6422 16356 6423
rect 16290 6370 16297 6422
rect 16349 6370 16356 6422
rect 16310 5911 16338 6370
rect 18149 5927 18202 5934
rect 16298 5910 16364 5911
rect 16298 5858 16305 5910
rect 16357 5858 16364 5910
rect 18201 5875 18202 5927
rect 18149 5868 18202 5875
rect 16310 5421 16338 5858
rect 16296 5420 16362 5421
rect 16296 5368 16303 5420
rect 16355 5368 16362 5420
rect 16296 5303 16349 5310
rect 16296 5296 16297 5303
rect 16202 5262 16297 5296
rect 16296 5251 16297 5262
rect 16296 5244 16349 5251
rect 16746 5239 16799 5246
rect 16798 5187 16799 5239
rect 16746 5180 16799 5187
rect 16439 5135 16492 5142
rect 16491 5083 16492 5135
rect 16439 5076 16492 5083
rect 16296 3383 16349 3390
rect 16348 3331 16349 3383
rect 16296 3324 16349 3331
rect 16308 2877 16336 3324
rect 16296 2825 16302 2877
rect 16354 2825 16360 2877
rect 16308 2688 16336 2825
rect 16049 2614 16083 2688
rect 16307 2654 16341 2688
rect 16451 2685 16479 5076
rect 16755 4859 16783 5180
rect 17030 5099 17096 5100
rect 17030 5047 17037 5099
rect 17089 5047 17096 5099
rect 16733 4858 16799 4859
rect 16733 4806 16740 4858
rect 16792 4806 16799 4858
rect 16647 4311 16654 4363
rect 16706 4311 16713 4363
rect 16660 3983 16688 4311
rect 16642 3931 16649 3983
rect 16701 3931 16708 3983
rect 16755 3499 16783 4806
rect 17047 4293 17075 5047
rect 18160 4859 18188 5868
rect 18313 5766 18319 5818
rect 18371 5766 18377 5818
rect 18313 5758 18377 5766
rect 18435 5810 18488 5817
rect 18435 5758 18436 5810
rect 18140 4858 18206 4859
rect 18140 4806 18147 4858
rect 18199 4806 18206 4858
rect 18160 4376 18188 4806
rect 18147 4369 18200 4376
rect 18199 4317 18200 4369
rect 18147 4310 18200 4317
rect 17031 4292 17097 4293
rect 17031 4240 17038 4292
rect 17090 4240 17097 4292
rect 18236 3931 18243 3983
rect 18295 3931 18302 3983
rect 18256 3547 18284 3931
rect 16744 3492 16797 3499
rect 18234 3495 18241 3547
rect 18293 3495 18300 3547
rect 16796 3440 16797 3492
rect 16744 3433 16797 3440
rect 18330 3353 18363 5758
rect 18435 5751 18488 5758
rect 18315 3301 18321 3353
rect 18373 3301 18379 3353
rect 18448 2954 18476 5751
rect 18592 5296 18625 6750
rect 20991 6733 21044 6740
rect 21043 6681 21044 6733
rect 20991 6674 21044 6681
rect 18685 6422 18751 6423
rect 18685 6370 18692 6422
rect 18744 6370 18751 6422
rect 18705 5910 18733 6370
rect 20540 5929 20593 5936
rect 18690 5909 18756 5910
rect 18690 5857 18697 5909
rect 18749 5857 18756 5909
rect 20592 5877 20593 5929
rect 20540 5870 20593 5877
rect 18705 5421 18733 5857
rect 18687 5420 18753 5421
rect 18687 5368 18694 5420
rect 18746 5368 18753 5420
rect 18684 5301 18737 5308
rect 18684 5296 18685 5301
rect 18592 5262 18685 5296
rect 18593 5261 18685 5262
rect 18684 5249 18685 5261
rect 18684 5242 18737 5249
rect 19136 5240 19189 5247
rect 19188 5188 19189 5240
rect 19136 5181 19189 5188
rect 18861 5124 18914 5131
rect 18913 5072 18914 5124
rect 18861 5065 18914 5072
rect 18604 4261 18657 4268
rect 18656 4209 18657 4261
rect 18604 4202 18657 4209
rect 18616 3086 18644 4202
rect 18691 3386 18744 3393
rect 18743 3334 18744 3386
rect 18691 3327 18744 3334
rect 18599 3018 18605 3086
rect 18657 3018 18663 3086
rect 18429 2902 18435 2954
rect 18487 2902 18494 2954
rect 17701 2756 17708 2808
rect 17760 2756 17766 2808
rect 16033 2562 16039 2614
rect 16091 2562 16097 2614
rect 16449 2613 16483 2685
rect 16434 2561 16440 2613
rect 16492 2561 16498 2613
rect 17301 2496 17307 2548
rect 17359 2496 17366 2548
rect 15679 2081 15685 2133
rect 15737 2081 15744 2133
rect 15520 1408 15576 1417
rect 15520 1343 15576 1352
rect 15595 874 15651 883
rect 15595 809 15651 818
rect 15308 -163 15315 -111
rect 15367 -163 15373 -111
rect 14506 -423 14562 -414
rect 14506 -488 14562 -479
rect 14695 -425 14751 -416
rect 14695 -490 14751 -481
rect 14900 -418 14956 -409
rect 14900 -483 14956 -474
rect 15091 -416 15147 -407
rect 15091 -481 15147 -472
rect 14384 -795 14438 -789
rect 14384 -847 14385 -795
rect 14437 -847 14438 -795
rect 14384 -853 14438 -847
rect 13611 -952 13667 -943
rect 13611 -1017 13667 -1008
rect 13807 -952 13863 -943
rect 13807 -1017 13863 -1008
rect 14237 -1109 14293 -1100
rect 14237 -1174 14293 -1165
rect 13429 -1261 13543 -1219
rect 14389 -1251 14431 -853
rect 14537 -1111 14593 -1102
rect 14537 -1176 14593 -1167
rect 14789 -1107 14845 -1098
rect 14789 -1172 14845 -1163
rect 15006 -1102 15062 -1093
rect 15006 -1167 15062 -1158
rect 15207 -1105 15263 -1096
rect 15207 -1170 15263 -1161
rect 13377 -1273 13429 -1267
rect 13655 -1279 13707 -1273
rect 14378 -1303 14384 -1251
rect 14436 -1303 14442 -1251
rect 13655 -1337 13707 -1331
rect 13169 -1390 13273 -1350
rect 13267 -1402 13273 -1390
rect 13327 -1402 13333 -1350
rect 13139 -1643 13195 -1634
rect 13139 -1708 13195 -1699
rect 13359 -1648 13415 -1639
rect 13359 -1713 13415 -1704
rect 13564 -1647 13620 -1638
rect 13564 -1712 13620 -1703
rect 13659 -1908 13701 -1337
rect 15322 -1404 15364 -163
rect 15547 -201 15553 -149
rect 15605 -201 15613 -149
rect 15400 -599 15452 -593
rect 15400 -657 15452 -651
rect 15311 -1405 15376 -1404
rect 15311 -1457 15317 -1405
rect 15369 -1457 15376 -1405
rect 15311 -1458 15376 -1457
rect 13785 -1641 13841 -1632
rect 13785 -1706 13841 -1697
rect 13990 -1648 14046 -1639
rect 13990 -1713 14046 -1704
rect 14199 -1647 14255 -1638
rect 14199 -1712 14255 -1703
rect 14416 -1647 14472 -1638
rect 14416 -1712 14472 -1703
rect 14630 -1642 14686 -1633
rect 14630 -1707 14686 -1698
rect 14825 -1644 14881 -1635
rect 14825 -1709 14881 -1700
rect 15020 -1647 15076 -1638
rect 15020 -1712 15076 -1703
rect 15222 -1644 15278 -1635
rect 15222 -1709 15278 -1700
rect 15404 -1908 15446 -657
rect 15559 -1348 15601 -201
rect 15689 -517 15731 2081
rect 15892 1715 15934 1735
rect 15880 1663 15886 1715
rect 15938 1663 15945 1715
rect 15793 1410 15849 1419
rect 15793 1345 15849 1354
rect 15799 876 15855 885
rect 15799 811 15855 820
rect 15768 -151 15822 -145
rect 15768 -203 15769 -151
rect 15821 -203 15822 -151
rect 15768 -209 15822 -203
rect 15683 -523 15735 -517
rect 15683 -581 15735 -575
rect 15774 -690 15816 -209
rect 15768 -696 15822 -690
rect 15768 -748 15769 -696
rect 15821 -748 15822 -696
rect 15768 -754 15822 -748
rect 15714 -959 15770 -950
rect 15714 -1024 15770 -1015
rect 15768 -1215 15820 -1209
rect 15892 -1219 15934 1663
rect 15996 1057 16002 1109
rect 16054 1057 16060 1109
rect 16002 525 16054 1057
rect 16122 874 16178 883
rect 16122 809 16178 818
rect 16769 691 16775 744
rect 16828 691 16834 744
rect 16769 690 16834 691
rect 15996 473 16002 525
rect 16054 473 16060 525
rect 16219 474 16226 526
rect 16278 474 16285 526
rect 16234 52 16271 474
rect 16220 0 16227 52
rect 16279 0 16286 52
rect 16100 -165 16107 -113
rect 16159 -165 16165 -113
rect 16014 -271 16070 -262
rect 16014 -336 16070 -327
rect 16113 -670 16155 -165
rect 16241 -266 16297 -257
rect 16241 -331 16297 -322
rect 16431 -264 16487 -255
rect 16431 -329 16487 -320
rect 16647 -273 16703 -264
rect 16647 -338 16703 -329
rect 16102 -723 16108 -670
rect 16160 -723 16167 -670
rect 16102 -724 16167 -723
rect 16781 -789 16823 690
rect 17145 270 17201 279
rect 17145 205 17201 214
rect 17313 38 17355 2496
rect 17480 475 17487 527
rect 17539 475 17546 527
rect 17397 267 17453 276
rect 17397 202 17453 211
rect 17495 53 17532 475
rect 17603 275 17659 284
rect 17603 210 17659 219
rect 17302 -15 17308 38
rect 17360 -15 17367 38
rect 17481 1 17488 53
rect 17540 1 17547 53
rect 17302 -16 17367 -15
rect 17715 -112 17757 2756
rect 18448 2690 18476 2902
rect 18616 2804 18644 3018
rect 18703 2808 18731 3327
rect 18614 2770 18648 2804
rect 18445 2656 18479 2690
rect 18448 2654 18476 2656
rect 18616 2654 18644 2770
rect 18685 2756 18691 2808
rect 18743 2756 18750 2808
rect 18701 2716 18735 2756
rect 18703 2654 18731 2716
rect 18873 2685 18901 5065
rect 19147 4859 19175 5181
rect 19422 5100 19488 5101
rect 19422 5048 19429 5100
rect 19481 5048 19488 5100
rect 19123 4858 19189 4859
rect 19123 4806 19130 4858
rect 19182 4806 19189 4858
rect 19034 4311 19041 4363
rect 19093 4311 19100 4363
rect 19049 3984 19077 4311
rect 19031 3932 19038 3984
rect 19090 3932 19097 3984
rect 19147 3500 19175 4806
rect 19440 4292 19468 5048
rect 20552 4859 20580 5870
rect 20835 5826 20888 5833
rect 20715 5795 20768 5802
rect 20767 5743 20768 5795
rect 20835 5774 20836 5826
rect 20835 5767 20888 5774
rect 20715 5736 20768 5743
rect 20537 4858 20603 4859
rect 20537 4806 20544 4858
rect 20596 4806 20603 4858
rect 20552 4372 20580 4806
rect 20538 4365 20591 4372
rect 20590 4313 20591 4365
rect 20538 4306 20591 4313
rect 19425 4291 19491 4292
rect 19425 4239 19432 4291
rect 19484 4239 19491 4291
rect 20623 3931 20630 3983
rect 20682 3931 20689 3983
rect 20643 3548 20671 3931
rect 19136 3493 19189 3500
rect 20623 3496 20630 3548
rect 20682 3496 20689 3548
rect 19188 3441 19189 3493
rect 19136 3434 19189 3441
rect 20722 3353 20755 5736
rect 20707 3301 20713 3353
rect 20765 3301 20771 3353
rect 20848 3149 20876 5767
rect 21000 5297 21033 6674
rect 23599 6466 23771 6476
rect 21080 6422 21146 6423
rect 21080 6370 21087 6422
rect 21139 6370 21146 6422
rect 23376 6422 23442 6423
rect 23376 6370 23383 6422
rect 23435 6370 23442 6422
rect 21100 5912 21128 6370
rect 23020 6117 23085 6122
rect 23020 6065 23026 6117
rect 23078 6065 23085 6117
rect 23020 6055 23085 6065
rect 22931 5927 22984 5934
rect 21085 5911 21151 5912
rect 21085 5859 21092 5911
rect 21144 5859 21151 5911
rect 22983 5875 22984 5927
rect 22931 5868 22984 5875
rect 21100 5417 21128 5859
rect 21081 5411 21134 5417
rect 21081 5359 21082 5411
rect 21081 5351 21134 5359
rect 21076 5302 21129 5309
rect 21076 5297 21077 5302
rect 21000 5263 21077 5297
rect 21076 5250 21077 5263
rect 21076 5243 21129 5250
rect 21530 5237 21583 5244
rect 21582 5185 21583 5237
rect 21530 5178 21583 5185
rect 21249 5132 21302 5139
rect 21301 5080 21302 5132
rect 21249 5073 21302 5080
rect 20996 4262 21049 4269
rect 21048 4210 21049 4262
rect 20996 4203 21049 4210
rect 21008 3149 21036 4203
rect 21080 3384 21133 3391
rect 21132 3332 21133 3384
rect 21080 3325 21133 3332
rect 20834 3097 20840 3149
rect 20892 3097 20898 3149
rect 20996 3097 21002 3149
rect 21054 3097 21060 3149
rect 19695 2961 19701 3013
rect 19753 2961 19759 3013
rect 18869 2481 18903 2685
rect 18857 2429 18863 2481
rect 18915 2429 18922 2481
rect 18070 2151 18076 2203
rect 18128 2151 18135 2203
rect 17886 269 17942 278
rect 17886 204 17942 213
rect 17701 -164 17708 -112
rect 17760 -164 17766 -112
rect 17136 -414 17192 -405
rect 17136 -479 17192 -470
rect 17326 -412 17382 -403
rect 17326 -477 17382 -468
rect 17520 -414 17576 -405
rect 17520 -479 17576 -470
rect 16776 -795 16830 -789
rect 16776 -847 16777 -795
rect 16829 -847 16830 -795
rect 16776 -853 16830 -847
rect 16015 -955 16071 -946
rect 16015 -1020 16071 -1011
rect 16221 -954 16277 -945
rect 16221 -1019 16277 -1010
rect 16431 -958 16487 -949
rect 16431 -1023 16487 -1014
rect 16642 -952 16698 -943
rect 16642 -1017 16698 -1008
rect 15820 -1261 15934 -1219
rect 16781 -1251 16823 -853
rect 17092 -1114 17148 -1105
rect 17092 -1179 17148 -1170
rect 17284 -1114 17340 -1105
rect 17284 -1179 17340 -1170
rect 17484 -1114 17540 -1105
rect 17484 -1179 17540 -1170
rect 15768 -1273 15820 -1267
rect 16048 -1279 16100 -1273
rect 16770 -1303 16776 -1251
rect 16828 -1303 16834 -1251
rect 16048 -1337 16100 -1331
rect 15559 -1388 15663 -1348
rect 15657 -1400 15663 -1388
rect 15717 -1400 15723 -1348
rect 15506 -1643 15562 -1634
rect 15506 -1708 15562 -1699
rect 15705 -1642 15761 -1633
rect 15705 -1707 15761 -1698
rect 15908 -1640 15964 -1631
rect 15908 -1705 15964 -1696
rect 16052 -1908 16094 -1337
rect 17715 -1405 17757 -164
rect 17939 -203 17945 -151
rect 17997 -203 18005 -151
rect 17831 -418 17887 -409
rect 17831 -483 17887 -474
rect 17793 -598 17845 -592
rect 17793 -656 17845 -650
rect 17704 -1458 17710 -1405
rect 17762 -1458 17769 -1405
rect 17704 -1459 17769 -1458
rect 16173 -1643 16229 -1634
rect 16173 -1708 16229 -1699
rect 16371 -1644 16427 -1635
rect 16371 -1709 16427 -1700
rect 16560 -1642 16616 -1633
rect 16560 -1707 16616 -1698
rect 16772 -1642 16828 -1633
rect 16772 -1707 16828 -1698
rect 16989 -1642 17045 -1633
rect 16989 -1707 17045 -1698
rect 17194 -1646 17250 -1637
rect 17194 -1711 17250 -1702
rect 17399 -1646 17455 -1637
rect 17399 -1711 17455 -1702
rect 17607 -1641 17663 -1632
rect 17607 -1706 17663 -1697
rect 17797 -1908 17839 -656
rect 17951 -1350 17993 -203
rect 18081 -517 18123 2151
rect 18273 1733 18279 1785
rect 18331 1733 18338 1785
rect 18184 270 18240 279
rect 18184 205 18240 214
rect 18159 -150 18213 -144
rect 18159 -202 18160 -150
rect 18212 -202 18213 -150
rect 18159 -208 18213 -202
rect 18075 -523 18127 -517
rect 18075 -581 18127 -575
rect 18165 -689 18207 -208
rect 18159 -695 18213 -689
rect 18159 -747 18160 -695
rect 18212 -747 18213 -695
rect 18159 -753 18213 -747
rect 18102 -1106 18158 -1097
rect 18102 -1171 18158 -1162
rect 18160 -1216 18212 -1210
rect 18284 -1220 18326 1733
rect 19161 691 19167 744
rect 19220 691 19226 744
rect 19161 690 19226 691
rect 18610 473 18617 525
rect 18669 473 18676 525
rect 18625 51 18662 473
rect 18611 -1 18618 51
rect 18670 -1 18677 51
rect 18492 -164 18499 -112
rect 18551 -164 18557 -112
rect 18505 -671 18547 -164
rect 18628 -270 18684 -261
rect 18628 -335 18684 -326
rect 18857 -267 18913 -258
rect 18857 -332 18913 -323
rect 19083 -262 19139 -253
rect 19083 -327 19139 -318
rect 18494 -724 18500 -671
rect 18552 -724 18559 -671
rect 18494 -725 18559 -724
rect 19173 -789 19215 690
rect 19705 37 19747 2961
rect 20092 2892 20099 2944
rect 20151 2892 20157 2944
rect 19873 475 19880 527
rect 19932 475 19939 527
rect 19888 53 19925 475
rect 20016 271 20072 280
rect 20016 206 20072 215
rect 19694 -16 19700 37
rect 19752 -16 19759 37
rect 19874 1 19881 53
rect 19933 1 19940 53
rect 19694 -17 19759 -16
rect 20106 -111 20148 2892
rect 20848 2685 20876 3097
rect 21008 2776 21036 3097
rect 21092 2944 21120 3325
rect 21261 3013 21289 5073
rect 21539 4859 21567 5178
rect 21811 5101 21877 5102
rect 21811 5049 21818 5101
rect 21870 5049 21877 5101
rect 21513 4858 21579 4859
rect 21513 4806 21520 4858
rect 21572 4806 21579 4858
rect 21437 4310 21444 4362
rect 21496 4310 21503 4362
rect 21458 3984 21486 4310
rect 21440 3932 21447 3984
rect 21499 3932 21506 3984
rect 21539 3501 21567 4806
rect 21832 4293 21860 5049
rect 22944 4859 22972 5868
rect 23038 5294 23071 6055
rect 23396 6054 23424 6370
rect 23599 6320 23609 6466
rect 23759 6320 23771 6466
rect 23599 6310 23771 6320
rect 23230 5826 23283 5833
rect 23106 5796 23159 5803
rect 23158 5744 23159 5796
rect 23230 5774 23231 5826
rect 23230 5767 23283 5774
rect 23106 5737 23159 5744
rect 23023 5242 23029 5294
rect 23081 5242 23087 5294
rect 22925 4858 22991 4859
rect 22925 4806 22932 4858
rect 22984 4806 22991 4858
rect 22944 4371 22972 4806
rect 22930 4364 22983 4371
rect 22982 4312 22983 4364
rect 22930 4305 22983 4312
rect 21811 4292 21877 4293
rect 21811 4240 21818 4292
rect 21870 4240 21877 4292
rect 23018 3932 23025 3984
rect 23077 3932 23084 3984
rect 23038 3548 23066 3932
rect 21529 3494 21582 3501
rect 23017 3496 23024 3548
rect 23076 3496 23083 3548
rect 21581 3442 21582 3494
rect 21529 3435 21582 3442
rect 23115 3353 23148 5737
rect 23098 3301 23104 3353
rect 23156 3301 23162 3353
rect 21245 2961 21251 3013
rect 21303 2961 21309 3013
rect 22486 2961 22493 3013
rect 22545 2961 22551 3013
rect 21076 2892 21082 2944
rect 21134 2892 21140 2944
rect 21092 2776 21120 2892
rect 21007 2742 21041 2776
rect 21090 2742 21124 2776
rect 20845 2651 20879 2685
rect 21008 2654 21036 2742
rect 21092 2654 21120 2742
rect 21261 2688 21289 2961
rect 21258 2654 21292 2688
rect 22083 2429 22089 2481
rect 22141 2429 22147 2481
rect 20462 2219 20468 2271
rect 20520 2219 20527 2271
rect 20226 273 20282 282
rect 20226 208 20282 217
rect 20093 -163 20100 -111
rect 20152 -163 20158 -111
rect 19311 -270 19367 -261
rect 19311 -335 19367 -326
rect 19547 -264 19603 -255
rect 19547 -329 19603 -320
rect 19739 -273 19795 -264
rect 19739 -338 19795 -329
rect 20014 -419 20070 -410
rect 20014 -484 20070 -475
rect 19167 -795 19221 -789
rect 19167 -847 19168 -795
rect 19220 -847 19221 -795
rect 19167 -855 19221 -847
rect 18522 -963 18578 -954
rect 18522 -1028 18578 -1019
rect 18779 -956 18835 -947
rect 18779 -1021 18835 -1012
rect 19029 -960 19085 -951
rect 19029 -1025 19085 -1016
rect 18212 -1262 18326 -1220
rect 19173 -1251 19215 -855
rect 19300 -955 19356 -946
rect 19300 -1020 19356 -1011
rect 19541 -952 19597 -943
rect 19541 -1017 19597 -1008
rect 19766 -956 19822 -947
rect 19766 -1021 19822 -1012
rect 20003 -1110 20059 -1101
rect 20003 -1175 20059 -1166
rect 18160 -1274 18212 -1268
rect 18440 -1279 18492 -1273
rect 19162 -1303 19168 -1251
rect 19220 -1303 19226 -1251
rect 18440 -1337 18492 -1331
rect 17951 -1390 18055 -1350
rect 18049 -1402 18055 -1390
rect 18109 -1402 18115 -1350
rect 17890 -1642 17946 -1633
rect 17890 -1707 17946 -1698
rect 18083 -1644 18139 -1635
rect 18083 -1709 18139 -1700
rect 18309 -1646 18365 -1637
rect 18309 -1711 18365 -1702
rect 18444 -1908 18486 -1337
rect 20106 -1405 20148 -163
rect 20331 -201 20337 -149
rect 20389 -201 20397 -149
rect 20218 -419 20274 -410
rect 20218 -484 20274 -475
rect 20184 -599 20236 -593
rect 20184 -657 20236 -651
rect 20095 -1458 20101 -1405
rect 20153 -1458 20160 -1405
rect 20095 -1459 20160 -1458
rect 18574 -1646 18630 -1637
rect 18574 -1711 18630 -1702
rect 18768 -1642 18824 -1633
rect 18768 -1707 18824 -1698
rect 18966 -1651 19022 -1642
rect 18966 -1716 19022 -1707
rect 19170 -1643 19226 -1634
rect 19170 -1708 19226 -1699
rect 19390 -1640 19446 -1631
rect 19390 -1705 19446 -1696
rect 19605 -1644 19661 -1635
rect 19605 -1709 19661 -1700
rect 19833 -1641 19889 -1632
rect 19833 -1706 19889 -1697
rect 20037 -1644 20093 -1635
rect 20037 -1709 20093 -1700
rect 20188 -1908 20230 -657
rect 20259 -1110 20315 -1101
rect 20259 -1175 20315 -1166
rect 20343 -1348 20385 -201
rect 20473 -517 20515 2219
rect 20666 1802 20672 1854
rect 20724 1802 20731 1854
rect 20577 271 20633 280
rect 20577 206 20633 215
rect 20551 -151 20605 -145
rect 20551 -203 20552 -151
rect 20604 -203 20605 -151
rect 20551 -209 20605 -203
rect 20467 -523 20519 -517
rect 20467 -581 20519 -575
rect 20557 -690 20599 -209
rect 20551 -696 20605 -690
rect 20551 -748 20552 -696
rect 20604 -748 20605 -696
rect 20551 -754 20605 -748
rect 20494 -1110 20550 -1101
rect 20494 -1175 20550 -1166
rect 20553 -1214 20605 -1208
rect 20677 -1218 20719 1802
rect 21552 691 21558 744
rect 21611 691 21617 744
rect 21552 690 21617 691
rect 21002 472 21009 524
rect 21061 472 21068 524
rect 20857 271 20913 280
rect 20857 206 20913 215
rect 21017 50 21054 472
rect 21174 270 21230 279
rect 21174 205 21230 214
rect 21003 -2 21010 50
rect 21062 -2 21069 50
rect 20884 -164 20891 -112
rect 20943 -164 20949 -112
rect 20783 -423 20839 -414
rect 20783 -488 20839 -479
rect 20897 -670 20939 -164
rect 21474 -273 21530 -264
rect 21474 -338 21530 -329
rect 21022 -421 21078 -412
rect 21022 -486 21078 -477
rect 21226 -421 21282 -412
rect 21226 -486 21282 -477
rect 20886 -723 20892 -670
rect 20944 -723 20951 -670
rect 20886 -724 20951 -723
rect 21564 -789 21606 690
rect 22094 37 22136 2429
rect 22262 475 22269 527
rect 22321 475 22328 527
rect 22277 53 22314 475
rect 22083 -16 22089 37
rect 22141 -16 22148 37
rect 22263 1 22270 53
rect 22322 1 22329 53
rect 22083 -17 22148 -16
rect 22499 -111 22541 2961
rect 23243 2685 23271 5767
rect 23395 5289 23428 6054
rect 23599 6040 23771 6050
rect 23599 5894 23609 6040
rect 23759 5894 23771 6040
rect 23933 6037 23963 7280
rect 24670 7275 24679 7331
rect 24735 7326 24744 7331
rect 24735 7322 25341 7326
rect 24735 7275 24775 7322
rect 24670 7271 24775 7275
rect 24671 7266 24775 7271
rect 24831 7266 24855 7322
rect 24911 7266 24935 7322
rect 24991 7266 25015 7322
rect 25071 7266 25095 7322
rect 25151 7266 25175 7322
rect 25231 7266 25341 7322
rect 24671 7260 25341 7266
rect 25403 7325 30311 7329
rect 25403 7269 25507 7325
rect 25563 7269 25587 7325
rect 25643 7269 25667 7325
rect 25723 7269 25747 7325
rect 25803 7269 25827 7325
rect 25883 7269 25907 7325
rect 25963 7269 26115 7325
rect 26171 7269 26195 7325
rect 26251 7269 26275 7325
rect 26331 7269 26355 7325
rect 26411 7269 26435 7325
rect 26491 7269 26515 7325
rect 26571 7269 26719 7325
rect 26775 7269 26799 7325
rect 26855 7269 26879 7325
rect 26935 7269 26959 7325
rect 27015 7269 27039 7325
rect 27095 7269 27119 7325
rect 27175 7269 27327 7325
rect 27383 7269 27407 7325
rect 27463 7269 27487 7325
rect 27543 7269 27567 7325
rect 27623 7269 27647 7325
rect 27703 7269 27727 7325
rect 27783 7269 27931 7325
rect 27987 7269 28011 7325
rect 28067 7269 28091 7325
rect 28147 7269 28171 7325
rect 28227 7269 28251 7325
rect 28307 7269 28331 7325
rect 28387 7269 28539 7325
rect 28595 7269 28619 7325
rect 28675 7269 28699 7325
rect 28755 7269 28779 7325
rect 28835 7269 28859 7325
rect 28915 7269 28939 7325
rect 28995 7269 29143 7325
rect 29199 7269 29223 7325
rect 29279 7269 29303 7325
rect 29359 7269 29383 7325
rect 29439 7269 29463 7325
rect 29519 7269 29543 7325
rect 29599 7269 29751 7325
rect 29807 7269 29831 7325
rect 29887 7269 29911 7325
rect 29967 7269 29991 7325
rect 30047 7269 30071 7325
rect 30127 7269 30151 7325
rect 30207 7269 30311 7325
rect 25403 7263 30311 7269
rect 30479 7269 30553 7273
rect 30479 7213 30488 7269
rect 30544 7213 30553 7269
rect 30479 7209 30553 7213
rect 30484 7125 30558 7129
rect 30484 7069 30493 7125
rect 30549 7069 30558 7125
rect 30484 7065 30558 7069
rect 30485 6973 30559 6977
rect 30485 6917 30494 6973
rect 30550 6917 30559 6973
rect 30485 6913 30559 6917
rect 30485 6803 30559 6807
rect 30485 6747 30494 6803
rect 30550 6747 30559 6803
rect 30485 6743 30559 6747
rect 24062 6726 24118 6735
rect 24062 6661 24118 6670
rect 24193 6725 24249 6734
rect 24193 6660 24249 6669
rect 24337 6726 24393 6735
rect 24337 6661 24393 6670
rect 30484 6646 30558 6650
rect 30484 6590 30493 6646
rect 30549 6590 30558 6646
rect 30484 6586 30558 6590
rect 24329 6361 24337 6413
rect 24389 6361 24395 6413
rect 30779 6412 30853 6416
rect 24329 6360 24395 6361
rect 30402 6404 30476 6408
rect 24347 6284 24393 6360
rect 30402 6348 30411 6404
rect 30467 6348 30476 6404
rect 30779 6356 30788 6412
rect 30844 6356 30853 6412
rect 30779 6352 30853 6356
rect 30979 6412 31053 6416
rect 30979 6356 30988 6412
rect 31044 6356 31053 6412
rect 30979 6352 31053 6356
rect 30402 6344 30476 6348
rect 24347 6238 24586 6284
rect 24080 6180 24136 6189
rect 24080 6115 24136 6124
rect 24200 6180 24256 6189
rect 24200 6115 24256 6124
rect 24343 6180 24399 6189
rect 24343 6115 24399 6124
rect 23914 5985 23921 6037
rect 23973 5985 23979 6037
rect 23914 5984 23979 5985
rect 23599 5884 23771 5894
rect 24343 5835 24408 5836
rect 23599 5814 23771 5824
rect 23599 5668 23609 5814
rect 23759 5668 23771 5814
rect 24343 5783 24349 5835
rect 24401 5832 24408 5835
rect 24540 5832 24586 6238
rect 25886 6145 25965 6146
rect 26113 6145 26192 6146
rect 27098 6145 27177 6146
rect 27325 6145 27404 6146
rect 28310 6145 28389 6146
rect 28537 6145 28616 6146
rect 29522 6145 29601 6146
rect 29749 6145 29828 6146
rect 25154 6142 25233 6143
rect 25151 6078 25161 6142
rect 25225 6078 25234 6142
rect 25883 6081 25893 6145
rect 25957 6081 25966 6145
rect 26112 6081 26121 6145
rect 26185 6081 26195 6145
rect 27095 6081 27105 6145
rect 27169 6081 27178 6145
rect 27324 6081 27333 6145
rect 27397 6081 27407 6145
rect 28307 6081 28317 6145
rect 28381 6081 28390 6145
rect 28536 6081 28545 6145
rect 28609 6081 28619 6145
rect 29519 6081 29529 6145
rect 29593 6081 29602 6145
rect 29748 6081 29757 6145
rect 29821 6081 29831 6145
rect 30490 6143 30564 6147
rect 30490 6087 30499 6143
rect 30555 6087 30564 6143
rect 30490 6083 30564 6087
rect 25508 5879 25517 5943
rect 25581 5879 25590 5943
rect 25508 5878 25590 5879
rect 26240 5879 26249 5943
rect 26313 5879 26322 5943
rect 26240 5878 26322 5879
rect 26458 5879 26467 5943
rect 26531 5879 26540 5943
rect 26458 5878 26540 5879
rect 27452 5879 27461 5943
rect 27525 5879 27534 5943
rect 27452 5878 27534 5879
rect 27670 5879 27679 5943
rect 27743 5879 27752 5943
rect 27670 5878 27752 5879
rect 28790 5879 28799 5943
rect 28863 5879 28872 5943
rect 28790 5878 28872 5879
rect 29008 5879 29017 5943
rect 29081 5879 29090 5943
rect 29008 5878 29090 5879
rect 29742 5879 29751 5943
rect 29815 5879 29824 5943
rect 30490 5940 30564 5944
rect 30490 5884 30499 5940
rect 30555 5884 30564 5940
rect 30490 5880 30564 5884
rect 29742 5878 29824 5879
rect 24830 5832 24837 5835
rect 24401 5786 24837 5832
rect 24401 5783 24408 5786
rect 24830 5783 24837 5786
rect 24889 5783 24895 5835
rect 24830 5782 24895 5783
rect 30590 5770 30664 5774
rect 30590 5714 30599 5770
rect 30655 5714 30664 5770
rect 30590 5710 30664 5714
rect 23599 5658 23771 5668
rect 30399 5678 30473 5682
rect 30399 5622 30408 5678
rect 30464 5622 30473 5678
rect 30399 5618 30473 5622
rect 23377 5237 23383 5289
rect 23435 5237 23441 5289
rect 23377 5236 23441 5237
rect 23615 5080 23787 5090
rect 23615 4934 23625 5080
rect 23775 4934 23787 5080
rect 23615 4924 23787 4934
rect 24656 4753 24730 4757
rect 24656 4697 24665 4753
rect 24721 4697 24730 4753
rect 24656 4693 24730 4697
rect 25191 4756 25523 4760
rect 25191 4700 25207 4756
rect 25263 4700 25287 4756
rect 25343 4700 25367 4756
rect 25423 4700 25447 4756
rect 25503 4700 25523 4756
rect 25191 4692 25523 4700
rect 25923 4756 26255 4760
rect 25923 4700 25939 4756
rect 25995 4700 26019 4756
rect 26075 4700 26099 4756
rect 26155 4700 26179 4756
rect 26235 4700 26255 4756
rect 25923 4692 26255 4700
rect 26525 4756 26857 4760
rect 26525 4700 26545 4756
rect 26601 4700 26625 4756
rect 26681 4700 26705 4756
rect 26761 4700 26785 4756
rect 26841 4700 26857 4756
rect 26525 4692 26857 4700
rect 27135 4756 27467 4760
rect 27135 4700 27151 4756
rect 27207 4700 27231 4756
rect 27287 4700 27311 4756
rect 27367 4700 27391 4756
rect 27447 4700 27467 4756
rect 27135 4692 27467 4700
rect 27737 4756 28069 4760
rect 27737 4700 27757 4756
rect 27813 4700 27837 4756
rect 27893 4700 27917 4756
rect 27973 4700 27997 4756
rect 28053 4700 28069 4756
rect 27737 4692 28069 4700
rect 28473 4756 28805 4760
rect 28473 4700 28489 4756
rect 28545 4700 28569 4756
rect 28625 4700 28649 4756
rect 28705 4700 28729 4756
rect 28785 4700 28805 4756
rect 28473 4692 28805 4700
rect 29075 4756 29407 4760
rect 29075 4700 29095 4756
rect 29151 4700 29175 4756
rect 29231 4700 29255 4756
rect 29311 4700 29335 4756
rect 29391 4700 29407 4756
rect 29075 4692 29407 4700
rect 29809 4756 30141 4760
rect 29809 4700 29829 4756
rect 29885 4700 29909 4756
rect 29965 4700 29989 4756
rect 30045 4700 30069 4756
rect 30125 4700 30141 4756
rect 29809 4692 30141 4700
rect 25616 4372 25622 4424
rect 25674 4372 25680 4424
rect 28010 4372 28016 4424
rect 28068 4372 28074 4424
rect 23386 4265 23439 4272
rect 23438 4213 23439 4265
rect 23386 4206 23439 4213
rect 23398 3503 23426 4206
rect 23595 4088 23767 4098
rect 23595 3942 23605 4088
rect 23755 3942 23767 4088
rect 25635 4087 25663 4372
rect 25703 4252 25712 4308
rect 25768 4252 25778 4308
rect 25703 4251 25778 4252
rect 25877 4251 25886 4307
rect 25942 4251 25952 4307
rect 26102 4253 26111 4309
rect 26167 4253 26177 4309
rect 26303 4255 26312 4311
rect 26368 4255 26378 4311
rect 26303 4254 26378 4255
rect 26102 4252 26177 4253
rect 26526 4253 26535 4309
rect 26591 4253 26601 4309
rect 26735 4258 26744 4314
rect 26800 4258 26810 4314
rect 26735 4257 26810 4258
rect 26526 4252 26601 4253
rect 25877 4250 25952 4251
rect 26963 4251 26972 4307
rect 27028 4251 27038 4307
rect 27153 4255 27162 4311
rect 27218 4255 27228 4311
rect 27358 4258 27367 4314
rect 27423 4258 27433 4314
rect 27358 4257 27433 4258
rect 27557 4258 27566 4314
rect 27622 4258 27632 4314
rect 27557 4257 27632 4258
rect 27153 4254 27228 4255
rect 27773 4253 27782 4309
rect 27838 4253 27848 4309
rect 27773 4252 27848 4253
rect 26963 4250 27038 4251
rect 25613 4081 25665 4087
rect 27061 4065 27070 4121
rect 27126 4065 27136 4121
rect 27061 4064 27136 4065
rect 25613 4023 25665 4029
rect 23595 3932 23767 3942
rect 23382 3497 23434 3503
rect 23382 3439 23434 3445
rect 23398 3013 23426 3439
rect 25635 3438 25663 4023
rect 27446 4014 27455 4070
rect 27511 4014 27521 4070
rect 28029 4045 28057 4372
rect 28161 4258 28170 4314
rect 28226 4258 28236 4314
rect 28161 4257 28236 4258
rect 28396 4253 28405 4309
rect 28461 4253 28471 4309
rect 28638 4255 28647 4311
rect 28703 4255 28713 4311
rect 28870 4256 28879 4312
rect 28935 4256 28945 4312
rect 29099 4259 29108 4315
rect 29164 4259 29174 4315
rect 29099 4258 29174 4259
rect 28870 4255 28945 4256
rect 28638 4254 28713 4255
rect 28396 4252 28471 4253
rect 29348 4251 29357 4307
rect 29413 4251 29423 4307
rect 29566 4255 29575 4311
rect 29631 4255 29641 4311
rect 29566 4254 29641 4255
rect 29348 4250 29423 4251
rect 29795 4251 29804 4307
rect 29860 4251 29870 4307
rect 30016 4253 30025 4309
rect 30081 4253 30091 4309
rect 30232 4258 30241 4314
rect 30297 4258 30307 4314
rect 30232 4257 30307 4258
rect 30016 4252 30091 4253
rect 29795 4250 29870 4251
rect 29456 4064 29465 4120
rect 29521 4064 29531 4120
rect 29456 4063 29531 4064
rect 27446 4013 27521 4014
rect 28005 4039 28057 4045
rect 29841 4015 29850 4071
rect 29906 4015 29916 4071
rect 29841 4014 29916 4015
rect 28005 3981 28057 3987
rect 25705 3669 25714 3725
rect 25770 3669 25780 3725
rect 25705 3668 25780 3669
rect 25880 3667 25889 3723
rect 25945 3667 25955 3723
rect 26077 3669 26086 3725
rect 26142 3669 26152 3725
rect 26296 3672 26305 3728
rect 26361 3672 26371 3728
rect 26296 3671 26371 3672
rect 26077 3668 26152 3669
rect 26528 3668 26537 3724
rect 26593 3668 26603 3724
rect 26528 3667 26603 3668
rect 26712 3675 26761 3731
rect 26817 3675 26827 3731
rect 25880 3666 25955 3667
rect 25608 3432 25663 3438
rect 23601 3410 23773 3420
rect 23601 3264 23611 3410
rect 23761 3264 23773 3410
rect 25660 3380 25663 3432
rect 25608 3374 25663 3380
rect 23601 3254 23773 3264
rect 24881 3103 24887 3155
rect 24940 3103 24946 3155
rect 23380 2961 23386 3013
rect 23438 2961 23444 3013
rect 23398 2760 23426 2961
rect 23395 2726 23429 2760
rect 23239 2549 23273 2685
rect 23398 2654 23426 2726
rect 24475 2564 24482 2616
rect 24534 2564 24540 2616
rect 23224 2497 23230 2549
rect 23282 2497 23288 2549
rect 22853 2290 22859 2342
rect 22911 2290 22918 2342
rect 22485 -163 22492 -111
rect 22544 -163 22550 -111
rect 21678 -268 21734 -259
rect 21678 -333 21734 -324
rect 21869 -273 21925 -264
rect 21869 -338 21925 -329
rect 22071 -274 22127 -265
rect 22071 -339 22127 -330
rect 22361 -273 22417 -264
rect 22361 -338 22417 -329
rect 21559 -795 21613 -789
rect 21559 -847 21560 -795
rect 21612 -847 21613 -795
rect 21559 -853 21613 -847
rect 21473 -958 21529 -949
rect 21473 -1023 21529 -1014
rect 20783 -1108 20839 -1099
rect 20783 -1173 20839 -1164
rect 20973 -1110 21029 -1101
rect 20973 -1175 21029 -1166
rect 21177 -1108 21233 -1099
rect 21177 -1173 21233 -1164
rect 20605 -1260 20719 -1218
rect 21565 -1250 21607 -853
rect 21674 -957 21730 -948
rect 21674 -1022 21730 -1013
rect 21892 -961 21948 -952
rect 21892 -1026 21948 -1017
rect 22099 -957 22155 -948
rect 22099 -1022 22155 -1013
rect 22304 -958 22360 -949
rect 22304 -1023 22360 -1014
rect 20553 -1272 20605 -1266
rect 20831 -1278 20883 -1272
rect 21554 -1302 21560 -1250
rect 21612 -1302 21618 -1250
rect 20831 -1336 20883 -1330
rect 20343 -1388 20447 -1348
rect 20441 -1400 20447 -1388
rect 20501 -1400 20507 -1348
rect 20275 -1642 20331 -1633
rect 20275 -1707 20331 -1698
rect 20468 -1641 20524 -1632
rect 20468 -1706 20524 -1697
rect 20665 -1646 20721 -1637
rect 20665 -1711 20721 -1702
rect 20835 -1908 20877 -1336
rect 22499 -1405 22541 -163
rect 22723 -203 22729 -151
rect 22781 -203 22789 -151
rect 22646 -274 22702 -265
rect 22646 -339 22702 -330
rect 22577 -600 22629 -594
rect 22577 -658 22629 -652
rect 22488 -1458 22494 -1405
rect 22546 -1458 22553 -1405
rect 22488 -1459 22553 -1458
rect 20921 -1643 20977 -1634
rect 20921 -1708 20977 -1699
rect 21160 -1647 21216 -1638
rect 21160 -1712 21216 -1703
rect 21393 -1651 21449 -1642
rect 21393 -1716 21449 -1707
rect 21614 -1646 21670 -1637
rect 21614 -1711 21670 -1702
rect 21805 -1646 21861 -1637
rect 21805 -1711 21861 -1702
rect 22033 -1644 22089 -1635
rect 22033 -1709 22089 -1700
rect 22230 -1649 22286 -1640
rect 22230 -1714 22286 -1705
rect 22442 -1649 22498 -1640
rect 22442 -1714 22498 -1705
rect 22581 -1908 22623 -658
rect 22651 -962 22707 -953
rect 22651 -1027 22707 -1018
rect 22735 -1350 22777 -203
rect 22865 -517 22907 2290
rect 23055 1872 23061 1924
rect 23113 1872 23120 1924
rect 22964 268 23020 277
rect 22964 203 23020 212
rect 22944 -150 22998 -144
rect 22944 -202 22945 -150
rect 22997 -202 22998 -150
rect 22944 -208 22998 -202
rect 22859 -523 22911 -517
rect 22859 -581 22911 -575
rect 22950 -689 22992 -208
rect 22944 -695 22998 -689
rect 22944 -747 22945 -695
rect 22997 -747 22998 -695
rect 22944 -753 22998 -747
rect 22963 -1102 23019 -1093
rect 22963 -1167 23019 -1158
rect 22944 -1214 22996 -1208
rect 23068 -1218 23110 1872
rect 23945 691 23951 744
rect 24004 691 24010 744
rect 23945 690 24010 691
rect 23394 473 23401 525
rect 23453 473 23460 525
rect 23259 268 23315 277
rect 23259 203 23315 212
rect 23409 51 23446 473
rect 23546 268 23602 277
rect 23546 203 23602 212
rect 23836 268 23892 277
rect 23836 203 23892 212
rect 23395 -1 23402 51
rect 23454 -1 23461 51
rect 23279 -164 23286 -112
rect 23338 -164 23344 -112
rect 23186 -413 23242 -404
rect 23186 -478 23242 -469
rect 23290 -671 23332 -164
rect 23419 -415 23475 -406
rect 23419 -480 23475 -471
rect 23626 -417 23682 -408
rect 23626 -482 23682 -473
rect 23835 -415 23891 -406
rect 23835 -480 23891 -471
rect 23279 -724 23285 -671
rect 23337 -724 23344 -671
rect 23279 -725 23344 -724
rect 23957 -789 23999 690
rect 24120 271 24176 280
rect 24120 206 24176 215
rect 24489 38 24531 2564
rect 24657 475 24664 527
rect 24716 475 24723 527
rect 24672 53 24709 475
rect 24478 -15 24484 38
rect 24536 -15 24543 38
rect 24658 1 24665 53
rect 24717 1 24724 53
rect 24478 -16 24543 -15
rect 24892 -111 24934 3103
rect 25635 2823 25663 3374
rect 26712 3622 26827 3675
rect 26964 3663 26973 3719
rect 27029 3663 27039 3719
rect 26964 3662 27039 3663
rect 27186 3659 27195 3715
rect 27251 3659 27261 3715
rect 27186 3658 27261 3659
rect 27408 3712 27496 3717
rect 27408 3656 27418 3712
rect 27474 3656 27496 3712
rect 27408 3636 27496 3656
rect 27619 3656 27628 3712
rect 27684 3656 27694 3712
rect 27619 3655 27694 3656
rect 27832 3656 27841 3712
rect 27897 3656 27907 3712
rect 27832 3655 27907 3656
rect 26712 3293 26756 3622
rect 27460 3357 27496 3636
rect 28029 3396 28057 3981
rect 28149 3649 28158 3705
rect 28214 3649 28224 3705
rect 28351 3652 28360 3708
rect 28416 3652 28426 3708
rect 28552 3653 28561 3709
rect 28617 3653 28627 3709
rect 28731 3654 28740 3710
rect 28796 3654 28806 3710
rect 28923 3658 28932 3714
rect 28988 3658 28998 3714
rect 28923 3657 28998 3658
rect 29096 3711 29184 3715
rect 28731 3653 28806 3654
rect 29096 3655 29117 3711
rect 29173 3655 29184 3711
rect 28552 3652 28627 3653
rect 28351 3651 28426 3652
rect 28149 3648 28224 3649
rect 28004 3390 28057 3396
rect 27449 3305 27455 3357
rect 27507 3305 27513 3357
rect 28056 3338 28057 3390
rect 28004 3332 28057 3338
rect 26691 3241 26697 3293
rect 26749 3276 26756 3293
rect 26749 3241 26755 3276
rect 26691 3240 26755 3241
rect 25732 3020 25741 3076
rect 25797 3020 25807 3076
rect 25948 3025 25957 3081
rect 26013 3025 26023 3081
rect 26154 3026 26163 3082
rect 26219 3026 26229 3082
rect 26154 3025 26229 3026
rect 25948 3024 26023 3025
rect 25732 3019 25807 3020
rect 26356 3018 26365 3074
rect 26421 3018 26431 3074
rect 26552 3020 26561 3076
rect 26617 3020 26627 3076
rect 26777 3022 26786 3078
rect 26842 3022 26852 3078
rect 26777 3021 26852 3022
rect 26552 3019 26627 3020
rect 26356 3017 26431 3018
rect 26992 3018 27001 3074
rect 27057 3018 27067 3074
rect 26992 3017 27067 3018
rect 27227 3018 27236 3074
rect 27292 3018 27302 3074
rect 27435 3021 27444 3077
rect 27500 3021 27510 3077
rect 27435 3020 27510 3021
rect 27677 3021 27686 3077
rect 27742 3021 27752 3077
rect 27875 3022 27884 3078
rect 27940 3022 27950 3078
rect 27875 3021 27950 3022
rect 27677 3020 27752 3021
rect 27227 3017 27302 3018
rect 25616 2817 25668 2823
rect 27066 2791 27075 2847
rect 27131 2791 27141 2847
rect 27066 2790 27141 2791
rect 25616 2759 25668 2765
rect 25247 2361 25253 2413
rect 25305 2361 25312 2413
rect 24880 -163 24887 -111
rect 24939 -163 24945 -111
rect 24401 -269 24457 -260
rect 24401 -334 24457 -325
rect 24595 -265 24651 -256
rect 24595 -330 24651 -321
rect 24784 -268 24840 -259
rect 24784 -333 24840 -324
rect 24115 -413 24171 -404
rect 24115 -478 24171 -469
rect 23951 -795 24005 -789
rect 23951 -847 23952 -795
rect 24004 -847 24005 -795
rect 23951 -853 24005 -847
rect 23205 -1106 23261 -1097
rect 23205 -1171 23261 -1162
rect 23405 -1107 23461 -1098
rect 23405 -1172 23461 -1163
rect 23595 -1099 23651 -1090
rect 23595 -1164 23651 -1155
rect 23816 -1101 23872 -1092
rect 23816 -1166 23872 -1157
rect 22996 -1260 23110 -1218
rect 23957 -1250 23999 -853
rect 24403 -958 24459 -949
rect 24403 -1023 24459 -1014
rect 24594 -955 24650 -946
rect 24594 -1020 24650 -1011
rect 24789 -953 24845 -944
rect 24789 -1018 24845 -1009
rect 24112 -1106 24168 -1097
rect 24112 -1171 24168 -1162
rect 22944 -1272 22996 -1266
rect 23224 -1279 23276 -1273
rect 23946 -1302 23952 -1250
rect 24004 -1302 24010 -1250
rect 23224 -1337 23276 -1331
rect 22735 -1390 22839 -1350
rect 22833 -1402 22839 -1390
rect 22893 -1402 22899 -1350
rect 22669 -1646 22725 -1637
rect 22669 -1711 22725 -1702
rect 22858 -1645 22914 -1636
rect 22858 -1710 22914 -1701
rect 23084 -1644 23140 -1635
rect 23084 -1709 23140 -1700
rect 23228 -1908 23270 -1337
rect 24892 -1405 24934 -163
rect 25115 -201 25121 -149
rect 25173 -201 25181 -149
rect 25007 -266 25063 -257
rect 25007 -331 25063 -322
rect 24970 -598 25022 -592
rect 24970 -656 25022 -650
rect 24881 -1458 24887 -1405
rect 24939 -1458 24946 -1405
rect 24881 -1459 24946 -1458
rect 23338 -1644 23394 -1635
rect 23338 -1709 23394 -1700
rect 23582 -1647 23638 -1638
rect 23582 -1712 23638 -1703
rect 23812 -1648 23868 -1639
rect 23812 -1713 23868 -1704
rect 24070 -1645 24126 -1636
rect 24070 -1710 24126 -1701
rect 24280 -1645 24336 -1636
rect 24280 -1710 24336 -1701
rect 24505 -1645 24561 -1636
rect 24505 -1710 24561 -1701
rect 24724 -1648 24780 -1639
rect 24724 -1713 24780 -1704
rect 24974 -1908 25016 -656
rect 25127 -1348 25169 -201
rect 25257 -517 25299 2361
rect 25635 2063 25663 2759
rect 27449 2732 27458 2788
rect 27514 2732 27524 2788
rect 28029 2780 28057 3332
rect 29096 3640 29184 3655
rect 29340 3654 29349 3710
rect 29405 3654 29415 3710
rect 29545 3656 29554 3712
rect 29610 3656 29620 3712
rect 29751 3658 29760 3714
rect 29816 3658 29826 3714
rect 29751 3657 29826 3658
rect 29856 3657 29862 3709
rect 29914 3657 29920 3709
rect 29959 3665 29968 3721
rect 30024 3665 30034 3721
rect 30181 3666 30190 3722
rect 30246 3666 30256 3722
rect 30181 3665 30256 3666
rect 29959 3664 30034 3665
rect 29545 3655 29620 3656
rect 29340 3653 29415 3654
rect 29096 3293 29140 3640
rect 29856 3358 29906 3657
rect 29842 3306 29848 3358
rect 29900 3306 29906 3358
rect 29086 3241 29092 3293
rect 29144 3241 29150 3293
rect 28182 3022 28191 3078
rect 28247 3022 28257 3078
rect 28407 3023 28416 3079
rect 28472 3023 28482 3079
rect 28407 3022 28482 3023
rect 28636 3022 28645 3078
rect 28701 3022 28711 3078
rect 28852 3026 28861 3082
rect 28917 3026 28927 3082
rect 29075 3029 29084 3085
rect 29140 3029 29150 3085
rect 29075 3028 29150 3029
rect 28852 3025 28927 3026
rect 29299 3025 29308 3081
rect 29364 3025 29374 3081
rect 29299 3024 29374 3025
rect 28182 3021 28257 3022
rect 28636 3021 28711 3022
rect 29526 3014 29535 3070
rect 29591 3014 29601 3070
rect 29526 3013 29601 3014
rect 29739 3013 29748 3069
rect 29804 3013 29814 3069
rect 29950 3017 29959 3073
rect 30015 3017 30025 3073
rect 30177 3018 30186 3074
rect 30242 3018 30252 3074
rect 30177 3017 30252 3018
rect 29950 3016 30025 3017
rect 29739 3012 29814 3013
rect 29458 2793 29467 2849
rect 29523 2793 29533 2849
rect 29458 2792 29533 2793
rect 27449 2731 27524 2732
rect 28003 2774 28057 2780
rect 28055 2722 28057 2774
rect 29835 2739 29844 2795
rect 29900 2739 29910 2795
rect 29835 2738 29910 2739
rect 28003 2716 28057 2722
rect 25758 2375 25767 2431
rect 25823 2375 25833 2431
rect 25983 2384 25992 2440
rect 26048 2384 26058 2440
rect 25983 2383 26058 2384
rect 26260 2381 26269 2437
rect 26325 2381 26335 2437
rect 26481 2384 26490 2440
rect 26546 2384 26556 2440
rect 26481 2383 26556 2384
rect 26697 2437 26765 2439
rect 26260 2380 26335 2381
rect 26697 2381 26735 2437
rect 26791 2381 26801 2437
rect 26952 2385 26961 2441
rect 27017 2385 27027 2441
rect 26952 2384 27027 2385
rect 27164 2383 27173 2439
rect 27229 2383 27239 2439
rect 27384 2389 27393 2445
rect 27449 2442 27459 2445
rect 27449 2389 27498 2442
rect 27622 2391 27631 2447
rect 27687 2391 27697 2447
rect 27835 2393 27844 2449
rect 27900 2393 27910 2449
rect 27835 2392 27910 2393
rect 27622 2390 27697 2391
rect 27384 2388 27498 2389
rect 27164 2382 27239 2383
rect 26697 2380 26801 2381
rect 25758 2374 25833 2375
rect 25611 2057 25663 2063
rect 26714 2013 26750 2380
rect 27453 2079 27498 2388
rect 28029 2093 28057 2716
rect 28222 2383 28231 2439
rect 28287 2383 28297 2439
rect 28569 2384 28578 2440
rect 28634 2384 28644 2440
rect 28986 2437 29303 2443
rect 28986 2435 29237 2437
rect 28569 2383 28644 2384
rect 28222 2382 28297 2383
rect 28805 2379 28814 2435
rect 28870 2379 28880 2435
rect 28805 2378 28880 2379
rect 28986 2379 28998 2435
rect 29054 2381 29237 2435
rect 29293 2381 29303 2437
rect 29054 2379 29303 2381
rect 28986 2368 29303 2379
rect 29431 2377 29440 2433
rect 29496 2377 29506 2433
rect 29431 2376 29506 2377
rect 29616 2374 29625 2430
rect 29681 2374 29691 2430
rect 29807 2376 29816 2432
rect 29872 2429 29882 2432
rect 29872 2376 29895 2429
rect 29998 2380 30007 2436
rect 30063 2380 30073 2436
rect 29998 2379 30073 2380
rect 29807 2375 29895 2376
rect 30184 2376 30193 2432
rect 30249 2376 30259 2432
rect 30184 2375 30259 2376
rect 29616 2373 29691 2374
rect 28004 2087 28057 2093
rect 27449 2078 27514 2079
rect 27449 2026 27455 2078
rect 27507 2026 27514 2078
rect 28056 2035 28057 2087
rect 28004 2029 28057 2035
rect 25611 1999 25663 2005
rect 25635 1998 25663 1999
rect 26697 1974 26706 2013
rect 26698 1961 26706 1974
rect 26758 1974 26765 2013
rect 28029 2011 28057 2029
rect 29107 2013 29143 2368
rect 29858 2080 29895 2375
rect 29841 2079 29905 2080
rect 29841 2027 29847 2079
rect 29899 2027 29905 2079
rect 26758 1961 26764 1974
rect 29089 1961 29096 2013
rect 29149 1961 29156 2013
rect 25631 1793 25640 1849
rect 25696 1793 25706 1849
rect 25631 1792 25706 1793
rect 25836 1789 25845 1845
rect 25901 1789 25911 1845
rect 26022 1794 26031 1850
rect 26087 1794 26097 1850
rect 26022 1793 26097 1794
rect 25836 1788 25911 1789
rect 26216 1787 26225 1843
rect 26281 1787 26291 1843
rect 26435 1792 26444 1848
rect 26500 1792 26510 1848
rect 26435 1791 26510 1792
rect 26645 1792 26654 1848
rect 26710 1792 26720 1848
rect 26645 1791 26720 1792
rect 26874 1789 26883 1845
rect 26939 1789 26949 1845
rect 26874 1788 26949 1789
rect 27120 1789 27129 1845
rect 27185 1789 27195 1845
rect 27120 1788 27195 1789
rect 27394 1789 27403 1845
rect 27459 1789 27469 1845
rect 27394 1788 27469 1789
rect 27669 1789 27678 1845
rect 27734 1789 27744 1845
rect 27669 1788 27744 1789
rect 27905 1789 27914 1845
rect 27970 1789 27980 1845
rect 28128 1792 28137 1848
rect 28193 1792 28203 1848
rect 28346 1795 28355 1851
rect 28411 1795 28421 1851
rect 28346 1794 28421 1795
rect 28128 1791 28203 1792
rect 27905 1788 27980 1789
rect 26216 1786 26291 1787
rect 28524 1786 28533 1842
rect 28589 1786 28599 1842
rect 28763 1788 28772 1844
rect 28828 1788 28838 1844
rect 28763 1787 28838 1788
rect 28960 1788 28969 1844
rect 29025 1788 29035 1844
rect 28960 1787 29035 1788
rect 29158 1788 29167 1844
rect 29223 1788 29233 1844
rect 29371 1789 29380 1845
rect 29436 1789 29446 1845
rect 29371 1788 29446 1789
rect 29594 1788 29603 1844
rect 29659 1788 29669 1844
rect 29791 1793 29800 1849
rect 29856 1793 29866 1849
rect 29791 1792 29866 1793
rect 30007 1791 30016 1847
rect 30072 1791 30082 1847
rect 30007 1790 30082 1791
rect 30216 1791 30225 1847
rect 30281 1791 30291 1847
rect 30216 1790 30291 1791
rect 29158 1787 29233 1788
rect 29594 1787 29669 1788
rect 28524 1785 28599 1786
rect 25251 -523 25303 -517
rect 25251 -581 25303 -575
rect 25236 -958 25292 -949
rect 25236 -1023 25292 -1014
rect 25127 -1388 25231 -1348
rect 25225 -1400 25231 -1388
rect 25285 -1400 25291 -1348
rect 25070 -1644 25126 -1635
rect 25070 -1709 25126 -1700
rect 25269 -1647 25325 -1638
rect 25269 -1712 25325 -1703
<< via2 >>
rect 13954 13626 14010 13628
rect 13954 13574 13956 13626
rect 13956 13574 14008 13626
rect 14008 13574 14010 13626
rect 13954 13572 14010 13574
rect 14050 13617 14106 13619
rect 14050 13565 14054 13617
rect 14054 13565 14106 13617
rect 14050 13563 14106 13565
rect 14130 13617 14186 13619
rect 14130 13565 14134 13617
rect 14134 13565 14186 13617
rect 14130 13563 14186 13565
rect 14210 13617 14266 13619
rect 14210 13565 14214 13617
rect 14214 13565 14266 13617
rect 14210 13563 14266 13565
rect 14290 13617 14346 13619
rect 14290 13565 14294 13617
rect 14294 13565 14346 13617
rect 14290 13563 14346 13565
rect 14370 13617 14426 13619
rect 14370 13565 14374 13617
rect 14374 13565 14426 13617
rect 14370 13563 14426 13565
rect 14450 13617 14506 13619
rect 14450 13565 14454 13617
rect 14454 13565 14506 13617
rect 14450 13563 14506 13565
rect 14782 13620 14838 13622
rect 14782 13568 14786 13620
rect 14786 13568 14838 13620
rect 14782 13566 14838 13568
rect 14862 13620 14918 13622
rect 14862 13568 14866 13620
rect 14866 13568 14918 13620
rect 14862 13566 14918 13568
rect 14942 13620 14998 13622
rect 14942 13568 14946 13620
rect 14946 13568 14998 13620
rect 14942 13566 14998 13568
rect 15022 13620 15078 13622
rect 15022 13568 15026 13620
rect 15026 13568 15078 13620
rect 15022 13566 15078 13568
rect 15102 13620 15158 13622
rect 15102 13568 15106 13620
rect 15106 13568 15158 13620
rect 15102 13566 15158 13568
rect 15182 13620 15238 13622
rect 15182 13568 15186 13620
rect 15186 13568 15238 13620
rect 15182 13566 15238 13568
rect 15390 13620 15446 13622
rect 15390 13568 15442 13620
rect 15442 13568 15446 13620
rect 15390 13566 15446 13568
rect 15470 13620 15526 13622
rect 15470 13568 15522 13620
rect 15522 13568 15526 13620
rect 15470 13566 15526 13568
rect 15550 13620 15606 13622
rect 15550 13568 15602 13620
rect 15602 13568 15606 13620
rect 15550 13566 15606 13568
rect 15630 13620 15686 13622
rect 15630 13568 15682 13620
rect 15682 13568 15686 13620
rect 15630 13566 15686 13568
rect 15710 13620 15766 13622
rect 15710 13568 15762 13620
rect 15762 13568 15766 13620
rect 15710 13566 15766 13568
rect 15790 13620 15846 13622
rect 15790 13568 15842 13620
rect 15842 13568 15846 13620
rect 15790 13566 15846 13568
rect 15994 13620 16050 13622
rect 15994 13568 15998 13620
rect 15998 13568 16050 13620
rect 15994 13566 16050 13568
rect 16074 13620 16130 13622
rect 16074 13568 16078 13620
rect 16078 13568 16130 13620
rect 16074 13566 16130 13568
rect 16154 13620 16210 13622
rect 16154 13568 16158 13620
rect 16158 13568 16210 13620
rect 16154 13566 16210 13568
rect 16234 13620 16290 13622
rect 16234 13568 16238 13620
rect 16238 13568 16290 13620
rect 16234 13566 16290 13568
rect 16314 13620 16370 13622
rect 16314 13568 16318 13620
rect 16318 13568 16370 13620
rect 16314 13566 16370 13568
rect 16394 13620 16450 13622
rect 16394 13568 16398 13620
rect 16398 13568 16450 13620
rect 16394 13566 16450 13568
rect 16602 13620 16658 13622
rect 16602 13568 16654 13620
rect 16654 13568 16658 13620
rect 16602 13566 16658 13568
rect 16682 13620 16738 13622
rect 16682 13568 16734 13620
rect 16734 13568 16738 13620
rect 16682 13566 16738 13568
rect 16762 13620 16818 13622
rect 16762 13568 16814 13620
rect 16814 13568 16818 13620
rect 16762 13566 16818 13568
rect 16842 13620 16898 13622
rect 16842 13568 16894 13620
rect 16894 13568 16898 13620
rect 16842 13566 16898 13568
rect 16922 13620 16978 13622
rect 16922 13568 16974 13620
rect 16974 13568 16978 13620
rect 16922 13566 16978 13568
rect 17002 13620 17058 13622
rect 17002 13568 17054 13620
rect 17054 13568 17058 13620
rect 17002 13566 17058 13568
rect 17206 13620 17262 13622
rect 17206 13568 17210 13620
rect 17210 13568 17262 13620
rect 17206 13566 17262 13568
rect 17286 13620 17342 13622
rect 17286 13568 17290 13620
rect 17290 13568 17342 13620
rect 17286 13566 17342 13568
rect 17366 13620 17422 13622
rect 17366 13568 17370 13620
rect 17370 13568 17422 13620
rect 17366 13566 17422 13568
rect 17446 13620 17502 13622
rect 17446 13568 17450 13620
rect 17450 13568 17502 13620
rect 17446 13566 17502 13568
rect 17526 13620 17582 13622
rect 17526 13568 17530 13620
rect 17530 13568 17582 13620
rect 17526 13566 17582 13568
rect 17606 13620 17662 13622
rect 17606 13568 17610 13620
rect 17610 13568 17662 13620
rect 17606 13566 17662 13568
rect 17814 13620 17870 13622
rect 17814 13568 17866 13620
rect 17866 13568 17870 13620
rect 17814 13566 17870 13568
rect 17894 13620 17950 13622
rect 17894 13568 17946 13620
rect 17946 13568 17950 13620
rect 17894 13566 17950 13568
rect 17974 13620 18030 13622
rect 17974 13568 18026 13620
rect 18026 13568 18030 13620
rect 17974 13566 18030 13568
rect 18054 13620 18110 13622
rect 18054 13568 18106 13620
rect 18106 13568 18110 13620
rect 18054 13566 18110 13568
rect 18134 13620 18190 13622
rect 18134 13568 18186 13620
rect 18186 13568 18190 13620
rect 18134 13566 18190 13568
rect 18214 13620 18270 13622
rect 18214 13568 18266 13620
rect 18266 13568 18270 13620
rect 18214 13566 18270 13568
rect 18418 13620 18474 13622
rect 18418 13568 18422 13620
rect 18422 13568 18474 13620
rect 18418 13566 18474 13568
rect 18498 13620 18554 13622
rect 18498 13568 18502 13620
rect 18502 13568 18554 13620
rect 18498 13566 18554 13568
rect 18578 13620 18634 13622
rect 18578 13568 18582 13620
rect 18582 13568 18634 13620
rect 18578 13566 18634 13568
rect 18658 13620 18714 13622
rect 18658 13568 18662 13620
rect 18662 13568 18714 13620
rect 18658 13566 18714 13568
rect 18738 13620 18794 13622
rect 18738 13568 18742 13620
rect 18742 13568 18794 13620
rect 18738 13566 18794 13568
rect 18818 13620 18874 13622
rect 18818 13568 18822 13620
rect 18822 13568 18874 13620
rect 18818 13566 18874 13568
rect 19026 13620 19082 13622
rect 19026 13568 19078 13620
rect 19078 13568 19082 13620
rect 19026 13566 19082 13568
rect 19106 13620 19162 13622
rect 19106 13568 19158 13620
rect 19158 13568 19162 13620
rect 19106 13566 19162 13568
rect 19186 13620 19242 13622
rect 19186 13568 19238 13620
rect 19238 13568 19242 13620
rect 19186 13566 19242 13568
rect 19266 13620 19322 13622
rect 19266 13568 19318 13620
rect 19318 13568 19322 13620
rect 19266 13566 19322 13568
rect 19346 13620 19402 13622
rect 19346 13568 19398 13620
rect 19398 13568 19402 13620
rect 19346 13566 19402 13568
rect 19426 13620 19482 13622
rect 19426 13568 19478 13620
rect 19478 13568 19482 13620
rect 19426 13566 19482 13568
rect 19763 13564 19819 13566
rect 19763 13512 19765 13564
rect 19765 13512 19817 13564
rect 19817 13512 19819 13564
rect 19763 13510 19819 13512
rect 20240 13567 20296 13569
rect 20240 13515 20242 13567
rect 20242 13515 20294 13567
rect 20294 13515 20296 13567
rect 20240 13513 20296 13515
rect 20663 13626 20719 13628
rect 20663 13574 20665 13626
rect 20665 13574 20717 13626
rect 20717 13574 20719 13626
rect 20663 13572 20719 13574
rect 20759 13617 20815 13619
rect 20759 13565 20763 13617
rect 20763 13565 20815 13617
rect 20759 13563 20815 13565
rect 20839 13617 20895 13619
rect 20839 13565 20843 13617
rect 20843 13565 20895 13617
rect 20839 13563 20895 13565
rect 20919 13617 20975 13619
rect 20919 13565 20923 13617
rect 20923 13565 20975 13617
rect 20919 13563 20975 13565
rect 20999 13617 21055 13619
rect 20999 13565 21003 13617
rect 21003 13565 21055 13617
rect 20999 13563 21055 13565
rect 21079 13617 21135 13619
rect 21079 13565 21083 13617
rect 21083 13565 21135 13617
rect 21079 13563 21135 13565
rect 21159 13617 21215 13619
rect 21159 13565 21163 13617
rect 21163 13565 21215 13617
rect 21159 13563 21215 13565
rect 21491 13620 21547 13622
rect 21491 13568 21495 13620
rect 21495 13568 21547 13620
rect 21491 13566 21547 13568
rect 21571 13620 21627 13622
rect 21571 13568 21575 13620
rect 21575 13568 21627 13620
rect 21571 13566 21627 13568
rect 21651 13620 21707 13622
rect 21651 13568 21655 13620
rect 21655 13568 21707 13620
rect 21651 13566 21707 13568
rect 21731 13620 21787 13622
rect 21731 13568 21735 13620
rect 21735 13568 21787 13620
rect 21731 13566 21787 13568
rect 21811 13620 21867 13622
rect 21811 13568 21815 13620
rect 21815 13568 21867 13620
rect 21811 13566 21867 13568
rect 21891 13620 21947 13622
rect 21891 13568 21895 13620
rect 21895 13568 21947 13620
rect 21891 13566 21947 13568
rect 22099 13620 22155 13622
rect 22099 13568 22151 13620
rect 22151 13568 22155 13620
rect 22099 13566 22155 13568
rect 22179 13620 22235 13622
rect 22179 13568 22231 13620
rect 22231 13568 22235 13620
rect 22179 13566 22235 13568
rect 22259 13620 22315 13622
rect 22259 13568 22311 13620
rect 22311 13568 22315 13620
rect 22259 13566 22315 13568
rect 22339 13620 22395 13622
rect 22339 13568 22391 13620
rect 22391 13568 22395 13620
rect 22339 13566 22395 13568
rect 22419 13620 22475 13622
rect 22419 13568 22471 13620
rect 22471 13568 22475 13620
rect 22419 13566 22475 13568
rect 22499 13620 22555 13622
rect 22499 13568 22551 13620
rect 22551 13568 22555 13620
rect 22499 13566 22555 13568
rect 22703 13620 22759 13622
rect 22703 13568 22707 13620
rect 22707 13568 22759 13620
rect 22703 13566 22759 13568
rect 22783 13620 22839 13622
rect 22783 13568 22787 13620
rect 22787 13568 22839 13620
rect 22783 13566 22839 13568
rect 22863 13620 22919 13622
rect 22863 13568 22867 13620
rect 22867 13568 22919 13620
rect 22863 13566 22919 13568
rect 22943 13620 22999 13622
rect 22943 13568 22947 13620
rect 22947 13568 22999 13620
rect 22943 13566 22999 13568
rect 23023 13620 23079 13622
rect 23023 13568 23027 13620
rect 23027 13568 23079 13620
rect 23023 13566 23079 13568
rect 23103 13620 23159 13622
rect 23103 13568 23107 13620
rect 23107 13568 23159 13620
rect 23103 13566 23159 13568
rect 23311 13620 23367 13622
rect 23311 13568 23363 13620
rect 23363 13568 23367 13620
rect 23311 13566 23367 13568
rect 23391 13620 23447 13622
rect 23391 13568 23443 13620
rect 23443 13568 23447 13620
rect 23391 13566 23447 13568
rect 23471 13620 23527 13622
rect 23471 13568 23523 13620
rect 23523 13568 23527 13620
rect 23471 13566 23527 13568
rect 23551 13620 23607 13622
rect 23551 13568 23603 13620
rect 23603 13568 23607 13620
rect 23551 13566 23607 13568
rect 23631 13620 23687 13622
rect 23631 13568 23683 13620
rect 23683 13568 23687 13620
rect 23631 13566 23687 13568
rect 23711 13620 23767 13622
rect 23711 13568 23763 13620
rect 23763 13568 23767 13620
rect 23711 13566 23767 13568
rect 23915 13620 23971 13622
rect 23915 13568 23919 13620
rect 23919 13568 23971 13620
rect 23915 13566 23971 13568
rect 23995 13620 24051 13622
rect 23995 13568 23999 13620
rect 23999 13568 24051 13620
rect 23995 13566 24051 13568
rect 24075 13620 24131 13622
rect 24075 13568 24079 13620
rect 24079 13568 24131 13620
rect 24075 13566 24131 13568
rect 24155 13620 24211 13622
rect 24155 13568 24159 13620
rect 24159 13568 24211 13620
rect 24155 13566 24211 13568
rect 24235 13620 24291 13622
rect 24235 13568 24239 13620
rect 24239 13568 24291 13620
rect 24235 13566 24291 13568
rect 24315 13620 24371 13622
rect 24315 13568 24319 13620
rect 24319 13568 24371 13620
rect 24315 13566 24371 13568
rect 24523 13620 24579 13622
rect 24523 13568 24575 13620
rect 24575 13568 24579 13620
rect 24523 13566 24579 13568
rect 24603 13620 24659 13622
rect 24603 13568 24655 13620
rect 24655 13568 24659 13620
rect 24603 13566 24659 13568
rect 24683 13620 24739 13622
rect 24683 13568 24735 13620
rect 24735 13568 24739 13620
rect 24683 13566 24739 13568
rect 24763 13620 24819 13622
rect 24763 13568 24815 13620
rect 24815 13568 24819 13620
rect 24763 13566 24819 13568
rect 24843 13620 24899 13622
rect 24843 13568 24895 13620
rect 24895 13568 24899 13620
rect 24843 13566 24899 13568
rect 24923 13620 24979 13622
rect 24923 13568 24975 13620
rect 24975 13568 24979 13620
rect 24923 13566 24979 13568
rect 25127 13620 25183 13622
rect 25127 13568 25131 13620
rect 25131 13568 25183 13620
rect 25127 13566 25183 13568
rect 25207 13620 25263 13622
rect 25207 13568 25211 13620
rect 25211 13568 25263 13620
rect 25207 13566 25263 13568
rect 25287 13620 25343 13622
rect 25287 13568 25291 13620
rect 25291 13568 25343 13620
rect 25287 13566 25343 13568
rect 25367 13620 25423 13622
rect 25367 13568 25371 13620
rect 25371 13568 25423 13620
rect 25367 13566 25423 13568
rect 25447 13620 25503 13622
rect 25447 13568 25451 13620
rect 25451 13568 25503 13620
rect 25447 13566 25503 13568
rect 25527 13620 25583 13622
rect 25527 13568 25531 13620
rect 25531 13568 25583 13620
rect 25527 13566 25583 13568
rect 25735 13620 25791 13622
rect 25735 13568 25787 13620
rect 25787 13568 25791 13620
rect 25735 13566 25791 13568
rect 25815 13620 25871 13622
rect 25815 13568 25867 13620
rect 25867 13568 25871 13620
rect 25815 13566 25871 13568
rect 25895 13620 25951 13622
rect 25895 13568 25947 13620
rect 25947 13568 25951 13620
rect 25895 13566 25951 13568
rect 25975 13620 26031 13622
rect 25975 13568 26027 13620
rect 26027 13568 26031 13620
rect 25975 13566 26031 13568
rect 26055 13620 26111 13622
rect 26055 13568 26107 13620
rect 26107 13568 26111 13620
rect 26055 13566 26111 13568
rect 26135 13620 26191 13622
rect 26135 13568 26187 13620
rect 26187 13568 26191 13620
rect 26135 13566 26191 13568
rect 26472 13564 26528 13566
rect 26472 13512 26474 13564
rect 26474 13512 26526 13564
rect 26526 13512 26528 13564
rect 26472 13510 26528 13512
rect 19768 13420 19824 13422
rect 19768 13368 19770 13420
rect 19770 13368 19822 13420
rect 19822 13368 19824 13420
rect 19768 13366 19824 13368
rect 3066 13151 3122 13153
rect 3066 13099 3068 13151
rect 3068 13099 3120 13151
rect 3120 13099 3122 13151
rect 20229 13395 20285 13397
rect 20229 13343 20231 13395
rect 20231 13343 20283 13395
rect 20283 13343 20285 13395
rect 20229 13341 20285 13343
rect 26477 13420 26533 13422
rect 26477 13368 26479 13420
rect 26479 13368 26531 13420
rect 26531 13368 26533 13420
rect 26477 13366 26533 13368
rect 19769 13268 19825 13270
rect 19769 13216 19771 13268
rect 19771 13216 19823 13268
rect 19823 13216 19825 13268
rect 19769 13214 19825 13216
rect 26478 13268 26534 13270
rect 26478 13216 26480 13268
rect 26480 13216 26532 13268
rect 26532 13216 26534 13268
rect 26478 13214 26534 13216
rect 3066 13097 3122 13099
rect 3162 13142 3218 13144
rect 3162 13090 3166 13142
rect 3166 13090 3218 13142
rect 3162 13088 3218 13090
rect 3242 13142 3298 13144
rect 3242 13090 3246 13142
rect 3246 13090 3298 13142
rect 3242 13088 3298 13090
rect 3322 13142 3378 13144
rect 3322 13090 3326 13142
rect 3326 13090 3378 13142
rect 3322 13088 3378 13090
rect 3402 13142 3458 13144
rect 3402 13090 3406 13142
rect 3406 13090 3458 13142
rect 3402 13088 3458 13090
rect 3482 13142 3538 13144
rect 3482 13090 3486 13142
rect 3486 13090 3538 13142
rect 3482 13088 3538 13090
rect 3562 13142 3618 13144
rect 3562 13090 3566 13142
rect 3566 13090 3618 13142
rect 3562 13088 3618 13090
rect 3894 13145 3950 13147
rect 3894 13093 3898 13145
rect 3898 13093 3950 13145
rect 3894 13091 3950 13093
rect 3974 13145 4030 13147
rect 3974 13093 3978 13145
rect 3978 13093 4030 13145
rect 3974 13091 4030 13093
rect 4054 13145 4110 13147
rect 4054 13093 4058 13145
rect 4058 13093 4110 13145
rect 4054 13091 4110 13093
rect 4134 13145 4190 13147
rect 4134 13093 4138 13145
rect 4138 13093 4190 13145
rect 4134 13091 4190 13093
rect 4214 13145 4270 13147
rect 4214 13093 4218 13145
rect 4218 13093 4270 13145
rect 4214 13091 4270 13093
rect 4294 13145 4350 13147
rect 4294 13093 4298 13145
rect 4298 13093 4350 13145
rect 4294 13091 4350 13093
rect 4502 13145 4558 13147
rect 4502 13093 4554 13145
rect 4554 13093 4558 13145
rect 4502 13091 4558 13093
rect 4582 13145 4638 13147
rect 4582 13093 4634 13145
rect 4634 13093 4638 13145
rect 4582 13091 4638 13093
rect 4662 13145 4718 13147
rect 4662 13093 4714 13145
rect 4714 13093 4718 13145
rect 4662 13091 4718 13093
rect 4742 13145 4798 13147
rect 4742 13093 4794 13145
rect 4794 13093 4798 13145
rect 4742 13091 4798 13093
rect 4822 13145 4878 13147
rect 4822 13093 4874 13145
rect 4874 13093 4878 13145
rect 4822 13091 4878 13093
rect 4902 13145 4958 13147
rect 4902 13093 4954 13145
rect 4954 13093 4958 13145
rect 4902 13091 4958 13093
rect 5106 13145 5162 13147
rect 5106 13093 5110 13145
rect 5110 13093 5162 13145
rect 5106 13091 5162 13093
rect 5186 13145 5242 13147
rect 5186 13093 5190 13145
rect 5190 13093 5242 13145
rect 5186 13091 5242 13093
rect 5266 13145 5322 13147
rect 5266 13093 5270 13145
rect 5270 13093 5322 13145
rect 5266 13091 5322 13093
rect 5346 13145 5402 13147
rect 5346 13093 5350 13145
rect 5350 13093 5402 13145
rect 5346 13091 5402 13093
rect 5426 13145 5482 13147
rect 5426 13093 5430 13145
rect 5430 13093 5482 13145
rect 5426 13091 5482 13093
rect 5506 13145 5562 13147
rect 5506 13093 5510 13145
rect 5510 13093 5562 13145
rect 5506 13091 5562 13093
rect 5714 13145 5770 13147
rect 5714 13093 5766 13145
rect 5766 13093 5770 13145
rect 5714 13091 5770 13093
rect 5794 13145 5850 13147
rect 5794 13093 5846 13145
rect 5846 13093 5850 13145
rect 5794 13091 5850 13093
rect 5874 13145 5930 13147
rect 5874 13093 5926 13145
rect 5926 13093 5930 13145
rect 5874 13091 5930 13093
rect 5954 13145 6010 13147
rect 5954 13093 6006 13145
rect 6006 13093 6010 13145
rect 5954 13091 6010 13093
rect 6034 13145 6090 13147
rect 6034 13093 6086 13145
rect 6086 13093 6090 13145
rect 6034 13091 6090 13093
rect 6114 13145 6170 13147
rect 6114 13093 6166 13145
rect 6166 13093 6170 13145
rect 6114 13091 6170 13093
rect 6318 13145 6374 13147
rect 6318 13093 6322 13145
rect 6322 13093 6374 13145
rect 6318 13091 6374 13093
rect 6398 13145 6454 13147
rect 6398 13093 6402 13145
rect 6402 13093 6454 13145
rect 6398 13091 6454 13093
rect 6478 13145 6534 13147
rect 6478 13093 6482 13145
rect 6482 13093 6534 13145
rect 6478 13091 6534 13093
rect 6558 13145 6614 13147
rect 6558 13093 6562 13145
rect 6562 13093 6614 13145
rect 6558 13091 6614 13093
rect 6638 13145 6694 13147
rect 6638 13093 6642 13145
rect 6642 13093 6694 13145
rect 6638 13091 6694 13093
rect 6718 13145 6774 13147
rect 6718 13093 6722 13145
rect 6722 13093 6774 13145
rect 6718 13091 6774 13093
rect 6926 13145 6982 13147
rect 6926 13093 6978 13145
rect 6978 13093 6982 13145
rect 6926 13091 6982 13093
rect 7006 13145 7062 13147
rect 7006 13093 7058 13145
rect 7058 13093 7062 13145
rect 7006 13091 7062 13093
rect 7086 13145 7142 13147
rect 7086 13093 7138 13145
rect 7138 13093 7142 13145
rect 7086 13091 7142 13093
rect 7166 13145 7222 13147
rect 7166 13093 7218 13145
rect 7218 13093 7222 13145
rect 7166 13091 7222 13093
rect 7246 13145 7302 13147
rect 7246 13093 7298 13145
rect 7298 13093 7302 13145
rect 7246 13091 7302 13093
rect 7326 13145 7382 13147
rect 7326 13093 7378 13145
rect 7378 13093 7382 13145
rect 7326 13091 7382 13093
rect 7530 13145 7586 13147
rect 7530 13093 7534 13145
rect 7534 13093 7586 13145
rect 7530 13091 7586 13093
rect 7610 13145 7666 13147
rect 7610 13093 7614 13145
rect 7614 13093 7666 13145
rect 7610 13091 7666 13093
rect 7690 13145 7746 13147
rect 7690 13093 7694 13145
rect 7694 13093 7746 13145
rect 7690 13091 7746 13093
rect 7770 13145 7826 13147
rect 7770 13093 7774 13145
rect 7774 13093 7826 13145
rect 7770 13091 7826 13093
rect 7850 13145 7906 13147
rect 7850 13093 7854 13145
rect 7854 13093 7906 13145
rect 7850 13091 7906 13093
rect 7930 13145 7986 13147
rect 7930 13093 7934 13145
rect 7934 13093 7986 13145
rect 7930 13091 7986 13093
rect 8138 13145 8194 13147
rect 8138 13093 8190 13145
rect 8190 13093 8194 13145
rect 8138 13091 8194 13093
rect 8218 13145 8274 13147
rect 8218 13093 8270 13145
rect 8270 13093 8274 13145
rect 8218 13091 8274 13093
rect 8298 13145 8354 13147
rect 8298 13093 8350 13145
rect 8350 13093 8354 13145
rect 8298 13091 8354 13093
rect 8378 13145 8434 13147
rect 8378 13093 8430 13145
rect 8430 13093 8434 13145
rect 8378 13091 8434 13093
rect 8458 13145 8514 13147
rect 8458 13093 8510 13145
rect 8510 13093 8514 13145
rect 8458 13091 8514 13093
rect 8538 13145 8594 13147
rect 8538 13093 8590 13145
rect 8590 13093 8594 13145
rect 8538 13091 8594 13093
rect 20229 13203 20285 13205
rect 20229 13151 20231 13203
rect 20231 13151 20283 13203
rect 20283 13151 20285 13203
rect 20229 13149 20285 13151
rect 2449 12546 2505 12548
rect 2449 12494 2451 12546
rect 2451 12494 2503 12546
rect 2503 12494 2505 12546
rect 2449 12492 2505 12494
rect 2580 12545 2636 12547
rect 2580 12493 2582 12545
rect 2582 12493 2634 12545
rect 2634 12493 2636 12545
rect 2580 12491 2636 12493
rect 2724 12546 2780 12548
rect 2724 12494 2726 12546
rect 2726 12494 2778 12546
rect 2778 12494 2780 12546
rect 2724 12492 2780 12494
rect 8875 13089 8931 13091
rect 8875 13037 8877 13089
rect 8877 13037 8929 13089
rect 8929 13037 8931 13089
rect 8875 13035 8931 13037
rect 19769 13098 19825 13100
rect 19769 13046 19771 13098
rect 19771 13046 19823 13098
rect 19823 13046 19825 13098
rect 19769 13044 19825 13046
rect 26478 13098 26534 13100
rect 26478 13046 26480 13098
rect 26480 13046 26532 13098
rect 26532 13046 26534 13098
rect 26478 13044 26534 13046
rect 13337 13021 13393 13023
rect 13337 12969 13339 13021
rect 13339 12969 13391 13021
rect 13391 12969 13393 13021
rect 13337 12967 13393 12969
rect 13468 13020 13524 13022
rect 13468 12968 13470 13020
rect 13470 12968 13522 13020
rect 13522 12968 13524 13020
rect 13468 12966 13524 12968
rect 13612 13021 13668 13023
rect 13612 12969 13614 13021
rect 13614 12969 13666 13021
rect 13666 12969 13668 13021
rect 13612 12967 13668 12969
rect 20046 13021 20102 13023
rect 20046 12969 20048 13021
rect 20048 12969 20100 13021
rect 20100 12969 20102 13021
rect 20046 12967 20102 12969
rect 20177 13020 20233 13022
rect 20177 12968 20179 13020
rect 20179 12968 20231 13020
rect 20231 12968 20233 13020
rect 20177 12966 20233 12968
rect 20321 13021 20377 13023
rect 20321 12969 20323 13021
rect 20323 12969 20375 13021
rect 20375 12969 20377 13021
rect 20321 12967 20377 12969
rect 8880 12945 8936 12947
rect 8880 12893 8882 12945
rect 8882 12893 8934 12945
rect 8934 12893 8936 12945
rect 8880 12891 8936 12893
rect 19768 12941 19824 12943
rect 19768 12889 19770 12941
rect 19770 12889 19822 12941
rect 19822 12889 19824 12941
rect 19768 12887 19824 12889
rect 26477 12941 26533 12943
rect 26477 12889 26479 12941
rect 26479 12889 26531 12941
rect 26531 12889 26533 12941
rect 26477 12887 26533 12889
rect 8881 12793 8937 12795
rect 8881 12741 8883 12793
rect 8883 12741 8935 12793
rect 8935 12741 8937 12793
rect 8881 12739 8937 12741
rect 8881 12623 8937 12625
rect 8881 12571 8883 12623
rect 8883 12571 8935 12623
rect 8935 12571 8937 12623
rect 8881 12569 8937 12571
rect 19686 12699 19742 12701
rect 19686 12647 19688 12699
rect 19688 12647 19740 12699
rect 19740 12647 19742 12699
rect 19686 12645 19742 12647
rect 26395 12699 26451 12701
rect 26395 12647 26397 12699
rect 26397 12647 26449 12699
rect 26449 12647 26451 12699
rect 26395 12645 26451 12647
rect 10985 12554 11041 12556
rect 10985 12502 10987 12554
rect 10987 12502 11039 12554
rect 11039 12502 11041 12554
rect 10985 12500 11041 12502
rect 11172 12556 11228 12558
rect 11172 12504 11174 12556
rect 11174 12504 11226 12556
rect 11226 12504 11228 12556
rect 11172 12502 11228 12504
rect 11357 12558 11413 12560
rect 11357 12506 11359 12558
rect 11359 12506 11411 12558
rect 11411 12506 11413 12558
rect 11357 12504 11413 12506
rect 11542 12559 11598 12561
rect 11542 12507 11544 12559
rect 11544 12507 11596 12559
rect 11596 12507 11598 12559
rect 11542 12505 11598 12507
rect 11745 12561 11801 12563
rect 11745 12509 11747 12561
rect 11747 12509 11799 12561
rect 11799 12509 11801 12561
rect 11745 12507 11801 12509
rect 11930 12563 11986 12565
rect 11930 12511 11932 12563
rect 11932 12511 11984 12563
rect 11984 12511 11986 12563
rect 11930 12509 11986 12511
rect 12129 12565 12185 12567
rect 12129 12513 12131 12565
rect 12131 12513 12183 12565
rect 12183 12513 12185 12565
rect 12129 12511 12185 12513
rect 12331 12564 12387 12566
rect 12331 12512 12333 12564
rect 12333 12512 12385 12564
rect 12385 12512 12387 12564
rect 12331 12510 12387 12512
rect 12541 12567 12597 12569
rect 12541 12515 12543 12567
rect 12543 12515 12595 12567
rect 12595 12515 12597 12567
rect 12541 12513 12597 12515
rect 12765 12567 12821 12569
rect 12765 12515 12767 12567
rect 12767 12515 12819 12567
rect 12819 12515 12821 12567
rect 12765 12513 12821 12515
rect 12971 12566 13027 12568
rect 12971 12514 12973 12566
rect 12973 12514 13025 12566
rect 13025 12514 13027 12566
rect 12971 12512 13027 12514
rect 13192 12565 13248 12567
rect 13192 12513 13194 12565
rect 13194 12513 13246 12565
rect 13246 12513 13248 12565
rect 13192 12511 13248 12513
rect 13355 12475 13411 12477
rect 8880 12466 8936 12468
rect 8880 12414 8882 12466
rect 8882 12414 8934 12466
rect 8934 12414 8936 12466
rect 8880 12412 8936 12414
rect 13355 12423 13357 12475
rect 13357 12423 13409 12475
rect 13409 12423 13411 12475
rect 13355 12421 13411 12423
rect 13475 12475 13531 12477
rect 13475 12423 13477 12475
rect 13477 12423 13529 12475
rect 13529 12423 13531 12475
rect 13475 12421 13531 12423
rect 13618 12475 13674 12477
rect 13618 12423 13620 12475
rect 13620 12423 13672 12475
rect 13672 12423 13674 12475
rect 13618 12421 13674 12423
rect 8798 12224 8854 12226
rect 8798 12172 8800 12224
rect 8800 12172 8852 12224
rect 8852 12172 8854 12224
rect 8798 12170 8854 12172
rect 9175 12276 9231 12278
rect 9175 12224 9177 12276
rect 9177 12224 9229 12276
rect 9229 12224 9231 12276
rect 9175 12222 9231 12224
rect 2467 12000 2523 12002
rect 2467 11948 2469 12000
rect 2469 11948 2521 12000
rect 2521 11948 2523 12000
rect 2467 11946 2523 11948
rect 2587 12000 2643 12002
rect 2587 11948 2589 12000
rect 2589 11948 2641 12000
rect 2641 11948 2643 12000
rect 2587 11946 2643 11948
rect 2730 12000 2786 12002
rect 2730 11948 2732 12000
rect 2732 11948 2784 12000
rect 2784 11948 2786 12000
rect 2730 11946 2786 11948
rect 3548 11900 3612 11964
rect 4280 11903 4344 11967
rect 4508 11903 4572 11967
rect 5492 11903 5556 11967
rect 5720 11903 5784 11967
rect 6704 11903 6768 11967
rect 6932 11903 6996 11967
rect 7916 11903 7980 11967
rect 8144 11903 8208 11967
rect 8886 11963 8942 11965
rect 8886 11911 8888 11963
rect 8888 11911 8940 11963
rect 8940 11911 8942 11963
rect 8886 11909 8942 11911
rect 10916 11882 10972 11883
rect 10916 11829 10917 11882
rect 10917 11829 10970 11882
rect 10970 11829 10972 11882
rect 10916 11827 10972 11829
rect 11116 11885 11172 11886
rect 11116 11832 11117 11885
rect 11117 11832 11170 11885
rect 11170 11832 11172 11885
rect 11116 11830 11172 11832
rect 11352 11883 11408 11884
rect 11352 11830 11353 11883
rect 11353 11830 11406 11883
rect 11406 11830 11408 11883
rect 11352 11828 11408 11830
rect 3904 11701 3968 11765
rect 4636 11701 4700 11765
rect 4854 11701 4918 11765
rect 5848 11701 5912 11765
rect 6066 11701 6130 11765
rect 7186 11701 7250 11765
rect 7404 11701 7468 11765
rect 8138 11701 8202 11765
rect 8886 11760 8942 11762
rect 8886 11708 8888 11760
rect 8888 11708 8940 11760
rect 8940 11708 8942 11760
rect 8886 11706 8942 11708
rect 8795 11498 8851 11500
rect 8795 11446 8797 11498
rect 8797 11446 8849 11498
rect 8849 11446 8851 11498
rect 8795 11444 8851 11446
rect 9198 11519 9254 11521
rect 9198 11467 9200 11519
rect 9200 11467 9252 11519
rect 9252 11467 9254 11519
rect 9198 11465 9254 11467
rect 3052 10573 3108 10575
rect 3052 10521 3054 10573
rect 3054 10521 3106 10573
rect 3106 10521 3108 10573
rect 3052 10519 3108 10521
rect 3594 10576 3650 10578
rect 3594 10524 3596 10576
rect 3596 10524 3648 10576
rect 3648 10524 3650 10576
rect 3594 10522 3650 10524
rect 3674 10576 3730 10578
rect 3674 10524 3676 10576
rect 3676 10524 3728 10576
rect 3728 10524 3730 10576
rect 3674 10522 3730 10524
rect 3754 10576 3810 10578
rect 3754 10524 3756 10576
rect 3756 10524 3808 10576
rect 3808 10524 3810 10576
rect 3754 10522 3810 10524
rect 3834 10576 3890 10578
rect 3834 10524 3836 10576
rect 3836 10524 3888 10576
rect 3888 10524 3890 10576
rect 3834 10522 3890 10524
rect 4326 10576 4382 10578
rect 4326 10524 4328 10576
rect 4328 10524 4380 10576
rect 4380 10524 4382 10576
rect 4326 10522 4382 10524
rect 4406 10576 4462 10578
rect 4406 10524 4408 10576
rect 4408 10524 4460 10576
rect 4460 10524 4462 10576
rect 4406 10522 4462 10524
rect 4486 10576 4542 10578
rect 4486 10524 4488 10576
rect 4488 10524 4540 10576
rect 4540 10524 4542 10576
rect 4486 10522 4542 10524
rect 4566 10576 4622 10578
rect 4566 10524 4568 10576
rect 4568 10524 4620 10576
rect 4620 10524 4622 10576
rect 4566 10522 4622 10524
rect 4932 10576 4988 10578
rect 4932 10524 4934 10576
rect 4934 10524 4986 10576
rect 4986 10524 4988 10576
rect 4932 10522 4988 10524
rect 5012 10576 5068 10578
rect 5012 10524 5014 10576
rect 5014 10524 5066 10576
rect 5066 10524 5068 10576
rect 5012 10522 5068 10524
rect 5092 10576 5148 10578
rect 5092 10524 5094 10576
rect 5094 10524 5146 10576
rect 5146 10524 5148 10576
rect 5092 10522 5148 10524
rect 5172 10576 5228 10578
rect 5172 10524 5174 10576
rect 5174 10524 5226 10576
rect 5226 10524 5228 10576
rect 5172 10522 5228 10524
rect 5538 10576 5594 10578
rect 5538 10524 5540 10576
rect 5540 10524 5592 10576
rect 5592 10524 5594 10576
rect 5538 10522 5594 10524
rect 5618 10576 5674 10578
rect 5618 10524 5620 10576
rect 5620 10524 5672 10576
rect 5672 10524 5674 10576
rect 5618 10522 5674 10524
rect 5698 10576 5754 10578
rect 5698 10524 5700 10576
rect 5700 10524 5752 10576
rect 5752 10524 5754 10576
rect 5698 10522 5754 10524
rect 5778 10576 5834 10578
rect 5778 10524 5780 10576
rect 5780 10524 5832 10576
rect 5832 10524 5834 10576
rect 5778 10522 5834 10524
rect 6144 10576 6200 10578
rect 6144 10524 6146 10576
rect 6146 10524 6198 10576
rect 6198 10524 6200 10576
rect 6144 10522 6200 10524
rect 6224 10576 6280 10578
rect 6224 10524 6226 10576
rect 6226 10524 6278 10576
rect 6278 10524 6280 10576
rect 6224 10522 6280 10524
rect 6304 10576 6360 10578
rect 6304 10524 6306 10576
rect 6306 10524 6358 10576
rect 6358 10524 6360 10576
rect 6304 10522 6360 10524
rect 6384 10576 6440 10578
rect 6384 10524 6386 10576
rect 6386 10524 6438 10576
rect 6438 10524 6440 10576
rect 6384 10522 6440 10524
rect 6876 10576 6932 10578
rect 6876 10524 6878 10576
rect 6878 10524 6930 10576
rect 6930 10524 6932 10576
rect 6876 10522 6932 10524
rect 6956 10576 7012 10578
rect 6956 10524 6958 10576
rect 6958 10524 7010 10576
rect 7010 10524 7012 10576
rect 6956 10522 7012 10524
rect 7036 10576 7092 10578
rect 7036 10524 7038 10576
rect 7038 10524 7090 10576
rect 7090 10524 7092 10576
rect 7036 10522 7092 10524
rect 7116 10576 7172 10578
rect 7116 10524 7118 10576
rect 7118 10524 7170 10576
rect 7170 10524 7172 10576
rect 7116 10522 7172 10524
rect 7482 10576 7538 10578
rect 7482 10524 7484 10576
rect 7484 10524 7536 10576
rect 7536 10524 7538 10576
rect 7482 10522 7538 10524
rect 7562 10576 7618 10578
rect 7562 10524 7564 10576
rect 7564 10524 7616 10576
rect 7616 10524 7618 10576
rect 7562 10522 7618 10524
rect 7642 10576 7698 10578
rect 7642 10524 7644 10576
rect 7644 10524 7696 10576
rect 7696 10524 7698 10576
rect 7642 10522 7698 10524
rect 7722 10576 7778 10578
rect 7722 10524 7724 10576
rect 7724 10524 7776 10576
rect 7776 10524 7778 10576
rect 7722 10522 7778 10524
rect 8216 10576 8272 10578
rect 8216 10524 8218 10576
rect 8218 10524 8270 10576
rect 8270 10524 8272 10576
rect 8216 10522 8272 10524
rect 8296 10576 8352 10578
rect 8296 10524 8298 10576
rect 8298 10524 8350 10576
rect 8350 10524 8352 10576
rect 8296 10522 8352 10524
rect 8376 10576 8432 10578
rect 8376 10524 8378 10576
rect 8378 10524 8430 10576
rect 8430 10524 8432 10576
rect 8376 10522 8432 10524
rect 8456 10576 8512 10578
rect 8456 10524 8458 10576
rect 8458 10524 8510 10576
rect 8510 10524 8512 10576
rect 8456 10522 8512 10524
rect 3052 10125 3108 10127
rect 3052 10073 3054 10125
rect 3054 10073 3106 10125
rect 3106 10073 3108 10125
rect 3052 10071 3108 10073
rect 3594 10122 3650 10124
rect 3594 10070 3596 10122
rect 3596 10070 3648 10122
rect 3648 10070 3650 10122
rect 3594 10068 3650 10070
rect 3674 10122 3730 10124
rect 3674 10070 3676 10122
rect 3676 10070 3728 10122
rect 3728 10070 3730 10122
rect 3674 10068 3730 10070
rect 3754 10122 3810 10124
rect 3754 10070 3756 10122
rect 3756 10070 3808 10122
rect 3808 10070 3810 10122
rect 3754 10068 3810 10070
rect 3834 10122 3890 10124
rect 3834 10070 3836 10122
rect 3836 10070 3888 10122
rect 3888 10070 3890 10122
rect 3834 10068 3890 10070
rect 4326 10122 4382 10124
rect 4326 10070 4328 10122
rect 4328 10070 4380 10122
rect 4380 10070 4382 10122
rect 4326 10068 4382 10070
rect 4406 10122 4462 10124
rect 4406 10070 4408 10122
rect 4408 10070 4460 10122
rect 4460 10070 4462 10122
rect 4406 10068 4462 10070
rect 4486 10122 4542 10124
rect 4486 10070 4488 10122
rect 4488 10070 4540 10122
rect 4540 10070 4542 10122
rect 4486 10068 4542 10070
rect 4566 10122 4622 10124
rect 4566 10070 4568 10122
rect 4568 10070 4620 10122
rect 4620 10070 4622 10122
rect 4566 10068 4622 10070
rect 4932 10122 4988 10124
rect 4932 10070 4934 10122
rect 4934 10070 4986 10122
rect 4986 10070 4988 10122
rect 4932 10068 4988 10070
rect 5012 10122 5068 10124
rect 5012 10070 5014 10122
rect 5014 10070 5066 10122
rect 5066 10070 5068 10122
rect 5012 10068 5068 10070
rect 5092 10122 5148 10124
rect 5092 10070 5094 10122
rect 5094 10070 5146 10122
rect 5146 10070 5148 10122
rect 5092 10068 5148 10070
rect 5172 10122 5228 10124
rect 5172 10070 5174 10122
rect 5174 10070 5226 10122
rect 5226 10070 5228 10122
rect 5172 10068 5228 10070
rect 5538 10122 5594 10124
rect 5538 10070 5540 10122
rect 5540 10070 5592 10122
rect 5592 10070 5594 10122
rect 5538 10068 5594 10070
rect 5618 10122 5674 10124
rect 5618 10070 5620 10122
rect 5620 10070 5672 10122
rect 5672 10070 5674 10122
rect 5618 10068 5674 10070
rect 5698 10122 5754 10124
rect 5698 10070 5700 10122
rect 5700 10070 5752 10122
rect 5752 10070 5754 10122
rect 5698 10068 5754 10070
rect 5778 10122 5834 10124
rect 5778 10070 5780 10122
rect 5780 10070 5832 10122
rect 5832 10070 5834 10122
rect 5778 10068 5834 10070
rect 6144 10122 6200 10124
rect 6144 10070 6146 10122
rect 6146 10070 6198 10122
rect 6198 10070 6200 10122
rect 6144 10068 6200 10070
rect 6224 10122 6280 10124
rect 6224 10070 6226 10122
rect 6226 10070 6278 10122
rect 6278 10070 6280 10122
rect 6224 10068 6280 10070
rect 6304 10122 6360 10124
rect 6304 10070 6306 10122
rect 6306 10070 6358 10122
rect 6358 10070 6360 10122
rect 6304 10068 6360 10070
rect 6384 10122 6440 10124
rect 6384 10070 6386 10122
rect 6386 10070 6438 10122
rect 6438 10070 6440 10122
rect 6384 10068 6440 10070
rect 6876 10122 6932 10124
rect 6876 10070 6878 10122
rect 6878 10070 6930 10122
rect 6930 10070 6932 10122
rect 6876 10068 6932 10070
rect 6956 10122 7012 10124
rect 6956 10070 6958 10122
rect 6958 10070 7010 10122
rect 7010 10070 7012 10122
rect 6956 10068 7012 10070
rect 7036 10122 7092 10124
rect 7036 10070 7038 10122
rect 7038 10070 7090 10122
rect 7090 10070 7092 10122
rect 7036 10068 7092 10070
rect 7116 10122 7172 10124
rect 7116 10070 7118 10122
rect 7118 10070 7170 10122
rect 7170 10070 7172 10122
rect 7116 10068 7172 10070
rect 7482 10122 7538 10124
rect 7482 10070 7484 10122
rect 7484 10070 7536 10122
rect 7536 10070 7538 10122
rect 7482 10068 7538 10070
rect 7562 10122 7618 10124
rect 7562 10070 7564 10122
rect 7564 10070 7616 10122
rect 7616 10070 7618 10122
rect 7562 10068 7618 10070
rect 7642 10122 7698 10124
rect 7642 10070 7644 10122
rect 7644 10070 7696 10122
rect 7696 10070 7698 10122
rect 7642 10068 7698 10070
rect 7722 10122 7778 10124
rect 7722 10070 7724 10122
rect 7724 10070 7776 10122
rect 7776 10070 7778 10122
rect 7722 10068 7778 10070
rect 8216 10122 8272 10124
rect 8216 10070 8218 10122
rect 8218 10070 8270 10122
rect 8270 10070 8272 10122
rect 8216 10068 8272 10070
rect 8296 10122 8352 10124
rect 8296 10070 8298 10122
rect 8298 10070 8350 10122
rect 8350 10070 8352 10122
rect 8296 10068 8352 10070
rect 8376 10122 8432 10124
rect 8376 10070 8378 10122
rect 8378 10070 8430 10122
rect 8430 10070 8432 10122
rect 8376 10068 8432 10070
rect 8456 10122 8512 10124
rect 8456 10070 8458 10122
rect 8458 10070 8510 10122
rect 8510 10070 8512 10122
rect 8456 10068 8512 10070
rect 8795 9200 8851 9202
rect 8795 9148 8797 9200
rect 8797 9148 8849 9200
rect 8849 9148 8851 9200
rect 8795 9146 8851 9148
rect 9223 9159 9279 9161
rect 9223 9107 9225 9159
rect 9225 9107 9277 9159
rect 9277 9107 9279 9159
rect 9223 9105 9279 9107
rect 9700 9159 9756 9161
rect 9700 9107 9702 9159
rect 9702 9107 9754 9159
rect 9754 9107 9756 9159
rect 9700 9105 9756 9107
rect 10120 9148 10176 9150
rect 10120 9096 10122 9148
rect 10122 9096 10174 9148
rect 10174 9096 10176 9148
rect 10120 9094 10176 9096
rect 2467 8698 2523 8700
rect 2467 8646 2469 8698
rect 2469 8646 2521 8698
rect 2521 8646 2523 8698
rect 2467 8644 2523 8646
rect 2587 8698 2643 8700
rect 2587 8646 2589 8698
rect 2589 8646 2641 8698
rect 2641 8646 2643 8698
rect 2587 8644 2643 8646
rect 2730 8698 2786 8700
rect 2730 8646 2732 8698
rect 2732 8646 2784 8698
rect 2784 8646 2786 8698
rect 2730 8644 2786 8646
rect 3904 8881 3968 8945
rect 4636 8881 4700 8945
rect 4854 8881 4918 8945
rect 5848 8881 5912 8945
rect 6066 8881 6130 8945
rect 7186 8881 7250 8945
rect 7404 8881 7468 8945
rect 8138 8881 8202 8945
rect 8886 8938 8942 8940
rect 8886 8886 8888 8938
rect 8888 8886 8940 8938
rect 8940 8886 8942 8938
rect 8886 8884 8942 8886
rect 11785 11877 11841 11878
rect 11785 11824 11786 11877
rect 11786 11824 11839 11877
rect 11839 11824 11841 11877
rect 11785 11822 11841 11824
rect 11986 11878 12042 11879
rect 11986 11825 11987 11878
rect 11987 11825 12040 11878
rect 12040 11825 12042 11878
rect 11986 11823 12042 11825
rect 12172 11876 12228 11877
rect 12172 11823 12173 11876
rect 12173 11823 12226 11876
rect 12226 11823 12228 11876
rect 12172 11821 12228 11823
rect 12363 11879 12419 11880
rect 12363 11826 12364 11879
rect 12364 11826 12417 11879
rect 12417 11826 12419 11879
rect 12363 11824 12419 11826
rect 12576 11878 12632 11879
rect 12576 11825 12577 11878
rect 12577 11825 12630 11878
rect 12630 11825 12632 11878
rect 12576 11823 12632 11825
rect 20064 12475 20120 12477
rect 14436 12375 14500 12439
rect 15168 12378 15232 12442
rect 15396 12378 15460 12442
rect 16380 12378 16444 12442
rect 16608 12378 16672 12442
rect 17592 12378 17656 12442
rect 17820 12378 17884 12442
rect 18804 12378 18868 12442
rect 19032 12378 19096 12442
rect 19774 12438 19830 12440
rect 19774 12386 19776 12438
rect 19776 12386 19828 12438
rect 19828 12386 19830 12438
rect 19774 12384 19830 12386
rect 20064 12423 20066 12475
rect 20066 12423 20118 12475
rect 20118 12423 20120 12475
rect 20064 12421 20120 12423
rect 20184 12475 20240 12477
rect 20184 12423 20186 12475
rect 20186 12423 20238 12475
rect 20238 12423 20240 12475
rect 20184 12421 20240 12423
rect 20327 12475 20383 12477
rect 20327 12423 20329 12475
rect 20329 12423 20381 12475
rect 20381 12423 20383 12475
rect 20327 12421 20383 12423
rect 14792 12176 14856 12240
rect 15524 12176 15588 12240
rect 15742 12176 15806 12240
rect 16736 12176 16800 12240
rect 16954 12176 17018 12240
rect 18074 12176 18138 12240
rect 18292 12176 18356 12240
rect 19026 12176 19090 12240
rect 19774 12235 19830 12237
rect 19774 12183 19776 12235
rect 19776 12183 19828 12235
rect 19828 12183 19830 12235
rect 19774 12181 19830 12183
rect 21145 12375 21209 12439
rect 21877 12378 21941 12442
rect 22105 12378 22169 12442
rect 23089 12378 23153 12442
rect 23317 12378 23381 12442
rect 24301 12378 24365 12442
rect 24529 12378 24593 12442
rect 25513 12378 25577 12442
rect 25741 12378 25805 12442
rect 26483 12438 26539 12440
rect 26483 12386 26485 12438
rect 26485 12386 26537 12438
rect 26537 12386 26539 12438
rect 26483 12384 26539 12386
rect 21501 12176 21565 12240
rect 22233 12176 22297 12240
rect 22451 12176 22515 12240
rect 23445 12176 23509 12240
rect 23663 12176 23727 12240
rect 24783 12176 24847 12240
rect 25001 12176 25065 12240
rect 25735 12176 25799 12240
rect 26483 12235 26539 12237
rect 26483 12183 26485 12235
rect 26485 12183 26537 12235
rect 26537 12183 26539 12235
rect 26483 12181 26539 12183
rect 10933 11257 10989 11259
rect 10933 11205 10935 11257
rect 10935 11205 10987 11257
rect 10987 11205 10989 11257
rect 10933 11203 10989 11205
rect 11121 11254 11177 11256
rect 11121 11202 11123 11254
rect 11123 11202 11175 11254
rect 11175 11202 11177 11254
rect 11121 11200 11177 11202
rect 11318 11252 11374 11254
rect 11318 11200 11320 11252
rect 11320 11200 11372 11252
rect 11372 11200 11374 11252
rect 11318 11198 11374 11200
rect 13314 11594 13381 11595
rect 13314 11538 13317 11594
rect 13317 11538 13377 11594
rect 13377 11538 13381 11594
rect 13314 11537 13381 11538
rect 13940 11048 13996 11050
rect 13940 10996 13942 11048
rect 13942 10996 13994 11048
rect 13994 10996 13996 11048
rect 13940 10994 13996 10996
rect 19683 11973 19739 11975
rect 19683 11921 19685 11973
rect 19685 11921 19737 11973
rect 19737 11921 19739 11973
rect 19683 11919 19739 11921
rect 14482 11051 14538 11053
rect 14482 10999 14484 11051
rect 14484 10999 14536 11051
rect 14536 10999 14538 11051
rect 14482 10997 14538 10999
rect 14562 11051 14618 11053
rect 14562 10999 14564 11051
rect 14564 10999 14616 11051
rect 14616 10999 14618 11051
rect 14562 10997 14618 10999
rect 14642 11051 14698 11053
rect 14642 10999 14644 11051
rect 14644 10999 14696 11051
rect 14696 10999 14698 11051
rect 14642 10997 14698 10999
rect 14722 11051 14778 11053
rect 14722 10999 14724 11051
rect 14724 10999 14776 11051
rect 14776 10999 14778 11051
rect 14722 10997 14778 10999
rect 15214 11051 15270 11053
rect 15214 10999 15216 11051
rect 15216 10999 15268 11051
rect 15268 10999 15270 11051
rect 15214 10997 15270 10999
rect 15294 11051 15350 11053
rect 15294 10999 15296 11051
rect 15296 10999 15348 11051
rect 15348 10999 15350 11051
rect 15294 10997 15350 10999
rect 15374 11051 15430 11053
rect 15374 10999 15376 11051
rect 15376 10999 15428 11051
rect 15428 10999 15430 11051
rect 15374 10997 15430 10999
rect 15454 11051 15510 11053
rect 15454 10999 15456 11051
rect 15456 10999 15508 11051
rect 15508 10999 15510 11051
rect 15454 10997 15510 10999
rect 15820 11051 15876 11053
rect 15820 10999 15822 11051
rect 15822 10999 15874 11051
rect 15874 10999 15876 11051
rect 15820 10997 15876 10999
rect 15900 11051 15956 11053
rect 15900 10999 15902 11051
rect 15902 10999 15954 11051
rect 15954 10999 15956 11051
rect 15900 10997 15956 10999
rect 15980 11051 16036 11053
rect 15980 10999 15982 11051
rect 15982 10999 16034 11051
rect 16034 10999 16036 11051
rect 15980 10997 16036 10999
rect 16060 11051 16116 11053
rect 16060 10999 16062 11051
rect 16062 10999 16114 11051
rect 16114 10999 16116 11051
rect 16060 10997 16116 10999
rect 16426 11051 16482 11053
rect 16426 10999 16428 11051
rect 16428 10999 16480 11051
rect 16480 10999 16482 11051
rect 16426 10997 16482 10999
rect 16506 11051 16562 11053
rect 16506 10999 16508 11051
rect 16508 10999 16560 11051
rect 16560 10999 16562 11051
rect 16506 10997 16562 10999
rect 16586 11051 16642 11053
rect 16586 10999 16588 11051
rect 16588 10999 16640 11051
rect 16640 10999 16642 11051
rect 16586 10997 16642 10999
rect 16666 11051 16722 11053
rect 16666 10999 16668 11051
rect 16668 10999 16720 11051
rect 16720 10999 16722 11051
rect 16666 10997 16722 10999
rect 17032 11051 17088 11053
rect 17032 10999 17034 11051
rect 17034 10999 17086 11051
rect 17086 10999 17088 11051
rect 17032 10997 17088 10999
rect 17112 11051 17168 11053
rect 17112 10999 17114 11051
rect 17114 10999 17166 11051
rect 17166 10999 17168 11051
rect 17112 10997 17168 10999
rect 17192 11051 17248 11053
rect 17192 10999 17194 11051
rect 17194 10999 17246 11051
rect 17246 10999 17248 11051
rect 17192 10997 17248 10999
rect 17272 11051 17328 11053
rect 17272 10999 17274 11051
rect 17274 10999 17326 11051
rect 17326 10999 17328 11051
rect 17272 10997 17328 10999
rect 17764 11051 17820 11053
rect 17764 10999 17766 11051
rect 17766 10999 17818 11051
rect 17818 10999 17820 11051
rect 17764 10997 17820 10999
rect 17844 11051 17900 11053
rect 17844 10999 17846 11051
rect 17846 10999 17898 11051
rect 17898 10999 17900 11051
rect 17844 10997 17900 10999
rect 17924 11051 17980 11053
rect 17924 10999 17926 11051
rect 17926 10999 17978 11051
rect 17978 10999 17980 11051
rect 17924 10997 17980 10999
rect 18004 11051 18060 11053
rect 18004 10999 18006 11051
rect 18006 10999 18058 11051
rect 18058 10999 18060 11051
rect 18004 10997 18060 10999
rect 18370 11051 18426 11053
rect 18370 10999 18372 11051
rect 18372 10999 18424 11051
rect 18424 10999 18426 11051
rect 18370 10997 18426 10999
rect 18450 11051 18506 11053
rect 18450 10999 18452 11051
rect 18452 10999 18504 11051
rect 18504 10999 18506 11051
rect 18450 10997 18506 10999
rect 18530 11051 18586 11053
rect 18530 10999 18532 11051
rect 18532 10999 18584 11051
rect 18584 10999 18586 11051
rect 18530 10997 18586 10999
rect 18610 11051 18666 11053
rect 18610 10999 18612 11051
rect 18612 10999 18664 11051
rect 18664 10999 18666 11051
rect 18610 10997 18666 10999
rect 19104 11051 19160 11053
rect 19104 10999 19106 11051
rect 19106 10999 19158 11051
rect 19158 10999 19160 11051
rect 19104 10997 19160 10999
rect 19184 11051 19240 11053
rect 19184 10999 19186 11051
rect 19186 10999 19238 11051
rect 19238 10999 19240 11051
rect 19184 10997 19240 10999
rect 19264 11051 19320 11053
rect 19264 10999 19266 11051
rect 19266 10999 19318 11051
rect 19318 10999 19320 11051
rect 19264 10997 19320 10999
rect 19344 11051 19400 11053
rect 19344 10999 19346 11051
rect 19346 10999 19398 11051
rect 19398 10999 19400 11051
rect 19344 10997 19400 10999
rect 20649 11048 20705 11050
rect 20649 10996 20651 11048
rect 20651 10996 20703 11048
rect 20703 10996 20705 11048
rect 20649 10994 20705 10996
rect 26392 11973 26448 11975
rect 26392 11921 26394 11973
rect 26394 11921 26446 11973
rect 26446 11921 26448 11973
rect 26392 11919 26448 11921
rect 21191 11051 21247 11053
rect 21191 10999 21193 11051
rect 21193 10999 21245 11051
rect 21245 10999 21247 11051
rect 21191 10997 21247 10999
rect 21271 11051 21327 11053
rect 21271 10999 21273 11051
rect 21273 10999 21325 11051
rect 21325 10999 21327 11051
rect 21271 10997 21327 10999
rect 21351 11051 21407 11053
rect 21351 10999 21353 11051
rect 21353 10999 21405 11051
rect 21405 10999 21407 11051
rect 21351 10997 21407 10999
rect 21431 11051 21487 11053
rect 21431 10999 21433 11051
rect 21433 10999 21485 11051
rect 21485 10999 21487 11051
rect 21431 10997 21487 10999
rect 21923 11051 21979 11053
rect 21923 10999 21925 11051
rect 21925 10999 21977 11051
rect 21977 10999 21979 11051
rect 21923 10997 21979 10999
rect 22003 11051 22059 11053
rect 22003 10999 22005 11051
rect 22005 10999 22057 11051
rect 22057 10999 22059 11051
rect 22003 10997 22059 10999
rect 22083 11051 22139 11053
rect 22083 10999 22085 11051
rect 22085 10999 22137 11051
rect 22137 10999 22139 11051
rect 22083 10997 22139 10999
rect 22163 11051 22219 11053
rect 22163 10999 22165 11051
rect 22165 10999 22217 11051
rect 22217 10999 22219 11051
rect 22163 10997 22219 10999
rect 22529 11051 22585 11053
rect 22529 10999 22531 11051
rect 22531 10999 22583 11051
rect 22583 10999 22585 11051
rect 22529 10997 22585 10999
rect 22609 11051 22665 11053
rect 22609 10999 22611 11051
rect 22611 10999 22663 11051
rect 22663 10999 22665 11051
rect 22609 10997 22665 10999
rect 22689 11051 22745 11053
rect 22689 10999 22691 11051
rect 22691 10999 22743 11051
rect 22743 10999 22745 11051
rect 22689 10997 22745 10999
rect 22769 11051 22825 11053
rect 22769 10999 22771 11051
rect 22771 10999 22823 11051
rect 22823 10999 22825 11051
rect 22769 10997 22825 10999
rect 23135 11051 23191 11053
rect 23135 10999 23137 11051
rect 23137 10999 23189 11051
rect 23189 10999 23191 11051
rect 23135 10997 23191 10999
rect 23215 11051 23271 11053
rect 23215 10999 23217 11051
rect 23217 10999 23269 11051
rect 23269 10999 23271 11051
rect 23215 10997 23271 10999
rect 23295 11051 23351 11053
rect 23295 10999 23297 11051
rect 23297 10999 23349 11051
rect 23349 10999 23351 11051
rect 23295 10997 23351 10999
rect 23375 11051 23431 11053
rect 23375 10999 23377 11051
rect 23377 10999 23429 11051
rect 23429 10999 23431 11051
rect 23375 10997 23431 10999
rect 23741 11051 23797 11053
rect 23741 10999 23743 11051
rect 23743 10999 23795 11051
rect 23795 10999 23797 11051
rect 23741 10997 23797 10999
rect 23821 11051 23877 11053
rect 23821 10999 23823 11051
rect 23823 10999 23875 11051
rect 23875 10999 23877 11051
rect 23821 10997 23877 10999
rect 23901 11051 23957 11053
rect 23901 10999 23903 11051
rect 23903 10999 23955 11051
rect 23955 10999 23957 11051
rect 23901 10997 23957 10999
rect 23981 11051 24037 11053
rect 23981 10999 23983 11051
rect 23983 10999 24035 11051
rect 24035 10999 24037 11051
rect 23981 10997 24037 10999
rect 24473 11051 24529 11053
rect 24473 10999 24475 11051
rect 24475 10999 24527 11051
rect 24527 10999 24529 11051
rect 24473 10997 24529 10999
rect 24553 11051 24609 11053
rect 24553 10999 24555 11051
rect 24555 10999 24607 11051
rect 24607 10999 24609 11051
rect 24553 10997 24609 10999
rect 24633 11051 24689 11053
rect 24633 10999 24635 11051
rect 24635 10999 24687 11051
rect 24687 10999 24689 11051
rect 24633 10997 24689 10999
rect 24713 11051 24769 11053
rect 24713 10999 24715 11051
rect 24715 10999 24767 11051
rect 24767 10999 24769 11051
rect 24713 10997 24769 10999
rect 25079 11051 25135 11053
rect 25079 10999 25081 11051
rect 25081 10999 25133 11051
rect 25133 10999 25135 11051
rect 25079 10997 25135 10999
rect 25159 11051 25215 11053
rect 25159 10999 25161 11051
rect 25161 10999 25213 11051
rect 25213 10999 25215 11051
rect 25159 10997 25215 10999
rect 25239 11051 25295 11053
rect 25239 10999 25241 11051
rect 25241 10999 25293 11051
rect 25293 10999 25295 11051
rect 25239 10997 25295 10999
rect 25319 11051 25375 11053
rect 25319 10999 25321 11051
rect 25321 10999 25373 11051
rect 25373 10999 25375 11051
rect 25319 10997 25375 10999
rect 25813 11051 25869 11053
rect 25813 10999 25815 11051
rect 25815 10999 25867 11051
rect 25867 10999 25869 11051
rect 25813 10997 25869 10999
rect 25893 11051 25949 11053
rect 25893 10999 25895 11051
rect 25895 10999 25947 11051
rect 25947 10999 25949 11051
rect 25893 10997 25949 10999
rect 25973 11051 26029 11053
rect 25973 10999 25975 11051
rect 25975 10999 26027 11051
rect 26027 10999 26029 11051
rect 25973 10997 26029 10999
rect 26053 11051 26109 11053
rect 26053 10999 26055 11051
rect 26055 10999 26107 11051
rect 26107 10999 26109 11051
rect 26053 10997 26109 10999
rect 13779 10110 13835 10112
rect 13779 10058 13781 10110
rect 13781 10058 13833 10110
rect 13833 10058 13835 10110
rect 13779 10056 13835 10058
rect 13859 10110 13915 10112
rect 13859 10058 13861 10110
rect 13861 10058 13913 10110
rect 13913 10058 13915 10110
rect 13859 10056 13915 10058
rect 13939 10110 13995 10112
rect 13939 10058 13941 10110
rect 13941 10058 13993 10110
rect 13993 10058 13995 10110
rect 13939 10056 13995 10058
rect 14019 10110 14075 10112
rect 14019 10058 14021 10110
rect 14021 10058 14073 10110
rect 14073 10058 14075 10110
rect 14019 10056 14075 10058
rect 14513 10110 14569 10112
rect 14513 10058 14515 10110
rect 14515 10058 14567 10110
rect 14567 10058 14569 10110
rect 14513 10056 14569 10058
rect 14593 10110 14649 10112
rect 14593 10058 14595 10110
rect 14595 10058 14647 10110
rect 14647 10058 14649 10110
rect 14593 10056 14649 10058
rect 14673 10110 14729 10112
rect 14673 10058 14675 10110
rect 14675 10058 14727 10110
rect 14727 10058 14729 10110
rect 14673 10056 14729 10058
rect 14753 10110 14809 10112
rect 14753 10058 14755 10110
rect 14755 10058 14807 10110
rect 14807 10058 14809 10110
rect 14753 10056 14809 10058
rect 15119 10110 15175 10112
rect 15119 10058 15121 10110
rect 15121 10058 15173 10110
rect 15173 10058 15175 10110
rect 15119 10056 15175 10058
rect 15199 10110 15255 10112
rect 15199 10058 15201 10110
rect 15201 10058 15253 10110
rect 15253 10058 15255 10110
rect 15199 10056 15255 10058
rect 15279 10110 15335 10112
rect 15279 10058 15281 10110
rect 15281 10058 15333 10110
rect 15333 10058 15335 10110
rect 15279 10056 15335 10058
rect 15359 10110 15415 10112
rect 15359 10058 15361 10110
rect 15361 10058 15413 10110
rect 15413 10058 15415 10110
rect 15359 10056 15415 10058
rect 15851 10110 15907 10112
rect 15851 10058 15853 10110
rect 15853 10058 15905 10110
rect 15905 10058 15907 10110
rect 15851 10056 15907 10058
rect 15931 10110 15987 10112
rect 15931 10058 15933 10110
rect 15933 10058 15985 10110
rect 15985 10058 15987 10110
rect 15931 10056 15987 10058
rect 16011 10110 16067 10112
rect 16011 10058 16013 10110
rect 16013 10058 16065 10110
rect 16065 10058 16067 10110
rect 16011 10056 16067 10058
rect 16091 10110 16147 10112
rect 16091 10058 16093 10110
rect 16093 10058 16145 10110
rect 16145 10058 16147 10110
rect 16091 10056 16147 10058
rect 16457 10110 16513 10112
rect 16457 10058 16459 10110
rect 16459 10058 16511 10110
rect 16511 10058 16513 10110
rect 16457 10056 16513 10058
rect 16537 10110 16593 10112
rect 16537 10058 16539 10110
rect 16539 10058 16591 10110
rect 16591 10058 16593 10110
rect 16537 10056 16593 10058
rect 16617 10110 16673 10112
rect 16617 10058 16619 10110
rect 16619 10058 16671 10110
rect 16671 10058 16673 10110
rect 16617 10056 16673 10058
rect 16697 10110 16753 10112
rect 16697 10058 16699 10110
rect 16699 10058 16751 10110
rect 16751 10058 16753 10110
rect 16697 10056 16753 10058
rect 17063 10110 17119 10112
rect 17063 10058 17065 10110
rect 17065 10058 17117 10110
rect 17117 10058 17119 10110
rect 17063 10056 17119 10058
rect 17143 10110 17199 10112
rect 17143 10058 17145 10110
rect 17145 10058 17197 10110
rect 17197 10058 17199 10110
rect 17143 10056 17199 10058
rect 17223 10110 17279 10112
rect 17223 10058 17225 10110
rect 17225 10058 17277 10110
rect 17277 10058 17279 10110
rect 17223 10056 17279 10058
rect 17303 10110 17359 10112
rect 17303 10058 17305 10110
rect 17305 10058 17357 10110
rect 17357 10058 17359 10110
rect 17303 10056 17359 10058
rect 17669 10110 17725 10112
rect 17669 10058 17671 10110
rect 17671 10058 17723 10110
rect 17723 10058 17725 10110
rect 17669 10056 17725 10058
rect 17749 10110 17805 10112
rect 17749 10058 17751 10110
rect 17751 10058 17803 10110
rect 17803 10058 17805 10110
rect 17749 10056 17805 10058
rect 17829 10110 17885 10112
rect 17829 10058 17831 10110
rect 17831 10058 17883 10110
rect 17883 10058 17885 10110
rect 17829 10056 17885 10058
rect 17909 10110 17965 10112
rect 17909 10058 17911 10110
rect 17911 10058 17963 10110
rect 17963 10058 17965 10110
rect 17909 10056 17965 10058
rect 18401 10110 18457 10112
rect 18401 10058 18403 10110
rect 18403 10058 18455 10110
rect 18455 10058 18457 10110
rect 18401 10056 18457 10058
rect 18481 10110 18537 10112
rect 18481 10058 18483 10110
rect 18483 10058 18535 10110
rect 18535 10058 18537 10110
rect 18481 10056 18537 10058
rect 18561 10110 18617 10112
rect 18561 10058 18563 10110
rect 18563 10058 18615 10110
rect 18615 10058 18617 10110
rect 18561 10056 18617 10058
rect 18641 10110 18697 10112
rect 18641 10058 18643 10110
rect 18643 10058 18695 10110
rect 18695 10058 18697 10110
rect 18641 10056 18697 10058
rect 10496 9156 10552 9158
rect 10496 9104 10498 9156
rect 10498 9104 10550 9156
rect 10550 9104 10552 9156
rect 10496 9102 10552 9104
rect 3548 8682 3612 8746
rect 4280 8679 4344 8743
rect 4508 8679 4572 8743
rect 5492 8679 5556 8743
rect 5720 8679 5784 8743
rect 6704 8679 6768 8743
rect 6932 8679 6996 8743
rect 7916 8679 7980 8743
rect 8144 8679 8208 8743
rect 8886 8735 8942 8737
rect 8886 8683 8888 8735
rect 8888 8683 8940 8735
rect 8940 8683 8942 8735
rect 8886 8681 8942 8683
rect 8798 8474 8854 8476
rect 8798 8422 8800 8474
rect 8800 8422 8852 8474
rect 8852 8422 8854 8474
rect 8798 8420 8854 8422
rect 9208 8448 9264 8450
rect 9208 8396 9210 8448
rect 9210 8396 9262 8448
rect 9262 8396 9264 8448
rect 9208 8394 9264 8396
rect 2449 8152 2505 8154
rect 2449 8100 2451 8152
rect 2451 8100 2503 8152
rect 2503 8100 2505 8152
rect 2449 8098 2505 8100
rect 2580 8153 2636 8155
rect 2580 8101 2582 8153
rect 2582 8101 2634 8153
rect 2634 8101 2636 8153
rect 2580 8099 2636 8101
rect 2724 8152 2780 8154
rect 2724 8100 2726 8152
rect 2726 8100 2778 8152
rect 2778 8100 2780 8152
rect 2724 8098 2780 8100
rect 8880 8232 8936 8234
rect 8880 8180 8882 8232
rect 8882 8180 8934 8232
rect 8934 8180 8936 8232
rect 8880 8178 8936 8180
rect 8881 8075 8937 8077
rect 8881 8023 8883 8075
rect 8883 8023 8935 8075
rect 8935 8023 8937 8075
rect 8881 8021 8937 8023
rect 9470 8449 9526 8451
rect 9470 8397 9472 8449
rect 9472 8397 9524 8449
rect 9524 8397 9526 8449
rect 9470 8395 9526 8397
rect 9742 8449 9798 8451
rect 9742 8397 9744 8449
rect 9744 8397 9796 8449
rect 9796 8397 9798 8449
rect 9742 8395 9798 8397
rect 10069 8449 10125 8451
rect 10069 8397 10071 8449
rect 10071 8397 10123 8449
rect 10123 8397 10125 8449
rect 10069 8395 10125 8397
rect 10450 8449 10506 8451
rect 10450 8397 10452 8449
rect 10452 8397 10504 8449
rect 10504 8397 10506 8449
rect 10450 8395 10506 8397
rect 10844 9156 10900 9158
rect 10844 9104 10846 9156
rect 10846 9104 10898 9156
rect 10898 9104 10900 9156
rect 10844 9102 10900 9104
rect 11102 9162 11158 9164
rect 11102 9110 11104 9162
rect 11104 9110 11156 9162
rect 11156 9110 11158 9162
rect 11102 9108 11158 9110
rect 11328 9162 11384 9164
rect 11328 9110 11330 9162
rect 11330 9110 11382 9162
rect 11382 9110 11384 9162
rect 11328 9108 11384 9110
rect 11587 9165 11643 9167
rect 11587 9113 11589 9165
rect 11589 9113 11641 9165
rect 11641 9113 11643 9165
rect 11587 9111 11643 9113
rect 12194 9127 12250 9129
rect 12194 9075 12196 9127
rect 12196 9075 12248 9127
rect 12248 9075 12250 9127
rect 12194 9073 12250 9075
rect 12426 9128 12482 9130
rect 12426 9076 12428 9128
rect 12428 9076 12480 9128
rect 12480 9076 12482 9128
rect 12426 9074 12482 9076
rect 12862 9134 12918 9136
rect 12862 9082 12864 9134
rect 12864 9082 12916 9134
rect 12916 9082 12918 9134
rect 12862 9080 12918 9082
rect 13097 9136 13153 9138
rect 13097 9084 13099 9136
rect 13099 9084 13151 9136
rect 13151 9084 13153 9136
rect 13097 9082 13153 9084
rect 13440 9188 13496 9190
rect 13440 9136 13442 9188
rect 13442 9136 13494 9188
rect 13494 9136 13496 9188
rect 13440 9134 13496 9136
rect 19183 10113 19239 10115
rect 19183 10061 19185 10113
rect 19185 10061 19237 10113
rect 19237 10061 19239 10113
rect 19183 10059 19239 10061
rect 20488 10110 20544 10112
rect 20488 10058 20490 10110
rect 20490 10058 20542 10110
rect 20542 10058 20544 10110
rect 20488 10056 20544 10058
rect 20568 10110 20624 10112
rect 20568 10058 20570 10110
rect 20570 10058 20622 10110
rect 20622 10058 20624 10110
rect 20568 10056 20624 10058
rect 20648 10110 20704 10112
rect 20648 10058 20650 10110
rect 20650 10058 20702 10110
rect 20702 10058 20704 10110
rect 20648 10056 20704 10058
rect 20728 10110 20784 10112
rect 20728 10058 20730 10110
rect 20730 10058 20782 10110
rect 20782 10058 20784 10110
rect 20728 10056 20784 10058
rect 21222 10110 21278 10112
rect 21222 10058 21224 10110
rect 21224 10058 21276 10110
rect 21276 10058 21278 10110
rect 21222 10056 21278 10058
rect 21302 10110 21358 10112
rect 21302 10058 21304 10110
rect 21304 10058 21356 10110
rect 21356 10058 21358 10110
rect 21302 10056 21358 10058
rect 21382 10110 21438 10112
rect 21382 10058 21384 10110
rect 21384 10058 21436 10110
rect 21436 10058 21438 10110
rect 21382 10056 21438 10058
rect 21462 10110 21518 10112
rect 21462 10058 21464 10110
rect 21464 10058 21516 10110
rect 21516 10058 21518 10110
rect 21462 10056 21518 10058
rect 21828 10110 21884 10112
rect 21828 10058 21830 10110
rect 21830 10058 21882 10110
rect 21882 10058 21884 10110
rect 21828 10056 21884 10058
rect 21908 10110 21964 10112
rect 21908 10058 21910 10110
rect 21910 10058 21962 10110
rect 21962 10058 21964 10110
rect 21908 10056 21964 10058
rect 21988 10110 22044 10112
rect 21988 10058 21990 10110
rect 21990 10058 22042 10110
rect 22042 10058 22044 10110
rect 21988 10056 22044 10058
rect 22068 10110 22124 10112
rect 22068 10058 22070 10110
rect 22070 10058 22122 10110
rect 22122 10058 22124 10110
rect 22068 10056 22124 10058
rect 22560 10110 22616 10112
rect 22560 10058 22562 10110
rect 22562 10058 22614 10110
rect 22614 10058 22616 10110
rect 22560 10056 22616 10058
rect 22640 10110 22696 10112
rect 22640 10058 22642 10110
rect 22642 10058 22694 10110
rect 22694 10058 22696 10110
rect 22640 10056 22696 10058
rect 22720 10110 22776 10112
rect 22720 10058 22722 10110
rect 22722 10058 22774 10110
rect 22774 10058 22776 10110
rect 22720 10056 22776 10058
rect 22800 10110 22856 10112
rect 22800 10058 22802 10110
rect 22802 10058 22854 10110
rect 22854 10058 22856 10110
rect 22800 10056 22856 10058
rect 23166 10110 23222 10112
rect 23166 10058 23168 10110
rect 23168 10058 23220 10110
rect 23220 10058 23222 10110
rect 23166 10056 23222 10058
rect 23246 10110 23302 10112
rect 23246 10058 23248 10110
rect 23248 10058 23300 10110
rect 23300 10058 23302 10110
rect 23246 10056 23302 10058
rect 23326 10110 23382 10112
rect 23326 10058 23328 10110
rect 23328 10058 23380 10110
rect 23380 10058 23382 10110
rect 23326 10056 23382 10058
rect 23406 10110 23462 10112
rect 23406 10058 23408 10110
rect 23408 10058 23460 10110
rect 23460 10058 23462 10110
rect 23406 10056 23462 10058
rect 23772 10110 23828 10112
rect 23772 10058 23774 10110
rect 23774 10058 23826 10110
rect 23826 10058 23828 10110
rect 23772 10056 23828 10058
rect 23852 10110 23908 10112
rect 23852 10058 23854 10110
rect 23854 10058 23906 10110
rect 23906 10058 23908 10110
rect 23852 10056 23908 10058
rect 23932 10110 23988 10112
rect 23932 10058 23934 10110
rect 23934 10058 23986 10110
rect 23986 10058 23988 10110
rect 23932 10056 23988 10058
rect 24012 10110 24068 10112
rect 24012 10058 24014 10110
rect 24014 10058 24066 10110
rect 24066 10058 24068 10110
rect 24012 10056 24068 10058
rect 24378 10110 24434 10112
rect 24378 10058 24380 10110
rect 24380 10058 24432 10110
rect 24432 10058 24434 10110
rect 24378 10056 24434 10058
rect 24458 10110 24514 10112
rect 24458 10058 24460 10110
rect 24460 10058 24512 10110
rect 24512 10058 24514 10110
rect 24458 10056 24514 10058
rect 24538 10110 24594 10112
rect 24538 10058 24540 10110
rect 24540 10058 24592 10110
rect 24592 10058 24594 10110
rect 24538 10056 24594 10058
rect 24618 10110 24674 10112
rect 24618 10058 24620 10110
rect 24620 10058 24672 10110
rect 24672 10058 24674 10110
rect 24618 10056 24674 10058
rect 25110 10110 25166 10112
rect 25110 10058 25112 10110
rect 25112 10058 25164 10110
rect 25164 10058 25166 10110
rect 25110 10056 25166 10058
rect 25190 10110 25246 10112
rect 25190 10058 25192 10110
rect 25192 10058 25244 10110
rect 25244 10058 25246 10110
rect 25190 10056 25246 10058
rect 25270 10110 25326 10112
rect 25270 10058 25272 10110
rect 25272 10058 25324 10110
rect 25324 10058 25326 10110
rect 25270 10056 25326 10058
rect 25350 10110 25406 10112
rect 25350 10058 25352 10110
rect 25352 10058 25404 10110
rect 25404 10058 25406 10110
rect 25350 10056 25406 10058
rect 20149 9188 20205 9190
rect 20149 9136 20151 9188
rect 20151 9136 20203 9188
rect 20203 9136 20205 9188
rect 20149 9134 20205 9136
rect 25892 10113 25948 10115
rect 25892 10061 25894 10113
rect 25894 10061 25946 10113
rect 25946 10061 25948 10113
rect 25892 10059 25948 10061
rect 13349 8926 13405 8928
rect 13349 8874 13351 8926
rect 13351 8874 13403 8926
rect 13403 8874 13405 8926
rect 13349 8872 13405 8874
rect 14089 8869 14153 8933
rect 14823 8869 14887 8933
rect 15041 8869 15105 8933
rect 16161 8869 16225 8933
rect 16379 8869 16443 8933
rect 17373 8869 17437 8933
rect 17591 8869 17655 8933
rect 18323 8869 18387 8933
rect 10827 8449 10883 8451
rect 10827 8397 10829 8449
rect 10829 8397 10881 8449
rect 10881 8397 10883 8449
rect 10827 8395 10883 8397
rect 13349 8723 13405 8725
rect 13349 8671 13351 8723
rect 13351 8671 13403 8723
rect 13403 8671 13405 8723
rect 13349 8669 13405 8671
rect 14083 8667 14147 8731
rect 14311 8667 14375 8731
rect 15295 8667 15359 8731
rect 15523 8667 15587 8731
rect 16507 8667 16571 8731
rect 16735 8667 16799 8731
rect 17719 8667 17783 8731
rect 17947 8667 18011 8731
rect 18679 8670 18743 8734
rect 12722 8509 12778 8510
rect 12722 8456 12723 8509
rect 12723 8456 12776 8509
rect 12776 8456 12778 8509
rect 12722 8454 12778 8456
rect 12227 8439 12283 8440
rect 12227 8386 12228 8439
rect 12228 8386 12281 8439
rect 12281 8386 12283 8439
rect 12227 8384 12283 8386
rect 12584 8366 12640 8367
rect 12584 8313 12585 8366
rect 12585 8313 12638 8366
rect 12638 8313 12640 8366
rect 12584 8311 12640 8313
rect 12768 8363 12824 8364
rect 12768 8310 12769 8363
rect 12769 8310 12822 8363
rect 12822 8310 12824 8363
rect 12768 8308 12824 8310
rect 8881 7905 8937 7907
rect 8881 7853 8883 7905
rect 8883 7853 8935 7905
rect 8935 7853 8937 7905
rect 8881 7851 8937 7853
rect 8880 7753 8936 7755
rect 8880 7701 8882 7753
rect 8882 7701 8934 7753
rect 8934 7701 8936 7753
rect 8880 7699 8936 7701
rect 10144 7723 10200 7725
rect 10144 7671 10146 7723
rect 10146 7671 10198 7723
rect 10198 7671 10200 7723
rect 10144 7669 10200 7671
rect 10392 7723 10448 7725
rect 10392 7671 10394 7723
rect 10394 7671 10446 7723
rect 10446 7671 10448 7723
rect 10392 7669 10448 7671
rect 3162 7556 3218 7558
rect 3066 7547 3122 7549
rect 3066 7495 3068 7547
rect 3068 7495 3120 7547
rect 3120 7495 3122 7547
rect 3162 7504 3166 7556
rect 3166 7504 3218 7556
rect 3162 7502 3218 7504
rect 3242 7556 3298 7558
rect 3242 7504 3246 7556
rect 3246 7504 3298 7556
rect 3242 7502 3298 7504
rect 3322 7556 3378 7558
rect 3322 7504 3326 7556
rect 3326 7504 3378 7556
rect 3322 7502 3378 7504
rect 3402 7556 3458 7558
rect 3402 7504 3406 7556
rect 3406 7504 3458 7556
rect 3402 7502 3458 7504
rect 3482 7556 3538 7558
rect 3482 7504 3486 7556
rect 3486 7504 3538 7556
rect 3482 7502 3538 7504
rect 3562 7556 3618 7558
rect 3562 7504 3566 7556
rect 3566 7504 3618 7556
rect 3562 7502 3618 7504
rect 3894 7553 3950 7555
rect 3894 7501 3898 7553
rect 3898 7501 3950 7553
rect 3894 7499 3950 7501
rect 3974 7553 4030 7555
rect 3974 7501 3978 7553
rect 3978 7501 4030 7553
rect 3974 7499 4030 7501
rect 4054 7553 4110 7555
rect 4054 7501 4058 7553
rect 4058 7501 4110 7553
rect 4054 7499 4110 7501
rect 4134 7553 4190 7555
rect 4134 7501 4138 7553
rect 4138 7501 4190 7553
rect 4134 7499 4190 7501
rect 4214 7553 4270 7555
rect 4214 7501 4218 7553
rect 4218 7501 4270 7553
rect 4214 7499 4270 7501
rect 4294 7553 4350 7555
rect 4294 7501 4298 7553
rect 4298 7501 4350 7553
rect 4294 7499 4350 7501
rect 4502 7553 4558 7555
rect 4502 7501 4554 7553
rect 4554 7501 4558 7553
rect 4502 7499 4558 7501
rect 4582 7553 4638 7555
rect 4582 7501 4634 7553
rect 4634 7501 4638 7553
rect 4582 7499 4638 7501
rect 4662 7553 4718 7555
rect 4662 7501 4714 7553
rect 4714 7501 4718 7553
rect 4662 7499 4718 7501
rect 4742 7553 4798 7555
rect 4742 7501 4794 7553
rect 4794 7501 4798 7553
rect 4742 7499 4798 7501
rect 4822 7553 4878 7555
rect 4822 7501 4874 7553
rect 4874 7501 4878 7553
rect 4822 7499 4878 7501
rect 4902 7553 4958 7555
rect 4902 7501 4954 7553
rect 4954 7501 4958 7553
rect 4902 7499 4958 7501
rect 5106 7553 5162 7555
rect 5106 7501 5110 7553
rect 5110 7501 5162 7553
rect 5106 7499 5162 7501
rect 5186 7553 5242 7555
rect 5186 7501 5190 7553
rect 5190 7501 5242 7553
rect 5186 7499 5242 7501
rect 5266 7553 5322 7555
rect 5266 7501 5270 7553
rect 5270 7501 5322 7553
rect 5266 7499 5322 7501
rect 5346 7553 5402 7555
rect 5346 7501 5350 7553
rect 5350 7501 5402 7553
rect 5346 7499 5402 7501
rect 5426 7553 5482 7555
rect 5426 7501 5430 7553
rect 5430 7501 5482 7553
rect 5426 7499 5482 7501
rect 5506 7553 5562 7555
rect 5506 7501 5510 7553
rect 5510 7501 5562 7553
rect 5506 7499 5562 7501
rect 5714 7553 5770 7555
rect 5714 7501 5766 7553
rect 5766 7501 5770 7553
rect 5714 7499 5770 7501
rect 5794 7553 5850 7555
rect 5794 7501 5846 7553
rect 5846 7501 5850 7553
rect 5794 7499 5850 7501
rect 5874 7553 5930 7555
rect 5874 7501 5926 7553
rect 5926 7501 5930 7553
rect 5874 7499 5930 7501
rect 5954 7553 6010 7555
rect 5954 7501 6006 7553
rect 6006 7501 6010 7553
rect 5954 7499 6010 7501
rect 6034 7553 6090 7555
rect 6034 7501 6086 7553
rect 6086 7501 6090 7553
rect 6034 7499 6090 7501
rect 6114 7553 6170 7555
rect 6114 7501 6166 7553
rect 6166 7501 6170 7553
rect 6114 7499 6170 7501
rect 6318 7553 6374 7555
rect 6318 7501 6322 7553
rect 6322 7501 6374 7553
rect 6318 7499 6374 7501
rect 6398 7553 6454 7555
rect 6398 7501 6402 7553
rect 6402 7501 6454 7553
rect 6398 7499 6454 7501
rect 6478 7553 6534 7555
rect 6478 7501 6482 7553
rect 6482 7501 6534 7553
rect 6478 7499 6534 7501
rect 6558 7553 6614 7555
rect 6558 7501 6562 7553
rect 6562 7501 6614 7553
rect 6558 7499 6614 7501
rect 6638 7553 6694 7555
rect 6638 7501 6642 7553
rect 6642 7501 6694 7553
rect 6638 7499 6694 7501
rect 6718 7553 6774 7555
rect 6718 7501 6722 7553
rect 6722 7501 6774 7553
rect 6718 7499 6774 7501
rect 6926 7553 6982 7555
rect 6926 7501 6978 7553
rect 6978 7501 6982 7553
rect 6926 7499 6982 7501
rect 7006 7553 7062 7555
rect 7006 7501 7058 7553
rect 7058 7501 7062 7553
rect 7006 7499 7062 7501
rect 7086 7553 7142 7555
rect 7086 7501 7138 7553
rect 7138 7501 7142 7553
rect 7086 7499 7142 7501
rect 7166 7553 7222 7555
rect 7166 7501 7218 7553
rect 7218 7501 7222 7553
rect 7166 7499 7222 7501
rect 7246 7553 7302 7555
rect 7246 7501 7298 7553
rect 7298 7501 7302 7553
rect 7246 7499 7302 7501
rect 7326 7553 7382 7555
rect 7326 7501 7378 7553
rect 7378 7501 7382 7553
rect 7326 7499 7382 7501
rect 7530 7553 7586 7555
rect 7530 7501 7534 7553
rect 7534 7501 7586 7553
rect 7530 7499 7586 7501
rect 7610 7553 7666 7555
rect 7610 7501 7614 7553
rect 7614 7501 7666 7553
rect 7610 7499 7666 7501
rect 7690 7553 7746 7555
rect 7690 7501 7694 7553
rect 7694 7501 7746 7553
rect 7690 7499 7746 7501
rect 7770 7553 7826 7555
rect 7770 7501 7774 7553
rect 7774 7501 7826 7553
rect 7770 7499 7826 7501
rect 7850 7553 7906 7555
rect 7850 7501 7854 7553
rect 7854 7501 7906 7553
rect 7850 7499 7906 7501
rect 7930 7553 7986 7555
rect 7930 7501 7934 7553
rect 7934 7501 7986 7553
rect 7930 7499 7986 7501
rect 8138 7553 8194 7555
rect 8138 7501 8190 7553
rect 8190 7501 8194 7553
rect 8138 7499 8194 7501
rect 8218 7553 8274 7555
rect 8218 7501 8270 7553
rect 8270 7501 8274 7553
rect 8218 7499 8274 7501
rect 8298 7553 8354 7555
rect 8298 7501 8350 7553
rect 8350 7501 8354 7553
rect 8298 7499 8354 7501
rect 8378 7553 8434 7555
rect 8378 7501 8430 7553
rect 8430 7501 8434 7553
rect 8378 7499 8434 7501
rect 8458 7553 8514 7555
rect 8458 7501 8510 7553
rect 8510 7501 8514 7553
rect 8458 7499 8514 7501
rect 8538 7553 8594 7555
rect 8538 7501 8590 7553
rect 8590 7501 8594 7553
rect 8538 7499 8594 7501
rect 8875 7609 8931 7611
rect 8875 7557 8877 7609
rect 8877 7557 8929 7609
rect 8929 7557 8931 7609
rect 8875 7555 8931 7557
rect 3066 7493 3122 7495
rect 10689 7723 10745 7725
rect 10689 7671 10691 7723
rect 10691 7671 10743 7723
rect 10743 7671 10745 7723
rect 10689 7669 10745 7671
rect 11033 7725 11089 7727
rect 11033 7673 11035 7725
rect 11035 7673 11087 7725
rect 11087 7673 11089 7725
rect 11033 7671 11089 7673
rect 11352 7725 11408 7727
rect 11352 7673 11354 7725
rect 11354 7673 11406 7725
rect 11406 7673 11408 7725
rect 11352 7671 11408 7673
rect 20058 8926 20114 8928
rect 20058 8874 20060 8926
rect 20060 8874 20112 8926
rect 20112 8874 20114 8926
rect 20058 8872 20114 8874
rect 20798 8869 20862 8933
rect 21532 8869 21596 8933
rect 21750 8869 21814 8933
rect 22870 8869 22934 8933
rect 23088 8869 23152 8933
rect 24082 8869 24146 8933
rect 24300 8869 24364 8933
rect 25032 8869 25096 8933
rect 19505 8686 19561 8688
rect 19505 8634 19507 8686
rect 19507 8634 19559 8686
rect 19559 8634 19561 8686
rect 19505 8632 19561 8634
rect 19648 8686 19704 8688
rect 19648 8634 19650 8686
rect 19650 8634 19702 8686
rect 19702 8634 19704 8686
rect 19648 8632 19704 8634
rect 19768 8686 19824 8688
rect 19768 8634 19770 8686
rect 19770 8634 19822 8686
rect 19822 8634 19824 8686
rect 20058 8723 20114 8725
rect 20058 8671 20060 8723
rect 20060 8671 20112 8723
rect 20112 8671 20114 8723
rect 20058 8669 20114 8671
rect 20792 8667 20856 8731
rect 21020 8667 21084 8731
rect 22004 8667 22068 8731
rect 22232 8667 22296 8731
rect 23216 8667 23280 8731
rect 23444 8667 23508 8731
rect 24428 8667 24492 8731
rect 24656 8667 24720 8731
rect 25388 8670 25452 8734
rect 19768 8632 19824 8634
rect 26214 8686 26270 8688
rect 26214 8634 26216 8686
rect 26216 8634 26268 8686
rect 26268 8634 26270 8686
rect 26214 8632 26270 8634
rect 26357 8686 26413 8688
rect 26357 8634 26359 8686
rect 26359 8634 26411 8686
rect 26411 8634 26413 8686
rect 26357 8632 26413 8634
rect 26477 8686 26533 8688
rect 26477 8634 26479 8686
rect 26479 8634 26531 8686
rect 26531 8634 26533 8686
rect 26477 8632 26533 8634
rect 13096 8509 13152 8510
rect 13096 8456 13097 8509
rect 13097 8456 13150 8509
rect 13150 8456 13152 8509
rect 13096 8454 13152 8456
rect 13437 8462 13493 8464
rect 13437 8410 13439 8462
rect 13439 8410 13491 8462
rect 13491 8410 13493 8462
rect 13437 8408 13493 8410
rect 20146 8462 20202 8464
rect 20146 8410 20148 8462
rect 20148 8410 20200 8462
rect 20200 8410 20202 8462
rect 20146 8408 20202 8410
rect 13070 8357 13126 8358
rect 13070 8304 13071 8357
rect 13071 8304 13124 8357
rect 13124 8304 13126 8357
rect 13070 8302 13126 8304
rect 13355 8220 13411 8222
rect 13355 8168 13357 8220
rect 13357 8168 13409 8220
rect 13409 8168 13411 8220
rect 13355 8166 13411 8168
rect 20064 8220 20120 8222
rect 20064 8168 20066 8220
rect 20066 8168 20118 8220
rect 20118 8168 20120 8220
rect 20064 8166 20120 8168
rect 19511 8140 19567 8142
rect 19511 8088 19513 8140
rect 19513 8088 19565 8140
rect 19565 8088 19567 8140
rect 19511 8086 19567 8088
rect 19655 8141 19711 8143
rect 19655 8089 19657 8141
rect 19657 8089 19709 8141
rect 19709 8089 19711 8141
rect 19655 8087 19711 8089
rect 19786 8140 19842 8142
rect 19786 8088 19788 8140
rect 19788 8088 19840 8140
rect 19840 8088 19842 8140
rect 19786 8086 19842 8088
rect 26220 8140 26276 8142
rect 26220 8088 26222 8140
rect 26222 8088 26274 8140
rect 26274 8088 26276 8140
rect 26220 8086 26276 8088
rect 26364 8141 26420 8143
rect 26364 8089 26366 8141
rect 26366 8089 26418 8141
rect 26418 8089 26420 8141
rect 26364 8087 26420 8089
rect 26495 8140 26551 8142
rect 26495 8088 26497 8140
rect 26497 8088 26549 8140
rect 26549 8088 26551 8140
rect 26495 8086 26551 8088
rect 13354 8063 13410 8065
rect 13354 8011 13356 8063
rect 13356 8011 13408 8063
rect 13408 8011 13410 8063
rect 13354 8009 13410 8011
rect 20063 8063 20119 8065
rect 20063 8011 20065 8063
rect 20065 8011 20117 8063
rect 20117 8011 20119 8063
rect 20063 8009 20119 8011
rect 19641 7991 19697 7993
rect 19641 7939 19643 7991
rect 19643 7939 19695 7991
rect 19695 7939 19697 7991
rect 19641 7937 19697 7939
rect 12938 7929 12994 7931
rect 12938 7877 12940 7929
rect 12940 7877 12992 7929
rect 12992 7877 12994 7929
rect 12938 7875 12994 7877
rect 13354 7893 13410 7895
rect 13354 7841 13356 7893
rect 13356 7841 13408 7893
rect 13408 7841 13410 7893
rect 13354 7839 13410 7841
rect 20063 7893 20119 7895
rect 20063 7841 20065 7893
rect 20065 7841 20117 7893
rect 20117 7841 20119 7893
rect 20063 7839 20119 7841
rect 11964 7734 12020 7736
rect 11964 7682 11966 7734
rect 11966 7682 12018 7734
rect 12018 7682 12020 7734
rect 11964 7680 12020 7682
rect 12218 7738 12274 7740
rect 12218 7686 12220 7738
rect 12220 7686 12272 7738
rect 12272 7686 12274 7738
rect 12218 7684 12274 7686
rect 12930 7709 12986 7711
rect 12930 7657 12932 7709
rect 12932 7657 12984 7709
rect 12984 7657 12986 7709
rect 12930 7655 12986 7657
rect 13355 7741 13411 7743
rect 13355 7689 13357 7741
rect 13357 7689 13409 7741
rect 13409 7689 13411 7741
rect 13355 7687 13411 7689
rect 19641 7795 19697 7797
rect 19641 7743 19643 7795
rect 19643 7743 19695 7795
rect 19695 7743 19697 7795
rect 19641 7741 19697 7743
rect 20064 7741 20120 7743
rect 20064 7689 20066 7741
rect 20066 7689 20118 7741
rect 20118 7689 20120 7741
rect 20064 7687 20120 7689
rect 11974 7589 12030 7591
rect 11974 7537 11976 7589
rect 11976 7537 12028 7589
rect 12028 7537 12030 7589
rect 11974 7535 12030 7537
rect 12226 7592 12282 7594
rect 12226 7540 12228 7592
rect 12228 7540 12280 7592
rect 12280 7540 12282 7592
rect 12226 7538 12282 7540
rect 13360 7597 13416 7599
rect 13360 7545 13362 7597
rect 13362 7545 13414 7597
rect 13414 7545 13416 7597
rect 13360 7543 13416 7545
rect 19641 7620 19697 7622
rect 19641 7568 19643 7620
rect 19643 7568 19695 7620
rect 19695 7568 19697 7620
rect 19641 7566 19697 7568
rect 13697 7541 13753 7543
rect 13697 7489 13701 7541
rect 13701 7489 13753 7541
rect 13697 7487 13753 7489
rect 13777 7541 13833 7543
rect 13777 7489 13781 7541
rect 13781 7489 13833 7541
rect 13777 7487 13833 7489
rect 13857 7541 13913 7543
rect 13857 7489 13861 7541
rect 13861 7489 13913 7541
rect 13857 7487 13913 7489
rect 13937 7541 13993 7543
rect 13937 7489 13941 7541
rect 13941 7489 13993 7541
rect 13937 7487 13993 7489
rect 14017 7541 14073 7543
rect 14017 7489 14021 7541
rect 14021 7489 14073 7541
rect 14017 7487 14073 7489
rect 14097 7541 14153 7543
rect 14097 7489 14101 7541
rect 14101 7489 14153 7541
rect 14097 7487 14153 7489
rect 14305 7541 14361 7543
rect 14305 7489 14357 7541
rect 14357 7489 14361 7541
rect 14305 7487 14361 7489
rect 14385 7541 14441 7543
rect 14385 7489 14437 7541
rect 14437 7489 14441 7541
rect 14385 7487 14441 7489
rect 14465 7541 14521 7543
rect 14465 7489 14517 7541
rect 14517 7489 14521 7541
rect 14465 7487 14521 7489
rect 14545 7541 14601 7543
rect 14545 7489 14597 7541
rect 14597 7489 14601 7541
rect 14545 7487 14601 7489
rect 14625 7541 14681 7543
rect 14625 7489 14677 7541
rect 14677 7489 14681 7541
rect 14625 7487 14681 7489
rect 14705 7541 14761 7543
rect 14705 7489 14757 7541
rect 14757 7489 14761 7541
rect 14705 7487 14761 7489
rect 14909 7541 14965 7543
rect 14909 7489 14913 7541
rect 14913 7489 14965 7541
rect 14909 7487 14965 7489
rect 14989 7541 15045 7543
rect 14989 7489 14993 7541
rect 14993 7489 15045 7541
rect 14989 7487 15045 7489
rect 15069 7541 15125 7543
rect 15069 7489 15073 7541
rect 15073 7489 15125 7541
rect 15069 7487 15125 7489
rect 15149 7541 15205 7543
rect 15149 7489 15153 7541
rect 15153 7489 15205 7541
rect 15149 7487 15205 7489
rect 15229 7541 15285 7543
rect 15229 7489 15233 7541
rect 15233 7489 15285 7541
rect 15229 7487 15285 7489
rect 15309 7541 15365 7543
rect 15309 7489 15313 7541
rect 15313 7489 15365 7541
rect 15309 7487 15365 7489
rect 15517 7541 15573 7543
rect 15517 7489 15569 7541
rect 15569 7489 15573 7541
rect 15517 7487 15573 7489
rect 15597 7541 15653 7543
rect 15597 7489 15649 7541
rect 15649 7489 15653 7541
rect 15597 7487 15653 7489
rect 15677 7541 15733 7543
rect 15677 7489 15729 7541
rect 15729 7489 15733 7541
rect 15677 7487 15733 7489
rect 15757 7541 15813 7543
rect 15757 7489 15809 7541
rect 15809 7489 15813 7541
rect 15757 7487 15813 7489
rect 15837 7541 15893 7543
rect 15837 7489 15889 7541
rect 15889 7489 15893 7541
rect 15837 7487 15893 7489
rect 15917 7541 15973 7543
rect 15917 7489 15969 7541
rect 15969 7489 15973 7541
rect 15917 7487 15973 7489
rect 16121 7541 16177 7543
rect 16121 7489 16125 7541
rect 16125 7489 16177 7541
rect 16121 7487 16177 7489
rect 16201 7541 16257 7543
rect 16201 7489 16205 7541
rect 16205 7489 16257 7541
rect 16201 7487 16257 7489
rect 16281 7541 16337 7543
rect 16281 7489 16285 7541
rect 16285 7489 16337 7541
rect 16281 7487 16337 7489
rect 16361 7541 16417 7543
rect 16361 7489 16365 7541
rect 16365 7489 16417 7541
rect 16361 7487 16417 7489
rect 16441 7541 16497 7543
rect 16441 7489 16445 7541
rect 16445 7489 16497 7541
rect 16441 7487 16497 7489
rect 16521 7541 16577 7543
rect 16521 7489 16525 7541
rect 16525 7489 16577 7541
rect 16521 7487 16577 7489
rect 16729 7541 16785 7543
rect 16729 7489 16781 7541
rect 16781 7489 16785 7541
rect 16729 7487 16785 7489
rect 16809 7541 16865 7543
rect 16809 7489 16861 7541
rect 16861 7489 16865 7541
rect 16809 7487 16865 7489
rect 16889 7541 16945 7543
rect 16889 7489 16941 7541
rect 16941 7489 16945 7541
rect 16889 7487 16945 7489
rect 16969 7541 17025 7543
rect 16969 7489 17021 7541
rect 17021 7489 17025 7541
rect 16969 7487 17025 7489
rect 17049 7541 17105 7543
rect 17049 7489 17101 7541
rect 17101 7489 17105 7541
rect 17049 7487 17105 7489
rect 17129 7541 17185 7543
rect 17129 7489 17181 7541
rect 17181 7489 17185 7541
rect 17129 7487 17185 7489
rect 17333 7541 17389 7543
rect 17333 7489 17337 7541
rect 17337 7489 17389 7541
rect 17333 7487 17389 7489
rect 17413 7541 17469 7543
rect 17413 7489 17417 7541
rect 17417 7489 17469 7541
rect 17413 7487 17469 7489
rect 17493 7541 17549 7543
rect 17493 7489 17497 7541
rect 17497 7489 17549 7541
rect 17493 7487 17549 7489
rect 17573 7541 17629 7543
rect 17573 7489 17577 7541
rect 17577 7489 17629 7541
rect 17573 7487 17629 7489
rect 17653 7541 17709 7543
rect 17653 7489 17657 7541
rect 17657 7489 17709 7541
rect 17653 7487 17709 7489
rect 17733 7541 17789 7543
rect 17733 7489 17737 7541
rect 17737 7489 17789 7541
rect 17733 7487 17789 7489
rect 17941 7541 17997 7543
rect 17941 7489 17993 7541
rect 17993 7489 17997 7541
rect 17941 7487 17997 7489
rect 18021 7541 18077 7543
rect 18021 7489 18073 7541
rect 18073 7489 18077 7541
rect 18021 7487 18077 7489
rect 18101 7541 18157 7543
rect 18101 7489 18153 7541
rect 18153 7489 18157 7541
rect 18101 7487 18157 7489
rect 18181 7541 18237 7543
rect 18181 7489 18233 7541
rect 18233 7489 18237 7541
rect 18181 7487 18237 7489
rect 18261 7541 18317 7543
rect 18261 7489 18313 7541
rect 18313 7489 18317 7541
rect 18261 7487 18317 7489
rect 18341 7541 18397 7543
rect 18341 7489 18393 7541
rect 18393 7489 18397 7541
rect 18341 7487 18397 7489
rect 18673 7544 18729 7546
rect 18673 7492 18725 7544
rect 18725 7492 18729 7544
rect 18673 7490 18729 7492
rect 18753 7544 18809 7546
rect 18753 7492 18805 7544
rect 18805 7492 18809 7544
rect 18753 7490 18809 7492
rect 18833 7544 18889 7546
rect 18833 7492 18885 7544
rect 18885 7492 18889 7544
rect 18833 7490 18889 7492
rect 18913 7544 18969 7546
rect 18913 7492 18965 7544
rect 18965 7492 18969 7544
rect 18913 7490 18969 7492
rect 18993 7544 19049 7546
rect 18993 7492 19045 7544
rect 19045 7492 19049 7544
rect 18993 7490 19049 7492
rect 19073 7544 19129 7546
rect 19073 7492 19125 7544
rect 19125 7492 19129 7544
rect 20069 7597 20125 7599
rect 20069 7545 20071 7597
rect 20071 7545 20123 7597
rect 20123 7545 20125 7597
rect 20069 7543 20125 7545
rect 19073 7490 19129 7492
rect 19169 7535 19225 7537
rect 19169 7483 19171 7535
rect 19171 7483 19223 7535
rect 19223 7483 19225 7535
rect 19169 7481 19225 7483
rect 20406 7541 20462 7543
rect 20406 7489 20410 7541
rect 20410 7489 20462 7541
rect 20406 7487 20462 7489
rect 20486 7541 20542 7543
rect 20486 7489 20490 7541
rect 20490 7489 20542 7541
rect 20486 7487 20542 7489
rect 20566 7541 20622 7543
rect 20566 7489 20570 7541
rect 20570 7489 20622 7541
rect 20566 7487 20622 7489
rect 20646 7541 20702 7543
rect 20646 7489 20650 7541
rect 20650 7489 20702 7541
rect 20646 7487 20702 7489
rect 20726 7541 20782 7543
rect 20726 7489 20730 7541
rect 20730 7489 20782 7541
rect 20726 7487 20782 7489
rect 20806 7541 20862 7543
rect 20806 7489 20810 7541
rect 20810 7489 20862 7541
rect 20806 7487 20862 7489
rect 21014 7541 21070 7543
rect 21014 7489 21066 7541
rect 21066 7489 21070 7541
rect 21014 7487 21070 7489
rect 21094 7541 21150 7543
rect 21094 7489 21146 7541
rect 21146 7489 21150 7541
rect 21094 7487 21150 7489
rect 21174 7541 21230 7543
rect 21174 7489 21226 7541
rect 21226 7489 21230 7541
rect 21174 7487 21230 7489
rect 21254 7541 21310 7543
rect 21254 7489 21306 7541
rect 21306 7489 21310 7541
rect 21254 7487 21310 7489
rect 21334 7541 21390 7543
rect 21334 7489 21386 7541
rect 21386 7489 21390 7541
rect 21334 7487 21390 7489
rect 21414 7541 21470 7543
rect 21414 7489 21466 7541
rect 21466 7489 21470 7541
rect 21414 7487 21470 7489
rect 21618 7541 21674 7543
rect 21618 7489 21622 7541
rect 21622 7489 21674 7541
rect 21618 7487 21674 7489
rect 21698 7541 21754 7543
rect 21698 7489 21702 7541
rect 21702 7489 21754 7541
rect 21698 7487 21754 7489
rect 21778 7541 21834 7543
rect 21778 7489 21782 7541
rect 21782 7489 21834 7541
rect 21778 7487 21834 7489
rect 21858 7541 21914 7543
rect 21858 7489 21862 7541
rect 21862 7489 21914 7541
rect 21858 7487 21914 7489
rect 21938 7541 21994 7543
rect 21938 7489 21942 7541
rect 21942 7489 21994 7541
rect 21938 7487 21994 7489
rect 22018 7541 22074 7543
rect 22018 7489 22022 7541
rect 22022 7489 22074 7541
rect 22018 7487 22074 7489
rect 22226 7541 22282 7543
rect 22226 7489 22278 7541
rect 22278 7489 22282 7541
rect 22226 7487 22282 7489
rect 22306 7541 22362 7543
rect 22306 7489 22358 7541
rect 22358 7489 22362 7541
rect 22306 7487 22362 7489
rect 22386 7541 22442 7543
rect 22386 7489 22438 7541
rect 22438 7489 22442 7541
rect 22386 7487 22442 7489
rect 22466 7541 22522 7543
rect 22466 7489 22518 7541
rect 22518 7489 22522 7541
rect 22466 7487 22522 7489
rect 22546 7541 22602 7543
rect 22546 7489 22598 7541
rect 22598 7489 22602 7541
rect 22546 7487 22602 7489
rect 22626 7541 22682 7543
rect 22626 7489 22678 7541
rect 22678 7489 22682 7541
rect 22626 7487 22682 7489
rect 22830 7541 22886 7543
rect 22830 7489 22834 7541
rect 22834 7489 22886 7541
rect 22830 7487 22886 7489
rect 22910 7541 22966 7543
rect 22910 7489 22914 7541
rect 22914 7489 22966 7541
rect 22910 7487 22966 7489
rect 22990 7541 23046 7543
rect 22990 7489 22994 7541
rect 22994 7489 23046 7541
rect 22990 7487 23046 7489
rect 23070 7541 23126 7543
rect 23070 7489 23074 7541
rect 23074 7489 23126 7541
rect 23070 7487 23126 7489
rect 23150 7541 23206 7543
rect 23150 7489 23154 7541
rect 23154 7489 23206 7541
rect 23150 7487 23206 7489
rect 23230 7541 23286 7543
rect 23230 7489 23234 7541
rect 23234 7489 23286 7541
rect 23230 7487 23286 7489
rect 23438 7541 23494 7543
rect 23438 7489 23490 7541
rect 23490 7489 23494 7541
rect 23438 7487 23494 7489
rect 23518 7541 23574 7543
rect 23518 7489 23570 7541
rect 23570 7489 23574 7541
rect 23518 7487 23574 7489
rect 23598 7541 23654 7543
rect 23598 7489 23650 7541
rect 23650 7489 23654 7541
rect 23598 7487 23654 7489
rect 23678 7541 23734 7543
rect 23678 7489 23730 7541
rect 23730 7489 23734 7541
rect 23678 7487 23734 7489
rect 23758 7541 23814 7543
rect 23758 7489 23810 7541
rect 23810 7489 23814 7541
rect 23758 7487 23814 7489
rect 23838 7541 23894 7543
rect 23838 7489 23890 7541
rect 23890 7489 23894 7541
rect 23838 7487 23894 7489
rect 24042 7541 24098 7543
rect 24042 7489 24046 7541
rect 24046 7489 24098 7541
rect 24042 7487 24098 7489
rect 24122 7541 24178 7543
rect 24122 7489 24126 7541
rect 24126 7489 24178 7541
rect 24122 7487 24178 7489
rect 24202 7541 24258 7543
rect 24202 7489 24206 7541
rect 24206 7489 24258 7541
rect 24202 7487 24258 7489
rect 24282 7541 24338 7543
rect 24282 7489 24286 7541
rect 24286 7489 24338 7541
rect 24282 7487 24338 7489
rect 24362 7541 24418 7543
rect 24362 7489 24366 7541
rect 24366 7489 24418 7541
rect 24362 7487 24418 7489
rect 24442 7541 24498 7543
rect 24442 7489 24446 7541
rect 24446 7489 24498 7541
rect 24442 7487 24498 7489
rect 24650 7541 24706 7543
rect 24650 7489 24702 7541
rect 24702 7489 24706 7541
rect 24650 7487 24706 7489
rect 24730 7541 24786 7543
rect 24730 7489 24782 7541
rect 24782 7489 24786 7541
rect 24730 7487 24786 7489
rect 24810 7541 24866 7543
rect 24810 7489 24862 7541
rect 24862 7489 24866 7541
rect 24810 7487 24866 7489
rect 24890 7541 24946 7543
rect 24890 7489 24942 7541
rect 24942 7489 24946 7541
rect 24890 7487 24946 7489
rect 24970 7541 25026 7543
rect 24970 7489 25022 7541
rect 25022 7489 25026 7541
rect 24970 7487 25026 7489
rect 25050 7541 25106 7543
rect 25050 7489 25102 7541
rect 25102 7489 25106 7541
rect 25050 7487 25106 7489
rect 25382 7544 25438 7546
rect 25382 7492 25434 7544
rect 25434 7492 25438 7544
rect 25382 7490 25438 7492
rect 25462 7544 25518 7546
rect 25462 7492 25514 7544
rect 25514 7492 25518 7544
rect 25462 7490 25518 7492
rect 25542 7544 25598 7546
rect 25542 7492 25594 7544
rect 25594 7492 25598 7544
rect 25542 7490 25598 7492
rect 25622 7544 25678 7546
rect 25622 7492 25674 7544
rect 25674 7492 25678 7544
rect 25622 7490 25678 7492
rect 25702 7544 25758 7546
rect 25702 7492 25754 7544
rect 25754 7492 25758 7544
rect 25702 7490 25758 7492
rect 25782 7544 25838 7546
rect 25782 7492 25834 7544
rect 25834 7492 25838 7544
rect 25782 7490 25838 7492
rect 25878 7535 25934 7537
rect 25878 7483 25880 7535
rect 25880 7483 25932 7535
rect 25932 7483 25934 7535
rect 25878 7481 25934 7483
rect 8626 1411 8682 1413
rect 8626 1359 8628 1411
rect 8628 1359 8680 1411
rect 8680 1359 8682 1411
rect 8626 1357 8682 1359
rect 8592 267 8648 269
rect 8592 215 8594 267
rect 8594 215 8646 267
rect 8646 215 8648 267
rect 8592 213 8648 215
rect 8620 -1109 8676 -1107
rect 8620 -1161 8622 -1109
rect 8622 -1161 8674 -1109
rect 8674 -1161 8676 -1109
rect 8620 -1163 8676 -1161
rect 10891 6934 11041 7080
rect 11203 6918 11353 7064
rect 10955 5974 11105 6120
rect 11261 5986 11411 6132
rect 10787 5346 10937 5492
rect 10823 4500 10973 4646
rect 11175 4504 11325 4650
rect 11621 4504 11771 4650
rect 10905 3646 11055 3792
rect 11255 3654 11405 3800
rect 12187 4508 12337 4654
rect 12853 4508 13003 4654
rect 13235 4492 13385 4638
rect 8828 1413 8884 1415
rect 8828 1361 8830 1413
rect 8830 1361 8882 1413
rect 8882 1361 8884 1413
rect 8828 1359 8884 1361
rect 9039 1411 9095 1413
rect 9039 1359 9041 1411
rect 9041 1359 9093 1411
rect 9093 1359 9095 1411
rect 9039 1357 9095 1359
rect 9229 1411 9285 1413
rect 9229 1359 9231 1411
rect 9231 1359 9283 1411
rect 9283 1359 9285 1411
rect 9229 1357 9285 1359
rect 9437 1413 9493 1415
rect 9437 1361 9439 1413
rect 9439 1361 9491 1413
rect 9491 1361 9493 1413
rect 9437 1359 9493 1361
rect 9639 1413 9695 1415
rect 9639 1361 9641 1413
rect 9641 1361 9693 1413
rect 9693 1361 9695 1413
rect 9639 1359 9695 1361
rect 9838 1415 9894 1417
rect 9838 1363 9840 1415
rect 9840 1363 9892 1415
rect 9892 1363 9894 1415
rect 9838 1361 9894 1363
rect 10033 1412 10089 1414
rect 10033 1360 10035 1412
rect 10035 1360 10087 1412
rect 10087 1360 10089 1412
rect 10033 1358 10089 1360
rect 9744 872 9800 874
rect 9744 820 9746 872
rect 9746 820 9798 872
rect 9798 820 9800 872
rect 9744 818 9800 820
rect 9963 876 10019 878
rect 9963 824 9965 876
rect 9965 824 10017 876
rect 10017 824 10019 876
rect 9963 822 10019 824
rect 8832 265 8888 267
rect 8832 213 8834 265
rect 8834 213 8886 265
rect 8886 213 8888 265
rect 8832 211 8888 213
rect 9154 264 9210 266
rect 9154 212 9156 264
rect 9156 212 9208 264
rect 9208 212 9210 264
rect 9154 210 9210 212
rect 9372 265 9428 267
rect 9372 213 9374 265
rect 9374 213 9426 265
rect 9426 213 9428 265
rect 9372 211 9428 213
rect 8838 -416 8894 -414
rect 8838 -468 8840 -416
rect 8840 -468 8892 -416
rect 8892 -468 8894 -416
rect 8838 -470 8894 -468
rect 9040 -420 9096 -418
rect 9040 -472 9042 -420
rect 9042 -472 9094 -420
rect 9094 -472 9096 -420
rect 9040 -474 9096 -472
rect 9229 -423 9285 -421
rect 9229 -475 9231 -423
rect 9231 -475 9283 -423
rect 9283 -475 9285 -423
rect 9229 -477 9285 -475
rect 9458 -422 9514 -420
rect 9458 -474 9460 -422
rect 9460 -474 9512 -422
rect 9512 -474 9514 -422
rect 9458 -476 9514 -474
rect 10234 1414 10290 1416
rect 10234 1362 10236 1414
rect 10236 1362 10288 1414
rect 10288 1362 10290 1414
rect 10234 1360 10290 1362
rect 10451 1412 10507 1414
rect 10451 1360 10453 1412
rect 10453 1360 10505 1412
rect 10505 1360 10507 1412
rect 10451 1358 10507 1360
rect 10246 876 10302 878
rect 10246 824 10248 876
rect 10248 824 10300 876
rect 10300 824 10302 876
rect 10246 822 10302 824
rect 10455 876 10511 878
rect 10455 824 10457 876
rect 10457 824 10509 876
rect 10509 824 10511 876
rect 10455 822 10511 824
rect 10725 1415 10781 1417
rect 10725 1363 10727 1415
rect 10727 1363 10779 1415
rect 10779 1363 10781 1415
rect 10725 1361 10781 1363
rect 10726 874 10782 876
rect 10726 822 10728 874
rect 10728 822 10780 874
rect 10780 822 10782 874
rect 10726 820 10782 822
rect 9783 -271 9839 -269
rect 9783 -323 9785 -271
rect 9785 -323 9837 -271
rect 9837 -323 9839 -271
rect 9783 -325 9839 -323
rect 10000 -271 10056 -269
rect 10000 -323 10002 -271
rect 10002 -323 10054 -271
rect 10054 -323 10056 -271
rect 10000 -325 10056 -323
rect 10219 -271 10275 -269
rect 10219 -323 10221 -271
rect 10221 -323 10273 -271
rect 10273 -323 10275 -271
rect 10219 -325 10275 -323
rect 10432 -275 10488 -273
rect 10432 -327 10434 -275
rect 10434 -327 10486 -275
rect 10486 -327 10488 -275
rect 10432 -329 10488 -327
rect 8853 -1113 8909 -1111
rect 8853 -1165 8855 -1113
rect 8855 -1165 8907 -1113
rect 8907 -1165 8909 -1113
rect 8853 -1167 8909 -1165
rect 9068 -1106 9124 -1104
rect 9068 -1158 9070 -1106
rect 9070 -1158 9122 -1106
rect 9122 -1158 9124 -1106
rect 9068 -1160 9124 -1158
rect 9286 -1109 9342 -1107
rect 9286 -1161 9288 -1109
rect 9288 -1161 9340 -1109
rect 9340 -1161 9342 -1109
rect 9286 -1163 9342 -1161
rect 9502 -1108 9558 -1106
rect 9502 -1160 9504 -1108
rect 9504 -1160 9556 -1108
rect 9556 -1160 9558 -1108
rect 9502 -1162 9558 -1160
rect 9994 -953 10050 -951
rect 9765 -965 9821 -963
rect 9765 -1017 9767 -965
rect 9767 -1017 9819 -965
rect 9819 -1017 9821 -965
rect 9994 -1005 9996 -953
rect 9996 -1005 10048 -953
rect 10048 -1005 10050 -953
rect 9994 -1007 10050 -1005
rect 10213 -963 10269 -961
rect 10213 -1015 10215 -963
rect 10215 -1015 10267 -963
rect 10267 -1015 10269 -963
rect 9765 -1019 9821 -1017
rect 10213 -1017 10269 -1015
rect 10405 -959 10461 -957
rect 10405 -1011 10407 -959
rect 10407 -1011 10459 -959
rect 10459 -1011 10461 -959
rect 10405 -1013 10461 -1011
rect 10643 -275 10699 -273
rect 10643 -327 10645 -275
rect 10645 -327 10697 -275
rect 10697 -327 10699 -275
rect 10643 -329 10699 -327
rect 8994 -1641 9050 -1639
rect 8994 -1693 8996 -1641
rect 8996 -1693 9048 -1641
rect 9048 -1693 9050 -1641
rect 8994 -1695 9050 -1693
rect 9193 -1644 9249 -1642
rect 9193 -1696 9195 -1644
rect 9195 -1696 9247 -1644
rect 9247 -1696 9249 -1644
rect 9193 -1698 9249 -1696
rect 9404 -1644 9460 -1642
rect 9404 -1696 9406 -1644
rect 9406 -1696 9458 -1644
rect 9458 -1696 9460 -1644
rect 9404 -1698 9460 -1696
rect 9610 -1644 9666 -1642
rect 9610 -1696 9612 -1644
rect 9612 -1696 9664 -1644
rect 9664 -1696 9666 -1644
rect 9610 -1698 9666 -1696
rect 9838 -1646 9894 -1644
rect 9838 -1698 9840 -1646
rect 9840 -1698 9892 -1646
rect 9892 -1698 9894 -1646
rect 9838 -1700 9894 -1698
rect 10082 -1646 10138 -1644
rect 10082 -1698 10084 -1646
rect 10084 -1698 10136 -1646
rect 10136 -1698 10138 -1646
rect 10082 -1700 10138 -1698
rect 10312 -1644 10368 -1642
rect 10312 -1696 10314 -1644
rect 10314 -1696 10366 -1644
rect 10366 -1696 10368 -1644
rect 10312 -1698 10368 -1696
rect 10518 -1644 10574 -1642
rect 10518 -1696 10520 -1644
rect 10520 -1696 10572 -1644
rect 10572 -1696 10574 -1644
rect 10518 -1698 10574 -1696
rect 11002 1408 11058 1410
rect 11002 1356 11004 1408
rect 11004 1356 11056 1408
rect 11056 1356 11058 1408
rect 11002 1354 11058 1356
rect 10899 -961 10955 -959
rect 10899 -1013 10901 -961
rect 10901 -1013 10953 -961
rect 10953 -1013 10955 -961
rect 10899 -1015 10955 -1013
rect 11225 1411 11281 1413
rect 11225 1359 11227 1411
rect 11227 1359 11279 1411
rect 11279 1359 11281 1411
rect 11225 1357 11281 1359
rect 11457 1410 11513 1412
rect 11457 1358 11459 1410
rect 11459 1358 11511 1410
rect 11511 1358 11513 1410
rect 11457 1356 11513 1358
rect 11276 269 11332 271
rect 11276 217 11278 269
rect 11278 217 11330 269
rect 11330 217 11332 269
rect 11276 215 11332 217
rect 11601 271 11657 273
rect 11601 219 11603 271
rect 11603 219 11655 271
rect 11655 219 11657 271
rect 11601 217 11657 219
rect 11869 271 11925 273
rect 11869 219 11871 271
rect 11871 219 11923 271
rect 11923 219 11925 271
rect 11869 217 11925 219
rect 11227 -419 11283 -417
rect 11227 -471 11229 -419
rect 11229 -471 11281 -419
rect 11281 -471 11283 -419
rect 11227 -473 11283 -471
rect 11442 -422 11498 -420
rect 11442 -474 11444 -422
rect 11444 -474 11496 -422
rect 11496 -474 11498 -422
rect 11442 -476 11498 -474
rect 11640 -425 11696 -423
rect 11640 -477 11642 -425
rect 11642 -477 11694 -425
rect 11694 -477 11696 -425
rect 11640 -479 11696 -477
rect 11835 -415 11891 -413
rect 11835 -467 11837 -415
rect 11837 -467 11889 -415
rect 11889 -467 11891 -415
rect 11835 -469 11891 -467
rect 12135 271 12191 273
rect 12135 219 12137 271
rect 12137 219 12189 271
rect 12189 219 12191 271
rect 12135 217 12191 219
rect 12375 269 12431 271
rect 12375 217 12377 269
rect 12377 217 12429 269
rect 12429 217 12431 269
rect 12375 215 12431 217
rect 12801 872 12857 874
rect 12801 820 12803 872
rect 12803 820 12855 872
rect 12855 820 12857 872
rect 12801 818 12857 820
rect 13093 1407 13149 1409
rect 13093 1355 13095 1407
rect 13095 1355 13147 1407
rect 13147 1355 13149 1407
rect 13093 1353 13149 1355
rect 13050 875 13106 877
rect 13050 823 13052 875
rect 13052 823 13104 875
rect 13104 823 13106 875
rect 13050 821 13106 823
rect 12767 -275 12823 -273
rect 12767 -327 12769 -275
rect 12769 -327 12821 -275
rect 12821 -327 12823 -275
rect 12767 -329 12823 -327
rect 12115 -417 12171 -415
rect 12115 -469 12117 -417
rect 12117 -469 12169 -417
rect 12169 -469 12171 -417
rect 12115 -471 12171 -469
rect 12334 -419 12390 -417
rect 12334 -471 12336 -419
rect 12336 -471 12388 -419
rect 12388 -471 12390 -419
rect 12334 -473 12390 -471
rect 11223 -1112 11279 -1110
rect 11223 -1164 11225 -1112
rect 11225 -1164 11277 -1112
rect 11277 -1164 11279 -1112
rect 11223 -1166 11279 -1164
rect 11413 -1112 11469 -1110
rect 11413 -1164 11415 -1112
rect 11415 -1164 11467 -1112
rect 11467 -1164 11469 -1112
rect 11413 -1166 11469 -1164
rect 11623 -1109 11679 -1107
rect 11623 -1161 11625 -1109
rect 11625 -1161 11677 -1109
rect 11677 -1161 11679 -1109
rect 11623 -1163 11679 -1161
rect 11840 -1112 11896 -1110
rect 11840 -1164 11842 -1112
rect 11842 -1164 11894 -1112
rect 11894 -1164 11896 -1112
rect 11840 -1166 11896 -1164
rect 12691 -962 12747 -960
rect 12691 -1014 12693 -962
rect 12693 -1014 12745 -962
rect 12745 -1014 12747 -962
rect 12691 -1016 12747 -1014
rect 12135 -1109 12191 -1107
rect 12135 -1161 12137 -1109
rect 12137 -1161 12189 -1109
rect 12189 -1161 12191 -1109
rect 12135 -1163 12191 -1161
rect 12359 -1104 12415 -1102
rect 12359 -1156 12361 -1104
rect 12361 -1156 12413 -1104
rect 12413 -1156 12415 -1104
rect 12359 -1158 12415 -1156
rect 10736 -1639 10792 -1637
rect 10736 -1691 10738 -1639
rect 10738 -1691 10790 -1639
rect 10790 -1691 10792 -1639
rect 10736 -1693 10792 -1691
rect 10939 -1645 10995 -1643
rect 10939 -1697 10941 -1645
rect 10941 -1697 10993 -1645
rect 10993 -1697 10995 -1645
rect 10939 -1699 10995 -1697
rect 11147 -1642 11203 -1640
rect 11147 -1694 11149 -1642
rect 11149 -1694 11201 -1642
rect 11201 -1694 11203 -1642
rect 11147 -1696 11203 -1694
rect 13045 -276 13101 -274
rect 13045 -328 13047 -276
rect 13047 -328 13099 -276
rect 13099 -328 13101 -276
rect 13045 -330 13101 -328
rect 11410 -1646 11466 -1644
rect 11410 -1698 11412 -1646
rect 11412 -1698 11464 -1646
rect 11464 -1698 11466 -1646
rect 11410 -1700 11466 -1698
rect 11618 -1645 11674 -1643
rect 11618 -1697 11620 -1645
rect 11620 -1697 11672 -1645
rect 11672 -1697 11674 -1645
rect 11618 -1699 11674 -1697
rect 11828 -1648 11884 -1646
rect 11828 -1700 11830 -1648
rect 11830 -1700 11882 -1648
rect 11882 -1700 11884 -1648
rect 11828 -1702 11884 -1700
rect 12028 -1642 12084 -1640
rect 12028 -1694 12030 -1642
rect 12030 -1694 12082 -1642
rect 12082 -1694 12084 -1642
rect 12028 -1696 12084 -1694
rect 12231 -1645 12287 -1643
rect 12231 -1697 12233 -1645
rect 12233 -1697 12285 -1645
rect 12285 -1697 12287 -1645
rect 12231 -1699 12287 -1697
rect 12441 -1645 12497 -1643
rect 12441 -1697 12443 -1645
rect 12443 -1697 12495 -1645
rect 12495 -1697 12497 -1645
rect 12441 -1699 12497 -1697
rect 12642 -1644 12698 -1642
rect 12642 -1696 12644 -1644
rect 12644 -1696 12696 -1644
rect 12696 -1696 12698 -1644
rect 12642 -1698 12698 -1696
rect 12858 -1643 12914 -1641
rect 12858 -1695 12860 -1643
rect 12860 -1695 12912 -1643
rect 12912 -1695 12914 -1643
rect 12858 -1697 12914 -1695
rect 13084 -964 13140 -962
rect 13084 -1016 13086 -964
rect 13086 -1016 13138 -964
rect 13138 -1016 13140 -964
rect 13084 -1018 13140 -1016
rect 13401 1408 13457 1410
rect 13401 1356 13403 1408
rect 13403 1356 13455 1408
rect 13455 1356 13457 1408
rect 13401 1354 13457 1356
rect 13394 861 13450 863
rect 13394 809 13396 861
rect 13396 809 13448 861
rect 13448 809 13450 861
rect 13394 807 13450 809
rect 13281 -956 13337 -954
rect 13281 -1008 13283 -956
rect 13283 -1008 13335 -956
rect 13335 -1008 13337 -956
rect 13281 -1010 13337 -1008
rect 13601 1409 13657 1411
rect 13601 1357 13603 1409
rect 13603 1357 13655 1409
rect 13655 1357 13657 1409
rect 13601 1355 13657 1357
rect 13820 1408 13876 1410
rect 13820 1356 13822 1408
rect 13822 1356 13874 1408
rect 13874 1356 13876 1408
rect 13820 1354 13876 1356
rect 14066 1407 14122 1409
rect 14066 1355 14068 1407
rect 14068 1355 14120 1407
rect 14120 1355 14122 1407
rect 14066 1353 14122 1355
rect 14274 1409 14330 1411
rect 14274 1357 14276 1409
rect 14276 1357 14328 1409
rect 14328 1357 14330 1409
rect 14274 1355 14330 1357
rect 14476 1410 14532 1412
rect 14476 1358 14478 1410
rect 14478 1358 14530 1410
rect 14530 1358 14532 1410
rect 14476 1356 14532 1358
rect 14669 1409 14725 1411
rect 14669 1357 14671 1409
rect 14671 1357 14723 1409
rect 14723 1357 14725 1409
rect 14669 1355 14725 1357
rect 13648 867 13704 869
rect 13648 815 13650 867
rect 13650 815 13702 867
rect 13702 815 13704 867
rect 13648 813 13704 815
rect 13877 867 13933 869
rect 13877 815 13879 867
rect 13879 815 13931 867
rect 13931 815 13933 867
rect 13877 813 13933 815
rect 14169 272 14225 274
rect 14169 220 14171 272
rect 14171 220 14223 272
rect 14223 220 14225 272
rect 14169 218 14225 220
rect 13617 -271 13673 -269
rect 13617 -323 13619 -271
rect 13619 -323 13671 -271
rect 13671 -323 13673 -271
rect 13617 -325 13673 -323
rect 13856 -271 13912 -269
rect 13856 -323 13858 -271
rect 13858 -323 13910 -271
rect 13910 -323 13912 -271
rect 13856 -325 13912 -323
rect 14155 -422 14211 -420
rect 14155 -474 14157 -422
rect 14157 -474 14209 -422
rect 14209 -474 14211 -422
rect 14155 -476 14211 -474
rect 14535 275 14591 277
rect 14535 223 14537 275
rect 14537 223 14589 275
rect 14589 223 14591 275
rect 14535 221 14591 223
rect 14779 275 14835 277
rect 14779 223 14781 275
rect 14781 223 14833 275
rect 14833 223 14835 275
rect 14779 221 14835 223
rect 15041 1408 15097 1410
rect 15041 1356 15043 1408
rect 15043 1356 15095 1408
rect 15095 1356 15097 1408
rect 15041 1354 15097 1356
rect 15230 1406 15286 1408
rect 15230 1354 15232 1406
rect 15232 1354 15284 1406
rect 15284 1354 15286 1406
rect 15230 1352 15286 1354
rect 15202 266 15258 268
rect 15202 214 15204 266
rect 15204 214 15256 266
rect 15256 214 15258 266
rect 15202 212 15258 214
rect 15520 1406 15576 1408
rect 15520 1354 15522 1406
rect 15522 1354 15574 1406
rect 15574 1354 15576 1406
rect 15520 1352 15576 1354
rect 15595 872 15651 874
rect 15595 820 15597 872
rect 15597 820 15649 872
rect 15649 820 15651 872
rect 15595 818 15651 820
rect 14506 -425 14562 -423
rect 14506 -477 14508 -425
rect 14508 -477 14560 -425
rect 14560 -477 14562 -425
rect 14506 -479 14562 -477
rect 14695 -427 14751 -425
rect 14695 -479 14697 -427
rect 14697 -479 14749 -427
rect 14749 -479 14751 -427
rect 14695 -481 14751 -479
rect 14900 -420 14956 -418
rect 14900 -472 14902 -420
rect 14902 -472 14954 -420
rect 14954 -472 14956 -420
rect 14900 -474 14956 -472
rect 15091 -418 15147 -416
rect 15091 -470 15093 -418
rect 15093 -470 15145 -418
rect 15145 -470 15147 -418
rect 15091 -472 15147 -470
rect 13611 -954 13667 -952
rect 13611 -1006 13613 -954
rect 13613 -1006 13665 -954
rect 13665 -1006 13667 -954
rect 13611 -1008 13667 -1006
rect 13807 -954 13863 -952
rect 13807 -1006 13809 -954
rect 13809 -1006 13861 -954
rect 13861 -1006 13863 -954
rect 13807 -1008 13863 -1006
rect 14237 -1111 14293 -1109
rect 14237 -1163 14239 -1111
rect 14239 -1163 14291 -1111
rect 14291 -1163 14293 -1111
rect 14237 -1165 14293 -1163
rect 14537 -1113 14593 -1111
rect 14537 -1165 14539 -1113
rect 14539 -1165 14591 -1113
rect 14591 -1165 14593 -1113
rect 14537 -1167 14593 -1165
rect 14789 -1109 14845 -1107
rect 14789 -1161 14791 -1109
rect 14791 -1161 14843 -1109
rect 14843 -1161 14845 -1109
rect 14789 -1163 14845 -1161
rect 15006 -1104 15062 -1102
rect 15006 -1156 15008 -1104
rect 15008 -1156 15060 -1104
rect 15060 -1156 15062 -1104
rect 15006 -1158 15062 -1156
rect 15207 -1107 15263 -1105
rect 15207 -1159 15209 -1107
rect 15209 -1159 15261 -1107
rect 15261 -1159 15263 -1107
rect 15207 -1161 15263 -1159
rect 13139 -1645 13195 -1643
rect 13139 -1697 13141 -1645
rect 13141 -1697 13193 -1645
rect 13193 -1697 13195 -1645
rect 13139 -1699 13195 -1697
rect 13359 -1650 13415 -1648
rect 13359 -1702 13361 -1650
rect 13361 -1702 13413 -1650
rect 13413 -1702 13415 -1650
rect 13359 -1704 13415 -1702
rect 13564 -1649 13620 -1647
rect 13564 -1701 13566 -1649
rect 13566 -1701 13618 -1649
rect 13618 -1701 13620 -1649
rect 13564 -1703 13620 -1701
rect 13785 -1643 13841 -1641
rect 13785 -1695 13787 -1643
rect 13787 -1695 13839 -1643
rect 13839 -1695 13841 -1643
rect 13785 -1697 13841 -1695
rect 13990 -1650 14046 -1648
rect 13990 -1702 13992 -1650
rect 13992 -1702 14044 -1650
rect 14044 -1702 14046 -1650
rect 13990 -1704 14046 -1702
rect 14199 -1649 14255 -1647
rect 14199 -1701 14201 -1649
rect 14201 -1701 14253 -1649
rect 14253 -1701 14255 -1649
rect 14199 -1703 14255 -1701
rect 14416 -1649 14472 -1647
rect 14416 -1701 14418 -1649
rect 14418 -1701 14470 -1649
rect 14470 -1701 14472 -1649
rect 14416 -1703 14472 -1701
rect 14630 -1644 14686 -1642
rect 14630 -1696 14632 -1644
rect 14632 -1696 14684 -1644
rect 14684 -1696 14686 -1644
rect 14630 -1698 14686 -1696
rect 14825 -1646 14881 -1644
rect 14825 -1698 14827 -1646
rect 14827 -1698 14879 -1646
rect 14879 -1698 14881 -1646
rect 14825 -1700 14881 -1698
rect 15020 -1649 15076 -1647
rect 15020 -1701 15022 -1649
rect 15022 -1701 15074 -1649
rect 15074 -1701 15076 -1649
rect 15020 -1703 15076 -1701
rect 15222 -1646 15278 -1644
rect 15222 -1698 15224 -1646
rect 15224 -1698 15276 -1646
rect 15276 -1698 15278 -1646
rect 15222 -1700 15278 -1698
rect 15793 1408 15849 1410
rect 15793 1356 15795 1408
rect 15795 1356 15847 1408
rect 15847 1356 15849 1408
rect 15793 1354 15849 1356
rect 15799 874 15855 876
rect 15799 822 15801 874
rect 15801 822 15853 874
rect 15853 822 15855 874
rect 15799 820 15855 822
rect 15714 -961 15770 -959
rect 15714 -1013 15716 -961
rect 15716 -1013 15768 -961
rect 15768 -1013 15770 -961
rect 15714 -1015 15770 -1013
rect 16122 872 16178 874
rect 16122 820 16124 872
rect 16124 820 16176 872
rect 16176 820 16178 872
rect 16122 818 16178 820
rect 16014 -273 16070 -271
rect 16014 -325 16016 -273
rect 16016 -325 16068 -273
rect 16068 -325 16070 -273
rect 16014 -327 16070 -325
rect 16241 -268 16297 -266
rect 16241 -320 16243 -268
rect 16243 -320 16295 -268
rect 16295 -320 16297 -268
rect 16241 -322 16297 -320
rect 16431 -266 16487 -264
rect 16431 -318 16433 -266
rect 16433 -318 16485 -266
rect 16485 -318 16487 -266
rect 16431 -320 16487 -318
rect 16647 -275 16703 -273
rect 16647 -327 16649 -275
rect 16649 -327 16701 -275
rect 16701 -327 16703 -275
rect 16647 -329 16703 -327
rect 17145 268 17201 270
rect 17145 216 17147 268
rect 17147 216 17199 268
rect 17199 216 17201 268
rect 17145 214 17201 216
rect 17397 265 17453 267
rect 17397 213 17399 265
rect 17399 213 17451 265
rect 17451 213 17453 265
rect 17397 211 17453 213
rect 17603 273 17659 275
rect 17603 221 17605 273
rect 17605 221 17657 273
rect 17657 221 17659 273
rect 17603 219 17659 221
rect 17886 267 17942 269
rect 17886 215 17888 267
rect 17888 215 17940 267
rect 17940 215 17942 267
rect 17886 213 17942 215
rect 17136 -416 17192 -414
rect 17136 -468 17138 -416
rect 17138 -468 17190 -416
rect 17190 -468 17192 -416
rect 17136 -470 17192 -468
rect 17326 -414 17382 -412
rect 17326 -466 17328 -414
rect 17328 -466 17380 -414
rect 17380 -466 17382 -414
rect 17326 -468 17382 -466
rect 17520 -416 17576 -414
rect 17520 -468 17522 -416
rect 17522 -468 17574 -416
rect 17574 -468 17576 -416
rect 17520 -470 17576 -468
rect 16015 -957 16071 -955
rect 16015 -1009 16017 -957
rect 16017 -1009 16069 -957
rect 16069 -1009 16071 -957
rect 16015 -1011 16071 -1009
rect 16221 -956 16277 -954
rect 16221 -1008 16223 -956
rect 16223 -1008 16275 -956
rect 16275 -1008 16277 -956
rect 16221 -1010 16277 -1008
rect 16431 -960 16487 -958
rect 16431 -1012 16433 -960
rect 16433 -1012 16485 -960
rect 16485 -1012 16487 -960
rect 16431 -1014 16487 -1012
rect 16642 -954 16698 -952
rect 16642 -1006 16644 -954
rect 16644 -1006 16696 -954
rect 16696 -1006 16698 -954
rect 16642 -1008 16698 -1006
rect 17092 -1116 17148 -1114
rect 17092 -1168 17094 -1116
rect 17094 -1168 17146 -1116
rect 17146 -1168 17148 -1116
rect 17092 -1170 17148 -1168
rect 17284 -1116 17340 -1114
rect 17284 -1168 17286 -1116
rect 17286 -1168 17338 -1116
rect 17338 -1168 17340 -1116
rect 17284 -1170 17340 -1168
rect 17484 -1116 17540 -1114
rect 17484 -1168 17486 -1116
rect 17486 -1168 17538 -1116
rect 17538 -1168 17540 -1116
rect 17484 -1170 17540 -1168
rect 15506 -1645 15562 -1643
rect 15506 -1697 15508 -1645
rect 15508 -1697 15560 -1645
rect 15560 -1697 15562 -1645
rect 15506 -1699 15562 -1697
rect 15705 -1644 15761 -1642
rect 15705 -1696 15707 -1644
rect 15707 -1696 15759 -1644
rect 15759 -1696 15761 -1644
rect 15705 -1698 15761 -1696
rect 15908 -1642 15964 -1640
rect 15908 -1694 15910 -1642
rect 15910 -1694 15962 -1642
rect 15962 -1694 15964 -1642
rect 15908 -1696 15964 -1694
rect 17831 -420 17887 -418
rect 17831 -472 17833 -420
rect 17833 -472 17885 -420
rect 17885 -472 17887 -420
rect 17831 -474 17887 -472
rect 16173 -1645 16229 -1643
rect 16173 -1697 16175 -1645
rect 16175 -1697 16227 -1645
rect 16227 -1697 16229 -1645
rect 16173 -1699 16229 -1697
rect 16371 -1646 16427 -1644
rect 16371 -1698 16373 -1646
rect 16373 -1698 16425 -1646
rect 16425 -1698 16427 -1646
rect 16371 -1700 16427 -1698
rect 16560 -1644 16616 -1642
rect 16560 -1696 16562 -1644
rect 16562 -1696 16614 -1644
rect 16614 -1696 16616 -1644
rect 16560 -1698 16616 -1696
rect 16772 -1644 16828 -1642
rect 16772 -1696 16774 -1644
rect 16774 -1696 16826 -1644
rect 16826 -1696 16828 -1644
rect 16772 -1698 16828 -1696
rect 16989 -1644 17045 -1642
rect 16989 -1696 16991 -1644
rect 16991 -1696 17043 -1644
rect 17043 -1696 17045 -1644
rect 16989 -1698 17045 -1696
rect 17194 -1648 17250 -1646
rect 17194 -1700 17196 -1648
rect 17196 -1700 17248 -1648
rect 17248 -1700 17250 -1648
rect 17194 -1702 17250 -1700
rect 17399 -1648 17455 -1646
rect 17399 -1700 17401 -1648
rect 17401 -1700 17453 -1648
rect 17453 -1700 17455 -1648
rect 17399 -1702 17455 -1700
rect 17607 -1643 17663 -1641
rect 17607 -1695 17609 -1643
rect 17609 -1695 17661 -1643
rect 17661 -1695 17663 -1643
rect 17607 -1697 17663 -1695
rect 18184 268 18240 270
rect 18184 216 18186 268
rect 18186 216 18238 268
rect 18238 216 18240 268
rect 18184 214 18240 216
rect 18102 -1108 18158 -1106
rect 18102 -1160 18104 -1108
rect 18104 -1160 18156 -1108
rect 18156 -1160 18158 -1108
rect 18102 -1162 18158 -1160
rect 18628 -272 18684 -270
rect 18628 -324 18630 -272
rect 18630 -324 18682 -272
rect 18682 -324 18684 -272
rect 18628 -326 18684 -324
rect 18857 -269 18913 -267
rect 18857 -321 18859 -269
rect 18859 -321 18911 -269
rect 18911 -321 18913 -269
rect 18857 -323 18913 -321
rect 19083 -264 19139 -262
rect 19083 -316 19085 -264
rect 19085 -316 19137 -264
rect 19137 -316 19139 -264
rect 19083 -318 19139 -316
rect 20016 269 20072 271
rect 20016 217 20018 269
rect 20018 217 20070 269
rect 20070 217 20072 269
rect 20016 215 20072 217
rect 23609 6320 23759 6466
rect 20226 271 20282 273
rect 20226 219 20228 271
rect 20228 219 20280 271
rect 20280 219 20282 271
rect 20226 217 20282 219
rect 19311 -272 19367 -270
rect 19311 -324 19313 -272
rect 19313 -324 19365 -272
rect 19365 -324 19367 -272
rect 19311 -326 19367 -324
rect 19547 -266 19603 -264
rect 19547 -318 19549 -266
rect 19549 -318 19601 -266
rect 19601 -318 19603 -266
rect 19547 -320 19603 -318
rect 19739 -275 19795 -273
rect 19739 -327 19741 -275
rect 19741 -327 19793 -275
rect 19793 -327 19795 -275
rect 19739 -329 19795 -327
rect 20014 -421 20070 -419
rect 20014 -473 20016 -421
rect 20016 -473 20068 -421
rect 20068 -473 20070 -421
rect 20014 -475 20070 -473
rect 18522 -965 18578 -963
rect 18522 -1017 18524 -965
rect 18524 -1017 18576 -965
rect 18576 -1017 18578 -965
rect 18522 -1019 18578 -1017
rect 18779 -958 18835 -956
rect 18779 -1010 18781 -958
rect 18781 -1010 18833 -958
rect 18833 -1010 18835 -958
rect 18779 -1012 18835 -1010
rect 19029 -962 19085 -960
rect 19029 -1014 19031 -962
rect 19031 -1014 19083 -962
rect 19083 -1014 19085 -962
rect 19029 -1016 19085 -1014
rect 19300 -957 19356 -955
rect 19300 -1009 19302 -957
rect 19302 -1009 19354 -957
rect 19354 -1009 19356 -957
rect 19300 -1011 19356 -1009
rect 19541 -954 19597 -952
rect 19541 -1006 19543 -954
rect 19543 -1006 19595 -954
rect 19595 -1006 19597 -954
rect 19541 -1008 19597 -1006
rect 19766 -958 19822 -956
rect 19766 -1010 19768 -958
rect 19768 -1010 19820 -958
rect 19820 -1010 19822 -958
rect 19766 -1012 19822 -1010
rect 20003 -1112 20059 -1110
rect 20003 -1164 20005 -1112
rect 20005 -1164 20057 -1112
rect 20057 -1164 20059 -1112
rect 20003 -1166 20059 -1164
rect 17890 -1644 17946 -1642
rect 17890 -1696 17892 -1644
rect 17892 -1696 17944 -1644
rect 17944 -1696 17946 -1644
rect 17890 -1698 17946 -1696
rect 18083 -1646 18139 -1644
rect 18083 -1698 18085 -1646
rect 18085 -1698 18137 -1646
rect 18137 -1698 18139 -1646
rect 18083 -1700 18139 -1698
rect 18309 -1648 18365 -1646
rect 18309 -1700 18311 -1648
rect 18311 -1700 18363 -1648
rect 18363 -1700 18365 -1648
rect 18309 -1702 18365 -1700
rect 20218 -421 20274 -419
rect 20218 -473 20220 -421
rect 20220 -473 20272 -421
rect 20272 -473 20274 -421
rect 20218 -475 20274 -473
rect 18574 -1648 18630 -1646
rect 18574 -1700 18576 -1648
rect 18576 -1700 18628 -1648
rect 18628 -1700 18630 -1648
rect 18574 -1702 18630 -1700
rect 18768 -1644 18824 -1642
rect 18768 -1696 18770 -1644
rect 18770 -1696 18822 -1644
rect 18822 -1696 18824 -1644
rect 18768 -1698 18824 -1696
rect 18966 -1653 19022 -1651
rect 18966 -1705 18968 -1653
rect 18968 -1705 19020 -1653
rect 19020 -1705 19022 -1653
rect 18966 -1707 19022 -1705
rect 19170 -1645 19226 -1643
rect 19170 -1697 19172 -1645
rect 19172 -1697 19224 -1645
rect 19224 -1697 19226 -1645
rect 19170 -1699 19226 -1697
rect 19390 -1642 19446 -1640
rect 19390 -1694 19392 -1642
rect 19392 -1694 19444 -1642
rect 19444 -1694 19446 -1642
rect 19390 -1696 19446 -1694
rect 19605 -1646 19661 -1644
rect 19605 -1698 19607 -1646
rect 19607 -1698 19659 -1646
rect 19659 -1698 19661 -1646
rect 19605 -1700 19661 -1698
rect 19833 -1643 19889 -1641
rect 19833 -1695 19835 -1643
rect 19835 -1695 19887 -1643
rect 19887 -1695 19889 -1643
rect 19833 -1697 19889 -1695
rect 20037 -1646 20093 -1644
rect 20037 -1698 20039 -1646
rect 20039 -1698 20091 -1646
rect 20091 -1698 20093 -1646
rect 20037 -1700 20093 -1698
rect 20259 -1112 20315 -1110
rect 20259 -1164 20261 -1112
rect 20261 -1164 20313 -1112
rect 20313 -1164 20315 -1112
rect 20259 -1166 20315 -1164
rect 20577 269 20633 271
rect 20577 217 20579 269
rect 20579 217 20631 269
rect 20631 217 20633 269
rect 20577 215 20633 217
rect 20494 -1112 20550 -1110
rect 20494 -1164 20496 -1112
rect 20496 -1164 20548 -1112
rect 20548 -1164 20550 -1112
rect 20494 -1166 20550 -1164
rect 20857 269 20913 271
rect 20857 217 20859 269
rect 20859 217 20911 269
rect 20911 217 20913 269
rect 20857 215 20913 217
rect 21174 268 21230 270
rect 21174 216 21176 268
rect 21176 216 21228 268
rect 21228 216 21230 268
rect 21174 214 21230 216
rect 20783 -425 20839 -423
rect 20783 -477 20785 -425
rect 20785 -477 20837 -425
rect 20837 -477 20839 -425
rect 20783 -479 20839 -477
rect 21474 -275 21530 -273
rect 21474 -327 21476 -275
rect 21476 -327 21528 -275
rect 21528 -327 21530 -275
rect 21474 -329 21530 -327
rect 21022 -423 21078 -421
rect 21022 -475 21024 -423
rect 21024 -475 21076 -423
rect 21076 -475 21078 -423
rect 21022 -477 21078 -475
rect 21226 -423 21282 -421
rect 21226 -475 21228 -423
rect 21228 -475 21280 -423
rect 21280 -475 21282 -423
rect 21226 -477 21282 -475
rect 23609 5894 23759 6040
rect 24679 7329 24735 7331
rect 24679 7277 24681 7329
rect 24681 7277 24733 7329
rect 24733 7277 24735 7329
rect 24679 7275 24735 7277
rect 24775 7320 24831 7322
rect 24775 7268 24779 7320
rect 24779 7268 24831 7320
rect 24775 7266 24831 7268
rect 24855 7320 24911 7322
rect 24855 7268 24859 7320
rect 24859 7268 24911 7320
rect 24855 7266 24911 7268
rect 24935 7320 24991 7322
rect 24935 7268 24939 7320
rect 24939 7268 24991 7320
rect 24935 7266 24991 7268
rect 25015 7320 25071 7322
rect 25015 7268 25019 7320
rect 25019 7268 25071 7320
rect 25015 7266 25071 7268
rect 25095 7320 25151 7322
rect 25095 7268 25099 7320
rect 25099 7268 25151 7320
rect 25095 7266 25151 7268
rect 25175 7320 25231 7322
rect 25175 7268 25179 7320
rect 25179 7268 25231 7320
rect 25175 7266 25231 7268
rect 25507 7323 25563 7325
rect 25507 7271 25511 7323
rect 25511 7271 25563 7323
rect 25507 7269 25563 7271
rect 25587 7323 25643 7325
rect 25587 7271 25591 7323
rect 25591 7271 25643 7323
rect 25587 7269 25643 7271
rect 25667 7323 25723 7325
rect 25667 7271 25671 7323
rect 25671 7271 25723 7323
rect 25667 7269 25723 7271
rect 25747 7323 25803 7325
rect 25747 7271 25751 7323
rect 25751 7271 25803 7323
rect 25747 7269 25803 7271
rect 25827 7323 25883 7325
rect 25827 7271 25831 7323
rect 25831 7271 25883 7323
rect 25827 7269 25883 7271
rect 25907 7323 25963 7325
rect 25907 7271 25911 7323
rect 25911 7271 25963 7323
rect 25907 7269 25963 7271
rect 26115 7323 26171 7325
rect 26115 7271 26167 7323
rect 26167 7271 26171 7323
rect 26115 7269 26171 7271
rect 26195 7323 26251 7325
rect 26195 7271 26247 7323
rect 26247 7271 26251 7323
rect 26195 7269 26251 7271
rect 26275 7323 26331 7325
rect 26275 7271 26327 7323
rect 26327 7271 26331 7323
rect 26275 7269 26331 7271
rect 26355 7323 26411 7325
rect 26355 7271 26407 7323
rect 26407 7271 26411 7323
rect 26355 7269 26411 7271
rect 26435 7323 26491 7325
rect 26435 7271 26487 7323
rect 26487 7271 26491 7323
rect 26435 7269 26491 7271
rect 26515 7323 26571 7325
rect 26515 7271 26567 7323
rect 26567 7271 26571 7323
rect 26515 7269 26571 7271
rect 26719 7323 26775 7325
rect 26719 7271 26723 7323
rect 26723 7271 26775 7323
rect 26719 7269 26775 7271
rect 26799 7323 26855 7325
rect 26799 7271 26803 7323
rect 26803 7271 26855 7323
rect 26799 7269 26855 7271
rect 26879 7323 26935 7325
rect 26879 7271 26883 7323
rect 26883 7271 26935 7323
rect 26879 7269 26935 7271
rect 26959 7323 27015 7325
rect 26959 7271 26963 7323
rect 26963 7271 27015 7323
rect 26959 7269 27015 7271
rect 27039 7323 27095 7325
rect 27039 7271 27043 7323
rect 27043 7271 27095 7323
rect 27039 7269 27095 7271
rect 27119 7323 27175 7325
rect 27119 7271 27123 7323
rect 27123 7271 27175 7323
rect 27119 7269 27175 7271
rect 27327 7323 27383 7325
rect 27327 7271 27379 7323
rect 27379 7271 27383 7323
rect 27327 7269 27383 7271
rect 27407 7323 27463 7325
rect 27407 7271 27459 7323
rect 27459 7271 27463 7323
rect 27407 7269 27463 7271
rect 27487 7323 27543 7325
rect 27487 7271 27539 7323
rect 27539 7271 27543 7323
rect 27487 7269 27543 7271
rect 27567 7323 27623 7325
rect 27567 7271 27619 7323
rect 27619 7271 27623 7323
rect 27567 7269 27623 7271
rect 27647 7323 27703 7325
rect 27647 7271 27699 7323
rect 27699 7271 27703 7323
rect 27647 7269 27703 7271
rect 27727 7323 27783 7325
rect 27727 7271 27779 7323
rect 27779 7271 27783 7323
rect 27727 7269 27783 7271
rect 27931 7323 27987 7325
rect 27931 7271 27935 7323
rect 27935 7271 27987 7323
rect 27931 7269 27987 7271
rect 28011 7323 28067 7325
rect 28011 7271 28015 7323
rect 28015 7271 28067 7323
rect 28011 7269 28067 7271
rect 28091 7323 28147 7325
rect 28091 7271 28095 7323
rect 28095 7271 28147 7323
rect 28091 7269 28147 7271
rect 28171 7323 28227 7325
rect 28171 7271 28175 7323
rect 28175 7271 28227 7323
rect 28171 7269 28227 7271
rect 28251 7323 28307 7325
rect 28251 7271 28255 7323
rect 28255 7271 28307 7323
rect 28251 7269 28307 7271
rect 28331 7323 28387 7325
rect 28331 7271 28335 7323
rect 28335 7271 28387 7323
rect 28331 7269 28387 7271
rect 28539 7323 28595 7325
rect 28539 7271 28591 7323
rect 28591 7271 28595 7323
rect 28539 7269 28595 7271
rect 28619 7323 28675 7325
rect 28619 7271 28671 7323
rect 28671 7271 28675 7323
rect 28619 7269 28675 7271
rect 28699 7323 28755 7325
rect 28699 7271 28751 7323
rect 28751 7271 28755 7323
rect 28699 7269 28755 7271
rect 28779 7323 28835 7325
rect 28779 7271 28831 7323
rect 28831 7271 28835 7323
rect 28779 7269 28835 7271
rect 28859 7323 28915 7325
rect 28859 7271 28911 7323
rect 28911 7271 28915 7323
rect 28859 7269 28915 7271
rect 28939 7323 28995 7325
rect 28939 7271 28991 7323
rect 28991 7271 28995 7323
rect 28939 7269 28995 7271
rect 29143 7323 29199 7325
rect 29143 7271 29147 7323
rect 29147 7271 29199 7323
rect 29143 7269 29199 7271
rect 29223 7323 29279 7325
rect 29223 7271 29227 7323
rect 29227 7271 29279 7323
rect 29223 7269 29279 7271
rect 29303 7323 29359 7325
rect 29303 7271 29307 7323
rect 29307 7271 29359 7323
rect 29303 7269 29359 7271
rect 29383 7323 29439 7325
rect 29383 7271 29387 7323
rect 29387 7271 29439 7323
rect 29383 7269 29439 7271
rect 29463 7323 29519 7325
rect 29463 7271 29467 7323
rect 29467 7271 29519 7323
rect 29463 7269 29519 7271
rect 29543 7323 29599 7325
rect 29543 7271 29547 7323
rect 29547 7271 29599 7323
rect 29543 7269 29599 7271
rect 29751 7323 29807 7325
rect 29751 7271 29803 7323
rect 29803 7271 29807 7323
rect 29751 7269 29807 7271
rect 29831 7323 29887 7325
rect 29831 7271 29883 7323
rect 29883 7271 29887 7323
rect 29831 7269 29887 7271
rect 29911 7323 29967 7325
rect 29911 7271 29963 7323
rect 29963 7271 29967 7323
rect 29911 7269 29967 7271
rect 29991 7323 30047 7325
rect 29991 7271 30043 7323
rect 30043 7271 30047 7323
rect 29991 7269 30047 7271
rect 30071 7323 30127 7325
rect 30071 7271 30123 7323
rect 30123 7271 30127 7323
rect 30071 7269 30127 7271
rect 30151 7323 30207 7325
rect 30151 7271 30203 7323
rect 30203 7271 30207 7323
rect 30151 7269 30207 7271
rect 30488 7267 30544 7269
rect 30488 7215 30490 7267
rect 30490 7215 30542 7267
rect 30542 7215 30544 7267
rect 30488 7213 30544 7215
rect 30493 7123 30549 7125
rect 30493 7071 30495 7123
rect 30495 7071 30547 7123
rect 30547 7071 30549 7123
rect 30493 7069 30549 7071
rect 30494 6971 30550 6973
rect 30494 6919 30496 6971
rect 30496 6919 30548 6971
rect 30548 6919 30550 6971
rect 30494 6917 30550 6919
rect 30494 6801 30550 6803
rect 30494 6749 30496 6801
rect 30496 6749 30548 6801
rect 30548 6749 30550 6801
rect 30494 6747 30550 6749
rect 24062 6724 24118 6726
rect 24062 6672 24064 6724
rect 24064 6672 24116 6724
rect 24116 6672 24118 6724
rect 24062 6670 24118 6672
rect 24193 6723 24249 6725
rect 24193 6671 24195 6723
rect 24195 6671 24247 6723
rect 24247 6671 24249 6723
rect 24193 6669 24249 6671
rect 24337 6724 24393 6726
rect 24337 6672 24339 6724
rect 24339 6672 24391 6724
rect 24391 6672 24393 6724
rect 24337 6670 24393 6672
rect 30493 6644 30549 6646
rect 30493 6592 30495 6644
rect 30495 6592 30547 6644
rect 30547 6592 30549 6644
rect 30493 6590 30549 6592
rect 30411 6402 30467 6404
rect 30411 6350 30413 6402
rect 30413 6350 30465 6402
rect 30465 6350 30467 6402
rect 30411 6348 30467 6350
rect 30788 6410 30844 6412
rect 30788 6358 30790 6410
rect 30790 6358 30842 6410
rect 30842 6358 30844 6410
rect 30788 6356 30844 6358
rect 30988 6410 31044 6412
rect 30988 6358 30990 6410
rect 30990 6358 31042 6410
rect 31042 6358 31044 6410
rect 30988 6356 31044 6358
rect 24080 6178 24136 6180
rect 24080 6126 24082 6178
rect 24082 6126 24134 6178
rect 24134 6126 24136 6178
rect 24080 6124 24136 6126
rect 24200 6178 24256 6180
rect 24200 6126 24202 6178
rect 24202 6126 24254 6178
rect 24254 6126 24256 6178
rect 24200 6124 24256 6126
rect 24343 6178 24399 6180
rect 24343 6126 24345 6178
rect 24345 6126 24397 6178
rect 24397 6126 24399 6178
rect 24343 6124 24399 6126
rect 23609 5668 23759 5814
rect 25161 6078 25225 6142
rect 25893 6081 25957 6145
rect 26121 6081 26185 6145
rect 27105 6081 27169 6145
rect 27333 6081 27397 6145
rect 28317 6081 28381 6145
rect 28545 6081 28609 6145
rect 29529 6081 29593 6145
rect 29757 6081 29821 6145
rect 30499 6141 30555 6143
rect 30499 6089 30501 6141
rect 30501 6089 30553 6141
rect 30553 6089 30555 6141
rect 30499 6087 30555 6089
rect 25517 5879 25581 5943
rect 26249 5879 26313 5943
rect 26467 5879 26531 5943
rect 27461 5879 27525 5943
rect 27679 5879 27743 5943
rect 28799 5879 28863 5943
rect 29017 5879 29081 5943
rect 29751 5879 29815 5943
rect 30499 5938 30555 5940
rect 30499 5886 30501 5938
rect 30501 5886 30553 5938
rect 30553 5886 30555 5938
rect 30499 5884 30555 5886
rect 30599 5768 30655 5770
rect 30599 5716 30601 5768
rect 30601 5716 30653 5768
rect 30653 5716 30655 5768
rect 30599 5714 30655 5716
rect 30408 5676 30464 5678
rect 30408 5624 30410 5676
rect 30410 5624 30462 5676
rect 30462 5624 30464 5676
rect 30408 5622 30464 5624
rect 23625 4934 23775 5080
rect 24665 4751 24721 4753
rect 24665 4699 24667 4751
rect 24667 4699 24719 4751
rect 24719 4699 24721 4751
rect 24665 4697 24721 4699
rect 25207 4754 25263 4756
rect 25207 4702 25209 4754
rect 25209 4702 25261 4754
rect 25261 4702 25263 4754
rect 25207 4700 25263 4702
rect 25287 4754 25343 4756
rect 25287 4702 25289 4754
rect 25289 4702 25341 4754
rect 25341 4702 25343 4754
rect 25287 4700 25343 4702
rect 25367 4754 25423 4756
rect 25367 4702 25369 4754
rect 25369 4702 25421 4754
rect 25421 4702 25423 4754
rect 25367 4700 25423 4702
rect 25447 4754 25503 4756
rect 25447 4702 25449 4754
rect 25449 4702 25501 4754
rect 25501 4702 25503 4754
rect 25447 4700 25503 4702
rect 25939 4754 25995 4756
rect 25939 4702 25941 4754
rect 25941 4702 25993 4754
rect 25993 4702 25995 4754
rect 25939 4700 25995 4702
rect 26019 4754 26075 4756
rect 26019 4702 26021 4754
rect 26021 4702 26073 4754
rect 26073 4702 26075 4754
rect 26019 4700 26075 4702
rect 26099 4754 26155 4756
rect 26099 4702 26101 4754
rect 26101 4702 26153 4754
rect 26153 4702 26155 4754
rect 26099 4700 26155 4702
rect 26179 4754 26235 4756
rect 26179 4702 26181 4754
rect 26181 4702 26233 4754
rect 26233 4702 26235 4754
rect 26179 4700 26235 4702
rect 26545 4754 26601 4756
rect 26545 4702 26547 4754
rect 26547 4702 26599 4754
rect 26599 4702 26601 4754
rect 26545 4700 26601 4702
rect 26625 4754 26681 4756
rect 26625 4702 26627 4754
rect 26627 4702 26679 4754
rect 26679 4702 26681 4754
rect 26625 4700 26681 4702
rect 26705 4754 26761 4756
rect 26705 4702 26707 4754
rect 26707 4702 26759 4754
rect 26759 4702 26761 4754
rect 26705 4700 26761 4702
rect 26785 4754 26841 4756
rect 26785 4702 26787 4754
rect 26787 4702 26839 4754
rect 26839 4702 26841 4754
rect 26785 4700 26841 4702
rect 27151 4754 27207 4756
rect 27151 4702 27153 4754
rect 27153 4702 27205 4754
rect 27205 4702 27207 4754
rect 27151 4700 27207 4702
rect 27231 4754 27287 4756
rect 27231 4702 27233 4754
rect 27233 4702 27285 4754
rect 27285 4702 27287 4754
rect 27231 4700 27287 4702
rect 27311 4754 27367 4756
rect 27311 4702 27313 4754
rect 27313 4702 27365 4754
rect 27365 4702 27367 4754
rect 27311 4700 27367 4702
rect 27391 4754 27447 4756
rect 27391 4702 27393 4754
rect 27393 4702 27445 4754
rect 27445 4702 27447 4754
rect 27391 4700 27447 4702
rect 27757 4754 27813 4756
rect 27757 4702 27759 4754
rect 27759 4702 27811 4754
rect 27811 4702 27813 4754
rect 27757 4700 27813 4702
rect 27837 4754 27893 4756
rect 27837 4702 27839 4754
rect 27839 4702 27891 4754
rect 27891 4702 27893 4754
rect 27837 4700 27893 4702
rect 27917 4754 27973 4756
rect 27917 4702 27919 4754
rect 27919 4702 27971 4754
rect 27971 4702 27973 4754
rect 27917 4700 27973 4702
rect 27997 4754 28053 4756
rect 27997 4702 27999 4754
rect 27999 4702 28051 4754
rect 28051 4702 28053 4754
rect 27997 4700 28053 4702
rect 28489 4754 28545 4756
rect 28489 4702 28491 4754
rect 28491 4702 28543 4754
rect 28543 4702 28545 4754
rect 28489 4700 28545 4702
rect 28569 4754 28625 4756
rect 28569 4702 28571 4754
rect 28571 4702 28623 4754
rect 28623 4702 28625 4754
rect 28569 4700 28625 4702
rect 28649 4754 28705 4756
rect 28649 4702 28651 4754
rect 28651 4702 28703 4754
rect 28703 4702 28705 4754
rect 28649 4700 28705 4702
rect 28729 4754 28785 4756
rect 28729 4702 28731 4754
rect 28731 4702 28783 4754
rect 28783 4702 28785 4754
rect 28729 4700 28785 4702
rect 29095 4754 29151 4756
rect 29095 4702 29097 4754
rect 29097 4702 29149 4754
rect 29149 4702 29151 4754
rect 29095 4700 29151 4702
rect 29175 4754 29231 4756
rect 29175 4702 29177 4754
rect 29177 4702 29229 4754
rect 29229 4702 29231 4754
rect 29175 4700 29231 4702
rect 29255 4754 29311 4756
rect 29255 4702 29257 4754
rect 29257 4702 29309 4754
rect 29309 4702 29311 4754
rect 29255 4700 29311 4702
rect 29335 4754 29391 4756
rect 29335 4702 29337 4754
rect 29337 4702 29389 4754
rect 29389 4702 29391 4754
rect 29335 4700 29391 4702
rect 29829 4754 29885 4756
rect 29829 4702 29831 4754
rect 29831 4702 29883 4754
rect 29883 4702 29885 4754
rect 29829 4700 29885 4702
rect 29909 4754 29965 4756
rect 29909 4702 29911 4754
rect 29911 4702 29963 4754
rect 29963 4702 29965 4754
rect 29909 4700 29965 4702
rect 29989 4754 30045 4756
rect 29989 4702 29991 4754
rect 29991 4702 30043 4754
rect 30043 4702 30045 4754
rect 29989 4700 30045 4702
rect 30069 4754 30125 4756
rect 30069 4702 30071 4754
rect 30071 4702 30123 4754
rect 30123 4702 30125 4754
rect 30069 4700 30125 4702
rect 23605 3942 23755 4088
rect 25712 4306 25768 4308
rect 25712 4254 25714 4306
rect 25714 4254 25766 4306
rect 25766 4254 25768 4306
rect 25712 4252 25768 4254
rect 25886 4305 25942 4307
rect 25886 4253 25888 4305
rect 25888 4253 25940 4305
rect 25940 4253 25942 4305
rect 25886 4251 25942 4253
rect 26111 4307 26167 4309
rect 26111 4255 26113 4307
rect 26113 4255 26165 4307
rect 26165 4255 26167 4307
rect 26111 4253 26167 4255
rect 26312 4309 26368 4311
rect 26312 4257 26314 4309
rect 26314 4257 26366 4309
rect 26366 4257 26368 4309
rect 26312 4255 26368 4257
rect 26535 4307 26591 4309
rect 26535 4255 26537 4307
rect 26537 4255 26589 4307
rect 26589 4255 26591 4307
rect 26535 4253 26591 4255
rect 26744 4312 26800 4314
rect 26744 4260 26746 4312
rect 26746 4260 26798 4312
rect 26798 4260 26800 4312
rect 26744 4258 26800 4260
rect 26972 4305 27028 4307
rect 26972 4253 26974 4305
rect 26974 4253 27026 4305
rect 27026 4253 27028 4305
rect 26972 4251 27028 4253
rect 27162 4309 27218 4311
rect 27162 4257 27164 4309
rect 27164 4257 27216 4309
rect 27216 4257 27218 4309
rect 27162 4255 27218 4257
rect 27367 4312 27423 4314
rect 27367 4260 27369 4312
rect 27369 4260 27421 4312
rect 27421 4260 27423 4312
rect 27367 4258 27423 4260
rect 27566 4312 27622 4314
rect 27566 4260 27568 4312
rect 27568 4260 27620 4312
rect 27620 4260 27622 4312
rect 27566 4258 27622 4260
rect 27782 4307 27838 4309
rect 27782 4255 27784 4307
rect 27784 4255 27836 4307
rect 27836 4255 27838 4307
rect 27782 4253 27838 4255
rect 27070 4119 27126 4121
rect 27070 4067 27072 4119
rect 27072 4067 27124 4119
rect 27124 4067 27126 4119
rect 27070 4065 27126 4067
rect 27455 4068 27511 4070
rect 27455 4016 27457 4068
rect 27457 4016 27509 4068
rect 27509 4016 27511 4068
rect 27455 4014 27511 4016
rect 28170 4312 28226 4314
rect 28170 4260 28172 4312
rect 28172 4260 28224 4312
rect 28224 4260 28226 4312
rect 28170 4258 28226 4260
rect 28405 4307 28461 4309
rect 28405 4255 28407 4307
rect 28407 4255 28459 4307
rect 28459 4255 28461 4307
rect 28405 4253 28461 4255
rect 28647 4309 28703 4311
rect 28647 4257 28649 4309
rect 28649 4257 28701 4309
rect 28701 4257 28703 4309
rect 28647 4255 28703 4257
rect 28879 4310 28935 4312
rect 28879 4258 28881 4310
rect 28881 4258 28933 4310
rect 28933 4258 28935 4310
rect 28879 4256 28935 4258
rect 29108 4313 29164 4315
rect 29108 4261 29110 4313
rect 29110 4261 29162 4313
rect 29162 4261 29164 4313
rect 29108 4259 29164 4261
rect 29357 4305 29413 4307
rect 29357 4253 29359 4305
rect 29359 4253 29411 4305
rect 29411 4253 29413 4305
rect 29357 4251 29413 4253
rect 29575 4309 29631 4311
rect 29575 4257 29577 4309
rect 29577 4257 29629 4309
rect 29629 4257 29631 4309
rect 29575 4255 29631 4257
rect 29804 4305 29860 4307
rect 29804 4253 29806 4305
rect 29806 4253 29858 4305
rect 29858 4253 29860 4305
rect 29804 4251 29860 4253
rect 30025 4307 30081 4309
rect 30025 4255 30027 4307
rect 30027 4255 30079 4307
rect 30079 4255 30081 4307
rect 30025 4253 30081 4255
rect 30241 4312 30297 4314
rect 30241 4260 30243 4312
rect 30243 4260 30295 4312
rect 30295 4260 30297 4312
rect 30241 4258 30297 4260
rect 29465 4118 29521 4120
rect 29465 4066 29467 4118
rect 29467 4066 29519 4118
rect 29519 4066 29521 4118
rect 29465 4064 29521 4066
rect 29850 4069 29906 4071
rect 29850 4017 29852 4069
rect 29852 4017 29904 4069
rect 29904 4017 29906 4069
rect 29850 4015 29906 4017
rect 25714 3723 25770 3725
rect 25714 3671 25716 3723
rect 25716 3671 25768 3723
rect 25768 3671 25770 3723
rect 25714 3669 25770 3671
rect 25889 3721 25945 3723
rect 25889 3669 25891 3721
rect 25891 3669 25943 3721
rect 25943 3669 25945 3721
rect 25889 3667 25945 3669
rect 26086 3723 26142 3725
rect 26086 3671 26088 3723
rect 26088 3671 26140 3723
rect 26140 3671 26142 3723
rect 26086 3669 26142 3671
rect 26305 3726 26361 3728
rect 26305 3674 26307 3726
rect 26307 3674 26359 3726
rect 26359 3674 26361 3726
rect 26305 3672 26361 3674
rect 26537 3722 26593 3724
rect 26537 3670 26539 3722
rect 26539 3670 26591 3722
rect 26591 3670 26593 3722
rect 26537 3668 26593 3670
rect 26761 3729 26817 3731
rect 26761 3677 26763 3729
rect 26763 3677 26815 3729
rect 26815 3677 26817 3729
rect 26761 3675 26817 3677
rect 23611 3264 23761 3410
rect 21678 -270 21734 -268
rect 21678 -322 21680 -270
rect 21680 -322 21732 -270
rect 21732 -322 21734 -270
rect 21678 -324 21734 -322
rect 21869 -275 21925 -273
rect 21869 -327 21871 -275
rect 21871 -327 21923 -275
rect 21923 -327 21925 -275
rect 21869 -329 21925 -327
rect 22071 -276 22127 -274
rect 22071 -328 22073 -276
rect 22073 -328 22125 -276
rect 22125 -328 22127 -276
rect 22071 -330 22127 -328
rect 22361 -275 22417 -273
rect 22361 -327 22363 -275
rect 22363 -327 22415 -275
rect 22415 -327 22417 -275
rect 22361 -329 22417 -327
rect 21473 -960 21529 -958
rect 21473 -1012 21475 -960
rect 21475 -1012 21527 -960
rect 21527 -1012 21529 -960
rect 21473 -1014 21529 -1012
rect 20783 -1110 20839 -1108
rect 20783 -1162 20785 -1110
rect 20785 -1162 20837 -1110
rect 20837 -1162 20839 -1110
rect 20783 -1164 20839 -1162
rect 20973 -1112 21029 -1110
rect 20973 -1164 20975 -1112
rect 20975 -1164 21027 -1112
rect 21027 -1164 21029 -1112
rect 20973 -1166 21029 -1164
rect 21177 -1110 21233 -1108
rect 21177 -1162 21179 -1110
rect 21179 -1162 21231 -1110
rect 21231 -1162 21233 -1110
rect 21177 -1164 21233 -1162
rect 21674 -959 21730 -957
rect 21674 -1011 21676 -959
rect 21676 -1011 21728 -959
rect 21728 -1011 21730 -959
rect 21674 -1013 21730 -1011
rect 21892 -963 21948 -961
rect 21892 -1015 21894 -963
rect 21894 -1015 21946 -963
rect 21946 -1015 21948 -963
rect 21892 -1017 21948 -1015
rect 22099 -959 22155 -957
rect 22099 -1011 22101 -959
rect 22101 -1011 22153 -959
rect 22153 -1011 22155 -959
rect 22099 -1013 22155 -1011
rect 22304 -960 22360 -958
rect 22304 -1012 22306 -960
rect 22306 -1012 22358 -960
rect 22358 -1012 22360 -960
rect 22304 -1014 22360 -1012
rect 20275 -1644 20331 -1642
rect 20275 -1696 20277 -1644
rect 20277 -1696 20329 -1644
rect 20329 -1696 20331 -1644
rect 20275 -1698 20331 -1696
rect 20468 -1643 20524 -1641
rect 20468 -1695 20470 -1643
rect 20470 -1695 20522 -1643
rect 20522 -1695 20524 -1643
rect 20468 -1697 20524 -1695
rect 20665 -1648 20721 -1646
rect 20665 -1700 20667 -1648
rect 20667 -1700 20719 -1648
rect 20719 -1700 20721 -1648
rect 20665 -1702 20721 -1700
rect 22646 -276 22702 -274
rect 22646 -328 22648 -276
rect 22648 -328 22700 -276
rect 22700 -328 22702 -276
rect 22646 -330 22702 -328
rect 20921 -1645 20977 -1643
rect 20921 -1697 20923 -1645
rect 20923 -1697 20975 -1645
rect 20975 -1697 20977 -1645
rect 20921 -1699 20977 -1697
rect 21160 -1649 21216 -1647
rect 21160 -1701 21162 -1649
rect 21162 -1701 21214 -1649
rect 21214 -1701 21216 -1649
rect 21160 -1703 21216 -1701
rect 21393 -1653 21449 -1651
rect 21393 -1705 21395 -1653
rect 21395 -1705 21447 -1653
rect 21447 -1705 21449 -1653
rect 21393 -1707 21449 -1705
rect 21614 -1648 21670 -1646
rect 21614 -1700 21616 -1648
rect 21616 -1700 21668 -1648
rect 21668 -1700 21670 -1648
rect 21614 -1702 21670 -1700
rect 21805 -1648 21861 -1646
rect 21805 -1700 21807 -1648
rect 21807 -1700 21859 -1648
rect 21859 -1700 21861 -1648
rect 21805 -1702 21861 -1700
rect 22033 -1646 22089 -1644
rect 22033 -1698 22035 -1646
rect 22035 -1698 22087 -1646
rect 22087 -1698 22089 -1646
rect 22033 -1700 22089 -1698
rect 22230 -1651 22286 -1649
rect 22230 -1703 22232 -1651
rect 22232 -1703 22284 -1651
rect 22284 -1703 22286 -1651
rect 22230 -1705 22286 -1703
rect 22442 -1651 22498 -1649
rect 22442 -1703 22444 -1651
rect 22444 -1703 22496 -1651
rect 22496 -1703 22498 -1651
rect 22442 -1705 22498 -1703
rect 22651 -964 22707 -962
rect 22651 -1016 22653 -964
rect 22653 -1016 22705 -964
rect 22705 -1016 22707 -964
rect 22651 -1018 22707 -1016
rect 22964 266 23020 268
rect 22964 214 22966 266
rect 22966 214 23018 266
rect 23018 214 23020 266
rect 22964 212 23020 214
rect 22963 -1104 23019 -1102
rect 22963 -1156 22965 -1104
rect 22965 -1156 23017 -1104
rect 23017 -1156 23019 -1104
rect 22963 -1158 23019 -1156
rect 23259 266 23315 268
rect 23259 214 23261 266
rect 23261 214 23313 266
rect 23313 214 23315 266
rect 23259 212 23315 214
rect 23546 266 23602 268
rect 23546 214 23548 266
rect 23548 214 23600 266
rect 23600 214 23602 266
rect 23546 212 23602 214
rect 23836 266 23892 268
rect 23836 214 23838 266
rect 23838 214 23890 266
rect 23890 214 23892 266
rect 23836 212 23892 214
rect 23186 -415 23242 -413
rect 23186 -467 23188 -415
rect 23188 -467 23240 -415
rect 23240 -467 23242 -415
rect 23186 -469 23242 -467
rect 23419 -417 23475 -415
rect 23419 -469 23421 -417
rect 23421 -469 23473 -417
rect 23473 -469 23475 -417
rect 23419 -471 23475 -469
rect 23626 -419 23682 -417
rect 23626 -471 23628 -419
rect 23628 -471 23680 -419
rect 23680 -471 23682 -419
rect 23626 -473 23682 -471
rect 23835 -417 23891 -415
rect 23835 -469 23837 -417
rect 23837 -469 23889 -417
rect 23889 -469 23891 -417
rect 23835 -471 23891 -469
rect 24120 269 24176 271
rect 24120 217 24122 269
rect 24122 217 24174 269
rect 24174 217 24176 269
rect 24120 215 24176 217
rect 26973 3717 27029 3719
rect 26973 3665 26975 3717
rect 26975 3665 27027 3717
rect 27027 3665 27029 3717
rect 26973 3663 27029 3665
rect 27195 3713 27251 3715
rect 27195 3661 27197 3713
rect 27197 3661 27249 3713
rect 27249 3661 27251 3713
rect 27195 3659 27251 3661
rect 27418 3710 27474 3712
rect 27418 3658 27420 3710
rect 27420 3658 27472 3710
rect 27472 3658 27474 3710
rect 27418 3656 27474 3658
rect 27628 3710 27684 3712
rect 27628 3658 27630 3710
rect 27630 3658 27682 3710
rect 27682 3658 27684 3710
rect 27628 3656 27684 3658
rect 27841 3710 27897 3712
rect 27841 3658 27843 3710
rect 27843 3658 27895 3710
rect 27895 3658 27897 3710
rect 27841 3656 27897 3658
rect 28158 3703 28214 3705
rect 28158 3651 28160 3703
rect 28160 3651 28212 3703
rect 28212 3651 28214 3703
rect 28158 3649 28214 3651
rect 28360 3706 28416 3708
rect 28360 3654 28362 3706
rect 28362 3654 28414 3706
rect 28414 3654 28416 3706
rect 28360 3652 28416 3654
rect 28561 3707 28617 3709
rect 28561 3655 28563 3707
rect 28563 3655 28615 3707
rect 28615 3655 28617 3707
rect 28561 3653 28617 3655
rect 28740 3708 28796 3710
rect 28740 3656 28742 3708
rect 28742 3656 28794 3708
rect 28794 3656 28796 3708
rect 28740 3654 28796 3656
rect 28932 3712 28988 3714
rect 28932 3660 28934 3712
rect 28934 3660 28986 3712
rect 28986 3660 28988 3712
rect 28932 3658 28988 3660
rect 29117 3709 29173 3711
rect 29117 3657 29119 3709
rect 29119 3657 29171 3709
rect 29171 3657 29173 3709
rect 29117 3655 29173 3657
rect 25741 3074 25797 3076
rect 25741 3022 25743 3074
rect 25743 3022 25795 3074
rect 25795 3022 25797 3074
rect 25741 3020 25797 3022
rect 25957 3079 26013 3081
rect 25957 3027 25959 3079
rect 25959 3027 26011 3079
rect 26011 3027 26013 3079
rect 25957 3025 26013 3027
rect 26163 3080 26219 3082
rect 26163 3028 26165 3080
rect 26165 3028 26217 3080
rect 26217 3028 26219 3080
rect 26163 3026 26219 3028
rect 26365 3072 26421 3074
rect 26365 3020 26367 3072
rect 26367 3020 26419 3072
rect 26419 3020 26421 3072
rect 26365 3018 26421 3020
rect 26561 3074 26617 3076
rect 26561 3022 26563 3074
rect 26563 3022 26615 3074
rect 26615 3022 26617 3074
rect 26561 3020 26617 3022
rect 26786 3076 26842 3078
rect 26786 3024 26788 3076
rect 26788 3024 26840 3076
rect 26840 3024 26842 3076
rect 26786 3022 26842 3024
rect 27001 3072 27057 3074
rect 27001 3020 27003 3072
rect 27003 3020 27055 3072
rect 27055 3020 27057 3072
rect 27001 3018 27057 3020
rect 27236 3072 27292 3074
rect 27236 3020 27238 3072
rect 27238 3020 27290 3072
rect 27290 3020 27292 3072
rect 27236 3018 27292 3020
rect 27444 3075 27500 3077
rect 27444 3023 27446 3075
rect 27446 3023 27498 3075
rect 27498 3023 27500 3075
rect 27444 3021 27500 3023
rect 27686 3075 27742 3077
rect 27686 3023 27688 3075
rect 27688 3023 27740 3075
rect 27740 3023 27742 3075
rect 27686 3021 27742 3023
rect 27884 3076 27940 3078
rect 27884 3024 27886 3076
rect 27886 3024 27938 3076
rect 27938 3024 27940 3076
rect 27884 3022 27940 3024
rect 27075 2845 27131 2847
rect 27075 2793 27077 2845
rect 27077 2793 27129 2845
rect 27129 2793 27131 2845
rect 27075 2791 27131 2793
rect 24401 -271 24457 -269
rect 24401 -323 24403 -271
rect 24403 -323 24455 -271
rect 24455 -323 24457 -271
rect 24401 -325 24457 -323
rect 24595 -267 24651 -265
rect 24595 -319 24597 -267
rect 24597 -319 24649 -267
rect 24649 -319 24651 -267
rect 24595 -321 24651 -319
rect 24784 -270 24840 -268
rect 24784 -322 24786 -270
rect 24786 -322 24838 -270
rect 24838 -322 24840 -270
rect 24784 -324 24840 -322
rect 24115 -415 24171 -413
rect 24115 -467 24117 -415
rect 24117 -467 24169 -415
rect 24169 -467 24171 -415
rect 24115 -469 24171 -467
rect 23205 -1108 23261 -1106
rect 23205 -1160 23207 -1108
rect 23207 -1160 23259 -1108
rect 23259 -1160 23261 -1108
rect 23205 -1162 23261 -1160
rect 23405 -1109 23461 -1107
rect 23405 -1161 23407 -1109
rect 23407 -1161 23459 -1109
rect 23459 -1161 23461 -1109
rect 23405 -1163 23461 -1161
rect 23595 -1101 23651 -1099
rect 23595 -1153 23597 -1101
rect 23597 -1153 23649 -1101
rect 23649 -1153 23651 -1101
rect 23595 -1155 23651 -1153
rect 23816 -1103 23872 -1101
rect 23816 -1155 23818 -1103
rect 23818 -1155 23870 -1103
rect 23870 -1155 23872 -1103
rect 23816 -1157 23872 -1155
rect 24403 -960 24459 -958
rect 24403 -1012 24405 -960
rect 24405 -1012 24457 -960
rect 24457 -1012 24459 -960
rect 24403 -1014 24459 -1012
rect 24594 -957 24650 -955
rect 24594 -1009 24596 -957
rect 24596 -1009 24648 -957
rect 24648 -1009 24650 -957
rect 24594 -1011 24650 -1009
rect 24789 -955 24845 -953
rect 24789 -1007 24791 -955
rect 24791 -1007 24843 -955
rect 24843 -1007 24845 -955
rect 24789 -1009 24845 -1007
rect 24112 -1108 24168 -1106
rect 24112 -1160 24114 -1108
rect 24114 -1160 24166 -1108
rect 24166 -1160 24168 -1108
rect 24112 -1162 24168 -1160
rect 22669 -1648 22725 -1646
rect 22669 -1700 22671 -1648
rect 22671 -1700 22723 -1648
rect 22723 -1700 22725 -1648
rect 22669 -1702 22725 -1700
rect 22858 -1647 22914 -1645
rect 22858 -1699 22860 -1647
rect 22860 -1699 22912 -1647
rect 22912 -1699 22914 -1647
rect 22858 -1701 22914 -1699
rect 23084 -1646 23140 -1644
rect 23084 -1698 23086 -1646
rect 23086 -1698 23138 -1646
rect 23138 -1698 23140 -1646
rect 23084 -1700 23140 -1698
rect 25007 -268 25063 -266
rect 25007 -320 25009 -268
rect 25009 -320 25061 -268
rect 25061 -320 25063 -268
rect 25007 -322 25063 -320
rect 23338 -1646 23394 -1644
rect 23338 -1698 23340 -1646
rect 23340 -1698 23392 -1646
rect 23392 -1698 23394 -1646
rect 23338 -1700 23394 -1698
rect 23582 -1649 23638 -1647
rect 23582 -1701 23584 -1649
rect 23584 -1701 23636 -1649
rect 23636 -1701 23638 -1649
rect 23582 -1703 23638 -1701
rect 23812 -1650 23868 -1648
rect 23812 -1702 23814 -1650
rect 23814 -1702 23866 -1650
rect 23866 -1702 23868 -1650
rect 23812 -1704 23868 -1702
rect 24070 -1647 24126 -1645
rect 24070 -1699 24072 -1647
rect 24072 -1699 24124 -1647
rect 24124 -1699 24126 -1647
rect 24070 -1701 24126 -1699
rect 24280 -1647 24336 -1645
rect 24280 -1699 24282 -1647
rect 24282 -1699 24334 -1647
rect 24334 -1699 24336 -1647
rect 24280 -1701 24336 -1699
rect 24505 -1647 24561 -1645
rect 24505 -1699 24507 -1647
rect 24507 -1699 24559 -1647
rect 24559 -1699 24561 -1647
rect 24505 -1701 24561 -1699
rect 24724 -1650 24780 -1648
rect 24724 -1702 24726 -1650
rect 24726 -1702 24778 -1650
rect 24778 -1702 24780 -1650
rect 24724 -1704 24780 -1702
rect 27458 2786 27514 2788
rect 27458 2734 27460 2786
rect 27460 2734 27512 2786
rect 27512 2734 27514 2786
rect 27458 2732 27514 2734
rect 29349 3708 29405 3710
rect 29349 3656 29351 3708
rect 29351 3656 29403 3708
rect 29403 3656 29405 3708
rect 29349 3654 29405 3656
rect 29554 3710 29610 3712
rect 29554 3658 29556 3710
rect 29556 3658 29608 3710
rect 29608 3658 29610 3710
rect 29554 3656 29610 3658
rect 29760 3712 29816 3714
rect 29760 3660 29762 3712
rect 29762 3660 29814 3712
rect 29814 3660 29816 3712
rect 29760 3658 29816 3660
rect 29968 3719 30024 3721
rect 29968 3667 29970 3719
rect 29970 3667 30022 3719
rect 30022 3667 30024 3719
rect 29968 3665 30024 3667
rect 30190 3720 30246 3722
rect 30190 3668 30192 3720
rect 30192 3668 30244 3720
rect 30244 3668 30246 3720
rect 30190 3666 30246 3668
rect 28191 3076 28247 3078
rect 28191 3024 28193 3076
rect 28193 3024 28245 3076
rect 28245 3024 28247 3076
rect 28191 3022 28247 3024
rect 28416 3077 28472 3079
rect 28416 3025 28418 3077
rect 28418 3025 28470 3077
rect 28470 3025 28472 3077
rect 28416 3023 28472 3025
rect 28645 3076 28701 3078
rect 28645 3024 28647 3076
rect 28647 3024 28699 3076
rect 28699 3024 28701 3076
rect 28645 3022 28701 3024
rect 28861 3080 28917 3082
rect 28861 3028 28863 3080
rect 28863 3028 28915 3080
rect 28915 3028 28917 3080
rect 28861 3026 28917 3028
rect 29084 3083 29140 3085
rect 29084 3031 29086 3083
rect 29086 3031 29138 3083
rect 29138 3031 29140 3083
rect 29084 3029 29140 3031
rect 29308 3079 29364 3081
rect 29308 3027 29310 3079
rect 29310 3027 29362 3079
rect 29362 3027 29364 3079
rect 29308 3025 29364 3027
rect 29535 3068 29591 3070
rect 29535 3016 29537 3068
rect 29537 3016 29589 3068
rect 29589 3016 29591 3068
rect 29535 3014 29591 3016
rect 29748 3067 29804 3069
rect 29748 3015 29750 3067
rect 29750 3015 29802 3067
rect 29802 3015 29804 3067
rect 29748 3013 29804 3015
rect 29959 3071 30015 3073
rect 29959 3019 29961 3071
rect 29961 3019 30013 3071
rect 30013 3019 30015 3071
rect 29959 3017 30015 3019
rect 30186 3072 30242 3074
rect 30186 3020 30188 3072
rect 30188 3020 30240 3072
rect 30240 3020 30242 3072
rect 30186 3018 30242 3020
rect 29467 2847 29523 2849
rect 29467 2795 29469 2847
rect 29469 2795 29521 2847
rect 29521 2795 29523 2847
rect 29467 2793 29523 2795
rect 29844 2793 29900 2795
rect 29844 2741 29846 2793
rect 29846 2741 29898 2793
rect 29898 2741 29900 2793
rect 29844 2739 29900 2741
rect 25767 2429 25823 2431
rect 25767 2377 25769 2429
rect 25769 2377 25821 2429
rect 25821 2377 25823 2429
rect 25767 2375 25823 2377
rect 25992 2438 26048 2440
rect 25992 2386 25994 2438
rect 25994 2386 26046 2438
rect 26046 2386 26048 2438
rect 25992 2384 26048 2386
rect 26269 2435 26325 2437
rect 26269 2383 26271 2435
rect 26271 2383 26323 2435
rect 26323 2383 26325 2435
rect 26269 2381 26325 2383
rect 26490 2438 26546 2440
rect 26490 2386 26492 2438
rect 26492 2386 26544 2438
rect 26544 2386 26546 2438
rect 26490 2384 26546 2386
rect 26735 2435 26791 2437
rect 26735 2383 26737 2435
rect 26737 2383 26789 2435
rect 26789 2383 26791 2435
rect 26735 2381 26791 2383
rect 26961 2439 27017 2441
rect 26961 2387 26963 2439
rect 26963 2387 27015 2439
rect 27015 2387 27017 2439
rect 26961 2385 27017 2387
rect 27173 2437 27229 2439
rect 27173 2385 27175 2437
rect 27175 2385 27227 2437
rect 27227 2385 27229 2437
rect 27173 2383 27229 2385
rect 27393 2443 27449 2445
rect 27393 2391 27395 2443
rect 27395 2391 27447 2443
rect 27447 2391 27449 2443
rect 27393 2389 27449 2391
rect 27631 2445 27687 2447
rect 27631 2393 27633 2445
rect 27633 2393 27685 2445
rect 27685 2393 27687 2445
rect 27631 2391 27687 2393
rect 27844 2447 27900 2449
rect 27844 2395 27846 2447
rect 27846 2395 27898 2447
rect 27898 2395 27900 2447
rect 27844 2393 27900 2395
rect 28231 2437 28287 2439
rect 28231 2385 28233 2437
rect 28233 2385 28285 2437
rect 28285 2385 28287 2437
rect 28231 2383 28287 2385
rect 28578 2438 28634 2440
rect 28578 2386 28580 2438
rect 28580 2386 28632 2438
rect 28632 2386 28634 2438
rect 28578 2384 28634 2386
rect 29237 2435 29293 2437
rect 28814 2433 28870 2435
rect 28814 2381 28816 2433
rect 28816 2381 28868 2433
rect 28868 2381 28870 2433
rect 28814 2379 28870 2381
rect 28998 2433 29054 2435
rect 28998 2381 29000 2433
rect 29000 2381 29052 2433
rect 29052 2381 29054 2433
rect 29237 2383 29239 2435
rect 29239 2383 29291 2435
rect 29291 2383 29293 2435
rect 29237 2381 29293 2383
rect 28998 2379 29054 2381
rect 29440 2431 29496 2433
rect 29440 2379 29442 2431
rect 29442 2379 29494 2431
rect 29494 2379 29496 2431
rect 29440 2377 29496 2379
rect 29625 2428 29681 2430
rect 29625 2376 29627 2428
rect 29627 2376 29679 2428
rect 29679 2376 29681 2428
rect 29625 2374 29681 2376
rect 29816 2430 29872 2432
rect 29816 2378 29818 2430
rect 29818 2378 29870 2430
rect 29870 2378 29872 2430
rect 29816 2376 29872 2378
rect 30007 2434 30063 2436
rect 30007 2382 30009 2434
rect 30009 2382 30061 2434
rect 30061 2382 30063 2434
rect 30007 2380 30063 2382
rect 30193 2430 30249 2432
rect 30193 2378 30195 2430
rect 30195 2378 30247 2430
rect 30247 2378 30249 2430
rect 30193 2376 30249 2378
rect 25640 1847 25696 1849
rect 25640 1795 25642 1847
rect 25642 1795 25694 1847
rect 25694 1795 25696 1847
rect 25640 1793 25696 1795
rect 25845 1843 25901 1845
rect 25845 1791 25847 1843
rect 25847 1791 25899 1843
rect 25899 1791 25901 1843
rect 25845 1789 25901 1791
rect 26031 1848 26087 1850
rect 26031 1796 26033 1848
rect 26033 1796 26085 1848
rect 26085 1796 26087 1848
rect 26031 1794 26087 1796
rect 26225 1841 26281 1843
rect 26225 1789 26227 1841
rect 26227 1789 26279 1841
rect 26279 1789 26281 1841
rect 26225 1787 26281 1789
rect 26444 1846 26500 1848
rect 26444 1794 26446 1846
rect 26446 1794 26498 1846
rect 26498 1794 26500 1846
rect 26444 1792 26500 1794
rect 26654 1846 26710 1848
rect 26654 1794 26656 1846
rect 26656 1794 26708 1846
rect 26708 1794 26710 1846
rect 26654 1792 26710 1794
rect 26883 1843 26939 1845
rect 26883 1791 26885 1843
rect 26885 1791 26937 1843
rect 26937 1791 26939 1843
rect 26883 1789 26939 1791
rect 27129 1843 27185 1845
rect 27129 1791 27131 1843
rect 27131 1791 27183 1843
rect 27183 1791 27185 1843
rect 27129 1789 27185 1791
rect 27403 1843 27459 1845
rect 27403 1791 27405 1843
rect 27405 1791 27457 1843
rect 27457 1791 27459 1843
rect 27403 1789 27459 1791
rect 27678 1843 27734 1845
rect 27678 1791 27680 1843
rect 27680 1791 27732 1843
rect 27732 1791 27734 1843
rect 27678 1789 27734 1791
rect 27914 1843 27970 1845
rect 27914 1791 27916 1843
rect 27916 1791 27968 1843
rect 27968 1791 27970 1843
rect 27914 1789 27970 1791
rect 28137 1846 28193 1848
rect 28137 1794 28139 1846
rect 28139 1794 28191 1846
rect 28191 1794 28193 1846
rect 28137 1792 28193 1794
rect 28355 1849 28411 1851
rect 28355 1797 28357 1849
rect 28357 1797 28409 1849
rect 28409 1797 28411 1849
rect 28355 1795 28411 1797
rect 28533 1840 28589 1842
rect 28533 1788 28535 1840
rect 28535 1788 28587 1840
rect 28587 1788 28589 1840
rect 28533 1786 28589 1788
rect 28772 1842 28828 1844
rect 28772 1790 28774 1842
rect 28774 1790 28826 1842
rect 28826 1790 28828 1842
rect 28772 1788 28828 1790
rect 28969 1842 29025 1844
rect 28969 1790 28971 1842
rect 28971 1790 29023 1842
rect 29023 1790 29025 1842
rect 28969 1788 29025 1790
rect 29167 1842 29223 1844
rect 29167 1790 29169 1842
rect 29169 1790 29221 1842
rect 29221 1790 29223 1842
rect 29167 1788 29223 1790
rect 29380 1843 29436 1845
rect 29380 1791 29382 1843
rect 29382 1791 29434 1843
rect 29434 1791 29436 1843
rect 29380 1789 29436 1791
rect 29603 1842 29659 1844
rect 29603 1790 29605 1842
rect 29605 1790 29657 1842
rect 29657 1790 29659 1842
rect 29603 1788 29659 1790
rect 29800 1847 29856 1849
rect 29800 1795 29802 1847
rect 29802 1795 29854 1847
rect 29854 1795 29856 1847
rect 29800 1793 29856 1795
rect 30016 1845 30072 1847
rect 30016 1793 30018 1845
rect 30018 1793 30070 1845
rect 30070 1793 30072 1845
rect 30016 1791 30072 1793
rect 30225 1845 30281 1847
rect 30225 1793 30227 1845
rect 30227 1793 30279 1845
rect 30279 1793 30281 1845
rect 30225 1791 30281 1793
rect 25236 -960 25292 -958
rect 25236 -1012 25238 -960
rect 25238 -1012 25290 -960
rect 25290 -1012 25292 -960
rect 25236 -1014 25292 -1012
rect 25070 -1646 25126 -1644
rect 25070 -1698 25072 -1646
rect 25072 -1698 25124 -1646
rect 25124 -1698 25126 -1646
rect 25070 -1700 25126 -1698
rect 25269 -1649 25325 -1647
rect 25269 -1701 25271 -1649
rect 25271 -1701 25323 -1649
rect 25323 -1701 25325 -1649
rect 25269 -1703 25325 -1701
<< metal3 >>
rect 13919 13632 14045 13642
rect 13919 13568 13950 13632
rect 14014 13624 14045 13632
rect 20628 13632 20754 13642
rect 14675 13625 19589 13627
rect 14014 13622 14615 13624
rect 14014 13568 14047 13622
rect 13919 13559 14047 13568
rect 13943 13558 14047 13559
rect 14111 13558 14127 13622
rect 14191 13558 14207 13622
rect 14271 13558 14287 13622
rect 14351 13558 14367 13622
rect 14431 13558 14447 13622
rect 14511 13558 14615 13622
rect 14675 13561 14779 13625
rect 14843 13561 14859 13625
rect 14923 13561 14939 13625
rect 15003 13561 15019 13625
rect 15083 13561 15099 13625
rect 15163 13561 15179 13625
rect 15243 13561 15385 13625
rect 15449 13561 15465 13625
rect 15529 13561 15545 13625
rect 15609 13561 15625 13625
rect 15689 13561 15705 13625
rect 15769 13561 15785 13625
rect 15849 13561 15991 13625
rect 16055 13561 16071 13625
rect 16135 13561 16151 13625
rect 16215 13561 16231 13625
rect 16295 13561 16311 13625
rect 16375 13561 16391 13625
rect 16455 13561 16597 13625
rect 16661 13561 16677 13625
rect 16741 13561 16757 13625
rect 16821 13561 16837 13625
rect 16901 13561 16917 13625
rect 16981 13561 16997 13625
rect 17061 13561 17203 13625
rect 17267 13561 17283 13625
rect 17347 13561 17363 13625
rect 17427 13561 17443 13625
rect 17507 13561 17523 13625
rect 17587 13561 17603 13625
rect 17667 13561 17809 13625
rect 17873 13561 17889 13625
rect 17953 13561 17969 13625
rect 18033 13561 18049 13625
rect 18113 13561 18129 13625
rect 18193 13561 18209 13625
rect 18273 13561 18415 13625
rect 18479 13561 18495 13625
rect 18559 13561 18575 13625
rect 18639 13561 18655 13625
rect 18719 13561 18735 13625
rect 18799 13561 18815 13625
rect 18879 13561 19021 13625
rect 19085 13561 19101 13625
rect 19165 13561 19181 13625
rect 19245 13561 19261 13625
rect 19325 13561 19341 13625
rect 19405 13561 19421 13625
rect 19485 13561 19589 13625
rect 14675 13559 19589 13561
rect 19728 13570 19854 13580
rect 13943 13556 14615 13558
rect 13943 13402 14009 13492
rect 13943 13338 13944 13402
rect 14008 13338 14009 13402
rect 13943 13322 14009 13338
rect 13943 13258 13944 13322
rect 14008 13258 14009 13322
rect 13943 13242 14009 13258
rect 13943 13178 13944 13242
rect 14008 13178 14009 13242
rect 3031 13157 3157 13167
rect 3031 13093 3062 13157
rect 3126 13149 3157 13157
rect 13943 13162 14009 13178
rect 3787 13150 8701 13152
rect 3126 13147 3727 13149
rect 3126 13093 3159 13147
rect 3031 13084 3159 13093
rect 3055 13083 3159 13084
rect 3223 13083 3239 13147
rect 3303 13083 3319 13147
rect 3383 13083 3399 13147
rect 3463 13083 3479 13147
rect 3543 13083 3559 13147
rect 3623 13083 3727 13147
rect 3787 13086 3891 13150
rect 3955 13086 3971 13150
rect 4035 13086 4051 13150
rect 4115 13086 4131 13150
rect 4195 13086 4211 13150
rect 4275 13086 4291 13150
rect 4355 13086 4497 13150
rect 4561 13086 4577 13150
rect 4641 13086 4657 13150
rect 4721 13086 4737 13150
rect 4801 13086 4817 13150
rect 4881 13086 4897 13150
rect 4961 13086 5103 13150
rect 5167 13086 5183 13150
rect 5247 13086 5263 13150
rect 5327 13086 5343 13150
rect 5407 13086 5423 13150
rect 5487 13086 5503 13150
rect 5567 13086 5709 13150
rect 5773 13086 5789 13150
rect 5853 13086 5869 13150
rect 5933 13086 5949 13150
rect 6013 13086 6029 13150
rect 6093 13086 6109 13150
rect 6173 13086 6315 13150
rect 6379 13086 6395 13150
rect 6459 13086 6475 13150
rect 6539 13086 6555 13150
rect 6619 13086 6635 13150
rect 6699 13086 6715 13150
rect 6779 13086 6921 13150
rect 6985 13086 7001 13150
rect 7065 13086 7081 13150
rect 7145 13086 7161 13150
rect 7225 13086 7241 13150
rect 7305 13086 7321 13150
rect 7385 13086 7527 13150
rect 7591 13086 7607 13150
rect 7671 13086 7687 13150
rect 7751 13086 7767 13150
rect 7831 13086 7847 13150
rect 7911 13086 7927 13150
rect 7991 13086 8133 13150
rect 8197 13086 8213 13150
rect 8277 13086 8293 13150
rect 8357 13086 8373 13150
rect 8437 13086 8453 13150
rect 8517 13086 8533 13150
rect 8597 13086 8701 13150
rect 3787 13084 8701 13086
rect 8840 13095 8966 13105
rect 3055 13081 3727 13083
rect 3055 12927 3121 13017
rect 3055 12863 3056 12927
rect 3120 12863 3121 12927
rect 3055 12847 3121 12863
rect 3055 12783 3056 12847
rect 3120 12783 3121 12847
rect 3055 12767 3121 12783
rect 3055 12703 3056 12767
rect 3120 12703 3121 12767
rect 3055 12687 3121 12703
rect 3055 12623 3056 12687
rect 3120 12623 3121 12687
rect 3055 12607 3121 12623
rect 2430 12566 2548 12567
rect 2679 12566 2823 12567
rect 2430 12552 2823 12566
rect 2430 12488 2445 12552
rect 2509 12551 2720 12552
rect 2509 12488 2576 12551
rect 2430 12487 2576 12488
rect 2640 12488 2720 12551
rect 2784 12488 2823 12552
rect 2640 12487 2823 12488
rect 2430 12471 2823 12487
rect 3055 12543 3056 12607
rect 3120 12543 3121 12607
rect 3055 12527 3121 12543
rect 2535 12470 2679 12471
rect 3055 12463 3056 12527
rect 3120 12463 3121 12527
rect 3055 12447 3121 12463
rect 3055 12383 3056 12447
rect 3120 12383 3121 12447
rect 3055 12367 3121 12383
rect 3055 12303 3056 12367
rect 3120 12303 3121 12367
rect 3055 12287 3121 12303
rect 3055 12223 3056 12287
rect 3120 12223 3121 12287
rect 3055 12207 3121 12223
rect 3055 12143 3056 12207
rect 3120 12143 3121 12207
rect 2570 12021 2662 12022
rect 2456 12006 2829 12021
rect 2456 11942 2463 12006
rect 2527 11942 2583 12006
rect 2647 11942 2726 12006
rect 2790 11942 2829 12006
rect 2456 11925 2829 11942
rect 3055 11989 3121 12143
rect 3181 11989 3241 13021
rect 3301 12051 3361 13081
rect 3421 11989 3481 13021
rect 3541 12051 3601 13081
rect 3661 12927 3727 13017
rect 3661 12863 3662 12927
rect 3726 12863 3727 12927
rect 3661 12847 3727 12863
rect 3661 12783 3662 12847
rect 3726 12783 3727 12847
rect 3661 12767 3727 12783
rect 3661 12703 3662 12767
rect 3726 12703 3727 12767
rect 3661 12687 3727 12703
rect 3661 12623 3662 12687
rect 3726 12623 3727 12687
rect 3661 12607 3727 12623
rect 3661 12543 3662 12607
rect 3726 12543 3727 12607
rect 3661 12527 3727 12543
rect 3661 12463 3662 12527
rect 3726 12463 3727 12527
rect 3661 12447 3727 12463
rect 3661 12383 3662 12447
rect 3726 12383 3727 12447
rect 3661 12367 3727 12383
rect 3661 12303 3662 12367
rect 3726 12303 3727 12367
rect 3661 12287 3727 12303
rect 3661 12223 3662 12287
rect 3726 12223 3727 12287
rect 3661 12207 3727 12223
rect 3661 12143 3662 12207
rect 3726 12143 3727 12207
rect 3661 11989 3727 12143
rect 3055 11987 3727 11989
rect 3055 11923 3159 11987
rect 3223 11923 3239 11987
rect 3303 11923 3319 11987
rect 3383 11923 3399 11987
rect 3463 11923 3479 11987
rect 3543 11964 3559 11987
rect 3543 11923 3548 11964
rect 3623 11923 3727 11987
rect 3787 12930 3853 13020
rect 3787 12866 3788 12930
rect 3852 12866 3853 12930
rect 3787 12850 3853 12866
rect 3787 12786 3788 12850
rect 3852 12786 3853 12850
rect 3787 12770 3853 12786
rect 3787 12706 3788 12770
rect 3852 12706 3853 12770
rect 3787 12690 3853 12706
rect 3787 12626 3788 12690
rect 3852 12626 3853 12690
rect 3787 12610 3853 12626
rect 3787 12546 3788 12610
rect 3852 12546 3853 12610
rect 3787 12530 3853 12546
rect 3787 12466 3788 12530
rect 3852 12466 3853 12530
rect 3787 12450 3853 12466
rect 3787 12386 3788 12450
rect 3852 12386 3853 12450
rect 3787 12370 3853 12386
rect 3787 12306 3788 12370
rect 3852 12306 3853 12370
rect 3787 12290 3853 12306
rect 3787 12226 3788 12290
rect 3852 12226 3853 12290
rect 3787 12210 3853 12226
rect 3787 12146 3788 12210
rect 3852 12146 3853 12210
rect 3787 11992 3853 12146
rect 3913 11992 3973 13024
rect 4033 12054 4093 13084
rect 4153 11992 4213 13024
rect 4273 12054 4333 13084
rect 4393 12930 4459 13020
rect 4393 12866 4394 12930
rect 4458 12866 4459 12930
rect 4393 12850 4459 12866
rect 4393 12786 4394 12850
rect 4458 12786 4459 12850
rect 4393 12770 4459 12786
rect 4393 12706 4394 12770
rect 4458 12706 4459 12770
rect 4393 12690 4459 12706
rect 4393 12626 4394 12690
rect 4458 12626 4459 12690
rect 4393 12610 4459 12626
rect 4393 12546 4394 12610
rect 4458 12546 4459 12610
rect 4393 12530 4459 12546
rect 4393 12466 4394 12530
rect 4458 12466 4459 12530
rect 4393 12450 4459 12466
rect 4393 12386 4394 12450
rect 4458 12386 4459 12450
rect 4393 12370 4459 12386
rect 4393 12306 4394 12370
rect 4458 12306 4459 12370
rect 4393 12290 4459 12306
rect 4393 12226 4394 12290
rect 4458 12226 4459 12290
rect 4393 12210 4459 12226
rect 4393 12146 4394 12210
rect 4458 12146 4459 12210
rect 4393 11992 4459 12146
rect 4519 12054 4579 13084
rect 4639 11992 4699 13024
rect 4759 12054 4819 13084
rect 4879 11992 4939 13024
rect 4999 12930 5065 13020
rect 4999 12866 5000 12930
rect 5064 12866 5065 12930
rect 4999 12850 5065 12866
rect 4999 12786 5000 12850
rect 5064 12786 5065 12850
rect 4999 12770 5065 12786
rect 4999 12706 5000 12770
rect 5064 12706 5065 12770
rect 4999 12690 5065 12706
rect 4999 12626 5000 12690
rect 5064 12626 5065 12690
rect 4999 12610 5065 12626
rect 4999 12546 5000 12610
rect 5064 12546 5065 12610
rect 4999 12530 5065 12546
rect 4999 12466 5000 12530
rect 5064 12466 5065 12530
rect 4999 12450 5065 12466
rect 4999 12386 5000 12450
rect 5064 12386 5065 12450
rect 4999 12370 5065 12386
rect 4999 12306 5000 12370
rect 5064 12306 5065 12370
rect 4999 12290 5065 12306
rect 4999 12226 5000 12290
rect 5064 12226 5065 12290
rect 4999 12210 5065 12226
rect 4999 12146 5000 12210
rect 5064 12146 5065 12210
rect 4999 11992 5065 12146
rect 5125 11992 5185 13024
rect 5245 12054 5305 13084
rect 5365 11992 5425 13024
rect 5485 12054 5545 13084
rect 5605 12930 5671 13020
rect 5605 12866 5606 12930
rect 5670 12866 5671 12930
rect 5605 12850 5671 12866
rect 5605 12786 5606 12850
rect 5670 12786 5671 12850
rect 5605 12770 5671 12786
rect 5605 12706 5606 12770
rect 5670 12706 5671 12770
rect 5605 12690 5671 12706
rect 5605 12626 5606 12690
rect 5670 12626 5671 12690
rect 5605 12610 5671 12626
rect 5605 12546 5606 12610
rect 5670 12546 5671 12610
rect 5605 12530 5671 12546
rect 5605 12466 5606 12530
rect 5670 12466 5671 12530
rect 5605 12450 5671 12466
rect 5605 12386 5606 12450
rect 5670 12386 5671 12450
rect 5605 12370 5671 12386
rect 5605 12306 5606 12370
rect 5670 12306 5671 12370
rect 5605 12290 5671 12306
rect 5605 12226 5606 12290
rect 5670 12226 5671 12290
rect 5605 12210 5671 12226
rect 5605 12146 5606 12210
rect 5670 12146 5671 12210
rect 5605 11992 5671 12146
rect 5731 12054 5791 13084
rect 5851 11992 5911 13024
rect 5971 12054 6031 13084
rect 6091 11992 6151 13024
rect 6211 12930 6277 13020
rect 6211 12866 6212 12930
rect 6276 12866 6277 12930
rect 6211 12850 6277 12866
rect 6211 12786 6212 12850
rect 6276 12786 6277 12850
rect 6211 12770 6277 12786
rect 6211 12706 6212 12770
rect 6276 12706 6277 12770
rect 6211 12690 6277 12706
rect 6211 12626 6212 12690
rect 6276 12626 6277 12690
rect 6211 12610 6277 12626
rect 6211 12546 6212 12610
rect 6276 12546 6277 12610
rect 6211 12530 6277 12546
rect 6211 12466 6212 12530
rect 6276 12466 6277 12530
rect 6211 12450 6277 12466
rect 6211 12386 6212 12450
rect 6276 12386 6277 12450
rect 6211 12370 6277 12386
rect 6211 12306 6212 12370
rect 6276 12306 6277 12370
rect 6211 12290 6277 12306
rect 6211 12226 6212 12290
rect 6276 12226 6277 12290
rect 6211 12210 6277 12226
rect 6211 12146 6212 12210
rect 6276 12146 6277 12210
rect 6211 11992 6277 12146
rect 6337 11992 6397 13024
rect 6457 12054 6517 13084
rect 6577 11992 6637 13024
rect 6697 12054 6757 13084
rect 6817 12930 6883 13020
rect 6817 12866 6818 12930
rect 6882 12866 6883 12930
rect 6817 12850 6883 12866
rect 6817 12786 6818 12850
rect 6882 12786 6883 12850
rect 6817 12770 6883 12786
rect 6817 12706 6818 12770
rect 6882 12706 6883 12770
rect 6817 12690 6883 12706
rect 6817 12626 6818 12690
rect 6882 12626 6883 12690
rect 6817 12610 6883 12626
rect 6817 12546 6818 12610
rect 6882 12546 6883 12610
rect 6817 12530 6883 12546
rect 6817 12466 6818 12530
rect 6882 12466 6883 12530
rect 6817 12450 6883 12466
rect 6817 12386 6818 12450
rect 6882 12386 6883 12450
rect 6817 12370 6883 12386
rect 6817 12306 6818 12370
rect 6882 12306 6883 12370
rect 6817 12290 6883 12306
rect 6817 12226 6818 12290
rect 6882 12226 6883 12290
rect 6817 12210 6883 12226
rect 6817 12146 6818 12210
rect 6882 12146 6883 12210
rect 6817 11992 6883 12146
rect 6943 12054 7003 13084
rect 7063 11992 7123 13024
rect 7183 12054 7243 13084
rect 7303 11992 7363 13024
rect 7423 12930 7489 13020
rect 7423 12866 7424 12930
rect 7488 12866 7489 12930
rect 7423 12850 7489 12866
rect 7423 12786 7424 12850
rect 7488 12786 7489 12850
rect 7423 12770 7489 12786
rect 7423 12706 7424 12770
rect 7488 12706 7489 12770
rect 7423 12690 7489 12706
rect 7423 12626 7424 12690
rect 7488 12626 7489 12690
rect 7423 12610 7489 12626
rect 7423 12546 7424 12610
rect 7488 12546 7489 12610
rect 7423 12530 7489 12546
rect 7423 12466 7424 12530
rect 7488 12466 7489 12530
rect 7423 12450 7489 12466
rect 7423 12386 7424 12450
rect 7488 12386 7489 12450
rect 7423 12370 7489 12386
rect 7423 12306 7424 12370
rect 7488 12306 7489 12370
rect 7423 12290 7489 12306
rect 7423 12226 7424 12290
rect 7488 12226 7489 12290
rect 7423 12210 7489 12226
rect 7423 12146 7424 12210
rect 7488 12146 7489 12210
rect 7423 11992 7489 12146
rect 7549 11992 7609 13024
rect 7669 12054 7729 13084
rect 7789 11992 7849 13024
rect 7909 12054 7969 13084
rect 8029 12930 8095 13020
rect 8029 12866 8030 12930
rect 8094 12866 8095 12930
rect 8029 12850 8095 12866
rect 8029 12786 8030 12850
rect 8094 12786 8095 12850
rect 8029 12770 8095 12786
rect 8029 12706 8030 12770
rect 8094 12706 8095 12770
rect 8029 12690 8095 12706
rect 8029 12626 8030 12690
rect 8094 12626 8095 12690
rect 8029 12610 8095 12626
rect 8029 12546 8030 12610
rect 8094 12546 8095 12610
rect 8029 12530 8095 12546
rect 8029 12466 8030 12530
rect 8094 12466 8095 12530
rect 8029 12450 8095 12466
rect 8029 12386 8030 12450
rect 8094 12386 8095 12450
rect 8029 12370 8095 12386
rect 8029 12306 8030 12370
rect 8094 12306 8095 12370
rect 8029 12290 8095 12306
rect 8029 12226 8030 12290
rect 8094 12226 8095 12290
rect 8029 12210 8095 12226
rect 8029 12146 8030 12210
rect 8094 12146 8095 12210
rect 8029 11992 8095 12146
rect 8155 12054 8215 13084
rect 8275 11992 8335 13024
rect 8395 12054 8455 13084
rect 8840 13031 8871 13095
rect 8935 13031 8966 13095
rect 13943 13098 13944 13162
rect 14008 13098 14009 13162
rect 13943 13082 14009 13098
rect 8515 11992 8575 13024
rect 8840 13021 8966 13031
rect 13318 13041 13436 13042
rect 13567 13041 13711 13042
rect 13318 13027 13711 13041
rect 8635 12930 8701 13020
rect 13318 12963 13333 13027
rect 13397 13026 13608 13027
rect 13397 12963 13464 13026
rect 13318 12962 13464 12963
rect 13528 12963 13608 13026
rect 13672 12963 13711 13027
rect 13528 12962 13711 12963
rect 8635 12866 8636 12930
rect 8700 12866 8701 12930
rect 8845 12951 8971 12961
rect 8845 12887 8876 12951
rect 8940 12887 8971 12951
rect 13318 12946 13711 12962
rect 13943 13018 13944 13082
rect 14008 13018 14009 13082
rect 13943 13002 14009 13018
rect 13423 12945 13567 12946
rect 8845 12877 8971 12887
rect 13943 12938 13944 13002
rect 14008 12938 14009 13002
rect 13943 12922 14009 12938
rect 8635 12850 8701 12866
rect 8635 12786 8636 12850
rect 8700 12786 8701 12850
rect 13943 12858 13944 12922
rect 14008 12858 14009 12922
rect 13943 12842 14009 12858
rect 8635 12770 8701 12786
rect 8635 12706 8636 12770
rect 8700 12706 8701 12770
rect 8846 12799 8972 12809
rect 8846 12735 8877 12799
rect 8941 12735 8972 12799
rect 8846 12725 8972 12735
rect 13943 12778 13944 12842
rect 14008 12778 14009 12842
rect 13943 12762 14009 12778
rect 8635 12690 8701 12706
rect 8635 12626 8636 12690
rect 8700 12626 8701 12690
rect 13943 12698 13944 12762
rect 14008 12698 14009 12762
rect 13943 12682 14009 12698
rect 8635 12610 8701 12626
rect 8635 12546 8636 12610
rect 8700 12546 8701 12610
rect 8846 12629 8972 12639
rect 8846 12565 8877 12629
rect 8941 12565 8972 12629
rect 13943 12618 13944 12682
rect 14008 12618 14009 12682
rect 8846 12555 8972 12565
rect 10951 12560 11076 12570
rect 8635 12530 8701 12546
rect 8635 12466 8636 12530
rect 8700 12466 8701 12530
rect 10951 12496 10981 12560
rect 11045 12496 11076 12560
rect 10951 12486 11076 12496
rect 11138 12562 11263 12572
rect 11138 12498 11168 12562
rect 11232 12498 11263 12562
rect 11138 12488 11263 12498
rect 11323 12564 11448 12574
rect 11323 12500 11353 12564
rect 11417 12500 11448 12564
rect 11323 12490 11448 12500
rect 11508 12565 11633 12575
rect 11508 12501 11538 12565
rect 11602 12501 11633 12565
rect 11508 12491 11633 12501
rect 11711 12567 11836 12577
rect 11711 12503 11741 12567
rect 11805 12503 11836 12567
rect 11711 12493 11836 12503
rect 11896 12569 12021 12579
rect 11896 12505 11926 12569
rect 11990 12505 12021 12569
rect 11896 12495 12021 12505
rect 12095 12571 12220 12581
rect 12095 12507 12125 12571
rect 12189 12507 12220 12571
rect 12095 12497 12220 12507
rect 12297 12570 12422 12580
rect 12297 12506 12327 12570
rect 12391 12506 12422 12570
rect 12297 12496 12422 12506
rect 12507 12573 12632 12583
rect 12507 12509 12537 12573
rect 12601 12509 12632 12573
rect 12507 12499 12632 12509
rect 12731 12573 12856 12583
rect 12731 12509 12761 12573
rect 12825 12509 12856 12573
rect 12731 12499 12856 12509
rect 12937 12572 13062 12582
rect 12937 12508 12967 12572
rect 13031 12508 13062 12572
rect 12937 12498 13062 12508
rect 13158 12571 13283 12581
rect 13158 12507 13188 12571
rect 13252 12507 13283 12571
rect 13158 12497 13283 12507
rect 13458 12496 13550 12497
rect 8635 12450 8701 12466
rect 8635 12386 8636 12450
rect 8700 12386 8701 12450
rect 8845 12472 8971 12482
rect 8845 12408 8876 12472
rect 8940 12408 8971 12472
rect 8845 12398 8971 12408
rect 13344 12481 13717 12496
rect 13344 12417 13351 12481
rect 13415 12417 13471 12481
rect 13535 12417 13614 12481
rect 13678 12417 13717 12481
rect 13344 12400 13717 12417
rect 13943 12464 14009 12618
rect 14069 12464 14129 13496
rect 14189 12526 14249 13556
rect 14309 12464 14369 13496
rect 14429 12526 14489 13556
rect 14549 13402 14615 13492
rect 14549 13338 14550 13402
rect 14614 13338 14615 13402
rect 14549 13322 14615 13338
rect 14549 13258 14550 13322
rect 14614 13258 14615 13322
rect 14549 13242 14615 13258
rect 14549 13178 14550 13242
rect 14614 13178 14615 13242
rect 14549 13162 14615 13178
rect 14549 13098 14550 13162
rect 14614 13098 14615 13162
rect 14549 13082 14615 13098
rect 14549 13018 14550 13082
rect 14614 13018 14615 13082
rect 14549 13002 14615 13018
rect 14549 12938 14550 13002
rect 14614 12938 14615 13002
rect 14549 12922 14615 12938
rect 14549 12858 14550 12922
rect 14614 12858 14615 12922
rect 14549 12842 14615 12858
rect 14549 12778 14550 12842
rect 14614 12778 14615 12842
rect 14549 12762 14615 12778
rect 14549 12698 14550 12762
rect 14614 12698 14615 12762
rect 14549 12682 14615 12698
rect 14549 12618 14550 12682
rect 14614 12618 14615 12682
rect 14549 12464 14615 12618
rect 13943 12462 14615 12464
rect 13943 12398 14047 12462
rect 14111 12398 14127 12462
rect 14191 12398 14207 12462
rect 14271 12398 14287 12462
rect 14351 12398 14367 12462
rect 14431 12439 14447 12462
rect 14431 12398 14436 12439
rect 14511 12398 14615 12462
rect 14675 13405 14741 13495
rect 14675 13341 14676 13405
rect 14740 13341 14741 13405
rect 14675 13325 14741 13341
rect 14675 13261 14676 13325
rect 14740 13261 14741 13325
rect 14675 13245 14741 13261
rect 14675 13181 14676 13245
rect 14740 13181 14741 13245
rect 14675 13165 14741 13181
rect 14675 13101 14676 13165
rect 14740 13101 14741 13165
rect 14675 13085 14741 13101
rect 14675 13021 14676 13085
rect 14740 13021 14741 13085
rect 14675 13005 14741 13021
rect 14675 12941 14676 13005
rect 14740 12941 14741 13005
rect 14675 12925 14741 12941
rect 14675 12861 14676 12925
rect 14740 12861 14741 12925
rect 14675 12845 14741 12861
rect 14675 12781 14676 12845
rect 14740 12781 14741 12845
rect 14675 12765 14741 12781
rect 14675 12701 14676 12765
rect 14740 12701 14741 12765
rect 14675 12685 14741 12701
rect 14675 12621 14676 12685
rect 14740 12621 14741 12685
rect 14675 12467 14741 12621
rect 14801 12467 14861 13499
rect 14921 12529 14981 13559
rect 15041 12467 15101 13499
rect 15161 12529 15221 13559
rect 15281 13405 15347 13495
rect 15281 13341 15282 13405
rect 15346 13341 15347 13405
rect 15281 13325 15347 13341
rect 15281 13261 15282 13325
rect 15346 13261 15347 13325
rect 15281 13245 15347 13261
rect 15281 13181 15282 13245
rect 15346 13181 15347 13245
rect 15281 13165 15347 13181
rect 15281 13101 15282 13165
rect 15346 13101 15347 13165
rect 15281 13085 15347 13101
rect 15281 13021 15282 13085
rect 15346 13021 15347 13085
rect 15281 13005 15347 13021
rect 15281 12941 15282 13005
rect 15346 12941 15347 13005
rect 15281 12925 15347 12941
rect 15281 12861 15282 12925
rect 15346 12861 15347 12925
rect 15281 12845 15347 12861
rect 15281 12781 15282 12845
rect 15346 12781 15347 12845
rect 15281 12765 15347 12781
rect 15281 12701 15282 12765
rect 15346 12701 15347 12765
rect 15281 12685 15347 12701
rect 15281 12621 15282 12685
rect 15346 12621 15347 12685
rect 15281 12467 15347 12621
rect 15407 12529 15467 13559
rect 15527 12467 15587 13499
rect 15647 12529 15707 13559
rect 15767 12467 15827 13499
rect 15887 13405 15953 13495
rect 15887 13341 15888 13405
rect 15952 13341 15953 13405
rect 15887 13325 15953 13341
rect 15887 13261 15888 13325
rect 15952 13261 15953 13325
rect 15887 13245 15953 13261
rect 15887 13181 15888 13245
rect 15952 13181 15953 13245
rect 15887 13165 15953 13181
rect 15887 13101 15888 13165
rect 15952 13101 15953 13165
rect 15887 13085 15953 13101
rect 15887 13021 15888 13085
rect 15952 13021 15953 13085
rect 15887 13005 15953 13021
rect 15887 12941 15888 13005
rect 15952 12941 15953 13005
rect 15887 12925 15953 12941
rect 15887 12861 15888 12925
rect 15952 12861 15953 12925
rect 15887 12845 15953 12861
rect 15887 12781 15888 12845
rect 15952 12781 15953 12845
rect 15887 12765 15953 12781
rect 15887 12701 15888 12765
rect 15952 12701 15953 12765
rect 15887 12685 15953 12701
rect 15887 12621 15888 12685
rect 15952 12621 15953 12685
rect 15887 12467 15953 12621
rect 16013 12467 16073 13499
rect 16133 12529 16193 13559
rect 16253 12467 16313 13499
rect 16373 12529 16433 13559
rect 16493 13405 16559 13495
rect 16493 13341 16494 13405
rect 16558 13341 16559 13405
rect 16493 13325 16559 13341
rect 16493 13261 16494 13325
rect 16558 13261 16559 13325
rect 16493 13245 16559 13261
rect 16493 13181 16494 13245
rect 16558 13181 16559 13245
rect 16493 13165 16559 13181
rect 16493 13101 16494 13165
rect 16558 13101 16559 13165
rect 16493 13085 16559 13101
rect 16493 13021 16494 13085
rect 16558 13021 16559 13085
rect 16493 13005 16559 13021
rect 16493 12941 16494 13005
rect 16558 12941 16559 13005
rect 16493 12925 16559 12941
rect 16493 12861 16494 12925
rect 16558 12861 16559 12925
rect 16493 12845 16559 12861
rect 16493 12781 16494 12845
rect 16558 12781 16559 12845
rect 16493 12765 16559 12781
rect 16493 12701 16494 12765
rect 16558 12701 16559 12765
rect 16493 12685 16559 12701
rect 16493 12621 16494 12685
rect 16558 12621 16559 12685
rect 16493 12467 16559 12621
rect 16619 12529 16679 13559
rect 16739 12467 16799 13499
rect 16859 12529 16919 13559
rect 16979 12467 17039 13499
rect 17099 13405 17165 13495
rect 17099 13341 17100 13405
rect 17164 13341 17165 13405
rect 17099 13325 17165 13341
rect 17099 13261 17100 13325
rect 17164 13261 17165 13325
rect 17099 13245 17165 13261
rect 17099 13181 17100 13245
rect 17164 13181 17165 13245
rect 17099 13165 17165 13181
rect 17099 13101 17100 13165
rect 17164 13101 17165 13165
rect 17099 13085 17165 13101
rect 17099 13021 17100 13085
rect 17164 13021 17165 13085
rect 17099 13005 17165 13021
rect 17099 12941 17100 13005
rect 17164 12941 17165 13005
rect 17099 12925 17165 12941
rect 17099 12861 17100 12925
rect 17164 12861 17165 12925
rect 17099 12845 17165 12861
rect 17099 12781 17100 12845
rect 17164 12781 17165 12845
rect 17099 12765 17165 12781
rect 17099 12701 17100 12765
rect 17164 12701 17165 12765
rect 17099 12685 17165 12701
rect 17099 12621 17100 12685
rect 17164 12621 17165 12685
rect 17099 12467 17165 12621
rect 17225 12467 17285 13499
rect 17345 12529 17405 13559
rect 17465 12467 17525 13499
rect 17585 12529 17645 13559
rect 17705 13405 17771 13495
rect 17705 13341 17706 13405
rect 17770 13341 17771 13405
rect 17705 13325 17771 13341
rect 17705 13261 17706 13325
rect 17770 13261 17771 13325
rect 17705 13245 17771 13261
rect 17705 13181 17706 13245
rect 17770 13181 17771 13245
rect 17705 13165 17771 13181
rect 17705 13101 17706 13165
rect 17770 13101 17771 13165
rect 17705 13085 17771 13101
rect 17705 13021 17706 13085
rect 17770 13021 17771 13085
rect 17705 13005 17771 13021
rect 17705 12941 17706 13005
rect 17770 12941 17771 13005
rect 17705 12925 17771 12941
rect 17705 12861 17706 12925
rect 17770 12861 17771 12925
rect 17705 12845 17771 12861
rect 17705 12781 17706 12845
rect 17770 12781 17771 12845
rect 17705 12765 17771 12781
rect 17705 12701 17706 12765
rect 17770 12701 17771 12765
rect 17705 12685 17771 12701
rect 17705 12621 17706 12685
rect 17770 12621 17771 12685
rect 17705 12467 17771 12621
rect 17831 12529 17891 13559
rect 17951 12467 18011 13499
rect 18071 12529 18131 13559
rect 18191 12467 18251 13499
rect 18311 13405 18377 13495
rect 18311 13341 18312 13405
rect 18376 13341 18377 13405
rect 18311 13325 18377 13341
rect 18311 13261 18312 13325
rect 18376 13261 18377 13325
rect 18311 13245 18377 13261
rect 18311 13181 18312 13245
rect 18376 13181 18377 13245
rect 18311 13165 18377 13181
rect 18311 13101 18312 13165
rect 18376 13101 18377 13165
rect 18311 13085 18377 13101
rect 18311 13021 18312 13085
rect 18376 13021 18377 13085
rect 18311 13005 18377 13021
rect 18311 12941 18312 13005
rect 18376 12941 18377 13005
rect 18311 12925 18377 12941
rect 18311 12861 18312 12925
rect 18376 12861 18377 12925
rect 18311 12845 18377 12861
rect 18311 12781 18312 12845
rect 18376 12781 18377 12845
rect 18311 12765 18377 12781
rect 18311 12701 18312 12765
rect 18376 12701 18377 12765
rect 18311 12685 18377 12701
rect 18311 12621 18312 12685
rect 18376 12621 18377 12685
rect 18311 12467 18377 12621
rect 18437 12467 18497 13499
rect 18557 12529 18617 13559
rect 18677 12467 18737 13499
rect 18797 12529 18857 13559
rect 18917 13405 18983 13495
rect 18917 13341 18918 13405
rect 18982 13341 18983 13405
rect 18917 13325 18983 13341
rect 18917 13261 18918 13325
rect 18982 13261 18983 13325
rect 18917 13245 18983 13261
rect 18917 13181 18918 13245
rect 18982 13181 18983 13245
rect 18917 13165 18983 13181
rect 18917 13101 18918 13165
rect 18982 13101 18983 13165
rect 18917 13085 18983 13101
rect 18917 13021 18918 13085
rect 18982 13021 18983 13085
rect 18917 13005 18983 13021
rect 18917 12941 18918 13005
rect 18982 12941 18983 13005
rect 18917 12925 18983 12941
rect 18917 12861 18918 12925
rect 18982 12861 18983 12925
rect 18917 12845 18983 12861
rect 18917 12781 18918 12845
rect 18982 12781 18983 12845
rect 18917 12765 18983 12781
rect 18917 12701 18918 12765
rect 18982 12701 18983 12765
rect 18917 12685 18983 12701
rect 18917 12621 18918 12685
rect 18982 12621 18983 12685
rect 18917 12467 18983 12621
rect 19043 12529 19103 13559
rect 19163 12467 19223 13499
rect 19283 12529 19343 13559
rect 19728 13506 19759 13570
rect 19823 13506 19854 13570
rect 19403 12467 19463 13499
rect 19728 13496 19854 13506
rect 20205 13573 20331 13583
rect 20205 13509 20236 13573
rect 20300 13509 20331 13573
rect 20628 13568 20659 13632
rect 20723 13624 20754 13632
rect 21384 13625 26298 13627
rect 20723 13622 21324 13624
rect 20723 13568 20756 13622
rect 20628 13559 20756 13568
rect 20652 13558 20756 13559
rect 20820 13558 20836 13622
rect 20900 13558 20916 13622
rect 20980 13558 20996 13622
rect 21060 13558 21076 13622
rect 21140 13558 21156 13622
rect 21220 13558 21324 13622
rect 21384 13561 21488 13625
rect 21552 13561 21568 13625
rect 21632 13561 21648 13625
rect 21712 13561 21728 13625
rect 21792 13561 21808 13625
rect 21872 13561 21888 13625
rect 21952 13561 22094 13625
rect 22158 13561 22174 13625
rect 22238 13561 22254 13625
rect 22318 13561 22334 13625
rect 22398 13561 22414 13625
rect 22478 13561 22494 13625
rect 22558 13561 22700 13625
rect 22764 13561 22780 13625
rect 22844 13561 22860 13625
rect 22924 13561 22940 13625
rect 23004 13561 23020 13625
rect 23084 13561 23100 13625
rect 23164 13561 23306 13625
rect 23370 13561 23386 13625
rect 23450 13561 23466 13625
rect 23530 13561 23546 13625
rect 23610 13561 23626 13625
rect 23690 13561 23706 13625
rect 23770 13561 23912 13625
rect 23976 13561 23992 13625
rect 24056 13561 24072 13625
rect 24136 13561 24152 13625
rect 24216 13561 24232 13625
rect 24296 13561 24312 13625
rect 24376 13561 24518 13625
rect 24582 13561 24598 13625
rect 24662 13561 24678 13625
rect 24742 13561 24758 13625
rect 24822 13561 24838 13625
rect 24902 13561 24918 13625
rect 24982 13561 25124 13625
rect 25188 13561 25204 13625
rect 25268 13561 25284 13625
rect 25348 13561 25364 13625
rect 25428 13561 25444 13625
rect 25508 13561 25524 13625
rect 25588 13561 25730 13625
rect 25794 13561 25810 13625
rect 25874 13561 25890 13625
rect 25954 13561 25970 13625
rect 26034 13561 26050 13625
rect 26114 13561 26130 13625
rect 26194 13561 26298 13625
rect 21384 13559 26298 13561
rect 26437 13570 26563 13580
rect 20652 13556 21324 13558
rect 20205 13499 20331 13509
rect 19523 13405 19589 13495
rect 19523 13341 19524 13405
rect 19588 13341 19589 13405
rect 19733 13426 19859 13436
rect 19733 13362 19764 13426
rect 19828 13362 19859 13426
rect 19733 13352 19859 13362
rect 20194 13401 20320 13411
rect 19523 13325 19589 13341
rect 20194 13337 20225 13401
rect 20289 13337 20320 13401
rect 20194 13327 20320 13337
rect 20652 13402 20718 13492
rect 20652 13338 20653 13402
rect 20717 13338 20718 13402
rect 19523 13261 19524 13325
rect 19588 13261 19589 13325
rect 20652 13322 20718 13338
rect 19523 13245 19589 13261
rect 19523 13181 19524 13245
rect 19588 13181 19589 13245
rect 19734 13274 19860 13284
rect 19734 13210 19765 13274
rect 19829 13210 19860 13274
rect 20652 13258 20653 13322
rect 20717 13258 20718 13322
rect 20652 13242 20718 13258
rect 19734 13200 19860 13210
rect 20194 13209 20320 13219
rect 19523 13165 19589 13181
rect 19523 13101 19524 13165
rect 19588 13101 19589 13165
rect 20194 13145 20225 13209
rect 20289 13145 20320 13209
rect 20194 13135 20320 13145
rect 20652 13178 20653 13242
rect 20717 13178 20718 13242
rect 20652 13162 20718 13178
rect 19523 13085 19589 13101
rect 19523 13021 19524 13085
rect 19588 13021 19589 13085
rect 19734 13104 19860 13114
rect 19734 13040 19765 13104
rect 19829 13040 19860 13104
rect 20652 13098 20653 13162
rect 20717 13098 20718 13162
rect 20652 13082 20718 13098
rect 19734 13030 19860 13040
rect 20027 13041 20145 13042
rect 20276 13041 20420 13042
rect 19523 13005 19589 13021
rect 19523 12941 19524 13005
rect 19588 12941 19589 13005
rect 20027 13027 20420 13041
rect 20027 12963 20042 13027
rect 20106 13026 20317 13027
rect 20106 12963 20173 13026
rect 20027 12962 20173 12963
rect 20237 12963 20317 13026
rect 20381 12963 20420 13027
rect 20237 12962 20420 12963
rect 19523 12925 19589 12941
rect 19523 12861 19524 12925
rect 19588 12861 19589 12925
rect 19733 12947 19859 12957
rect 19733 12883 19764 12947
rect 19828 12883 19859 12947
rect 20027 12946 20420 12962
rect 20652 13018 20653 13082
rect 20717 13018 20718 13082
rect 20652 13002 20718 13018
rect 20132 12945 20276 12946
rect 19733 12873 19859 12883
rect 20652 12938 20653 13002
rect 20717 12938 20718 13002
rect 20652 12922 20718 12938
rect 19523 12845 19589 12861
rect 19523 12781 19524 12845
rect 19588 12781 19589 12845
rect 19523 12765 19589 12781
rect 19523 12701 19524 12765
rect 19588 12701 19589 12765
rect 20652 12858 20653 12922
rect 20717 12858 20718 12922
rect 20652 12842 20718 12858
rect 20652 12778 20653 12842
rect 20717 12778 20718 12842
rect 20652 12762 20718 12778
rect 19523 12685 19589 12701
rect 19523 12621 19524 12685
rect 19588 12621 19589 12685
rect 19651 12705 19777 12715
rect 19651 12641 19682 12705
rect 19746 12641 19777 12705
rect 19651 12631 19777 12641
rect 20652 12698 20653 12762
rect 20717 12698 20718 12762
rect 20652 12682 20718 12698
rect 19523 12467 19589 12621
rect 20652 12618 20653 12682
rect 20717 12618 20718 12682
rect 20167 12496 20259 12497
rect 14675 12465 19589 12467
rect 14675 12401 14779 12465
rect 14843 12401 14859 12465
rect 14923 12401 14939 12465
rect 15003 12401 15019 12465
rect 15083 12401 15099 12465
rect 15163 12442 15179 12465
rect 15163 12401 15168 12442
rect 15243 12401 15385 12465
rect 15449 12442 15465 12465
rect 15460 12401 15465 12442
rect 15529 12401 15545 12465
rect 15609 12401 15625 12465
rect 15689 12401 15705 12465
rect 15769 12401 15785 12465
rect 15849 12401 15991 12465
rect 16055 12401 16071 12465
rect 16135 12401 16151 12465
rect 16215 12401 16231 12465
rect 16295 12401 16311 12465
rect 16375 12442 16391 12465
rect 16375 12401 16380 12442
rect 16455 12401 16597 12465
rect 16661 12442 16677 12465
rect 16672 12401 16677 12442
rect 16741 12401 16757 12465
rect 16821 12401 16837 12465
rect 16901 12401 16917 12465
rect 16981 12401 16997 12465
rect 17061 12401 17203 12465
rect 17267 12401 17283 12465
rect 17347 12401 17363 12465
rect 17427 12401 17443 12465
rect 17507 12401 17523 12465
rect 17587 12442 17603 12465
rect 17587 12401 17592 12442
rect 17667 12401 17809 12465
rect 17873 12442 17889 12465
rect 17884 12401 17889 12442
rect 17953 12401 17969 12465
rect 18033 12401 18049 12465
rect 18113 12401 18129 12465
rect 18193 12401 18209 12465
rect 18273 12401 18415 12465
rect 18479 12401 18495 12465
rect 18559 12401 18575 12465
rect 18639 12401 18655 12465
rect 18719 12401 18735 12465
rect 18799 12442 18815 12465
rect 18799 12401 18804 12442
rect 18879 12401 19021 12465
rect 19085 12442 19101 12465
rect 19096 12401 19101 12442
rect 19165 12401 19181 12465
rect 19245 12401 19261 12465
rect 19325 12401 19341 12465
rect 19405 12401 19421 12465
rect 19485 12401 19589 12465
rect 20053 12481 20426 12496
rect 14675 12399 15168 12401
rect 13943 12396 14436 12398
rect 8635 12370 8701 12386
rect 14426 12375 14436 12396
rect 14500 12396 14615 12398
rect 14500 12375 14509 12396
rect 14426 12370 14509 12375
rect 15158 12378 15168 12399
rect 15232 12399 15396 12401
rect 15232 12378 15241 12399
rect 15158 12373 15241 12378
rect 15387 12378 15396 12399
rect 15460 12399 16380 12401
rect 15460 12378 15470 12399
rect 15387 12373 15470 12378
rect 16370 12378 16380 12399
rect 16444 12399 16608 12401
rect 16444 12378 16453 12399
rect 16370 12373 16453 12378
rect 16599 12378 16608 12399
rect 16672 12399 17592 12401
rect 16672 12378 16682 12399
rect 16599 12373 16682 12378
rect 17582 12378 17592 12399
rect 17656 12399 17820 12401
rect 17656 12378 17665 12399
rect 17582 12373 17665 12378
rect 17811 12378 17820 12399
rect 17884 12399 18804 12401
rect 17884 12378 17894 12399
rect 17811 12373 17894 12378
rect 18794 12378 18804 12399
rect 18868 12399 19032 12401
rect 18868 12378 18877 12399
rect 18794 12373 18877 12378
rect 19023 12378 19032 12399
rect 19096 12399 19589 12401
rect 19739 12444 19865 12454
rect 19096 12378 19106 12399
rect 19023 12373 19106 12378
rect 19739 12380 19770 12444
rect 19834 12380 19865 12444
rect 20053 12417 20060 12481
rect 20124 12417 20180 12481
rect 20244 12417 20323 12481
rect 20387 12417 20426 12481
rect 20053 12400 20426 12417
rect 20652 12464 20718 12618
rect 20778 12464 20838 13496
rect 20898 12526 20958 13556
rect 21018 12464 21078 13496
rect 21138 12526 21198 13556
rect 21258 13402 21324 13492
rect 21258 13338 21259 13402
rect 21323 13338 21324 13402
rect 21258 13322 21324 13338
rect 21258 13258 21259 13322
rect 21323 13258 21324 13322
rect 21258 13242 21324 13258
rect 21258 13178 21259 13242
rect 21323 13178 21324 13242
rect 21258 13162 21324 13178
rect 21258 13098 21259 13162
rect 21323 13098 21324 13162
rect 21258 13082 21324 13098
rect 21258 13018 21259 13082
rect 21323 13018 21324 13082
rect 21258 13002 21324 13018
rect 21258 12938 21259 13002
rect 21323 12938 21324 13002
rect 21258 12922 21324 12938
rect 21258 12858 21259 12922
rect 21323 12858 21324 12922
rect 21258 12842 21324 12858
rect 21258 12778 21259 12842
rect 21323 12778 21324 12842
rect 21258 12762 21324 12778
rect 21258 12698 21259 12762
rect 21323 12698 21324 12762
rect 21258 12682 21324 12698
rect 21258 12618 21259 12682
rect 21323 12618 21324 12682
rect 21258 12464 21324 12618
rect 20652 12462 21324 12464
rect 20652 12398 20756 12462
rect 20820 12398 20836 12462
rect 20900 12398 20916 12462
rect 20980 12398 20996 12462
rect 21060 12398 21076 12462
rect 21140 12439 21156 12462
rect 21140 12398 21145 12439
rect 21220 12398 21324 12462
rect 21384 13405 21450 13495
rect 21384 13341 21385 13405
rect 21449 13341 21450 13405
rect 21384 13325 21450 13341
rect 21384 13261 21385 13325
rect 21449 13261 21450 13325
rect 21384 13245 21450 13261
rect 21384 13181 21385 13245
rect 21449 13181 21450 13245
rect 21384 13165 21450 13181
rect 21384 13101 21385 13165
rect 21449 13101 21450 13165
rect 21384 13085 21450 13101
rect 21384 13021 21385 13085
rect 21449 13021 21450 13085
rect 21384 13005 21450 13021
rect 21384 12941 21385 13005
rect 21449 12941 21450 13005
rect 21384 12925 21450 12941
rect 21384 12861 21385 12925
rect 21449 12861 21450 12925
rect 21384 12845 21450 12861
rect 21384 12781 21385 12845
rect 21449 12781 21450 12845
rect 21384 12765 21450 12781
rect 21384 12701 21385 12765
rect 21449 12701 21450 12765
rect 21384 12685 21450 12701
rect 21384 12621 21385 12685
rect 21449 12621 21450 12685
rect 21384 12467 21450 12621
rect 21510 12467 21570 13499
rect 21630 12529 21690 13559
rect 21750 12467 21810 13499
rect 21870 12529 21930 13559
rect 21990 13405 22056 13495
rect 21990 13341 21991 13405
rect 22055 13341 22056 13405
rect 21990 13325 22056 13341
rect 21990 13261 21991 13325
rect 22055 13261 22056 13325
rect 21990 13245 22056 13261
rect 21990 13181 21991 13245
rect 22055 13181 22056 13245
rect 21990 13165 22056 13181
rect 21990 13101 21991 13165
rect 22055 13101 22056 13165
rect 21990 13085 22056 13101
rect 21990 13021 21991 13085
rect 22055 13021 22056 13085
rect 21990 13005 22056 13021
rect 21990 12941 21991 13005
rect 22055 12941 22056 13005
rect 21990 12925 22056 12941
rect 21990 12861 21991 12925
rect 22055 12861 22056 12925
rect 21990 12845 22056 12861
rect 21990 12781 21991 12845
rect 22055 12781 22056 12845
rect 21990 12765 22056 12781
rect 21990 12701 21991 12765
rect 22055 12701 22056 12765
rect 21990 12685 22056 12701
rect 21990 12621 21991 12685
rect 22055 12621 22056 12685
rect 21990 12467 22056 12621
rect 22116 12529 22176 13559
rect 22236 12467 22296 13499
rect 22356 12529 22416 13559
rect 22476 12467 22536 13499
rect 22596 13405 22662 13495
rect 22596 13341 22597 13405
rect 22661 13341 22662 13405
rect 22596 13325 22662 13341
rect 22596 13261 22597 13325
rect 22661 13261 22662 13325
rect 22596 13245 22662 13261
rect 22596 13181 22597 13245
rect 22661 13181 22662 13245
rect 22596 13165 22662 13181
rect 22596 13101 22597 13165
rect 22661 13101 22662 13165
rect 22596 13085 22662 13101
rect 22596 13021 22597 13085
rect 22661 13021 22662 13085
rect 22596 13005 22662 13021
rect 22596 12941 22597 13005
rect 22661 12941 22662 13005
rect 22596 12925 22662 12941
rect 22596 12861 22597 12925
rect 22661 12861 22662 12925
rect 22596 12845 22662 12861
rect 22596 12781 22597 12845
rect 22661 12781 22662 12845
rect 22596 12765 22662 12781
rect 22596 12701 22597 12765
rect 22661 12701 22662 12765
rect 22596 12685 22662 12701
rect 22596 12621 22597 12685
rect 22661 12621 22662 12685
rect 22596 12467 22662 12621
rect 22722 12467 22782 13499
rect 22842 12529 22902 13559
rect 22962 12467 23022 13499
rect 23082 12529 23142 13559
rect 23202 13405 23268 13495
rect 23202 13341 23203 13405
rect 23267 13341 23268 13405
rect 23202 13325 23268 13341
rect 23202 13261 23203 13325
rect 23267 13261 23268 13325
rect 23202 13245 23268 13261
rect 23202 13181 23203 13245
rect 23267 13181 23268 13245
rect 23202 13165 23268 13181
rect 23202 13101 23203 13165
rect 23267 13101 23268 13165
rect 23202 13085 23268 13101
rect 23202 13021 23203 13085
rect 23267 13021 23268 13085
rect 23202 13005 23268 13021
rect 23202 12941 23203 13005
rect 23267 12941 23268 13005
rect 23202 12925 23268 12941
rect 23202 12861 23203 12925
rect 23267 12861 23268 12925
rect 23202 12845 23268 12861
rect 23202 12781 23203 12845
rect 23267 12781 23268 12845
rect 23202 12765 23268 12781
rect 23202 12701 23203 12765
rect 23267 12701 23268 12765
rect 23202 12685 23268 12701
rect 23202 12621 23203 12685
rect 23267 12621 23268 12685
rect 23202 12467 23268 12621
rect 23328 12529 23388 13559
rect 23448 12467 23508 13499
rect 23568 12529 23628 13559
rect 23688 12467 23748 13499
rect 23808 13405 23874 13495
rect 23808 13341 23809 13405
rect 23873 13341 23874 13405
rect 23808 13325 23874 13341
rect 23808 13261 23809 13325
rect 23873 13261 23874 13325
rect 23808 13245 23874 13261
rect 23808 13181 23809 13245
rect 23873 13181 23874 13245
rect 23808 13165 23874 13181
rect 23808 13101 23809 13165
rect 23873 13101 23874 13165
rect 23808 13085 23874 13101
rect 23808 13021 23809 13085
rect 23873 13021 23874 13085
rect 23808 13005 23874 13021
rect 23808 12941 23809 13005
rect 23873 12941 23874 13005
rect 23808 12925 23874 12941
rect 23808 12861 23809 12925
rect 23873 12861 23874 12925
rect 23808 12845 23874 12861
rect 23808 12781 23809 12845
rect 23873 12781 23874 12845
rect 23808 12765 23874 12781
rect 23808 12701 23809 12765
rect 23873 12701 23874 12765
rect 23808 12685 23874 12701
rect 23808 12621 23809 12685
rect 23873 12621 23874 12685
rect 23808 12467 23874 12621
rect 23934 12467 23994 13499
rect 24054 12529 24114 13559
rect 24174 12467 24234 13499
rect 24294 12529 24354 13559
rect 24414 13405 24480 13495
rect 24414 13341 24415 13405
rect 24479 13341 24480 13405
rect 24414 13325 24480 13341
rect 24414 13261 24415 13325
rect 24479 13261 24480 13325
rect 24414 13245 24480 13261
rect 24414 13181 24415 13245
rect 24479 13181 24480 13245
rect 24414 13165 24480 13181
rect 24414 13101 24415 13165
rect 24479 13101 24480 13165
rect 24414 13085 24480 13101
rect 24414 13021 24415 13085
rect 24479 13021 24480 13085
rect 24414 13005 24480 13021
rect 24414 12941 24415 13005
rect 24479 12941 24480 13005
rect 24414 12925 24480 12941
rect 24414 12861 24415 12925
rect 24479 12861 24480 12925
rect 24414 12845 24480 12861
rect 24414 12781 24415 12845
rect 24479 12781 24480 12845
rect 24414 12765 24480 12781
rect 24414 12701 24415 12765
rect 24479 12701 24480 12765
rect 24414 12685 24480 12701
rect 24414 12621 24415 12685
rect 24479 12621 24480 12685
rect 24414 12467 24480 12621
rect 24540 12529 24600 13559
rect 24660 12467 24720 13499
rect 24780 12529 24840 13559
rect 24900 12467 24960 13499
rect 25020 13405 25086 13495
rect 25020 13341 25021 13405
rect 25085 13341 25086 13405
rect 25020 13325 25086 13341
rect 25020 13261 25021 13325
rect 25085 13261 25086 13325
rect 25020 13245 25086 13261
rect 25020 13181 25021 13245
rect 25085 13181 25086 13245
rect 25020 13165 25086 13181
rect 25020 13101 25021 13165
rect 25085 13101 25086 13165
rect 25020 13085 25086 13101
rect 25020 13021 25021 13085
rect 25085 13021 25086 13085
rect 25020 13005 25086 13021
rect 25020 12941 25021 13005
rect 25085 12941 25086 13005
rect 25020 12925 25086 12941
rect 25020 12861 25021 12925
rect 25085 12861 25086 12925
rect 25020 12845 25086 12861
rect 25020 12781 25021 12845
rect 25085 12781 25086 12845
rect 25020 12765 25086 12781
rect 25020 12701 25021 12765
rect 25085 12701 25086 12765
rect 25020 12685 25086 12701
rect 25020 12621 25021 12685
rect 25085 12621 25086 12685
rect 25020 12467 25086 12621
rect 25146 12467 25206 13499
rect 25266 12529 25326 13559
rect 25386 12467 25446 13499
rect 25506 12529 25566 13559
rect 25626 13405 25692 13495
rect 25626 13341 25627 13405
rect 25691 13341 25692 13405
rect 25626 13325 25692 13341
rect 25626 13261 25627 13325
rect 25691 13261 25692 13325
rect 25626 13245 25692 13261
rect 25626 13181 25627 13245
rect 25691 13181 25692 13245
rect 25626 13165 25692 13181
rect 25626 13101 25627 13165
rect 25691 13101 25692 13165
rect 25626 13085 25692 13101
rect 25626 13021 25627 13085
rect 25691 13021 25692 13085
rect 25626 13005 25692 13021
rect 25626 12941 25627 13005
rect 25691 12941 25692 13005
rect 25626 12925 25692 12941
rect 25626 12861 25627 12925
rect 25691 12861 25692 12925
rect 25626 12845 25692 12861
rect 25626 12781 25627 12845
rect 25691 12781 25692 12845
rect 25626 12765 25692 12781
rect 25626 12701 25627 12765
rect 25691 12701 25692 12765
rect 25626 12685 25692 12701
rect 25626 12621 25627 12685
rect 25691 12621 25692 12685
rect 25626 12467 25692 12621
rect 25752 12529 25812 13559
rect 25872 12467 25932 13499
rect 25992 12529 26052 13559
rect 26437 13506 26468 13570
rect 26532 13506 26563 13570
rect 26112 12467 26172 13499
rect 26437 13496 26563 13506
rect 26232 13405 26298 13495
rect 26232 13341 26233 13405
rect 26297 13341 26298 13405
rect 26442 13426 26568 13436
rect 26442 13362 26473 13426
rect 26537 13362 26568 13426
rect 26442 13352 26568 13362
rect 26232 13325 26298 13341
rect 26232 13261 26233 13325
rect 26297 13261 26298 13325
rect 26232 13245 26298 13261
rect 26232 13181 26233 13245
rect 26297 13181 26298 13245
rect 26443 13274 26569 13284
rect 26443 13210 26474 13274
rect 26538 13210 26569 13274
rect 26443 13200 26569 13210
rect 26232 13165 26298 13181
rect 26232 13101 26233 13165
rect 26297 13101 26298 13165
rect 26232 13085 26298 13101
rect 26232 13021 26233 13085
rect 26297 13021 26298 13085
rect 26443 13104 26569 13114
rect 26443 13040 26474 13104
rect 26538 13040 26569 13104
rect 26443 13030 26569 13040
rect 26232 13005 26298 13021
rect 26232 12941 26233 13005
rect 26297 12941 26298 13005
rect 26232 12925 26298 12941
rect 26232 12861 26233 12925
rect 26297 12861 26298 12925
rect 26442 12947 26568 12957
rect 26442 12883 26473 12947
rect 26537 12883 26568 12947
rect 26442 12873 26568 12883
rect 26232 12845 26298 12861
rect 26232 12781 26233 12845
rect 26297 12781 26298 12845
rect 26232 12765 26298 12781
rect 26232 12701 26233 12765
rect 26297 12701 26298 12765
rect 26232 12685 26298 12701
rect 26232 12621 26233 12685
rect 26297 12621 26298 12685
rect 26360 12705 26486 12715
rect 26360 12641 26391 12705
rect 26455 12641 26486 12705
rect 26360 12631 26486 12641
rect 26232 12467 26298 12621
rect 21384 12465 26298 12467
rect 21384 12401 21488 12465
rect 21552 12401 21568 12465
rect 21632 12401 21648 12465
rect 21712 12401 21728 12465
rect 21792 12401 21808 12465
rect 21872 12442 21888 12465
rect 21872 12401 21877 12442
rect 21952 12401 22094 12465
rect 22158 12442 22174 12465
rect 22169 12401 22174 12442
rect 22238 12401 22254 12465
rect 22318 12401 22334 12465
rect 22398 12401 22414 12465
rect 22478 12401 22494 12465
rect 22558 12401 22700 12465
rect 22764 12401 22780 12465
rect 22844 12401 22860 12465
rect 22924 12401 22940 12465
rect 23004 12401 23020 12465
rect 23084 12442 23100 12465
rect 23084 12401 23089 12442
rect 23164 12401 23306 12465
rect 23370 12442 23386 12465
rect 23381 12401 23386 12442
rect 23450 12401 23466 12465
rect 23530 12401 23546 12465
rect 23610 12401 23626 12465
rect 23690 12401 23706 12465
rect 23770 12401 23912 12465
rect 23976 12401 23992 12465
rect 24056 12401 24072 12465
rect 24136 12401 24152 12465
rect 24216 12401 24232 12465
rect 24296 12442 24312 12465
rect 24296 12401 24301 12442
rect 24376 12401 24518 12465
rect 24582 12442 24598 12465
rect 24593 12401 24598 12442
rect 24662 12401 24678 12465
rect 24742 12401 24758 12465
rect 24822 12401 24838 12465
rect 24902 12401 24918 12465
rect 24982 12401 25124 12465
rect 25188 12401 25204 12465
rect 25268 12401 25284 12465
rect 25348 12401 25364 12465
rect 25428 12401 25444 12465
rect 25508 12442 25524 12465
rect 25508 12401 25513 12442
rect 25588 12401 25730 12465
rect 25794 12442 25810 12465
rect 25805 12401 25810 12442
rect 25874 12401 25890 12465
rect 25954 12401 25970 12465
rect 26034 12401 26050 12465
rect 26114 12401 26130 12465
rect 26194 12401 26298 12465
rect 21384 12399 21877 12401
rect 20652 12396 21145 12398
rect 19739 12370 19865 12380
rect 21135 12375 21145 12396
rect 21209 12396 21324 12398
rect 21209 12375 21218 12396
rect 21135 12370 21218 12375
rect 21867 12378 21877 12399
rect 21941 12399 22105 12401
rect 21941 12378 21950 12399
rect 21867 12373 21950 12378
rect 22096 12378 22105 12399
rect 22169 12399 23089 12401
rect 22169 12378 22179 12399
rect 22096 12373 22179 12378
rect 23079 12378 23089 12399
rect 23153 12399 23317 12401
rect 23153 12378 23162 12399
rect 23079 12373 23162 12378
rect 23308 12378 23317 12399
rect 23381 12399 24301 12401
rect 23381 12378 23391 12399
rect 23308 12373 23391 12378
rect 24291 12378 24301 12399
rect 24365 12399 24529 12401
rect 24365 12378 24374 12399
rect 24291 12373 24374 12378
rect 24520 12378 24529 12399
rect 24593 12399 25513 12401
rect 24593 12378 24603 12399
rect 24520 12373 24603 12378
rect 25503 12378 25513 12399
rect 25577 12399 25741 12401
rect 25577 12378 25586 12399
rect 25503 12373 25586 12378
rect 25732 12378 25741 12399
rect 25805 12399 26298 12401
rect 26448 12444 26574 12454
rect 25805 12378 25815 12399
rect 25732 12373 25815 12378
rect 26448 12380 26479 12444
rect 26543 12380 26574 12444
rect 26448 12370 26574 12380
rect 8635 12306 8636 12370
rect 8700 12306 8701 12370
rect 8635 12290 8701 12306
rect 8635 12226 8636 12290
rect 8700 12226 8701 12290
rect 9141 12282 9266 12292
rect 8635 12210 8701 12226
rect 8635 12146 8636 12210
rect 8700 12146 8701 12210
rect 8763 12230 8889 12240
rect 8763 12166 8794 12230
rect 8858 12166 8889 12230
rect 9141 12218 9171 12282
rect 9235 12218 9266 12282
rect 14783 12240 14865 12246
rect 14783 12219 14792 12240
rect 9141 12209 9266 12218
rect 14294 12217 14792 12219
rect 14856 12219 14865 12240
rect 15515 12240 15597 12246
rect 15515 12219 15524 12240
rect 14856 12217 14966 12219
rect 8763 12156 8889 12166
rect 8635 11992 8701 12146
rect 3787 11990 8701 11992
rect 3787 11926 3891 11990
rect 3955 11926 3971 11990
rect 4035 11926 4051 11990
rect 4115 11926 4131 11990
rect 4195 11926 4211 11990
rect 4275 11967 4291 11990
rect 4275 11926 4280 11967
rect 4355 11926 4497 11990
rect 4561 11967 4577 11990
rect 4572 11926 4577 11967
rect 4641 11926 4657 11990
rect 4721 11926 4737 11990
rect 4801 11926 4817 11990
rect 4881 11926 4897 11990
rect 4961 11926 5103 11990
rect 5167 11926 5183 11990
rect 5247 11926 5263 11990
rect 5327 11926 5343 11990
rect 5407 11926 5423 11990
rect 5487 11967 5503 11990
rect 5487 11926 5492 11967
rect 5567 11926 5709 11990
rect 5773 11967 5789 11990
rect 5784 11926 5789 11967
rect 5853 11926 5869 11990
rect 5933 11926 5949 11990
rect 6013 11926 6029 11990
rect 6093 11926 6109 11990
rect 6173 11926 6315 11990
rect 6379 11926 6395 11990
rect 6459 11926 6475 11990
rect 6539 11926 6555 11990
rect 6619 11926 6635 11990
rect 6699 11967 6715 11990
rect 6699 11926 6704 11967
rect 6779 11926 6921 11990
rect 6985 11967 7001 11990
rect 6996 11926 7001 11967
rect 7065 11926 7081 11990
rect 7145 11926 7161 11990
rect 7225 11926 7241 11990
rect 7305 11926 7321 11990
rect 7385 11926 7527 11990
rect 7591 11926 7607 11990
rect 7671 11926 7687 11990
rect 7751 11926 7767 11990
rect 7831 11926 7847 11990
rect 7911 11967 7927 11990
rect 7911 11926 7916 11967
rect 7991 11926 8133 11990
rect 8197 11967 8213 11990
rect 8208 11926 8213 11967
rect 8277 11926 8293 11990
rect 8357 11926 8373 11990
rect 8437 11926 8453 11990
rect 8517 11926 8533 11990
rect 8597 11926 8701 11990
rect 14294 12153 14398 12217
rect 14462 12153 14478 12217
rect 14542 12153 14558 12217
rect 14622 12153 14638 12217
rect 14702 12153 14718 12217
rect 14782 12176 14792 12217
rect 14782 12153 14798 12176
rect 14862 12153 14966 12217
rect 14294 12151 14966 12153
rect 14294 11997 14360 12151
rect 3787 11924 4280 11926
rect 3055 11921 3548 11923
rect 3538 11900 3548 11921
rect 3612 11921 3727 11923
rect 3612 11900 3621 11921
rect 3538 11895 3621 11900
rect 4270 11903 4280 11924
rect 4344 11924 4508 11926
rect 4344 11903 4353 11924
rect 4270 11898 4353 11903
rect 4499 11903 4508 11924
rect 4572 11924 5492 11926
rect 4572 11903 4582 11924
rect 4499 11898 4582 11903
rect 5482 11903 5492 11924
rect 5556 11924 5720 11926
rect 5556 11903 5565 11924
rect 5482 11898 5565 11903
rect 5711 11903 5720 11924
rect 5784 11924 6704 11926
rect 5784 11903 5794 11924
rect 5711 11898 5794 11903
rect 6694 11903 6704 11924
rect 6768 11924 6932 11926
rect 6768 11903 6777 11924
rect 6694 11898 6777 11903
rect 6923 11903 6932 11924
rect 6996 11924 7916 11926
rect 6996 11903 7006 11924
rect 6923 11898 7006 11903
rect 7906 11903 7916 11924
rect 7980 11924 8144 11926
rect 7980 11903 7989 11924
rect 7906 11898 7989 11903
rect 8135 11903 8144 11924
rect 8208 11924 8701 11926
rect 8851 11969 8977 11979
rect 8208 11903 8218 11924
rect 8135 11898 8218 11903
rect 8851 11905 8882 11969
rect 8946 11905 8977 11969
rect 8851 11895 8977 11905
rect 14294 11933 14295 11997
rect 14359 11933 14360 11997
rect 14294 11917 14360 11933
rect 10886 11885 11007 11894
rect 10886 11821 10913 11885
rect 10977 11821 11007 11885
rect 10886 11812 11007 11821
rect 11086 11888 11207 11897
rect 11086 11824 11113 11888
rect 11177 11824 11207 11888
rect 11086 11815 11207 11824
rect 11322 11886 11443 11895
rect 11322 11822 11349 11886
rect 11413 11822 11443 11886
rect 11322 11813 11443 11822
rect 11755 11880 11876 11889
rect 11755 11816 11782 11880
rect 11846 11816 11876 11880
rect 11755 11807 11876 11816
rect 11956 11881 12077 11890
rect 11956 11817 11983 11881
rect 12047 11817 12077 11881
rect 11956 11808 12077 11817
rect 12142 11879 12263 11888
rect 12142 11815 12169 11879
rect 12233 11815 12263 11879
rect 12142 11806 12263 11815
rect 12333 11882 12454 11891
rect 12333 11818 12360 11882
rect 12424 11818 12454 11882
rect 12333 11809 12454 11818
rect 12546 11881 12667 11890
rect 12546 11817 12573 11881
rect 12637 11817 12667 11881
rect 12546 11808 12667 11817
rect 14294 11853 14295 11917
rect 14359 11853 14360 11917
rect 14294 11837 14360 11853
rect 3895 11765 3977 11771
rect 3895 11744 3904 11765
rect 3406 11742 3904 11744
rect 3968 11744 3977 11765
rect 4627 11765 4709 11771
rect 4627 11744 4636 11765
rect 3968 11742 4078 11744
rect 3406 11678 3510 11742
rect 3574 11678 3590 11742
rect 3654 11678 3670 11742
rect 3734 11678 3750 11742
rect 3814 11678 3830 11742
rect 3894 11701 3904 11742
rect 3894 11678 3910 11701
rect 3974 11678 4078 11742
rect 3406 11676 4078 11678
rect 3406 11522 3472 11676
rect 3406 11458 3407 11522
rect 3471 11458 3472 11522
rect 3406 11442 3472 11458
rect 3406 11378 3407 11442
rect 3471 11378 3472 11442
rect 3406 11362 3472 11378
rect 3406 11298 3407 11362
rect 3471 11298 3472 11362
rect 3406 11282 3472 11298
rect 3406 11218 3407 11282
rect 3471 11218 3472 11282
rect 3406 11202 3472 11218
rect 3406 11138 3407 11202
rect 3471 11138 3472 11202
rect 3406 11122 3472 11138
rect 3406 11058 3407 11122
rect 3471 11058 3472 11122
rect 3406 11042 3472 11058
rect 3406 10978 3407 11042
rect 3471 10978 3472 11042
rect 3406 10962 3472 10978
rect 3406 10898 3407 10962
rect 3471 10898 3472 10962
rect 3406 10882 3472 10898
rect 3406 10818 3407 10882
rect 3471 10818 3472 10882
rect 3406 10802 3472 10818
rect 3406 10738 3407 10802
rect 3471 10738 3472 10802
rect 3406 10648 3472 10738
rect 3532 10644 3592 11676
rect 3018 10579 3143 10589
rect 3652 10584 3712 11614
rect 3772 10644 3832 11676
rect 3892 10584 3952 11614
rect 4012 11522 4078 11676
rect 4012 11458 4013 11522
rect 4077 11458 4078 11522
rect 4012 11442 4078 11458
rect 4012 11378 4013 11442
rect 4077 11378 4078 11442
rect 4012 11362 4078 11378
rect 4012 11298 4013 11362
rect 4077 11298 4078 11362
rect 4012 11282 4078 11298
rect 4012 11218 4013 11282
rect 4077 11218 4078 11282
rect 4012 11202 4078 11218
rect 4012 11138 4013 11202
rect 4077 11138 4078 11202
rect 4012 11122 4078 11138
rect 4012 11058 4013 11122
rect 4077 11058 4078 11122
rect 4012 11042 4078 11058
rect 4012 10978 4013 11042
rect 4077 10978 4078 11042
rect 4012 10962 4078 10978
rect 4012 10898 4013 10962
rect 4077 10898 4078 10962
rect 4012 10882 4078 10898
rect 4012 10818 4013 10882
rect 4077 10818 4078 10882
rect 4012 10802 4078 10818
rect 4012 10738 4013 10802
rect 4077 10738 4078 10802
rect 4012 10648 4078 10738
rect 4138 11742 4636 11744
rect 4700 11744 4709 11765
rect 4845 11765 4927 11771
rect 4845 11744 4854 11765
rect 4700 11742 4854 11744
rect 4918 11744 4927 11765
rect 5839 11765 5921 11771
rect 5839 11744 5848 11765
rect 4918 11742 5848 11744
rect 5912 11744 5921 11765
rect 6057 11765 6139 11771
rect 6057 11744 6066 11765
rect 5912 11742 6066 11744
rect 6130 11744 6139 11765
rect 7177 11765 7259 11771
rect 7177 11744 7186 11765
rect 6130 11742 6628 11744
rect 4138 11678 4242 11742
rect 4306 11678 4322 11742
rect 4386 11678 4402 11742
rect 4466 11678 4482 11742
rect 4546 11678 4562 11742
rect 4626 11701 4636 11742
rect 4626 11678 4642 11701
rect 4706 11678 4848 11742
rect 4918 11701 4928 11742
rect 4912 11678 4928 11701
rect 4992 11678 5008 11742
rect 5072 11678 5088 11742
rect 5152 11678 5168 11742
rect 5232 11678 5248 11742
rect 5312 11678 5454 11742
rect 5518 11678 5534 11742
rect 5598 11678 5614 11742
rect 5678 11678 5694 11742
rect 5758 11678 5774 11742
rect 5838 11701 5848 11742
rect 5838 11678 5854 11701
rect 5918 11678 6060 11742
rect 6130 11701 6140 11742
rect 6124 11678 6140 11701
rect 6204 11678 6220 11742
rect 6284 11678 6300 11742
rect 6364 11678 6380 11742
rect 6444 11678 6460 11742
rect 6524 11678 6628 11742
rect 4138 11676 6628 11678
rect 4138 11522 4204 11676
rect 4138 11458 4139 11522
rect 4203 11458 4204 11522
rect 4138 11442 4204 11458
rect 4138 11378 4139 11442
rect 4203 11378 4204 11442
rect 4138 11362 4204 11378
rect 4138 11298 4139 11362
rect 4203 11298 4204 11362
rect 4138 11282 4204 11298
rect 4138 11218 4139 11282
rect 4203 11218 4204 11282
rect 4138 11202 4204 11218
rect 4138 11138 4139 11202
rect 4203 11138 4204 11202
rect 4138 11122 4204 11138
rect 4138 11058 4139 11122
rect 4203 11058 4204 11122
rect 4138 11042 4204 11058
rect 4138 10978 4139 11042
rect 4203 10978 4204 11042
rect 4138 10962 4204 10978
rect 4138 10898 4139 10962
rect 4203 10898 4204 10962
rect 4138 10882 4204 10898
rect 4138 10818 4139 10882
rect 4203 10818 4204 10882
rect 4138 10802 4204 10818
rect 4138 10738 4139 10802
rect 4203 10738 4204 10802
rect 4138 10648 4204 10738
rect 4264 10644 4324 11676
rect 4384 10584 4444 11614
rect 4504 10644 4564 11676
rect 4624 10584 4684 11614
rect 4744 11522 4810 11676
rect 4744 11458 4745 11522
rect 4809 11458 4810 11522
rect 4744 11442 4810 11458
rect 4744 11378 4745 11442
rect 4809 11378 4810 11442
rect 4744 11362 4810 11378
rect 4744 11298 4745 11362
rect 4809 11298 4810 11362
rect 4744 11282 4810 11298
rect 4744 11218 4745 11282
rect 4809 11218 4810 11282
rect 4744 11202 4810 11218
rect 4744 11138 4745 11202
rect 4809 11138 4810 11202
rect 4744 11122 4810 11138
rect 4744 11058 4745 11122
rect 4809 11058 4810 11122
rect 4744 11042 4810 11058
rect 4744 10978 4745 11042
rect 4809 10978 4810 11042
rect 4744 10962 4810 10978
rect 4744 10898 4745 10962
rect 4809 10898 4810 10962
rect 4744 10882 4810 10898
rect 4744 10818 4745 10882
rect 4809 10818 4810 10882
rect 4744 10802 4810 10818
rect 4744 10738 4745 10802
rect 4809 10738 4810 10802
rect 4744 10648 4810 10738
rect 4870 10584 4930 11614
rect 4990 10644 5050 11676
rect 5110 10584 5170 11614
rect 5230 10644 5290 11676
rect 5350 11522 5416 11676
rect 5350 11458 5351 11522
rect 5415 11458 5416 11522
rect 5350 11442 5416 11458
rect 5350 11378 5351 11442
rect 5415 11378 5416 11442
rect 5350 11362 5416 11378
rect 5350 11298 5351 11362
rect 5415 11298 5416 11362
rect 5350 11282 5416 11298
rect 5350 11218 5351 11282
rect 5415 11218 5416 11282
rect 5350 11202 5416 11218
rect 5350 11138 5351 11202
rect 5415 11138 5416 11202
rect 5350 11122 5416 11138
rect 5350 11058 5351 11122
rect 5415 11058 5416 11122
rect 5350 11042 5416 11058
rect 5350 10978 5351 11042
rect 5415 10978 5416 11042
rect 5350 10962 5416 10978
rect 5350 10898 5351 10962
rect 5415 10898 5416 10962
rect 5350 10882 5416 10898
rect 5350 10818 5351 10882
rect 5415 10818 5416 10882
rect 5350 10802 5416 10818
rect 5350 10738 5351 10802
rect 5415 10738 5416 10802
rect 5350 10648 5416 10738
rect 5476 10644 5536 11676
rect 5596 10584 5656 11614
rect 5716 10644 5776 11676
rect 5836 10584 5896 11614
rect 5956 11522 6022 11676
rect 5956 11458 5957 11522
rect 6021 11458 6022 11522
rect 5956 11442 6022 11458
rect 5956 11378 5957 11442
rect 6021 11378 6022 11442
rect 5956 11362 6022 11378
rect 5956 11298 5957 11362
rect 6021 11298 6022 11362
rect 5956 11282 6022 11298
rect 5956 11218 5957 11282
rect 6021 11218 6022 11282
rect 5956 11202 6022 11218
rect 5956 11138 5957 11202
rect 6021 11138 6022 11202
rect 5956 11122 6022 11138
rect 5956 11058 5957 11122
rect 6021 11058 6022 11122
rect 5956 11042 6022 11058
rect 5956 10978 5957 11042
rect 6021 10978 6022 11042
rect 5956 10962 6022 10978
rect 5956 10898 5957 10962
rect 6021 10898 6022 10962
rect 5956 10882 6022 10898
rect 5956 10818 5957 10882
rect 6021 10818 6022 10882
rect 5956 10802 6022 10818
rect 5956 10738 5957 10802
rect 6021 10738 6022 10802
rect 5956 10648 6022 10738
rect 6082 10584 6142 11614
rect 6202 10644 6262 11676
rect 6322 10584 6382 11614
rect 6442 10644 6502 11676
rect 6562 11522 6628 11676
rect 6562 11458 6563 11522
rect 6627 11458 6628 11522
rect 6562 11442 6628 11458
rect 6562 11378 6563 11442
rect 6627 11378 6628 11442
rect 6562 11362 6628 11378
rect 6562 11298 6563 11362
rect 6627 11298 6628 11362
rect 6562 11282 6628 11298
rect 6562 11218 6563 11282
rect 6627 11218 6628 11282
rect 6562 11202 6628 11218
rect 6562 11138 6563 11202
rect 6627 11138 6628 11202
rect 6562 11122 6628 11138
rect 6562 11058 6563 11122
rect 6627 11058 6628 11122
rect 6562 11042 6628 11058
rect 6562 10978 6563 11042
rect 6627 10978 6628 11042
rect 6562 10962 6628 10978
rect 6562 10898 6563 10962
rect 6627 10898 6628 10962
rect 6562 10882 6628 10898
rect 6562 10818 6563 10882
rect 6627 10818 6628 10882
rect 6562 10802 6628 10818
rect 6562 10738 6563 10802
rect 6627 10738 6628 10802
rect 6562 10648 6628 10738
rect 6688 11742 7186 11744
rect 7250 11744 7259 11765
rect 7395 11765 7477 11771
rect 7395 11744 7404 11765
rect 7250 11742 7404 11744
rect 7468 11744 7477 11765
rect 8129 11765 8211 11771
rect 8129 11744 8138 11765
rect 7468 11742 7966 11744
rect 6688 11678 6792 11742
rect 6856 11678 6872 11742
rect 6936 11678 6952 11742
rect 7016 11678 7032 11742
rect 7096 11678 7112 11742
rect 7176 11701 7186 11742
rect 7176 11678 7192 11701
rect 7256 11678 7398 11742
rect 7468 11701 7478 11742
rect 7462 11678 7478 11701
rect 7542 11678 7558 11742
rect 7622 11678 7638 11742
rect 7702 11678 7718 11742
rect 7782 11678 7798 11742
rect 7862 11678 7966 11742
rect 6688 11676 7966 11678
rect 6688 11522 6754 11676
rect 6688 11458 6689 11522
rect 6753 11458 6754 11522
rect 6688 11442 6754 11458
rect 6688 11378 6689 11442
rect 6753 11378 6754 11442
rect 6688 11362 6754 11378
rect 6688 11298 6689 11362
rect 6753 11298 6754 11362
rect 6688 11282 6754 11298
rect 6688 11218 6689 11282
rect 6753 11218 6754 11282
rect 6688 11202 6754 11218
rect 6688 11138 6689 11202
rect 6753 11138 6754 11202
rect 6688 11122 6754 11138
rect 6688 11058 6689 11122
rect 6753 11058 6754 11122
rect 6688 11042 6754 11058
rect 6688 10978 6689 11042
rect 6753 10978 6754 11042
rect 6688 10962 6754 10978
rect 6688 10898 6689 10962
rect 6753 10898 6754 10962
rect 6688 10882 6754 10898
rect 6688 10818 6689 10882
rect 6753 10818 6754 10882
rect 6688 10802 6754 10818
rect 6688 10738 6689 10802
rect 6753 10738 6754 10802
rect 6688 10648 6754 10738
rect 6814 10644 6874 11676
rect 6934 10584 6994 11614
rect 7054 10644 7114 11676
rect 7174 10584 7234 11614
rect 7294 11522 7360 11676
rect 7294 11458 7295 11522
rect 7359 11458 7360 11522
rect 7294 11442 7360 11458
rect 7294 11378 7295 11442
rect 7359 11378 7360 11442
rect 7294 11362 7360 11378
rect 7294 11298 7295 11362
rect 7359 11298 7360 11362
rect 7294 11282 7360 11298
rect 7294 11218 7295 11282
rect 7359 11218 7360 11282
rect 7294 11202 7360 11218
rect 7294 11138 7295 11202
rect 7359 11138 7360 11202
rect 7294 11122 7360 11138
rect 7294 11058 7295 11122
rect 7359 11058 7360 11122
rect 7294 11042 7360 11058
rect 7294 10978 7295 11042
rect 7359 10978 7360 11042
rect 7294 10962 7360 10978
rect 7294 10898 7295 10962
rect 7359 10898 7360 10962
rect 7294 10882 7360 10898
rect 7294 10818 7295 10882
rect 7359 10818 7360 10882
rect 7294 10802 7360 10818
rect 7294 10738 7295 10802
rect 7359 10738 7360 10802
rect 7294 10648 7360 10738
rect 7420 10584 7480 11614
rect 7540 10644 7600 11676
rect 7660 10584 7720 11614
rect 7780 10644 7840 11676
rect 7900 11522 7966 11676
rect 7900 11458 7901 11522
rect 7965 11458 7966 11522
rect 7900 11442 7966 11458
rect 7900 11378 7901 11442
rect 7965 11378 7966 11442
rect 7900 11362 7966 11378
rect 7900 11298 7901 11362
rect 7965 11298 7966 11362
rect 7900 11282 7966 11298
rect 7900 11218 7901 11282
rect 7965 11218 7966 11282
rect 7900 11202 7966 11218
rect 7900 11138 7901 11202
rect 7965 11138 7966 11202
rect 7900 11122 7966 11138
rect 7900 11058 7901 11122
rect 7965 11058 7966 11122
rect 7900 11042 7966 11058
rect 7900 10978 7901 11042
rect 7965 10978 7966 11042
rect 7900 10962 7966 10978
rect 7900 10898 7901 10962
rect 7965 10898 7966 10962
rect 7900 10882 7966 10898
rect 7900 10818 7901 10882
rect 7965 10818 7966 10882
rect 7900 10802 7966 10818
rect 7900 10738 7901 10802
rect 7965 10738 7966 10802
rect 7900 10648 7966 10738
rect 8028 11742 8138 11744
rect 8202 11744 8211 11765
rect 8851 11766 8977 11776
rect 8202 11742 8700 11744
rect 8028 11678 8132 11742
rect 8202 11701 8212 11742
rect 8196 11678 8212 11701
rect 8276 11678 8292 11742
rect 8356 11678 8372 11742
rect 8436 11678 8452 11742
rect 8516 11678 8532 11742
rect 8596 11678 8700 11742
rect 8851 11702 8882 11766
rect 8946 11702 8977 11766
rect 8851 11692 8977 11702
rect 14294 11773 14295 11837
rect 14359 11773 14360 11837
rect 14294 11757 14360 11773
rect 14294 11693 14295 11757
rect 14359 11693 14360 11757
rect 8877 11691 8951 11692
rect 8028 11676 8700 11678
rect 8028 11522 8094 11676
rect 8028 11458 8029 11522
rect 8093 11458 8094 11522
rect 8028 11442 8094 11458
rect 8028 11378 8029 11442
rect 8093 11378 8094 11442
rect 8028 11362 8094 11378
rect 8028 11298 8029 11362
rect 8093 11298 8094 11362
rect 8028 11282 8094 11298
rect 8028 11218 8029 11282
rect 8093 11218 8094 11282
rect 8028 11202 8094 11218
rect 8028 11138 8029 11202
rect 8093 11138 8094 11202
rect 8028 11122 8094 11138
rect 8028 11058 8029 11122
rect 8093 11058 8094 11122
rect 8028 11042 8094 11058
rect 8028 10978 8029 11042
rect 8093 10978 8094 11042
rect 8028 10962 8094 10978
rect 8028 10898 8029 10962
rect 8093 10898 8094 10962
rect 8028 10882 8094 10898
rect 8028 10818 8029 10882
rect 8093 10818 8094 10882
rect 8028 10802 8094 10818
rect 8028 10738 8029 10802
rect 8093 10738 8094 10802
rect 8028 10648 8094 10738
rect 8154 10584 8214 11614
rect 8274 10644 8334 11676
rect 8394 10584 8454 11614
rect 8514 10644 8574 11676
rect 8634 11522 8700 11676
rect 14294 11677 14360 11693
rect 13261 11601 13425 11628
rect 13261 11595 13318 11601
rect 13261 11537 13314 11595
rect 13383 11537 13425 11601
rect 8634 11458 8635 11522
rect 8699 11458 8700 11522
rect 9164 11525 9289 11535
rect 8634 11442 8700 11458
rect 8634 11378 8635 11442
rect 8699 11378 8700 11442
rect 8761 11504 8886 11514
rect 8761 11440 8791 11504
rect 8855 11440 8886 11504
rect 9164 11461 9194 11525
rect 9258 11461 9289 11525
rect 13261 11506 13425 11537
rect 14294 11613 14295 11677
rect 14359 11613 14360 11677
rect 14294 11597 14360 11613
rect 14294 11533 14295 11597
rect 14359 11533 14360 11597
rect 14294 11517 14360 11533
rect 9164 11452 9289 11461
rect 14294 11453 14295 11517
rect 14359 11453 14360 11517
rect 8761 11430 8886 11440
rect 14294 11437 14360 11453
rect 8634 11362 8700 11378
rect 8634 11298 8635 11362
rect 8699 11298 8700 11362
rect 8634 11282 8700 11298
rect 8634 11218 8635 11282
rect 8699 11218 8700 11282
rect 14294 11373 14295 11437
rect 14359 11373 14360 11437
rect 14294 11357 14360 11373
rect 14294 11293 14295 11357
rect 14359 11293 14360 11357
rect 14294 11277 14360 11293
rect 8634 11202 8700 11218
rect 8634 11138 8635 11202
rect 8699 11138 8700 11202
rect 10899 11263 11024 11273
rect 10899 11199 10929 11263
rect 10993 11199 11024 11263
rect 10899 11189 11024 11199
rect 11087 11260 11212 11270
rect 11087 11196 11117 11260
rect 11181 11196 11212 11260
rect 11087 11186 11212 11196
rect 11284 11258 11409 11268
rect 11284 11194 11314 11258
rect 11378 11194 11409 11258
rect 11284 11184 11409 11194
rect 14294 11213 14295 11277
rect 14359 11213 14360 11277
rect 8634 11122 8700 11138
rect 14294 11123 14360 11213
rect 8634 11058 8635 11122
rect 8699 11058 8700 11122
rect 14420 11119 14480 12151
rect 8634 11042 8700 11058
rect 8634 10978 8635 11042
rect 8699 10978 8700 11042
rect 13906 11054 14031 11064
rect 14540 11059 14600 12089
rect 14660 11119 14720 12151
rect 14780 11059 14840 12089
rect 14900 11997 14966 12151
rect 14900 11933 14901 11997
rect 14965 11933 14966 11997
rect 14900 11917 14966 11933
rect 14900 11853 14901 11917
rect 14965 11853 14966 11917
rect 14900 11837 14966 11853
rect 14900 11773 14901 11837
rect 14965 11773 14966 11837
rect 14900 11757 14966 11773
rect 14900 11693 14901 11757
rect 14965 11693 14966 11757
rect 14900 11677 14966 11693
rect 14900 11613 14901 11677
rect 14965 11613 14966 11677
rect 14900 11597 14966 11613
rect 14900 11533 14901 11597
rect 14965 11533 14966 11597
rect 14900 11517 14966 11533
rect 14900 11453 14901 11517
rect 14965 11453 14966 11517
rect 14900 11437 14966 11453
rect 14900 11373 14901 11437
rect 14965 11373 14966 11437
rect 14900 11357 14966 11373
rect 14900 11293 14901 11357
rect 14965 11293 14966 11357
rect 14900 11277 14966 11293
rect 14900 11213 14901 11277
rect 14965 11213 14966 11277
rect 14900 11123 14966 11213
rect 15026 12217 15524 12219
rect 15588 12219 15597 12240
rect 15733 12240 15815 12246
rect 15733 12219 15742 12240
rect 15588 12217 15742 12219
rect 15806 12219 15815 12240
rect 16727 12240 16809 12246
rect 16727 12219 16736 12240
rect 15806 12217 16736 12219
rect 16800 12219 16809 12240
rect 16945 12240 17027 12246
rect 16945 12219 16954 12240
rect 16800 12217 16954 12219
rect 17018 12219 17027 12240
rect 18065 12240 18147 12246
rect 18065 12219 18074 12240
rect 17018 12217 17516 12219
rect 15026 12153 15130 12217
rect 15194 12153 15210 12217
rect 15274 12153 15290 12217
rect 15354 12153 15370 12217
rect 15434 12153 15450 12217
rect 15514 12176 15524 12217
rect 15514 12153 15530 12176
rect 15594 12153 15736 12217
rect 15806 12176 15816 12217
rect 15800 12153 15816 12176
rect 15880 12153 15896 12217
rect 15960 12153 15976 12217
rect 16040 12153 16056 12217
rect 16120 12153 16136 12217
rect 16200 12153 16342 12217
rect 16406 12153 16422 12217
rect 16486 12153 16502 12217
rect 16566 12153 16582 12217
rect 16646 12153 16662 12217
rect 16726 12176 16736 12217
rect 16726 12153 16742 12176
rect 16806 12153 16948 12217
rect 17018 12176 17028 12217
rect 17012 12153 17028 12176
rect 17092 12153 17108 12217
rect 17172 12153 17188 12217
rect 17252 12153 17268 12217
rect 17332 12153 17348 12217
rect 17412 12153 17516 12217
rect 15026 12151 17516 12153
rect 15026 11997 15092 12151
rect 15026 11933 15027 11997
rect 15091 11933 15092 11997
rect 15026 11917 15092 11933
rect 15026 11853 15027 11917
rect 15091 11853 15092 11917
rect 15026 11837 15092 11853
rect 15026 11773 15027 11837
rect 15091 11773 15092 11837
rect 15026 11757 15092 11773
rect 15026 11693 15027 11757
rect 15091 11693 15092 11757
rect 15026 11677 15092 11693
rect 15026 11613 15027 11677
rect 15091 11613 15092 11677
rect 15026 11597 15092 11613
rect 15026 11533 15027 11597
rect 15091 11533 15092 11597
rect 15026 11517 15092 11533
rect 15026 11453 15027 11517
rect 15091 11453 15092 11517
rect 15026 11437 15092 11453
rect 15026 11373 15027 11437
rect 15091 11373 15092 11437
rect 15026 11357 15092 11373
rect 15026 11293 15027 11357
rect 15091 11293 15092 11357
rect 15026 11277 15092 11293
rect 15026 11213 15027 11277
rect 15091 11213 15092 11277
rect 15026 11123 15092 11213
rect 15152 11119 15212 12151
rect 15272 11059 15332 12089
rect 15392 11119 15452 12151
rect 15512 11059 15572 12089
rect 15632 11997 15698 12151
rect 15632 11933 15633 11997
rect 15697 11933 15698 11997
rect 15632 11917 15698 11933
rect 15632 11853 15633 11917
rect 15697 11853 15698 11917
rect 15632 11837 15698 11853
rect 15632 11773 15633 11837
rect 15697 11773 15698 11837
rect 15632 11757 15698 11773
rect 15632 11693 15633 11757
rect 15697 11693 15698 11757
rect 15632 11677 15698 11693
rect 15632 11613 15633 11677
rect 15697 11613 15698 11677
rect 15632 11597 15698 11613
rect 15632 11533 15633 11597
rect 15697 11533 15698 11597
rect 15632 11517 15698 11533
rect 15632 11453 15633 11517
rect 15697 11453 15698 11517
rect 15632 11437 15698 11453
rect 15632 11373 15633 11437
rect 15697 11373 15698 11437
rect 15632 11357 15698 11373
rect 15632 11293 15633 11357
rect 15697 11293 15698 11357
rect 15632 11277 15698 11293
rect 15632 11213 15633 11277
rect 15697 11213 15698 11277
rect 15632 11123 15698 11213
rect 15758 11059 15818 12089
rect 15878 11119 15938 12151
rect 15998 11059 16058 12089
rect 16118 11119 16178 12151
rect 16238 11997 16304 12151
rect 16238 11933 16239 11997
rect 16303 11933 16304 11997
rect 16238 11917 16304 11933
rect 16238 11853 16239 11917
rect 16303 11853 16304 11917
rect 16238 11837 16304 11853
rect 16238 11773 16239 11837
rect 16303 11773 16304 11837
rect 16238 11757 16304 11773
rect 16238 11693 16239 11757
rect 16303 11693 16304 11757
rect 16238 11677 16304 11693
rect 16238 11613 16239 11677
rect 16303 11613 16304 11677
rect 16238 11597 16304 11613
rect 16238 11533 16239 11597
rect 16303 11533 16304 11597
rect 16238 11517 16304 11533
rect 16238 11453 16239 11517
rect 16303 11453 16304 11517
rect 16238 11437 16304 11453
rect 16238 11373 16239 11437
rect 16303 11373 16304 11437
rect 16238 11357 16304 11373
rect 16238 11293 16239 11357
rect 16303 11293 16304 11357
rect 16238 11277 16304 11293
rect 16238 11213 16239 11277
rect 16303 11213 16304 11277
rect 16238 11123 16304 11213
rect 16364 11119 16424 12151
rect 16484 11059 16544 12089
rect 16604 11119 16664 12151
rect 16724 11059 16784 12089
rect 16844 11997 16910 12151
rect 16844 11933 16845 11997
rect 16909 11933 16910 11997
rect 16844 11917 16910 11933
rect 16844 11853 16845 11917
rect 16909 11853 16910 11917
rect 16844 11837 16910 11853
rect 16844 11773 16845 11837
rect 16909 11773 16910 11837
rect 16844 11757 16910 11773
rect 16844 11693 16845 11757
rect 16909 11693 16910 11757
rect 16844 11677 16910 11693
rect 16844 11613 16845 11677
rect 16909 11613 16910 11677
rect 16844 11597 16910 11613
rect 16844 11533 16845 11597
rect 16909 11533 16910 11597
rect 16844 11517 16910 11533
rect 16844 11453 16845 11517
rect 16909 11453 16910 11517
rect 16844 11437 16910 11453
rect 16844 11373 16845 11437
rect 16909 11373 16910 11437
rect 16844 11357 16910 11373
rect 16844 11293 16845 11357
rect 16909 11293 16910 11357
rect 16844 11277 16910 11293
rect 16844 11213 16845 11277
rect 16909 11213 16910 11277
rect 16844 11123 16910 11213
rect 16970 11059 17030 12089
rect 17090 11119 17150 12151
rect 17210 11059 17270 12089
rect 17330 11119 17390 12151
rect 17450 11997 17516 12151
rect 17450 11933 17451 11997
rect 17515 11933 17516 11997
rect 17450 11917 17516 11933
rect 17450 11853 17451 11917
rect 17515 11853 17516 11917
rect 17450 11837 17516 11853
rect 17450 11773 17451 11837
rect 17515 11773 17516 11837
rect 17450 11757 17516 11773
rect 17450 11693 17451 11757
rect 17515 11693 17516 11757
rect 17450 11677 17516 11693
rect 17450 11613 17451 11677
rect 17515 11613 17516 11677
rect 17450 11597 17516 11613
rect 17450 11533 17451 11597
rect 17515 11533 17516 11597
rect 17450 11517 17516 11533
rect 17450 11453 17451 11517
rect 17515 11453 17516 11517
rect 17450 11437 17516 11453
rect 17450 11373 17451 11437
rect 17515 11373 17516 11437
rect 17450 11357 17516 11373
rect 17450 11293 17451 11357
rect 17515 11293 17516 11357
rect 17450 11277 17516 11293
rect 17450 11213 17451 11277
rect 17515 11213 17516 11277
rect 17450 11123 17516 11213
rect 17576 12217 18074 12219
rect 18138 12219 18147 12240
rect 18283 12240 18365 12246
rect 18283 12219 18292 12240
rect 18138 12217 18292 12219
rect 18356 12219 18365 12240
rect 19017 12240 19099 12246
rect 19017 12219 19026 12240
rect 18356 12217 18854 12219
rect 17576 12153 17680 12217
rect 17744 12153 17760 12217
rect 17824 12153 17840 12217
rect 17904 12153 17920 12217
rect 17984 12153 18000 12217
rect 18064 12176 18074 12217
rect 18064 12153 18080 12176
rect 18144 12153 18286 12217
rect 18356 12176 18366 12217
rect 18350 12153 18366 12176
rect 18430 12153 18446 12217
rect 18510 12153 18526 12217
rect 18590 12153 18606 12217
rect 18670 12153 18686 12217
rect 18750 12153 18854 12217
rect 17576 12151 18854 12153
rect 17576 11997 17642 12151
rect 17576 11933 17577 11997
rect 17641 11933 17642 11997
rect 17576 11917 17642 11933
rect 17576 11853 17577 11917
rect 17641 11853 17642 11917
rect 17576 11837 17642 11853
rect 17576 11773 17577 11837
rect 17641 11773 17642 11837
rect 17576 11757 17642 11773
rect 17576 11693 17577 11757
rect 17641 11693 17642 11757
rect 17576 11677 17642 11693
rect 17576 11613 17577 11677
rect 17641 11613 17642 11677
rect 17576 11597 17642 11613
rect 17576 11533 17577 11597
rect 17641 11533 17642 11597
rect 17576 11517 17642 11533
rect 17576 11453 17577 11517
rect 17641 11453 17642 11517
rect 17576 11437 17642 11453
rect 17576 11373 17577 11437
rect 17641 11373 17642 11437
rect 17576 11357 17642 11373
rect 17576 11293 17577 11357
rect 17641 11293 17642 11357
rect 17576 11277 17642 11293
rect 17576 11213 17577 11277
rect 17641 11213 17642 11277
rect 17576 11123 17642 11213
rect 17702 11119 17762 12151
rect 17822 11059 17882 12089
rect 17942 11119 18002 12151
rect 18062 11059 18122 12089
rect 18182 11997 18248 12151
rect 18182 11933 18183 11997
rect 18247 11933 18248 11997
rect 18182 11917 18248 11933
rect 18182 11853 18183 11917
rect 18247 11853 18248 11917
rect 18182 11837 18248 11853
rect 18182 11773 18183 11837
rect 18247 11773 18248 11837
rect 18182 11757 18248 11773
rect 18182 11693 18183 11757
rect 18247 11693 18248 11757
rect 18182 11677 18248 11693
rect 18182 11613 18183 11677
rect 18247 11613 18248 11677
rect 18182 11597 18248 11613
rect 18182 11533 18183 11597
rect 18247 11533 18248 11597
rect 18182 11517 18248 11533
rect 18182 11453 18183 11517
rect 18247 11453 18248 11517
rect 18182 11437 18248 11453
rect 18182 11373 18183 11437
rect 18247 11373 18248 11437
rect 18182 11357 18248 11373
rect 18182 11293 18183 11357
rect 18247 11293 18248 11357
rect 18182 11277 18248 11293
rect 18182 11213 18183 11277
rect 18247 11213 18248 11277
rect 18182 11123 18248 11213
rect 18308 11059 18368 12089
rect 18428 11119 18488 12151
rect 18548 11059 18608 12089
rect 18668 11119 18728 12151
rect 18788 11997 18854 12151
rect 18788 11933 18789 11997
rect 18853 11933 18854 11997
rect 18788 11917 18854 11933
rect 18788 11853 18789 11917
rect 18853 11853 18854 11917
rect 18788 11837 18854 11853
rect 18788 11773 18789 11837
rect 18853 11773 18854 11837
rect 18788 11757 18854 11773
rect 18788 11693 18789 11757
rect 18853 11693 18854 11757
rect 18788 11677 18854 11693
rect 18788 11613 18789 11677
rect 18853 11613 18854 11677
rect 18788 11597 18854 11613
rect 18788 11533 18789 11597
rect 18853 11533 18854 11597
rect 18788 11517 18854 11533
rect 18788 11453 18789 11517
rect 18853 11453 18854 11517
rect 18788 11437 18854 11453
rect 18788 11373 18789 11437
rect 18853 11373 18854 11437
rect 18788 11357 18854 11373
rect 18788 11293 18789 11357
rect 18853 11293 18854 11357
rect 18788 11277 18854 11293
rect 18788 11213 18789 11277
rect 18853 11213 18854 11277
rect 18788 11123 18854 11213
rect 18916 12217 19026 12219
rect 19090 12219 19099 12240
rect 19739 12241 19865 12251
rect 19090 12217 19588 12219
rect 18916 12153 19020 12217
rect 19090 12176 19100 12217
rect 19084 12153 19100 12176
rect 19164 12153 19180 12217
rect 19244 12153 19260 12217
rect 19324 12153 19340 12217
rect 19404 12153 19420 12217
rect 19484 12153 19588 12217
rect 19739 12177 19770 12241
rect 19834 12177 19865 12241
rect 21492 12240 21574 12246
rect 21492 12219 21501 12240
rect 19739 12167 19865 12177
rect 21003 12217 21501 12219
rect 21565 12219 21574 12240
rect 22224 12240 22306 12246
rect 22224 12219 22233 12240
rect 21565 12217 21675 12219
rect 19765 12166 19839 12167
rect 18916 12151 19588 12153
rect 18916 11997 18982 12151
rect 18916 11933 18917 11997
rect 18981 11933 18982 11997
rect 18916 11917 18982 11933
rect 18916 11853 18917 11917
rect 18981 11853 18982 11917
rect 18916 11837 18982 11853
rect 18916 11773 18917 11837
rect 18981 11773 18982 11837
rect 18916 11757 18982 11773
rect 18916 11693 18917 11757
rect 18981 11693 18982 11757
rect 18916 11677 18982 11693
rect 18916 11613 18917 11677
rect 18981 11613 18982 11677
rect 18916 11597 18982 11613
rect 18916 11533 18917 11597
rect 18981 11533 18982 11597
rect 18916 11517 18982 11533
rect 18916 11453 18917 11517
rect 18981 11453 18982 11517
rect 18916 11437 18982 11453
rect 18916 11373 18917 11437
rect 18981 11373 18982 11437
rect 18916 11357 18982 11373
rect 18916 11293 18917 11357
rect 18981 11293 18982 11357
rect 18916 11277 18982 11293
rect 18916 11213 18917 11277
rect 18981 11213 18982 11277
rect 18916 11123 18982 11213
rect 19042 11059 19102 12089
rect 19162 11119 19222 12151
rect 19282 11059 19342 12089
rect 19402 11119 19462 12151
rect 19522 11997 19588 12151
rect 19522 11933 19523 11997
rect 19587 11933 19588 11997
rect 21003 12153 21107 12217
rect 21171 12153 21187 12217
rect 21251 12153 21267 12217
rect 21331 12153 21347 12217
rect 21411 12153 21427 12217
rect 21491 12176 21501 12217
rect 21491 12153 21507 12176
rect 21571 12153 21675 12217
rect 21003 12151 21675 12153
rect 21003 11997 21069 12151
rect 19522 11917 19588 11933
rect 19522 11853 19523 11917
rect 19587 11853 19588 11917
rect 19649 11979 19774 11989
rect 19649 11915 19679 11979
rect 19743 11915 19774 11979
rect 19649 11905 19774 11915
rect 21003 11933 21004 11997
rect 21068 11933 21069 11997
rect 21003 11917 21069 11933
rect 19522 11837 19588 11853
rect 19522 11773 19523 11837
rect 19587 11773 19588 11837
rect 19522 11757 19588 11773
rect 19522 11693 19523 11757
rect 19587 11693 19588 11757
rect 19522 11677 19588 11693
rect 19522 11613 19523 11677
rect 19587 11613 19588 11677
rect 19522 11597 19588 11613
rect 19522 11533 19523 11597
rect 19587 11533 19588 11597
rect 19522 11517 19588 11533
rect 19522 11453 19523 11517
rect 19587 11453 19588 11517
rect 19522 11437 19588 11453
rect 19522 11373 19523 11437
rect 19587 11373 19588 11437
rect 19522 11357 19588 11373
rect 19522 11293 19523 11357
rect 19587 11293 19588 11357
rect 19522 11277 19588 11293
rect 19522 11213 19523 11277
rect 19587 11213 19588 11277
rect 19522 11123 19588 11213
rect 21003 11853 21004 11917
rect 21068 11853 21069 11917
rect 21003 11837 21069 11853
rect 21003 11773 21004 11837
rect 21068 11773 21069 11837
rect 21003 11757 21069 11773
rect 21003 11693 21004 11757
rect 21068 11693 21069 11757
rect 21003 11677 21069 11693
rect 21003 11613 21004 11677
rect 21068 11613 21069 11677
rect 21003 11597 21069 11613
rect 21003 11533 21004 11597
rect 21068 11533 21069 11597
rect 21003 11517 21069 11533
rect 21003 11453 21004 11517
rect 21068 11453 21069 11517
rect 21003 11437 21069 11453
rect 21003 11373 21004 11437
rect 21068 11373 21069 11437
rect 21003 11357 21069 11373
rect 21003 11293 21004 11357
rect 21068 11293 21069 11357
rect 21003 11277 21069 11293
rect 21003 11213 21004 11277
rect 21068 11213 21069 11277
rect 21003 11123 21069 11213
rect 21129 11119 21189 12151
rect 13906 10990 13936 11054
rect 14000 10990 14031 11054
rect 14294 11057 14966 11059
rect 14294 10993 14478 11057
rect 14542 10993 14558 11057
rect 14622 10993 14638 11057
rect 14702 10993 14718 11057
rect 14782 10993 14966 11057
rect 14294 10991 14966 10993
rect 15026 11057 17516 11059
rect 15026 10993 15210 11057
rect 15274 10993 15290 11057
rect 15354 10993 15370 11057
rect 15434 10993 15450 11057
rect 15514 10993 15816 11057
rect 15880 10993 15896 11057
rect 15960 10993 15976 11057
rect 16040 10993 16056 11057
rect 16120 10993 16422 11057
rect 16486 10993 16502 11057
rect 16566 10993 16582 11057
rect 16646 10993 16662 11057
rect 16726 10993 17028 11057
rect 17092 10993 17108 11057
rect 17172 10993 17188 11057
rect 17252 10993 17268 11057
rect 17332 10993 17516 11057
rect 15026 10991 17516 10993
rect 17576 11057 18854 11059
rect 17576 10993 17760 11057
rect 17824 10993 17840 11057
rect 17904 10993 17920 11057
rect 17984 10993 18000 11057
rect 18064 10993 18366 11057
rect 18430 10993 18446 11057
rect 18510 10993 18526 11057
rect 18590 10993 18606 11057
rect 18670 10993 18854 11057
rect 17576 10991 18854 10993
rect 18916 11057 19588 11059
rect 18916 10993 19100 11057
rect 19164 10993 19180 11057
rect 19244 10993 19260 11057
rect 19324 10993 19340 11057
rect 19404 10993 19588 11057
rect 18916 10991 19588 10993
rect 20615 11054 20740 11064
rect 21249 11059 21309 12089
rect 21369 11119 21429 12151
rect 21489 11059 21549 12089
rect 21609 11997 21675 12151
rect 21609 11933 21610 11997
rect 21674 11933 21675 11997
rect 21609 11917 21675 11933
rect 21609 11853 21610 11917
rect 21674 11853 21675 11917
rect 21609 11837 21675 11853
rect 21609 11773 21610 11837
rect 21674 11773 21675 11837
rect 21609 11757 21675 11773
rect 21609 11693 21610 11757
rect 21674 11693 21675 11757
rect 21609 11677 21675 11693
rect 21609 11613 21610 11677
rect 21674 11613 21675 11677
rect 21609 11597 21675 11613
rect 21609 11533 21610 11597
rect 21674 11533 21675 11597
rect 21609 11517 21675 11533
rect 21609 11453 21610 11517
rect 21674 11453 21675 11517
rect 21609 11437 21675 11453
rect 21609 11373 21610 11437
rect 21674 11373 21675 11437
rect 21609 11357 21675 11373
rect 21609 11293 21610 11357
rect 21674 11293 21675 11357
rect 21609 11277 21675 11293
rect 21609 11213 21610 11277
rect 21674 11213 21675 11277
rect 21609 11123 21675 11213
rect 21735 12217 22233 12219
rect 22297 12219 22306 12240
rect 22442 12240 22524 12246
rect 22442 12219 22451 12240
rect 22297 12217 22451 12219
rect 22515 12219 22524 12240
rect 23436 12240 23518 12246
rect 23436 12219 23445 12240
rect 22515 12217 23445 12219
rect 23509 12219 23518 12240
rect 23654 12240 23736 12246
rect 23654 12219 23663 12240
rect 23509 12217 23663 12219
rect 23727 12219 23736 12240
rect 24774 12240 24856 12246
rect 24774 12219 24783 12240
rect 23727 12217 24225 12219
rect 21735 12153 21839 12217
rect 21903 12153 21919 12217
rect 21983 12153 21999 12217
rect 22063 12153 22079 12217
rect 22143 12153 22159 12217
rect 22223 12176 22233 12217
rect 22223 12153 22239 12176
rect 22303 12153 22445 12217
rect 22515 12176 22525 12217
rect 22509 12153 22525 12176
rect 22589 12153 22605 12217
rect 22669 12153 22685 12217
rect 22749 12153 22765 12217
rect 22829 12153 22845 12217
rect 22909 12153 23051 12217
rect 23115 12153 23131 12217
rect 23195 12153 23211 12217
rect 23275 12153 23291 12217
rect 23355 12153 23371 12217
rect 23435 12176 23445 12217
rect 23435 12153 23451 12176
rect 23515 12153 23657 12217
rect 23727 12176 23737 12217
rect 23721 12153 23737 12176
rect 23801 12153 23817 12217
rect 23881 12153 23897 12217
rect 23961 12153 23977 12217
rect 24041 12153 24057 12217
rect 24121 12153 24225 12217
rect 21735 12151 24225 12153
rect 21735 11997 21801 12151
rect 21735 11933 21736 11997
rect 21800 11933 21801 11997
rect 21735 11917 21801 11933
rect 21735 11853 21736 11917
rect 21800 11853 21801 11917
rect 21735 11837 21801 11853
rect 21735 11773 21736 11837
rect 21800 11773 21801 11837
rect 21735 11757 21801 11773
rect 21735 11693 21736 11757
rect 21800 11693 21801 11757
rect 21735 11677 21801 11693
rect 21735 11613 21736 11677
rect 21800 11613 21801 11677
rect 21735 11597 21801 11613
rect 21735 11533 21736 11597
rect 21800 11533 21801 11597
rect 21735 11517 21801 11533
rect 21735 11453 21736 11517
rect 21800 11453 21801 11517
rect 21735 11437 21801 11453
rect 21735 11373 21736 11437
rect 21800 11373 21801 11437
rect 21735 11357 21801 11373
rect 21735 11293 21736 11357
rect 21800 11293 21801 11357
rect 21735 11277 21801 11293
rect 21735 11213 21736 11277
rect 21800 11213 21801 11277
rect 21735 11123 21801 11213
rect 21861 11119 21921 12151
rect 21981 11059 22041 12089
rect 22101 11119 22161 12151
rect 22221 11059 22281 12089
rect 22341 11997 22407 12151
rect 22341 11933 22342 11997
rect 22406 11933 22407 11997
rect 22341 11917 22407 11933
rect 22341 11853 22342 11917
rect 22406 11853 22407 11917
rect 22341 11837 22407 11853
rect 22341 11773 22342 11837
rect 22406 11773 22407 11837
rect 22341 11757 22407 11773
rect 22341 11693 22342 11757
rect 22406 11693 22407 11757
rect 22341 11677 22407 11693
rect 22341 11613 22342 11677
rect 22406 11613 22407 11677
rect 22341 11597 22407 11613
rect 22341 11533 22342 11597
rect 22406 11533 22407 11597
rect 22341 11517 22407 11533
rect 22341 11453 22342 11517
rect 22406 11453 22407 11517
rect 22341 11437 22407 11453
rect 22341 11373 22342 11437
rect 22406 11373 22407 11437
rect 22341 11357 22407 11373
rect 22341 11293 22342 11357
rect 22406 11293 22407 11357
rect 22341 11277 22407 11293
rect 22341 11213 22342 11277
rect 22406 11213 22407 11277
rect 22341 11123 22407 11213
rect 22467 11059 22527 12089
rect 22587 11119 22647 12151
rect 22707 11059 22767 12089
rect 22827 11119 22887 12151
rect 22947 11997 23013 12151
rect 22947 11933 22948 11997
rect 23012 11933 23013 11997
rect 22947 11917 23013 11933
rect 22947 11853 22948 11917
rect 23012 11853 23013 11917
rect 22947 11837 23013 11853
rect 22947 11773 22948 11837
rect 23012 11773 23013 11837
rect 22947 11757 23013 11773
rect 22947 11693 22948 11757
rect 23012 11693 23013 11757
rect 22947 11677 23013 11693
rect 22947 11613 22948 11677
rect 23012 11613 23013 11677
rect 22947 11597 23013 11613
rect 22947 11533 22948 11597
rect 23012 11533 23013 11597
rect 22947 11517 23013 11533
rect 22947 11453 22948 11517
rect 23012 11453 23013 11517
rect 22947 11437 23013 11453
rect 22947 11373 22948 11437
rect 23012 11373 23013 11437
rect 22947 11357 23013 11373
rect 22947 11293 22948 11357
rect 23012 11293 23013 11357
rect 22947 11277 23013 11293
rect 22947 11213 22948 11277
rect 23012 11213 23013 11277
rect 22947 11123 23013 11213
rect 23073 11119 23133 12151
rect 23193 11059 23253 12089
rect 23313 11119 23373 12151
rect 23433 11059 23493 12089
rect 23553 11997 23619 12151
rect 23553 11933 23554 11997
rect 23618 11933 23619 11997
rect 23553 11917 23619 11933
rect 23553 11853 23554 11917
rect 23618 11853 23619 11917
rect 23553 11837 23619 11853
rect 23553 11773 23554 11837
rect 23618 11773 23619 11837
rect 23553 11757 23619 11773
rect 23553 11693 23554 11757
rect 23618 11693 23619 11757
rect 23553 11677 23619 11693
rect 23553 11613 23554 11677
rect 23618 11613 23619 11677
rect 23553 11597 23619 11613
rect 23553 11533 23554 11597
rect 23618 11533 23619 11597
rect 23553 11517 23619 11533
rect 23553 11453 23554 11517
rect 23618 11453 23619 11517
rect 23553 11437 23619 11453
rect 23553 11373 23554 11437
rect 23618 11373 23619 11437
rect 23553 11357 23619 11373
rect 23553 11293 23554 11357
rect 23618 11293 23619 11357
rect 23553 11277 23619 11293
rect 23553 11213 23554 11277
rect 23618 11213 23619 11277
rect 23553 11123 23619 11213
rect 23679 11059 23739 12089
rect 23799 11119 23859 12151
rect 23919 11059 23979 12089
rect 24039 11119 24099 12151
rect 24159 11997 24225 12151
rect 24159 11933 24160 11997
rect 24224 11933 24225 11997
rect 24159 11917 24225 11933
rect 24159 11853 24160 11917
rect 24224 11853 24225 11917
rect 24159 11837 24225 11853
rect 24159 11773 24160 11837
rect 24224 11773 24225 11837
rect 24159 11757 24225 11773
rect 24159 11693 24160 11757
rect 24224 11693 24225 11757
rect 24159 11677 24225 11693
rect 24159 11613 24160 11677
rect 24224 11613 24225 11677
rect 24159 11597 24225 11613
rect 24159 11533 24160 11597
rect 24224 11533 24225 11597
rect 24159 11517 24225 11533
rect 24159 11453 24160 11517
rect 24224 11453 24225 11517
rect 24159 11437 24225 11453
rect 24159 11373 24160 11437
rect 24224 11373 24225 11437
rect 24159 11357 24225 11373
rect 24159 11293 24160 11357
rect 24224 11293 24225 11357
rect 24159 11277 24225 11293
rect 24159 11213 24160 11277
rect 24224 11213 24225 11277
rect 24159 11123 24225 11213
rect 24285 12217 24783 12219
rect 24847 12219 24856 12240
rect 24992 12240 25074 12246
rect 24992 12219 25001 12240
rect 24847 12217 25001 12219
rect 25065 12219 25074 12240
rect 25726 12240 25808 12246
rect 25726 12219 25735 12240
rect 25065 12217 25563 12219
rect 24285 12153 24389 12217
rect 24453 12153 24469 12217
rect 24533 12153 24549 12217
rect 24613 12153 24629 12217
rect 24693 12153 24709 12217
rect 24773 12176 24783 12217
rect 24773 12153 24789 12176
rect 24853 12153 24995 12217
rect 25065 12176 25075 12217
rect 25059 12153 25075 12176
rect 25139 12153 25155 12217
rect 25219 12153 25235 12217
rect 25299 12153 25315 12217
rect 25379 12153 25395 12217
rect 25459 12153 25563 12217
rect 24285 12151 25563 12153
rect 24285 11997 24351 12151
rect 24285 11933 24286 11997
rect 24350 11933 24351 11997
rect 24285 11917 24351 11933
rect 24285 11853 24286 11917
rect 24350 11853 24351 11917
rect 24285 11837 24351 11853
rect 24285 11773 24286 11837
rect 24350 11773 24351 11837
rect 24285 11757 24351 11773
rect 24285 11693 24286 11757
rect 24350 11693 24351 11757
rect 24285 11677 24351 11693
rect 24285 11613 24286 11677
rect 24350 11613 24351 11677
rect 24285 11597 24351 11613
rect 24285 11533 24286 11597
rect 24350 11533 24351 11597
rect 24285 11517 24351 11533
rect 24285 11453 24286 11517
rect 24350 11453 24351 11517
rect 24285 11437 24351 11453
rect 24285 11373 24286 11437
rect 24350 11373 24351 11437
rect 24285 11357 24351 11373
rect 24285 11293 24286 11357
rect 24350 11293 24351 11357
rect 24285 11277 24351 11293
rect 24285 11213 24286 11277
rect 24350 11213 24351 11277
rect 24285 11123 24351 11213
rect 24411 11119 24471 12151
rect 24531 11059 24591 12089
rect 24651 11119 24711 12151
rect 24771 11059 24831 12089
rect 24891 11997 24957 12151
rect 24891 11933 24892 11997
rect 24956 11933 24957 11997
rect 24891 11917 24957 11933
rect 24891 11853 24892 11917
rect 24956 11853 24957 11917
rect 24891 11837 24957 11853
rect 24891 11773 24892 11837
rect 24956 11773 24957 11837
rect 24891 11757 24957 11773
rect 24891 11693 24892 11757
rect 24956 11693 24957 11757
rect 24891 11677 24957 11693
rect 24891 11613 24892 11677
rect 24956 11613 24957 11677
rect 24891 11597 24957 11613
rect 24891 11533 24892 11597
rect 24956 11533 24957 11597
rect 24891 11517 24957 11533
rect 24891 11453 24892 11517
rect 24956 11453 24957 11517
rect 24891 11437 24957 11453
rect 24891 11373 24892 11437
rect 24956 11373 24957 11437
rect 24891 11357 24957 11373
rect 24891 11293 24892 11357
rect 24956 11293 24957 11357
rect 24891 11277 24957 11293
rect 24891 11213 24892 11277
rect 24956 11213 24957 11277
rect 24891 11123 24957 11213
rect 25017 11059 25077 12089
rect 25137 11119 25197 12151
rect 25257 11059 25317 12089
rect 25377 11119 25437 12151
rect 25497 11997 25563 12151
rect 25497 11933 25498 11997
rect 25562 11933 25563 11997
rect 25497 11917 25563 11933
rect 25497 11853 25498 11917
rect 25562 11853 25563 11917
rect 25497 11837 25563 11853
rect 25497 11773 25498 11837
rect 25562 11773 25563 11837
rect 25497 11757 25563 11773
rect 25497 11693 25498 11757
rect 25562 11693 25563 11757
rect 25497 11677 25563 11693
rect 25497 11613 25498 11677
rect 25562 11613 25563 11677
rect 25497 11597 25563 11613
rect 25497 11533 25498 11597
rect 25562 11533 25563 11597
rect 25497 11517 25563 11533
rect 25497 11453 25498 11517
rect 25562 11453 25563 11517
rect 25497 11437 25563 11453
rect 25497 11373 25498 11437
rect 25562 11373 25563 11437
rect 25497 11357 25563 11373
rect 25497 11293 25498 11357
rect 25562 11293 25563 11357
rect 25497 11277 25563 11293
rect 25497 11213 25498 11277
rect 25562 11213 25563 11277
rect 25497 11123 25563 11213
rect 25625 12217 25735 12219
rect 25799 12219 25808 12240
rect 26448 12241 26574 12251
rect 25799 12217 26297 12219
rect 25625 12153 25729 12217
rect 25799 12176 25809 12217
rect 25793 12153 25809 12176
rect 25873 12153 25889 12217
rect 25953 12153 25969 12217
rect 26033 12153 26049 12217
rect 26113 12153 26129 12217
rect 26193 12153 26297 12217
rect 26448 12177 26479 12241
rect 26543 12177 26574 12241
rect 26448 12167 26574 12177
rect 26474 12166 26548 12167
rect 25625 12151 26297 12153
rect 25625 11997 25691 12151
rect 25625 11933 25626 11997
rect 25690 11933 25691 11997
rect 25625 11917 25691 11933
rect 25625 11853 25626 11917
rect 25690 11853 25691 11917
rect 25625 11837 25691 11853
rect 25625 11773 25626 11837
rect 25690 11773 25691 11837
rect 25625 11757 25691 11773
rect 25625 11693 25626 11757
rect 25690 11693 25691 11757
rect 25625 11677 25691 11693
rect 25625 11613 25626 11677
rect 25690 11613 25691 11677
rect 25625 11597 25691 11613
rect 25625 11533 25626 11597
rect 25690 11533 25691 11597
rect 25625 11517 25691 11533
rect 25625 11453 25626 11517
rect 25690 11453 25691 11517
rect 25625 11437 25691 11453
rect 25625 11373 25626 11437
rect 25690 11373 25691 11437
rect 25625 11357 25691 11373
rect 25625 11293 25626 11357
rect 25690 11293 25691 11357
rect 25625 11277 25691 11293
rect 25625 11213 25626 11277
rect 25690 11213 25691 11277
rect 25625 11123 25691 11213
rect 25751 11059 25811 12089
rect 25871 11119 25931 12151
rect 25991 11059 26051 12089
rect 26111 11119 26171 12151
rect 26231 11997 26297 12151
rect 26231 11933 26232 11997
rect 26296 11933 26297 11997
rect 26231 11917 26297 11933
rect 26231 11853 26232 11917
rect 26296 11853 26297 11917
rect 26358 11979 26483 11989
rect 26358 11915 26388 11979
rect 26452 11915 26483 11979
rect 26358 11905 26483 11915
rect 26231 11837 26297 11853
rect 26231 11773 26232 11837
rect 26296 11773 26297 11837
rect 26231 11757 26297 11773
rect 26231 11693 26232 11757
rect 26296 11693 26297 11757
rect 26231 11677 26297 11693
rect 26231 11613 26232 11677
rect 26296 11613 26297 11677
rect 26231 11597 26297 11613
rect 26231 11533 26232 11597
rect 26296 11533 26297 11597
rect 26231 11517 26297 11533
rect 26231 11453 26232 11517
rect 26296 11453 26297 11517
rect 26231 11437 26297 11453
rect 26231 11373 26232 11437
rect 26296 11373 26297 11437
rect 26231 11357 26297 11373
rect 26231 11293 26232 11357
rect 26296 11293 26297 11357
rect 26231 11277 26297 11293
rect 26231 11213 26232 11277
rect 26296 11213 26297 11277
rect 26231 11123 26297 11213
rect 13906 10980 14031 10990
rect 20615 10990 20645 11054
rect 20709 10990 20740 11054
rect 21003 11057 21675 11059
rect 21003 10993 21187 11057
rect 21251 10993 21267 11057
rect 21331 10993 21347 11057
rect 21411 10993 21427 11057
rect 21491 10993 21675 11057
rect 21003 10991 21675 10993
rect 21735 11057 24225 11059
rect 21735 10993 21919 11057
rect 21983 10993 21999 11057
rect 22063 10993 22079 11057
rect 22143 10993 22159 11057
rect 22223 10993 22525 11057
rect 22589 10993 22605 11057
rect 22669 10993 22685 11057
rect 22749 10993 22765 11057
rect 22829 10993 23131 11057
rect 23195 10993 23211 11057
rect 23275 10993 23291 11057
rect 23355 10993 23371 11057
rect 23435 10993 23737 11057
rect 23801 10993 23817 11057
rect 23881 10993 23897 11057
rect 23961 10993 23977 11057
rect 24041 10993 24225 11057
rect 21735 10991 24225 10993
rect 24285 11057 25563 11059
rect 24285 10993 24469 11057
rect 24533 10993 24549 11057
rect 24613 10993 24629 11057
rect 24693 10993 24709 11057
rect 24773 10993 25075 11057
rect 25139 10993 25155 11057
rect 25219 10993 25235 11057
rect 25299 10993 25315 11057
rect 25379 10993 25563 11057
rect 24285 10991 25563 10993
rect 25625 11057 26297 11059
rect 25625 10993 25809 11057
rect 25873 10993 25889 11057
rect 25953 10993 25969 11057
rect 26033 10993 26049 11057
rect 26113 10993 26297 11057
rect 25625 10991 26297 10993
rect 20615 10980 20740 10990
rect 8634 10962 8700 10978
rect 8634 10898 8635 10962
rect 8699 10898 8700 10962
rect 8634 10882 8700 10898
rect 8634 10818 8635 10882
rect 8699 10818 8700 10882
rect 8634 10802 8700 10818
rect 8634 10738 8635 10802
rect 8699 10738 8700 10802
rect 8634 10648 8700 10738
rect 3018 10515 3048 10579
rect 3112 10515 3143 10579
rect 3406 10582 4078 10584
rect 3406 10518 3590 10582
rect 3654 10518 3670 10582
rect 3734 10518 3750 10582
rect 3814 10518 3830 10582
rect 3894 10518 4078 10582
rect 3406 10516 4078 10518
rect 4138 10582 6628 10584
rect 4138 10518 4322 10582
rect 4386 10518 4402 10582
rect 4466 10518 4482 10582
rect 4546 10518 4562 10582
rect 4626 10518 4928 10582
rect 4992 10518 5008 10582
rect 5072 10518 5088 10582
rect 5152 10518 5168 10582
rect 5232 10518 5534 10582
rect 5598 10518 5614 10582
rect 5678 10518 5694 10582
rect 5758 10518 5774 10582
rect 5838 10518 6140 10582
rect 6204 10518 6220 10582
rect 6284 10518 6300 10582
rect 6364 10518 6380 10582
rect 6444 10518 6628 10582
rect 4138 10516 6628 10518
rect 6688 10582 7966 10584
rect 6688 10518 6872 10582
rect 6936 10518 6952 10582
rect 7016 10518 7032 10582
rect 7096 10518 7112 10582
rect 7176 10518 7478 10582
rect 7542 10518 7558 10582
rect 7622 10518 7638 10582
rect 7702 10518 7718 10582
rect 7782 10518 7966 10582
rect 6688 10516 7966 10518
rect 8028 10582 8700 10584
rect 8028 10518 8212 10582
rect 8276 10518 8292 10582
rect 8356 10518 8372 10582
rect 8436 10518 8452 10582
rect 8516 10518 8700 10582
rect 8028 10516 8700 10518
rect 3018 10505 3143 10515
rect 3018 10131 3143 10141
rect 3018 10067 3048 10131
rect 3112 10067 3143 10131
rect 3018 10057 3143 10067
rect 3406 10128 4078 10130
rect 3406 10064 3590 10128
rect 3654 10064 3670 10128
rect 3734 10064 3750 10128
rect 3814 10064 3830 10128
rect 3894 10064 4078 10128
rect 3406 10062 4078 10064
rect 4138 10128 6628 10130
rect 4138 10064 4322 10128
rect 4386 10064 4402 10128
rect 4466 10064 4482 10128
rect 4546 10064 4562 10128
rect 4626 10064 4928 10128
rect 4992 10064 5008 10128
rect 5072 10064 5088 10128
rect 5152 10064 5168 10128
rect 5232 10064 5534 10128
rect 5598 10064 5614 10128
rect 5678 10064 5694 10128
rect 5758 10064 5774 10128
rect 5838 10064 6140 10128
rect 6204 10064 6220 10128
rect 6284 10064 6300 10128
rect 6364 10064 6380 10128
rect 6444 10064 6628 10128
rect 4138 10062 6628 10064
rect 6688 10128 7966 10130
rect 6688 10064 6872 10128
rect 6936 10064 6952 10128
rect 7016 10064 7032 10128
rect 7096 10064 7112 10128
rect 7176 10064 7478 10128
rect 7542 10064 7558 10128
rect 7622 10064 7638 10128
rect 7702 10064 7718 10128
rect 7782 10064 7966 10128
rect 6688 10062 7966 10064
rect 8028 10128 8700 10130
rect 8028 10064 8212 10128
rect 8276 10064 8292 10128
rect 8356 10064 8372 10128
rect 8436 10064 8452 10128
rect 8516 10064 8700 10128
rect 19148 10119 19273 10129
rect 8028 10062 8700 10064
rect 13591 10116 14263 10118
rect 3406 9908 3472 9998
rect 3406 9844 3407 9908
rect 3471 9844 3472 9908
rect 3406 9828 3472 9844
rect 3406 9764 3407 9828
rect 3471 9764 3472 9828
rect 3406 9748 3472 9764
rect 3406 9684 3407 9748
rect 3471 9684 3472 9748
rect 3406 9668 3472 9684
rect 3406 9604 3407 9668
rect 3471 9604 3472 9668
rect 3406 9588 3472 9604
rect 3406 9524 3407 9588
rect 3471 9524 3472 9588
rect 3406 9508 3472 9524
rect 3406 9444 3407 9508
rect 3471 9444 3472 9508
rect 3406 9428 3472 9444
rect 3406 9364 3407 9428
rect 3471 9364 3472 9428
rect 3406 9348 3472 9364
rect 3406 9284 3407 9348
rect 3471 9284 3472 9348
rect 3406 9268 3472 9284
rect 3406 9204 3407 9268
rect 3471 9204 3472 9268
rect 3406 9188 3472 9204
rect 3406 9124 3407 9188
rect 3471 9124 3472 9188
rect 3406 8970 3472 9124
rect 3532 8970 3592 10002
rect 3652 9032 3712 10062
rect 3772 8970 3832 10002
rect 3892 9032 3952 10062
rect 4012 9908 4078 9998
rect 4012 9844 4013 9908
rect 4077 9844 4078 9908
rect 4012 9828 4078 9844
rect 4012 9764 4013 9828
rect 4077 9764 4078 9828
rect 4012 9748 4078 9764
rect 4012 9684 4013 9748
rect 4077 9684 4078 9748
rect 4012 9668 4078 9684
rect 4012 9604 4013 9668
rect 4077 9604 4078 9668
rect 4012 9588 4078 9604
rect 4012 9524 4013 9588
rect 4077 9524 4078 9588
rect 4012 9508 4078 9524
rect 4012 9444 4013 9508
rect 4077 9444 4078 9508
rect 4012 9428 4078 9444
rect 4012 9364 4013 9428
rect 4077 9364 4078 9428
rect 4012 9348 4078 9364
rect 4012 9284 4013 9348
rect 4077 9284 4078 9348
rect 4012 9268 4078 9284
rect 4012 9204 4013 9268
rect 4077 9204 4078 9268
rect 4012 9188 4078 9204
rect 4012 9124 4013 9188
rect 4077 9124 4078 9188
rect 4012 8970 4078 9124
rect 3406 8968 4078 8970
rect 3406 8904 3510 8968
rect 3574 8904 3590 8968
rect 3654 8904 3670 8968
rect 3734 8904 3750 8968
rect 3814 8904 3830 8968
rect 3894 8945 3910 8968
rect 3894 8904 3904 8945
rect 3974 8904 4078 8968
rect 3406 8902 3904 8904
rect 3895 8881 3904 8902
rect 3968 8902 4078 8904
rect 4138 9908 4204 9998
rect 4138 9844 4139 9908
rect 4203 9844 4204 9908
rect 4138 9828 4204 9844
rect 4138 9764 4139 9828
rect 4203 9764 4204 9828
rect 4138 9748 4204 9764
rect 4138 9684 4139 9748
rect 4203 9684 4204 9748
rect 4138 9668 4204 9684
rect 4138 9604 4139 9668
rect 4203 9604 4204 9668
rect 4138 9588 4204 9604
rect 4138 9524 4139 9588
rect 4203 9524 4204 9588
rect 4138 9508 4204 9524
rect 4138 9444 4139 9508
rect 4203 9444 4204 9508
rect 4138 9428 4204 9444
rect 4138 9364 4139 9428
rect 4203 9364 4204 9428
rect 4138 9348 4204 9364
rect 4138 9284 4139 9348
rect 4203 9284 4204 9348
rect 4138 9268 4204 9284
rect 4138 9204 4139 9268
rect 4203 9204 4204 9268
rect 4138 9188 4204 9204
rect 4138 9124 4139 9188
rect 4203 9124 4204 9188
rect 4138 8970 4204 9124
rect 4264 8970 4324 10002
rect 4384 9032 4444 10062
rect 4504 8970 4564 10002
rect 4624 9032 4684 10062
rect 4744 9908 4810 9998
rect 4744 9844 4745 9908
rect 4809 9844 4810 9908
rect 4744 9828 4810 9844
rect 4744 9764 4745 9828
rect 4809 9764 4810 9828
rect 4744 9748 4810 9764
rect 4744 9684 4745 9748
rect 4809 9684 4810 9748
rect 4744 9668 4810 9684
rect 4744 9604 4745 9668
rect 4809 9604 4810 9668
rect 4744 9588 4810 9604
rect 4744 9524 4745 9588
rect 4809 9524 4810 9588
rect 4744 9508 4810 9524
rect 4744 9444 4745 9508
rect 4809 9444 4810 9508
rect 4744 9428 4810 9444
rect 4744 9364 4745 9428
rect 4809 9364 4810 9428
rect 4744 9348 4810 9364
rect 4744 9284 4745 9348
rect 4809 9284 4810 9348
rect 4744 9268 4810 9284
rect 4744 9204 4745 9268
rect 4809 9204 4810 9268
rect 4744 9188 4810 9204
rect 4744 9124 4745 9188
rect 4809 9124 4810 9188
rect 4744 8970 4810 9124
rect 4870 9032 4930 10062
rect 4990 8970 5050 10002
rect 5110 9032 5170 10062
rect 5230 8970 5290 10002
rect 5350 9908 5416 9998
rect 5350 9844 5351 9908
rect 5415 9844 5416 9908
rect 5350 9828 5416 9844
rect 5350 9764 5351 9828
rect 5415 9764 5416 9828
rect 5350 9748 5416 9764
rect 5350 9684 5351 9748
rect 5415 9684 5416 9748
rect 5350 9668 5416 9684
rect 5350 9604 5351 9668
rect 5415 9604 5416 9668
rect 5350 9588 5416 9604
rect 5350 9524 5351 9588
rect 5415 9524 5416 9588
rect 5350 9508 5416 9524
rect 5350 9444 5351 9508
rect 5415 9444 5416 9508
rect 5350 9428 5416 9444
rect 5350 9364 5351 9428
rect 5415 9364 5416 9428
rect 5350 9348 5416 9364
rect 5350 9284 5351 9348
rect 5415 9284 5416 9348
rect 5350 9268 5416 9284
rect 5350 9204 5351 9268
rect 5415 9204 5416 9268
rect 5350 9188 5416 9204
rect 5350 9124 5351 9188
rect 5415 9124 5416 9188
rect 5350 8970 5416 9124
rect 5476 8970 5536 10002
rect 5596 9032 5656 10062
rect 5716 8970 5776 10002
rect 5836 9032 5896 10062
rect 5956 9908 6022 9998
rect 5956 9844 5957 9908
rect 6021 9844 6022 9908
rect 5956 9828 6022 9844
rect 5956 9764 5957 9828
rect 6021 9764 6022 9828
rect 5956 9748 6022 9764
rect 5956 9684 5957 9748
rect 6021 9684 6022 9748
rect 5956 9668 6022 9684
rect 5956 9604 5957 9668
rect 6021 9604 6022 9668
rect 5956 9588 6022 9604
rect 5956 9524 5957 9588
rect 6021 9524 6022 9588
rect 5956 9508 6022 9524
rect 5956 9444 5957 9508
rect 6021 9444 6022 9508
rect 5956 9428 6022 9444
rect 5956 9364 5957 9428
rect 6021 9364 6022 9428
rect 5956 9348 6022 9364
rect 5956 9284 5957 9348
rect 6021 9284 6022 9348
rect 5956 9268 6022 9284
rect 5956 9204 5957 9268
rect 6021 9204 6022 9268
rect 5956 9188 6022 9204
rect 5956 9124 5957 9188
rect 6021 9124 6022 9188
rect 5956 8970 6022 9124
rect 6082 9032 6142 10062
rect 6202 8970 6262 10002
rect 6322 9032 6382 10062
rect 6442 8970 6502 10002
rect 6562 9908 6628 9998
rect 6562 9844 6563 9908
rect 6627 9844 6628 9908
rect 6562 9828 6628 9844
rect 6562 9764 6563 9828
rect 6627 9764 6628 9828
rect 6562 9748 6628 9764
rect 6562 9684 6563 9748
rect 6627 9684 6628 9748
rect 6562 9668 6628 9684
rect 6562 9604 6563 9668
rect 6627 9604 6628 9668
rect 6562 9588 6628 9604
rect 6562 9524 6563 9588
rect 6627 9524 6628 9588
rect 6562 9508 6628 9524
rect 6562 9444 6563 9508
rect 6627 9444 6628 9508
rect 6562 9428 6628 9444
rect 6562 9364 6563 9428
rect 6627 9364 6628 9428
rect 6562 9348 6628 9364
rect 6562 9284 6563 9348
rect 6627 9284 6628 9348
rect 6562 9268 6628 9284
rect 6562 9204 6563 9268
rect 6627 9204 6628 9268
rect 6562 9188 6628 9204
rect 6562 9124 6563 9188
rect 6627 9124 6628 9188
rect 6562 8970 6628 9124
rect 4138 8968 6628 8970
rect 4138 8904 4242 8968
rect 4306 8904 4322 8968
rect 4386 8904 4402 8968
rect 4466 8904 4482 8968
rect 4546 8904 4562 8968
rect 4626 8945 4642 8968
rect 4626 8904 4636 8945
rect 4706 8904 4848 8968
rect 4912 8945 4928 8968
rect 4918 8904 4928 8945
rect 4992 8904 5008 8968
rect 5072 8904 5088 8968
rect 5152 8904 5168 8968
rect 5232 8904 5248 8968
rect 5312 8904 5454 8968
rect 5518 8904 5534 8968
rect 5598 8904 5614 8968
rect 5678 8904 5694 8968
rect 5758 8904 5774 8968
rect 5838 8945 5854 8968
rect 5838 8904 5848 8945
rect 5918 8904 6060 8968
rect 6124 8945 6140 8968
rect 6130 8904 6140 8945
rect 6204 8904 6220 8968
rect 6284 8904 6300 8968
rect 6364 8904 6380 8968
rect 6444 8904 6460 8968
rect 6524 8904 6628 8968
rect 4138 8902 4636 8904
rect 3968 8881 3977 8902
rect 3895 8875 3977 8881
rect 4627 8881 4636 8902
rect 4700 8902 4854 8904
rect 4700 8881 4709 8902
rect 4627 8875 4709 8881
rect 4845 8881 4854 8902
rect 4918 8902 5848 8904
rect 4918 8881 4927 8902
rect 4845 8875 4927 8881
rect 5839 8881 5848 8902
rect 5912 8902 6066 8904
rect 5912 8881 5921 8902
rect 5839 8875 5921 8881
rect 6057 8881 6066 8902
rect 6130 8902 6628 8904
rect 6688 9908 6754 9998
rect 6688 9844 6689 9908
rect 6753 9844 6754 9908
rect 6688 9828 6754 9844
rect 6688 9764 6689 9828
rect 6753 9764 6754 9828
rect 6688 9748 6754 9764
rect 6688 9684 6689 9748
rect 6753 9684 6754 9748
rect 6688 9668 6754 9684
rect 6688 9604 6689 9668
rect 6753 9604 6754 9668
rect 6688 9588 6754 9604
rect 6688 9524 6689 9588
rect 6753 9524 6754 9588
rect 6688 9508 6754 9524
rect 6688 9444 6689 9508
rect 6753 9444 6754 9508
rect 6688 9428 6754 9444
rect 6688 9364 6689 9428
rect 6753 9364 6754 9428
rect 6688 9348 6754 9364
rect 6688 9284 6689 9348
rect 6753 9284 6754 9348
rect 6688 9268 6754 9284
rect 6688 9204 6689 9268
rect 6753 9204 6754 9268
rect 6688 9188 6754 9204
rect 6688 9124 6689 9188
rect 6753 9124 6754 9188
rect 6688 8970 6754 9124
rect 6814 8970 6874 10002
rect 6934 9032 6994 10062
rect 7054 8970 7114 10002
rect 7174 9032 7234 10062
rect 7294 9908 7360 9998
rect 7294 9844 7295 9908
rect 7359 9844 7360 9908
rect 7294 9828 7360 9844
rect 7294 9764 7295 9828
rect 7359 9764 7360 9828
rect 7294 9748 7360 9764
rect 7294 9684 7295 9748
rect 7359 9684 7360 9748
rect 7294 9668 7360 9684
rect 7294 9604 7295 9668
rect 7359 9604 7360 9668
rect 7294 9588 7360 9604
rect 7294 9524 7295 9588
rect 7359 9524 7360 9588
rect 7294 9508 7360 9524
rect 7294 9444 7295 9508
rect 7359 9444 7360 9508
rect 7294 9428 7360 9444
rect 7294 9364 7295 9428
rect 7359 9364 7360 9428
rect 7294 9348 7360 9364
rect 7294 9284 7295 9348
rect 7359 9284 7360 9348
rect 7294 9268 7360 9284
rect 7294 9204 7295 9268
rect 7359 9204 7360 9268
rect 7294 9188 7360 9204
rect 7294 9124 7295 9188
rect 7359 9124 7360 9188
rect 7294 8970 7360 9124
rect 7420 9032 7480 10062
rect 7540 8970 7600 10002
rect 7660 9032 7720 10062
rect 7780 8970 7840 10002
rect 7900 9908 7966 9998
rect 7900 9844 7901 9908
rect 7965 9844 7966 9908
rect 7900 9828 7966 9844
rect 7900 9764 7901 9828
rect 7965 9764 7966 9828
rect 7900 9748 7966 9764
rect 7900 9684 7901 9748
rect 7965 9684 7966 9748
rect 7900 9668 7966 9684
rect 7900 9604 7901 9668
rect 7965 9604 7966 9668
rect 7900 9588 7966 9604
rect 7900 9524 7901 9588
rect 7965 9524 7966 9588
rect 7900 9508 7966 9524
rect 7900 9444 7901 9508
rect 7965 9444 7966 9508
rect 7900 9428 7966 9444
rect 7900 9364 7901 9428
rect 7965 9364 7966 9428
rect 7900 9348 7966 9364
rect 7900 9284 7901 9348
rect 7965 9284 7966 9348
rect 7900 9268 7966 9284
rect 7900 9204 7901 9268
rect 7965 9204 7966 9268
rect 7900 9188 7966 9204
rect 7900 9124 7901 9188
rect 7965 9124 7966 9188
rect 7900 8970 7966 9124
rect 6688 8968 7966 8970
rect 6688 8904 6792 8968
rect 6856 8904 6872 8968
rect 6936 8904 6952 8968
rect 7016 8904 7032 8968
rect 7096 8904 7112 8968
rect 7176 8945 7192 8968
rect 7176 8904 7186 8945
rect 7256 8904 7398 8968
rect 7462 8945 7478 8968
rect 7468 8904 7478 8945
rect 7542 8904 7558 8968
rect 7622 8904 7638 8968
rect 7702 8904 7718 8968
rect 7782 8904 7798 8968
rect 7862 8904 7966 8968
rect 6688 8902 7186 8904
rect 6130 8881 6139 8902
rect 6057 8875 6139 8881
rect 7177 8881 7186 8902
rect 7250 8902 7404 8904
rect 7250 8881 7259 8902
rect 7177 8875 7259 8881
rect 7395 8881 7404 8902
rect 7468 8902 7966 8904
rect 8028 9908 8094 9998
rect 8028 9844 8029 9908
rect 8093 9844 8094 9908
rect 8028 9828 8094 9844
rect 8028 9764 8029 9828
rect 8093 9764 8094 9828
rect 8028 9748 8094 9764
rect 8028 9684 8029 9748
rect 8093 9684 8094 9748
rect 8028 9668 8094 9684
rect 8028 9604 8029 9668
rect 8093 9604 8094 9668
rect 8028 9588 8094 9604
rect 8028 9524 8029 9588
rect 8093 9524 8094 9588
rect 8028 9508 8094 9524
rect 8028 9444 8029 9508
rect 8093 9444 8094 9508
rect 8028 9428 8094 9444
rect 8028 9364 8029 9428
rect 8093 9364 8094 9428
rect 8028 9348 8094 9364
rect 8028 9284 8029 9348
rect 8093 9284 8094 9348
rect 8028 9268 8094 9284
rect 8028 9204 8029 9268
rect 8093 9204 8094 9268
rect 8028 9188 8094 9204
rect 8028 9124 8029 9188
rect 8093 9124 8094 9188
rect 8028 8970 8094 9124
rect 8154 9032 8214 10062
rect 8274 8970 8334 10002
rect 8394 9032 8454 10062
rect 13591 10052 13775 10116
rect 13839 10052 13855 10116
rect 13919 10052 13935 10116
rect 13999 10052 14015 10116
rect 14079 10052 14263 10116
rect 13591 10050 14263 10052
rect 14325 10116 15603 10118
rect 14325 10052 14509 10116
rect 14573 10052 14589 10116
rect 14653 10052 14669 10116
rect 14733 10052 14749 10116
rect 14813 10052 15115 10116
rect 15179 10052 15195 10116
rect 15259 10052 15275 10116
rect 15339 10052 15355 10116
rect 15419 10052 15603 10116
rect 14325 10050 15603 10052
rect 15663 10116 18153 10118
rect 15663 10052 15847 10116
rect 15911 10052 15927 10116
rect 15991 10052 16007 10116
rect 16071 10052 16087 10116
rect 16151 10052 16453 10116
rect 16517 10052 16533 10116
rect 16597 10052 16613 10116
rect 16677 10052 16693 10116
rect 16757 10052 17059 10116
rect 17123 10052 17139 10116
rect 17203 10052 17219 10116
rect 17283 10052 17299 10116
rect 17363 10052 17665 10116
rect 17729 10052 17745 10116
rect 17809 10052 17825 10116
rect 17889 10052 17905 10116
rect 17969 10052 18153 10116
rect 15663 10050 18153 10052
rect 18213 10116 18885 10118
rect 18213 10052 18397 10116
rect 18461 10052 18477 10116
rect 18541 10052 18557 10116
rect 18621 10052 18637 10116
rect 18701 10052 18885 10116
rect 18213 10050 18885 10052
rect 19148 10055 19179 10119
rect 19243 10055 19273 10119
rect 25857 10119 25982 10129
rect 8514 8970 8574 10002
rect 8634 9908 8700 9998
rect 8634 9844 8635 9908
rect 8699 9844 8700 9908
rect 8634 9828 8700 9844
rect 8634 9764 8635 9828
rect 8699 9764 8700 9828
rect 8634 9748 8700 9764
rect 8634 9684 8635 9748
rect 8699 9684 8700 9748
rect 8634 9668 8700 9684
rect 8634 9604 8635 9668
rect 8699 9604 8700 9668
rect 8634 9588 8700 9604
rect 8634 9524 8635 9588
rect 8699 9524 8700 9588
rect 8634 9508 8700 9524
rect 8634 9444 8635 9508
rect 8699 9444 8700 9508
rect 8634 9428 8700 9444
rect 8634 9364 8635 9428
rect 8699 9364 8700 9428
rect 8634 9348 8700 9364
rect 8634 9284 8635 9348
rect 8699 9284 8700 9348
rect 8634 9268 8700 9284
rect 8634 9204 8635 9268
rect 8699 9204 8700 9268
rect 13591 9896 13657 9986
rect 13591 9832 13592 9896
rect 13656 9832 13657 9896
rect 13591 9816 13657 9832
rect 13591 9752 13592 9816
rect 13656 9752 13657 9816
rect 13591 9736 13657 9752
rect 13591 9672 13592 9736
rect 13656 9672 13657 9736
rect 13591 9656 13657 9672
rect 13591 9592 13592 9656
rect 13656 9592 13657 9656
rect 13591 9576 13657 9592
rect 13591 9512 13592 9576
rect 13656 9512 13657 9576
rect 13591 9496 13657 9512
rect 13591 9432 13592 9496
rect 13656 9432 13657 9496
rect 13591 9416 13657 9432
rect 13591 9352 13592 9416
rect 13656 9352 13657 9416
rect 13591 9336 13657 9352
rect 13591 9272 13592 9336
rect 13656 9272 13657 9336
rect 13591 9256 13657 9272
rect 8634 9188 8700 9204
rect 8634 9124 8635 9188
rect 8699 9124 8700 9188
rect 8761 9206 8886 9216
rect 8761 9142 8791 9206
rect 8855 9142 8886 9206
rect 13405 9194 13530 9204
rect 8761 9132 8886 9142
rect 9189 9165 9314 9175
rect 8634 8970 8700 9124
rect 9189 9101 9219 9165
rect 9283 9101 9314 9165
rect 9189 9092 9314 9101
rect 9666 9165 9791 9175
rect 9666 9101 9696 9165
rect 9760 9101 9791 9165
rect 9666 9092 9791 9101
rect 10086 9154 10211 9164
rect 10086 9090 10116 9154
rect 10180 9090 10211 9154
rect 10086 9081 10211 9090
rect 10462 9162 10587 9172
rect 10462 9098 10492 9162
rect 10556 9098 10587 9162
rect 10462 9089 10587 9098
rect 10810 9162 10935 9172
rect 10810 9098 10840 9162
rect 10904 9098 10935 9162
rect 10810 9089 10935 9098
rect 11068 9168 11193 9178
rect 11068 9104 11098 9168
rect 11162 9104 11193 9168
rect 11068 9095 11193 9104
rect 11294 9168 11419 9178
rect 11294 9104 11324 9168
rect 11388 9104 11419 9168
rect 11294 9095 11419 9104
rect 11553 9171 11678 9181
rect 11553 9107 11583 9171
rect 11647 9107 11678 9171
rect 11553 9098 11678 9107
rect 12160 9133 12285 9143
rect 12160 9069 12190 9133
rect 12254 9069 12285 9133
rect 12160 9059 12285 9069
rect 12392 9134 12517 9144
rect 12392 9070 12422 9134
rect 12486 9070 12517 9134
rect 12392 9060 12517 9070
rect 12828 9140 12953 9150
rect 12828 9076 12858 9140
rect 12922 9076 12953 9140
rect 12828 9066 12953 9076
rect 13063 9142 13188 9152
rect 13063 9078 13093 9142
rect 13157 9078 13188 9142
rect 13405 9130 13436 9194
rect 13500 9130 13530 9194
rect 13405 9120 13530 9130
rect 13591 9192 13592 9256
rect 13656 9192 13657 9256
rect 13591 9176 13657 9192
rect 13063 9068 13188 9078
rect 13591 9112 13592 9176
rect 13656 9112 13657 9176
rect 8028 8968 8700 8970
rect 8028 8904 8132 8968
rect 8196 8945 8212 8968
rect 8202 8904 8212 8945
rect 8276 8904 8292 8968
rect 8356 8904 8372 8968
rect 8436 8904 8452 8968
rect 8516 8904 8532 8968
rect 8596 8904 8700 8968
rect 13591 8958 13657 9112
rect 13717 8958 13777 9990
rect 13837 9020 13897 10050
rect 13957 8958 14017 9990
rect 14077 9020 14137 10050
rect 14197 9896 14263 9986
rect 14197 9832 14198 9896
rect 14262 9832 14263 9896
rect 14197 9816 14263 9832
rect 14197 9752 14198 9816
rect 14262 9752 14263 9816
rect 14197 9736 14263 9752
rect 14197 9672 14198 9736
rect 14262 9672 14263 9736
rect 14197 9656 14263 9672
rect 14197 9592 14198 9656
rect 14262 9592 14263 9656
rect 14197 9576 14263 9592
rect 14197 9512 14198 9576
rect 14262 9512 14263 9576
rect 14197 9496 14263 9512
rect 14197 9432 14198 9496
rect 14262 9432 14263 9496
rect 14197 9416 14263 9432
rect 14197 9352 14198 9416
rect 14262 9352 14263 9416
rect 14197 9336 14263 9352
rect 14197 9272 14198 9336
rect 14262 9272 14263 9336
rect 14197 9256 14263 9272
rect 14197 9192 14198 9256
rect 14262 9192 14263 9256
rect 14197 9176 14263 9192
rect 14197 9112 14198 9176
rect 14262 9112 14263 9176
rect 14197 8958 14263 9112
rect 13591 8956 14263 8958
rect 8877 8954 8951 8955
rect 8028 8902 8138 8904
rect 7468 8881 7477 8902
rect 7395 8875 7477 8881
rect 8129 8881 8138 8902
rect 8202 8902 8700 8904
rect 8851 8944 8977 8954
rect 8202 8881 8211 8902
rect 8129 8875 8211 8881
rect 8851 8880 8882 8944
rect 8946 8880 8977 8944
rect 13340 8942 13414 8943
rect 8851 8870 8977 8880
rect 13314 8932 13440 8942
rect 13314 8868 13345 8932
rect 13409 8868 13440 8932
rect 13591 8892 13695 8956
rect 13759 8892 13775 8956
rect 13839 8892 13855 8956
rect 13919 8892 13935 8956
rect 13999 8892 14015 8956
rect 14079 8933 14095 8956
rect 14079 8892 14089 8933
rect 14159 8892 14263 8956
rect 13591 8890 14089 8892
rect 13314 8858 13440 8868
rect 14080 8869 14089 8890
rect 14153 8890 14263 8892
rect 14325 9896 14391 9986
rect 14325 9832 14326 9896
rect 14390 9832 14391 9896
rect 14325 9816 14391 9832
rect 14325 9752 14326 9816
rect 14390 9752 14391 9816
rect 14325 9736 14391 9752
rect 14325 9672 14326 9736
rect 14390 9672 14391 9736
rect 14325 9656 14391 9672
rect 14325 9592 14326 9656
rect 14390 9592 14391 9656
rect 14325 9576 14391 9592
rect 14325 9512 14326 9576
rect 14390 9512 14391 9576
rect 14325 9496 14391 9512
rect 14325 9432 14326 9496
rect 14390 9432 14391 9496
rect 14325 9416 14391 9432
rect 14325 9352 14326 9416
rect 14390 9352 14391 9416
rect 14325 9336 14391 9352
rect 14325 9272 14326 9336
rect 14390 9272 14391 9336
rect 14325 9256 14391 9272
rect 14325 9192 14326 9256
rect 14390 9192 14391 9256
rect 14325 9176 14391 9192
rect 14325 9112 14326 9176
rect 14390 9112 14391 9176
rect 14325 8958 14391 9112
rect 14451 8958 14511 9990
rect 14571 9020 14631 10050
rect 14691 8958 14751 9990
rect 14811 9020 14871 10050
rect 14931 9896 14997 9986
rect 14931 9832 14932 9896
rect 14996 9832 14997 9896
rect 14931 9816 14997 9832
rect 14931 9752 14932 9816
rect 14996 9752 14997 9816
rect 14931 9736 14997 9752
rect 14931 9672 14932 9736
rect 14996 9672 14997 9736
rect 14931 9656 14997 9672
rect 14931 9592 14932 9656
rect 14996 9592 14997 9656
rect 14931 9576 14997 9592
rect 14931 9512 14932 9576
rect 14996 9512 14997 9576
rect 14931 9496 14997 9512
rect 14931 9432 14932 9496
rect 14996 9432 14997 9496
rect 14931 9416 14997 9432
rect 14931 9352 14932 9416
rect 14996 9352 14997 9416
rect 14931 9336 14997 9352
rect 14931 9272 14932 9336
rect 14996 9272 14997 9336
rect 14931 9256 14997 9272
rect 14931 9192 14932 9256
rect 14996 9192 14997 9256
rect 14931 9176 14997 9192
rect 14931 9112 14932 9176
rect 14996 9112 14997 9176
rect 14931 8958 14997 9112
rect 15057 9020 15117 10050
rect 15177 8958 15237 9990
rect 15297 9020 15357 10050
rect 15417 8958 15477 9990
rect 15537 9896 15603 9986
rect 15537 9832 15538 9896
rect 15602 9832 15603 9896
rect 15537 9816 15603 9832
rect 15537 9752 15538 9816
rect 15602 9752 15603 9816
rect 15537 9736 15603 9752
rect 15537 9672 15538 9736
rect 15602 9672 15603 9736
rect 15537 9656 15603 9672
rect 15537 9592 15538 9656
rect 15602 9592 15603 9656
rect 15537 9576 15603 9592
rect 15537 9512 15538 9576
rect 15602 9512 15603 9576
rect 15537 9496 15603 9512
rect 15537 9432 15538 9496
rect 15602 9432 15603 9496
rect 15537 9416 15603 9432
rect 15537 9352 15538 9416
rect 15602 9352 15603 9416
rect 15537 9336 15603 9352
rect 15537 9272 15538 9336
rect 15602 9272 15603 9336
rect 15537 9256 15603 9272
rect 15537 9192 15538 9256
rect 15602 9192 15603 9256
rect 15537 9176 15603 9192
rect 15537 9112 15538 9176
rect 15602 9112 15603 9176
rect 15537 8958 15603 9112
rect 14325 8956 15603 8958
rect 14325 8892 14429 8956
rect 14493 8892 14509 8956
rect 14573 8892 14589 8956
rect 14653 8892 14669 8956
rect 14733 8892 14749 8956
rect 14813 8933 14829 8956
rect 14813 8892 14823 8933
rect 14893 8892 15035 8956
rect 15099 8933 15115 8956
rect 15105 8892 15115 8933
rect 15179 8892 15195 8956
rect 15259 8892 15275 8956
rect 15339 8892 15355 8956
rect 15419 8892 15435 8956
rect 15499 8892 15603 8956
rect 14325 8890 14823 8892
rect 14153 8869 14162 8890
rect 14080 8863 14162 8869
rect 14814 8869 14823 8890
rect 14887 8890 15041 8892
rect 14887 8869 14896 8890
rect 14814 8863 14896 8869
rect 15032 8869 15041 8890
rect 15105 8890 15603 8892
rect 15663 9896 15729 9986
rect 15663 9832 15664 9896
rect 15728 9832 15729 9896
rect 15663 9816 15729 9832
rect 15663 9752 15664 9816
rect 15728 9752 15729 9816
rect 15663 9736 15729 9752
rect 15663 9672 15664 9736
rect 15728 9672 15729 9736
rect 15663 9656 15729 9672
rect 15663 9592 15664 9656
rect 15728 9592 15729 9656
rect 15663 9576 15729 9592
rect 15663 9512 15664 9576
rect 15728 9512 15729 9576
rect 15663 9496 15729 9512
rect 15663 9432 15664 9496
rect 15728 9432 15729 9496
rect 15663 9416 15729 9432
rect 15663 9352 15664 9416
rect 15728 9352 15729 9416
rect 15663 9336 15729 9352
rect 15663 9272 15664 9336
rect 15728 9272 15729 9336
rect 15663 9256 15729 9272
rect 15663 9192 15664 9256
rect 15728 9192 15729 9256
rect 15663 9176 15729 9192
rect 15663 9112 15664 9176
rect 15728 9112 15729 9176
rect 15663 8958 15729 9112
rect 15789 8958 15849 9990
rect 15909 9020 15969 10050
rect 16029 8958 16089 9990
rect 16149 9020 16209 10050
rect 16269 9896 16335 9986
rect 16269 9832 16270 9896
rect 16334 9832 16335 9896
rect 16269 9816 16335 9832
rect 16269 9752 16270 9816
rect 16334 9752 16335 9816
rect 16269 9736 16335 9752
rect 16269 9672 16270 9736
rect 16334 9672 16335 9736
rect 16269 9656 16335 9672
rect 16269 9592 16270 9656
rect 16334 9592 16335 9656
rect 16269 9576 16335 9592
rect 16269 9512 16270 9576
rect 16334 9512 16335 9576
rect 16269 9496 16335 9512
rect 16269 9432 16270 9496
rect 16334 9432 16335 9496
rect 16269 9416 16335 9432
rect 16269 9352 16270 9416
rect 16334 9352 16335 9416
rect 16269 9336 16335 9352
rect 16269 9272 16270 9336
rect 16334 9272 16335 9336
rect 16269 9256 16335 9272
rect 16269 9192 16270 9256
rect 16334 9192 16335 9256
rect 16269 9176 16335 9192
rect 16269 9112 16270 9176
rect 16334 9112 16335 9176
rect 16269 8958 16335 9112
rect 16395 9020 16455 10050
rect 16515 8958 16575 9990
rect 16635 9020 16695 10050
rect 16755 8958 16815 9990
rect 16875 9896 16941 9986
rect 16875 9832 16876 9896
rect 16940 9832 16941 9896
rect 16875 9816 16941 9832
rect 16875 9752 16876 9816
rect 16940 9752 16941 9816
rect 16875 9736 16941 9752
rect 16875 9672 16876 9736
rect 16940 9672 16941 9736
rect 16875 9656 16941 9672
rect 16875 9592 16876 9656
rect 16940 9592 16941 9656
rect 16875 9576 16941 9592
rect 16875 9512 16876 9576
rect 16940 9512 16941 9576
rect 16875 9496 16941 9512
rect 16875 9432 16876 9496
rect 16940 9432 16941 9496
rect 16875 9416 16941 9432
rect 16875 9352 16876 9416
rect 16940 9352 16941 9416
rect 16875 9336 16941 9352
rect 16875 9272 16876 9336
rect 16940 9272 16941 9336
rect 16875 9256 16941 9272
rect 16875 9192 16876 9256
rect 16940 9192 16941 9256
rect 16875 9176 16941 9192
rect 16875 9112 16876 9176
rect 16940 9112 16941 9176
rect 16875 8958 16941 9112
rect 17001 8958 17061 9990
rect 17121 9020 17181 10050
rect 17241 8958 17301 9990
rect 17361 9020 17421 10050
rect 17481 9896 17547 9986
rect 17481 9832 17482 9896
rect 17546 9832 17547 9896
rect 17481 9816 17547 9832
rect 17481 9752 17482 9816
rect 17546 9752 17547 9816
rect 17481 9736 17547 9752
rect 17481 9672 17482 9736
rect 17546 9672 17547 9736
rect 17481 9656 17547 9672
rect 17481 9592 17482 9656
rect 17546 9592 17547 9656
rect 17481 9576 17547 9592
rect 17481 9512 17482 9576
rect 17546 9512 17547 9576
rect 17481 9496 17547 9512
rect 17481 9432 17482 9496
rect 17546 9432 17547 9496
rect 17481 9416 17547 9432
rect 17481 9352 17482 9416
rect 17546 9352 17547 9416
rect 17481 9336 17547 9352
rect 17481 9272 17482 9336
rect 17546 9272 17547 9336
rect 17481 9256 17547 9272
rect 17481 9192 17482 9256
rect 17546 9192 17547 9256
rect 17481 9176 17547 9192
rect 17481 9112 17482 9176
rect 17546 9112 17547 9176
rect 17481 8958 17547 9112
rect 17607 9020 17667 10050
rect 17727 8958 17787 9990
rect 17847 9020 17907 10050
rect 17967 8958 18027 9990
rect 18087 9896 18153 9986
rect 18087 9832 18088 9896
rect 18152 9832 18153 9896
rect 18087 9816 18153 9832
rect 18087 9752 18088 9816
rect 18152 9752 18153 9816
rect 18087 9736 18153 9752
rect 18087 9672 18088 9736
rect 18152 9672 18153 9736
rect 18087 9656 18153 9672
rect 18087 9592 18088 9656
rect 18152 9592 18153 9656
rect 18087 9576 18153 9592
rect 18087 9512 18088 9576
rect 18152 9512 18153 9576
rect 18087 9496 18153 9512
rect 18087 9432 18088 9496
rect 18152 9432 18153 9496
rect 18087 9416 18153 9432
rect 18087 9352 18088 9416
rect 18152 9352 18153 9416
rect 18087 9336 18153 9352
rect 18087 9272 18088 9336
rect 18152 9272 18153 9336
rect 18087 9256 18153 9272
rect 18087 9192 18088 9256
rect 18152 9192 18153 9256
rect 18087 9176 18153 9192
rect 18087 9112 18088 9176
rect 18152 9112 18153 9176
rect 18087 8958 18153 9112
rect 15663 8956 18153 8958
rect 15663 8892 15767 8956
rect 15831 8892 15847 8956
rect 15911 8892 15927 8956
rect 15991 8892 16007 8956
rect 16071 8892 16087 8956
rect 16151 8933 16167 8956
rect 16151 8892 16161 8933
rect 16231 8892 16373 8956
rect 16437 8933 16453 8956
rect 16443 8892 16453 8933
rect 16517 8892 16533 8956
rect 16597 8892 16613 8956
rect 16677 8892 16693 8956
rect 16757 8892 16773 8956
rect 16837 8892 16979 8956
rect 17043 8892 17059 8956
rect 17123 8892 17139 8956
rect 17203 8892 17219 8956
rect 17283 8892 17299 8956
rect 17363 8933 17379 8956
rect 17363 8892 17373 8933
rect 17443 8892 17585 8956
rect 17649 8933 17665 8956
rect 17655 8892 17665 8933
rect 17729 8892 17745 8956
rect 17809 8892 17825 8956
rect 17889 8892 17905 8956
rect 17969 8892 17985 8956
rect 18049 8892 18153 8956
rect 15663 8890 16161 8892
rect 15105 8869 15114 8890
rect 15032 8863 15114 8869
rect 16152 8869 16161 8890
rect 16225 8890 16379 8892
rect 16225 8869 16234 8890
rect 16152 8863 16234 8869
rect 16370 8869 16379 8890
rect 16443 8890 17373 8892
rect 16443 8869 16452 8890
rect 16370 8863 16452 8869
rect 17364 8869 17373 8890
rect 17437 8890 17591 8892
rect 17437 8869 17446 8890
rect 17364 8863 17446 8869
rect 17582 8869 17591 8890
rect 17655 8890 18153 8892
rect 18213 9896 18279 9986
rect 18213 9832 18214 9896
rect 18278 9832 18279 9896
rect 18213 9816 18279 9832
rect 18213 9752 18214 9816
rect 18278 9752 18279 9816
rect 18213 9736 18279 9752
rect 18213 9672 18214 9736
rect 18278 9672 18279 9736
rect 18213 9656 18279 9672
rect 18213 9592 18214 9656
rect 18278 9592 18279 9656
rect 18213 9576 18279 9592
rect 18213 9512 18214 9576
rect 18278 9512 18279 9576
rect 18213 9496 18279 9512
rect 18213 9432 18214 9496
rect 18278 9432 18279 9496
rect 18213 9416 18279 9432
rect 18213 9352 18214 9416
rect 18278 9352 18279 9416
rect 18213 9336 18279 9352
rect 18213 9272 18214 9336
rect 18278 9272 18279 9336
rect 18213 9256 18279 9272
rect 18213 9192 18214 9256
rect 18278 9192 18279 9256
rect 18213 9176 18279 9192
rect 18213 9112 18214 9176
rect 18278 9112 18279 9176
rect 18213 8958 18279 9112
rect 18339 9020 18399 10050
rect 18459 8958 18519 9990
rect 18579 9020 18639 10050
rect 19148 10045 19273 10055
rect 20300 10116 20972 10118
rect 20300 10052 20484 10116
rect 20548 10052 20564 10116
rect 20628 10052 20644 10116
rect 20708 10052 20724 10116
rect 20788 10052 20972 10116
rect 20300 10050 20972 10052
rect 21034 10116 22312 10118
rect 21034 10052 21218 10116
rect 21282 10052 21298 10116
rect 21362 10052 21378 10116
rect 21442 10052 21458 10116
rect 21522 10052 21824 10116
rect 21888 10052 21904 10116
rect 21968 10052 21984 10116
rect 22048 10052 22064 10116
rect 22128 10052 22312 10116
rect 21034 10050 22312 10052
rect 22372 10116 24862 10118
rect 22372 10052 22556 10116
rect 22620 10052 22636 10116
rect 22700 10052 22716 10116
rect 22780 10052 22796 10116
rect 22860 10052 23162 10116
rect 23226 10052 23242 10116
rect 23306 10052 23322 10116
rect 23386 10052 23402 10116
rect 23466 10052 23768 10116
rect 23832 10052 23848 10116
rect 23912 10052 23928 10116
rect 23992 10052 24008 10116
rect 24072 10052 24374 10116
rect 24438 10052 24454 10116
rect 24518 10052 24534 10116
rect 24598 10052 24614 10116
rect 24678 10052 24862 10116
rect 22372 10050 24862 10052
rect 24922 10116 25594 10118
rect 24922 10052 25106 10116
rect 25170 10052 25186 10116
rect 25250 10052 25266 10116
rect 25330 10052 25346 10116
rect 25410 10052 25594 10116
rect 24922 10050 25594 10052
rect 25857 10055 25888 10119
rect 25952 10055 25982 10119
rect 18699 8958 18759 9990
rect 18819 9896 18885 9986
rect 18819 9832 18820 9896
rect 18884 9832 18885 9896
rect 18819 9816 18885 9832
rect 18819 9752 18820 9816
rect 18884 9752 18885 9816
rect 18819 9736 18885 9752
rect 18819 9672 18820 9736
rect 18884 9672 18885 9736
rect 18819 9656 18885 9672
rect 18819 9592 18820 9656
rect 18884 9592 18885 9656
rect 18819 9576 18885 9592
rect 18819 9512 18820 9576
rect 18884 9512 18885 9576
rect 18819 9496 18885 9512
rect 18819 9432 18820 9496
rect 18884 9432 18885 9496
rect 18819 9416 18885 9432
rect 18819 9352 18820 9416
rect 18884 9352 18885 9416
rect 18819 9336 18885 9352
rect 18819 9272 18820 9336
rect 18884 9272 18885 9336
rect 18819 9256 18885 9272
rect 18819 9192 18820 9256
rect 18884 9192 18885 9256
rect 20300 9896 20366 9986
rect 20300 9832 20301 9896
rect 20365 9832 20366 9896
rect 20300 9816 20366 9832
rect 20300 9752 20301 9816
rect 20365 9752 20366 9816
rect 20300 9736 20366 9752
rect 20300 9672 20301 9736
rect 20365 9672 20366 9736
rect 20300 9656 20366 9672
rect 20300 9592 20301 9656
rect 20365 9592 20366 9656
rect 20300 9576 20366 9592
rect 20300 9512 20301 9576
rect 20365 9512 20366 9576
rect 20300 9496 20366 9512
rect 20300 9432 20301 9496
rect 20365 9432 20366 9496
rect 20300 9416 20366 9432
rect 20300 9352 20301 9416
rect 20365 9352 20366 9416
rect 20300 9336 20366 9352
rect 20300 9272 20301 9336
rect 20365 9272 20366 9336
rect 20300 9256 20366 9272
rect 18819 9176 18885 9192
rect 18819 9112 18820 9176
rect 18884 9112 18885 9176
rect 20114 9194 20239 9204
rect 20114 9130 20145 9194
rect 20209 9130 20239 9194
rect 20114 9120 20239 9130
rect 20300 9192 20301 9256
rect 20365 9192 20366 9256
rect 20300 9176 20366 9192
rect 18819 8958 18885 9112
rect 18213 8956 18885 8958
rect 18213 8892 18317 8956
rect 18381 8933 18397 8956
rect 18387 8892 18397 8933
rect 18461 8892 18477 8956
rect 18541 8892 18557 8956
rect 18621 8892 18637 8956
rect 18701 8892 18717 8956
rect 18781 8892 18885 8956
rect 20300 9112 20301 9176
rect 20365 9112 20366 9176
rect 20300 8958 20366 9112
rect 20426 8958 20486 9990
rect 20546 9020 20606 10050
rect 20666 8958 20726 9990
rect 20786 9020 20846 10050
rect 20906 9896 20972 9986
rect 20906 9832 20907 9896
rect 20971 9832 20972 9896
rect 20906 9816 20972 9832
rect 20906 9752 20907 9816
rect 20971 9752 20972 9816
rect 20906 9736 20972 9752
rect 20906 9672 20907 9736
rect 20971 9672 20972 9736
rect 20906 9656 20972 9672
rect 20906 9592 20907 9656
rect 20971 9592 20972 9656
rect 20906 9576 20972 9592
rect 20906 9512 20907 9576
rect 20971 9512 20972 9576
rect 20906 9496 20972 9512
rect 20906 9432 20907 9496
rect 20971 9432 20972 9496
rect 20906 9416 20972 9432
rect 20906 9352 20907 9416
rect 20971 9352 20972 9416
rect 20906 9336 20972 9352
rect 20906 9272 20907 9336
rect 20971 9272 20972 9336
rect 20906 9256 20972 9272
rect 20906 9192 20907 9256
rect 20971 9192 20972 9256
rect 20906 9176 20972 9192
rect 20906 9112 20907 9176
rect 20971 9112 20972 9176
rect 20906 8958 20972 9112
rect 20300 8956 20972 8958
rect 20049 8942 20123 8943
rect 18213 8890 18323 8892
rect 17655 8869 17664 8890
rect 17582 8863 17664 8869
rect 18314 8869 18323 8890
rect 18387 8890 18885 8892
rect 20023 8932 20149 8942
rect 18387 8869 18396 8890
rect 18314 8863 18396 8869
rect 20023 8868 20054 8932
rect 20118 8868 20149 8932
rect 20300 8892 20404 8956
rect 20468 8892 20484 8956
rect 20548 8892 20564 8956
rect 20628 8892 20644 8956
rect 20708 8892 20724 8956
rect 20788 8933 20804 8956
rect 20788 8892 20798 8933
rect 20868 8892 20972 8956
rect 20300 8890 20798 8892
rect 20023 8858 20149 8868
rect 20789 8869 20798 8890
rect 20862 8890 20972 8892
rect 21034 9896 21100 9986
rect 21034 9832 21035 9896
rect 21099 9832 21100 9896
rect 21034 9816 21100 9832
rect 21034 9752 21035 9816
rect 21099 9752 21100 9816
rect 21034 9736 21100 9752
rect 21034 9672 21035 9736
rect 21099 9672 21100 9736
rect 21034 9656 21100 9672
rect 21034 9592 21035 9656
rect 21099 9592 21100 9656
rect 21034 9576 21100 9592
rect 21034 9512 21035 9576
rect 21099 9512 21100 9576
rect 21034 9496 21100 9512
rect 21034 9432 21035 9496
rect 21099 9432 21100 9496
rect 21034 9416 21100 9432
rect 21034 9352 21035 9416
rect 21099 9352 21100 9416
rect 21034 9336 21100 9352
rect 21034 9272 21035 9336
rect 21099 9272 21100 9336
rect 21034 9256 21100 9272
rect 21034 9192 21035 9256
rect 21099 9192 21100 9256
rect 21034 9176 21100 9192
rect 21034 9112 21035 9176
rect 21099 9112 21100 9176
rect 21034 8958 21100 9112
rect 21160 8958 21220 9990
rect 21280 9020 21340 10050
rect 21400 8958 21460 9990
rect 21520 9020 21580 10050
rect 21640 9896 21706 9986
rect 21640 9832 21641 9896
rect 21705 9832 21706 9896
rect 21640 9816 21706 9832
rect 21640 9752 21641 9816
rect 21705 9752 21706 9816
rect 21640 9736 21706 9752
rect 21640 9672 21641 9736
rect 21705 9672 21706 9736
rect 21640 9656 21706 9672
rect 21640 9592 21641 9656
rect 21705 9592 21706 9656
rect 21640 9576 21706 9592
rect 21640 9512 21641 9576
rect 21705 9512 21706 9576
rect 21640 9496 21706 9512
rect 21640 9432 21641 9496
rect 21705 9432 21706 9496
rect 21640 9416 21706 9432
rect 21640 9352 21641 9416
rect 21705 9352 21706 9416
rect 21640 9336 21706 9352
rect 21640 9272 21641 9336
rect 21705 9272 21706 9336
rect 21640 9256 21706 9272
rect 21640 9192 21641 9256
rect 21705 9192 21706 9256
rect 21640 9176 21706 9192
rect 21640 9112 21641 9176
rect 21705 9112 21706 9176
rect 21640 8958 21706 9112
rect 21766 9020 21826 10050
rect 21886 8958 21946 9990
rect 22006 9020 22066 10050
rect 22126 8958 22186 9990
rect 22246 9896 22312 9986
rect 22246 9832 22247 9896
rect 22311 9832 22312 9896
rect 22246 9816 22312 9832
rect 22246 9752 22247 9816
rect 22311 9752 22312 9816
rect 22246 9736 22312 9752
rect 22246 9672 22247 9736
rect 22311 9672 22312 9736
rect 22246 9656 22312 9672
rect 22246 9592 22247 9656
rect 22311 9592 22312 9656
rect 22246 9576 22312 9592
rect 22246 9512 22247 9576
rect 22311 9512 22312 9576
rect 22246 9496 22312 9512
rect 22246 9432 22247 9496
rect 22311 9432 22312 9496
rect 22246 9416 22312 9432
rect 22246 9352 22247 9416
rect 22311 9352 22312 9416
rect 22246 9336 22312 9352
rect 22246 9272 22247 9336
rect 22311 9272 22312 9336
rect 22246 9256 22312 9272
rect 22246 9192 22247 9256
rect 22311 9192 22312 9256
rect 22246 9176 22312 9192
rect 22246 9112 22247 9176
rect 22311 9112 22312 9176
rect 22246 8958 22312 9112
rect 21034 8956 22312 8958
rect 21034 8892 21138 8956
rect 21202 8892 21218 8956
rect 21282 8892 21298 8956
rect 21362 8892 21378 8956
rect 21442 8892 21458 8956
rect 21522 8933 21538 8956
rect 21522 8892 21532 8933
rect 21602 8892 21744 8956
rect 21808 8933 21824 8956
rect 21814 8892 21824 8933
rect 21888 8892 21904 8956
rect 21968 8892 21984 8956
rect 22048 8892 22064 8956
rect 22128 8892 22144 8956
rect 22208 8892 22312 8956
rect 21034 8890 21532 8892
rect 20862 8869 20871 8890
rect 20789 8863 20871 8869
rect 21523 8869 21532 8890
rect 21596 8890 21750 8892
rect 21596 8869 21605 8890
rect 21523 8863 21605 8869
rect 21741 8869 21750 8890
rect 21814 8890 22312 8892
rect 22372 9896 22438 9986
rect 22372 9832 22373 9896
rect 22437 9832 22438 9896
rect 22372 9816 22438 9832
rect 22372 9752 22373 9816
rect 22437 9752 22438 9816
rect 22372 9736 22438 9752
rect 22372 9672 22373 9736
rect 22437 9672 22438 9736
rect 22372 9656 22438 9672
rect 22372 9592 22373 9656
rect 22437 9592 22438 9656
rect 22372 9576 22438 9592
rect 22372 9512 22373 9576
rect 22437 9512 22438 9576
rect 22372 9496 22438 9512
rect 22372 9432 22373 9496
rect 22437 9432 22438 9496
rect 22372 9416 22438 9432
rect 22372 9352 22373 9416
rect 22437 9352 22438 9416
rect 22372 9336 22438 9352
rect 22372 9272 22373 9336
rect 22437 9272 22438 9336
rect 22372 9256 22438 9272
rect 22372 9192 22373 9256
rect 22437 9192 22438 9256
rect 22372 9176 22438 9192
rect 22372 9112 22373 9176
rect 22437 9112 22438 9176
rect 22372 8958 22438 9112
rect 22498 8958 22558 9990
rect 22618 9020 22678 10050
rect 22738 8958 22798 9990
rect 22858 9020 22918 10050
rect 22978 9896 23044 9986
rect 22978 9832 22979 9896
rect 23043 9832 23044 9896
rect 22978 9816 23044 9832
rect 22978 9752 22979 9816
rect 23043 9752 23044 9816
rect 22978 9736 23044 9752
rect 22978 9672 22979 9736
rect 23043 9672 23044 9736
rect 22978 9656 23044 9672
rect 22978 9592 22979 9656
rect 23043 9592 23044 9656
rect 22978 9576 23044 9592
rect 22978 9512 22979 9576
rect 23043 9512 23044 9576
rect 22978 9496 23044 9512
rect 22978 9432 22979 9496
rect 23043 9432 23044 9496
rect 22978 9416 23044 9432
rect 22978 9352 22979 9416
rect 23043 9352 23044 9416
rect 22978 9336 23044 9352
rect 22978 9272 22979 9336
rect 23043 9272 23044 9336
rect 22978 9256 23044 9272
rect 22978 9192 22979 9256
rect 23043 9192 23044 9256
rect 22978 9176 23044 9192
rect 22978 9112 22979 9176
rect 23043 9112 23044 9176
rect 22978 8958 23044 9112
rect 23104 9020 23164 10050
rect 23224 8958 23284 9990
rect 23344 9020 23404 10050
rect 23464 8958 23524 9990
rect 23584 9896 23650 9986
rect 23584 9832 23585 9896
rect 23649 9832 23650 9896
rect 23584 9816 23650 9832
rect 23584 9752 23585 9816
rect 23649 9752 23650 9816
rect 23584 9736 23650 9752
rect 23584 9672 23585 9736
rect 23649 9672 23650 9736
rect 23584 9656 23650 9672
rect 23584 9592 23585 9656
rect 23649 9592 23650 9656
rect 23584 9576 23650 9592
rect 23584 9512 23585 9576
rect 23649 9512 23650 9576
rect 23584 9496 23650 9512
rect 23584 9432 23585 9496
rect 23649 9432 23650 9496
rect 23584 9416 23650 9432
rect 23584 9352 23585 9416
rect 23649 9352 23650 9416
rect 23584 9336 23650 9352
rect 23584 9272 23585 9336
rect 23649 9272 23650 9336
rect 23584 9256 23650 9272
rect 23584 9192 23585 9256
rect 23649 9192 23650 9256
rect 23584 9176 23650 9192
rect 23584 9112 23585 9176
rect 23649 9112 23650 9176
rect 23584 8958 23650 9112
rect 23710 8958 23770 9990
rect 23830 9020 23890 10050
rect 23950 8958 24010 9990
rect 24070 9020 24130 10050
rect 24190 9896 24256 9986
rect 24190 9832 24191 9896
rect 24255 9832 24256 9896
rect 24190 9816 24256 9832
rect 24190 9752 24191 9816
rect 24255 9752 24256 9816
rect 24190 9736 24256 9752
rect 24190 9672 24191 9736
rect 24255 9672 24256 9736
rect 24190 9656 24256 9672
rect 24190 9592 24191 9656
rect 24255 9592 24256 9656
rect 24190 9576 24256 9592
rect 24190 9512 24191 9576
rect 24255 9512 24256 9576
rect 24190 9496 24256 9512
rect 24190 9432 24191 9496
rect 24255 9432 24256 9496
rect 24190 9416 24256 9432
rect 24190 9352 24191 9416
rect 24255 9352 24256 9416
rect 24190 9336 24256 9352
rect 24190 9272 24191 9336
rect 24255 9272 24256 9336
rect 24190 9256 24256 9272
rect 24190 9192 24191 9256
rect 24255 9192 24256 9256
rect 24190 9176 24256 9192
rect 24190 9112 24191 9176
rect 24255 9112 24256 9176
rect 24190 8958 24256 9112
rect 24316 9020 24376 10050
rect 24436 8958 24496 9990
rect 24556 9020 24616 10050
rect 24676 8958 24736 9990
rect 24796 9896 24862 9986
rect 24796 9832 24797 9896
rect 24861 9832 24862 9896
rect 24796 9816 24862 9832
rect 24796 9752 24797 9816
rect 24861 9752 24862 9816
rect 24796 9736 24862 9752
rect 24796 9672 24797 9736
rect 24861 9672 24862 9736
rect 24796 9656 24862 9672
rect 24796 9592 24797 9656
rect 24861 9592 24862 9656
rect 24796 9576 24862 9592
rect 24796 9512 24797 9576
rect 24861 9512 24862 9576
rect 24796 9496 24862 9512
rect 24796 9432 24797 9496
rect 24861 9432 24862 9496
rect 24796 9416 24862 9432
rect 24796 9352 24797 9416
rect 24861 9352 24862 9416
rect 24796 9336 24862 9352
rect 24796 9272 24797 9336
rect 24861 9272 24862 9336
rect 24796 9256 24862 9272
rect 24796 9192 24797 9256
rect 24861 9192 24862 9256
rect 24796 9176 24862 9192
rect 24796 9112 24797 9176
rect 24861 9112 24862 9176
rect 24796 8958 24862 9112
rect 22372 8956 24862 8958
rect 22372 8892 22476 8956
rect 22540 8892 22556 8956
rect 22620 8892 22636 8956
rect 22700 8892 22716 8956
rect 22780 8892 22796 8956
rect 22860 8933 22876 8956
rect 22860 8892 22870 8933
rect 22940 8892 23082 8956
rect 23146 8933 23162 8956
rect 23152 8892 23162 8933
rect 23226 8892 23242 8956
rect 23306 8892 23322 8956
rect 23386 8892 23402 8956
rect 23466 8892 23482 8956
rect 23546 8892 23688 8956
rect 23752 8892 23768 8956
rect 23832 8892 23848 8956
rect 23912 8892 23928 8956
rect 23992 8892 24008 8956
rect 24072 8933 24088 8956
rect 24072 8892 24082 8933
rect 24152 8892 24294 8956
rect 24358 8933 24374 8956
rect 24364 8892 24374 8933
rect 24438 8892 24454 8956
rect 24518 8892 24534 8956
rect 24598 8892 24614 8956
rect 24678 8892 24694 8956
rect 24758 8892 24862 8956
rect 22372 8890 22870 8892
rect 21814 8869 21823 8890
rect 21741 8863 21823 8869
rect 22861 8869 22870 8890
rect 22934 8890 23088 8892
rect 22934 8869 22943 8890
rect 22861 8863 22943 8869
rect 23079 8869 23088 8890
rect 23152 8890 24082 8892
rect 23152 8869 23161 8890
rect 23079 8863 23161 8869
rect 24073 8869 24082 8890
rect 24146 8890 24300 8892
rect 24146 8869 24155 8890
rect 24073 8863 24155 8869
rect 24291 8869 24300 8890
rect 24364 8890 24862 8892
rect 24922 9896 24988 9986
rect 24922 9832 24923 9896
rect 24987 9832 24988 9896
rect 24922 9816 24988 9832
rect 24922 9752 24923 9816
rect 24987 9752 24988 9816
rect 24922 9736 24988 9752
rect 24922 9672 24923 9736
rect 24987 9672 24988 9736
rect 24922 9656 24988 9672
rect 24922 9592 24923 9656
rect 24987 9592 24988 9656
rect 24922 9576 24988 9592
rect 24922 9512 24923 9576
rect 24987 9512 24988 9576
rect 24922 9496 24988 9512
rect 24922 9432 24923 9496
rect 24987 9432 24988 9496
rect 24922 9416 24988 9432
rect 24922 9352 24923 9416
rect 24987 9352 24988 9416
rect 24922 9336 24988 9352
rect 24922 9272 24923 9336
rect 24987 9272 24988 9336
rect 24922 9256 24988 9272
rect 24922 9192 24923 9256
rect 24987 9192 24988 9256
rect 24922 9176 24988 9192
rect 24922 9112 24923 9176
rect 24987 9112 24988 9176
rect 24922 8958 24988 9112
rect 25048 9020 25108 10050
rect 25168 8958 25228 9990
rect 25288 9020 25348 10050
rect 25857 10045 25982 10055
rect 25408 8958 25468 9990
rect 25528 9896 25594 9986
rect 25528 9832 25529 9896
rect 25593 9832 25594 9896
rect 25528 9816 25594 9832
rect 25528 9752 25529 9816
rect 25593 9752 25594 9816
rect 25528 9736 25594 9752
rect 25528 9672 25529 9736
rect 25593 9672 25594 9736
rect 25528 9656 25594 9672
rect 25528 9592 25529 9656
rect 25593 9592 25594 9656
rect 25528 9576 25594 9592
rect 25528 9512 25529 9576
rect 25593 9512 25594 9576
rect 25528 9496 25594 9512
rect 25528 9432 25529 9496
rect 25593 9432 25594 9496
rect 25528 9416 25594 9432
rect 25528 9352 25529 9416
rect 25593 9352 25594 9416
rect 25528 9336 25594 9352
rect 25528 9272 25529 9336
rect 25593 9272 25594 9336
rect 25528 9256 25594 9272
rect 25528 9192 25529 9256
rect 25593 9192 25594 9256
rect 25528 9176 25594 9192
rect 25528 9112 25529 9176
rect 25593 9112 25594 9176
rect 25528 8958 25594 9112
rect 24922 8956 25594 8958
rect 24922 8892 25026 8956
rect 25090 8933 25106 8956
rect 25096 8892 25106 8933
rect 25170 8892 25186 8956
rect 25250 8892 25266 8956
rect 25330 8892 25346 8956
rect 25410 8892 25426 8956
rect 25490 8892 25594 8956
rect 24922 8890 25032 8892
rect 24364 8869 24373 8890
rect 24291 8863 24373 8869
rect 25023 8869 25032 8890
rect 25096 8890 25594 8892
rect 25096 8869 25105 8890
rect 25023 8863 25105 8869
rect 3538 8746 3621 8751
rect 3538 8725 3548 8746
rect 3055 8723 3548 8725
rect 3612 8725 3621 8746
rect 4270 8743 4353 8748
rect 3612 8723 3727 8725
rect 2456 8704 2829 8721
rect 2456 8640 2463 8704
rect 2527 8640 2583 8704
rect 2647 8640 2726 8704
rect 2790 8640 2829 8704
rect 2456 8625 2829 8640
rect 3055 8659 3159 8723
rect 3223 8659 3239 8723
rect 3303 8659 3319 8723
rect 3383 8659 3399 8723
rect 3463 8659 3479 8723
rect 3543 8682 3548 8723
rect 3543 8659 3559 8682
rect 3623 8659 3727 8723
rect 4270 8722 4280 8743
rect 3055 8657 3727 8659
rect 2570 8624 2662 8625
rect 3055 8503 3121 8657
rect 3055 8439 3056 8503
rect 3120 8439 3121 8503
rect 3055 8423 3121 8439
rect 3055 8359 3056 8423
rect 3120 8359 3121 8423
rect 3055 8343 3121 8359
rect 3055 8279 3056 8343
rect 3120 8279 3121 8343
rect 3055 8263 3121 8279
rect 3055 8199 3056 8263
rect 3120 8199 3121 8263
rect 3055 8183 3121 8199
rect 2535 8175 2679 8176
rect 2430 8159 2823 8175
rect 2430 8158 2576 8159
rect 2430 8094 2445 8158
rect 2509 8095 2576 8158
rect 2640 8158 2823 8159
rect 2640 8095 2720 8158
rect 2509 8094 2720 8095
rect 2784 8094 2823 8158
rect 2430 8080 2823 8094
rect 2430 8079 2548 8080
rect 2679 8079 2823 8080
rect 3055 8119 3056 8183
rect 3120 8119 3121 8183
rect 3055 8103 3121 8119
rect 3055 8039 3056 8103
rect 3120 8039 3121 8103
rect 3055 8023 3121 8039
rect 3055 7959 3056 8023
rect 3120 7959 3121 8023
rect 3055 7943 3121 7959
rect 3055 7879 3056 7943
rect 3120 7879 3121 7943
rect 3055 7863 3121 7879
rect 3055 7799 3056 7863
rect 3120 7799 3121 7863
rect 3055 7783 3121 7799
rect 3055 7719 3056 7783
rect 3120 7719 3121 7783
rect 3055 7629 3121 7719
rect 3181 7625 3241 8657
rect 3301 7565 3361 8595
rect 3421 7625 3481 8657
rect 3541 7565 3601 8595
rect 3661 8503 3727 8657
rect 3661 8439 3662 8503
rect 3726 8439 3727 8503
rect 3661 8423 3727 8439
rect 3661 8359 3662 8423
rect 3726 8359 3727 8423
rect 3661 8343 3727 8359
rect 3661 8279 3662 8343
rect 3726 8279 3727 8343
rect 3661 8263 3727 8279
rect 3661 8199 3662 8263
rect 3726 8199 3727 8263
rect 3661 8183 3727 8199
rect 3661 8119 3662 8183
rect 3726 8119 3727 8183
rect 3661 8103 3727 8119
rect 3661 8039 3662 8103
rect 3726 8039 3727 8103
rect 3661 8023 3727 8039
rect 3661 7959 3662 8023
rect 3726 7959 3727 8023
rect 3661 7943 3727 7959
rect 3661 7879 3662 7943
rect 3726 7879 3727 7943
rect 3661 7863 3727 7879
rect 3661 7799 3662 7863
rect 3726 7799 3727 7863
rect 3661 7783 3727 7799
rect 3661 7719 3662 7783
rect 3726 7719 3727 7783
rect 3661 7629 3727 7719
rect 3787 8720 4280 8722
rect 4344 8722 4353 8743
rect 4499 8743 4582 8748
rect 4499 8722 4508 8743
rect 4344 8720 4508 8722
rect 4572 8722 4582 8743
rect 5482 8743 5565 8748
rect 5482 8722 5492 8743
rect 4572 8720 5492 8722
rect 5556 8722 5565 8743
rect 5711 8743 5794 8748
rect 5711 8722 5720 8743
rect 5556 8720 5720 8722
rect 5784 8722 5794 8743
rect 6694 8743 6777 8748
rect 6694 8722 6704 8743
rect 5784 8720 6704 8722
rect 6768 8722 6777 8743
rect 6923 8743 7006 8748
rect 6923 8722 6932 8743
rect 6768 8720 6932 8722
rect 6996 8722 7006 8743
rect 7906 8743 7989 8748
rect 7906 8722 7916 8743
rect 6996 8720 7916 8722
rect 7980 8722 7989 8743
rect 8135 8743 8218 8748
rect 8135 8722 8144 8743
rect 7980 8720 8144 8722
rect 8208 8722 8218 8743
rect 8851 8741 8977 8751
rect 8208 8720 8701 8722
rect 3787 8656 3891 8720
rect 3955 8656 3971 8720
rect 4035 8656 4051 8720
rect 4115 8656 4131 8720
rect 4195 8656 4211 8720
rect 4275 8679 4280 8720
rect 4275 8656 4291 8679
rect 4355 8656 4497 8720
rect 4572 8679 4577 8720
rect 4561 8656 4577 8679
rect 4641 8656 4657 8720
rect 4721 8656 4737 8720
rect 4801 8656 4817 8720
rect 4881 8656 4897 8720
rect 4961 8656 5103 8720
rect 5167 8656 5183 8720
rect 5247 8656 5263 8720
rect 5327 8656 5343 8720
rect 5407 8656 5423 8720
rect 5487 8679 5492 8720
rect 5487 8656 5503 8679
rect 5567 8656 5709 8720
rect 5784 8679 5789 8720
rect 5773 8656 5789 8679
rect 5853 8656 5869 8720
rect 5933 8656 5949 8720
rect 6013 8656 6029 8720
rect 6093 8656 6109 8720
rect 6173 8656 6315 8720
rect 6379 8656 6395 8720
rect 6459 8656 6475 8720
rect 6539 8656 6555 8720
rect 6619 8656 6635 8720
rect 6699 8679 6704 8720
rect 6699 8656 6715 8679
rect 6779 8656 6921 8720
rect 6996 8679 7001 8720
rect 6985 8656 7001 8679
rect 7065 8656 7081 8720
rect 7145 8656 7161 8720
rect 7225 8656 7241 8720
rect 7305 8656 7321 8720
rect 7385 8656 7527 8720
rect 7591 8656 7607 8720
rect 7671 8656 7687 8720
rect 7751 8656 7767 8720
rect 7831 8656 7847 8720
rect 7911 8679 7916 8720
rect 7911 8656 7927 8679
rect 7991 8656 8133 8720
rect 8208 8679 8213 8720
rect 8197 8656 8213 8679
rect 8277 8656 8293 8720
rect 8357 8656 8373 8720
rect 8437 8656 8453 8720
rect 8517 8656 8533 8720
rect 8597 8656 8701 8720
rect 8851 8677 8882 8741
rect 8946 8677 8977 8741
rect 8851 8667 8977 8677
rect 13314 8729 13440 8739
rect 3787 8654 8701 8656
rect 13314 8665 13345 8729
rect 13409 8665 13440 8729
rect 14073 8731 14156 8736
rect 14073 8710 14083 8731
rect 13314 8655 13440 8665
rect 13590 8708 14083 8710
rect 14147 8710 14156 8731
rect 14302 8731 14385 8736
rect 14302 8710 14311 8731
rect 14147 8708 14311 8710
rect 14375 8710 14385 8731
rect 15285 8731 15368 8736
rect 15285 8710 15295 8731
rect 14375 8708 15295 8710
rect 15359 8710 15368 8731
rect 15514 8731 15597 8736
rect 15514 8710 15523 8731
rect 15359 8708 15523 8710
rect 15587 8710 15597 8731
rect 16497 8731 16580 8736
rect 16497 8710 16507 8731
rect 15587 8708 16507 8710
rect 16571 8710 16580 8731
rect 16726 8731 16809 8736
rect 16726 8710 16735 8731
rect 16571 8708 16735 8710
rect 16799 8710 16809 8731
rect 17709 8731 17792 8736
rect 17709 8710 17719 8731
rect 16799 8708 17719 8710
rect 17783 8710 17792 8731
rect 17938 8731 18021 8736
rect 17938 8710 17947 8731
rect 17783 8708 17947 8710
rect 18011 8710 18021 8731
rect 18670 8734 18753 8739
rect 18670 8713 18679 8734
rect 18564 8711 18679 8713
rect 18743 8713 18753 8734
rect 20023 8729 20149 8739
rect 18743 8711 19236 8713
rect 18011 8708 18504 8710
rect 3787 8500 3853 8654
rect 3787 8436 3788 8500
rect 3852 8436 3853 8500
rect 3787 8420 3853 8436
rect 3787 8356 3788 8420
rect 3852 8356 3853 8420
rect 3787 8340 3853 8356
rect 3787 8276 3788 8340
rect 3852 8276 3853 8340
rect 3787 8260 3853 8276
rect 3787 8196 3788 8260
rect 3852 8196 3853 8260
rect 3787 8180 3853 8196
rect 3787 8116 3788 8180
rect 3852 8116 3853 8180
rect 3787 8100 3853 8116
rect 3787 8036 3788 8100
rect 3852 8036 3853 8100
rect 3787 8020 3853 8036
rect 3787 7956 3788 8020
rect 3852 7956 3853 8020
rect 3787 7940 3853 7956
rect 3787 7876 3788 7940
rect 3852 7876 3853 7940
rect 3787 7860 3853 7876
rect 3787 7796 3788 7860
rect 3852 7796 3853 7860
rect 3787 7780 3853 7796
rect 3787 7716 3788 7780
rect 3852 7716 3853 7780
rect 3787 7626 3853 7716
rect 3913 7622 3973 8654
rect 3055 7563 3727 7565
rect 3055 7562 3159 7563
rect 3031 7553 3159 7562
rect 3031 7489 3062 7553
rect 3126 7499 3159 7553
rect 3223 7499 3239 7563
rect 3303 7499 3319 7563
rect 3383 7499 3399 7563
rect 3463 7499 3479 7563
rect 3543 7499 3559 7563
rect 3623 7499 3727 7563
rect 4033 7562 4093 8592
rect 4153 7622 4213 8654
rect 4273 7562 4333 8592
rect 4393 8500 4459 8654
rect 4393 8436 4394 8500
rect 4458 8436 4459 8500
rect 4393 8420 4459 8436
rect 4393 8356 4394 8420
rect 4458 8356 4459 8420
rect 4393 8340 4459 8356
rect 4393 8276 4394 8340
rect 4458 8276 4459 8340
rect 4393 8260 4459 8276
rect 4393 8196 4394 8260
rect 4458 8196 4459 8260
rect 4393 8180 4459 8196
rect 4393 8116 4394 8180
rect 4458 8116 4459 8180
rect 4393 8100 4459 8116
rect 4393 8036 4394 8100
rect 4458 8036 4459 8100
rect 4393 8020 4459 8036
rect 4393 7956 4394 8020
rect 4458 7956 4459 8020
rect 4393 7940 4459 7956
rect 4393 7876 4394 7940
rect 4458 7876 4459 7940
rect 4393 7860 4459 7876
rect 4393 7796 4394 7860
rect 4458 7796 4459 7860
rect 4393 7780 4459 7796
rect 4393 7716 4394 7780
rect 4458 7716 4459 7780
rect 4393 7626 4459 7716
rect 4519 7562 4579 8592
rect 4639 7622 4699 8654
rect 4759 7562 4819 8592
rect 4879 7622 4939 8654
rect 4999 8500 5065 8654
rect 4999 8436 5000 8500
rect 5064 8436 5065 8500
rect 4999 8420 5065 8436
rect 4999 8356 5000 8420
rect 5064 8356 5065 8420
rect 4999 8340 5065 8356
rect 4999 8276 5000 8340
rect 5064 8276 5065 8340
rect 4999 8260 5065 8276
rect 4999 8196 5000 8260
rect 5064 8196 5065 8260
rect 4999 8180 5065 8196
rect 4999 8116 5000 8180
rect 5064 8116 5065 8180
rect 4999 8100 5065 8116
rect 4999 8036 5000 8100
rect 5064 8036 5065 8100
rect 4999 8020 5065 8036
rect 4999 7956 5000 8020
rect 5064 7956 5065 8020
rect 4999 7940 5065 7956
rect 4999 7876 5000 7940
rect 5064 7876 5065 7940
rect 4999 7860 5065 7876
rect 4999 7796 5000 7860
rect 5064 7796 5065 7860
rect 4999 7780 5065 7796
rect 4999 7716 5000 7780
rect 5064 7716 5065 7780
rect 4999 7626 5065 7716
rect 5125 7622 5185 8654
rect 5245 7562 5305 8592
rect 5365 7622 5425 8654
rect 5485 7562 5545 8592
rect 5605 8500 5671 8654
rect 5605 8436 5606 8500
rect 5670 8436 5671 8500
rect 5605 8420 5671 8436
rect 5605 8356 5606 8420
rect 5670 8356 5671 8420
rect 5605 8340 5671 8356
rect 5605 8276 5606 8340
rect 5670 8276 5671 8340
rect 5605 8260 5671 8276
rect 5605 8196 5606 8260
rect 5670 8196 5671 8260
rect 5605 8180 5671 8196
rect 5605 8116 5606 8180
rect 5670 8116 5671 8180
rect 5605 8100 5671 8116
rect 5605 8036 5606 8100
rect 5670 8036 5671 8100
rect 5605 8020 5671 8036
rect 5605 7956 5606 8020
rect 5670 7956 5671 8020
rect 5605 7940 5671 7956
rect 5605 7876 5606 7940
rect 5670 7876 5671 7940
rect 5605 7860 5671 7876
rect 5605 7796 5606 7860
rect 5670 7796 5671 7860
rect 5605 7780 5671 7796
rect 5605 7716 5606 7780
rect 5670 7716 5671 7780
rect 5605 7626 5671 7716
rect 5731 7562 5791 8592
rect 5851 7622 5911 8654
rect 5971 7562 6031 8592
rect 6091 7622 6151 8654
rect 6211 8500 6277 8654
rect 6211 8436 6212 8500
rect 6276 8436 6277 8500
rect 6211 8420 6277 8436
rect 6211 8356 6212 8420
rect 6276 8356 6277 8420
rect 6211 8340 6277 8356
rect 6211 8276 6212 8340
rect 6276 8276 6277 8340
rect 6211 8260 6277 8276
rect 6211 8196 6212 8260
rect 6276 8196 6277 8260
rect 6211 8180 6277 8196
rect 6211 8116 6212 8180
rect 6276 8116 6277 8180
rect 6211 8100 6277 8116
rect 6211 8036 6212 8100
rect 6276 8036 6277 8100
rect 6211 8020 6277 8036
rect 6211 7956 6212 8020
rect 6276 7956 6277 8020
rect 6211 7940 6277 7956
rect 6211 7876 6212 7940
rect 6276 7876 6277 7940
rect 6211 7860 6277 7876
rect 6211 7796 6212 7860
rect 6276 7796 6277 7860
rect 6211 7780 6277 7796
rect 6211 7716 6212 7780
rect 6276 7716 6277 7780
rect 6211 7626 6277 7716
rect 6337 7622 6397 8654
rect 6457 7562 6517 8592
rect 6577 7622 6637 8654
rect 6697 7562 6757 8592
rect 6817 8500 6883 8654
rect 6817 8436 6818 8500
rect 6882 8436 6883 8500
rect 6817 8420 6883 8436
rect 6817 8356 6818 8420
rect 6882 8356 6883 8420
rect 6817 8340 6883 8356
rect 6817 8276 6818 8340
rect 6882 8276 6883 8340
rect 6817 8260 6883 8276
rect 6817 8196 6818 8260
rect 6882 8196 6883 8260
rect 6817 8180 6883 8196
rect 6817 8116 6818 8180
rect 6882 8116 6883 8180
rect 6817 8100 6883 8116
rect 6817 8036 6818 8100
rect 6882 8036 6883 8100
rect 6817 8020 6883 8036
rect 6817 7956 6818 8020
rect 6882 7956 6883 8020
rect 6817 7940 6883 7956
rect 6817 7876 6818 7940
rect 6882 7876 6883 7940
rect 6817 7860 6883 7876
rect 6817 7796 6818 7860
rect 6882 7796 6883 7860
rect 6817 7780 6883 7796
rect 6817 7716 6818 7780
rect 6882 7716 6883 7780
rect 6817 7626 6883 7716
rect 6943 7562 7003 8592
rect 7063 7622 7123 8654
rect 7183 7562 7243 8592
rect 7303 7622 7363 8654
rect 7423 8500 7489 8654
rect 7423 8436 7424 8500
rect 7488 8436 7489 8500
rect 7423 8420 7489 8436
rect 7423 8356 7424 8420
rect 7488 8356 7489 8420
rect 7423 8340 7489 8356
rect 7423 8276 7424 8340
rect 7488 8276 7489 8340
rect 7423 8260 7489 8276
rect 7423 8196 7424 8260
rect 7488 8196 7489 8260
rect 7423 8180 7489 8196
rect 7423 8116 7424 8180
rect 7488 8116 7489 8180
rect 7423 8100 7489 8116
rect 7423 8036 7424 8100
rect 7488 8036 7489 8100
rect 7423 8020 7489 8036
rect 7423 7956 7424 8020
rect 7488 7956 7489 8020
rect 7423 7940 7489 7956
rect 7423 7876 7424 7940
rect 7488 7876 7489 7940
rect 7423 7860 7489 7876
rect 7423 7796 7424 7860
rect 7488 7796 7489 7860
rect 7423 7780 7489 7796
rect 7423 7716 7424 7780
rect 7488 7716 7489 7780
rect 7423 7626 7489 7716
rect 7549 7622 7609 8654
rect 7669 7562 7729 8592
rect 7789 7622 7849 8654
rect 7909 7562 7969 8592
rect 8029 8500 8095 8654
rect 8029 8436 8030 8500
rect 8094 8436 8095 8500
rect 8029 8420 8095 8436
rect 8029 8356 8030 8420
rect 8094 8356 8095 8420
rect 8029 8340 8095 8356
rect 8029 8276 8030 8340
rect 8094 8276 8095 8340
rect 8029 8260 8095 8276
rect 8029 8196 8030 8260
rect 8094 8196 8095 8260
rect 8029 8180 8095 8196
rect 8029 8116 8030 8180
rect 8094 8116 8095 8180
rect 8029 8100 8095 8116
rect 8029 8036 8030 8100
rect 8094 8036 8095 8100
rect 8029 8020 8095 8036
rect 8029 7956 8030 8020
rect 8094 7956 8095 8020
rect 8029 7940 8095 7956
rect 8029 7876 8030 7940
rect 8094 7876 8095 7940
rect 8029 7860 8095 7876
rect 8029 7796 8030 7860
rect 8094 7796 8095 7860
rect 8029 7780 8095 7796
rect 8029 7716 8030 7780
rect 8094 7716 8095 7780
rect 8029 7626 8095 7716
rect 8155 7562 8215 8592
rect 8275 7622 8335 8654
rect 8395 7562 8455 8592
rect 8515 7622 8575 8654
rect 8635 8500 8701 8654
rect 13590 8644 13694 8708
rect 13758 8644 13774 8708
rect 13838 8644 13854 8708
rect 13918 8644 13934 8708
rect 13998 8644 14014 8708
rect 14078 8667 14083 8708
rect 14078 8644 14094 8667
rect 14158 8644 14300 8708
rect 14375 8667 14380 8708
rect 14364 8644 14380 8667
rect 14444 8644 14460 8708
rect 14524 8644 14540 8708
rect 14604 8644 14620 8708
rect 14684 8644 14700 8708
rect 14764 8644 14906 8708
rect 14970 8644 14986 8708
rect 15050 8644 15066 8708
rect 15130 8644 15146 8708
rect 15210 8644 15226 8708
rect 15290 8667 15295 8708
rect 15290 8644 15306 8667
rect 15370 8644 15512 8708
rect 15587 8667 15592 8708
rect 15576 8644 15592 8667
rect 15656 8644 15672 8708
rect 15736 8644 15752 8708
rect 15816 8644 15832 8708
rect 15896 8644 15912 8708
rect 15976 8644 16118 8708
rect 16182 8644 16198 8708
rect 16262 8644 16278 8708
rect 16342 8644 16358 8708
rect 16422 8644 16438 8708
rect 16502 8667 16507 8708
rect 16502 8644 16518 8667
rect 16582 8644 16724 8708
rect 16799 8667 16804 8708
rect 16788 8644 16804 8667
rect 16868 8644 16884 8708
rect 16948 8644 16964 8708
rect 17028 8644 17044 8708
rect 17108 8644 17124 8708
rect 17188 8644 17330 8708
rect 17394 8644 17410 8708
rect 17474 8644 17490 8708
rect 17554 8644 17570 8708
rect 17634 8644 17650 8708
rect 17714 8667 17719 8708
rect 17714 8644 17730 8667
rect 17794 8644 17936 8708
rect 18011 8667 18016 8708
rect 18000 8644 18016 8667
rect 18080 8644 18096 8708
rect 18160 8644 18176 8708
rect 18240 8644 18256 8708
rect 18320 8644 18336 8708
rect 18400 8644 18504 8708
rect 13590 8642 18504 8644
rect 8635 8436 8636 8500
rect 8700 8436 8701 8500
rect 12692 8512 12813 8521
rect 8635 8420 8701 8436
rect 8635 8356 8636 8420
rect 8700 8356 8701 8420
rect 8763 8480 8889 8490
rect 8763 8416 8794 8480
rect 8858 8416 8889 8480
rect 8763 8406 8889 8416
rect 9171 8454 9297 8464
rect 9171 8390 9204 8454
rect 9268 8390 9297 8454
rect 9171 8381 9297 8390
rect 9433 8455 9559 8465
rect 9433 8391 9466 8455
rect 9530 8391 9559 8455
rect 9433 8383 9559 8391
rect 9705 8455 9831 8465
rect 9705 8391 9738 8455
rect 9802 8391 9831 8455
rect 9705 8383 9831 8391
rect 10032 8455 10158 8465
rect 10032 8391 10065 8455
rect 10129 8391 10158 8455
rect 10032 8383 10158 8391
rect 10413 8455 10539 8465
rect 10413 8391 10446 8455
rect 10510 8391 10539 8455
rect 10413 8383 10539 8391
rect 10790 8455 10916 8463
rect 10790 8391 10823 8455
rect 10887 8391 10916 8455
rect 10790 8383 10916 8391
rect 12197 8442 12318 8451
rect 9190 8380 9280 8381
rect 12197 8378 12224 8442
rect 12288 8378 12318 8442
rect 12692 8448 12719 8512
rect 12783 8448 12813 8512
rect 12692 8439 12813 8448
rect 13066 8512 13187 8521
rect 13066 8448 13093 8512
rect 13157 8448 13187 8512
rect 13590 8488 13656 8642
rect 13066 8439 13187 8448
rect 13402 8468 13528 8478
rect 13402 8404 13433 8468
rect 13497 8404 13528 8468
rect 13402 8394 13528 8404
rect 13590 8424 13591 8488
rect 13655 8424 13656 8488
rect 13590 8408 13656 8424
rect 12197 8369 12318 8378
rect 12554 8369 12675 8378
rect 8635 8340 8701 8356
rect 8635 8276 8636 8340
rect 8700 8276 8701 8340
rect 12554 8305 12581 8369
rect 12645 8305 12675 8369
rect 12554 8296 12675 8305
rect 12738 8366 12859 8375
rect 12738 8302 12765 8366
rect 12829 8302 12859 8366
rect 12738 8293 12859 8302
rect 13040 8360 13161 8369
rect 13040 8296 13067 8360
rect 13131 8296 13161 8360
rect 13040 8287 13161 8296
rect 13590 8344 13591 8408
rect 13655 8344 13656 8408
rect 13590 8328 13656 8344
rect 8635 8260 8701 8276
rect 8635 8196 8636 8260
rect 8700 8196 8701 8260
rect 13590 8264 13591 8328
rect 13655 8264 13656 8328
rect 13590 8248 13656 8264
rect 8635 8180 8701 8196
rect 8635 8116 8636 8180
rect 8700 8116 8701 8180
rect 8845 8238 8971 8248
rect 8845 8174 8876 8238
rect 8940 8174 8971 8238
rect 8845 8164 8971 8174
rect 13320 8226 13446 8236
rect 13320 8162 13351 8226
rect 13415 8162 13446 8226
rect 13320 8152 13446 8162
rect 13590 8184 13591 8248
rect 13655 8184 13656 8248
rect 13590 8168 13656 8184
rect 8635 8100 8701 8116
rect 8635 8036 8636 8100
rect 8700 8036 8701 8100
rect 13590 8104 13591 8168
rect 13655 8104 13656 8168
rect 8635 8020 8701 8036
rect 8635 7956 8636 8020
rect 8700 7956 8701 8020
rect 8846 8081 8972 8091
rect 8846 8017 8877 8081
rect 8941 8017 8972 8081
rect 13590 8088 13656 8104
rect 8846 8007 8972 8017
rect 13319 8069 13445 8079
rect 13319 8005 13350 8069
rect 13414 8005 13445 8069
rect 13319 7995 13445 8005
rect 13590 8024 13591 8088
rect 13655 8024 13656 8088
rect 13590 8008 13656 8024
rect 8635 7940 8701 7956
rect 8635 7876 8636 7940
rect 8700 7876 8701 7940
rect 12903 7935 13029 7945
rect 8635 7860 8701 7876
rect 8635 7796 8636 7860
rect 8700 7796 8701 7860
rect 8846 7911 8972 7921
rect 8846 7847 8877 7911
rect 8941 7847 8972 7911
rect 12903 7871 12934 7935
rect 12998 7871 13029 7935
rect 13590 7944 13591 8008
rect 13655 7944 13656 8008
rect 13590 7928 13656 7944
rect 12903 7861 13029 7871
rect 13319 7899 13445 7909
rect 8846 7837 8972 7847
rect 13319 7835 13350 7899
rect 13414 7835 13445 7899
rect 13319 7825 13445 7835
rect 13590 7864 13591 7928
rect 13655 7864 13656 7928
rect 13590 7848 13656 7864
rect 8635 7780 8701 7796
rect 8635 7716 8636 7780
rect 8700 7716 8701 7780
rect 13590 7784 13591 7848
rect 13655 7784 13656 7848
rect 8635 7626 8701 7716
rect 8845 7759 8971 7769
rect 8845 7695 8876 7759
rect 8940 7695 8971 7759
rect 13590 7768 13656 7784
rect 8845 7685 8971 7695
rect 10110 7729 10235 7739
rect 10110 7665 10140 7729
rect 10204 7665 10235 7729
rect 10110 7655 10235 7665
rect 10358 7729 10483 7739
rect 10358 7665 10388 7729
rect 10452 7665 10483 7729
rect 10358 7655 10483 7665
rect 10655 7729 10780 7739
rect 10655 7665 10685 7729
rect 10749 7665 10780 7729
rect 10655 7655 10780 7665
rect 10999 7731 11124 7741
rect 10999 7667 11029 7731
rect 11093 7667 11124 7731
rect 10999 7657 11124 7667
rect 11318 7731 11443 7741
rect 11318 7667 11348 7731
rect 11412 7667 11443 7731
rect 11318 7657 11443 7667
rect 11930 7740 12055 7750
rect 11930 7676 11960 7740
rect 12024 7676 12055 7740
rect 11930 7666 12055 7676
rect 12184 7744 12309 7754
rect 12184 7680 12214 7744
rect 12278 7680 12309 7744
rect 13320 7747 13446 7757
rect 12184 7670 12309 7680
rect 12895 7715 13021 7725
rect 12895 7651 12926 7715
rect 12990 7651 13021 7715
rect 13320 7683 13351 7747
rect 13415 7683 13446 7747
rect 13320 7673 13446 7683
rect 13590 7704 13591 7768
rect 13655 7704 13656 7768
rect 12895 7641 13021 7651
rect 8840 7615 8966 7625
rect 3126 7497 3727 7499
rect 3787 7560 8701 7562
rect 3126 7489 3157 7497
rect 3787 7496 3891 7560
rect 3955 7496 3971 7560
rect 4035 7496 4051 7560
rect 4115 7496 4131 7560
rect 4195 7496 4211 7560
rect 4275 7496 4291 7560
rect 4355 7496 4497 7560
rect 4561 7496 4577 7560
rect 4641 7496 4657 7560
rect 4721 7496 4737 7560
rect 4801 7496 4817 7560
rect 4881 7496 4897 7560
rect 4961 7496 5103 7560
rect 5167 7496 5183 7560
rect 5247 7496 5263 7560
rect 5327 7496 5343 7560
rect 5407 7496 5423 7560
rect 5487 7496 5503 7560
rect 5567 7496 5709 7560
rect 5773 7496 5789 7560
rect 5853 7496 5869 7560
rect 5933 7496 5949 7560
rect 6013 7496 6029 7560
rect 6093 7496 6109 7560
rect 6173 7496 6315 7560
rect 6379 7496 6395 7560
rect 6459 7496 6475 7560
rect 6539 7496 6555 7560
rect 6619 7496 6635 7560
rect 6699 7496 6715 7560
rect 6779 7496 6921 7560
rect 6985 7496 7001 7560
rect 7065 7496 7081 7560
rect 7145 7496 7161 7560
rect 7225 7496 7241 7560
rect 7305 7496 7321 7560
rect 7385 7496 7527 7560
rect 7591 7496 7607 7560
rect 7671 7496 7687 7560
rect 7751 7496 7767 7560
rect 7831 7496 7847 7560
rect 7911 7496 7927 7560
rect 7991 7496 8133 7560
rect 8197 7496 8213 7560
rect 8277 7496 8293 7560
rect 8357 7496 8373 7560
rect 8437 7496 8453 7560
rect 8517 7496 8533 7560
rect 8597 7496 8701 7560
rect 8840 7551 8871 7615
rect 8935 7551 8966 7615
rect 13590 7614 13656 7704
rect 8840 7541 8966 7551
rect 11940 7595 12065 7605
rect 11940 7531 11970 7595
rect 12034 7531 12065 7595
rect 11940 7521 12065 7531
rect 12192 7598 12317 7607
rect 12192 7534 12222 7598
rect 12286 7534 12317 7598
rect 12192 7524 12317 7534
rect 13325 7603 13451 7613
rect 13716 7610 13776 8642
rect 13325 7539 13356 7603
rect 13420 7539 13451 7603
rect 13836 7550 13896 8580
rect 13956 7610 14016 8642
rect 14076 7550 14136 8580
rect 14196 8488 14262 8642
rect 14196 8424 14197 8488
rect 14261 8424 14262 8488
rect 14196 8408 14262 8424
rect 14196 8344 14197 8408
rect 14261 8344 14262 8408
rect 14196 8328 14262 8344
rect 14196 8264 14197 8328
rect 14261 8264 14262 8328
rect 14196 8248 14262 8264
rect 14196 8184 14197 8248
rect 14261 8184 14262 8248
rect 14196 8168 14262 8184
rect 14196 8104 14197 8168
rect 14261 8104 14262 8168
rect 14196 8088 14262 8104
rect 14196 8024 14197 8088
rect 14261 8024 14262 8088
rect 14196 8008 14262 8024
rect 14196 7944 14197 8008
rect 14261 7944 14262 8008
rect 14196 7928 14262 7944
rect 14196 7864 14197 7928
rect 14261 7864 14262 7928
rect 14196 7848 14262 7864
rect 14196 7784 14197 7848
rect 14261 7784 14262 7848
rect 14196 7768 14262 7784
rect 14196 7704 14197 7768
rect 14261 7704 14262 7768
rect 14196 7614 14262 7704
rect 14322 7550 14382 8580
rect 14442 7610 14502 8642
rect 14562 7550 14622 8580
rect 14682 7610 14742 8642
rect 14802 8488 14868 8642
rect 14802 8424 14803 8488
rect 14867 8424 14868 8488
rect 14802 8408 14868 8424
rect 14802 8344 14803 8408
rect 14867 8344 14868 8408
rect 14802 8328 14868 8344
rect 14802 8264 14803 8328
rect 14867 8264 14868 8328
rect 14802 8248 14868 8264
rect 14802 8184 14803 8248
rect 14867 8184 14868 8248
rect 14802 8168 14868 8184
rect 14802 8104 14803 8168
rect 14867 8104 14868 8168
rect 14802 8088 14868 8104
rect 14802 8024 14803 8088
rect 14867 8024 14868 8088
rect 14802 8008 14868 8024
rect 14802 7944 14803 8008
rect 14867 7944 14868 8008
rect 14802 7928 14868 7944
rect 14802 7864 14803 7928
rect 14867 7864 14868 7928
rect 14802 7848 14868 7864
rect 14802 7784 14803 7848
rect 14867 7784 14868 7848
rect 14802 7768 14868 7784
rect 14802 7704 14803 7768
rect 14867 7704 14868 7768
rect 14802 7614 14868 7704
rect 14928 7610 14988 8642
rect 15048 7550 15108 8580
rect 15168 7610 15228 8642
rect 15288 7550 15348 8580
rect 15408 8488 15474 8642
rect 15408 8424 15409 8488
rect 15473 8424 15474 8488
rect 15408 8408 15474 8424
rect 15408 8344 15409 8408
rect 15473 8344 15474 8408
rect 15408 8328 15474 8344
rect 15408 8264 15409 8328
rect 15473 8264 15474 8328
rect 15408 8248 15474 8264
rect 15408 8184 15409 8248
rect 15473 8184 15474 8248
rect 15408 8168 15474 8184
rect 15408 8104 15409 8168
rect 15473 8104 15474 8168
rect 15408 8088 15474 8104
rect 15408 8024 15409 8088
rect 15473 8024 15474 8088
rect 15408 8008 15474 8024
rect 15408 7944 15409 8008
rect 15473 7944 15474 8008
rect 15408 7928 15474 7944
rect 15408 7864 15409 7928
rect 15473 7864 15474 7928
rect 15408 7848 15474 7864
rect 15408 7784 15409 7848
rect 15473 7784 15474 7848
rect 15408 7768 15474 7784
rect 15408 7704 15409 7768
rect 15473 7704 15474 7768
rect 15408 7614 15474 7704
rect 15534 7550 15594 8580
rect 15654 7610 15714 8642
rect 15774 7550 15834 8580
rect 15894 7610 15954 8642
rect 16014 8488 16080 8642
rect 16014 8424 16015 8488
rect 16079 8424 16080 8488
rect 16014 8408 16080 8424
rect 16014 8344 16015 8408
rect 16079 8344 16080 8408
rect 16014 8328 16080 8344
rect 16014 8264 16015 8328
rect 16079 8264 16080 8328
rect 16014 8248 16080 8264
rect 16014 8184 16015 8248
rect 16079 8184 16080 8248
rect 16014 8168 16080 8184
rect 16014 8104 16015 8168
rect 16079 8104 16080 8168
rect 16014 8088 16080 8104
rect 16014 8024 16015 8088
rect 16079 8024 16080 8088
rect 16014 8008 16080 8024
rect 16014 7944 16015 8008
rect 16079 7944 16080 8008
rect 16014 7928 16080 7944
rect 16014 7864 16015 7928
rect 16079 7864 16080 7928
rect 16014 7848 16080 7864
rect 16014 7784 16015 7848
rect 16079 7784 16080 7848
rect 16014 7768 16080 7784
rect 16014 7704 16015 7768
rect 16079 7704 16080 7768
rect 16014 7614 16080 7704
rect 16140 7610 16200 8642
rect 16260 7550 16320 8580
rect 16380 7610 16440 8642
rect 16500 7550 16560 8580
rect 16620 8488 16686 8642
rect 16620 8424 16621 8488
rect 16685 8424 16686 8488
rect 16620 8408 16686 8424
rect 16620 8344 16621 8408
rect 16685 8344 16686 8408
rect 16620 8328 16686 8344
rect 16620 8264 16621 8328
rect 16685 8264 16686 8328
rect 16620 8248 16686 8264
rect 16620 8184 16621 8248
rect 16685 8184 16686 8248
rect 16620 8168 16686 8184
rect 16620 8104 16621 8168
rect 16685 8104 16686 8168
rect 16620 8088 16686 8104
rect 16620 8024 16621 8088
rect 16685 8024 16686 8088
rect 16620 8008 16686 8024
rect 16620 7944 16621 8008
rect 16685 7944 16686 8008
rect 16620 7928 16686 7944
rect 16620 7864 16621 7928
rect 16685 7864 16686 7928
rect 16620 7848 16686 7864
rect 16620 7784 16621 7848
rect 16685 7784 16686 7848
rect 16620 7768 16686 7784
rect 16620 7704 16621 7768
rect 16685 7704 16686 7768
rect 16620 7614 16686 7704
rect 16746 7550 16806 8580
rect 16866 7610 16926 8642
rect 16986 7550 17046 8580
rect 17106 7610 17166 8642
rect 17226 8488 17292 8642
rect 17226 8424 17227 8488
rect 17291 8424 17292 8488
rect 17226 8408 17292 8424
rect 17226 8344 17227 8408
rect 17291 8344 17292 8408
rect 17226 8328 17292 8344
rect 17226 8264 17227 8328
rect 17291 8264 17292 8328
rect 17226 8248 17292 8264
rect 17226 8184 17227 8248
rect 17291 8184 17292 8248
rect 17226 8168 17292 8184
rect 17226 8104 17227 8168
rect 17291 8104 17292 8168
rect 17226 8088 17292 8104
rect 17226 8024 17227 8088
rect 17291 8024 17292 8088
rect 17226 8008 17292 8024
rect 17226 7944 17227 8008
rect 17291 7944 17292 8008
rect 17226 7928 17292 7944
rect 17226 7864 17227 7928
rect 17291 7864 17292 7928
rect 17226 7848 17292 7864
rect 17226 7784 17227 7848
rect 17291 7784 17292 7848
rect 17226 7768 17292 7784
rect 17226 7704 17227 7768
rect 17291 7704 17292 7768
rect 17226 7614 17292 7704
rect 17352 7610 17412 8642
rect 17472 7550 17532 8580
rect 17592 7610 17652 8642
rect 17712 7550 17772 8580
rect 17832 8488 17898 8642
rect 17832 8424 17833 8488
rect 17897 8424 17898 8488
rect 17832 8408 17898 8424
rect 17832 8344 17833 8408
rect 17897 8344 17898 8408
rect 17832 8328 17898 8344
rect 17832 8264 17833 8328
rect 17897 8264 17898 8328
rect 17832 8248 17898 8264
rect 17832 8184 17833 8248
rect 17897 8184 17898 8248
rect 17832 8168 17898 8184
rect 17832 8104 17833 8168
rect 17897 8104 17898 8168
rect 17832 8088 17898 8104
rect 17832 8024 17833 8088
rect 17897 8024 17898 8088
rect 17832 8008 17898 8024
rect 17832 7944 17833 8008
rect 17897 7944 17898 8008
rect 17832 7928 17898 7944
rect 17832 7864 17833 7928
rect 17897 7864 17898 7928
rect 17832 7848 17898 7864
rect 17832 7784 17833 7848
rect 17897 7784 17898 7848
rect 17832 7768 17898 7784
rect 17832 7704 17833 7768
rect 17897 7704 17898 7768
rect 17832 7614 17898 7704
rect 17958 7550 18018 8580
rect 18078 7610 18138 8642
rect 18198 7550 18258 8580
rect 18318 7610 18378 8642
rect 18438 8488 18504 8642
rect 18438 8424 18439 8488
rect 18503 8424 18504 8488
rect 18438 8408 18504 8424
rect 18438 8344 18439 8408
rect 18503 8344 18504 8408
rect 18438 8328 18504 8344
rect 18438 8264 18439 8328
rect 18503 8264 18504 8328
rect 18438 8248 18504 8264
rect 18438 8184 18439 8248
rect 18503 8184 18504 8248
rect 18438 8168 18504 8184
rect 18438 8104 18439 8168
rect 18503 8104 18504 8168
rect 18438 8088 18504 8104
rect 18438 8024 18439 8088
rect 18503 8024 18504 8088
rect 18438 8008 18504 8024
rect 18438 7944 18439 8008
rect 18503 7944 18504 8008
rect 18438 7928 18504 7944
rect 18438 7864 18439 7928
rect 18503 7864 18504 7928
rect 18438 7848 18504 7864
rect 18438 7784 18439 7848
rect 18503 7784 18504 7848
rect 18438 7768 18504 7784
rect 18438 7704 18439 7768
rect 18503 7704 18504 7768
rect 18438 7614 18504 7704
rect 18564 8647 18668 8711
rect 18743 8670 18748 8711
rect 18732 8647 18748 8670
rect 18812 8647 18828 8711
rect 18892 8647 18908 8711
rect 18972 8647 18988 8711
rect 19052 8647 19068 8711
rect 19132 8647 19236 8711
rect 18564 8645 19236 8647
rect 18564 8491 18630 8645
rect 18564 8427 18565 8491
rect 18629 8427 18630 8491
rect 18564 8411 18630 8427
rect 18564 8347 18565 8411
rect 18629 8347 18630 8411
rect 18564 8331 18630 8347
rect 18564 8267 18565 8331
rect 18629 8267 18630 8331
rect 18564 8251 18630 8267
rect 18564 8187 18565 8251
rect 18629 8187 18630 8251
rect 18564 8171 18630 8187
rect 18564 8107 18565 8171
rect 18629 8107 18630 8171
rect 18564 8091 18630 8107
rect 18564 8027 18565 8091
rect 18629 8027 18630 8091
rect 18564 8011 18630 8027
rect 18564 7947 18565 8011
rect 18629 7947 18630 8011
rect 18564 7931 18630 7947
rect 18564 7867 18565 7931
rect 18629 7867 18630 7931
rect 18564 7851 18630 7867
rect 18564 7787 18565 7851
rect 18629 7787 18630 7851
rect 18564 7771 18630 7787
rect 18564 7707 18565 7771
rect 18629 7707 18630 7771
rect 18564 7617 18630 7707
rect 18690 7553 18750 8583
rect 18810 7613 18870 8645
rect 18930 7553 18990 8583
rect 19050 7613 19110 8645
rect 19170 8491 19236 8645
rect 19462 8692 19835 8709
rect 19462 8628 19501 8692
rect 19565 8628 19644 8692
rect 19708 8628 19764 8692
rect 19828 8628 19835 8692
rect 20023 8665 20054 8729
rect 20118 8665 20149 8729
rect 20782 8731 20865 8736
rect 20782 8710 20792 8731
rect 20023 8655 20149 8665
rect 20299 8708 20792 8710
rect 20856 8710 20865 8731
rect 21011 8731 21094 8736
rect 21011 8710 21020 8731
rect 20856 8708 21020 8710
rect 21084 8710 21094 8731
rect 21994 8731 22077 8736
rect 21994 8710 22004 8731
rect 21084 8708 22004 8710
rect 22068 8710 22077 8731
rect 22223 8731 22306 8736
rect 22223 8710 22232 8731
rect 22068 8708 22232 8710
rect 22296 8710 22306 8731
rect 23206 8731 23289 8736
rect 23206 8710 23216 8731
rect 22296 8708 23216 8710
rect 23280 8710 23289 8731
rect 23435 8731 23518 8736
rect 23435 8710 23444 8731
rect 23280 8708 23444 8710
rect 23508 8710 23518 8731
rect 24418 8731 24501 8736
rect 24418 8710 24428 8731
rect 23508 8708 24428 8710
rect 24492 8710 24501 8731
rect 24647 8731 24730 8736
rect 24647 8710 24656 8731
rect 24492 8708 24656 8710
rect 24720 8710 24730 8731
rect 25379 8734 25462 8739
rect 25379 8713 25388 8734
rect 25273 8711 25388 8713
rect 25452 8713 25462 8734
rect 25452 8711 25945 8713
rect 24720 8708 25213 8710
rect 19462 8613 19835 8628
rect 20299 8644 20403 8708
rect 20467 8644 20483 8708
rect 20547 8644 20563 8708
rect 20627 8644 20643 8708
rect 20707 8644 20723 8708
rect 20787 8667 20792 8708
rect 20787 8644 20803 8667
rect 20867 8644 21009 8708
rect 21084 8667 21089 8708
rect 21073 8644 21089 8667
rect 21153 8644 21169 8708
rect 21233 8644 21249 8708
rect 21313 8644 21329 8708
rect 21393 8644 21409 8708
rect 21473 8644 21615 8708
rect 21679 8644 21695 8708
rect 21759 8644 21775 8708
rect 21839 8644 21855 8708
rect 21919 8644 21935 8708
rect 21999 8667 22004 8708
rect 21999 8644 22015 8667
rect 22079 8644 22221 8708
rect 22296 8667 22301 8708
rect 22285 8644 22301 8667
rect 22365 8644 22381 8708
rect 22445 8644 22461 8708
rect 22525 8644 22541 8708
rect 22605 8644 22621 8708
rect 22685 8644 22827 8708
rect 22891 8644 22907 8708
rect 22971 8644 22987 8708
rect 23051 8644 23067 8708
rect 23131 8644 23147 8708
rect 23211 8667 23216 8708
rect 23211 8644 23227 8667
rect 23291 8644 23433 8708
rect 23508 8667 23513 8708
rect 23497 8644 23513 8667
rect 23577 8644 23593 8708
rect 23657 8644 23673 8708
rect 23737 8644 23753 8708
rect 23817 8644 23833 8708
rect 23897 8644 24039 8708
rect 24103 8644 24119 8708
rect 24183 8644 24199 8708
rect 24263 8644 24279 8708
rect 24343 8644 24359 8708
rect 24423 8667 24428 8708
rect 24423 8644 24439 8667
rect 24503 8644 24645 8708
rect 24720 8667 24725 8708
rect 24709 8644 24725 8667
rect 24789 8644 24805 8708
rect 24869 8644 24885 8708
rect 24949 8644 24965 8708
rect 25029 8644 25045 8708
rect 25109 8644 25213 8708
rect 20299 8642 25213 8644
rect 19629 8612 19721 8613
rect 19170 8427 19171 8491
rect 19235 8427 19236 8491
rect 20299 8488 20365 8642
rect 19170 8411 19236 8427
rect 19170 8347 19171 8411
rect 19235 8347 19236 8411
rect 20111 8468 20237 8478
rect 20111 8404 20142 8468
rect 20206 8404 20237 8468
rect 20111 8394 20237 8404
rect 20299 8424 20300 8488
rect 20364 8424 20365 8488
rect 20299 8408 20365 8424
rect 19170 8331 19236 8347
rect 19170 8267 19171 8331
rect 19235 8267 19236 8331
rect 19170 8251 19236 8267
rect 19170 8187 19171 8251
rect 19235 8187 19236 8251
rect 20299 8344 20300 8408
rect 20364 8344 20365 8408
rect 20299 8328 20365 8344
rect 20299 8264 20300 8328
rect 20364 8264 20365 8328
rect 20299 8248 20365 8264
rect 19170 8171 19236 8187
rect 19170 8107 19171 8171
rect 19235 8107 19236 8171
rect 20029 8226 20155 8236
rect 19612 8163 19756 8164
rect 19170 8091 19236 8107
rect 19170 8027 19171 8091
rect 19235 8027 19236 8091
rect 19468 8147 19861 8163
rect 20029 8162 20060 8226
rect 20124 8162 20155 8226
rect 20029 8152 20155 8162
rect 20299 8184 20300 8248
rect 20364 8184 20365 8248
rect 20299 8168 20365 8184
rect 19468 8146 19651 8147
rect 19468 8082 19507 8146
rect 19571 8083 19651 8146
rect 19715 8146 19861 8147
rect 19715 8083 19782 8146
rect 19571 8082 19782 8083
rect 19846 8082 19861 8146
rect 19468 8068 19861 8082
rect 20299 8104 20300 8168
rect 20364 8104 20365 8168
rect 20299 8088 20365 8104
rect 19468 8067 19612 8068
rect 19743 8067 19861 8068
rect 20028 8069 20154 8079
rect 19170 8011 19236 8027
rect 19170 7947 19171 8011
rect 19235 7947 19236 8011
rect 19170 7931 19236 7947
rect 19170 7867 19171 7931
rect 19235 7867 19236 7931
rect 19606 7997 19732 8007
rect 19606 7933 19637 7997
rect 19701 7933 19732 7997
rect 20028 8005 20059 8069
rect 20123 8005 20154 8069
rect 20028 7995 20154 8005
rect 20299 8024 20300 8088
rect 20364 8024 20365 8088
rect 20299 8008 20365 8024
rect 19606 7923 19732 7933
rect 20299 7944 20300 8008
rect 20364 7944 20365 8008
rect 20299 7928 20365 7944
rect 19170 7851 19236 7867
rect 19170 7787 19171 7851
rect 19235 7787 19236 7851
rect 20028 7899 20154 7909
rect 20028 7835 20059 7899
rect 20123 7835 20154 7899
rect 20028 7825 20154 7835
rect 20299 7864 20300 7928
rect 20364 7864 20365 7928
rect 20299 7848 20365 7864
rect 19170 7771 19236 7787
rect 19170 7707 19171 7771
rect 19235 7707 19236 7771
rect 19606 7801 19732 7811
rect 19606 7737 19637 7801
rect 19701 7737 19732 7801
rect 20299 7784 20300 7848
rect 20364 7784 20365 7848
rect 20299 7768 20365 7784
rect 19606 7727 19732 7737
rect 20029 7747 20155 7757
rect 19170 7617 19236 7707
rect 20029 7683 20060 7747
rect 20124 7683 20155 7747
rect 20029 7673 20155 7683
rect 20299 7704 20300 7768
rect 20364 7704 20365 7768
rect 19606 7626 19732 7636
rect 19606 7562 19637 7626
rect 19701 7562 19732 7626
rect 20299 7614 20365 7704
rect 18564 7551 19236 7553
rect 19606 7552 19732 7562
rect 20034 7603 20160 7613
rect 20425 7610 20485 8642
rect 13325 7529 13451 7539
rect 13590 7548 18504 7550
rect 3787 7494 8701 7496
rect 3031 7479 3157 7489
rect 13590 7484 13694 7548
rect 13758 7484 13774 7548
rect 13838 7484 13854 7548
rect 13918 7484 13934 7548
rect 13998 7484 14014 7548
rect 14078 7484 14094 7548
rect 14158 7484 14300 7548
rect 14364 7484 14380 7548
rect 14444 7484 14460 7548
rect 14524 7484 14540 7548
rect 14604 7484 14620 7548
rect 14684 7484 14700 7548
rect 14764 7484 14906 7548
rect 14970 7484 14986 7548
rect 15050 7484 15066 7548
rect 15130 7484 15146 7548
rect 15210 7484 15226 7548
rect 15290 7484 15306 7548
rect 15370 7484 15512 7548
rect 15576 7484 15592 7548
rect 15656 7484 15672 7548
rect 15736 7484 15752 7548
rect 15816 7484 15832 7548
rect 15896 7484 15912 7548
rect 15976 7484 16118 7548
rect 16182 7484 16198 7548
rect 16262 7484 16278 7548
rect 16342 7484 16358 7548
rect 16422 7484 16438 7548
rect 16502 7484 16518 7548
rect 16582 7484 16724 7548
rect 16788 7484 16804 7548
rect 16868 7484 16884 7548
rect 16948 7484 16964 7548
rect 17028 7484 17044 7548
rect 17108 7484 17124 7548
rect 17188 7484 17330 7548
rect 17394 7484 17410 7548
rect 17474 7484 17490 7548
rect 17554 7484 17570 7548
rect 17634 7484 17650 7548
rect 17714 7484 17730 7548
rect 17794 7484 17936 7548
rect 18000 7484 18016 7548
rect 18080 7484 18096 7548
rect 18160 7484 18176 7548
rect 18240 7484 18256 7548
rect 18320 7484 18336 7548
rect 18400 7484 18504 7548
rect 18564 7487 18668 7551
rect 18732 7487 18748 7551
rect 18812 7487 18828 7551
rect 18892 7487 18908 7551
rect 18972 7487 18988 7551
rect 19052 7487 19068 7551
rect 19132 7550 19236 7551
rect 19132 7541 19260 7550
rect 19132 7487 19165 7541
rect 18564 7485 19165 7487
rect 13590 7482 18504 7484
rect 19134 7477 19165 7485
rect 19229 7477 19260 7541
rect 20034 7539 20065 7603
rect 20129 7539 20160 7603
rect 20545 7550 20605 8580
rect 20665 7610 20725 8642
rect 20785 7550 20845 8580
rect 20905 8488 20971 8642
rect 20905 8424 20906 8488
rect 20970 8424 20971 8488
rect 20905 8408 20971 8424
rect 20905 8344 20906 8408
rect 20970 8344 20971 8408
rect 20905 8328 20971 8344
rect 20905 8264 20906 8328
rect 20970 8264 20971 8328
rect 20905 8248 20971 8264
rect 20905 8184 20906 8248
rect 20970 8184 20971 8248
rect 20905 8168 20971 8184
rect 20905 8104 20906 8168
rect 20970 8104 20971 8168
rect 20905 8088 20971 8104
rect 20905 8024 20906 8088
rect 20970 8024 20971 8088
rect 20905 8008 20971 8024
rect 20905 7944 20906 8008
rect 20970 7944 20971 8008
rect 20905 7928 20971 7944
rect 20905 7864 20906 7928
rect 20970 7864 20971 7928
rect 20905 7848 20971 7864
rect 20905 7784 20906 7848
rect 20970 7784 20971 7848
rect 20905 7768 20971 7784
rect 20905 7704 20906 7768
rect 20970 7704 20971 7768
rect 20905 7614 20971 7704
rect 21031 7550 21091 8580
rect 21151 7610 21211 8642
rect 21271 7550 21331 8580
rect 21391 7610 21451 8642
rect 21511 8488 21577 8642
rect 21511 8424 21512 8488
rect 21576 8424 21577 8488
rect 21511 8408 21577 8424
rect 21511 8344 21512 8408
rect 21576 8344 21577 8408
rect 21511 8328 21577 8344
rect 21511 8264 21512 8328
rect 21576 8264 21577 8328
rect 21511 8248 21577 8264
rect 21511 8184 21512 8248
rect 21576 8184 21577 8248
rect 21511 8168 21577 8184
rect 21511 8104 21512 8168
rect 21576 8104 21577 8168
rect 21511 8088 21577 8104
rect 21511 8024 21512 8088
rect 21576 8024 21577 8088
rect 21511 8008 21577 8024
rect 21511 7944 21512 8008
rect 21576 7944 21577 8008
rect 21511 7928 21577 7944
rect 21511 7864 21512 7928
rect 21576 7864 21577 7928
rect 21511 7848 21577 7864
rect 21511 7784 21512 7848
rect 21576 7784 21577 7848
rect 21511 7768 21577 7784
rect 21511 7704 21512 7768
rect 21576 7704 21577 7768
rect 21511 7614 21577 7704
rect 21637 7610 21697 8642
rect 21757 7550 21817 8580
rect 21877 7610 21937 8642
rect 21997 7550 22057 8580
rect 22117 8488 22183 8642
rect 22117 8424 22118 8488
rect 22182 8424 22183 8488
rect 22117 8408 22183 8424
rect 22117 8344 22118 8408
rect 22182 8344 22183 8408
rect 22117 8328 22183 8344
rect 22117 8264 22118 8328
rect 22182 8264 22183 8328
rect 22117 8248 22183 8264
rect 22117 8184 22118 8248
rect 22182 8184 22183 8248
rect 22117 8168 22183 8184
rect 22117 8104 22118 8168
rect 22182 8104 22183 8168
rect 22117 8088 22183 8104
rect 22117 8024 22118 8088
rect 22182 8024 22183 8088
rect 22117 8008 22183 8024
rect 22117 7944 22118 8008
rect 22182 7944 22183 8008
rect 22117 7928 22183 7944
rect 22117 7864 22118 7928
rect 22182 7864 22183 7928
rect 22117 7848 22183 7864
rect 22117 7784 22118 7848
rect 22182 7784 22183 7848
rect 22117 7768 22183 7784
rect 22117 7704 22118 7768
rect 22182 7704 22183 7768
rect 22117 7614 22183 7704
rect 22243 7550 22303 8580
rect 22363 7610 22423 8642
rect 22483 7550 22543 8580
rect 22603 7610 22663 8642
rect 22723 8488 22789 8642
rect 22723 8424 22724 8488
rect 22788 8424 22789 8488
rect 22723 8408 22789 8424
rect 22723 8344 22724 8408
rect 22788 8344 22789 8408
rect 22723 8328 22789 8344
rect 22723 8264 22724 8328
rect 22788 8264 22789 8328
rect 22723 8248 22789 8264
rect 22723 8184 22724 8248
rect 22788 8184 22789 8248
rect 22723 8168 22789 8184
rect 22723 8104 22724 8168
rect 22788 8104 22789 8168
rect 22723 8088 22789 8104
rect 22723 8024 22724 8088
rect 22788 8024 22789 8088
rect 22723 8008 22789 8024
rect 22723 7944 22724 8008
rect 22788 7944 22789 8008
rect 22723 7928 22789 7944
rect 22723 7864 22724 7928
rect 22788 7864 22789 7928
rect 22723 7848 22789 7864
rect 22723 7784 22724 7848
rect 22788 7784 22789 7848
rect 22723 7768 22789 7784
rect 22723 7704 22724 7768
rect 22788 7704 22789 7768
rect 22723 7614 22789 7704
rect 22849 7610 22909 8642
rect 22969 7550 23029 8580
rect 23089 7610 23149 8642
rect 23209 7550 23269 8580
rect 23329 8488 23395 8642
rect 23329 8424 23330 8488
rect 23394 8424 23395 8488
rect 23329 8408 23395 8424
rect 23329 8344 23330 8408
rect 23394 8344 23395 8408
rect 23329 8328 23395 8344
rect 23329 8264 23330 8328
rect 23394 8264 23395 8328
rect 23329 8248 23395 8264
rect 23329 8184 23330 8248
rect 23394 8184 23395 8248
rect 23329 8168 23395 8184
rect 23329 8104 23330 8168
rect 23394 8104 23395 8168
rect 23329 8088 23395 8104
rect 23329 8024 23330 8088
rect 23394 8024 23395 8088
rect 23329 8008 23395 8024
rect 23329 7944 23330 8008
rect 23394 7944 23395 8008
rect 23329 7928 23395 7944
rect 23329 7864 23330 7928
rect 23394 7864 23395 7928
rect 23329 7848 23395 7864
rect 23329 7784 23330 7848
rect 23394 7784 23395 7848
rect 23329 7768 23395 7784
rect 23329 7704 23330 7768
rect 23394 7704 23395 7768
rect 23329 7614 23395 7704
rect 23455 7550 23515 8580
rect 23575 7610 23635 8642
rect 23695 7550 23755 8580
rect 23815 7610 23875 8642
rect 23935 8488 24001 8642
rect 23935 8424 23936 8488
rect 24000 8424 24001 8488
rect 23935 8408 24001 8424
rect 23935 8344 23936 8408
rect 24000 8344 24001 8408
rect 23935 8328 24001 8344
rect 23935 8264 23936 8328
rect 24000 8264 24001 8328
rect 23935 8248 24001 8264
rect 23935 8184 23936 8248
rect 24000 8184 24001 8248
rect 23935 8168 24001 8184
rect 23935 8104 23936 8168
rect 24000 8104 24001 8168
rect 23935 8088 24001 8104
rect 23935 8024 23936 8088
rect 24000 8024 24001 8088
rect 23935 8008 24001 8024
rect 23935 7944 23936 8008
rect 24000 7944 24001 8008
rect 23935 7928 24001 7944
rect 23935 7864 23936 7928
rect 24000 7864 24001 7928
rect 23935 7848 24001 7864
rect 23935 7784 23936 7848
rect 24000 7784 24001 7848
rect 23935 7768 24001 7784
rect 23935 7704 23936 7768
rect 24000 7704 24001 7768
rect 23935 7614 24001 7704
rect 24061 7610 24121 8642
rect 24181 7550 24241 8580
rect 24301 7610 24361 8642
rect 24421 7550 24481 8580
rect 24541 8488 24607 8642
rect 24541 8424 24542 8488
rect 24606 8424 24607 8488
rect 24541 8408 24607 8424
rect 24541 8344 24542 8408
rect 24606 8344 24607 8408
rect 24541 8328 24607 8344
rect 24541 8264 24542 8328
rect 24606 8264 24607 8328
rect 24541 8248 24607 8264
rect 24541 8184 24542 8248
rect 24606 8184 24607 8248
rect 24541 8168 24607 8184
rect 24541 8104 24542 8168
rect 24606 8104 24607 8168
rect 24541 8088 24607 8104
rect 24541 8024 24542 8088
rect 24606 8024 24607 8088
rect 24541 8008 24607 8024
rect 24541 7944 24542 8008
rect 24606 7944 24607 8008
rect 24541 7928 24607 7944
rect 24541 7864 24542 7928
rect 24606 7864 24607 7928
rect 24541 7848 24607 7864
rect 24541 7784 24542 7848
rect 24606 7784 24607 7848
rect 24541 7768 24607 7784
rect 24541 7704 24542 7768
rect 24606 7704 24607 7768
rect 24541 7614 24607 7704
rect 24667 7550 24727 8580
rect 24787 7610 24847 8642
rect 24907 7550 24967 8580
rect 25027 7610 25087 8642
rect 25147 8488 25213 8642
rect 25147 8424 25148 8488
rect 25212 8424 25213 8488
rect 25147 8408 25213 8424
rect 25147 8344 25148 8408
rect 25212 8344 25213 8408
rect 25147 8328 25213 8344
rect 25147 8264 25148 8328
rect 25212 8264 25213 8328
rect 25147 8248 25213 8264
rect 25147 8184 25148 8248
rect 25212 8184 25213 8248
rect 25147 8168 25213 8184
rect 25147 8104 25148 8168
rect 25212 8104 25213 8168
rect 25147 8088 25213 8104
rect 25147 8024 25148 8088
rect 25212 8024 25213 8088
rect 25147 8008 25213 8024
rect 25147 7944 25148 8008
rect 25212 7944 25213 8008
rect 25147 7928 25213 7944
rect 25147 7864 25148 7928
rect 25212 7864 25213 7928
rect 25147 7848 25213 7864
rect 25147 7784 25148 7848
rect 25212 7784 25213 7848
rect 25147 7768 25213 7784
rect 25147 7704 25148 7768
rect 25212 7704 25213 7768
rect 25147 7614 25213 7704
rect 25273 8647 25377 8711
rect 25452 8670 25457 8711
rect 25441 8647 25457 8670
rect 25521 8647 25537 8711
rect 25601 8647 25617 8711
rect 25681 8647 25697 8711
rect 25761 8647 25777 8711
rect 25841 8647 25945 8711
rect 25273 8645 25945 8647
rect 25273 8491 25339 8645
rect 25273 8427 25274 8491
rect 25338 8427 25339 8491
rect 25273 8411 25339 8427
rect 25273 8347 25274 8411
rect 25338 8347 25339 8411
rect 25273 8331 25339 8347
rect 25273 8267 25274 8331
rect 25338 8267 25339 8331
rect 25273 8251 25339 8267
rect 25273 8187 25274 8251
rect 25338 8187 25339 8251
rect 25273 8171 25339 8187
rect 25273 8107 25274 8171
rect 25338 8107 25339 8171
rect 25273 8091 25339 8107
rect 25273 8027 25274 8091
rect 25338 8027 25339 8091
rect 25273 8011 25339 8027
rect 25273 7947 25274 8011
rect 25338 7947 25339 8011
rect 25273 7931 25339 7947
rect 25273 7867 25274 7931
rect 25338 7867 25339 7931
rect 25273 7851 25339 7867
rect 25273 7787 25274 7851
rect 25338 7787 25339 7851
rect 25273 7771 25339 7787
rect 25273 7707 25274 7771
rect 25338 7707 25339 7771
rect 25273 7617 25339 7707
rect 25399 7553 25459 8583
rect 25519 7613 25579 8645
rect 25639 7553 25699 8583
rect 25759 7613 25819 8645
rect 25879 8491 25945 8645
rect 26171 8692 26544 8709
rect 26171 8628 26210 8692
rect 26274 8628 26353 8692
rect 26417 8628 26473 8692
rect 26537 8628 26544 8692
rect 26171 8613 26544 8628
rect 26338 8612 26430 8613
rect 25879 8427 25880 8491
rect 25944 8427 25945 8491
rect 25879 8411 25945 8427
rect 25879 8347 25880 8411
rect 25944 8347 25945 8411
rect 25879 8331 25945 8347
rect 25879 8267 25880 8331
rect 25944 8267 25945 8331
rect 25879 8251 25945 8267
rect 25879 8187 25880 8251
rect 25944 8187 25945 8251
rect 25879 8171 25945 8187
rect 25879 8107 25880 8171
rect 25944 8107 25945 8171
rect 26321 8163 26465 8164
rect 25879 8091 25945 8107
rect 25879 8027 25880 8091
rect 25944 8027 25945 8091
rect 26177 8147 26570 8163
rect 26177 8146 26360 8147
rect 26177 8082 26216 8146
rect 26280 8083 26360 8146
rect 26424 8146 26570 8147
rect 26424 8083 26491 8146
rect 26280 8082 26491 8083
rect 26555 8082 26570 8146
rect 26177 8068 26570 8082
rect 26177 8067 26321 8068
rect 26452 8067 26570 8068
rect 25879 8011 25945 8027
rect 25879 7947 25880 8011
rect 25944 7947 25945 8011
rect 25879 7931 25945 7947
rect 25879 7867 25880 7931
rect 25944 7867 25945 7931
rect 25879 7851 25945 7867
rect 25879 7787 25880 7851
rect 25944 7787 25945 7851
rect 25879 7771 25945 7787
rect 25879 7707 25880 7771
rect 25944 7707 25945 7771
rect 25879 7617 25945 7707
rect 25273 7551 25945 7553
rect 20034 7529 20160 7539
rect 20299 7548 25213 7550
rect 20299 7484 20403 7548
rect 20467 7484 20483 7548
rect 20547 7484 20563 7548
rect 20627 7484 20643 7548
rect 20707 7484 20723 7548
rect 20787 7484 20803 7548
rect 20867 7484 21009 7548
rect 21073 7484 21089 7548
rect 21153 7484 21169 7548
rect 21233 7484 21249 7548
rect 21313 7484 21329 7548
rect 21393 7484 21409 7548
rect 21473 7484 21615 7548
rect 21679 7484 21695 7548
rect 21759 7484 21775 7548
rect 21839 7484 21855 7548
rect 21919 7484 21935 7548
rect 21999 7484 22015 7548
rect 22079 7484 22221 7548
rect 22285 7484 22301 7548
rect 22365 7484 22381 7548
rect 22445 7484 22461 7548
rect 22525 7484 22541 7548
rect 22605 7484 22621 7548
rect 22685 7484 22827 7548
rect 22891 7484 22907 7548
rect 22971 7484 22987 7548
rect 23051 7484 23067 7548
rect 23131 7484 23147 7548
rect 23211 7484 23227 7548
rect 23291 7484 23433 7548
rect 23497 7484 23513 7548
rect 23577 7484 23593 7548
rect 23657 7484 23673 7548
rect 23737 7484 23753 7548
rect 23817 7484 23833 7548
rect 23897 7484 24039 7548
rect 24103 7484 24119 7548
rect 24183 7484 24199 7548
rect 24263 7484 24279 7548
rect 24343 7484 24359 7548
rect 24423 7484 24439 7548
rect 24503 7484 24645 7548
rect 24709 7484 24725 7548
rect 24789 7484 24805 7548
rect 24869 7484 24885 7548
rect 24949 7484 24965 7548
rect 25029 7484 25045 7548
rect 25109 7484 25213 7548
rect 25273 7487 25377 7551
rect 25441 7487 25457 7551
rect 25521 7487 25537 7551
rect 25601 7487 25617 7551
rect 25681 7487 25697 7551
rect 25761 7487 25777 7551
rect 25841 7550 25945 7551
rect 25841 7541 25969 7550
rect 25841 7487 25874 7541
rect 25273 7485 25874 7487
rect 20299 7482 25213 7484
rect 19134 7467 19260 7477
rect 25843 7477 25874 7485
rect 25938 7477 25969 7541
rect 25843 7467 25969 7477
rect 24644 7335 24770 7345
rect 24644 7271 24675 7335
rect 24739 7327 24770 7335
rect 25400 7328 30314 7330
rect 24739 7325 25340 7327
rect 24739 7271 24772 7325
rect 24644 7262 24772 7271
rect 24668 7261 24772 7262
rect 24836 7261 24852 7325
rect 24916 7261 24932 7325
rect 24996 7261 25012 7325
rect 25076 7261 25092 7325
rect 25156 7261 25172 7325
rect 25236 7261 25340 7325
rect 25400 7264 25504 7328
rect 25568 7264 25584 7328
rect 25648 7264 25664 7328
rect 25728 7264 25744 7328
rect 25808 7264 25824 7328
rect 25888 7264 25904 7328
rect 25968 7264 26110 7328
rect 26174 7264 26190 7328
rect 26254 7264 26270 7328
rect 26334 7264 26350 7328
rect 26414 7264 26430 7328
rect 26494 7264 26510 7328
rect 26574 7264 26716 7328
rect 26780 7264 26796 7328
rect 26860 7264 26876 7328
rect 26940 7264 26956 7328
rect 27020 7264 27036 7328
rect 27100 7264 27116 7328
rect 27180 7264 27322 7328
rect 27386 7264 27402 7328
rect 27466 7264 27482 7328
rect 27546 7264 27562 7328
rect 27626 7264 27642 7328
rect 27706 7264 27722 7328
rect 27786 7264 27928 7328
rect 27992 7264 28008 7328
rect 28072 7264 28088 7328
rect 28152 7264 28168 7328
rect 28232 7264 28248 7328
rect 28312 7264 28328 7328
rect 28392 7264 28534 7328
rect 28598 7264 28614 7328
rect 28678 7264 28694 7328
rect 28758 7264 28774 7328
rect 28838 7264 28854 7328
rect 28918 7264 28934 7328
rect 28998 7264 29140 7328
rect 29204 7264 29220 7328
rect 29284 7264 29300 7328
rect 29364 7264 29380 7328
rect 29444 7264 29460 7328
rect 29524 7264 29540 7328
rect 29604 7264 29746 7328
rect 29810 7264 29826 7328
rect 29890 7264 29906 7328
rect 29970 7264 29986 7328
rect 30050 7264 30066 7328
rect 30130 7264 30146 7328
rect 30210 7264 30314 7328
rect 25400 7262 30314 7264
rect 30453 7273 30579 7283
rect 24668 7259 25340 7261
rect 24668 7105 24734 7195
rect 10881 7080 11053 7090
rect 10881 6934 10891 7080
rect 11041 6934 11053 7080
rect 10881 6924 11053 6934
rect 11193 7064 11365 7074
rect 11193 6918 11203 7064
rect 11353 6918 11365 7064
rect 11193 6908 11365 6918
rect 24668 7041 24669 7105
rect 24733 7041 24734 7105
rect 24668 7025 24734 7041
rect 24668 6961 24669 7025
rect 24733 6961 24734 7025
rect 24668 6945 24734 6961
rect 24668 6881 24669 6945
rect 24733 6881 24734 6945
rect 24668 6865 24734 6881
rect 24668 6801 24669 6865
rect 24733 6801 24734 6865
rect 24668 6785 24734 6801
rect 24043 6744 24161 6745
rect 24292 6744 24436 6745
rect 24043 6730 24436 6744
rect 24043 6666 24058 6730
rect 24122 6729 24333 6730
rect 24122 6666 24189 6729
rect 24043 6665 24189 6666
rect 24253 6666 24333 6729
rect 24397 6666 24436 6730
rect 24253 6665 24436 6666
rect 24043 6649 24436 6665
rect 24668 6721 24669 6785
rect 24733 6721 24734 6785
rect 24668 6705 24734 6721
rect 24148 6648 24292 6649
rect 24668 6641 24669 6705
rect 24733 6641 24734 6705
rect 24668 6625 24734 6641
rect 24668 6561 24669 6625
rect 24733 6561 24734 6625
rect 24668 6545 24734 6561
rect 24668 6481 24669 6545
rect 24733 6481 24734 6545
rect 23599 6466 23771 6476
rect 23599 6320 23609 6466
rect 23759 6320 23771 6466
rect 23599 6310 23771 6320
rect 24668 6465 24734 6481
rect 24668 6401 24669 6465
rect 24733 6401 24734 6465
rect 24668 6385 24734 6401
rect 24668 6321 24669 6385
rect 24733 6321 24734 6385
rect 24183 6199 24275 6200
rect 24069 6184 24442 6199
rect 11251 6132 11423 6142
rect 10945 6120 11117 6130
rect 10945 5974 10955 6120
rect 11105 5974 11117 6120
rect 11251 5986 11261 6132
rect 11411 5986 11423 6132
rect 24069 6120 24076 6184
rect 24140 6120 24196 6184
rect 24260 6120 24339 6184
rect 24403 6120 24442 6184
rect 24069 6103 24442 6120
rect 24668 6167 24734 6321
rect 24794 6167 24854 7199
rect 24914 6229 24974 7259
rect 25034 6167 25094 7199
rect 25154 6229 25214 7259
rect 25274 7105 25340 7195
rect 25274 7041 25275 7105
rect 25339 7041 25340 7105
rect 25274 7025 25340 7041
rect 25274 6961 25275 7025
rect 25339 6961 25340 7025
rect 25274 6945 25340 6961
rect 25274 6881 25275 6945
rect 25339 6881 25340 6945
rect 25274 6865 25340 6881
rect 25274 6801 25275 6865
rect 25339 6801 25340 6865
rect 25274 6785 25340 6801
rect 25274 6721 25275 6785
rect 25339 6721 25340 6785
rect 25274 6705 25340 6721
rect 25274 6641 25275 6705
rect 25339 6641 25340 6705
rect 25274 6625 25340 6641
rect 25274 6561 25275 6625
rect 25339 6561 25340 6625
rect 25274 6545 25340 6561
rect 25274 6481 25275 6545
rect 25339 6481 25340 6545
rect 25274 6465 25340 6481
rect 25274 6401 25275 6465
rect 25339 6401 25340 6465
rect 25274 6385 25340 6401
rect 25274 6321 25275 6385
rect 25339 6321 25340 6385
rect 25274 6167 25340 6321
rect 24668 6165 25340 6167
rect 24668 6101 24772 6165
rect 24836 6101 24852 6165
rect 24916 6101 24932 6165
rect 24996 6101 25012 6165
rect 25076 6101 25092 6165
rect 25156 6142 25172 6165
rect 25156 6101 25161 6142
rect 25236 6101 25340 6165
rect 25400 7108 25466 7198
rect 25400 7044 25401 7108
rect 25465 7044 25466 7108
rect 25400 7028 25466 7044
rect 25400 6964 25401 7028
rect 25465 6964 25466 7028
rect 25400 6948 25466 6964
rect 25400 6884 25401 6948
rect 25465 6884 25466 6948
rect 25400 6868 25466 6884
rect 25400 6804 25401 6868
rect 25465 6804 25466 6868
rect 25400 6788 25466 6804
rect 25400 6724 25401 6788
rect 25465 6724 25466 6788
rect 25400 6708 25466 6724
rect 25400 6644 25401 6708
rect 25465 6644 25466 6708
rect 25400 6628 25466 6644
rect 25400 6564 25401 6628
rect 25465 6564 25466 6628
rect 25400 6548 25466 6564
rect 25400 6484 25401 6548
rect 25465 6484 25466 6548
rect 25400 6468 25466 6484
rect 25400 6404 25401 6468
rect 25465 6404 25466 6468
rect 25400 6388 25466 6404
rect 25400 6324 25401 6388
rect 25465 6324 25466 6388
rect 25400 6170 25466 6324
rect 25526 6170 25586 7202
rect 25646 6232 25706 7262
rect 25766 6170 25826 7202
rect 25886 6232 25946 7262
rect 26006 7108 26072 7198
rect 26006 7044 26007 7108
rect 26071 7044 26072 7108
rect 26006 7028 26072 7044
rect 26006 6964 26007 7028
rect 26071 6964 26072 7028
rect 26006 6948 26072 6964
rect 26006 6884 26007 6948
rect 26071 6884 26072 6948
rect 26006 6868 26072 6884
rect 26006 6804 26007 6868
rect 26071 6804 26072 6868
rect 26006 6788 26072 6804
rect 26006 6724 26007 6788
rect 26071 6724 26072 6788
rect 26006 6708 26072 6724
rect 26006 6644 26007 6708
rect 26071 6644 26072 6708
rect 26006 6628 26072 6644
rect 26006 6564 26007 6628
rect 26071 6564 26072 6628
rect 26006 6548 26072 6564
rect 26006 6484 26007 6548
rect 26071 6484 26072 6548
rect 26006 6468 26072 6484
rect 26006 6404 26007 6468
rect 26071 6404 26072 6468
rect 26006 6388 26072 6404
rect 26006 6324 26007 6388
rect 26071 6324 26072 6388
rect 26006 6170 26072 6324
rect 26132 6232 26192 7262
rect 26252 6170 26312 7202
rect 26372 6232 26432 7262
rect 26492 6170 26552 7202
rect 26612 7108 26678 7198
rect 26612 7044 26613 7108
rect 26677 7044 26678 7108
rect 26612 7028 26678 7044
rect 26612 6964 26613 7028
rect 26677 6964 26678 7028
rect 26612 6948 26678 6964
rect 26612 6884 26613 6948
rect 26677 6884 26678 6948
rect 26612 6868 26678 6884
rect 26612 6804 26613 6868
rect 26677 6804 26678 6868
rect 26612 6788 26678 6804
rect 26612 6724 26613 6788
rect 26677 6724 26678 6788
rect 26612 6708 26678 6724
rect 26612 6644 26613 6708
rect 26677 6644 26678 6708
rect 26612 6628 26678 6644
rect 26612 6564 26613 6628
rect 26677 6564 26678 6628
rect 26612 6548 26678 6564
rect 26612 6484 26613 6548
rect 26677 6484 26678 6548
rect 26612 6468 26678 6484
rect 26612 6404 26613 6468
rect 26677 6404 26678 6468
rect 26612 6388 26678 6404
rect 26612 6324 26613 6388
rect 26677 6324 26678 6388
rect 26612 6170 26678 6324
rect 26738 6170 26798 7202
rect 26858 6232 26918 7262
rect 26978 6170 27038 7202
rect 27098 6232 27158 7262
rect 27218 7108 27284 7198
rect 27218 7044 27219 7108
rect 27283 7044 27284 7108
rect 27218 7028 27284 7044
rect 27218 6964 27219 7028
rect 27283 6964 27284 7028
rect 27218 6948 27284 6964
rect 27218 6884 27219 6948
rect 27283 6884 27284 6948
rect 27218 6868 27284 6884
rect 27218 6804 27219 6868
rect 27283 6804 27284 6868
rect 27218 6788 27284 6804
rect 27218 6724 27219 6788
rect 27283 6724 27284 6788
rect 27218 6708 27284 6724
rect 27218 6644 27219 6708
rect 27283 6644 27284 6708
rect 27218 6628 27284 6644
rect 27218 6564 27219 6628
rect 27283 6564 27284 6628
rect 27218 6548 27284 6564
rect 27218 6484 27219 6548
rect 27283 6484 27284 6548
rect 27218 6468 27284 6484
rect 27218 6404 27219 6468
rect 27283 6404 27284 6468
rect 27218 6388 27284 6404
rect 27218 6324 27219 6388
rect 27283 6324 27284 6388
rect 27218 6170 27284 6324
rect 27344 6232 27404 7262
rect 27464 6170 27524 7202
rect 27584 6232 27644 7262
rect 27704 6170 27764 7202
rect 27824 7108 27890 7198
rect 27824 7044 27825 7108
rect 27889 7044 27890 7108
rect 27824 7028 27890 7044
rect 27824 6964 27825 7028
rect 27889 6964 27890 7028
rect 27824 6948 27890 6964
rect 27824 6884 27825 6948
rect 27889 6884 27890 6948
rect 27824 6868 27890 6884
rect 27824 6804 27825 6868
rect 27889 6804 27890 6868
rect 27824 6788 27890 6804
rect 27824 6724 27825 6788
rect 27889 6724 27890 6788
rect 27824 6708 27890 6724
rect 27824 6644 27825 6708
rect 27889 6644 27890 6708
rect 27824 6628 27890 6644
rect 27824 6564 27825 6628
rect 27889 6564 27890 6628
rect 27824 6548 27890 6564
rect 27824 6484 27825 6548
rect 27889 6484 27890 6548
rect 27824 6468 27890 6484
rect 27824 6404 27825 6468
rect 27889 6404 27890 6468
rect 27824 6388 27890 6404
rect 27824 6324 27825 6388
rect 27889 6324 27890 6388
rect 27824 6170 27890 6324
rect 27950 6170 28010 7202
rect 28070 6232 28130 7262
rect 28190 6170 28250 7202
rect 28310 6232 28370 7262
rect 28430 7108 28496 7198
rect 28430 7044 28431 7108
rect 28495 7044 28496 7108
rect 28430 7028 28496 7044
rect 28430 6964 28431 7028
rect 28495 6964 28496 7028
rect 28430 6948 28496 6964
rect 28430 6884 28431 6948
rect 28495 6884 28496 6948
rect 28430 6868 28496 6884
rect 28430 6804 28431 6868
rect 28495 6804 28496 6868
rect 28430 6788 28496 6804
rect 28430 6724 28431 6788
rect 28495 6724 28496 6788
rect 28430 6708 28496 6724
rect 28430 6644 28431 6708
rect 28495 6644 28496 6708
rect 28430 6628 28496 6644
rect 28430 6564 28431 6628
rect 28495 6564 28496 6628
rect 28430 6548 28496 6564
rect 28430 6484 28431 6548
rect 28495 6484 28496 6548
rect 28430 6468 28496 6484
rect 28430 6404 28431 6468
rect 28495 6404 28496 6468
rect 28430 6388 28496 6404
rect 28430 6324 28431 6388
rect 28495 6324 28496 6388
rect 28430 6170 28496 6324
rect 28556 6232 28616 7262
rect 28676 6170 28736 7202
rect 28796 6232 28856 7262
rect 28916 6170 28976 7202
rect 29036 7108 29102 7198
rect 29036 7044 29037 7108
rect 29101 7044 29102 7108
rect 29036 7028 29102 7044
rect 29036 6964 29037 7028
rect 29101 6964 29102 7028
rect 29036 6948 29102 6964
rect 29036 6884 29037 6948
rect 29101 6884 29102 6948
rect 29036 6868 29102 6884
rect 29036 6804 29037 6868
rect 29101 6804 29102 6868
rect 29036 6788 29102 6804
rect 29036 6724 29037 6788
rect 29101 6724 29102 6788
rect 29036 6708 29102 6724
rect 29036 6644 29037 6708
rect 29101 6644 29102 6708
rect 29036 6628 29102 6644
rect 29036 6564 29037 6628
rect 29101 6564 29102 6628
rect 29036 6548 29102 6564
rect 29036 6484 29037 6548
rect 29101 6484 29102 6548
rect 29036 6468 29102 6484
rect 29036 6404 29037 6468
rect 29101 6404 29102 6468
rect 29036 6388 29102 6404
rect 29036 6324 29037 6388
rect 29101 6324 29102 6388
rect 29036 6170 29102 6324
rect 29162 6170 29222 7202
rect 29282 6232 29342 7262
rect 29402 6170 29462 7202
rect 29522 6232 29582 7262
rect 29642 7108 29708 7198
rect 29642 7044 29643 7108
rect 29707 7044 29708 7108
rect 29642 7028 29708 7044
rect 29642 6964 29643 7028
rect 29707 6964 29708 7028
rect 29642 6948 29708 6964
rect 29642 6884 29643 6948
rect 29707 6884 29708 6948
rect 29642 6868 29708 6884
rect 29642 6804 29643 6868
rect 29707 6804 29708 6868
rect 29642 6788 29708 6804
rect 29642 6724 29643 6788
rect 29707 6724 29708 6788
rect 29642 6708 29708 6724
rect 29642 6644 29643 6708
rect 29707 6644 29708 6708
rect 29642 6628 29708 6644
rect 29642 6564 29643 6628
rect 29707 6564 29708 6628
rect 29642 6548 29708 6564
rect 29642 6484 29643 6548
rect 29707 6484 29708 6548
rect 29642 6468 29708 6484
rect 29642 6404 29643 6468
rect 29707 6404 29708 6468
rect 29642 6388 29708 6404
rect 29642 6324 29643 6388
rect 29707 6324 29708 6388
rect 29642 6170 29708 6324
rect 29768 6232 29828 7262
rect 29888 6170 29948 7202
rect 30008 6232 30068 7262
rect 30453 7209 30484 7273
rect 30548 7209 30579 7273
rect 30128 6170 30188 7202
rect 30453 7199 30579 7209
rect 30248 7108 30314 7198
rect 30248 7044 30249 7108
rect 30313 7044 30314 7108
rect 30458 7129 30584 7139
rect 30458 7065 30489 7129
rect 30553 7065 30584 7129
rect 30458 7055 30584 7065
rect 30248 7028 30314 7044
rect 30248 6964 30249 7028
rect 30313 6964 30314 7028
rect 30248 6948 30314 6964
rect 30248 6884 30249 6948
rect 30313 6884 30314 6948
rect 30459 6977 30585 6987
rect 30459 6913 30490 6977
rect 30554 6913 30585 6977
rect 30459 6903 30585 6913
rect 30248 6868 30314 6884
rect 30248 6804 30249 6868
rect 30313 6804 30314 6868
rect 30248 6788 30314 6804
rect 30248 6724 30249 6788
rect 30313 6724 30314 6788
rect 30459 6807 30585 6817
rect 30459 6743 30490 6807
rect 30554 6743 30585 6807
rect 30459 6733 30585 6743
rect 30248 6708 30314 6724
rect 30248 6644 30249 6708
rect 30313 6644 30314 6708
rect 30248 6628 30314 6644
rect 30248 6564 30249 6628
rect 30313 6564 30314 6628
rect 30458 6650 30584 6660
rect 30458 6586 30489 6650
rect 30553 6586 30584 6650
rect 30458 6576 30584 6586
rect 30248 6548 30314 6564
rect 30248 6484 30249 6548
rect 30313 6484 30314 6548
rect 30248 6468 30314 6484
rect 30248 6404 30249 6468
rect 30313 6404 30314 6468
rect 30248 6388 30314 6404
rect 30248 6324 30249 6388
rect 30313 6324 30314 6388
rect 30376 6408 30502 6418
rect 30376 6344 30407 6408
rect 30471 6344 30502 6408
rect 30376 6334 30502 6344
rect 30753 6416 30879 6426
rect 30753 6352 30784 6416
rect 30848 6352 30879 6416
rect 30753 6342 30879 6352
rect 30953 6416 31079 6426
rect 30953 6352 30984 6416
rect 31048 6352 31079 6416
rect 30953 6342 31079 6352
rect 30248 6170 30314 6324
rect 25400 6168 30314 6170
rect 25400 6104 25504 6168
rect 25568 6104 25584 6168
rect 25648 6104 25664 6168
rect 25728 6104 25744 6168
rect 25808 6104 25824 6168
rect 25888 6145 25904 6168
rect 25888 6104 25893 6145
rect 25968 6104 26110 6168
rect 26174 6145 26190 6168
rect 26185 6104 26190 6145
rect 26254 6104 26270 6168
rect 26334 6104 26350 6168
rect 26414 6104 26430 6168
rect 26494 6104 26510 6168
rect 26574 6104 26716 6168
rect 26780 6104 26796 6168
rect 26860 6104 26876 6168
rect 26940 6104 26956 6168
rect 27020 6104 27036 6168
rect 27100 6145 27116 6168
rect 27100 6104 27105 6145
rect 27180 6104 27322 6168
rect 27386 6145 27402 6168
rect 27397 6104 27402 6145
rect 27466 6104 27482 6168
rect 27546 6104 27562 6168
rect 27626 6104 27642 6168
rect 27706 6104 27722 6168
rect 27786 6104 27928 6168
rect 27992 6104 28008 6168
rect 28072 6104 28088 6168
rect 28152 6104 28168 6168
rect 28232 6104 28248 6168
rect 28312 6145 28328 6168
rect 28312 6104 28317 6145
rect 28392 6104 28534 6168
rect 28598 6145 28614 6168
rect 28609 6104 28614 6145
rect 28678 6104 28694 6168
rect 28758 6104 28774 6168
rect 28838 6104 28854 6168
rect 28918 6104 28934 6168
rect 28998 6104 29140 6168
rect 29204 6104 29220 6168
rect 29284 6104 29300 6168
rect 29364 6104 29380 6168
rect 29444 6104 29460 6168
rect 29524 6145 29540 6168
rect 29524 6104 29529 6145
rect 29604 6104 29746 6168
rect 29810 6145 29826 6168
rect 29821 6104 29826 6145
rect 29890 6104 29906 6168
rect 29970 6104 29986 6168
rect 30050 6104 30066 6168
rect 30130 6104 30146 6168
rect 30210 6104 30314 6168
rect 25400 6102 25893 6104
rect 24668 6099 25161 6101
rect 25151 6078 25161 6099
rect 25225 6099 25340 6101
rect 25225 6078 25234 6099
rect 25151 6073 25234 6078
rect 25883 6081 25893 6102
rect 25957 6102 26121 6104
rect 25957 6081 25966 6102
rect 25883 6076 25966 6081
rect 26112 6081 26121 6102
rect 26185 6102 27105 6104
rect 26185 6081 26195 6102
rect 26112 6076 26195 6081
rect 27095 6081 27105 6102
rect 27169 6102 27333 6104
rect 27169 6081 27178 6102
rect 27095 6076 27178 6081
rect 27324 6081 27333 6102
rect 27397 6102 28317 6104
rect 27397 6081 27407 6102
rect 27324 6076 27407 6081
rect 28307 6081 28317 6102
rect 28381 6102 28545 6104
rect 28381 6081 28390 6102
rect 28307 6076 28390 6081
rect 28536 6081 28545 6102
rect 28609 6102 29529 6104
rect 28609 6081 28619 6102
rect 28536 6076 28619 6081
rect 29519 6081 29529 6102
rect 29593 6102 29757 6104
rect 29593 6081 29602 6102
rect 29519 6076 29602 6081
rect 29748 6081 29757 6102
rect 29821 6102 30314 6104
rect 30464 6147 30590 6157
rect 29821 6081 29831 6102
rect 29748 6076 29831 6081
rect 30464 6083 30495 6147
rect 30559 6083 30590 6147
rect 30464 6073 30590 6083
rect 11251 5976 11423 5986
rect 23599 6040 23771 6050
rect 10945 5964 11117 5974
rect 23599 5894 23609 6040
rect 23759 5894 23771 6040
rect 25508 5943 25590 5949
rect 25508 5922 25517 5943
rect 23599 5884 23771 5894
rect 25019 5920 25517 5922
rect 25581 5922 25590 5943
rect 26240 5943 26322 5949
rect 26240 5922 26249 5943
rect 25581 5920 25691 5922
rect 25019 5856 25123 5920
rect 25187 5856 25203 5920
rect 25267 5856 25283 5920
rect 25347 5856 25363 5920
rect 25427 5856 25443 5920
rect 25507 5879 25517 5920
rect 25507 5856 25523 5879
rect 25587 5856 25691 5920
rect 25019 5854 25691 5856
rect 23599 5814 23771 5824
rect 23599 5668 23609 5814
rect 23759 5668 23771 5814
rect 23599 5658 23771 5668
rect 25019 5700 25085 5854
rect 25019 5636 25020 5700
rect 25084 5636 25085 5700
rect 25019 5620 25085 5636
rect 25019 5556 25020 5620
rect 25084 5556 25085 5620
rect 25019 5540 25085 5556
rect 10777 5492 10949 5502
rect 10777 5346 10787 5492
rect 10937 5346 10949 5492
rect 10777 5336 10949 5346
rect 25019 5476 25020 5540
rect 25084 5476 25085 5540
rect 25019 5460 25085 5476
rect 25019 5396 25020 5460
rect 25084 5396 25085 5460
rect 25019 5380 25085 5396
rect 25019 5316 25020 5380
rect 25084 5316 25085 5380
rect 25019 5300 25085 5316
rect 25019 5236 25020 5300
rect 25084 5236 25085 5300
rect 25019 5220 25085 5236
rect 25019 5156 25020 5220
rect 25084 5156 25085 5220
rect 25019 5140 25085 5156
rect 23615 5080 23787 5090
rect 23615 4934 23625 5080
rect 23775 4934 23787 5080
rect 23615 4924 23787 4934
rect 25019 5076 25020 5140
rect 25084 5076 25085 5140
rect 25019 5060 25085 5076
rect 25019 4996 25020 5060
rect 25084 4996 25085 5060
rect 25019 4980 25085 4996
rect 25019 4916 25020 4980
rect 25084 4916 25085 4980
rect 25019 4826 25085 4916
rect 25145 4822 25205 5854
rect 24631 4757 24756 4767
rect 25265 4762 25325 5792
rect 25385 4822 25445 5854
rect 25505 4762 25565 5792
rect 25625 5700 25691 5854
rect 25625 5636 25626 5700
rect 25690 5636 25691 5700
rect 25625 5620 25691 5636
rect 25625 5556 25626 5620
rect 25690 5556 25691 5620
rect 25625 5540 25691 5556
rect 25625 5476 25626 5540
rect 25690 5476 25691 5540
rect 25625 5460 25691 5476
rect 25625 5396 25626 5460
rect 25690 5396 25691 5460
rect 25625 5380 25691 5396
rect 25625 5316 25626 5380
rect 25690 5316 25691 5380
rect 25625 5300 25691 5316
rect 25625 5236 25626 5300
rect 25690 5236 25691 5300
rect 25625 5220 25691 5236
rect 25625 5156 25626 5220
rect 25690 5156 25691 5220
rect 25625 5140 25691 5156
rect 25625 5076 25626 5140
rect 25690 5076 25691 5140
rect 25625 5060 25691 5076
rect 25625 4996 25626 5060
rect 25690 4996 25691 5060
rect 25625 4980 25691 4996
rect 25625 4916 25626 4980
rect 25690 4916 25691 4980
rect 25625 4826 25691 4916
rect 25751 5920 26249 5922
rect 26313 5922 26322 5943
rect 26458 5943 26540 5949
rect 26458 5922 26467 5943
rect 26313 5920 26467 5922
rect 26531 5922 26540 5943
rect 27452 5943 27534 5949
rect 27452 5922 27461 5943
rect 26531 5920 27461 5922
rect 27525 5922 27534 5943
rect 27670 5943 27752 5949
rect 27670 5922 27679 5943
rect 27525 5920 27679 5922
rect 27743 5922 27752 5943
rect 28790 5943 28872 5949
rect 28790 5922 28799 5943
rect 27743 5920 28241 5922
rect 25751 5856 25855 5920
rect 25919 5856 25935 5920
rect 25999 5856 26015 5920
rect 26079 5856 26095 5920
rect 26159 5856 26175 5920
rect 26239 5879 26249 5920
rect 26239 5856 26255 5879
rect 26319 5856 26461 5920
rect 26531 5879 26541 5920
rect 26525 5856 26541 5879
rect 26605 5856 26621 5920
rect 26685 5856 26701 5920
rect 26765 5856 26781 5920
rect 26845 5856 26861 5920
rect 26925 5856 27067 5920
rect 27131 5856 27147 5920
rect 27211 5856 27227 5920
rect 27291 5856 27307 5920
rect 27371 5856 27387 5920
rect 27451 5879 27461 5920
rect 27451 5856 27467 5879
rect 27531 5856 27673 5920
rect 27743 5879 27753 5920
rect 27737 5856 27753 5879
rect 27817 5856 27833 5920
rect 27897 5856 27913 5920
rect 27977 5856 27993 5920
rect 28057 5856 28073 5920
rect 28137 5856 28241 5920
rect 25751 5854 28241 5856
rect 25751 5700 25817 5854
rect 25751 5636 25752 5700
rect 25816 5636 25817 5700
rect 25751 5620 25817 5636
rect 25751 5556 25752 5620
rect 25816 5556 25817 5620
rect 25751 5540 25817 5556
rect 25751 5476 25752 5540
rect 25816 5476 25817 5540
rect 25751 5460 25817 5476
rect 25751 5396 25752 5460
rect 25816 5396 25817 5460
rect 25751 5380 25817 5396
rect 25751 5316 25752 5380
rect 25816 5316 25817 5380
rect 25751 5300 25817 5316
rect 25751 5236 25752 5300
rect 25816 5236 25817 5300
rect 25751 5220 25817 5236
rect 25751 5156 25752 5220
rect 25816 5156 25817 5220
rect 25751 5140 25817 5156
rect 25751 5076 25752 5140
rect 25816 5076 25817 5140
rect 25751 5060 25817 5076
rect 25751 4996 25752 5060
rect 25816 4996 25817 5060
rect 25751 4980 25817 4996
rect 25751 4916 25752 4980
rect 25816 4916 25817 4980
rect 25751 4826 25817 4916
rect 25877 4822 25937 5854
rect 25997 4762 26057 5792
rect 26117 4822 26177 5854
rect 26237 4762 26297 5792
rect 26357 5700 26423 5854
rect 26357 5636 26358 5700
rect 26422 5636 26423 5700
rect 26357 5620 26423 5636
rect 26357 5556 26358 5620
rect 26422 5556 26423 5620
rect 26357 5540 26423 5556
rect 26357 5476 26358 5540
rect 26422 5476 26423 5540
rect 26357 5460 26423 5476
rect 26357 5396 26358 5460
rect 26422 5396 26423 5460
rect 26357 5380 26423 5396
rect 26357 5316 26358 5380
rect 26422 5316 26423 5380
rect 26357 5300 26423 5316
rect 26357 5236 26358 5300
rect 26422 5236 26423 5300
rect 26357 5220 26423 5236
rect 26357 5156 26358 5220
rect 26422 5156 26423 5220
rect 26357 5140 26423 5156
rect 26357 5076 26358 5140
rect 26422 5076 26423 5140
rect 26357 5060 26423 5076
rect 26357 4996 26358 5060
rect 26422 4996 26423 5060
rect 26357 4980 26423 4996
rect 26357 4916 26358 4980
rect 26422 4916 26423 4980
rect 26357 4826 26423 4916
rect 26483 4762 26543 5792
rect 26603 4822 26663 5854
rect 26723 4762 26783 5792
rect 26843 4822 26903 5854
rect 26963 5700 27029 5854
rect 26963 5636 26964 5700
rect 27028 5636 27029 5700
rect 26963 5620 27029 5636
rect 26963 5556 26964 5620
rect 27028 5556 27029 5620
rect 26963 5540 27029 5556
rect 26963 5476 26964 5540
rect 27028 5476 27029 5540
rect 26963 5460 27029 5476
rect 26963 5396 26964 5460
rect 27028 5396 27029 5460
rect 26963 5380 27029 5396
rect 26963 5316 26964 5380
rect 27028 5316 27029 5380
rect 26963 5300 27029 5316
rect 26963 5236 26964 5300
rect 27028 5236 27029 5300
rect 26963 5220 27029 5236
rect 26963 5156 26964 5220
rect 27028 5156 27029 5220
rect 26963 5140 27029 5156
rect 26963 5076 26964 5140
rect 27028 5076 27029 5140
rect 26963 5060 27029 5076
rect 26963 4996 26964 5060
rect 27028 4996 27029 5060
rect 26963 4980 27029 4996
rect 26963 4916 26964 4980
rect 27028 4916 27029 4980
rect 26963 4826 27029 4916
rect 27089 4822 27149 5854
rect 27209 4762 27269 5792
rect 27329 4822 27389 5854
rect 27449 4762 27509 5792
rect 27569 5700 27635 5854
rect 27569 5636 27570 5700
rect 27634 5636 27635 5700
rect 27569 5620 27635 5636
rect 27569 5556 27570 5620
rect 27634 5556 27635 5620
rect 27569 5540 27635 5556
rect 27569 5476 27570 5540
rect 27634 5476 27635 5540
rect 27569 5460 27635 5476
rect 27569 5396 27570 5460
rect 27634 5396 27635 5460
rect 27569 5380 27635 5396
rect 27569 5316 27570 5380
rect 27634 5316 27635 5380
rect 27569 5300 27635 5316
rect 27569 5236 27570 5300
rect 27634 5236 27635 5300
rect 27569 5220 27635 5236
rect 27569 5156 27570 5220
rect 27634 5156 27635 5220
rect 27569 5140 27635 5156
rect 27569 5076 27570 5140
rect 27634 5076 27635 5140
rect 27569 5060 27635 5076
rect 27569 4996 27570 5060
rect 27634 4996 27635 5060
rect 27569 4980 27635 4996
rect 27569 4916 27570 4980
rect 27634 4916 27635 4980
rect 27569 4826 27635 4916
rect 27695 4762 27755 5792
rect 27815 4822 27875 5854
rect 27935 4762 27995 5792
rect 28055 4822 28115 5854
rect 28175 5700 28241 5854
rect 28175 5636 28176 5700
rect 28240 5636 28241 5700
rect 28175 5620 28241 5636
rect 28175 5556 28176 5620
rect 28240 5556 28241 5620
rect 28175 5540 28241 5556
rect 28175 5476 28176 5540
rect 28240 5476 28241 5540
rect 28175 5460 28241 5476
rect 28175 5396 28176 5460
rect 28240 5396 28241 5460
rect 28175 5380 28241 5396
rect 28175 5316 28176 5380
rect 28240 5316 28241 5380
rect 28175 5300 28241 5316
rect 28175 5236 28176 5300
rect 28240 5236 28241 5300
rect 28175 5220 28241 5236
rect 28175 5156 28176 5220
rect 28240 5156 28241 5220
rect 28175 5140 28241 5156
rect 28175 5076 28176 5140
rect 28240 5076 28241 5140
rect 28175 5060 28241 5076
rect 28175 4996 28176 5060
rect 28240 4996 28241 5060
rect 28175 4980 28241 4996
rect 28175 4916 28176 4980
rect 28240 4916 28241 4980
rect 28175 4826 28241 4916
rect 28301 5920 28799 5922
rect 28863 5922 28872 5943
rect 29008 5943 29090 5949
rect 29008 5922 29017 5943
rect 28863 5920 29017 5922
rect 29081 5922 29090 5943
rect 29742 5943 29824 5949
rect 29742 5922 29751 5943
rect 29081 5920 29579 5922
rect 28301 5856 28405 5920
rect 28469 5856 28485 5920
rect 28549 5856 28565 5920
rect 28629 5856 28645 5920
rect 28709 5856 28725 5920
rect 28789 5879 28799 5920
rect 28789 5856 28805 5879
rect 28869 5856 29011 5920
rect 29081 5879 29091 5920
rect 29075 5856 29091 5879
rect 29155 5856 29171 5920
rect 29235 5856 29251 5920
rect 29315 5856 29331 5920
rect 29395 5856 29411 5920
rect 29475 5856 29579 5920
rect 28301 5854 29579 5856
rect 28301 5700 28367 5854
rect 28301 5636 28302 5700
rect 28366 5636 28367 5700
rect 28301 5620 28367 5636
rect 28301 5556 28302 5620
rect 28366 5556 28367 5620
rect 28301 5540 28367 5556
rect 28301 5476 28302 5540
rect 28366 5476 28367 5540
rect 28301 5460 28367 5476
rect 28301 5396 28302 5460
rect 28366 5396 28367 5460
rect 28301 5380 28367 5396
rect 28301 5316 28302 5380
rect 28366 5316 28367 5380
rect 28301 5300 28367 5316
rect 28301 5236 28302 5300
rect 28366 5236 28367 5300
rect 28301 5220 28367 5236
rect 28301 5156 28302 5220
rect 28366 5156 28367 5220
rect 28301 5140 28367 5156
rect 28301 5076 28302 5140
rect 28366 5076 28367 5140
rect 28301 5060 28367 5076
rect 28301 4996 28302 5060
rect 28366 4996 28367 5060
rect 28301 4980 28367 4996
rect 28301 4916 28302 4980
rect 28366 4916 28367 4980
rect 28301 4826 28367 4916
rect 28427 4822 28487 5854
rect 28547 4762 28607 5792
rect 28667 4822 28727 5854
rect 28787 4762 28847 5792
rect 28907 5700 28973 5854
rect 28907 5636 28908 5700
rect 28972 5636 28973 5700
rect 28907 5620 28973 5636
rect 28907 5556 28908 5620
rect 28972 5556 28973 5620
rect 28907 5540 28973 5556
rect 28907 5476 28908 5540
rect 28972 5476 28973 5540
rect 28907 5460 28973 5476
rect 28907 5396 28908 5460
rect 28972 5396 28973 5460
rect 28907 5380 28973 5396
rect 28907 5316 28908 5380
rect 28972 5316 28973 5380
rect 28907 5300 28973 5316
rect 28907 5236 28908 5300
rect 28972 5236 28973 5300
rect 28907 5220 28973 5236
rect 28907 5156 28908 5220
rect 28972 5156 28973 5220
rect 28907 5140 28973 5156
rect 28907 5076 28908 5140
rect 28972 5076 28973 5140
rect 28907 5060 28973 5076
rect 28907 4996 28908 5060
rect 28972 4996 28973 5060
rect 28907 4980 28973 4996
rect 28907 4916 28908 4980
rect 28972 4916 28973 4980
rect 28907 4826 28973 4916
rect 29033 4762 29093 5792
rect 29153 4822 29213 5854
rect 29273 4762 29333 5792
rect 29393 4822 29453 5854
rect 29513 5700 29579 5854
rect 29513 5636 29514 5700
rect 29578 5636 29579 5700
rect 29513 5620 29579 5636
rect 29513 5556 29514 5620
rect 29578 5556 29579 5620
rect 29513 5540 29579 5556
rect 29513 5476 29514 5540
rect 29578 5476 29579 5540
rect 29513 5460 29579 5476
rect 29513 5396 29514 5460
rect 29578 5396 29579 5460
rect 29513 5380 29579 5396
rect 29513 5316 29514 5380
rect 29578 5316 29579 5380
rect 29513 5300 29579 5316
rect 29513 5236 29514 5300
rect 29578 5236 29579 5300
rect 29513 5220 29579 5236
rect 29513 5156 29514 5220
rect 29578 5156 29579 5220
rect 29513 5140 29579 5156
rect 29513 5076 29514 5140
rect 29578 5076 29579 5140
rect 29513 5060 29579 5076
rect 29513 4996 29514 5060
rect 29578 4996 29579 5060
rect 29513 4980 29579 4996
rect 29513 4916 29514 4980
rect 29578 4916 29579 4980
rect 29513 4826 29579 4916
rect 29641 5920 29751 5922
rect 29815 5922 29824 5943
rect 30464 5944 30590 5954
rect 29815 5920 30313 5922
rect 29641 5856 29745 5920
rect 29815 5879 29825 5920
rect 29809 5856 29825 5879
rect 29889 5856 29905 5920
rect 29969 5856 29985 5920
rect 30049 5856 30065 5920
rect 30129 5856 30145 5920
rect 30209 5856 30313 5920
rect 30464 5880 30495 5944
rect 30559 5880 30590 5944
rect 30464 5870 30590 5880
rect 30490 5869 30564 5870
rect 29641 5854 30313 5856
rect 29641 5700 29707 5854
rect 29641 5636 29642 5700
rect 29706 5636 29707 5700
rect 29641 5620 29707 5636
rect 29641 5556 29642 5620
rect 29706 5556 29707 5620
rect 29641 5540 29707 5556
rect 29641 5476 29642 5540
rect 29706 5476 29707 5540
rect 29641 5460 29707 5476
rect 29641 5396 29642 5460
rect 29706 5396 29707 5460
rect 29641 5380 29707 5396
rect 29641 5316 29642 5380
rect 29706 5316 29707 5380
rect 29641 5300 29707 5316
rect 29641 5236 29642 5300
rect 29706 5236 29707 5300
rect 29641 5220 29707 5236
rect 29641 5156 29642 5220
rect 29706 5156 29707 5220
rect 29641 5140 29707 5156
rect 29641 5076 29642 5140
rect 29706 5076 29707 5140
rect 29641 5060 29707 5076
rect 29641 4996 29642 5060
rect 29706 4996 29707 5060
rect 29641 4980 29707 4996
rect 29641 4916 29642 4980
rect 29706 4916 29707 4980
rect 29641 4826 29707 4916
rect 29767 4762 29827 5792
rect 29887 4822 29947 5854
rect 30007 4762 30067 5792
rect 30127 4822 30187 5854
rect 30247 5700 30313 5854
rect 30565 5774 30690 5784
rect 30565 5710 30595 5774
rect 30659 5710 30690 5774
rect 30565 5700 30690 5710
rect 30247 5636 30248 5700
rect 30312 5636 30313 5700
rect 30247 5620 30313 5636
rect 30247 5556 30248 5620
rect 30312 5556 30313 5620
rect 30374 5682 30499 5692
rect 30374 5618 30404 5682
rect 30468 5618 30499 5682
rect 30374 5608 30499 5618
rect 30247 5540 30313 5556
rect 30247 5476 30248 5540
rect 30312 5476 30313 5540
rect 30247 5460 30313 5476
rect 30247 5396 30248 5460
rect 30312 5396 30313 5460
rect 30247 5380 30313 5396
rect 30247 5316 30248 5380
rect 30312 5316 30313 5380
rect 30247 5300 30313 5316
rect 30247 5236 30248 5300
rect 30312 5236 30313 5300
rect 30247 5220 30313 5236
rect 30247 5156 30248 5220
rect 30312 5156 30313 5220
rect 30247 5140 30313 5156
rect 30247 5076 30248 5140
rect 30312 5076 30313 5140
rect 30247 5060 30313 5076
rect 30247 4996 30248 5060
rect 30312 4996 30313 5060
rect 30247 4980 30313 4996
rect 30247 4916 30248 4980
rect 30312 4916 30313 4980
rect 30247 4826 30313 4916
rect 24631 4693 24661 4757
rect 24725 4693 24756 4757
rect 25019 4760 25691 4762
rect 25019 4696 25203 4760
rect 25267 4696 25283 4760
rect 25347 4696 25363 4760
rect 25427 4696 25443 4760
rect 25507 4696 25691 4760
rect 25019 4694 25691 4696
rect 25751 4760 28241 4762
rect 25751 4696 25935 4760
rect 25999 4696 26015 4760
rect 26079 4696 26095 4760
rect 26159 4696 26175 4760
rect 26239 4696 26541 4760
rect 26605 4696 26621 4760
rect 26685 4696 26701 4760
rect 26765 4696 26781 4760
rect 26845 4696 27147 4760
rect 27211 4696 27227 4760
rect 27291 4696 27307 4760
rect 27371 4696 27387 4760
rect 27451 4696 27753 4760
rect 27817 4696 27833 4760
rect 27897 4696 27913 4760
rect 27977 4696 27993 4760
rect 28057 4696 28241 4760
rect 25751 4694 28241 4696
rect 28301 4760 29579 4762
rect 28301 4696 28485 4760
rect 28549 4696 28565 4760
rect 28629 4696 28645 4760
rect 28709 4696 28725 4760
rect 28789 4696 29091 4760
rect 29155 4696 29171 4760
rect 29235 4696 29251 4760
rect 29315 4696 29331 4760
rect 29395 4696 29579 4760
rect 28301 4694 29579 4696
rect 29641 4760 30313 4762
rect 29641 4696 29825 4760
rect 29889 4696 29905 4760
rect 29969 4696 29985 4760
rect 30049 4696 30065 4760
rect 30129 4696 30313 4760
rect 29641 4694 30313 4696
rect 24631 4683 24756 4693
rect 10813 4646 10985 4656
rect 10813 4500 10823 4646
rect 10973 4500 10985 4646
rect 10813 4490 10985 4500
rect 11165 4650 11337 4660
rect 11165 4504 11175 4650
rect 11325 4504 11337 4650
rect 11165 4494 11337 4504
rect 11611 4650 11783 4660
rect 11611 4504 11621 4650
rect 11771 4504 11783 4650
rect 11611 4494 11783 4504
rect 12177 4654 12349 4664
rect 12177 4508 12187 4654
rect 12337 4508 12349 4654
rect 12177 4498 12349 4508
rect 12843 4654 13015 4664
rect 12843 4508 12853 4654
rect 13003 4508 13015 4654
rect 12843 4498 13015 4508
rect 13225 4638 13397 4648
rect 13225 4492 13235 4638
rect 13385 4492 13397 4638
rect 13225 4482 13397 4492
rect 25685 4312 25799 4325
rect 25685 4248 25708 4312
rect 25772 4248 25799 4312
rect 25685 4238 25799 4248
rect 25859 4311 25973 4324
rect 25859 4247 25882 4311
rect 25946 4247 25973 4311
rect 25859 4237 25973 4247
rect 26084 4313 26198 4326
rect 26084 4249 26107 4313
rect 26171 4249 26198 4313
rect 26084 4239 26198 4249
rect 26285 4315 26399 4328
rect 26285 4251 26308 4315
rect 26372 4251 26399 4315
rect 26285 4241 26399 4251
rect 26508 4313 26622 4326
rect 26508 4249 26531 4313
rect 26595 4249 26622 4313
rect 26508 4239 26622 4249
rect 26717 4318 26831 4331
rect 26717 4254 26740 4318
rect 26804 4254 26831 4318
rect 26717 4244 26831 4254
rect 26945 4311 27059 4324
rect 26945 4247 26968 4311
rect 27032 4247 27059 4311
rect 26945 4237 27059 4247
rect 27135 4315 27249 4328
rect 27135 4251 27158 4315
rect 27222 4251 27249 4315
rect 27135 4241 27249 4251
rect 27340 4318 27454 4331
rect 27340 4254 27363 4318
rect 27427 4254 27454 4318
rect 27340 4244 27454 4254
rect 27539 4318 27653 4331
rect 27539 4254 27562 4318
rect 27626 4254 27653 4318
rect 27539 4244 27653 4254
rect 27755 4313 27869 4326
rect 27755 4249 27778 4313
rect 27842 4249 27869 4313
rect 27755 4239 27869 4249
rect 28143 4318 28257 4331
rect 28143 4254 28166 4318
rect 28230 4254 28257 4318
rect 28143 4244 28257 4254
rect 28378 4313 28492 4326
rect 28378 4249 28401 4313
rect 28465 4249 28492 4313
rect 28378 4239 28492 4249
rect 28620 4315 28734 4328
rect 28620 4251 28643 4315
rect 28707 4251 28734 4315
rect 28620 4241 28734 4251
rect 28852 4316 28966 4329
rect 28852 4252 28875 4316
rect 28939 4252 28966 4316
rect 28852 4242 28966 4252
rect 29081 4319 29195 4332
rect 29081 4255 29104 4319
rect 29168 4255 29195 4319
rect 29081 4245 29195 4255
rect 29330 4311 29444 4324
rect 29330 4247 29353 4311
rect 29417 4247 29444 4311
rect 29330 4237 29444 4247
rect 29548 4315 29662 4328
rect 29548 4251 29571 4315
rect 29635 4251 29662 4315
rect 29548 4241 29662 4251
rect 29777 4311 29891 4324
rect 29777 4247 29800 4311
rect 29864 4247 29891 4311
rect 29777 4237 29891 4247
rect 29998 4313 30112 4326
rect 29998 4249 30021 4313
rect 30085 4249 30112 4313
rect 29998 4239 30112 4249
rect 30214 4318 30328 4331
rect 30214 4254 30237 4318
rect 30301 4254 30328 4318
rect 30214 4244 30328 4254
rect 27043 4125 27157 4138
rect 23595 4088 23767 4098
rect 23595 3942 23605 4088
rect 23755 3942 23767 4088
rect 27043 4061 27066 4125
rect 27130 4061 27157 4125
rect 29438 4124 29552 4137
rect 27043 4051 27157 4061
rect 27428 4074 27542 4087
rect 27428 4010 27451 4074
rect 27515 4010 27542 4074
rect 29438 4060 29461 4124
rect 29525 4060 29552 4124
rect 29438 4050 29552 4060
rect 29823 4075 29937 4088
rect 27428 4000 27542 4010
rect 29823 4011 29846 4075
rect 29910 4011 29937 4075
rect 29823 4001 29937 4011
rect 23595 3932 23767 3942
rect 10895 3792 11067 3802
rect 10895 3646 10905 3792
rect 11055 3646 11067 3792
rect 10895 3636 11067 3646
rect 11245 3800 11417 3810
rect 11245 3654 11255 3800
rect 11405 3654 11417 3800
rect 25687 3729 25801 3742
rect 25687 3665 25710 3729
rect 25774 3665 25801 3729
rect 25687 3655 25801 3665
rect 25862 3727 25976 3740
rect 25862 3663 25885 3727
rect 25949 3663 25976 3727
rect 11245 3644 11417 3654
rect 25862 3653 25976 3663
rect 26059 3729 26173 3742
rect 26059 3665 26082 3729
rect 26146 3665 26173 3729
rect 26059 3655 26173 3665
rect 26278 3732 26392 3745
rect 26278 3668 26301 3732
rect 26365 3668 26392 3732
rect 26278 3658 26392 3668
rect 26510 3728 26624 3741
rect 26510 3664 26533 3728
rect 26597 3664 26624 3728
rect 26510 3654 26624 3664
rect 26734 3735 26848 3748
rect 26734 3671 26757 3735
rect 26821 3671 26848 3735
rect 26734 3661 26848 3671
rect 26946 3723 27060 3736
rect 26946 3659 26969 3723
rect 27033 3659 27060 3723
rect 26946 3649 27060 3659
rect 27168 3719 27282 3732
rect 27168 3655 27191 3719
rect 27255 3655 27282 3719
rect 27168 3645 27282 3655
rect 27391 3716 27505 3729
rect 27391 3652 27414 3716
rect 27478 3652 27505 3716
rect 27391 3642 27505 3652
rect 27601 3716 27715 3729
rect 27601 3652 27624 3716
rect 27688 3652 27715 3716
rect 27601 3642 27715 3652
rect 27814 3716 27928 3729
rect 27814 3652 27837 3716
rect 27901 3652 27928 3716
rect 27814 3642 27928 3652
rect 28131 3709 28245 3722
rect 28131 3645 28154 3709
rect 28218 3645 28245 3709
rect 28131 3635 28245 3645
rect 28333 3712 28447 3725
rect 28333 3648 28356 3712
rect 28420 3648 28447 3712
rect 28333 3638 28447 3648
rect 28534 3713 28648 3726
rect 28534 3649 28557 3713
rect 28621 3649 28648 3713
rect 28534 3639 28648 3649
rect 28713 3714 28827 3727
rect 28713 3650 28736 3714
rect 28800 3650 28827 3714
rect 28713 3640 28827 3650
rect 28905 3718 29019 3731
rect 28905 3654 28928 3718
rect 28992 3654 29019 3718
rect 28905 3644 29019 3654
rect 29090 3715 29204 3728
rect 29090 3651 29113 3715
rect 29177 3651 29204 3715
rect 29090 3641 29204 3651
rect 29322 3714 29436 3727
rect 29322 3650 29345 3714
rect 29409 3650 29436 3714
rect 29322 3640 29436 3650
rect 29527 3716 29641 3729
rect 29527 3652 29550 3716
rect 29614 3652 29641 3716
rect 29527 3642 29641 3652
rect 29733 3718 29847 3731
rect 29733 3654 29756 3718
rect 29820 3654 29847 3718
rect 29733 3644 29847 3654
rect 29941 3725 30055 3738
rect 29941 3661 29964 3725
rect 30028 3661 30055 3725
rect 29941 3651 30055 3661
rect 30163 3726 30277 3739
rect 30163 3662 30186 3726
rect 30250 3662 30277 3726
rect 30163 3652 30277 3662
rect 23601 3410 23773 3420
rect 23601 3264 23611 3410
rect 23761 3264 23773 3410
rect 23601 3254 23773 3264
rect 25714 3080 25828 3093
rect 25714 3016 25737 3080
rect 25801 3016 25828 3080
rect 25714 3006 25828 3016
rect 25930 3085 26044 3098
rect 25930 3021 25953 3085
rect 26017 3021 26044 3085
rect 25930 3011 26044 3021
rect 26136 3086 26250 3099
rect 26136 3022 26159 3086
rect 26223 3022 26250 3086
rect 26136 3012 26250 3022
rect 26338 3078 26452 3091
rect 26338 3014 26361 3078
rect 26425 3014 26452 3078
rect 26338 3004 26452 3014
rect 26534 3080 26648 3093
rect 26534 3016 26557 3080
rect 26621 3016 26648 3080
rect 26534 3006 26648 3016
rect 26759 3082 26873 3095
rect 26759 3018 26782 3082
rect 26846 3018 26873 3082
rect 26759 3008 26873 3018
rect 26974 3078 27088 3091
rect 26974 3014 26997 3078
rect 27061 3014 27088 3078
rect 26974 3004 27088 3014
rect 27209 3078 27323 3091
rect 27209 3014 27232 3078
rect 27296 3014 27323 3078
rect 27209 3004 27323 3014
rect 27417 3081 27531 3094
rect 27417 3017 27440 3081
rect 27504 3017 27531 3081
rect 27417 3007 27531 3017
rect 27659 3081 27773 3094
rect 27659 3017 27682 3081
rect 27746 3017 27773 3081
rect 27659 3007 27773 3017
rect 27857 3082 27971 3095
rect 27857 3018 27880 3082
rect 27944 3018 27971 3082
rect 27857 3008 27971 3018
rect 28164 3082 28278 3095
rect 28164 3018 28187 3082
rect 28251 3018 28278 3082
rect 28164 3008 28278 3018
rect 28389 3083 28503 3096
rect 28389 3019 28412 3083
rect 28476 3019 28503 3083
rect 28389 3009 28503 3019
rect 28618 3082 28732 3095
rect 28618 3018 28641 3082
rect 28705 3018 28732 3082
rect 28618 3008 28732 3018
rect 28834 3086 28948 3099
rect 28834 3022 28857 3086
rect 28921 3022 28948 3086
rect 28834 3012 28948 3022
rect 29057 3089 29171 3102
rect 29057 3025 29080 3089
rect 29144 3025 29171 3089
rect 29057 3015 29171 3025
rect 29281 3085 29395 3098
rect 29281 3021 29304 3085
rect 29368 3021 29395 3085
rect 29281 3011 29395 3021
rect 29508 3074 29622 3087
rect 29508 3010 29531 3074
rect 29595 3010 29622 3074
rect 29508 3000 29622 3010
rect 29721 3073 29835 3086
rect 29721 3009 29744 3073
rect 29808 3009 29835 3073
rect 29721 2999 29835 3009
rect 29932 3077 30046 3090
rect 29932 3013 29955 3077
rect 30019 3013 30046 3077
rect 29932 3003 30046 3013
rect 30159 3078 30273 3091
rect 30159 3014 30182 3078
rect 30246 3014 30273 3078
rect 30159 3004 30273 3014
rect 27048 2851 27162 2864
rect 27048 2787 27071 2851
rect 27135 2787 27162 2851
rect 29440 2853 29554 2866
rect 27048 2777 27162 2787
rect 27431 2792 27545 2805
rect 27431 2728 27454 2792
rect 27518 2728 27545 2792
rect 29440 2789 29463 2853
rect 29527 2789 29554 2853
rect 29440 2779 29554 2789
rect 29817 2799 29931 2812
rect 27431 2718 27545 2728
rect 29817 2735 29840 2799
rect 29904 2735 29931 2799
rect 29817 2725 29931 2735
rect 25740 2435 25854 2448
rect 25740 2371 25763 2435
rect 25827 2371 25854 2435
rect 25740 2361 25854 2371
rect 25965 2444 26079 2457
rect 25965 2380 25988 2444
rect 26052 2380 26079 2444
rect 25965 2370 26079 2380
rect 26242 2441 26356 2454
rect 26242 2377 26265 2441
rect 26329 2377 26356 2441
rect 26242 2367 26356 2377
rect 26463 2444 26577 2457
rect 26463 2380 26486 2444
rect 26550 2380 26577 2444
rect 26463 2370 26577 2380
rect 26708 2441 26822 2454
rect 26708 2377 26731 2441
rect 26795 2377 26822 2441
rect 26708 2367 26822 2377
rect 26934 2445 27048 2458
rect 26934 2381 26957 2445
rect 27021 2381 27048 2445
rect 26934 2371 27048 2381
rect 27146 2443 27260 2456
rect 27146 2379 27169 2443
rect 27233 2379 27260 2443
rect 27146 2369 27260 2379
rect 27366 2449 27480 2462
rect 27366 2385 27389 2449
rect 27453 2385 27480 2449
rect 27366 2375 27480 2385
rect 27604 2451 27718 2464
rect 27604 2387 27627 2451
rect 27691 2387 27718 2451
rect 27604 2377 27718 2387
rect 27817 2453 27931 2466
rect 27817 2389 27840 2453
rect 27904 2389 27931 2453
rect 27817 2379 27931 2389
rect 28204 2443 28318 2456
rect 28204 2379 28227 2443
rect 28291 2379 28318 2443
rect 28204 2369 28318 2379
rect 28551 2444 28665 2457
rect 28551 2380 28574 2444
rect 28638 2380 28665 2444
rect 28551 2370 28665 2380
rect 28787 2439 28901 2452
rect 28787 2375 28810 2439
rect 28874 2375 28901 2439
rect 28787 2365 28901 2375
rect 28971 2439 29085 2452
rect 28971 2375 28994 2439
rect 29058 2375 29085 2439
rect 28971 2365 29085 2375
rect 29210 2441 29324 2454
rect 29210 2377 29233 2441
rect 29297 2377 29324 2441
rect 29210 2367 29324 2377
rect 29413 2437 29527 2450
rect 29413 2373 29436 2437
rect 29500 2373 29527 2437
rect 29413 2363 29527 2373
rect 29598 2434 29712 2447
rect 29598 2370 29621 2434
rect 29685 2370 29712 2434
rect 29598 2360 29712 2370
rect 29789 2436 29903 2449
rect 29789 2372 29812 2436
rect 29876 2372 29903 2436
rect 29789 2362 29903 2372
rect 29980 2440 30094 2453
rect 29980 2376 30003 2440
rect 30067 2376 30094 2440
rect 29980 2366 30094 2376
rect 30166 2436 30280 2449
rect 30166 2372 30189 2436
rect 30253 2372 30280 2436
rect 30166 2362 30280 2372
rect 25613 1853 25727 1866
rect 25613 1789 25636 1853
rect 25700 1789 25727 1853
rect 25613 1779 25727 1789
rect 25818 1849 25932 1862
rect 25818 1785 25841 1849
rect 25905 1785 25932 1849
rect 25818 1775 25932 1785
rect 26004 1854 26118 1867
rect 26004 1790 26027 1854
rect 26091 1790 26118 1854
rect 26004 1780 26118 1790
rect 26198 1847 26312 1860
rect 26198 1783 26221 1847
rect 26285 1783 26312 1847
rect 26198 1773 26312 1783
rect 26417 1852 26531 1865
rect 26417 1788 26440 1852
rect 26504 1788 26531 1852
rect 26417 1778 26531 1788
rect 26627 1852 26741 1865
rect 26627 1788 26650 1852
rect 26714 1788 26741 1852
rect 26627 1778 26741 1788
rect 26856 1849 26970 1862
rect 26856 1785 26879 1849
rect 26943 1785 26970 1849
rect 26856 1775 26970 1785
rect 27102 1849 27216 1862
rect 27102 1785 27125 1849
rect 27189 1785 27216 1849
rect 27102 1775 27216 1785
rect 27376 1849 27490 1862
rect 27376 1785 27399 1849
rect 27463 1785 27490 1849
rect 27376 1775 27490 1785
rect 27651 1849 27765 1862
rect 27651 1785 27674 1849
rect 27738 1785 27765 1849
rect 27651 1775 27765 1785
rect 27887 1849 28001 1862
rect 27887 1785 27910 1849
rect 27974 1785 28001 1849
rect 27887 1775 28001 1785
rect 28110 1852 28224 1865
rect 28110 1788 28133 1852
rect 28197 1788 28224 1852
rect 28110 1778 28224 1788
rect 28328 1855 28442 1868
rect 28328 1791 28351 1855
rect 28415 1791 28442 1855
rect 28328 1781 28442 1791
rect 28506 1846 28620 1859
rect 28506 1782 28529 1846
rect 28593 1782 28620 1846
rect 28506 1772 28620 1782
rect 28745 1848 28859 1861
rect 28745 1784 28768 1848
rect 28832 1784 28859 1848
rect 28745 1774 28859 1784
rect 28942 1848 29056 1861
rect 28942 1784 28965 1848
rect 29029 1784 29056 1848
rect 28942 1774 29056 1784
rect 29140 1848 29254 1861
rect 29140 1784 29163 1848
rect 29227 1784 29254 1848
rect 29140 1774 29254 1784
rect 29353 1849 29467 1862
rect 29353 1785 29376 1849
rect 29440 1785 29467 1849
rect 29353 1775 29467 1785
rect 29576 1848 29690 1861
rect 29576 1784 29599 1848
rect 29663 1784 29690 1848
rect 29576 1774 29690 1784
rect 29773 1853 29887 1866
rect 29773 1789 29796 1853
rect 29860 1789 29887 1853
rect 29773 1779 29887 1789
rect 29989 1851 30103 1864
rect 29989 1787 30012 1851
rect 30076 1787 30103 1851
rect 29989 1777 30103 1787
rect 30198 1851 30312 1864
rect 30198 1787 30221 1851
rect 30285 1787 30312 1851
rect 30198 1777 30312 1787
rect 8591 1417 8720 1428
rect 8591 1353 8622 1417
rect 8686 1353 8720 1417
rect 8591 1342 8720 1353
rect 8793 1419 8922 1430
rect 8793 1355 8824 1419
rect 8888 1355 8922 1419
rect 8793 1344 8922 1355
rect 9004 1417 9133 1428
rect 9004 1353 9035 1417
rect 9099 1353 9133 1417
rect 9004 1342 9133 1353
rect 9194 1417 9323 1428
rect 9194 1353 9225 1417
rect 9289 1353 9323 1417
rect 9194 1342 9323 1353
rect 9402 1419 9531 1430
rect 9402 1355 9433 1419
rect 9497 1355 9531 1419
rect 9402 1344 9531 1355
rect 9604 1419 9733 1430
rect 9604 1355 9635 1419
rect 9699 1355 9733 1419
rect 9604 1344 9733 1355
rect 9803 1421 9932 1432
rect 9803 1357 9834 1421
rect 9898 1357 9932 1421
rect 9803 1346 9932 1357
rect 9998 1418 10127 1429
rect 9998 1354 10029 1418
rect 10093 1354 10127 1418
rect 9998 1343 10127 1354
rect 10199 1420 10328 1431
rect 10199 1356 10230 1420
rect 10294 1356 10328 1420
rect 10199 1345 10328 1356
rect 10416 1418 10545 1429
rect 10416 1354 10447 1418
rect 10511 1354 10545 1418
rect 10416 1343 10545 1354
rect 10690 1421 10819 1432
rect 10690 1357 10721 1421
rect 10785 1357 10819 1421
rect 10690 1346 10819 1357
rect 10967 1414 11096 1425
rect 10967 1350 10998 1414
rect 11062 1350 11096 1414
rect 10967 1339 11096 1350
rect 11190 1417 11319 1428
rect 11190 1353 11221 1417
rect 11285 1353 11319 1417
rect 11190 1342 11319 1353
rect 11422 1416 11551 1427
rect 11422 1352 11453 1416
rect 11517 1352 11551 1416
rect 11422 1341 11551 1352
rect 13058 1413 13187 1424
rect 13058 1349 13089 1413
rect 13153 1349 13187 1413
rect 13058 1338 13187 1349
rect 13366 1414 13495 1425
rect 13366 1350 13397 1414
rect 13461 1350 13495 1414
rect 13366 1339 13495 1350
rect 13566 1415 13695 1426
rect 13566 1351 13597 1415
rect 13661 1351 13695 1415
rect 13566 1340 13695 1351
rect 13785 1414 13914 1425
rect 13785 1350 13816 1414
rect 13880 1350 13914 1414
rect 13785 1339 13914 1350
rect 14031 1413 14160 1424
rect 14031 1349 14062 1413
rect 14126 1349 14160 1413
rect 14031 1338 14160 1349
rect 14239 1415 14368 1426
rect 14239 1351 14270 1415
rect 14334 1351 14368 1415
rect 14239 1340 14368 1351
rect 14441 1416 14570 1427
rect 14441 1352 14472 1416
rect 14536 1352 14570 1416
rect 14441 1341 14570 1352
rect 14634 1415 14763 1426
rect 14634 1351 14665 1415
rect 14729 1351 14763 1415
rect 14634 1340 14763 1351
rect 15006 1414 15135 1425
rect 15006 1350 15037 1414
rect 15101 1350 15135 1414
rect 15006 1339 15135 1350
rect 15195 1412 15324 1423
rect 15195 1348 15226 1412
rect 15290 1348 15324 1412
rect 15195 1337 15324 1348
rect 15485 1412 15614 1423
rect 15485 1348 15516 1412
rect 15580 1348 15614 1412
rect 15485 1337 15614 1348
rect 15758 1414 15887 1425
rect 15758 1350 15789 1414
rect 15853 1350 15887 1414
rect 15758 1339 15887 1350
rect 9709 878 9838 889
rect 9709 814 9740 878
rect 9804 814 9838 878
rect 9709 803 9838 814
rect 9928 882 10057 893
rect 9928 818 9959 882
rect 10023 818 10057 882
rect 9928 807 10057 818
rect 10211 882 10340 893
rect 10211 818 10242 882
rect 10306 818 10340 882
rect 10211 807 10340 818
rect 10420 882 10549 893
rect 10420 818 10451 882
rect 10515 818 10549 882
rect 10420 807 10549 818
rect 10691 880 10820 891
rect 10691 816 10722 880
rect 10786 816 10820 880
rect 10691 805 10820 816
rect 12766 878 12895 889
rect 12766 814 12797 878
rect 12861 814 12895 878
rect 12766 803 12895 814
rect 13015 881 13144 892
rect 13015 817 13046 881
rect 13110 817 13144 881
rect 13015 806 13144 817
rect 13359 867 13488 878
rect 13359 803 13390 867
rect 13454 803 13488 867
rect 13359 792 13488 803
rect 13613 873 13742 884
rect 13613 809 13644 873
rect 13708 809 13742 873
rect 13613 798 13742 809
rect 13842 873 13971 884
rect 13842 809 13873 873
rect 13937 809 13971 873
rect 13842 798 13971 809
rect 15560 878 15689 889
rect 15560 814 15591 878
rect 15655 814 15689 878
rect 15560 803 15689 814
rect 15764 880 15893 891
rect 15764 816 15795 880
rect 15859 816 15893 880
rect 15764 805 15893 816
rect 16087 878 16216 889
rect 16087 814 16118 878
rect 16182 814 16216 878
rect 16087 803 16216 814
rect 8557 273 8686 284
rect 8557 209 8588 273
rect 8652 209 8686 273
rect 8557 198 8686 209
rect 8797 271 8926 282
rect 8797 207 8828 271
rect 8892 207 8926 271
rect 8797 196 8926 207
rect 9119 270 9248 281
rect 9119 206 9150 270
rect 9214 206 9248 270
rect 9119 195 9248 206
rect 9337 271 9466 282
rect 9337 207 9368 271
rect 9432 207 9466 271
rect 9337 196 9466 207
rect 11241 275 11370 286
rect 11241 211 11272 275
rect 11336 211 11370 275
rect 11241 200 11370 211
rect 11566 277 11695 288
rect 11566 213 11597 277
rect 11661 213 11695 277
rect 11566 202 11695 213
rect 11834 277 11963 288
rect 11834 213 11865 277
rect 11929 213 11963 277
rect 11834 202 11963 213
rect 12100 277 12229 288
rect 12100 213 12131 277
rect 12195 213 12229 277
rect 12100 202 12229 213
rect 12340 275 12469 286
rect 12340 211 12371 275
rect 12435 211 12469 275
rect 12340 200 12469 211
rect 14134 278 14263 289
rect 14134 214 14165 278
rect 14229 214 14263 278
rect 14134 203 14263 214
rect 14500 281 14629 292
rect 14500 217 14531 281
rect 14595 217 14629 281
rect 14500 206 14629 217
rect 14744 281 14873 292
rect 14744 217 14775 281
rect 14839 217 14873 281
rect 14744 206 14873 217
rect 15167 272 15296 283
rect 15167 208 15198 272
rect 15262 208 15296 272
rect 15167 197 15296 208
rect 17110 274 17239 285
rect 17110 210 17141 274
rect 17205 210 17239 274
rect 17110 199 17239 210
rect 17362 271 17491 282
rect 17362 207 17393 271
rect 17457 207 17491 271
rect 17362 196 17491 207
rect 17568 279 17697 290
rect 17568 215 17599 279
rect 17663 215 17697 279
rect 17568 204 17697 215
rect 17851 273 17980 284
rect 17851 209 17882 273
rect 17946 209 17980 273
rect 17851 198 17980 209
rect 18149 274 18278 285
rect 18149 210 18180 274
rect 18244 210 18278 274
rect 18149 199 18278 210
rect 19981 275 20110 286
rect 19981 211 20012 275
rect 20076 211 20110 275
rect 19981 200 20110 211
rect 20191 277 20320 288
rect 20191 213 20222 277
rect 20286 213 20320 277
rect 20191 202 20320 213
rect 20542 275 20671 286
rect 20542 211 20573 275
rect 20637 211 20671 275
rect 20542 200 20671 211
rect 20822 275 20951 286
rect 20822 211 20853 275
rect 20917 211 20951 275
rect 20822 200 20951 211
rect 21139 274 21268 285
rect 21139 210 21170 274
rect 21234 210 21268 274
rect 21139 199 21268 210
rect 22929 272 23058 283
rect 22929 208 22960 272
rect 23024 208 23058 272
rect 22929 197 23058 208
rect 23224 272 23353 283
rect 23224 208 23255 272
rect 23319 208 23353 272
rect 23224 197 23353 208
rect 23511 272 23640 283
rect 23511 208 23542 272
rect 23606 208 23640 272
rect 23511 197 23640 208
rect 23801 272 23930 283
rect 23801 208 23832 272
rect 23896 208 23930 272
rect 23801 197 23930 208
rect 24085 275 24214 286
rect 24085 211 24116 275
rect 24180 211 24214 275
rect 24085 200 24214 211
rect 9748 -265 9877 -254
rect 9748 -329 9779 -265
rect 9843 -329 9877 -265
rect 9748 -340 9877 -329
rect 9965 -265 10094 -254
rect 9965 -329 9996 -265
rect 10060 -329 10094 -265
rect 9965 -340 10094 -329
rect 10184 -265 10313 -254
rect 10184 -329 10215 -265
rect 10279 -329 10313 -265
rect 10184 -340 10313 -329
rect 10397 -269 10526 -258
rect 10397 -333 10428 -269
rect 10492 -333 10526 -269
rect 10397 -344 10526 -333
rect 10608 -269 10737 -258
rect 10608 -333 10639 -269
rect 10703 -333 10737 -269
rect 10608 -344 10737 -333
rect 12732 -269 12861 -258
rect 12732 -333 12763 -269
rect 12827 -333 12861 -269
rect 12732 -344 12861 -333
rect 13010 -270 13139 -259
rect 13010 -334 13041 -270
rect 13105 -334 13139 -270
rect 13010 -345 13139 -334
rect 13582 -265 13711 -254
rect 13582 -329 13613 -265
rect 13677 -329 13711 -265
rect 13582 -340 13711 -329
rect 13821 -265 13950 -254
rect 13821 -329 13852 -265
rect 13916 -329 13950 -265
rect 13821 -340 13950 -329
rect 15979 -267 16108 -256
rect 15979 -331 16010 -267
rect 16074 -331 16108 -267
rect 15979 -342 16108 -331
rect 16206 -262 16335 -251
rect 16206 -326 16237 -262
rect 16301 -326 16335 -262
rect 16206 -337 16335 -326
rect 16396 -260 16525 -249
rect 16396 -324 16427 -260
rect 16491 -324 16525 -260
rect 16396 -335 16525 -324
rect 16612 -269 16741 -258
rect 16612 -333 16643 -269
rect 16707 -333 16741 -269
rect 16612 -344 16741 -333
rect 18593 -266 18722 -255
rect 18593 -330 18624 -266
rect 18688 -330 18722 -266
rect 18593 -341 18722 -330
rect 18822 -263 18951 -252
rect 18822 -327 18853 -263
rect 18917 -327 18951 -263
rect 18822 -338 18951 -327
rect 19048 -258 19177 -247
rect 19048 -322 19079 -258
rect 19143 -322 19177 -258
rect 19048 -333 19177 -322
rect 19276 -266 19405 -255
rect 19276 -330 19307 -266
rect 19371 -330 19405 -266
rect 19276 -341 19405 -330
rect 19512 -260 19641 -249
rect 19512 -324 19543 -260
rect 19607 -324 19641 -260
rect 19512 -335 19641 -324
rect 19704 -269 19833 -258
rect 19704 -333 19735 -269
rect 19799 -333 19833 -269
rect 19704 -344 19833 -333
rect 21439 -269 21568 -258
rect 21439 -333 21470 -269
rect 21534 -333 21568 -269
rect 21439 -344 21568 -333
rect 21643 -264 21772 -253
rect 21643 -328 21674 -264
rect 21738 -328 21772 -264
rect 21643 -339 21772 -328
rect 21834 -269 21963 -258
rect 21834 -333 21865 -269
rect 21929 -333 21963 -269
rect 21834 -344 21963 -333
rect 22036 -270 22165 -259
rect 22036 -334 22067 -270
rect 22131 -334 22165 -270
rect 22036 -345 22165 -334
rect 22326 -269 22455 -258
rect 22326 -333 22357 -269
rect 22421 -333 22455 -269
rect 22326 -344 22455 -333
rect 22611 -270 22740 -259
rect 22611 -334 22642 -270
rect 22706 -334 22740 -270
rect 22611 -345 22740 -334
rect 24366 -265 24495 -254
rect 24366 -329 24397 -265
rect 24461 -329 24495 -265
rect 24366 -340 24495 -329
rect 24560 -261 24689 -250
rect 24560 -325 24591 -261
rect 24655 -325 24689 -261
rect 24560 -336 24689 -325
rect 24749 -264 24878 -253
rect 24749 -328 24780 -264
rect 24844 -328 24878 -264
rect 24749 -339 24878 -328
rect 24972 -262 25101 -251
rect 24972 -326 25003 -262
rect 25067 -326 25101 -262
rect 24972 -337 25101 -326
rect 8803 -410 8932 -399
rect 8803 -474 8834 -410
rect 8898 -474 8932 -410
rect 8803 -485 8932 -474
rect 9005 -414 9134 -403
rect 9005 -478 9036 -414
rect 9100 -478 9134 -414
rect 9005 -489 9134 -478
rect 9194 -417 9323 -406
rect 9194 -481 9225 -417
rect 9289 -481 9323 -417
rect 9194 -492 9323 -481
rect 9423 -416 9552 -405
rect 9423 -480 9454 -416
rect 9518 -480 9552 -416
rect 9423 -491 9552 -480
rect 11192 -413 11321 -402
rect 11192 -477 11223 -413
rect 11287 -477 11321 -413
rect 11192 -488 11321 -477
rect 11407 -416 11536 -405
rect 11407 -480 11438 -416
rect 11502 -480 11536 -416
rect 11407 -491 11536 -480
rect 11605 -419 11734 -408
rect 11605 -483 11636 -419
rect 11700 -483 11734 -419
rect 11605 -494 11734 -483
rect 11800 -409 11929 -398
rect 11800 -473 11831 -409
rect 11895 -473 11929 -409
rect 11800 -484 11929 -473
rect 12080 -411 12209 -400
rect 12080 -475 12111 -411
rect 12175 -475 12209 -411
rect 12080 -486 12209 -475
rect 12299 -413 12428 -402
rect 12299 -477 12330 -413
rect 12394 -477 12428 -413
rect 12299 -488 12428 -477
rect 14120 -416 14249 -405
rect 14120 -480 14151 -416
rect 14215 -480 14249 -416
rect 14120 -491 14249 -480
rect 14471 -419 14600 -408
rect 14471 -483 14502 -419
rect 14566 -483 14600 -419
rect 14471 -494 14600 -483
rect 14660 -421 14789 -410
rect 14660 -485 14691 -421
rect 14755 -485 14789 -421
rect 14660 -496 14789 -485
rect 14865 -414 14994 -403
rect 14865 -478 14896 -414
rect 14960 -478 14994 -414
rect 14865 -489 14994 -478
rect 15056 -412 15185 -401
rect 15056 -476 15087 -412
rect 15151 -476 15185 -412
rect 15056 -487 15185 -476
rect 17101 -410 17230 -399
rect 17101 -474 17132 -410
rect 17196 -474 17230 -410
rect 17101 -485 17230 -474
rect 17291 -408 17420 -397
rect 17291 -472 17322 -408
rect 17386 -472 17420 -408
rect 17291 -483 17420 -472
rect 17485 -410 17614 -399
rect 17485 -474 17516 -410
rect 17580 -474 17614 -410
rect 17485 -485 17614 -474
rect 17796 -414 17925 -403
rect 17796 -478 17827 -414
rect 17891 -478 17925 -414
rect 17796 -489 17925 -478
rect 19979 -415 20108 -404
rect 19979 -479 20010 -415
rect 20074 -479 20108 -415
rect 19979 -490 20108 -479
rect 20183 -415 20312 -404
rect 20183 -479 20214 -415
rect 20278 -479 20312 -415
rect 20183 -490 20312 -479
rect 20748 -419 20877 -408
rect 20748 -483 20779 -419
rect 20843 -483 20877 -419
rect 20748 -494 20877 -483
rect 20987 -417 21116 -406
rect 20987 -481 21018 -417
rect 21082 -481 21116 -417
rect 20987 -492 21116 -481
rect 21191 -417 21320 -406
rect 21191 -481 21222 -417
rect 21286 -481 21320 -417
rect 21191 -492 21320 -481
rect 23151 -409 23280 -398
rect 23151 -473 23182 -409
rect 23246 -473 23280 -409
rect 23151 -484 23280 -473
rect 23384 -411 23513 -400
rect 23384 -475 23415 -411
rect 23479 -475 23513 -411
rect 23384 -486 23513 -475
rect 23591 -413 23720 -402
rect 23591 -477 23622 -413
rect 23686 -477 23720 -413
rect 23591 -488 23720 -477
rect 23800 -411 23929 -400
rect 23800 -475 23831 -411
rect 23895 -475 23929 -411
rect 23800 -486 23929 -475
rect 24080 -409 24209 -398
rect 24080 -473 24111 -409
rect 24175 -473 24209 -409
rect 24080 -484 24209 -473
rect 9959 -947 10088 -936
rect 9730 -959 9859 -948
rect 9730 -1023 9761 -959
rect 9825 -1023 9859 -959
rect 9959 -1011 9990 -947
rect 10054 -1011 10088 -947
rect 9959 -1022 10088 -1011
rect 10178 -957 10307 -946
rect 10178 -1021 10209 -957
rect 10273 -1021 10307 -957
rect 9730 -1034 9859 -1023
rect 10178 -1032 10307 -1021
rect 10370 -953 10499 -942
rect 10370 -1017 10401 -953
rect 10465 -1017 10499 -953
rect 10370 -1028 10499 -1017
rect 10864 -955 10993 -944
rect 10864 -1019 10895 -955
rect 10959 -1019 10993 -955
rect 10864 -1030 10993 -1019
rect 12656 -956 12785 -945
rect 12656 -1020 12687 -956
rect 12751 -1020 12785 -956
rect 12656 -1031 12785 -1020
rect 13049 -958 13178 -947
rect 13049 -1022 13080 -958
rect 13144 -1022 13178 -958
rect 13049 -1033 13178 -1022
rect 13246 -950 13375 -939
rect 13246 -1014 13277 -950
rect 13341 -1014 13375 -950
rect 13246 -1025 13375 -1014
rect 13576 -948 13705 -937
rect 13576 -1012 13607 -948
rect 13671 -1012 13705 -948
rect 13576 -1023 13705 -1012
rect 13772 -948 13901 -937
rect 13772 -1012 13803 -948
rect 13867 -1012 13901 -948
rect 13772 -1023 13901 -1012
rect 15679 -955 15808 -944
rect 15679 -1019 15710 -955
rect 15774 -1019 15808 -955
rect 15679 -1030 15808 -1019
rect 15980 -951 16109 -940
rect 15980 -1015 16011 -951
rect 16075 -1015 16109 -951
rect 15980 -1026 16109 -1015
rect 16186 -950 16315 -939
rect 16186 -1014 16217 -950
rect 16281 -1014 16315 -950
rect 16186 -1025 16315 -1014
rect 16396 -954 16525 -943
rect 16396 -1018 16427 -954
rect 16491 -1018 16525 -954
rect 16396 -1029 16525 -1018
rect 16607 -948 16736 -937
rect 16607 -1012 16638 -948
rect 16702 -1012 16736 -948
rect 16607 -1023 16736 -1012
rect 18487 -959 18616 -948
rect 18487 -1023 18518 -959
rect 18582 -1023 18616 -959
rect 18487 -1034 18616 -1023
rect 18744 -952 18873 -941
rect 18744 -1016 18775 -952
rect 18839 -1016 18873 -952
rect 18744 -1027 18873 -1016
rect 18994 -956 19123 -945
rect 18994 -1020 19025 -956
rect 19089 -1020 19123 -956
rect 18994 -1031 19123 -1020
rect 19265 -951 19394 -940
rect 19265 -1015 19296 -951
rect 19360 -1015 19394 -951
rect 19265 -1026 19394 -1015
rect 19506 -948 19635 -937
rect 19506 -1012 19537 -948
rect 19601 -1012 19635 -948
rect 19506 -1023 19635 -1012
rect 19731 -952 19860 -941
rect 19731 -1016 19762 -952
rect 19826 -1016 19860 -952
rect 19731 -1027 19860 -1016
rect 21438 -954 21567 -943
rect 21438 -1018 21469 -954
rect 21533 -1018 21567 -954
rect 21438 -1029 21567 -1018
rect 21639 -953 21768 -942
rect 21639 -1017 21670 -953
rect 21734 -1017 21768 -953
rect 21639 -1028 21768 -1017
rect 21857 -957 21986 -946
rect 21857 -1021 21888 -957
rect 21952 -1021 21986 -957
rect 21857 -1032 21986 -1021
rect 22064 -953 22193 -942
rect 22064 -1017 22095 -953
rect 22159 -1017 22193 -953
rect 22064 -1028 22193 -1017
rect 22269 -954 22398 -943
rect 22269 -1018 22300 -954
rect 22364 -1018 22398 -954
rect 22269 -1029 22398 -1018
rect 22616 -958 22745 -947
rect 22616 -1022 22647 -958
rect 22711 -1022 22745 -958
rect 22616 -1033 22745 -1022
rect 24368 -954 24497 -943
rect 24368 -1018 24399 -954
rect 24463 -1018 24497 -954
rect 24368 -1029 24497 -1018
rect 24559 -951 24688 -940
rect 24559 -1015 24590 -951
rect 24654 -1015 24688 -951
rect 24559 -1026 24688 -1015
rect 24754 -949 24883 -938
rect 24754 -1013 24785 -949
rect 24849 -1013 24883 -949
rect 24754 -1024 24883 -1013
rect 25201 -954 25330 -943
rect 25201 -1018 25232 -954
rect 25296 -1018 25330 -954
rect 25201 -1029 25330 -1018
rect 8585 -1103 8714 -1092
rect 8585 -1167 8616 -1103
rect 8680 -1167 8714 -1103
rect 8585 -1178 8714 -1167
rect 8818 -1107 8947 -1096
rect 8818 -1171 8849 -1107
rect 8913 -1171 8947 -1107
rect 8818 -1182 8947 -1171
rect 9033 -1100 9162 -1089
rect 9033 -1164 9064 -1100
rect 9128 -1164 9162 -1100
rect 9033 -1175 9162 -1164
rect 9251 -1103 9380 -1092
rect 9251 -1167 9282 -1103
rect 9346 -1167 9380 -1103
rect 9251 -1178 9380 -1167
rect 9467 -1102 9596 -1091
rect 9467 -1166 9498 -1102
rect 9562 -1166 9596 -1102
rect 9467 -1177 9596 -1166
rect 11188 -1106 11317 -1095
rect 11188 -1170 11219 -1106
rect 11283 -1170 11317 -1106
rect 11188 -1181 11317 -1170
rect 11378 -1106 11507 -1095
rect 11378 -1170 11409 -1106
rect 11473 -1170 11507 -1106
rect 11378 -1181 11507 -1170
rect 11588 -1103 11717 -1092
rect 11588 -1167 11619 -1103
rect 11683 -1167 11717 -1103
rect 11588 -1178 11717 -1167
rect 11805 -1106 11934 -1095
rect 11805 -1170 11836 -1106
rect 11900 -1170 11934 -1106
rect 11805 -1181 11934 -1170
rect 12100 -1103 12229 -1092
rect 12100 -1167 12131 -1103
rect 12195 -1167 12229 -1103
rect 12100 -1178 12229 -1167
rect 12324 -1098 12453 -1087
rect 12324 -1162 12355 -1098
rect 12419 -1162 12453 -1098
rect 12324 -1173 12453 -1162
rect 14202 -1105 14331 -1094
rect 14202 -1169 14233 -1105
rect 14297 -1169 14331 -1105
rect 14202 -1180 14331 -1169
rect 14502 -1107 14631 -1096
rect 14502 -1171 14533 -1107
rect 14597 -1171 14631 -1107
rect 14502 -1182 14631 -1171
rect 14754 -1103 14883 -1092
rect 14754 -1167 14785 -1103
rect 14849 -1167 14883 -1103
rect 14754 -1178 14883 -1167
rect 14971 -1098 15100 -1087
rect 14971 -1162 15002 -1098
rect 15066 -1162 15100 -1098
rect 14971 -1173 15100 -1162
rect 15172 -1101 15301 -1090
rect 15172 -1165 15203 -1101
rect 15267 -1165 15301 -1101
rect 15172 -1176 15301 -1165
rect 17057 -1110 17186 -1099
rect 17057 -1174 17088 -1110
rect 17152 -1174 17186 -1110
rect 17057 -1185 17186 -1174
rect 17249 -1110 17378 -1099
rect 17249 -1174 17280 -1110
rect 17344 -1174 17378 -1110
rect 17249 -1185 17378 -1174
rect 17449 -1110 17578 -1099
rect 17449 -1174 17480 -1110
rect 17544 -1174 17578 -1110
rect 17449 -1185 17578 -1174
rect 18067 -1102 18196 -1091
rect 18067 -1166 18098 -1102
rect 18162 -1166 18196 -1102
rect 18067 -1177 18196 -1166
rect 19968 -1106 20097 -1095
rect 19968 -1170 19999 -1106
rect 20063 -1170 20097 -1106
rect 19968 -1181 20097 -1170
rect 20224 -1106 20353 -1095
rect 20224 -1170 20255 -1106
rect 20319 -1170 20353 -1106
rect 20224 -1181 20353 -1170
rect 20459 -1106 20588 -1095
rect 20459 -1170 20490 -1106
rect 20554 -1170 20588 -1106
rect 20459 -1181 20588 -1170
rect 20748 -1104 20877 -1093
rect 20748 -1168 20779 -1104
rect 20843 -1168 20877 -1104
rect 20748 -1179 20877 -1168
rect 20938 -1106 21067 -1095
rect 20938 -1170 20969 -1106
rect 21033 -1170 21067 -1106
rect 20938 -1181 21067 -1170
rect 21142 -1104 21271 -1093
rect 21142 -1168 21173 -1104
rect 21237 -1168 21271 -1104
rect 21142 -1179 21271 -1168
rect 22928 -1098 23057 -1087
rect 22928 -1162 22959 -1098
rect 23023 -1162 23057 -1098
rect 22928 -1173 23057 -1162
rect 23170 -1102 23299 -1091
rect 23170 -1166 23201 -1102
rect 23265 -1166 23299 -1102
rect 23170 -1177 23299 -1166
rect 23370 -1103 23499 -1092
rect 23370 -1167 23401 -1103
rect 23465 -1167 23499 -1103
rect 23370 -1178 23499 -1167
rect 23560 -1095 23689 -1084
rect 23560 -1159 23591 -1095
rect 23655 -1159 23689 -1095
rect 23560 -1170 23689 -1159
rect 23781 -1097 23910 -1086
rect 23781 -1161 23812 -1097
rect 23876 -1161 23910 -1097
rect 23781 -1172 23910 -1161
rect 24077 -1102 24206 -1091
rect 24077 -1166 24108 -1102
rect 24172 -1166 24206 -1102
rect 24077 -1177 24206 -1166
rect 8959 -1635 9088 -1624
rect 8959 -1699 8990 -1635
rect 9054 -1699 9088 -1635
rect 8959 -1710 9088 -1699
rect 9158 -1638 9287 -1627
rect 9158 -1702 9189 -1638
rect 9253 -1702 9287 -1638
rect 9158 -1713 9287 -1702
rect 9369 -1638 9498 -1627
rect 9369 -1702 9400 -1638
rect 9464 -1702 9498 -1638
rect 9369 -1713 9498 -1702
rect 9575 -1638 9704 -1627
rect 9575 -1702 9606 -1638
rect 9670 -1702 9704 -1638
rect 9575 -1713 9704 -1702
rect 9803 -1640 9932 -1629
rect 9803 -1704 9834 -1640
rect 9898 -1704 9932 -1640
rect 9803 -1715 9932 -1704
rect 10047 -1640 10176 -1629
rect 10047 -1704 10078 -1640
rect 10142 -1704 10176 -1640
rect 10047 -1715 10176 -1704
rect 10277 -1638 10406 -1627
rect 10277 -1702 10308 -1638
rect 10372 -1702 10406 -1638
rect 10277 -1713 10406 -1702
rect 10483 -1638 10612 -1627
rect 10483 -1702 10514 -1638
rect 10578 -1702 10612 -1638
rect 10483 -1713 10612 -1702
rect 10701 -1633 10830 -1622
rect 10701 -1697 10732 -1633
rect 10796 -1697 10830 -1633
rect 10701 -1708 10830 -1697
rect 10904 -1639 11033 -1628
rect 10904 -1703 10935 -1639
rect 10999 -1703 11033 -1639
rect 10904 -1714 11033 -1703
rect 11112 -1636 11241 -1625
rect 11112 -1700 11143 -1636
rect 11207 -1700 11241 -1636
rect 11112 -1711 11241 -1700
rect 11375 -1640 11504 -1629
rect 11375 -1704 11406 -1640
rect 11470 -1704 11504 -1640
rect 11375 -1715 11504 -1704
rect 11583 -1639 11712 -1628
rect 11583 -1703 11614 -1639
rect 11678 -1703 11712 -1639
rect 11583 -1714 11712 -1703
rect 11793 -1642 11922 -1631
rect 11793 -1706 11824 -1642
rect 11888 -1706 11922 -1642
rect 11793 -1717 11922 -1706
rect 11993 -1636 12122 -1625
rect 11993 -1700 12024 -1636
rect 12088 -1700 12122 -1636
rect 11993 -1711 12122 -1700
rect 12196 -1639 12325 -1628
rect 12196 -1703 12227 -1639
rect 12291 -1703 12325 -1639
rect 12196 -1714 12325 -1703
rect 12406 -1639 12535 -1628
rect 12406 -1703 12437 -1639
rect 12501 -1703 12535 -1639
rect 12406 -1714 12535 -1703
rect 12607 -1638 12736 -1627
rect 12607 -1702 12638 -1638
rect 12702 -1702 12736 -1638
rect 12607 -1713 12736 -1702
rect 12823 -1637 12952 -1626
rect 12823 -1701 12854 -1637
rect 12918 -1701 12952 -1637
rect 12823 -1712 12952 -1701
rect 13104 -1639 13233 -1628
rect 13104 -1703 13135 -1639
rect 13199 -1703 13233 -1639
rect 13104 -1714 13233 -1703
rect 13324 -1644 13453 -1633
rect 13324 -1708 13355 -1644
rect 13419 -1708 13453 -1644
rect 13324 -1719 13453 -1708
rect 13529 -1643 13658 -1632
rect 13529 -1707 13560 -1643
rect 13624 -1707 13658 -1643
rect 13529 -1718 13658 -1707
rect 13750 -1637 13879 -1626
rect 13750 -1701 13781 -1637
rect 13845 -1701 13879 -1637
rect 13750 -1712 13879 -1701
rect 13955 -1644 14084 -1633
rect 13955 -1708 13986 -1644
rect 14050 -1708 14084 -1644
rect 13955 -1719 14084 -1708
rect 14164 -1643 14293 -1632
rect 14164 -1707 14195 -1643
rect 14259 -1707 14293 -1643
rect 14164 -1718 14293 -1707
rect 14381 -1643 14510 -1632
rect 14381 -1707 14412 -1643
rect 14476 -1707 14510 -1643
rect 14381 -1718 14510 -1707
rect 14595 -1638 14724 -1627
rect 14595 -1702 14626 -1638
rect 14690 -1702 14724 -1638
rect 14595 -1713 14724 -1702
rect 14790 -1640 14919 -1629
rect 14790 -1704 14821 -1640
rect 14885 -1704 14919 -1640
rect 14790 -1715 14919 -1704
rect 14985 -1643 15114 -1632
rect 14985 -1707 15016 -1643
rect 15080 -1707 15114 -1643
rect 14985 -1718 15114 -1707
rect 15187 -1640 15316 -1629
rect 15187 -1704 15218 -1640
rect 15282 -1704 15316 -1640
rect 15187 -1715 15316 -1704
rect 15471 -1639 15600 -1628
rect 15471 -1703 15502 -1639
rect 15566 -1703 15600 -1639
rect 15471 -1714 15600 -1703
rect 15670 -1638 15799 -1627
rect 15670 -1702 15701 -1638
rect 15765 -1702 15799 -1638
rect 15670 -1713 15799 -1702
rect 15873 -1636 16002 -1625
rect 15873 -1700 15904 -1636
rect 15968 -1700 16002 -1636
rect 15873 -1711 16002 -1700
rect 16138 -1639 16267 -1628
rect 16138 -1703 16169 -1639
rect 16233 -1703 16267 -1639
rect 16138 -1714 16267 -1703
rect 16336 -1640 16465 -1629
rect 16336 -1704 16367 -1640
rect 16431 -1704 16465 -1640
rect 16336 -1715 16465 -1704
rect 16525 -1638 16654 -1627
rect 16525 -1702 16556 -1638
rect 16620 -1702 16654 -1638
rect 16525 -1713 16654 -1702
rect 16737 -1638 16866 -1627
rect 16737 -1702 16768 -1638
rect 16832 -1702 16866 -1638
rect 16737 -1713 16866 -1702
rect 16954 -1638 17083 -1627
rect 16954 -1702 16985 -1638
rect 17049 -1702 17083 -1638
rect 16954 -1713 17083 -1702
rect 17159 -1642 17288 -1631
rect 17159 -1706 17190 -1642
rect 17254 -1706 17288 -1642
rect 17159 -1717 17288 -1706
rect 17364 -1642 17493 -1631
rect 17364 -1706 17395 -1642
rect 17459 -1706 17493 -1642
rect 17364 -1717 17493 -1706
rect 17572 -1637 17701 -1626
rect 17572 -1701 17603 -1637
rect 17667 -1701 17701 -1637
rect 17572 -1712 17701 -1701
rect 17855 -1638 17984 -1627
rect 17855 -1702 17886 -1638
rect 17950 -1702 17984 -1638
rect 17855 -1713 17984 -1702
rect 18048 -1640 18177 -1629
rect 18048 -1704 18079 -1640
rect 18143 -1704 18177 -1640
rect 18048 -1715 18177 -1704
rect 18274 -1642 18403 -1631
rect 18274 -1706 18305 -1642
rect 18369 -1706 18403 -1642
rect 18274 -1717 18403 -1706
rect 18539 -1642 18668 -1631
rect 18539 -1706 18570 -1642
rect 18634 -1706 18668 -1642
rect 18539 -1717 18668 -1706
rect 18733 -1638 18862 -1627
rect 18733 -1702 18764 -1638
rect 18828 -1702 18862 -1638
rect 18733 -1713 18862 -1702
rect 18931 -1647 19060 -1636
rect 18931 -1711 18962 -1647
rect 19026 -1711 19060 -1647
rect 18931 -1722 19060 -1711
rect 19135 -1639 19264 -1628
rect 19135 -1703 19166 -1639
rect 19230 -1703 19264 -1639
rect 19135 -1714 19264 -1703
rect 19355 -1636 19484 -1625
rect 19355 -1700 19386 -1636
rect 19450 -1700 19484 -1636
rect 19355 -1711 19484 -1700
rect 19570 -1640 19699 -1629
rect 19570 -1704 19601 -1640
rect 19665 -1704 19699 -1640
rect 19570 -1715 19699 -1704
rect 19798 -1637 19927 -1626
rect 19798 -1701 19829 -1637
rect 19893 -1701 19927 -1637
rect 19798 -1712 19927 -1701
rect 20002 -1640 20131 -1629
rect 20002 -1704 20033 -1640
rect 20097 -1704 20131 -1640
rect 20002 -1715 20131 -1704
rect 20240 -1638 20369 -1627
rect 20240 -1702 20271 -1638
rect 20335 -1702 20369 -1638
rect 20240 -1713 20369 -1702
rect 20433 -1637 20562 -1626
rect 20433 -1701 20464 -1637
rect 20528 -1701 20562 -1637
rect 20433 -1712 20562 -1701
rect 20630 -1642 20759 -1631
rect 20630 -1706 20661 -1642
rect 20725 -1706 20759 -1642
rect 20630 -1717 20759 -1706
rect 20886 -1639 21015 -1628
rect 20886 -1703 20917 -1639
rect 20981 -1703 21015 -1639
rect 20886 -1714 21015 -1703
rect 21125 -1643 21254 -1632
rect 21125 -1707 21156 -1643
rect 21220 -1707 21254 -1643
rect 21125 -1718 21254 -1707
rect 21358 -1647 21487 -1636
rect 21358 -1711 21389 -1647
rect 21453 -1711 21487 -1647
rect 21358 -1722 21487 -1711
rect 21579 -1642 21708 -1631
rect 21579 -1706 21610 -1642
rect 21674 -1706 21708 -1642
rect 21579 -1717 21708 -1706
rect 21770 -1642 21899 -1631
rect 21770 -1706 21801 -1642
rect 21865 -1706 21899 -1642
rect 21770 -1717 21899 -1706
rect 21998 -1640 22127 -1629
rect 21998 -1704 22029 -1640
rect 22093 -1704 22127 -1640
rect 21998 -1715 22127 -1704
rect 22195 -1645 22324 -1634
rect 22195 -1709 22226 -1645
rect 22290 -1709 22324 -1645
rect 22195 -1720 22324 -1709
rect 22407 -1645 22536 -1634
rect 22407 -1709 22438 -1645
rect 22502 -1709 22536 -1645
rect 22407 -1720 22536 -1709
rect 22634 -1642 22763 -1631
rect 22634 -1706 22665 -1642
rect 22729 -1706 22763 -1642
rect 22634 -1717 22763 -1706
rect 22823 -1641 22952 -1630
rect 22823 -1705 22854 -1641
rect 22918 -1705 22952 -1641
rect 22823 -1716 22952 -1705
rect 23049 -1640 23178 -1629
rect 23049 -1704 23080 -1640
rect 23144 -1704 23178 -1640
rect 23049 -1715 23178 -1704
rect 23303 -1640 23432 -1629
rect 23303 -1704 23334 -1640
rect 23398 -1704 23432 -1640
rect 23303 -1715 23432 -1704
rect 23547 -1643 23676 -1632
rect 23547 -1707 23578 -1643
rect 23642 -1707 23676 -1643
rect 23547 -1718 23676 -1707
rect 23777 -1644 23906 -1633
rect 23777 -1708 23808 -1644
rect 23872 -1708 23906 -1644
rect 23777 -1719 23906 -1708
rect 24035 -1641 24164 -1630
rect 24035 -1705 24066 -1641
rect 24130 -1705 24164 -1641
rect 24035 -1716 24164 -1705
rect 24245 -1641 24374 -1630
rect 24245 -1705 24276 -1641
rect 24340 -1705 24374 -1641
rect 24245 -1716 24374 -1705
rect 24470 -1641 24599 -1630
rect 24470 -1705 24501 -1641
rect 24565 -1705 24599 -1641
rect 24470 -1716 24599 -1705
rect 24689 -1644 24818 -1633
rect 24689 -1708 24720 -1644
rect 24784 -1708 24818 -1644
rect 24689 -1719 24818 -1708
rect 25035 -1640 25164 -1629
rect 25035 -1704 25066 -1640
rect 25130 -1704 25164 -1640
rect 25035 -1715 25164 -1704
rect 25234 -1643 25363 -1632
rect 25234 -1707 25265 -1643
rect 25329 -1707 25363 -1643
rect 25234 -1718 25363 -1707
<< via3 >>
rect 13950 13628 14014 13632
rect 13950 13572 13954 13628
rect 13954 13572 14010 13628
rect 14010 13572 14014 13628
rect 13950 13568 14014 13572
rect 14047 13619 14111 13622
rect 14047 13563 14050 13619
rect 14050 13563 14106 13619
rect 14106 13563 14111 13619
rect 14047 13558 14111 13563
rect 14127 13619 14191 13622
rect 14127 13563 14130 13619
rect 14130 13563 14186 13619
rect 14186 13563 14191 13619
rect 14127 13558 14191 13563
rect 14207 13619 14271 13622
rect 14207 13563 14210 13619
rect 14210 13563 14266 13619
rect 14266 13563 14271 13619
rect 14207 13558 14271 13563
rect 14287 13619 14351 13622
rect 14287 13563 14290 13619
rect 14290 13563 14346 13619
rect 14346 13563 14351 13619
rect 14287 13558 14351 13563
rect 14367 13619 14431 13622
rect 14367 13563 14370 13619
rect 14370 13563 14426 13619
rect 14426 13563 14431 13619
rect 14367 13558 14431 13563
rect 14447 13619 14511 13622
rect 14447 13563 14450 13619
rect 14450 13563 14506 13619
rect 14506 13563 14511 13619
rect 14447 13558 14511 13563
rect 14779 13622 14843 13625
rect 14779 13566 14782 13622
rect 14782 13566 14838 13622
rect 14838 13566 14843 13622
rect 14779 13561 14843 13566
rect 14859 13622 14923 13625
rect 14859 13566 14862 13622
rect 14862 13566 14918 13622
rect 14918 13566 14923 13622
rect 14859 13561 14923 13566
rect 14939 13622 15003 13625
rect 14939 13566 14942 13622
rect 14942 13566 14998 13622
rect 14998 13566 15003 13622
rect 14939 13561 15003 13566
rect 15019 13622 15083 13625
rect 15019 13566 15022 13622
rect 15022 13566 15078 13622
rect 15078 13566 15083 13622
rect 15019 13561 15083 13566
rect 15099 13622 15163 13625
rect 15099 13566 15102 13622
rect 15102 13566 15158 13622
rect 15158 13566 15163 13622
rect 15099 13561 15163 13566
rect 15179 13622 15243 13625
rect 15179 13566 15182 13622
rect 15182 13566 15238 13622
rect 15238 13566 15243 13622
rect 15179 13561 15243 13566
rect 15385 13622 15449 13625
rect 15385 13566 15390 13622
rect 15390 13566 15446 13622
rect 15446 13566 15449 13622
rect 15385 13561 15449 13566
rect 15465 13622 15529 13625
rect 15465 13566 15470 13622
rect 15470 13566 15526 13622
rect 15526 13566 15529 13622
rect 15465 13561 15529 13566
rect 15545 13622 15609 13625
rect 15545 13566 15550 13622
rect 15550 13566 15606 13622
rect 15606 13566 15609 13622
rect 15545 13561 15609 13566
rect 15625 13622 15689 13625
rect 15625 13566 15630 13622
rect 15630 13566 15686 13622
rect 15686 13566 15689 13622
rect 15625 13561 15689 13566
rect 15705 13622 15769 13625
rect 15705 13566 15710 13622
rect 15710 13566 15766 13622
rect 15766 13566 15769 13622
rect 15705 13561 15769 13566
rect 15785 13622 15849 13625
rect 15785 13566 15790 13622
rect 15790 13566 15846 13622
rect 15846 13566 15849 13622
rect 15785 13561 15849 13566
rect 15991 13622 16055 13625
rect 15991 13566 15994 13622
rect 15994 13566 16050 13622
rect 16050 13566 16055 13622
rect 15991 13561 16055 13566
rect 16071 13622 16135 13625
rect 16071 13566 16074 13622
rect 16074 13566 16130 13622
rect 16130 13566 16135 13622
rect 16071 13561 16135 13566
rect 16151 13622 16215 13625
rect 16151 13566 16154 13622
rect 16154 13566 16210 13622
rect 16210 13566 16215 13622
rect 16151 13561 16215 13566
rect 16231 13622 16295 13625
rect 16231 13566 16234 13622
rect 16234 13566 16290 13622
rect 16290 13566 16295 13622
rect 16231 13561 16295 13566
rect 16311 13622 16375 13625
rect 16311 13566 16314 13622
rect 16314 13566 16370 13622
rect 16370 13566 16375 13622
rect 16311 13561 16375 13566
rect 16391 13622 16455 13625
rect 16391 13566 16394 13622
rect 16394 13566 16450 13622
rect 16450 13566 16455 13622
rect 16391 13561 16455 13566
rect 16597 13622 16661 13625
rect 16597 13566 16602 13622
rect 16602 13566 16658 13622
rect 16658 13566 16661 13622
rect 16597 13561 16661 13566
rect 16677 13622 16741 13625
rect 16677 13566 16682 13622
rect 16682 13566 16738 13622
rect 16738 13566 16741 13622
rect 16677 13561 16741 13566
rect 16757 13622 16821 13625
rect 16757 13566 16762 13622
rect 16762 13566 16818 13622
rect 16818 13566 16821 13622
rect 16757 13561 16821 13566
rect 16837 13622 16901 13625
rect 16837 13566 16842 13622
rect 16842 13566 16898 13622
rect 16898 13566 16901 13622
rect 16837 13561 16901 13566
rect 16917 13622 16981 13625
rect 16917 13566 16922 13622
rect 16922 13566 16978 13622
rect 16978 13566 16981 13622
rect 16917 13561 16981 13566
rect 16997 13622 17061 13625
rect 16997 13566 17002 13622
rect 17002 13566 17058 13622
rect 17058 13566 17061 13622
rect 16997 13561 17061 13566
rect 17203 13622 17267 13625
rect 17203 13566 17206 13622
rect 17206 13566 17262 13622
rect 17262 13566 17267 13622
rect 17203 13561 17267 13566
rect 17283 13622 17347 13625
rect 17283 13566 17286 13622
rect 17286 13566 17342 13622
rect 17342 13566 17347 13622
rect 17283 13561 17347 13566
rect 17363 13622 17427 13625
rect 17363 13566 17366 13622
rect 17366 13566 17422 13622
rect 17422 13566 17427 13622
rect 17363 13561 17427 13566
rect 17443 13622 17507 13625
rect 17443 13566 17446 13622
rect 17446 13566 17502 13622
rect 17502 13566 17507 13622
rect 17443 13561 17507 13566
rect 17523 13622 17587 13625
rect 17523 13566 17526 13622
rect 17526 13566 17582 13622
rect 17582 13566 17587 13622
rect 17523 13561 17587 13566
rect 17603 13622 17667 13625
rect 17603 13566 17606 13622
rect 17606 13566 17662 13622
rect 17662 13566 17667 13622
rect 17603 13561 17667 13566
rect 17809 13622 17873 13625
rect 17809 13566 17814 13622
rect 17814 13566 17870 13622
rect 17870 13566 17873 13622
rect 17809 13561 17873 13566
rect 17889 13622 17953 13625
rect 17889 13566 17894 13622
rect 17894 13566 17950 13622
rect 17950 13566 17953 13622
rect 17889 13561 17953 13566
rect 17969 13622 18033 13625
rect 17969 13566 17974 13622
rect 17974 13566 18030 13622
rect 18030 13566 18033 13622
rect 17969 13561 18033 13566
rect 18049 13622 18113 13625
rect 18049 13566 18054 13622
rect 18054 13566 18110 13622
rect 18110 13566 18113 13622
rect 18049 13561 18113 13566
rect 18129 13622 18193 13625
rect 18129 13566 18134 13622
rect 18134 13566 18190 13622
rect 18190 13566 18193 13622
rect 18129 13561 18193 13566
rect 18209 13622 18273 13625
rect 18209 13566 18214 13622
rect 18214 13566 18270 13622
rect 18270 13566 18273 13622
rect 18209 13561 18273 13566
rect 18415 13622 18479 13625
rect 18415 13566 18418 13622
rect 18418 13566 18474 13622
rect 18474 13566 18479 13622
rect 18415 13561 18479 13566
rect 18495 13622 18559 13625
rect 18495 13566 18498 13622
rect 18498 13566 18554 13622
rect 18554 13566 18559 13622
rect 18495 13561 18559 13566
rect 18575 13622 18639 13625
rect 18575 13566 18578 13622
rect 18578 13566 18634 13622
rect 18634 13566 18639 13622
rect 18575 13561 18639 13566
rect 18655 13622 18719 13625
rect 18655 13566 18658 13622
rect 18658 13566 18714 13622
rect 18714 13566 18719 13622
rect 18655 13561 18719 13566
rect 18735 13622 18799 13625
rect 18735 13566 18738 13622
rect 18738 13566 18794 13622
rect 18794 13566 18799 13622
rect 18735 13561 18799 13566
rect 18815 13622 18879 13625
rect 18815 13566 18818 13622
rect 18818 13566 18874 13622
rect 18874 13566 18879 13622
rect 18815 13561 18879 13566
rect 19021 13622 19085 13625
rect 19021 13566 19026 13622
rect 19026 13566 19082 13622
rect 19082 13566 19085 13622
rect 19021 13561 19085 13566
rect 19101 13622 19165 13625
rect 19101 13566 19106 13622
rect 19106 13566 19162 13622
rect 19162 13566 19165 13622
rect 19101 13561 19165 13566
rect 19181 13622 19245 13625
rect 19181 13566 19186 13622
rect 19186 13566 19242 13622
rect 19242 13566 19245 13622
rect 19181 13561 19245 13566
rect 19261 13622 19325 13625
rect 19261 13566 19266 13622
rect 19266 13566 19322 13622
rect 19322 13566 19325 13622
rect 19261 13561 19325 13566
rect 19341 13622 19405 13625
rect 19341 13566 19346 13622
rect 19346 13566 19402 13622
rect 19402 13566 19405 13622
rect 19341 13561 19405 13566
rect 19421 13622 19485 13625
rect 19421 13566 19426 13622
rect 19426 13566 19482 13622
rect 19482 13566 19485 13622
rect 19421 13561 19485 13566
rect 13944 13338 14008 13402
rect 13944 13258 14008 13322
rect 13944 13178 14008 13242
rect 3062 13153 3126 13157
rect 3062 13097 3066 13153
rect 3066 13097 3122 13153
rect 3122 13097 3126 13153
rect 3062 13093 3126 13097
rect 3159 13144 3223 13147
rect 3159 13088 3162 13144
rect 3162 13088 3218 13144
rect 3218 13088 3223 13144
rect 3159 13083 3223 13088
rect 3239 13144 3303 13147
rect 3239 13088 3242 13144
rect 3242 13088 3298 13144
rect 3298 13088 3303 13144
rect 3239 13083 3303 13088
rect 3319 13144 3383 13147
rect 3319 13088 3322 13144
rect 3322 13088 3378 13144
rect 3378 13088 3383 13144
rect 3319 13083 3383 13088
rect 3399 13144 3463 13147
rect 3399 13088 3402 13144
rect 3402 13088 3458 13144
rect 3458 13088 3463 13144
rect 3399 13083 3463 13088
rect 3479 13144 3543 13147
rect 3479 13088 3482 13144
rect 3482 13088 3538 13144
rect 3538 13088 3543 13144
rect 3479 13083 3543 13088
rect 3559 13144 3623 13147
rect 3559 13088 3562 13144
rect 3562 13088 3618 13144
rect 3618 13088 3623 13144
rect 3559 13083 3623 13088
rect 3891 13147 3955 13150
rect 3891 13091 3894 13147
rect 3894 13091 3950 13147
rect 3950 13091 3955 13147
rect 3891 13086 3955 13091
rect 3971 13147 4035 13150
rect 3971 13091 3974 13147
rect 3974 13091 4030 13147
rect 4030 13091 4035 13147
rect 3971 13086 4035 13091
rect 4051 13147 4115 13150
rect 4051 13091 4054 13147
rect 4054 13091 4110 13147
rect 4110 13091 4115 13147
rect 4051 13086 4115 13091
rect 4131 13147 4195 13150
rect 4131 13091 4134 13147
rect 4134 13091 4190 13147
rect 4190 13091 4195 13147
rect 4131 13086 4195 13091
rect 4211 13147 4275 13150
rect 4211 13091 4214 13147
rect 4214 13091 4270 13147
rect 4270 13091 4275 13147
rect 4211 13086 4275 13091
rect 4291 13147 4355 13150
rect 4291 13091 4294 13147
rect 4294 13091 4350 13147
rect 4350 13091 4355 13147
rect 4291 13086 4355 13091
rect 4497 13147 4561 13150
rect 4497 13091 4502 13147
rect 4502 13091 4558 13147
rect 4558 13091 4561 13147
rect 4497 13086 4561 13091
rect 4577 13147 4641 13150
rect 4577 13091 4582 13147
rect 4582 13091 4638 13147
rect 4638 13091 4641 13147
rect 4577 13086 4641 13091
rect 4657 13147 4721 13150
rect 4657 13091 4662 13147
rect 4662 13091 4718 13147
rect 4718 13091 4721 13147
rect 4657 13086 4721 13091
rect 4737 13147 4801 13150
rect 4737 13091 4742 13147
rect 4742 13091 4798 13147
rect 4798 13091 4801 13147
rect 4737 13086 4801 13091
rect 4817 13147 4881 13150
rect 4817 13091 4822 13147
rect 4822 13091 4878 13147
rect 4878 13091 4881 13147
rect 4817 13086 4881 13091
rect 4897 13147 4961 13150
rect 4897 13091 4902 13147
rect 4902 13091 4958 13147
rect 4958 13091 4961 13147
rect 4897 13086 4961 13091
rect 5103 13147 5167 13150
rect 5103 13091 5106 13147
rect 5106 13091 5162 13147
rect 5162 13091 5167 13147
rect 5103 13086 5167 13091
rect 5183 13147 5247 13150
rect 5183 13091 5186 13147
rect 5186 13091 5242 13147
rect 5242 13091 5247 13147
rect 5183 13086 5247 13091
rect 5263 13147 5327 13150
rect 5263 13091 5266 13147
rect 5266 13091 5322 13147
rect 5322 13091 5327 13147
rect 5263 13086 5327 13091
rect 5343 13147 5407 13150
rect 5343 13091 5346 13147
rect 5346 13091 5402 13147
rect 5402 13091 5407 13147
rect 5343 13086 5407 13091
rect 5423 13147 5487 13150
rect 5423 13091 5426 13147
rect 5426 13091 5482 13147
rect 5482 13091 5487 13147
rect 5423 13086 5487 13091
rect 5503 13147 5567 13150
rect 5503 13091 5506 13147
rect 5506 13091 5562 13147
rect 5562 13091 5567 13147
rect 5503 13086 5567 13091
rect 5709 13147 5773 13150
rect 5709 13091 5714 13147
rect 5714 13091 5770 13147
rect 5770 13091 5773 13147
rect 5709 13086 5773 13091
rect 5789 13147 5853 13150
rect 5789 13091 5794 13147
rect 5794 13091 5850 13147
rect 5850 13091 5853 13147
rect 5789 13086 5853 13091
rect 5869 13147 5933 13150
rect 5869 13091 5874 13147
rect 5874 13091 5930 13147
rect 5930 13091 5933 13147
rect 5869 13086 5933 13091
rect 5949 13147 6013 13150
rect 5949 13091 5954 13147
rect 5954 13091 6010 13147
rect 6010 13091 6013 13147
rect 5949 13086 6013 13091
rect 6029 13147 6093 13150
rect 6029 13091 6034 13147
rect 6034 13091 6090 13147
rect 6090 13091 6093 13147
rect 6029 13086 6093 13091
rect 6109 13147 6173 13150
rect 6109 13091 6114 13147
rect 6114 13091 6170 13147
rect 6170 13091 6173 13147
rect 6109 13086 6173 13091
rect 6315 13147 6379 13150
rect 6315 13091 6318 13147
rect 6318 13091 6374 13147
rect 6374 13091 6379 13147
rect 6315 13086 6379 13091
rect 6395 13147 6459 13150
rect 6395 13091 6398 13147
rect 6398 13091 6454 13147
rect 6454 13091 6459 13147
rect 6395 13086 6459 13091
rect 6475 13147 6539 13150
rect 6475 13091 6478 13147
rect 6478 13091 6534 13147
rect 6534 13091 6539 13147
rect 6475 13086 6539 13091
rect 6555 13147 6619 13150
rect 6555 13091 6558 13147
rect 6558 13091 6614 13147
rect 6614 13091 6619 13147
rect 6555 13086 6619 13091
rect 6635 13147 6699 13150
rect 6635 13091 6638 13147
rect 6638 13091 6694 13147
rect 6694 13091 6699 13147
rect 6635 13086 6699 13091
rect 6715 13147 6779 13150
rect 6715 13091 6718 13147
rect 6718 13091 6774 13147
rect 6774 13091 6779 13147
rect 6715 13086 6779 13091
rect 6921 13147 6985 13150
rect 6921 13091 6926 13147
rect 6926 13091 6982 13147
rect 6982 13091 6985 13147
rect 6921 13086 6985 13091
rect 7001 13147 7065 13150
rect 7001 13091 7006 13147
rect 7006 13091 7062 13147
rect 7062 13091 7065 13147
rect 7001 13086 7065 13091
rect 7081 13147 7145 13150
rect 7081 13091 7086 13147
rect 7086 13091 7142 13147
rect 7142 13091 7145 13147
rect 7081 13086 7145 13091
rect 7161 13147 7225 13150
rect 7161 13091 7166 13147
rect 7166 13091 7222 13147
rect 7222 13091 7225 13147
rect 7161 13086 7225 13091
rect 7241 13147 7305 13150
rect 7241 13091 7246 13147
rect 7246 13091 7302 13147
rect 7302 13091 7305 13147
rect 7241 13086 7305 13091
rect 7321 13147 7385 13150
rect 7321 13091 7326 13147
rect 7326 13091 7382 13147
rect 7382 13091 7385 13147
rect 7321 13086 7385 13091
rect 7527 13147 7591 13150
rect 7527 13091 7530 13147
rect 7530 13091 7586 13147
rect 7586 13091 7591 13147
rect 7527 13086 7591 13091
rect 7607 13147 7671 13150
rect 7607 13091 7610 13147
rect 7610 13091 7666 13147
rect 7666 13091 7671 13147
rect 7607 13086 7671 13091
rect 7687 13147 7751 13150
rect 7687 13091 7690 13147
rect 7690 13091 7746 13147
rect 7746 13091 7751 13147
rect 7687 13086 7751 13091
rect 7767 13147 7831 13150
rect 7767 13091 7770 13147
rect 7770 13091 7826 13147
rect 7826 13091 7831 13147
rect 7767 13086 7831 13091
rect 7847 13147 7911 13150
rect 7847 13091 7850 13147
rect 7850 13091 7906 13147
rect 7906 13091 7911 13147
rect 7847 13086 7911 13091
rect 7927 13147 7991 13150
rect 7927 13091 7930 13147
rect 7930 13091 7986 13147
rect 7986 13091 7991 13147
rect 7927 13086 7991 13091
rect 8133 13147 8197 13150
rect 8133 13091 8138 13147
rect 8138 13091 8194 13147
rect 8194 13091 8197 13147
rect 8133 13086 8197 13091
rect 8213 13147 8277 13150
rect 8213 13091 8218 13147
rect 8218 13091 8274 13147
rect 8274 13091 8277 13147
rect 8213 13086 8277 13091
rect 8293 13147 8357 13150
rect 8293 13091 8298 13147
rect 8298 13091 8354 13147
rect 8354 13091 8357 13147
rect 8293 13086 8357 13091
rect 8373 13147 8437 13150
rect 8373 13091 8378 13147
rect 8378 13091 8434 13147
rect 8434 13091 8437 13147
rect 8373 13086 8437 13091
rect 8453 13147 8517 13150
rect 8453 13091 8458 13147
rect 8458 13091 8514 13147
rect 8514 13091 8517 13147
rect 8453 13086 8517 13091
rect 8533 13147 8597 13150
rect 8533 13091 8538 13147
rect 8538 13091 8594 13147
rect 8594 13091 8597 13147
rect 8533 13086 8597 13091
rect 3056 12863 3120 12927
rect 3056 12783 3120 12847
rect 3056 12703 3120 12767
rect 3056 12623 3120 12687
rect 2445 12548 2509 12552
rect 2445 12492 2449 12548
rect 2449 12492 2505 12548
rect 2505 12492 2509 12548
rect 2445 12488 2509 12492
rect 2576 12547 2640 12551
rect 2576 12491 2580 12547
rect 2580 12491 2636 12547
rect 2636 12491 2640 12547
rect 2576 12487 2640 12491
rect 2720 12548 2784 12552
rect 2720 12492 2724 12548
rect 2724 12492 2780 12548
rect 2780 12492 2784 12548
rect 2720 12488 2784 12492
rect 3056 12543 3120 12607
rect 3056 12463 3120 12527
rect 3056 12383 3120 12447
rect 3056 12303 3120 12367
rect 3056 12223 3120 12287
rect 3056 12143 3120 12207
rect 2463 12002 2527 12006
rect 2463 11946 2467 12002
rect 2467 11946 2523 12002
rect 2523 11946 2527 12002
rect 2463 11942 2527 11946
rect 2583 12002 2647 12006
rect 2583 11946 2587 12002
rect 2587 11946 2643 12002
rect 2643 11946 2647 12002
rect 2583 11942 2647 11946
rect 2726 12002 2790 12006
rect 2726 11946 2730 12002
rect 2730 11946 2786 12002
rect 2786 11946 2790 12002
rect 2726 11942 2790 11946
rect 3662 12863 3726 12927
rect 3662 12783 3726 12847
rect 3662 12703 3726 12767
rect 3662 12623 3726 12687
rect 3662 12543 3726 12607
rect 3662 12463 3726 12527
rect 3662 12383 3726 12447
rect 3662 12303 3726 12367
rect 3662 12223 3726 12287
rect 3662 12143 3726 12207
rect 3159 11923 3223 11987
rect 3239 11923 3303 11987
rect 3319 11923 3383 11987
rect 3399 11923 3463 11987
rect 3479 11923 3543 11987
rect 3559 11964 3623 11987
rect 3559 11923 3612 11964
rect 3612 11923 3623 11964
rect 3788 12866 3852 12930
rect 3788 12786 3852 12850
rect 3788 12706 3852 12770
rect 3788 12626 3852 12690
rect 3788 12546 3852 12610
rect 3788 12466 3852 12530
rect 3788 12386 3852 12450
rect 3788 12306 3852 12370
rect 3788 12226 3852 12290
rect 3788 12146 3852 12210
rect 4394 12866 4458 12930
rect 4394 12786 4458 12850
rect 4394 12706 4458 12770
rect 4394 12626 4458 12690
rect 4394 12546 4458 12610
rect 4394 12466 4458 12530
rect 4394 12386 4458 12450
rect 4394 12306 4458 12370
rect 4394 12226 4458 12290
rect 4394 12146 4458 12210
rect 5000 12866 5064 12930
rect 5000 12786 5064 12850
rect 5000 12706 5064 12770
rect 5000 12626 5064 12690
rect 5000 12546 5064 12610
rect 5000 12466 5064 12530
rect 5000 12386 5064 12450
rect 5000 12306 5064 12370
rect 5000 12226 5064 12290
rect 5000 12146 5064 12210
rect 5606 12866 5670 12930
rect 5606 12786 5670 12850
rect 5606 12706 5670 12770
rect 5606 12626 5670 12690
rect 5606 12546 5670 12610
rect 5606 12466 5670 12530
rect 5606 12386 5670 12450
rect 5606 12306 5670 12370
rect 5606 12226 5670 12290
rect 5606 12146 5670 12210
rect 6212 12866 6276 12930
rect 6212 12786 6276 12850
rect 6212 12706 6276 12770
rect 6212 12626 6276 12690
rect 6212 12546 6276 12610
rect 6212 12466 6276 12530
rect 6212 12386 6276 12450
rect 6212 12306 6276 12370
rect 6212 12226 6276 12290
rect 6212 12146 6276 12210
rect 6818 12866 6882 12930
rect 6818 12786 6882 12850
rect 6818 12706 6882 12770
rect 6818 12626 6882 12690
rect 6818 12546 6882 12610
rect 6818 12466 6882 12530
rect 6818 12386 6882 12450
rect 6818 12306 6882 12370
rect 6818 12226 6882 12290
rect 6818 12146 6882 12210
rect 7424 12866 7488 12930
rect 7424 12786 7488 12850
rect 7424 12706 7488 12770
rect 7424 12626 7488 12690
rect 7424 12546 7488 12610
rect 7424 12466 7488 12530
rect 7424 12386 7488 12450
rect 7424 12306 7488 12370
rect 7424 12226 7488 12290
rect 7424 12146 7488 12210
rect 8030 12866 8094 12930
rect 8030 12786 8094 12850
rect 8030 12706 8094 12770
rect 8030 12626 8094 12690
rect 8030 12546 8094 12610
rect 8030 12466 8094 12530
rect 8030 12386 8094 12450
rect 8030 12306 8094 12370
rect 8030 12226 8094 12290
rect 8030 12146 8094 12210
rect 8871 13091 8935 13095
rect 8871 13035 8875 13091
rect 8875 13035 8931 13091
rect 8931 13035 8935 13091
rect 8871 13031 8935 13035
rect 13944 13098 14008 13162
rect 13333 13023 13397 13027
rect 13333 12967 13337 13023
rect 13337 12967 13393 13023
rect 13393 12967 13397 13023
rect 13333 12963 13397 12967
rect 13464 13022 13528 13026
rect 13464 12966 13468 13022
rect 13468 12966 13524 13022
rect 13524 12966 13528 13022
rect 13464 12962 13528 12966
rect 13608 13023 13672 13027
rect 13608 12967 13612 13023
rect 13612 12967 13668 13023
rect 13668 12967 13672 13023
rect 13608 12963 13672 12967
rect 8636 12866 8700 12930
rect 8876 12947 8940 12951
rect 8876 12891 8880 12947
rect 8880 12891 8936 12947
rect 8936 12891 8940 12947
rect 8876 12887 8940 12891
rect 13944 13018 14008 13082
rect 13944 12938 14008 13002
rect 8636 12786 8700 12850
rect 13944 12858 14008 12922
rect 8636 12706 8700 12770
rect 8877 12795 8941 12799
rect 8877 12739 8881 12795
rect 8881 12739 8937 12795
rect 8937 12739 8941 12795
rect 8877 12735 8941 12739
rect 13944 12778 14008 12842
rect 8636 12626 8700 12690
rect 13944 12698 14008 12762
rect 8636 12546 8700 12610
rect 8877 12625 8941 12629
rect 8877 12569 8881 12625
rect 8881 12569 8937 12625
rect 8937 12569 8941 12625
rect 8877 12565 8941 12569
rect 13944 12618 14008 12682
rect 8636 12466 8700 12530
rect 10981 12556 11045 12560
rect 10981 12500 10985 12556
rect 10985 12500 11041 12556
rect 11041 12500 11045 12556
rect 10981 12496 11045 12500
rect 11168 12558 11232 12562
rect 11168 12502 11172 12558
rect 11172 12502 11228 12558
rect 11228 12502 11232 12558
rect 11168 12498 11232 12502
rect 11353 12560 11417 12564
rect 11353 12504 11357 12560
rect 11357 12504 11413 12560
rect 11413 12504 11417 12560
rect 11353 12500 11417 12504
rect 11538 12561 11602 12565
rect 11538 12505 11542 12561
rect 11542 12505 11598 12561
rect 11598 12505 11602 12561
rect 11538 12501 11602 12505
rect 11741 12563 11805 12567
rect 11741 12507 11745 12563
rect 11745 12507 11801 12563
rect 11801 12507 11805 12563
rect 11741 12503 11805 12507
rect 11926 12565 11990 12569
rect 11926 12509 11930 12565
rect 11930 12509 11986 12565
rect 11986 12509 11990 12565
rect 11926 12505 11990 12509
rect 12125 12567 12189 12571
rect 12125 12511 12129 12567
rect 12129 12511 12185 12567
rect 12185 12511 12189 12567
rect 12125 12507 12189 12511
rect 12327 12566 12391 12570
rect 12327 12510 12331 12566
rect 12331 12510 12387 12566
rect 12387 12510 12391 12566
rect 12327 12506 12391 12510
rect 12537 12569 12601 12573
rect 12537 12513 12541 12569
rect 12541 12513 12597 12569
rect 12597 12513 12601 12569
rect 12537 12509 12601 12513
rect 12761 12569 12825 12573
rect 12761 12513 12765 12569
rect 12765 12513 12821 12569
rect 12821 12513 12825 12569
rect 12761 12509 12825 12513
rect 12967 12568 13031 12572
rect 12967 12512 12971 12568
rect 12971 12512 13027 12568
rect 13027 12512 13031 12568
rect 12967 12508 13031 12512
rect 13188 12567 13252 12571
rect 13188 12511 13192 12567
rect 13192 12511 13248 12567
rect 13248 12511 13252 12567
rect 13188 12507 13252 12511
rect 8636 12386 8700 12450
rect 8876 12468 8940 12472
rect 8876 12412 8880 12468
rect 8880 12412 8936 12468
rect 8936 12412 8940 12468
rect 8876 12408 8940 12412
rect 13351 12477 13415 12481
rect 13351 12421 13355 12477
rect 13355 12421 13411 12477
rect 13411 12421 13415 12477
rect 13351 12417 13415 12421
rect 13471 12477 13535 12481
rect 13471 12421 13475 12477
rect 13475 12421 13531 12477
rect 13531 12421 13535 12477
rect 13471 12417 13535 12421
rect 13614 12477 13678 12481
rect 13614 12421 13618 12477
rect 13618 12421 13674 12477
rect 13674 12421 13678 12477
rect 13614 12417 13678 12421
rect 14550 13338 14614 13402
rect 14550 13258 14614 13322
rect 14550 13178 14614 13242
rect 14550 13098 14614 13162
rect 14550 13018 14614 13082
rect 14550 12938 14614 13002
rect 14550 12858 14614 12922
rect 14550 12778 14614 12842
rect 14550 12698 14614 12762
rect 14550 12618 14614 12682
rect 14047 12398 14111 12462
rect 14127 12398 14191 12462
rect 14207 12398 14271 12462
rect 14287 12398 14351 12462
rect 14367 12398 14431 12462
rect 14447 12439 14511 12462
rect 14447 12398 14500 12439
rect 14500 12398 14511 12439
rect 14676 13341 14740 13405
rect 14676 13261 14740 13325
rect 14676 13181 14740 13245
rect 14676 13101 14740 13165
rect 14676 13021 14740 13085
rect 14676 12941 14740 13005
rect 14676 12861 14740 12925
rect 14676 12781 14740 12845
rect 14676 12701 14740 12765
rect 14676 12621 14740 12685
rect 15282 13341 15346 13405
rect 15282 13261 15346 13325
rect 15282 13181 15346 13245
rect 15282 13101 15346 13165
rect 15282 13021 15346 13085
rect 15282 12941 15346 13005
rect 15282 12861 15346 12925
rect 15282 12781 15346 12845
rect 15282 12701 15346 12765
rect 15282 12621 15346 12685
rect 15888 13341 15952 13405
rect 15888 13261 15952 13325
rect 15888 13181 15952 13245
rect 15888 13101 15952 13165
rect 15888 13021 15952 13085
rect 15888 12941 15952 13005
rect 15888 12861 15952 12925
rect 15888 12781 15952 12845
rect 15888 12701 15952 12765
rect 15888 12621 15952 12685
rect 16494 13341 16558 13405
rect 16494 13261 16558 13325
rect 16494 13181 16558 13245
rect 16494 13101 16558 13165
rect 16494 13021 16558 13085
rect 16494 12941 16558 13005
rect 16494 12861 16558 12925
rect 16494 12781 16558 12845
rect 16494 12701 16558 12765
rect 16494 12621 16558 12685
rect 17100 13341 17164 13405
rect 17100 13261 17164 13325
rect 17100 13181 17164 13245
rect 17100 13101 17164 13165
rect 17100 13021 17164 13085
rect 17100 12941 17164 13005
rect 17100 12861 17164 12925
rect 17100 12781 17164 12845
rect 17100 12701 17164 12765
rect 17100 12621 17164 12685
rect 17706 13341 17770 13405
rect 17706 13261 17770 13325
rect 17706 13181 17770 13245
rect 17706 13101 17770 13165
rect 17706 13021 17770 13085
rect 17706 12941 17770 13005
rect 17706 12861 17770 12925
rect 17706 12781 17770 12845
rect 17706 12701 17770 12765
rect 17706 12621 17770 12685
rect 18312 13341 18376 13405
rect 18312 13261 18376 13325
rect 18312 13181 18376 13245
rect 18312 13101 18376 13165
rect 18312 13021 18376 13085
rect 18312 12941 18376 13005
rect 18312 12861 18376 12925
rect 18312 12781 18376 12845
rect 18312 12701 18376 12765
rect 18312 12621 18376 12685
rect 18918 13341 18982 13405
rect 18918 13261 18982 13325
rect 18918 13181 18982 13245
rect 18918 13101 18982 13165
rect 18918 13021 18982 13085
rect 18918 12941 18982 13005
rect 18918 12861 18982 12925
rect 18918 12781 18982 12845
rect 18918 12701 18982 12765
rect 18918 12621 18982 12685
rect 19759 13566 19823 13570
rect 19759 13510 19763 13566
rect 19763 13510 19819 13566
rect 19819 13510 19823 13566
rect 19759 13506 19823 13510
rect 20236 13569 20300 13573
rect 20236 13513 20240 13569
rect 20240 13513 20296 13569
rect 20296 13513 20300 13569
rect 20236 13509 20300 13513
rect 20659 13628 20723 13632
rect 20659 13572 20663 13628
rect 20663 13572 20719 13628
rect 20719 13572 20723 13628
rect 20659 13568 20723 13572
rect 20756 13619 20820 13622
rect 20756 13563 20759 13619
rect 20759 13563 20815 13619
rect 20815 13563 20820 13619
rect 20756 13558 20820 13563
rect 20836 13619 20900 13622
rect 20836 13563 20839 13619
rect 20839 13563 20895 13619
rect 20895 13563 20900 13619
rect 20836 13558 20900 13563
rect 20916 13619 20980 13622
rect 20916 13563 20919 13619
rect 20919 13563 20975 13619
rect 20975 13563 20980 13619
rect 20916 13558 20980 13563
rect 20996 13619 21060 13622
rect 20996 13563 20999 13619
rect 20999 13563 21055 13619
rect 21055 13563 21060 13619
rect 20996 13558 21060 13563
rect 21076 13619 21140 13622
rect 21076 13563 21079 13619
rect 21079 13563 21135 13619
rect 21135 13563 21140 13619
rect 21076 13558 21140 13563
rect 21156 13619 21220 13622
rect 21156 13563 21159 13619
rect 21159 13563 21215 13619
rect 21215 13563 21220 13619
rect 21156 13558 21220 13563
rect 21488 13622 21552 13625
rect 21488 13566 21491 13622
rect 21491 13566 21547 13622
rect 21547 13566 21552 13622
rect 21488 13561 21552 13566
rect 21568 13622 21632 13625
rect 21568 13566 21571 13622
rect 21571 13566 21627 13622
rect 21627 13566 21632 13622
rect 21568 13561 21632 13566
rect 21648 13622 21712 13625
rect 21648 13566 21651 13622
rect 21651 13566 21707 13622
rect 21707 13566 21712 13622
rect 21648 13561 21712 13566
rect 21728 13622 21792 13625
rect 21728 13566 21731 13622
rect 21731 13566 21787 13622
rect 21787 13566 21792 13622
rect 21728 13561 21792 13566
rect 21808 13622 21872 13625
rect 21808 13566 21811 13622
rect 21811 13566 21867 13622
rect 21867 13566 21872 13622
rect 21808 13561 21872 13566
rect 21888 13622 21952 13625
rect 21888 13566 21891 13622
rect 21891 13566 21947 13622
rect 21947 13566 21952 13622
rect 21888 13561 21952 13566
rect 22094 13622 22158 13625
rect 22094 13566 22099 13622
rect 22099 13566 22155 13622
rect 22155 13566 22158 13622
rect 22094 13561 22158 13566
rect 22174 13622 22238 13625
rect 22174 13566 22179 13622
rect 22179 13566 22235 13622
rect 22235 13566 22238 13622
rect 22174 13561 22238 13566
rect 22254 13622 22318 13625
rect 22254 13566 22259 13622
rect 22259 13566 22315 13622
rect 22315 13566 22318 13622
rect 22254 13561 22318 13566
rect 22334 13622 22398 13625
rect 22334 13566 22339 13622
rect 22339 13566 22395 13622
rect 22395 13566 22398 13622
rect 22334 13561 22398 13566
rect 22414 13622 22478 13625
rect 22414 13566 22419 13622
rect 22419 13566 22475 13622
rect 22475 13566 22478 13622
rect 22414 13561 22478 13566
rect 22494 13622 22558 13625
rect 22494 13566 22499 13622
rect 22499 13566 22555 13622
rect 22555 13566 22558 13622
rect 22494 13561 22558 13566
rect 22700 13622 22764 13625
rect 22700 13566 22703 13622
rect 22703 13566 22759 13622
rect 22759 13566 22764 13622
rect 22700 13561 22764 13566
rect 22780 13622 22844 13625
rect 22780 13566 22783 13622
rect 22783 13566 22839 13622
rect 22839 13566 22844 13622
rect 22780 13561 22844 13566
rect 22860 13622 22924 13625
rect 22860 13566 22863 13622
rect 22863 13566 22919 13622
rect 22919 13566 22924 13622
rect 22860 13561 22924 13566
rect 22940 13622 23004 13625
rect 22940 13566 22943 13622
rect 22943 13566 22999 13622
rect 22999 13566 23004 13622
rect 22940 13561 23004 13566
rect 23020 13622 23084 13625
rect 23020 13566 23023 13622
rect 23023 13566 23079 13622
rect 23079 13566 23084 13622
rect 23020 13561 23084 13566
rect 23100 13622 23164 13625
rect 23100 13566 23103 13622
rect 23103 13566 23159 13622
rect 23159 13566 23164 13622
rect 23100 13561 23164 13566
rect 23306 13622 23370 13625
rect 23306 13566 23311 13622
rect 23311 13566 23367 13622
rect 23367 13566 23370 13622
rect 23306 13561 23370 13566
rect 23386 13622 23450 13625
rect 23386 13566 23391 13622
rect 23391 13566 23447 13622
rect 23447 13566 23450 13622
rect 23386 13561 23450 13566
rect 23466 13622 23530 13625
rect 23466 13566 23471 13622
rect 23471 13566 23527 13622
rect 23527 13566 23530 13622
rect 23466 13561 23530 13566
rect 23546 13622 23610 13625
rect 23546 13566 23551 13622
rect 23551 13566 23607 13622
rect 23607 13566 23610 13622
rect 23546 13561 23610 13566
rect 23626 13622 23690 13625
rect 23626 13566 23631 13622
rect 23631 13566 23687 13622
rect 23687 13566 23690 13622
rect 23626 13561 23690 13566
rect 23706 13622 23770 13625
rect 23706 13566 23711 13622
rect 23711 13566 23767 13622
rect 23767 13566 23770 13622
rect 23706 13561 23770 13566
rect 23912 13622 23976 13625
rect 23912 13566 23915 13622
rect 23915 13566 23971 13622
rect 23971 13566 23976 13622
rect 23912 13561 23976 13566
rect 23992 13622 24056 13625
rect 23992 13566 23995 13622
rect 23995 13566 24051 13622
rect 24051 13566 24056 13622
rect 23992 13561 24056 13566
rect 24072 13622 24136 13625
rect 24072 13566 24075 13622
rect 24075 13566 24131 13622
rect 24131 13566 24136 13622
rect 24072 13561 24136 13566
rect 24152 13622 24216 13625
rect 24152 13566 24155 13622
rect 24155 13566 24211 13622
rect 24211 13566 24216 13622
rect 24152 13561 24216 13566
rect 24232 13622 24296 13625
rect 24232 13566 24235 13622
rect 24235 13566 24291 13622
rect 24291 13566 24296 13622
rect 24232 13561 24296 13566
rect 24312 13622 24376 13625
rect 24312 13566 24315 13622
rect 24315 13566 24371 13622
rect 24371 13566 24376 13622
rect 24312 13561 24376 13566
rect 24518 13622 24582 13625
rect 24518 13566 24523 13622
rect 24523 13566 24579 13622
rect 24579 13566 24582 13622
rect 24518 13561 24582 13566
rect 24598 13622 24662 13625
rect 24598 13566 24603 13622
rect 24603 13566 24659 13622
rect 24659 13566 24662 13622
rect 24598 13561 24662 13566
rect 24678 13622 24742 13625
rect 24678 13566 24683 13622
rect 24683 13566 24739 13622
rect 24739 13566 24742 13622
rect 24678 13561 24742 13566
rect 24758 13622 24822 13625
rect 24758 13566 24763 13622
rect 24763 13566 24819 13622
rect 24819 13566 24822 13622
rect 24758 13561 24822 13566
rect 24838 13622 24902 13625
rect 24838 13566 24843 13622
rect 24843 13566 24899 13622
rect 24899 13566 24902 13622
rect 24838 13561 24902 13566
rect 24918 13622 24982 13625
rect 24918 13566 24923 13622
rect 24923 13566 24979 13622
rect 24979 13566 24982 13622
rect 24918 13561 24982 13566
rect 25124 13622 25188 13625
rect 25124 13566 25127 13622
rect 25127 13566 25183 13622
rect 25183 13566 25188 13622
rect 25124 13561 25188 13566
rect 25204 13622 25268 13625
rect 25204 13566 25207 13622
rect 25207 13566 25263 13622
rect 25263 13566 25268 13622
rect 25204 13561 25268 13566
rect 25284 13622 25348 13625
rect 25284 13566 25287 13622
rect 25287 13566 25343 13622
rect 25343 13566 25348 13622
rect 25284 13561 25348 13566
rect 25364 13622 25428 13625
rect 25364 13566 25367 13622
rect 25367 13566 25423 13622
rect 25423 13566 25428 13622
rect 25364 13561 25428 13566
rect 25444 13622 25508 13625
rect 25444 13566 25447 13622
rect 25447 13566 25503 13622
rect 25503 13566 25508 13622
rect 25444 13561 25508 13566
rect 25524 13622 25588 13625
rect 25524 13566 25527 13622
rect 25527 13566 25583 13622
rect 25583 13566 25588 13622
rect 25524 13561 25588 13566
rect 25730 13622 25794 13625
rect 25730 13566 25735 13622
rect 25735 13566 25791 13622
rect 25791 13566 25794 13622
rect 25730 13561 25794 13566
rect 25810 13622 25874 13625
rect 25810 13566 25815 13622
rect 25815 13566 25871 13622
rect 25871 13566 25874 13622
rect 25810 13561 25874 13566
rect 25890 13622 25954 13625
rect 25890 13566 25895 13622
rect 25895 13566 25951 13622
rect 25951 13566 25954 13622
rect 25890 13561 25954 13566
rect 25970 13622 26034 13625
rect 25970 13566 25975 13622
rect 25975 13566 26031 13622
rect 26031 13566 26034 13622
rect 25970 13561 26034 13566
rect 26050 13622 26114 13625
rect 26050 13566 26055 13622
rect 26055 13566 26111 13622
rect 26111 13566 26114 13622
rect 26050 13561 26114 13566
rect 26130 13622 26194 13625
rect 26130 13566 26135 13622
rect 26135 13566 26191 13622
rect 26191 13566 26194 13622
rect 26130 13561 26194 13566
rect 19524 13341 19588 13405
rect 19764 13422 19828 13426
rect 19764 13366 19768 13422
rect 19768 13366 19824 13422
rect 19824 13366 19828 13422
rect 19764 13362 19828 13366
rect 20225 13397 20289 13401
rect 20225 13341 20229 13397
rect 20229 13341 20285 13397
rect 20285 13341 20289 13397
rect 20225 13337 20289 13341
rect 20653 13338 20717 13402
rect 19524 13261 19588 13325
rect 19524 13181 19588 13245
rect 19765 13270 19829 13274
rect 19765 13214 19769 13270
rect 19769 13214 19825 13270
rect 19825 13214 19829 13270
rect 19765 13210 19829 13214
rect 20653 13258 20717 13322
rect 19524 13101 19588 13165
rect 20225 13205 20289 13209
rect 20225 13149 20229 13205
rect 20229 13149 20285 13205
rect 20285 13149 20289 13205
rect 20225 13145 20289 13149
rect 20653 13178 20717 13242
rect 19524 13021 19588 13085
rect 19765 13100 19829 13104
rect 19765 13044 19769 13100
rect 19769 13044 19825 13100
rect 19825 13044 19829 13100
rect 19765 13040 19829 13044
rect 20653 13098 20717 13162
rect 19524 12941 19588 13005
rect 20042 13023 20106 13027
rect 20042 12967 20046 13023
rect 20046 12967 20102 13023
rect 20102 12967 20106 13023
rect 20042 12963 20106 12967
rect 20173 13022 20237 13026
rect 20173 12966 20177 13022
rect 20177 12966 20233 13022
rect 20233 12966 20237 13022
rect 20173 12962 20237 12966
rect 20317 13023 20381 13027
rect 20317 12967 20321 13023
rect 20321 12967 20377 13023
rect 20377 12967 20381 13023
rect 20317 12963 20381 12967
rect 19524 12861 19588 12925
rect 19764 12943 19828 12947
rect 19764 12887 19768 12943
rect 19768 12887 19824 12943
rect 19824 12887 19828 12943
rect 19764 12883 19828 12887
rect 20653 13018 20717 13082
rect 20653 12938 20717 13002
rect 19524 12781 19588 12845
rect 19524 12701 19588 12765
rect 20653 12858 20717 12922
rect 20653 12778 20717 12842
rect 19524 12621 19588 12685
rect 19682 12701 19746 12705
rect 19682 12645 19686 12701
rect 19686 12645 19742 12701
rect 19742 12645 19746 12701
rect 19682 12641 19746 12645
rect 20653 12698 20717 12762
rect 20653 12618 20717 12682
rect 14779 12401 14843 12465
rect 14859 12401 14923 12465
rect 14939 12401 15003 12465
rect 15019 12401 15083 12465
rect 15099 12401 15163 12465
rect 15179 12442 15243 12465
rect 15179 12401 15232 12442
rect 15232 12401 15243 12442
rect 15385 12442 15449 12465
rect 15385 12401 15396 12442
rect 15396 12401 15449 12442
rect 15465 12401 15529 12465
rect 15545 12401 15609 12465
rect 15625 12401 15689 12465
rect 15705 12401 15769 12465
rect 15785 12401 15849 12465
rect 15991 12401 16055 12465
rect 16071 12401 16135 12465
rect 16151 12401 16215 12465
rect 16231 12401 16295 12465
rect 16311 12401 16375 12465
rect 16391 12442 16455 12465
rect 16391 12401 16444 12442
rect 16444 12401 16455 12442
rect 16597 12442 16661 12465
rect 16597 12401 16608 12442
rect 16608 12401 16661 12442
rect 16677 12401 16741 12465
rect 16757 12401 16821 12465
rect 16837 12401 16901 12465
rect 16917 12401 16981 12465
rect 16997 12401 17061 12465
rect 17203 12401 17267 12465
rect 17283 12401 17347 12465
rect 17363 12401 17427 12465
rect 17443 12401 17507 12465
rect 17523 12401 17587 12465
rect 17603 12442 17667 12465
rect 17603 12401 17656 12442
rect 17656 12401 17667 12442
rect 17809 12442 17873 12465
rect 17809 12401 17820 12442
rect 17820 12401 17873 12442
rect 17889 12401 17953 12465
rect 17969 12401 18033 12465
rect 18049 12401 18113 12465
rect 18129 12401 18193 12465
rect 18209 12401 18273 12465
rect 18415 12401 18479 12465
rect 18495 12401 18559 12465
rect 18575 12401 18639 12465
rect 18655 12401 18719 12465
rect 18735 12401 18799 12465
rect 18815 12442 18879 12465
rect 18815 12401 18868 12442
rect 18868 12401 18879 12442
rect 19021 12442 19085 12465
rect 19021 12401 19032 12442
rect 19032 12401 19085 12442
rect 19101 12401 19165 12465
rect 19181 12401 19245 12465
rect 19261 12401 19325 12465
rect 19341 12401 19405 12465
rect 19421 12401 19485 12465
rect 19770 12440 19834 12444
rect 19770 12384 19774 12440
rect 19774 12384 19830 12440
rect 19830 12384 19834 12440
rect 19770 12380 19834 12384
rect 20060 12477 20124 12481
rect 20060 12421 20064 12477
rect 20064 12421 20120 12477
rect 20120 12421 20124 12477
rect 20060 12417 20124 12421
rect 20180 12477 20244 12481
rect 20180 12421 20184 12477
rect 20184 12421 20240 12477
rect 20240 12421 20244 12477
rect 20180 12417 20244 12421
rect 20323 12477 20387 12481
rect 20323 12421 20327 12477
rect 20327 12421 20383 12477
rect 20383 12421 20387 12477
rect 20323 12417 20387 12421
rect 21259 13338 21323 13402
rect 21259 13258 21323 13322
rect 21259 13178 21323 13242
rect 21259 13098 21323 13162
rect 21259 13018 21323 13082
rect 21259 12938 21323 13002
rect 21259 12858 21323 12922
rect 21259 12778 21323 12842
rect 21259 12698 21323 12762
rect 21259 12618 21323 12682
rect 20756 12398 20820 12462
rect 20836 12398 20900 12462
rect 20916 12398 20980 12462
rect 20996 12398 21060 12462
rect 21076 12398 21140 12462
rect 21156 12439 21220 12462
rect 21156 12398 21209 12439
rect 21209 12398 21220 12439
rect 21385 13341 21449 13405
rect 21385 13261 21449 13325
rect 21385 13181 21449 13245
rect 21385 13101 21449 13165
rect 21385 13021 21449 13085
rect 21385 12941 21449 13005
rect 21385 12861 21449 12925
rect 21385 12781 21449 12845
rect 21385 12701 21449 12765
rect 21385 12621 21449 12685
rect 21991 13341 22055 13405
rect 21991 13261 22055 13325
rect 21991 13181 22055 13245
rect 21991 13101 22055 13165
rect 21991 13021 22055 13085
rect 21991 12941 22055 13005
rect 21991 12861 22055 12925
rect 21991 12781 22055 12845
rect 21991 12701 22055 12765
rect 21991 12621 22055 12685
rect 22597 13341 22661 13405
rect 22597 13261 22661 13325
rect 22597 13181 22661 13245
rect 22597 13101 22661 13165
rect 22597 13021 22661 13085
rect 22597 12941 22661 13005
rect 22597 12861 22661 12925
rect 22597 12781 22661 12845
rect 22597 12701 22661 12765
rect 22597 12621 22661 12685
rect 23203 13341 23267 13405
rect 23203 13261 23267 13325
rect 23203 13181 23267 13245
rect 23203 13101 23267 13165
rect 23203 13021 23267 13085
rect 23203 12941 23267 13005
rect 23203 12861 23267 12925
rect 23203 12781 23267 12845
rect 23203 12701 23267 12765
rect 23203 12621 23267 12685
rect 23809 13341 23873 13405
rect 23809 13261 23873 13325
rect 23809 13181 23873 13245
rect 23809 13101 23873 13165
rect 23809 13021 23873 13085
rect 23809 12941 23873 13005
rect 23809 12861 23873 12925
rect 23809 12781 23873 12845
rect 23809 12701 23873 12765
rect 23809 12621 23873 12685
rect 24415 13341 24479 13405
rect 24415 13261 24479 13325
rect 24415 13181 24479 13245
rect 24415 13101 24479 13165
rect 24415 13021 24479 13085
rect 24415 12941 24479 13005
rect 24415 12861 24479 12925
rect 24415 12781 24479 12845
rect 24415 12701 24479 12765
rect 24415 12621 24479 12685
rect 25021 13341 25085 13405
rect 25021 13261 25085 13325
rect 25021 13181 25085 13245
rect 25021 13101 25085 13165
rect 25021 13021 25085 13085
rect 25021 12941 25085 13005
rect 25021 12861 25085 12925
rect 25021 12781 25085 12845
rect 25021 12701 25085 12765
rect 25021 12621 25085 12685
rect 25627 13341 25691 13405
rect 25627 13261 25691 13325
rect 25627 13181 25691 13245
rect 25627 13101 25691 13165
rect 25627 13021 25691 13085
rect 25627 12941 25691 13005
rect 25627 12861 25691 12925
rect 25627 12781 25691 12845
rect 25627 12701 25691 12765
rect 25627 12621 25691 12685
rect 26468 13566 26532 13570
rect 26468 13510 26472 13566
rect 26472 13510 26528 13566
rect 26528 13510 26532 13566
rect 26468 13506 26532 13510
rect 26233 13341 26297 13405
rect 26473 13422 26537 13426
rect 26473 13366 26477 13422
rect 26477 13366 26533 13422
rect 26533 13366 26537 13422
rect 26473 13362 26537 13366
rect 26233 13261 26297 13325
rect 26233 13181 26297 13245
rect 26474 13270 26538 13274
rect 26474 13214 26478 13270
rect 26478 13214 26534 13270
rect 26534 13214 26538 13270
rect 26474 13210 26538 13214
rect 26233 13101 26297 13165
rect 26233 13021 26297 13085
rect 26474 13100 26538 13104
rect 26474 13044 26478 13100
rect 26478 13044 26534 13100
rect 26534 13044 26538 13100
rect 26474 13040 26538 13044
rect 26233 12941 26297 13005
rect 26233 12861 26297 12925
rect 26473 12943 26537 12947
rect 26473 12887 26477 12943
rect 26477 12887 26533 12943
rect 26533 12887 26537 12943
rect 26473 12883 26537 12887
rect 26233 12781 26297 12845
rect 26233 12701 26297 12765
rect 26233 12621 26297 12685
rect 26391 12701 26455 12705
rect 26391 12645 26395 12701
rect 26395 12645 26451 12701
rect 26451 12645 26455 12701
rect 26391 12641 26455 12645
rect 21488 12401 21552 12465
rect 21568 12401 21632 12465
rect 21648 12401 21712 12465
rect 21728 12401 21792 12465
rect 21808 12401 21872 12465
rect 21888 12442 21952 12465
rect 21888 12401 21941 12442
rect 21941 12401 21952 12442
rect 22094 12442 22158 12465
rect 22094 12401 22105 12442
rect 22105 12401 22158 12442
rect 22174 12401 22238 12465
rect 22254 12401 22318 12465
rect 22334 12401 22398 12465
rect 22414 12401 22478 12465
rect 22494 12401 22558 12465
rect 22700 12401 22764 12465
rect 22780 12401 22844 12465
rect 22860 12401 22924 12465
rect 22940 12401 23004 12465
rect 23020 12401 23084 12465
rect 23100 12442 23164 12465
rect 23100 12401 23153 12442
rect 23153 12401 23164 12442
rect 23306 12442 23370 12465
rect 23306 12401 23317 12442
rect 23317 12401 23370 12442
rect 23386 12401 23450 12465
rect 23466 12401 23530 12465
rect 23546 12401 23610 12465
rect 23626 12401 23690 12465
rect 23706 12401 23770 12465
rect 23912 12401 23976 12465
rect 23992 12401 24056 12465
rect 24072 12401 24136 12465
rect 24152 12401 24216 12465
rect 24232 12401 24296 12465
rect 24312 12442 24376 12465
rect 24312 12401 24365 12442
rect 24365 12401 24376 12442
rect 24518 12442 24582 12465
rect 24518 12401 24529 12442
rect 24529 12401 24582 12442
rect 24598 12401 24662 12465
rect 24678 12401 24742 12465
rect 24758 12401 24822 12465
rect 24838 12401 24902 12465
rect 24918 12401 24982 12465
rect 25124 12401 25188 12465
rect 25204 12401 25268 12465
rect 25284 12401 25348 12465
rect 25364 12401 25428 12465
rect 25444 12401 25508 12465
rect 25524 12442 25588 12465
rect 25524 12401 25577 12442
rect 25577 12401 25588 12442
rect 25730 12442 25794 12465
rect 25730 12401 25741 12442
rect 25741 12401 25794 12442
rect 25810 12401 25874 12465
rect 25890 12401 25954 12465
rect 25970 12401 26034 12465
rect 26050 12401 26114 12465
rect 26130 12401 26194 12465
rect 26479 12440 26543 12444
rect 26479 12384 26483 12440
rect 26483 12384 26539 12440
rect 26539 12384 26543 12440
rect 26479 12380 26543 12384
rect 8636 12306 8700 12370
rect 8636 12226 8700 12290
rect 8636 12146 8700 12210
rect 8794 12226 8858 12230
rect 8794 12170 8798 12226
rect 8798 12170 8854 12226
rect 8854 12170 8858 12226
rect 8794 12166 8858 12170
rect 9171 12278 9235 12282
rect 9171 12222 9175 12278
rect 9175 12222 9231 12278
rect 9231 12222 9235 12278
rect 9171 12218 9235 12222
rect 3891 11926 3955 11990
rect 3971 11926 4035 11990
rect 4051 11926 4115 11990
rect 4131 11926 4195 11990
rect 4211 11926 4275 11990
rect 4291 11967 4355 11990
rect 4291 11926 4344 11967
rect 4344 11926 4355 11967
rect 4497 11967 4561 11990
rect 4497 11926 4508 11967
rect 4508 11926 4561 11967
rect 4577 11926 4641 11990
rect 4657 11926 4721 11990
rect 4737 11926 4801 11990
rect 4817 11926 4881 11990
rect 4897 11926 4961 11990
rect 5103 11926 5167 11990
rect 5183 11926 5247 11990
rect 5263 11926 5327 11990
rect 5343 11926 5407 11990
rect 5423 11926 5487 11990
rect 5503 11967 5567 11990
rect 5503 11926 5556 11967
rect 5556 11926 5567 11967
rect 5709 11967 5773 11990
rect 5709 11926 5720 11967
rect 5720 11926 5773 11967
rect 5789 11926 5853 11990
rect 5869 11926 5933 11990
rect 5949 11926 6013 11990
rect 6029 11926 6093 11990
rect 6109 11926 6173 11990
rect 6315 11926 6379 11990
rect 6395 11926 6459 11990
rect 6475 11926 6539 11990
rect 6555 11926 6619 11990
rect 6635 11926 6699 11990
rect 6715 11967 6779 11990
rect 6715 11926 6768 11967
rect 6768 11926 6779 11967
rect 6921 11967 6985 11990
rect 6921 11926 6932 11967
rect 6932 11926 6985 11967
rect 7001 11926 7065 11990
rect 7081 11926 7145 11990
rect 7161 11926 7225 11990
rect 7241 11926 7305 11990
rect 7321 11926 7385 11990
rect 7527 11926 7591 11990
rect 7607 11926 7671 11990
rect 7687 11926 7751 11990
rect 7767 11926 7831 11990
rect 7847 11926 7911 11990
rect 7927 11967 7991 11990
rect 7927 11926 7980 11967
rect 7980 11926 7991 11967
rect 8133 11967 8197 11990
rect 8133 11926 8144 11967
rect 8144 11926 8197 11967
rect 8213 11926 8277 11990
rect 8293 11926 8357 11990
rect 8373 11926 8437 11990
rect 8453 11926 8517 11990
rect 8533 11926 8597 11990
rect 14398 12153 14462 12217
rect 14478 12153 14542 12217
rect 14558 12153 14622 12217
rect 14638 12153 14702 12217
rect 14718 12153 14782 12217
rect 14798 12176 14856 12217
rect 14856 12176 14862 12217
rect 14798 12153 14862 12176
rect 8882 11965 8946 11969
rect 8882 11909 8886 11965
rect 8886 11909 8942 11965
rect 8942 11909 8946 11965
rect 8882 11905 8946 11909
rect 14295 11933 14359 11997
rect 10913 11883 10977 11885
rect 10913 11827 10916 11883
rect 10916 11827 10972 11883
rect 10972 11827 10977 11883
rect 10913 11821 10977 11827
rect 11113 11886 11177 11888
rect 11113 11830 11116 11886
rect 11116 11830 11172 11886
rect 11172 11830 11177 11886
rect 11113 11824 11177 11830
rect 11349 11884 11413 11886
rect 11349 11828 11352 11884
rect 11352 11828 11408 11884
rect 11408 11828 11413 11884
rect 11349 11822 11413 11828
rect 11782 11878 11846 11880
rect 11782 11822 11785 11878
rect 11785 11822 11841 11878
rect 11841 11822 11846 11878
rect 11782 11816 11846 11822
rect 11983 11879 12047 11881
rect 11983 11823 11986 11879
rect 11986 11823 12042 11879
rect 12042 11823 12047 11879
rect 11983 11817 12047 11823
rect 12169 11877 12233 11879
rect 12169 11821 12172 11877
rect 12172 11821 12228 11877
rect 12228 11821 12233 11877
rect 12169 11815 12233 11821
rect 12360 11880 12424 11882
rect 12360 11824 12363 11880
rect 12363 11824 12419 11880
rect 12419 11824 12424 11880
rect 12360 11818 12424 11824
rect 12573 11879 12637 11881
rect 12573 11823 12576 11879
rect 12576 11823 12632 11879
rect 12632 11823 12637 11879
rect 12573 11817 12637 11823
rect 14295 11853 14359 11917
rect 3510 11678 3574 11742
rect 3590 11678 3654 11742
rect 3670 11678 3734 11742
rect 3750 11678 3814 11742
rect 3830 11678 3894 11742
rect 3910 11701 3968 11742
rect 3968 11701 3974 11742
rect 3910 11678 3974 11701
rect 3407 11458 3471 11522
rect 3407 11378 3471 11442
rect 3407 11298 3471 11362
rect 3407 11218 3471 11282
rect 3407 11138 3471 11202
rect 3407 11058 3471 11122
rect 3407 10978 3471 11042
rect 3407 10898 3471 10962
rect 3407 10818 3471 10882
rect 3407 10738 3471 10802
rect 4013 11458 4077 11522
rect 4013 11378 4077 11442
rect 4013 11298 4077 11362
rect 4013 11218 4077 11282
rect 4013 11138 4077 11202
rect 4013 11058 4077 11122
rect 4013 10978 4077 11042
rect 4013 10898 4077 10962
rect 4013 10818 4077 10882
rect 4013 10738 4077 10802
rect 4242 11678 4306 11742
rect 4322 11678 4386 11742
rect 4402 11678 4466 11742
rect 4482 11678 4546 11742
rect 4562 11678 4626 11742
rect 4642 11701 4700 11742
rect 4700 11701 4706 11742
rect 4642 11678 4706 11701
rect 4848 11701 4854 11742
rect 4854 11701 4912 11742
rect 4848 11678 4912 11701
rect 4928 11678 4992 11742
rect 5008 11678 5072 11742
rect 5088 11678 5152 11742
rect 5168 11678 5232 11742
rect 5248 11678 5312 11742
rect 5454 11678 5518 11742
rect 5534 11678 5598 11742
rect 5614 11678 5678 11742
rect 5694 11678 5758 11742
rect 5774 11678 5838 11742
rect 5854 11701 5912 11742
rect 5912 11701 5918 11742
rect 5854 11678 5918 11701
rect 6060 11701 6066 11742
rect 6066 11701 6124 11742
rect 6060 11678 6124 11701
rect 6140 11678 6204 11742
rect 6220 11678 6284 11742
rect 6300 11678 6364 11742
rect 6380 11678 6444 11742
rect 6460 11678 6524 11742
rect 4139 11458 4203 11522
rect 4139 11378 4203 11442
rect 4139 11298 4203 11362
rect 4139 11218 4203 11282
rect 4139 11138 4203 11202
rect 4139 11058 4203 11122
rect 4139 10978 4203 11042
rect 4139 10898 4203 10962
rect 4139 10818 4203 10882
rect 4139 10738 4203 10802
rect 4745 11458 4809 11522
rect 4745 11378 4809 11442
rect 4745 11298 4809 11362
rect 4745 11218 4809 11282
rect 4745 11138 4809 11202
rect 4745 11058 4809 11122
rect 4745 10978 4809 11042
rect 4745 10898 4809 10962
rect 4745 10818 4809 10882
rect 4745 10738 4809 10802
rect 5351 11458 5415 11522
rect 5351 11378 5415 11442
rect 5351 11298 5415 11362
rect 5351 11218 5415 11282
rect 5351 11138 5415 11202
rect 5351 11058 5415 11122
rect 5351 10978 5415 11042
rect 5351 10898 5415 10962
rect 5351 10818 5415 10882
rect 5351 10738 5415 10802
rect 5957 11458 6021 11522
rect 5957 11378 6021 11442
rect 5957 11298 6021 11362
rect 5957 11218 6021 11282
rect 5957 11138 6021 11202
rect 5957 11058 6021 11122
rect 5957 10978 6021 11042
rect 5957 10898 6021 10962
rect 5957 10818 6021 10882
rect 5957 10738 6021 10802
rect 6563 11458 6627 11522
rect 6563 11378 6627 11442
rect 6563 11298 6627 11362
rect 6563 11218 6627 11282
rect 6563 11138 6627 11202
rect 6563 11058 6627 11122
rect 6563 10978 6627 11042
rect 6563 10898 6627 10962
rect 6563 10818 6627 10882
rect 6563 10738 6627 10802
rect 6792 11678 6856 11742
rect 6872 11678 6936 11742
rect 6952 11678 7016 11742
rect 7032 11678 7096 11742
rect 7112 11678 7176 11742
rect 7192 11701 7250 11742
rect 7250 11701 7256 11742
rect 7192 11678 7256 11701
rect 7398 11701 7404 11742
rect 7404 11701 7462 11742
rect 7398 11678 7462 11701
rect 7478 11678 7542 11742
rect 7558 11678 7622 11742
rect 7638 11678 7702 11742
rect 7718 11678 7782 11742
rect 7798 11678 7862 11742
rect 6689 11458 6753 11522
rect 6689 11378 6753 11442
rect 6689 11298 6753 11362
rect 6689 11218 6753 11282
rect 6689 11138 6753 11202
rect 6689 11058 6753 11122
rect 6689 10978 6753 11042
rect 6689 10898 6753 10962
rect 6689 10818 6753 10882
rect 6689 10738 6753 10802
rect 7295 11458 7359 11522
rect 7295 11378 7359 11442
rect 7295 11298 7359 11362
rect 7295 11218 7359 11282
rect 7295 11138 7359 11202
rect 7295 11058 7359 11122
rect 7295 10978 7359 11042
rect 7295 10898 7359 10962
rect 7295 10818 7359 10882
rect 7295 10738 7359 10802
rect 7901 11458 7965 11522
rect 7901 11378 7965 11442
rect 7901 11298 7965 11362
rect 7901 11218 7965 11282
rect 7901 11138 7965 11202
rect 7901 11058 7965 11122
rect 7901 10978 7965 11042
rect 7901 10898 7965 10962
rect 7901 10818 7965 10882
rect 7901 10738 7965 10802
rect 8132 11701 8138 11742
rect 8138 11701 8196 11742
rect 8132 11678 8196 11701
rect 8212 11678 8276 11742
rect 8292 11678 8356 11742
rect 8372 11678 8436 11742
rect 8452 11678 8516 11742
rect 8532 11678 8596 11742
rect 8882 11762 8946 11766
rect 8882 11706 8886 11762
rect 8886 11706 8942 11762
rect 8942 11706 8946 11762
rect 8882 11702 8946 11706
rect 14295 11773 14359 11837
rect 14295 11693 14359 11757
rect 8029 11458 8093 11522
rect 8029 11378 8093 11442
rect 8029 11298 8093 11362
rect 8029 11218 8093 11282
rect 8029 11138 8093 11202
rect 8029 11058 8093 11122
rect 8029 10978 8093 11042
rect 8029 10898 8093 10962
rect 8029 10818 8093 10882
rect 8029 10738 8093 10802
rect 13318 11595 13383 11601
rect 13318 11537 13381 11595
rect 13381 11537 13383 11595
rect 8635 11458 8699 11522
rect 8635 11378 8699 11442
rect 8791 11500 8855 11504
rect 8791 11444 8795 11500
rect 8795 11444 8851 11500
rect 8851 11444 8855 11500
rect 8791 11440 8855 11444
rect 9194 11521 9258 11525
rect 9194 11465 9198 11521
rect 9198 11465 9254 11521
rect 9254 11465 9258 11521
rect 9194 11461 9258 11465
rect 14295 11613 14359 11677
rect 14295 11533 14359 11597
rect 14295 11453 14359 11517
rect 8635 11298 8699 11362
rect 8635 11218 8699 11282
rect 14295 11373 14359 11437
rect 14295 11293 14359 11357
rect 8635 11138 8699 11202
rect 10929 11259 10993 11263
rect 10929 11203 10933 11259
rect 10933 11203 10989 11259
rect 10989 11203 10993 11259
rect 10929 11199 10993 11203
rect 11117 11256 11181 11260
rect 11117 11200 11121 11256
rect 11121 11200 11177 11256
rect 11177 11200 11181 11256
rect 11117 11196 11181 11200
rect 11314 11254 11378 11258
rect 11314 11198 11318 11254
rect 11318 11198 11374 11254
rect 11374 11198 11378 11254
rect 11314 11194 11378 11198
rect 14295 11213 14359 11277
rect 8635 11058 8699 11122
rect 8635 10978 8699 11042
rect 14901 11933 14965 11997
rect 14901 11853 14965 11917
rect 14901 11773 14965 11837
rect 14901 11693 14965 11757
rect 14901 11613 14965 11677
rect 14901 11533 14965 11597
rect 14901 11453 14965 11517
rect 14901 11373 14965 11437
rect 14901 11293 14965 11357
rect 14901 11213 14965 11277
rect 15130 12153 15194 12217
rect 15210 12153 15274 12217
rect 15290 12153 15354 12217
rect 15370 12153 15434 12217
rect 15450 12153 15514 12217
rect 15530 12176 15588 12217
rect 15588 12176 15594 12217
rect 15530 12153 15594 12176
rect 15736 12176 15742 12217
rect 15742 12176 15800 12217
rect 15736 12153 15800 12176
rect 15816 12153 15880 12217
rect 15896 12153 15960 12217
rect 15976 12153 16040 12217
rect 16056 12153 16120 12217
rect 16136 12153 16200 12217
rect 16342 12153 16406 12217
rect 16422 12153 16486 12217
rect 16502 12153 16566 12217
rect 16582 12153 16646 12217
rect 16662 12153 16726 12217
rect 16742 12176 16800 12217
rect 16800 12176 16806 12217
rect 16742 12153 16806 12176
rect 16948 12176 16954 12217
rect 16954 12176 17012 12217
rect 16948 12153 17012 12176
rect 17028 12153 17092 12217
rect 17108 12153 17172 12217
rect 17188 12153 17252 12217
rect 17268 12153 17332 12217
rect 17348 12153 17412 12217
rect 15027 11933 15091 11997
rect 15027 11853 15091 11917
rect 15027 11773 15091 11837
rect 15027 11693 15091 11757
rect 15027 11613 15091 11677
rect 15027 11533 15091 11597
rect 15027 11453 15091 11517
rect 15027 11373 15091 11437
rect 15027 11293 15091 11357
rect 15027 11213 15091 11277
rect 15633 11933 15697 11997
rect 15633 11853 15697 11917
rect 15633 11773 15697 11837
rect 15633 11693 15697 11757
rect 15633 11613 15697 11677
rect 15633 11533 15697 11597
rect 15633 11453 15697 11517
rect 15633 11373 15697 11437
rect 15633 11293 15697 11357
rect 15633 11213 15697 11277
rect 16239 11933 16303 11997
rect 16239 11853 16303 11917
rect 16239 11773 16303 11837
rect 16239 11693 16303 11757
rect 16239 11613 16303 11677
rect 16239 11533 16303 11597
rect 16239 11453 16303 11517
rect 16239 11373 16303 11437
rect 16239 11293 16303 11357
rect 16239 11213 16303 11277
rect 16845 11933 16909 11997
rect 16845 11853 16909 11917
rect 16845 11773 16909 11837
rect 16845 11693 16909 11757
rect 16845 11613 16909 11677
rect 16845 11533 16909 11597
rect 16845 11453 16909 11517
rect 16845 11373 16909 11437
rect 16845 11293 16909 11357
rect 16845 11213 16909 11277
rect 17451 11933 17515 11997
rect 17451 11853 17515 11917
rect 17451 11773 17515 11837
rect 17451 11693 17515 11757
rect 17451 11613 17515 11677
rect 17451 11533 17515 11597
rect 17451 11453 17515 11517
rect 17451 11373 17515 11437
rect 17451 11293 17515 11357
rect 17451 11213 17515 11277
rect 17680 12153 17744 12217
rect 17760 12153 17824 12217
rect 17840 12153 17904 12217
rect 17920 12153 17984 12217
rect 18000 12153 18064 12217
rect 18080 12176 18138 12217
rect 18138 12176 18144 12217
rect 18080 12153 18144 12176
rect 18286 12176 18292 12217
rect 18292 12176 18350 12217
rect 18286 12153 18350 12176
rect 18366 12153 18430 12217
rect 18446 12153 18510 12217
rect 18526 12153 18590 12217
rect 18606 12153 18670 12217
rect 18686 12153 18750 12217
rect 17577 11933 17641 11997
rect 17577 11853 17641 11917
rect 17577 11773 17641 11837
rect 17577 11693 17641 11757
rect 17577 11613 17641 11677
rect 17577 11533 17641 11597
rect 17577 11453 17641 11517
rect 17577 11373 17641 11437
rect 17577 11293 17641 11357
rect 17577 11213 17641 11277
rect 18183 11933 18247 11997
rect 18183 11853 18247 11917
rect 18183 11773 18247 11837
rect 18183 11693 18247 11757
rect 18183 11613 18247 11677
rect 18183 11533 18247 11597
rect 18183 11453 18247 11517
rect 18183 11373 18247 11437
rect 18183 11293 18247 11357
rect 18183 11213 18247 11277
rect 18789 11933 18853 11997
rect 18789 11853 18853 11917
rect 18789 11773 18853 11837
rect 18789 11693 18853 11757
rect 18789 11613 18853 11677
rect 18789 11533 18853 11597
rect 18789 11453 18853 11517
rect 18789 11373 18853 11437
rect 18789 11293 18853 11357
rect 18789 11213 18853 11277
rect 19020 12176 19026 12217
rect 19026 12176 19084 12217
rect 19020 12153 19084 12176
rect 19100 12153 19164 12217
rect 19180 12153 19244 12217
rect 19260 12153 19324 12217
rect 19340 12153 19404 12217
rect 19420 12153 19484 12217
rect 19770 12237 19834 12241
rect 19770 12181 19774 12237
rect 19774 12181 19830 12237
rect 19830 12181 19834 12237
rect 19770 12177 19834 12181
rect 18917 11933 18981 11997
rect 18917 11853 18981 11917
rect 18917 11773 18981 11837
rect 18917 11693 18981 11757
rect 18917 11613 18981 11677
rect 18917 11533 18981 11597
rect 18917 11453 18981 11517
rect 18917 11373 18981 11437
rect 18917 11293 18981 11357
rect 18917 11213 18981 11277
rect 19523 11933 19587 11997
rect 21107 12153 21171 12217
rect 21187 12153 21251 12217
rect 21267 12153 21331 12217
rect 21347 12153 21411 12217
rect 21427 12153 21491 12217
rect 21507 12176 21565 12217
rect 21565 12176 21571 12217
rect 21507 12153 21571 12176
rect 19523 11853 19587 11917
rect 19679 11975 19743 11979
rect 19679 11919 19683 11975
rect 19683 11919 19739 11975
rect 19739 11919 19743 11975
rect 19679 11915 19743 11919
rect 21004 11933 21068 11997
rect 19523 11773 19587 11837
rect 19523 11693 19587 11757
rect 19523 11613 19587 11677
rect 19523 11533 19587 11597
rect 19523 11453 19587 11517
rect 19523 11373 19587 11437
rect 19523 11293 19587 11357
rect 19523 11213 19587 11277
rect 21004 11853 21068 11917
rect 21004 11773 21068 11837
rect 21004 11693 21068 11757
rect 21004 11613 21068 11677
rect 21004 11533 21068 11597
rect 21004 11453 21068 11517
rect 21004 11373 21068 11437
rect 21004 11293 21068 11357
rect 21004 11213 21068 11277
rect 13936 11050 14000 11054
rect 13936 10994 13940 11050
rect 13940 10994 13996 11050
rect 13996 10994 14000 11050
rect 13936 10990 14000 10994
rect 14478 11053 14542 11057
rect 14478 10997 14482 11053
rect 14482 10997 14538 11053
rect 14538 10997 14542 11053
rect 14478 10993 14542 10997
rect 14558 11053 14622 11057
rect 14558 10997 14562 11053
rect 14562 10997 14618 11053
rect 14618 10997 14622 11053
rect 14558 10993 14622 10997
rect 14638 11053 14702 11057
rect 14638 10997 14642 11053
rect 14642 10997 14698 11053
rect 14698 10997 14702 11053
rect 14638 10993 14702 10997
rect 14718 11053 14782 11057
rect 14718 10997 14722 11053
rect 14722 10997 14778 11053
rect 14778 10997 14782 11053
rect 14718 10993 14782 10997
rect 15210 11053 15274 11057
rect 15210 10997 15214 11053
rect 15214 10997 15270 11053
rect 15270 10997 15274 11053
rect 15210 10993 15274 10997
rect 15290 11053 15354 11057
rect 15290 10997 15294 11053
rect 15294 10997 15350 11053
rect 15350 10997 15354 11053
rect 15290 10993 15354 10997
rect 15370 11053 15434 11057
rect 15370 10997 15374 11053
rect 15374 10997 15430 11053
rect 15430 10997 15434 11053
rect 15370 10993 15434 10997
rect 15450 11053 15514 11057
rect 15450 10997 15454 11053
rect 15454 10997 15510 11053
rect 15510 10997 15514 11053
rect 15450 10993 15514 10997
rect 15816 11053 15880 11057
rect 15816 10997 15820 11053
rect 15820 10997 15876 11053
rect 15876 10997 15880 11053
rect 15816 10993 15880 10997
rect 15896 11053 15960 11057
rect 15896 10997 15900 11053
rect 15900 10997 15956 11053
rect 15956 10997 15960 11053
rect 15896 10993 15960 10997
rect 15976 11053 16040 11057
rect 15976 10997 15980 11053
rect 15980 10997 16036 11053
rect 16036 10997 16040 11053
rect 15976 10993 16040 10997
rect 16056 11053 16120 11057
rect 16056 10997 16060 11053
rect 16060 10997 16116 11053
rect 16116 10997 16120 11053
rect 16056 10993 16120 10997
rect 16422 11053 16486 11057
rect 16422 10997 16426 11053
rect 16426 10997 16482 11053
rect 16482 10997 16486 11053
rect 16422 10993 16486 10997
rect 16502 11053 16566 11057
rect 16502 10997 16506 11053
rect 16506 10997 16562 11053
rect 16562 10997 16566 11053
rect 16502 10993 16566 10997
rect 16582 11053 16646 11057
rect 16582 10997 16586 11053
rect 16586 10997 16642 11053
rect 16642 10997 16646 11053
rect 16582 10993 16646 10997
rect 16662 11053 16726 11057
rect 16662 10997 16666 11053
rect 16666 10997 16722 11053
rect 16722 10997 16726 11053
rect 16662 10993 16726 10997
rect 17028 11053 17092 11057
rect 17028 10997 17032 11053
rect 17032 10997 17088 11053
rect 17088 10997 17092 11053
rect 17028 10993 17092 10997
rect 17108 11053 17172 11057
rect 17108 10997 17112 11053
rect 17112 10997 17168 11053
rect 17168 10997 17172 11053
rect 17108 10993 17172 10997
rect 17188 11053 17252 11057
rect 17188 10997 17192 11053
rect 17192 10997 17248 11053
rect 17248 10997 17252 11053
rect 17188 10993 17252 10997
rect 17268 11053 17332 11057
rect 17268 10997 17272 11053
rect 17272 10997 17328 11053
rect 17328 10997 17332 11053
rect 17268 10993 17332 10997
rect 17760 11053 17824 11057
rect 17760 10997 17764 11053
rect 17764 10997 17820 11053
rect 17820 10997 17824 11053
rect 17760 10993 17824 10997
rect 17840 11053 17904 11057
rect 17840 10997 17844 11053
rect 17844 10997 17900 11053
rect 17900 10997 17904 11053
rect 17840 10993 17904 10997
rect 17920 11053 17984 11057
rect 17920 10997 17924 11053
rect 17924 10997 17980 11053
rect 17980 10997 17984 11053
rect 17920 10993 17984 10997
rect 18000 11053 18064 11057
rect 18000 10997 18004 11053
rect 18004 10997 18060 11053
rect 18060 10997 18064 11053
rect 18000 10993 18064 10997
rect 18366 11053 18430 11057
rect 18366 10997 18370 11053
rect 18370 10997 18426 11053
rect 18426 10997 18430 11053
rect 18366 10993 18430 10997
rect 18446 11053 18510 11057
rect 18446 10997 18450 11053
rect 18450 10997 18506 11053
rect 18506 10997 18510 11053
rect 18446 10993 18510 10997
rect 18526 11053 18590 11057
rect 18526 10997 18530 11053
rect 18530 10997 18586 11053
rect 18586 10997 18590 11053
rect 18526 10993 18590 10997
rect 18606 11053 18670 11057
rect 18606 10997 18610 11053
rect 18610 10997 18666 11053
rect 18666 10997 18670 11053
rect 18606 10993 18670 10997
rect 19100 11053 19164 11057
rect 19100 10997 19104 11053
rect 19104 10997 19160 11053
rect 19160 10997 19164 11053
rect 19100 10993 19164 10997
rect 19180 11053 19244 11057
rect 19180 10997 19184 11053
rect 19184 10997 19240 11053
rect 19240 10997 19244 11053
rect 19180 10993 19244 10997
rect 19260 11053 19324 11057
rect 19260 10997 19264 11053
rect 19264 10997 19320 11053
rect 19320 10997 19324 11053
rect 19260 10993 19324 10997
rect 19340 11053 19404 11057
rect 19340 10997 19344 11053
rect 19344 10997 19400 11053
rect 19400 10997 19404 11053
rect 19340 10993 19404 10997
rect 21610 11933 21674 11997
rect 21610 11853 21674 11917
rect 21610 11773 21674 11837
rect 21610 11693 21674 11757
rect 21610 11613 21674 11677
rect 21610 11533 21674 11597
rect 21610 11453 21674 11517
rect 21610 11373 21674 11437
rect 21610 11293 21674 11357
rect 21610 11213 21674 11277
rect 21839 12153 21903 12217
rect 21919 12153 21983 12217
rect 21999 12153 22063 12217
rect 22079 12153 22143 12217
rect 22159 12153 22223 12217
rect 22239 12176 22297 12217
rect 22297 12176 22303 12217
rect 22239 12153 22303 12176
rect 22445 12176 22451 12217
rect 22451 12176 22509 12217
rect 22445 12153 22509 12176
rect 22525 12153 22589 12217
rect 22605 12153 22669 12217
rect 22685 12153 22749 12217
rect 22765 12153 22829 12217
rect 22845 12153 22909 12217
rect 23051 12153 23115 12217
rect 23131 12153 23195 12217
rect 23211 12153 23275 12217
rect 23291 12153 23355 12217
rect 23371 12153 23435 12217
rect 23451 12176 23509 12217
rect 23509 12176 23515 12217
rect 23451 12153 23515 12176
rect 23657 12176 23663 12217
rect 23663 12176 23721 12217
rect 23657 12153 23721 12176
rect 23737 12153 23801 12217
rect 23817 12153 23881 12217
rect 23897 12153 23961 12217
rect 23977 12153 24041 12217
rect 24057 12153 24121 12217
rect 21736 11933 21800 11997
rect 21736 11853 21800 11917
rect 21736 11773 21800 11837
rect 21736 11693 21800 11757
rect 21736 11613 21800 11677
rect 21736 11533 21800 11597
rect 21736 11453 21800 11517
rect 21736 11373 21800 11437
rect 21736 11293 21800 11357
rect 21736 11213 21800 11277
rect 22342 11933 22406 11997
rect 22342 11853 22406 11917
rect 22342 11773 22406 11837
rect 22342 11693 22406 11757
rect 22342 11613 22406 11677
rect 22342 11533 22406 11597
rect 22342 11453 22406 11517
rect 22342 11373 22406 11437
rect 22342 11293 22406 11357
rect 22342 11213 22406 11277
rect 22948 11933 23012 11997
rect 22948 11853 23012 11917
rect 22948 11773 23012 11837
rect 22948 11693 23012 11757
rect 22948 11613 23012 11677
rect 22948 11533 23012 11597
rect 22948 11453 23012 11517
rect 22948 11373 23012 11437
rect 22948 11293 23012 11357
rect 22948 11213 23012 11277
rect 23554 11933 23618 11997
rect 23554 11853 23618 11917
rect 23554 11773 23618 11837
rect 23554 11693 23618 11757
rect 23554 11613 23618 11677
rect 23554 11533 23618 11597
rect 23554 11453 23618 11517
rect 23554 11373 23618 11437
rect 23554 11293 23618 11357
rect 23554 11213 23618 11277
rect 24160 11933 24224 11997
rect 24160 11853 24224 11917
rect 24160 11773 24224 11837
rect 24160 11693 24224 11757
rect 24160 11613 24224 11677
rect 24160 11533 24224 11597
rect 24160 11453 24224 11517
rect 24160 11373 24224 11437
rect 24160 11293 24224 11357
rect 24160 11213 24224 11277
rect 24389 12153 24453 12217
rect 24469 12153 24533 12217
rect 24549 12153 24613 12217
rect 24629 12153 24693 12217
rect 24709 12153 24773 12217
rect 24789 12176 24847 12217
rect 24847 12176 24853 12217
rect 24789 12153 24853 12176
rect 24995 12176 25001 12217
rect 25001 12176 25059 12217
rect 24995 12153 25059 12176
rect 25075 12153 25139 12217
rect 25155 12153 25219 12217
rect 25235 12153 25299 12217
rect 25315 12153 25379 12217
rect 25395 12153 25459 12217
rect 24286 11933 24350 11997
rect 24286 11853 24350 11917
rect 24286 11773 24350 11837
rect 24286 11693 24350 11757
rect 24286 11613 24350 11677
rect 24286 11533 24350 11597
rect 24286 11453 24350 11517
rect 24286 11373 24350 11437
rect 24286 11293 24350 11357
rect 24286 11213 24350 11277
rect 24892 11933 24956 11997
rect 24892 11853 24956 11917
rect 24892 11773 24956 11837
rect 24892 11693 24956 11757
rect 24892 11613 24956 11677
rect 24892 11533 24956 11597
rect 24892 11453 24956 11517
rect 24892 11373 24956 11437
rect 24892 11293 24956 11357
rect 24892 11213 24956 11277
rect 25498 11933 25562 11997
rect 25498 11853 25562 11917
rect 25498 11773 25562 11837
rect 25498 11693 25562 11757
rect 25498 11613 25562 11677
rect 25498 11533 25562 11597
rect 25498 11453 25562 11517
rect 25498 11373 25562 11437
rect 25498 11293 25562 11357
rect 25498 11213 25562 11277
rect 25729 12176 25735 12217
rect 25735 12176 25793 12217
rect 25729 12153 25793 12176
rect 25809 12153 25873 12217
rect 25889 12153 25953 12217
rect 25969 12153 26033 12217
rect 26049 12153 26113 12217
rect 26129 12153 26193 12217
rect 26479 12237 26543 12241
rect 26479 12181 26483 12237
rect 26483 12181 26539 12237
rect 26539 12181 26543 12237
rect 26479 12177 26543 12181
rect 25626 11933 25690 11997
rect 25626 11853 25690 11917
rect 25626 11773 25690 11837
rect 25626 11693 25690 11757
rect 25626 11613 25690 11677
rect 25626 11533 25690 11597
rect 25626 11453 25690 11517
rect 25626 11373 25690 11437
rect 25626 11293 25690 11357
rect 25626 11213 25690 11277
rect 26232 11933 26296 11997
rect 26232 11853 26296 11917
rect 26388 11975 26452 11979
rect 26388 11919 26392 11975
rect 26392 11919 26448 11975
rect 26448 11919 26452 11975
rect 26388 11915 26452 11919
rect 26232 11773 26296 11837
rect 26232 11693 26296 11757
rect 26232 11613 26296 11677
rect 26232 11533 26296 11597
rect 26232 11453 26296 11517
rect 26232 11373 26296 11437
rect 26232 11293 26296 11357
rect 26232 11213 26296 11277
rect 20645 11050 20709 11054
rect 20645 10994 20649 11050
rect 20649 10994 20705 11050
rect 20705 10994 20709 11050
rect 20645 10990 20709 10994
rect 21187 11053 21251 11057
rect 21187 10997 21191 11053
rect 21191 10997 21247 11053
rect 21247 10997 21251 11053
rect 21187 10993 21251 10997
rect 21267 11053 21331 11057
rect 21267 10997 21271 11053
rect 21271 10997 21327 11053
rect 21327 10997 21331 11053
rect 21267 10993 21331 10997
rect 21347 11053 21411 11057
rect 21347 10997 21351 11053
rect 21351 10997 21407 11053
rect 21407 10997 21411 11053
rect 21347 10993 21411 10997
rect 21427 11053 21491 11057
rect 21427 10997 21431 11053
rect 21431 10997 21487 11053
rect 21487 10997 21491 11053
rect 21427 10993 21491 10997
rect 21919 11053 21983 11057
rect 21919 10997 21923 11053
rect 21923 10997 21979 11053
rect 21979 10997 21983 11053
rect 21919 10993 21983 10997
rect 21999 11053 22063 11057
rect 21999 10997 22003 11053
rect 22003 10997 22059 11053
rect 22059 10997 22063 11053
rect 21999 10993 22063 10997
rect 22079 11053 22143 11057
rect 22079 10997 22083 11053
rect 22083 10997 22139 11053
rect 22139 10997 22143 11053
rect 22079 10993 22143 10997
rect 22159 11053 22223 11057
rect 22159 10997 22163 11053
rect 22163 10997 22219 11053
rect 22219 10997 22223 11053
rect 22159 10993 22223 10997
rect 22525 11053 22589 11057
rect 22525 10997 22529 11053
rect 22529 10997 22585 11053
rect 22585 10997 22589 11053
rect 22525 10993 22589 10997
rect 22605 11053 22669 11057
rect 22605 10997 22609 11053
rect 22609 10997 22665 11053
rect 22665 10997 22669 11053
rect 22605 10993 22669 10997
rect 22685 11053 22749 11057
rect 22685 10997 22689 11053
rect 22689 10997 22745 11053
rect 22745 10997 22749 11053
rect 22685 10993 22749 10997
rect 22765 11053 22829 11057
rect 22765 10997 22769 11053
rect 22769 10997 22825 11053
rect 22825 10997 22829 11053
rect 22765 10993 22829 10997
rect 23131 11053 23195 11057
rect 23131 10997 23135 11053
rect 23135 10997 23191 11053
rect 23191 10997 23195 11053
rect 23131 10993 23195 10997
rect 23211 11053 23275 11057
rect 23211 10997 23215 11053
rect 23215 10997 23271 11053
rect 23271 10997 23275 11053
rect 23211 10993 23275 10997
rect 23291 11053 23355 11057
rect 23291 10997 23295 11053
rect 23295 10997 23351 11053
rect 23351 10997 23355 11053
rect 23291 10993 23355 10997
rect 23371 11053 23435 11057
rect 23371 10997 23375 11053
rect 23375 10997 23431 11053
rect 23431 10997 23435 11053
rect 23371 10993 23435 10997
rect 23737 11053 23801 11057
rect 23737 10997 23741 11053
rect 23741 10997 23797 11053
rect 23797 10997 23801 11053
rect 23737 10993 23801 10997
rect 23817 11053 23881 11057
rect 23817 10997 23821 11053
rect 23821 10997 23877 11053
rect 23877 10997 23881 11053
rect 23817 10993 23881 10997
rect 23897 11053 23961 11057
rect 23897 10997 23901 11053
rect 23901 10997 23957 11053
rect 23957 10997 23961 11053
rect 23897 10993 23961 10997
rect 23977 11053 24041 11057
rect 23977 10997 23981 11053
rect 23981 10997 24037 11053
rect 24037 10997 24041 11053
rect 23977 10993 24041 10997
rect 24469 11053 24533 11057
rect 24469 10997 24473 11053
rect 24473 10997 24529 11053
rect 24529 10997 24533 11053
rect 24469 10993 24533 10997
rect 24549 11053 24613 11057
rect 24549 10997 24553 11053
rect 24553 10997 24609 11053
rect 24609 10997 24613 11053
rect 24549 10993 24613 10997
rect 24629 11053 24693 11057
rect 24629 10997 24633 11053
rect 24633 10997 24689 11053
rect 24689 10997 24693 11053
rect 24629 10993 24693 10997
rect 24709 11053 24773 11057
rect 24709 10997 24713 11053
rect 24713 10997 24769 11053
rect 24769 10997 24773 11053
rect 24709 10993 24773 10997
rect 25075 11053 25139 11057
rect 25075 10997 25079 11053
rect 25079 10997 25135 11053
rect 25135 10997 25139 11053
rect 25075 10993 25139 10997
rect 25155 11053 25219 11057
rect 25155 10997 25159 11053
rect 25159 10997 25215 11053
rect 25215 10997 25219 11053
rect 25155 10993 25219 10997
rect 25235 11053 25299 11057
rect 25235 10997 25239 11053
rect 25239 10997 25295 11053
rect 25295 10997 25299 11053
rect 25235 10993 25299 10997
rect 25315 11053 25379 11057
rect 25315 10997 25319 11053
rect 25319 10997 25375 11053
rect 25375 10997 25379 11053
rect 25315 10993 25379 10997
rect 25809 11053 25873 11057
rect 25809 10997 25813 11053
rect 25813 10997 25869 11053
rect 25869 10997 25873 11053
rect 25809 10993 25873 10997
rect 25889 11053 25953 11057
rect 25889 10997 25893 11053
rect 25893 10997 25949 11053
rect 25949 10997 25953 11053
rect 25889 10993 25953 10997
rect 25969 11053 26033 11057
rect 25969 10997 25973 11053
rect 25973 10997 26029 11053
rect 26029 10997 26033 11053
rect 25969 10993 26033 10997
rect 26049 11053 26113 11057
rect 26049 10997 26053 11053
rect 26053 10997 26109 11053
rect 26109 10997 26113 11053
rect 26049 10993 26113 10997
rect 8635 10898 8699 10962
rect 8635 10818 8699 10882
rect 8635 10738 8699 10802
rect 3048 10575 3112 10579
rect 3048 10519 3052 10575
rect 3052 10519 3108 10575
rect 3108 10519 3112 10575
rect 3048 10515 3112 10519
rect 3590 10578 3654 10582
rect 3590 10522 3594 10578
rect 3594 10522 3650 10578
rect 3650 10522 3654 10578
rect 3590 10518 3654 10522
rect 3670 10578 3734 10582
rect 3670 10522 3674 10578
rect 3674 10522 3730 10578
rect 3730 10522 3734 10578
rect 3670 10518 3734 10522
rect 3750 10578 3814 10582
rect 3750 10522 3754 10578
rect 3754 10522 3810 10578
rect 3810 10522 3814 10578
rect 3750 10518 3814 10522
rect 3830 10578 3894 10582
rect 3830 10522 3834 10578
rect 3834 10522 3890 10578
rect 3890 10522 3894 10578
rect 3830 10518 3894 10522
rect 4322 10578 4386 10582
rect 4322 10522 4326 10578
rect 4326 10522 4382 10578
rect 4382 10522 4386 10578
rect 4322 10518 4386 10522
rect 4402 10578 4466 10582
rect 4402 10522 4406 10578
rect 4406 10522 4462 10578
rect 4462 10522 4466 10578
rect 4402 10518 4466 10522
rect 4482 10578 4546 10582
rect 4482 10522 4486 10578
rect 4486 10522 4542 10578
rect 4542 10522 4546 10578
rect 4482 10518 4546 10522
rect 4562 10578 4626 10582
rect 4562 10522 4566 10578
rect 4566 10522 4622 10578
rect 4622 10522 4626 10578
rect 4562 10518 4626 10522
rect 4928 10578 4992 10582
rect 4928 10522 4932 10578
rect 4932 10522 4988 10578
rect 4988 10522 4992 10578
rect 4928 10518 4992 10522
rect 5008 10578 5072 10582
rect 5008 10522 5012 10578
rect 5012 10522 5068 10578
rect 5068 10522 5072 10578
rect 5008 10518 5072 10522
rect 5088 10578 5152 10582
rect 5088 10522 5092 10578
rect 5092 10522 5148 10578
rect 5148 10522 5152 10578
rect 5088 10518 5152 10522
rect 5168 10578 5232 10582
rect 5168 10522 5172 10578
rect 5172 10522 5228 10578
rect 5228 10522 5232 10578
rect 5168 10518 5232 10522
rect 5534 10578 5598 10582
rect 5534 10522 5538 10578
rect 5538 10522 5594 10578
rect 5594 10522 5598 10578
rect 5534 10518 5598 10522
rect 5614 10578 5678 10582
rect 5614 10522 5618 10578
rect 5618 10522 5674 10578
rect 5674 10522 5678 10578
rect 5614 10518 5678 10522
rect 5694 10578 5758 10582
rect 5694 10522 5698 10578
rect 5698 10522 5754 10578
rect 5754 10522 5758 10578
rect 5694 10518 5758 10522
rect 5774 10578 5838 10582
rect 5774 10522 5778 10578
rect 5778 10522 5834 10578
rect 5834 10522 5838 10578
rect 5774 10518 5838 10522
rect 6140 10578 6204 10582
rect 6140 10522 6144 10578
rect 6144 10522 6200 10578
rect 6200 10522 6204 10578
rect 6140 10518 6204 10522
rect 6220 10578 6284 10582
rect 6220 10522 6224 10578
rect 6224 10522 6280 10578
rect 6280 10522 6284 10578
rect 6220 10518 6284 10522
rect 6300 10578 6364 10582
rect 6300 10522 6304 10578
rect 6304 10522 6360 10578
rect 6360 10522 6364 10578
rect 6300 10518 6364 10522
rect 6380 10578 6444 10582
rect 6380 10522 6384 10578
rect 6384 10522 6440 10578
rect 6440 10522 6444 10578
rect 6380 10518 6444 10522
rect 6872 10578 6936 10582
rect 6872 10522 6876 10578
rect 6876 10522 6932 10578
rect 6932 10522 6936 10578
rect 6872 10518 6936 10522
rect 6952 10578 7016 10582
rect 6952 10522 6956 10578
rect 6956 10522 7012 10578
rect 7012 10522 7016 10578
rect 6952 10518 7016 10522
rect 7032 10578 7096 10582
rect 7032 10522 7036 10578
rect 7036 10522 7092 10578
rect 7092 10522 7096 10578
rect 7032 10518 7096 10522
rect 7112 10578 7176 10582
rect 7112 10522 7116 10578
rect 7116 10522 7172 10578
rect 7172 10522 7176 10578
rect 7112 10518 7176 10522
rect 7478 10578 7542 10582
rect 7478 10522 7482 10578
rect 7482 10522 7538 10578
rect 7538 10522 7542 10578
rect 7478 10518 7542 10522
rect 7558 10578 7622 10582
rect 7558 10522 7562 10578
rect 7562 10522 7618 10578
rect 7618 10522 7622 10578
rect 7558 10518 7622 10522
rect 7638 10578 7702 10582
rect 7638 10522 7642 10578
rect 7642 10522 7698 10578
rect 7698 10522 7702 10578
rect 7638 10518 7702 10522
rect 7718 10578 7782 10582
rect 7718 10522 7722 10578
rect 7722 10522 7778 10578
rect 7778 10522 7782 10578
rect 7718 10518 7782 10522
rect 8212 10578 8276 10582
rect 8212 10522 8216 10578
rect 8216 10522 8272 10578
rect 8272 10522 8276 10578
rect 8212 10518 8276 10522
rect 8292 10578 8356 10582
rect 8292 10522 8296 10578
rect 8296 10522 8352 10578
rect 8352 10522 8356 10578
rect 8292 10518 8356 10522
rect 8372 10578 8436 10582
rect 8372 10522 8376 10578
rect 8376 10522 8432 10578
rect 8432 10522 8436 10578
rect 8372 10518 8436 10522
rect 8452 10578 8516 10582
rect 8452 10522 8456 10578
rect 8456 10522 8512 10578
rect 8512 10522 8516 10578
rect 8452 10518 8516 10522
rect 3048 10127 3112 10131
rect 3048 10071 3052 10127
rect 3052 10071 3108 10127
rect 3108 10071 3112 10127
rect 3048 10067 3112 10071
rect 3590 10124 3654 10128
rect 3590 10068 3594 10124
rect 3594 10068 3650 10124
rect 3650 10068 3654 10124
rect 3590 10064 3654 10068
rect 3670 10124 3734 10128
rect 3670 10068 3674 10124
rect 3674 10068 3730 10124
rect 3730 10068 3734 10124
rect 3670 10064 3734 10068
rect 3750 10124 3814 10128
rect 3750 10068 3754 10124
rect 3754 10068 3810 10124
rect 3810 10068 3814 10124
rect 3750 10064 3814 10068
rect 3830 10124 3894 10128
rect 3830 10068 3834 10124
rect 3834 10068 3890 10124
rect 3890 10068 3894 10124
rect 3830 10064 3894 10068
rect 4322 10124 4386 10128
rect 4322 10068 4326 10124
rect 4326 10068 4382 10124
rect 4382 10068 4386 10124
rect 4322 10064 4386 10068
rect 4402 10124 4466 10128
rect 4402 10068 4406 10124
rect 4406 10068 4462 10124
rect 4462 10068 4466 10124
rect 4402 10064 4466 10068
rect 4482 10124 4546 10128
rect 4482 10068 4486 10124
rect 4486 10068 4542 10124
rect 4542 10068 4546 10124
rect 4482 10064 4546 10068
rect 4562 10124 4626 10128
rect 4562 10068 4566 10124
rect 4566 10068 4622 10124
rect 4622 10068 4626 10124
rect 4562 10064 4626 10068
rect 4928 10124 4992 10128
rect 4928 10068 4932 10124
rect 4932 10068 4988 10124
rect 4988 10068 4992 10124
rect 4928 10064 4992 10068
rect 5008 10124 5072 10128
rect 5008 10068 5012 10124
rect 5012 10068 5068 10124
rect 5068 10068 5072 10124
rect 5008 10064 5072 10068
rect 5088 10124 5152 10128
rect 5088 10068 5092 10124
rect 5092 10068 5148 10124
rect 5148 10068 5152 10124
rect 5088 10064 5152 10068
rect 5168 10124 5232 10128
rect 5168 10068 5172 10124
rect 5172 10068 5228 10124
rect 5228 10068 5232 10124
rect 5168 10064 5232 10068
rect 5534 10124 5598 10128
rect 5534 10068 5538 10124
rect 5538 10068 5594 10124
rect 5594 10068 5598 10124
rect 5534 10064 5598 10068
rect 5614 10124 5678 10128
rect 5614 10068 5618 10124
rect 5618 10068 5674 10124
rect 5674 10068 5678 10124
rect 5614 10064 5678 10068
rect 5694 10124 5758 10128
rect 5694 10068 5698 10124
rect 5698 10068 5754 10124
rect 5754 10068 5758 10124
rect 5694 10064 5758 10068
rect 5774 10124 5838 10128
rect 5774 10068 5778 10124
rect 5778 10068 5834 10124
rect 5834 10068 5838 10124
rect 5774 10064 5838 10068
rect 6140 10124 6204 10128
rect 6140 10068 6144 10124
rect 6144 10068 6200 10124
rect 6200 10068 6204 10124
rect 6140 10064 6204 10068
rect 6220 10124 6284 10128
rect 6220 10068 6224 10124
rect 6224 10068 6280 10124
rect 6280 10068 6284 10124
rect 6220 10064 6284 10068
rect 6300 10124 6364 10128
rect 6300 10068 6304 10124
rect 6304 10068 6360 10124
rect 6360 10068 6364 10124
rect 6300 10064 6364 10068
rect 6380 10124 6444 10128
rect 6380 10068 6384 10124
rect 6384 10068 6440 10124
rect 6440 10068 6444 10124
rect 6380 10064 6444 10068
rect 6872 10124 6936 10128
rect 6872 10068 6876 10124
rect 6876 10068 6932 10124
rect 6932 10068 6936 10124
rect 6872 10064 6936 10068
rect 6952 10124 7016 10128
rect 6952 10068 6956 10124
rect 6956 10068 7012 10124
rect 7012 10068 7016 10124
rect 6952 10064 7016 10068
rect 7032 10124 7096 10128
rect 7032 10068 7036 10124
rect 7036 10068 7092 10124
rect 7092 10068 7096 10124
rect 7032 10064 7096 10068
rect 7112 10124 7176 10128
rect 7112 10068 7116 10124
rect 7116 10068 7172 10124
rect 7172 10068 7176 10124
rect 7112 10064 7176 10068
rect 7478 10124 7542 10128
rect 7478 10068 7482 10124
rect 7482 10068 7538 10124
rect 7538 10068 7542 10124
rect 7478 10064 7542 10068
rect 7558 10124 7622 10128
rect 7558 10068 7562 10124
rect 7562 10068 7618 10124
rect 7618 10068 7622 10124
rect 7558 10064 7622 10068
rect 7638 10124 7702 10128
rect 7638 10068 7642 10124
rect 7642 10068 7698 10124
rect 7698 10068 7702 10124
rect 7638 10064 7702 10068
rect 7718 10124 7782 10128
rect 7718 10068 7722 10124
rect 7722 10068 7778 10124
rect 7778 10068 7782 10124
rect 7718 10064 7782 10068
rect 8212 10124 8276 10128
rect 8212 10068 8216 10124
rect 8216 10068 8272 10124
rect 8272 10068 8276 10124
rect 8212 10064 8276 10068
rect 8292 10124 8356 10128
rect 8292 10068 8296 10124
rect 8296 10068 8352 10124
rect 8352 10068 8356 10124
rect 8292 10064 8356 10068
rect 8372 10124 8436 10128
rect 8372 10068 8376 10124
rect 8376 10068 8432 10124
rect 8432 10068 8436 10124
rect 8372 10064 8436 10068
rect 8452 10124 8516 10128
rect 8452 10068 8456 10124
rect 8456 10068 8512 10124
rect 8512 10068 8516 10124
rect 8452 10064 8516 10068
rect 3407 9844 3471 9908
rect 3407 9764 3471 9828
rect 3407 9684 3471 9748
rect 3407 9604 3471 9668
rect 3407 9524 3471 9588
rect 3407 9444 3471 9508
rect 3407 9364 3471 9428
rect 3407 9284 3471 9348
rect 3407 9204 3471 9268
rect 3407 9124 3471 9188
rect 4013 9844 4077 9908
rect 4013 9764 4077 9828
rect 4013 9684 4077 9748
rect 4013 9604 4077 9668
rect 4013 9524 4077 9588
rect 4013 9444 4077 9508
rect 4013 9364 4077 9428
rect 4013 9284 4077 9348
rect 4013 9204 4077 9268
rect 4013 9124 4077 9188
rect 3510 8904 3574 8968
rect 3590 8904 3654 8968
rect 3670 8904 3734 8968
rect 3750 8904 3814 8968
rect 3830 8904 3894 8968
rect 3910 8945 3974 8968
rect 3910 8904 3968 8945
rect 3968 8904 3974 8945
rect 4139 9844 4203 9908
rect 4139 9764 4203 9828
rect 4139 9684 4203 9748
rect 4139 9604 4203 9668
rect 4139 9524 4203 9588
rect 4139 9444 4203 9508
rect 4139 9364 4203 9428
rect 4139 9284 4203 9348
rect 4139 9204 4203 9268
rect 4139 9124 4203 9188
rect 4745 9844 4809 9908
rect 4745 9764 4809 9828
rect 4745 9684 4809 9748
rect 4745 9604 4809 9668
rect 4745 9524 4809 9588
rect 4745 9444 4809 9508
rect 4745 9364 4809 9428
rect 4745 9284 4809 9348
rect 4745 9204 4809 9268
rect 4745 9124 4809 9188
rect 5351 9844 5415 9908
rect 5351 9764 5415 9828
rect 5351 9684 5415 9748
rect 5351 9604 5415 9668
rect 5351 9524 5415 9588
rect 5351 9444 5415 9508
rect 5351 9364 5415 9428
rect 5351 9284 5415 9348
rect 5351 9204 5415 9268
rect 5351 9124 5415 9188
rect 5957 9844 6021 9908
rect 5957 9764 6021 9828
rect 5957 9684 6021 9748
rect 5957 9604 6021 9668
rect 5957 9524 6021 9588
rect 5957 9444 6021 9508
rect 5957 9364 6021 9428
rect 5957 9284 6021 9348
rect 5957 9204 6021 9268
rect 5957 9124 6021 9188
rect 6563 9844 6627 9908
rect 6563 9764 6627 9828
rect 6563 9684 6627 9748
rect 6563 9604 6627 9668
rect 6563 9524 6627 9588
rect 6563 9444 6627 9508
rect 6563 9364 6627 9428
rect 6563 9284 6627 9348
rect 6563 9204 6627 9268
rect 6563 9124 6627 9188
rect 4242 8904 4306 8968
rect 4322 8904 4386 8968
rect 4402 8904 4466 8968
rect 4482 8904 4546 8968
rect 4562 8904 4626 8968
rect 4642 8945 4706 8968
rect 4642 8904 4700 8945
rect 4700 8904 4706 8945
rect 4848 8945 4912 8968
rect 4848 8904 4854 8945
rect 4854 8904 4912 8945
rect 4928 8904 4992 8968
rect 5008 8904 5072 8968
rect 5088 8904 5152 8968
rect 5168 8904 5232 8968
rect 5248 8904 5312 8968
rect 5454 8904 5518 8968
rect 5534 8904 5598 8968
rect 5614 8904 5678 8968
rect 5694 8904 5758 8968
rect 5774 8904 5838 8968
rect 5854 8945 5918 8968
rect 5854 8904 5912 8945
rect 5912 8904 5918 8945
rect 6060 8945 6124 8968
rect 6060 8904 6066 8945
rect 6066 8904 6124 8945
rect 6140 8904 6204 8968
rect 6220 8904 6284 8968
rect 6300 8904 6364 8968
rect 6380 8904 6444 8968
rect 6460 8904 6524 8968
rect 6689 9844 6753 9908
rect 6689 9764 6753 9828
rect 6689 9684 6753 9748
rect 6689 9604 6753 9668
rect 6689 9524 6753 9588
rect 6689 9444 6753 9508
rect 6689 9364 6753 9428
rect 6689 9284 6753 9348
rect 6689 9204 6753 9268
rect 6689 9124 6753 9188
rect 7295 9844 7359 9908
rect 7295 9764 7359 9828
rect 7295 9684 7359 9748
rect 7295 9604 7359 9668
rect 7295 9524 7359 9588
rect 7295 9444 7359 9508
rect 7295 9364 7359 9428
rect 7295 9284 7359 9348
rect 7295 9204 7359 9268
rect 7295 9124 7359 9188
rect 7901 9844 7965 9908
rect 7901 9764 7965 9828
rect 7901 9684 7965 9748
rect 7901 9604 7965 9668
rect 7901 9524 7965 9588
rect 7901 9444 7965 9508
rect 7901 9364 7965 9428
rect 7901 9284 7965 9348
rect 7901 9204 7965 9268
rect 7901 9124 7965 9188
rect 6792 8904 6856 8968
rect 6872 8904 6936 8968
rect 6952 8904 7016 8968
rect 7032 8904 7096 8968
rect 7112 8904 7176 8968
rect 7192 8945 7256 8968
rect 7192 8904 7250 8945
rect 7250 8904 7256 8945
rect 7398 8945 7462 8968
rect 7398 8904 7404 8945
rect 7404 8904 7462 8945
rect 7478 8904 7542 8968
rect 7558 8904 7622 8968
rect 7638 8904 7702 8968
rect 7718 8904 7782 8968
rect 7798 8904 7862 8968
rect 8029 9844 8093 9908
rect 8029 9764 8093 9828
rect 8029 9684 8093 9748
rect 8029 9604 8093 9668
rect 8029 9524 8093 9588
rect 8029 9444 8093 9508
rect 8029 9364 8093 9428
rect 8029 9284 8093 9348
rect 8029 9204 8093 9268
rect 8029 9124 8093 9188
rect 13775 10112 13839 10116
rect 13775 10056 13779 10112
rect 13779 10056 13835 10112
rect 13835 10056 13839 10112
rect 13775 10052 13839 10056
rect 13855 10112 13919 10116
rect 13855 10056 13859 10112
rect 13859 10056 13915 10112
rect 13915 10056 13919 10112
rect 13855 10052 13919 10056
rect 13935 10112 13999 10116
rect 13935 10056 13939 10112
rect 13939 10056 13995 10112
rect 13995 10056 13999 10112
rect 13935 10052 13999 10056
rect 14015 10112 14079 10116
rect 14015 10056 14019 10112
rect 14019 10056 14075 10112
rect 14075 10056 14079 10112
rect 14015 10052 14079 10056
rect 14509 10112 14573 10116
rect 14509 10056 14513 10112
rect 14513 10056 14569 10112
rect 14569 10056 14573 10112
rect 14509 10052 14573 10056
rect 14589 10112 14653 10116
rect 14589 10056 14593 10112
rect 14593 10056 14649 10112
rect 14649 10056 14653 10112
rect 14589 10052 14653 10056
rect 14669 10112 14733 10116
rect 14669 10056 14673 10112
rect 14673 10056 14729 10112
rect 14729 10056 14733 10112
rect 14669 10052 14733 10056
rect 14749 10112 14813 10116
rect 14749 10056 14753 10112
rect 14753 10056 14809 10112
rect 14809 10056 14813 10112
rect 14749 10052 14813 10056
rect 15115 10112 15179 10116
rect 15115 10056 15119 10112
rect 15119 10056 15175 10112
rect 15175 10056 15179 10112
rect 15115 10052 15179 10056
rect 15195 10112 15259 10116
rect 15195 10056 15199 10112
rect 15199 10056 15255 10112
rect 15255 10056 15259 10112
rect 15195 10052 15259 10056
rect 15275 10112 15339 10116
rect 15275 10056 15279 10112
rect 15279 10056 15335 10112
rect 15335 10056 15339 10112
rect 15275 10052 15339 10056
rect 15355 10112 15419 10116
rect 15355 10056 15359 10112
rect 15359 10056 15415 10112
rect 15415 10056 15419 10112
rect 15355 10052 15419 10056
rect 15847 10112 15911 10116
rect 15847 10056 15851 10112
rect 15851 10056 15907 10112
rect 15907 10056 15911 10112
rect 15847 10052 15911 10056
rect 15927 10112 15991 10116
rect 15927 10056 15931 10112
rect 15931 10056 15987 10112
rect 15987 10056 15991 10112
rect 15927 10052 15991 10056
rect 16007 10112 16071 10116
rect 16007 10056 16011 10112
rect 16011 10056 16067 10112
rect 16067 10056 16071 10112
rect 16007 10052 16071 10056
rect 16087 10112 16151 10116
rect 16087 10056 16091 10112
rect 16091 10056 16147 10112
rect 16147 10056 16151 10112
rect 16087 10052 16151 10056
rect 16453 10112 16517 10116
rect 16453 10056 16457 10112
rect 16457 10056 16513 10112
rect 16513 10056 16517 10112
rect 16453 10052 16517 10056
rect 16533 10112 16597 10116
rect 16533 10056 16537 10112
rect 16537 10056 16593 10112
rect 16593 10056 16597 10112
rect 16533 10052 16597 10056
rect 16613 10112 16677 10116
rect 16613 10056 16617 10112
rect 16617 10056 16673 10112
rect 16673 10056 16677 10112
rect 16613 10052 16677 10056
rect 16693 10112 16757 10116
rect 16693 10056 16697 10112
rect 16697 10056 16753 10112
rect 16753 10056 16757 10112
rect 16693 10052 16757 10056
rect 17059 10112 17123 10116
rect 17059 10056 17063 10112
rect 17063 10056 17119 10112
rect 17119 10056 17123 10112
rect 17059 10052 17123 10056
rect 17139 10112 17203 10116
rect 17139 10056 17143 10112
rect 17143 10056 17199 10112
rect 17199 10056 17203 10112
rect 17139 10052 17203 10056
rect 17219 10112 17283 10116
rect 17219 10056 17223 10112
rect 17223 10056 17279 10112
rect 17279 10056 17283 10112
rect 17219 10052 17283 10056
rect 17299 10112 17363 10116
rect 17299 10056 17303 10112
rect 17303 10056 17359 10112
rect 17359 10056 17363 10112
rect 17299 10052 17363 10056
rect 17665 10112 17729 10116
rect 17665 10056 17669 10112
rect 17669 10056 17725 10112
rect 17725 10056 17729 10112
rect 17665 10052 17729 10056
rect 17745 10112 17809 10116
rect 17745 10056 17749 10112
rect 17749 10056 17805 10112
rect 17805 10056 17809 10112
rect 17745 10052 17809 10056
rect 17825 10112 17889 10116
rect 17825 10056 17829 10112
rect 17829 10056 17885 10112
rect 17885 10056 17889 10112
rect 17825 10052 17889 10056
rect 17905 10112 17969 10116
rect 17905 10056 17909 10112
rect 17909 10056 17965 10112
rect 17965 10056 17969 10112
rect 17905 10052 17969 10056
rect 18397 10112 18461 10116
rect 18397 10056 18401 10112
rect 18401 10056 18457 10112
rect 18457 10056 18461 10112
rect 18397 10052 18461 10056
rect 18477 10112 18541 10116
rect 18477 10056 18481 10112
rect 18481 10056 18537 10112
rect 18537 10056 18541 10112
rect 18477 10052 18541 10056
rect 18557 10112 18621 10116
rect 18557 10056 18561 10112
rect 18561 10056 18617 10112
rect 18617 10056 18621 10112
rect 18557 10052 18621 10056
rect 18637 10112 18701 10116
rect 18637 10056 18641 10112
rect 18641 10056 18697 10112
rect 18697 10056 18701 10112
rect 18637 10052 18701 10056
rect 19179 10115 19243 10119
rect 19179 10059 19183 10115
rect 19183 10059 19239 10115
rect 19239 10059 19243 10115
rect 19179 10055 19243 10059
rect 8635 9844 8699 9908
rect 8635 9764 8699 9828
rect 8635 9684 8699 9748
rect 8635 9604 8699 9668
rect 8635 9524 8699 9588
rect 8635 9444 8699 9508
rect 8635 9364 8699 9428
rect 8635 9284 8699 9348
rect 8635 9204 8699 9268
rect 13592 9832 13656 9896
rect 13592 9752 13656 9816
rect 13592 9672 13656 9736
rect 13592 9592 13656 9656
rect 13592 9512 13656 9576
rect 13592 9432 13656 9496
rect 13592 9352 13656 9416
rect 13592 9272 13656 9336
rect 8635 9124 8699 9188
rect 8791 9202 8855 9206
rect 8791 9146 8795 9202
rect 8795 9146 8851 9202
rect 8851 9146 8855 9202
rect 8791 9142 8855 9146
rect 9219 9161 9283 9165
rect 9219 9105 9223 9161
rect 9223 9105 9279 9161
rect 9279 9105 9283 9161
rect 9219 9101 9283 9105
rect 9696 9161 9760 9165
rect 9696 9105 9700 9161
rect 9700 9105 9756 9161
rect 9756 9105 9760 9161
rect 9696 9101 9760 9105
rect 10116 9150 10180 9154
rect 10116 9094 10120 9150
rect 10120 9094 10176 9150
rect 10176 9094 10180 9150
rect 10116 9090 10180 9094
rect 10492 9158 10556 9162
rect 10492 9102 10496 9158
rect 10496 9102 10552 9158
rect 10552 9102 10556 9158
rect 10492 9098 10556 9102
rect 10840 9158 10904 9162
rect 10840 9102 10844 9158
rect 10844 9102 10900 9158
rect 10900 9102 10904 9158
rect 10840 9098 10904 9102
rect 11098 9164 11162 9168
rect 11098 9108 11102 9164
rect 11102 9108 11158 9164
rect 11158 9108 11162 9164
rect 11098 9104 11162 9108
rect 11324 9164 11388 9168
rect 11324 9108 11328 9164
rect 11328 9108 11384 9164
rect 11384 9108 11388 9164
rect 11324 9104 11388 9108
rect 11583 9167 11647 9171
rect 11583 9111 11587 9167
rect 11587 9111 11643 9167
rect 11643 9111 11647 9167
rect 11583 9107 11647 9111
rect 12190 9129 12254 9133
rect 12190 9073 12194 9129
rect 12194 9073 12250 9129
rect 12250 9073 12254 9129
rect 12190 9069 12254 9073
rect 12422 9130 12486 9134
rect 12422 9074 12426 9130
rect 12426 9074 12482 9130
rect 12482 9074 12486 9130
rect 12422 9070 12486 9074
rect 12858 9136 12922 9140
rect 12858 9080 12862 9136
rect 12862 9080 12918 9136
rect 12918 9080 12922 9136
rect 12858 9076 12922 9080
rect 13093 9138 13157 9142
rect 13093 9082 13097 9138
rect 13097 9082 13153 9138
rect 13153 9082 13157 9138
rect 13093 9078 13157 9082
rect 13436 9190 13500 9194
rect 13436 9134 13440 9190
rect 13440 9134 13496 9190
rect 13496 9134 13500 9190
rect 13436 9130 13500 9134
rect 13592 9192 13656 9256
rect 13592 9112 13656 9176
rect 8132 8945 8196 8968
rect 8132 8904 8138 8945
rect 8138 8904 8196 8945
rect 8212 8904 8276 8968
rect 8292 8904 8356 8968
rect 8372 8904 8436 8968
rect 8452 8904 8516 8968
rect 8532 8904 8596 8968
rect 14198 9832 14262 9896
rect 14198 9752 14262 9816
rect 14198 9672 14262 9736
rect 14198 9592 14262 9656
rect 14198 9512 14262 9576
rect 14198 9432 14262 9496
rect 14198 9352 14262 9416
rect 14198 9272 14262 9336
rect 14198 9192 14262 9256
rect 14198 9112 14262 9176
rect 8882 8940 8946 8944
rect 8882 8884 8886 8940
rect 8886 8884 8942 8940
rect 8942 8884 8946 8940
rect 8882 8880 8946 8884
rect 13345 8928 13409 8932
rect 13345 8872 13349 8928
rect 13349 8872 13405 8928
rect 13405 8872 13409 8928
rect 13345 8868 13409 8872
rect 13695 8892 13759 8956
rect 13775 8892 13839 8956
rect 13855 8892 13919 8956
rect 13935 8892 13999 8956
rect 14015 8892 14079 8956
rect 14095 8933 14159 8956
rect 14095 8892 14153 8933
rect 14153 8892 14159 8933
rect 14326 9832 14390 9896
rect 14326 9752 14390 9816
rect 14326 9672 14390 9736
rect 14326 9592 14390 9656
rect 14326 9512 14390 9576
rect 14326 9432 14390 9496
rect 14326 9352 14390 9416
rect 14326 9272 14390 9336
rect 14326 9192 14390 9256
rect 14326 9112 14390 9176
rect 14932 9832 14996 9896
rect 14932 9752 14996 9816
rect 14932 9672 14996 9736
rect 14932 9592 14996 9656
rect 14932 9512 14996 9576
rect 14932 9432 14996 9496
rect 14932 9352 14996 9416
rect 14932 9272 14996 9336
rect 14932 9192 14996 9256
rect 14932 9112 14996 9176
rect 15538 9832 15602 9896
rect 15538 9752 15602 9816
rect 15538 9672 15602 9736
rect 15538 9592 15602 9656
rect 15538 9512 15602 9576
rect 15538 9432 15602 9496
rect 15538 9352 15602 9416
rect 15538 9272 15602 9336
rect 15538 9192 15602 9256
rect 15538 9112 15602 9176
rect 14429 8892 14493 8956
rect 14509 8892 14573 8956
rect 14589 8892 14653 8956
rect 14669 8892 14733 8956
rect 14749 8892 14813 8956
rect 14829 8933 14893 8956
rect 14829 8892 14887 8933
rect 14887 8892 14893 8933
rect 15035 8933 15099 8956
rect 15035 8892 15041 8933
rect 15041 8892 15099 8933
rect 15115 8892 15179 8956
rect 15195 8892 15259 8956
rect 15275 8892 15339 8956
rect 15355 8892 15419 8956
rect 15435 8892 15499 8956
rect 15664 9832 15728 9896
rect 15664 9752 15728 9816
rect 15664 9672 15728 9736
rect 15664 9592 15728 9656
rect 15664 9512 15728 9576
rect 15664 9432 15728 9496
rect 15664 9352 15728 9416
rect 15664 9272 15728 9336
rect 15664 9192 15728 9256
rect 15664 9112 15728 9176
rect 16270 9832 16334 9896
rect 16270 9752 16334 9816
rect 16270 9672 16334 9736
rect 16270 9592 16334 9656
rect 16270 9512 16334 9576
rect 16270 9432 16334 9496
rect 16270 9352 16334 9416
rect 16270 9272 16334 9336
rect 16270 9192 16334 9256
rect 16270 9112 16334 9176
rect 16876 9832 16940 9896
rect 16876 9752 16940 9816
rect 16876 9672 16940 9736
rect 16876 9592 16940 9656
rect 16876 9512 16940 9576
rect 16876 9432 16940 9496
rect 16876 9352 16940 9416
rect 16876 9272 16940 9336
rect 16876 9192 16940 9256
rect 16876 9112 16940 9176
rect 17482 9832 17546 9896
rect 17482 9752 17546 9816
rect 17482 9672 17546 9736
rect 17482 9592 17546 9656
rect 17482 9512 17546 9576
rect 17482 9432 17546 9496
rect 17482 9352 17546 9416
rect 17482 9272 17546 9336
rect 17482 9192 17546 9256
rect 17482 9112 17546 9176
rect 18088 9832 18152 9896
rect 18088 9752 18152 9816
rect 18088 9672 18152 9736
rect 18088 9592 18152 9656
rect 18088 9512 18152 9576
rect 18088 9432 18152 9496
rect 18088 9352 18152 9416
rect 18088 9272 18152 9336
rect 18088 9192 18152 9256
rect 18088 9112 18152 9176
rect 15767 8892 15831 8956
rect 15847 8892 15911 8956
rect 15927 8892 15991 8956
rect 16007 8892 16071 8956
rect 16087 8892 16151 8956
rect 16167 8933 16231 8956
rect 16167 8892 16225 8933
rect 16225 8892 16231 8933
rect 16373 8933 16437 8956
rect 16373 8892 16379 8933
rect 16379 8892 16437 8933
rect 16453 8892 16517 8956
rect 16533 8892 16597 8956
rect 16613 8892 16677 8956
rect 16693 8892 16757 8956
rect 16773 8892 16837 8956
rect 16979 8892 17043 8956
rect 17059 8892 17123 8956
rect 17139 8892 17203 8956
rect 17219 8892 17283 8956
rect 17299 8892 17363 8956
rect 17379 8933 17443 8956
rect 17379 8892 17437 8933
rect 17437 8892 17443 8933
rect 17585 8933 17649 8956
rect 17585 8892 17591 8933
rect 17591 8892 17649 8933
rect 17665 8892 17729 8956
rect 17745 8892 17809 8956
rect 17825 8892 17889 8956
rect 17905 8892 17969 8956
rect 17985 8892 18049 8956
rect 18214 9832 18278 9896
rect 18214 9752 18278 9816
rect 18214 9672 18278 9736
rect 18214 9592 18278 9656
rect 18214 9512 18278 9576
rect 18214 9432 18278 9496
rect 18214 9352 18278 9416
rect 18214 9272 18278 9336
rect 18214 9192 18278 9256
rect 18214 9112 18278 9176
rect 20484 10112 20548 10116
rect 20484 10056 20488 10112
rect 20488 10056 20544 10112
rect 20544 10056 20548 10112
rect 20484 10052 20548 10056
rect 20564 10112 20628 10116
rect 20564 10056 20568 10112
rect 20568 10056 20624 10112
rect 20624 10056 20628 10112
rect 20564 10052 20628 10056
rect 20644 10112 20708 10116
rect 20644 10056 20648 10112
rect 20648 10056 20704 10112
rect 20704 10056 20708 10112
rect 20644 10052 20708 10056
rect 20724 10112 20788 10116
rect 20724 10056 20728 10112
rect 20728 10056 20784 10112
rect 20784 10056 20788 10112
rect 20724 10052 20788 10056
rect 21218 10112 21282 10116
rect 21218 10056 21222 10112
rect 21222 10056 21278 10112
rect 21278 10056 21282 10112
rect 21218 10052 21282 10056
rect 21298 10112 21362 10116
rect 21298 10056 21302 10112
rect 21302 10056 21358 10112
rect 21358 10056 21362 10112
rect 21298 10052 21362 10056
rect 21378 10112 21442 10116
rect 21378 10056 21382 10112
rect 21382 10056 21438 10112
rect 21438 10056 21442 10112
rect 21378 10052 21442 10056
rect 21458 10112 21522 10116
rect 21458 10056 21462 10112
rect 21462 10056 21518 10112
rect 21518 10056 21522 10112
rect 21458 10052 21522 10056
rect 21824 10112 21888 10116
rect 21824 10056 21828 10112
rect 21828 10056 21884 10112
rect 21884 10056 21888 10112
rect 21824 10052 21888 10056
rect 21904 10112 21968 10116
rect 21904 10056 21908 10112
rect 21908 10056 21964 10112
rect 21964 10056 21968 10112
rect 21904 10052 21968 10056
rect 21984 10112 22048 10116
rect 21984 10056 21988 10112
rect 21988 10056 22044 10112
rect 22044 10056 22048 10112
rect 21984 10052 22048 10056
rect 22064 10112 22128 10116
rect 22064 10056 22068 10112
rect 22068 10056 22124 10112
rect 22124 10056 22128 10112
rect 22064 10052 22128 10056
rect 22556 10112 22620 10116
rect 22556 10056 22560 10112
rect 22560 10056 22616 10112
rect 22616 10056 22620 10112
rect 22556 10052 22620 10056
rect 22636 10112 22700 10116
rect 22636 10056 22640 10112
rect 22640 10056 22696 10112
rect 22696 10056 22700 10112
rect 22636 10052 22700 10056
rect 22716 10112 22780 10116
rect 22716 10056 22720 10112
rect 22720 10056 22776 10112
rect 22776 10056 22780 10112
rect 22716 10052 22780 10056
rect 22796 10112 22860 10116
rect 22796 10056 22800 10112
rect 22800 10056 22856 10112
rect 22856 10056 22860 10112
rect 22796 10052 22860 10056
rect 23162 10112 23226 10116
rect 23162 10056 23166 10112
rect 23166 10056 23222 10112
rect 23222 10056 23226 10112
rect 23162 10052 23226 10056
rect 23242 10112 23306 10116
rect 23242 10056 23246 10112
rect 23246 10056 23302 10112
rect 23302 10056 23306 10112
rect 23242 10052 23306 10056
rect 23322 10112 23386 10116
rect 23322 10056 23326 10112
rect 23326 10056 23382 10112
rect 23382 10056 23386 10112
rect 23322 10052 23386 10056
rect 23402 10112 23466 10116
rect 23402 10056 23406 10112
rect 23406 10056 23462 10112
rect 23462 10056 23466 10112
rect 23402 10052 23466 10056
rect 23768 10112 23832 10116
rect 23768 10056 23772 10112
rect 23772 10056 23828 10112
rect 23828 10056 23832 10112
rect 23768 10052 23832 10056
rect 23848 10112 23912 10116
rect 23848 10056 23852 10112
rect 23852 10056 23908 10112
rect 23908 10056 23912 10112
rect 23848 10052 23912 10056
rect 23928 10112 23992 10116
rect 23928 10056 23932 10112
rect 23932 10056 23988 10112
rect 23988 10056 23992 10112
rect 23928 10052 23992 10056
rect 24008 10112 24072 10116
rect 24008 10056 24012 10112
rect 24012 10056 24068 10112
rect 24068 10056 24072 10112
rect 24008 10052 24072 10056
rect 24374 10112 24438 10116
rect 24374 10056 24378 10112
rect 24378 10056 24434 10112
rect 24434 10056 24438 10112
rect 24374 10052 24438 10056
rect 24454 10112 24518 10116
rect 24454 10056 24458 10112
rect 24458 10056 24514 10112
rect 24514 10056 24518 10112
rect 24454 10052 24518 10056
rect 24534 10112 24598 10116
rect 24534 10056 24538 10112
rect 24538 10056 24594 10112
rect 24594 10056 24598 10112
rect 24534 10052 24598 10056
rect 24614 10112 24678 10116
rect 24614 10056 24618 10112
rect 24618 10056 24674 10112
rect 24674 10056 24678 10112
rect 24614 10052 24678 10056
rect 25106 10112 25170 10116
rect 25106 10056 25110 10112
rect 25110 10056 25166 10112
rect 25166 10056 25170 10112
rect 25106 10052 25170 10056
rect 25186 10112 25250 10116
rect 25186 10056 25190 10112
rect 25190 10056 25246 10112
rect 25246 10056 25250 10112
rect 25186 10052 25250 10056
rect 25266 10112 25330 10116
rect 25266 10056 25270 10112
rect 25270 10056 25326 10112
rect 25326 10056 25330 10112
rect 25266 10052 25330 10056
rect 25346 10112 25410 10116
rect 25346 10056 25350 10112
rect 25350 10056 25406 10112
rect 25406 10056 25410 10112
rect 25346 10052 25410 10056
rect 25888 10115 25952 10119
rect 25888 10059 25892 10115
rect 25892 10059 25948 10115
rect 25948 10059 25952 10115
rect 25888 10055 25952 10059
rect 18820 9832 18884 9896
rect 18820 9752 18884 9816
rect 18820 9672 18884 9736
rect 18820 9592 18884 9656
rect 18820 9512 18884 9576
rect 18820 9432 18884 9496
rect 18820 9352 18884 9416
rect 18820 9272 18884 9336
rect 18820 9192 18884 9256
rect 20301 9832 20365 9896
rect 20301 9752 20365 9816
rect 20301 9672 20365 9736
rect 20301 9592 20365 9656
rect 20301 9512 20365 9576
rect 20301 9432 20365 9496
rect 20301 9352 20365 9416
rect 20301 9272 20365 9336
rect 18820 9112 18884 9176
rect 20145 9190 20209 9194
rect 20145 9134 20149 9190
rect 20149 9134 20205 9190
rect 20205 9134 20209 9190
rect 20145 9130 20209 9134
rect 20301 9192 20365 9256
rect 18317 8933 18381 8956
rect 18317 8892 18323 8933
rect 18323 8892 18381 8933
rect 18397 8892 18461 8956
rect 18477 8892 18541 8956
rect 18557 8892 18621 8956
rect 18637 8892 18701 8956
rect 18717 8892 18781 8956
rect 20301 9112 20365 9176
rect 20907 9832 20971 9896
rect 20907 9752 20971 9816
rect 20907 9672 20971 9736
rect 20907 9592 20971 9656
rect 20907 9512 20971 9576
rect 20907 9432 20971 9496
rect 20907 9352 20971 9416
rect 20907 9272 20971 9336
rect 20907 9192 20971 9256
rect 20907 9112 20971 9176
rect 20054 8928 20118 8932
rect 20054 8872 20058 8928
rect 20058 8872 20114 8928
rect 20114 8872 20118 8928
rect 20054 8868 20118 8872
rect 20404 8892 20468 8956
rect 20484 8892 20548 8956
rect 20564 8892 20628 8956
rect 20644 8892 20708 8956
rect 20724 8892 20788 8956
rect 20804 8933 20868 8956
rect 20804 8892 20862 8933
rect 20862 8892 20868 8933
rect 21035 9832 21099 9896
rect 21035 9752 21099 9816
rect 21035 9672 21099 9736
rect 21035 9592 21099 9656
rect 21035 9512 21099 9576
rect 21035 9432 21099 9496
rect 21035 9352 21099 9416
rect 21035 9272 21099 9336
rect 21035 9192 21099 9256
rect 21035 9112 21099 9176
rect 21641 9832 21705 9896
rect 21641 9752 21705 9816
rect 21641 9672 21705 9736
rect 21641 9592 21705 9656
rect 21641 9512 21705 9576
rect 21641 9432 21705 9496
rect 21641 9352 21705 9416
rect 21641 9272 21705 9336
rect 21641 9192 21705 9256
rect 21641 9112 21705 9176
rect 22247 9832 22311 9896
rect 22247 9752 22311 9816
rect 22247 9672 22311 9736
rect 22247 9592 22311 9656
rect 22247 9512 22311 9576
rect 22247 9432 22311 9496
rect 22247 9352 22311 9416
rect 22247 9272 22311 9336
rect 22247 9192 22311 9256
rect 22247 9112 22311 9176
rect 21138 8892 21202 8956
rect 21218 8892 21282 8956
rect 21298 8892 21362 8956
rect 21378 8892 21442 8956
rect 21458 8892 21522 8956
rect 21538 8933 21602 8956
rect 21538 8892 21596 8933
rect 21596 8892 21602 8933
rect 21744 8933 21808 8956
rect 21744 8892 21750 8933
rect 21750 8892 21808 8933
rect 21824 8892 21888 8956
rect 21904 8892 21968 8956
rect 21984 8892 22048 8956
rect 22064 8892 22128 8956
rect 22144 8892 22208 8956
rect 22373 9832 22437 9896
rect 22373 9752 22437 9816
rect 22373 9672 22437 9736
rect 22373 9592 22437 9656
rect 22373 9512 22437 9576
rect 22373 9432 22437 9496
rect 22373 9352 22437 9416
rect 22373 9272 22437 9336
rect 22373 9192 22437 9256
rect 22373 9112 22437 9176
rect 22979 9832 23043 9896
rect 22979 9752 23043 9816
rect 22979 9672 23043 9736
rect 22979 9592 23043 9656
rect 22979 9512 23043 9576
rect 22979 9432 23043 9496
rect 22979 9352 23043 9416
rect 22979 9272 23043 9336
rect 22979 9192 23043 9256
rect 22979 9112 23043 9176
rect 23585 9832 23649 9896
rect 23585 9752 23649 9816
rect 23585 9672 23649 9736
rect 23585 9592 23649 9656
rect 23585 9512 23649 9576
rect 23585 9432 23649 9496
rect 23585 9352 23649 9416
rect 23585 9272 23649 9336
rect 23585 9192 23649 9256
rect 23585 9112 23649 9176
rect 24191 9832 24255 9896
rect 24191 9752 24255 9816
rect 24191 9672 24255 9736
rect 24191 9592 24255 9656
rect 24191 9512 24255 9576
rect 24191 9432 24255 9496
rect 24191 9352 24255 9416
rect 24191 9272 24255 9336
rect 24191 9192 24255 9256
rect 24191 9112 24255 9176
rect 24797 9832 24861 9896
rect 24797 9752 24861 9816
rect 24797 9672 24861 9736
rect 24797 9592 24861 9656
rect 24797 9512 24861 9576
rect 24797 9432 24861 9496
rect 24797 9352 24861 9416
rect 24797 9272 24861 9336
rect 24797 9192 24861 9256
rect 24797 9112 24861 9176
rect 22476 8892 22540 8956
rect 22556 8892 22620 8956
rect 22636 8892 22700 8956
rect 22716 8892 22780 8956
rect 22796 8892 22860 8956
rect 22876 8933 22940 8956
rect 22876 8892 22934 8933
rect 22934 8892 22940 8933
rect 23082 8933 23146 8956
rect 23082 8892 23088 8933
rect 23088 8892 23146 8933
rect 23162 8892 23226 8956
rect 23242 8892 23306 8956
rect 23322 8892 23386 8956
rect 23402 8892 23466 8956
rect 23482 8892 23546 8956
rect 23688 8892 23752 8956
rect 23768 8892 23832 8956
rect 23848 8892 23912 8956
rect 23928 8892 23992 8956
rect 24008 8892 24072 8956
rect 24088 8933 24152 8956
rect 24088 8892 24146 8933
rect 24146 8892 24152 8933
rect 24294 8933 24358 8956
rect 24294 8892 24300 8933
rect 24300 8892 24358 8933
rect 24374 8892 24438 8956
rect 24454 8892 24518 8956
rect 24534 8892 24598 8956
rect 24614 8892 24678 8956
rect 24694 8892 24758 8956
rect 24923 9832 24987 9896
rect 24923 9752 24987 9816
rect 24923 9672 24987 9736
rect 24923 9592 24987 9656
rect 24923 9512 24987 9576
rect 24923 9432 24987 9496
rect 24923 9352 24987 9416
rect 24923 9272 24987 9336
rect 24923 9192 24987 9256
rect 24923 9112 24987 9176
rect 25529 9832 25593 9896
rect 25529 9752 25593 9816
rect 25529 9672 25593 9736
rect 25529 9592 25593 9656
rect 25529 9512 25593 9576
rect 25529 9432 25593 9496
rect 25529 9352 25593 9416
rect 25529 9272 25593 9336
rect 25529 9192 25593 9256
rect 25529 9112 25593 9176
rect 25026 8933 25090 8956
rect 25026 8892 25032 8933
rect 25032 8892 25090 8933
rect 25106 8892 25170 8956
rect 25186 8892 25250 8956
rect 25266 8892 25330 8956
rect 25346 8892 25410 8956
rect 25426 8892 25490 8956
rect 2463 8700 2527 8704
rect 2463 8644 2467 8700
rect 2467 8644 2523 8700
rect 2523 8644 2527 8700
rect 2463 8640 2527 8644
rect 2583 8700 2647 8704
rect 2583 8644 2587 8700
rect 2587 8644 2643 8700
rect 2643 8644 2647 8700
rect 2583 8640 2647 8644
rect 2726 8700 2790 8704
rect 2726 8644 2730 8700
rect 2730 8644 2786 8700
rect 2786 8644 2790 8700
rect 2726 8640 2790 8644
rect 3159 8659 3223 8723
rect 3239 8659 3303 8723
rect 3319 8659 3383 8723
rect 3399 8659 3463 8723
rect 3479 8659 3543 8723
rect 3559 8682 3612 8723
rect 3612 8682 3623 8723
rect 3559 8659 3623 8682
rect 3056 8439 3120 8503
rect 3056 8359 3120 8423
rect 3056 8279 3120 8343
rect 3056 8199 3120 8263
rect 2445 8154 2509 8158
rect 2445 8098 2449 8154
rect 2449 8098 2505 8154
rect 2505 8098 2509 8154
rect 2445 8094 2509 8098
rect 2576 8155 2640 8159
rect 2576 8099 2580 8155
rect 2580 8099 2636 8155
rect 2636 8099 2640 8155
rect 2576 8095 2640 8099
rect 2720 8154 2784 8158
rect 2720 8098 2724 8154
rect 2724 8098 2780 8154
rect 2780 8098 2784 8154
rect 2720 8094 2784 8098
rect 3056 8119 3120 8183
rect 3056 8039 3120 8103
rect 3056 7959 3120 8023
rect 3056 7879 3120 7943
rect 3056 7799 3120 7863
rect 3056 7719 3120 7783
rect 3662 8439 3726 8503
rect 3662 8359 3726 8423
rect 3662 8279 3726 8343
rect 3662 8199 3726 8263
rect 3662 8119 3726 8183
rect 3662 8039 3726 8103
rect 3662 7959 3726 8023
rect 3662 7879 3726 7943
rect 3662 7799 3726 7863
rect 3662 7719 3726 7783
rect 3891 8656 3955 8720
rect 3971 8656 4035 8720
rect 4051 8656 4115 8720
rect 4131 8656 4195 8720
rect 4211 8656 4275 8720
rect 4291 8679 4344 8720
rect 4344 8679 4355 8720
rect 4291 8656 4355 8679
rect 4497 8679 4508 8720
rect 4508 8679 4561 8720
rect 4497 8656 4561 8679
rect 4577 8656 4641 8720
rect 4657 8656 4721 8720
rect 4737 8656 4801 8720
rect 4817 8656 4881 8720
rect 4897 8656 4961 8720
rect 5103 8656 5167 8720
rect 5183 8656 5247 8720
rect 5263 8656 5327 8720
rect 5343 8656 5407 8720
rect 5423 8656 5487 8720
rect 5503 8679 5556 8720
rect 5556 8679 5567 8720
rect 5503 8656 5567 8679
rect 5709 8679 5720 8720
rect 5720 8679 5773 8720
rect 5709 8656 5773 8679
rect 5789 8656 5853 8720
rect 5869 8656 5933 8720
rect 5949 8656 6013 8720
rect 6029 8656 6093 8720
rect 6109 8656 6173 8720
rect 6315 8656 6379 8720
rect 6395 8656 6459 8720
rect 6475 8656 6539 8720
rect 6555 8656 6619 8720
rect 6635 8656 6699 8720
rect 6715 8679 6768 8720
rect 6768 8679 6779 8720
rect 6715 8656 6779 8679
rect 6921 8679 6932 8720
rect 6932 8679 6985 8720
rect 6921 8656 6985 8679
rect 7001 8656 7065 8720
rect 7081 8656 7145 8720
rect 7161 8656 7225 8720
rect 7241 8656 7305 8720
rect 7321 8656 7385 8720
rect 7527 8656 7591 8720
rect 7607 8656 7671 8720
rect 7687 8656 7751 8720
rect 7767 8656 7831 8720
rect 7847 8656 7911 8720
rect 7927 8679 7980 8720
rect 7980 8679 7991 8720
rect 7927 8656 7991 8679
rect 8133 8679 8144 8720
rect 8144 8679 8197 8720
rect 8133 8656 8197 8679
rect 8213 8656 8277 8720
rect 8293 8656 8357 8720
rect 8373 8656 8437 8720
rect 8453 8656 8517 8720
rect 8533 8656 8597 8720
rect 8882 8737 8946 8741
rect 8882 8681 8886 8737
rect 8886 8681 8942 8737
rect 8942 8681 8946 8737
rect 8882 8677 8946 8681
rect 13345 8725 13409 8729
rect 13345 8669 13349 8725
rect 13349 8669 13405 8725
rect 13405 8669 13409 8725
rect 13345 8665 13409 8669
rect 3788 8436 3852 8500
rect 3788 8356 3852 8420
rect 3788 8276 3852 8340
rect 3788 8196 3852 8260
rect 3788 8116 3852 8180
rect 3788 8036 3852 8100
rect 3788 7956 3852 8020
rect 3788 7876 3852 7940
rect 3788 7796 3852 7860
rect 3788 7716 3852 7780
rect 3159 7558 3223 7563
rect 3062 7549 3126 7553
rect 3062 7493 3066 7549
rect 3066 7493 3122 7549
rect 3122 7493 3126 7549
rect 3159 7502 3162 7558
rect 3162 7502 3218 7558
rect 3218 7502 3223 7558
rect 3159 7499 3223 7502
rect 3239 7558 3303 7563
rect 3239 7502 3242 7558
rect 3242 7502 3298 7558
rect 3298 7502 3303 7558
rect 3239 7499 3303 7502
rect 3319 7558 3383 7563
rect 3319 7502 3322 7558
rect 3322 7502 3378 7558
rect 3378 7502 3383 7558
rect 3319 7499 3383 7502
rect 3399 7558 3463 7563
rect 3399 7502 3402 7558
rect 3402 7502 3458 7558
rect 3458 7502 3463 7558
rect 3399 7499 3463 7502
rect 3479 7558 3543 7563
rect 3479 7502 3482 7558
rect 3482 7502 3538 7558
rect 3538 7502 3543 7558
rect 3479 7499 3543 7502
rect 3559 7558 3623 7563
rect 3559 7502 3562 7558
rect 3562 7502 3618 7558
rect 3618 7502 3623 7558
rect 3559 7499 3623 7502
rect 4394 8436 4458 8500
rect 4394 8356 4458 8420
rect 4394 8276 4458 8340
rect 4394 8196 4458 8260
rect 4394 8116 4458 8180
rect 4394 8036 4458 8100
rect 4394 7956 4458 8020
rect 4394 7876 4458 7940
rect 4394 7796 4458 7860
rect 4394 7716 4458 7780
rect 5000 8436 5064 8500
rect 5000 8356 5064 8420
rect 5000 8276 5064 8340
rect 5000 8196 5064 8260
rect 5000 8116 5064 8180
rect 5000 8036 5064 8100
rect 5000 7956 5064 8020
rect 5000 7876 5064 7940
rect 5000 7796 5064 7860
rect 5000 7716 5064 7780
rect 5606 8436 5670 8500
rect 5606 8356 5670 8420
rect 5606 8276 5670 8340
rect 5606 8196 5670 8260
rect 5606 8116 5670 8180
rect 5606 8036 5670 8100
rect 5606 7956 5670 8020
rect 5606 7876 5670 7940
rect 5606 7796 5670 7860
rect 5606 7716 5670 7780
rect 6212 8436 6276 8500
rect 6212 8356 6276 8420
rect 6212 8276 6276 8340
rect 6212 8196 6276 8260
rect 6212 8116 6276 8180
rect 6212 8036 6276 8100
rect 6212 7956 6276 8020
rect 6212 7876 6276 7940
rect 6212 7796 6276 7860
rect 6212 7716 6276 7780
rect 6818 8436 6882 8500
rect 6818 8356 6882 8420
rect 6818 8276 6882 8340
rect 6818 8196 6882 8260
rect 6818 8116 6882 8180
rect 6818 8036 6882 8100
rect 6818 7956 6882 8020
rect 6818 7876 6882 7940
rect 6818 7796 6882 7860
rect 6818 7716 6882 7780
rect 7424 8436 7488 8500
rect 7424 8356 7488 8420
rect 7424 8276 7488 8340
rect 7424 8196 7488 8260
rect 7424 8116 7488 8180
rect 7424 8036 7488 8100
rect 7424 7956 7488 8020
rect 7424 7876 7488 7940
rect 7424 7796 7488 7860
rect 7424 7716 7488 7780
rect 8030 8436 8094 8500
rect 8030 8356 8094 8420
rect 8030 8276 8094 8340
rect 8030 8196 8094 8260
rect 8030 8116 8094 8180
rect 8030 8036 8094 8100
rect 8030 7956 8094 8020
rect 8030 7876 8094 7940
rect 8030 7796 8094 7860
rect 8030 7716 8094 7780
rect 13694 8644 13758 8708
rect 13774 8644 13838 8708
rect 13854 8644 13918 8708
rect 13934 8644 13998 8708
rect 14014 8644 14078 8708
rect 14094 8667 14147 8708
rect 14147 8667 14158 8708
rect 14094 8644 14158 8667
rect 14300 8667 14311 8708
rect 14311 8667 14364 8708
rect 14300 8644 14364 8667
rect 14380 8644 14444 8708
rect 14460 8644 14524 8708
rect 14540 8644 14604 8708
rect 14620 8644 14684 8708
rect 14700 8644 14764 8708
rect 14906 8644 14970 8708
rect 14986 8644 15050 8708
rect 15066 8644 15130 8708
rect 15146 8644 15210 8708
rect 15226 8644 15290 8708
rect 15306 8667 15359 8708
rect 15359 8667 15370 8708
rect 15306 8644 15370 8667
rect 15512 8667 15523 8708
rect 15523 8667 15576 8708
rect 15512 8644 15576 8667
rect 15592 8644 15656 8708
rect 15672 8644 15736 8708
rect 15752 8644 15816 8708
rect 15832 8644 15896 8708
rect 15912 8644 15976 8708
rect 16118 8644 16182 8708
rect 16198 8644 16262 8708
rect 16278 8644 16342 8708
rect 16358 8644 16422 8708
rect 16438 8644 16502 8708
rect 16518 8667 16571 8708
rect 16571 8667 16582 8708
rect 16518 8644 16582 8667
rect 16724 8667 16735 8708
rect 16735 8667 16788 8708
rect 16724 8644 16788 8667
rect 16804 8644 16868 8708
rect 16884 8644 16948 8708
rect 16964 8644 17028 8708
rect 17044 8644 17108 8708
rect 17124 8644 17188 8708
rect 17330 8644 17394 8708
rect 17410 8644 17474 8708
rect 17490 8644 17554 8708
rect 17570 8644 17634 8708
rect 17650 8644 17714 8708
rect 17730 8667 17783 8708
rect 17783 8667 17794 8708
rect 17730 8644 17794 8667
rect 17936 8667 17947 8708
rect 17947 8667 18000 8708
rect 17936 8644 18000 8667
rect 18016 8644 18080 8708
rect 18096 8644 18160 8708
rect 18176 8644 18240 8708
rect 18256 8644 18320 8708
rect 18336 8644 18400 8708
rect 8636 8436 8700 8500
rect 8636 8356 8700 8420
rect 8794 8476 8858 8480
rect 8794 8420 8798 8476
rect 8798 8420 8854 8476
rect 8854 8420 8858 8476
rect 8794 8416 8858 8420
rect 9204 8450 9268 8454
rect 9204 8394 9208 8450
rect 9208 8394 9264 8450
rect 9264 8394 9268 8450
rect 9204 8390 9268 8394
rect 9466 8451 9530 8455
rect 9466 8395 9470 8451
rect 9470 8395 9526 8451
rect 9526 8395 9530 8451
rect 9466 8391 9530 8395
rect 9738 8451 9802 8455
rect 9738 8395 9742 8451
rect 9742 8395 9798 8451
rect 9798 8395 9802 8451
rect 9738 8391 9802 8395
rect 10065 8451 10129 8455
rect 10065 8395 10069 8451
rect 10069 8395 10125 8451
rect 10125 8395 10129 8451
rect 10065 8391 10129 8395
rect 10446 8451 10510 8455
rect 10446 8395 10450 8451
rect 10450 8395 10506 8451
rect 10506 8395 10510 8451
rect 10446 8391 10510 8395
rect 10823 8451 10887 8455
rect 10823 8395 10827 8451
rect 10827 8395 10883 8451
rect 10883 8395 10887 8451
rect 10823 8391 10887 8395
rect 12224 8440 12288 8442
rect 12224 8384 12227 8440
rect 12227 8384 12283 8440
rect 12283 8384 12288 8440
rect 12224 8378 12288 8384
rect 12719 8510 12783 8512
rect 12719 8454 12722 8510
rect 12722 8454 12778 8510
rect 12778 8454 12783 8510
rect 12719 8448 12783 8454
rect 13093 8510 13157 8512
rect 13093 8454 13096 8510
rect 13096 8454 13152 8510
rect 13152 8454 13157 8510
rect 13093 8448 13157 8454
rect 13433 8464 13497 8468
rect 13433 8408 13437 8464
rect 13437 8408 13493 8464
rect 13493 8408 13497 8464
rect 13433 8404 13497 8408
rect 13591 8424 13655 8488
rect 8636 8276 8700 8340
rect 12581 8367 12645 8369
rect 12581 8311 12584 8367
rect 12584 8311 12640 8367
rect 12640 8311 12645 8367
rect 12581 8305 12645 8311
rect 12765 8364 12829 8366
rect 12765 8308 12768 8364
rect 12768 8308 12824 8364
rect 12824 8308 12829 8364
rect 12765 8302 12829 8308
rect 13067 8358 13131 8360
rect 13067 8302 13070 8358
rect 13070 8302 13126 8358
rect 13126 8302 13131 8358
rect 13067 8296 13131 8302
rect 13591 8344 13655 8408
rect 8636 8196 8700 8260
rect 13591 8264 13655 8328
rect 8636 8116 8700 8180
rect 8876 8234 8940 8238
rect 8876 8178 8880 8234
rect 8880 8178 8936 8234
rect 8936 8178 8940 8234
rect 8876 8174 8940 8178
rect 13351 8222 13415 8226
rect 13351 8166 13355 8222
rect 13355 8166 13411 8222
rect 13411 8166 13415 8222
rect 13351 8162 13415 8166
rect 13591 8184 13655 8248
rect 8636 8036 8700 8100
rect 13591 8104 13655 8168
rect 8636 7956 8700 8020
rect 8877 8077 8941 8081
rect 8877 8021 8881 8077
rect 8881 8021 8937 8077
rect 8937 8021 8941 8077
rect 8877 8017 8941 8021
rect 13350 8065 13414 8069
rect 13350 8009 13354 8065
rect 13354 8009 13410 8065
rect 13410 8009 13414 8065
rect 13350 8005 13414 8009
rect 13591 8024 13655 8088
rect 8636 7876 8700 7940
rect 8636 7796 8700 7860
rect 8877 7907 8941 7911
rect 8877 7851 8881 7907
rect 8881 7851 8937 7907
rect 8937 7851 8941 7907
rect 8877 7847 8941 7851
rect 12934 7931 12998 7935
rect 12934 7875 12938 7931
rect 12938 7875 12994 7931
rect 12994 7875 12998 7931
rect 12934 7871 12998 7875
rect 13591 7944 13655 8008
rect 13350 7895 13414 7899
rect 13350 7839 13354 7895
rect 13354 7839 13410 7895
rect 13410 7839 13414 7895
rect 13350 7835 13414 7839
rect 13591 7864 13655 7928
rect 8636 7716 8700 7780
rect 13591 7784 13655 7848
rect 8876 7755 8940 7759
rect 8876 7699 8880 7755
rect 8880 7699 8936 7755
rect 8936 7699 8940 7755
rect 8876 7695 8940 7699
rect 10140 7725 10204 7729
rect 10140 7669 10144 7725
rect 10144 7669 10200 7725
rect 10200 7669 10204 7725
rect 10140 7665 10204 7669
rect 10388 7725 10452 7729
rect 10388 7669 10392 7725
rect 10392 7669 10448 7725
rect 10448 7669 10452 7725
rect 10388 7665 10452 7669
rect 10685 7725 10749 7729
rect 10685 7669 10689 7725
rect 10689 7669 10745 7725
rect 10745 7669 10749 7725
rect 10685 7665 10749 7669
rect 11029 7727 11093 7731
rect 11029 7671 11033 7727
rect 11033 7671 11089 7727
rect 11089 7671 11093 7727
rect 11029 7667 11093 7671
rect 11348 7727 11412 7731
rect 11348 7671 11352 7727
rect 11352 7671 11408 7727
rect 11408 7671 11412 7727
rect 11348 7667 11412 7671
rect 11960 7736 12024 7740
rect 11960 7680 11964 7736
rect 11964 7680 12020 7736
rect 12020 7680 12024 7736
rect 11960 7676 12024 7680
rect 12214 7740 12278 7744
rect 12214 7684 12218 7740
rect 12218 7684 12274 7740
rect 12274 7684 12278 7740
rect 12214 7680 12278 7684
rect 12926 7711 12990 7715
rect 12926 7655 12930 7711
rect 12930 7655 12986 7711
rect 12986 7655 12990 7711
rect 12926 7651 12990 7655
rect 13351 7743 13415 7747
rect 13351 7687 13355 7743
rect 13355 7687 13411 7743
rect 13411 7687 13415 7743
rect 13351 7683 13415 7687
rect 13591 7704 13655 7768
rect 3062 7489 3126 7493
rect 3891 7555 3955 7560
rect 3891 7499 3894 7555
rect 3894 7499 3950 7555
rect 3950 7499 3955 7555
rect 3891 7496 3955 7499
rect 3971 7555 4035 7560
rect 3971 7499 3974 7555
rect 3974 7499 4030 7555
rect 4030 7499 4035 7555
rect 3971 7496 4035 7499
rect 4051 7555 4115 7560
rect 4051 7499 4054 7555
rect 4054 7499 4110 7555
rect 4110 7499 4115 7555
rect 4051 7496 4115 7499
rect 4131 7555 4195 7560
rect 4131 7499 4134 7555
rect 4134 7499 4190 7555
rect 4190 7499 4195 7555
rect 4131 7496 4195 7499
rect 4211 7555 4275 7560
rect 4211 7499 4214 7555
rect 4214 7499 4270 7555
rect 4270 7499 4275 7555
rect 4211 7496 4275 7499
rect 4291 7555 4355 7560
rect 4291 7499 4294 7555
rect 4294 7499 4350 7555
rect 4350 7499 4355 7555
rect 4291 7496 4355 7499
rect 4497 7555 4561 7560
rect 4497 7499 4502 7555
rect 4502 7499 4558 7555
rect 4558 7499 4561 7555
rect 4497 7496 4561 7499
rect 4577 7555 4641 7560
rect 4577 7499 4582 7555
rect 4582 7499 4638 7555
rect 4638 7499 4641 7555
rect 4577 7496 4641 7499
rect 4657 7555 4721 7560
rect 4657 7499 4662 7555
rect 4662 7499 4718 7555
rect 4718 7499 4721 7555
rect 4657 7496 4721 7499
rect 4737 7555 4801 7560
rect 4737 7499 4742 7555
rect 4742 7499 4798 7555
rect 4798 7499 4801 7555
rect 4737 7496 4801 7499
rect 4817 7555 4881 7560
rect 4817 7499 4822 7555
rect 4822 7499 4878 7555
rect 4878 7499 4881 7555
rect 4817 7496 4881 7499
rect 4897 7555 4961 7560
rect 4897 7499 4902 7555
rect 4902 7499 4958 7555
rect 4958 7499 4961 7555
rect 4897 7496 4961 7499
rect 5103 7555 5167 7560
rect 5103 7499 5106 7555
rect 5106 7499 5162 7555
rect 5162 7499 5167 7555
rect 5103 7496 5167 7499
rect 5183 7555 5247 7560
rect 5183 7499 5186 7555
rect 5186 7499 5242 7555
rect 5242 7499 5247 7555
rect 5183 7496 5247 7499
rect 5263 7555 5327 7560
rect 5263 7499 5266 7555
rect 5266 7499 5322 7555
rect 5322 7499 5327 7555
rect 5263 7496 5327 7499
rect 5343 7555 5407 7560
rect 5343 7499 5346 7555
rect 5346 7499 5402 7555
rect 5402 7499 5407 7555
rect 5343 7496 5407 7499
rect 5423 7555 5487 7560
rect 5423 7499 5426 7555
rect 5426 7499 5482 7555
rect 5482 7499 5487 7555
rect 5423 7496 5487 7499
rect 5503 7555 5567 7560
rect 5503 7499 5506 7555
rect 5506 7499 5562 7555
rect 5562 7499 5567 7555
rect 5503 7496 5567 7499
rect 5709 7555 5773 7560
rect 5709 7499 5714 7555
rect 5714 7499 5770 7555
rect 5770 7499 5773 7555
rect 5709 7496 5773 7499
rect 5789 7555 5853 7560
rect 5789 7499 5794 7555
rect 5794 7499 5850 7555
rect 5850 7499 5853 7555
rect 5789 7496 5853 7499
rect 5869 7555 5933 7560
rect 5869 7499 5874 7555
rect 5874 7499 5930 7555
rect 5930 7499 5933 7555
rect 5869 7496 5933 7499
rect 5949 7555 6013 7560
rect 5949 7499 5954 7555
rect 5954 7499 6010 7555
rect 6010 7499 6013 7555
rect 5949 7496 6013 7499
rect 6029 7555 6093 7560
rect 6029 7499 6034 7555
rect 6034 7499 6090 7555
rect 6090 7499 6093 7555
rect 6029 7496 6093 7499
rect 6109 7555 6173 7560
rect 6109 7499 6114 7555
rect 6114 7499 6170 7555
rect 6170 7499 6173 7555
rect 6109 7496 6173 7499
rect 6315 7555 6379 7560
rect 6315 7499 6318 7555
rect 6318 7499 6374 7555
rect 6374 7499 6379 7555
rect 6315 7496 6379 7499
rect 6395 7555 6459 7560
rect 6395 7499 6398 7555
rect 6398 7499 6454 7555
rect 6454 7499 6459 7555
rect 6395 7496 6459 7499
rect 6475 7555 6539 7560
rect 6475 7499 6478 7555
rect 6478 7499 6534 7555
rect 6534 7499 6539 7555
rect 6475 7496 6539 7499
rect 6555 7555 6619 7560
rect 6555 7499 6558 7555
rect 6558 7499 6614 7555
rect 6614 7499 6619 7555
rect 6555 7496 6619 7499
rect 6635 7555 6699 7560
rect 6635 7499 6638 7555
rect 6638 7499 6694 7555
rect 6694 7499 6699 7555
rect 6635 7496 6699 7499
rect 6715 7555 6779 7560
rect 6715 7499 6718 7555
rect 6718 7499 6774 7555
rect 6774 7499 6779 7555
rect 6715 7496 6779 7499
rect 6921 7555 6985 7560
rect 6921 7499 6926 7555
rect 6926 7499 6982 7555
rect 6982 7499 6985 7555
rect 6921 7496 6985 7499
rect 7001 7555 7065 7560
rect 7001 7499 7006 7555
rect 7006 7499 7062 7555
rect 7062 7499 7065 7555
rect 7001 7496 7065 7499
rect 7081 7555 7145 7560
rect 7081 7499 7086 7555
rect 7086 7499 7142 7555
rect 7142 7499 7145 7555
rect 7081 7496 7145 7499
rect 7161 7555 7225 7560
rect 7161 7499 7166 7555
rect 7166 7499 7222 7555
rect 7222 7499 7225 7555
rect 7161 7496 7225 7499
rect 7241 7555 7305 7560
rect 7241 7499 7246 7555
rect 7246 7499 7302 7555
rect 7302 7499 7305 7555
rect 7241 7496 7305 7499
rect 7321 7555 7385 7560
rect 7321 7499 7326 7555
rect 7326 7499 7382 7555
rect 7382 7499 7385 7555
rect 7321 7496 7385 7499
rect 7527 7555 7591 7560
rect 7527 7499 7530 7555
rect 7530 7499 7586 7555
rect 7586 7499 7591 7555
rect 7527 7496 7591 7499
rect 7607 7555 7671 7560
rect 7607 7499 7610 7555
rect 7610 7499 7666 7555
rect 7666 7499 7671 7555
rect 7607 7496 7671 7499
rect 7687 7555 7751 7560
rect 7687 7499 7690 7555
rect 7690 7499 7746 7555
rect 7746 7499 7751 7555
rect 7687 7496 7751 7499
rect 7767 7555 7831 7560
rect 7767 7499 7770 7555
rect 7770 7499 7826 7555
rect 7826 7499 7831 7555
rect 7767 7496 7831 7499
rect 7847 7555 7911 7560
rect 7847 7499 7850 7555
rect 7850 7499 7906 7555
rect 7906 7499 7911 7555
rect 7847 7496 7911 7499
rect 7927 7555 7991 7560
rect 7927 7499 7930 7555
rect 7930 7499 7986 7555
rect 7986 7499 7991 7555
rect 7927 7496 7991 7499
rect 8133 7555 8197 7560
rect 8133 7499 8138 7555
rect 8138 7499 8194 7555
rect 8194 7499 8197 7555
rect 8133 7496 8197 7499
rect 8213 7555 8277 7560
rect 8213 7499 8218 7555
rect 8218 7499 8274 7555
rect 8274 7499 8277 7555
rect 8213 7496 8277 7499
rect 8293 7555 8357 7560
rect 8293 7499 8298 7555
rect 8298 7499 8354 7555
rect 8354 7499 8357 7555
rect 8293 7496 8357 7499
rect 8373 7555 8437 7560
rect 8373 7499 8378 7555
rect 8378 7499 8434 7555
rect 8434 7499 8437 7555
rect 8373 7496 8437 7499
rect 8453 7555 8517 7560
rect 8453 7499 8458 7555
rect 8458 7499 8514 7555
rect 8514 7499 8517 7555
rect 8453 7496 8517 7499
rect 8533 7555 8597 7560
rect 8533 7499 8538 7555
rect 8538 7499 8594 7555
rect 8594 7499 8597 7555
rect 8533 7496 8597 7499
rect 8871 7611 8935 7615
rect 8871 7555 8875 7611
rect 8875 7555 8931 7611
rect 8931 7555 8935 7611
rect 8871 7551 8935 7555
rect 11970 7591 12034 7595
rect 11970 7535 11974 7591
rect 11974 7535 12030 7591
rect 12030 7535 12034 7591
rect 11970 7531 12034 7535
rect 12222 7594 12286 7598
rect 12222 7538 12226 7594
rect 12226 7538 12282 7594
rect 12282 7538 12286 7594
rect 12222 7534 12286 7538
rect 13356 7599 13420 7603
rect 13356 7543 13360 7599
rect 13360 7543 13416 7599
rect 13416 7543 13420 7599
rect 13356 7539 13420 7543
rect 14197 8424 14261 8488
rect 14197 8344 14261 8408
rect 14197 8264 14261 8328
rect 14197 8184 14261 8248
rect 14197 8104 14261 8168
rect 14197 8024 14261 8088
rect 14197 7944 14261 8008
rect 14197 7864 14261 7928
rect 14197 7784 14261 7848
rect 14197 7704 14261 7768
rect 14803 8424 14867 8488
rect 14803 8344 14867 8408
rect 14803 8264 14867 8328
rect 14803 8184 14867 8248
rect 14803 8104 14867 8168
rect 14803 8024 14867 8088
rect 14803 7944 14867 8008
rect 14803 7864 14867 7928
rect 14803 7784 14867 7848
rect 14803 7704 14867 7768
rect 15409 8424 15473 8488
rect 15409 8344 15473 8408
rect 15409 8264 15473 8328
rect 15409 8184 15473 8248
rect 15409 8104 15473 8168
rect 15409 8024 15473 8088
rect 15409 7944 15473 8008
rect 15409 7864 15473 7928
rect 15409 7784 15473 7848
rect 15409 7704 15473 7768
rect 16015 8424 16079 8488
rect 16015 8344 16079 8408
rect 16015 8264 16079 8328
rect 16015 8184 16079 8248
rect 16015 8104 16079 8168
rect 16015 8024 16079 8088
rect 16015 7944 16079 8008
rect 16015 7864 16079 7928
rect 16015 7784 16079 7848
rect 16015 7704 16079 7768
rect 16621 8424 16685 8488
rect 16621 8344 16685 8408
rect 16621 8264 16685 8328
rect 16621 8184 16685 8248
rect 16621 8104 16685 8168
rect 16621 8024 16685 8088
rect 16621 7944 16685 8008
rect 16621 7864 16685 7928
rect 16621 7784 16685 7848
rect 16621 7704 16685 7768
rect 17227 8424 17291 8488
rect 17227 8344 17291 8408
rect 17227 8264 17291 8328
rect 17227 8184 17291 8248
rect 17227 8104 17291 8168
rect 17227 8024 17291 8088
rect 17227 7944 17291 8008
rect 17227 7864 17291 7928
rect 17227 7784 17291 7848
rect 17227 7704 17291 7768
rect 17833 8424 17897 8488
rect 17833 8344 17897 8408
rect 17833 8264 17897 8328
rect 17833 8184 17897 8248
rect 17833 8104 17897 8168
rect 17833 8024 17897 8088
rect 17833 7944 17897 8008
rect 17833 7864 17897 7928
rect 17833 7784 17897 7848
rect 17833 7704 17897 7768
rect 18439 8424 18503 8488
rect 18439 8344 18503 8408
rect 18439 8264 18503 8328
rect 18439 8184 18503 8248
rect 18439 8104 18503 8168
rect 18439 8024 18503 8088
rect 18439 7944 18503 8008
rect 18439 7864 18503 7928
rect 18439 7784 18503 7848
rect 18439 7704 18503 7768
rect 18668 8670 18679 8711
rect 18679 8670 18732 8711
rect 18668 8647 18732 8670
rect 18748 8647 18812 8711
rect 18828 8647 18892 8711
rect 18908 8647 18972 8711
rect 18988 8647 19052 8711
rect 19068 8647 19132 8711
rect 18565 8427 18629 8491
rect 18565 8347 18629 8411
rect 18565 8267 18629 8331
rect 18565 8187 18629 8251
rect 18565 8107 18629 8171
rect 18565 8027 18629 8091
rect 18565 7947 18629 8011
rect 18565 7867 18629 7931
rect 18565 7787 18629 7851
rect 18565 7707 18629 7771
rect 19501 8688 19565 8692
rect 19501 8632 19505 8688
rect 19505 8632 19561 8688
rect 19561 8632 19565 8688
rect 19501 8628 19565 8632
rect 19644 8688 19708 8692
rect 19644 8632 19648 8688
rect 19648 8632 19704 8688
rect 19704 8632 19708 8688
rect 19644 8628 19708 8632
rect 19764 8688 19828 8692
rect 19764 8632 19768 8688
rect 19768 8632 19824 8688
rect 19824 8632 19828 8688
rect 19764 8628 19828 8632
rect 20054 8725 20118 8729
rect 20054 8669 20058 8725
rect 20058 8669 20114 8725
rect 20114 8669 20118 8725
rect 20054 8665 20118 8669
rect 20403 8644 20467 8708
rect 20483 8644 20547 8708
rect 20563 8644 20627 8708
rect 20643 8644 20707 8708
rect 20723 8644 20787 8708
rect 20803 8667 20856 8708
rect 20856 8667 20867 8708
rect 20803 8644 20867 8667
rect 21009 8667 21020 8708
rect 21020 8667 21073 8708
rect 21009 8644 21073 8667
rect 21089 8644 21153 8708
rect 21169 8644 21233 8708
rect 21249 8644 21313 8708
rect 21329 8644 21393 8708
rect 21409 8644 21473 8708
rect 21615 8644 21679 8708
rect 21695 8644 21759 8708
rect 21775 8644 21839 8708
rect 21855 8644 21919 8708
rect 21935 8644 21999 8708
rect 22015 8667 22068 8708
rect 22068 8667 22079 8708
rect 22015 8644 22079 8667
rect 22221 8667 22232 8708
rect 22232 8667 22285 8708
rect 22221 8644 22285 8667
rect 22301 8644 22365 8708
rect 22381 8644 22445 8708
rect 22461 8644 22525 8708
rect 22541 8644 22605 8708
rect 22621 8644 22685 8708
rect 22827 8644 22891 8708
rect 22907 8644 22971 8708
rect 22987 8644 23051 8708
rect 23067 8644 23131 8708
rect 23147 8644 23211 8708
rect 23227 8667 23280 8708
rect 23280 8667 23291 8708
rect 23227 8644 23291 8667
rect 23433 8667 23444 8708
rect 23444 8667 23497 8708
rect 23433 8644 23497 8667
rect 23513 8644 23577 8708
rect 23593 8644 23657 8708
rect 23673 8644 23737 8708
rect 23753 8644 23817 8708
rect 23833 8644 23897 8708
rect 24039 8644 24103 8708
rect 24119 8644 24183 8708
rect 24199 8644 24263 8708
rect 24279 8644 24343 8708
rect 24359 8644 24423 8708
rect 24439 8667 24492 8708
rect 24492 8667 24503 8708
rect 24439 8644 24503 8667
rect 24645 8667 24656 8708
rect 24656 8667 24709 8708
rect 24645 8644 24709 8667
rect 24725 8644 24789 8708
rect 24805 8644 24869 8708
rect 24885 8644 24949 8708
rect 24965 8644 25029 8708
rect 25045 8644 25109 8708
rect 19171 8427 19235 8491
rect 19171 8347 19235 8411
rect 20142 8464 20206 8468
rect 20142 8408 20146 8464
rect 20146 8408 20202 8464
rect 20202 8408 20206 8464
rect 20142 8404 20206 8408
rect 20300 8424 20364 8488
rect 19171 8267 19235 8331
rect 19171 8187 19235 8251
rect 20300 8344 20364 8408
rect 20300 8264 20364 8328
rect 19171 8107 19235 8171
rect 19171 8027 19235 8091
rect 20060 8222 20124 8226
rect 20060 8166 20064 8222
rect 20064 8166 20120 8222
rect 20120 8166 20124 8222
rect 20060 8162 20124 8166
rect 20300 8184 20364 8248
rect 19507 8142 19571 8146
rect 19507 8086 19511 8142
rect 19511 8086 19567 8142
rect 19567 8086 19571 8142
rect 19507 8082 19571 8086
rect 19651 8143 19715 8147
rect 19651 8087 19655 8143
rect 19655 8087 19711 8143
rect 19711 8087 19715 8143
rect 19651 8083 19715 8087
rect 19782 8142 19846 8146
rect 19782 8086 19786 8142
rect 19786 8086 19842 8142
rect 19842 8086 19846 8142
rect 19782 8082 19846 8086
rect 20300 8104 20364 8168
rect 19171 7947 19235 8011
rect 19171 7867 19235 7931
rect 19637 7993 19701 7997
rect 19637 7937 19641 7993
rect 19641 7937 19697 7993
rect 19697 7937 19701 7993
rect 19637 7933 19701 7937
rect 20059 8065 20123 8069
rect 20059 8009 20063 8065
rect 20063 8009 20119 8065
rect 20119 8009 20123 8065
rect 20059 8005 20123 8009
rect 20300 8024 20364 8088
rect 20300 7944 20364 8008
rect 19171 7787 19235 7851
rect 20059 7895 20123 7899
rect 20059 7839 20063 7895
rect 20063 7839 20119 7895
rect 20119 7839 20123 7895
rect 20059 7835 20123 7839
rect 20300 7864 20364 7928
rect 19171 7707 19235 7771
rect 19637 7797 19701 7801
rect 19637 7741 19641 7797
rect 19641 7741 19697 7797
rect 19697 7741 19701 7797
rect 19637 7737 19701 7741
rect 20300 7784 20364 7848
rect 20060 7743 20124 7747
rect 20060 7687 20064 7743
rect 20064 7687 20120 7743
rect 20120 7687 20124 7743
rect 20060 7683 20124 7687
rect 20300 7704 20364 7768
rect 19637 7622 19701 7626
rect 19637 7566 19641 7622
rect 19641 7566 19697 7622
rect 19697 7566 19701 7622
rect 19637 7562 19701 7566
rect 13694 7543 13758 7548
rect 13694 7487 13697 7543
rect 13697 7487 13753 7543
rect 13753 7487 13758 7543
rect 13694 7484 13758 7487
rect 13774 7543 13838 7548
rect 13774 7487 13777 7543
rect 13777 7487 13833 7543
rect 13833 7487 13838 7543
rect 13774 7484 13838 7487
rect 13854 7543 13918 7548
rect 13854 7487 13857 7543
rect 13857 7487 13913 7543
rect 13913 7487 13918 7543
rect 13854 7484 13918 7487
rect 13934 7543 13998 7548
rect 13934 7487 13937 7543
rect 13937 7487 13993 7543
rect 13993 7487 13998 7543
rect 13934 7484 13998 7487
rect 14014 7543 14078 7548
rect 14014 7487 14017 7543
rect 14017 7487 14073 7543
rect 14073 7487 14078 7543
rect 14014 7484 14078 7487
rect 14094 7543 14158 7548
rect 14094 7487 14097 7543
rect 14097 7487 14153 7543
rect 14153 7487 14158 7543
rect 14094 7484 14158 7487
rect 14300 7543 14364 7548
rect 14300 7487 14305 7543
rect 14305 7487 14361 7543
rect 14361 7487 14364 7543
rect 14300 7484 14364 7487
rect 14380 7543 14444 7548
rect 14380 7487 14385 7543
rect 14385 7487 14441 7543
rect 14441 7487 14444 7543
rect 14380 7484 14444 7487
rect 14460 7543 14524 7548
rect 14460 7487 14465 7543
rect 14465 7487 14521 7543
rect 14521 7487 14524 7543
rect 14460 7484 14524 7487
rect 14540 7543 14604 7548
rect 14540 7487 14545 7543
rect 14545 7487 14601 7543
rect 14601 7487 14604 7543
rect 14540 7484 14604 7487
rect 14620 7543 14684 7548
rect 14620 7487 14625 7543
rect 14625 7487 14681 7543
rect 14681 7487 14684 7543
rect 14620 7484 14684 7487
rect 14700 7543 14764 7548
rect 14700 7487 14705 7543
rect 14705 7487 14761 7543
rect 14761 7487 14764 7543
rect 14700 7484 14764 7487
rect 14906 7543 14970 7548
rect 14906 7487 14909 7543
rect 14909 7487 14965 7543
rect 14965 7487 14970 7543
rect 14906 7484 14970 7487
rect 14986 7543 15050 7548
rect 14986 7487 14989 7543
rect 14989 7487 15045 7543
rect 15045 7487 15050 7543
rect 14986 7484 15050 7487
rect 15066 7543 15130 7548
rect 15066 7487 15069 7543
rect 15069 7487 15125 7543
rect 15125 7487 15130 7543
rect 15066 7484 15130 7487
rect 15146 7543 15210 7548
rect 15146 7487 15149 7543
rect 15149 7487 15205 7543
rect 15205 7487 15210 7543
rect 15146 7484 15210 7487
rect 15226 7543 15290 7548
rect 15226 7487 15229 7543
rect 15229 7487 15285 7543
rect 15285 7487 15290 7543
rect 15226 7484 15290 7487
rect 15306 7543 15370 7548
rect 15306 7487 15309 7543
rect 15309 7487 15365 7543
rect 15365 7487 15370 7543
rect 15306 7484 15370 7487
rect 15512 7543 15576 7548
rect 15512 7487 15517 7543
rect 15517 7487 15573 7543
rect 15573 7487 15576 7543
rect 15512 7484 15576 7487
rect 15592 7543 15656 7548
rect 15592 7487 15597 7543
rect 15597 7487 15653 7543
rect 15653 7487 15656 7543
rect 15592 7484 15656 7487
rect 15672 7543 15736 7548
rect 15672 7487 15677 7543
rect 15677 7487 15733 7543
rect 15733 7487 15736 7543
rect 15672 7484 15736 7487
rect 15752 7543 15816 7548
rect 15752 7487 15757 7543
rect 15757 7487 15813 7543
rect 15813 7487 15816 7543
rect 15752 7484 15816 7487
rect 15832 7543 15896 7548
rect 15832 7487 15837 7543
rect 15837 7487 15893 7543
rect 15893 7487 15896 7543
rect 15832 7484 15896 7487
rect 15912 7543 15976 7548
rect 15912 7487 15917 7543
rect 15917 7487 15973 7543
rect 15973 7487 15976 7543
rect 15912 7484 15976 7487
rect 16118 7543 16182 7548
rect 16118 7487 16121 7543
rect 16121 7487 16177 7543
rect 16177 7487 16182 7543
rect 16118 7484 16182 7487
rect 16198 7543 16262 7548
rect 16198 7487 16201 7543
rect 16201 7487 16257 7543
rect 16257 7487 16262 7543
rect 16198 7484 16262 7487
rect 16278 7543 16342 7548
rect 16278 7487 16281 7543
rect 16281 7487 16337 7543
rect 16337 7487 16342 7543
rect 16278 7484 16342 7487
rect 16358 7543 16422 7548
rect 16358 7487 16361 7543
rect 16361 7487 16417 7543
rect 16417 7487 16422 7543
rect 16358 7484 16422 7487
rect 16438 7543 16502 7548
rect 16438 7487 16441 7543
rect 16441 7487 16497 7543
rect 16497 7487 16502 7543
rect 16438 7484 16502 7487
rect 16518 7543 16582 7548
rect 16518 7487 16521 7543
rect 16521 7487 16577 7543
rect 16577 7487 16582 7543
rect 16518 7484 16582 7487
rect 16724 7543 16788 7548
rect 16724 7487 16729 7543
rect 16729 7487 16785 7543
rect 16785 7487 16788 7543
rect 16724 7484 16788 7487
rect 16804 7543 16868 7548
rect 16804 7487 16809 7543
rect 16809 7487 16865 7543
rect 16865 7487 16868 7543
rect 16804 7484 16868 7487
rect 16884 7543 16948 7548
rect 16884 7487 16889 7543
rect 16889 7487 16945 7543
rect 16945 7487 16948 7543
rect 16884 7484 16948 7487
rect 16964 7543 17028 7548
rect 16964 7487 16969 7543
rect 16969 7487 17025 7543
rect 17025 7487 17028 7543
rect 16964 7484 17028 7487
rect 17044 7543 17108 7548
rect 17044 7487 17049 7543
rect 17049 7487 17105 7543
rect 17105 7487 17108 7543
rect 17044 7484 17108 7487
rect 17124 7543 17188 7548
rect 17124 7487 17129 7543
rect 17129 7487 17185 7543
rect 17185 7487 17188 7543
rect 17124 7484 17188 7487
rect 17330 7543 17394 7548
rect 17330 7487 17333 7543
rect 17333 7487 17389 7543
rect 17389 7487 17394 7543
rect 17330 7484 17394 7487
rect 17410 7543 17474 7548
rect 17410 7487 17413 7543
rect 17413 7487 17469 7543
rect 17469 7487 17474 7543
rect 17410 7484 17474 7487
rect 17490 7543 17554 7548
rect 17490 7487 17493 7543
rect 17493 7487 17549 7543
rect 17549 7487 17554 7543
rect 17490 7484 17554 7487
rect 17570 7543 17634 7548
rect 17570 7487 17573 7543
rect 17573 7487 17629 7543
rect 17629 7487 17634 7543
rect 17570 7484 17634 7487
rect 17650 7543 17714 7548
rect 17650 7487 17653 7543
rect 17653 7487 17709 7543
rect 17709 7487 17714 7543
rect 17650 7484 17714 7487
rect 17730 7543 17794 7548
rect 17730 7487 17733 7543
rect 17733 7487 17789 7543
rect 17789 7487 17794 7543
rect 17730 7484 17794 7487
rect 17936 7543 18000 7548
rect 17936 7487 17941 7543
rect 17941 7487 17997 7543
rect 17997 7487 18000 7543
rect 17936 7484 18000 7487
rect 18016 7543 18080 7548
rect 18016 7487 18021 7543
rect 18021 7487 18077 7543
rect 18077 7487 18080 7543
rect 18016 7484 18080 7487
rect 18096 7543 18160 7548
rect 18096 7487 18101 7543
rect 18101 7487 18157 7543
rect 18157 7487 18160 7543
rect 18096 7484 18160 7487
rect 18176 7543 18240 7548
rect 18176 7487 18181 7543
rect 18181 7487 18237 7543
rect 18237 7487 18240 7543
rect 18176 7484 18240 7487
rect 18256 7543 18320 7548
rect 18256 7487 18261 7543
rect 18261 7487 18317 7543
rect 18317 7487 18320 7543
rect 18256 7484 18320 7487
rect 18336 7543 18400 7548
rect 18336 7487 18341 7543
rect 18341 7487 18397 7543
rect 18397 7487 18400 7543
rect 18336 7484 18400 7487
rect 18668 7546 18732 7551
rect 18668 7490 18673 7546
rect 18673 7490 18729 7546
rect 18729 7490 18732 7546
rect 18668 7487 18732 7490
rect 18748 7546 18812 7551
rect 18748 7490 18753 7546
rect 18753 7490 18809 7546
rect 18809 7490 18812 7546
rect 18748 7487 18812 7490
rect 18828 7546 18892 7551
rect 18828 7490 18833 7546
rect 18833 7490 18889 7546
rect 18889 7490 18892 7546
rect 18828 7487 18892 7490
rect 18908 7546 18972 7551
rect 18908 7490 18913 7546
rect 18913 7490 18969 7546
rect 18969 7490 18972 7546
rect 18908 7487 18972 7490
rect 18988 7546 19052 7551
rect 18988 7490 18993 7546
rect 18993 7490 19049 7546
rect 19049 7490 19052 7546
rect 18988 7487 19052 7490
rect 19068 7546 19132 7551
rect 19068 7490 19073 7546
rect 19073 7490 19129 7546
rect 19129 7490 19132 7546
rect 19068 7487 19132 7490
rect 19165 7537 19229 7541
rect 19165 7481 19169 7537
rect 19169 7481 19225 7537
rect 19225 7481 19229 7537
rect 19165 7477 19229 7481
rect 20065 7599 20129 7603
rect 20065 7543 20069 7599
rect 20069 7543 20125 7599
rect 20125 7543 20129 7599
rect 20065 7539 20129 7543
rect 20906 8424 20970 8488
rect 20906 8344 20970 8408
rect 20906 8264 20970 8328
rect 20906 8184 20970 8248
rect 20906 8104 20970 8168
rect 20906 8024 20970 8088
rect 20906 7944 20970 8008
rect 20906 7864 20970 7928
rect 20906 7784 20970 7848
rect 20906 7704 20970 7768
rect 21512 8424 21576 8488
rect 21512 8344 21576 8408
rect 21512 8264 21576 8328
rect 21512 8184 21576 8248
rect 21512 8104 21576 8168
rect 21512 8024 21576 8088
rect 21512 7944 21576 8008
rect 21512 7864 21576 7928
rect 21512 7784 21576 7848
rect 21512 7704 21576 7768
rect 22118 8424 22182 8488
rect 22118 8344 22182 8408
rect 22118 8264 22182 8328
rect 22118 8184 22182 8248
rect 22118 8104 22182 8168
rect 22118 8024 22182 8088
rect 22118 7944 22182 8008
rect 22118 7864 22182 7928
rect 22118 7784 22182 7848
rect 22118 7704 22182 7768
rect 22724 8424 22788 8488
rect 22724 8344 22788 8408
rect 22724 8264 22788 8328
rect 22724 8184 22788 8248
rect 22724 8104 22788 8168
rect 22724 8024 22788 8088
rect 22724 7944 22788 8008
rect 22724 7864 22788 7928
rect 22724 7784 22788 7848
rect 22724 7704 22788 7768
rect 23330 8424 23394 8488
rect 23330 8344 23394 8408
rect 23330 8264 23394 8328
rect 23330 8184 23394 8248
rect 23330 8104 23394 8168
rect 23330 8024 23394 8088
rect 23330 7944 23394 8008
rect 23330 7864 23394 7928
rect 23330 7784 23394 7848
rect 23330 7704 23394 7768
rect 23936 8424 24000 8488
rect 23936 8344 24000 8408
rect 23936 8264 24000 8328
rect 23936 8184 24000 8248
rect 23936 8104 24000 8168
rect 23936 8024 24000 8088
rect 23936 7944 24000 8008
rect 23936 7864 24000 7928
rect 23936 7784 24000 7848
rect 23936 7704 24000 7768
rect 24542 8424 24606 8488
rect 24542 8344 24606 8408
rect 24542 8264 24606 8328
rect 24542 8184 24606 8248
rect 24542 8104 24606 8168
rect 24542 8024 24606 8088
rect 24542 7944 24606 8008
rect 24542 7864 24606 7928
rect 24542 7784 24606 7848
rect 24542 7704 24606 7768
rect 25148 8424 25212 8488
rect 25148 8344 25212 8408
rect 25148 8264 25212 8328
rect 25148 8184 25212 8248
rect 25148 8104 25212 8168
rect 25148 8024 25212 8088
rect 25148 7944 25212 8008
rect 25148 7864 25212 7928
rect 25148 7784 25212 7848
rect 25148 7704 25212 7768
rect 25377 8670 25388 8711
rect 25388 8670 25441 8711
rect 25377 8647 25441 8670
rect 25457 8647 25521 8711
rect 25537 8647 25601 8711
rect 25617 8647 25681 8711
rect 25697 8647 25761 8711
rect 25777 8647 25841 8711
rect 25274 8427 25338 8491
rect 25274 8347 25338 8411
rect 25274 8267 25338 8331
rect 25274 8187 25338 8251
rect 25274 8107 25338 8171
rect 25274 8027 25338 8091
rect 25274 7947 25338 8011
rect 25274 7867 25338 7931
rect 25274 7787 25338 7851
rect 25274 7707 25338 7771
rect 26210 8688 26274 8692
rect 26210 8632 26214 8688
rect 26214 8632 26270 8688
rect 26270 8632 26274 8688
rect 26210 8628 26274 8632
rect 26353 8688 26417 8692
rect 26353 8632 26357 8688
rect 26357 8632 26413 8688
rect 26413 8632 26417 8688
rect 26353 8628 26417 8632
rect 26473 8688 26537 8692
rect 26473 8632 26477 8688
rect 26477 8632 26533 8688
rect 26533 8632 26537 8688
rect 26473 8628 26537 8632
rect 25880 8427 25944 8491
rect 25880 8347 25944 8411
rect 25880 8267 25944 8331
rect 25880 8187 25944 8251
rect 25880 8107 25944 8171
rect 25880 8027 25944 8091
rect 26216 8142 26280 8146
rect 26216 8086 26220 8142
rect 26220 8086 26276 8142
rect 26276 8086 26280 8142
rect 26216 8082 26280 8086
rect 26360 8143 26424 8147
rect 26360 8087 26364 8143
rect 26364 8087 26420 8143
rect 26420 8087 26424 8143
rect 26360 8083 26424 8087
rect 26491 8142 26555 8146
rect 26491 8086 26495 8142
rect 26495 8086 26551 8142
rect 26551 8086 26555 8142
rect 26491 8082 26555 8086
rect 25880 7947 25944 8011
rect 25880 7867 25944 7931
rect 25880 7787 25944 7851
rect 25880 7707 25944 7771
rect 20403 7543 20467 7548
rect 20403 7487 20406 7543
rect 20406 7487 20462 7543
rect 20462 7487 20467 7543
rect 20403 7484 20467 7487
rect 20483 7543 20547 7548
rect 20483 7487 20486 7543
rect 20486 7487 20542 7543
rect 20542 7487 20547 7543
rect 20483 7484 20547 7487
rect 20563 7543 20627 7548
rect 20563 7487 20566 7543
rect 20566 7487 20622 7543
rect 20622 7487 20627 7543
rect 20563 7484 20627 7487
rect 20643 7543 20707 7548
rect 20643 7487 20646 7543
rect 20646 7487 20702 7543
rect 20702 7487 20707 7543
rect 20643 7484 20707 7487
rect 20723 7543 20787 7548
rect 20723 7487 20726 7543
rect 20726 7487 20782 7543
rect 20782 7487 20787 7543
rect 20723 7484 20787 7487
rect 20803 7543 20867 7548
rect 20803 7487 20806 7543
rect 20806 7487 20862 7543
rect 20862 7487 20867 7543
rect 20803 7484 20867 7487
rect 21009 7543 21073 7548
rect 21009 7487 21014 7543
rect 21014 7487 21070 7543
rect 21070 7487 21073 7543
rect 21009 7484 21073 7487
rect 21089 7543 21153 7548
rect 21089 7487 21094 7543
rect 21094 7487 21150 7543
rect 21150 7487 21153 7543
rect 21089 7484 21153 7487
rect 21169 7543 21233 7548
rect 21169 7487 21174 7543
rect 21174 7487 21230 7543
rect 21230 7487 21233 7543
rect 21169 7484 21233 7487
rect 21249 7543 21313 7548
rect 21249 7487 21254 7543
rect 21254 7487 21310 7543
rect 21310 7487 21313 7543
rect 21249 7484 21313 7487
rect 21329 7543 21393 7548
rect 21329 7487 21334 7543
rect 21334 7487 21390 7543
rect 21390 7487 21393 7543
rect 21329 7484 21393 7487
rect 21409 7543 21473 7548
rect 21409 7487 21414 7543
rect 21414 7487 21470 7543
rect 21470 7487 21473 7543
rect 21409 7484 21473 7487
rect 21615 7543 21679 7548
rect 21615 7487 21618 7543
rect 21618 7487 21674 7543
rect 21674 7487 21679 7543
rect 21615 7484 21679 7487
rect 21695 7543 21759 7548
rect 21695 7487 21698 7543
rect 21698 7487 21754 7543
rect 21754 7487 21759 7543
rect 21695 7484 21759 7487
rect 21775 7543 21839 7548
rect 21775 7487 21778 7543
rect 21778 7487 21834 7543
rect 21834 7487 21839 7543
rect 21775 7484 21839 7487
rect 21855 7543 21919 7548
rect 21855 7487 21858 7543
rect 21858 7487 21914 7543
rect 21914 7487 21919 7543
rect 21855 7484 21919 7487
rect 21935 7543 21999 7548
rect 21935 7487 21938 7543
rect 21938 7487 21994 7543
rect 21994 7487 21999 7543
rect 21935 7484 21999 7487
rect 22015 7543 22079 7548
rect 22015 7487 22018 7543
rect 22018 7487 22074 7543
rect 22074 7487 22079 7543
rect 22015 7484 22079 7487
rect 22221 7543 22285 7548
rect 22221 7487 22226 7543
rect 22226 7487 22282 7543
rect 22282 7487 22285 7543
rect 22221 7484 22285 7487
rect 22301 7543 22365 7548
rect 22301 7487 22306 7543
rect 22306 7487 22362 7543
rect 22362 7487 22365 7543
rect 22301 7484 22365 7487
rect 22381 7543 22445 7548
rect 22381 7487 22386 7543
rect 22386 7487 22442 7543
rect 22442 7487 22445 7543
rect 22381 7484 22445 7487
rect 22461 7543 22525 7548
rect 22461 7487 22466 7543
rect 22466 7487 22522 7543
rect 22522 7487 22525 7543
rect 22461 7484 22525 7487
rect 22541 7543 22605 7548
rect 22541 7487 22546 7543
rect 22546 7487 22602 7543
rect 22602 7487 22605 7543
rect 22541 7484 22605 7487
rect 22621 7543 22685 7548
rect 22621 7487 22626 7543
rect 22626 7487 22682 7543
rect 22682 7487 22685 7543
rect 22621 7484 22685 7487
rect 22827 7543 22891 7548
rect 22827 7487 22830 7543
rect 22830 7487 22886 7543
rect 22886 7487 22891 7543
rect 22827 7484 22891 7487
rect 22907 7543 22971 7548
rect 22907 7487 22910 7543
rect 22910 7487 22966 7543
rect 22966 7487 22971 7543
rect 22907 7484 22971 7487
rect 22987 7543 23051 7548
rect 22987 7487 22990 7543
rect 22990 7487 23046 7543
rect 23046 7487 23051 7543
rect 22987 7484 23051 7487
rect 23067 7543 23131 7548
rect 23067 7487 23070 7543
rect 23070 7487 23126 7543
rect 23126 7487 23131 7543
rect 23067 7484 23131 7487
rect 23147 7543 23211 7548
rect 23147 7487 23150 7543
rect 23150 7487 23206 7543
rect 23206 7487 23211 7543
rect 23147 7484 23211 7487
rect 23227 7543 23291 7548
rect 23227 7487 23230 7543
rect 23230 7487 23286 7543
rect 23286 7487 23291 7543
rect 23227 7484 23291 7487
rect 23433 7543 23497 7548
rect 23433 7487 23438 7543
rect 23438 7487 23494 7543
rect 23494 7487 23497 7543
rect 23433 7484 23497 7487
rect 23513 7543 23577 7548
rect 23513 7487 23518 7543
rect 23518 7487 23574 7543
rect 23574 7487 23577 7543
rect 23513 7484 23577 7487
rect 23593 7543 23657 7548
rect 23593 7487 23598 7543
rect 23598 7487 23654 7543
rect 23654 7487 23657 7543
rect 23593 7484 23657 7487
rect 23673 7543 23737 7548
rect 23673 7487 23678 7543
rect 23678 7487 23734 7543
rect 23734 7487 23737 7543
rect 23673 7484 23737 7487
rect 23753 7543 23817 7548
rect 23753 7487 23758 7543
rect 23758 7487 23814 7543
rect 23814 7487 23817 7543
rect 23753 7484 23817 7487
rect 23833 7543 23897 7548
rect 23833 7487 23838 7543
rect 23838 7487 23894 7543
rect 23894 7487 23897 7543
rect 23833 7484 23897 7487
rect 24039 7543 24103 7548
rect 24039 7487 24042 7543
rect 24042 7487 24098 7543
rect 24098 7487 24103 7543
rect 24039 7484 24103 7487
rect 24119 7543 24183 7548
rect 24119 7487 24122 7543
rect 24122 7487 24178 7543
rect 24178 7487 24183 7543
rect 24119 7484 24183 7487
rect 24199 7543 24263 7548
rect 24199 7487 24202 7543
rect 24202 7487 24258 7543
rect 24258 7487 24263 7543
rect 24199 7484 24263 7487
rect 24279 7543 24343 7548
rect 24279 7487 24282 7543
rect 24282 7487 24338 7543
rect 24338 7487 24343 7543
rect 24279 7484 24343 7487
rect 24359 7543 24423 7548
rect 24359 7487 24362 7543
rect 24362 7487 24418 7543
rect 24418 7487 24423 7543
rect 24359 7484 24423 7487
rect 24439 7543 24503 7548
rect 24439 7487 24442 7543
rect 24442 7487 24498 7543
rect 24498 7487 24503 7543
rect 24439 7484 24503 7487
rect 24645 7543 24709 7548
rect 24645 7487 24650 7543
rect 24650 7487 24706 7543
rect 24706 7487 24709 7543
rect 24645 7484 24709 7487
rect 24725 7543 24789 7548
rect 24725 7487 24730 7543
rect 24730 7487 24786 7543
rect 24786 7487 24789 7543
rect 24725 7484 24789 7487
rect 24805 7543 24869 7548
rect 24805 7487 24810 7543
rect 24810 7487 24866 7543
rect 24866 7487 24869 7543
rect 24805 7484 24869 7487
rect 24885 7543 24949 7548
rect 24885 7487 24890 7543
rect 24890 7487 24946 7543
rect 24946 7487 24949 7543
rect 24885 7484 24949 7487
rect 24965 7543 25029 7548
rect 24965 7487 24970 7543
rect 24970 7487 25026 7543
rect 25026 7487 25029 7543
rect 24965 7484 25029 7487
rect 25045 7543 25109 7548
rect 25045 7487 25050 7543
rect 25050 7487 25106 7543
rect 25106 7487 25109 7543
rect 25045 7484 25109 7487
rect 25377 7546 25441 7551
rect 25377 7490 25382 7546
rect 25382 7490 25438 7546
rect 25438 7490 25441 7546
rect 25377 7487 25441 7490
rect 25457 7546 25521 7551
rect 25457 7490 25462 7546
rect 25462 7490 25518 7546
rect 25518 7490 25521 7546
rect 25457 7487 25521 7490
rect 25537 7546 25601 7551
rect 25537 7490 25542 7546
rect 25542 7490 25598 7546
rect 25598 7490 25601 7546
rect 25537 7487 25601 7490
rect 25617 7546 25681 7551
rect 25617 7490 25622 7546
rect 25622 7490 25678 7546
rect 25678 7490 25681 7546
rect 25617 7487 25681 7490
rect 25697 7546 25761 7551
rect 25697 7490 25702 7546
rect 25702 7490 25758 7546
rect 25758 7490 25761 7546
rect 25697 7487 25761 7490
rect 25777 7546 25841 7551
rect 25777 7490 25782 7546
rect 25782 7490 25838 7546
rect 25838 7490 25841 7546
rect 25777 7487 25841 7490
rect 25874 7537 25938 7541
rect 25874 7481 25878 7537
rect 25878 7481 25934 7537
rect 25934 7481 25938 7537
rect 25874 7477 25938 7481
rect 24675 7331 24739 7335
rect 24675 7275 24679 7331
rect 24679 7275 24735 7331
rect 24735 7275 24739 7331
rect 24675 7271 24739 7275
rect 24772 7322 24836 7325
rect 24772 7266 24775 7322
rect 24775 7266 24831 7322
rect 24831 7266 24836 7322
rect 24772 7261 24836 7266
rect 24852 7322 24916 7325
rect 24852 7266 24855 7322
rect 24855 7266 24911 7322
rect 24911 7266 24916 7322
rect 24852 7261 24916 7266
rect 24932 7322 24996 7325
rect 24932 7266 24935 7322
rect 24935 7266 24991 7322
rect 24991 7266 24996 7322
rect 24932 7261 24996 7266
rect 25012 7322 25076 7325
rect 25012 7266 25015 7322
rect 25015 7266 25071 7322
rect 25071 7266 25076 7322
rect 25012 7261 25076 7266
rect 25092 7322 25156 7325
rect 25092 7266 25095 7322
rect 25095 7266 25151 7322
rect 25151 7266 25156 7322
rect 25092 7261 25156 7266
rect 25172 7322 25236 7325
rect 25172 7266 25175 7322
rect 25175 7266 25231 7322
rect 25231 7266 25236 7322
rect 25172 7261 25236 7266
rect 25504 7325 25568 7328
rect 25504 7269 25507 7325
rect 25507 7269 25563 7325
rect 25563 7269 25568 7325
rect 25504 7264 25568 7269
rect 25584 7325 25648 7328
rect 25584 7269 25587 7325
rect 25587 7269 25643 7325
rect 25643 7269 25648 7325
rect 25584 7264 25648 7269
rect 25664 7325 25728 7328
rect 25664 7269 25667 7325
rect 25667 7269 25723 7325
rect 25723 7269 25728 7325
rect 25664 7264 25728 7269
rect 25744 7325 25808 7328
rect 25744 7269 25747 7325
rect 25747 7269 25803 7325
rect 25803 7269 25808 7325
rect 25744 7264 25808 7269
rect 25824 7325 25888 7328
rect 25824 7269 25827 7325
rect 25827 7269 25883 7325
rect 25883 7269 25888 7325
rect 25824 7264 25888 7269
rect 25904 7325 25968 7328
rect 25904 7269 25907 7325
rect 25907 7269 25963 7325
rect 25963 7269 25968 7325
rect 25904 7264 25968 7269
rect 26110 7325 26174 7328
rect 26110 7269 26115 7325
rect 26115 7269 26171 7325
rect 26171 7269 26174 7325
rect 26110 7264 26174 7269
rect 26190 7325 26254 7328
rect 26190 7269 26195 7325
rect 26195 7269 26251 7325
rect 26251 7269 26254 7325
rect 26190 7264 26254 7269
rect 26270 7325 26334 7328
rect 26270 7269 26275 7325
rect 26275 7269 26331 7325
rect 26331 7269 26334 7325
rect 26270 7264 26334 7269
rect 26350 7325 26414 7328
rect 26350 7269 26355 7325
rect 26355 7269 26411 7325
rect 26411 7269 26414 7325
rect 26350 7264 26414 7269
rect 26430 7325 26494 7328
rect 26430 7269 26435 7325
rect 26435 7269 26491 7325
rect 26491 7269 26494 7325
rect 26430 7264 26494 7269
rect 26510 7325 26574 7328
rect 26510 7269 26515 7325
rect 26515 7269 26571 7325
rect 26571 7269 26574 7325
rect 26510 7264 26574 7269
rect 26716 7325 26780 7328
rect 26716 7269 26719 7325
rect 26719 7269 26775 7325
rect 26775 7269 26780 7325
rect 26716 7264 26780 7269
rect 26796 7325 26860 7328
rect 26796 7269 26799 7325
rect 26799 7269 26855 7325
rect 26855 7269 26860 7325
rect 26796 7264 26860 7269
rect 26876 7325 26940 7328
rect 26876 7269 26879 7325
rect 26879 7269 26935 7325
rect 26935 7269 26940 7325
rect 26876 7264 26940 7269
rect 26956 7325 27020 7328
rect 26956 7269 26959 7325
rect 26959 7269 27015 7325
rect 27015 7269 27020 7325
rect 26956 7264 27020 7269
rect 27036 7325 27100 7328
rect 27036 7269 27039 7325
rect 27039 7269 27095 7325
rect 27095 7269 27100 7325
rect 27036 7264 27100 7269
rect 27116 7325 27180 7328
rect 27116 7269 27119 7325
rect 27119 7269 27175 7325
rect 27175 7269 27180 7325
rect 27116 7264 27180 7269
rect 27322 7325 27386 7328
rect 27322 7269 27327 7325
rect 27327 7269 27383 7325
rect 27383 7269 27386 7325
rect 27322 7264 27386 7269
rect 27402 7325 27466 7328
rect 27402 7269 27407 7325
rect 27407 7269 27463 7325
rect 27463 7269 27466 7325
rect 27402 7264 27466 7269
rect 27482 7325 27546 7328
rect 27482 7269 27487 7325
rect 27487 7269 27543 7325
rect 27543 7269 27546 7325
rect 27482 7264 27546 7269
rect 27562 7325 27626 7328
rect 27562 7269 27567 7325
rect 27567 7269 27623 7325
rect 27623 7269 27626 7325
rect 27562 7264 27626 7269
rect 27642 7325 27706 7328
rect 27642 7269 27647 7325
rect 27647 7269 27703 7325
rect 27703 7269 27706 7325
rect 27642 7264 27706 7269
rect 27722 7325 27786 7328
rect 27722 7269 27727 7325
rect 27727 7269 27783 7325
rect 27783 7269 27786 7325
rect 27722 7264 27786 7269
rect 27928 7325 27992 7328
rect 27928 7269 27931 7325
rect 27931 7269 27987 7325
rect 27987 7269 27992 7325
rect 27928 7264 27992 7269
rect 28008 7325 28072 7328
rect 28008 7269 28011 7325
rect 28011 7269 28067 7325
rect 28067 7269 28072 7325
rect 28008 7264 28072 7269
rect 28088 7325 28152 7328
rect 28088 7269 28091 7325
rect 28091 7269 28147 7325
rect 28147 7269 28152 7325
rect 28088 7264 28152 7269
rect 28168 7325 28232 7328
rect 28168 7269 28171 7325
rect 28171 7269 28227 7325
rect 28227 7269 28232 7325
rect 28168 7264 28232 7269
rect 28248 7325 28312 7328
rect 28248 7269 28251 7325
rect 28251 7269 28307 7325
rect 28307 7269 28312 7325
rect 28248 7264 28312 7269
rect 28328 7325 28392 7328
rect 28328 7269 28331 7325
rect 28331 7269 28387 7325
rect 28387 7269 28392 7325
rect 28328 7264 28392 7269
rect 28534 7325 28598 7328
rect 28534 7269 28539 7325
rect 28539 7269 28595 7325
rect 28595 7269 28598 7325
rect 28534 7264 28598 7269
rect 28614 7325 28678 7328
rect 28614 7269 28619 7325
rect 28619 7269 28675 7325
rect 28675 7269 28678 7325
rect 28614 7264 28678 7269
rect 28694 7325 28758 7328
rect 28694 7269 28699 7325
rect 28699 7269 28755 7325
rect 28755 7269 28758 7325
rect 28694 7264 28758 7269
rect 28774 7325 28838 7328
rect 28774 7269 28779 7325
rect 28779 7269 28835 7325
rect 28835 7269 28838 7325
rect 28774 7264 28838 7269
rect 28854 7325 28918 7328
rect 28854 7269 28859 7325
rect 28859 7269 28915 7325
rect 28915 7269 28918 7325
rect 28854 7264 28918 7269
rect 28934 7325 28998 7328
rect 28934 7269 28939 7325
rect 28939 7269 28995 7325
rect 28995 7269 28998 7325
rect 28934 7264 28998 7269
rect 29140 7325 29204 7328
rect 29140 7269 29143 7325
rect 29143 7269 29199 7325
rect 29199 7269 29204 7325
rect 29140 7264 29204 7269
rect 29220 7325 29284 7328
rect 29220 7269 29223 7325
rect 29223 7269 29279 7325
rect 29279 7269 29284 7325
rect 29220 7264 29284 7269
rect 29300 7325 29364 7328
rect 29300 7269 29303 7325
rect 29303 7269 29359 7325
rect 29359 7269 29364 7325
rect 29300 7264 29364 7269
rect 29380 7325 29444 7328
rect 29380 7269 29383 7325
rect 29383 7269 29439 7325
rect 29439 7269 29444 7325
rect 29380 7264 29444 7269
rect 29460 7325 29524 7328
rect 29460 7269 29463 7325
rect 29463 7269 29519 7325
rect 29519 7269 29524 7325
rect 29460 7264 29524 7269
rect 29540 7325 29604 7328
rect 29540 7269 29543 7325
rect 29543 7269 29599 7325
rect 29599 7269 29604 7325
rect 29540 7264 29604 7269
rect 29746 7325 29810 7328
rect 29746 7269 29751 7325
rect 29751 7269 29807 7325
rect 29807 7269 29810 7325
rect 29746 7264 29810 7269
rect 29826 7325 29890 7328
rect 29826 7269 29831 7325
rect 29831 7269 29887 7325
rect 29887 7269 29890 7325
rect 29826 7264 29890 7269
rect 29906 7325 29970 7328
rect 29906 7269 29911 7325
rect 29911 7269 29967 7325
rect 29967 7269 29970 7325
rect 29906 7264 29970 7269
rect 29986 7325 30050 7328
rect 29986 7269 29991 7325
rect 29991 7269 30047 7325
rect 30047 7269 30050 7325
rect 29986 7264 30050 7269
rect 30066 7325 30130 7328
rect 30066 7269 30071 7325
rect 30071 7269 30127 7325
rect 30127 7269 30130 7325
rect 30066 7264 30130 7269
rect 30146 7325 30210 7328
rect 30146 7269 30151 7325
rect 30151 7269 30207 7325
rect 30207 7269 30210 7325
rect 30146 7264 30210 7269
rect 10891 6934 11041 7080
rect 11203 6918 11353 7064
rect 24669 7041 24733 7105
rect 24669 6961 24733 7025
rect 24669 6881 24733 6945
rect 24669 6801 24733 6865
rect 24058 6726 24122 6730
rect 24058 6670 24062 6726
rect 24062 6670 24118 6726
rect 24118 6670 24122 6726
rect 24058 6666 24122 6670
rect 24189 6725 24253 6729
rect 24189 6669 24193 6725
rect 24193 6669 24249 6725
rect 24249 6669 24253 6725
rect 24189 6665 24253 6669
rect 24333 6726 24397 6730
rect 24333 6670 24337 6726
rect 24337 6670 24393 6726
rect 24393 6670 24397 6726
rect 24333 6666 24397 6670
rect 24669 6721 24733 6785
rect 24669 6641 24733 6705
rect 24669 6561 24733 6625
rect 24669 6481 24733 6545
rect 23609 6320 23759 6466
rect 24669 6401 24733 6465
rect 24669 6321 24733 6385
rect 10955 5974 11105 6120
rect 11261 5986 11411 6132
rect 24076 6180 24140 6184
rect 24076 6124 24080 6180
rect 24080 6124 24136 6180
rect 24136 6124 24140 6180
rect 24076 6120 24140 6124
rect 24196 6180 24260 6184
rect 24196 6124 24200 6180
rect 24200 6124 24256 6180
rect 24256 6124 24260 6180
rect 24196 6120 24260 6124
rect 24339 6180 24403 6184
rect 24339 6124 24343 6180
rect 24343 6124 24399 6180
rect 24399 6124 24403 6180
rect 24339 6120 24403 6124
rect 25275 7041 25339 7105
rect 25275 6961 25339 7025
rect 25275 6881 25339 6945
rect 25275 6801 25339 6865
rect 25275 6721 25339 6785
rect 25275 6641 25339 6705
rect 25275 6561 25339 6625
rect 25275 6481 25339 6545
rect 25275 6401 25339 6465
rect 25275 6321 25339 6385
rect 24772 6101 24836 6165
rect 24852 6101 24916 6165
rect 24932 6101 24996 6165
rect 25012 6101 25076 6165
rect 25092 6101 25156 6165
rect 25172 6142 25236 6165
rect 25172 6101 25225 6142
rect 25225 6101 25236 6142
rect 25401 7044 25465 7108
rect 25401 6964 25465 7028
rect 25401 6884 25465 6948
rect 25401 6804 25465 6868
rect 25401 6724 25465 6788
rect 25401 6644 25465 6708
rect 25401 6564 25465 6628
rect 25401 6484 25465 6548
rect 25401 6404 25465 6468
rect 25401 6324 25465 6388
rect 26007 7044 26071 7108
rect 26007 6964 26071 7028
rect 26007 6884 26071 6948
rect 26007 6804 26071 6868
rect 26007 6724 26071 6788
rect 26007 6644 26071 6708
rect 26007 6564 26071 6628
rect 26007 6484 26071 6548
rect 26007 6404 26071 6468
rect 26007 6324 26071 6388
rect 26613 7044 26677 7108
rect 26613 6964 26677 7028
rect 26613 6884 26677 6948
rect 26613 6804 26677 6868
rect 26613 6724 26677 6788
rect 26613 6644 26677 6708
rect 26613 6564 26677 6628
rect 26613 6484 26677 6548
rect 26613 6404 26677 6468
rect 26613 6324 26677 6388
rect 27219 7044 27283 7108
rect 27219 6964 27283 7028
rect 27219 6884 27283 6948
rect 27219 6804 27283 6868
rect 27219 6724 27283 6788
rect 27219 6644 27283 6708
rect 27219 6564 27283 6628
rect 27219 6484 27283 6548
rect 27219 6404 27283 6468
rect 27219 6324 27283 6388
rect 27825 7044 27889 7108
rect 27825 6964 27889 7028
rect 27825 6884 27889 6948
rect 27825 6804 27889 6868
rect 27825 6724 27889 6788
rect 27825 6644 27889 6708
rect 27825 6564 27889 6628
rect 27825 6484 27889 6548
rect 27825 6404 27889 6468
rect 27825 6324 27889 6388
rect 28431 7044 28495 7108
rect 28431 6964 28495 7028
rect 28431 6884 28495 6948
rect 28431 6804 28495 6868
rect 28431 6724 28495 6788
rect 28431 6644 28495 6708
rect 28431 6564 28495 6628
rect 28431 6484 28495 6548
rect 28431 6404 28495 6468
rect 28431 6324 28495 6388
rect 29037 7044 29101 7108
rect 29037 6964 29101 7028
rect 29037 6884 29101 6948
rect 29037 6804 29101 6868
rect 29037 6724 29101 6788
rect 29037 6644 29101 6708
rect 29037 6564 29101 6628
rect 29037 6484 29101 6548
rect 29037 6404 29101 6468
rect 29037 6324 29101 6388
rect 29643 7044 29707 7108
rect 29643 6964 29707 7028
rect 29643 6884 29707 6948
rect 29643 6804 29707 6868
rect 29643 6724 29707 6788
rect 29643 6644 29707 6708
rect 29643 6564 29707 6628
rect 29643 6484 29707 6548
rect 29643 6404 29707 6468
rect 29643 6324 29707 6388
rect 30484 7269 30548 7273
rect 30484 7213 30488 7269
rect 30488 7213 30544 7269
rect 30544 7213 30548 7269
rect 30484 7209 30548 7213
rect 30249 7044 30313 7108
rect 30489 7125 30553 7129
rect 30489 7069 30493 7125
rect 30493 7069 30549 7125
rect 30549 7069 30553 7125
rect 30489 7065 30553 7069
rect 30249 6964 30313 7028
rect 30249 6884 30313 6948
rect 30490 6973 30554 6977
rect 30490 6917 30494 6973
rect 30494 6917 30550 6973
rect 30550 6917 30554 6973
rect 30490 6913 30554 6917
rect 30249 6804 30313 6868
rect 30249 6724 30313 6788
rect 30490 6803 30554 6807
rect 30490 6747 30494 6803
rect 30494 6747 30550 6803
rect 30550 6747 30554 6803
rect 30490 6743 30554 6747
rect 30249 6644 30313 6708
rect 30249 6564 30313 6628
rect 30489 6646 30553 6650
rect 30489 6590 30493 6646
rect 30493 6590 30549 6646
rect 30549 6590 30553 6646
rect 30489 6586 30553 6590
rect 30249 6484 30313 6548
rect 30249 6404 30313 6468
rect 30249 6324 30313 6388
rect 30407 6404 30471 6408
rect 30407 6348 30411 6404
rect 30411 6348 30467 6404
rect 30467 6348 30471 6404
rect 30407 6344 30471 6348
rect 30784 6412 30848 6416
rect 30784 6356 30788 6412
rect 30788 6356 30844 6412
rect 30844 6356 30848 6412
rect 30784 6352 30848 6356
rect 30984 6412 31048 6416
rect 30984 6356 30988 6412
rect 30988 6356 31044 6412
rect 31044 6356 31048 6412
rect 30984 6352 31048 6356
rect 25504 6104 25568 6168
rect 25584 6104 25648 6168
rect 25664 6104 25728 6168
rect 25744 6104 25808 6168
rect 25824 6104 25888 6168
rect 25904 6145 25968 6168
rect 25904 6104 25957 6145
rect 25957 6104 25968 6145
rect 26110 6145 26174 6168
rect 26110 6104 26121 6145
rect 26121 6104 26174 6145
rect 26190 6104 26254 6168
rect 26270 6104 26334 6168
rect 26350 6104 26414 6168
rect 26430 6104 26494 6168
rect 26510 6104 26574 6168
rect 26716 6104 26780 6168
rect 26796 6104 26860 6168
rect 26876 6104 26940 6168
rect 26956 6104 27020 6168
rect 27036 6104 27100 6168
rect 27116 6145 27180 6168
rect 27116 6104 27169 6145
rect 27169 6104 27180 6145
rect 27322 6145 27386 6168
rect 27322 6104 27333 6145
rect 27333 6104 27386 6145
rect 27402 6104 27466 6168
rect 27482 6104 27546 6168
rect 27562 6104 27626 6168
rect 27642 6104 27706 6168
rect 27722 6104 27786 6168
rect 27928 6104 27992 6168
rect 28008 6104 28072 6168
rect 28088 6104 28152 6168
rect 28168 6104 28232 6168
rect 28248 6104 28312 6168
rect 28328 6145 28392 6168
rect 28328 6104 28381 6145
rect 28381 6104 28392 6145
rect 28534 6145 28598 6168
rect 28534 6104 28545 6145
rect 28545 6104 28598 6145
rect 28614 6104 28678 6168
rect 28694 6104 28758 6168
rect 28774 6104 28838 6168
rect 28854 6104 28918 6168
rect 28934 6104 28998 6168
rect 29140 6104 29204 6168
rect 29220 6104 29284 6168
rect 29300 6104 29364 6168
rect 29380 6104 29444 6168
rect 29460 6104 29524 6168
rect 29540 6145 29604 6168
rect 29540 6104 29593 6145
rect 29593 6104 29604 6145
rect 29746 6145 29810 6168
rect 29746 6104 29757 6145
rect 29757 6104 29810 6145
rect 29826 6104 29890 6168
rect 29906 6104 29970 6168
rect 29986 6104 30050 6168
rect 30066 6104 30130 6168
rect 30146 6104 30210 6168
rect 30495 6143 30559 6147
rect 30495 6087 30499 6143
rect 30499 6087 30555 6143
rect 30555 6087 30559 6143
rect 30495 6083 30559 6087
rect 23609 5894 23759 6040
rect 25123 5856 25187 5920
rect 25203 5856 25267 5920
rect 25283 5856 25347 5920
rect 25363 5856 25427 5920
rect 25443 5856 25507 5920
rect 25523 5879 25581 5920
rect 25581 5879 25587 5920
rect 25523 5856 25587 5879
rect 23609 5668 23759 5814
rect 25020 5636 25084 5700
rect 25020 5556 25084 5620
rect 10787 5346 10937 5492
rect 25020 5476 25084 5540
rect 25020 5396 25084 5460
rect 25020 5316 25084 5380
rect 25020 5236 25084 5300
rect 25020 5156 25084 5220
rect 23625 4934 23775 5080
rect 25020 5076 25084 5140
rect 25020 4996 25084 5060
rect 25020 4916 25084 4980
rect 25626 5636 25690 5700
rect 25626 5556 25690 5620
rect 25626 5476 25690 5540
rect 25626 5396 25690 5460
rect 25626 5316 25690 5380
rect 25626 5236 25690 5300
rect 25626 5156 25690 5220
rect 25626 5076 25690 5140
rect 25626 4996 25690 5060
rect 25626 4916 25690 4980
rect 25855 5856 25919 5920
rect 25935 5856 25999 5920
rect 26015 5856 26079 5920
rect 26095 5856 26159 5920
rect 26175 5856 26239 5920
rect 26255 5879 26313 5920
rect 26313 5879 26319 5920
rect 26255 5856 26319 5879
rect 26461 5879 26467 5920
rect 26467 5879 26525 5920
rect 26461 5856 26525 5879
rect 26541 5856 26605 5920
rect 26621 5856 26685 5920
rect 26701 5856 26765 5920
rect 26781 5856 26845 5920
rect 26861 5856 26925 5920
rect 27067 5856 27131 5920
rect 27147 5856 27211 5920
rect 27227 5856 27291 5920
rect 27307 5856 27371 5920
rect 27387 5856 27451 5920
rect 27467 5879 27525 5920
rect 27525 5879 27531 5920
rect 27467 5856 27531 5879
rect 27673 5879 27679 5920
rect 27679 5879 27737 5920
rect 27673 5856 27737 5879
rect 27753 5856 27817 5920
rect 27833 5856 27897 5920
rect 27913 5856 27977 5920
rect 27993 5856 28057 5920
rect 28073 5856 28137 5920
rect 25752 5636 25816 5700
rect 25752 5556 25816 5620
rect 25752 5476 25816 5540
rect 25752 5396 25816 5460
rect 25752 5316 25816 5380
rect 25752 5236 25816 5300
rect 25752 5156 25816 5220
rect 25752 5076 25816 5140
rect 25752 4996 25816 5060
rect 25752 4916 25816 4980
rect 26358 5636 26422 5700
rect 26358 5556 26422 5620
rect 26358 5476 26422 5540
rect 26358 5396 26422 5460
rect 26358 5316 26422 5380
rect 26358 5236 26422 5300
rect 26358 5156 26422 5220
rect 26358 5076 26422 5140
rect 26358 4996 26422 5060
rect 26358 4916 26422 4980
rect 26964 5636 27028 5700
rect 26964 5556 27028 5620
rect 26964 5476 27028 5540
rect 26964 5396 27028 5460
rect 26964 5316 27028 5380
rect 26964 5236 27028 5300
rect 26964 5156 27028 5220
rect 26964 5076 27028 5140
rect 26964 4996 27028 5060
rect 26964 4916 27028 4980
rect 27570 5636 27634 5700
rect 27570 5556 27634 5620
rect 27570 5476 27634 5540
rect 27570 5396 27634 5460
rect 27570 5316 27634 5380
rect 27570 5236 27634 5300
rect 27570 5156 27634 5220
rect 27570 5076 27634 5140
rect 27570 4996 27634 5060
rect 27570 4916 27634 4980
rect 28176 5636 28240 5700
rect 28176 5556 28240 5620
rect 28176 5476 28240 5540
rect 28176 5396 28240 5460
rect 28176 5316 28240 5380
rect 28176 5236 28240 5300
rect 28176 5156 28240 5220
rect 28176 5076 28240 5140
rect 28176 4996 28240 5060
rect 28176 4916 28240 4980
rect 28405 5856 28469 5920
rect 28485 5856 28549 5920
rect 28565 5856 28629 5920
rect 28645 5856 28709 5920
rect 28725 5856 28789 5920
rect 28805 5879 28863 5920
rect 28863 5879 28869 5920
rect 28805 5856 28869 5879
rect 29011 5879 29017 5920
rect 29017 5879 29075 5920
rect 29011 5856 29075 5879
rect 29091 5856 29155 5920
rect 29171 5856 29235 5920
rect 29251 5856 29315 5920
rect 29331 5856 29395 5920
rect 29411 5856 29475 5920
rect 28302 5636 28366 5700
rect 28302 5556 28366 5620
rect 28302 5476 28366 5540
rect 28302 5396 28366 5460
rect 28302 5316 28366 5380
rect 28302 5236 28366 5300
rect 28302 5156 28366 5220
rect 28302 5076 28366 5140
rect 28302 4996 28366 5060
rect 28302 4916 28366 4980
rect 28908 5636 28972 5700
rect 28908 5556 28972 5620
rect 28908 5476 28972 5540
rect 28908 5396 28972 5460
rect 28908 5316 28972 5380
rect 28908 5236 28972 5300
rect 28908 5156 28972 5220
rect 28908 5076 28972 5140
rect 28908 4996 28972 5060
rect 28908 4916 28972 4980
rect 29514 5636 29578 5700
rect 29514 5556 29578 5620
rect 29514 5476 29578 5540
rect 29514 5396 29578 5460
rect 29514 5316 29578 5380
rect 29514 5236 29578 5300
rect 29514 5156 29578 5220
rect 29514 5076 29578 5140
rect 29514 4996 29578 5060
rect 29514 4916 29578 4980
rect 29745 5879 29751 5920
rect 29751 5879 29809 5920
rect 29745 5856 29809 5879
rect 29825 5856 29889 5920
rect 29905 5856 29969 5920
rect 29985 5856 30049 5920
rect 30065 5856 30129 5920
rect 30145 5856 30209 5920
rect 30495 5940 30559 5944
rect 30495 5884 30499 5940
rect 30499 5884 30555 5940
rect 30555 5884 30559 5940
rect 30495 5880 30559 5884
rect 29642 5636 29706 5700
rect 29642 5556 29706 5620
rect 29642 5476 29706 5540
rect 29642 5396 29706 5460
rect 29642 5316 29706 5380
rect 29642 5236 29706 5300
rect 29642 5156 29706 5220
rect 29642 5076 29706 5140
rect 29642 4996 29706 5060
rect 29642 4916 29706 4980
rect 30595 5770 30659 5774
rect 30595 5714 30599 5770
rect 30599 5714 30655 5770
rect 30655 5714 30659 5770
rect 30595 5710 30659 5714
rect 30248 5636 30312 5700
rect 30248 5556 30312 5620
rect 30404 5678 30468 5682
rect 30404 5622 30408 5678
rect 30408 5622 30464 5678
rect 30464 5622 30468 5678
rect 30404 5618 30468 5622
rect 30248 5476 30312 5540
rect 30248 5396 30312 5460
rect 30248 5316 30312 5380
rect 30248 5236 30312 5300
rect 30248 5156 30312 5220
rect 30248 5076 30312 5140
rect 30248 4996 30312 5060
rect 30248 4916 30312 4980
rect 24661 4753 24725 4757
rect 24661 4697 24665 4753
rect 24665 4697 24721 4753
rect 24721 4697 24725 4753
rect 24661 4693 24725 4697
rect 25203 4756 25267 4760
rect 25203 4700 25207 4756
rect 25207 4700 25263 4756
rect 25263 4700 25267 4756
rect 25203 4696 25267 4700
rect 25283 4756 25347 4760
rect 25283 4700 25287 4756
rect 25287 4700 25343 4756
rect 25343 4700 25347 4756
rect 25283 4696 25347 4700
rect 25363 4756 25427 4760
rect 25363 4700 25367 4756
rect 25367 4700 25423 4756
rect 25423 4700 25427 4756
rect 25363 4696 25427 4700
rect 25443 4756 25507 4760
rect 25443 4700 25447 4756
rect 25447 4700 25503 4756
rect 25503 4700 25507 4756
rect 25443 4696 25507 4700
rect 25935 4756 25999 4760
rect 25935 4700 25939 4756
rect 25939 4700 25995 4756
rect 25995 4700 25999 4756
rect 25935 4696 25999 4700
rect 26015 4756 26079 4760
rect 26015 4700 26019 4756
rect 26019 4700 26075 4756
rect 26075 4700 26079 4756
rect 26015 4696 26079 4700
rect 26095 4756 26159 4760
rect 26095 4700 26099 4756
rect 26099 4700 26155 4756
rect 26155 4700 26159 4756
rect 26095 4696 26159 4700
rect 26175 4756 26239 4760
rect 26175 4700 26179 4756
rect 26179 4700 26235 4756
rect 26235 4700 26239 4756
rect 26175 4696 26239 4700
rect 26541 4756 26605 4760
rect 26541 4700 26545 4756
rect 26545 4700 26601 4756
rect 26601 4700 26605 4756
rect 26541 4696 26605 4700
rect 26621 4756 26685 4760
rect 26621 4700 26625 4756
rect 26625 4700 26681 4756
rect 26681 4700 26685 4756
rect 26621 4696 26685 4700
rect 26701 4756 26765 4760
rect 26701 4700 26705 4756
rect 26705 4700 26761 4756
rect 26761 4700 26765 4756
rect 26701 4696 26765 4700
rect 26781 4756 26845 4760
rect 26781 4700 26785 4756
rect 26785 4700 26841 4756
rect 26841 4700 26845 4756
rect 26781 4696 26845 4700
rect 27147 4756 27211 4760
rect 27147 4700 27151 4756
rect 27151 4700 27207 4756
rect 27207 4700 27211 4756
rect 27147 4696 27211 4700
rect 27227 4756 27291 4760
rect 27227 4700 27231 4756
rect 27231 4700 27287 4756
rect 27287 4700 27291 4756
rect 27227 4696 27291 4700
rect 27307 4756 27371 4760
rect 27307 4700 27311 4756
rect 27311 4700 27367 4756
rect 27367 4700 27371 4756
rect 27307 4696 27371 4700
rect 27387 4756 27451 4760
rect 27387 4700 27391 4756
rect 27391 4700 27447 4756
rect 27447 4700 27451 4756
rect 27387 4696 27451 4700
rect 27753 4756 27817 4760
rect 27753 4700 27757 4756
rect 27757 4700 27813 4756
rect 27813 4700 27817 4756
rect 27753 4696 27817 4700
rect 27833 4756 27897 4760
rect 27833 4700 27837 4756
rect 27837 4700 27893 4756
rect 27893 4700 27897 4756
rect 27833 4696 27897 4700
rect 27913 4756 27977 4760
rect 27913 4700 27917 4756
rect 27917 4700 27973 4756
rect 27973 4700 27977 4756
rect 27913 4696 27977 4700
rect 27993 4756 28057 4760
rect 27993 4700 27997 4756
rect 27997 4700 28053 4756
rect 28053 4700 28057 4756
rect 27993 4696 28057 4700
rect 28485 4756 28549 4760
rect 28485 4700 28489 4756
rect 28489 4700 28545 4756
rect 28545 4700 28549 4756
rect 28485 4696 28549 4700
rect 28565 4756 28629 4760
rect 28565 4700 28569 4756
rect 28569 4700 28625 4756
rect 28625 4700 28629 4756
rect 28565 4696 28629 4700
rect 28645 4756 28709 4760
rect 28645 4700 28649 4756
rect 28649 4700 28705 4756
rect 28705 4700 28709 4756
rect 28645 4696 28709 4700
rect 28725 4756 28789 4760
rect 28725 4700 28729 4756
rect 28729 4700 28785 4756
rect 28785 4700 28789 4756
rect 28725 4696 28789 4700
rect 29091 4756 29155 4760
rect 29091 4700 29095 4756
rect 29095 4700 29151 4756
rect 29151 4700 29155 4756
rect 29091 4696 29155 4700
rect 29171 4756 29235 4760
rect 29171 4700 29175 4756
rect 29175 4700 29231 4756
rect 29231 4700 29235 4756
rect 29171 4696 29235 4700
rect 29251 4756 29315 4760
rect 29251 4700 29255 4756
rect 29255 4700 29311 4756
rect 29311 4700 29315 4756
rect 29251 4696 29315 4700
rect 29331 4756 29395 4760
rect 29331 4700 29335 4756
rect 29335 4700 29391 4756
rect 29391 4700 29395 4756
rect 29331 4696 29395 4700
rect 29825 4756 29889 4760
rect 29825 4700 29829 4756
rect 29829 4700 29885 4756
rect 29885 4700 29889 4756
rect 29825 4696 29889 4700
rect 29905 4756 29969 4760
rect 29905 4700 29909 4756
rect 29909 4700 29965 4756
rect 29965 4700 29969 4756
rect 29905 4696 29969 4700
rect 29985 4756 30049 4760
rect 29985 4700 29989 4756
rect 29989 4700 30045 4756
rect 30045 4700 30049 4756
rect 29985 4696 30049 4700
rect 30065 4756 30129 4760
rect 30065 4700 30069 4756
rect 30069 4700 30125 4756
rect 30125 4700 30129 4756
rect 30065 4696 30129 4700
rect 10823 4500 10973 4646
rect 11175 4504 11325 4650
rect 11621 4504 11771 4650
rect 12187 4508 12337 4654
rect 12853 4508 13003 4654
rect 13235 4492 13385 4638
rect 25708 4308 25772 4312
rect 25708 4252 25712 4308
rect 25712 4252 25768 4308
rect 25768 4252 25772 4308
rect 25708 4248 25772 4252
rect 25882 4307 25946 4311
rect 25882 4251 25886 4307
rect 25886 4251 25942 4307
rect 25942 4251 25946 4307
rect 25882 4247 25946 4251
rect 26107 4309 26171 4313
rect 26107 4253 26111 4309
rect 26111 4253 26167 4309
rect 26167 4253 26171 4309
rect 26107 4249 26171 4253
rect 26308 4311 26372 4315
rect 26308 4255 26312 4311
rect 26312 4255 26368 4311
rect 26368 4255 26372 4311
rect 26308 4251 26372 4255
rect 26531 4309 26595 4313
rect 26531 4253 26535 4309
rect 26535 4253 26591 4309
rect 26591 4253 26595 4309
rect 26531 4249 26595 4253
rect 26740 4314 26804 4318
rect 26740 4258 26744 4314
rect 26744 4258 26800 4314
rect 26800 4258 26804 4314
rect 26740 4254 26804 4258
rect 26968 4307 27032 4311
rect 26968 4251 26972 4307
rect 26972 4251 27028 4307
rect 27028 4251 27032 4307
rect 26968 4247 27032 4251
rect 27158 4311 27222 4315
rect 27158 4255 27162 4311
rect 27162 4255 27218 4311
rect 27218 4255 27222 4311
rect 27158 4251 27222 4255
rect 27363 4314 27427 4318
rect 27363 4258 27367 4314
rect 27367 4258 27423 4314
rect 27423 4258 27427 4314
rect 27363 4254 27427 4258
rect 27562 4314 27626 4318
rect 27562 4258 27566 4314
rect 27566 4258 27622 4314
rect 27622 4258 27626 4314
rect 27562 4254 27626 4258
rect 27778 4309 27842 4313
rect 27778 4253 27782 4309
rect 27782 4253 27838 4309
rect 27838 4253 27842 4309
rect 27778 4249 27842 4253
rect 28166 4314 28230 4318
rect 28166 4258 28170 4314
rect 28170 4258 28226 4314
rect 28226 4258 28230 4314
rect 28166 4254 28230 4258
rect 28401 4309 28465 4313
rect 28401 4253 28405 4309
rect 28405 4253 28461 4309
rect 28461 4253 28465 4309
rect 28401 4249 28465 4253
rect 28643 4311 28707 4315
rect 28643 4255 28647 4311
rect 28647 4255 28703 4311
rect 28703 4255 28707 4311
rect 28643 4251 28707 4255
rect 28875 4312 28939 4316
rect 28875 4256 28879 4312
rect 28879 4256 28935 4312
rect 28935 4256 28939 4312
rect 28875 4252 28939 4256
rect 29104 4315 29168 4319
rect 29104 4259 29108 4315
rect 29108 4259 29164 4315
rect 29164 4259 29168 4315
rect 29104 4255 29168 4259
rect 29353 4307 29417 4311
rect 29353 4251 29357 4307
rect 29357 4251 29413 4307
rect 29413 4251 29417 4307
rect 29353 4247 29417 4251
rect 29571 4311 29635 4315
rect 29571 4255 29575 4311
rect 29575 4255 29631 4311
rect 29631 4255 29635 4311
rect 29571 4251 29635 4255
rect 29800 4307 29864 4311
rect 29800 4251 29804 4307
rect 29804 4251 29860 4307
rect 29860 4251 29864 4307
rect 29800 4247 29864 4251
rect 30021 4309 30085 4313
rect 30021 4253 30025 4309
rect 30025 4253 30081 4309
rect 30081 4253 30085 4309
rect 30021 4249 30085 4253
rect 30237 4314 30301 4318
rect 30237 4258 30241 4314
rect 30241 4258 30297 4314
rect 30297 4258 30301 4314
rect 30237 4254 30301 4258
rect 23605 3942 23755 4088
rect 27066 4121 27130 4125
rect 27066 4065 27070 4121
rect 27070 4065 27126 4121
rect 27126 4065 27130 4121
rect 27066 4061 27130 4065
rect 27451 4070 27515 4074
rect 27451 4014 27455 4070
rect 27455 4014 27511 4070
rect 27511 4014 27515 4070
rect 27451 4010 27515 4014
rect 29461 4120 29525 4124
rect 29461 4064 29465 4120
rect 29465 4064 29521 4120
rect 29521 4064 29525 4120
rect 29461 4060 29525 4064
rect 29846 4071 29910 4075
rect 29846 4015 29850 4071
rect 29850 4015 29906 4071
rect 29906 4015 29910 4071
rect 29846 4011 29910 4015
rect 10905 3646 11055 3792
rect 11255 3654 11405 3800
rect 25710 3725 25774 3729
rect 25710 3669 25714 3725
rect 25714 3669 25770 3725
rect 25770 3669 25774 3725
rect 25710 3665 25774 3669
rect 25885 3723 25949 3727
rect 25885 3667 25889 3723
rect 25889 3667 25945 3723
rect 25945 3667 25949 3723
rect 25885 3663 25949 3667
rect 26082 3725 26146 3729
rect 26082 3669 26086 3725
rect 26086 3669 26142 3725
rect 26142 3669 26146 3725
rect 26082 3665 26146 3669
rect 26301 3728 26365 3732
rect 26301 3672 26305 3728
rect 26305 3672 26361 3728
rect 26361 3672 26365 3728
rect 26301 3668 26365 3672
rect 26533 3724 26597 3728
rect 26533 3668 26537 3724
rect 26537 3668 26593 3724
rect 26593 3668 26597 3724
rect 26533 3664 26597 3668
rect 26757 3731 26821 3735
rect 26757 3675 26761 3731
rect 26761 3675 26817 3731
rect 26817 3675 26821 3731
rect 26757 3671 26821 3675
rect 26969 3719 27033 3723
rect 26969 3663 26973 3719
rect 26973 3663 27029 3719
rect 27029 3663 27033 3719
rect 26969 3659 27033 3663
rect 27191 3715 27255 3719
rect 27191 3659 27195 3715
rect 27195 3659 27251 3715
rect 27251 3659 27255 3715
rect 27191 3655 27255 3659
rect 27414 3712 27478 3716
rect 27414 3656 27418 3712
rect 27418 3656 27474 3712
rect 27474 3656 27478 3712
rect 27414 3652 27478 3656
rect 27624 3712 27688 3716
rect 27624 3656 27628 3712
rect 27628 3656 27684 3712
rect 27684 3656 27688 3712
rect 27624 3652 27688 3656
rect 27837 3712 27901 3716
rect 27837 3656 27841 3712
rect 27841 3656 27897 3712
rect 27897 3656 27901 3712
rect 27837 3652 27901 3656
rect 28154 3705 28218 3709
rect 28154 3649 28158 3705
rect 28158 3649 28214 3705
rect 28214 3649 28218 3705
rect 28154 3645 28218 3649
rect 28356 3708 28420 3712
rect 28356 3652 28360 3708
rect 28360 3652 28416 3708
rect 28416 3652 28420 3708
rect 28356 3648 28420 3652
rect 28557 3709 28621 3713
rect 28557 3653 28561 3709
rect 28561 3653 28617 3709
rect 28617 3653 28621 3709
rect 28557 3649 28621 3653
rect 28736 3710 28800 3714
rect 28736 3654 28740 3710
rect 28740 3654 28796 3710
rect 28796 3654 28800 3710
rect 28736 3650 28800 3654
rect 28928 3714 28992 3718
rect 28928 3658 28932 3714
rect 28932 3658 28988 3714
rect 28988 3658 28992 3714
rect 28928 3654 28992 3658
rect 29113 3711 29177 3715
rect 29113 3655 29117 3711
rect 29117 3655 29173 3711
rect 29173 3655 29177 3711
rect 29113 3651 29177 3655
rect 29345 3710 29409 3714
rect 29345 3654 29349 3710
rect 29349 3654 29405 3710
rect 29405 3654 29409 3710
rect 29345 3650 29409 3654
rect 29550 3712 29614 3716
rect 29550 3656 29554 3712
rect 29554 3656 29610 3712
rect 29610 3656 29614 3712
rect 29550 3652 29614 3656
rect 29756 3714 29820 3718
rect 29756 3658 29760 3714
rect 29760 3658 29816 3714
rect 29816 3658 29820 3714
rect 29756 3654 29820 3658
rect 29964 3721 30028 3725
rect 29964 3665 29968 3721
rect 29968 3665 30024 3721
rect 30024 3665 30028 3721
rect 29964 3661 30028 3665
rect 30186 3722 30250 3726
rect 30186 3666 30190 3722
rect 30190 3666 30246 3722
rect 30246 3666 30250 3722
rect 30186 3662 30250 3666
rect 23611 3264 23761 3410
rect 25737 3076 25801 3080
rect 25737 3020 25741 3076
rect 25741 3020 25797 3076
rect 25797 3020 25801 3076
rect 25737 3016 25801 3020
rect 25953 3081 26017 3085
rect 25953 3025 25957 3081
rect 25957 3025 26013 3081
rect 26013 3025 26017 3081
rect 25953 3021 26017 3025
rect 26159 3082 26223 3086
rect 26159 3026 26163 3082
rect 26163 3026 26219 3082
rect 26219 3026 26223 3082
rect 26159 3022 26223 3026
rect 26361 3074 26425 3078
rect 26361 3018 26365 3074
rect 26365 3018 26421 3074
rect 26421 3018 26425 3074
rect 26361 3014 26425 3018
rect 26557 3076 26621 3080
rect 26557 3020 26561 3076
rect 26561 3020 26617 3076
rect 26617 3020 26621 3076
rect 26557 3016 26621 3020
rect 26782 3078 26846 3082
rect 26782 3022 26786 3078
rect 26786 3022 26842 3078
rect 26842 3022 26846 3078
rect 26782 3018 26846 3022
rect 26997 3074 27061 3078
rect 26997 3018 27001 3074
rect 27001 3018 27057 3074
rect 27057 3018 27061 3074
rect 26997 3014 27061 3018
rect 27232 3074 27296 3078
rect 27232 3018 27236 3074
rect 27236 3018 27292 3074
rect 27292 3018 27296 3074
rect 27232 3014 27296 3018
rect 27440 3077 27504 3081
rect 27440 3021 27444 3077
rect 27444 3021 27500 3077
rect 27500 3021 27504 3077
rect 27440 3017 27504 3021
rect 27682 3077 27746 3081
rect 27682 3021 27686 3077
rect 27686 3021 27742 3077
rect 27742 3021 27746 3077
rect 27682 3017 27746 3021
rect 27880 3078 27944 3082
rect 27880 3022 27884 3078
rect 27884 3022 27940 3078
rect 27940 3022 27944 3078
rect 27880 3018 27944 3022
rect 28187 3078 28251 3082
rect 28187 3022 28191 3078
rect 28191 3022 28247 3078
rect 28247 3022 28251 3078
rect 28187 3018 28251 3022
rect 28412 3079 28476 3083
rect 28412 3023 28416 3079
rect 28416 3023 28472 3079
rect 28472 3023 28476 3079
rect 28412 3019 28476 3023
rect 28641 3078 28705 3082
rect 28641 3022 28645 3078
rect 28645 3022 28701 3078
rect 28701 3022 28705 3078
rect 28641 3018 28705 3022
rect 28857 3082 28921 3086
rect 28857 3026 28861 3082
rect 28861 3026 28917 3082
rect 28917 3026 28921 3082
rect 28857 3022 28921 3026
rect 29080 3085 29144 3089
rect 29080 3029 29084 3085
rect 29084 3029 29140 3085
rect 29140 3029 29144 3085
rect 29080 3025 29144 3029
rect 29304 3081 29368 3085
rect 29304 3025 29308 3081
rect 29308 3025 29364 3081
rect 29364 3025 29368 3081
rect 29304 3021 29368 3025
rect 29531 3070 29595 3074
rect 29531 3014 29535 3070
rect 29535 3014 29591 3070
rect 29591 3014 29595 3070
rect 29531 3010 29595 3014
rect 29744 3069 29808 3073
rect 29744 3013 29748 3069
rect 29748 3013 29804 3069
rect 29804 3013 29808 3069
rect 29744 3009 29808 3013
rect 29955 3073 30019 3077
rect 29955 3017 29959 3073
rect 29959 3017 30015 3073
rect 30015 3017 30019 3073
rect 29955 3013 30019 3017
rect 30182 3074 30246 3078
rect 30182 3018 30186 3074
rect 30186 3018 30242 3074
rect 30242 3018 30246 3074
rect 30182 3014 30246 3018
rect 27071 2847 27135 2851
rect 27071 2791 27075 2847
rect 27075 2791 27131 2847
rect 27131 2791 27135 2847
rect 27071 2787 27135 2791
rect 27454 2788 27518 2792
rect 27454 2732 27458 2788
rect 27458 2732 27514 2788
rect 27514 2732 27518 2788
rect 27454 2728 27518 2732
rect 29463 2849 29527 2853
rect 29463 2793 29467 2849
rect 29467 2793 29523 2849
rect 29523 2793 29527 2849
rect 29463 2789 29527 2793
rect 29840 2795 29904 2799
rect 29840 2739 29844 2795
rect 29844 2739 29900 2795
rect 29900 2739 29904 2795
rect 29840 2735 29904 2739
rect 25763 2431 25827 2435
rect 25763 2375 25767 2431
rect 25767 2375 25823 2431
rect 25823 2375 25827 2431
rect 25763 2371 25827 2375
rect 25988 2440 26052 2444
rect 25988 2384 25992 2440
rect 25992 2384 26048 2440
rect 26048 2384 26052 2440
rect 25988 2380 26052 2384
rect 26265 2437 26329 2441
rect 26265 2381 26269 2437
rect 26269 2381 26325 2437
rect 26325 2381 26329 2437
rect 26265 2377 26329 2381
rect 26486 2440 26550 2444
rect 26486 2384 26490 2440
rect 26490 2384 26546 2440
rect 26546 2384 26550 2440
rect 26486 2380 26550 2384
rect 26731 2437 26795 2441
rect 26731 2381 26735 2437
rect 26735 2381 26791 2437
rect 26791 2381 26795 2437
rect 26731 2377 26795 2381
rect 26957 2441 27021 2445
rect 26957 2385 26961 2441
rect 26961 2385 27017 2441
rect 27017 2385 27021 2441
rect 26957 2381 27021 2385
rect 27169 2439 27233 2443
rect 27169 2383 27173 2439
rect 27173 2383 27229 2439
rect 27229 2383 27233 2439
rect 27169 2379 27233 2383
rect 27389 2445 27453 2449
rect 27389 2389 27393 2445
rect 27393 2389 27449 2445
rect 27449 2389 27453 2445
rect 27389 2385 27453 2389
rect 27627 2447 27691 2451
rect 27627 2391 27631 2447
rect 27631 2391 27687 2447
rect 27687 2391 27691 2447
rect 27627 2387 27691 2391
rect 27840 2449 27904 2453
rect 27840 2393 27844 2449
rect 27844 2393 27900 2449
rect 27900 2393 27904 2449
rect 27840 2389 27904 2393
rect 28227 2439 28291 2443
rect 28227 2383 28231 2439
rect 28231 2383 28287 2439
rect 28287 2383 28291 2439
rect 28227 2379 28291 2383
rect 28574 2440 28638 2444
rect 28574 2384 28578 2440
rect 28578 2384 28634 2440
rect 28634 2384 28638 2440
rect 28574 2380 28638 2384
rect 28810 2435 28874 2439
rect 28810 2379 28814 2435
rect 28814 2379 28870 2435
rect 28870 2379 28874 2435
rect 28810 2375 28874 2379
rect 28994 2435 29058 2439
rect 28994 2379 28998 2435
rect 28998 2379 29054 2435
rect 29054 2379 29058 2435
rect 28994 2375 29058 2379
rect 29233 2437 29297 2441
rect 29233 2381 29237 2437
rect 29237 2381 29293 2437
rect 29293 2381 29297 2437
rect 29233 2377 29297 2381
rect 29436 2433 29500 2437
rect 29436 2377 29440 2433
rect 29440 2377 29496 2433
rect 29496 2377 29500 2433
rect 29436 2373 29500 2377
rect 29621 2430 29685 2434
rect 29621 2374 29625 2430
rect 29625 2374 29681 2430
rect 29681 2374 29685 2430
rect 29621 2370 29685 2374
rect 29812 2432 29876 2436
rect 29812 2376 29816 2432
rect 29816 2376 29872 2432
rect 29872 2376 29876 2432
rect 29812 2372 29876 2376
rect 30003 2436 30067 2440
rect 30003 2380 30007 2436
rect 30007 2380 30063 2436
rect 30063 2380 30067 2436
rect 30003 2376 30067 2380
rect 30189 2432 30253 2436
rect 30189 2376 30193 2432
rect 30193 2376 30249 2432
rect 30249 2376 30253 2432
rect 30189 2372 30253 2376
rect 25636 1849 25700 1853
rect 25636 1793 25640 1849
rect 25640 1793 25696 1849
rect 25696 1793 25700 1849
rect 25636 1789 25700 1793
rect 25841 1845 25905 1849
rect 25841 1789 25845 1845
rect 25845 1789 25901 1845
rect 25901 1789 25905 1845
rect 25841 1785 25905 1789
rect 26027 1850 26091 1854
rect 26027 1794 26031 1850
rect 26031 1794 26087 1850
rect 26087 1794 26091 1850
rect 26027 1790 26091 1794
rect 26221 1843 26285 1847
rect 26221 1787 26225 1843
rect 26225 1787 26281 1843
rect 26281 1787 26285 1843
rect 26221 1783 26285 1787
rect 26440 1848 26504 1852
rect 26440 1792 26444 1848
rect 26444 1792 26500 1848
rect 26500 1792 26504 1848
rect 26440 1788 26504 1792
rect 26650 1848 26714 1852
rect 26650 1792 26654 1848
rect 26654 1792 26710 1848
rect 26710 1792 26714 1848
rect 26650 1788 26714 1792
rect 26879 1845 26943 1849
rect 26879 1789 26883 1845
rect 26883 1789 26939 1845
rect 26939 1789 26943 1845
rect 26879 1785 26943 1789
rect 27125 1845 27189 1849
rect 27125 1789 27129 1845
rect 27129 1789 27185 1845
rect 27185 1789 27189 1845
rect 27125 1785 27189 1789
rect 27399 1845 27463 1849
rect 27399 1789 27403 1845
rect 27403 1789 27459 1845
rect 27459 1789 27463 1845
rect 27399 1785 27463 1789
rect 27674 1845 27738 1849
rect 27674 1789 27678 1845
rect 27678 1789 27734 1845
rect 27734 1789 27738 1845
rect 27674 1785 27738 1789
rect 27910 1845 27974 1849
rect 27910 1789 27914 1845
rect 27914 1789 27970 1845
rect 27970 1789 27974 1845
rect 27910 1785 27974 1789
rect 28133 1848 28197 1852
rect 28133 1792 28137 1848
rect 28137 1792 28193 1848
rect 28193 1792 28197 1848
rect 28133 1788 28197 1792
rect 28351 1851 28415 1855
rect 28351 1795 28355 1851
rect 28355 1795 28411 1851
rect 28411 1795 28415 1851
rect 28351 1791 28415 1795
rect 28529 1842 28593 1846
rect 28529 1786 28533 1842
rect 28533 1786 28589 1842
rect 28589 1786 28593 1842
rect 28529 1782 28593 1786
rect 28768 1844 28832 1848
rect 28768 1788 28772 1844
rect 28772 1788 28828 1844
rect 28828 1788 28832 1844
rect 28768 1784 28832 1788
rect 28965 1844 29029 1848
rect 28965 1788 28969 1844
rect 28969 1788 29025 1844
rect 29025 1788 29029 1844
rect 28965 1784 29029 1788
rect 29163 1844 29227 1848
rect 29163 1788 29167 1844
rect 29167 1788 29223 1844
rect 29223 1788 29227 1844
rect 29163 1784 29227 1788
rect 29376 1845 29440 1849
rect 29376 1789 29380 1845
rect 29380 1789 29436 1845
rect 29436 1789 29440 1845
rect 29376 1785 29440 1789
rect 29599 1844 29663 1848
rect 29599 1788 29603 1844
rect 29603 1788 29659 1844
rect 29659 1788 29663 1844
rect 29599 1784 29663 1788
rect 29796 1849 29860 1853
rect 29796 1793 29800 1849
rect 29800 1793 29856 1849
rect 29856 1793 29860 1849
rect 29796 1789 29860 1793
rect 30012 1847 30076 1851
rect 30012 1791 30016 1847
rect 30016 1791 30072 1847
rect 30072 1791 30076 1847
rect 30012 1787 30076 1791
rect 30221 1847 30285 1851
rect 30221 1791 30225 1847
rect 30225 1791 30281 1847
rect 30281 1791 30285 1847
rect 30221 1787 30285 1791
rect 8622 1413 8686 1417
rect 8622 1357 8626 1413
rect 8626 1357 8682 1413
rect 8682 1357 8686 1413
rect 8622 1353 8686 1357
rect 8824 1415 8888 1419
rect 8824 1359 8828 1415
rect 8828 1359 8884 1415
rect 8884 1359 8888 1415
rect 8824 1355 8888 1359
rect 9035 1413 9099 1417
rect 9035 1357 9039 1413
rect 9039 1357 9095 1413
rect 9095 1357 9099 1413
rect 9035 1353 9099 1357
rect 9225 1413 9289 1417
rect 9225 1357 9229 1413
rect 9229 1357 9285 1413
rect 9285 1357 9289 1413
rect 9225 1353 9289 1357
rect 9433 1415 9497 1419
rect 9433 1359 9437 1415
rect 9437 1359 9493 1415
rect 9493 1359 9497 1415
rect 9433 1355 9497 1359
rect 9635 1415 9699 1419
rect 9635 1359 9639 1415
rect 9639 1359 9695 1415
rect 9695 1359 9699 1415
rect 9635 1355 9699 1359
rect 9834 1417 9898 1421
rect 9834 1361 9838 1417
rect 9838 1361 9894 1417
rect 9894 1361 9898 1417
rect 9834 1357 9898 1361
rect 10029 1414 10093 1418
rect 10029 1358 10033 1414
rect 10033 1358 10089 1414
rect 10089 1358 10093 1414
rect 10029 1354 10093 1358
rect 10230 1416 10294 1420
rect 10230 1360 10234 1416
rect 10234 1360 10290 1416
rect 10290 1360 10294 1416
rect 10230 1356 10294 1360
rect 10447 1414 10511 1418
rect 10447 1358 10451 1414
rect 10451 1358 10507 1414
rect 10507 1358 10511 1414
rect 10447 1354 10511 1358
rect 10721 1417 10785 1421
rect 10721 1361 10725 1417
rect 10725 1361 10781 1417
rect 10781 1361 10785 1417
rect 10721 1357 10785 1361
rect 10998 1410 11062 1414
rect 10998 1354 11002 1410
rect 11002 1354 11058 1410
rect 11058 1354 11062 1410
rect 10998 1350 11062 1354
rect 11221 1413 11285 1417
rect 11221 1357 11225 1413
rect 11225 1357 11281 1413
rect 11281 1357 11285 1413
rect 11221 1353 11285 1357
rect 11453 1412 11517 1416
rect 11453 1356 11457 1412
rect 11457 1356 11513 1412
rect 11513 1356 11517 1412
rect 11453 1352 11517 1356
rect 13089 1409 13153 1413
rect 13089 1353 13093 1409
rect 13093 1353 13149 1409
rect 13149 1353 13153 1409
rect 13089 1349 13153 1353
rect 13397 1410 13461 1414
rect 13397 1354 13401 1410
rect 13401 1354 13457 1410
rect 13457 1354 13461 1410
rect 13397 1350 13461 1354
rect 13597 1411 13661 1415
rect 13597 1355 13601 1411
rect 13601 1355 13657 1411
rect 13657 1355 13661 1411
rect 13597 1351 13661 1355
rect 13816 1410 13880 1414
rect 13816 1354 13820 1410
rect 13820 1354 13876 1410
rect 13876 1354 13880 1410
rect 13816 1350 13880 1354
rect 14062 1409 14126 1413
rect 14062 1353 14066 1409
rect 14066 1353 14122 1409
rect 14122 1353 14126 1409
rect 14062 1349 14126 1353
rect 14270 1411 14334 1415
rect 14270 1355 14274 1411
rect 14274 1355 14330 1411
rect 14330 1355 14334 1411
rect 14270 1351 14334 1355
rect 14472 1412 14536 1416
rect 14472 1356 14476 1412
rect 14476 1356 14532 1412
rect 14532 1356 14536 1412
rect 14472 1352 14536 1356
rect 14665 1411 14729 1415
rect 14665 1355 14669 1411
rect 14669 1355 14725 1411
rect 14725 1355 14729 1411
rect 14665 1351 14729 1355
rect 15037 1410 15101 1414
rect 15037 1354 15041 1410
rect 15041 1354 15097 1410
rect 15097 1354 15101 1410
rect 15037 1350 15101 1354
rect 15226 1408 15290 1412
rect 15226 1352 15230 1408
rect 15230 1352 15286 1408
rect 15286 1352 15290 1408
rect 15226 1348 15290 1352
rect 15516 1408 15580 1412
rect 15516 1352 15520 1408
rect 15520 1352 15576 1408
rect 15576 1352 15580 1408
rect 15516 1348 15580 1352
rect 15789 1410 15853 1414
rect 15789 1354 15793 1410
rect 15793 1354 15849 1410
rect 15849 1354 15853 1410
rect 15789 1350 15853 1354
rect 9740 874 9804 878
rect 9740 818 9744 874
rect 9744 818 9800 874
rect 9800 818 9804 874
rect 9740 814 9804 818
rect 9959 878 10023 882
rect 9959 822 9963 878
rect 9963 822 10019 878
rect 10019 822 10023 878
rect 9959 818 10023 822
rect 10242 878 10306 882
rect 10242 822 10246 878
rect 10246 822 10302 878
rect 10302 822 10306 878
rect 10242 818 10306 822
rect 10451 878 10515 882
rect 10451 822 10455 878
rect 10455 822 10511 878
rect 10511 822 10515 878
rect 10451 818 10515 822
rect 10722 876 10786 880
rect 10722 820 10726 876
rect 10726 820 10782 876
rect 10782 820 10786 876
rect 10722 816 10786 820
rect 12797 874 12861 878
rect 12797 818 12801 874
rect 12801 818 12857 874
rect 12857 818 12861 874
rect 12797 814 12861 818
rect 13046 877 13110 881
rect 13046 821 13050 877
rect 13050 821 13106 877
rect 13106 821 13110 877
rect 13046 817 13110 821
rect 13390 863 13454 867
rect 13390 807 13394 863
rect 13394 807 13450 863
rect 13450 807 13454 863
rect 13390 803 13454 807
rect 13644 869 13708 873
rect 13644 813 13648 869
rect 13648 813 13704 869
rect 13704 813 13708 869
rect 13644 809 13708 813
rect 13873 869 13937 873
rect 13873 813 13877 869
rect 13877 813 13933 869
rect 13933 813 13937 869
rect 13873 809 13937 813
rect 15591 874 15655 878
rect 15591 818 15595 874
rect 15595 818 15651 874
rect 15651 818 15655 874
rect 15591 814 15655 818
rect 15795 876 15859 880
rect 15795 820 15799 876
rect 15799 820 15855 876
rect 15855 820 15859 876
rect 15795 816 15859 820
rect 16118 874 16182 878
rect 16118 818 16122 874
rect 16122 818 16178 874
rect 16178 818 16182 874
rect 16118 814 16182 818
rect 8588 269 8652 273
rect 8588 213 8592 269
rect 8592 213 8648 269
rect 8648 213 8652 269
rect 8588 209 8652 213
rect 8828 267 8892 271
rect 8828 211 8832 267
rect 8832 211 8888 267
rect 8888 211 8892 267
rect 8828 207 8892 211
rect 9150 266 9214 270
rect 9150 210 9154 266
rect 9154 210 9210 266
rect 9210 210 9214 266
rect 9150 206 9214 210
rect 9368 267 9432 271
rect 9368 211 9372 267
rect 9372 211 9428 267
rect 9428 211 9432 267
rect 9368 207 9432 211
rect 11272 271 11336 275
rect 11272 215 11276 271
rect 11276 215 11332 271
rect 11332 215 11336 271
rect 11272 211 11336 215
rect 11597 273 11661 277
rect 11597 217 11601 273
rect 11601 217 11657 273
rect 11657 217 11661 273
rect 11597 213 11661 217
rect 11865 273 11929 277
rect 11865 217 11869 273
rect 11869 217 11925 273
rect 11925 217 11929 273
rect 11865 213 11929 217
rect 12131 273 12195 277
rect 12131 217 12135 273
rect 12135 217 12191 273
rect 12191 217 12195 273
rect 12131 213 12195 217
rect 12371 271 12435 275
rect 12371 215 12375 271
rect 12375 215 12431 271
rect 12431 215 12435 271
rect 12371 211 12435 215
rect 14165 274 14229 278
rect 14165 218 14169 274
rect 14169 218 14225 274
rect 14225 218 14229 274
rect 14165 214 14229 218
rect 14531 277 14595 281
rect 14531 221 14535 277
rect 14535 221 14591 277
rect 14591 221 14595 277
rect 14531 217 14595 221
rect 14775 277 14839 281
rect 14775 221 14779 277
rect 14779 221 14835 277
rect 14835 221 14839 277
rect 14775 217 14839 221
rect 15198 268 15262 272
rect 15198 212 15202 268
rect 15202 212 15258 268
rect 15258 212 15262 268
rect 15198 208 15262 212
rect 17141 270 17205 274
rect 17141 214 17145 270
rect 17145 214 17201 270
rect 17201 214 17205 270
rect 17141 210 17205 214
rect 17393 267 17457 271
rect 17393 211 17397 267
rect 17397 211 17453 267
rect 17453 211 17457 267
rect 17393 207 17457 211
rect 17599 275 17663 279
rect 17599 219 17603 275
rect 17603 219 17659 275
rect 17659 219 17663 275
rect 17599 215 17663 219
rect 17882 269 17946 273
rect 17882 213 17886 269
rect 17886 213 17942 269
rect 17942 213 17946 269
rect 17882 209 17946 213
rect 18180 270 18244 274
rect 18180 214 18184 270
rect 18184 214 18240 270
rect 18240 214 18244 270
rect 18180 210 18244 214
rect 20012 271 20076 275
rect 20012 215 20016 271
rect 20016 215 20072 271
rect 20072 215 20076 271
rect 20012 211 20076 215
rect 20222 273 20286 277
rect 20222 217 20226 273
rect 20226 217 20282 273
rect 20282 217 20286 273
rect 20222 213 20286 217
rect 20573 271 20637 275
rect 20573 215 20577 271
rect 20577 215 20633 271
rect 20633 215 20637 271
rect 20573 211 20637 215
rect 20853 271 20917 275
rect 20853 215 20857 271
rect 20857 215 20913 271
rect 20913 215 20917 271
rect 20853 211 20917 215
rect 21170 270 21234 274
rect 21170 214 21174 270
rect 21174 214 21230 270
rect 21230 214 21234 270
rect 21170 210 21234 214
rect 22960 268 23024 272
rect 22960 212 22964 268
rect 22964 212 23020 268
rect 23020 212 23024 268
rect 22960 208 23024 212
rect 23255 268 23319 272
rect 23255 212 23259 268
rect 23259 212 23315 268
rect 23315 212 23319 268
rect 23255 208 23319 212
rect 23542 268 23606 272
rect 23542 212 23546 268
rect 23546 212 23602 268
rect 23602 212 23606 268
rect 23542 208 23606 212
rect 23832 268 23896 272
rect 23832 212 23836 268
rect 23836 212 23892 268
rect 23892 212 23896 268
rect 23832 208 23896 212
rect 24116 271 24180 275
rect 24116 215 24120 271
rect 24120 215 24176 271
rect 24176 215 24180 271
rect 24116 211 24180 215
rect 9779 -269 9843 -265
rect 9779 -325 9783 -269
rect 9783 -325 9839 -269
rect 9839 -325 9843 -269
rect 9779 -329 9843 -325
rect 9996 -269 10060 -265
rect 9996 -325 10000 -269
rect 10000 -325 10056 -269
rect 10056 -325 10060 -269
rect 9996 -329 10060 -325
rect 10215 -269 10279 -265
rect 10215 -325 10219 -269
rect 10219 -325 10275 -269
rect 10275 -325 10279 -269
rect 10215 -329 10279 -325
rect 10428 -273 10492 -269
rect 10428 -329 10432 -273
rect 10432 -329 10488 -273
rect 10488 -329 10492 -273
rect 10428 -333 10492 -329
rect 10639 -273 10703 -269
rect 10639 -329 10643 -273
rect 10643 -329 10699 -273
rect 10699 -329 10703 -273
rect 10639 -333 10703 -329
rect 12763 -273 12827 -269
rect 12763 -329 12767 -273
rect 12767 -329 12823 -273
rect 12823 -329 12827 -273
rect 12763 -333 12827 -329
rect 13041 -274 13105 -270
rect 13041 -330 13045 -274
rect 13045 -330 13101 -274
rect 13101 -330 13105 -274
rect 13041 -334 13105 -330
rect 13613 -269 13677 -265
rect 13613 -325 13617 -269
rect 13617 -325 13673 -269
rect 13673 -325 13677 -269
rect 13613 -329 13677 -325
rect 13852 -269 13916 -265
rect 13852 -325 13856 -269
rect 13856 -325 13912 -269
rect 13912 -325 13916 -269
rect 13852 -329 13916 -325
rect 16010 -271 16074 -267
rect 16010 -327 16014 -271
rect 16014 -327 16070 -271
rect 16070 -327 16074 -271
rect 16010 -331 16074 -327
rect 16237 -266 16301 -262
rect 16237 -322 16241 -266
rect 16241 -322 16297 -266
rect 16297 -322 16301 -266
rect 16237 -326 16301 -322
rect 16427 -264 16491 -260
rect 16427 -320 16431 -264
rect 16431 -320 16487 -264
rect 16487 -320 16491 -264
rect 16427 -324 16491 -320
rect 16643 -273 16707 -269
rect 16643 -329 16647 -273
rect 16647 -329 16703 -273
rect 16703 -329 16707 -273
rect 16643 -333 16707 -329
rect 18624 -270 18688 -266
rect 18624 -326 18628 -270
rect 18628 -326 18684 -270
rect 18684 -326 18688 -270
rect 18624 -330 18688 -326
rect 18853 -267 18917 -263
rect 18853 -323 18857 -267
rect 18857 -323 18913 -267
rect 18913 -323 18917 -267
rect 18853 -327 18917 -323
rect 19079 -262 19143 -258
rect 19079 -318 19083 -262
rect 19083 -318 19139 -262
rect 19139 -318 19143 -262
rect 19079 -322 19143 -318
rect 19307 -270 19371 -266
rect 19307 -326 19311 -270
rect 19311 -326 19367 -270
rect 19367 -326 19371 -270
rect 19307 -330 19371 -326
rect 19543 -264 19607 -260
rect 19543 -320 19547 -264
rect 19547 -320 19603 -264
rect 19603 -320 19607 -264
rect 19543 -324 19607 -320
rect 19735 -273 19799 -269
rect 19735 -329 19739 -273
rect 19739 -329 19795 -273
rect 19795 -329 19799 -273
rect 19735 -333 19799 -329
rect 21470 -273 21534 -269
rect 21470 -329 21474 -273
rect 21474 -329 21530 -273
rect 21530 -329 21534 -273
rect 21470 -333 21534 -329
rect 21674 -268 21738 -264
rect 21674 -324 21678 -268
rect 21678 -324 21734 -268
rect 21734 -324 21738 -268
rect 21674 -328 21738 -324
rect 21865 -273 21929 -269
rect 21865 -329 21869 -273
rect 21869 -329 21925 -273
rect 21925 -329 21929 -273
rect 21865 -333 21929 -329
rect 22067 -274 22131 -270
rect 22067 -330 22071 -274
rect 22071 -330 22127 -274
rect 22127 -330 22131 -274
rect 22067 -334 22131 -330
rect 22357 -273 22421 -269
rect 22357 -329 22361 -273
rect 22361 -329 22417 -273
rect 22417 -329 22421 -273
rect 22357 -333 22421 -329
rect 22642 -274 22706 -270
rect 22642 -330 22646 -274
rect 22646 -330 22702 -274
rect 22702 -330 22706 -274
rect 22642 -334 22706 -330
rect 24397 -269 24461 -265
rect 24397 -325 24401 -269
rect 24401 -325 24457 -269
rect 24457 -325 24461 -269
rect 24397 -329 24461 -325
rect 24591 -265 24655 -261
rect 24591 -321 24595 -265
rect 24595 -321 24651 -265
rect 24651 -321 24655 -265
rect 24591 -325 24655 -321
rect 24780 -268 24844 -264
rect 24780 -324 24784 -268
rect 24784 -324 24840 -268
rect 24840 -324 24844 -268
rect 24780 -328 24844 -324
rect 25003 -266 25067 -262
rect 25003 -322 25007 -266
rect 25007 -322 25063 -266
rect 25063 -322 25067 -266
rect 25003 -326 25067 -322
rect 8834 -414 8898 -410
rect 8834 -470 8838 -414
rect 8838 -470 8894 -414
rect 8894 -470 8898 -414
rect 8834 -474 8898 -470
rect 9036 -418 9100 -414
rect 9036 -474 9040 -418
rect 9040 -474 9096 -418
rect 9096 -474 9100 -418
rect 9036 -478 9100 -474
rect 9225 -421 9289 -417
rect 9225 -477 9229 -421
rect 9229 -477 9285 -421
rect 9285 -477 9289 -421
rect 9225 -481 9289 -477
rect 9454 -420 9518 -416
rect 9454 -476 9458 -420
rect 9458 -476 9514 -420
rect 9514 -476 9518 -420
rect 9454 -480 9518 -476
rect 11223 -417 11287 -413
rect 11223 -473 11227 -417
rect 11227 -473 11283 -417
rect 11283 -473 11287 -417
rect 11223 -477 11287 -473
rect 11438 -420 11502 -416
rect 11438 -476 11442 -420
rect 11442 -476 11498 -420
rect 11498 -476 11502 -420
rect 11438 -480 11502 -476
rect 11636 -423 11700 -419
rect 11636 -479 11640 -423
rect 11640 -479 11696 -423
rect 11696 -479 11700 -423
rect 11636 -483 11700 -479
rect 11831 -413 11895 -409
rect 11831 -469 11835 -413
rect 11835 -469 11891 -413
rect 11891 -469 11895 -413
rect 11831 -473 11895 -469
rect 12111 -415 12175 -411
rect 12111 -471 12115 -415
rect 12115 -471 12171 -415
rect 12171 -471 12175 -415
rect 12111 -475 12175 -471
rect 12330 -417 12394 -413
rect 12330 -473 12334 -417
rect 12334 -473 12390 -417
rect 12390 -473 12394 -417
rect 12330 -477 12394 -473
rect 14151 -420 14215 -416
rect 14151 -476 14155 -420
rect 14155 -476 14211 -420
rect 14211 -476 14215 -420
rect 14151 -480 14215 -476
rect 14502 -423 14566 -419
rect 14502 -479 14506 -423
rect 14506 -479 14562 -423
rect 14562 -479 14566 -423
rect 14502 -483 14566 -479
rect 14691 -425 14755 -421
rect 14691 -481 14695 -425
rect 14695 -481 14751 -425
rect 14751 -481 14755 -425
rect 14691 -485 14755 -481
rect 14896 -418 14960 -414
rect 14896 -474 14900 -418
rect 14900 -474 14956 -418
rect 14956 -474 14960 -418
rect 14896 -478 14960 -474
rect 15087 -416 15151 -412
rect 15087 -472 15091 -416
rect 15091 -472 15147 -416
rect 15147 -472 15151 -416
rect 15087 -476 15151 -472
rect 17132 -414 17196 -410
rect 17132 -470 17136 -414
rect 17136 -470 17192 -414
rect 17192 -470 17196 -414
rect 17132 -474 17196 -470
rect 17322 -412 17386 -408
rect 17322 -468 17326 -412
rect 17326 -468 17382 -412
rect 17382 -468 17386 -412
rect 17322 -472 17386 -468
rect 17516 -414 17580 -410
rect 17516 -470 17520 -414
rect 17520 -470 17576 -414
rect 17576 -470 17580 -414
rect 17516 -474 17580 -470
rect 17827 -418 17891 -414
rect 17827 -474 17831 -418
rect 17831 -474 17887 -418
rect 17887 -474 17891 -418
rect 17827 -478 17891 -474
rect 20010 -419 20074 -415
rect 20010 -475 20014 -419
rect 20014 -475 20070 -419
rect 20070 -475 20074 -419
rect 20010 -479 20074 -475
rect 20214 -419 20278 -415
rect 20214 -475 20218 -419
rect 20218 -475 20274 -419
rect 20274 -475 20278 -419
rect 20214 -479 20278 -475
rect 20779 -423 20843 -419
rect 20779 -479 20783 -423
rect 20783 -479 20839 -423
rect 20839 -479 20843 -423
rect 20779 -483 20843 -479
rect 21018 -421 21082 -417
rect 21018 -477 21022 -421
rect 21022 -477 21078 -421
rect 21078 -477 21082 -421
rect 21018 -481 21082 -477
rect 21222 -421 21286 -417
rect 21222 -477 21226 -421
rect 21226 -477 21282 -421
rect 21282 -477 21286 -421
rect 21222 -481 21286 -477
rect 23182 -413 23246 -409
rect 23182 -469 23186 -413
rect 23186 -469 23242 -413
rect 23242 -469 23246 -413
rect 23182 -473 23246 -469
rect 23415 -415 23479 -411
rect 23415 -471 23419 -415
rect 23419 -471 23475 -415
rect 23475 -471 23479 -415
rect 23415 -475 23479 -471
rect 23622 -417 23686 -413
rect 23622 -473 23626 -417
rect 23626 -473 23682 -417
rect 23682 -473 23686 -417
rect 23622 -477 23686 -473
rect 23831 -415 23895 -411
rect 23831 -471 23835 -415
rect 23835 -471 23891 -415
rect 23891 -471 23895 -415
rect 23831 -475 23895 -471
rect 24111 -413 24175 -409
rect 24111 -469 24115 -413
rect 24115 -469 24171 -413
rect 24171 -469 24175 -413
rect 24111 -473 24175 -469
rect 9761 -963 9825 -959
rect 9761 -1019 9765 -963
rect 9765 -1019 9821 -963
rect 9821 -1019 9825 -963
rect 9761 -1023 9825 -1019
rect 9990 -951 10054 -947
rect 9990 -1007 9994 -951
rect 9994 -1007 10050 -951
rect 10050 -1007 10054 -951
rect 9990 -1011 10054 -1007
rect 10209 -961 10273 -957
rect 10209 -1017 10213 -961
rect 10213 -1017 10269 -961
rect 10269 -1017 10273 -961
rect 10209 -1021 10273 -1017
rect 10401 -957 10465 -953
rect 10401 -1013 10405 -957
rect 10405 -1013 10461 -957
rect 10461 -1013 10465 -957
rect 10401 -1017 10465 -1013
rect 10895 -959 10959 -955
rect 10895 -1015 10899 -959
rect 10899 -1015 10955 -959
rect 10955 -1015 10959 -959
rect 10895 -1019 10959 -1015
rect 12687 -960 12751 -956
rect 12687 -1016 12691 -960
rect 12691 -1016 12747 -960
rect 12747 -1016 12751 -960
rect 12687 -1020 12751 -1016
rect 13080 -962 13144 -958
rect 13080 -1018 13084 -962
rect 13084 -1018 13140 -962
rect 13140 -1018 13144 -962
rect 13080 -1022 13144 -1018
rect 13277 -954 13341 -950
rect 13277 -1010 13281 -954
rect 13281 -1010 13337 -954
rect 13337 -1010 13341 -954
rect 13277 -1014 13341 -1010
rect 13607 -952 13671 -948
rect 13607 -1008 13611 -952
rect 13611 -1008 13667 -952
rect 13667 -1008 13671 -952
rect 13607 -1012 13671 -1008
rect 13803 -952 13867 -948
rect 13803 -1008 13807 -952
rect 13807 -1008 13863 -952
rect 13863 -1008 13867 -952
rect 13803 -1012 13867 -1008
rect 15710 -959 15774 -955
rect 15710 -1015 15714 -959
rect 15714 -1015 15770 -959
rect 15770 -1015 15774 -959
rect 15710 -1019 15774 -1015
rect 16011 -955 16075 -951
rect 16011 -1011 16015 -955
rect 16015 -1011 16071 -955
rect 16071 -1011 16075 -955
rect 16011 -1015 16075 -1011
rect 16217 -954 16281 -950
rect 16217 -1010 16221 -954
rect 16221 -1010 16277 -954
rect 16277 -1010 16281 -954
rect 16217 -1014 16281 -1010
rect 16427 -958 16491 -954
rect 16427 -1014 16431 -958
rect 16431 -1014 16487 -958
rect 16487 -1014 16491 -958
rect 16427 -1018 16491 -1014
rect 16638 -952 16702 -948
rect 16638 -1008 16642 -952
rect 16642 -1008 16698 -952
rect 16698 -1008 16702 -952
rect 16638 -1012 16702 -1008
rect 18518 -963 18582 -959
rect 18518 -1019 18522 -963
rect 18522 -1019 18578 -963
rect 18578 -1019 18582 -963
rect 18518 -1023 18582 -1019
rect 18775 -956 18839 -952
rect 18775 -1012 18779 -956
rect 18779 -1012 18835 -956
rect 18835 -1012 18839 -956
rect 18775 -1016 18839 -1012
rect 19025 -960 19089 -956
rect 19025 -1016 19029 -960
rect 19029 -1016 19085 -960
rect 19085 -1016 19089 -960
rect 19025 -1020 19089 -1016
rect 19296 -955 19360 -951
rect 19296 -1011 19300 -955
rect 19300 -1011 19356 -955
rect 19356 -1011 19360 -955
rect 19296 -1015 19360 -1011
rect 19537 -952 19601 -948
rect 19537 -1008 19541 -952
rect 19541 -1008 19597 -952
rect 19597 -1008 19601 -952
rect 19537 -1012 19601 -1008
rect 19762 -956 19826 -952
rect 19762 -1012 19766 -956
rect 19766 -1012 19822 -956
rect 19822 -1012 19826 -956
rect 19762 -1016 19826 -1012
rect 21469 -958 21533 -954
rect 21469 -1014 21473 -958
rect 21473 -1014 21529 -958
rect 21529 -1014 21533 -958
rect 21469 -1018 21533 -1014
rect 21670 -957 21734 -953
rect 21670 -1013 21674 -957
rect 21674 -1013 21730 -957
rect 21730 -1013 21734 -957
rect 21670 -1017 21734 -1013
rect 21888 -961 21952 -957
rect 21888 -1017 21892 -961
rect 21892 -1017 21948 -961
rect 21948 -1017 21952 -961
rect 21888 -1021 21952 -1017
rect 22095 -957 22159 -953
rect 22095 -1013 22099 -957
rect 22099 -1013 22155 -957
rect 22155 -1013 22159 -957
rect 22095 -1017 22159 -1013
rect 22300 -958 22364 -954
rect 22300 -1014 22304 -958
rect 22304 -1014 22360 -958
rect 22360 -1014 22364 -958
rect 22300 -1018 22364 -1014
rect 22647 -962 22711 -958
rect 22647 -1018 22651 -962
rect 22651 -1018 22707 -962
rect 22707 -1018 22711 -962
rect 22647 -1022 22711 -1018
rect 24399 -958 24463 -954
rect 24399 -1014 24403 -958
rect 24403 -1014 24459 -958
rect 24459 -1014 24463 -958
rect 24399 -1018 24463 -1014
rect 24590 -955 24654 -951
rect 24590 -1011 24594 -955
rect 24594 -1011 24650 -955
rect 24650 -1011 24654 -955
rect 24590 -1015 24654 -1011
rect 24785 -953 24849 -949
rect 24785 -1009 24789 -953
rect 24789 -1009 24845 -953
rect 24845 -1009 24849 -953
rect 24785 -1013 24849 -1009
rect 25232 -958 25296 -954
rect 25232 -1014 25236 -958
rect 25236 -1014 25292 -958
rect 25292 -1014 25296 -958
rect 25232 -1018 25296 -1014
rect 8616 -1107 8680 -1103
rect 8616 -1163 8620 -1107
rect 8620 -1163 8676 -1107
rect 8676 -1163 8680 -1107
rect 8616 -1167 8680 -1163
rect 8849 -1111 8913 -1107
rect 8849 -1167 8853 -1111
rect 8853 -1167 8909 -1111
rect 8909 -1167 8913 -1111
rect 8849 -1171 8913 -1167
rect 9064 -1104 9128 -1100
rect 9064 -1160 9068 -1104
rect 9068 -1160 9124 -1104
rect 9124 -1160 9128 -1104
rect 9064 -1164 9128 -1160
rect 9282 -1107 9346 -1103
rect 9282 -1163 9286 -1107
rect 9286 -1163 9342 -1107
rect 9342 -1163 9346 -1107
rect 9282 -1167 9346 -1163
rect 9498 -1106 9562 -1102
rect 9498 -1162 9502 -1106
rect 9502 -1162 9558 -1106
rect 9558 -1162 9562 -1106
rect 9498 -1166 9562 -1162
rect 11219 -1110 11283 -1106
rect 11219 -1166 11223 -1110
rect 11223 -1166 11279 -1110
rect 11279 -1166 11283 -1110
rect 11219 -1170 11283 -1166
rect 11409 -1110 11473 -1106
rect 11409 -1166 11413 -1110
rect 11413 -1166 11469 -1110
rect 11469 -1166 11473 -1110
rect 11409 -1170 11473 -1166
rect 11619 -1107 11683 -1103
rect 11619 -1163 11623 -1107
rect 11623 -1163 11679 -1107
rect 11679 -1163 11683 -1107
rect 11619 -1167 11683 -1163
rect 11836 -1110 11900 -1106
rect 11836 -1166 11840 -1110
rect 11840 -1166 11896 -1110
rect 11896 -1166 11900 -1110
rect 11836 -1170 11900 -1166
rect 12131 -1107 12195 -1103
rect 12131 -1163 12135 -1107
rect 12135 -1163 12191 -1107
rect 12191 -1163 12195 -1107
rect 12131 -1167 12195 -1163
rect 12355 -1102 12419 -1098
rect 12355 -1158 12359 -1102
rect 12359 -1158 12415 -1102
rect 12415 -1158 12419 -1102
rect 12355 -1162 12419 -1158
rect 14233 -1109 14297 -1105
rect 14233 -1165 14237 -1109
rect 14237 -1165 14293 -1109
rect 14293 -1165 14297 -1109
rect 14233 -1169 14297 -1165
rect 14533 -1111 14597 -1107
rect 14533 -1167 14537 -1111
rect 14537 -1167 14593 -1111
rect 14593 -1167 14597 -1111
rect 14533 -1171 14597 -1167
rect 14785 -1107 14849 -1103
rect 14785 -1163 14789 -1107
rect 14789 -1163 14845 -1107
rect 14845 -1163 14849 -1107
rect 14785 -1167 14849 -1163
rect 15002 -1102 15066 -1098
rect 15002 -1158 15006 -1102
rect 15006 -1158 15062 -1102
rect 15062 -1158 15066 -1102
rect 15002 -1162 15066 -1158
rect 15203 -1105 15267 -1101
rect 15203 -1161 15207 -1105
rect 15207 -1161 15263 -1105
rect 15263 -1161 15267 -1105
rect 15203 -1165 15267 -1161
rect 17088 -1114 17152 -1110
rect 17088 -1170 17092 -1114
rect 17092 -1170 17148 -1114
rect 17148 -1170 17152 -1114
rect 17088 -1174 17152 -1170
rect 17280 -1114 17344 -1110
rect 17280 -1170 17284 -1114
rect 17284 -1170 17340 -1114
rect 17340 -1170 17344 -1114
rect 17280 -1174 17344 -1170
rect 17480 -1114 17544 -1110
rect 17480 -1170 17484 -1114
rect 17484 -1170 17540 -1114
rect 17540 -1170 17544 -1114
rect 17480 -1174 17544 -1170
rect 18098 -1106 18162 -1102
rect 18098 -1162 18102 -1106
rect 18102 -1162 18158 -1106
rect 18158 -1162 18162 -1106
rect 18098 -1166 18162 -1162
rect 19999 -1110 20063 -1106
rect 19999 -1166 20003 -1110
rect 20003 -1166 20059 -1110
rect 20059 -1166 20063 -1110
rect 19999 -1170 20063 -1166
rect 20255 -1110 20319 -1106
rect 20255 -1166 20259 -1110
rect 20259 -1166 20315 -1110
rect 20315 -1166 20319 -1110
rect 20255 -1170 20319 -1166
rect 20490 -1110 20554 -1106
rect 20490 -1166 20494 -1110
rect 20494 -1166 20550 -1110
rect 20550 -1166 20554 -1110
rect 20490 -1170 20554 -1166
rect 20779 -1108 20843 -1104
rect 20779 -1164 20783 -1108
rect 20783 -1164 20839 -1108
rect 20839 -1164 20843 -1108
rect 20779 -1168 20843 -1164
rect 20969 -1110 21033 -1106
rect 20969 -1166 20973 -1110
rect 20973 -1166 21029 -1110
rect 21029 -1166 21033 -1110
rect 20969 -1170 21033 -1166
rect 21173 -1108 21237 -1104
rect 21173 -1164 21177 -1108
rect 21177 -1164 21233 -1108
rect 21233 -1164 21237 -1108
rect 21173 -1168 21237 -1164
rect 22959 -1102 23023 -1098
rect 22959 -1158 22963 -1102
rect 22963 -1158 23019 -1102
rect 23019 -1158 23023 -1102
rect 22959 -1162 23023 -1158
rect 23201 -1106 23265 -1102
rect 23201 -1162 23205 -1106
rect 23205 -1162 23261 -1106
rect 23261 -1162 23265 -1106
rect 23201 -1166 23265 -1162
rect 23401 -1107 23465 -1103
rect 23401 -1163 23405 -1107
rect 23405 -1163 23461 -1107
rect 23461 -1163 23465 -1107
rect 23401 -1167 23465 -1163
rect 23591 -1099 23655 -1095
rect 23591 -1155 23595 -1099
rect 23595 -1155 23651 -1099
rect 23651 -1155 23655 -1099
rect 23591 -1159 23655 -1155
rect 23812 -1101 23876 -1097
rect 23812 -1157 23816 -1101
rect 23816 -1157 23872 -1101
rect 23872 -1157 23876 -1101
rect 23812 -1161 23876 -1157
rect 24108 -1106 24172 -1102
rect 24108 -1162 24112 -1106
rect 24112 -1162 24168 -1106
rect 24168 -1162 24172 -1106
rect 24108 -1166 24172 -1162
rect 8990 -1639 9054 -1635
rect 8990 -1695 8994 -1639
rect 8994 -1695 9050 -1639
rect 9050 -1695 9054 -1639
rect 8990 -1699 9054 -1695
rect 9189 -1642 9253 -1638
rect 9189 -1698 9193 -1642
rect 9193 -1698 9249 -1642
rect 9249 -1698 9253 -1642
rect 9189 -1702 9253 -1698
rect 9400 -1642 9464 -1638
rect 9400 -1698 9404 -1642
rect 9404 -1698 9460 -1642
rect 9460 -1698 9464 -1642
rect 9400 -1702 9464 -1698
rect 9606 -1642 9670 -1638
rect 9606 -1698 9610 -1642
rect 9610 -1698 9666 -1642
rect 9666 -1698 9670 -1642
rect 9606 -1702 9670 -1698
rect 9834 -1644 9898 -1640
rect 9834 -1700 9838 -1644
rect 9838 -1700 9894 -1644
rect 9894 -1700 9898 -1644
rect 9834 -1704 9898 -1700
rect 10078 -1644 10142 -1640
rect 10078 -1700 10082 -1644
rect 10082 -1700 10138 -1644
rect 10138 -1700 10142 -1644
rect 10078 -1704 10142 -1700
rect 10308 -1642 10372 -1638
rect 10308 -1698 10312 -1642
rect 10312 -1698 10368 -1642
rect 10368 -1698 10372 -1642
rect 10308 -1702 10372 -1698
rect 10514 -1642 10578 -1638
rect 10514 -1698 10518 -1642
rect 10518 -1698 10574 -1642
rect 10574 -1698 10578 -1642
rect 10514 -1702 10578 -1698
rect 10732 -1637 10796 -1633
rect 10732 -1693 10736 -1637
rect 10736 -1693 10792 -1637
rect 10792 -1693 10796 -1637
rect 10732 -1697 10796 -1693
rect 10935 -1643 10999 -1639
rect 10935 -1699 10939 -1643
rect 10939 -1699 10995 -1643
rect 10995 -1699 10999 -1643
rect 10935 -1703 10999 -1699
rect 11143 -1640 11207 -1636
rect 11143 -1696 11147 -1640
rect 11147 -1696 11203 -1640
rect 11203 -1696 11207 -1640
rect 11143 -1700 11207 -1696
rect 11406 -1644 11470 -1640
rect 11406 -1700 11410 -1644
rect 11410 -1700 11466 -1644
rect 11466 -1700 11470 -1644
rect 11406 -1704 11470 -1700
rect 11614 -1643 11678 -1639
rect 11614 -1699 11618 -1643
rect 11618 -1699 11674 -1643
rect 11674 -1699 11678 -1643
rect 11614 -1703 11678 -1699
rect 11824 -1646 11888 -1642
rect 11824 -1702 11828 -1646
rect 11828 -1702 11884 -1646
rect 11884 -1702 11888 -1646
rect 11824 -1706 11888 -1702
rect 12024 -1640 12088 -1636
rect 12024 -1696 12028 -1640
rect 12028 -1696 12084 -1640
rect 12084 -1696 12088 -1640
rect 12024 -1700 12088 -1696
rect 12227 -1643 12291 -1639
rect 12227 -1699 12231 -1643
rect 12231 -1699 12287 -1643
rect 12287 -1699 12291 -1643
rect 12227 -1703 12291 -1699
rect 12437 -1643 12501 -1639
rect 12437 -1699 12441 -1643
rect 12441 -1699 12497 -1643
rect 12497 -1699 12501 -1643
rect 12437 -1703 12501 -1699
rect 12638 -1642 12702 -1638
rect 12638 -1698 12642 -1642
rect 12642 -1698 12698 -1642
rect 12698 -1698 12702 -1642
rect 12638 -1702 12702 -1698
rect 12854 -1641 12918 -1637
rect 12854 -1697 12858 -1641
rect 12858 -1697 12914 -1641
rect 12914 -1697 12918 -1641
rect 12854 -1701 12918 -1697
rect 13135 -1643 13199 -1639
rect 13135 -1699 13139 -1643
rect 13139 -1699 13195 -1643
rect 13195 -1699 13199 -1643
rect 13135 -1703 13199 -1699
rect 13355 -1648 13419 -1644
rect 13355 -1704 13359 -1648
rect 13359 -1704 13415 -1648
rect 13415 -1704 13419 -1648
rect 13355 -1708 13419 -1704
rect 13560 -1647 13624 -1643
rect 13560 -1703 13564 -1647
rect 13564 -1703 13620 -1647
rect 13620 -1703 13624 -1647
rect 13560 -1707 13624 -1703
rect 13781 -1641 13845 -1637
rect 13781 -1697 13785 -1641
rect 13785 -1697 13841 -1641
rect 13841 -1697 13845 -1641
rect 13781 -1701 13845 -1697
rect 13986 -1648 14050 -1644
rect 13986 -1704 13990 -1648
rect 13990 -1704 14046 -1648
rect 14046 -1704 14050 -1648
rect 13986 -1708 14050 -1704
rect 14195 -1647 14259 -1643
rect 14195 -1703 14199 -1647
rect 14199 -1703 14255 -1647
rect 14255 -1703 14259 -1647
rect 14195 -1707 14259 -1703
rect 14412 -1647 14476 -1643
rect 14412 -1703 14416 -1647
rect 14416 -1703 14472 -1647
rect 14472 -1703 14476 -1647
rect 14412 -1707 14476 -1703
rect 14626 -1642 14690 -1638
rect 14626 -1698 14630 -1642
rect 14630 -1698 14686 -1642
rect 14686 -1698 14690 -1642
rect 14626 -1702 14690 -1698
rect 14821 -1644 14885 -1640
rect 14821 -1700 14825 -1644
rect 14825 -1700 14881 -1644
rect 14881 -1700 14885 -1644
rect 14821 -1704 14885 -1700
rect 15016 -1647 15080 -1643
rect 15016 -1703 15020 -1647
rect 15020 -1703 15076 -1647
rect 15076 -1703 15080 -1647
rect 15016 -1707 15080 -1703
rect 15218 -1644 15282 -1640
rect 15218 -1700 15222 -1644
rect 15222 -1700 15278 -1644
rect 15278 -1700 15282 -1644
rect 15218 -1704 15282 -1700
rect 15502 -1643 15566 -1639
rect 15502 -1699 15506 -1643
rect 15506 -1699 15562 -1643
rect 15562 -1699 15566 -1643
rect 15502 -1703 15566 -1699
rect 15701 -1642 15765 -1638
rect 15701 -1698 15705 -1642
rect 15705 -1698 15761 -1642
rect 15761 -1698 15765 -1642
rect 15701 -1702 15765 -1698
rect 15904 -1640 15968 -1636
rect 15904 -1696 15908 -1640
rect 15908 -1696 15964 -1640
rect 15964 -1696 15968 -1640
rect 15904 -1700 15968 -1696
rect 16169 -1643 16233 -1639
rect 16169 -1699 16173 -1643
rect 16173 -1699 16229 -1643
rect 16229 -1699 16233 -1643
rect 16169 -1703 16233 -1699
rect 16367 -1644 16431 -1640
rect 16367 -1700 16371 -1644
rect 16371 -1700 16427 -1644
rect 16427 -1700 16431 -1644
rect 16367 -1704 16431 -1700
rect 16556 -1642 16620 -1638
rect 16556 -1698 16560 -1642
rect 16560 -1698 16616 -1642
rect 16616 -1698 16620 -1642
rect 16556 -1702 16620 -1698
rect 16768 -1642 16832 -1638
rect 16768 -1698 16772 -1642
rect 16772 -1698 16828 -1642
rect 16828 -1698 16832 -1642
rect 16768 -1702 16832 -1698
rect 16985 -1642 17049 -1638
rect 16985 -1698 16989 -1642
rect 16989 -1698 17045 -1642
rect 17045 -1698 17049 -1642
rect 16985 -1702 17049 -1698
rect 17190 -1646 17254 -1642
rect 17190 -1702 17194 -1646
rect 17194 -1702 17250 -1646
rect 17250 -1702 17254 -1646
rect 17190 -1706 17254 -1702
rect 17395 -1646 17459 -1642
rect 17395 -1702 17399 -1646
rect 17399 -1702 17455 -1646
rect 17455 -1702 17459 -1646
rect 17395 -1706 17459 -1702
rect 17603 -1641 17667 -1637
rect 17603 -1697 17607 -1641
rect 17607 -1697 17663 -1641
rect 17663 -1697 17667 -1641
rect 17603 -1701 17667 -1697
rect 17886 -1642 17950 -1638
rect 17886 -1698 17890 -1642
rect 17890 -1698 17946 -1642
rect 17946 -1698 17950 -1642
rect 17886 -1702 17950 -1698
rect 18079 -1644 18143 -1640
rect 18079 -1700 18083 -1644
rect 18083 -1700 18139 -1644
rect 18139 -1700 18143 -1644
rect 18079 -1704 18143 -1700
rect 18305 -1646 18369 -1642
rect 18305 -1702 18309 -1646
rect 18309 -1702 18365 -1646
rect 18365 -1702 18369 -1646
rect 18305 -1706 18369 -1702
rect 18570 -1646 18634 -1642
rect 18570 -1702 18574 -1646
rect 18574 -1702 18630 -1646
rect 18630 -1702 18634 -1646
rect 18570 -1706 18634 -1702
rect 18764 -1642 18828 -1638
rect 18764 -1698 18768 -1642
rect 18768 -1698 18824 -1642
rect 18824 -1698 18828 -1642
rect 18764 -1702 18828 -1698
rect 18962 -1651 19026 -1647
rect 18962 -1707 18966 -1651
rect 18966 -1707 19022 -1651
rect 19022 -1707 19026 -1651
rect 18962 -1711 19026 -1707
rect 19166 -1643 19230 -1639
rect 19166 -1699 19170 -1643
rect 19170 -1699 19226 -1643
rect 19226 -1699 19230 -1643
rect 19166 -1703 19230 -1699
rect 19386 -1640 19450 -1636
rect 19386 -1696 19390 -1640
rect 19390 -1696 19446 -1640
rect 19446 -1696 19450 -1640
rect 19386 -1700 19450 -1696
rect 19601 -1644 19665 -1640
rect 19601 -1700 19605 -1644
rect 19605 -1700 19661 -1644
rect 19661 -1700 19665 -1644
rect 19601 -1704 19665 -1700
rect 19829 -1641 19893 -1637
rect 19829 -1697 19833 -1641
rect 19833 -1697 19889 -1641
rect 19889 -1697 19893 -1641
rect 19829 -1701 19893 -1697
rect 20033 -1644 20097 -1640
rect 20033 -1700 20037 -1644
rect 20037 -1700 20093 -1644
rect 20093 -1700 20097 -1644
rect 20033 -1704 20097 -1700
rect 20271 -1642 20335 -1638
rect 20271 -1698 20275 -1642
rect 20275 -1698 20331 -1642
rect 20331 -1698 20335 -1642
rect 20271 -1702 20335 -1698
rect 20464 -1641 20528 -1637
rect 20464 -1697 20468 -1641
rect 20468 -1697 20524 -1641
rect 20524 -1697 20528 -1641
rect 20464 -1701 20528 -1697
rect 20661 -1646 20725 -1642
rect 20661 -1702 20665 -1646
rect 20665 -1702 20721 -1646
rect 20721 -1702 20725 -1646
rect 20661 -1706 20725 -1702
rect 20917 -1643 20981 -1639
rect 20917 -1699 20921 -1643
rect 20921 -1699 20977 -1643
rect 20977 -1699 20981 -1643
rect 20917 -1703 20981 -1699
rect 21156 -1647 21220 -1643
rect 21156 -1703 21160 -1647
rect 21160 -1703 21216 -1647
rect 21216 -1703 21220 -1647
rect 21156 -1707 21220 -1703
rect 21389 -1651 21453 -1647
rect 21389 -1707 21393 -1651
rect 21393 -1707 21449 -1651
rect 21449 -1707 21453 -1651
rect 21389 -1711 21453 -1707
rect 21610 -1646 21674 -1642
rect 21610 -1702 21614 -1646
rect 21614 -1702 21670 -1646
rect 21670 -1702 21674 -1646
rect 21610 -1706 21674 -1702
rect 21801 -1646 21865 -1642
rect 21801 -1702 21805 -1646
rect 21805 -1702 21861 -1646
rect 21861 -1702 21865 -1646
rect 21801 -1706 21865 -1702
rect 22029 -1644 22093 -1640
rect 22029 -1700 22033 -1644
rect 22033 -1700 22089 -1644
rect 22089 -1700 22093 -1644
rect 22029 -1704 22093 -1700
rect 22226 -1649 22290 -1645
rect 22226 -1705 22230 -1649
rect 22230 -1705 22286 -1649
rect 22286 -1705 22290 -1649
rect 22226 -1709 22290 -1705
rect 22438 -1649 22502 -1645
rect 22438 -1705 22442 -1649
rect 22442 -1705 22498 -1649
rect 22498 -1705 22502 -1649
rect 22438 -1709 22502 -1705
rect 22665 -1646 22729 -1642
rect 22665 -1702 22669 -1646
rect 22669 -1702 22725 -1646
rect 22725 -1702 22729 -1646
rect 22665 -1706 22729 -1702
rect 22854 -1645 22918 -1641
rect 22854 -1701 22858 -1645
rect 22858 -1701 22914 -1645
rect 22914 -1701 22918 -1645
rect 22854 -1705 22918 -1701
rect 23080 -1644 23144 -1640
rect 23080 -1700 23084 -1644
rect 23084 -1700 23140 -1644
rect 23140 -1700 23144 -1644
rect 23080 -1704 23144 -1700
rect 23334 -1644 23398 -1640
rect 23334 -1700 23338 -1644
rect 23338 -1700 23394 -1644
rect 23394 -1700 23398 -1644
rect 23334 -1704 23398 -1700
rect 23578 -1647 23642 -1643
rect 23578 -1703 23582 -1647
rect 23582 -1703 23638 -1647
rect 23638 -1703 23642 -1647
rect 23578 -1707 23642 -1703
rect 23808 -1648 23872 -1644
rect 23808 -1704 23812 -1648
rect 23812 -1704 23868 -1648
rect 23868 -1704 23872 -1648
rect 23808 -1708 23872 -1704
rect 24066 -1645 24130 -1641
rect 24066 -1701 24070 -1645
rect 24070 -1701 24126 -1645
rect 24126 -1701 24130 -1645
rect 24066 -1705 24130 -1701
rect 24276 -1645 24340 -1641
rect 24276 -1701 24280 -1645
rect 24280 -1701 24336 -1645
rect 24336 -1701 24340 -1645
rect 24276 -1705 24340 -1701
rect 24501 -1645 24565 -1641
rect 24501 -1701 24505 -1645
rect 24505 -1701 24561 -1645
rect 24561 -1701 24565 -1645
rect 24501 -1705 24565 -1701
rect 24720 -1648 24784 -1644
rect 24720 -1704 24724 -1648
rect 24724 -1704 24780 -1648
rect 24780 -1704 24784 -1648
rect 24720 -1708 24784 -1704
rect 25066 -1644 25130 -1640
rect 25066 -1700 25070 -1644
rect 25070 -1700 25126 -1644
rect 25126 -1700 25130 -1644
rect 25066 -1704 25130 -1700
rect 25265 -1647 25329 -1643
rect 25265 -1703 25269 -1647
rect 25269 -1703 25325 -1647
rect 25325 -1703 25329 -1647
rect 25265 -1707 25329 -1703
<< metal4 >>
rect 13318 13748 27105 13749
rect 13318 13747 27155 13748
rect 10645 13632 27155 13747
rect 10645 13568 13950 13632
rect 14014 13626 20659 13632
rect 14014 13625 19967 13626
rect 14014 13622 14779 13625
rect 14014 13568 14047 13622
rect 10645 13559 14047 13568
rect 3031 13162 3157 13167
rect 2064 13159 9079 13162
rect 10645 13159 13736 13559
rect 13943 13558 14047 13559
rect 14111 13558 14127 13622
rect 14191 13558 14207 13622
rect 14271 13558 14287 13622
rect 14351 13558 14367 13622
rect 14431 13558 14447 13622
rect 14511 13561 14779 13622
rect 14843 13561 14859 13625
rect 14923 13561 14939 13625
rect 15003 13561 15019 13625
rect 15083 13561 15099 13625
rect 15163 13561 15179 13625
rect 15243 13561 15385 13625
rect 15449 13561 15465 13625
rect 15529 13561 15545 13625
rect 15609 13561 15625 13625
rect 15689 13561 15705 13625
rect 15769 13561 15785 13625
rect 15849 13561 15991 13625
rect 16055 13561 16071 13625
rect 16135 13561 16151 13625
rect 16215 13561 16231 13625
rect 16295 13561 16311 13625
rect 16375 13561 16391 13625
rect 16455 13561 16597 13625
rect 16661 13561 16677 13625
rect 16741 13561 16757 13625
rect 16821 13561 16837 13625
rect 16901 13561 16917 13625
rect 16981 13561 16997 13625
rect 17061 13561 17203 13625
rect 17267 13561 17283 13625
rect 17347 13561 17363 13625
rect 17427 13561 17443 13625
rect 17507 13561 17523 13625
rect 17587 13561 17603 13625
rect 17667 13561 17809 13625
rect 17873 13561 17889 13625
rect 17953 13561 17969 13625
rect 18033 13561 18049 13625
rect 18113 13561 18129 13625
rect 18193 13561 18209 13625
rect 18273 13561 18415 13625
rect 18479 13561 18495 13625
rect 18559 13561 18575 13625
rect 18639 13561 18655 13625
rect 18719 13561 18735 13625
rect 18799 13561 18815 13625
rect 18879 13561 19021 13625
rect 19085 13561 19101 13625
rect 19165 13561 19181 13625
rect 19245 13561 19261 13625
rect 19325 13561 19341 13625
rect 19405 13561 19421 13625
rect 19485 13570 19967 13625
rect 19485 13561 19759 13570
rect 14511 13559 19759 13561
rect 14511 13558 14616 13559
rect 13943 13557 14616 13558
rect 13943 13556 14615 13557
rect 2064 13157 13736 13159
rect 2064 13093 3062 13157
rect 3126 13150 13736 13157
rect 3126 13147 3891 13150
rect 3126 13093 3159 13147
rect 2064 13084 3159 13093
rect 2064 12552 2848 13084
rect 3055 13083 3159 13084
rect 3223 13083 3239 13147
rect 3303 13083 3319 13147
rect 3383 13083 3399 13147
rect 3463 13083 3479 13147
rect 3543 13083 3559 13147
rect 3623 13086 3891 13147
rect 3955 13086 3971 13150
rect 4035 13086 4051 13150
rect 4115 13086 4131 13150
rect 4195 13086 4211 13150
rect 4275 13086 4291 13150
rect 4355 13086 4497 13150
rect 4561 13086 4577 13150
rect 4641 13086 4657 13150
rect 4721 13086 4737 13150
rect 4801 13086 4817 13150
rect 4881 13086 4897 13150
rect 4961 13086 5103 13150
rect 5167 13086 5183 13150
rect 5247 13086 5263 13150
rect 5327 13086 5343 13150
rect 5407 13086 5423 13150
rect 5487 13086 5503 13150
rect 5567 13086 5709 13150
rect 5773 13086 5789 13150
rect 5853 13086 5869 13150
rect 5933 13086 5949 13150
rect 6013 13086 6029 13150
rect 6093 13086 6109 13150
rect 6173 13086 6315 13150
rect 6379 13086 6395 13150
rect 6459 13086 6475 13150
rect 6539 13086 6555 13150
rect 6619 13086 6635 13150
rect 6699 13086 6715 13150
rect 6779 13086 6921 13150
rect 6985 13086 7001 13150
rect 7065 13086 7081 13150
rect 7145 13086 7161 13150
rect 7225 13086 7241 13150
rect 7305 13086 7321 13150
rect 7385 13086 7527 13150
rect 7591 13086 7607 13150
rect 7671 13086 7687 13150
rect 7751 13086 7767 13150
rect 7831 13086 7847 13150
rect 7911 13086 7927 13150
rect 7991 13086 8133 13150
rect 8197 13086 8213 13150
rect 8277 13086 8293 13150
rect 8357 13086 8373 13150
rect 8437 13086 8453 13150
rect 8517 13086 8533 13150
rect 8597 13095 13736 13150
rect 8597 13086 8871 13095
rect 3623 13084 8871 13086
rect 3623 13083 3728 13084
rect 3055 13082 3728 13083
rect 3055 13081 3727 13082
rect 2064 8094 2370 12552
rect 2430 12488 2445 12552
rect 2509 12551 2720 12552
rect 2509 12488 2576 12551
rect 2430 12487 2576 12488
rect 2640 12488 2720 12551
rect 2784 12546 2848 12552
rect 3055 12927 3121 13017
rect 3055 12863 3056 12927
rect 3120 12863 3121 12927
rect 3055 12847 3121 12863
rect 3055 12783 3056 12847
rect 3120 12783 3121 12847
rect 3055 12767 3121 12783
rect 3055 12703 3056 12767
rect 3120 12703 3121 12767
rect 3055 12687 3121 12703
rect 3055 12623 3056 12687
rect 3120 12623 3121 12687
rect 3055 12607 3121 12623
rect 2784 12488 2847 12546
rect 2640 12487 2847 12488
rect 2430 12469 2847 12487
rect 3055 12543 3056 12607
rect 3120 12543 3121 12607
rect 3055 12527 3121 12543
rect 3055 12463 3056 12527
rect 3120 12463 3121 12527
rect 3055 12447 3121 12463
rect 3055 12383 3056 12447
rect 3120 12383 3121 12447
rect 3055 12367 3121 12383
rect 3055 12303 3056 12367
rect 3120 12303 3121 12367
rect 3055 12287 3121 12303
rect 3055 12223 3056 12287
rect 3120 12223 3121 12287
rect 3055 12207 3121 12223
rect 3055 12143 3056 12207
rect 3120 12143 3121 12207
rect 2456 12006 2833 12021
rect 2456 11942 2463 12006
rect 2527 11942 2583 12006
rect 2647 11942 2726 12006
rect 2790 11942 2833 12006
rect 3055 11989 3121 12143
rect 3181 12051 3241 13081
rect 3301 11989 3361 13021
rect 3421 12051 3481 13081
rect 3541 11989 3601 13021
rect 3661 12927 3727 13017
rect 3661 12863 3662 12927
rect 3726 12863 3727 12927
rect 3661 12847 3727 12863
rect 3661 12783 3662 12847
rect 3726 12783 3727 12847
rect 3661 12767 3727 12783
rect 3661 12703 3662 12767
rect 3726 12703 3727 12767
rect 3661 12687 3727 12703
rect 3661 12623 3662 12687
rect 3726 12623 3727 12687
rect 3661 12607 3727 12623
rect 3661 12543 3662 12607
rect 3726 12543 3727 12607
rect 3661 12527 3727 12543
rect 3661 12463 3662 12527
rect 3726 12463 3727 12527
rect 3661 12447 3727 12463
rect 3661 12383 3662 12447
rect 3726 12383 3727 12447
rect 3661 12367 3727 12383
rect 3661 12303 3662 12367
rect 3726 12303 3727 12367
rect 3661 12287 3727 12303
rect 3661 12223 3662 12287
rect 3726 12223 3727 12287
rect 3661 12207 3727 12223
rect 3661 12143 3662 12207
rect 3726 12143 3727 12207
rect 3661 11989 3727 12143
rect 3055 11987 3727 11989
rect 2458 10583 2834 11942
rect 3055 11923 3159 11987
rect 3223 11923 3239 11987
rect 3303 11923 3319 11987
rect 3383 11923 3399 11987
rect 3463 11923 3479 11987
rect 3543 11923 3559 11987
rect 3623 11923 3727 11987
rect 3787 12930 3853 13020
rect 3787 12866 3788 12930
rect 3852 12866 3853 12930
rect 3787 12850 3853 12866
rect 3787 12786 3788 12850
rect 3852 12786 3853 12850
rect 3787 12770 3853 12786
rect 3787 12706 3788 12770
rect 3852 12706 3853 12770
rect 3787 12690 3853 12706
rect 3787 12626 3788 12690
rect 3852 12626 3853 12690
rect 3787 12610 3853 12626
rect 3787 12546 3788 12610
rect 3852 12546 3853 12610
rect 3787 12530 3853 12546
rect 3787 12466 3788 12530
rect 3852 12466 3853 12530
rect 3787 12450 3853 12466
rect 3787 12386 3788 12450
rect 3852 12386 3853 12450
rect 3787 12370 3853 12386
rect 3787 12306 3788 12370
rect 3852 12306 3853 12370
rect 3787 12290 3853 12306
rect 3787 12226 3788 12290
rect 3852 12226 3853 12290
rect 3787 12210 3853 12226
rect 3787 12146 3788 12210
rect 3852 12146 3853 12210
rect 3787 11992 3853 12146
rect 3913 12054 3973 13084
rect 4033 11992 4093 13024
rect 4153 12054 4213 13084
rect 4273 11992 4333 13024
rect 4393 12930 4459 13020
rect 4393 12866 4394 12930
rect 4458 12866 4459 12930
rect 4393 12850 4459 12866
rect 4393 12786 4394 12850
rect 4458 12786 4459 12850
rect 4393 12770 4459 12786
rect 4393 12706 4394 12770
rect 4458 12706 4459 12770
rect 4393 12690 4459 12706
rect 4393 12626 4394 12690
rect 4458 12626 4459 12690
rect 4393 12610 4459 12626
rect 4393 12546 4394 12610
rect 4458 12546 4459 12610
rect 4393 12530 4459 12546
rect 4393 12466 4394 12530
rect 4458 12466 4459 12530
rect 4393 12450 4459 12466
rect 4393 12386 4394 12450
rect 4458 12386 4459 12450
rect 4393 12370 4459 12386
rect 4393 12306 4394 12370
rect 4458 12306 4459 12370
rect 4393 12290 4459 12306
rect 4393 12226 4394 12290
rect 4458 12226 4459 12290
rect 4393 12210 4459 12226
rect 4393 12146 4394 12210
rect 4458 12146 4459 12210
rect 4393 11992 4459 12146
rect 4519 11992 4579 13024
rect 4639 12054 4699 13084
rect 4759 11992 4819 13024
rect 4879 12054 4939 13084
rect 4999 12930 5065 13020
rect 4999 12866 5000 12930
rect 5064 12866 5065 12930
rect 4999 12850 5065 12866
rect 4999 12786 5000 12850
rect 5064 12786 5065 12850
rect 4999 12770 5065 12786
rect 4999 12706 5000 12770
rect 5064 12706 5065 12770
rect 4999 12690 5065 12706
rect 4999 12626 5000 12690
rect 5064 12626 5065 12690
rect 4999 12610 5065 12626
rect 4999 12546 5000 12610
rect 5064 12546 5065 12610
rect 4999 12530 5065 12546
rect 4999 12466 5000 12530
rect 5064 12466 5065 12530
rect 4999 12450 5065 12466
rect 4999 12386 5000 12450
rect 5064 12386 5065 12450
rect 4999 12370 5065 12386
rect 4999 12306 5000 12370
rect 5064 12306 5065 12370
rect 4999 12290 5065 12306
rect 4999 12226 5000 12290
rect 5064 12226 5065 12290
rect 4999 12210 5065 12226
rect 4999 12146 5000 12210
rect 5064 12146 5065 12210
rect 4999 11992 5065 12146
rect 5125 12054 5185 13084
rect 5245 11992 5305 13024
rect 5365 12054 5425 13084
rect 5485 11992 5545 13024
rect 5605 12930 5671 13020
rect 5605 12866 5606 12930
rect 5670 12866 5671 12930
rect 5605 12850 5671 12866
rect 5605 12786 5606 12850
rect 5670 12786 5671 12850
rect 5605 12770 5671 12786
rect 5605 12706 5606 12770
rect 5670 12706 5671 12770
rect 5605 12690 5671 12706
rect 5605 12626 5606 12690
rect 5670 12626 5671 12690
rect 5605 12610 5671 12626
rect 5605 12546 5606 12610
rect 5670 12546 5671 12610
rect 5605 12530 5671 12546
rect 5605 12466 5606 12530
rect 5670 12466 5671 12530
rect 5605 12450 5671 12466
rect 5605 12386 5606 12450
rect 5670 12386 5671 12450
rect 5605 12370 5671 12386
rect 5605 12306 5606 12370
rect 5670 12306 5671 12370
rect 5605 12290 5671 12306
rect 5605 12226 5606 12290
rect 5670 12226 5671 12290
rect 5605 12210 5671 12226
rect 5605 12146 5606 12210
rect 5670 12146 5671 12210
rect 5605 11992 5671 12146
rect 5731 11992 5791 13024
rect 5851 12054 5911 13084
rect 5971 11992 6031 13024
rect 6091 12054 6151 13084
rect 6211 12930 6277 13020
rect 6211 12866 6212 12930
rect 6276 12866 6277 12930
rect 6211 12850 6277 12866
rect 6211 12786 6212 12850
rect 6276 12786 6277 12850
rect 6211 12770 6277 12786
rect 6211 12706 6212 12770
rect 6276 12706 6277 12770
rect 6211 12690 6277 12706
rect 6211 12626 6212 12690
rect 6276 12626 6277 12690
rect 6211 12610 6277 12626
rect 6211 12546 6212 12610
rect 6276 12546 6277 12610
rect 6211 12530 6277 12546
rect 6211 12466 6212 12530
rect 6276 12466 6277 12530
rect 6211 12450 6277 12466
rect 6211 12386 6212 12450
rect 6276 12386 6277 12450
rect 6211 12370 6277 12386
rect 6211 12306 6212 12370
rect 6276 12306 6277 12370
rect 6211 12290 6277 12306
rect 6211 12226 6212 12290
rect 6276 12226 6277 12290
rect 6211 12210 6277 12226
rect 6211 12146 6212 12210
rect 6276 12146 6277 12210
rect 6211 11992 6277 12146
rect 6337 12054 6397 13084
rect 6457 11992 6517 13024
rect 6577 12054 6637 13084
rect 6697 11992 6757 13024
rect 6817 12930 6883 13020
rect 6817 12866 6818 12930
rect 6882 12866 6883 12930
rect 6817 12850 6883 12866
rect 6817 12786 6818 12850
rect 6882 12786 6883 12850
rect 6817 12770 6883 12786
rect 6817 12706 6818 12770
rect 6882 12706 6883 12770
rect 6817 12690 6883 12706
rect 6817 12626 6818 12690
rect 6882 12626 6883 12690
rect 6817 12610 6883 12626
rect 6817 12546 6818 12610
rect 6882 12546 6883 12610
rect 6817 12530 6883 12546
rect 6817 12466 6818 12530
rect 6882 12466 6883 12530
rect 6817 12450 6883 12466
rect 6817 12386 6818 12450
rect 6882 12386 6883 12450
rect 6817 12370 6883 12386
rect 6817 12306 6818 12370
rect 6882 12306 6883 12370
rect 6817 12290 6883 12306
rect 6817 12226 6818 12290
rect 6882 12226 6883 12290
rect 6817 12210 6883 12226
rect 6817 12146 6818 12210
rect 6882 12146 6883 12210
rect 6817 11992 6883 12146
rect 6943 11992 7003 13024
rect 7063 12054 7123 13084
rect 7183 11992 7243 13024
rect 7303 12054 7363 13084
rect 7423 12930 7489 13020
rect 7423 12866 7424 12930
rect 7488 12866 7489 12930
rect 7423 12850 7489 12866
rect 7423 12786 7424 12850
rect 7488 12786 7489 12850
rect 7423 12770 7489 12786
rect 7423 12706 7424 12770
rect 7488 12706 7489 12770
rect 7423 12690 7489 12706
rect 7423 12626 7424 12690
rect 7488 12626 7489 12690
rect 7423 12610 7489 12626
rect 7423 12546 7424 12610
rect 7488 12546 7489 12610
rect 7423 12530 7489 12546
rect 7423 12466 7424 12530
rect 7488 12466 7489 12530
rect 7423 12450 7489 12466
rect 7423 12386 7424 12450
rect 7488 12386 7489 12450
rect 7423 12370 7489 12386
rect 7423 12306 7424 12370
rect 7488 12306 7489 12370
rect 7423 12290 7489 12306
rect 7423 12226 7424 12290
rect 7488 12226 7489 12290
rect 7423 12210 7489 12226
rect 7423 12146 7424 12210
rect 7488 12146 7489 12210
rect 7423 11992 7489 12146
rect 7549 12054 7609 13084
rect 7669 11992 7729 13024
rect 7789 12054 7849 13084
rect 7909 11992 7969 13024
rect 8029 12930 8095 13020
rect 8029 12866 8030 12930
rect 8094 12866 8095 12930
rect 8029 12850 8095 12866
rect 8029 12786 8030 12850
rect 8094 12786 8095 12850
rect 8029 12770 8095 12786
rect 8029 12706 8030 12770
rect 8094 12706 8095 12770
rect 8029 12690 8095 12706
rect 8029 12626 8030 12690
rect 8094 12626 8095 12690
rect 8029 12610 8095 12626
rect 8029 12546 8030 12610
rect 8094 12546 8095 12610
rect 8029 12530 8095 12546
rect 8029 12466 8030 12530
rect 8094 12466 8095 12530
rect 8029 12450 8095 12466
rect 8029 12386 8030 12450
rect 8094 12386 8095 12450
rect 8029 12370 8095 12386
rect 8029 12306 8030 12370
rect 8094 12306 8095 12370
rect 8029 12290 8095 12306
rect 8029 12226 8030 12290
rect 8094 12226 8095 12290
rect 8029 12210 8095 12226
rect 8029 12146 8030 12210
rect 8094 12146 8095 12210
rect 8029 11992 8095 12146
rect 8155 11992 8215 13024
rect 8275 12054 8335 13084
rect 8395 11992 8455 13024
rect 8515 12054 8575 13084
rect 8761 13031 8871 13084
rect 8935 13031 13736 13095
rect 8761 13027 13736 13031
rect 8635 12930 8701 13020
rect 8635 12866 8636 12930
rect 8700 12866 8701 12930
rect 8635 12850 8701 12866
rect 8635 12786 8636 12850
rect 8700 12786 8701 12850
rect 8635 12770 8701 12786
rect 8635 12706 8636 12770
rect 8700 12706 8701 12770
rect 8635 12690 8701 12706
rect 8635 12626 8636 12690
rect 8700 12626 8701 12690
rect 8635 12610 8701 12626
rect 8635 12546 8636 12610
rect 8700 12546 8701 12610
rect 8635 12530 8701 12546
rect 8635 12466 8636 12530
rect 8700 12466 8701 12530
rect 8635 12450 8701 12466
rect 8635 12386 8636 12450
rect 8700 12386 8701 12450
rect 8635 12370 8701 12386
rect 8635 12306 8636 12370
rect 8700 12306 8701 12370
rect 8635 12290 8701 12306
rect 8635 12226 8636 12290
rect 8700 12226 8701 12290
rect 8635 12210 8701 12226
rect 8635 12146 8636 12210
rect 8700 12146 8701 12210
rect 8761 12963 13333 13027
rect 13397 13026 13608 13027
rect 13397 12963 13464 13026
rect 8761 12962 13464 12963
rect 13528 12963 13608 13026
rect 13672 13021 13736 13027
rect 13943 13402 14009 13492
rect 13943 13338 13944 13402
rect 14008 13338 14009 13402
rect 13943 13322 14009 13338
rect 13943 13258 13944 13322
rect 14008 13258 14009 13322
rect 13943 13242 14009 13258
rect 13943 13178 13944 13242
rect 14008 13178 14009 13242
rect 13943 13162 14009 13178
rect 13943 13098 13944 13162
rect 14008 13098 14009 13162
rect 13943 13082 14009 13098
rect 13672 12963 13735 13021
rect 13528 12962 13735 12963
rect 8761 12951 13735 12962
rect 8761 12887 8876 12951
rect 8940 12944 13735 12951
rect 13943 13018 13944 13082
rect 14008 13018 14009 13082
rect 13943 13002 14009 13018
rect 8940 12887 13437 12944
rect 8761 12799 13437 12887
rect 8761 12735 8877 12799
rect 8941 12760 13437 12799
rect 13943 12938 13944 13002
rect 14008 12938 14009 13002
rect 13943 12922 14009 12938
rect 13943 12858 13944 12922
rect 14008 12858 14009 12922
rect 13943 12842 14009 12858
rect 13943 12778 13944 12842
rect 14008 12778 14009 12842
rect 13943 12762 14009 12778
rect 8941 12735 10819 12760
rect 8761 12629 10819 12735
rect 13943 12698 13944 12762
rect 14008 12698 14009 12762
rect 13943 12682 14009 12698
rect 8761 12565 8877 12629
rect 8941 12571 10819 12629
rect 8941 12565 9079 12571
rect 8761 12472 9079 12565
rect 8761 12408 8876 12472
rect 8940 12408 9079 12472
rect 8761 12383 9079 12408
rect 8761 12282 9335 12383
rect 8761 12230 9171 12282
rect 8761 12166 8794 12230
rect 8858 12218 9171 12230
rect 9235 12218 9335 12282
rect 8858 12188 9335 12218
rect 8858 12166 9079 12188
rect 8761 12154 9079 12166
rect 8635 11992 8701 12146
rect 3787 11990 8701 11992
rect 3787 11926 3891 11990
rect 3955 11926 3971 11990
rect 4035 11926 4051 11990
rect 4115 11926 4131 11990
rect 4195 11926 4211 11990
rect 4275 11926 4291 11990
rect 4355 11926 4497 11990
rect 4561 11926 4577 11990
rect 4641 11926 4657 11990
rect 4721 11926 4737 11990
rect 4801 11926 4817 11990
rect 4881 11926 4897 11990
rect 4961 11926 5103 11990
rect 5167 11926 5183 11990
rect 5247 11926 5263 11990
rect 5327 11926 5343 11990
rect 5407 11926 5423 11990
rect 5487 11926 5503 11990
rect 5567 11926 5709 11990
rect 5773 11926 5789 11990
rect 5853 11926 5869 11990
rect 5933 11926 5949 11990
rect 6013 11926 6029 11990
rect 6093 11926 6109 11990
rect 6173 11926 6315 11990
rect 6379 11926 6395 11990
rect 6459 11926 6475 11990
rect 6539 11926 6555 11990
rect 6619 11926 6635 11990
rect 6699 11926 6715 11990
rect 6779 11926 6921 11990
rect 6985 11926 7001 11990
rect 7065 11926 7081 11990
rect 7145 11926 7161 11990
rect 7225 11926 7241 11990
rect 7305 11926 7321 11990
rect 7385 11926 7527 11990
rect 7591 11926 7607 11990
rect 7671 11926 7687 11990
rect 7751 11926 7767 11990
rect 7831 11926 7847 11990
rect 7911 11926 7927 11990
rect 7991 11926 8133 11990
rect 8197 11926 8213 11990
rect 8277 11926 8293 11990
rect 8357 11926 8373 11990
rect 8437 11926 8453 11990
rect 8517 11926 8533 11990
rect 8597 11926 8701 11990
rect 3787 11924 8701 11926
rect 8761 11969 8959 11979
rect 3055 11921 3727 11923
rect 8761 11905 8882 11969
rect 8946 11905 8959 11969
rect 8761 11895 8959 11905
rect 3406 11742 4078 11744
rect 3406 11678 3510 11742
rect 3574 11678 3590 11742
rect 3654 11678 3670 11742
rect 3734 11678 3750 11742
rect 3814 11678 3830 11742
rect 3894 11678 3910 11742
rect 3974 11678 4078 11742
rect 3406 11676 4078 11678
rect 3406 11522 3472 11676
rect 3406 11458 3407 11522
rect 3471 11458 3472 11522
rect 3406 11442 3472 11458
rect 3406 11378 3407 11442
rect 3471 11378 3472 11442
rect 3406 11362 3472 11378
rect 3406 11298 3407 11362
rect 3471 11298 3472 11362
rect 3406 11282 3472 11298
rect 3406 11218 3407 11282
rect 3471 11218 3472 11282
rect 3406 11202 3472 11218
rect 3406 11138 3407 11202
rect 3471 11138 3472 11202
rect 3406 11122 3472 11138
rect 3406 11058 3407 11122
rect 3471 11058 3472 11122
rect 3406 11042 3472 11058
rect 3406 10978 3407 11042
rect 3471 10978 3472 11042
rect 3406 10962 3472 10978
rect 3406 10898 3407 10962
rect 3471 10898 3472 10962
rect 3406 10882 3472 10898
rect 3406 10818 3407 10882
rect 3471 10818 3472 10882
rect 3406 10802 3472 10818
rect 3406 10738 3407 10802
rect 3471 10738 3472 10802
rect 3406 10648 3472 10738
rect 3018 10583 3143 10589
rect 3532 10584 3592 11614
rect 3652 10644 3712 11676
rect 3772 10584 3832 11614
rect 3892 10644 3952 11676
rect 4012 11522 4078 11676
rect 4012 11458 4013 11522
rect 4077 11458 4078 11522
rect 4012 11442 4078 11458
rect 4012 11378 4013 11442
rect 4077 11378 4078 11442
rect 4012 11362 4078 11378
rect 4012 11298 4013 11362
rect 4077 11298 4078 11362
rect 4012 11282 4078 11298
rect 4012 11218 4013 11282
rect 4077 11218 4078 11282
rect 4012 11202 4078 11218
rect 4012 11138 4013 11202
rect 4077 11138 4078 11202
rect 4012 11122 4078 11138
rect 4012 11058 4013 11122
rect 4077 11058 4078 11122
rect 4012 11042 4078 11058
rect 4012 10978 4013 11042
rect 4077 10978 4078 11042
rect 4012 10962 4078 10978
rect 4012 10898 4013 10962
rect 4077 10898 4078 10962
rect 4012 10882 4078 10898
rect 4012 10818 4013 10882
rect 4077 10818 4078 10882
rect 4012 10802 4078 10818
rect 4012 10738 4013 10802
rect 4077 10738 4078 10802
rect 4012 10648 4078 10738
rect 4138 11742 6628 11744
rect 4138 11678 4242 11742
rect 4306 11678 4322 11742
rect 4386 11678 4402 11742
rect 4466 11678 4482 11742
rect 4546 11678 4562 11742
rect 4626 11678 4642 11742
rect 4706 11678 4848 11742
rect 4912 11678 4928 11742
rect 4992 11678 5008 11742
rect 5072 11678 5088 11742
rect 5152 11678 5168 11742
rect 5232 11678 5248 11742
rect 5312 11678 5454 11742
rect 5518 11678 5534 11742
rect 5598 11678 5614 11742
rect 5678 11678 5694 11742
rect 5758 11678 5774 11742
rect 5838 11678 5854 11742
rect 5918 11678 6060 11742
rect 6124 11678 6140 11742
rect 6204 11678 6220 11742
rect 6284 11678 6300 11742
rect 6364 11678 6380 11742
rect 6444 11678 6460 11742
rect 6524 11678 6628 11742
rect 4138 11676 6628 11678
rect 4138 11522 4204 11676
rect 4138 11458 4139 11522
rect 4203 11458 4204 11522
rect 4138 11442 4204 11458
rect 4138 11378 4139 11442
rect 4203 11378 4204 11442
rect 4138 11362 4204 11378
rect 4138 11298 4139 11362
rect 4203 11298 4204 11362
rect 4138 11282 4204 11298
rect 4138 11218 4139 11282
rect 4203 11218 4204 11282
rect 4138 11202 4204 11218
rect 4138 11138 4139 11202
rect 4203 11138 4204 11202
rect 4138 11122 4204 11138
rect 4138 11058 4139 11122
rect 4203 11058 4204 11122
rect 4138 11042 4204 11058
rect 4138 10978 4139 11042
rect 4203 10978 4204 11042
rect 4138 10962 4204 10978
rect 4138 10898 4139 10962
rect 4203 10898 4204 10962
rect 4138 10882 4204 10898
rect 4138 10818 4139 10882
rect 4203 10818 4204 10882
rect 4138 10802 4204 10818
rect 4138 10738 4139 10802
rect 4203 10738 4204 10802
rect 4138 10648 4204 10738
rect 4264 10584 4324 11614
rect 4384 10644 4444 11676
rect 4504 10584 4564 11614
rect 4624 10644 4684 11676
rect 4744 11522 4810 11676
rect 4744 11458 4745 11522
rect 4809 11458 4810 11522
rect 4744 11442 4810 11458
rect 4744 11378 4745 11442
rect 4809 11378 4810 11442
rect 4744 11362 4810 11378
rect 4744 11298 4745 11362
rect 4809 11298 4810 11362
rect 4744 11282 4810 11298
rect 4744 11218 4745 11282
rect 4809 11218 4810 11282
rect 4744 11202 4810 11218
rect 4744 11138 4745 11202
rect 4809 11138 4810 11202
rect 4744 11122 4810 11138
rect 4744 11058 4745 11122
rect 4809 11058 4810 11122
rect 4744 11042 4810 11058
rect 4744 10978 4745 11042
rect 4809 10978 4810 11042
rect 4744 10962 4810 10978
rect 4744 10898 4745 10962
rect 4809 10898 4810 10962
rect 4744 10882 4810 10898
rect 4744 10818 4745 10882
rect 4809 10818 4810 10882
rect 4744 10802 4810 10818
rect 4744 10738 4745 10802
rect 4809 10738 4810 10802
rect 4744 10648 4810 10738
rect 4870 10644 4930 11676
rect 4990 10584 5050 11614
rect 5110 10644 5170 11676
rect 5230 10584 5290 11614
rect 5350 11522 5416 11676
rect 5350 11458 5351 11522
rect 5415 11458 5416 11522
rect 5350 11442 5416 11458
rect 5350 11378 5351 11442
rect 5415 11378 5416 11442
rect 5350 11362 5416 11378
rect 5350 11298 5351 11362
rect 5415 11298 5416 11362
rect 5350 11282 5416 11298
rect 5350 11218 5351 11282
rect 5415 11218 5416 11282
rect 5350 11202 5416 11218
rect 5350 11138 5351 11202
rect 5415 11138 5416 11202
rect 5350 11122 5416 11138
rect 5350 11058 5351 11122
rect 5415 11058 5416 11122
rect 5350 11042 5416 11058
rect 5350 10978 5351 11042
rect 5415 10978 5416 11042
rect 5350 10962 5416 10978
rect 5350 10898 5351 10962
rect 5415 10898 5416 10962
rect 5350 10882 5416 10898
rect 5350 10818 5351 10882
rect 5415 10818 5416 10882
rect 5350 10802 5416 10818
rect 5350 10738 5351 10802
rect 5415 10738 5416 10802
rect 5350 10648 5416 10738
rect 5476 10584 5536 11614
rect 5596 10644 5656 11676
rect 5716 10584 5776 11614
rect 5836 10644 5896 11676
rect 5956 11522 6022 11676
rect 5956 11458 5957 11522
rect 6021 11458 6022 11522
rect 5956 11442 6022 11458
rect 5956 11378 5957 11442
rect 6021 11378 6022 11442
rect 5956 11362 6022 11378
rect 5956 11298 5957 11362
rect 6021 11298 6022 11362
rect 5956 11282 6022 11298
rect 5956 11218 5957 11282
rect 6021 11218 6022 11282
rect 5956 11202 6022 11218
rect 5956 11138 5957 11202
rect 6021 11138 6022 11202
rect 5956 11122 6022 11138
rect 5956 11058 5957 11122
rect 6021 11058 6022 11122
rect 5956 11042 6022 11058
rect 5956 10978 5957 11042
rect 6021 10978 6022 11042
rect 5956 10962 6022 10978
rect 5956 10898 5957 10962
rect 6021 10898 6022 10962
rect 5956 10882 6022 10898
rect 5956 10818 5957 10882
rect 6021 10818 6022 10882
rect 5956 10802 6022 10818
rect 5956 10738 5957 10802
rect 6021 10738 6022 10802
rect 5956 10648 6022 10738
rect 6082 10644 6142 11676
rect 6202 10584 6262 11614
rect 6322 10644 6382 11676
rect 6442 10584 6502 11614
rect 6562 11522 6628 11676
rect 6562 11458 6563 11522
rect 6627 11458 6628 11522
rect 6562 11442 6628 11458
rect 6562 11378 6563 11442
rect 6627 11378 6628 11442
rect 6562 11362 6628 11378
rect 6562 11298 6563 11362
rect 6627 11298 6628 11362
rect 6562 11282 6628 11298
rect 6562 11218 6563 11282
rect 6627 11218 6628 11282
rect 6562 11202 6628 11218
rect 6562 11138 6563 11202
rect 6627 11138 6628 11202
rect 6562 11122 6628 11138
rect 6562 11058 6563 11122
rect 6627 11058 6628 11122
rect 6562 11042 6628 11058
rect 6562 10978 6563 11042
rect 6627 10978 6628 11042
rect 6562 10962 6628 10978
rect 6562 10898 6563 10962
rect 6627 10898 6628 10962
rect 6562 10882 6628 10898
rect 6562 10818 6563 10882
rect 6627 10818 6628 10882
rect 6562 10802 6628 10818
rect 6562 10738 6563 10802
rect 6627 10738 6628 10802
rect 6562 10648 6628 10738
rect 6688 11742 7966 11744
rect 6688 11678 6792 11742
rect 6856 11678 6872 11742
rect 6936 11678 6952 11742
rect 7016 11678 7032 11742
rect 7096 11678 7112 11742
rect 7176 11678 7192 11742
rect 7256 11678 7398 11742
rect 7462 11678 7478 11742
rect 7542 11678 7558 11742
rect 7622 11678 7638 11742
rect 7702 11678 7718 11742
rect 7782 11678 7798 11742
rect 7862 11678 7966 11742
rect 6688 11676 7966 11678
rect 6688 11522 6754 11676
rect 6688 11458 6689 11522
rect 6753 11458 6754 11522
rect 6688 11442 6754 11458
rect 6688 11378 6689 11442
rect 6753 11378 6754 11442
rect 6688 11362 6754 11378
rect 6688 11298 6689 11362
rect 6753 11298 6754 11362
rect 6688 11282 6754 11298
rect 6688 11218 6689 11282
rect 6753 11218 6754 11282
rect 6688 11202 6754 11218
rect 6688 11138 6689 11202
rect 6753 11138 6754 11202
rect 6688 11122 6754 11138
rect 6688 11058 6689 11122
rect 6753 11058 6754 11122
rect 6688 11042 6754 11058
rect 6688 10978 6689 11042
rect 6753 10978 6754 11042
rect 6688 10962 6754 10978
rect 6688 10898 6689 10962
rect 6753 10898 6754 10962
rect 6688 10882 6754 10898
rect 6688 10818 6689 10882
rect 6753 10818 6754 10882
rect 6688 10802 6754 10818
rect 6688 10738 6689 10802
rect 6753 10738 6754 10802
rect 6688 10648 6754 10738
rect 6814 10584 6874 11614
rect 6934 10644 6994 11676
rect 7054 10584 7114 11614
rect 7174 10644 7234 11676
rect 7294 11522 7360 11676
rect 7294 11458 7295 11522
rect 7359 11458 7360 11522
rect 7294 11442 7360 11458
rect 7294 11378 7295 11442
rect 7359 11378 7360 11442
rect 7294 11362 7360 11378
rect 7294 11298 7295 11362
rect 7359 11298 7360 11362
rect 7294 11282 7360 11298
rect 7294 11218 7295 11282
rect 7359 11218 7360 11282
rect 7294 11202 7360 11218
rect 7294 11138 7295 11202
rect 7359 11138 7360 11202
rect 7294 11122 7360 11138
rect 7294 11058 7295 11122
rect 7359 11058 7360 11122
rect 7294 11042 7360 11058
rect 7294 10978 7295 11042
rect 7359 10978 7360 11042
rect 7294 10962 7360 10978
rect 7294 10898 7295 10962
rect 7359 10898 7360 10962
rect 7294 10882 7360 10898
rect 7294 10818 7295 10882
rect 7359 10818 7360 10882
rect 7294 10802 7360 10818
rect 7294 10738 7295 10802
rect 7359 10738 7360 10802
rect 7294 10648 7360 10738
rect 7420 10644 7480 11676
rect 7540 10584 7600 11614
rect 7660 10644 7720 11676
rect 7780 10584 7840 11614
rect 7900 11522 7966 11676
rect 7900 11458 7901 11522
rect 7965 11458 7966 11522
rect 7900 11442 7966 11458
rect 7900 11378 7901 11442
rect 7965 11378 7966 11442
rect 7900 11362 7966 11378
rect 7900 11298 7901 11362
rect 7965 11298 7966 11362
rect 7900 11282 7966 11298
rect 7900 11218 7901 11282
rect 7965 11218 7966 11282
rect 7900 11202 7966 11218
rect 7900 11138 7901 11202
rect 7965 11138 7966 11202
rect 7900 11122 7966 11138
rect 7900 11058 7901 11122
rect 7965 11058 7966 11122
rect 7900 11042 7966 11058
rect 7900 10978 7901 11042
rect 7965 10978 7966 11042
rect 7900 10962 7966 10978
rect 7900 10898 7901 10962
rect 7965 10898 7966 10962
rect 7900 10882 7966 10898
rect 7900 10818 7901 10882
rect 7965 10818 7966 10882
rect 7900 10802 7966 10818
rect 7900 10738 7901 10802
rect 7965 10738 7966 10802
rect 7900 10648 7966 10738
rect 8028 11742 8700 11744
rect 8028 11678 8132 11742
rect 8196 11678 8212 11742
rect 8276 11678 8292 11742
rect 8356 11678 8372 11742
rect 8436 11678 8452 11742
rect 8516 11678 8532 11742
rect 8596 11678 8700 11742
rect 8028 11676 8700 11678
rect 8028 11522 8094 11676
rect 8028 11458 8029 11522
rect 8093 11458 8094 11522
rect 8028 11442 8094 11458
rect 8028 11378 8029 11442
rect 8093 11378 8094 11442
rect 8028 11362 8094 11378
rect 8028 11298 8029 11362
rect 8093 11298 8094 11362
rect 8028 11282 8094 11298
rect 8028 11218 8029 11282
rect 8093 11218 8094 11282
rect 8028 11202 8094 11218
rect 8028 11138 8029 11202
rect 8093 11138 8094 11202
rect 8028 11122 8094 11138
rect 8028 11058 8029 11122
rect 8093 11058 8094 11122
rect 8028 11042 8094 11058
rect 8028 10978 8029 11042
rect 8093 10978 8094 11042
rect 8028 10962 8094 10978
rect 8028 10898 8029 10962
rect 8093 10898 8094 10962
rect 8028 10882 8094 10898
rect 8028 10818 8029 10882
rect 8093 10818 8094 10882
rect 8028 10802 8094 10818
rect 8028 10738 8029 10802
rect 8093 10738 8094 10802
rect 8028 10648 8094 10738
rect 8154 10644 8214 11676
rect 8274 10584 8334 11614
rect 8394 10644 8454 11676
rect 8514 10584 8574 11614
rect 8634 11522 8700 11676
rect 8634 11458 8635 11522
rect 8699 11458 8700 11522
rect 8634 11442 8700 11458
rect 8634 11378 8635 11442
rect 8699 11378 8700 11442
rect 8634 11362 8700 11378
rect 8634 11298 8635 11362
rect 8699 11298 8700 11362
rect 8634 11282 8700 11298
rect 8634 11218 8635 11282
rect 8699 11218 8700 11282
rect 8634 11202 8700 11218
rect 8634 11138 8635 11202
rect 8699 11138 8700 11202
rect 8634 11122 8700 11138
rect 8634 11058 8635 11122
rect 8699 11058 8700 11122
rect 8634 11042 8700 11058
rect 8634 10978 8635 11042
rect 8699 10978 8700 11042
rect 8634 10962 8700 10978
rect 8634 10898 8635 10962
rect 8699 10898 8700 10962
rect 8634 10882 8700 10898
rect 8634 10818 8635 10882
rect 8699 10818 8700 10882
rect 8634 10802 8700 10818
rect 8634 10738 8635 10802
rect 8699 10738 8700 10802
rect 8634 10648 8700 10738
rect 8761 11573 8821 11895
rect 9019 11776 9079 12154
rect 8881 11766 9079 11776
rect 8881 11702 8882 11766
rect 8946 11702 9079 11766
rect 8881 11692 9079 11702
rect 10646 12091 10819 12571
rect 10883 12573 13694 12680
rect 10883 12571 12537 12573
rect 10883 12569 12125 12571
rect 10883 12567 11926 12569
rect 10883 12565 11741 12567
rect 10883 12564 11538 12565
rect 10883 12562 11353 12564
rect 10883 12560 11168 12562
rect 10883 12496 10981 12560
rect 11045 12498 11168 12560
rect 11232 12500 11353 12562
rect 11417 12501 11538 12564
rect 11602 12503 11741 12565
rect 11805 12505 11926 12567
rect 11990 12507 12125 12569
rect 12189 12570 12537 12571
rect 12189 12507 12327 12570
rect 11990 12506 12327 12507
rect 12391 12509 12537 12570
rect 12601 12509 12761 12573
rect 12825 12572 13694 12573
rect 12825 12509 12967 12572
rect 12391 12508 12967 12509
rect 13031 12571 13694 12572
rect 13031 12508 13188 12571
rect 12391 12507 13188 12508
rect 13252 12507 13694 12571
rect 12391 12506 13694 12507
rect 11990 12505 13694 12506
rect 11805 12503 13694 12505
rect 11602 12501 13694 12503
rect 11417 12500 13694 12501
rect 11232 12498 13694 12500
rect 11045 12496 13694 12498
rect 13943 12618 13944 12682
rect 14008 12618 14009 12682
rect 10883 12481 13721 12496
rect 10883 12417 13351 12481
rect 13415 12417 13471 12481
rect 13535 12417 13614 12481
rect 13678 12417 13721 12481
rect 13943 12464 14009 12618
rect 14069 12526 14129 13556
rect 14189 12464 14249 13496
rect 14309 12526 14369 13556
rect 14429 12464 14489 13496
rect 14549 13402 14615 13492
rect 14549 13338 14550 13402
rect 14614 13338 14615 13402
rect 14549 13322 14615 13338
rect 14549 13258 14550 13322
rect 14614 13258 14615 13322
rect 14549 13242 14615 13258
rect 14549 13178 14550 13242
rect 14614 13178 14615 13242
rect 14549 13162 14615 13178
rect 14549 13098 14550 13162
rect 14614 13098 14615 13162
rect 14549 13082 14615 13098
rect 14549 13018 14550 13082
rect 14614 13018 14615 13082
rect 14549 13002 14615 13018
rect 14549 12938 14550 13002
rect 14614 12938 14615 13002
rect 14549 12922 14615 12938
rect 14549 12858 14550 12922
rect 14614 12858 14615 12922
rect 14549 12842 14615 12858
rect 14549 12778 14550 12842
rect 14614 12778 14615 12842
rect 14549 12762 14615 12778
rect 14549 12698 14550 12762
rect 14614 12698 14615 12762
rect 14549 12682 14615 12698
rect 14549 12618 14550 12682
rect 14614 12618 14615 12682
rect 14549 12464 14615 12618
rect 13943 12462 14615 12464
rect 10883 12172 13722 12417
rect 13943 12398 14047 12462
rect 14111 12398 14127 12462
rect 14191 12398 14207 12462
rect 14271 12398 14287 12462
rect 14351 12398 14367 12462
rect 14431 12398 14447 12462
rect 14511 12398 14615 12462
rect 14675 13405 14741 13495
rect 14675 13341 14676 13405
rect 14740 13341 14741 13405
rect 14675 13325 14741 13341
rect 14675 13261 14676 13325
rect 14740 13261 14741 13325
rect 14675 13245 14741 13261
rect 14675 13181 14676 13245
rect 14740 13181 14741 13245
rect 14675 13165 14741 13181
rect 14675 13101 14676 13165
rect 14740 13101 14741 13165
rect 14675 13085 14741 13101
rect 14675 13021 14676 13085
rect 14740 13021 14741 13085
rect 14675 13005 14741 13021
rect 14675 12941 14676 13005
rect 14740 12941 14741 13005
rect 14675 12925 14741 12941
rect 14675 12861 14676 12925
rect 14740 12861 14741 12925
rect 14675 12845 14741 12861
rect 14675 12781 14676 12845
rect 14740 12781 14741 12845
rect 14675 12765 14741 12781
rect 14675 12701 14676 12765
rect 14740 12701 14741 12765
rect 14675 12685 14741 12701
rect 14675 12621 14676 12685
rect 14740 12621 14741 12685
rect 14675 12467 14741 12621
rect 14801 12529 14861 13559
rect 14921 12467 14981 13499
rect 15041 12529 15101 13559
rect 15161 12467 15221 13499
rect 15281 13405 15347 13495
rect 15281 13341 15282 13405
rect 15346 13341 15347 13405
rect 15281 13325 15347 13341
rect 15281 13261 15282 13325
rect 15346 13261 15347 13325
rect 15281 13245 15347 13261
rect 15281 13181 15282 13245
rect 15346 13181 15347 13245
rect 15281 13165 15347 13181
rect 15281 13101 15282 13165
rect 15346 13101 15347 13165
rect 15281 13085 15347 13101
rect 15281 13021 15282 13085
rect 15346 13021 15347 13085
rect 15281 13005 15347 13021
rect 15281 12941 15282 13005
rect 15346 12941 15347 13005
rect 15281 12925 15347 12941
rect 15281 12861 15282 12925
rect 15346 12861 15347 12925
rect 15281 12845 15347 12861
rect 15281 12781 15282 12845
rect 15346 12781 15347 12845
rect 15281 12765 15347 12781
rect 15281 12701 15282 12765
rect 15346 12701 15347 12765
rect 15281 12685 15347 12701
rect 15281 12621 15282 12685
rect 15346 12621 15347 12685
rect 15281 12467 15347 12621
rect 15407 12467 15467 13499
rect 15527 12529 15587 13559
rect 15647 12467 15707 13499
rect 15767 12529 15827 13559
rect 15887 13405 15953 13495
rect 15887 13341 15888 13405
rect 15952 13341 15953 13405
rect 15887 13325 15953 13341
rect 15887 13261 15888 13325
rect 15952 13261 15953 13325
rect 15887 13245 15953 13261
rect 15887 13181 15888 13245
rect 15952 13181 15953 13245
rect 15887 13165 15953 13181
rect 15887 13101 15888 13165
rect 15952 13101 15953 13165
rect 15887 13085 15953 13101
rect 15887 13021 15888 13085
rect 15952 13021 15953 13085
rect 15887 13005 15953 13021
rect 15887 12941 15888 13005
rect 15952 12941 15953 13005
rect 15887 12925 15953 12941
rect 15887 12861 15888 12925
rect 15952 12861 15953 12925
rect 15887 12845 15953 12861
rect 15887 12781 15888 12845
rect 15952 12781 15953 12845
rect 15887 12765 15953 12781
rect 15887 12701 15888 12765
rect 15952 12701 15953 12765
rect 15887 12685 15953 12701
rect 15887 12621 15888 12685
rect 15952 12621 15953 12685
rect 15887 12467 15953 12621
rect 16013 12529 16073 13559
rect 16133 12467 16193 13499
rect 16253 12529 16313 13559
rect 16373 12467 16433 13499
rect 16493 13405 16559 13495
rect 16493 13341 16494 13405
rect 16558 13341 16559 13405
rect 16493 13325 16559 13341
rect 16493 13261 16494 13325
rect 16558 13261 16559 13325
rect 16493 13245 16559 13261
rect 16493 13181 16494 13245
rect 16558 13181 16559 13245
rect 16493 13165 16559 13181
rect 16493 13101 16494 13165
rect 16558 13101 16559 13165
rect 16493 13085 16559 13101
rect 16493 13021 16494 13085
rect 16558 13021 16559 13085
rect 16493 13005 16559 13021
rect 16493 12941 16494 13005
rect 16558 12941 16559 13005
rect 16493 12925 16559 12941
rect 16493 12861 16494 12925
rect 16558 12861 16559 12925
rect 16493 12845 16559 12861
rect 16493 12781 16494 12845
rect 16558 12781 16559 12845
rect 16493 12765 16559 12781
rect 16493 12701 16494 12765
rect 16558 12701 16559 12765
rect 16493 12685 16559 12701
rect 16493 12621 16494 12685
rect 16558 12621 16559 12685
rect 16493 12467 16559 12621
rect 16619 12467 16679 13499
rect 16739 12529 16799 13559
rect 16859 12467 16919 13499
rect 16979 12529 17039 13559
rect 17099 13405 17165 13495
rect 17099 13341 17100 13405
rect 17164 13341 17165 13405
rect 17099 13325 17165 13341
rect 17099 13261 17100 13325
rect 17164 13261 17165 13325
rect 17099 13245 17165 13261
rect 17099 13181 17100 13245
rect 17164 13181 17165 13245
rect 17099 13165 17165 13181
rect 17099 13101 17100 13165
rect 17164 13101 17165 13165
rect 17099 13085 17165 13101
rect 17099 13021 17100 13085
rect 17164 13021 17165 13085
rect 17099 13005 17165 13021
rect 17099 12941 17100 13005
rect 17164 12941 17165 13005
rect 17099 12925 17165 12941
rect 17099 12861 17100 12925
rect 17164 12861 17165 12925
rect 17099 12845 17165 12861
rect 17099 12781 17100 12845
rect 17164 12781 17165 12845
rect 17099 12765 17165 12781
rect 17099 12701 17100 12765
rect 17164 12701 17165 12765
rect 17099 12685 17165 12701
rect 17099 12621 17100 12685
rect 17164 12621 17165 12685
rect 17099 12467 17165 12621
rect 17225 12529 17285 13559
rect 17345 12467 17405 13499
rect 17465 12529 17525 13559
rect 17585 12467 17645 13499
rect 17705 13405 17771 13495
rect 17705 13341 17706 13405
rect 17770 13341 17771 13405
rect 17705 13325 17771 13341
rect 17705 13261 17706 13325
rect 17770 13261 17771 13325
rect 17705 13245 17771 13261
rect 17705 13181 17706 13245
rect 17770 13181 17771 13245
rect 17705 13165 17771 13181
rect 17705 13101 17706 13165
rect 17770 13101 17771 13165
rect 17705 13085 17771 13101
rect 17705 13021 17706 13085
rect 17770 13021 17771 13085
rect 17705 13005 17771 13021
rect 17705 12941 17706 13005
rect 17770 12941 17771 13005
rect 17705 12925 17771 12941
rect 17705 12861 17706 12925
rect 17770 12861 17771 12925
rect 17705 12845 17771 12861
rect 17705 12781 17706 12845
rect 17770 12781 17771 12845
rect 17705 12765 17771 12781
rect 17705 12701 17706 12765
rect 17770 12701 17771 12765
rect 17705 12685 17771 12701
rect 17705 12621 17706 12685
rect 17770 12621 17771 12685
rect 17705 12467 17771 12621
rect 17831 12467 17891 13499
rect 17951 12529 18011 13559
rect 18071 12467 18131 13499
rect 18191 12529 18251 13559
rect 18311 13405 18377 13495
rect 18311 13341 18312 13405
rect 18376 13341 18377 13405
rect 18311 13325 18377 13341
rect 18311 13261 18312 13325
rect 18376 13261 18377 13325
rect 18311 13245 18377 13261
rect 18311 13181 18312 13245
rect 18376 13181 18377 13245
rect 18311 13165 18377 13181
rect 18311 13101 18312 13165
rect 18376 13101 18377 13165
rect 18311 13085 18377 13101
rect 18311 13021 18312 13085
rect 18376 13021 18377 13085
rect 18311 13005 18377 13021
rect 18311 12941 18312 13005
rect 18376 12941 18377 13005
rect 18311 12925 18377 12941
rect 18311 12861 18312 12925
rect 18376 12861 18377 12925
rect 18311 12845 18377 12861
rect 18311 12781 18312 12845
rect 18376 12781 18377 12845
rect 18311 12765 18377 12781
rect 18311 12701 18312 12765
rect 18376 12701 18377 12765
rect 18311 12685 18377 12701
rect 18311 12621 18312 12685
rect 18376 12621 18377 12685
rect 18311 12467 18377 12621
rect 18437 12529 18497 13559
rect 18557 12467 18617 13499
rect 18677 12529 18737 13559
rect 18797 12467 18857 13499
rect 18917 13405 18983 13495
rect 18917 13341 18918 13405
rect 18982 13341 18983 13405
rect 18917 13325 18983 13341
rect 18917 13261 18918 13325
rect 18982 13261 18983 13325
rect 18917 13245 18983 13261
rect 18917 13181 18918 13245
rect 18982 13181 18983 13245
rect 18917 13165 18983 13181
rect 18917 13101 18918 13165
rect 18982 13101 18983 13165
rect 18917 13085 18983 13101
rect 18917 13021 18918 13085
rect 18982 13021 18983 13085
rect 18917 13005 18983 13021
rect 18917 12941 18918 13005
rect 18982 12941 18983 13005
rect 18917 12925 18983 12941
rect 18917 12861 18918 12925
rect 18982 12861 18983 12925
rect 18917 12845 18983 12861
rect 18917 12781 18918 12845
rect 18982 12781 18983 12845
rect 18917 12765 18983 12781
rect 18917 12701 18918 12765
rect 18982 12701 18983 12765
rect 18917 12685 18983 12701
rect 18917 12621 18918 12685
rect 18982 12621 18983 12685
rect 18917 12467 18983 12621
rect 19043 12467 19103 13499
rect 19163 12529 19223 13559
rect 19283 12467 19343 13499
rect 19403 12529 19463 13559
rect 19649 13506 19759 13559
rect 19823 13506 19967 13570
rect 19523 13405 19589 13495
rect 19523 13341 19524 13405
rect 19588 13341 19589 13405
rect 19523 13325 19589 13341
rect 19523 13261 19524 13325
rect 19588 13261 19589 13325
rect 19523 13245 19589 13261
rect 19523 13181 19524 13245
rect 19588 13181 19589 13245
rect 19523 13165 19589 13181
rect 19523 13101 19524 13165
rect 19588 13101 19589 13165
rect 19523 13085 19589 13101
rect 19523 13021 19524 13085
rect 19588 13021 19589 13085
rect 19523 13005 19589 13021
rect 19523 12941 19524 13005
rect 19588 12941 19589 13005
rect 19523 12925 19589 12941
rect 19523 12861 19524 12925
rect 19588 12861 19589 12925
rect 19523 12845 19589 12861
rect 19523 12781 19524 12845
rect 19588 12781 19589 12845
rect 19523 12765 19589 12781
rect 19523 12701 19524 12765
rect 19588 12701 19589 12765
rect 19523 12685 19589 12701
rect 19523 12621 19524 12685
rect 19588 12621 19589 12685
rect 19649 13426 19967 13506
rect 19649 13362 19764 13426
rect 19828 13362 19967 13426
rect 19649 13274 19967 13362
rect 19649 13210 19765 13274
rect 19829 13210 19967 13274
rect 19649 13104 19967 13210
rect 19649 13040 19765 13104
rect 19829 13040 19967 13104
rect 19649 12947 19967 13040
rect 19649 12883 19764 12947
rect 19828 12883 19967 12947
rect 20027 13573 20659 13626
rect 20027 13509 20236 13573
rect 20300 13568 20659 13573
rect 20723 13625 27155 13632
rect 20723 13622 21488 13625
rect 20723 13568 20756 13622
rect 20300 13559 20756 13568
rect 20300 13509 20445 13559
rect 20652 13558 20756 13559
rect 20820 13558 20836 13622
rect 20900 13558 20916 13622
rect 20980 13558 20996 13622
rect 21060 13558 21076 13622
rect 21140 13558 21156 13622
rect 21220 13561 21488 13622
rect 21552 13561 21568 13625
rect 21632 13561 21648 13625
rect 21712 13561 21728 13625
rect 21792 13561 21808 13625
rect 21872 13561 21888 13625
rect 21952 13561 22094 13625
rect 22158 13561 22174 13625
rect 22238 13561 22254 13625
rect 22318 13561 22334 13625
rect 22398 13561 22414 13625
rect 22478 13561 22494 13625
rect 22558 13561 22700 13625
rect 22764 13561 22780 13625
rect 22844 13561 22860 13625
rect 22924 13561 22940 13625
rect 23004 13561 23020 13625
rect 23084 13561 23100 13625
rect 23164 13561 23306 13625
rect 23370 13561 23386 13625
rect 23450 13561 23466 13625
rect 23530 13561 23546 13625
rect 23610 13561 23626 13625
rect 23690 13561 23706 13625
rect 23770 13561 23912 13625
rect 23976 13561 23992 13625
rect 24056 13561 24072 13625
rect 24136 13561 24152 13625
rect 24216 13561 24232 13625
rect 24296 13561 24312 13625
rect 24376 13561 24518 13625
rect 24582 13561 24598 13625
rect 24662 13561 24678 13625
rect 24742 13561 24758 13625
rect 24822 13561 24838 13625
rect 24902 13561 24918 13625
rect 24982 13561 25124 13625
rect 25188 13561 25204 13625
rect 25268 13561 25284 13625
rect 25348 13561 25364 13625
rect 25428 13561 25444 13625
rect 25508 13561 25524 13625
rect 25588 13561 25730 13625
rect 25794 13561 25810 13625
rect 25874 13561 25890 13625
rect 25954 13561 25970 13625
rect 26034 13561 26050 13625
rect 26114 13561 26130 13625
rect 26194 13570 26676 13625
rect 26194 13561 26468 13570
rect 21220 13559 26468 13561
rect 21220 13558 21325 13559
rect 20652 13557 21325 13558
rect 20652 13556 21324 13557
rect 20027 13401 20445 13509
rect 20027 13337 20225 13401
rect 20289 13337 20445 13401
rect 20027 13209 20445 13337
rect 20027 13145 20225 13209
rect 20289 13145 20445 13209
rect 20027 13027 20445 13145
rect 20027 12963 20042 13027
rect 20106 13026 20317 13027
rect 20106 12963 20173 13026
rect 20027 12962 20173 12963
rect 20237 12963 20317 13026
rect 20381 13021 20445 13027
rect 20652 13402 20718 13492
rect 20652 13338 20653 13402
rect 20717 13338 20718 13402
rect 20652 13322 20718 13338
rect 20652 13258 20653 13322
rect 20717 13258 20718 13322
rect 20652 13242 20718 13258
rect 20652 13178 20653 13242
rect 20717 13178 20718 13242
rect 20652 13162 20718 13178
rect 20652 13098 20653 13162
rect 20717 13098 20718 13162
rect 20652 13082 20718 13098
rect 20381 12963 20444 13021
rect 20237 12962 20444 12963
rect 20027 12944 20444 12962
rect 20652 13018 20653 13082
rect 20717 13018 20718 13082
rect 20652 13002 20718 13018
rect 19649 12705 19967 12883
rect 19649 12641 19682 12705
rect 19746 12641 19967 12705
rect 19649 12629 19967 12641
rect 19523 12467 19589 12621
rect 14675 12465 19589 12467
rect 14675 12401 14779 12465
rect 14843 12401 14859 12465
rect 14923 12401 14939 12465
rect 15003 12401 15019 12465
rect 15083 12401 15099 12465
rect 15163 12401 15179 12465
rect 15243 12401 15385 12465
rect 15449 12401 15465 12465
rect 15529 12401 15545 12465
rect 15609 12401 15625 12465
rect 15689 12401 15705 12465
rect 15769 12401 15785 12465
rect 15849 12401 15991 12465
rect 16055 12401 16071 12465
rect 16135 12401 16151 12465
rect 16215 12401 16231 12465
rect 16295 12401 16311 12465
rect 16375 12401 16391 12465
rect 16455 12401 16597 12465
rect 16661 12401 16677 12465
rect 16741 12401 16757 12465
rect 16821 12401 16837 12465
rect 16901 12401 16917 12465
rect 16981 12401 16997 12465
rect 17061 12401 17203 12465
rect 17267 12401 17283 12465
rect 17347 12401 17363 12465
rect 17427 12401 17443 12465
rect 17507 12401 17523 12465
rect 17587 12401 17603 12465
rect 17667 12401 17809 12465
rect 17873 12401 17889 12465
rect 17953 12401 17969 12465
rect 18033 12401 18049 12465
rect 18113 12401 18129 12465
rect 18193 12401 18209 12465
rect 18273 12401 18415 12465
rect 18479 12401 18495 12465
rect 18559 12401 18575 12465
rect 18639 12401 18655 12465
rect 18719 12401 18735 12465
rect 18799 12401 18815 12465
rect 18879 12401 19021 12465
rect 19085 12401 19101 12465
rect 19165 12401 19181 12465
rect 19245 12401 19261 12465
rect 19325 12401 19341 12465
rect 19405 12401 19421 12465
rect 19485 12401 19589 12465
rect 14675 12399 19589 12401
rect 19649 12444 19847 12454
rect 13943 12396 14615 12398
rect 19649 12380 19770 12444
rect 19834 12380 19847 12444
rect 19649 12370 19847 12380
rect 10646 11888 13067 12091
rect 10646 11885 11113 11888
rect 10646 11821 10913 11885
rect 10977 11824 11113 11885
rect 11177 11886 13067 11888
rect 11177 11824 11349 11886
rect 10977 11822 11349 11824
rect 11413 11882 13067 11886
rect 11413 11881 12360 11882
rect 11413 11880 11983 11881
rect 11413 11822 11782 11880
rect 10977 11821 11782 11822
rect 10646 11816 11782 11821
rect 11846 11817 11983 11880
rect 12047 11879 12360 11881
rect 12047 11817 12169 11879
rect 11846 11816 12169 11817
rect 10646 11815 12169 11816
rect 12233 11818 12360 11879
rect 12424 11881 13067 11882
rect 12424 11818 12573 11881
rect 12233 11817 12573 11818
rect 12637 11817 13067 11881
rect 12233 11815 13067 11817
rect 10646 11599 13067 11815
rect 13215 11601 13722 12172
rect 8761 11525 9342 11573
rect 8761 11504 9194 11525
rect 8761 11440 8791 11504
rect 8855 11461 9194 11504
rect 9258 11461 9342 11525
rect 8855 11440 9342 11461
rect 8761 11398 9342 11440
rect 13215 11537 13318 11601
rect 13383 11537 13722 11601
rect 3406 10583 4078 10584
rect 4138 10583 6628 10584
rect 6688 10583 7966 10584
rect 8028 10583 8700 10584
rect 8761 10583 9079 11398
rect 13215 11322 13722 11537
rect 11374 11301 13722 11322
rect 2458 10582 9079 10583
rect 2458 10579 3590 10582
rect 2458 10515 3048 10579
rect 3112 10518 3590 10579
rect 3654 10518 3670 10582
rect 3734 10518 3750 10582
rect 3814 10518 3830 10582
rect 3894 10518 4322 10582
rect 4386 10518 4402 10582
rect 4466 10518 4482 10582
rect 4546 10518 4562 10582
rect 4626 10518 4928 10582
rect 4992 10518 5008 10582
rect 5072 10518 5088 10582
rect 5152 10518 5168 10582
rect 5232 10518 5534 10582
rect 5598 10518 5614 10582
rect 5678 10518 5694 10582
rect 5758 10518 5774 10582
rect 5838 10518 6140 10582
rect 6204 10518 6220 10582
rect 6284 10518 6300 10582
rect 6364 10518 6380 10582
rect 6444 10518 6872 10582
rect 6936 10518 6952 10582
rect 7016 10518 7032 10582
rect 7096 10518 7112 10582
rect 7176 10518 7478 10582
rect 7542 10518 7558 10582
rect 7622 10518 7638 10582
rect 7702 10518 7718 10582
rect 7782 10518 8212 10582
rect 8276 10518 8292 10582
rect 8356 10518 8372 10582
rect 8436 10518 8452 10582
rect 8516 10518 9079 10582
rect 3112 10515 9079 10518
rect 2458 10505 9079 10515
rect 10878 11263 13722 11301
rect 10878 11199 10929 11263
rect 10993 11260 13722 11263
rect 10993 11199 11117 11260
rect 10878 11196 11117 11199
rect 11181 11258 13722 11260
rect 11181 11196 11314 11258
rect 10878 11194 11314 11196
rect 11378 11194 13722 11258
rect 10878 11058 13722 11194
rect 14294 12217 14966 12219
rect 14294 12153 14398 12217
rect 14462 12153 14478 12217
rect 14542 12153 14558 12217
rect 14622 12153 14638 12217
rect 14702 12153 14718 12217
rect 14782 12153 14798 12217
rect 14862 12153 14966 12217
rect 14294 12151 14966 12153
rect 14294 11997 14360 12151
rect 14294 11933 14295 11997
rect 14359 11933 14360 11997
rect 14294 11917 14360 11933
rect 14294 11853 14295 11917
rect 14359 11853 14360 11917
rect 14294 11837 14360 11853
rect 14294 11773 14295 11837
rect 14359 11773 14360 11837
rect 14294 11757 14360 11773
rect 14294 11693 14295 11757
rect 14359 11693 14360 11757
rect 14294 11677 14360 11693
rect 14294 11613 14295 11677
rect 14359 11613 14360 11677
rect 14294 11597 14360 11613
rect 14294 11533 14295 11597
rect 14359 11533 14360 11597
rect 14294 11517 14360 11533
rect 14294 11453 14295 11517
rect 14359 11453 14360 11517
rect 14294 11437 14360 11453
rect 14294 11373 14295 11437
rect 14359 11373 14360 11437
rect 14294 11357 14360 11373
rect 14294 11293 14295 11357
rect 14359 11293 14360 11357
rect 14294 11277 14360 11293
rect 14294 11213 14295 11277
rect 14359 11213 14360 11277
rect 14294 11123 14360 11213
rect 13906 11058 14031 11064
rect 14420 11059 14480 12089
rect 14540 11119 14600 12151
rect 14660 11059 14720 12089
rect 14780 11119 14840 12151
rect 14900 11997 14966 12151
rect 14900 11933 14901 11997
rect 14965 11933 14966 11997
rect 14900 11917 14966 11933
rect 14900 11853 14901 11917
rect 14965 11853 14966 11917
rect 14900 11837 14966 11853
rect 14900 11773 14901 11837
rect 14965 11773 14966 11837
rect 14900 11757 14966 11773
rect 14900 11693 14901 11757
rect 14965 11693 14966 11757
rect 14900 11677 14966 11693
rect 14900 11613 14901 11677
rect 14965 11613 14966 11677
rect 14900 11597 14966 11613
rect 14900 11533 14901 11597
rect 14965 11533 14966 11597
rect 14900 11517 14966 11533
rect 14900 11453 14901 11517
rect 14965 11453 14966 11517
rect 14900 11437 14966 11453
rect 14900 11373 14901 11437
rect 14965 11373 14966 11437
rect 14900 11357 14966 11373
rect 14900 11293 14901 11357
rect 14965 11293 14966 11357
rect 14900 11277 14966 11293
rect 14900 11213 14901 11277
rect 14965 11213 14966 11277
rect 14900 11123 14966 11213
rect 15026 12217 17516 12219
rect 15026 12153 15130 12217
rect 15194 12153 15210 12217
rect 15274 12153 15290 12217
rect 15354 12153 15370 12217
rect 15434 12153 15450 12217
rect 15514 12153 15530 12217
rect 15594 12153 15736 12217
rect 15800 12153 15816 12217
rect 15880 12153 15896 12217
rect 15960 12153 15976 12217
rect 16040 12153 16056 12217
rect 16120 12153 16136 12217
rect 16200 12153 16342 12217
rect 16406 12153 16422 12217
rect 16486 12153 16502 12217
rect 16566 12153 16582 12217
rect 16646 12153 16662 12217
rect 16726 12153 16742 12217
rect 16806 12153 16948 12217
rect 17012 12153 17028 12217
rect 17092 12153 17108 12217
rect 17172 12153 17188 12217
rect 17252 12153 17268 12217
rect 17332 12153 17348 12217
rect 17412 12153 17516 12217
rect 15026 12151 17516 12153
rect 15026 11997 15092 12151
rect 15026 11933 15027 11997
rect 15091 11933 15092 11997
rect 15026 11917 15092 11933
rect 15026 11853 15027 11917
rect 15091 11853 15092 11917
rect 15026 11837 15092 11853
rect 15026 11773 15027 11837
rect 15091 11773 15092 11837
rect 15026 11757 15092 11773
rect 15026 11693 15027 11757
rect 15091 11693 15092 11757
rect 15026 11677 15092 11693
rect 15026 11613 15027 11677
rect 15091 11613 15092 11677
rect 15026 11597 15092 11613
rect 15026 11533 15027 11597
rect 15091 11533 15092 11597
rect 15026 11517 15092 11533
rect 15026 11453 15027 11517
rect 15091 11453 15092 11517
rect 15026 11437 15092 11453
rect 15026 11373 15027 11437
rect 15091 11373 15092 11437
rect 15026 11357 15092 11373
rect 15026 11293 15027 11357
rect 15091 11293 15092 11357
rect 15026 11277 15092 11293
rect 15026 11213 15027 11277
rect 15091 11213 15092 11277
rect 15026 11123 15092 11213
rect 15152 11059 15212 12089
rect 15272 11119 15332 12151
rect 15392 11059 15452 12089
rect 15512 11119 15572 12151
rect 15632 11997 15698 12151
rect 15632 11933 15633 11997
rect 15697 11933 15698 11997
rect 15632 11917 15698 11933
rect 15632 11853 15633 11917
rect 15697 11853 15698 11917
rect 15632 11837 15698 11853
rect 15632 11773 15633 11837
rect 15697 11773 15698 11837
rect 15632 11757 15698 11773
rect 15632 11693 15633 11757
rect 15697 11693 15698 11757
rect 15632 11677 15698 11693
rect 15632 11613 15633 11677
rect 15697 11613 15698 11677
rect 15632 11597 15698 11613
rect 15632 11533 15633 11597
rect 15697 11533 15698 11597
rect 15632 11517 15698 11533
rect 15632 11453 15633 11517
rect 15697 11453 15698 11517
rect 15632 11437 15698 11453
rect 15632 11373 15633 11437
rect 15697 11373 15698 11437
rect 15632 11357 15698 11373
rect 15632 11293 15633 11357
rect 15697 11293 15698 11357
rect 15632 11277 15698 11293
rect 15632 11213 15633 11277
rect 15697 11213 15698 11277
rect 15632 11123 15698 11213
rect 15758 11119 15818 12151
rect 15878 11059 15938 12089
rect 15998 11119 16058 12151
rect 16118 11059 16178 12089
rect 16238 11997 16304 12151
rect 16238 11933 16239 11997
rect 16303 11933 16304 11997
rect 16238 11917 16304 11933
rect 16238 11853 16239 11917
rect 16303 11853 16304 11917
rect 16238 11837 16304 11853
rect 16238 11773 16239 11837
rect 16303 11773 16304 11837
rect 16238 11757 16304 11773
rect 16238 11693 16239 11757
rect 16303 11693 16304 11757
rect 16238 11677 16304 11693
rect 16238 11613 16239 11677
rect 16303 11613 16304 11677
rect 16238 11597 16304 11613
rect 16238 11533 16239 11597
rect 16303 11533 16304 11597
rect 16238 11517 16304 11533
rect 16238 11453 16239 11517
rect 16303 11453 16304 11517
rect 16238 11437 16304 11453
rect 16238 11373 16239 11437
rect 16303 11373 16304 11437
rect 16238 11357 16304 11373
rect 16238 11293 16239 11357
rect 16303 11293 16304 11357
rect 16238 11277 16304 11293
rect 16238 11213 16239 11277
rect 16303 11213 16304 11277
rect 16238 11123 16304 11213
rect 16364 11059 16424 12089
rect 16484 11119 16544 12151
rect 16604 11059 16664 12089
rect 16724 11119 16784 12151
rect 16844 11997 16910 12151
rect 16844 11933 16845 11997
rect 16909 11933 16910 11997
rect 16844 11917 16910 11933
rect 16844 11853 16845 11917
rect 16909 11853 16910 11917
rect 16844 11837 16910 11853
rect 16844 11773 16845 11837
rect 16909 11773 16910 11837
rect 16844 11757 16910 11773
rect 16844 11693 16845 11757
rect 16909 11693 16910 11757
rect 16844 11677 16910 11693
rect 16844 11613 16845 11677
rect 16909 11613 16910 11677
rect 16844 11597 16910 11613
rect 16844 11533 16845 11597
rect 16909 11533 16910 11597
rect 16844 11517 16910 11533
rect 16844 11453 16845 11517
rect 16909 11453 16910 11517
rect 16844 11437 16910 11453
rect 16844 11373 16845 11437
rect 16909 11373 16910 11437
rect 16844 11357 16910 11373
rect 16844 11293 16845 11357
rect 16909 11293 16910 11357
rect 16844 11277 16910 11293
rect 16844 11213 16845 11277
rect 16909 11213 16910 11277
rect 16844 11123 16910 11213
rect 16970 11119 17030 12151
rect 17090 11059 17150 12089
rect 17210 11119 17270 12151
rect 17330 11059 17390 12089
rect 17450 11997 17516 12151
rect 17450 11933 17451 11997
rect 17515 11933 17516 11997
rect 17450 11917 17516 11933
rect 17450 11853 17451 11917
rect 17515 11853 17516 11917
rect 17450 11837 17516 11853
rect 17450 11773 17451 11837
rect 17515 11773 17516 11837
rect 17450 11757 17516 11773
rect 17450 11693 17451 11757
rect 17515 11693 17516 11757
rect 17450 11677 17516 11693
rect 17450 11613 17451 11677
rect 17515 11613 17516 11677
rect 17450 11597 17516 11613
rect 17450 11533 17451 11597
rect 17515 11533 17516 11597
rect 17450 11517 17516 11533
rect 17450 11453 17451 11517
rect 17515 11453 17516 11517
rect 17450 11437 17516 11453
rect 17450 11373 17451 11437
rect 17515 11373 17516 11437
rect 17450 11357 17516 11373
rect 17450 11293 17451 11357
rect 17515 11293 17516 11357
rect 17450 11277 17516 11293
rect 17450 11213 17451 11277
rect 17515 11213 17516 11277
rect 17450 11123 17516 11213
rect 17576 12217 18854 12219
rect 17576 12153 17680 12217
rect 17744 12153 17760 12217
rect 17824 12153 17840 12217
rect 17904 12153 17920 12217
rect 17984 12153 18000 12217
rect 18064 12153 18080 12217
rect 18144 12153 18286 12217
rect 18350 12153 18366 12217
rect 18430 12153 18446 12217
rect 18510 12153 18526 12217
rect 18590 12153 18606 12217
rect 18670 12153 18686 12217
rect 18750 12153 18854 12217
rect 17576 12151 18854 12153
rect 17576 11997 17642 12151
rect 17576 11933 17577 11997
rect 17641 11933 17642 11997
rect 17576 11917 17642 11933
rect 17576 11853 17577 11917
rect 17641 11853 17642 11917
rect 17576 11837 17642 11853
rect 17576 11773 17577 11837
rect 17641 11773 17642 11837
rect 17576 11757 17642 11773
rect 17576 11693 17577 11757
rect 17641 11693 17642 11757
rect 17576 11677 17642 11693
rect 17576 11613 17577 11677
rect 17641 11613 17642 11677
rect 17576 11597 17642 11613
rect 17576 11533 17577 11597
rect 17641 11533 17642 11597
rect 17576 11517 17642 11533
rect 17576 11453 17577 11517
rect 17641 11453 17642 11517
rect 17576 11437 17642 11453
rect 17576 11373 17577 11437
rect 17641 11373 17642 11437
rect 17576 11357 17642 11373
rect 17576 11293 17577 11357
rect 17641 11293 17642 11357
rect 17576 11277 17642 11293
rect 17576 11213 17577 11277
rect 17641 11213 17642 11277
rect 17576 11123 17642 11213
rect 17702 11059 17762 12089
rect 17822 11119 17882 12151
rect 17942 11059 18002 12089
rect 18062 11119 18122 12151
rect 18182 11997 18248 12151
rect 18182 11933 18183 11997
rect 18247 11933 18248 11997
rect 18182 11917 18248 11933
rect 18182 11853 18183 11917
rect 18247 11853 18248 11917
rect 18182 11837 18248 11853
rect 18182 11773 18183 11837
rect 18247 11773 18248 11837
rect 18182 11757 18248 11773
rect 18182 11693 18183 11757
rect 18247 11693 18248 11757
rect 18182 11677 18248 11693
rect 18182 11613 18183 11677
rect 18247 11613 18248 11677
rect 18182 11597 18248 11613
rect 18182 11533 18183 11597
rect 18247 11533 18248 11597
rect 18182 11517 18248 11533
rect 18182 11453 18183 11517
rect 18247 11453 18248 11517
rect 18182 11437 18248 11453
rect 18182 11373 18183 11437
rect 18247 11373 18248 11437
rect 18182 11357 18248 11373
rect 18182 11293 18183 11357
rect 18247 11293 18248 11357
rect 18182 11277 18248 11293
rect 18182 11213 18183 11277
rect 18247 11213 18248 11277
rect 18182 11123 18248 11213
rect 18308 11119 18368 12151
rect 18428 11059 18488 12089
rect 18548 11119 18608 12151
rect 18668 11059 18728 12089
rect 18788 11997 18854 12151
rect 18788 11933 18789 11997
rect 18853 11933 18854 11997
rect 18788 11917 18854 11933
rect 18788 11853 18789 11917
rect 18853 11853 18854 11917
rect 18788 11837 18854 11853
rect 18788 11773 18789 11837
rect 18853 11773 18854 11837
rect 18788 11757 18854 11773
rect 18788 11693 18789 11757
rect 18853 11693 18854 11757
rect 18788 11677 18854 11693
rect 18788 11613 18789 11677
rect 18853 11613 18854 11677
rect 18788 11597 18854 11613
rect 18788 11533 18789 11597
rect 18853 11533 18854 11597
rect 18788 11517 18854 11533
rect 18788 11453 18789 11517
rect 18853 11453 18854 11517
rect 18788 11437 18854 11453
rect 18788 11373 18789 11437
rect 18853 11373 18854 11437
rect 18788 11357 18854 11373
rect 18788 11293 18789 11357
rect 18853 11293 18854 11357
rect 18788 11277 18854 11293
rect 18788 11213 18789 11277
rect 18853 11213 18854 11277
rect 18788 11123 18854 11213
rect 18916 12217 19588 12219
rect 18916 12153 19020 12217
rect 19084 12153 19100 12217
rect 19164 12153 19180 12217
rect 19244 12153 19260 12217
rect 19324 12153 19340 12217
rect 19404 12153 19420 12217
rect 19484 12153 19588 12217
rect 18916 12151 19588 12153
rect 18916 11997 18982 12151
rect 18916 11933 18917 11997
rect 18981 11933 18982 11997
rect 18916 11917 18982 11933
rect 18916 11853 18917 11917
rect 18981 11853 18982 11917
rect 18916 11837 18982 11853
rect 18916 11773 18917 11837
rect 18981 11773 18982 11837
rect 18916 11757 18982 11773
rect 18916 11693 18917 11757
rect 18981 11693 18982 11757
rect 18916 11677 18982 11693
rect 18916 11613 18917 11677
rect 18981 11613 18982 11677
rect 18916 11597 18982 11613
rect 18916 11533 18917 11597
rect 18981 11533 18982 11597
rect 18916 11517 18982 11533
rect 18916 11453 18917 11517
rect 18981 11453 18982 11517
rect 18916 11437 18982 11453
rect 18916 11373 18917 11437
rect 18981 11373 18982 11437
rect 18916 11357 18982 11373
rect 18916 11293 18917 11357
rect 18981 11293 18982 11357
rect 18916 11277 18982 11293
rect 18916 11213 18917 11277
rect 18981 11213 18982 11277
rect 18916 11123 18982 11213
rect 19042 11119 19102 12151
rect 19162 11059 19222 12089
rect 19282 11119 19342 12151
rect 19402 11059 19462 12089
rect 19522 11997 19588 12151
rect 19522 11933 19523 11997
rect 19587 11933 19588 11997
rect 19522 11917 19588 11933
rect 19522 11853 19523 11917
rect 19587 11853 19588 11917
rect 19522 11837 19588 11853
rect 19522 11773 19523 11837
rect 19587 11773 19588 11837
rect 19522 11757 19588 11773
rect 19522 11693 19523 11757
rect 19587 11693 19588 11757
rect 19522 11677 19588 11693
rect 19522 11613 19523 11677
rect 19587 11613 19588 11677
rect 19522 11597 19588 11613
rect 19522 11533 19523 11597
rect 19587 11533 19588 11597
rect 19522 11517 19588 11533
rect 19522 11453 19523 11517
rect 19587 11453 19588 11517
rect 19522 11437 19588 11453
rect 19522 11373 19523 11437
rect 19587 11373 19588 11437
rect 19522 11357 19588 11373
rect 19522 11293 19523 11357
rect 19587 11293 19588 11357
rect 19522 11277 19588 11293
rect 19522 11213 19523 11277
rect 19587 11213 19588 11277
rect 19522 11123 19588 11213
rect 19649 11989 19709 12370
rect 19907 12251 19967 12629
rect 20652 12938 20653 13002
rect 20717 12938 20718 13002
rect 20652 12922 20718 12938
rect 20652 12858 20653 12922
rect 20717 12858 20718 12922
rect 20652 12842 20718 12858
rect 20652 12778 20653 12842
rect 20717 12778 20718 12842
rect 20652 12762 20718 12778
rect 20652 12698 20653 12762
rect 20717 12698 20718 12762
rect 20652 12682 20718 12698
rect 20652 12618 20653 12682
rect 20717 12618 20718 12682
rect 20053 12481 20430 12496
rect 20053 12417 20060 12481
rect 20124 12417 20180 12481
rect 20244 12417 20323 12481
rect 20387 12417 20430 12481
rect 20652 12464 20718 12618
rect 20778 12526 20838 13556
rect 20898 12464 20958 13496
rect 21018 12526 21078 13556
rect 21138 12464 21198 13496
rect 21258 13402 21324 13492
rect 21258 13338 21259 13402
rect 21323 13338 21324 13402
rect 21258 13322 21324 13338
rect 21258 13258 21259 13322
rect 21323 13258 21324 13322
rect 21258 13242 21324 13258
rect 21258 13178 21259 13242
rect 21323 13178 21324 13242
rect 21258 13162 21324 13178
rect 21258 13098 21259 13162
rect 21323 13098 21324 13162
rect 21258 13082 21324 13098
rect 21258 13018 21259 13082
rect 21323 13018 21324 13082
rect 21258 13002 21324 13018
rect 21258 12938 21259 13002
rect 21323 12938 21324 13002
rect 21258 12922 21324 12938
rect 21258 12858 21259 12922
rect 21323 12858 21324 12922
rect 21258 12842 21324 12858
rect 21258 12778 21259 12842
rect 21323 12778 21324 12842
rect 21258 12762 21324 12778
rect 21258 12698 21259 12762
rect 21323 12698 21324 12762
rect 21258 12682 21324 12698
rect 21258 12618 21259 12682
rect 21323 12618 21324 12682
rect 21258 12464 21324 12618
rect 20652 12462 21324 12464
rect 19769 12241 19967 12251
rect 19769 12177 19770 12241
rect 19834 12177 19967 12241
rect 19769 12167 19967 12177
rect 19649 11979 19967 11989
rect 19649 11915 19679 11979
rect 19743 11915 19967 11979
rect 14294 11058 14966 11059
rect 15026 11058 17516 11059
rect 17576 11058 18854 11059
rect 18916 11058 19588 11059
rect 19649 11058 19967 11915
rect 10878 11057 19967 11058
rect 10878 11054 14478 11057
rect 10878 10990 13936 11054
rect 14000 10993 14478 11054
rect 14542 10993 14558 11057
rect 14622 10993 14638 11057
rect 14702 10993 14718 11057
rect 14782 10993 15210 11057
rect 15274 10993 15290 11057
rect 15354 10993 15370 11057
rect 15434 10993 15450 11057
rect 15514 10993 15816 11057
rect 15880 10993 15896 11057
rect 15960 10993 15976 11057
rect 16040 10993 16056 11057
rect 16120 10993 16422 11057
rect 16486 10993 16502 11057
rect 16566 10993 16582 11057
rect 16646 10993 16662 11057
rect 16726 10993 17028 11057
rect 17092 10993 17108 11057
rect 17172 10993 17188 11057
rect 17252 10993 17268 11057
rect 17332 10993 17760 11057
rect 17824 10993 17840 11057
rect 17904 10993 17920 11057
rect 17984 10993 18000 11057
rect 18064 10993 18366 11057
rect 18430 10993 18446 11057
rect 18510 10993 18526 11057
rect 18590 10993 18606 11057
rect 18670 10993 19100 11057
rect 19164 10993 19180 11057
rect 19244 10993 19260 11057
rect 19324 10993 19340 11057
rect 19404 11044 19967 11057
rect 20055 11058 20431 12417
rect 20652 12398 20756 12462
rect 20820 12398 20836 12462
rect 20900 12398 20916 12462
rect 20980 12398 20996 12462
rect 21060 12398 21076 12462
rect 21140 12398 21156 12462
rect 21220 12398 21324 12462
rect 21384 13405 21450 13495
rect 21384 13341 21385 13405
rect 21449 13341 21450 13405
rect 21384 13325 21450 13341
rect 21384 13261 21385 13325
rect 21449 13261 21450 13325
rect 21384 13245 21450 13261
rect 21384 13181 21385 13245
rect 21449 13181 21450 13245
rect 21384 13165 21450 13181
rect 21384 13101 21385 13165
rect 21449 13101 21450 13165
rect 21384 13085 21450 13101
rect 21384 13021 21385 13085
rect 21449 13021 21450 13085
rect 21384 13005 21450 13021
rect 21384 12941 21385 13005
rect 21449 12941 21450 13005
rect 21384 12925 21450 12941
rect 21384 12861 21385 12925
rect 21449 12861 21450 12925
rect 21384 12845 21450 12861
rect 21384 12781 21385 12845
rect 21449 12781 21450 12845
rect 21384 12765 21450 12781
rect 21384 12701 21385 12765
rect 21449 12701 21450 12765
rect 21384 12685 21450 12701
rect 21384 12621 21385 12685
rect 21449 12621 21450 12685
rect 21384 12467 21450 12621
rect 21510 12529 21570 13559
rect 21630 12467 21690 13499
rect 21750 12529 21810 13559
rect 21870 12467 21930 13499
rect 21990 13405 22056 13495
rect 21990 13341 21991 13405
rect 22055 13341 22056 13405
rect 21990 13325 22056 13341
rect 21990 13261 21991 13325
rect 22055 13261 22056 13325
rect 21990 13245 22056 13261
rect 21990 13181 21991 13245
rect 22055 13181 22056 13245
rect 21990 13165 22056 13181
rect 21990 13101 21991 13165
rect 22055 13101 22056 13165
rect 21990 13085 22056 13101
rect 21990 13021 21991 13085
rect 22055 13021 22056 13085
rect 21990 13005 22056 13021
rect 21990 12941 21991 13005
rect 22055 12941 22056 13005
rect 21990 12925 22056 12941
rect 21990 12861 21991 12925
rect 22055 12861 22056 12925
rect 21990 12845 22056 12861
rect 21990 12781 21991 12845
rect 22055 12781 22056 12845
rect 21990 12765 22056 12781
rect 21990 12701 21991 12765
rect 22055 12701 22056 12765
rect 21990 12685 22056 12701
rect 21990 12621 21991 12685
rect 22055 12621 22056 12685
rect 21990 12467 22056 12621
rect 22116 12467 22176 13499
rect 22236 12529 22296 13559
rect 22356 12467 22416 13499
rect 22476 12529 22536 13559
rect 22596 13405 22662 13495
rect 22596 13341 22597 13405
rect 22661 13341 22662 13405
rect 22596 13325 22662 13341
rect 22596 13261 22597 13325
rect 22661 13261 22662 13325
rect 22596 13245 22662 13261
rect 22596 13181 22597 13245
rect 22661 13181 22662 13245
rect 22596 13165 22662 13181
rect 22596 13101 22597 13165
rect 22661 13101 22662 13165
rect 22596 13085 22662 13101
rect 22596 13021 22597 13085
rect 22661 13021 22662 13085
rect 22596 13005 22662 13021
rect 22596 12941 22597 13005
rect 22661 12941 22662 13005
rect 22596 12925 22662 12941
rect 22596 12861 22597 12925
rect 22661 12861 22662 12925
rect 22596 12845 22662 12861
rect 22596 12781 22597 12845
rect 22661 12781 22662 12845
rect 22596 12765 22662 12781
rect 22596 12701 22597 12765
rect 22661 12701 22662 12765
rect 22596 12685 22662 12701
rect 22596 12621 22597 12685
rect 22661 12621 22662 12685
rect 22596 12467 22662 12621
rect 22722 12529 22782 13559
rect 22842 12467 22902 13499
rect 22962 12529 23022 13559
rect 23082 12467 23142 13499
rect 23202 13405 23268 13495
rect 23202 13341 23203 13405
rect 23267 13341 23268 13405
rect 23202 13325 23268 13341
rect 23202 13261 23203 13325
rect 23267 13261 23268 13325
rect 23202 13245 23268 13261
rect 23202 13181 23203 13245
rect 23267 13181 23268 13245
rect 23202 13165 23268 13181
rect 23202 13101 23203 13165
rect 23267 13101 23268 13165
rect 23202 13085 23268 13101
rect 23202 13021 23203 13085
rect 23267 13021 23268 13085
rect 23202 13005 23268 13021
rect 23202 12941 23203 13005
rect 23267 12941 23268 13005
rect 23202 12925 23268 12941
rect 23202 12861 23203 12925
rect 23267 12861 23268 12925
rect 23202 12845 23268 12861
rect 23202 12781 23203 12845
rect 23267 12781 23268 12845
rect 23202 12765 23268 12781
rect 23202 12701 23203 12765
rect 23267 12701 23268 12765
rect 23202 12685 23268 12701
rect 23202 12621 23203 12685
rect 23267 12621 23268 12685
rect 23202 12467 23268 12621
rect 23328 12467 23388 13499
rect 23448 12529 23508 13559
rect 23568 12467 23628 13499
rect 23688 12529 23748 13559
rect 23808 13405 23874 13495
rect 23808 13341 23809 13405
rect 23873 13341 23874 13405
rect 23808 13325 23874 13341
rect 23808 13261 23809 13325
rect 23873 13261 23874 13325
rect 23808 13245 23874 13261
rect 23808 13181 23809 13245
rect 23873 13181 23874 13245
rect 23808 13165 23874 13181
rect 23808 13101 23809 13165
rect 23873 13101 23874 13165
rect 23808 13085 23874 13101
rect 23808 13021 23809 13085
rect 23873 13021 23874 13085
rect 23808 13005 23874 13021
rect 23808 12941 23809 13005
rect 23873 12941 23874 13005
rect 23808 12925 23874 12941
rect 23808 12861 23809 12925
rect 23873 12861 23874 12925
rect 23808 12845 23874 12861
rect 23808 12781 23809 12845
rect 23873 12781 23874 12845
rect 23808 12765 23874 12781
rect 23808 12701 23809 12765
rect 23873 12701 23874 12765
rect 23808 12685 23874 12701
rect 23808 12621 23809 12685
rect 23873 12621 23874 12685
rect 23808 12467 23874 12621
rect 23934 12529 23994 13559
rect 24054 12467 24114 13499
rect 24174 12529 24234 13559
rect 24294 12467 24354 13499
rect 24414 13405 24480 13495
rect 24414 13341 24415 13405
rect 24479 13341 24480 13405
rect 24414 13325 24480 13341
rect 24414 13261 24415 13325
rect 24479 13261 24480 13325
rect 24414 13245 24480 13261
rect 24414 13181 24415 13245
rect 24479 13181 24480 13245
rect 24414 13165 24480 13181
rect 24414 13101 24415 13165
rect 24479 13101 24480 13165
rect 24414 13085 24480 13101
rect 24414 13021 24415 13085
rect 24479 13021 24480 13085
rect 24414 13005 24480 13021
rect 24414 12941 24415 13005
rect 24479 12941 24480 13005
rect 24414 12925 24480 12941
rect 24414 12861 24415 12925
rect 24479 12861 24480 12925
rect 24414 12845 24480 12861
rect 24414 12781 24415 12845
rect 24479 12781 24480 12845
rect 24414 12765 24480 12781
rect 24414 12701 24415 12765
rect 24479 12701 24480 12765
rect 24414 12685 24480 12701
rect 24414 12621 24415 12685
rect 24479 12621 24480 12685
rect 24414 12467 24480 12621
rect 24540 12467 24600 13499
rect 24660 12529 24720 13559
rect 24780 12467 24840 13499
rect 24900 12529 24960 13559
rect 25020 13405 25086 13495
rect 25020 13341 25021 13405
rect 25085 13341 25086 13405
rect 25020 13325 25086 13341
rect 25020 13261 25021 13325
rect 25085 13261 25086 13325
rect 25020 13245 25086 13261
rect 25020 13181 25021 13245
rect 25085 13181 25086 13245
rect 25020 13165 25086 13181
rect 25020 13101 25021 13165
rect 25085 13101 25086 13165
rect 25020 13085 25086 13101
rect 25020 13021 25021 13085
rect 25085 13021 25086 13085
rect 25020 13005 25086 13021
rect 25020 12941 25021 13005
rect 25085 12941 25086 13005
rect 25020 12925 25086 12941
rect 25020 12861 25021 12925
rect 25085 12861 25086 12925
rect 25020 12845 25086 12861
rect 25020 12781 25021 12845
rect 25085 12781 25086 12845
rect 25020 12765 25086 12781
rect 25020 12701 25021 12765
rect 25085 12701 25086 12765
rect 25020 12685 25086 12701
rect 25020 12621 25021 12685
rect 25085 12621 25086 12685
rect 25020 12467 25086 12621
rect 25146 12529 25206 13559
rect 25266 12467 25326 13499
rect 25386 12529 25446 13559
rect 25506 12467 25566 13499
rect 25626 13405 25692 13495
rect 25626 13341 25627 13405
rect 25691 13341 25692 13405
rect 25626 13325 25692 13341
rect 25626 13261 25627 13325
rect 25691 13261 25692 13325
rect 25626 13245 25692 13261
rect 25626 13181 25627 13245
rect 25691 13181 25692 13245
rect 25626 13165 25692 13181
rect 25626 13101 25627 13165
rect 25691 13101 25692 13165
rect 25626 13085 25692 13101
rect 25626 13021 25627 13085
rect 25691 13021 25692 13085
rect 25626 13005 25692 13021
rect 25626 12941 25627 13005
rect 25691 12941 25692 13005
rect 25626 12925 25692 12941
rect 25626 12861 25627 12925
rect 25691 12861 25692 12925
rect 25626 12845 25692 12861
rect 25626 12781 25627 12845
rect 25691 12781 25692 12845
rect 25626 12765 25692 12781
rect 25626 12701 25627 12765
rect 25691 12701 25692 12765
rect 25626 12685 25692 12701
rect 25626 12621 25627 12685
rect 25691 12621 25692 12685
rect 25626 12467 25692 12621
rect 25752 12467 25812 13499
rect 25872 12529 25932 13559
rect 25992 12467 26052 13499
rect 26112 12529 26172 13559
rect 26358 13506 26468 13559
rect 26532 13506 26676 13570
rect 26232 13405 26298 13495
rect 26232 13341 26233 13405
rect 26297 13341 26298 13405
rect 26232 13325 26298 13341
rect 26232 13261 26233 13325
rect 26297 13261 26298 13325
rect 26232 13245 26298 13261
rect 26232 13181 26233 13245
rect 26297 13181 26298 13245
rect 26232 13165 26298 13181
rect 26232 13101 26233 13165
rect 26297 13101 26298 13165
rect 26232 13085 26298 13101
rect 26232 13021 26233 13085
rect 26297 13021 26298 13085
rect 26232 13005 26298 13021
rect 26232 12941 26233 13005
rect 26297 12941 26298 13005
rect 26232 12925 26298 12941
rect 26232 12861 26233 12925
rect 26297 12861 26298 12925
rect 26232 12845 26298 12861
rect 26232 12781 26233 12845
rect 26297 12781 26298 12845
rect 26232 12765 26298 12781
rect 26232 12701 26233 12765
rect 26297 12701 26298 12765
rect 26232 12685 26298 12701
rect 26232 12621 26233 12685
rect 26297 12621 26298 12685
rect 26358 13426 26676 13506
rect 26358 13362 26473 13426
rect 26537 13362 26676 13426
rect 26358 13274 26676 13362
rect 26358 13210 26474 13274
rect 26538 13210 26676 13274
rect 26358 13104 26676 13210
rect 26358 13040 26474 13104
rect 26538 13040 26676 13104
rect 26358 12947 26676 13040
rect 26358 12883 26473 12947
rect 26537 12883 26676 12947
rect 26358 12705 26676 12883
rect 26358 12641 26391 12705
rect 26455 12641 26676 12705
rect 26358 12629 26676 12641
rect 26232 12467 26298 12621
rect 21384 12465 26298 12467
rect 21384 12401 21488 12465
rect 21552 12401 21568 12465
rect 21632 12401 21648 12465
rect 21712 12401 21728 12465
rect 21792 12401 21808 12465
rect 21872 12401 21888 12465
rect 21952 12401 22094 12465
rect 22158 12401 22174 12465
rect 22238 12401 22254 12465
rect 22318 12401 22334 12465
rect 22398 12401 22414 12465
rect 22478 12401 22494 12465
rect 22558 12401 22700 12465
rect 22764 12401 22780 12465
rect 22844 12401 22860 12465
rect 22924 12401 22940 12465
rect 23004 12401 23020 12465
rect 23084 12401 23100 12465
rect 23164 12401 23306 12465
rect 23370 12401 23386 12465
rect 23450 12401 23466 12465
rect 23530 12401 23546 12465
rect 23610 12401 23626 12465
rect 23690 12401 23706 12465
rect 23770 12401 23912 12465
rect 23976 12401 23992 12465
rect 24056 12401 24072 12465
rect 24136 12401 24152 12465
rect 24216 12401 24232 12465
rect 24296 12401 24312 12465
rect 24376 12401 24518 12465
rect 24582 12401 24598 12465
rect 24662 12401 24678 12465
rect 24742 12401 24758 12465
rect 24822 12401 24838 12465
rect 24902 12401 24918 12465
rect 24982 12401 25124 12465
rect 25188 12401 25204 12465
rect 25268 12401 25284 12465
rect 25348 12401 25364 12465
rect 25428 12401 25444 12465
rect 25508 12401 25524 12465
rect 25588 12401 25730 12465
rect 25794 12401 25810 12465
rect 25874 12401 25890 12465
rect 25954 12401 25970 12465
rect 26034 12401 26050 12465
rect 26114 12401 26130 12465
rect 26194 12401 26298 12465
rect 21384 12399 26298 12401
rect 26358 12444 26556 12454
rect 20652 12396 21324 12398
rect 26358 12380 26479 12444
rect 26543 12380 26556 12444
rect 26358 12370 26556 12380
rect 21003 12217 21675 12219
rect 21003 12153 21107 12217
rect 21171 12153 21187 12217
rect 21251 12153 21267 12217
rect 21331 12153 21347 12217
rect 21411 12153 21427 12217
rect 21491 12153 21507 12217
rect 21571 12153 21675 12217
rect 21003 12151 21675 12153
rect 21003 11997 21069 12151
rect 21003 11933 21004 11997
rect 21068 11933 21069 11997
rect 21003 11917 21069 11933
rect 21003 11853 21004 11917
rect 21068 11853 21069 11917
rect 21003 11837 21069 11853
rect 21003 11773 21004 11837
rect 21068 11773 21069 11837
rect 21003 11757 21069 11773
rect 21003 11693 21004 11757
rect 21068 11693 21069 11757
rect 21003 11677 21069 11693
rect 21003 11613 21004 11677
rect 21068 11613 21069 11677
rect 21003 11597 21069 11613
rect 21003 11533 21004 11597
rect 21068 11533 21069 11597
rect 21003 11517 21069 11533
rect 21003 11453 21004 11517
rect 21068 11453 21069 11517
rect 21003 11437 21069 11453
rect 21003 11373 21004 11437
rect 21068 11373 21069 11437
rect 21003 11357 21069 11373
rect 21003 11293 21004 11357
rect 21068 11293 21069 11357
rect 21003 11277 21069 11293
rect 21003 11213 21004 11277
rect 21068 11213 21069 11277
rect 21003 11123 21069 11213
rect 20615 11058 20740 11064
rect 21129 11059 21189 12089
rect 21249 11119 21309 12151
rect 21369 11059 21429 12089
rect 21489 11119 21549 12151
rect 21609 11997 21675 12151
rect 21609 11933 21610 11997
rect 21674 11933 21675 11997
rect 21609 11917 21675 11933
rect 21609 11853 21610 11917
rect 21674 11853 21675 11917
rect 21609 11837 21675 11853
rect 21609 11773 21610 11837
rect 21674 11773 21675 11837
rect 21609 11757 21675 11773
rect 21609 11693 21610 11757
rect 21674 11693 21675 11757
rect 21609 11677 21675 11693
rect 21609 11613 21610 11677
rect 21674 11613 21675 11677
rect 21609 11597 21675 11613
rect 21609 11533 21610 11597
rect 21674 11533 21675 11597
rect 21609 11517 21675 11533
rect 21609 11453 21610 11517
rect 21674 11453 21675 11517
rect 21609 11437 21675 11453
rect 21609 11373 21610 11437
rect 21674 11373 21675 11437
rect 21609 11357 21675 11373
rect 21609 11293 21610 11357
rect 21674 11293 21675 11357
rect 21609 11277 21675 11293
rect 21609 11213 21610 11277
rect 21674 11213 21675 11277
rect 21609 11123 21675 11213
rect 21735 12217 24225 12219
rect 21735 12153 21839 12217
rect 21903 12153 21919 12217
rect 21983 12153 21999 12217
rect 22063 12153 22079 12217
rect 22143 12153 22159 12217
rect 22223 12153 22239 12217
rect 22303 12153 22445 12217
rect 22509 12153 22525 12217
rect 22589 12153 22605 12217
rect 22669 12153 22685 12217
rect 22749 12153 22765 12217
rect 22829 12153 22845 12217
rect 22909 12153 23051 12217
rect 23115 12153 23131 12217
rect 23195 12153 23211 12217
rect 23275 12153 23291 12217
rect 23355 12153 23371 12217
rect 23435 12153 23451 12217
rect 23515 12153 23657 12217
rect 23721 12153 23737 12217
rect 23801 12153 23817 12217
rect 23881 12153 23897 12217
rect 23961 12153 23977 12217
rect 24041 12153 24057 12217
rect 24121 12153 24225 12217
rect 21735 12151 24225 12153
rect 21735 11997 21801 12151
rect 21735 11933 21736 11997
rect 21800 11933 21801 11997
rect 21735 11917 21801 11933
rect 21735 11853 21736 11917
rect 21800 11853 21801 11917
rect 21735 11837 21801 11853
rect 21735 11773 21736 11837
rect 21800 11773 21801 11837
rect 21735 11757 21801 11773
rect 21735 11693 21736 11757
rect 21800 11693 21801 11757
rect 21735 11677 21801 11693
rect 21735 11613 21736 11677
rect 21800 11613 21801 11677
rect 21735 11597 21801 11613
rect 21735 11533 21736 11597
rect 21800 11533 21801 11597
rect 21735 11517 21801 11533
rect 21735 11453 21736 11517
rect 21800 11453 21801 11517
rect 21735 11437 21801 11453
rect 21735 11373 21736 11437
rect 21800 11373 21801 11437
rect 21735 11357 21801 11373
rect 21735 11293 21736 11357
rect 21800 11293 21801 11357
rect 21735 11277 21801 11293
rect 21735 11213 21736 11277
rect 21800 11213 21801 11277
rect 21735 11123 21801 11213
rect 21861 11059 21921 12089
rect 21981 11119 22041 12151
rect 22101 11059 22161 12089
rect 22221 11119 22281 12151
rect 22341 11997 22407 12151
rect 22341 11933 22342 11997
rect 22406 11933 22407 11997
rect 22341 11917 22407 11933
rect 22341 11853 22342 11917
rect 22406 11853 22407 11917
rect 22341 11837 22407 11853
rect 22341 11773 22342 11837
rect 22406 11773 22407 11837
rect 22341 11757 22407 11773
rect 22341 11693 22342 11757
rect 22406 11693 22407 11757
rect 22341 11677 22407 11693
rect 22341 11613 22342 11677
rect 22406 11613 22407 11677
rect 22341 11597 22407 11613
rect 22341 11533 22342 11597
rect 22406 11533 22407 11597
rect 22341 11517 22407 11533
rect 22341 11453 22342 11517
rect 22406 11453 22407 11517
rect 22341 11437 22407 11453
rect 22341 11373 22342 11437
rect 22406 11373 22407 11437
rect 22341 11357 22407 11373
rect 22341 11293 22342 11357
rect 22406 11293 22407 11357
rect 22341 11277 22407 11293
rect 22341 11213 22342 11277
rect 22406 11213 22407 11277
rect 22341 11123 22407 11213
rect 22467 11119 22527 12151
rect 22587 11059 22647 12089
rect 22707 11119 22767 12151
rect 22827 11059 22887 12089
rect 22947 11997 23013 12151
rect 22947 11933 22948 11997
rect 23012 11933 23013 11997
rect 22947 11917 23013 11933
rect 22947 11853 22948 11917
rect 23012 11853 23013 11917
rect 22947 11837 23013 11853
rect 22947 11773 22948 11837
rect 23012 11773 23013 11837
rect 22947 11757 23013 11773
rect 22947 11693 22948 11757
rect 23012 11693 23013 11757
rect 22947 11677 23013 11693
rect 22947 11613 22948 11677
rect 23012 11613 23013 11677
rect 22947 11597 23013 11613
rect 22947 11533 22948 11597
rect 23012 11533 23013 11597
rect 22947 11517 23013 11533
rect 22947 11453 22948 11517
rect 23012 11453 23013 11517
rect 22947 11437 23013 11453
rect 22947 11373 22948 11437
rect 23012 11373 23013 11437
rect 22947 11357 23013 11373
rect 22947 11293 22948 11357
rect 23012 11293 23013 11357
rect 22947 11277 23013 11293
rect 22947 11213 22948 11277
rect 23012 11213 23013 11277
rect 22947 11123 23013 11213
rect 23073 11059 23133 12089
rect 23193 11119 23253 12151
rect 23313 11059 23373 12089
rect 23433 11119 23493 12151
rect 23553 11997 23619 12151
rect 23553 11933 23554 11997
rect 23618 11933 23619 11997
rect 23553 11917 23619 11933
rect 23553 11853 23554 11917
rect 23618 11853 23619 11917
rect 23553 11837 23619 11853
rect 23553 11773 23554 11837
rect 23618 11773 23619 11837
rect 23553 11757 23619 11773
rect 23553 11693 23554 11757
rect 23618 11693 23619 11757
rect 23553 11677 23619 11693
rect 23553 11613 23554 11677
rect 23618 11613 23619 11677
rect 23553 11597 23619 11613
rect 23553 11533 23554 11597
rect 23618 11533 23619 11597
rect 23553 11517 23619 11533
rect 23553 11453 23554 11517
rect 23618 11453 23619 11517
rect 23553 11437 23619 11453
rect 23553 11373 23554 11437
rect 23618 11373 23619 11437
rect 23553 11357 23619 11373
rect 23553 11293 23554 11357
rect 23618 11293 23619 11357
rect 23553 11277 23619 11293
rect 23553 11213 23554 11277
rect 23618 11213 23619 11277
rect 23553 11123 23619 11213
rect 23679 11119 23739 12151
rect 23799 11059 23859 12089
rect 23919 11119 23979 12151
rect 24039 11059 24099 12089
rect 24159 11997 24225 12151
rect 24159 11933 24160 11997
rect 24224 11933 24225 11997
rect 24159 11917 24225 11933
rect 24159 11853 24160 11917
rect 24224 11853 24225 11917
rect 24159 11837 24225 11853
rect 24159 11773 24160 11837
rect 24224 11773 24225 11837
rect 24159 11757 24225 11773
rect 24159 11693 24160 11757
rect 24224 11693 24225 11757
rect 24159 11677 24225 11693
rect 24159 11613 24160 11677
rect 24224 11613 24225 11677
rect 24159 11597 24225 11613
rect 24159 11533 24160 11597
rect 24224 11533 24225 11597
rect 24159 11517 24225 11533
rect 24159 11453 24160 11517
rect 24224 11453 24225 11517
rect 24159 11437 24225 11453
rect 24159 11373 24160 11437
rect 24224 11373 24225 11437
rect 24159 11357 24225 11373
rect 24159 11293 24160 11357
rect 24224 11293 24225 11357
rect 24159 11277 24225 11293
rect 24159 11213 24160 11277
rect 24224 11213 24225 11277
rect 24159 11123 24225 11213
rect 24285 12217 25563 12219
rect 24285 12153 24389 12217
rect 24453 12153 24469 12217
rect 24533 12153 24549 12217
rect 24613 12153 24629 12217
rect 24693 12153 24709 12217
rect 24773 12153 24789 12217
rect 24853 12153 24995 12217
rect 25059 12153 25075 12217
rect 25139 12153 25155 12217
rect 25219 12153 25235 12217
rect 25299 12153 25315 12217
rect 25379 12153 25395 12217
rect 25459 12153 25563 12217
rect 24285 12151 25563 12153
rect 24285 11997 24351 12151
rect 24285 11933 24286 11997
rect 24350 11933 24351 11997
rect 24285 11917 24351 11933
rect 24285 11853 24286 11917
rect 24350 11853 24351 11917
rect 24285 11837 24351 11853
rect 24285 11773 24286 11837
rect 24350 11773 24351 11837
rect 24285 11757 24351 11773
rect 24285 11693 24286 11757
rect 24350 11693 24351 11757
rect 24285 11677 24351 11693
rect 24285 11613 24286 11677
rect 24350 11613 24351 11677
rect 24285 11597 24351 11613
rect 24285 11533 24286 11597
rect 24350 11533 24351 11597
rect 24285 11517 24351 11533
rect 24285 11453 24286 11517
rect 24350 11453 24351 11517
rect 24285 11437 24351 11453
rect 24285 11373 24286 11437
rect 24350 11373 24351 11437
rect 24285 11357 24351 11373
rect 24285 11293 24286 11357
rect 24350 11293 24351 11357
rect 24285 11277 24351 11293
rect 24285 11213 24286 11277
rect 24350 11213 24351 11277
rect 24285 11123 24351 11213
rect 24411 11059 24471 12089
rect 24531 11119 24591 12151
rect 24651 11059 24711 12089
rect 24771 11119 24831 12151
rect 24891 11997 24957 12151
rect 24891 11933 24892 11997
rect 24956 11933 24957 11997
rect 24891 11917 24957 11933
rect 24891 11853 24892 11917
rect 24956 11853 24957 11917
rect 24891 11837 24957 11853
rect 24891 11773 24892 11837
rect 24956 11773 24957 11837
rect 24891 11757 24957 11773
rect 24891 11693 24892 11757
rect 24956 11693 24957 11757
rect 24891 11677 24957 11693
rect 24891 11613 24892 11677
rect 24956 11613 24957 11677
rect 24891 11597 24957 11613
rect 24891 11533 24892 11597
rect 24956 11533 24957 11597
rect 24891 11517 24957 11533
rect 24891 11453 24892 11517
rect 24956 11453 24957 11517
rect 24891 11437 24957 11453
rect 24891 11373 24892 11437
rect 24956 11373 24957 11437
rect 24891 11357 24957 11373
rect 24891 11293 24892 11357
rect 24956 11293 24957 11357
rect 24891 11277 24957 11293
rect 24891 11213 24892 11277
rect 24956 11213 24957 11277
rect 24891 11123 24957 11213
rect 25017 11119 25077 12151
rect 25137 11059 25197 12089
rect 25257 11119 25317 12151
rect 25377 11059 25437 12089
rect 25497 11997 25563 12151
rect 25497 11933 25498 11997
rect 25562 11933 25563 11997
rect 25497 11917 25563 11933
rect 25497 11853 25498 11917
rect 25562 11853 25563 11917
rect 25497 11837 25563 11853
rect 25497 11773 25498 11837
rect 25562 11773 25563 11837
rect 25497 11757 25563 11773
rect 25497 11693 25498 11757
rect 25562 11693 25563 11757
rect 25497 11677 25563 11693
rect 25497 11613 25498 11677
rect 25562 11613 25563 11677
rect 25497 11597 25563 11613
rect 25497 11533 25498 11597
rect 25562 11533 25563 11597
rect 25497 11517 25563 11533
rect 25497 11453 25498 11517
rect 25562 11453 25563 11517
rect 25497 11437 25563 11453
rect 25497 11373 25498 11437
rect 25562 11373 25563 11437
rect 25497 11357 25563 11373
rect 25497 11293 25498 11357
rect 25562 11293 25563 11357
rect 25497 11277 25563 11293
rect 25497 11213 25498 11277
rect 25562 11213 25563 11277
rect 25497 11123 25563 11213
rect 25625 12217 26297 12219
rect 25625 12153 25729 12217
rect 25793 12153 25809 12217
rect 25873 12153 25889 12217
rect 25953 12153 25969 12217
rect 26033 12153 26049 12217
rect 26113 12153 26129 12217
rect 26193 12153 26297 12217
rect 25625 12151 26297 12153
rect 25625 11997 25691 12151
rect 25625 11933 25626 11997
rect 25690 11933 25691 11997
rect 25625 11917 25691 11933
rect 25625 11853 25626 11917
rect 25690 11853 25691 11917
rect 25625 11837 25691 11853
rect 25625 11773 25626 11837
rect 25690 11773 25691 11837
rect 25625 11757 25691 11773
rect 25625 11693 25626 11757
rect 25690 11693 25691 11757
rect 25625 11677 25691 11693
rect 25625 11613 25626 11677
rect 25690 11613 25691 11677
rect 25625 11597 25691 11613
rect 25625 11533 25626 11597
rect 25690 11533 25691 11597
rect 25625 11517 25691 11533
rect 25625 11453 25626 11517
rect 25690 11453 25691 11517
rect 25625 11437 25691 11453
rect 25625 11373 25626 11437
rect 25690 11373 25691 11437
rect 25625 11357 25691 11373
rect 25625 11293 25626 11357
rect 25690 11293 25691 11357
rect 25625 11277 25691 11293
rect 25625 11213 25626 11277
rect 25690 11213 25691 11277
rect 25625 11123 25691 11213
rect 25751 11119 25811 12151
rect 25871 11059 25931 12089
rect 25991 11119 26051 12151
rect 26111 11059 26171 12089
rect 26231 11997 26297 12151
rect 26231 11933 26232 11997
rect 26296 11933 26297 11997
rect 26231 11917 26297 11933
rect 26231 11853 26232 11917
rect 26296 11853 26297 11917
rect 26231 11837 26297 11853
rect 26231 11773 26232 11837
rect 26296 11773 26297 11837
rect 26231 11757 26297 11773
rect 26231 11693 26232 11757
rect 26296 11693 26297 11757
rect 26231 11677 26297 11693
rect 26231 11613 26232 11677
rect 26296 11613 26297 11677
rect 26231 11597 26297 11613
rect 26231 11533 26232 11597
rect 26296 11533 26297 11597
rect 26231 11517 26297 11533
rect 26231 11453 26232 11517
rect 26296 11453 26297 11517
rect 26231 11437 26297 11453
rect 26231 11373 26232 11437
rect 26296 11373 26297 11437
rect 26231 11357 26297 11373
rect 26231 11293 26232 11357
rect 26296 11293 26297 11357
rect 26231 11277 26297 11293
rect 26231 11213 26232 11277
rect 26296 11213 26297 11277
rect 26231 11123 26297 11213
rect 26358 11989 26418 12370
rect 26616 12251 26676 12629
rect 26478 12241 26676 12251
rect 26478 12177 26479 12241
rect 26543 12177 26676 12241
rect 26478 12167 26676 12177
rect 26358 11979 26676 11989
rect 26358 11915 26388 11979
rect 26452 11915 26676 11979
rect 21003 11058 21675 11059
rect 21735 11058 24225 11059
rect 24285 11058 25563 11059
rect 25625 11058 26297 11059
rect 26358 11058 26676 11915
rect 20055 11057 26676 11058
rect 20055 11054 21187 11057
rect 20055 11044 20645 11054
rect 19404 10993 20645 11044
rect 14000 10990 20645 10993
rect 20709 10993 21187 11054
rect 21251 10993 21267 11057
rect 21331 10993 21347 11057
rect 21411 10993 21427 11057
rect 21491 10993 21919 11057
rect 21983 10993 21999 11057
rect 22063 10993 22079 11057
rect 22143 10993 22159 11057
rect 22223 10993 22525 11057
rect 22589 10993 22605 11057
rect 22669 10993 22685 11057
rect 22749 10993 22765 11057
rect 22829 10993 23131 11057
rect 23195 10993 23211 11057
rect 23275 10993 23291 11057
rect 23355 10993 23371 11057
rect 23435 10993 23737 11057
rect 23801 10993 23817 11057
rect 23881 10993 23897 11057
rect 23961 10993 23977 11057
rect 24041 10993 24469 11057
rect 24533 10993 24549 11057
rect 24613 10993 24629 11057
rect 24693 10993 24709 11057
rect 24773 10993 25075 11057
rect 25139 10993 25155 11057
rect 25219 10993 25235 11057
rect 25299 10993 25315 11057
rect 25379 10993 25809 11057
rect 25873 10993 25889 11057
rect 25953 10993 25969 11057
rect 26033 10993 26049 11057
rect 26113 10993 26676 11057
rect 20709 10990 26676 10993
rect 10878 10761 26676 10990
rect 2458 10141 9078 10505
rect 10878 10413 14145 10761
rect 2458 10131 9079 10141
rect 2458 10067 3048 10131
rect 3112 10128 9079 10131
rect 3112 10067 3590 10128
rect 2458 10064 3590 10067
rect 3654 10064 3670 10128
rect 3734 10064 3750 10128
rect 3814 10064 3830 10128
rect 3894 10064 4322 10128
rect 4386 10064 4402 10128
rect 4466 10064 4482 10128
rect 4546 10064 4562 10128
rect 4626 10064 4928 10128
rect 4992 10064 5008 10128
rect 5072 10064 5088 10128
rect 5152 10064 5168 10128
rect 5232 10064 5534 10128
rect 5598 10064 5614 10128
rect 5678 10064 5694 10128
rect 5758 10064 5774 10128
rect 5838 10064 6140 10128
rect 6204 10064 6220 10128
rect 6284 10064 6300 10128
rect 6364 10064 6380 10128
rect 6444 10064 6872 10128
rect 6936 10064 6952 10128
rect 7016 10064 7032 10128
rect 7096 10064 7112 10128
rect 7176 10064 7478 10128
rect 7542 10064 7558 10128
rect 7622 10064 7638 10128
rect 7702 10064 7718 10128
rect 7782 10064 8212 10128
rect 8276 10064 8292 10128
rect 8356 10064 8372 10128
rect 8436 10064 8452 10128
rect 8516 10064 9079 10128
rect 2458 10063 9079 10064
rect 2458 8704 2834 10063
rect 3018 10057 3143 10063
rect 3406 10062 4078 10063
rect 4138 10062 6628 10063
rect 6688 10062 7966 10063
rect 8028 10062 8700 10063
rect 3406 9908 3472 9998
rect 3406 9844 3407 9908
rect 3471 9844 3472 9908
rect 3406 9828 3472 9844
rect 3406 9764 3407 9828
rect 3471 9764 3472 9828
rect 3406 9748 3472 9764
rect 3406 9684 3407 9748
rect 3471 9684 3472 9748
rect 3406 9668 3472 9684
rect 3406 9604 3407 9668
rect 3471 9604 3472 9668
rect 3406 9588 3472 9604
rect 3406 9524 3407 9588
rect 3471 9524 3472 9588
rect 3406 9508 3472 9524
rect 3406 9444 3407 9508
rect 3471 9444 3472 9508
rect 3406 9428 3472 9444
rect 3406 9364 3407 9428
rect 3471 9364 3472 9428
rect 3406 9348 3472 9364
rect 3406 9284 3407 9348
rect 3471 9284 3472 9348
rect 3406 9268 3472 9284
rect 3406 9204 3407 9268
rect 3471 9204 3472 9268
rect 3406 9188 3472 9204
rect 3406 9124 3407 9188
rect 3471 9124 3472 9188
rect 3406 8970 3472 9124
rect 3532 9032 3592 10062
rect 3652 8970 3712 10002
rect 3772 9032 3832 10062
rect 3892 8970 3952 10002
rect 4012 9908 4078 9998
rect 4012 9844 4013 9908
rect 4077 9844 4078 9908
rect 4012 9828 4078 9844
rect 4012 9764 4013 9828
rect 4077 9764 4078 9828
rect 4012 9748 4078 9764
rect 4012 9684 4013 9748
rect 4077 9684 4078 9748
rect 4012 9668 4078 9684
rect 4012 9604 4013 9668
rect 4077 9604 4078 9668
rect 4012 9588 4078 9604
rect 4012 9524 4013 9588
rect 4077 9524 4078 9588
rect 4012 9508 4078 9524
rect 4012 9444 4013 9508
rect 4077 9444 4078 9508
rect 4012 9428 4078 9444
rect 4012 9364 4013 9428
rect 4077 9364 4078 9428
rect 4012 9348 4078 9364
rect 4012 9284 4013 9348
rect 4077 9284 4078 9348
rect 4012 9268 4078 9284
rect 4012 9204 4013 9268
rect 4077 9204 4078 9268
rect 4012 9188 4078 9204
rect 4012 9124 4013 9188
rect 4077 9124 4078 9188
rect 4012 8970 4078 9124
rect 3406 8968 4078 8970
rect 3406 8904 3510 8968
rect 3574 8904 3590 8968
rect 3654 8904 3670 8968
rect 3734 8904 3750 8968
rect 3814 8904 3830 8968
rect 3894 8904 3910 8968
rect 3974 8904 4078 8968
rect 3406 8902 4078 8904
rect 4138 9908 4204 9998
rect 4138 9844 4139 9908
rect 4203 9844 4204 9908
rect 4138 9828 4204 9844
rect 4138 9764 4139 9828
rect 4203 9764 4204 9828
rect 4138 9748 4204 9764
rect 4138 9684 4139 9748
rect 4203 9684 4204 9748
rect 4138 9668 4204 9684
rect 4138 9604 4139 9668
rect 4203 9604 4204 9668
rect 4138 9588 4204 9604
rect 4138 9524 4139 9588
rect 4203 9524 4204 9588
rect 4138 9508 4204 9524
rect 4138 9444 4139 9508
rect 4203 9444 4204 9508
rect 4138 9428 4204 9444
rect 4138 9364 4139 9428
rect 4203 9364 4204 9428
rect 4138 9348 4204 9364
rect 4138 9284 4139 9348
rect 4203 9284 4204 9348
rect 4138 9268 4204 9284
rect 4138 9204 4139 9268
rect 4203 9204 4204 9268
rect 4138 9188 4204 9204
rect 4138 9124 4139 9188
rect 4203 9124 4204 9188
rect 4138 8970 4204 9124
rect 4264 9032 4324 10062
rect 4384 8970 4444 10002
rect 4504 9032 4564 10062
rect 4624 8970 4684 10002
rect 4744 9908 4810 9998
rect 4744 9844 4745 9908
rect 4809 9844 4810 9908
rect 4744 9828 4810 9844
rect 4744 9764 4745 9828
rect 4809 9764 4810 9828
rect 4744 9748 4810 9764
rect 4744 9684 4745 9748
rect 4809 9684 4810 9748
rect 4744 9668 4810 9684
rect 4744 9604 4745 9668
rect 4809 9604 4810 9668
rect 4744 9588 4810 9604
rect 4744 9524 4745 9588
rect 4809 9524 4810 9588
rect 4744 9508 4810 9524
rect 4744 9444 4745 9508
rect 4809 9444 4810 9508
rect 4744 9428 4810 9444
rect 4744 9364 4745 9428
rect 4809 9364 4810 9428
rect 4744 9348 4810 9364
rect 4744 9284 4745 9348
rect 4809 9284 4810 9348
rect 4744 9268 4810 9284
rect 4744 9204 4745 9268
rect 4809 9204 4810 9268
rect 4744 9188 4810 9204
rect 4744 9124 4745 9188
rect 4809 9124 4810 9188
rect 4744 8970 4810 9124
rect 4870 8970 4930 10002
rect 4990 9032 5050 10062
rect 5110 8970 5170 10002
rect 5230 9032 5290 10062
rect 5350 9908 5416 9998
rect 5350 9844 5351 9908
rect 5415 9844 5416 9908
rect 5350 9828 5416 9844
rect 5350 9764 5351 9828
rect 5415 9764 5416 9828
rect 5350 9748 5416 9764
rect 5350 9684 5351 9748
rect 5415 9684 5416 9748
rect 5350 9668 5416 9684
rect 5350 9604 5351 9668
rect 5415 9604 5416 9668
rect 5350 9588 5416 9604
rect 5350 9524 5351 9588
rect 5415 9524 5416 9588
rect 5350 9508 5416 9524
rect 5350 9444 5351 9508
rect 5415 9444 5416 9508
rect 5350 9428 5416 9444
rect 5350 9364 5351 9428
rect 5415 9364 5416 9428
rect 5350 9348 5416 9364
rect 5350 9284 5351 9348
rect 5415 9284 5416 9348
rect 5350 9268 5416 9284
rect 5350 9204 5351 9268
rect 5415 9204 5416 9268
rect 5350 9188 5416 9204
rect 5350 9124 5351 9188
rect 5415 9124 5416 9188
rect 5350 8970 5416 9124
rect 5476 9032 5536 10062
rect 5596 8970 5656 10002
rect 5716 9032 5776 10062
rect 5836 8970 5896 10002
rect 5956 9908 6022 9998
rect 5956 9844 5957 9908
rect 6021 9844 6022 9908
rect 5956 9828 6022 9844
rect 5956 9764 5957 9828
rect 6021 9764 6022 9828
rect 5956 9748 6022 9764
rect 5956 9684 5957 9748
rect 6021 9684 6022 9748
rect 5956 9668 6022 9684
rect 5956 9604 5957 9668
rect 6021 9604 6022 9668
rect 5956 9588 6022 9604
rect 5956 9524 5957 9588
rect 6021 9524 6022 9588
rect 5956 9508 6022 9524
rect 5956 9444 5957 9508
rect 6021 9444 6022 9508
rect 5956 9428 6022 9444
rect 5956 9364 5957 9428
rect 6021 9364 6022 9428
rect 5956 9348 6022 9364
rect 5956 9284 5957 9348
rect 6021 9284 6022 9348
rect 5956 9268 6022 9284
rect 5956 9204 5957 9268
rect 6021 9204 6022 9268
rect 5956 9188 6022 9204
rect 5956 9124 5957 9188
rect 6021 9124 6022 9188
rect 5956 8970 6022 9124
rect 6082 8970 6142 10002
rect 6202 9032 6262 10062
rect 6322 8970 6382 10002
rect 6442 9032 6502 10062
rect 6562 9908 6628 9998
rect 6562 9844 6563 9908
rect 6627 9844 6628 9908
rect 6562 9828 6628 9844
rect 6562 9764 6563 9828
rect 6627 9764 6628 9828
rect 6562 9748 6628 9764
rect 6562 9684 6563 9748
rect 6627 9684 6628 9748
rect 6562 9668 6628 9684
rect 6562 9604 6563 9668
rect 6627 9604 6628 9668
rect 6562 9588 6628 9604
rect 6562 9524 6563 9588
rect 6627 9524 6628 9588
rect 6562 9508 6628 9524
rect 6562 9444 6563 9508
rect 6627 9444 6628 9508
rect 6562 9428 6628 9444
rect 6562 9364 6563 9428
rect 6627 9364 6628 9428
rect 6562 9348 6628 9364
rect 6562 9284 6563 9348
rect 6627 9284 6628 9348
rect 6562 9268 6628 9284
rect 6562 9204 6563 9268
rect 6627 9204 6628 9268
rect 6562 9188 6628 9204
rect 6562 9124 6563 9188
rect 6627 9124 6628 9188
rect 6562 8970 6628 9124
rect 4138 8968 6628 8970
rect 4138 8904 4242 8968
rect 4306 8904 4322 8968
rect 4386 8904 4402 8968
rect 4466 8904 4482 8968
rect 4546 8904 4562 8968
rect 4626 8904 4642 8968
rect 4706 8904 4848 8968
rect 4912 8904 4928 8968
rect 4992 8904 5008 8968
rect 5072 8904 5088 8968
rect 5152 8904 5168 8968
rect 5232 8904 5248 8968
rect 5312 8904 5454 8968
rect 5518 8904 5534 8968
rect 5598 8904 5614 8968
rect 5678 8904 5694 8968
rect 5758 8904 5774 8968
rect 5838 8904 5854 8968
rect 5918 8904 6060 8968
rect 6124 8904 6140 8968
rect 6204 8904 6220 8968
rect 6284 8904 6300 8968
rect 6364 8904 6380 8968
rect 6444 8904 6460 8968
rect 6524 8904 6628 8968
rect 4138 8902 6628 8904
rect 6688 9908 6754 9998
rect 6688 9844 6689 9908
rect 6753 9844 6754 9908
rect 6688 9828 6754 9844
rect 6688 9764 6689 9828
rect 6753 9764 6754 9828
rect 6688 9748 6754 9764
rect 6688 9684 6689 9748
rect 6753 9684 6754 9748
rect 6688 9668 6754 9684
rect 6688 9604 6689 9668
rect 6753 9604 6754 9668
rect 6688 9588 6754 9604
rect 6688 9524 6689 9588
rect 6753 9524 6754 9588
rect 6688 9508 6754 9524
rect 6688 9444 6689 9508
rect 6753 9444 6754 9508
rect 6688 9428 6754 9444
rect 6688 9364 6689 9428
rect 6753 9364 6754 9428
rect 6688 9348 6754 9364
rect 6688 9284 6689 9348
rect 6753 9284 6754 9348
rect 6688 9268 6754 9284
rect 6688 9204 6689 9268
rect 6753 9204 6754 9268
rect 6688 9188 6754 9204
rect 6688 9124 6689 9188
rect 6753 9124 6754 9188
rect 6688 8970 6754 9124
rect 6814 9032 6874 10062
rect 6934 8970 6994 10002
rect 7054 9032 7114 10062
rect 7174 8970 7234 10002
rect 7294 9908 7360 9998
rect 7294 9844 7295 9908
rect 7359 9844 7360 9908
rect 7294 9828 7360 9844
rect 7294 9764 7295 9828
rect 7359 9764 7360 9828
rect 7294 9748 7360 9764
rect 7294 9684 7295 9748
rect 7359 9684 7360 9748
rect 7294 9668 7360 9684
rect 7294 9604 7295 9668
rect 7359 9604 7360 9668
rect 7294 9588 7360 9604
rect 7294 9524 7295 9588
rect 7359 9524 7360 9588
rect 7294 9508 7360 9524
rect 7294 9444 7295 9508
rect 7359 9444 7360 9508
rect 7294 9428 7360 9444
rect 7294 9364 7295 9428
rect 7359 9364 7360 9428
rect 7294 9348 7360 9364
rect 7294 9284 7295 9348
rect 7359 9284 7360 9348
rect 7294 9268 7360 9284
rect 7294 9204 7295 9268
rect 7359 9204 7360 9268
rect 7294 9188 7360 9204
rect 7294 9124 7295 9188
rect 7359 9124 7360 9188
rect 7294 8970 7360 9124
rect 7420 8970 7480 10002
rect 7540 9032 7600 10062
rect 7660 8970 7720 10002
rect 7780 9032 7840 10062
rect 7900 9908 7966 9998
rect 7900 9844 7901 9908
rect 7965 9844 7966 9908
rect 7900 9828 7966 9844
rect 7900 9764 7901 9828
rect 7965 9764 7966 9828
rect 7900 9748 7966 9764
rect 7900 9684 7901 9748
rect 7965 9684 7966 9748
rect 7900 9668 7966 9684
rect 7900 9604 7901 9668
rect 7965 9604 7966 9668
rect 7900 9588 7966 9604
rect 7900 9524 7901 9588
rect 7965 9524 7966 9588
rect 7900 9508 7966 9524
rect 7900 9444 7901 9508
rect 7965 9444 7966 9508
rect 7900 9428 7966 9444
rect 7900 9364 7901 9428
rect 7965 9364 7966 9428
rect 7900 9348 7966 9364
rect 7900 9284 7901 9348
rect 7965 9284 7966 9348
rect 7900 9268 7966 9284
rect 7900 9204 7901 9268
rect 7965 9204 7966 9268
rect 7900 9188 7966 9204
rect 7900 9124 7901 9188
rect 7965 9124 7966 9188
rect 7900 8970 7966 9124
rect 6688 8968 7966 8970
rect 6688 8904 6792 8968
rect 6856 8904 6872 8968
rect 6936 8904 6952 8968
rect 7016 8904 7032 8968
rect 7096 8904 7112 8968
rect 7176 8904 7192 8968
rect 7256 8904 7398 8968
rect 7462 8904 7478 8968
rect 7542 8904 7558 8968
rect 7622 8904 7638 8968
rect 7702 8904 7718 8968
rect 7782 8904 7798 8968
rect 7862 8904 7966 8968
rect 6688 8902 7966 8904
rect 8028 9908 8094 9998
rect 8028 9844 8029 9908
rect 8093 9844 8094 9908
rect 8028 9828 8094 9844
rect 8028 9764 8029 9828
rect 8093 9764 8094 9828
rect 8028 9748 8094 9764
rect 8028 9684 8029 9748
rect 8093 9684 8094 9748
rect 8028 9668 8094 9684
rect 8028 9604 8029 9668
rect 8093 9604 8094 9668
rect 8028 9588 8094 9604
rect 8028 9524 8029 9588
rect 8093 9524 8094 9588
rect 8028 9508 8094 9524
rect 8028 9444 8029 9508
rect 8093 9444 8094 9508
rect 8028 9428 8094 9444
rect 8028 9364 8029 9428
rect 8093 9364 8094 9428
rect 8028 9348 8094 9364
rect 8028 9284 8029 9348
rect 8093 9284 8094 9348
rect 8028 9268 8094 9284
rect 8028 9204 8029 9268
rect 8093 9204 8094 9268
rect 8028 9188 8094 9204
rect 8028 9124 8029 9188
rect 8093 9124 8094 9188
rect 8028 8970 8094 9124
rect 8154 8970 8214 10002
rect 8274 9032 8334 10062
rect 8394 8970 8454 10002
rect 8514 9032 8574 10062
rect 8634 9908 8700 9998
rect 8634 9844 8635 9908
rect 8699 9844 8700 9908
rect 8634 9828 8700 9844
rect 8634 9764 8635 9828
rect 8699 9764 8700 9828
rect 8634 9748 8700 9764
rect 8634 9684 8635 9748
rect 8699 9684 8700 9748
rect 8634 9668 8700 9684
rect 8634 9604 8635 9668
rect 8699 9604 8700 9668
rect 8634 9588 8700 9604
rect 8634 9524 8635 9588
rect 8699 9524 8700 9588
rect 8634 9508 8700 9524
rect 8634 9444 8635 9508
rect 8699 9444 8700 9508
rect 8634 9428 8700 9444
rect 8634 9364 8635 9428
rect 8699 9364 8700 9428
rect 8634 9348 8700 9364
rect 8634 9284 8635 9348
rect 8699 9284 8700 9348
rect 8634 9268 8700 9284
rect 8634 9204 8635 9268
rect 8699 9204 8700 9268
rect 8634 9188 8700 9204
rect 8634 9124 8635 9188
rect 8699 9124 8700 9188
rect 8634 8970 8700 9124
rect 8028 8968 8700 8970
rect 8028 8904 8132 8968
rect 8196 8904 8212 8968
rect 8276 8904 8292 8968
rect 8356 8904 8372 8968
rect 8436 8904 8452 8968
rect 8516 8904 8532 8968
rect 8596 8904 8700 8968
rect 8028 8902 8700 8904
rect 8761 9339 9079 10063
rect 10878 10059 12863 10413
rect 13121 10377 14145 10413
rect 15449 10377 15984 10761
rect 17096 10377 17496 10761
rect 18991 10760 26676 10761
rect 18991 10397 20213 10760
rect 21350 10397 21939 10760
rect 22817 10397 23328 10760
rect 24323 10397 24853 10760
rect 25767 10397 26676 10760
rect 18991 10377 26676 10397
rect 13121 10119 26676 10377
rect 13121 10116 19179 10119
rect 13121 10059 13775 10116
rect 10878 10052 13775 10059
rect 13839 10052 13855 10116
rect 13919 10052 13935 10116
rect 13999 10052 14015 10116
rect 14079 10052 14509 10116
rect 14573 10052 14589 10116
rect 14653 10052 14669 10116
rect 14733 10052 14749 10116
rect 14813 10052 15115 10116
rect 15179 10052 15195 10116
rect 15259 10052 15275 10116
rect 15339 10052 15355 10116
rect 15419 10052 15847 10116
rect 15911 10052 15927 10116
rect 15991 10052 16007 10116
rect 16071 10052 16087 10116
rect 16151 10052 16453 10116
rect 16517 10052 16533 10116
rect 16597 10052 16613 10116
rect 16677 10052 16693 10116
rect 16757 10052 17059 10116
rect 17123 10052 17139 10116
rect 17203 10052 17219 10116
rect 17283 10052 17299 10116
rect 17363 10052 17665 10116
rect 17729 10052 17745 10116
rect 17809 10052 17825 10116
rect 17889 10052 17905 10116
rect 17969 10052 18397 10116
rect 18461 10052 18477 10116
rect 18541 10052 18557 10116
rect 18621 10052 18637 10116
rect 18701 10055 19179 10116
rect 19243 10116 25888 10119
rect 19243 10111 20484 10116
rect 19243 10055 19833 10111
rect 18701 10052 19833 10055
rect 10878 10051 19833 10052
rect 10878 9962 13530 10051
rect 13591 10050 14263 10051
rect 14325 10050 15603 10051
rect 15663 10050 18153 10051
rect 18213 10050 18885 10051
rect 10878 9608 12874 9962
rect 13132 9608 13530 9962
rect 10878 9486 13530 9608
rect 10878 9481 12886 9486
rect 11374 9339 12886 9481
rect 8761 9206 12886 9339
rect 8761 9142 8791 9206
rect 8855 9171 12886 9206
rect 8855 9168 11583 9171
rect 8855 9165 11098 9168
rect 8855 9142 9219 9165
rect 8761 9101 9219 9142
rect 9283 9101 9696 9165
rect 9760 9162 11098 9165
rect 9760 9154 10492 9162
rect 9760 9101 10116 9154
rect 8761 9090 10116 9101
rect 10180 9098 10492 9154
rect 10556 9098 10840 9162
rect 10904 9104 11098 9162
rect 11162 9104 11324 9168
rect 11388 9107 11583 9168
rect 11647 9150 12886 9171
rect 13144 9194 13530 9486
rect 13144 9152 13436 9194
rect 11647 9140 12954 9150
rect 11647 9134 12858 9140
rect 11647 9133 12422 9134
rect 11647 9107 12190 9133
rect 11388 9104 12190 9107
rect 10904 9098 12190 9104
rect 10180 9090 12190 9098
rect 8761 9080 12190 9090
rect 8761 8751 8821 9080
rect 11053 9069 12190 9080
rect 12254 9070 12422 9133
rect 12486 9076 12858 9134
rect 12922 9132 12954 9140
rect 13063 9142 13436 9152
rect 13063 9132 13093 9142
rect 12922 9078 13093 9132
rect 13157 9130 13436 9142
rect 13500 9130 13530 9194
rect 13157 9120 13530 9130
rect 13157 9078 13269 9120
rect 12922 9076 13269 9078
rect 12486 9070 13269 9076
rect 12254 9069 13269 9070
rect 11053 9022 13269 9069
rect 11053 8999 12195 9022
rect 8881 8944 9079 8954
rect 8881 8880 8882 8944
rect 8946 8880 9079 8944
rect 8881 8870 9079 8880
rect 8761 8741 8959 8751
rect 3055 8723 3727 8725
rect 2456 8640 2463 8704
rect 2527 8640 2583 8704
rect 2647 8640 2726 8704
rect 2790 8640 2833 8704
rect 2456 8625 2833 8640
rect 3055 8659 3159 8723
rect 3223 8659 3239 8723
rect 3303 8659 3319 8723
rect 3383 8659 3399 8723
rect 3463 8659 3479 8723
rect 3543 8659 3559 8723
rect 3623 8659 3727 8723
rect 3055 8657 3727 8659
rect 3055 8503 3121 8657
rect 3055 8439 3056 8503
rect 3120 8439 3121 8503
rect 3055 8423 3121 8439
rect 3055 8359 3056 8423
rect 3120 8359 3121 8423
rect 3055 8343 3121 8359
rect 3055 8279 3056 8343
rect 3120 8279 3121 8343
rect 3055 8263 3121 8279
rect 3055 8199 3056 8263
rect 3120 8199 3121 8263
rect 3055 8183 3121 8199
rect 2430 8159 2847 8177
rect 2430 8158 2576 8159
rect 2430 8094 2445 8158
rect 2509 8095 2576 8158
rect 2640 8158 2847 8159
rect 2640 8095 2720 8158
rect 2509 8094 2720 8095
rect 2784 8100 2847 8158
rect 3055 8119 3056 8183
rect 3120 8119 3121 8183
rect 3055 8103 3121 8119
rect 2784 8094 2848 8100
rect 2064 7562 2848 8094
rect 3055 8039 3056 8103
rect 3120 8039 3121 8103
rect 3055 8023 3121 8039
rect 3055 7959 3056 8023
rect 3120 7959 3121 8023
rect 3055 7943 3121 7959
rect 3055 7879 3056 7943
rect 3120 7879 3121 7943
rect 3055 7863 3121 7879
rect 3055 7799 3056 7863
rect 3120 7799 3121 7863
rect 3055 7783 3121 7799
rect 3055 7719 3056 7783
rect 3120 7719 3121 7783
rect 3055 7629 3121 7719
rect 3181 7565 3241 8595
rect 3301 7625 3361 8657
rect 3421 7565 3481 8595
rect 3541 7625 3601 8657
rect 3661 8503 3727 8657
rect 3661 8439 3662 8503
rect 3726 8439 3727 8503
rect 3661 8423 3727 8439
rect 3661 8359 3662 8423
rect 3726 8359 3727 8423
rect 3661 8343 3727 8359
rect 3661 8279 3662 8343
rect 3726 8279 3727 8343
rect 3661 8263 3727 8279
rect 3661 8199 3662 8263
rect 3726 8199 3727 8263
rect 3661 8183 3727 8199
rect 3661 8119 3662 8183
rect 3726 8119 3727 8183
rect 3661 8103 3727 8119
rect 3661 8039 3662 8103
rect 3726 8039 3727 8103
rect 3661 8023 3727 8039
rect 3661 7959 3662 8023
rect 3726 7959 3727 8023
rect 3661 7943 3727 7959
rect 3661 7879 3662 7943
rect 3726 7879 3727 7943
rect 3661 7863 3727 7879
rect 3661 7799 3662 7863
rect 3726 7799 3727 7863
rect 3661 7783 3727 7799
rect 3661 7719 3662 7783
rect 3726 7719 3727 7783
rect 3661 7629 3727 7719
rect 3787 8720 8701 8722
rect 3787 8656 3891 8720
rect 3955 8656 3971 8720
rect 4035 8656 4051 8720
rect 4115 8656 4131 8720
rect 4195 8656 4211 8720
rect 4275 8656 4291 8720
rect 4355 8656 4497 8720
rect 4561 8656 4577 8720
rect 4641 8656 4657 8720
rect 4721 8656 4737 8720
rect 4801 8656 4817 8720
rect 4881 8656 4897 8720
rect 4961 8656 5103 8720
rect 5167 8656 5183 8720
rect 5247 8656 5263 8720
rect 5327 8656 5343 8720
rect 5407 8656 5423 8720
rect 5487 8656 5503 8720
rect 5567 8656 5709 8720
rect 5773 8656 5789 8720
rect 5853 8656 5869 8720
rect 5933 8656 5949 8720
rect 6013 8656 6029 8720
rect 6093 8656 6109 8720
rect 6173 8656 6315 8720
rect 6379 8656 6395 8720
rect 6459 8656 6475 8720
rect 6539 8656 6555 8720
rect 6619 8656 6635 8720
rect 6699 8656 6715 8720
rect 6779 8656 6921 8720
rect 6985 8656 7001 8720
rect 7065 8656 7081 8720
rect 7145 8656 7161 8720
rect 7225 8656 7241 8720
rect 7305 8656 7321 8720
rect 7385 8656 7527 8720
rect 7591 8656 7607 8720
rect 7671 8656 7687 8720
rect 7751 8656 7767 8720
rect 7831 8656 7847 8720
rect 7911 8656 7927 8720
rect 7991 8656 8133 8720
rect 8197 8656 8213 8720
rect 8277 8656 8293 8720
rect 8357 8656 8373 8720
rect 8437 8656 8453 8720
rect 8517 8656 8533 8720
rect 8597 8656 8701 8720
rect 8761 8677 8882 8741
rect 8946 8677 8959 8741
rect 8761 8667 8959 8677
rect 3787 8654 8701 8656
rect 3787 8500 3853 8654
rect 3787 8436 3788 8500
rect 3852 8436 3853 8500
rect 3787 8420 3853 8436
rect 3787 8356 3788 8420
rect 3852 8356 3853 8420
rect 3787 8340 3853 8356
rect 3787 8276 3788 8340
rect 3852 8276 3853 8340
rect 3787 8260 3853 8276
rect 3787 8196 3788 8260
rect 3852 8196 3853 8260
rect 3787 8180 3853 8196
rect 3787 8116 3788 8180
rect 3852 8116 3853 8180
rect 3787 8100 3853 8116
rect 3787 8036 3788 8100
rect 3852 8036 3853 8100
rect 3787 8020 3853 8036
rect 3787 7956 3788 8020
rect 3852 7956 3853 8020
rect 3787 7940 3853 7956
rect 3787 7876 3788 7940
rect 3852 7876 3853 7940
rect 3787 7860 3853 7876
rect 3787 7796 3788 7860
rect 3852 7796 3853 7860
rect 3787 7780 3853 7796
rect 3787 7716 3788 7780
rect 3852 7716 3853 7780
rect 3787 7626 3853 7716
rect 3055 7564 3727 7565
rect 3055 7563 3728 7564
rect 3055 7562 3159 7563
rect 2064 7553 3159 7562
rect 2064 7489 3062 7553
rect 3126 7499 3159 7553
rect 3223 7499 3239 7563
rect 3303 7499 3319 7563
rect 3383 7499 3399 7563
rect 3463 7499 3479 7563
rect 3543 7499 3559 7563
rect 3623 7562 3728 7563
rect 3913 7562 3973 8592
rect 4033 7622 4093 8654
rect 4153 7562 4213 8592
rect 4273 7622 4333 8654
rect 4393 8500 4459 8654
rect 4393 8436 4394 8500
rect 4458 8436 4459 8500
rect 4393 8420 4459 8436
rect 4393 8356 4394 8420
rect 4458 8356 4459 8420
rect 4393 8340 4459 8356
rect 4393 8276 4394 8340
rect 4458 8276 4459 8340
rect 4393 8260 4459 8276
rect 4393 8196 4394 8260
rect 4458 8196 4459 8260
rect 4393 8180 4459 8196
rect 4393 8116 4394 8180
rect 4458 8116 4459 8180
rect 4393 8100 4459 8116
rect 4393 8036 4394 8100
rect 4458 8036 4459 8100
rect 4393 8020 4459 8036
rect 4393 7956 4394 8020
rect 4458 7956 4459 8020
rect 4393 7940 4459 7956
rect 4393 7876 4394 7940
rect 4458 7876 4459 7940
rect 4393 7860 4459 7876
rect 4393 7796 4394 7860
rect 4458 7796 4459 7860
rect 4393 7780 4459 7796
rect 4393 7716 4394 7780
rect 4458 7716 4459 7780
rect 4393 7626 4459 7716
rect 4519 7622 4579 8654
rect 4639 7562 4699 8592
rect 4759 7622 4819 8654
rect 4879 7562 4939 8592
rect 4999 8500 5065 8654
rect 4999 8436 5000 8500
rect 5064 8436 5065 8500
rect 4999 8420 5065 8436
rect 4999 8356 5000 8420
rect 5064 8356 5065 8420
rect 4999 8340 5065 8356
rect 4999 8276 5000 8340
rect 5064 8276 5065 8340
rect 4999 8260 5065 8276
rect 4999 8196 5000 8260
rect 5064 8196 5065 8260
rect 4999 8180 5065 8196
rect 4999 8116 5000 8180
rect 5064 8116 5065 8180
rect 4999 8100 5065 8116
rect 4999 8036 5000 8100
rect 5064 8036 5065 8100
rect 4999 8020 5065 8036
rect 4999 7956 5000 8020
rect 5064 7956 5065 8020
rect 4999 7940 5065 7956
rect 4999 7876 5000 7940
rect 5064 7876 5065 7940
rect 4999 7860 5065 7876
rect 4999 7796 5000 7860
rect 5064 7796 5065 7860
rect 4999 7780 5065 7796
rect 4999 7716 5000 7780
rect 5064 7716 5065 7780
rect 4999 7626 5065 7716
rect 5125 7562 5185 8592
rect 5245 7622 5305 8654
rect 5365 7562 5425 8592
rect 5485 7622 5545 8654
rect 5605 8500 5671 8654
rect 5605 8436 5606 8500
rect 5670 8436 5671 8500
rect 5605 8420 5671 8436
rect 5605 8356 5606 8420
rect 5670 8356 5671 8420
rect 5605 8340 5671 8356
rect 5605 8276 5606 8340
rect 5670 8276 5671 8340
rect 5605 8260 5671 8276
rect 5605 8196 5606 8260
rect 5670 8196 5671 8260
rect 5605 8180 5671 8196
rect 5605 8116 5606 8180
rect 5670 8116 5671 8180
rect 5605 8100 5671 8116
rect 5605 8036 5606 8100
rect 5670 8036 5671 8100
rect 5605 8020 5671 8036
rect 5605 7956 5606 8020
rect 5670 7956 5671 8020
rect 5605 7940 5671 7956
rect 5605 7876 5606 7940
rect 5670 7876 5671 7940
rect 5605 7860 5671 7876
rect 5605 7796 5606 7860
rect 5670 7796 5671 7860
rect 5605 7780 5671 7796
rect 5605 7716 5606 7780
rect 5670 7716 5671 7780
rect 5605 7626 5671 7716
rect 5731 7622 5791 8654
rect 5851 7562 5911 8592
rect 5971 7622 6031 8654
rect 6091 7562 6151 8592
rect 6211 8500 6277 8654
rect 6211 8436 6212 8500
rect 6276 8436 6277 8500
rect 6211 8420 6277 8436
rect 6211 8356 6212 8420
rect 6276 8356 6277 8420
rect 6211 8340 6277 8356
rect 6211 8276 6212 8340
rect 6276 8276 6277 8340
rect 6211 8260 6277 8276
rect 6211 8196 6212 8260
rect 6276 8196 6277 8260
rect 6211 8180 6277 8196
rect 6211 8116 6212 8180
rect 6276 8116 6277 8180
rect 6211 8100 6277 8116
rect 6211 8036 6212 8100
rect 6276 8036 6277 8100
rect 6211 8020 6277 8036
rect 6211 7956 6212 8020
rect 6276 7956 6277 8020
rect 6211 7940 6277 7956
rect 6211 7876 6212 7940
rect 6276 7876 6277 7940
rect 6211 7860 6277 7876
rect 6211 7796 6212 7860
rect 6276 7796 6277 7860
rect 6211 7780 6277 7796
rect 6211 7716 6212 7780
rect 6276 7716 6277 7780
rect 6211 7626 6277 7716
rect 6337 7562 6397 8592
rect 6457 7622 6517 8654
rect 6577 7562 6637 8592
rect 6697 7622 6757 8654
rect 6817 8500 6883 8654
rect 6817 8436 6818 8500
rect 6882 8436 6883 8500
rect 6817 8420 6883 8436
rect 6817 8356 6818 8420
rect 6882 8356 6883 8420
rect 6817 8340 6883 8356
rect 6817 8276 6818 8340
rect 6882 8276 6883 8340
rect 6817 8260 6883 8276
rect 6817 8196 6818 8260
rect 6882 8196 6883 8260
rect 6817 8180 6883 8196
rect 6817 8116 6818 8180
rect 6882 8116 6883 8180
rect 6817 8100 6883 8116
rect 6817 8036 6818 8100
rect 6882 8036 6883 8100
rect 6817 8020 6883 8036
rect 6817 7956 6818 8020
rect 6882 7956 6883 8020
rect 6817 7940 6883 7956
rect 6817 7876 6818 7940
rect 6882 7876 6883 7940
rect 6817 7860 6883 7876
rect 6817 7796 6818 7860
rect 6882 7796 6883 7860
rect 6817 7780 6883 7796
rect 6817 7716 6818 7780
rect 6882 7716 6883 7780
rect 6817 7626 6883 7716
rect 6943 7622 7003 8654
rect 7063 7562 7123 8592
rect 7183 7622 7243 8654
rect 7303 7562 7363 8592
rect 7423 8500 7489 8654
rect 7423 8436 7424 8500
rect 7488 8436 7489 8500
rect 7423 8420 7489 8436
rect 7423 8356 7424 8420
rect 7488 8356 7489 8420
rect 7423 8340 7489 8356
rect 7423 8276 7424 8340
rect 7488 8276 7489 8340
rect 7423 8260 7489 8276
rect 7423 8196 7424 8260
rect 7488 8196 7489 8260
rect 7423 8180 7489 8196
rect 7423 8116 7424 8180
rect 7488 8116 7489 8180
rect 7423 8100 7489 8116
rect 7423 8036 7424 8100
rect 7488 8036 7489 8100
rect 7423 8020 7489 8036
rect 7423 7956 7424 8020
rect 7488 7956 7489 8020
rect 7423 7940 7489 7956
rect 7423 7876 7424 7940
rect 7488 7876 7489 7940
rect 7423 7860 7489 7876
rect 7423 7796 7424 7860
rect 7488 7796 7489 7860
rect 7423 7780 7489 7796
rect 7423 7716 7424 7780
rect 7488 7716 7489 7780
rect 7423 7626 7489 7716
rect 7549 7562 7609 8592
rect 7669 7622 7729 8654
rect 7789 7562 7849 8592
rect 7909 7622 7969 8654
rect 8029 8500 8095 8654
rect 8029 8436 8030 8500
rect 8094 8436 8095 8500
rect 8029 8420 8095 8436
rect 8029 8356 8030 8420
rect 8094 8356 8095 8420
rect 8029 8340 8095 8356
rect 8029 8276 8030 8340
rect 8094 8276 8095 8340
rect 8029 8260 8095 8276
rect 8029 8196 8030 8260
rect 8094 8196 8095 8260
rect 8029 8180 8095 8196
rect 8029 8116 8030 8180
rect 8094 8116 8095 8180
rect 8029 8100 8095 8116
rect 8029 8036 8030 8100
rect 8094 8036 8095 8100
rect 8029 8020 8095 8036
rect 8029 7956 8030 8020
rect 8094 7956 8095 8020
rect 8029 7940 8095 7956
rect 8029 7876 8030 7940
rect 8094 7876 8095 7940
rect 8029 7860 8095 7876
rect 8029 7796 8030 7860
rect 8094 7796 8095 7860
rect 8029 7780 8095 7796
rect 8029 7716 8030 7780
rect 8094 7716 8095 7780
rect 8029 7626 8095 7716
rect 8155 7622 8215 8654
rect 8275 7562 8335 8592
rect 8395 7622 8455 8654
rect 8515 7562 8575 8592
rect 8635 8500 8701 8654
rect 9019 8564 9079 8870
rect 11053 8700 11710 8999
rect 8635 8436 8636 8500
rect 8700 8436 8701 8500
rect 8771 8492 10955 8564
rect 8635 8420 8701 8436
rect 8635 8356 8636 8420
rect 8700 8356 8701 8420
rect 8635 8340 8701 8356
rect 8635 8276 8636 8340
rect 8700 8276 8701 8340
rect 8635 8260 8701 8276
rect 8635 8196 8636 8260
rect 8700 8196 8701 8260
rect 8635 8180 8701 8196
rect 8635 8116 8636 8180
rect 8700 8116 8701 8180
rect 8635 8100 8701 8116
rect 8635 8036 8636 8100
rect 8700 8036 8701 8100
rect 8635 8020 8701 8036
rect 8635 7956 8636 8020
rect 8700 7956 8701 8020
rect 8635 7940 8701 7956
rect 8635 7876 8636 7940
rect 8700 7876 8701 7940
rect 8635 7860 8701 7876
rect 8635 7796 8636 7860
rect 8700 7796 8701 7860
rect 8635 7780 8701 7796
rect 8635 7716 8636 7780
rect 8700 7716 8701 7780
rect 8635 7626 8701 7716
rect 8761 8480 10955 8492
rect 8761 8416 8794 8480
rect 8858 8455 10955 8480
rect 8858 8454 9466 8455
rect 8858 8416 9204 8454
rect 8761 8390 9204 8416
rect 9268 8391 9466 8454
rect 9530 8391 9738 8455
rect 9802 8391 10065 8455
rect 10129 8391 10446 8455
rect 10510 8391 10823 8455
rect 10887 8391 10955 8455
rect 9268 8390 10955 8391
rect 8761 8278 10955 8390
rect 8761 8238 9079 8278
rect 8761 8174 8876 8238
rect 8940 8174 9079 8238
rect 8761 8081 9079 8174
rect 8761 8017 8877 8081
rect 8941 8017 9079 8081
rect 8761 7911 9079 8017
rect 8761 7847 8877 7911
rect 8941 7847 9079 7911
rect 8761 7759 9079 7847
rect 11053 8144 11246 8700
rect 11342 8144 11710 8700
rect 13069 8942 13228 8943
rect 13069 8932 13410 8942
rect 13069 8868 13345 8932
rect 13409 8868 13410 8932
rect 13069 8858 13410 8868
rect 13069 8615 13272 8858
rect 13470 8739 13530 9120
rect 13591 9896 13657 9986
rect 13591 9832 13592 9896
rect 13656 9832 13657 9896
rect 13591 9816 13657 9832
rect 13591 9752 13592 9816
rect 13656 9752 13657 9816
rect 13591 9736 13657 9752
rect 13591 9672 13592 9736
rect 13656 9672 13657 9736
rect 13591 9656 13657 9672
rect 13591 9592 13592 9656
rect 13656 9592 13657 9656
rect 13591 9576 13657 9592
rect 13591 9512 13592 9576
rect 13656 9512 13657 9576
rect 13591 9496 13657 9512
rect 13591 9432 13592 9496
rect 13656 9432 13657 9496
rect 13591 9416 13657 9432
rect 13591 9352 13592 9416
rect 13656 9352 13657 9416
rect 13591 9336 13657 9352
rect 13591 9272 13592 9336
rect 13656 9272 13657 9336
rect 13591 9256 13657 9272
rect 13591 9192 13592 9256
rect 13656 9192 13657 9256
rect 13591 9176 13657 9192
rect 13591 9112 13592 9176
rect 13656 9112 13657 9176
rect 13591 8958 13657 9112
rect 13717 9020 13777 10050
rect 13837 8958 13897 9990
rect 13957 9020 14017 10050
rect 14077 8958 14137 9990
rect 14197 9896 14263 9986
rect 14197 9832 14198 9896
rect 14262 9832 14263 9896
rect 14197 9816 14263 9832
rect 14197 9752 14198 9816
rect 14262 9752 14263 9816
rect 14197 9736 14263 9752
rect 14197 9672 14198 9736
rect 14262 9672 14263 9736
rect 14197 9656 14263 9672
rect 14197 9592 14198 9656
rect 14262 9592 14263 9656
rect 14197 9576 14263 9592
rect 14197 9512 14198 9576
rect 14262 9512 14263 9576
rect 14197 9496 14263 9512
rect 14197 9432 14198 9496
rect 14262 9432 14263 9496
rect 14197 9416 14263 9432
rect 14197 9352 14198 9416
rect 14262 9352 14263 9416
rect 14197 9336 14263 9352
rect 14197 9272 14198 9336
rect 14262 9272 14263 9336
rect 14197 9256 14263 9272
rect 14197 9192 14198 9256
rect 14262 9192 14263 9256
rect 14197 9176 14263 9192
rect 14197 9112 14198 9176
rect 14262 9112 14263 9176
rect 14197 8958 14263 9112
rect 13591 8956 14263 8958
rect 13591 8892 13695 8956
rect 13759 8892 13775 8956
rect 13839 8892 13855 8956
rect 13919 8892 13935 8956
rect 13999 8892 14015 8956
rect 14079 8892 14095 8956
rect 14159 8892 14263 8956
rect 13591 8890 14263 8892
rect 14325 9896 14391 9986
rect 14325 9832 14326 9896
rect 14390 9832 14391 9896
rect 14325 9816 14391 9832
rect 14325 9752 14326 9816
rect 14390 9752 14391 9816
rect 14325 9736 14391 9752
rect 14325 9672 14326 9736
rect 14390 9672 14391 9736
rect 14325 9656 14391 9672
rect 14325 9592 14326 9656
rect 14390 9592 14391 9656
rect 14325 9576 14391 9592
rect 14325 9512 14326 9576
rect 14390 9512 14391 9576
rect 14325 9496 14391 9512
rect 14325 9432 14326 9496
rect 14390 9432 14391 9496
rect 14325 9416 14391 9432
rect 14325 9352 14326 9416
rect 14390 9352 14391 9416
rect 14325 9336 14391 9352
rect 14325 9272 14326 9336
rect 14390 9272 14391 9336
rect 14325 9256 14391 9272
rect 14325 9192 14326 9256
rect 14390 9192 14391 9256
rect 14325 9176 14391 9192
rect 14325 9112 14326 9176
rect 14390 9112 14391 9176
rect 14325 8958 14391 9112
rect 14451 9020 14511 10050
rect 14571 8958 14631 9990
rect 14691 9020 14751 10050
rect 14811 8958 14871 9990
rect 14931 9896 14997 9986
rect 14931 9832 14932 9896
rect 14996 9832 14997 9896
rect 14931 9816 14997 9832
rect 14931 9752 14932 9816
rect 14996 9752 14997 9816
rect 14931 9736 14997 9752
rect 14931 9672 14932 9736
rect 14996 9672 14997 9736
rect 14931 9656 14997 9672
rect 14931 9592 14932 9656
rect 14996 9592 14997 9656
rect 14931 9576 14997 9592
rect 14931 9512 14932 9576
rect 14996 9512 14997 9576
rect 14931 9496 14997 9512
rect 14931 9432 14932 9496
rect 14996 9432 14997 9496
rect 14931 9416 14997 9432
rect 14931 9352 14932 9416
rect 14996 9352 14997 9416
rect 14931 9336 14997 9352
rect 14931 9272 14932 9336
rect 14996 9272 14997 9336
rect 14931 9256 14997 9272
rect 14931 9192 14932 9256
rect 14996 9192 14997 9256
rect 14931 9176 14997 9192
rect 14931 9112 14932 9176
rect 14996 9112 14997 9176
rect 14931 8958 14997 9112
rect 15057 8958 15117 9990
rect 15177 9020 15237 10050
rect 15297 8958 15357 9990
rect 15417 9020 15477 10050
rect 15537 9896 15603 9986
rect 15537 9832 15538 9896
rect 15602 9832 15603 9896
rect 15537 9816 15603 9832
rect 15537 9752 15538 9816
rect 15602 9752 15603 9816
rect 15537 9736 15603 9752
rect 15537 9672 15538 9736
rect 15602 9672 15603 9736
rect 15537 9656 15603 9672
rect 15537 9592 15538 9656
rect 15602 9592 15603 9656
rect 15537 9576 15603 9592
rect 15537 9512 15538 9576
rect 15602 9512 15603 9576
rect 15537 9496 15603 9512
rect 15537 9432 15538 9496
rect 15602 9432 15603 9496
rect 15537 9416 15603 9432
rect 15537 9352 15538 9416
rect 15602 9352 15603 9416
rect 15537 9336 15603 9352
rect 15537 9272 15538 9336
rect 15602 9272 15603 9336
rect 15537 9256 15603 9272
rect 15537 9192 15538 9256
rect 15602 9192 15603 9256
rect 15537 9176 15603 9192
rect 15537 9112 15538 9176
rect 15602 9112 15603 9176
rect 15537 8958 15603 9112
rect 14325 8956 15603 8958
rect 14325 8892 14429 8956
rect 14493 8892 14509 8956
rect 14573 8892 14589 8956
rect 14653 8892 14669 8956
rect 14733 8892 14749 8956
rect 14813 8892 14829 8956
rect 14893 8892 15035 8956
rect 15099 8892 15115 8956
rect 15179 8892 15195 8956
rect 15259 8892 15275 8956
rect 15339 8892 15355 8956
rect 15419 8892 15435 8956
rect 15499 8892 15603 8956
rect 14325 8890 15603 8892
rect 15663 9896 15729 9986
rect 15663 9832 15664 9896
rect 15728 9832 15729 9896
rect 15663 9816 15729 9832
rect 15663 9752 15664 9816
rect 15728 9752 15729 9816
rect 15663 9736 15729 9752
rect 15663 9672 15664 9736
rect 15728 9672 15729 9736
rect 15663 9656 15729 9672
rect 15663 9592 15664 9656
rect 15728 9592 15729 9656
rect 15663 9576 15729 9592
rect 15663 9512 15664 9576
rect 15728 9512 15729 9576
rect 15663 9496 15729 9512
rect 15663 9432 15664 9496
rect 15728 9432 15729 9496
rect 15663 9416 15729 9432
rect 15663 9352 15664 9416
rect 15728 9352 15729 9416
rect 15663 9336 15729 9352
rect 15663 9272 15664 9336
rect 15728 9272 15729 9336
rect 15663 9256 15729 9272
rect 15663 9192 15664 9256
rect 15728 9192 15729 9256
rect 15663 9176 15729 9192
rect 15663 9112 15664 9176
rect 15728 9112 15729 9176
rect 15663 8958 15729 9112
rect 15789 9020 15849 10050
rect 15909 8958 15969 9990
rect 16029 9020 16089 10050
rect 16149 8958 16209 9990
rect 16269 9896 16335 9986
rect 16269 9832 16270 9896
rect 16334 9832 16335 9896
rect 16269 9816 16335 9832
rect 16269 9752 16270 9816
rect 16334 9752 16335 9816
rect 16269 9736 16335 9752
rect 16269 9672 16270 9736
rect 16334 9672 16335 9736
rect 16269 9656 16335 9672
rect 16269 9592 16270 9656
rect 16334 9592 16335 9656
rect 16269 9576 16335 9592
rect 16269 9512 16270 9576
rect 16334 9512 16335 9576
rect 16269 9496 16335 9512
rect 16269 9432 16270 9496
rect 16334 9432 16335 9496
rect 16269 9416 16335 9432
rect 16269 9352 16270 9416
rect 16334 9352 16335 9416
rect 16269 9336 16335 9352
rect 16269 9272 16270 9336
rect 16334 9272 16335 9336
rect 16269 9256 16335 9272
rect 16269 9192 16270 9256
rect 16334 9192 16335 9256
rect 16269 9176 16335 9192
rect 16269 9112 16270 9176
rect 16334 9112 16335 9176
rect 16269 8958 16335 9112
rect 16395 8958 16455 9990
rect 16515 9020 16575 10050
rect 16635 8958 16695 9990
rect 16755 9020 16815 10050
rect 16875 9896 16941 9986
rect 16875 9832 16876 9896
rect 16940 9832 16941 9896
rect 16875 9816 16941 9832
rect 16875 9752 16876 9816
rect 16940 9752 16941 9816
rect 16875 9736 16941 9752
rect 16875 9672 16876 9736
rect 16940 9672 16941 9736
rect 16875 9656 16941 9672
rect 16875 9592 16876 9656
rect 16940 9592 16941 9656
rect 16875 9576 16941 9592
rect 16875 9512 16876 9576
rect 16940 9512 16941 9576
rect 16875 9496 16941 9512
rect 16875 9432 16876 9496
rect 16940 9432 16941 9496
rect 16875 9416 16941 9432
rect 16875 9352 16876 9416
rect 16940 9352 16941 9416
rect 16875 9336 16941 9352
rect 16875 9272 16876 9336
rect 16940 9272 16941 9336
rect 16875 9256 16941 9272
rect 16875 9192 16876 9256
rect 16940 9192 16941 9256
rect 16875 9176 16941 9192
rect 16875 9112 16876 9176
rect 16940 9112 16941 9176
rect 16875 8958 16941 9112
rect 17001 9020 17061 10050
rect 17121 8958 17181 9990
rect 17241 9020 17301 10050
rect 17361 8958 17421 9990
rect 17481 9896 17547 9986
rect 17481 9832 17482 9896
rect 17546 9832 17547 9896
rect 17481 9816 17547 9832
rect 17481 9752 17482 9816
rect 17546 9752 17547 9816
rect 17481 9736 17547 9752
rect 17481 9672 17482 9736
rect 17546 9672 17547 9736
rect 17481 9656 17547 9672
rect 17481 9592 17482 9656
rect 17546 9592 17547 9656
rect 17481 9576 17547 9592
rect 17481 9512 17482 9576
rect 17546 9512 17547 9576
rect 17481 9496 17547 9512
rect 17481 9432 17482 9496
rect 17546 9432 17547 9496
rect 17481 9416 17547 9432
rect 17481 9352 17482 9416
rect 17546 9352 17547 9416
rect 17481 9336 17547 9352
rect 17481 9272 17482 9336
rect 17546 9272 17547 9336
rect 17481 9256 17547 9272
rect 17481 9192 17482 9256
rect 17546 9192 17547 9256
rect 17481 9176 17547 9192
rect 17481 9112 17482 9176
rect 17546 9112 17547 9176
rect 17481 8958 17547 9112
rect 17607 8958 17667 9990
rect 17727 9020 17787 10050
rect 17847 8958 17907 9990
rect 17967 9020 18027 10050
rect 18087 9896 18153 9986
rect 18087 9832 18088 9896
rect 18152 9832 18153 9896
rect 18087 9816 18153 9832
rect 18087 9752 18088 9816
rect 18152 9752 18153 9816
rect 18087 9736 18153 9752
rect 18087 9672 18088 9736
rect 18152 9672 18153 9736
rect 18087 9656 18153 9672
rect 18087 9592 18088 9656
rect 18152 9592 18153 9656
rect 18087 9576 18153 9592
rect 18087 9512 18088 9576
rect 18152 9512 18153 9576
rect 18087 9496 18153 9512
rect 18087 9432 18088 9496
rect 18152 9432 18153 9496
rect 18087 9416 18153 9432
rect 18087 9352 18088 9416
rect 18152 9352 18153 9416
rect 18087 9336 18153 9352
rect 18087 9272 18088 9336
rect 18152 9272 18153 9336
rect 18087 9256 18153 9272
rect 18087 9192 18088 9256
rect 18152 9192 18153 9256
rect 18087 9176 18153 9192
rect 18087 9112 18088 9176
rect 18152 9112 18153 9176
rect 18087 8958 18153 9112
rect 15663 8956 18153 8958
rect 15663 8892 15767 8956
rect 15831 8892 15847 8956
rect 15911 8892 15927 8956
rect 15991 8892 16007 8956
rect 16071 8892 16087 8956
rect 16151 8892 16167 8956
rect 16231 8892 16373 8956
rect 16437 8892 16453 8956
rect 16517 8892 16533 8956
rect 16597 8892 16613 8956
rect 16677 8892 16693 8956
rect 16757 8892 16773 8956
rect 16837 8892 16979 8956
rect 17043 8892 17059 8956
rect 17123 8892 17139 8956
rect 17203 8892 17219 8956
rect 17283 8892 17299 8956
rect 17363 8892 17379 8956
rect 17443 8892 17585 8956
rect 17649 8892 17665 8956
rect 17729 8892 17745 8956
rect 17809 8892 17825 8956
rect 17889 8892 17905 8956
rect 17969 8892 17985 8956
rect 18049 8892 18153 8956
rect 15663 8890 18153 8892
rect 18213 9896 18279 9986
rect 18213 9832 18214 9896
rect 18278 9832 18279 9896
rect 18213 9816 18279 9832
rect 18213 9752 18214 9816
rect 18278 9752 18279 9816
rect 18213 9736 18279 9752
rect 18213 9672 18214 9736
rect 18278 9672 18279 9736
rect 18213 9656 18279 9672
rect 18213 9592 18214 9656
rect 18278 9592 18279 9656
rect 18213 9576 18279 9592
rect 18213 9512 18214 9576
rect 18278 9512 18279 9576
rect 18213 9496 18279 9512
rect 18213 9432 18214 9496
rect 18278 9432 18279 9496
rect 18213 9416 18279 9432
rect 18213 9352 18214 9416
rect 18278 9352 18279 9416
rect 18213 9336 18279 9352
rect 18213 9272 18214 9336
rect 18278 9272 18279 9336
rect 18213 9256 18279 9272
rect 18213 9192 18214 9256
rect 18278 9192 18279 9256
rect 18213 9176 18279 9192
rect 18213 9112 18214 9176
rect 18278 9112 18279 9176
rect 18213 8958 18279 9112
rect 18339 8958 18399 9990
rect 18459 9020 18519 10050
rect 18579 8958 18639 9990
rect 18699 9020 18759 10050
rect 19148 10045 19273 10051
rect 18819 9896 18885 9986
rect 18819 9832 18820 9896
rect 18884 9832 18885 9896
rect 18819 9816 18885 9832
rect 18819 9752 18820 9816
rect 18884 9752 18885 9816
rect 18819 9736 18885 9752
rect 18819 9672 18820 9736
rect 18884 9672 18885 9736
rect 18819 9656 18885 9672
rect 18819 9592 18820 9656
rect 18884 9592 18885 9656
rect 18819 9576 18885 9592
rect 18819 9512 18820 9576
rect 18884 9512 18885 9576
rect 18819 9496 18885 9512
rect 18819 9432 18820 9496
rect 18884 9432 18885 9496
rect 18819 9416 18885 9432
rect 18819 9352 18820 9416
rect 18884 9352 18885 9416
rect 18819 9336 18885 9352
rect 18819 9272 18820 9336
rect 18884 9272 18885 9336
rect 18819 9256 18885 9272
rect 18819 9192 18820 9256
rect 18884 9192 18885 9256
rect 18819 9176 18885 9192
rect 18819 9112 18820 9176
rect 18884 9112 18885 9176
rect 18819 8958 18885 9112
rect 18213 8956 18885 8958
rect 18213 8892 18317 8956
rect 18381 8892 18397 8956
rect 18461 8892 18477 8956
rect 18541 8892 18557 8956
rect 18621 8892 18637 8956
rect 18701 8892 18717 8956
rect 18781 8892 18885 8956
rect 18213 8890 18885 8892
rect 13332 8729 13530 8739
rect 13332 8665 13345 8729
rect 13409 8665 13530 8729
rect 18564 8711 19236 8713
rect 13332 8655 13530 8665
rect 13590 8708 18504 8710
rect 11782 8512 13272 8615
rect 11782 8448 12719 8512
rect 12783 8448 13093 8512
rect 13157 8480 13272 8512
rect 13590 8644 13694 8708
rect 13758 8644 13774 8708
rect 13838 8644 13854 8708
rect 13918 8644 13934 8708
rect 13998 8644 14014 8708
rect 14078 8644 14094 8708
rect 14158 8644 14300 8708
rect 14364 8644 14380 8708
rect 14444 8644 14460 8708
rect 14524 8644 14540 8708
rect 14604 8644 14620 8708
rect 14684 8644 14700 8708
rect 14764 8644 14906 8708
rect 14970 8644 14986 8708
rect 15050 8644 15066 8708
rect 15130 8644 15146 8708
rect 15210 8644 15226 8708
rect 15290 8644 15306 8708
rect 15370 8644 15512 8708
rect 15576 8644 15592 8708
rect 15656 8644 15672 8708
rect 15736 8644 15752 8708
rect 15816 8644 15832 8708
rect 15896 8644 15912 8708
rect 15976 8644 16118 8708
rect 16182 8644 16198 8708
rect 16262 8644 16278 8708
rect 16342 8644 16358 8708
rect 16422 8644 16438 8708
rect 16502 8644 16518 8708
rect 16582 8644 16724 8708
rect 16788 8644 16804 8708
rect 16868 8644 16884 8708
rect 16948 8644 16964 8708
rect 17028 8644 17044 8708
rect 17108 8644 17124 8708
rect 17188 8644 17330 8708
rect 17394 8644 17410 8708
rect 17474 8644 17490 8708
rect 17554 8644 17570 8708
rect 17634 8644 17650 8708
rect 17714 8644 17730 8708
rect 17794 8644 17936 8708
rect 18000 8644 18016 8708
rect 18080 8644 18096 8708
rect 18160 8644 18176 8708
rect 18240 8644 18256 8708
rect 18320 8644 18336 8708
rect 18400 8644 18504 8708
rect 13590 8642 18504 8644
rect 13590 8488 13656 8642
rect 13157 8468 13530 8480
rect 13157 8448 13433 8468
rect 11782 8442 13433 8448
rect 11782 8419 12224 8442
rect 11053 7909 11710 8144
rect 11786 8378 12224 8419
rect 12288 8404 13433 8442
rect 13497 8404 13530 8468
rect 12288 8378 13530 8404
rect 11786 8369 13530 8378
rect 11786 8305 12581 8369
rect 12645 8366 13530 8369
rect 12645 8305 12765 8366
rect 11786 8302 12765 8305
rect 12829 8360 13530 8366
rect 12829 8302 13067 8360
rect 11786 8296 13067 8302
rect 13131 8296 13530 8360
rect 11786 8226 13530 8296
rect 11786 8162 13351 8226
rect 13415 8162 13530 8226
rect 11786 8109 13530 8162
rect 12825 8069 13530 8109
rect 12825 8005 13350 8069
rect 13414 8005 13530 8069
rect 12825 7988 13530 8005
rect 12825 7935 13133 7988
rect 11053 7771 12582 7909
rect 8761 7695 8876 7759
rect 8940 7695 9079 7759
rect 8761 7615 9079 7695
rect 10054 7744 12582 7771
rect 10054 7740 12214 7744
rect 10054 7731 11960 7740
rect 10054 7729 11029 7731
rect 10054 7665 10140 7729
rect 10204 7665 10388 7729
rect 10452 7665 10685 7729
rect 10749 7667 11029 7729
rect 11093 7667 11348 7731
rect 11412 7676 11960 7731
rect 12024 7680 12214 7740
rect 12278 7680 12582 7744
rect 12024 7676 12582 7680
rect 11412 7667 12582 7676
rect 10749 7665 12582 7667
rect 10054 7656 12582 7665
rect 8761 7562 8871 7615
rect 3623 7560 8871 7562
rect 3623 7499 3891 7560
rect 3126 7496 3891 7499
rect 3955 7496 3971 7560
rect 4035 7496 4051 7560
rect 4115 7496 4131 7560
rect 4195 7496 4211 7560
rect 4275 7496 4291 7560
rect 4355 7496 4497 7560
rect 4561 7496 4577 7560
rect 4641 7496 4657 7560
rect 4721 7496 4737 7560
rect 4801 7496 4817 7560
rect 4881 7496 4897 7560
rect 4961 7496 5103 7560
rect 5167 7496 5183 7560
rect 5247 7496 5263 7560
rect 5327 7496 5343 7560
rect 5407 7496 5423 7560
rect 5487 7496 5503 7560
rect 5567 7496 5709 7560
rect 5773 7496 5789 7560
rect 5853 7496 5869 7560
rect 5933 7496 5949 7560
rect 6013 7496 6029 7560
rect 6093 7496 6109 7560
rect 6173 7496 6315 7560
rect 6379 7496 6395 7560
rect 6459 7496 6475 7560
rect 6539 7496 6555 7560
rect 6619 7496 6635 7560
rect 6699 7496 6715 7560
rect 6779 7496 6921 7560
rect 6985 7496 7001 7560
rect 7065 7496 7081 7560
rect 7145 7496 7161 7560
rect 7225 7496 7241 7560
rect 7305 7496 7321 7560
rect 7385 7496 7527 7560
rect 7591 7496 7607 7560
rect 7671 7496 7687 7560
rect 7751 7496 7767 7560
rect 7831 7496 7847 7560
rect 7911 7496 7927 7560
rect 7991 7496 8133 7560
rect 8197 7496 8213 7560
rect 8277 7496 8293 7560
rect 8357 7496 8373 7560
rect 8437 7496 8453 7560
rect 8517 7496 8533 7560
rect 8597 7551 8871 7560
rect 8935 7551 9079 7615
rect 8597 7496 9079 7551
rect 3126 7489 9079 7496
rect 2064 7484 9079 7489
rect 3031 7479 3157 7484
rect 10055 2874 10580 7656
rect 10655 7655 10781 7656
rect 11383 7598 12582 7656
rect 11383 7595 12222 7598
rect 11383 7531 11970 7595
rect 12034 7534 12222 7595
rect 12286 7534 12582 7598
rect 12825 7871 12934 7935
rect 12998 7871 13133 7935
rect 12825 7715 13133 7871
rect 12825 7651 12926 7715
rect 12990 7651 13133 7715
rect 12825 7558 13133 7651
rect 13211 7899 13530 7988
rect 13211 7835 13350 7899
rect 13414 7835 13530 7899
rect 13211 7747 13530 7835
rect 13211 7683 13351 7747
rect 13415 7683 13530 7747
rect 13211 7603 13530 7683
rect 13590 8424 13591 8488
rect 13655 8424 13656 8488
rect 13590 8408 13656 8424
rect 13590 8344 13591 8408
rect 13655 8344 13656 8408
rect 13590 8328 13656 8344
rect 13590 8264 13591 8328
rect 13655 8264 13656 8328
rect 13590 8248 13656 8264
rect 13590 8184 13591 8248
rect 13655 8184 13656 8248
rect 13590 8168 13656 8184
rect 13590 8104 13591 8168
rect 13655 8104 13656 8168
rect 13590 8088 13656 8104
rect 13590 8024 13591 8088
rect 13655 8024 13656 8088
rect 13590 8008 13656 8024
rect 13590 7944 13591 8008
rect 13655 7944 13656 8008
rect 13590 7928 13656 7944
rect 13590 7864 13591 7928
rect 13655 7864 13656 7928
rect 13590 7848 13656 7864
rect 13590 7784 13591 7848
rect 13655 7784 13656 7848
rect 13590 7768 13656 7784
rect 13590 7704 13591 7768
rect 13655 7704 13656 7768
rect 13590 7614 13656 7704
rect 13211 7558 13356 7603
rect 12825 7540 13356 7558
rect 12034 7531 12582 7534
rect 11383 7441 12582 7531
rect 12824 7539 13356 7540
rect 13420 7550 13530 7603
rect 13716 7550 13776 8580
rect 13836 7610 13896 8642
rect 13956 7550 14016 8580
rect 14076 7610 14136 8642
rect 14196 8488 14262 8642
rect 14196 8424 14197 8488
rect 14261 8424 14262 8488
rect 14196 8408 14262 8424
rect 14196 8344 14197 8408
rect 14261 8344 14262 8408
rect 14196 8328 14262 8344
rect 14196 8264 14197 8328
rect 14261 8264 14262 8328
rect 14196 8248 14262 8264
rect 14196 8184 14197 8248
rect 14261 8184 14262 8248
rect 14196 8168 14262 8184
rect 14196 8104 14197 8168
rect 14261 8104 14262 8168
rect 14196 8088 14262 8104
rect 14196 8024 14197 8088
rect 14261 8024 14262 8088
rect 14196 8008 14262 8024
rect 14196 7944 14197 8008
rect 14261 7944 14262 8008
rect 14196 7928 14262 7944
rect 14196 7864 14197 7928
rect 14261 7864 14262 7928
rect 14196 7848 14262 7864
rect 14196 7784 14197 7848
rect 14261 7784 14262 7848
rect 14196 7768 14262 7784
rect 14196 7704 14197 7768
rect 14261 7704 14262 7768
rect 14196 7614 14262 7704
rect 14322 7610 14382 8642
rect 14442 7550 14502 8580
rect 14562 7610 14622 8642
rect 14682 7550 14742 8580
rect 14802 8488 14868 8642
rect 14802 8424 14803 8488
rect 14867 8424 14868 8488
rect 14802 8408 14868 8424
rect 14802 8344 14803 8408
rect 14867 8344 14868 8408
rect 14802 8328 14868 8344
rect 14802 8264 14803 8328
rect 14867 8264 14868 8328
rect 14802 8248 14868 8264
rect 14802 8184 14803 8248
rect 14867 8184 14868 8248
rect 14802 8168 14868 8184
rect 14802 8104 14803 8168
rect 14867 8104 14868 8168
rect 14802 8088 14868 8104
rect 14802 8024 14803 8088
rect 14867 8024 14868 8088
rect 14802 8008 14868 8024
rect 14802 7944 14803 8008
rect 14867 7944 14868 8008
rect 14802 7928 14868 7944
rect 14802 7864 14803 7928
rect 14867 7864 14868 7928
rect 14802 7848 14868 7864
rect 14802 7784 14803 7848
rect 14867 7784 14868 7848
rect 14802 7768 14868 7784
rect 14802 7704 14803 7768
rect 14867 7704 14868 7768
rect 14802 7614 14868 7704
rect 14928 7550 14988 8580
rect 15048 7610 15108 8642
rect 15168 7550 15228 8580
rect 15288 7610 15348 8642
rect 15408 8488 15474 8642
rect 15408 8424 15409 8488
rect 15473 8424 15474 8488
rect 15408 8408 15474 8424
rect 15408 8344 15409 8408
rect 15473 8344 15474 8408
rect 15408 8328 15474 8344
rect 15408 8264 15409 8328
rect 15473 8264 15474 8328
rect 15408 8248 15474 8264
rect 15408 8184 15409 8248
rect 15473 8184 15474 8248
rect 15408 8168 15474 8184
rect 15408 8104 15409 8168
rect 15473 8104 15474 8168
rect 15408 8088 15474 8104
rect 15408 8024 15409 8088
rect 15473 8024 15474 8088
rect 15408 8008 15474 8024
rect 15408 7944 15409 8008
rect 15473 7944 15474 8008
rect 15408 7928 15474 7944
rect 15408 7864 15409 7928
rect 15473 7864 15474 7928
rect 15408 7848 15474 7864
rect 15408 7784 15409 7848
rect 15473 7784 15474 7848
rect 15408 7768 15474 7784
rect 15408 7704 15409 7768
rect 15473 7704 15474 7768
rect 15408 7614 15474 7704
rect 15534 7610 15594 8642
rect 15654 7550 15714 8580
rect 15774 7610 15834 8642
rect 15894 7550 15954 8580
rect 16014 8488 16080 8642
rect 16014 8424 16015 8488
rect 16079 8424 16080 8488
rect 16014 8408 16080 8424
rect 16014 8344 16015 8408
rect 16079 8344 16080 8408
rect 16014 8328 16080 8344
rect 16014 8264 16015 8328
rect 16079 8264 16080 8328
rect 16014 8248 16080 8264
rect 16014 8184 16015 8248
rect 16079 8184 16080 8248
rect 16014 8168 16080 8184
rect 16014 8104 16015 8168
rect 16079 8104 16080 8168
rect 16014 8088 16080 8104
rect 16014 8024 16015 8088
rect 16079 8024 16080 8088
rect 16014 8008 16080 8024
rect 16014 7944 16015 8008
rect 16079 7944 16080 8008
rect 16014 7928 16080 7944
rect 16014 7864 16015 7928
rect 16079 7864 16080 7928
rect 16014 7848 16080 7864
rect 16014 7784 16015 7848
rect 16079 7784 16080 7848
rect 16014 7768 16080 7784
rect 16014 7704 16015 7768
rect 16079 7704 16080 7768
rect 16014 7614 16080 7704
rect 16140 7550 16200 8580
rect 16260 7610 16320 8642
rect 16380 7550 16440 8580
rect 16500 7610 16560 8642
rect 16620 8488 16686 8642
rect 16620 8424 16621 8488
rect 16685 8424 16686 8488
rect 16620 8408 16686 8424
rect 16620 8344 16621 8408
rect 16685 8344 16686 8408
rect 16620 8328 16686 8344
rect 16620 8264 16621 8328
rect 16685 8264 16686 8328
rect 16620 8248 16686 8264
rect 16620 8184 16621 8248
rect 16685 8184 16686 8248
rect 16620 8168 16686 8184
rect 16620 8104 16621 8168
rect 16685 8104 16686 8168
rect 16620 8088 16686 8104
rect 16620 8024 16621 8088
rect 16685 8024 16686 8088
rect 16620 8008 16686 8024
rect 16620 7944 16621 8008
rect 16685 7944 16686 8008
rect 16620 7928 16686 7944
rect 16620 7864 16621 7928
rect 16685 7864 16686 7928
rect 16620 7848 16686 7864
rect 16620 7784 16621 7848
rect 16685 7784 16686 7848
rect 16620 7768 16686 7784
rect 16620 7704 16621 7768
rect 16685 7704 16686 7768
rect 16620 7614 16686 7704
rect 16746 7610 16806 8642
rect 16866 7550 16926 8580
rect 16986 7610 17046 8642
rect 17106 7550 17166 8580
rect 17226 8488 17292 8642
rect 17226 8424 17227 8488
rect 17291 8424 17292 8488
rect 17226 8408 17292 8424
rect 17226 8344 17227 8408
rect 17291 8344 17292 8408
rect 17226 8328 17292 8344
rect 17226 8264 17227 8328
rect 17291 8264 17292 8328
rect 17226 8248 17292 8264
rect 17226 8184 17227 8248
rect 17291 8184 17292 8248
rect 17226 8168 17292 8184
rect 17226 8104 17227 8168
rect 17291 8104 17292 8168
rect 17226 8088 17292 8104
rect 17226 8024 17227 8088
rect 17291 8024 17292 8088
rect 17226 8008 17292 8024
rect 17226 7944 17227 8008
rect 17291 7944 17292 8008
rect 17226 7928 17292 7944
rect 17226 7864 17227 7928
rect 17291 7864 17292 7928
rect 17226 7848 17292 7864
rect 17226 7784 17227 7848
rect 17291 7784 17292 7848
rect 17226 7768 17292 7784
rect 17226 7704 17227 7768
rect 17291 7704 17292 7768
rect 17226 7614 17292 7704
rect 17352 7550 17412 8580
rect 17472 7610 17532 8642
rect 17592 7550 17652 8580
rect 17712 7610 17772 8642
rect 17832 8488 17898 8642
rect 17832 8424 17833 8488
rect 17897 8424 17898 8488
rect 17832 8408 17898 8424
rect 17832 8344 17833 8408
rect 17897 8344 17898 8408
rect 17832 8328 17898 8344
rect 17832 8264 17833 8328
rect 17897 8264 17898 8328
rect 17832 8248 17898 8264
rect 17832 8184 17833 8248
rect 17897 8184 17898 8248
rect 17832 8168 17898 8184
rect 17832 8104 17833 8168
rect 17897 8104 17898 8168
rect 17832 8088 17898 8104
rect 17832 8024 17833 8088
rect 17897 8024 17898 8088
rect 17832 8008 17898 8024
rect 17832 7944 17833 8008
rect 17897 7944 17898 8008
rect 17832 7928 17898 7944
rect 17832 7864 17833 7928
rect 17897 7864 17898 7928
rect 17832 7848 17898 7864
rect 17832 7784 17833 7848
rect 17897 7784 17898 7848
rect 17832 7768 17898 7784
rect 17832 7704 17833 7768
rect 17897 7704 17898 7768
rect 17832 7614 17898 7704
rect 17958 7610 18018 8642
rect 18078 7550 18138 8580
rect 18198 7610 18258 8642
rect 18318 7550 18378 8580
rect 18438 8488 18504 8642
rect 18438 8424 18439 8488
rect 18503 8424 18504 8488
rect 18438 8408 18504 8424
rect 18438 8344 18439 8408
rect 18503 8344 18504 8408
rect 18438 8328 18504 8344
rect 18438 8264 18439 8328
rect 18503 8264 18504 8328
rect 18438 8248 18504 8264
rect 18438 8184 18439 8248
rect 18503 8184 18504 8248
rect 18438 8168 18504 8184
rect 18438 8104 18439 8168
rect 18503 8104 18504 8168
rect 18438 8088 18504 8104
rect 18438 8024 18439 8088
rect 18503 8024 18504 8088
rect 18438 8008 18504 8024
rect 18438 7944 18439 8008
rect 18503 7944 18504 8008
rect 18438 7928 18504 7944
rect 18438 7864 18439 7928
rect 18503 7864 18504 7928
rect 18438 7848 18504 7864
rect 18438 7784 18439 7848
rect 18503 7784 18504 7848
rect 18438 7768 18504 7784
rect 18438 7704 18439 7768
rect 18503 7704 18504 7768
rect 18438 7614 18504 7704
rect 18564 8647 18668 8711
rect 18732 8647 18748 8711
rect 18812 8647 18828 8711
rect 18892 8647 18908 8711
rect 18972 8647 18988 8711
rect 19052 8647 19068 8711
rect 19132 8647 19236 8711
rect 19457 8692 19833 10051
rect 19921 10052 20484 10111
rect 20548 10052 20564 10116
rect 20628 10052 20644 10116
rect 20708 10052 20724 10116
rect 20788 10052 21218 10116
rect 21282 10052 21298 10116
rect 21362 10052 21378 10116
rect 21442 10052 21458 10116
rect 21522 10052 21824 10116
rect 21888 10052 21904 10116
rect 21968 10052 21984 10116
rect 22048 10052 22064 10116
rect 22128 10052 22556 10116
rect 22620 10052 22636 10116
rect 22700 10052 22716 10116
rect 22780 10052 22796 10116
rect 22860 10052 23162 10116
rect 23226 10052 23242 10116
rect 23306 10052 23322 10116
rect 23386 10052 23402 10116
rect 23466 10052 23768 10116
rect 23832 10052 23848 10116
rect 23912 10052 23928 10116
rect 23992 10052 24008 10116
rect 24072 10052 24374 10116
rect 24438 10052 24454 10116
rect 24518 10052 24534 10116
rect 24598 10052 24614 10116
rect 24678 10052 25106 10116
rect 25170 10052 25186 10116
rect 25250 10052 25266 10116
rect 25330 10052 25346 10116
rect 25410 10055 25888 10116
rect 25952 10055 26676 10119
rect 25410 10052 26676 10055
rect 19921 10051 26676 10052
rect 19921 9194 20239 10051
rect 20300 10050 20972 10051
rect 21034 10050 22312 10051
rect 22372 10050 24862 10051
rect 24922 10050 25594 10051
rect 19921 9130 20145 9194
rect 20209 9130 20239 9194
rect 19921 9120 20239 9130
rect 19921 8932 20119 8942
rect 19921 8868 20054 8932
rect 20118 8868 20119 8932
rect 19921 8858 20119 8868
rect 18564 8645 19236 8647
rect 18564 8491 18630 8645
rect 18564 8427 18565 8491
rect 18629 8427 18630 8491
rect 18564 8411 18630 8427
rect 18564 8347 18565 8411
rect 18629 8347 18630 8411
rect 18564 8331 18630 8347
rect 18564 8267 18565 8331
rect 18629 8267 18630 8331
rect 18564 8251 18630 8267
rect 18564 8187 18565 8251
rect 18629 8187 18630 8251
rect 18564 8171 18630 8187
rect 18564 8107 18565 8171
rect 18629 8107 18630 8171
rect 18564 8091 18630 8107
rect 18564 8027 18565 8091
rect 18629 8027 18630 8091
rect 18564 8011 18630 8027
rect 18564 7947 18565 8011
rect 18629 7947 18630 8011
rect 18564 7931 18630 7947
rect 18564 7867 18565 7931
rect 18629 7867 18630 7931
rect 18564 7851 18630 7867
rect 18564 7787 18565 7851
rect 18629 7787 18630 7851
rect 18564 7771 18630 7787
rect 18564 7707 18565 7771
rect 18629 7707 18630 7771
rect 18564 7617 18630 7707
rect 18690 7613 18750 8645
rect 18810 7553 18870 8583
rect 18930 7613 18990 8645
rect 19050 7553 19110 8583
rect 19170 8491 19236 8645
rect 19458 8628 19501 8692
rect 19565 8628 19644 8692
rect 19708 8628 19764 8692
rect 19828 8628 19835 8692
rect 19458 8613 19835 8628
rect 19170 8427 19171 8491
rect 19235 8427 19236 8491
rect 19170 8411 19236 8427
rect 19170 8347 19171 8411
rect 19235 8347 19236 8411
rect 19170 8331 19236 8347
rect 19170 8267 19171 8331
rect 19235 8267 19236 8331
rect 19170 8251 19236 8267
rect 19170 8187 19171 8251
rect 19235 8187 19236 8251
rect 19170 8171 19236 8187
rect 19170 8107 19171 8171
rect 19235 8107 19236 8171
rect 19921 8480 19981 8858
rect 20179 8739 20239 9120
rect 20300 9896 20366 9986
rect 20300 9832 20301 9896
rect 20365 9832 20366 9896
rect 20300 9816 20366 9832
rect 20300 9752 20301 9816
rect 20365 9752 20366 9816
rect 20300 9736 20366 9752
rect 20300 9672 20301 9736
rect 20365 9672 20366 9736
rect 20300 9656 20366 9672
rect 20300 9592 20301 9656
rect 20365 9592 20366 9656
rect 20300 9576 20366 9592
rect 20300 9512 20301 9576
rect 20365 9512 20366 9576
rect 20300 9496 20366 9512
rect 20300 9432 20301 9496
rect 20365 9432 20366 9496
rect 20300 9416 20366 9432
rect 20300 9352 20301 9416
rect 20365 9352 20366 9416
rect 20300 9336 20366 9352
rect 20300 9272 20301 9336
rect 20365 9272 20366 9336
rect 20300 9256 20366 9272
rect 20300 9192 20301 9256
rect 20365 9192 20366 9256
rect 20300 9176 20366 9192
rect 20300 9112 20301 9176
rect 20365 9112 20366 9176
rect 20300 8958 20366 9112
rect 20426 9020 20486 10050
rect 20546 8958 20606 9990
rect 20666 9020 20726 10050
rect 20786 8958 20846 9990
rect 20906 9896 20972 9986
rect 20906 9832 20907 9896
rect 20971 9832 20972 9896
rect 20906 9816 20972 9832
rect 20906 9752 20907 9816
rect 20971 9752 20972 9816
rect 20906 9736 20972 9752
rect 20906 9672 20907 9736
rect 20971 9672 20972 9736
rect 20906 9656 20972 9672
rect 20906 9592 20907 9656
rect 20971 9592 20972 9656
rect 20906 9576 20972 9592
rect 20906 9512 20907 9576
rect 20971 9512 20972 9576
rect 20906 9496 20972 9512
rect 20906 9432 20907 9496
rect 20971 9432 20972 9496
rect 20906 9416 20972 9432
rect 20906 9352 20907 9416
rect 20971 9352 20972 9416
rect 20906 9336 20972 9352
rect 20906 9272 20907 9336
rect 20971 9272 20972 9336
rect 20906 9256 20972 9272
rect 20906 9192 20907 9256
rect 20971 9192 20972 9256
rect 20906 9176 20972 9192
rect 20906 9112 20907 9176
rect 20971 9112 20972 9176
rect 20906 8958 20972 9112
rect 20300 8956 20972 8958
rect 20300 8892 20404 8956
rect 20468 8892 20484 8956
rect 20548 8892 20564 8956
rect 20628 8892 20644 8956
rect 20708 8892 20724 8956
rect 20788 8892 20804 8956
rect 20868 8892 20972 8956
rect 20300 8890 20972 8892
rect 21034 9896 21100 9986
rect 21034 9832 21035 9896
rect 21099 9832 21100 9896
rect 21034 9816 21100 9832
rect 21034 9752 21035 9816
rect 21099 9752 21100 9816
rect 21034 9736 21100 9752
rect 21034 9672 21035 9736
rect 21099 9672 21100 9736
rect 21034 9656 21100 9672
rect 21034 9592 21035 9656
rect 21099 9592 21100 9656
rect 21034 9576 21100 9592
rect 21034 9512 21035 9576
rect 21099 9512 21100 9576
rect 21034 9496 21100 9512
rect 21034 9432 21035 9496
rect 21099 9432 21100 9496
rect 21034 9416 21100 9432
rect 21034 9352 21035 9416
rect 21099 9352 21100 9416
rect 21034 9336 21100 9352
rect 21034 9272 21035 9336
rect 21099 9272 21100 9336
rect 21034 9256 21100 9272
rect 21034 9192 21035 9256
rect 21099 9192 21100 9256
rect 21034 9176 21100 9192
rect 21034 9112 21035 9176
rect 21099 9112 21100 9176
rect 21034 8958 21100 9112
rect 21160 9020 21220 10050
rect 21280 8958 21340 9990
rect 21400 9020 21460 10050
rect 21520 8958 21580 9990
rect 21640 9896 21706 9986
rect 21640 9832 21641 9896
rect 21705 9832 21706 9896
rect 21640 9816 21706 9832
rect 21640 9752 21641 9816
rect 21705 9752 21706 9816
rect 21640 9736 21706 9752
rect 21640 9672 21641 9736
rect 21705 9672 21706 9736
rect 21640 9656 21706 9672
rect 21640 9592 21641 9656
rect 21705 9592 21706 9656
rect 21640 9576 21706 9592
rect 21640 9512 21641 9576
rect 21705 9512 21706 9576
rect 21640 9496 21706 9512
rect 21640 9432 21641 9496
rect 21705 9432 21706 9496
rect 21640 9416 21706 9432
rect 21640 9352 21641 9416
rect 21705 9352 21706 9416
rect 21640 9336 21706 9352
rect 21640 9272 21641 9336
rect 21705 9272 21706 9336
rect 21640 9256 21706 9272
rect 21640 9192 21641 9256
rect 21705 9192 21706 9256
rect 21640 9176 21706 9192
rect 21640 9112 21641 9176
rect 21705 9112 21706 9176
rect 21640 8958 21706 9112
rect 21766 8958 21826 9990
rect 21886 9020 21946 10050
rect 22006 8958 22066 9990
rect 22126 9020 22186 10050
rect 22246 9896 22312 9986
rect 22246 9832 22247 9896
rect 22311 9832 22312 9896
rect 22246 9816 22312 9832
rect 22246 9752 22247 9816
rect 22311 9752 22312 9816
rect 22246 9736 22312 9752
rect 22246 9672 22247 9736
rect 22311 9672 22312 9736
rect 22246 9656 22312 9672
rect 22246 9592 22247 9656
rect 22311 9592 22312 9656
rect 22246 9576 22312 9592
rect 22246 9512 22247 9576
rect 22311 9512 22312 9576
rect 22246 9496 22312 9512
rect 22246 9432 22247 9496
rect 22311 9432 22312 9496
rect 22246 9416 22312 9432
rect 22246 9352 22247 9416
rect 22311 9352 22312 9416
rect 22246 9336 22312 9352
rect 22246 9272 22247 9336
rect 22311 9272 22312 9336
rect 22246 9256 22312 9272
rect 22246 9192 22247 9256
rect 22311 9192 22312 9256
rect 22246 9176 22312 9192
rect 22246 9112 22247 9176
rect 22311 9112 22312 9176
rect 22246 8958 22312 9112
rect 21034 8956 22312 8958
rect 21034 8892 21138 8956
rect 21202 8892 21218 8956
rect 21282 8892 21298 8956
rect 21362 8892 21378 8956
rect 21442 8892 21458 8956
rect 21522 8892 21538 8956
rect 21602 8892 21744 8956
rect 21808 8892 21824 8956
rect 21888 8892 21904 8956
rect 21968 8892 21984 8956
rect 22048 8892 22064 8956
rect 22128 8892 22144 8956
rect 22208 8892 22312 8956
rect 21034 8890 22312 8892
rect 22372 9896 22438 9986
rect 22372 9832 22373 9896
rect 22437 9832 22438 9896
rect 22372 9816 22438 9832
rect 22372 9752 22373 9816
rect 22437 9752 22438 9816
rect 22372 9736 22438 9752
rect 22372 9672 22373 9736
rect 22437 9672 22438 9736
rect 22372 9656 22438 9672
rect 22372 9592 22373 9656
rect 22437 9592 22438 9656
rect 22372 9576 22438 9592
rect 22372 9512 22373 9576
rect 22437 9512 22438 9576
rect 22372 9496 22438 9512
rect 22372 9432 22373 9496
rect 22437 9432 22438 9496
rect 22372 9416 22438 9432
rect 22372 9352 22373 9416
rect 22437 9352 22438 9416
rect 22372 9336 22438 9352
rect 22372 9272 22373 9336
rect 22437 9272 22438 9336
rect 22372 9256 22438 9272
rect 22372 9192 22373 9256
rect 22437 9192 22438 9256
rect 22372 9176 22438 9192
rect 22372 9112 22373 9176
rect 22437 9112 22438 9176
rect 22372 8958 22438 9112
rect 22498 9020 22558 10050
rect 22618 8958 22678 9990
rect 22738 9020 22798 10050
rect 22858 8958 22918 9990
rect 22978 9896 23044 9986
rect 22978 9832 22979 9896
rect 23043 9832 23044 9896
rect 22978 9816 23044 9832
rect 22978 9752 22979 9816
rect 23043 9752 23044 9816
rect 22978 9736 23044 9752
rect 22978 9672 22979 9736
rect 23043 9672 23044 9736
rect 22978 9656 23044 9672
rect 22978 9592 22979 9656
rect 23043 9592 23044 9656
rect 22978 9576 23044 9592
rect 22978 9512 22979 9576
rect 23043 9512 23044 9576
rect 22978 9496 23044 9512
rect 22978 9432 22979 9496
rect 23043 9432 23044 9496
rect 22978 9416 23044 9432
rect 22978 9352 22979 9416
rect 23043 9352 23044 9416
rect 22978 9336 23044 9352
rect 22978 9272 22979 9336
rect 23043 9272 23044 9336
rect 22978 9256 23044 9272
rect 22978 9192 22979 9256
rect 23043 9192 23044 9256
rect 22978 9176 23044 9192
rect 22978 9112 22979 9176
rect 23043 9112 23044 9176
rect 22978 8958 23044 9112
rect 23104 8958 23164 9990
rect 23224 9020 23284 10050
rect 23344 8958 23404 9990
rect 23464 9020 23524 10050
rect 23584 9896 23650 9986
rect 23584 9832 23585 9896
rect 23649 9832 23650 9896
rect 23584 9816 23650 9832
rect 23584 9752 23585 9816
rect 23649 9752 23650 9816
rect 23584 9736 23650 9752
rect 23584 9672 23585 9736
rect 23649 9672 23650 9736
rect 23584 9656 23650 9672
rect 23584 9592 23585 9656
rect 23649 9592 23650 9656
rect 23584 9576 23650 9592
rect 23584 9512 23585 9576
rect 23649 9512 23650 9576
rect 23584 9496 23650 9512
rect 23584 9432 23585 9496
rect 23649 9432 23650 9496
rect 23584 9416 23650 9432
rect 23584 9352 23585 9416
rect 23649 9352 23650 9416
rect 23584 9336 23650 9352
rect 23584 9272 23585 9336
rect 23649 9272 23650 9336
rect 23584 9256 23650 9272
rect 23584 9192 23585 9256
rect 23649 9192 23650 9256
rect 23584 9176 23650 9192
rect 23584 9112 23585 9176
rect 23649 9112 23650 9176
rect 23584 8958 23650 9112
rect 23710 9020 23770 10050
rect 23830 8958 23890 9990
rect 23950 9020 24010 10050
rect 24070 8958 24130 9990
rect 24190 9896 24256 9986
rect 24190 9832 24191 9896
rect 24255 9832 24256 9896
rect 24190 9816 24256 9832
rect 24190 9752 24191 9816
rect 24255 9752 24256 9816
rect 24190 9736 24256 9752
rect 24190 9672 24191 9736
rect 24255 9672 24256 9736
rect 24190 9656 24256 9672
rect 24190 9592 24191 9656
rect 24255 9592 24256 9656
rect 24190 9576 24256 9592
rect 24190 9512 24191 9576
rect 24255 9512 24256 9576
rect 24190 9496 24256 9512
rect 24190 9432 24191 9496
rect 24255 9432 24256 9496
rect 24190 9416 24256 9432
rect 24190 9352 24191 9416
rect 24255 9352 24256 9416
rect 24190 9336 24256 9352
rect 24190 9272 24191 9336
rect 24255 9272 24256 9336
rect 24190 9256 24256 9272
rect 24190 9192 24191 9256
rect 24255 9192 24256 9256
rect 24190 9176 24256 9192
rect 24190 9112 24191 9176
rect 24255 9112 24256 9176
rect 24190 8958 24256 9112
rect 24316 8958 24376 9990
rect 24436 9020 24496 10050
rect 24556 8958 24616 9990
rect 24676 9020 24736 10050
rect 24796 9896 24862 9986
rect 24796 9832 24797 9896
rect 24861 9832 24862 9896
rect 24796 9816 24862 9832
rect 24796 9752 24797 9816
rect 24861 9752 24862 9816
rect 24796 9736 24862 9752
rect 24796 9672 24797 9736
rect 24861 9672 24862 9736
rect 24796 9656 24862 9672
rect 24796 9592 24797 9656
rect 24861 9592 24862 9656
rect 24796 9576 24862 9592
rect 24796 9512 24797 9576
rect 24861 9512 24862 9576
rect 24796 9496 24862 9512
rect 24796 9432 24797 9496
rect 24861 9432 24862 9496
rect 24796 9416 24862 9432
rect 24796 9352 24797 9416
rect 24861 9352 24862 9416
rect 24796 9336 24862 9352
rect 24796 9272 24797 9336
rect 24861 9272 24862 9336
rect 24796 9256 24862 9272
rect 24796 9192 24797 9256
rect 24861 9192 24862 9256
rect 24796 9176 24862 9192
rect 24796 9112 24797 9176
rect 24861 9112 24862 9176
rect 24796 8958 24862 9112
rect 22372 8956 24862 8958
rect 22372 8892 22476 8956
rect 22540 8892 22556 8956
rect 22620 8892 22636 8956
rect 22700 8892 22716 8956
rect 22780 8892 22796 8956
rect 22860 8892 22876 8956
rect 22940 8892 23082 8956
rect 23146 8892 23162 8956
rect 23226 8892 23242 8956
rect 23306 8892 23322 8956
rect 23386 8892 23402 8956
rect 23466 8892 23482 8956
rect 23546 8892 23688 8956
rect 23752 8892 23768 8956
rect 23832 8892 23848 8956
rect 23912 8892 23928 8956
rect 23992 8892 24008 8956
rect 24072 8892 24088 8956
rect 24152 8892 24294 8956
rect 24358 8892 24374 8956
rect 24438 8892 24454 8956
rect 24518 8892 24534 8956
rect 24598 8892 24614 8956
rect 24678 8892 24694 8956
rect 24758 8892 24862 8956
rect 22372 8890 24862 8892
rect 24922 9896 24988 9986
rect 24922 9832 24923 9896
rect 24987 9832 24988 9896
rect 24922 9816 24988 9832
rect 24922 9752 24923 9816
rect 24987 9752 24988 9816
rect 24922 9736 24988 9752
rect 24922 9672 24923 9736
rect 24987 9672 24988 9736
rect 24922 9656 24988 9672
rect 24922 9592 24923 9656
rect 24987 9592 24988 9656
rect 24922 9576 24988 9592
rect 24922 9512 24923 9576
rect 24987 9512 24988 9576
rect 24922 9496 24988 9512
rect 24922 9432 24923 9496
rect 24987 9432 24988 9496
rect 24922 9416 24988 9432
rect 24922 9352 24923 9416
rect 24987 9352 24988 9416
rect 24922 9336 24988 9352
rect 24922 9272 24923 9336
rect 24987 9272 24988 9336
rect 24922 9256 24988 9272
rect 24922 9192 24923 9256
rect 24987 9192 24988 9256
rect 24922 9176 24988 9192
rect 24922 9112 24923 9176
rect 24987 9112 24988 9176
rect 24922 8958 24988 9112
rect 25048 8958 25108 9990
rect 25168 9020 25228 10050
rect 25288 8958 25348 9990
rect 25408 9020 25468 10050
rect 25857 10045 25982 10051
rect 25528 9896 25594 9986
rect 25528 9832 25529 9896
rect 25593 9832 25594 9896
rect 25528 9816 25594 9832
rect 25528 9752 25529 9816
rect 25593 9752 25594 9816
rect 25528 9736 25594 9752
rect 25528 9672 25529 9736
rect 25593 9672 25594 9736
rect 25528 9656 25594 9672
rect 25528 9592 25529 9656
rect 25593 9592 25594 9656
rect 25528 9576 25594 9592
rect 25528 9512 25529 9576
rect 25593 9512 25594 9576
rect 25528 9496 25594 9512
rect 25528 9432 25529 9496
rect 25593 9432 25594 9496
rect 25528 9416 25594 9432
rect 25528 9352 25529 9416
rect 25593 9352 25594 9416
rect 25528 9336 25594 9352
rect 25528 9272 25529 9336
rect 25593 9272 25594 9336
rect 25528 9256 25594 9272
rect 25528 9192 25529 9256
rect 25593 9192 25594 9256
rect 25528 9176 25594 9192
rect 25528 9112 25529 9176
rect 25593 9112 25594 9176
rect 25528 8958 25594 9112
rect 24922 8956 25594 8958
rect 24922 8892 25026 8956
rect 25090 8892 25106 8956
rect 25170 8892 25186 8956
rect 25250 8892 25266 8956
rect 25330 8892 25346 8956
rect 25410 8892 25426 8956
rect 25490 8892 25594 8956
rect 24922 8890 25594 8892
rect 20041 8729 20239 8739
rect 20041 8665 20054 8729
rect 20118 8665 20239 8729
rect 25273 8711 25945 8713
rect 20041 8655 20239 8665
rect 20299 8708 25213 8710
rect 20299 8644 20403 8708
rect 20467 8644 20483 8708
rect 20547 8644 20563 8708
rect 20627 8644 20643 8708
rect 20707 8644 20723 8708
rect 20787 8644 20803 8708
rect 20867 8644 21009 8708
rect 21073 8644 21089 8708
rect 21153 8644 21169 8708
rect 21233 8644 21249 8708
rect 21313 8644 21329 8708
rect 21393 8644 21409 8708
rect 21473 8644 21615 8708
rect 21679 8644 21695 8708
rect 21759 8644 21775 8708
rect 21839 8644 21855 8708
rect 21919 8644 21935 8708
rect 21999 8644 22015 8708
rect 22079 8644 22221 8708
rect 22285 8644 22301 8708
rect 22365 8644 22381 8708
rect 22445 8644 22461 8708
rect 22525 8644 22541 8708
rect 22605 8644 22621 8708
rect 22685 8644 22827 8708
rect 22891 8644 22907 8708
rect 22971 8644 22987 8708
rect 23051 8644 23067 8708
rect 23131 8644 23147 8708
rect 23211 8644 23227 8708
rect 23291 8644 23433 8708
rect 23497 8644 23513 8708
rect 23577 8644 23593 8708
rect 23657 8644 23673 8708
rect 23737 8644 23753 8708
rect 23817 8644 23833 8708
rect 23897 8644 24039 8708
rect 24103 8644 24119 8708
rect 24183 8644 24199 8708
rect 24263 8644 24279 8708
rect 24343 8644 24359 8708
rect 24423 8644 24439 8708
rect 24503 8644 24645 8708
rect 24709 8644 24725 8708
rect 24789 8644 24805 8708
rect 24869 8644 24885 8708
rect 24949 8644 24965 8708
rect 25029 8644 25045 8708
rect 25109 8644 25213 8708
rect 20299 8642 25213 8644
rect 20299 8488 20365 8642
rect 19921 8468 20239 8480
rect 19921 8404 20142 8468
rect 20206 8404 20239 8468
rect 19921 8226 20239 8404
rect 19170 8091 19236 8107
rect 19170 8027 19171 8091
rect 19235 8027 19236 8091
rect 19444 8147 19861 8165
rect 19444 8146 19651 8147
rect 19444 8088 19507 8146
rect 19170 8011 19236 8027
rect 19170 7947 19171 8011
rect 19235 7947 19236 8011
rect 19170 7931 19236 7947
rect 19170 7867 19171 7931
rect 19235 7867 19236 7931
rect 19170 7851 19236 7867
rect 19170 7787 19171 7851
rect 19235 7787 19236 7851
rect 19170 7771 19236 7787
rect 19170 7707 19171 7771
rect 19235 7707 19236 7771
rect 19170 7617 19236 7707
rect 19443 8082 19507 8088
rect 19571 8083 19651 8146
rect 19715 8146 19861 8147
rect 19715 8083 19782 8146
rect 19571 8082 19782 8083
rect 19846 8082 19861 8146
rect 19443 7997 19861 8082
rect 19443 7933 19637 7997
rect 19701 7933 19861 7997
rect 19443 7801 19861 7933
rect 19443 7737 19637 7801
rect 19701 7737 19861 7801
rect 19443 7626 19861 7737
rect 19443 7562 19637 7626
rect 19701 7562 19861 7626
rect 18564 7552 19236 7553
rect 18563 7551 19236 7552
rect 18563 7550 18668 7551
rect 13420 7548 18668 7550
rect 13420 7539 13694 7548
rect 12824 7484 13694 7539
rect 13758 7484 13774 7548
rect 13838 7484 13854 7548
rect 13918 7484 13934 7548
rect 13998 7484 14014 7548
rect 14078 7484 14094 7548
rect 14158 7484 14300 7548
rect 14364 7484 14380 7548
rect 14444 7484 14460 7548
rect 14524 7484 14540 7548
rect 14604 7484 14620 7548
rect 14684 7484 14700 7548
rect 14764 7484 14906 7548
rect 14970 7484 14986 7548
rect 15050 7484 15066 7548
rect 15130 7484 15146 7548
rect 15210 7484 15226 7548
rect 15290 7484 15306 7548
rect 15370 7484 15512 7548
rect 15576 7484 15592 7548
rect 15656 7484 15672 7548
rect 15736 7484 15752 7548
rect 15816 7484 15832 7548
rect 15896 7484 15912 7548
rect 15976 7484 16118 7548
rect 16182 7484 16198 7548
rect 16262 7484 16278 7548
rect 16342 7484 16358 7548
rect 16422 7484 16438 7548
rect 16502 7484 16518 7548
rect 16582 7484 16724 7548
rect 16788 7484 16804 7548
rect 16868 7484 16884 7548
rect 16948 7484 16964 7548
rect 17028 7484 17044 7548
rect 17108 7484 17124 7548
rect 17188 7484 17330 7548
rect 17394 7484 17410 7548
rect 17474 7484 17490 7548
rect 17554 7484 17570 7548
rect 17634 7484 17650 7548
rect 17714 7484 17730 7548
rect 17794 7484 17936 7548
rect 18000 7484 18016 7548
rect 18080 7484 18096 7548
rect 18160 7484 18176 7548
rect 18240 7484 18256 7548
rect 18320 7484 18336 7548
rect 18400 7487 18668 7548
rect 18732 7487 18748 7551
rect 18812 7487 18828 7551
rect 18892 7487 18908 7551
rect 18972 7487 18988 7551
rect 19052 7487 19068 7551
rect 19132 7550 19236 7551
rect 19443 7550 19861 7562
rect 19132 7541 19861 7550
rect 19132 7487 19165 7541
rect 18400 7484 19165 7487
rect 12824 7477 19165 7484
rect 19229 7502 19861 7541
rect 19921 8162 20060 8226
rect 20124 8162 20239 8226
rect 19921 8069 20239 8162
rect 19921 8005 20059 8069
rect 20123 8005 20239 8069
rect 19921 7899 20239 8005
rect 19921 7835 20059 7899
rect 20123 7835 20239 7899
rect 19921 7747 20239 7835
rect 19921 7683 20060 7747
rect 20124 7683 20239 7747
rect 19921 7603 20239 7683
rect 20299 8424 20300 8488
rect 20364 8424 20365 8488
rect 20299 8408 20365 8424
rect 20299 8344 20300 8408
rect 20364 8344 20365 8408
rect 20299 8328 20365 8344
rect 20299 8264 20300 8328
rect 20364 8264 20365 8328
rect 20299 8248 20365 8264
rect 20299 8184 20300 8248
rect 20364 8184 20365 8248
rect 20299 8168 20365 8184
rect 20299 8104 20300 8168
rect 20364 8104 20365 8168
rect 20299 8088 20365 8104
rect 20299 8024 20300 8088
rect 20364 8024 20365 8088
rect 20299 8008 20365 8024
rect 20299 7944 20300 8008
rect 20364 7944 20365 8008
rect 20299 7928 20365 7944
rect 20299 7864 20300 7928
rect 20364 7864 20365 7928
rect 20299 7848 20365 7864
rect 20299 7784 20300 7848
rect 20364 7784 20365 7848
rect 20299 7768 20365 7784
rect 20299 7704 20300 7768
rect 20364 7704 20365 7768
rect 20299 7614 20365 7704
rect 19921 7539 20065 7603
rect 20129 7550 20239 7603
rect 20425 7550 20485 8580
rect 20545 7610 20605 8642
rect 20665 7550 20725 8580
rect 20785 7610 20845 8642
rect 20905 8488 20971 8642
rect 20905 8424 20906 8488
rect 20970 8424 20971 8488
rect 20905 8408 20971 8424
rect 20905 8344 20906 8408
rect 20970 8344 20971 8408
rect 20905 8328 20971 8344
rect 20905 8264 20906 8328
rect 20970 8264 20971 8328
rect 20905 8248 20971 8264
rect 20905 8184 20906 8248
rect 20970 8184 20971 8248
rect 20905 8168 20971 8184
rect 20905 8104 20906 8168
rect 20970 8104 20971 8168
rect 20905 8088 20971 8104
rect 20905 8024 20906 8088
rect 20970 8024 20971 8088
rect 20905 8008 20971 8024
rect 20905 7944 20906 8008
rect 20970 7944 20971 8008
rect 20905 7928 20971 7944
rect 20905 7864 20906 7928
rect 20970 7864 20971 7928
rect 20905 7848 20971 7864
rect 20905 7784 20906 7848
rect 20970 7784 20971 7848
rect 20905 7768 20971 7784
rect 20905 7704 20906 7768
rect 20970 7704 20971 7768
rect 20905 7614 20971 7704
rect 21031 7610 21091 8642
rect 21151 7550 21211 8580
rect 21271 7610 21331 8642
rect 21391 7550 21451 8580
rect 21511 8488 21577 8642
rect 21511 8424 21512 8488
rect 21576 8424 21577 8488
rect 21511 8408 21577 8424
rect 21511 8344 21512 8408
rect 21576 8344 21577 8408
rect 21511 8328 21577 8344
rect 21511 8264 21512 8328
rect 21576 8264 21577 8328
rect 21511 8248 21577 8264
rect 21511 8184 21512 8248
rect 21576 8184 21577 8248
rect 21511 8168 21577 8184
rect 21511 8104 21512 8168
rect 21576 8104 21577 8168
rect 21511 8088 21577 8104
rect 21511 8024 21512 8088
rect 21576 8024 21577 8088
rect 21511 8008 21577 8024
rect 21511 7944 21512 8008
rect 21576 7944 21577 8008
rect 21511 7928 21577 7944
rect 21511 7864 21512 7928
rect 21576 7864 21577 7928
rect 21511 7848 21577 7864
rect 21511 7784 21512 7848
rect 21576 7784 21577 7848
rect 21511 7768 21577 7784
rect 21511 7704 21512 7768
rect 21576 7704 21577 7768
rect 21511 7614 21577 7704
rect 21637 7550 21697 8580
rect 21757 7610 21817 8642
rect 21877 7550 21937 8580
rect 21997 7610 22057 8642
rect 22117 8488 22183 8642
rect 22117 8424 22118 8488
rect 22182 8424 22183 8488
rect 22117 8408 22183 8424
rect 22117 8344 22118 8408
rect 22182 8344 22183 8408
rect 22117 8328 22183 8344
rect 22117 8264 22118 8328
rect 22182 8264 22183 8328
rect 22117 8248 22183 8264
rect 22117 8184 22118 8248
rect 22182 8184 22183 8248
rect 22117 8168 22183 8184
rect 22117 8104 22118 8168
rect 22182 8104 22183 8168
rect 22117 8088 22183 8104
rect 22117 8024 22118 8088
rect 22182 8024 22183 8088
rect 22117 8008 22183 8024
rect 22117 7944 22118 8008
rect 22182 7944 22183 8008
rect 22117 7928 22183 7944
rect 22117 7864 22118 7928
rect 22182 7864 22183 7928
rect 22117 7848 22183 7864
rect 22117 7784 22118 7848
rect 22182 7784 22183 7848
rect 22117 7768 22183 7784
rect 22117 7704 22118 7768
rect 22182 7704 22183 7768
rect 22117 7614 22183 7704
rect 22243 7610 22303 8642
rect 22363 7550 22423 8580
rect 22483 7610 22543 8642
rect 22603 7550 22663 8580
rect 22723 8488 22789 8642
rect 22723 8424 22724 8488
rect 22788 8424 22789 8488
rect 22723 8408 22789 8424
rect 22723 8344 22724 8408
rect 22788 8344 22789 8408
rect 22723 8328 22789 8344
rect 22723 8264 22724 8328
rect 22788 8264 22789 8328
rect 22723 8248 22789 8264
rect 22723 8184 22724 8248
rect 22788 8184 22789 8248
rect 22723 8168 22789 8184
rect 22723 8104 22724 8168
rect 22788 8104 22789 8168
rect 22723 8088 22789 8104
rect 22723 8024 22724 8088
rect 22788 8024 22789 8088
rect 22723 8008 22789 8024
rect 22723 7944 22724 8008
rect 22788 7944 22789 8008
rect 22723 7928 22789 7944
rect 22723 7864 22724 7928
rect 22788 7864 22789 7928
rect 22723 7848 22789 7864
rect 22723 7784 22724 7848
rect 22788 7784 22789 7848
rect 22723 7768 22789 7784
rect 22723 7704 22724 7768
rect 22788 7704 22789 7768
rect 22723 7614 22789 7704
rect 22849 7550 22909 8580
rect 22969 7610 23029 8642
rect 23089 7550 23149 8580
rect 23209 7610 23269 8642
rect 23329 8488 23395 8642
rect 23329 8424 23330 8488
rect 23394 8424 23395 8488
rect 23329 8408 23395 8424
rect 23329 8344 23330 8408
rect 23394 8344 23395 8408
rect 23329 8328 23395 8344
rect 23329 8264 23330 8328
rect 23394 8264 23395 8328
rect 23329 8248 23395 8264
rect 23329 8184 23330 8248
rect 23394 8184 23395 8248
rect 23329 8168 23395 8184
rect 23329 8104 23330 8168
rect 23394 8104 23395 8168
rect 23329 8088 23395 8104
rect 23329 8024 23330 8088
rect 23394 8024 23395 8088
rect 23329 8008 23395 8024
rect 23329 7944 23330 8008
rect 23394 7944 23395 8008
rect 23329 7928 23395 7944
rect 23329 7864 23330 7928
rect 23394 7864 23395 7928
rect 23329 7848 23395 7864
rect 23329 7784 23330 7848
rect 23394 7784 23395 7848
rect 23329 7768 23395 7784
rect 23329 7704 23330 7768
rect 23394 7704 23395 7768
rect 23329 7614 23395 7704
rect 23455 7610 23515 8642
rect 23575 7550 23635 8580
rect 23695 7610 23755 8642
rect 23815 7550 23875 8580
rect 23935 8488 24001 8642
rect 23935 8424 23936 8488
rect 24000 8424 24001 8488
rect 23935 8408 24001 8424
rect 23935 8344 23936 8408
rect 24000 8344 24001 8408
rect 23935 8328 24001 8344
rect 23935 8264 23936 8328
rect 24000 8264 24001 8328
rect 23935 8248 24001 8264
rect 23935 8184 23936 8248
rect 24000 8184 24001 8248
rect 23935 8168 24001 8184
rect 23935 8104 23936 8168
rect 24000 8104 24001 8168
rect 23935 8088 24001 8104
rect 23935 8024 23936 8088
rect 24000 8024 24001 8088
rect 23935 8008 24001 8024
rect 23935 7944 23936 8008
rect 24000 7944 24001 8008
rect 23935 7928 24001 7944
rect 23935 7864 23936 7928
rect 24000 7864 24001 7928
rect 23935 7848 24001 7864
rect 23935 7784 23936 7848
rect 24000 7784 24001 7848
rect 23935 7768 24001 7784
rect 23935 7704 23936 7768
rect 24000 7704 24001 7768
rect 23935 7614 24001 7704
rect 24061 7550 24121 8580
rect 24181 7610 24241 8642
rect 24301 7550 24361 8580
rect 24421 7610 24481 8642
rect 24541 8488 24607 8642
rect 24541 8424 24542 8488
rect 24606 8424 24607 8488
rect 24541 8408 24607 8424
rect 24541 8344 24542 8408
rect 24606 8344 24607 8408
rect 24541 8328 24607 8344
rect 24541 8264 24542 8328
rect 24606 8264 24607 8328
rect 24541 8248 24607 8264
rect 24541 8184 24542 8248
rect 24606 8184 24607 8248
rect 24541 8168 24607 8184
rect 24541 8104 24542 8168
rect 24606 8104 24607 8168
rect 24541 8088 24607 8104
rect 24541 8024 24542 8088
rect 24606 8024 24607 8088
rect 24541 8008 24607 8024
rect 24541 7944 24542 8008
rect 24606 7944 24607 8008
rect 24541 7928 24607 7944
rect 24541 7864 24542 7928
rect 24606 7864 24607 7928
rect 24541 7848 24607 7864
rect 24541 7784 24542 7848
rect 24606 7784 24607 7848
rect 24541 7768 24607 7784
rect 24541 7704 24542 7768
rect 24606 7704 24607 7768
rect 24541 7614 24607 7704
rect 24667 7610 24727 8642
rect 24787 7550 24847 8580
rect 24907 7610 24967 8642
rect 25027 7550 25087 8580
rect 25147 8488 25213 8642
rect 25147 8424 25148 8488
rect 25212 8424 25213 8488
rect 25147 8408 25213 8424
rect 25147 8344 25148 8408
rect 25212 8344 25213 8408
rect 25147 8328 25213 8344
rect 25147 8264 25148 8328
rect 25212 8264 25213 8328
rect 25147 8248 25213 8264
rect 25147 8184 25148 8248
rect 25212 8184 25213 8248
rect 25147 8168 25213 8184
rect 25147 8104 25148 8168
rect 25212 8104 25213 8168
rect 25147 8088 25213 8104
rect 25147 8024 25148 8088
rect 25212 8024 25213 8088
rect 25147 8008 25213 8024
rect 25147 7944 25148 8008
rect 25212 7944 25213 8008
rect 25147 7928 25213 7944
rect 25147 7864 25148 7928
rect 25212 7864 25213 7928
rect 25147 7848 25213 7864
rect 25147 7784 25148 7848
rect 25212 7784 25213 7848
rect 25147 7768 25213 7784
rect 25147 7704 25148 7768
rect 25212 7704 25213 7768
rect 25147 7614 25213 7704
rect 25273 8647 25377 8711
rect 25441 8647 25457 8711
rect 25521 8647 25537 8711
rect 25601 8647 25617 8711
rect 25681 8647 25697 8711
rect 25761 8647 25777 8711
rect 25841 8647 25945 8711
rect 26166 8692 26676 10051
rect 25273 8645 25945 8647
rect 25273 8491 25339 8645
rect 25273 8427 25274 8491
rect 25338 8427 25339 8491
rect 25273 8411 25339 8427
rect 25273 8347 25274 8411
rect 25338 8347 25339 8411
rect 25273 8331 25339 8347
rect 25273 8267 25274 8331
rect 25338 8267 25339 8331
rect 25273 8251 25339 8267
rect 25273 8187 25274 8251
rect 25338 8187 25339 8251
rect 25273 8171 25339 8187
rect 25273 8107 25274 8171
rect 25338 8107 25339 8171
rect 25273 8091 25339 8107
rect 25273 8027 25274 8091
rect 25338 8027 25339 8091
rect 25273 8011 25339 8027
rect 25273 7947 25274 8011
rect 25338 7947 25339 8011
rect 25273 7931 25339 7947
rect 25273 7867 25274 7931
rect 25338 7867 25339 7931
rect 25273 7851 25339 7867
rect 25273 7787 25274 7851
rect 25338 7787 25339 7851
rect 25273 7771 25339 7787
rect 25273 7707 25274 7771
rect 25338 7707 25339 7771
rect 25273 7617 25339 7707
rect 25399 7613 25459 8645
rect 25519 7553 25579 8583
rect 25639 7613 25699 8645
rect 25759 7553 25819 8583
rect 25879 8491 25945 8645
rect 26167 8628 26210 8692
rect 26274 8628 26353 8692
rect 26417 8628 26473 8692
rect 26537 8689 26676 8692
rect 26537 8628 26544 8689
rect 26167 8613 26544 8628
rect 25879 8427 25880 8491
rect 25944 8427 25945 8491
rect 25879 8411 25945 8427
rect 25879 8347 25880 8411
rect 25944 8347 25945 8411
rect 25879 8331 25945 8347
rect 25879 8267 25880 8331
rect 25944 8267 25945 8331
rect 25879 8251 25945 8267
rect 25879 8187 25880 8251
rect 25944 8187 25945 8251
rect 25879 8171 25945 8187
rect 25879 8107 25880 8171
rect 25944 8107 25945 8171
rect 25879 8091 25945 8107
rect 25879 8027 25880 8091
rect 25944 8027 25945 8091
rect 26153 8147 26570 8165
rect 26153 8146 26360 8147
rect 26153 8088 26216 8146
rect 25879 8011 25945 8027
rect 25879 7947 25880 8011
rect 25944 7947 25945 8011
rect 25879 7931 25945 7947
rect 25879 7867 25880 7931
rect 25944 7867 25945 7931
rect 25879 7851 25945 7867
rect 25879 7787 25880 7851
rect 25944 7787 25945 7851
rect 25879 7771 25945 7787
rect 25879 7707 25880 7771
rect 25944 7707 25945 7771
rect 25879 7617 25945 7707
rect 26152 8082 26216 8088
rect 26280 8083 26360 8146
rect 26424 8146 26570 8147
rect 26424 8083 26491 8146
rect 26280 8082 26491 8083
rect 26555 8082 26570 8146
rect 25273 7552 25945 7553
rect 25272 7551 25945 7552
rect 25272 7550 25377 7551
rect 20129 7548 25377 7550
rect 20129 7539 20403 7548
rect 19921 7502 20403 7539
rect 19229 7484 20403 7502
rect 20467 7484 20483 7548
rect 20547 7484 20563 7548
rect 20627 7484 20643 7548
rect 20707 7484 20723 7548
rect 20787 7484 20803 7548
rect 20867 7484 21009 7548
rect 21073 7484 21089 7548
rect 21153 7484 21169 7548
rect 21233 7484 21249 7548
rect 21313 7484 21329 7548
rect 21393 7484 21409 7548
rect 21473 7484 21615 7548
rect 21679 7484 21695 7548
rect 21759 7484 21775 7548
rect 21839 7484 21855 7548
rect 21919 7484 21935 7548
rect 21999 7484 22015 7548
rect 22079 7484 22221 7548
rect 22285 7484 22301 7548
rect 22365 7484 22381 7548
rect 22445 7484 22461 7548
rect 22525 7484 22541 7548
rect 22605 7484 22621 7548
rect 22685 7484 22827 7548
rect 22891 7484 22907 7548
rect 22971 7484 22987 7548
rect 23051 7484 23067 7548
rect 23131 7484 23147 7548
rect 23211 7484 23227 7548
rect 23291 7484 23433 7548
rect 23497 7484 23513 7548
rect 23577 7484 23593 7548
rect 23657 7484 23673 7548
rect 23737 7484 23753 7548
rect 23817 7484 23833 7548
rect 23897 7484 24039 7548
rect 24103 7484 24119 7548
rect 24183 7484 24199 7548
rect 24263 7484 24279 7548
rect 24343 7484 24359 7548
rect 24423 7484 24439 7548
rect 24503 7484 24645 7548
rect 24709 7484 24725 7548
rect 24789 7484 24805 7548
rect 24869 7484 24885 7548
rect 24949 7484 24965 7548
rect 25029 7484 25045 7548
rect 25109 7487 25377 7548
rect 25441 7487 25457 7551
rect 25521 7487 25537 7551
rect 25601 7487 25617 7551
rect 25681 7487 25697 7551
rect 25761 7487 25777 7551
rect 25841 7550 25945 7551
rect 26152 7550 26570 8082
rect 25841 7541 26570 7550
rect 25841 7487 25874 7541
rect 25109 7484 25874 7487
rect 19229 7477 25874 7484
rect 25938 7502 26570 7541
rect 26756 7502 27155 13625
rect 25938 7477 27155 7502
rect 12824 7444 27155 7477
rect 12825 7437 27155 7444
rect 12825 7358 27157 7437
rect 12826 7292 13822 7358
rect 12826 7212 13488 7292
rect 13654 7212 13822 7292
rect 12826 7134 13822 7212
rect 24043 7340 27157 7358
rect 24043 7335 31248 7340
rect 24043 7271 24675 7335
rect 24739 7328 31248 7335
rect 24739 7325 25504 7328
rect 24739 7271 24772 7325
rect 24043 7262 24772 7271
rect 10753 7080 14359 7134
rect 10753 6934 10891 7080
rect 11041 7064 14359 7080
rect 11041 6934 11203 7064
rect 10753 6918 11203 6934
rect 11353 6918 14359 7064
rect 10753 6132 14359 6918
rect 10753 6120 11261 6132
rect 10753 5974 10955 6120
rect 11105 5986 11261 6120
rect 11411 5986 14359 6132
rect 11105 5974 14359 5986
rect 10753 5492 14359 5974
rect 10753 5346 10787 5492
rect 10937 5346 14359 5492
rect 10753 4654 14359 5346
rect 10753 4650 12187 4654
rect 10753 4646 11175 4650
rect 10753 4500 10823 4646
rect 10973 4504 11175 4646
rect 11325 4504 11621 4650
rect 11771 4508 12187 4650
rect 12337 4508 12853 4654
rect 13003 4638 14359 4654
rect 13003 4508 13235 4638
rect 11771 4504 13235 4508
rect 10973 4500 13235 4504
rect 10753 4492 13235 4500
rect 13385 4492 14359 4638
rect 10753 3800 14359 4492
rect 10753 3792 11255 3800
rect 10753 3646 10905 3792
rect 11055 3654 11255 3792
rect 11405 3654 14359 3800
rect 11055 3646 14359 3654
rect 10753 3212 14359 3646
rect 8122 2660 10580 2874
rect 10751 3164 14359 3212
rect 23357 7108 23859 7110
rect 23357 6466 23907 7108
rect 24043 6730 24461 7262
rect 24668 7261 24772 7262
rect 24836 7261 24852 7325
rect 24916 7261 24932 7325
rect 24996 7261 25012 7325
rect 25076 7261 25092 7325
rect 25156 7261 25172 7325
rect 25236 7264 25504 7325
rect 25568 7264 25584 7328
rect 25648 7264 25664 7328
rect 25728 7264 25744 7328
rect 25808 7264 25824 7328
rect 25888 7264 25904 7328
rect 25968 7264 26110 7328
rect 26174 7264 26190 7328
rect 26254 7264 26270 7328
rect 26334 7264 26350 7328
rect 26414 7264 26430 7328
rect 26494 7264 26510 7328
rect 26574 7264 26716 7328
rect 26780 7264 26796 7328
rect 26860 7264 26876 7328
rect 26940 7264 26956 7328
rect 27020 7264 27036 7328
rect 27100 7264 27116 7328
rect 27180 7264 27322 7328
rect 27386 7264 27402 7328
rect 27466 7264 27482 7328
rect 27546 7264 27562 7328
rect 27626 7264 27642 7328
rect 27706 7264 27722 7328
rect 27786 7264 27928 7328
rect 27992 7264 28008 7328
rect 28072 7264 28088 7328
rect 28152 7264 28168 7328
rect 28232 7264 28248 7328
rect 28312 7264 28328 7328
rect 28392 7264 28534 7328
rect 28598 7264 28614 7328
rect 28678 7264 28694 7328
rect 28758 7264 28774 7328
rect 28838 7264 28854 7328
rect 28918 7264 28934 7328
rect 28998 7264 29140 7328
rect 29204 7264 29220 7328
rect 29284 7264 29300 7328
rect 29364 7264 29380 7328
rect 29444 7264 29460 7328
rect 29524 7264 29540 7328
rect 29604 7264 29746 7328
rect 29810 7264 29826 7328
rect 29890 7264 29906 7328
rect 29970 7264 29986 7328
rect 30050 7264 30066 7328
rect 30130 7264 30146 7328
rect 30210 7273 31248 7328
rect 30210 7264 30484 7273
rect 25236 7262 30484 7264
rect 25236 7261 25341 7262
rect 24668 7260 25341 7261
rect 24668 7259 25340 7260
rect 24043 6666 24058 6730
rect 24122 6729 24333 6730
rect 24122 6666 24189 6729
rect 24043 6665 24189 6666
rect 24253 6666 24333 6729
rect 24397 6724 24461 6730
rect 24668 7105 24734 7195
rect 24668 7041 24669 7105
rect 24733 7041 24734 7105
rect 24668 7025 24734 7041
rect 24668 6961 24669 7025
rect 24733 6961 24734 7025
rect 24668 6945 24734 6961
rect 24668 6881 24669 6945
rect 24733 6881 24734 6945
rect 24668 6865 24734 6881
rect 24668 6801 24669 6865
rect 24733 6801 24734 6865
rect 24668 6785 24734 6801
rect 24397 6666 24460 6724
rect 24253 6665 24460 6666
rect 24043 6647 24460 6665
rect 24668 6721 24669 6785
rect 24733 6721 24734 6785
rect 24668 6705 24734 6721
rect 23357 6320 23609 6466
rect 23759 6320 23907 6466
rect 23357 6040 23907 6320
rect 24668 6641 24669 6705
rect 24733 6641 24734 6705
rect 24668 6625 24734 6641
rect 24668 6561 24669 6625
rect 24733 6561 24734 6625
rect 24668 6545 24734 6561
rect 24668 6481 24669 6545
rect 24733 6481 24734 6545
rect 24668 6465 24734 6481
rect 24668 6401 24669 6465
rect 24733 6401 24734 6465
rect 24668 6385 24734 6401
rect 24668 6321 24669 6385
rect 24733 6321 24734 6385
rect 24069 6184 24446 6199
rect 24069 6120 24076 6184
rect 24140 6120 24196 6184
rect 24260 6120 24339 6184
rect 24403 6120 24446 6184
rect 24668 6167 24734 6321
rect 24794 6229 24854 7259
rect 24914 6167 24974 7199
rect 25034 6229 25094 7259
rect 25154 6167 25214 7199
rect 25274 7105 25340 7195
rect 25274 7041 25275 7105
rect 25339 7041 25340 7105
rect 25274 7025 25340 7041
rect 25274 6961 25275 7025
rect 25339 6961 25340 7025
rect 25274 6945 25340 6961
rect 25274 6881 25275 6945
rect 25339 6881 25340 6945
rect 25274 6865 25340 6881
rect 25274 6801 25275 6865
rect 25339 6801 25340 6865
rect 25274 6785 25340 6801
rect 25274 6721 25275 6785
rect 25339 6721 25340 6785
rect 25274 6705 25340 6721
rect 25274 6641 25275 6705
rect 25339 6641 25340 6705
rect 25274 6625 25340 6641
rect 25274 6561 25275 6625
rect 25339 6561 25340 6625
rect 25274 6545 25340 6561
rect 25274 6481 25275 6545
rect 25339 6481 25340 6545
rect 25274 6465 25340 6481
rect 25274 6401 25275 6465
rect 25339 6401 25340 6465
rect 25274 6385 25340 6401
rect 25274 6321 25275 6385
rect 25339 6321 25340 6385
rect 25274 6167 25340 6321
rect 24668 6165 25340 6167
rect 23357 5894 23609 6040
rect 23759 5894 23907 6040
rect 23357 5814 23907 5894
rect 23357 5668 23609 5814
rect 23759 5668 23907 5814
rect 23357 5080 23907 5668
rect 23357 4934 23625 5080
rect 23775 4934 23907 5080
rect 23357 4546 23907 4934
rect 24071 4761 24447 6120
rect 24668 6101 24772 6165
rect 24836 6101 24852 6165
rect 24916 6101 24932 6165
rect 24996 6101 25012 6165
rect 25076 6101 25092 6165
rect 25156 6101 25172 6165
rect 25236 6101 25340 6165
rect 25400 7108 25466 7198
rect 25400 7044 25401 7108
rect 25465 7044 25466 7108
rect 25400 7028 25466 7044
rect 25400 6964 25401 7028
rect 25465 6964 25466 7028
rect 25400 6948 25466 6964
rect 25400 6884 25401 6948
rect 25465 6884 25466 6948
rect 25400 6868 25466 6884
rect 25400 6804 25401 6868
rect 25465 6804 25466 6868
rect 25400 6788 25466 6804
rect 25400 6724 25401 6788
rect 25465 6724 25466 6788
rect 25400 6708 25466 6724
rect 25400 6644 25401 6708
rect 25465 6644 25466 6708
rect 25400 6628 25466 6644
rect 25400 6564 25401 6628
rect 25465 6564 25466 6628
rect 25400 6548 25466 6564
rect 25400 6484 25401 6548
rect 25465 6484 25466 6548
rect 25400 6468 25466 6484
rect 25400 6404 25401 6468
rect 25465 6404 25466 6468
rect 25400 6388 25466 6404
rect 25400 6324 25401 6388
rect 25465 6324 25466 6388
rect 25400 6170 25466 6324
rect 25526 6232 25586 7262
rect 25646 6170 25706 7202
rect 25766 6232 25826 7262
rect 25886 6170 25946 7202
rect 26006 7108 26072 7198
rect 26006 7044 26007 7108
rect 26071 7044 26072 7108
rect 26006 7028 26072 7044
rect 26006 6964 26007 7028
rect 26071 6964 26072 7028
rect 26006 6948 26072 6964
rect 26006 6884 26007 6948
rect 26071 6884 26072 6948
rect 26006 6868 26072 6884
rect 26006 6804 26007 6868
rect 26071 6804 26072 6868
rect 26006 6788 26072 6804
rect 26006 6724 26007 6788
rect 26071 6724 26072 6788
rect 26006 6708 26072 6724
rect 26006 6644 26007 6708
rect 26071 6644 26072 6708
rect 26006 6628 26072 6644
rect 26006 6564 26007 6628
rect 26071 6564 26072 6628
rect 26006 6548 26072 6564
rect 26006 6484 26007 6548
rect 26071 6484 26072 6548
rect 26006 6468 26072 6484
rect 26006 6404 26007 6468
rect 26071 6404 26072 6468
rect 26006 6388 26072 6404
rect 26006 6324 26007 6388
rect 26071 6324 26072 6388
rect 26006 6170 26072 6324
rect 26132 6170 26192 7202
rect 26252 6232 26312 7262
rect 26372 6170 26432 7202
rect 26492 6232 26552 7262
rect 26612 7108 26678 7198
rect 26612 7044 26613 7108
rect 26677 7044 26678 7108
rect 26612 7028 26678 7044
rect 26612 6964 26613 7028
rect 26677 6964 26678 7028
rect 26612 6948 26678 6964
rect 26612 6884 26613 6948
rect 26677 6884 26678 6948
rect 26612 6868 26678 6884
rect 26612 6804 26613 6868
rect 26677 6804 26678 6868
rect 26612 6788 26678 6804
rect 26612 6724 26613 6788
rect 26677 6724 26678 6788
rect 26612 6708 26678 6724
rect 26612 6644 26613 6708
rect 26677 6644 26678 6708
rect 26612 6628 26678 6644
rect 26612 6564 26613 6628
rect 26677 6564 26678 6628
rect 26612 6548 26678 6564
rect 26612 6484 26613 6548
rect 26677 6484 26678 6548
rect 26612 6468 26678 6484
rect 26612 6404 26613 6468
rect 26677 6404 26678 6468
rect 26612 6388 26678 6404
rect 26612 6324 26613 6388
rect 26677 6324 26678 6388
rect 26612 6170 26678 6324
rect 26738 6232 26798 7262
rect 26858 6170 26918 7202
rect 26978 6232 27038 7262
rect 27098 6170 27158 7202
rect 27218 7108 27284 7198
rect 27218 7044 27219 7108
rect 27283 7044 27284 7108
rect 27218 7028 27284 7044
rect 27218 6964 27219 7028
rect 27283 6964 27284 7028
rect 27218 6948 27284 6964
rect 27218 6884 27219 6948
rect 27283 6884 27284 6948
rect 27218 6868 27284 6884
rect 27218 6804 27219 6868
rect 27283 6804 27284 6868
rect 27218 6788 27284 6804
rect 27218 6724 27219 6788
rect 27283 6724 27284 6788
rect 27218 6708 27284 6724
rect 27218 6644 27219 6708
rect 27283 6644 27284 6708
rect 27218 6628 27284 6644
rect 27218 6564 27219 6628
rect 27283 6564 27284 6628
rect 27218 6548 27284 6564
rect 27218 6484 27219 6548
rect 27283 6484 27284 6548
rect 27218 6468 27284 6484
rect 27218 6404 27219 6468
rect 27283 6404 27284 6468
rect 27218 6388 27284 6404
rect 27218 6324 27219 6388
rect 27283 6324 27284 6388
rect 27218 6170 27284 6324
rect 27344 6170 27404 7202
rect 27464 6232 27524 7262
rect 27584 6170 27644 7202
rect 27704 6232 27764 7262
rect 27824 7108 27890 7198
rect 27824 7044 27825 7108
rect 27889 7044 27890 7108
rect 27824 7028 27890 7044
rect 27824 6964 27825 7028
rect 27889 6964 27890 7028
rect 27824 6948 27890 6964
rect 27824 6884 27825 6948
rect 27889 6884 27890 6948
rect 27824 6868 27890 6884
rect 27824 6804 27825 6868
rect 27889 6804 27890 6868
rect 27824 6788 27890 6804
rect 27824 6724 27825 6788
rect 27889 6724 27890 6788
rect 27824 6708 27890 6724
rect 27824 6644 27825 6708
rect 27889 6644 27890 6708
rect 27824 6628 27890 6644
rect 27824 6564 27825 6628
rect 27889 6564 27890 6628
rect 27824 6548 27890 6564
rect 27824 6484 27825 6548
rect 27889 6484 27890 6548
rect 27824 6468 27890 6484
rect 27824 6404 27825 6468
rect 27889 6404 27890 6468
rect 27824 6388 27890 6404
rect 27824 6324 27825 6388
rect 27889 6324 27890 6388
rect 27824 6170 27890 6324
rect 27950 6232 28010 7262
rect 28070 6170 28130 7202
rect 28190 6232 28250 7262
rect 28310 6170 28370 7202
rect 28430 7108 28496 7198
rect 28430 7044 28431 7108
rect 28495 7044 28496 7108
rect 28430 7028 28496 7044
rect 28430 6964 28431 7028
rect 28495 6964 28496 7028
rect 28430 6948 28496 6964
rect 28430 6884 28431 6948
rect 28495 6884 28496 6948
rect 28430 6868 28496 6884
rect 28430 6804 28431 6868
rect 28495 6804 28496 6868
rect 28430 6788 28496 6804
rect 28430 6724 28431 6788
rect 28495 6724 28496 6788
rect 28430 6708 28496 6724
rect 28430 6644 28431 6708
rect 28495 6644 28496 6708
rect 28430 6628 28496 6644
rect 28430 6564 28431 6628
rect 28495 6564 28496 6628
rect 28430 6548 28496 6564
rect 28430 6484 28431 6548
rect 28495 6484 28496 6548
rect 28430 6468 28496 6484
rect 28430 6404 28431 6468
rect 28495 6404 28496 6468
rect 28430 6388 28496 6404
rect 28430 6324 28431 6388
rect 28495 6324 28496 6388
rect 28430 6170 28496 6324
rect 28556 6170 28616 7202
rect 28676 6232 28736 7262
rect 28796 6170 28856 7202
rect 28916 6232 28976 7262
rect 29036 7108 29102 7198
rect 29036 7044 29037 7108
rect 29101 7044 29102 7108
rect 29036 7028 29102 7044
rect 29036 6964 29037 7028
rect 29101 6964 29102 7028
rect 29036 6948 29102 6964
rect 29036 6884 29037 6948
rect 29101 6884 29102 6948
rect 29036 6868 29102 6884
rect 29036 6804 29037 6868
rect 29101 6804 29102 6868
rect 29036 6788 29102 6804
rect 29036 6724 29037 6788
rect 29101 6724 29102 6788
rect 29036 6708 29102 6724
rect 29036 6644 29037 6708
rect 29101 6644 29102 6708
rect 29036 6628 29102 6644
rect 29036 6564 29037 6628
rect 29101 6564 29102 6628
rect 29036 6548 29102 6564
rect 29036 6484 29037 6548
rect 29101 6484 29102 6548
rect 29036 6468 29102 6484
rect 29036 6404 29037 6468
rect 29101 6404 29102 6468
rect 29036 6388 29102 6404
rect 29036 6324 29037 6388
rect 29101 6324 29102 6388
rect 29036 6170 29102 6324
rect 29162 6232 29222 7262
rect 29282 6170 29342 7202
rect 29402 6232 29462 7262
rect 29522 6170 29582 7202
rect 29642 7108 29708 7198
rect 29642 7044 29643 7108
rect 29707 7044 29708 7108
rect 29642 7028 29708 7044
rect 29642 6964 29643 7028
rect 29707 6964 29708 7028
rect 29642 6948 29708 6964
rect 29642 6884 29643 6948
rect 29707 6884 29708 6948
rect 29642 6868 29708 6884
rect 29642 6804 29643 6868
rect 29707 6804 29708 6868
rect 29642 6788 29708 6804
rect 29642 6724 29643 6788
rect 29707 6724 29708 6788
rect 29642 6708 29708 6724
rect 29642 6644 29643 6708
rect 29707 6644 29708 6708
rect 29642 6628 29708 6644
rect 29642 6564 29643 6628
rect 29707 6564 29708 6628
rect 29642 6548 29708 6564
rect 29642 6484 29643 6548
rect 29707 6484 29708 6548
rect 29642 6468 29708 6484
rect 29642 6404 29643 6468
rect 29707 6404 29708 6468
rect 29642 6388 29708 6404
rect 29642 6324 29643 6388
rect 29707 6324 29708 6388
rect 29642 6170 29708 6324
rect 29768 6170 29828 7202
rect 29888 6232 29948 7262
rect 30008 6170 30068 7202
rect 30128 6232 30188 7262
rect 30374 7209 30484 7262
rect 30548 7209 31248 7273
rect 30248 7108 30314 7198
rect 30248 7044 30249 7108
rect 30313 7044 30314 7108
rect 30248 7028 30314 7044
rect 30248 6964 30249 7028
rect 30313 6964 30314 7028
rect 30248 6948 30314 6964
rect 30248 6884 30249 6948
rect 30313 6884 30314 6948
rect 30248 6868 30314 6884
rect 30248 6804 30249 6868
rect 30313 6804 30314 6868
rect 30248 6788 30314 6804
rect 30248 6724 30249 6788
rect 30313 6724 30314 6788
rect 30248 6708 30314 6724
rect 30248 6644 30249 6708
rect 30313 6644 30314 6708
rect 30248 6628 30314 6644
rect 30248 6564 30249 6628
rect 30313 6564 30314 6628
rect 30248 6548 30314 6564
rect 30248 6484 30249 6548
rect 30313 6484 30314 6548
rect 30248 6468 30314 6484
rect 30248 6404 30249 6468
rect 30313 6404 30314 6468
rect 30248 6388 30314 6404
rect 30248 6324 30249 6388
rect 30313 6324 30314 6388
rect 30374 7129 30700 7209
rect 30374 7065 30489 7129
rect 30553 7065 30700 7129
rect 30374 6977 30700 7065
rect 30374 6913 30490 6977
rect 30554 6934 30700 6977
rect 30797 6934 31248 7209
rect 30554 6913 31248 6934
rect 30374 6807 31248 6913
rect 30374 6743 30490 6807
rect 30554 6743 31248 6807
rect 30374 6650 31248 6743
rect 30374 6586 30489 6650
rect 30553 6586 31248 6650
rect 30374 6416 31248 6586
rect 30374 6408 30784 6416
rect 30374 6344 30407 6408
rect 30471 6353 30784 6408
rect 30471 6344 30692 6353
rect 30374 6332 30692 6344
rect 30248 6170 30314 6324
rect 25400 6168 30314 6170
rect 25400 6104 25504 6168
rect 25568 6104 25584 6168
rect 25648 6104 25664 6168
rect 25728 6104 25744 6168
rect 25808 6104 25824 6168
rect 25888 6104 25904 6168
rect 25968 6104 26110 6168
rect 26174 6104 26190 6168
rect 26254 6104 26270 6168
rect 26334 6104 26350 6168
rect 26414 6104 26430 6168
rect 26494 6104 26510 6168
rect 26574 6104 26716 6168
rect 26780 6104 26796 6168
rect 26860 6104 26876 6168
rect 26940 6104 26956 6168
rect 27020 6104 27036 6168
rect 27100 6104 27116 6168
rect 27180 6104 27322 6168
rect 27386 6104 27402 6168
rect 27466 6104 27482 6168
rect 27546 6104 27562 6168
rect 27626 6104 27642 6168
rect 27706 6104 27722 6168
rect 27786 6104 27928 6168
rect 27992 6104 28008 6168
rect 28072 6104 28088 6168
rect 28152 6104 28168 6168
rect 28232 6104 28248 6168
rect 28312 6104 28328 6168
rect 28392 6104 28534 6168
rect 28598 6104 28614 6168
rect 28678 6104 28694 6168
rect 28758 6104 28774 6168
rect 28838 6104 28854 6168
rect 28918 6104 28934 6168
rect 28998 6104 29140 6168
rect 29204 6104 29220 6168
rect 29284 6104 29300 6168
rect 29364 6104 29380 6168
rect 29444 6104 29460 6168
rect 29524 6104 29540 6168
rect 29604 6104 29746 6168
rect 29810 6104 29826 6168
rect 29890 6104 29906 6168
rect 29970 6104 29986 6168
rect 30050 6104 30066 6168
rect 30130 6104 30146 6168
rect 30210 6104 30314 6168
rect 25400 6102 30314 6104
rect 30374 6147 30572 6157
rect 24668 6099 25340 6101
rect 30374 6083 30495 6147
rect 30559 6083 30572 6147
rect 30374 6073 30572 6083
rect 25019 5920 25691 5922
rect 25019 5856 25123 5920
rect 25187 5856 25203 5920
rect 25267 5856 25283 5920
rect 25347 5856 25363 5920
rect 25427 5856 25443 5920
rect 25507 5856 25523 5920
rect 25587 5856 25691 5920
rect 25019 5854 25691 5856
rect 25019 5700 25085 5854
rect 25019 5636 25020 5700
rect 25084 5636 25085 5700
rect 25019 5620 25085 5636
rect 25019 5556 25020 5620
rect 25084 5556 25085 5620
rect 25019 5540 25085 5556
rect 25019 5476 25020 5540
rect 25084 5476 25085 5540
rect 25019 5460 25085 5476
rect 25019 5396 25020 5460
rect 25084 5396 25085 5460
rect 25019 5380 25085 5396
rect 25019 5316 25020 5380
rect 25084 5316 25085 5380
rect 25019 5300 25085 5316
rect 25019 5236 25020 5300
rect 25084 5236 25085 5300
rect 25019 5220 25085 5236
rect 25019 5156 25020 5220
rect 25084 5156 25085 5220
rect 25019 5140 25085 5156
rect 25019 5076 25020 5140
rect 25084 5076 25085 5140
rect 25019 5060 25085 5076
rect 25019 4996 25020 5060
rect 25084 4996 25085 5060
rect 25019 4980 25085 4996
rect 25019 4916 25020 4980
rect 25084 4916 25085 4980
rect 25019 4826 25085 4916
rect 24631 4761 24756 4767
rect 25145 4762 25205 5792
rect 25265 4822 25325 5854
rect 25385 4762 25445 5792
rect 25505 4822 25565 5854
rect 25625 5700 25691 5854
rect 25625 5636 25626 5700
rect 25690 5636 25691 5700
rect 25625 5620 25691 5636
rect 25625 5556 25626 5620
rect 25690 5556 25691 5620
rect 25625 5540 25691 5556
rect 25625 5476 25626 5540
rect 25690 5476 25691 5540
rect 25625 5460 25691 5476
rect 25625 5396 25626 5460
rect 25690 5396 25691 5460
rect 25625 5380 25691 5396
rect 25625 5316 25626 5380
rect 25690 5316 25691 5380
rect 25625 5300 25691 5316
rect 25625 5236 25626 5300
rect 25690 5236 25691 5300
rect 25625 5220 25691 5236
rect 25625 5156 25626 5220
rect 25690 5156 25691 5220
rect 25625 5140 25691 5156
rect 25625 5076 25626 5140
rect 25690 5076 25691 5140
rect 25625 5060 25691 5076
rect 25625 4996 25626 5060
rect 25690 4996 25691 5060
rect 25625 4980 25691 4996
rect 25625 4916 25626 4980
rect 25690 4916 25691 4980
rect 25625 4826 25691 4916
rect 25751 5920 28241 5922
rect 25751 5856 25855 5920
rect 25919 5856 25935 5920
rect 25999 5856 26015 5920
rect 26079 5856 26095 5920
rect 26159 5856 26175 5920
rect 26239 5856 26255 5920
rect 26319 5856 26461 5920
rect 26525 5856 26541 5920
rect 26605 5856 26621 5920
rect 26685 5856 26701 5920
rect 26765 5856 26781 5920
rect 26845 5856 26861 5920
rect 26925 5856 27067 5920
rect 27131 5856 27147 5920
rect 27211 5856 27227 5920
rect 27291 5856 27307 5920
rect 27371 5856 27387 5920
rect 27451 5856 27467 5920
rect 27531 5856 27673 5920
rect 27737 5856 27753 5920
rect 27817 5856 27833 5920
rect 27897 5856 27913 5920
rect 27977 5856 27993 5920
rect 28057 5856 28073 5920
rect 28137 5856 28241 5920
rect 25751 5854 28241 5856
rect 25751 5700 25817 5854
rect 25751 5636 25752 5700
rect 25816 5636 25817 5700
rect 25751 5620 25817 5636
rect 25751 5556 25752 5620
rect 25816 5556 25817 5620
rect 25751 5540 25817 5556
rect 25751 5476 25752 5540
rect 25816 5476 25817 5540
rect 25751 5460 25817 5476
rect 25751 5396 25752 5460
rect 25816 5396 25817 5460
rect 25751 5380 25817 5396
rect 25751 5316 25752 5380
rect 25816 5316 25817 5380
rect 25751 5300 25817 5316
rect 25751 5236 25752 5300
rect 25816 5236 25817 5300
rect 25751 5220 25817 5236
rect 25751 5156 25752 5220
rect 25816 5156 25817 5220
rect 25751 5140 25817 5156
rect 25751 5076 25752 5140
rect 25816 5076 25817 5140
rect 25751 5060 25817 5076
rect 25751 4996 25752 5060
rect 25816 4996 25817 5060
rect 25751 4980 25817 4996
rect 25751 4916 25752 4980
rect 25816 4916 25817 4980
rect 25751 4826 25817 4916
rect 25877 4762 25937 5792
rect 25997 4822 26057 5854
rect 26117 4762 26177 5792
rect 26237 4822 26297 5854
rect 26357 5700 26423 5854
rect 26357 5636 26358 5700
rect 26422 5636 26423 5700
rect 26357 5620 26423 5636
rect 26357 5556 26358 5620
rect 26422 5556 26423 5620
rect 26357 5540 26423 5556
rect 26357 5476 26358 5540
rect 26422 5476 26423 5540
rect 26357 5460 26423 5476
rect 26357 5396 26358 5460
rect 26422 5396 26423 5460
rect 26357 5380 26423 5396
rect 26357 5316 26358 5380
rect 26422 5316 26423 5380
rect 26357 5300 26423 5316
rect 26357 5236 26358 5300
rect 26422 5236 26423 5300
rect 26357 5220 26423 5236
rect 26357 5156 26358 5220
rect 26422 5156 26423 5220
rect 26357 5140 26423 5156
rect 26357 5076 26358 5140
rect 26422 5076 26423 5140
rect 26357 5060 26423 5076
rect 26357 4996 26358 5060
rect 26422 4996 26423 5060
rect 26357 4980 26423 4996
rect 26357 4916 26358 4980
rect 26422 4916 26423 4980
rect 26357 4826 26423 4916
rect 26483 4822 26543 5854
rect 26603 4762 26663 5792
rect 26723 4822 26783 5854
rect 26843 4762 26903 5792
rect 26963 5700 27029 5854
rect 26963 5636 26964 5700
rect 27028 5636 27029 5700
rect 26963 5620 27029 5636
rect 26963 5556 26964 5620
rect 27028 5556 27029 5620
rect 26963 5540 27029 5556
rect 26963 5476 26964 5540
rect 27028 5476 27029 5540
rect 26963 5460 27029 5476
rect 26963 5396 26964 5460
rect 27028 5396 27029 5460
rect 26963 5380 27029 5396
rect 26963 5316 26964 5380
rect 27028 5316 27029 5380
rect 26963 5300 27029 5316
rect 26963 5236 26964 5300
rect 27028 5236 27029 5300
rect 26963 5220 27029 5236
rect 26963 5156 26964 5220
rect 27028 5156 27029 5220
rect 26963 5140 27029 5156
rect 26963 5076 26964 5140
rect 27028 5076 27029 5140
rect 26963 5060 27029 5076
rect 26963 4996 26964 5060
rect 27028 4996 27029 5060
rect 26963 4980 27029 4996
rect 26963 4916 26964 4980
rect 27028 4916 27029 4980
rect 26963 4826 27029 4916
rect 27089 4762 27149 5792
rect 27209 4822 27269 5854
rect 27329 4762 27389 5792
rect 27449 4822 27509 5854
rect 27569 5700 27635 5854
rect 27569 5636 27570 5700
rect 27634 5636 27635 5700
rect 27569 5620 27635 5636
rect 27569 5556 27570 5620
rect 27634 5556 27635 5620
rect 27569 5540 27635 5556
rect 27569 5476 27570 5540
rect 27634 5476 27635 5540
rect 27569 5460 27635 5476
rect 27569 5396 27570 5460
rect 27634 5396 27635 5460
rect 27569 5380 27635 5396
rect 27569 5316 27570 5380
rect 27634 5316 27635 5380
rect 27569 5300 27635 5316
rect 27569 5236 27570 5300
rect 27634 5236 27635 5300
rect 27569 5220 27635 5236
rect 27569 5156 27570 5220
rect 27634 5156 27635 5220
rect 27569 5140 27635 5156
rect 27569 5076 27570 5140
rect 27634 5076 27635 5140
rect 27569 5060 27635 5076
rect 27569 4996 27570 5060
rect 27634 4996 27635 5060
rect 27569 4980 27635 4996
rect 27569 4916 27570 4980
rect 27634 4916 27635 4980
rect 27569 4826 27635 4916
rect 27695 4822 27755 5854
rect 27815 4762 27875 5792
rect 27935 4822 27995 5854
rect 28055 4762 28115 5792
rect 28175 5700 28241 5854
rect 28175 5636 28176 5700
rect 28240 5636 28241 5700
rect 28175 5620 28241 5636
rect 28175 5556 28176 5620
rect 28240 5556 28241 5620
rect 28175 5540 28241 5556
rect 28175 5476 28176 5540
rect 28240 5476 28241 5540
rect 28175 5460 28241 5476
rect 28175 5396 28176 5460
rect 28240 5396 28241 5460
rect 28175 5380 28241 5396
rect 28175 5316 28176 5380
rect 28240 5316 28241 5380
rect 28175 5300 28241 5316
rect 28175 5236 28176 5300
rect 28240 5236 28241 5300
rect 28175 5220 28241 5236
rect 28175 5156 28176 5220
rect 28240 5156 28241 5220
rect 28175 5140 28241 5156
rect 28175 5076 28176 5140
rect 28240 5076 28241 5140
rect 28175 5060 28241 5076
rect 28175 4996 28176 5060
rect 28240 4996 28241 5060
rect 28175 4980 28241 4996
rect 28175 4916 28176 4980
rect 28240 4916 28241 4980
rect 28175 4826 28241 4916
rect 28301 5920 29579 5922
rect 28301 5856 28405 5920
rect 28469 5856 28485 5920
rect 28549 5856 28565 5920
rect 28629 5856 28645 5920
rect 28709 5856 28725 5920
rect 28789 5856 28805 5920
rect 28869 5856 29011 5920
rect 29075 5856 29091 5920
rect 29155 5856 29171 5920
rect 29235 5856 29251 5920
rect 29315 5856 29331 5920
rect 29395 5856 29411 5920
rect 29475 5856 29579 5920
rect 28301 5854 29579 5856
rect 28301 5700 28367 5854
rect 28301 5636 28302 5700
rect 28366 5636 28367 5700
rect 28301 5620 28367 5636
rect 28301 5556 28302 5620
rect 28366 5556 28367 5620
rect 28301 5540 28367 5556
rect 28301 5476 28302 5540
rect 28366 5476 28367 5540
rect 28301 5460 28367 5476
rect 28301 5396 28302 5460
rect 28366 5396 28367 5460
rect 28301 5380 28367 5396
rect 28301 5316 28302 5380
rect 28366 5316 28367 5380
rect 28301 5300 28367 5316
rect 28301 5236 28302 5300
rect 28366 5236 28367 5300
rect 28301 5220 28367 5236
rect 28301 5156 28302 5220
rect 28366 5156 28367 5220
rect 28301 5140 28367 5156
rect 28301 5076 28302 5140
rect 28366 5076 28367 5140
rect 28301 5060 28367 5076
rect 28301 4996 28302 5060
rect 28366 4996 28367 5060
rect 28301 4980 28367 4996
rect 28301 4916 28302 4980
rect 28366 4916 28367 4980
rect 28301 4826 28367 4916
rect 28427 4762 28487 5792
rect 28547 4822 28607 5854
rect 28667 4762 28727 5792
rect 28787 4822 28847 5854
rect 28907 5700 28973 5854
rect 28907 5636 28908 5700
rect 28972 5636 28973 5700
rect 28907 5620 28973 5636
rect 28907 5556 28908 5620
rect 28972 5556 28973 5620
rect 28907 5540 28973 5556
rect 28907 5476 28908 5540
rect 28972 5476 28973 5540
rect 28907 5460 28973 5476
rect 28907 5396 28908 5460
rect 28972 5396 28973 5460
rect 28907 5380 28973 5396
rect 28907 5316 28908 5380
rect 28972 5316 28973 5380
rect 28907 5300 28973 5316
rect 28907 5236 28908 5300
rect 28972 5236 28973 5300
rect 28907 5220 28973 5236
rect 28907 5156 28908 5220
rect 28972 5156 28973 5220
rect 28907 5140 28973 5156
rect 28907 5076 28908 5140
rect 28972 5076 28973 5140
rect 28907 5060 28973 5076
rect 28907 4996 28908 5060
rect 28972 4996 28973 5060
rect 28907 4980 28973 4996
rect 28907 4916 28908 4980
rect 28972 4916 28973 4980
rect 28907 4826 28973 4916
rect 29033 4822 29093 5854
rect 29153 4762 29213 5792
rect 29273 4822 29333 5854
rect 29393 4762 29453 5792
rect 29513 5700 29579 5854
rect 29513 5636 29514 5700
rect 29578 5636 29579 5700
rect 29513 5620 29579 5636
rect 29513 5556 29514 5620
rect 29578 5556 29579 5620
rect 29513 5540 29579 5556
rect 29513 5476 29514 5540
rect 29578 5476 29579 5540
rect 29513 5460 29579 5476
rect 29513 5396 29514 5460
rect 29578 5396 29579 5460
rect 29513 5380 29579 5396
rect 29513 5316 29514 5380
rect 29578 5316 29579 5380
rect 29513 5300 29579 5316
rect 29513 5236 29514 5300
rect 29578 5236 29579 5300
rect 29513 5220 29579 5236
rect 29513 5156 29514 5220
rect 29578 5156 29579 5220
rect 29513 5140 29579 5156
rect 29513 5076 29514 5140
rect 29578 5076 29579 5140
rect 29513 5060 29579 5076
rect 29513 4996 29514 5060
rect 29578 4996 29579 5060
rect 29513 4980 29579 4996
rect 29513 4916 29514 4980
rect 29578 4916 29579 4980
rect 29513 4826 29579 4916
rect 29641 5920 30313 5922
rect 29641 5856 29745 5920
rect 29809 5856 29825 5920
rect 29889 5856 29905 5920
rect 29969 5856 29985 5920
rect 30049 5856 30065 5920
rect 30129 5856 30145 5920
rect 30209 5856 30313 5920
rect 29641 5854 30313 5856
rect 29641 5700 29707 5854
rect 29641 5636 29642 5700
rect 29706 5636 29707 5700
rect 29641 5620 29707 5636
rect 29641 5556 29642 5620
rect 29706 5556 29707 5620
rect 29641 5540 29707 5556
rect 29641 5476 29642 5540
rect 29706 5476 29707 5540
rect 29641 5460 29707 5476
rect 29641 5396 29642 5460
rect 29706 5396 29707 5460
rect 29641 5380 29707 5396
rect 29641 5316 29642 5380
rect 29706 5316 29707 5380
rect 29641 5300 29707 5316
rect 29641 5236 29642 5300
rect 29706 5236 29707 5300
rect 29641 5220 29707 5236
rect 29641 5156 29642 5220
rect 29706 5156 29707 5220
rect 29641 5140 29707 5156
rect 29641 5076 29642 5140
rect 29706 5076 29707 5140
rect 29641 5060 29707 5076
rect 29641 4996 29642 5060
rect 29706 4996 29707 5060
rect 29641 4980 29707 4996
rect 29641 4916 29642 4980
rect 29706 4916 29707 4980
rect 29641 4826 29707 4916
rect 29767 4822 29827 5854
rect 29887 4762 29947 5792
rect 30007 4822 30067 5854
rect 30127 4762 30187 5792
rect 30247 5700 30313 5854
rect 30247 5636 30248 5700
rect 30312 5636 30313 5700
rect 30247 5620 30313 5636
rect 30247 5556 30248 5620
rect 30312 5556 30313 5620
rect 30247 5540 30313 5556
rect 30247 5476 30248 5540
rect 30312 5476 30313 5540
rect 30247 5460 30313 5476
rect 30247 5396 30248 5460
rect 30312 5396 30313 5460
rect 30247 5380 30313 5396
rect 30247 5316 30248 5380
rect 30312 5316 30313 5380
rect 30247 5300 30313 5316
rect 30247 5236 30248 5300
rect 30312 5236 30313 5300
rect 30247 5220 30313 5236
rect 30247 5156 30248 5220
rect 30312 5156 30313 5220
rect 30247 5140 30313 5156
rect 30247 5076 30248 5140
rect 30312 5076 30313 5140
rect 30247 5060 30313 5076
rect 30247 4996 30248 5060
rect 30312 4996 30313 5060
rect 30247 4980 30313 4996
rect 30247 4916 30248 4980
rect 30312 4916 30313 4980
rect 30247 4826 30313 4916
rect 30374 5810 30434 6073
rect 30632 5954 30692 6332
rect 30494 5944 30692 5954
rect 30494 5880 30495 5944
rect 30559 5880 30692 5944
rect 30494 5870 30692 5880
rect 30752 6352 30784 6353
rect 30848 6352 30984 6416
rect 31048 6352 31248 6416
rect 30374 5774 30690 5810
rect 30374 5710 30595 5774
rect 30659 5710 30690 5774
rect 30374 5692 30690 5710
rect 30374 5682 30692 5692
rect 30374 5618 30404 5682
rect 30468 5618 30692 5682
rect 25019 4761 25691 4762
rect 25751 4761 28241 4762
rect 28301 4761 29579 4762
rect 29641 4761 30313 4762
rect 30374 4761 30692 5618
rect 24071 4760 30692 4761
rect 24071 4757 25203 4760
rect 24071 4693 24661 4757
rect 24725 4696 25203 4757
rect 25267 4696 25283 4760
rect 25347 4696 25363 4760
rect 25427 4696 25443 4760
rect 25507 4696 25935 4760
rect 25999 4696 26015 4760
rect 26079 4696 26095 4760
rect 26159 4696 26175 4760
rect 26239 4696 26541 4760
rect 26605 4696 26621 4760
rect 26685 4696 26701 4760
rect 26765 4696 26781 4760
rect 26845 4696 27147 4760
rect 27211 4696 27227 4760
rect 27291 4696 27307 4760
rect 27371 4696 27387 4760
rect 27451 4696 27753 4760
rect 27817 4696 27833 4760
rect 27897 4696 27913 4760
rect 27977 4696 27993 4760
rect 28057 4696 28485 4760
rect 28549 4696 28565 4760
rect 28629 4696 28645 4760
rect 28709 4696 28725 4760
rect 28789 4696 29091 4760
rect 29155 4696 29171 4760
rect 29235 4696 29251 4760
rect 29315 4696 29331 4760
rect 29395 4696 29825 4760
rect 29889 4696 29905 4760
rect 29969 4696 29985 4760
rect 30049 4696 30065 4760
rect 30129 4696 30692 4760
rect 24725 4693 30692 4696
rect 24071 4683 30692 4693
rect 24071 4546 30361 4683
rect 23357 4319 30361 4546
rect 23357 4318 29104 4319
rect 23357 4315 26740 4318
rect 23357 4313 26308 4315
rect 23357 4312 26107 4313
rect 23357 4248 25708 4312
rect 25772 4311 26107 4312
rect 25772 4248 25882 4311
rect 23357 4247 25882 4248
rect 25946 4249 26107 4311
rect 26171 4251 26308 4313
rect 26372 4313 26740 4315
rect 26372 4251 26531 4313
rect 26171 4249 26531 4251
rect 26595 4254 26740 4313
rect 26804 4315 27363 4318
rect 26804 4311 27158 4315
rect 26804 4254 26968 4311
rect 26595 4249 26968 4254
rect 25946 4247 26968 4249
rect 27032 4251 27158 4311
rect 27222 4254 27363 4315
rect 27427 4254 27562 4318
rect 27626 4313 28166 4318
rect 27626 4254 27778 4313
rect 27222 4251 27778 4254
rect 27032 4249 27778 4251
rect 27842 4254 28166 4313
rect 28230 4316 29104 4318
rect 28230 4315 28875 4316
rect 28230 4313 28643 4315
rect 28230 4254 28401 4313
rect 27842 4249 28401 4254
rect 28465 4251 28643 4313
rect 28707 4252 28875 4315
rect 28939 4255 29104 4316
rect 29168 4318 30361 4319
rect 29168 4315 30237 4318
rect 29168 4311 29571 4315
rect 29168 4255 29353 4311
rect 28939 4252 29353 4255
rect 28707 4251 29353 4252
rect 28465 4249 29353 4251
rect 27032 4247 29353 4249
rect 29417 4251 29571 4311
rect 29635 4313 30237 4315
rect 29635 4311 30021 4313
rect 29635 4251 29800 4311
rect 29417 4247 29800 4251
rect 29864 4249 30021 4311
rect 30085 4254 30237 4313
rect 30301 4254 30361 4318
rect 30085 4249 30361 4254
rect 29864 4247 30361 4249
rect 23357 4198 30361 4247
rect 23357 4088 24814 4198
rect 23357 3942 23605 4088
rect 23755 3942 24814 4088
rect 23357 3834 24814 3942
rect 24978 3834 25474 4198
rect 27043 4125 27157 4138
rect 27043 4068 27066 4125
rect 23357 3643 25474 3834
rect 23357 3431 24798 3643
rect 24978 3431 25474 3643
rect 25537 4061 27066 4068
rect 27130 4068 27157 4125
rect 29438 4124 29552 4137
rect 27428 4074 27542 4087
rect 27428 4068 27451 4074
rect 27130 4061 27451 4068
rect 25537 4010 27451 4061
rect 27515 4068 27542 4074
rect 29438 4068 29461 4124
rect 27515 4060 29461 4068
rect 29525 4068 29552 4124
rect 29823 4075 29937 4088
rect 29823 4068 29846 4075
rect 29525 4060 29846 4068
rect 27515 4011 29846 4060
rect 29910 4068 29937 4075
rect 30752 4068 31248 6352
rect 29910 4011 31250 4068
rect 27515 4010 31250 4011
rect 25537 3863 31250 4010
rect 25537 3735 31249 3863
rect 25537 3732 26757 3735
rect 25537 3729 26301 3732
rect 25537 3665 25710 3729
rect 25774 3727 26082 3729
rect 25774 3665 25885 3727
rect 25537 3663 25885 3665
rect 25949 3665 26082 3727
rect 26146 3668 26301 3729
rect 26365 3728 26757 3732
rect 26365 3668 26533 3728
rect 26146 3665 26533 3668
rect 25949 3664 26533 3665
rect 26597 3671 26757 3728
rect 26821 3726 31249 3735
rect 26821 3725 30186 3726
rect 26821 3723 29964 3725
rect 26821 3671 26969 3723
rect 26597 3664 26969 3671
rect 25949 3663 26969 3664
rect 25537 3659 26969 3663
rect 27033 3719 29964 3723
rect 27033 3659 27191 3719
rect 25537 3655 27191 3659
rect 27255 3718 29964 3719
rect 27255 3716 28928 3718
rect 27255 3655 27414 3716
rect 25537 3652 27414 3655
rect 27478 3652 27624 3716
rect 27688 3652 27837 3716
rect 27901 3714 28928 3716
rect 27901 3713 28736 3714
rect 27901 3712 28557 3713
rect 27901 3709 28356 3712
rect 27901 3652 28154 3709
rect 25537 3645 28154 3652
rect 28218 3648 28356 3709
rect 28420 3649 28557 3712
rect 28621 3650 28736 3713
rect 28800 3654 28928 3714
rect 28992 3716 29756 3718
rect 28992 3715 29550 3716
rect 28992 3654 29113 3715
rect 28800 3651 29113 3654
rect 29177 3714 29550 3715
rect 29177 3651 29345 3714
rect 28800 3650 29345 3651
rect 29409 3652 29550 3714
rect 29614 3654 29756 3716
rect 29820 3661 29964 3718
rect 30028 3662 30186 3725
rect 30250 3662 31249 3726
rect 30028 3661 31249 3662
rect 29820 3654 31249 3661
rect 29614 3652 31249 3654
rect 29409 3650 31249 3652
rect 28621 3649 31249 3650
rect 28420 3648 31249 3649
rect 28218 3645 31249 3648
rect 25537 3583 31249 3645
rect 23357 3421 25474 3431
rect 23357 3410 30400 3421
rect 23357 3264 23611 3410
rect 23761 3264 30400 3410
rect 8122 2503 10581 2660
rect 8122 -1451 8351 2503
rect 10751 2451 13822 3164
rect 23357 3152 30400 3264
rect 23435 3150 30400 3152
rect 23794 3120 30400 3150
rect 24978 3089 30400 3120
rect 24978 3086 29080 3089
rect 24978 3085 26159 3086
rect 24978 3080 25953 3085
rect 24978 3016 25737 3080
rect 25801 3021 25953 3080
rect 26017 3022 26159 3085
rect 26223 3083 28857 3086
rect 26223 3082 28412 3083
rect 26223 3080 26782 3082
rect 26223 3078 26557 3080
rect 26223 3022 26361 3078
rect 26017 3021 26361 3022
rect 25801 3016 26361 3021
rect 24978 3014 26361 3016
rect 26425 3016 26557 3078
rect 26621 3018 26782 3080
rect 26846 3081 27880 3082
rect 26846 3078 27440 3081
rect 26846 3018 26997 3078
rect 26621 3016 26997 3018
rect 26425 3014 26997 3016
rect 27061 3014 27232 3078
rect 27296 3017 27440 3078
rect 27504 3017 27682 3081
rect 27746 3018 27880 3081
rect 27944 3018 28187 3082
rect 28251 3019 28412 3082
rect 28476 3082 28857 3083
rect 28476 3019 28641 3082
rect 28251 3018 28641 3019
rect 28705 3022 28857 3082
rect 28921 3025 29080 3086
rect 29144 3085 30400 3089
rect 29144 3025 29304 3085
rect 28921 3022 29304 3025
rect 28705 3021 29304 3022
rect 29368 3078 30400 3085
rect 29368 3077 30182 3078
rect 29368 3074 29955 3077
rect 29368 3021 29531 3074
rect 28705 3018 29531 3021
rect 27746 3017 29531 3018
rect 27296 3014 29531 3017
rect 24978 3010 29531 3014
rect 29595 3073 29955 3074
rect 29595 3010 29744 3073
rect 24978 3009 29744 3010
rect 29808 3013 29955 3073
rect 30019 3014 30182 3077
rect 30246 3014 30400 3078
rect 30019 3013 30400 3014
rect 29808 3009 30400 3013
rect 24978 2936 30400 3009
rect 24978 2459 25474 2936
rect 27048 2851 27162 2864
rect 27048 2793 27071 2851
rect 10751 1476 13823 2451
rect 24345 2367 25474 2459
rect 24345 2207 24914 2367
rect 24978 2242 25474 2367
rect 25534 2787 27071 2793
rect 27135 2793 27162 2851
rect 29440 2853 29554 2866
rect 27431 2793 27545 2805
rect 29440 2793 29463 2853
rect 27135 2792 29463 2793
rect 27135 2787 27454 2792
rect 25534 2728 27454 2787
rect 27518 2789 29463 2792
rect 29527 2793 29554 2853
rect 29817 2799 29931 2812
rect 29817 2793 29840 2799
rect 29527 2789 29840 2793
rect 27518 2735 29840 2789
rect 29904 2793 29931 2799
rect 30752 2793 31248 3583
rect 29904 2735 31250 2793
rect 27518 2728 31250 2735
rect 25534 2611 31250 2728
rect 25534 2502 31249 2611
rect 25534 2453 31250 2502
rect 25534 2451 27840 2453
rect 25534 2449 27627 2451
rect 25534 2445 27389 2449
rect 25534 2444 26957 2445
rect 25534 2435 25988 2444
rect 25534 2371 25763 2435
rect 25827 2380 25988 2435
rect 26052 2441 26486 2444
rect 26052 2380 26265 2441
rect 25827 2377 26265 2380
rect 26329 2380 26486 2441
rect 26550 2441 26957 2444
rect 26550 2380 26731 2441
rect 26329 2377 26731 2380
rect 26795 2381 26957 2441
rect 27021 2443 27389 2445
rect 27021 2381 27169 2443
rect 26795 2379 27169 2381
rect 27233 2385 27389 2443
rect 27453 2387 27627 2449
rect 27691 2389 27840 2451
rect 27904 2444 31250 2453
rect 27904 2443 28574 2444
rect 27904 2389 28227 2443
rect 27691 2387 28227 2389
rect 27453 2385 28227 2387
rect 27233 2379 28227 2385
rect 28291 2380 28574 2443
rect 28638 2441 31250 2444
rect 28638 2439 29233 2441
rect 28638 2380 28810 2439
rect 28291 2379 28810 2380
rect 26795 2377 28810 2379
rect 25827 2375 28810 2377
rect 28874 2375 28994 2439
rect 29058 2377 29233 2439
rect 29297 2440 31250 2441
rect 29297 2437 30003 2440
rect 29297 2377 29436 2437
rect 29058 2375 29436 2377
rect 25827 2373 29436 2375
rect 29500 2436 30003 2437
rect 29500 2434 29812 2436
rect 29500 2373 29621 2434
rect 25827 2371 29621 2373
rect 25534 2370 29621 2371
rect 29685 2372 29812 2434
rect 29876 2376 30003 2436
rect 30067 2436 31250 2440
rect 30067 2376 30189 2436
rect 29876 2372 30189 2376
rect 30253 2372 31250 2436
rect 29685 2370 31250 2372
rect 25534 2308 31250 2370
rect 24978 2207 30402 2242
rect 24345 2044 30402 2207
rect 24342 1855 30402 2044
rect 24342 1854 28351 1855
rect 24342 1853 26027 1854
rect 24342 1789 25636 1853
rect 25700 1849 26027 1853
rect 25700 1789 25841 1849
rect 24342 1785 25841 1789
rect 25905 1790 26027 1849
rect 26091 1852 28351 1854
rect 26091 1847 26440 1852
rect 26091 1790 26221 1847
rect 25905 1785 26221 1790
rect 24342 1783 26221 1785
rect 26285 1788 26440 1847
rect 26504 1788 26650 1852
rect 26714 1849 28133 1852
rect 26714 1788 26879 1849
rect 26285 1785 26879 1788
rect 26943 1785 27125 1849
rect 27189 1785 27399 1849
rect 27463 1785 27674 1849
rect 27738 1785 27910 1849
rect 27974 1788 28133 1849
rect 28197 1791 28351 1852
rect 28415 1853 30402 1855
rect 28415 1849 29796 1853
rect 28415 1848 29376 1849
rect 28415 1846 28768 1848
rect 28415 1791 28529 1846
rect 28197 1788 28529 1791
rect 27974 1785 28529 1788
rect 26285 1783 28529 1785
rect 24342 1782 28529 1783
rect 28593 1784 28768 1846
rect 28832 1784 28965 1848
rect 29029 1784 29163 1848
rect 29227 1785 29376 1848
rect 29440 1848 29796 1849
rect 29440 1785 29599 1848
rect 29227 1784 29599 1785
rect 29663 1789 29796 1848
rect 29860 1851 30402 1853
rect 29860 1789 30012 1851
rect 29663 1787 30012 1789
rect 30076 1787 30221 1851
rect 30285 1787 30402 1851
rect 29663 1784 30402 1787
rect 28593 1782 30402 1784
rect 24342 1757 30402 1782
rect 24342 1532 25452 1757
rect 8431 1453 15853 1476
rect 8431 1421 24265 1453
rect 8431 1419 9834 1421
rect 8431 1417 8824 1419
rect 8431 1353 8622 1417
rect 8686 1355 8824 1417
rect 8888 1417 9433 1419
rect 8888 1355 9035 1417
rect 8686 1353 9035 1355
rect 9099 1353 9225 1417
rect 9289 1355 9433 1417
rect 9497 1355 9635 1419
rect 9699 1357 9834 1419
rect 9898 1420 10721 1421
rect 9898 1418 10230 1420
rect 9898 1357 10029 1418
rect 9699 1355 10029 1357
rect 9289 1354 10029 1355
rect 10093 1356 10230 1418
rect 10294 1418 10721 1420
rect 10294 1356 10447 1418
rect 10093 1354 10447 1356
rect 10511 1357 10721 1418
rect 10785 1417 24265 1421
rect 10785 1414 11221 1417
rect 10785 1357 10998 1414
rect 10511 1354 10998 1357
rect 9289 1353 10998 1354
rect 8431 1350 10998 1353
rect 11062 1353 11221 1414
rect 11285 1416 24265 1417
rect 11285 1353 11453 1416
rect 11062 1352 11453 1353
rect 11517 1415 14472 1416
rect 11517 1414 13597 1415
rect 11517 1413 13397 1414
rect 11517 1352 13089 1413
rect 11062 1350 13089 1352
rect 8431 1349 13089 1350
rect 13153 1350 13397 1413
rect 13461 1351 13597 1414
rect 13661 1414 14270 1415
rect 13661 1351 13816 1414
rect 13461 1350 13816 1351
rect 13880 1413 14270 1414
rect 13880 1350 14062 1413
rect 13153 1349 14062 1350
rect 14126 1351 14270 1413
rect 14334 1352 14472 1415
rect 14536 1415 24265 1416
rect 14536 1352 14665 1415
rect 14334 1351 14665 1352
rect 14729 1414 24265 1415
rect 14729 1351 15037 1414
rect 14126 1350 15037 1351
rect 15101 1412 15789 1414
rect 15101 1350 15226 1412
rect 14126 1349 15226 1350
rect 8431 1348 15226 1349
rect 15290 1348 15516 1412
rect 15580 1350 15789 1412
rect 15853 1350 24265 1414
rect 15580 1348 24265 1350
rect 8431 1156 24265 1348
rect 8431 273 9605 1156
rect 8431 209 8588 273
rect 8652 271 9605 273
rect 8652 209 8828 271
rect 8431 207 8828 209
rect 8892 270 9368 271
rect 8892 207 9150 270
rect 8431 206 9150 207
rect 9214 207 9368 270
rect 9432 207 9605 271
rect 9214 206 9605 207
rect 8431 -410 9605 206
rect 8431 -474 8834 -410
rect 8898 -414 9605 -410
rect 8898 -474 9036 -414
rect 8431 -478 9036 -474
rect 9100 -416 9605 -414
rect 9100 -417 9454 -416
rect 9100 -478 9225 -417
rect 8431 -481 9225 -478
rect 9289 -480 9454 -417
rect 9518 -480 9605 -416
rect 9289 -481 9605 -480
rect 8431 -1100 9605 -481
rect 8431 -1103 9064 -1100
rect 8431 -1167 8616 -1103
rect 8680 -1107 9064 -1103
rect 8680 -1167 8849 -1107
rect 8431 -1171 8849 -1167
rect 8913 -1164 9064 -1107
rect 9128 -1102 9605 -1100
rect 9128 -1103 9498 -1102
rect 9128 -1164 9282 -1103
rect 8913 -1167 9282 -1164
rect 9346 -1166 9498 -1103
rect 9562 -1166 9605 -1102
rect 9346 -1167 9605 -1166
rect 8913 -1171 9605 -1167
rect 8431 -1370 9605 -1171
rect 9685 882 11071 1075
rect 9685 878 9959 882
rect 9685 814 9740 878
rect 9804 818 9959 878
rect 10023 818 10242 882
rect 10306 818 10451 882
rect 10515 880 11071 882
rect 10515 818 10722 880
rect 9804 816 10722 818
rect 10786 816 11071 880
rect 9804 814 11071 816
rect 9685 -265 11071 814
rect 9685 -329 9779 -265
rect 9843 -329 9996 -265
rect 10060 -329 10215 -265
rect 10279 -269 11071 -265
rect 10279 -329 10428 -269
rect 9685 -333 10428 -329
rect 10492 -333 10639 -269
rect 10703 -333 11071 -269
rect 9685 -947 11071 -333
rect 9685 -959 9990 -947
rect 9685 -1023 9761 -959
rect 9825 -1011 9990 -959
rect 10054 -953 11071 -947
rect 10054 -957 10401 -953
rect 10054 -1011 10209 -957
rect 9825 -1021 10209 -1011
rect 10273 -1017 10401 -957
rect 10465 -955 11071 -953
rect 10465 -1017 10895 -955
rect 10273 -1019 10895 -1017
rect 10959 -1019 11071 -955
rect 10273 -1021 11071 -1019
rect 9825 -1023 11071 -1021
rect 9685 -1451 11071 -1023
rect 11151 277 12537 1156
rect 11151 275 11597 277
rect 11151 211 11272 275
rect 11336 213 11597 275
rect 11661 213 11865 277
rect 11929 213 12131 277
rect 12195 275 12537 277
rect 12195 213 12371 275
rect 11336 211 12371 213
rect 12435 211 12537 275
rect 11151 -409 12537 211
rect 11151 -413 11831 -409
rect 11151 -477 11223 -413
rect 11287 -416 11831 -413
rect 11287 -477 11438 -416
rect 11151 -480 11438 -477
rect 11502 -419 11831 -416
rect 11502 -480 11636 -419
rect 11151 -483 11636 -480
rect 11700 -473 11831 -419
rect 11895 -411 12537 -409
rect 11895 -473 12111 -411
rect 11700 -475 12111 -473
rect 12175 -413 12537 -411
rect 12175 -475 12330 -413
rect 11700 -477 12330 -475
rect 12394 -477 12537 -413
rect 11700 -483 12537 -477
rect 11151 -1098 12537 -483
rect 11151 -1103 12355 -1098
rect 11151 -1106 11619 -1103
rect 11151 -1170 11219 -1106
rect 11283 -1170 11409 -1106
rect 11473 -1167 11619 -1106
rect 11683 -1106 12131 -1103
rect 11683 -1167 11836 -1106
rect 11473 -1170 11836 -1167
rect 11900 -1167 12131 -1106
rect 12195 -1162 12355 -1103
rect 12419 -1162 12537 -1098
rect 12195 -1167 12537 -1162
rect 11900 -1170 12537 -1167
rect 11151 -1370 12537 -1170
rect 12617 881 14003 1075
rect 12617 878 13046 881
rect 12617 814 12797 878
rect 12861 817 13046 878
rect 13110 873 14003 881
rect 13110 867 13644 873
rect 13110 817 13390 867
rect 12861 814 13390 817
rect 12617 803 13390 814
rect 13454 809 13644 867
rect 13708 809 13873 873
rect 13937 809 14003 873
rect 13454 803 14003 809
rect 12617 -265 14003 803
rect 12617 -269 13613 -265
rect 12617 -333 12763 -269
rect 12827 -270 13613 -269
rect 12827 -333 13041 -270
rect 12617 -334 13041 -333
rect 13105 -329 13613 -270
rect 13677 -329 13852 -265
rect 13916 -329 14003 -265
rect 13105 -334 14003 -329
rect 12617 -948 14003 -334
rect 12617 -950 13607 -948
rect 12617 -956 13277 -950
rect 12617 -1020 12687 -956
rect 12751 -958 13277 -956
rect 12751 -1020 13080 -958
rect 12617 -1022 13080 -1020
rect 13144 -1014 13277 -958
rect 13341 -1012 13607 -950
rect 13671 -1012 13803 -948
rect 13867 -1012 14003 -948
rect 13341 -1014 14003 -1012
rect 13144 -1022 14003 -1014
rect 12617 -1451 14003 -1022
rect 14083 281 15469 1156
rect 14083 278 14531 281
rect 14083 214 14165 278
rect 14229 217 14531 278
rect 14595 217 14775 281
rect 14839 272 15469 281
rect 14839 217 15198 272
rect 14229 214 15198 217
rect 14083 208 15198 214
rect 15262 208 15469 272
rect 14083 -412 15469 208
rect 14083 -414 15087 -412
rect 14083 -416 14896 -414
rect 14083 -480 14151 -416
rect 14215 -419 14896 -416
rect 14215 -480 14502 -419
rect 14083 -483 14502 -480
rect 14566 -421 14896 -419
rect 14566 -483 14691 -421
rect 14083 -485 14691 -483
rect 14755 -478 14896 -421
rect 14960 -476 15087 -414
rect 15151 -476 15469 -412
rect 14960 -478 15469 -476
rect 14755 -485 15469 -478
rect 14083 -1098 15469 -485
rect 14083 -1103 15002 -1098
rect 14083 -1105 14785 -1103
rect 14083 -1169 14233 -1105
rect 14297 -1107 14785 -1105
rect 14297 -1169 14533 -1107
rect 14083 -1171 14533 -1169
rect 14597 -1167 14785 -1107
rect 14849 -1162 15002 -1103
rect 15066 -1101 15469 -1098
rect 15066 -1162 15203 -1101
rect 14849 -1165 15203 -1162
rect 15267 -1165 15469 -1101
rect 14849 -1167 15469 -1165
rect 14597 -1171 15469 -1167
rect 14083 -1371 15469 -1171
rect 15549 880 16935 1075
rect 15549 878 15795 880
rect 15549 814 15591 878
rect 15655 816 15795 878
rect 15859 878 16935 880
rect 15859 816 16118 878
rect 15655 814 16118 816
rect 16182 814 16935 878
rect 15549 -260 16935 814
rect 15549 -262 16427 -260
rect 15549 -267 16237 -262
rect 15549 -331 16010 -267
rect 16074 -326 16237 -267
rect 16301 -324 16427 -262
rect 16491 -269 16935 -260
rect 16491 -324 16643 -269
rect 16301 -326 16643 -324
rect 16074 -331 16643 -326
rect 15549 -333 16643 -331
rect 16707 -333 16935 -269
rect 15549 -948 16935 -333
rect 15549 -950 16638 -948
rect 15549 -951 16217 -950
rect 15549 -955 16011 -951
rect 15549 -1019 15710 -955
rect 15774 -1015 16011 -955
rect 16075 -1014 16217 -951
rect 16281 -954 16638 -950
rect 16281 -1014 16427 -954
rect 16075 -1015 16427 -1014
rect 15774 -1018 16427 -1015
rect 16491 -1012 16638 -954
rect 16702 -1012 16935 -948
rect 16491 -1018 16935 -1012
rect 15774 -1019 16935 -1018
rect 15549 -1451 16935 -1019
rect 17015 279 18401 1156
rect 17015 274 17599 279
rect 17015 210 17141 274
rect 17205 271 17599 274
rect 17205 210 17393 271
rect 17015 207 17393 210
rect 17457 215 17599 271
rect 17663 274 18401 279
rect 17663 273 18180 274
rect 17663 215 17882 273
rect 17457 209 17882 215
rect 17946 210 18180 273
rect 18244 210 18401 274
rect 17946 209 18401 210
rect 17457 207 18401 209
rect 17015 -408 18401 207
rect 17015 -410 17322 -408
rect 17015 -474 17132 -410
rect 17196 -472 17322 -410
rect 17386 -410 18401 -408
rect 17386 -472 17516 -410
rect 17196 -474 17516 -472
rect 17580 -414 18401 -410
rect 17580 -474 17827 -414
rect 17015 -478 17827 -474
rect 17891 -478 18401 -414
rect 17015 -1102 18401 -478
rect 17015 -1110 18098 -1102
rect 17015 -1174 17088 -1110
rect 17152 -1174 17280 -1110
rect 17344 -1174 17480 -1110
rect 17544 -1166 18098 -1110
rect 18162 -1166 18401 -1102
rect 17544 -1174 18401 -1166
rect 17015 -1370 18401 -1174
rect 18481 -258 19867 1076
rect 18481 -263 19079 -258
rect 18481 -266 18853 -263
rect 18481 -330 18624 -266
rect 18688 -327 18853 -266
rect 18917 -322 19079 -263
rect 19143 -260 19867 -258
rect 19143 -266 19543 -260
rect 19143 -322 19307 -266
rect 18917 -327 19307 -322
rect 18688 -330 19307 -327
rect 19371 -324 19543 -266
rect 19607 -269 19867 -260
rect 19607 -324 19735 -269
rect 19371 -330 19735 -324
rect 18481 -333 19735 -330
rect 19799 -333 19867 -269
rect 18481 -948 19867 -333
rect 18481 -951 19537 -948
rect 18481 -952 19296 -951
rect 18481 -959 18775 -952
rect 18481 -1023 18518 -959
rect 18582 -1016 18775 -959
rect 18839 -956 19296 -952
rect 18839 -1016 19025 -956
rect 18582 -1020 19025 -1016
rect 19089 -1015 19296 -956
rect 19360 -1012 19537 -951
rect 19601 -952 19867 -948
rect 19601 -1012 19762 -952
rect 19360 -1015 19762 -1012
rect 19089 -1016 19762 -1015
rect 19826 -1016 19867 -952
rect 19089 -1020 19867 -1016
rect 18582 -1023 19867 -1020
rect 18481 -1451 19867 -1023
rect 19947 277 21333 1156
rect 19947 275 20222 277
rect 19947 211 20012 275
rect 20076 213 20222 275
rect 20286 275 21333 277
rect 20286 213 20573 275
rect 20076 211 20573 213
rect 20637 211 20853 275
rect 20917 274 21333 275
rect 20917 211 21170 274
rect 19947 210 21170 211
rect 21234 210 21333 274
rect 19947 -415 21333 210
rect 19947 -479 20010 -415
rect 20074 -479 20214 -415
rect 20278 -417 21333 -415
rect 20278 -419 21018 -417
rect 20278 -479 20779 -419
rect 19947 -483 20779 -479
rect 20843 -481 21018 -419
rect 21082 -481 21222 -417
rect 21286 -481 21333 -417
rect 20843 -483 21333 -481
rect 19947 -1104 21333 -483
rect 19947 -1106 20779 -1104
rect 19947 -1170 19999 -1106
rect 20063 -1170 20255 -1106
rect 20319 -1170 20490 -1106
rect 20554 -1168 20779 -1106
rect 20843 -1106 21173 -1104
rect 20843 -1168 20969 -1106
rect 20554 -1170 20969 -1168
rect 21033 -1168 21173 -1106
rect 21237 -1168 21333 -1104
rect 21033 -1170 21333 -1168
rect 19947 -1370 21333 -1170
rect 21413 -264 22799 1075
rect 21413 -269 21674 -264
rect 21413 -333 21470 -269
rect 21534 -328 21674 -269
rect 21738 -269 22799 -264
rect 21738 -328 21865 -269
rect 21534 -333 21865 -328
rect 21929 -270 22357 -269
rect 21929 -333 22067 -270
rect 21413 -334 22067 -333
rect 22131 -333 22357 -270
rect 22421 -270 22799 -269
rect 22421 -333 22642 -270
rect 22131 -334 22642 -333
rect 22706 -334 22799 -270
rect 21413 -953 22799 -334
rect 21413 -954 21670 -953
rect 21413 -1018 21469 -954
rect 21533 -1017 21670 -954
rect 21734 -957 22095 -953
rect 21734 -1017 21888 -957
rect 21533 -1018 21888 -1017
rect 21413 -1021 21888 -1018
rect 21952 -1017 22095 -957
rect 22159 -954 22799 -953
rect 22159 -1017 22300 -954
rect 21952 -1018 22300 -1017
rect 22364 -958 22799 -954
rect 22364 -1018 22647 -958
rect 21952 -1021 22647 -1018
rect 21413 -1022 22647 -1021
rect 22711 -1022 22799 -958
rect 21413 -1451 22799 -1022
rect 22879 275 24265 1156
rect 24346 1446 25452 1532
rect 24346 1138 24410 1446
rect 24500 1138 25452 1446
rect 24346 1075 25452 1138
rect 22879 272 24116 275
rect 22879 208 22960 272
rect 23024 208 23255 272
rect 23319 208 23542 272
rect 23606 208 23832 272
rect 23896 211 24116 272
rect 24180 211 24265 275
rect 23896 208 24265 211
rect 22879 -409 24265 208
rect 22879 -473 23182 -409
rect 23246 -411 24111 -409
rect 23246 -473 23415 -411
rect 22879 -475 23415 -473
rect 23479 -413 23831 -411
rect 23479 -475 23622 -413
rect 22879 -477 23622 -475
rect 23686 -475 23831 -413
rect 23895 -473 24111 -411
rect 24175 -473 24265 -409
rect 23895 -475 24265 -473
rect 23686 -477 24265 -475
rect 22879 -1095 24265 -477
rect 22879 -1098 23591 -1095
rect 22879 -1162 22959 -1098
rect 23023 -1102 23591 -1098
rect 23023 -1162 23201 -1102
rect 22879 -1166 23201 -1162
rect 23265 -1103 23591 -1102
rect 23265 -1166 23401 -1103
rect 22879 -1167 23401 -1166
rect 23465 -1159 23591 -1103
rect 23655 -1097 24265 -1095
rect 23655 -1159 23812 -1097
rect 23465 -1161 23812 -1159
rect 23876 -1102 24265 -1097
rect 23876 -1161 24108 -1102
rect 23465 -1166 24108 -1161
rect 24172 -1166 24265 -1102
rect 23465 -1167 24265 -1166
rect 22879 -1370 24265 -1167
rect 24345 902 25452 1075
rect 24345 -261 25451 902
rect 24345 -265 24591 -261
rect 24345 -329 24397 -265
rect 24461 -325 24591 -265
rect 24655 -262 25451 -261
rect 24655 -264 25003 -262
rect 24655 -325 24780 -264
rect 24461 -328 24780 -325
rect 24844 -326 25003 -264
rect 25067 -326 25451 -262
rect 24844 -328 25451 -326
rect 24461 -329 25451 -328
rect 24345 -949 25451 -329
rect 24345 -951 24785 -949
rect 24345 -954 24590 -951
rect 24345 -1018 24399 -954
rect 24463 -1015 24590 -954
rect 24654 -1013 24785 -951
rect 24849 -954 25451 -949
rect 24849 -1013 25232 -954
rect 24654 -1015 25232 -1013
rect 24463 -1018 25232 -1015
rect 25296 -1018 25451 -954
rect 24345 -1451 25451 -1018
rect 8122 -1633 25451 -1451
rect 8122 -1635 10732 -1633
rect 8122 -1699 8990 -1635
rect 9054 -1638 10732 -1635
rect 9054 -1699 9189 -1638
rect 8122 -1702 9189 -1699
rect 9253 -1702 9400 -1638
rect 9464 -1702 9606 -1638
rect 9670 -1640 10308 -1638
rect 9670 -1702 9834 -1640
rect 8122 -1704 9834 -1702
rect 9898 -1704 10078 -1640
rect 10142 -1702 10308 -1640
rect 10372 -1702 10514 -1638
rect 10578 -1697 10732 -1638
rect 10796 -1636 25451 -1633
rect 10796 -1639 11143 -1636
rect 10796 -1697 10935 -1639
rect 10578 -1702 10935 -1697
rect 10142 -1703 10935 -1702
rect 10999 -1700 11143 -1639
rect 11207 -1639 12024 -1636
rect 11207 -1640 11614 -1639
rect 11207 -1700 11406 -1640
rect 10999 -1703 11406 -1700
rect 10142 -1704 11406 -1703
rect 11470 -1703 11614 -1640
rect 11678 -1642 12024 -1639
rect 11678 -1703 11824 -1642
rect 11470 -1704 11824 -1703
rect 8122 -1706 11824 -1704
rect 11888 -1700 12024 -1642
rect 12088 -1637 15904 -1636
rect 12088 -1638 12854 -1637
rect 12088 -1639 12638 -1638
rect 12088 -1700 12227 -1639
rect 11888 -1703 12227 -1700
rect 12291 -1703 12437 -1639
rect 12501 -1702 12638 -1639
rect 12702 -1701 12854 -1638
rect 12918 -1639 13781 -1637
rect 12918 -1701 13135 -1639
rect 12702 -1702 13135 -1701
rect 12501 -1703 13135 -1702
rect 13199 -1643 13781 -1639
rect 13199 -1644 13560 -1643
rect 13199 -1703 13355 -1644
rect 11888 -1706 13355 -1703
rect 8122 -1708 13355 -1706
rect 13419 -1707 13560 -1644
rect 13624 -1701 13781 -1643
rect 13845 -1638 15904 -1637
rect 13845 -1643 14626 -1638
rect 13845 -1644 14195 -1643
rect 13845 -1701 13986 -1644
rect 13624 -1707 13986 -1701
rect 13419 -1708 13986 -1707
rect 14050 -1707 14195 -1644
rect 14259 -1707 14412 -1643
rect 14476 -1702 14626 -1643
rect 14690 -1639 15701 -1638
rect 14690 -1640 15502 -1639
rect 14690 -1702 14821 -1640
rect 14476 -1704 14821 -1702
rect 14885 -1643 15218 -1640
rect 14885 -1704 15016 -1643
rect 14476 -1707 15016 -1704
rect 15080 -1704 15218 -1643
rect 15282 -1703 15502 -1640
rect 15566 -1702 15701 -1639
rect 15765 -1700 15904 -1638
rect 15968 -1637 19386 -1636
rect 15968 -1638 17603 -1637
rect 15968 -1639 16556 -1638
rect 15968 -1700 16169 -1639
rect 15765 -1702 16169 -1700
rect 15566 -1703 16169 -1702
rect 16233 -1640 16556 -1639
rect 16233 -1703 16367 -1640
rect 15282 -1704 16367 -1703
rect 16431 -1702 16556 -1640
rect 16620 -1702 16768 -1638
rect 16832 -1702 16985 -1638
rect 17049 -1642 17603 -1638
rect 17049 -1702 17190 -1642
rect 16431 -1704 17190 -1702
rect 15080 -1706 17190 -1704
rect 17254 -1706 17395 -1642
rect 17459 -1701 17603 -1642
rect 17667 -1638 19386 -1637
rect 17667 -1701 17886 -1638
rect 17459 -1702 17886 -1701
rect 17950 -1640 18764 -1638
rect 17950 -1702 18079 -1640
rect 17459 -1704 18079 -1702
rect 18143 -1642 18764 -1640
rect 18143 -1704 18305 -1642
rect 17459 -1706 18305 -1704
rect 18369 -1706 18570 -1642
rect 18634 -1702 18764 -1642
rect 18828 -1639 19386 -1638
rect 18828 -1647 19166 -1639
rect 18828 -1702 18962 -1647
rect 18634 -1706 18962 -1702
rect 15080 -1707 18962 -1706
rect 14050 -1708 18962 -1707
rect 8122 -1711 18962 -1708
rect 19026 -1703 19166 -1647
rect 19230 -1700 19386 -1639
rect 19450 -1637 25451 -1636
rect 19450 -1640 19829 -1637
rect 19450 -1700 19601 -1640
rect 19230 -1703 19601 -1700
rect 19026 -1704 19601 -1703
rect 19665 -1701 19829 -1640
rect 19893 -1638 20464 -1637
rect 19893 -1640 20271 -1638
rect 19893 -1701 20033 -1640
rect 19665 -1704 20033 -1701
rect 20097 -1702 20271 -1640
rect 20335 -1701 20464 -1638
rect 20528 -1639 25451 -1637
rect 20528 -1642 20917 -1639
rect 20528 -1701 20661 -1642
rect 20335 -1702 20661 -1701
rect 20097 -1704 20661 -1702
rect 19026 -1706 20661 -1704
rect 20725 -1703 20917 -1642
rect 20981 -1640 25451 -1639
rect 20981 -1642 22029 -1640
rect 20981 -1643 21610 -1642
rect 20981 -1703 21156 -1643
rect 20725 -1706 21156 -1703
rect 19026 -1707 21156 -1706
rect 21220 -1647 21610 -1643
rect 21220 -1707 21389 -1647
rect 19026 -1711 21389 -1707
rect 21453 -1706 21610 -1647
rect 21674 -1706 21801 -1642
rect 21865 -1704 22029 -1642
rect 22093 -1641 23080 -1640
rect 22093 -1642 22854 -1641
rect 22093 -1645 22665 -1642
rect 22093 -1704 22226 -1645
rect 21865 -1706 22226 -1704
rect 21453 -1709 22226 -1706
rect 22290 -1709 22438 -1645
rect 22502 -1706 22665 -1645
rect 22729 -1705 22854 -1642
rect 22918 -1704 23080 -1641
rect 23144 -1704 23334 -1640
rect 23398 -1641 25066 -1640
rect 23398 -1643 24066 -1641
rect 23398 -1704 23578 -1643
rect 22918 -1705 23578 -1704
rect 22729 -1706 23578 -1705
rect 22502 -1707 23578 -1706
rect 23642 -1644 24066 -1643
rect 23642 -1707 23808 -1644
rect 22502 -1708 23808 -1707
rect 23872 -1705 24066 -1644
rect 24130 -1705 24276 -1641
rect 24340 -1705 24501 -1641
rect 24565 -1644 25066 -1641
rect 24565 -1705 24720 -1644
rect 23872 -1708 24720 -1705
rect 24784 -1704 25066 -1644
rect 25130 -1643 25451 -1640
rect 25130 -1704 25265 -1643
rect 24784 -1707 25265 -1704
rect 25329 -1707 25451 -1643
rect 24784 -1708 25451 -1707
rect 22502 -1709 25451 -1708
rect 21453 -1711 25451 -1709
rect 8122 -1771 25451 -1711
<< labels >>
flabel metal1 10933 3942 10967 3977 0 FreeSans 320 0 0 0 comp_result
port 55 nsew
flabel metal2 10001 2976 10029 6744 0 FreeSans 320 0 0 0 sar_clk
port 8 nsew
flabel metal2 11750 7806 11802 7855 0 FreeSans 320 0 0 0 sample_clk_b
port 7 nsew
flabel metal1 11827 8983 11873 9018 0 FreeSans 320 0 0 0 sample_clk
port 6 nsew
flabel metal1 10869 12169 10912 12233 0 FreeSans 320 0 0 0 ext_clk
port 4 nsew
flabel metal1 2330 11810 2393 11857 0 FreeSans 320 0 0 0 ready
port 1 nsew
flabel metal4 12826 2361 13488 7539 0 FreeSans 1600 0 0 0 VDD
port 10 nsew
flabel metal4 10055 2503 10580 7673 0 FreeSans 1600 0 0 0 VSS
port 9 nsew
flabel metal1 10922 6824 10956 6858 0 FreeSans 320 0 0 0 sel_bit[0]
port 11 nsew
flabel metal1 10927 6687 10962 6722 0 FreeSans 320 0 0 0 sel_bit[1]
port 12 nsew
flabel metal1 30455 3815 30764 3863 0 FreeSans 320 0 0 0 sar_result[0]
port 20 nsew
flabel metal1 30445 4145 30754 4193 0 FreeSans 320 0 0 0 sar_result[1]
port 13 nsew
flabel metal1 30447 3516 30756 3564 0 FreeSans 320 0 0 0 sar_result[2]
port 14 nsew
flabel metal1 30461 3174 30770 3222 0 FreeSans 320 0 0 0 sar_result[3]
port 15 nsew
flabel metal1 30450 2864 30759 2912 0 FreeSans 320 0 0 0 sar_result[5]
port 16 nsew
flabel metal1 30456 2533 30765 2581 0 FreeSans 320 0 0 0 sar_result[4]
port 17 nsew
flabel metal1 30453 2237 30762 2285 0 FreeSans 320 0 0 0 sar_result[6]
port 18 nsew
flabel metal1 30451 1893 30760 1941 0 FreeSans 320 0 0 0 sar_result[7]
port 19 nsew
flabel metal1 13479 10913 13504 10941 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[2]
port 21 nsew
flabel metal1 13481 10857 13506 10885 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[1]
port 22 nsew
flabel metal1 13483 10801 13508 10829 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[0]
port 23 nsew
flabel metal1 13484 10745 13509 10773 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[6]
port 24 nsew
flabel metal1 13486 10689 13511 10717 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[5]
port 25 nsew
flabel metal1 13485 10633 13510 10661 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[4]
port 26 nsew
flabel metal1 13473 10493 13505 10605 0 FreeSans 320 0 0 0 sample_delay_offset
port 35 nsew
flabel metal1 13198 12668 13224 12702 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[3]
port 36 nsew
flabel metal1 19914 12668 19940 12702 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[7]
port 37 nsew
flabel metal1 26659 8407 26685 8441 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[11]
port 38 nsew
flabel metal1 19956 8407 19982 8441 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[15]
port 39 nsew
flabel metal1 2930 10449 4871 10477 0 FreeSans 320 0 0 0 async_setb_delay_cap_ctrl_code[2]
port 40 nsew
flabel metal1 2931 10393 7297 10421 0 FreeSans 320 0 0 0 async_setb_delay_cap_ctrl_code[1]
port 41 nsew
flabel metal1 2929 10337 8154 10365 0 FreeSans 320 0 0 0 async_setb_delay_cap_ctrl_code[0]
port 42 nsew
flabel metal1 2928 10281 8154 10309 0 FreeSans 320 0 0 0 async_resetb_delay_cap_ctrl_code[0]
port 43 nsew
flabel metal1 2932 10225 7297 10253 0 FreeSans 320 0 0 0 async_resetb_delay_cap_ctrl_code[1]
port 44 nsew
flabel metal1 2930 10169 4871 10197 0 FreeSans 320 0 0 0 async_resetb_delay_cap_ctrl_code[2]
port 45 nsew
flabel metal1 2324 12193 2356 12227 0 FreeSans 320 0 0 0 async_setb_delay_cap_ctrl_code[3]
port 46 nsew
flabel metal1 2324 8419 2366 8453 0 FreeSans 320 0 0 0 async_resetb_delay_cap_ctrl_code[3]
port 47 nsew
flabel metal2 2737 9041 2790 11605 0 FreeSans 320 0 0 0 async_delay_offset
port 48 nsew
flabel metal1 23937 6371 24075 6405 0 FreeSans 320 0 0 0 retimer_delay_code[3]
port 50 nsew
flabel metal1 25545 4635 26484 4663 0 FreeSans 320 0 0 0 retimer_delay_code[2]
port 51 nsew
flabel metal1 25545 4579 28910 4607 0 FreeSans 320 0 0 0 retimer_delay_code[1]
port 52 nsew
flabel metal1 25545 4523 29767 4551 0 FreeSans 320 0 0 0 retimer_delay_code[0]
port 54 nsew
flabel metal2 8716 -1261 8758 2925 0 FreeSans 320 0 0 0 vss_sw[7]
port 56 nsew
flabel metal2 8798 1577 8840 2925 0 FreeSans 320 0 0 0 vss_sw[6]
port 57 nsew
flabel metal2 8882 1647 8924 2925 0 FreeSans 320 0 0 0 vss_sw[5]
port 58 nsew
flabel metal2 8970 1716 9012 2925 0 FreeSans 320 0 0 0 vss_sw[4]
port 59 nsew
flabel metal2 9057 1786 9099 2925 0 FreeSans 320 0 0 0 vss_sw[3]
port 60 nsew
flabel metal2 9143 1855 9185 2925 0 FreeSans 320 0 0 0 vss_sw[2]
port 61 nsew
flabel metal2 9229 1925 9271 2925 0 FreeSans 320 0 0 0 vss_sw[1]
port 62 nsew
flabel metal2 9316 1995 9358 2925 0 FreeSans 320 0 0 0 vdd_sw[7]
port 63 nsew
flabel metal2 9402 2065 9444 2925 0 FreeSans 320 0 0 0 vdd_sw[6]
port 64 nsew
flabel metal2 9488 2134 9530 2925 0 FreeSans 320 0 0 0 vdd_sw[5]
port 65 nsew
flabel metal2 9575 2204 9617 2925 0 FreeSans 320 0 0 0 vdd_sw[4]
port 66 nsew
flabel metal2 9660 2274 9702 2925 0 FreeSans 320 0 0 0 vdd_sw[3]
port 67 nsew
flabel metal2 9747 2343 9789 2925 0 FreeSans 320 0 0 0 vdd_sw[2]
port 68 nsew
flabel metal2 9834 2412 9876 2925 0 FreeSans 320 0 0 0 vdd_sw[1]
port 69 nsew
flabel metal2 8876 -1908 8918 -1331 0 FreeSans 320 0 0 0 vss_sw_b[7]
port 70 nsew
flabel metal2 11268 -1908 11310 -1331 0 FreeSans 320 0 0 0 vss_sw_b[6]
port 71 nsew
flabel metal2 13659 -1908 13701 -1331 0 FreeSans 320 0 0 0 vss_sw_b[5]
port 72 nsew
flabel metal2 16052 -1908 16094 -1331 0 FreeSans 320 0 0 0 vss_sw_b[4]
port 73 nsew
flabel metal2 18444 -1908 18486 -1331 0 FreeSans 320 0 0 0 vss_sw_b[3]
port 74 nsew
flabel metal2 20835 -1908 20877 -1330 0 FreeSans 320 0 0 0 vss_sw_b[2]
port 75 nsew
flabel metal2 23228 -1908 23270 -1331 0 FreeSans 320 0 0 0 vss_sw_b[1]
port 76 nsew
flabel metal2 24974 -1908 25016 -650 0 FreeSans 320 0 0 0 vdd_sw_b[1]
port 77 nsew
flabel metal2 22581 -1908 22623 -652 0 FreeSans 320 0 0 0 vdd_sw_b[2]
port 78 nsew
flabel metal2 20188 -1908 20230 -651 0 FreeSans 320 0 0 0 vdd_sw_b[3]
port 79 nsew
flabel metal2 17797 -1908 17839 -650 0 FreeSans 320 0 0 0 vdd_sw_b[4]
port 80 nsew
flabel metal2 15404 -1908 15446 -651 0 FreeSans 320 0 0 0 vdd_sw_b[5]
port 81 nsew
flabel metal2 13013 -1908 13055 -651 0 FreeSans 320 0 0 0 vdd_sw_b[6]
port 82 nsew
flabel metal2 10621 -1908 10663 -652 0 FreeSans 320 0 0 0 vdd_sw_b[7]
port 83 nsew
flabel space 10504 -1881 10546 -625 0 FreeSans 320 0 0 0 vdd_sw_b[7]
port 84 nsew
flabel metal1 13484 10382 13510 10408 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[9]
port 88 nsew
flabel metal1 13486 10326 13512 10352 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[8]
port 89 nsew
flabel metal1 13482 10270 13508 10296 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[14]
port 90 nsew
flabel metal1 13486 10214 13512 10240 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[13]
port 91 nsew
flabel metal1 13484 10158 13510 10184 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[12]
port 92 nsew
flabel metal1 13482 10438 13506 10464 0 FreeSans 320 0 0 0 sample_delay_cap_ctrl_code[10]
port 93 nsew
flabel metal1 24237 5786 24349 5834 0 FreeSans 320 0 0 0 retimer_eob_delay_offset
port 49 nsew
flabel metal4 24071 4683 24447 6120 0 FreeSans 320 0 0 0 x5.VSS
flabel metal4 24043 6730 24461 7340 0 FreeSans 320 0 0 0 x5.VDD
flabel metal1 23974 5988 24071 6035 0 FreeSans 320 0 0 0 x5.eob
flabel metal1 25545 4635 26484 4663 0 FreeSans 320 0 0 0 x5.delay_code[2]
flabel metal1 25545 4579 28910 4607 0 FreeSans 320 0 0 0 x5.delay_code[1]
flabel metal1 25545 4523 29767 4551 0 FreeSans 320 0 0 0 x5.delay_code[0]
flabel metal1 23937 6371 23991 6405 0 FreeSans 320 0 0 0 x5.delay_code[3]
flabel metal1 25504 3949 25549 3997 0 FreeSans 320 0 0 0 x5.sar_logic[0]
flabel metal1 25496 4155 25541 4203 0 FreeSans 320 0 0 0 x5.sar_logic[1]
flabel metal1 25514 3308 25559 3356 0 FreeSans 320 0 0 0 x5.sar_logic[2]
flabel metal1 25505 2671 25550 2719 0 FreeSans 320 0 0 0 x5.sar_logic[4]
flabel metal1 25504 2874 25549 2922 0 FreeSans 320 0 0 0 x5.sar_logic[5]
flabel metal1 30414 4145 30459 4193 0 FreeSans 320 0 0 0 x5.sar_retimer[1]
flabel metal1 30414 3815 30459 3863 0 FreeSans 320 0 0 0 x5.sar_retimer[0]
flabel metal1 30419 3174 30464 3222 0 FreeSans 320 0 0 0 x5.sar_retimer[3]
flabel metal1 30414 3516 30459 3564 0 FreeSans 320 0 0 0 x5.sar_retimer[2]
flabel metal1 30410 2864 30455 2912 0 FreeSans 320 0 0 0 x5.sar_retimer[5]
flabel metal1 30413 2533 30458 2581 0 FreeSans 320 0 0 0 x5.sar_retimer[4]
flabel metal1 30412 1893 30457 1941 0 FreeSans 320 0 0 0 x5.sar_retimer[7]
flabel metal1 30416 2237 30461 2285 0 FreeSans 320 0 0 0 x5.sar_retimer[6]
flabel metal1 25517 3174 25562 3222 0 FreeSans 320 0 0 0 x5.sar_logic[3]
flabel metal1 25492 2093 25537 2141 0 FreeSans 320 0 0 0 x5.sar_logic[6]
flabel metal1 25489 1894 25534 1942 0 FreeSans 320 0 0 0 x5.sar_logic[7]
flabel metal1 24237 5786 24349 5834 0 FreeSans 320 0 0 0 x5.delay_offset
flabel locali 27440 4016 27515 4062 0 FreeSans 400 0 0 0 x5.x1[0].RESET_B
flabel locali 25607 4264 25641 4298 3 FreeSans 400 0 0 0 x5.x1[0].VGND
flabel locali 25607 4026 25641 4060 0 FreeSans 400 0 0 0 x5.x1[0].CLK
flabel locali 25607 3958 25641 3992 0 FreeSans 400 0 0 0 x5.x1[0].CLK
flabel locali 26343 4094 26377 4128 0 FreeSans 400 0 0 0 x5.x1[0].SET_B
flabel locali 27905 4162 27939 4196 0 FreeSans 400 0 0 0 x5.x1[0].Q
flabel locali 27905 3890 27939 3924 0 FreeSans 400 0 0 0 x5.x1[0].Q
flabel locali 27905 3822 27939 3856 0 FreeSans 400 0 0 0 x5.x1[0].Q
flabel locali 25607 3720 25641 3754 3 FreeSans 400 0 0 0 x5.x1[0].VPWR
flabel locali 25975 4026 26009 4060 0 FreeSans 200 0 0 0 x5.x1[0].D
flabel locali 25975 3958 26009 3992 0 FreeSans 200 0 0 0 x5.x1[0].D
flabel locali 27625 3822 27659 3856 0 FreeSans 400 0 0 0 x5.x1[0].Q_N
flabel locali 27625 3890 27659 3924 0 FreeSans 400 0 0 0 x5.x1[0].Q_N
flabel locali 27625 4162 27659 4196 0 FreeSans 400 0 0 0 x5.x1[0].Q_N
flabel metal1 25607 4264 25641 4298 0 FreeSans 200 0 0 0 x5.x1[0].VGND
flabel metal1 25607 3720 25641 3754 0 FreeSans 200 0 0 0 x5.x1[0].VPWR
flabel nwell 25607 3720 25641 3754 3 FreeSans 400 0 0 0 x5.x1[0].VPB
flabel nwell 25624 3737 25624 3737 0 FreeSans 200 0 0 0 x5.x1[0].VPB
flabel pwell 25607 4264 25641 4298 3 FreeSans 400 0 0 0 x5.x1[0].VNB
flabel pwell 25624 4281 25624 4281 0 FreeSans 200 0 0 0 x5.x1[0].VNB
rlabel comment 25577 4281 25577 4281 2 x5.x1[0].dfbbp_1
rlabel locali 27069 4068 27144 4134 5 x5.x1[0].SET_B
rlabel metal1 27067 4088 27125 4097 5 x5.x1[0].SET_B
rlabel metal1 27067 4125 27125 4134 5 x5.x1[0].SET_B
rlabel metal1 26331 4088 26389 4097 5 x5.x1[0].SET_B
rlabel metal1 26331 4097 27125 4125 5 x5.x1[0].SET_B
rlabel metal1 26331 4125 26389 4134 5 x5.x1[0].SET_B
rlabel metal1 25577 4233 27969 4329 5 x5.x1[0].VGND
rlabel metal1 25577 3689 27969 3785 5 x5.x1[0].VPWR
flabel locali 29832 4016 29907 4062 0 FreeSans 400 0 0 0 x5.x1[1].RESET_B
flabel locali 27999 4264 28033 4298 3 FreeSans 400 0 0 0 x5.x1[1].VGND
flabel locali 27999 4026 28033 4060 0 FreeSans 400 0 0 0 x5.x1[1].CLK
flabel locali 27999 3958 28033 3992 0 FreeSans 400 0 0 0 x5.x1[1].CLK
flabel locali 28735 4094 28769 4128 0 FreeSans 400 0 0 0 x5.x1[1].SET_B
flabel locali 30297 4162 30331 4196 0 FreeSans 400 0 0 0 x5.x1[1].Q
flabel locali 30297 3890 30331 3924 0 FreeSans 400 0 0 0 x5.x1[1].Q
flabel locali 30297 3822 30331 3856 0 FreeSans 400 0 0 0 x5.x1[1].Q
flabel locali 27999 3720 28033 3754 3 FreeSans 400 0 0 0 x5.x1[1].VPWR
flabel locali 28367 4026 28401 4060 0 FreeSans 200 0 0 0 x5.x1[1].D
flabel locali 28367 3958 28401 3992 0 FreeSans 200 0 0 0 x5.x1[1].D
flabel locali 30017 3822 30051 3856 0 FreeSans 400 0 0 0 x5.x1[1].Q_N
flabel locali 30017 3890 30051 3924 0 FreeSans 400 0 0 0 x5.x1[1].Q_N
flabel locali 30017 4162 30051 4196 0 FreeSans 400 0 0 0 x5.x1[1].Q_N
flabel metal1 27999 4264 28033 4298 0 FreeSans 200 0 0 0 x5.x1[1].VGND
flabel metal1 27999 3720 28033 3754 0 FreeSans 200 0 0 0 x5.x1[1].VPWR
flabel nwell 27999 3720 28033 3754 3 FreeSans 400 0 0 0 x5.x1[1].VPB
flabel nwell 28016 3737 28016 3737 0 FreeSans 200 0 0 0 x5.x1[1].VPB
flabel pwell 27999 4264 28033 4298 3 FreeSans 400 0 0 0 x5.x1[1].VNB
flabel pwell 28016 4281 28016 4281 0 FreeSans 200 0 0 0 x5.x1[1].VNB
rlabel comment 27969 4281 27969 4281 2 x5.x1[1].dfbbp_1
rlabel locali 29461 4068 29536 4134 5 x5.x1[1].SET_B
rlabel metal1 29459 4088 29517 4097 5 x5.x1[1].SET_B
rlabel metal1 29459 4125 29517 4134 5 x5.x1[1].SET_B
rlabel metal1 28723 4088 28781 4097 5 x5.x1[1].SET_B
rlabel metal1 28723 4097 29517 4125 5 x5.x1[1].SET_B
rlabel metal1 28723 4125 28781 4134 5 x5.x1[1].SET_B
rlabel metal1 27969 4233 30361 4329 5 x5.x1[1].VGND
rlabel metal1 27969 3689 30361 3785 5 x5.x1[1].VPWR
flabel locali 27440 3316 27515 3362 0 FreeSans 400 0 0 0 x5.x1[2].RESET_B
flabel locali 25607 3080 25641 3114 3 FreeSans 400 0 0 0 x5.x1[2].VGND
flabel locali 25607 3318 25641 3352 0 FreeSans 400 0 0 0 x5.x1[2].CLK
flabel locali 25607 3386 25641 3420 0 FreeSans 400 0 0 0 x5.x1[2].CLK
flabel locali 26343 3250 26377 3284 0 FreeSans 400 0 0 0 x5.x1[2].SET_B
flabel locali 27905 3182 27939 3216 0 FreeSans 400 0 0 0 x5.x1[2].Q
flabel locali 27905 3454 27939 3488 0 FreeSans 400 0 0 0 x5.x1[2].Q
flabel locali 27905 3522 27939 3556 0 FreeSans 400 0 0 0 x5.x1[2].Q
flabel locali 25607 3624 25641 3658 3 FreeSans 400 0 0 0 x5.x1[2].VPWR
flabel locali 25975 3318 26009 3352 0 FreeSans 200 0 0 0 x5.x1[2].D
flabel locali 25975 3386 26009 3420 0 FreeSans 200 0 0 0 x5.x1[2].D
flabel locali 27625 3522 27659 3556 0 FreeSans 400 0 0 0 x5.x1[2].Q_N
flabel locali 27625 3454 27659 3488 0 FreeSans 400 0 0 0 x5.x1[2].Q_N
flabel locali 27625 3182 27659 3216 0 FreeSans 400 0 0 0 x5.x1[2].Q_N
flabel metal1 25607 3080 25641 3114 0 FreeSans 200 0 0 0 x5.x1[2].VGND
flabel metal1 25607 3624 25641 3658 0 FreeSans 200 0 0 0 x5.x1[2].VPWR
flabel nwell 25607 3624 25641 3658 3 FreeSans 400 0 0 0 x5.x1[2].VPB
flabel nwell 25624 3641 25624 3641 0 FreeSans 200 0 0 0 x5.x1[2].VPB
flabel pwell 25607 3080 25641 3114 3 FreeSans 400 0 0 0 x5.x1[2].VNB
flabel pwell 25624 3097 25624 3097 0 FreeSans 200 0 0 0 x5.x1[2].VNB
rlabel comment 25577 3097 25577 3097 4 x5.x1[2].dfbbp_1
rlabel locali 27069 3244 27144 3310 1 x5.x1[2].SET_B
rlabel metal1 27067 3281 27125 3290 1 x5.x1[2].SET_B
rlabel metal1 27067 3244 27125 3253 1 x5.x1[2].SET_B
rlabel metal1 26331 3281 26389 3290 1 x5.x1[2].SET_B
rlabel metal1 26331 3253 27125 3281 1 x5.x1[2].SET_B
rlabel metal1 26331 3244 26389 3253 1 x5.x1[2].SET_B
rlabel metal1 25577 3049 27969 3145 1 x5.x1[2].VGND
rlabel metal1 25577 3593 27969 3689 1 x5.x1[2].VPWR
flabel locali 29832 3316 29907 3362 0 FreeSans 400 0 0 0 x5.x1[3].RESET_B
flabel locali 27999 3080 28033 3114 3 FreeSans 400 0 0 0 x5.x1[3].VGND
flabel locali 27999 3318 28033 3352 0 FreeSans 400 0 0 0 x5.x1[3].CLK
flabel locali 27999 3386 28033 3420 0 FreeSans 400 0 0 0 x5.x1[3].CLK
flabel locali 28735 3250 28769 3284 0 FreeSans 400 0 0 0 x5.x1[3].SET_B
flabel locali 30297 3182 30331 3216 0 FreeSans 400 0 0 0 x5.x1[3].Q
flabel locali 30297 3454 30331 3488 0 FreeSans 400 0 0 0 x5.x1[3].Q
flabel locali 30297 3522 30331 3556 0 FreeSans 400 0 0 0 x5.x1[3].Q
flabel locali 27999 3624 28033 3658 3 FreeSans 400 0 0 0 x5.x1[3].VPWR
flabel locali 28367 3318 28401 3352 0 FreeSans 200 0 0 0 x5.x1[3].D
flabel locali 28367 3386 28401 3420 0 FreeSans 200 0 0 0 x5.x1[3].D
flabel locali 30017 3522 30051 3556 0 FreeSans 400 0 0 0 x5.x1[3].Q_N
flabel locali 30017 3454 30051 3488 0 FreeSans 400 0 0 0 x5.x1[3].Q_N
flabel locali 30017 3182 30051 3216 0 FreeSans 400 0 0 0 x5.x1[3].Q_N
flabel metal1 27999 3080 28033 3114 0 FreeSans 200 0 0 0 x5.x1[3].VGND
flabel metal1 27999 3624 28033 3658 0 FreeSans 200 0 0 0 x5.x1[3].VPWR
flabel nwell 27999 3624 28033 3658 3 FreeSans 400 0 0 0 x5.x1[3].VPB
flabel nwell 28016 3641 28016 3641 0 FreeSans 200 0 0 0 x5.x1[3].VPB
flabel pwell 27999 3080 28033 3114 3 FreeSans 400 0 0 0 x5.x1[3].VNB
flabel pwell 28016 3097 28016 3097 0 FreeSans 200 0 0 0 x5.x1[3].VNB
rlabel comment 27969 3097 27969 3097 4 x5.x1[3].dfbbp_1
rlabel locali 29461 3244 29536 3310 1 x5.x1[3].SET_B
rlabel metal1 29459 3281 29517 3290 1 x5.x1[3].SET_B
rlabel metal1 29459 3244 29517 3253 1 x5.x1[3].SET_B
rlabel metal1 28723 3281 28781 3290 1 x5.x1[3].SET_B
rlabel metal1 28723 3253 29517 3281 1 x5.x1[3].SET_B
rlabel metal1 28723 3244 28781 3253 1 x5.x1[3].SET_B
rlabel metal1 27969 3049 30361 3145 1 x5.x1[3].VGND
rlabel metal1 27969 3593 30361 3689 1 x5.x1[3].VPWR
flabel locali 27440 2736 27515 2782 0 FreeSans 400 0 0 0 x5.x1[4].RESET_B
flabel locali 25607 2984 25641 3018 3 FreeSans 400 0 0 0 x5.x1[4].VGND
flabel locali 25607 2746 25641 2780 0 FreeSans 400 0 0 0 x5.x1[4].CLK
flabel locali 25607 2678 25641 2712 0 FreeSans 400 0 0 0 x5.x1[4].CLK
flabel locali 26343 2814 26377 2848 0 FreeSans 400 0 0 0 x5.x1[4].SET_B
flabel locali 27905 2882 27939 2916 0 FreeSans 400 0 0 0 x5.x1[4].Q
flabel locali 27905 2610 27939 2644 0 FreeSans 400 0 0 0 x5.x1[4].Q
flabel locali 27905 2542 27939 2576 0 FreeSans 400 0 0 0 x5.x1[4].Q
flabel locali 25607 2440 25641 2474 3 FreeSans 400 0 0 0 x5.x1[4].VPWR
flabel locali 25975 2746 26009 2780 0 FreeSans 200 0 0 0 x5.x1[4].D
flabel locali 25975 2678 26009 2712 0 FreeSans 200 0 0 0 x5.x1[4].D
flabel locali 27625 2542 27659 2576 0 FreeSans 400 0 0 0 x5.x1[4].Q_N
flabel locali 27625 2610 27659 2644 0 FreeSans 400 0 0 0 x5.x1[4].Q_N
flabel locali 27625 2882 27659 2916 0 FreeSans 400 0 0 0 x5.x1[4].Q_N
flabel metal1 25607 2984 25641 3018 0 FreeSans 200 0 0 0 x5.x1[4].VGND
flabel metal1 25607 2440 25641 2474 0 FreeSans 200 0 0 0 x5.x1[4].VPWR
flabel nwell 25607 2440 25641 2474 3 FreeSans 400 0 0 0 x5.x1[4].VPB
flabel nwell 25624 2457 25624 2457 0 FreeSans 200 0 0 0 x5.x1[4].VPB
flabel pwell 25607 2984 25641 3018 3 FreeSans 400 0 0 0 x5.x1[4].VNB
flabel pwell 25624 3001 25624 3001 0 FreeSans 200 0 0 0 x5.x1[4].VNB
rlabel comment 25577 3001 25577 3001 2 x5.x1[4].dfbbp_1
rlabel locali 27069 2788 27144 2854 5 x5.x1[4].SET_B
rlabel metal1 27067 2808 27125 2817 5 x5.x1[4].SET_B
rlabel metal1 27067 2845 27125 2854 5 x5.x1[4].SET_B
rlabel metal1 26331 2808 26389 2817 5 x5.x1[4].SET_B
rlabel metal1 26331 2817 27125 2845 5 x5.x1[4].SET_B
rlabel metal1 26331 2845 26389 2854 5 x5.x1[4].SET_B
rlabel metal1 25577 2953 27969 3049 5 x5.x1[4].VGND
rlabel metal1 25577 2409 27969 2505 5 x5.x1[4].VPWR
flabel locali 29832 2736 29907 2782 0 FreeSans 400 0 0 0 x5.x1[5].RESET_B
flabel locali 27999 2984 28033 3018 3 FreeSans 400 0 0 0 x5.x1[5].VGND
flabel locali 27999 2746 28033 2780 0 FreeSans 400 0 0 0 x5.x1[5].CLK
flabel locali 27999 2678 28033 2712 0 FreeSans 400 0 0 0 x5.x1[5].CLK
flabel locali 28735 2814 28769 2848 0 FreeSans 400 0 0 0 x5.x1[5].SET_B
flabel locali 30297 2882 30331 2916 0 FreeSans 400 0 0 0 x5.x1[5].Q
flabel locali 30297 2610 30331 2644 0 FreeSans 400 0 0 0 x5.x1[5].Q
flabel locali 30297 2542 30331 2576 0 FreeSans 400 0 0 0 x5.x1[5].Q
flabel locali 27999 2440 28033 2474 3 FreeSans 400 0 0 0 x5.x1[5].VPWR
flabel locali 28367 2746 28401 2780 0 FreeSans 200 0 0 0 x5.x1[5].D
flabel locali 28367 2678 28401 2712 0 FreeSans 200 0 0 0 x5.x1[5].D
flabel locali 30017 2542 30051 2576 0 FreeSans 400 0 0 0 x5.x1[5].Q_N
flabel locali 30017 2610 30051 2644 0 FreeSans 400 0 0 0 x5.x1[5].Q_N
flabel locali 30017 2882 30051 2916 0 FreeSans 400 0 0 0 x5.x1[5].Q_N
flabel metal1 27999 2984 28033 3018 0 FreeSans 200 0 0 0 x5.x1[5].VGND
flabel metal1 27999 2440 28033 2474 0 FreeSans 200 0 0 0 x5.x1[5].VPWR
flabel nwell 27999 2440 28033 2474 3 FreeSans 400 0 0 0 x5.x1[5].VPB
flabel nwell 28016 2457 28016 2457 0 FreeSans 200 0 0 0 x5.x1[5].VPB
flabel pwell 27999 2984 28033 3018 3 FreeSans 400 0 0 0 x5.x1[5].VNB
flabel pwell 28016 3001 28016 3001 0 FreeSans 200 0 0 0 x5.x1[5].VNB
rlabel comment 27969 3001 27969 3001 2 x5.x1[5].dfbbp_1
rlabel locali 29461 2788 29536 2854 5 x5.x1[5].SET_B
rlabel metal1 29459 2808 29517 2817 5 x5.x1[5].SET_B
rlabel metal1 29459 2845 29517 2854 5 x5.x1[5].SET_B
rlabel metal1 28723 2808 28781 2817 5 x5.x1[5].SET_B
rlabel metal1 28723 2817 29517 2845 5 x5.x1[5].SET_B
rlabel metal1 28723 2845 28781 2854 5 x5.x1[5].SET_B
rlabel metal1 27969 2953 30361 3049 5 x5.x1[5].VGND
rlabel metal1 27969 2409 30361 2505 5 x5.x1[5].VPWR
flabel locali 27440 2036 27515 2082 0 FreeSans 400 0 0 0 x5.x1[6].RESET_B
flabel locali 25607 1800 25641 1834 3 FreeSans 400 0 0 0 x5.x1[6].VGND
flabel locali 25607 2038 25641 2072 0 FreeSans 400 0 0 0 x5.x1[6].CLK
flabel locali 25607 2106 25641 2140 0 FreeSans 400 0 0 0 x5.x1[6].CLK
flabel locali 26343 1970 26377 2004 0 FreeSans 400 0 0 0 x5.x1[6].SET_B
flabel locali 27905 1902 27939 1936 0 FreeSans 400 0 0 0 x5.x1[6].Q
flabel locali 27905 2174 27939 2208 0 FreeSans 400 0 0 0 x5.x1[6].Q
flabel locali 27905 2242 27939 2276 0 FreeSans 400 0 0 0 x5.x1[6].Q
flabel locali 25607 2344 25641 2378 3 FreeSans 400 0 0 0 x5.x1[6].VPWR
flabel locali 25975 2038 26009 2072 0 FreeSans 200 0 0 0 x5.x1[6].D
flabel locali 25975 2106 26009 2140 0 FreeSans 200 0 0 0 x5.x1[6].D
flabel locali 27625 2242 27659 2276 0 FreeSans 400 0 0 0 x5.x1[6].Q_N
flabel locali 27625 2174 27659 2208 0 FreeSans 400 0 0 0 x5.x1[6].Q_N
flabel locali 27625 1902 27659 1936 0 FreeSans 400 0 0 0 x5.x1[6].Q_N
flabel metal1 25607 1800 25641 1834 0 FreeSans 200 0 0 0 x5.x1[6].VGND
flabel metal1 25607 2344 25641 2378 0 FreeSans 200 0 0 0 x5.x1[6].VPWR
flabel nwell 25607 2344 25641 2378 3 FreeSans 400 0 0 0 x5.x1[6].VPB
flabel nwell 25624 2361 25624 2361 0 FreeSans 200 0 0 0 x5.x1[6].VPB
flabel pwell 25607 1800 25641 1834 3 FreeSans 400 0 0 0 x5.x1[6].VNB
flabel pwell 25624 1817 25624 1817 0 FreeSans 200 0 0 0 x5.x1[6].VNB
rlabel comment 25577 1817 25577 1817 4 x5.x1[6].dfbbp_1
rlabel locali 27069 1964 27144 2030 1 x5.x1[6].SET_B
rlabel metal1 27067 2001 27125 2010 1 x5.x1[6].SET_B
rlabel metal1 27067 1964 27125 1973 1 x5.x1[6].SET_B
rlabel metal1 26331 2001 26389 2010 1 x5.x1[6].SET_B
rlabel metal1 26331 1973 27125 2001 1 x5.x1[6].SET_B
rlabel metal1 26331 1964 26389 1973 1 x5.x1[6].SET_B
rlabel metal1 25577 1769 27969 1865 1 x5.x1[6].VGND
rlabel metal1 25577 2313 27969 2409 1 x5.x1[6].VPWR
flabel locali 29832 2036 29907 2082 0 FreeSans 400 0 0 0 x5.x1[7].RESET_B
flabel locali 27999 1800 28033 1834 3 FreeSans 400 0 0 0 x5.x1[7].VGND
flabel locali 27999 2038 28033 2072 0 FreeSans 400 0 0 0 x5.x1[7].CLK
flabel locali 27999 2106 28033 2140 0 FreeSans 400 0 0 0 x5.x1[7].CLK
flabel locali 28735 1970 28769 2004 0 FreeSans 400 0 0 0 x5.x1[7].SET_B
flabel locali 30297 1902 30331 1936 0 FreeSans 400 0 0 0 x5.x1[7].Q
flabel locali 30297 2174 30331 2208 0 FreeSans 400 0 0 0 x5.x1[7].Q
flabel locali 30297 2242 30331 2276 0 FreeSans 400 0 0 0 x5.x1[7].Q
flabel locali 27999 2344 28033 2378 3 FreeSans 400 0 0 0 x5.x1[7].VPWR
flabel locali 28367 2038 28401 2072 0 FreeSans 200 0 0 0 x5.x1[7].D
flabel locali 28367 2106 28401 2140 0 FreeSans 200 0 0 0 x5.x1[7].D
flabel locali 30017 2242 30051 2276 0 FreeSans 400 0 0 0 x5.x1[7].Q_N
flabel locali 30017 2174 30051 2208 0 FreeSans 400 0 0 0 x5.x1[7].Q_N
flabel locali 30017 1902 30051 1936 0 FreeSans 400 0 0 0 x5.x1[7].Q_N
flabel metal1 27999 1800 28033 1834 0 FreeSans 200 0 0 0 x5.x1[7].VGND
flabel metal1 27999 2344 28033 2378 0 FreeSans 200 0 0 0 x5.x1[7].VPWR
flabel nwell 27999 2344 28033 2378 3 FreeSans 400 0 0 0 x5.x1[7].VPB
flabel nwell 28016 2361 28016 2361 0 FreeSans 200 0 0 0 x5.x1[7].VPB
flabel pwell 27999 1800 28033 1834 3 FreeSans 400 0 0 0 x5.x1[7].VNB
flabel pwell 28016 1817 28016 1817 0 FreeSans 200 0 0 0 x5.x1[7].VNB
rlabel comment 27969 1817 27969 1817 4 x5.x1[7].dfbbp_1
rlabel locali 29461 1964 29536 2030 1 x5.x1[7].SET_B
rlabel metal1 29459 2001 29517 2010 1 x5.x1[7].SET_B
rlabel metal1 29459 1964 29517 1973 1 x5.x1[7].SET_B
rlabel metal1 28723 2001 28781 2010 1 x5.x1[7].SET_B
rlabel metal1 28723 1973 29517 2001 1 x5.x1[7].SET_B
rlabel metal1 28723 1964 28781 1973 1 x5.x1[7].SET_B
rlabel metal1 27969 1769 30361 1865 1 x5.x1[7].VGND
rlabel metal1 27969 2313 30361 2409 1 x5.x1[7].VPWR
flabel metal1 23974 5988 24642 6035 0 FreeSans 320 0 0 0 x5.x2.IN
flabel metal1 30450 5986 30632 6032 0 FreeSans 320 0 0 0 x5.x2.OUT
flabel metal1 23937 6371 24075 6405 0 FreeSans 320 0 0 0 x5.x2.code[3]
flabel metal1 28852 4660 28910 5837 0 FreeSans 320 0 0 0 x5.x2.code[1]
flabel metal1 26426 4660 26484 5837 0 FreeSans 320 0 0 0 x5.x2.code[2]
flabel metal4 24043 6730 24461 7340 0 FreeSans 320 0 0 0 x5.x2.VDD
flabel metal4 24071 4683 24447 6120 0 FreeSans 320 0 0 0 x5.x2.VSS
flabel metal2 24401 5786 24837 5832 0 FreeSans 320 0 0 0 x5.x2.code_offset
flabel metal1 29708 4659 29767 5840 0 FreeSans 320 0 0 0 x5.x2.code[0]
flabel metal1 24585 6441 24619 6475 0 FreeSans 320 0 0 0 x5.x2.x8.input_stack
flabel nwell 24629 7224 24663 7284 0 FreeSans 320 0 0 0 x5.x2.x8.vdd
flabel metal1 24623 6522 24669 6534 0 FreeSans 320 0 0 0 x5.x2.x8.output_stack
flabel poly 24562 5784 24664 5814 0 FreeSans 320 0 0 0 x5.x2.x9.input_stack
flabel metal1 24676 4731 24710 4791 0 FreeSans 320 0 0 0 x5.x2.x9.vss
flabel metal1 24670 5757 24716 5769 0 FreeSans 320 0 0 0 x5.x2.x9.output_stack
flabel locali 24163 6441 24197 6475 0 FreeSans 340 0 0 0 x5.x2.x10.Y
flabel locali 24163 6373 24197 6407 0 FreeSans 340 0 0 0 x5.x2.x10.Y
flabel locali 24071 6373 24105 6407 0 FreeSans 340 0 0 0 x5.x2.x10.A
flabel metal1 24028 6135 24062 6169 0 FreeSans 200 0 0 0 x5.x2.x10.VGND
flabel metal1 24028 6679 24062 6713 0 FreeSans 200 0 0 0 x5.x2.x10.VPWR
rlabel comment 23999 6152 23999 6152 4 x5.x2.x10.inv_1
rlabel metal1 23999 6104 24275 6200 1 x5.x2.x10.VGND
rlabel metal1 23999 6648 24275 6744 1 x5.x2.x10.VPWR
flabel pwell 24028 6135 24062 6169 0 FreeSans 200 0 0 0 x5.x2.x10.VNB
flabel nwell 24028 6679 24062 6713 0 FreeSans 200 0 0 0 x5.x2.x10.VPB
flabel locali 24261 6441 24295 6475 0 FreeSans 340 0 0 0 x5.x2.x11.Y
flabel locali 24261 6373 24295 6407 0 FreeSans 340 0 0 0 x5.x2.x11.Y
flabel locali 24353 6373 24387 6407 0 FreeSans 340 0 0 0 x5.x2.x11.A
flabel metal1 24396 6135 24430 6169 0 FreeSans 200 0 0 0 x5.x2.x11.VGND
flabel metal1 24396 6679 24430 6713 0 FreeSans 200 0 0 0 x5.x2.x11.VPWR
rlabel comment 24459 6152 24459 6152 6 x5.x2.x11.inv_1
rlabel metal1 24183 6104 24459 6200 1 x5.x2.x11.VGND
rlabel metal1 24183 6648 24459 6744 1 x5.x2.x11.VPWR
flabel pwell 24396 6135 24430 6169 0 FreeSans 200 0 0 0 x5.x2.x11.VNB
flabel nwell 24396 6679 24430 6713 0 FreeSans 200 0 0 0 x5.x2.x11.VPB
flabel metal1 25227 6198 25261 6232 0 FreeSans 320 0 0 0 x5.x2.x6.SW
flabel nwell 24671 7260 25341 7328 0 FreeSans 320 0 0 0 x5.x2.x6.VDD
flabel pdiff 25259 6067 25317 6151 0 FreeSans 320 0 0 0 x5.x2.x6.delay_signal
flabel metal4 24671 7259 24772 7328 0 FreeSans 320 0 0 0 x5.x2.x6.VDD
flabel via3 24772 6101 24836 6165 0 FreeSans 320 0 0 0 x5.x2.x6.floating
flabel viali 25580 5797 25614 5831 0 FreeSans 320 0 0 0 x5.x2.x7.SW
flabel ndiff 25612 5869 25670 5953 0 FreeSans 320 0 0 0 x5.x2.x7.delay_signal
flabel metal4 25019 4692 25691 4760 0 FreeSans 320 0 0 0 x5.x2.x7.VSS
flabel via3 25123 5856 25187 5920 0 FreeSans 320 0 0 0 x5.x2.x7.floating
flabel viali 26312 5797 26346 5831 0 FreeSans 320 0 0 0 x5.x2.x4[3].SW
flabel ndiff 26344 5869 26402 5953 0 FreeSans 320 0 0 0 x5.x2.x4[3].delay_signal
flabel metal4 25751 4692 26423 4760 0 FreeSans 320 0 0 0 x5.x2.x4[3].VSS
flabel via3 25855 5856 25919 5920 0 FreeSans 320 0 0 0 x5.x2.x4[3].floating
flabel metal1 26085 6201 26119 6235 0 FreeSans 320 0 0 0 x5.x2.x5[6].SW
flabel nwell 26005 7263 26675 7331 0 FreeSans 320 0 0 0 x5.x2.x5[6].VDD
flabel pdiff 26029 6070 26087 6154 0 FreeSans 320 0 0 0 x5.x2.x5[6].delay_signal
flabel metal4 26574 7262 26675 7331 0 FreeSans 320 0 0 0 x5.x2.x5[6].VDD
flabel via3 26510 6104 26574 6168 0 FreeSans 320 0 0 0 x5.x2.x5[6].floating
flabel metal1 25959 6201 25993 6235 0 FreeSans 320 0 0 0 x5.x2.x5[7].SW
flabel nwell 25403 7263 26073 7331 0 FreeSans 320 0 0 0 x5.x2.x5[7].VDD
flabel pdiff 25991 6070 26049 6154 0 FreeSans 320 0 0 0 x5.x2.x5[7].delay_signal
flabel metal4 25403 7262 25504 7331 0 FreeSans 320 0 0 0 x5.x2.x5[7].VDD
flabel via3 25504 6104 25568 6168 0 FreeSans 320 0 0 0 x5.x2.x5[7].floating
flabel viali 26434 5797 26468 5831 0 FreeSans 320 0 0 0 x5.x2.x4[2].SW
flabel ndiff 26378 5869 26436 5953 0 FreeSans 320 0 0 0 x5.x2.x4[2].delay_signal
flabel metal4 26357 4692 27029 4760 0 FreeSans 320 0 0 0 x5.x2.x4[2].VSS
flabel via3 26861 5856 26925 5920 0 FreeSans 320 0 0 0 x5.x2.x4[2].floating
flabel metal1 27171 6201 27205 6235 0 FreeSans 320 0 0 0 x5.x2.x5[5].SW
flabel nwell 26615 7263 27285 7331 0 FreeSans 320 0 0 0 x5.x2.x5[5].VDD
flabel pdiff 27203 6070 27261 6154 0 FreeSans 320 0 0 0 x5.x2.x5[5].delay_signal
flabel metal4 26615 7262 26716 7331 0 FreeSans 320 0 0 0 x5.x2.x5[5].VDD
flabel via3 26716 6104 26780 6168 0 FreeSans 320 0 0 0 x5.x2.x5[5].floating
flabel viali 27524 5797 27558 5831 0 FreeSans 320 0 0 0 x5.x2.x4[1].SW
flabel ndiff 27556 5869 27614 5953 0 FreeSans 320 0 0 0 x5.x2.x4[1].delay_signal
flabel metal4 26963 4692 27635 4760 0 FreeSans 320 0 0 0 x5.x2.x4[1].VSS
flabel via3 27067 5856 27131 5920 0 FreeSans 320 0 0 0 x5.x2.x4[1].floating
flabel metal1 27297 6201 27331 6235 0 FreeSans 320 0 0 0 x5.x2.x5[4].SW
flabel nwell 27217 7263 27887 7331 0 FreeSans 320 0 0 0 x5.x2.x5[4].VDD
flabel pdiff 27241 6070 27299 6154 0 FreeSans 320 0 0 0 x5.x2.x5[4].delay_signal
flabel metal4 27786 7262 27887 7331 0 FreeSans 320 0 0 0 x5.x2.x5[4].VDD
flabel via3 27722 6104 27786 6168 0 FreeSans 320 0 0 0 x5.x2.x5[4].floating
flabel viali 27646 5797 27680 5831 0 FreeSans 320 0 0 0 x5.x2.x4[0].SW
flabel ndiff 27590 5869 27648 5953 0 FreeSans 320 0 0 0 x5.x2.x4[0].delay_signal
flabel metal4 27569 4692 28241 4760 0 FreeSans 320 0 0 0 x5.x2.x4[0].VSS
flabel via3 28073 5856 28137 5920 0 FreeSans 320 0 0 0 x5.x2.x4[0].floating
flabel metal1 28383 6201 28417 6235 0 FreeSans 320 0 0 0 x5.x2.x5[3].SW
flabel nwell 27827 7263 28497 7331 0 FreeSans 320 0 0 0 x5.x2.x5[3].VDD
flabel pdiff 28415 6070 28473 6154 0 FreeSans 320 0 0 0 x5.x2.x5[3].delay_signal
flabel metal4 27827 7262 27928 7331 0 FreeSans 320 0 0 0 x5.x2.x5[3].VDD
flabel via3 27928 6104 27992 6168 0 FreeSans 320 0 0 0 x5.x2.x5[3].floating
flabel viali 28862 5797 28896 5831 0 FreeSans 320 0 0 0 x5.x2.x3[1].SW
flabel ndiff 28894 5869 28952 5953 0 FreeSans 320 0 0 0 x5.x2.x3[1].delay_signal
flabel metal4 28301 4692 28973 4760 0 FreeSans 320 0 0 0 x5.x2.x3[1].VSS
flabel via3 28405 5856 28469 5920 0 FreeSans 320 0 0 0 x5.x2.x3[1].floating
flabel metal1 28509 6201 28543 6235 0 FreeSans 320 0 0 0 x5.x2.x5[2].SW
flabel nwell 28429 7263 29099 7331 0 FreeSans 320 0 0 0 x5.x2.x5[2].VDD
flabel pdiff 28453 6070 28511 6154 0 FreeSans 320 0 0 0 x5.x2.x5[2].delay_signal
flabel metal4 28998 7262 29099 7331 0 FreeSans 320 0 0 0 x5.x2.x5[2].VDD
flabel via3 28934 6104 28998 6168 0 FreeSans 320 0 0 0 x5.x2.x5[2].floating
flabel viali 28984 5797 29018 5831 0 FreeSans 320 0 0 0 x5.x2.x3[0].SW
flabel ndiff 28928 5869 28986 5953 0 FreeSans 320 0 0 0 x5.x2.x3[0].delay_signal
flabel metal4 28907 4692 29579 4760 0 FreeSans 320 0 0 0 x5.x2.x3[0].VSS
flabel via3 29411 5856 29475 5920 0 FreeSans 320 0 0 0 x5.x2.x3[0].floating
flabel metal1 29595 6201 29629 6235 0 FreeSans 320 0 0 0 x5.x2.x5[1].SW
flabel nwell 29039 7263 29709 7331 0 FreeSans 320 0 0 0 x5.x2.x5[1].VDD
flabel pdiff 29627 6070 29685 6154 0 FreeSans 320 0 0 0 x5.x2.x5[1].delay_signal
flabel metal4 29039 7262 29140 7331 0 FreeSans 320 0 0 0 x5.x2.x5[1].VDD
flabel via3 29140 6104 29204 6168 0 FreeSans 320 0 0 0 x5.x2.x5[1].floating
flabel viali 29718 5797 29752 5831 0 FreeSans 320 0 0 0 x5.x2.x2.SW
flabel ndiff 29662 5869 29720 5953 0 FreeSans 320 0 0 0 x5.x2.x2.delay_signal
flabel metal4 29641 4692 30313 4760 0 FreeSans 320 0 0 0 x5.x2.x2.VSS
flabel via3 30145 5856 30209 5920 0 FreeSans 320 0 0 0 x5.x2.x2.floating
flabel metal1 29721 6201 29755 6235 0 FreeSans 320 0 0 0 x5.x2.x5[0].SW
flabel nwell 29641 7263 30311 7331 0 FreeSans 320 0 0 0 x5.x2.x5[0].VDD
flabel pdiff 29665 6070 29723 6154 0 FreeSans 320 0 0 0 x5.x2.x5[0].delay_signal
flabel metal4 30210 7262 30311 7331 0 FreeSans 320 0 0 0 x5.x2.x5[0].VDD
flabel via3 30146 6104 30210 6168 0 FreeSans 320 0 0 0 x5.x2.x5[0].floating
flabel metal1 30708 6302 30742 6336 0 FreeSans 200 0 0 0 x5.x3.VPWR
flabel metal1 30708 5758 30742 5792 0 FreeSans 200 0 0 0 x5.x3.VGND
flabel locali 30708 6302 30742 6336 0 FreeSans 200 0 0 0 x5.x3.VPWR
flabel locali 30708 5758 30742 5792 0 FreeSans 200 0 0 0 x5.x3.VGND
flabel locali 30891 5860 30925 5894 0 FreeSans 200 0 0 0 x5.x3.X
flabel locali 30891 6132 30925 6166 0 FreeSans 200 0 0 0 x5.x3.X
flabel locali 30891 6200 30925 6234 0 FreeSans 200 0 0 0 x5.x3.X
flabel locali 30708 5996 30742 6030 0 FreeSans 200 0 0 0 x5.x3.A
flabel nwell 30708 6302 30742 6336 0 FreeSans 200 0 0 0 x5.x3.VPB
flabel pwell 30708 5758 30742 5792 0 FreeSans 200 0 0 0 x5.x3.VNB
rlabel comment 30679 5775 30679 5775 4 x5.x3.buf_2
rlabel metal1 30679 5727 31047 5823 1 x5.x3.VGND
rlabel metal1 30679 6271 31047 6367 1 x5.x3.VPWR
flabel metal2 18284 -1221 18326 1735 0 FreeSans 320 0 0 0 x4.VSS_SW[3]
flabel metal2 15892 -1220 15934 1735 0 FreeSans 320 0 0 0 x4.VSS_SW[4]
flabel metal2 13501 -1220 13543 1735 0 FreeSans 320 0 0 0 x4.VSS_SW[5]
flabel metal2 22865 -503 22907 1735 0 FreeSans 320 0 0 0 x4.VDD_SW[2]
flabel metal2 20473 -503 20515 1735 0 FreeSans 320 0 0 0 x4.VDD_SW[3]
flabel metal2 18081 -503 18123 1735 0 FreeSans 320 0 0 0 x4.VDD_SW[4]
flabel metal2 15689 -503 15731 1735 0 FreeSans 320 0 0 0 x4.VDD_SW[5]
flabel metal2 13297 -503 13339 1735 0 FreeSans 320 0 0 0 x4.VDD_SW[6]
flabel metal2 22499 -111 22541 1735 0 FreeSans 320 0 0 0 x4.D[2]
flabel metal2 20106 -111 20148 1735 0 FreeSans 320 0 0 0 x4.D[3]
flabel metal2 17715 -112 17757 1735 0 FreeSans 320 0 0 0 x4.D[4]
flabel metal2 15322 -111 15364 1735 0 FreeSans 320 0 0 0 x4.D[5]
flabel metal2 12931 -112 12973 1735 0 FreeSans 320 0 0 0 x4.D[6]
flabel metal2 22094 37 22136 1735 0 FreeSans 320 0 0 0 x4.check[1]
flabel metal2 19705 37 19747 1735 0 FreeSans 320 0 0 0 x4.check[2]
flabel metal2 17313 38 17355 1735 0 FreeSans 320 0 0 0 x4.check[3]
flabel metal2 14919 37 14961 1735 0 FreeSans 320 0 0 0 x4.check[4]
flabel metal2 12529 37 12571 1735 0 FreeSans 320 0 0 0 x4.check[5]
flabel metal2 25257 -503 25299 1735 0 FreeSans 320 0 0 0 x4.VDD_SW[1]
flabel metal2 10137 38 10179 1735 0 FreeSans 320 0 0 0 x4.check[6]
flabel metal2 10539 -112 10581 1735 0 FreeSans 320 0 0 0 x4.D[7]
flabel metal2 10905 -503 10947 1735 0 FreeSans 320 0 0 0 x4.VDD_SW[7]
flabel metal2 11108 -1220 11150 1735 0 FreeSans 320 0 0 0 x4.VSS_SW[6]
flabel metal2 8716 -1220 8758 1735 0 FreeSans 320 0 0 0 x4.VSS_SW[7]
rlabel comment 12961 845 12961 845 4 x4.buf_1
rlabel comment 13789 845 13789 845 4 x4.buf_16
rlabel comment 13237 845 13237 845 4 x4.buf_4
rlabel comment 8851 -297 8851 -297 4 x4.buf_4
rlabel comment 9403 -297 9403 -297 4 x4.buf_16
rlabel comment 8575 -297 8575 -297 4 x4.buf_1
rlabel comment 11703 -297 11703 -297 4 x4.buf_4
rlabel comment 12255 -297 12255 -297 4 x4.buf_16
rlabel comment 11427 -297 11427 -297 4 x4.buf_1
rlabel comment 14791 -297 14791 -297 4 x4.buf_1
rlabel comment 15619 -297 15619 -297 4 x4.buf_16
rlabel comment 15067 -297 15067 -297 4 x4.buf_4
rlabel comment 17643 -297 17643 -297 4 x4.buf_1
rlabel comment 18471 -297 18471 -297 4 x4.buf_16
rlabel comment 17919 -297 17919 -297 4 x4.buf_4
rlabel comment 20557 -297 20557 -297 4 x4.buf_1
rlabel comment 21385 -297 21385 -297 4 x4.buf_16
rlabel comment 20833 -297 20833 -297 4 x4.buf_4
rlabel comment 22305 -297 22305 -297 4 x4.buf_1
rlabel comment 23133 -297 23133 -297 4 x4.buf_16
rlabel comment 22581 -297 22581 -297 4 x4.buf_4
flabel metal2 24974 -1887 25016 -650 0 FreeSans 320 0 0 0 x4.VDD_SW_b[1]
flabel metal2 22581 -1887 22623 -652 0 FreeSans 320 0 0 0 x4.VDD_SW_b[2]
flabel metal2 20188 -1887 20230 -651 0 FreeSans 320 0 0 0 x4.VDD_SW_b[3]
flabel metal2 17797 -1887 17839 -650 0 FreeSans 320 0 0 0 x4.VDD_SW_b[4]
flabel metal2 13013 -1887 13055 -651 0 FreeSans 320 0 0 0 x4.VDD_SW_b[6]
flabel metal2 10621 -1887 10663 -652 0 FreeSans 320 0 0 0 x4.VDD_SW_b[7]
rlabel comment 8851 -985 8851 -985 4 x4.buf_4
rlabel comment 9403 -985 9403 -985 4 x4.buf_16
rlabel comment 8575 -985 8575 -985 4 x4.buf_1
rlabel comment 11427 -985 11427 -985 4 x4.buf_1
rlabel comment 12255 -985 12255 -985 4 x4.buf_16
rlabel comment 11703 -985 11703 -985 4 x4.buf_4
rlabel comment 14555 -985 14555 -985 4 x4.buf_4
rlabel comment 15107 -985 15107 -985 4 x4.buf_16
rlabel comment 14279 -985 14279 -985 4 x4.buf_1
rlabel comment 17131 -985 17131 -985 4 x4.buf_1
rlabel comment 17959 -985 17959 -985 4 x4.buf_16
rlabel comment 17407 -985 17407 -985 4 x4.buf_4
rlabel comment 19983 -985 19983 -985 4 x4.buf_1
rlabel comment 20811 -985 20811 -985 4 x4.buf_16
rlabel comment 20259 -985 20259 -985 4 x4.buf_4
rlabel comment 22835 -985 22835 -985 4 x4.buf_1
rlabel comment 23663 -985 23663 -985 4 x4.buf_16
rlabel comment 23111 -985 23111 -985 4 x4.buf_4
flabel metal2 23228 -1908 23270 -1331 0 FreeSans 320 0 0 0 x4.VSS_SW_b[1]
flabel metal2 20835 -1908 20877 -1330 0 FreeSans 320 0 0 0 x4.VSS_SW_b[2]
flabel metal2 18444 -1908 18486 -1331 0 FreeSans 320 0 0 0 x4.VSS_SW_b[3]
flabel metal2 16052 -1908 16094 -1331 0 FreeSans 320 0 0 0 x4.VSS_SW_b[4]
flabel metal2 13659 -1908 13701 -1331 0 FreeSans 320 0 0 0 x4.VSS_SW_b[5]
flabel metal2 11268 -1908 11310 -1331 0 FreeSans 320 0 0 0 x4.VSS_SW_b[6]
flabel metal2 8876 -1908 8918 -1331 0 FreeSans 320 0 0 0 x4.VSS_SW_b[7]
flabel metal2 23068 -1219 23110 1735 0 FreeSans 320 0 0 0 x4.VSS_SW[1]
flabel metal2 20677 -1219 20719 1735 0 FreeSans 320 0 0 0 x4.VSS_SW[2]
flabel metal1 8449 961 12877 995 0 FreeSans 320 0 0 0 x4.ready
flabel metal1 8449 1157 8541 1191 0 FreeSans 320 0 0 0 x4.reset
flabel metal2 15404 -1887 15446 -651 0 FreeSans 320 0 0 0 x4.VDD_SW_b[5]
flabel metal4 20981 -1640 25451 -1451 0 FreeSans 1600 0 0 0 x4.VSS
flabel metal2 24489 38 24531 1735 0 FreeSans 320 0 0 0 x4.check[0]
flabel metal2 24892 -111 24934 1735 0 FreeSans 320 0 0 0 x4.D[1]
flabel metal4 15853 1156 24265 1453 0 FreeSans 1600 0 0 0 x4.VDD
flabel locali 23416 -1453 23450 -1419 0 FreeSans 400 0 0 0 x4.x35.RESET_B
flabel locali 25256 -1691 25290 -1657 7 FreeSans 400 0 0 0 x4.x35.VGND
flabel locali 25256 -1453 25290 -1419 0 FreeSans 400 0 0 0 x4.x35.CLK_N
flabel locali 25256 -1385 25290 -1351 0 FreeSans 400 0 0 0 x4.x35.CLK_N
flabel locali 24520 -1521 24554 -1487 0 FreeSans 400 0 0 0 x4.x35.SET_B
flabel locali 22956 -1589 22990 -1555 0 FreeSans 400 0 0 0 x4.x35.Q
flabel locali 22956 -1317 22990 -1283 0 FreeSans 400 0 0 0 x4.x35.Q
flabel locali 22956 -1249 22990 -1215 0 FreeSans 400 0 0 0 x4.x35.Q
flabel locali 25256 -1147 25290 -1113 7 FreeSans 400 0 0 0 x4.x35.VPWR
flabel locali 24888 -1453 24922 -1419 0 FreeSans 200 0 0 0 x4.x35.D
flabel locali 24888 -1385 24922 -1351 0 FreeSans 200 0 0 0 x4.x35.D
flabel locali 23232 -1249 23266 -1215 0 FreeSans 400 0 0 0 x4.x35.Q_N
flabel locali 23232 -1317 23266 -1283 0 FreeSans 400 0 0 0 x4.x35.Q_N
flabel locali 23232 -1589 23266 -1555 0 FreeSans 400 0 0 0 x4.x35.Q_N
flabel metal1 25256 -1691 25290 -1657 0 FreeSans 200 0 0 0 x4.x35.VGND
flabel metal1 25256 -1147 25290 -1113 0 FreeSans 200 0 0 0 x4.x35.VPWR
flabel nwell 25256 -1147 25290 -1113 7 FreeSans 400 0 0 0 x4.x35.VPB
flabel nwell 25273 -1130 25273 -1130 0 FreeSans 200 0 0 0 x4.x35.VPB
flabel pwell 25256 -1691 25290 -1657 7 FreeSans 400 0 0 0 x4.x35.VNB
flabel pwell 25273 -1674 25273 -1674 0 FreeSans 200 0 0 0 x4.x35.VNB
rlabel comment 25319 -1674 25319 -1674 6 x4.x35.dfbbn_1
rlabel locali 23754 -1527 23863 -1461 1 x4.x35.SET_B
rlabel metal1 23758 -1490 23816 -1481 1 x4.x35.SET_B
rlabel metal1 23758 -1527 23816 -1518 1 x4.x35.SET_B
rlabel metal1 24508 -1490 24566 -1481 1 x4.x35.SET_B
rlabel metal1 23758 -1518 24566 -1490 1 x4.x35.SET_B
rlabel metal1 24508 -1527 24566 -1518 1 x4.x35.SET_B
rlabel metal1 22927 -1722 25319 -1626 1 x4.x35.VGND
rlabel metal1 22927 -1178 25319 -1082 1 x4.x35.VPWR
flabel locali 24796 -764 24830 -730 0 FreeSans 400 0 0 0 x4.x34.RESET_B
flabel locali 22956 -1002 22990 -968 3 FreeSans 400 0 0 0 x4.x34.VGND
flabel locali 22956 -764 22990 -730 0 FreeSans 400 0 0 0 x4.x34.CLK_N
flabel locali 22956 -696 22990 -662 0 FreeSans 400 0 0 0 x4.x34.CLK_N
flabel locali 23692 -832 23726 -798 0 FreeSans 400 0 0 0 x4.x34.SET_B
flabel locali 25256 -900 25290 -866 0 FreeSans 400 0 0 0 x4.x34.Q
flabel locali 25256 -628 25290 -594 0 FreeSans 400 0 0 0 x4.x34.Q
flabel locali 25256 -560 25290 -526 0 FreeSans 400 0 0 0 x4.x34.Q
flabel locali 22956 -458 22990 -424 3 FreeSans 400 0 0 0 x4.x34.VPWR
flabel locali 23324 -764 23358 -730 0 FreeSans 200 0 0 0 x4.x34.D
flabel locali 23324 -696 23358 -662 0 FreeSans 200 0 0 0 x4.x34.D
flabel locali 24980 -560 25014 -526 0 FreeSans 400 0 0 0 x4.x34.Q_N
flabel locali 24980 -628 25014 -594 0 FreeSans 400 0 0 0 x4.x34.Q_N
flabel locali 24980 -900 25014 -866 0 FreeSans 400 0 0 0 x4.x34.Q_N
flabel metal1 22956 -1002 22990 -968 0 FreeSans 200 0 0 0 x4.x34.VGND
flabel metal1 22956 -458 22990 -424 0 FreeSans 200 0 0 0 x4.x34.VPWR
flabel nwell 22956 -458 22990 -424 3 FreeSans 400 0 0 0 x4.x34.VPB
flabel nwell 22973 -441 22973 -441 0 FreeSans 200 0 0 0 x4.x34.VPB
flabel pwell 22956 -1002 22990 -968 3 FreeSans 400 0 0 0 x4.x34.VNB
flabel pwell 22973 -985 22973 -985 0 FreeSans 200 0 0 0 x4.x34.VNB
rlabel comment 22927 -985 22927 -985 4 x4.x34.dfbbn_1
rlabel locali 24383 -838 24492 -772 1 x4.x34.SET_B
rlabel metal1 24430 -801 24488 -792 1 x4.x34.SET_B
rlabel metal1 24430 -838 24488 -829 1 x4.x34.SET_B
rlabel metal1 23680 -801 23738 -792 1 x4.x34.SET_B
rlabel metal1 23680 -829 24488 -801 1 x4.x34.SET_B
rlabel metal1 23680 -838 23738 -829 1 x4.x34.SET_B
rlabel metal1 22927 -1033 25319 -937 1 x4.x34.VGND
rlabel metal1 22927 -489 25319 -393 1 x4.x34.VPWR
flabel locali 21024 -1453 21058 -1419 0 FreeSans 400 0 0 0 x4.x32.RESET_B
flabel locali 22864 -1691 22898 -1657 7 FreeSans 400 0 0 0 x4.x32.VGND
flabel locali 22864 -1453 22898 -1419 0 FreeSans 400 0 0 0 x4.x32.CLK_N
flabel locali 22864 -1385 22898 -1351 0 FreeSans 400 0 0 0 x4.x32.CLK_N
flabel locali 22128 -1521 22162 -1487 0 FreeSans 400 0 0 0 x4.x32.SET_B
flabel locali 20564 -1589 20598 -1555 0 FreeSans 400 0 0 0 x4.x32.Q
flabel locali 20564 -1317 20598 -1283 0 FreeSans 400 0 0 0 x4.x32.Q
flabel locali 20564 -1249 20598 -1215 0 FreeSans 400 0 0 0 x4.x32.Q
flabel locali 22864 -1147 22898 -1113 7 FreeSans 400 0 0 0 x4.x32.VPWR
flabel locali 22496 -1453 22530 -1419 0 FreeSans 200 0 0 0 x4.x32.D
flabel locali 22496 -1385 22530 -1351 0 FreeSans 200 0 0 0 x4.x32.D
flabel locali 20840 -1249 20874 -1215 0 FreeSans 400 0 0 0 x4.x32.Q_N
flabel locali 20840 -1317 20874 -1283 0 FreeSans 400 0 0 0 x4.x32.Q_N
flabel locali 20840 -1589 20874 -1555 0 FreeSans 400 0 0 0 x4.x32.Q_N
flabel metal1 22864 -1691 22898 -1657 0 FreeSans 200 0 0 0 x4.x32.VGND
flabel metal1 22864 -1147 22898 -1113 0 FreeSans 200 0 0 0 x4.x32.VPWR
flabel nwell 22864 -1147 22898 -1113 7 FreeSans 400 0 0 0 x4.x32.VPB
flabel nwell 22881 -1130 22881 -1130 0 FreeSans 200 0 0 0 x4.x32.VPB
flabel pwell 22864 -1691 22898 -1657 7 FreeSans 400 0 0 0 x4.x32.VNB
flabel pwell 22881 -1674 22881 -1674 0 FreeSans 200 0 0 0 x4.x32.VNB
rlabel comment 22927 -1674 22927 -1674 6 x4.x32.dfbbn_1
rlabel locali 21362 -1527 21471 -1461 1 x4.x32.SET_B
rlabel metal1 21366 -1490 21424 -1481 1 x4.x32.SET_B
rlabel metal1 21366 -1527 21424 -1518 1 x4.x32.SET_B
rlabel metal1 22116 -1490 22174 -1481 1 x4.x32.SET_B
rlabel metal1 21366 -1518 22174 -1490 1 x4.x32.SET_B
rlabel metal1 22116 -1527 22174 -1518 1 x4.x32.SET_B
rlabel metal1 20535 -1722 22927 -1626 1 x4.x32.VGND
rlabel metal1 20535 -1178 22927 -1082 1 x4.x32.VPWR
flabel locali 22404 -764 22438 -730 0 FreeSans 400 0 0 0 x4.x31.RESET_B
flabel locali 20564 -1002 20598 -968 3 FreeSans 400 0 0 0 x4.x31.VGND
flabel locali 20564 -764 20598 -730 0 FreeSans 400 0 0 0 x4.x31.CLK_N
flabel locali 20564 -696 20598 -662 0 FreeSans 400 0 0 0 x4.x31.CLK_N
flabel locali 21300 -832 21334 -798 0 FreeSans 400 0 0 0 x4.x31.SET_B
flabel locali 22864 -900 22898 -866 0 FreeSans 400 0 0 0 x4.x31.Q
flabel locali 22864 -628 22898 -594 0 FreeSans 400 0 0 0 x4.x31.Q
flabel locali 22864 -560 22898 -526 0 FreeSans 400 0 0 0 x4.x31.Q
flabel locali 20564 -458 20598 -424 3 FreeSans 400 0 0 0 x4.x31.VPWR
flabel locali 20932 -764 20966 -730 0 FreeSans 200 0 0 0 x4.x31.D
flabel locali 20932 -696 20966 -662 0 FreeSans 200 0 0 0 x4.x31.D
flabel locali 22588 -560 22622 -526 0 FreeSans 400 0 0 0 x4.x31.Q_N
flabel locali 22588 -628 22622 -594 0 FreeSans 400 0 0 0 x4.x31.Q_N
flabel locali 22588 -900 22622 -866 0 FreeSans 400 0 0 0 x4.x31.Q_N
flabel metal1 20564 -1002 20598 -968 0 FreeSans 200 0 0 0 x4.x31.VGND
flabel metal1 20564 -458 20598 -424 0 FreeSans 200 0 0 0 x4.x31.VPWR
flabel nwell 20564 -458 20598 -424 3 FreeSans 400 0 0 0 x4.x31.VPB
flabel nwell 20581 -441 20581 -441 0 FreeSans 200 0 0 0 x4.x31.VPB
flabel pwell 20564 -1002 20598 -968 3 FreeSans 400 0 0 0 x4.x31.VNB
flabel pwell 20581 -985 20581 -985 0 FreeSans 200 0 0 0 x4.x31.VNB
rlabel comment 20535 -985 20535 -985 4 x4.x31.dfbbn_1
rlabel locali 21991 -838 22100 -772 1 x4.x31.SET_B
rlabel metal1 22038 -801 22096 -792 1 x4.x31.SET_B
rlabel metal1 22038 -838 22096 -829 1 x4.x31.SET_B
rlabel metal1 21288 -801 21346 -792 1 x4.x31.SET_B
rlabel metal1 21288 -829 22096 -801 1 x4.x31.SET_B
rlabel metal1 21288 -838 21346 -829 1 x4.x31.SET_B
rlabel metal1 20535 -1033 22927 -937 1 x4.x31.VGND
rlabel metal1 20535 -489 22927 -393 1 x4.x31.VPWR
flabel locali 14187 1066 14221 1100 0 FreeSans 200 0 0 0 x4.x30.A
flabel locali 14095 1066 14129 1100 0 FreeSans 200 0 0 0 x4.x30.A
flabel locali 15750 1066 15784 1100 0 FreeSans 200 0 0 0 x4.x30.X
flabel locali 15750 1134 15784 1168 0 FreeSans 200 0 0 0 x4.x30.X
flabel pwell 13819 828 13853 862 0 FreeSans 200 0 0 0 x4.x30.VNB
flabel nwell 13819 1372 13853 1406 0 FreeSans 200 0 0 0 x4.x30.VPB
flabel metal1 13819 828 13853 862 0 FreeSans 200 0 0 0 x4.x30.VGND
flabel metal1 13819 1372 13853 1406 0 FreeSans 200 0 0 0 x4.x30.VPWR
rlabel comment 13789 845 13789 845 4 x4.x30.buf_16
rlabel metal1 13789 797 15813 893 1 x4.x30.VGND
rlabel metal1 13789 1341 15813 1437 1 x4.x30.VPWR
flabel locali 18632 -1453 18666 -1419 0 FreeSans 400 0 0 0 x4.x29.RESET_B
flabel locali 20472 -1691 20506 -1657 7 FreeSans 400 0 0 0 x4.x29.VGND
flabel locali 20472 -1453 20506 -1419 0 FreeSans 400 0 0 0 x4.x29.CLK_N
flabel locali 20472 -1385 20506 -1351 0 FreeSans 400 0 0 0 x4.x29.CLK_N
flabel locali 19736 -1521 19770 -1487 0 FreeSans 400 0 0 0 x4.x29.SET_B
flabel locali 18172 -1589 18206 -1555 0 FreeSans 400 0 0 0 x4.x29.Q
flabel locali 18172 -1317 18206 -1283 0 FreeSans 400 0 0 0 x4.x29.Q
flabel locali 18172 -1249 18206 -1215 0 FreeSans 400 0 0 0 x4.x29.Q
flabel locali 20472 -1147 20506 -1113 7 FreeSans 400 0 0 0 x4.x29.VPWR
flabel locali 20104 -1453 20138 -1419 0 FreeSans 200 0 0 0 x4.x29.D
flabel locali 20104 -1385 20138 -1351 0 FreeSans 200 0 0 0 x4.x29.D
flabel locali 18448 -1249 18482 -1215 0 FreeSans 400 0 0 0 x4.x29.Q_N
flabel locali 18448 -1317 18482 -1283 0 FreeSans 400 0 0 0 x4.x29.Q_N
flabel locali 18448 -1589 18482 -1555 0 FreeSans 400 0 0 0 x4.x29.Q_N
flabel metal1 20472 -1691 20506 -1657 0 FreeSans 200 0 0 0 x4.x29.VGND
flabel metal1 20472 -1147 20506 -1113 0 FreeSans 200 0 0 0 x4.x29.VPWR
flabel nwell 20472 -1147 20506 -1113 7 FreeSans 400 0 0 0 x4.x29.VPB
flabel nwell 20489 -1130 20489 -1130 0 FreeSans 200 0 0 0 x4.x29.VPB
flabel pwell 20472 -1691 20506 -1657 7 FreeSans 400 0 0 0 x4.x29.VNB
flabel pwell 20489 -1674 20489 -1674 0 FreeSans 200 0 0 0 x4.x29.VNB
rlabel comment 20535 -1674 20535 -1674 6 x4.x29.dfbbn_1
rlabel locali 18970 -1527 19079 -1461 1 x4.x29.SET_B
rlabel metal1 18974 -1490 19032 -1481 1 x4.x29.SET_B
rlabel metal1 18974 -1527 19032 -1518 1 x4.x29.SET_B
rlabel metal1 19724 -1490 19782 -1481 1 x4.x29.SET_B
rlabel metal1 18974 -1518 19782 -1490 1 x4.x29.SET_B
rlabel metal1 19724 -1527 19782 -1518 1 x4.x29.SET_B
rlabel metal1 18143 -1722 20535 -1626 1 x4.x29.VGND
rlabel metal1 18143 -1178 20535 -1082 1 x4.x29.VPWR
flabel locali 20012 -764 20046 -730 0 FreeSans 400 0 0 0 x4.x28.RESET_B
flabel locali 18172 -1002 18206 -968 3 FreeSans 400 0 0 0 x4.x28.VGND
flabel locali 18172 -764 18206 -730 0 FreeSans 400 0 0 0 x4.x28.CLK_N
flabel locali 18172 -696 18206 -662 0 FreeSans 400 0 0 0 x4.x28.CLK_N
flabel locali 18908 -832 18942 -798 0 FreeSans 400 0 0 0 x4.x28.SET_B
flabel locali 20472 -900 20506 -866 0 FreeSans 400 0 0 0 x4.x28.Q
flabel locali 20472 -628 20506 -594 0 FreeSans 400 0 0 0 x4.x28.Q
flabel locali 20472 -560 20506 -526 0 FreeSans 400 0 0 0 x4.x28.Q
flabel locali 18172 -458 18206 -424 3 FreeSans 400 0 0 0 x4.x28.VPWR
flabel locali 18540 -764 18574 -730 0 FreeSans 200 0 0 0 x4.x28.D
flabel locali 18540 -696 18574 -662 0 FreeSans 200 0 0 0 x4.x28.D
flabel locali 20196 -560 20230 -526 0 FreeSans 400 0 0 0 x4.x28.Q_N
flabel locali 20196 -628 20230 -594 0 FreeSans 400 0 0 0 x4.x28.Q_N
flabel locali 20196 -900 20230 -866 0 FreeSans 400 0 0 0 x4.x28.Q_N
flabel metal1 18172 -1002 18206 -968 0 FreeSans 200 0 0 0 x4.x28.VGND
flabel metal1 18172 -458 18206 -424 0 FreeSans 200 0 0 0 x4.x28.VPWR
flabel nwell 18172 -458 18206 -424 3 FreeSans 400 0 0 0 x4.x28.VPB
flabel nwell 18189 -441 18189 -441 0 FreeSans 200 0 0 0 x4.x28.VPB
flabel pwell 18172 -1002 18206 -968 3 FreeSans 400 0 0 0 x4.x28.VNB
flabel pwell 18189 -985 18189 -985 0 FreeSans 200 0 0 0 x4.x28.VNB
rlabel comment 18143 -985 18143 -985 4 x4.x28.dfbbn_1
rlabel locali 19599 -838 19708 -772 1 x4.x28.SET_B
rlabel metal1 19646 -801 19704 -792 1 x4.x28.SET_B
rlabel metal1 19646 -838 19704 -829 1 x4.x28.SET_B
rlabel metal1 18896 -801 18954 -792 1 x4.x28.SET_B
rlabel metal1 18896 -829 19704 -801 1 x4.x28.SET_B
rlabel metal1 18896 -838 18954 -829 1 x4.x28.SET_B
rlabel metal1 18143 -1033 20535 -937 1 x4.x28.VGND
rlabel metal1 18143 -489 20535 -393 1 x4.x28.VPWR
flabel metal1 13267 1372 13301 1406 0 FreeSans 200 0 0 0 x4.x27.VPWR
flabel metal1 13267 828 13301 862 0 FreeSans 200 0 0 0 x4.x27.VGND
flabel locali 13543 1066 13577 1100 0 FreeSans 200 0 0 0 x4.x27.X
flabel locali 13543 1134 13577 1168 0 FreeSans 200 0 0 0 x4.x27.X
flabel locali 13543 998 13577 1032 0 FreeSans 200 0 0 0 x4.x27.X
flabel locali 13267 1372 13301 1406 0 FreeSans 200 0 0 0 x4.x27.VPWR
flabel locali 13267 828 13301 862 0 FreeSans 200 0 0 0 x4.x27.VGND
flabel locali 13267 1066 13301 1100 0 FreeSans 200 0 0 0 x4.x27.A
flabel nwell 13267 1372 13301 1406 0 FreeSans 200 0 0 0 x4.x27.VPB
flabel pwell 13267 828 13301 862 0 FreeSans 200 0 0 0 x4.x27.VNB
rlabel comment 13237 845 13237 845 4 x4.x27.buf_4
rlabel metal1 13237 797 13789 893 1 x4.x27.VGND
rlabel metal1 13237 1341 13789 1437 1 x4.x27.VPWR
flabel locali 16240 -1453 16274 -1419 0 FreeSans 400 0 0 0 x4.x26.RESET_B
flabel locali 18080 -1691 18114 -1657 7 FreeSans 400 0 0 0 x4.x26.VGND
flabel locali 18080 -1453 18114 -1419 0 FreeSans 400 0 0 0 x4.x26.CLK_N
flabel locali 18080 -1385 18114 -1351 0 FreeSans 400 0 0 0 x4.x26.CLK_N
flabel locali 17344 -1521 17378 -1487 0 FreeSans 400 0 0 0 x4.x26.SET_B
flabel locali 15780 -1589 15814 -1555 0 FreeSans 400 0 0 0 x4.x26.Q
flabel locali 15780 -1317 15814 -1283 0 FreeSans 400 0 0 0 x4.x26.Q
flabel locali 15780 -1249 15814 -1215 0 FreeSans 400 0 0 0 x4.x26.Q
flabel locali 18080 -1147 18114 -1113 7 FreeSans 400 0 0 0 x4.x26.VPWR
flabel locali 17712 -1453 17746 -1419 0 FreeSans 200 0 0 0 x4.x26.D
flabel locali 17712 -1385 17746 -1351 0 FreeSans 200 0 0 0 x4.x26.D
flabel locali 16056 -1249 16090 -1215 0 FreeSans 400 0 0 0 x4.x26.Q_N
flabel locali 16056 -1317 16090 -1283 0 FreeSans 400 0 0 0 x4.x26.Q_N
flabel locali 16056 -1589 16090 -1555 0 FreeSans 400 0 0 0 x4.x26.Q_N
flabel metal1 18080 -1691 18114 -1657 0 FreeSans 200 0 0 0 x4.x26.VGND
flabel metal1 18080 -1147 18114 -1113 0 FreeSans 200 0 0 0 x4.x26.VPWR
flabel nwell 18080 -1147 18114 -1113 7 FreeSans 400 0 0 0 x4.x26.VPB
flabel nwell 18097 -1130 18097 -1130 0 FreeSans 200 0 0 0 x4.x26.VPB
flabel pwell 18080 -1691 18114 -1657 7 FreeSans 400 0 0 0 x4.x26.VNB
flabel pwell 18097 -1674 18097 -1674 0 FreeSans 200 0 0 0 x4.x26.VNB
rlabel comment 18143 -1674 18143 -1674 6 x4.x26.dfbbn_1
rlabel locali 16578 -1527 16687 -1461 1 x4.x26.SET_B
rlabel metal1 16582 -1490 16640 -1481 1 x4.x26.SET_B
rlabel metal1 16582 -1527 16640 -1518 1 x4.x26.SET_B
rlabel metal1 17332 -1490 17390 -1481 1 x4.x26.SET_B
rlabel metal1 16582 -1518 17390 -1490 1 x4.x26.SET_B
rlabel metal1 17332 -1527 17390 -1518 1 x4.x26.SET_B
rlabel metal1 15751 -1722 18143 -1626 1 x4.x26.VGND
rlabel metal1 15751 -1178 18143 -1082 1 x4.x26.VPWR
flabel locali 17620 -764 17654 -730 0 FreeSans 400 0 0 0 x4.x25.RESET_B
flabel locali 15780 -1002 15814 -968 3 FreeSans 400 0 0 0 x4.x25.VGND
flabel locali 15780 -764 15814 -730 0 FreeSans 400 0 0 0 x4.x25.CLK_N
flabel locali 15780 -696 15814 -662 0 FreeSans 400 0 0 0 x4.x25.CLK_N
flabel locali 16516 -832 16550 -798 0 FreeSans 400 0 0 0 x4.x25.SET_B
flabel locali 18080 -900 18114 -866 0 FreeSans 400 0 0 0 x4.x25.Q
flabel locali 18080 -628 18114 -594 0 FreeSans 400 0 0 0 x4.x25.Q
flabel locali 18080 -560 18114 -526 0 FreeSans 400 0 0 0 x4.x25.Q
flabel locali 15780 -458 15814 -424 3 FreeSans 400 0 0 0 x4.x25.VPWR
flabel locali 16148 -764 16182 -730 0 FreeSans 200 0 0 0 x4.x25.D
flabel locali 16148 -696 16182 -662 0 FreeSans 200 0 0 0 x4.x25.D
flabel locali 17804 -560 17838 -526 0 FreeSans 400 0 0 0 x4.x25.Q_N
flabel locali 17804 -628 17838 -594 0 FreeSans 400 0 0 0 x4.x25.Q_N
flabel locali 17804 -900 17838 -866 0 FreeSans 400 0 0 0 x4.x25.Q_N
flabel metal1 15780 -1002 15814 -968 0 FreeSans 200 0 0 0 x4.x25.VGND
flabel metal1 15780 -458 15814 -424 0 FreeSans 200 0 0 0 x4.x25.VPWR
flabel nwell 15780 -458 15814 -424 3 FreeSans 400 0 0 0 x4.x25.VPB
flabel nwell 15797 -441 15797 -441 0 FreeSans 200 0 0 0 x4.x25.VPB
flabel pwell 15780 -1002 15814 -968 3 FreeSans 400 0 0 0 x4.x25.VNB
flabel pwell 15797 -985 15797 -985 0 FreeSans 200 0 0 0 x4.x25.VNB
rlabel comment 15751 -985 15751 -985 4 x4.x25.dfbbn_1
rlabel locali 17207 -838 17316 -772 1 x4.x25.SET_B
rlabel metal1 17254 -801 17312 -792 1 x4.x25.SET_B
rlabel metal1 17254 -838 17312 -829 1 x4.x25.SET_B
rlabel metal1 16504 -801 16562 -792 1 x4.x25.SET_B
rlabel metal1 16504 -829 17312 -801 1 x4.x25.SET_B
rlabel metal1 16504 -838 16562 -829 1 x4.x25.SET_B
rlabel metal1 15751 -1033 18143 -937 1 x4.x25.VGND
rlabel metal1 15751 -489 18143 -393 1 x4.x25.VPWR
flabel locali 13848 -1453 13882 -1419 0 FreeSans 400 0 0 0 x4.x24.RESET_B
flabel locali 15688 -1691 15722 -1657 7 FreeSans 400 0 0 0 x4.x24.VGND
flabel locali 15688 -1453 15722 -1419 0 FreeSans 400 0 0 0 x4.x24.CLK_N
flabel locali 15688 -1385 15722 -1351 0 FreeSans 400 0 0 0 x4.x24.CLK_N
flabel locali 14952 -1521 14986 -1487 0 FreeSans 400 0 0 0 x4.x24.SET_B
flabel locali 13388 -1589 13422 -1555 0 FreeSans 400 0 0 0 x4.x24.Q
flabel locali 13388 -1317 13422 -1283 0 FreeSans 400 0 0 0 x4.x24.Q
flabel locali 13388 -1249 13422 -1215 0 FreeSans 400 0 0 0 x4.x24.Q
flabel locali 15688 -1147 15722 -1113 7 FreeSans 400 0 0 0 x4.x24.VPWR
flabel locali 15320 -1453 15354 -1419 0 FreeSans 200 0 0 0 x4.x24.D
flabel locali 15320 -1385 15354 -1351 0 FreeSans 200 0 0 0 x4.x24.D
flabel locali 13664 -1249 13698 -1215 0 FreeSans 400 0 0 0 x4.x24.Q_N
flabel locali 13664 -1317 13698 -1283 0 FreeSans 400 0 0 0 x4.x24.Q_N
flabel locali 13664 -1589 13698 -1555 0 FreeSans 400 0 0 0 x4.x24.Q_N
flabel metal1 15688 -1691 15722 -1657 0 FreeSans 200 0 0 0 x4.x24.VGND
flabel metal1 15688 -1147 15722 -1113 0 FreeSans 200 0 0 0 x4.x24.VPWR
flabel nwell 15688 -1147 15722 -1113 7 FreeSans 400 0 0 0 x4.x24.VPB
flabel nwell 15705 -1130 15705 -1130 0 FreeSans 200 0 0 0 x4.x24.VPB
flabel pwell 15688 -1691 15722 -1657 7 FreeSans 400 0 0 0 x4.x24.VNB
flabel pwell 15705 -1674 15705 -1674 0 FreeSans 200 0 0 0 x4.x24.VNB
rlabel comment 15751 -1674 15751 -1674 6 x4.x24.dfbbn_1
rlabel locali 14186 -1527 14295 -1461 1 x4.x24.SET_B
rlabel metal1 14190 -1490 14248 -1481 1 x4.x24.SET_B
rlabel metal1 14190 -1527 14248 -1518 1 x4.x24.SET_B
rlabel metal1 14940 -1490 14998 -1481 1 x4.x24.SET_B
rlabel metal1 14190 -1518 14998 -1490 1 x4.x24.SET_B
rlabel metal1 14940 -1527 14998 -1518 1 x4.x24.SET_B
rlabel metal1 13359 -1722 15751 -1626 1 x4.x24.VGND
rlabel metal1 13359 -1178 15751 -1082 1 x4.x24.VPWR
flabel locali 15228 -764 15262 -730 0 FreeSans 400 0 0 0 x4.x23.RESET_B
flabel locali 13388 -1002 13422 -968 3 FreeSans 400 0 0 0 x4.x23.VGND
flabel locali 13388 -764 13422 -730 0 FreeSans 400 0 0 0 x4.x23.CLK_N
flabel locali 13388 -696 13422 -662 0 FreeSans 400 0 0 0 x4.x23.CLK_N
flabel locali 14124 -832 14158 -798 0 FreeSans 400 0 0 0 x4.x23.SET_B
flabel locali 15688 -900 15722 -866 0 FreeSans 400 0 0 0 x4.x23.Q
flabel locali 15688 -628 15722 -594 0 FreeSans 400 0 0 0 x4.x23.Q
flabel locali 15688 -560 15722 -526 0 FreeSans 400 0 0 0 x4.x23.Q
flabel locali 13388 -458 13422 -424 3 FreeSans 400 0 0 0 x4.x23.VPWR
flabel locali 13756 -764 13790 -730 0 FreeSans 200 0 0 0 x4.x23.D
flabel locali 13756 -696 13790 -662 0 FreeSans 200 0 0 0 x4.x23.D
flabel locali 15412 -560 15446 -526 0 FreeSans 400 0 0 0 x4.x23.Q_N
flabel locali 15412 -628 15446 -594 0 FreeSans 400 0 0 0 x4.x23.Q_N
flabel locali 15412 -900 15446 -866 0 FreeSans 400 0 0 0 x4.x23.Q_N
flabel metal1 13388 -1002 13422 -968 0 FreeSans 200 0 0 0 x4.x23.VGND
flabel metal1 13388 -458 13422 -424 0 FreeSans 200 0 0 0 x4.x23.VPWR
flabel nwell 13388 -458 13422 -424 3 FreeSans 400 0 0 0 x4.x23.VPB
flabel nwell 13405 -441 13405 -441 0 FreeSans 200 0 0 0 x4.x23.VPB
flabel pwell 13388 -1002 13422 -968 3 FreeSans 400 0 0 0 x4.x23.VNB
flabel pwell 13405 -985 13405 -985 0 FreeSans 200 0 0 0 x4.x23.VNB
rlabel comment 13359 -985 13359 -985 4 x4.x23.dfbbn_1
rlabel locali 14815 -838 14924 -772 1 x4.x23.SET_B
rlabel metal1 14862 -801 14920 -792 1 x4.x23.SET_B
rlabel metal1 14862 -838 14920 -829 1 x4.x23.SET_B
rlabel metal1 14112 -801 14170 -792 1 x4.x23.SET_B
rlabel metal1 14112 -829 14920 -801 1 x4.x23.SET_B
rlabel metal1 14112 -838 14170 -829 1 x4.x23.SET_B
rlabel metal1 13359 -1033 15751 -937 1 x4.x23.VGND
rlabel metal1 13359 -489 15751 -393 1 x4.x23.VPWR
flabel metal1 12992 828 13026 862 0 FreeSans 200 0 0 0 x4.x22.VGND
flabel metal1 12990 1372 13024 1406 0 FreeSans 200 0 0 0 x4.x22.VPWR
flabel locali 12990 1372 13024 1406 0 FreeSans 200 0 0 0 x4.x22.VPWR
flabel locali 12992 828 13026 862 0 FreeSans 200 0 0 0 x4.x22.VGND
flabel locali 13172 930 13206 964 0 FreeSans 200 0 0 0 x4.x22.X
flabel locali 13172 1202 13206 1236 0 FreeSans 200 0 0 0 x4.x22.X
flabel locali 13172 1270 13206 1304 0 FreeSans 200 0 0 0 x4.x22.X
flabel locali 12990 1066 13024 1100 0 FreeSans 200 0 0 0 x4.x22.A
flabel nwell 12990 1372 13024 1406 0 FreeSans 200 0 0 0 x4.x22.VPB
flabel pwell 12992 828 13026 862 0 FreeSans 200 0 0 0 x4.x22.VNB
rlabel comment 12961 845 12961 845 4 x4.x22.buf_1
rlabel metal1 12961 797 13237 893 1 x4.x22.VGND
rlabel metal1 12961 1341 13237 1437 1 x4.x22.VPWR
flabel locali 11456 -1453 11490 -1419 0 FreeSans 400 0 0 0 x4.x21.RESET_B
flabel locali 13296 -1691 13330 -1657 7 FreeSans 400 0 0 0 x4.x21.VGND
flabel locali 13296 -1453 13330 -1419 0 FreeSans 400 0 0 0 x4.x21.CLK_N
flabel locali 13296 -1385 13330 -1351 0 FreeSans 400 0 0 0 x4.x21.CLK_N
flabel locali 12560 -1521 12594 -1487 0 FreeSans 400 0 0 0 x4.x21.SET_B
flabel locali 10996 -1589 11030 -1555 0 FreeSans 400 0 0 0 x4.x21.Q
flabel locali 10996 -1317 11030 -1283 0 FreeSans 400 0 0 0 x4.x21.Q
flabel locali 10996 -1249 11030 -1215 0 FreeSans 400 0 0 0 x4.x21.Q
flabel locali 13296 -1147 13330 -1113 7 FreeSans 400 0 0 0 x4.x21.VPWR
flabel locali 12928 -1453 12962 -1419 0 FreeSans 200 0 0 0 x4.x21.D
flabel locali 12928 -1385 12962 -1351 0 FreeSans 200 0 0 0 x4.x21.D
flabel locali 11272 -1249 11306 -1215 0 FreeSans 400 0 0 0 x4.x21.Q_N
flabel locali 11272 -1317 11306 -1283 0 FreeSans 400 0 0 0 x4.x21.Q_N
flabel locali 11272 -1589 11306 -1555 0 FreeSans 400 0 0 0 x4.x21.Q_N
flabel metal1 13296 -1691 13330 -1657 0 FreeSans 200 0 0 0 x4.x21.VGND
flabel metal1 13296 -1147 13330 -1113 0 FreeSans 200 0 0 0 x4.x21.VPWR
flabel nwell 13296 -1147 13330 -1113 7 FreeSans 400 0 0 0 x4.x21.VPB
flabel nwell 13313 -1130 13313 -1130 0 FreeSans 200 0 0 0 x4.x21.VPB
flabel pwell 13296 -1691 13330 -1657 7 FreeSans 400 0 0 0 x4.x21.VNB
flabel pwell 13313 -1674 13313 -1674 0 FreeSans 200 0 0 0 x4.x21.VNB
rlabel comment 13359 -1674 13359 -1674 6 x4.x21.dfbbn_1
rlabel locali 11794 -1527 11903 -1461 1 x4.x21.SET_B
rlabel metal1 11798 -1490 11856 -1481 1 x4.x21.SET_B
rlabel metal1 11798 -1527 11856 -1518 1 x4.x21.SET_B
rlabel metal1 12548 -1490 12606 -1481 1 x4.x21.SET_B
rlabel metal1 11798 -1518 12606 -1490 1 x4.x21.SET_B
rlabel metal1 12548 -1527 12606 -1518 1 x4.x21.SET_B
rlabel metal1 10967 -1722 13359 -1626 1 x4.x21.VGND
rlabel metal1 10967 -1178 13359 -1082 1 x4.x21.VPWR
flabel metal1 25125 -314 25159 -280 0 FreeSans 200 0 0 0 x4.x20.VGND
flabel metal1 25125 230 25159 264 0 FreeSans 200 0 0 0 x4.x20.VPWR
flabel locali 24481 -8 24515 26 0 FreeSans 250 0 0 0 x4.x20.S
flabel locali 24573 -8 24607 26 0 FreeSans 250 0 0 0 x4.x20.S
flabel locali 24665 -144 24699 -110 0 FreeSans 250 0 0 0 x4.x20.A1
flabel locali 24665 -76 24699 -42 0 FreeSans 250 0 0 0 x4.x20.A1
flabel locali 24757 -76 24791 -42 0 FreeSans 250 0 0 0 x4.x20.A0
flabel locali 25125 -212 25159 -178 0 FreeSans 250 0 0 0 x4.x20.X
flabel locali 25125 60 25159 94 0 FreeSans 250 0 0 0 x4.x20.X
flabel locali 25125 128 25159 162 0 FreeSans 250 0 0 0 x4.x20.X
flabel nwell 25081 230 25115 264 0 FreeSans 250 0 0 0 x4.x20.VPB
flabel pwell 25071 -314 25105 -280 0 FreeSans 250 0 0 0 x4.x20.VNB
rlabel comment 25189 -297 25189 -297 6 x4.x20.mux2_1
rlabel metal1 24361 -345 25189 -249 1 x4.x20.VGND
rlabel metal1 24361 199 25189 295 1 x4.x20.VPWR
flabel locali 12836 -764 12870 -730 0 FreeSans 400 0 0 0 x4.x19.RESET_B
flabel locali 10996 -1002 11030 -968 3 FreeSans 400 0 0 0 x4.x19.VGND
flabel locali 10996 -764 11030 -730 0 FreeSans 400 0 0 0 x4.x19.CLK_N
flabel locali 10996 -696 11030 -662 0 FreeSans 400 0 0 0 x4.x19.CLK_N
flabel locali 11732 -832 11766 -798 0 FreeSans 400 0 0 0 x4.x19.SET_B
flabel locali 13296 -900 13330 -866 0 FreeSans 400 0 0 0 x4.x19.Q
flabel locali 13296 -628 13330 -594 0 FreeSans 400 0 0 0 x4.x19.Q
flabel locali 13296 -560 13330 -526 0 FreeSans 400 0 0 0 x4.x19.Q
flabel locali 10996 -458 11030 -424 3 FreeSans 400 0 0 0 x4.x19.VPWR
flabel locali 11364 -764 11398 -730 0 FreeSans 200 0 0 0 x4.x19.D
flabel locali 11364 -696 11398 -662 0 FreeSans 200 0 0 0 x4.x19.D
flabel locali 13020 -560 13054 -526 0 FreeSans 400 0 0 0 x4.x19.Q_N
flabel locali 13020 -628 13054 -594 0 FreeSans 400 0 0 0 x4.x19.Q_N
flabel locali 13020 -900 13054 -866 0 FreeSans 400 0 0 0 x4.x19.Q_N
flabel metal1 10996 -1002 11030 -968 0 FreeSans 200 0 0 0 x4.x19.VGND
flabel metal1 10996 -458 11030 -424 0 FreeSans 200 0 0 0 x4.x19.VPWR
flabel nwell 10996 -458 11030 -424 3 FreeSans 400 0 0 0 x4.x19.VPB
flabel nwell 11013 -441 11013 -441 0 FreeSans 200 0 0 0 x4.x19.VPB
flabel pwell 10996 -1002 11030 -968 3 FreeSans 400 0 0 0 x4.x19.VNB
flabel pwell 11013 -985 11013 -985 0 FreeSans 200 0 0 0 x4.x19.VNB
rlabel comment 10967 -985 10967 -985 4 x4.x19.dfbbn_1
rlabel locali 12423 -838 12532 -772 1 x4.x19.SET_B
rlabel metal1 12470 -801 12528 -792 1 x4.x19.SET_B
rlabel metal1 12470 -838 12528 -829 1 x4.x19.SET_B
rlabel metal1 11720 -801 11778 -792 1 x4.x19.SET_B
rlabel metal1 11720 -829 12528 -801 1 x4.x19.SET_B
rlabel metal1 11720 -838 11778 -829 1 x4.x19.SET_B
rlabel metal1 10967 -1033 13359 -937 1 x4.x19.VGND
rlabel metal1 10967 -489 13359 -393 1 x4.x19.VPWR
flabel metal1 22957 -314 22991 -280 0 FreeSans 200 0 0 0 x4.x18.VGND
flabel metal1 22957 230 22991 264 0 FreeSans 200 0 0 0 x4.x18.VPWR
flabel locali 23601 -8 23635 26 0 FreeSans 250 0 0 0 x4.x18.S
flabel locali 23509 -8 23543 26 0 FreeSans 250 0 0 0 x4.x18.S
flabel locali 23417 -144 23451 -110 0 FreeSans 250 0 0 0 x4.x18.A1
flabel locali 23417 -76 23451 -42 0 FreeSans 250 0 0 0 x4.x18.A1
flabel locali 23325 -76 23359 -42 0 FreeSans 250 0 0 0 x4.x18.A0
flabel locali 22957 -212 22991 -178 0 FreeSans 250 0 0 0 x4.x18.X
flabel locali 22957 60 22991 94 0 FreeSans 250 0 0 0 x4.x18.X
flabel locali 22957 128 22991 162 0 FreeSans 250 0 0 0 x4.x18.X
flabel nwell 23001 230 23035 264 0 FreeSans 250 0 0 0 x4.x18.VPB
flabel pwell 23011 -314 23045 -280 0 FreeSans 250 0 0 0 x4.x18.VNB
rlabel comment 22927 -297 22927 -297 4 x4.x18.mux2_1
rlabel metal1 22927 -345 23755 -249 1 x4.x18.VGND
rlabel metal1 22927 199 23755 295 1 x4.x18.VPWR
flabel metal1 22731 -314 22765 -280 0 FreeSans 200 0 0 0 x4.x17.VGND
flabel metal1 22731 230 22765 264 0 FreeSans 200 0 0 0 x4.x17.VPWR
flabel locali 22087 -8 22121 26 0 FreeSans 250 0 0 0 x4.x17.S
flabel locali 22179 -8 22213 26 0 FreeSans 250 0 0 0 x4.x17.S
flabel locali 22271 -144 22305 -110 0 FreeSans 250 0 0 0 x4.x17.A1
flabel locali 22271 -76 22305 -42 0 FreeSans 250 0 0 0 x4.x17.A1
flabel locali 22363 -76 22397 -42 0 FreeSans 250 0 0 0 x4.x17.A0
flabel locali 22731 -212 22765 -178 0 FreeSans 250 0 0 0 x4.x17.X
flabel locali 22731 60 22765 94 0 FreeSans 250 0 0 0 x4.x17.X
flabel locali 22731 128 22765 162 0 FreeSans 250 0 0 0 x4.x17.X
flabel nwell 22687 230 22721 264 0 FreeSans 250 0 0 0 x4.x17.VPB
flabel pwell 22677 -314 22711 -280 0 FreeSans 250 0 0 0 x4.x17.VNB
rlabel comment 22795 -297 22795 -297 6 x4.x17.mux2_1
rlabel metal1 21967 -345 22795 -249 1 x4.x17.VGND
rlabel metal1 21967 199 22795 295 1 x4.x17.VPWR
flabel metal1 20565 -314 20599 -280 0 FreeSans 200 0 0 0 x4.x16.VGND
flabel metal1 20565 230 20599 264 0 FreeSans 200 0 0 0 x4.x16.VPWR
flabel locali 21209 -8 21243 26 0 FreeSans 250 0 0 0 x4.x16.S
flabel locali 21117 -8 21151 26 0 FreeSans 250 0 0 0 x4.x16.S
flabel locali 21025 -144 21059 -110 0 FreeSans 250 0 0 0 x4.x16.A1
flabel locali 21025 -76 21059 -42 0 FreeSans 250 0 0 0 x4.x16.A1
flabel locali 20933 -76 20967 -42 0 FreeSans 250 0 0 0 x4.x16.A0
flabel locali 20565 -212 20599 -178 0 FreeSans 250 0 0 0 x4.x16.X
flabel locali 20565 60 20599 94 0 FreeSans 250 0 0 0 x4.x16.X
flabel locali 20565 128 20599 162 0 FreeSans 250 0 0 0 x4.x16.X
flabel nwell 20609 230 20643 264 0 FreeSans 250 0 0 0 x4.x16.VPB
flabel pwell 20619 -314 20653 -280 0 FreeSans 250 0 0 0 x4.x16.VNB
rlabel comment 20535 -297 20535 -297 4 x4.x16.mux2_1
rlabel metal1 20535 -345 21363 -249 1 x4.x16.VGND
rlabel metal1 20535 199 21363 295 1 x4.x16.VPWR
flabel metal1 20341 -314 20375 -280 0 FreeSans 200 0 0 0 x4.x15.VGND
flabel metal1 20341 230 20375 264 0 FreeSans 200 0 0 0 x4.x15.VPWR
flabel locali 19697 -8 19731 26 0 FreeSans 250 0 0 0 x4.x15.S
flabel locali 19789 -8 19823 26 0 FreeSans 250 0 0 0 x4.x15.S
flabel locali 19881 -144 19915 -110 0 FreeSans 250 0 0 0 x4.x15.A1
flabel locali 19881 -76 19915 -42 0 FreeSans 250 0 0 0 x4.x15.A1
flabel locali 19973 -76 20007 -42 0 FreeSans 250 0 0 0 x4.x15.A0
flabel locali 20341 -212 20375 -178 0 FreeSans 250 0 0 0 x4.x15.X
flabel locali 20341 60 20375 94 0 FreeSans 250 0 0 0 x4.x15.X
flabel locali 20341 128 20375 162 0 FreeSans 250 0 0 0 x4.x15.X
flabel nwell 20297 230 20331 264 0 FreeSans 250 0 0 0 x4.x15.VPB
flabel pwell 20287 -314 20321 -280 0 FreeSans 250 0 0 0 x4.x15.VNB
rlabel comment 20405 -297 20405 -297 6 x4.x15.mux2_1
rlabel metal1 19577 -345 20405 -249 1 x4.x15.VGND
rlabel metal1 19577 199 20405 295 1 x4.x15.VPWR
flabel metal1 18173 -314 18207 -280 0 FreeSans 200 0 0 0 x4.x14.VGND
flabel metal1 18173 230 18207 264 0 FreeSans 200 0 0 0 x4.x14.VPWR
flabel locali 18817 -8 18851 26 0 FreeSans 250 0 0 0 x4.x14.S
flabel locali 18725 -8 18759 26 0 FreeSans 250 0 0 0 x4.x14.S
flabel locali 18633 -144 18667 -110 0 FreeSans 250 0 0 0 x4.x14.A1
flabel locali 18633 -76 18667 -42 0 FreeSans 250 0 0 0 x4.x14.A1
flabel locali 18541 -76 18575 -42 0 FreeSans 250 0 0 0 x4.x14.A0
flabel locali 18173 -212 18207 -178 0 FreeSans 250 0 0 0 x4.x14.X
flabel locali 18173 60 18207 94 0 FreeSans 250 0 0 0 x4.x14.X
flabel locali 18173 128 18207 162 0 FreeSans 250 0 0 0 x4.x14.X
flabel nwell 18217 230 18251 264 0 FreeSans 250 0 0 0 x4.x14.VPB
flabel pwell 18227 -314 18261 -280 0 FreeSans 250 0 0 0 x4.x14.VNB
rlabel comment 18143 -297 18143 -297 4 x4.x14.mux2_1
rlabel metal1 18143 -345 18971 -249 1 x4.x14.VGND
rlabel metal1 18143 199 18971 295 1 x4.x14.VPWR
flabel metal1 17949 -314 17983 -280 0 FreeSans 200 0 0 0 x4.x13.VGND
flabel metal1 17949 230 17983 264 0 FreeSans 200 0 0 0 x4.x13.VPWR
flabel locali 17305 -8 17339 26 0 FreeSans 250 0 0 0 x4.x13.S
flabel locali 17397 -8 17431 26 0 FreeSans 250 0 0 0 x4.x13.S
flabel locali 17489 -144 17523 -110 0 FreeSans 250 0 0 0 x4.x13.A1
flabel locali 17489 -76 17523 -42 0 FreeSans 250 0 0 0 x4.x13.A1
flabel locali 17581 -76 17615 -42 0 FreeSans 250 0 0 0 x4.x13.A0
flabel locali 17949 -212 17983 -178 0 FreeSans 250 0 0 0 x4.x13.X
flabel locali 17949 60 17983 94 0 FreeSans 250 0 0 0 x4.x13.X
flabel locali 17949 128 17983 162 0 FreeSans 250 0 0 0 x4.x13.X
flabel nwell 17905 230 17939 264 0 FreeSans 250 0 0 0 x4.x13.VPB
flabel pwell 17895 -314 17929 -280 0 FreeSans 250 0 0 0 x4.x13.VNB
rlabel comment 18013 -297 18013 -297 6 x4.x13.mux2_1
rlabel metal1 17185 -345 18013 -249 1 x4.x13.VGND
rlabel metal1 17185 199 18013 295 1 x4.x13.VPWR
flabel metal1 15781 -314 15815 -280 0 FreeSans 200 0 0 0 x4.x12.VGND
flabel metal1 15781 230 15815 264 0 FreeSans 200 0 0 0 x4.x12.VPWR
flabel locali 16425 -8 16459 26 0 FreeSans 250 0 0 0 x4.x12.S
flabel locali 16333 -8 16367 26 0 FreeSans 250 0 0 0 x4.x12.S
flabel locali 16241 -144 16275 -110 0 FreeSans 250 0 0 0 x4.x12.A1
flabel locali 16241 -76 16275 -42 0 FreeSans 250 0 0 0 x4.x12.A1
flabel locali 16149 -76 16183 -42 0 FreeSans 250 0 0 0 x4.x12.A0
flabel locali 15781 -212 15815 -178 0 FreeSans 250 0 0 0 x4.x12.X
flabel locali 15781 60 15815 94 0 FreeSans 250 0 0 0 x4.x12.X
flabel locali 15781 128 15815 162 0 FreeSans 250 0 0 0 x4.x12.X
flabel nwell 15825 230 15859 264 0 FreeSans 250 0 0 0 x4.x12.VPB
flabel pwell 15835 -314 15869 -280 0 FreeSans 250 0 0 0 x4.x12.VNB
rlabel comment 15751 -297 15751 -297 4 x4.x12.mux2_1
rlabel metal1 15751 -345 16579 -249 1 x4.x12.VGND
rlabel metal1 15751 199 16579 295 1 x4.x12.VPWR
flabel metal1 15555 -314 15589 -280 0 FreeSans 200 0 0 0 x4.x11.VGND
flabel metal1 15555 230 15589 264 0 FreeSans 200 0 0 0 x4.x11.VPWR
flabel locali 14911 -8 14945 26 0 FreeSans 250 0 0 0 x4.x11.S
flabel locali 15003 -8 15037 26 0 FreeSans 250 0 0 0 x4.x11.S
flabel locali 15095 -144 15129 -110 0 FreeSans 250 0 0 0 x4.x11.A1
flabel locali 15095 -76 15129 -42 0 FreeSans 250 0 0 0 x4.x11.A1
flabel locali 15187 -76 15221 -42 0 FreeSans 250 0 0 0 x4.x11.A0
flabel locali 15555 -212 15589 -178 0 FreeSans 250 0 0 0 x4.x11.X
flabel locali 15555 60 15589 94 0 FreeSans 250 0 0 0 x4.x11.X
flabel locali 15555 128 15589 162 0 FreeSans 250 0 0 0 x4.x11.X
flabel nwell 15511 230 15545 264 0 FreeSans 250 0 0 0 x4.x11.VPB
flabel pwell 15501 -314 15535 -280 0 FreeSans 250 0 0 0 x4.x11.VNB
rlabel comment 15619 -297 15619 -297 6 x4.x11.mux2_1
rlabel metal1 14791 -345 15619 -249 1 x4.x11.VGND
rlabel metal1 14791 199 15619 295 1 x4.x11.VPWR
flabel metal1 13389 -314 13423 -280 0 FreeSans 200 0 0 0 x4.x10.VGND
flabel metal1 13389 230 13423 264 0 FreeSans 200 0 0 0 x4.x10.VPWR
flabel locali 14033 -8 14067 26 0 FreeSans 250 0 0 0 x4.x10.S
flabel locali 13941 -8 13975 26 0 FreeSans 250 0 0 0 x4.x10.S
flabel locali 13849 -144 13883 -110 0 FreeSans 250 0 0 0 x4.x10.A1
flabel locali 13849 -76 13883 -42 0 FreeSans 250 0 0 0 x4.x10.A1
flabel locali 13757 -76 13791 -42 0 FreeSans 250 0 0 0 x4.x10.A0
flabel locali 13389 -212 13423 -178 0 FreeSans 250 0 0 0 x4.x10.X
flabel locali 13389 60 13423 94 0 FreeSans 250 0 0 0 x4.x10.X
flabel locali 13389 128 13423 162 0 FreeSans 250 0 0 0 x4.x10.X
flabel nwell 13433 230 13467 264 0 FreeSans 250 0 0 0 x4.x10.VPB
flabel pwell 13443 -314 13477 -280 0 FreeSans 250 0 0 0 x4.x10.VNB
rlabel comment 13359 -297 13359 -297 4 x4.x10.mux2_1
rlabel metal1 13359 -345 14187 -249 1 x4.x10.VGND
rlabel metal1 13359 199 14187 295 1 x4.x10.VPWR
flabel metal1 13165 -314 13199 -280 0 FreeSans 200 0 0 0 x4.x9.VGND
flabel metal1 13165 230 13199 264 0 FreeSans 200 0 0 0 x4.x9.VPWR
flabel locali 12521 -8 12555 26 0 FreeSans 250 0 0 0 x4.x9.S
flabel locali 12613 -8 12647 26 0 FreeSans 250 0 0 0 x4.x9.S
flabel locali 12705 -144 12739 -110 0 FreeSans 250 0 0 0 x4.x9.A1
flabel locali 12705 -76 12739 -42 0 FreeSans 250 0 0 0 x4.x9.A1
flabel locali 12797 -76 12831 -42 0 FreeSans 250 0 0 0 x4.x9.A0
flabel locali 13165 -212 13199 -178 0 FreeSans 250 0 0 0 x4.x9.X
flabel locali 13165 60 13199 94 0 FreeSans 250 0 0 0 x4.x9.X
flabel locali 13165 128 13199 162 0 FreeSans 250 0 0 0 x4.x9.X
flabel nwell 13121 230 13155 264 0 FreeSans 250 0 0 0 x4.x9.VPB
flabel pwell 13111 -314 13145 -280 0 FreeSans 250 0 0 0 x4.x9.VNB
rlabel comment 13229 -297 13229 -297 6 x4.x9.mux2_1
rlabel metal1 12401 -345 13229 -249 1 x4.x9.VGND
rlabel metal1 12401 199 13229 295 1 x4.x9.VPWR
flabel metal1 10997 -314 11031 -280 0 FreeSans 200 0 0 0 x4.x8.VGND
flabel metal1 10997 230 11031 264 0 FreeSans 200 0 0 0 x4.x8.VPWR
flabel locali 11641 -8 11675 26 0 FreeSans 250 0 0 0 x4.x8.S
flabel locali 11549 -8 11583 26 0 FreeSans 250 0 0 0 x4.x8.S
flabel locali 11457 -144 11491 -110 0 FreeSans 250 0 0 0 x4.x8.A1
flabel locali 11457 -76 11491 -42 0 FreeSans 250 0 0 0 x4.x8.A1
flabel locali 11365 -76 11399 -42 0 FreeSans 250 0 0 0 x4.x8.A0
flabel locali 10997 -212 11031 -178 0 FreeSans 250 0 0 0 x4.x8.X
flabel locali 10997 60 11031 94 0 FreeSans 250 0 0 0 x4.x8.X
flabel locali 10997 128 11031 162 0 FreeSans 250 0 0 0 x4.x8.X
flabel nwell 11041 230 11075 264 0 FreeSans 250 0 0 0 x4.x8.VPB
flabel pwell 11051 -314 11085 -280 0 FreeSans 250 0 0 0 x4.x8.VNB
rlabel comment 10967 -297 10967 -297 4 x4.x8.mux2_1
rlabel metal1 10967 -345 11795 -249 1 x4.x8.VGND
rlabel metal1 10967 199 11795 295 1 x4.x8.VPWR
flabel metal1 10773 -314 10807 -280 0 FreeSans 200 0 0 0 x4.x7.VGND
flabel metal1 10773 230 10807 264 0 FreeSans 200 0 0 0 x4.x7.VPWR
flabel locali 10129 -8 10163 26 0 FreeSans 250 0 0 0 x4.x7.S
flabel locali 10221 -8 10255 26 0 FreeSans 250 0 0 0 x4.x7.S
flabel locali 10313 -144 10347 -110 0 FreeSans 250 0 0 0 x4.x7.A1
flabel locali 10313 -76 10347 -42 0 FreeSans 250 0 0 0 x4.x7.A1
flabel locali 10405 -76 10439 -42 0 FreeSans 250 0 0 0 x4.x7.A0
flabel locali 10773 -212 10807 -178 0 FreeSans 250 0 0 0 x4.x7.X
flabel locali 10773 60 10807 94 0 FreeSans 250 0 0 0 x4.x7.X
flabel locali 10773 128 10807 162 0 FreeSans 250 0 0 0 x4.x7.X
flabel nwell 10729 230 10763 264 0 FreeSans 250 0 0 0 x4.x7.VPB
flabel pwell 10719 -314 10753 -280 0 FreeSans 250 0 0 0 x4.x7.VNB
rlabel comment 10837 -297 10837 -297 6 x4.x7.mux2_1
rlabel metal1 10009 -345 10837 -249 1 x4.x7.VGND
rlabel metal1 10009 199 10837 295 1 x4.x7.VPWR
flabel metal1 8605 -314 8639 -280 0 FreeSans 200 0 0 0 x4.x6.VGND
flabel metal1 8605 230 8639 264 0 FreeSans 200 0 0 0 x4.x6.VPWR
flabel locali 9249 -8 9283 26 0 FreeSans 250 0 0 0 x4.x6.S
flabel locali 9157 -8 9191 26 0 FreeSans 250 0 0 0 x4.x6.S
flabel locali 9065 -144 9099 -110 0 FreeSans 250 0 0 0 x4.x6.A1
flabel locali 9065 -76 9099 -42 0 FreeSans 250 0 0 0 x4.x6.A1
flabel locali 8973 -76 9007 -42 0 FreeSans 250 0 0 0 x4.x6.A0
flabel locali 8605 -212 8639 -178 0 FreeSans 250 0 0 0 x4.x6.X
flabel locali 8605 60 8639 94 0 FreeSans 250 0 0 0 x4.x6.X
flabel locali 8605 128 8639 162 0 FreeSans 250 0 0 0 x4.x6.X
flabel nwell 8649 230 8683 264 0 FreeSans 250 0 0 0 x4.x6.VPB
flabel pwell 8659 -314 8693 -280 0 FreeSans 250 0 0 0 x4.x6.VNB
rlabel comment 8575 -297 8575 -297 4 x4.x6.mux2_1
rlabel metal1 8575 -345 9403 -249 1 x4.x6.VGND
rlabel metal1 8575 199 9403 295 1 x4.x6.VPWR
flabel locali 9064 -1453 9098 -1419 0 FreeSans 400 0 0 0 x4.x5.RESET_B
flabel locali 10904 -1691 10938 -1657 7 FreeSans 400 0 0 0 x4.x5.VGND
flabel locali 10904 -1453 10938 -1419 0 FreeSans 400 0 0 0 x4.x5.CLK_N
flabel locali 10904 -1385 10938 -1351 0 FreeSans 400 0 0 0 x4.x5.CLK_N
flabel locali 10168 -1521 10202 -1487 0 FreeSans 400 0 0 0 x4.x5.SET_B
flabel locali 8604 -1589 8638 -1555 0 FreeSans 400 0 0 0 x4.x5.Q
flabel locali 8604 -1317 8638 -1283 0 FreeSans 400 0 0 0 x4.x5.Q
flabel locali 8604 -1249 8638 -1215 0 FreeSans 400 0 0 0 x4.x5.Q
flabel locali 10904 -1147 10938 -1113 7 FreeSans 400 0 0 0 x4.x5.VPWR
flabel locali 10536 -1453 10570 -1419 0 FreeSans 200 0 0 0 x4.x5.D
flabel locali 10536 -1385 10570 -1351 0 FreeSans 200 0 0 0 x4.x5.D
flabel locali 8880 -1249 8914 -1215 0 FreeSans 400 0 0 0 x4.x5.Q_N
flabel locali 8880 -1317 8914 -1283 0 FreeSans 400 0 0 0 x4.x5.Q_N
flabel locali 8880 -1589 8914 -1555 0 FreeSans 400 0 0 0 x4.x5.Q_N
flabel metal1 10904 -1691 10938 -1657 0 FreeSans 200 0 0 0 x4.x5.VGND
flabel metal1 10904 -1147 10938 -1113 0 FreeSans 200 0 0 0 x4.x5.VPWR
flabel nwell 10904 -1147 10938 -1113 7 FreeSans 400 0 0 0 x4.x5.VPB
flabel nwell 10921 -1130 10921 -1130 0 FreeSans 200 0 0 0 x4.x5.VPB
flabel pwell 10904 -1691 10938 -1657 7 FreeSans 400 0 0 0 x4.x5.VNB
flabel pwell 10921 -1674 10921 -1674 0 FreeSans 200 0 0 0 x4.x5.VNB
rlabel comment 10967 -1674 10967 -1674 6 x4.x5.dfbbn_1
rlabel locali 9402 -1527 9511 -1461 1 x4.x5.SET_B
rlabel metal1 9406 -1490 9464 -1481 1 x4.x5.SET_B
rlabel metal1 9406 -1527 9464 -1518 1 x4.x5.SET_B
rlabel metal1 10156 -1490 10214 -1481 1 x4.x5.SET_B
rlabel metal1 9406 -1518 10214 -1490 1 x4.x5.SET_B
rlabel metal1 10156 -1527 10214 -1518 1 x4.x5.SET_B
rlabel metal1 8575 -1722 10967 -1626 1 x4.x5.VGND
rlabel metal1 8575 -1178 10967 -1082 1 x4.x5.VPWR
flabel metal1 8883 1372 8917 1406 0 FreeSans 200 0 0 0 x4.x3.VPWR
flabel metal1 8883 828 8917 862 0 FreeSans 200 0 0 0 x4.x3.VGND
flabel locali 9159 1066 9193 1100 0 FreeSans 200 0 0 0 x4.x3.X
flabel locali 9159 1134 9193 1168 0 FreeSans 200 0 0 0 x4.x3.X
flabel locali 9159 998 9193 1032 0 FreeSans 200 0 0 0 x4.x3.X
flabel locali 8883 1372 8917 1406 0 FreeSans 200 0 0 0 x4.x3.VPWR
flabel locali 8883 828 8917 862 0 FreeSans 200 0 0 0 x4.x3.VGND
flabel locali 8883 1066 8917 1100 0 FreeSans 200 0 0 0 x4.x3.A
flabel nwell 8883 1372 8917 1406 0 FreeSans 200 0 0 0 x4.x3.VPB
flabel pwell 8883 828 8917 862 0 FreeSans 200 0 0 0 x4.x3.VNB
rlabel comment 8853 845 8853 845 4 x4.x3.buf_4
rlabel metal1 8853 797 9405 893 1 x4.x3.VGND
rlabel metal1 8853 1341 9405 1437 1 x4.x3.VPWR
flabel locali 9803 1066 9837 1100 0 FreeSans 200 0 0 0 x4.x2.A
flabel locali 9711 1066 9745 1100 0 FreeSans 200 0 0 0 x4.x2.A
flabel locali 11366 1066 11400 1100 0 FreeSans 200 0 0 0 x4.x2.X
flabel locali 11366 1134 11400 1168 0 FreeSans 200 0 0 0 x4.x2.X
flabel pwell 9435 828 9469 862 0 FreeSans 200 0 0 0 x4.x2.VNB
flabel nwell 9435 1372 9469 1406 0 FreeSans 200 0 0 0 x4.x2.VPB
flabel metal1 9435 828 9469 862 0 FreeSans 200 0 0 0 x4.x2.VGND
flabel metal1 9435 1372 9469 1406 0 FreeSans 200 0 0 0 x4.x2.VPWR
rlabel comment 9405 845 9405 845 4 x4.x2.buf_16
rlabel metal1 9405 797 11429 893 1 x4.x2.VGND
rlabel metal1 9405 1341 11429 1437 1 x4.x2.VPWR
flabel metal1 8608 828 8642 862 0 FreeSans 200 0 0 0 x4.x1.VGND
flabel metal1 8606 1372 8640 1406 0 FreeSans 200 0 0 0 x4.x1.VPWR
flabel locali 8606 1372 8640 1406 0 FreeSans 200 0 0 0 x4.x1.VPWR
flabel locali 8608 828 8642 862 0 FreeSans 200 0 0 0 x4.x1.VGND
flabel locali 8788 930 8822 964 0 FreeSans 200 0 0 0 x4.x1.X
flabel locali 8788 1202 8822 1236 0 FreeSans 200 0 0 0 x4.x1.X
flabel locali 8788 1270 8822 1304 0 FreeSans 200 0 0 0 x4.x1.X
flabel locali 8606 1066 8640 1100 0 FreeSans 200 0 0 0 x4.x1.A
flabel nwell 8606 1372 8640 1406 0 FreeSans 200 0 0 0 x4.x1.VPB
flabel pwell 8608 828 8642 862 0 FreeSans 200 0 0 0 x4.x1.VNB
rlabel comment 8577 845 8577 845 4 x4.x1.buf_1
rlabel metal1 8577 797 8853 893 1 x4.x1.VGND
rlabel metal1 8577 1341 8853 1437 1 x4.x1.VPWR
flabel locali 10444 -764 10478 -730 0 FreeSans 400 0 0 0 x4.sky130_fd_sc_hd__dfbbn_1_0.RESET_B
flabel locali 8604 -1002 8638 -968 3 FreeSans 400 0 0 0 x4.sky130_fd_sc_hd__dfbbn_1_0.VGND
flabel locali 8604 -764 8638 -730 0 FreeSans 400 0 0 0 x4.sky130_fd_sc_hd__dfbbn_1_0.CLK_N
flabel locali 8604 -696 8638 -662 0 FreeSans 400 0 0 0 x4.sky130_fd_sc_hd__dfbbn_1_0.CLK_N
flabel locali 9340 -832 9374 -798 0 FreeSans 400 0 0 0 x4.sky130_fd_sc_hd__dfbbn_1_0.SET_B
flabel locali 10904 -900 10938 -866 0 FreeSans 400 0 0 0 x4.sky130_fd_sc_hd__dfbbn_1_0.Q
flabel locali 10904 -628 10938 -594 0 FreeSans 400 0 0 0 x4.sky130_fd_sc_hd__dfbbn_1_0.Q
flabel locali 10904 -560 10938 -526 0 FreeSans 400 0 0 0 x4.sky130_fd_sc_hd__dfbbn_1_0.Q
flabel locali 8604 -458 8638 -424 3 FreeSans 400 0 0 0 x4.sky130_fd_sc_hd__dfbbn_1_0.VPWR
flabel locali 8972 -764 9006 -730 0 FreeSans 200 0 0 0 x4.sky130_fd_sc_hd__dfbbn_1_0.D
flabel locali 8972 -696 9006 -662 0 FreeSans 200 0 0 0 x4.sky130_fd_sc_hd__dfbbn_1_0.D
flabel locali 10628 -560 10662 -526 0 FreeSans 400 0 0 0 x4.sky130_fd_sc_hd__dfbbn_1_0.Q_N
flabel locali 10628 -628 10662 -594 0 FreeSans 400 0 0 0 x4.sky130_fd_sc_hd__dfbbn_1_0.Q_N
flabel locali 10628 -900 10662 -866 0 FreeSans 400 0 0 0 x4.sky130_fd_sc_hd__dfbbn_1_0.Q_N
flabel metal1 8604 -1002 8638 -968 0 FreeSans 200 0 0 0 x4.sky130_fd_sc_hd__dfbbn_1_0.VGND
flabel metal1 8604 -458 8638 -424 0 FreeSans 200 0 0 0 x4.sky130_fd_sc_hd__dfbbn_1_0.VPWR
flabel nwell 8604 -458 8638 -424 3 FreeSans 400 0 0 0 x4.sky130_fd_sc_hd__dfbbn_1_0.VPB
flabel nwell 8621 -441 8621 -441 0 FreeSans 200 0 0 0 x4.sky130_fd_sc_hd__dfbbn_1_0.VPB
flabel pwell 8604 -1002 8638 -968 3 FreeSans 400 0 0 0 x4.sky130_fd_sc_hd__dfbbn_1_0.VNB
flabel pwell 8621 -985 8621 -985 0 FreeSans 200 0 0 0 x4.sky130_fd_sc_hd__dfbbn_1_0.VNB
rlabel comment 8575 -985 8575 -985 4 x4.sky130_fd_sc_hd__dfbbn_1_0.dfbbn_1
rlabel locali 10031 -838 10140 -772 1 x4.sky130_fd_sc_hd__dfbbn_1_0.SET_B
rlabel metal1 10078 -801 10136 -792 1 x4.sky130_fd_sc_hd__dfbbn_1_0.SET_B
rlabel metal1 10078 -838 10136 -829 1 x4.sky130_fd_sc_hd__dfbbn_1_0.SET_B
rlabel metal1 9328 -801 9386 -792 1 x4.sky130_fd_sc_hd__dfbbn_1_0.SET_B
rlabel metal1 9328 -829 10136 -801 1 x4.sky130_fd_sc_hd__dfbbn_1_0.SET_B
rlabel metal1 9328 -838 9386 -829 1 x4.sky130_fd_sc_hd__dfbbn_1_0.SET_B
rlabel metal1 8575 -1033 10967 -937 1 x4.sky130_fd_sc_hd__dfbbn_1_0.VGND
rlabel metal1 8575 -489 10967 -393 1 x4.sky130_fd_sc_hd__dfbbn_1_0.VPWR
flabel metal2 11521 2656 11555 2690 0 FreeSans 480 0 0 0 x3.D[7]
flabel metal2 13913 2656 13947 2690 0 FreeSans 480 0 0 0 x3.D[6]
flabel metal2 16307 2654 16341 2688 0 FreeSans 480 0 0 0 x3.D[5]
flabel metal2 18445 2656 18479 2690 0 FreeSans 480 0 0 0 x3.check[5]
flabel metal2 18869 2651 18903 2685 0 FreeSans 480 0 0 0 x3.check[1]
flabel metal2 20845 2651 20879 2685 0 FreeSans 480 0 0 0 x3.check[4]
flabel metal2 21258 2654 21292 2688 0 FreeSans 480 0 0 0 x3.check[2]
flabel metal2 23239 2651 23273 2685 0 FreeSans 480 0 0 0 x3.check[3]
flabel metal2 21090 2742 21124 2776 0 FreeSans 480 0 0 0 x3.D[3]
flabel metal2 21007 2742 21041 2776 0 FreeSans 480 0 0 0 x3.D[1]
flabel metal2 16049 2654 16083 2688 0 FreeSans 480 0 0 0 x3.check[6]
flabel metal2 18701 2716 18735 2750 0 FreeSans 480 0 0 0 x3.D[4]
flabel metal2 18614 2770 18648 2804 0 FreeSans 480 0 0 0 x3.D[0]
flabel metal2 23395 2726 23429 2760 0 FreeSans 480 0 0 0 x3.D[2]
flabel metal2 16449 2651 16483 2685 0 FreeSans 480 0 0 0 x3.check[0]
flabel metal1 10933 5194 10967 5228 0 FreeSans 480 0 0 0 x3.reset
flabel metal1 10931 4320 10965 4354 0 FreeSans 480 0 0 0 x3.eob
flabel metal1 10933 3943 10967 3977 0 FreeSans 480 0 0 0 x3.comparator_out
flabel metal1 10925 6754 10959 6788 0 FreeSans 480 0 0 0 x3.clk_sar
flabel metal1 10927 6688 10961 6722 0 FreeSans 480 0 0 0 x3.sel_bit[1]
flabel metal1 10922 6824 10956 6858 0 FreeSans 480 0 0 0 x3.sel_bit[0]
flabel metal4 23357 6466 23907 7108 0 FreeSans 320 0 0 0 x3.VSS
flabel metal4 10753 6132 14359 6918 0 FreeSans 320 0 0 0 x3.VDD
flabel locali 13795 4387 13829 4421 0 FreeSans 340 0 0 0 x3.x77.Y
flabel locali 13795 4319 13829 4353 0 FreeSans 340 0 0 0 x3.x77.Y
flabel locali 13703 4319 13737 4353 0 FreeSans 340 0 0 0 x3.x77.A
flabel metal1 13660 4081 13694 4115 0 FreeSans 200 0 0 0 x3.x77.VGND
flabel metal1 13660 4625 13694 4659 0 FreeSans 200 0 0 0 x3.x77.VPWR
rlabel comment 13631 4098 13631 4098 4 x3.x77.inv_1
rlabel metal1 13631 4050 13907 4146 1 x3.x77.VGND
rlabel metal1 13631 4594 13907 4690 1 x3.x77.VPWR
flabel pwell 13660 4081 13694 4115 0 FreeSans 200 0 0 0 x3.x77.VNB
flabel nwell 13660 4625 13694 4659 0 FreeSans 200 0 0 0 x3.x77.VPB
flabel locali 15751 4317 15826 4363 0 FreeSans 400 0 0 0 x3.x75.RESET_B
flabel locali 13918 4081 13952 4115 3 FreeSans 400 0 0 0 x3.x75.VGND
flabel locali 13918 4319 13952 4353 0 FreeSans 400 0 0 0 x3.x75.CLK
flabel locali 13918 4387 13952 4421 0 FreeSans 400 0 0 0 x3.x75.CLK
flabel locali 14654 4251 14688 4285 0 FreeSans 400 0 0 0 x3.x75.SET_B
flabel locali 16216 4183 16250 4217 0 FreeSans 400 0 0 0 x3.x75.Q
flabel locali 16216 4455 16250 4489 0 FreeSans 400 0 0 0 x3.x75.Q
flabel locali 16216 4523 16250 4557 0 FreeSans 400 0 0 0 x3.x75.Q
flabel locali 13918 4625 13952 4659 3 FreeSans 400 0 0 0 x3.x75.VPWR
flabel locali 14286 4319 14320 4353 0 FreeSans 200 0 0 0 x3.x75.D
flabel locali 14286 4387 14320 4421 0 FreeSans 200 0 0 0 x3.x75.D
flabel locali 15936 4523 15970 4557 0 FreeSans 400 0 0 0 x3.x75.Q_N
flabel locali 15936 4455 15970 4489 0 FreeSans 400 0 0 0 x3.x75.Q_N
flabel locali 15936 4183 15970 4217 0 FreeSans 400 0 0 0 x3.x75.Q_N
flabel metal1 13918 4081 13952 4115 0 FreeSans 200 0 0 0 x3.x75.VGND
flabel metal1 13918 4625 13952 4659 0 FreeSans 200 0 0 0 x3.x75.VPWR
flabel nwell 13918 4625 13952 4659 3 FreeSans 400 0 0 0 x3.x75.VPB
flabel nwell 13935 4642 13935 4642 0 FreeSans 200 0 0 0 x3.x75.VPB
flabel pwell 13918 4081 13952 4115 3 FreeSans 400 0 0 0 x3.x75.VNB
flabel pwell 13935 4098 13935 4098 0 FreeSans 200 0 0 0 x3.x75.VNB
rlabel comment 13888 4098 13888 4098 4 x3.x75.dfbbp_1
rlabel locali 15380 4245 15455 4311 1 x3.x75.SET_B
rlabel metal1 15378 4282 15436 4291 1 x3.x75.SET_B
rlabel metal1 15378 4245 15436 4254 1 x3.x75.SET_B
rlabel metal1 14642 4282 14700 4291 1 x3.x75.SET_B
rlabel metal1 14642 4254 15436 4282 1 x3.x75.SET_B
rlabel metal1 14642 4245 14700 4254 1 x3.x75.SET_B
rlabel metal1 13888 4050 16280 4146 1 x3.x75.VGND
rlabel metal1 13888 4594 16280 4690 1 x3.x75.VPWR
flabel locali 18143 4317 18218 4363 0 FreeSans 400 0 0 0 x3.x72.RESET_B
flabel locali 16310 4081 16344 4115 3 FreeSans 400 0 0 0 x3.x72.VGND
flabel locali 16310 4319 16344 4353 0 FreeSans 400 0 0 0 x3.x72.CLK
flabel locali 16310 4387 16344 4421 0 FreeSans 400 0 0 0 x3.x72.CLK
flabel locali 17046 4251 17080 4285 0 FreeSans 400 0 0 0 x3.x72.SET_B
flabel locali 18608 4183 18642 4217 0 FreeSans 400 0 0 0 x3.x72.Q
flabel locali 18608 4455 18642 4489 0 FreeSans 400 0 0 0 x3.x72.Q
flabel locali 18608 4523 18642 4557 0 FreeSans 400 0 0 0 x3.x72.Q
flabel locali 16310 4625 16344 4659 3 FreeSans 400 0 0 0 x3.x72.VPWR
flabel locali 16678 4319 16712 4353 0 FreeSans 200 0 0 0 x3.x72.D
flabel locali 16678 4387 16712 4421 0 FreeSans 200 0 0 0 x3.x72.D
flabel locali 18328 4523 18362 4557 0 FreeSans 400 0 0 0 x3.x72.Q_N
flabel locali 18328 4455 18362 4489 0 FreeSans 400 0 0 0 x3.x72.Q_N
flabel locali 18328 4183 18362 4217 0 FreeSans 400 0 0 0 x3.x72.Q_N
flabel metal1 16310 4081 16344 4115 0 FreeSans 200 0 0 0 x3.x72.VGND
flabel metal1 16310 4625 16344 4659 0 FreeSans 200 0 0 0 x3.x72.VPWR
flabel nwell 16310 4625 16344 4659 3 FreeSans 400 0 0 0 x3.x72.VPB
flabel nwell 16327 4642 16327 4642 0 FreeSans 200 0 0 0 x3.x72.VPB
flabel pwell 16310 4081 16344 4115 3 FreeSans 400 0 0 0 x3.x72.VNB
flabel pwell 16327 4098 16327 4098 0 FreeSans 200 0 0 0 x3.x72.VNB
rlabel comment 16280 4098 16280 4098 4 x3.x72.dfbbp_1
rlabel locali 17772 4245 17847 4311 1 x3.x72.SET_B
rlabel metal1 17770 4282 17828 4291 1 x3.x72.SET_B
rlabel metal1 17770 4245 17828 4254 1 x3.x72.SET_B
rlabel metal1 17034 4282 17092 4291 1 x3.x72.SET_B
rlabel metal1 17034 4254 17828 4282 1 x3.x72.SET_B
rlabel metal1 17034 4245 17092 4254 1 x3.x72.SET_B
rlabel metal1 16280 4050 18672 4146 1 x3.x72.VGND
rlabel metal1 16280 4594 18672 4690 1 x3.x72.VPWR
flabel locali 20535 4317 20610 4363 0 FreeSans 400 0 0 0 x3.x69.RESET_B
flabel locali 18702 4081 18736 4115 3 FreeSans 400 0 0 0 x3.x69.VGND
flabel locali 18702 4319 18736 4353 0 FreeSans 400 0 0 0 x3.x69.CLK
flabel locali 18702 4387 18736 4421 0 FreeSans 400 0 0 0 x3.x69.CLK
flabel locali 19438 4251 19472 4285 0 FreeSans 400 0 0 0 x3.x69.SET_B
flabel locali 21000 4183 21034 4217 0 FreeSans 400 0 0 0 x3.x69.Q
flabel locali 21000 4455 21034 4489 0 FreeSans 400 0 0 0 x3.x69.Q
flabel locali 21000 4523 21034 4557 0 FreeSans 400 0 0 0 x3.x69.Q
flabel locali 18702 4625 18736 4659 3 FreeSans 400 0 0 0 x3.x69.VPWR
flabel locali 19070 4319 19104 4353 0 FreeSans 200 0 0 0 x3.x69.D
flabel locali 19070 4387 19104 4421 0 FreeSans 200 0 0 0 x3.x69.D
flabel locali 20720 4523 20754 4557 0 FreeSans 400 0 0 0 x3.x69.Q_N
flabel locali 20720 4455 20754 4489 0 FreeSans 400 0 0 0 x3.x69.Q_N
flabel locali 20720 4183 20754 4217 0 FreeSans 400 0 0 0 x3.x69.Q_N
flabel metal1 18702 4081 18736 4115 0 FreeSans 200 0 0 0 x3.x69.VGND
flabel metal1 18702 4625 18736 4659 0 FreeSans 200 0 0 0 x3.x69.VPWR
flabel nwell 18702 4625 18736 4659 3 FreeSans 400 0 0 0 x3.x69.VPB
flabel nwell 18719 4642 18719 4642 0 FreeSans 200 0 0 0 x3.x69.VPB
flabel pwell 18702 4081 18736 4115 3 FreeSans 400 0 0 0 x3.x69.VNB
flabel pwell 18719 4098 18719 4098 0 FreeSans 200 0 0 0 x3.x69.VNB
rlabel comment 18672 4098 18672 4098 4 x3.x69.dfbbp_1
rlabel locali 20164 4245 20239 4311 1 x3.x69.SET_B
rlabel metal1 20162 4282 20220 4291 1 x3.x69.SET_B
rlabel metal1 20162 4245 20220 4254 1 x3.x69.SET_B
rlabel metal1 19426 4282 19484 4291 1 x3.x69.SET_B
rlabel metal1 19426 4254 20220 4282 1 x3.x69.SET_B
rlabel metal1 19426 4245 19484 4254 1 x3.x69.SET_B
rlabel metal1 18672 4050 21064 4146 1 x3.x69.VGND
rlabel metal1 18672 4594 21064 4690 1 x3.x69.VPWR
flabel locali 22927 4317 23002 4363 0 FreeSans 400 0 0 0 x3.x66.RESET_B
flabel locali 21094 4081 21128 4115 3 FreeSans 400 0 0 0 x3.x66.VGND
flabel locali 21094 4319 21128 4353 0 FreeSans 400 0 0 0 x3.x66.CLK
flabel locali 21094 4387 21128 4421 0 FreeSans 400 0 0 0 x3.x66.CLK
flabel locali 21830 4251 21864 4285 0 FreeSans 400 0 0 0 x3.x66.SET_B
flabel locali 23392 4183 23426 4217 0 FreeSans 400 0 0 0 x3.x66.Q
flabel locali 23392 4455 23426 4489 0 FreeSans 400 0 0 0 x3.x66.Q
flabel locali 23392 4523 23426 4557 0 FreeSans 400 0 0 0 x3.x66.Q
flabel locali 21094 4625 21128 4659 3 FreeSans 400 0 0 0 x3.x66.VPWR
flabel locali 21462 4319 21496 4353 0 FreeSans 200 0 0 0 x3.x66.D
flabel locali 21462 4387 21496 4421 0 FreeSans 200 0 0 0 x3.x66.D
flabel locali 23112 4523 23146 4557 0 FreeSans 400 0 0 0 x3.x66.Q_N
flabel locali 23112 4455 23146 4489 0 FreeSans 400 0 0 0 x3.x66.Q_N
flabel locali 23112 4183 23146 4217 0 FreeSans 400 0 0 0 x3.x66.Q_N
flabel metal1 21094 4081 21128 4115 0 FreeSans 200 0 0 0 x3.x66.VGND
flabel metal1 21094 4625 21128 4659 0 FreeSans 200 0 0 0 x3.x66.VPWR
flabel nwell 21094 4625 21128 4659 3 FreeSans 400 0 0 0 x3.x66.VPB
flabel nwell 21111 4642 21111 4642 0 FreeSans 200 0 0 0 x3.x66.VPB
flabel pwell 21094 4081 21128 4115 3 FreeSans 400 0 0 0 x3.x66.VNB
flabel pwell 21111 4098 21111 4098 0 FreeSans 200 0 0 0 x3.x66.VNB
rlabel comment 21064 4098 21064 4098 4 x3.x66.dfbbp_1
rlabel locali 22556 4245 22631 4311 1 x3.x66.SET_B
rlabel metal1 22554 4282 22612 4291 1 x3.x66.SET_B
rlabel metal1 22554 4245 22612 4254 1 x3.x66.SET_B
rlabel metal1 21818 4282 21876 4291 1 x3.x66.SET_B
rlabel metal1 21818 4254 22612 4282 1 x3.x66.SET_B
rlabel metal1 21818 4245 21876 4254 1 x3.x66.SET_B
rlabel metal1 21064 4050 23456 4146 1 x3.x66.VGND
rlabel metal1 21064 4594 23456 4690 1 x3.x66.VPWR
flabel locali 21518 3444 21593 3490 0 FreeSans 400 0 0 0 x3.x63.RESET_B
flabel locali 23392 3208 23426 3242 7 FreeSans 400 0 0 0 x3.x63.VGND
flabel locali 23392 3446 23426 3480 0 FreeSans 400 0 0 0 x3.x63.CLK
flabel locali 23392 3514 23426 3548 0 FreeSans 400 0 0 0 x3.x63.CLK
flabel locali 22656 3378 22690 3412 0 FreeSans 400 0 0 0 x3.x63.SET_B
flabel locali 21094 3310 21128 3344 0 FreeSans 400 0 0 0 x3.x63.Q
flabel locali 21094 3582 21128 3616 0 FreeSans 400 0 0 0 x3.x63.Q
flabel locali 21094 3650 21128 3684 0 FreeSans 400 0 0 0 x3.x63.Q
flabel locali 23392 3752 23426 3786 7 FreeSans 400 0 0 0 x3.x63.VPWR
flabel locali 23024 3446 23058 3480 0 FreeSans 200 0 0 0 x3.x63.D
flabel locali 23024 3514 23058 3548 0 FreeSans 200 0 0 0 x3.x63.D
flabel locali 21374 3650 21408 3684 0 FreeSans 400 0 0 0 x3.x63.Q_N
flabel locali 21374 3582 21408 3616 0 FreeSans 400 0 0 0 x3.x63.Q_N
flabel locali 21374 3310 21408 3344 0 FreeSans 400 0 0 0 x3.x63.Q_N
flabel metal1 23392 3208 23426 3242 0 FreeSans 200 0 0 0 x3.x63.VGND
flabel metal1 23392 3752 23426 3786 0 FreeSans 200 0 0 0 x3.x63.VPWR
flabel nwell 23392 3752 23426 3786 7 FreeSans 400 0 0 0 x3.x63.VPB
flabel nwell 23409 3769 23409 3769 0 FreeSans 200 0 0 0 x3.x63.VPB
flabel pwell 23392 3208 23426 3242 7 FreeSans 400 0 0 0 x3.x63.VNB
flabel pwell 23409 3225 23409 3225 0 FreeSans 200 0 0 0 x3.x63.VNB
rlabel comment 23456 3225 23456 3225 6 x3.x63.dfbbp_1
rlabel locali 21889 3372 21964 3438 1 x3.x63.SET_B
rlabel metal1 21908 3409 21966 3418 1 x3.x63.SET_B
rlabel metal1 21908 3372 21966 3381 1 x3.x63.SET_B
rlabel metal1 22644 3409 22702 3418 1 x3.x63.SET_B
rlabel metal1 21908 3381 22702 3409 1 x3.x63.SET_B
rlabel metal1 22644 3372 22702 3381 1 x3.x63.SET_B
rlabel metal1 21064 3177 23456 3273 1 x3.x63.VGND
rlabel metal1 21064 3721 23456 3817 1 x3.x63.VPWR
flabel locali 19126 3444 19201 3490 0 FreeSans 400 0 0 0 x3.x60.RESET_B
flabel locali 21000 3208 21034 3242 7 FreeSans 400 0 0 0 x3.x60.VGND
flabel locali 21000 3446 21034 3480 0 FreeSans 400 0 0 0 x3.x60.CLK
flabel locali 21000 3514 21034 3548 0 FreeSans 400 0 0 0 x3.x60.CLK
flabel locali 20264 3378 20298 3412 0 FreeSans 400 0 0 0 x3.x60.SET_B
flabel locali 18702 3310 18736 3344 0 FreeSans 400 0 0 0 x3.x60.Q
flabel locali 18702 3582 18736 3616 0 FreeSans 400 0 0 0 x3.x60.Q
flabel locali 18702 3650 18736 3684 0 FreeSans 400 0 0 0 x3.x60.Q
flabel locali 21000 3752 21034 3786 7 FreeSans 400 0 0 0 x3.x60.VPWR
flabel locali 20632 3446 20666 3480 0 FreeSans 200 0 0 0 x3.x60.D
flabel locali 20632 3514 20666 3548 0 FreeSans 200 0 0 0 x3.x60.D
flabel locali 18982 3650 19016 3684 0 FreeSans 400 0 0 0 x3.x60.Q_N
flabel locali 18982 3582 19016 3616 0 FreeSans 400 0 0 0 x3.x60.Q_N
flabel locali 18982 3310 19016 3344 0 FreeSans 400 0 0 0 x3.x60.Q_N
flabel metal1 21000 3208 21034 3242 0 FreeSans 200 0 0 0 x3.x60.VGND
flabel metal1 21000 3752 21034 3786 0 FreeSans 200 0 0 0 x3.x60.VPWR
flabel nwell 21000 3752 21034 3786 7 FreeSans 400 0 0 0 x3.x60.VPB
flabel nwell 21017 3769 21017 3769 0 FreeSans 200 0 0 0 x3.x60.VPB
flabel pwell 21000 3208 21034 3242 7 FreeSans 400 0 0 0 x3.x60.VNB
flabel pwell 21017 3225 21017 3225 0 FreeSans 200 0 0 0 x3.x60.VNB
rlabel comment 21064 3225 21064 3225 6 x3.x60.dfbbp_1
rlabel locali 19497 3372 19572 3438 1 x3.x60.SET_B
rlabel metal1 19516 3409 19574 3418 1 x3.x60.SET_B
rlabel metal1 19516 3372 19574 3381 1 x3.x60.SET_B
rlabel metal1 20252 3409 20310 3418 1 x3.x60.SET_B
rlabel metal1 19516 3381 20310 3409 1 x3.x60.SET_B
rlabel metal1 20252 3372 20310 3381 1 x3.x60.SET_B
rlabel metal1 18672 3177 21064 3273 1 x3.x60.VGND
rlabel metal1 18672 3721 21064 3817 1 x3.x60.VPWR
flabel locali 16734 3444 16809 3490 0 FreeSans 400 0 0 0 x3.x57.RESET_B
flabel locali 18608 3208 18642 3242 7 FreeSans 400 0 0 0 x3.x57.VGND
flabel locali 18608 3446 18642 3480 0 FreeSans 400 0 0 0 x3.x57.CLK
flabel locali 18608 3514 18642 3548 0 FreeSans 400 0 0 0 x3.x57.CLK
flabel locali 17872 3378 17906 3412 0 FreeSans 400 0 0 0 x3.x57.SET_B
flabel locali 16310 3310 16344 3344 0 FreeSans 400 0 0 0 x3.x57.Q
flabel locali 16310 3582 16344 3616 0 FreeSans 400 0 0 0 x3.x57.Q
flabel locali 16310 3650 16344 3684 0 FreeSans 400 0 0 0 x3.x57.Q
flabel locali 18608 3752 18642 3786 7 FreeSans 400 0 0 0 x3.x57.VPWR
flabel locali 18240 3446 18274 3480 0 FreeSans 200 0 0 0 x3.x57.D
flabel locali 18240 3514 18274 3548 0 FreeSans 200 0 0 0 x3.x57.D
flabel locali 16590 3650 16624 3684 0 FreeSans 400 0 0 0 x3.x57.Q_N
flabel locali 16590 3582 16624 3616 0 FreeSans 400 0 0 0 x3.x57.Q_N
flabel locali 16590 3310 16624 3344 0 FreeSans 400 0 0 0 x3.x57.Q_N
flabel metal1 18608 3208 18642 3242 0 FreeSans 200 0 0 0 x3.x57.VGND
flabel metal1 18608 3752 18642 3786 0 FreeSans 200 0 0 0 x3.x57.VPWR
flabel nwell 18608 3752 18642 3786 7 FreeSans 400 0 0 0 x3.x57.VPB
flabel nwell 18625 3769 18625 3769 0 FreeSans 200 0 0 0 x3.x57.VPB
flabel pwell 18608 3208 18642 3242 7 FreeSans 400 0 0 0 x3.x57.VNB
flabel pwell 18625 3225 18625 3225 0 FreeSans 200 0 0 0 x3.x57.VNB
rlabel comment 18672 3225 18672 3225 6 x3.x57.dfbbp_1
rlabel locali 17105 3372 17180 3438 1 x3.x57.SET_B
rlabel metal1 17124 3409 17182 3418 1 x3.x57.SET_B
rlabel metal1 17124 3372 17182 3381 1 x3.x57.SET_B
rlabel metal1 17860 3409 17918 3418 1 x3.x57.SET_B
rlabel metal1 17124 3381 17918 3409 1 x3.x57.SET_B
rlabel metal1 17860 3372 17918 3381 1 x3.x57.SET_B
rlabel metal1 16280 3177 18672 3273 1 x3.x57.VGND
rlabel metal1 16280 3721 18672 3817 1 x3.x57.VPWR
flabel locali 14342 3444 14417 3490 0 FreeSans 400 0 0 0 x3.x54.RESET_B
flabel locali 16216 3208 16250 3242 7 FreeSans 400 0 0 0 x3.x54.VGND
flabel locali 16216 3446 16250 3480 0 FreeSans 400 0 0 0 x3.x54.CLK
flabel locali 16216 3514 16250 3548 0 FreeSans 400 0 0 0 x3.x54.CLK
flabel locali 15480 3378 15514 3412 0 FreeSans 400 0 0 0 x3.x54.SET_B
flabel locali 13918 3310 13952 3344 0 FreeSans 400 0 0 0 x3.x54.Q
flabel locali 13918 3582 13952 3616 0 FreeSans 400 0 0 0 x3.x54.Q
flabel locali 13918 3650 13952 3684 0 FreeSans 400 0 0 0 x3.x54.Q
flabel locali 16216 3752 16250 3786 7 FreeSans 400 0 0 0 x3.x54.VPWR
flabel locali 15848 3446 15882 3480 0 FreeSans 200 0 0 0 x3.x54.D
flabel locali 15848 3514 15882 3548 0 FreeSans 200 0 0 0 x3.x54.D
flabel locali 14198 3650 14232 3684 0 FreeSans 400 0 0 0 x3.x54.Q_N
flabel locali 14198 3582 14232 3616 0 FreeSans 400 0 0 0 x3.x54.Q_N
flabel locali 14198 3310 14232 3344 0 FreeSans 400 0 0 0 x3.x54.Q_N
flabel metal1 16216 3208 16250 3242 0 FreeSans 200 0 0 0 x3.x54.VGND
flabel metal1 16216 3752 16250 3786 0 FreeSans 200 0 0 0 x3.x54.VPWR
flabel nwell 16216 3752 16250 3786 7 FreeSans 400 0 0 0 x3.x54.VPB
flabel nwell 16233 3769 16233 3769 0 FreeSans 200 0 0 0 x3.x54.VPB
flabel pwell 16216 3208 16250 3242 7 FreeSans 400 0 0 0 x3.x54.VNB
flabel pwell 16233 3225 16233 3225 0 FreeSans 200 0 0 0 x3.x54.VNB
rlabel comment 16280 3225 16280 3225 6 x3.x54.dfbbp_1
rlabel locali 14713 3372 14788 3438 1 x3.x54.SET_B
rlabel metal1 14732 3409 14790 3418 1 x3.x54.SET_B
rlabel metal1 14732 3372 14790 3381 1 x3.x54.SET_B
rlabel metal1 15468 3409 15526 3418 1 x3.x54.SET_B
rlabel metal1 14732 3381 15526 3409 1 x3.x54.SET_B
rlabel metal1 15468 3372 15526 3381 1 x3.x54.SET_B
rlabel metal1 13888 3177 16280 3273 1 x3.x54.VGND
rlabel metal1 13888 3721 16280 3817 1 x3.x54.VPWR
flabel locali 11950 3444 12025 3490 0 FreeSans 400 0 0 0 x3.x51.RESET_B
flabel locali 13824 3208 13858 3242 7 FreeSans 400 0 0 0 x3.x51.VGND
flabel locali 13824 3446 13858 3480 0 FreeSans 400 0 0 0 x3.x51.CLK
flabel locali 13824 3514 13858 3548 0 FreeSans 400 0 0 0 x3.x51.CLK
flabel locali 13088 3378 13122 3412 0 FreeSans 400 0 0 0 x3.x51.SET_B
flabel locali 11526 3310 11560 3344 0 FreeSans 400 0 0 0 x3.x51.Q
flabel locali 11526 3582 11560 3616 0 FreeSans 400 0 0 0 x3.x51.Q
flabel locali 11526 3650 11560 3684 0 FreeSans 400 0 0 0 x3.x51.Q
flabel locali 13824 3752 13858 3786 7 FreeSans 400 0 0 0 x3.x51.VPWR
flabel locali 13456 3446 13490 3480 0 FreeSans 200 0 0 0 x3.x51.D
flabel locali 13456 3514 13490 3548 0 FreeSans 200 0 0 0 x3.x51.D
flabel locali 11806 3650 11840 3684 0 FreeSans 400 0 0 0 x3.x51.Q_N
flabel locali 11806 3582 11840 3616 0 FreeSans 400 0 0 0 x3.x51.Q_N
flabel locali 11806 3310 11840 3344 0 FreeSans 400 0 0 0 x3.x51.Q_N
flabel metal1 13824 3208 13858 3242 0 FreeSans 200 0 0 0 x3.x51.VGND
flabel metal1 13824 3752 13858 3786 0 FreeSans 200 0 0 0 x3.x51.VPWR
flabel nwell 13824 3752 13858 3786 7 FreeSans 400 0 0 0 x3.x51.VPB
flabel nwell 13841 3769 13841 3769 0 FreeSans 200 0 0 0 x3.x51.VPB
flabel pwell 13824 3208 13858 3242 7 FreeSans 400 0 0 0 x3.x51.VNB
flabel pwell 13841 3225 13841 3225 0 FreeSans 200 0 0 0 x3.x51.VNB
rlabel comment 13888 3225 13888 3225 6 x3.x51.dfbbp_1
rlabel locali 12321 3372 12396 3438 1 x3.x51.SET_B
rlabel metal1 12340 3409 12398 3418 1 x3.x51.SET_B
rlabel metal1 12340 3372 12398 3381 1 x3.x51.SET_B
rlabel metal1 13076 3409 13134 3418 1 x3.x51.SET_B
rlabel metal1 12340 3381 13134 3409 1 x3.x51.SET_B
rlabel metal1 13076 3372 13134 3381 1 x3.x51.SET_B
rlabel metal1 11496 3177 13888 3273 1 x3.x51.VGND
rlabel metal1 11496 3721 13888 3817 1 x3.x51.VPWR
flabel locali 14343 5190 14418 5236 0 FreeSans 400 0 0 0 x3.x48.RESET_B
flabel locali 16217 4954 16251 4988 7 FreeSans 400 0 0 0 x3.x48.VGND
flabel locali 16217 5192 16251 5226 0 FreeSans 400 0 0 0 x3.x48.CLK
flabel locali 16217 5260 16251 5294 0 FreeSans 400 0 0 0 x3.x48.CLK
flabel locali 15481 5124 15515 5158 0 FreeSans 400 0 0 0 x3.x48.SET_B
flabel locali 13919 5056 13953 5090 0 FreeSans 400 0 0 0 x3.x48.Q
flabel locali 13919 5328 13953 5362 0 FreeSans 400 0 0 0 x3.x48.Q
flabel locali 13919 5396 13953 5430 0 FreeSans 400 0 0 0 x3.x48.Q
flabel locali 16217 5498 16251 5532 7 FreeSans 400 0 0 0 x3.x48.VPWR
flabel locali 15849 5192 15883 5226 0 FreeSans 200 0 0 0 x3.x48.D
flabel locali 15849 5260 15883 5294 0 FreeSans 200 0 0 0 x3.x48.D
flabel locali 14199 5396 14233 5430 0 FreeSans 400 0 0 0 x3.x48.Q_N
flabel locali 14199 5328 14233 5362 0 FreeSans 400 0 0 0 x3.x48.Q_N
flabel locali 14199 5056 14233 5090 0 FreeSans 400 0 0 0 x3.x48.Q_N
flabel metal1 16217 4954 16251 4988 0 FreeSans 200 0 0 0 x3.x48.VGND
flabel metal1 16217 5498 16251 5532 0 FreeSans 200 0 0 0 x3.x48.VPWR
flabel nwell 16217 5498 16251 5532 7 FreeSans 400 0 0 0 x3.x48.VPB
flabel nwell 16234 5515 16234 5515 0 FreeSans 200 0 0 0 x3.x48.VPB
flabel pwell 16217 4954 16251 4988 7 FreeSans 400 0 0 0 x3.x48.VNB
flabel pwell 16234 4971 16234 4971 0 FreeSans 200 0 0 0 x3.x48.VNB
rlabel comment 16281 4971 16281 4971 6 x3.x48.dfbbp_1
rlabel locali 14714 5118 14789 5184 1 x3.x48.SET_B
rlabel metal1 14733 5155 14791 5164 1 x3.x48.SET_B
rlabel metal1 14733 5118 14791 5127 1 x3.x48.SET_B
rlabel metal1 15469 5155 15527 5164 1 x3.x48.SET_B
rlabel metal1 14733 5127 15527 5155 1 x3.x48.SET_B
rlabel metal1 15469 5118 15527 5127 1 x3.x48.SET_B
rlabel metal1 13889 4923 16281 5019 1 x3.x48.VGND
rlabel metal1 13889 5467 16281 5563 1 x3.x48.VPWR
flabel locali 16735 5190 16810 5236 0 FreeSans 400 0 0 0 x3.x45.RESET_B
flabel locali 18609 4954 18643 4988 7 FreeSans 400 0 0 0 x3.x45.VGND
flabel locali 18609 5192 18643 5226 0 FreeSans 400 0 0 0 x3.x45.CLK
flabel locali 18609 5260 18643 5294 0 FreeSans 400 0 0 0 x3.x45.CLK
flabel locali 17873 5124 17907 5158 0 FreeSans 400 0 0 0 x3.x45.SET_B
flabel locali 16311 5056 16345 5090 0 FreeSans 400 0 0 0 x3.x45.Q
flabel locali 16311 5328 16345 5362 0 FreeSans 400 0 0 0 x3.x45.Q
flabel locali 16311 5396 16345 5430 0 FreeSans 400 0 0 0 x3.x45.Q
flabel locali 18609 5498 18643 5532 7 FreeSans 400 0 0 0 x3.x45.VPWR
flabel locali 18241 5192 18275 5226 0 FreeSans 200 0 0 0 x3.x45.D
flabel locali 18241 5260 18275 5294 0 FreeSans 200 0 0 0 x3.x45.D
flabel locali 16591 5396 16625 5430 0 FreeSans 400 0 0 0 x3.x45.Q_N
flabel locali 16591 5328 16625 5362 0 FreeSans 400 0 0 0 x3.x45.Q_N
flabel locali 16591 5056 16625 5090 0 FreeSans 400 0 0 0 x3.x45.Q_N
flabel metal1 18609 4954 18643 4988 0 FreeSans 200 0 0 0 x3.x45.VGND
flabel metal1 18609 5498 18643 5532 0 FreeSans 200 0 0 0 x3.x45.VPWR
flabel nwell 18609 5498 18643 5532 7 FreeSans 400 0 0 0 x3.x45.VPB
flabel nwell 18626 5515 18626 5515 0 FreeSans 200 0 0 0 x3.x45.VPB
flabel pwell 18609 4954 18643 4988 7 FreeSans 400 0 0 0 x3.x45.VNB
flabel pwell 18626 4971 18626 4971 0 FreeSans 200 0 0 0 x3.x45.VNB
rlabel comment 18673 4971 18673 4971 6 x3.x45.dfbbp_1
rlabel locali 17106 5118 17181 5184 1 x3.x45.SET_B
rlabel metal1 17125 5155 17183 5164 1 x3.x45.SET_B
rlabel metal1 17125 5118 17183 5127 1 x3.x45.SET_B
rlabel metal1 17861 5155 17919 5164 1 x3.x45.SET_B
rlabel metal1 17125 5127 17919 5155 1 x3.x45.SET_B
rlabel metal1 17861 5118 17919 5127 1 x3.x45.SET_B
rlabel metal1 16281 4923 18673 5019 1 x3.x45.VGND
rlabel metal1 16281 5467 18673 5563 1 x3.x45.VPWR
flabel locali 19127 5190 19202 5236 0 FreeSans 400 0 0 0 x3.x42.RESET_B
flabel locali 21001 4954 21035 4988 7 FreeSans 400 0 0 0 x3.x42.VGND
flabel locali 21001 5192 21035 5226 0 FreeSans 400 0 0 0 x3.x42.CLK
flabel locali 21001 5260 21035 5294 0 FreeSans 400 0 0 0 x3.x42.CLK
flabel locali 20265 5124 20299 5158 0 FreeSans 400 0 0 0 x3.x42.SET_B
flabel locali 18703 5056 18737 5090 0 FreeSans 400 0 0 0 x3.x42.Q
flabel locali 18703 5328 18737 5362 0 FreeSans 400 0 0 0 x3.x42.Q
flabel locali 18703 5396 18737 5430 0 FreeSans 400 0 0 0 x3.x42.Q
flabel locali 21001 5498 21035 5532 7 FreeSans 400 0 0 0 x3.x42.VPWR
flabel locali 20633 5192 20667 5226 0 FreeSans 200 0 0 0 x3.x42.D
flabel locali 20633 5260 20667 5294 0 FreeSans 200 0 0 0 x3.x42.D
flabel locali 18983 5396 19017 5430 0 FreeSans 400 0 0 0 x3.x42.Q_N
flabel locali 18983 5328 19017 5362 0 FreeSans 400 0 0 0 x3.x42.Q_N
flabel locali 18983 5056 19017 5090 0 FreeSans 400 0 0 0 x3.x42.Q_N
flabel metal1 21001 4954 21035 4988 0 FreeSans 200 0 0 0 x3.x42.VGND
flabel metal1 21001 5498 21035 5532 0 FreeSans 200 0 0 0 x3.x42.VPWR
flabel nwell 21001 5498 21035 5532 7 FreeSans 400 0 0 0 x3.x42.VPB
flabel nwell 21018 5515 21018 5515 0 FreeSans 200 0 0 0 x3.x42.VPB
flabel pwell 21001 4954 21035 4988 7 FreeSans 400 0 0 0 x3.x42.VNB
flabel pwell 21018 4971 21018 4971 0 FreeSans 200 0 0 0 x3.x42.VNB
rlabel comment 21065 4971 21065 4971 6 x3.x42.dfbbp_1
rlabel locali 19498 5118 19573 5184 1 x3.x42.SET_B
rlabel metal1 19517 5155 19575 5164 1 x3.x42.SET_B
rlabel metal1 19517 5118 19575 5127 1 x3.x42.SET_B
rlabel metal1 20253 5155 20311 5164 1 x3.x42.SET_B
rlabel metal1 19517 5127 20311 5155 1 x3.x42.SET_B
rlabel metal1 20253 5118 20311 5127 1 x3.x42.SET_B
rlabel metal1 18673 4923 21065 5019 1 x3.x42.VGND
rlabel metal1 18673 5467 21065 5563 1 x3.x42.VPWR
flabel locali 21519 5190 21594 5236 0 FreeSans 400 0 0 0 x3.x39.RESET_B
flabel locali 23393 4954 23427 4988 7 FreeSans 400 0 0 0 x3.x39.VGND
flabel locali 23393 5192 23427 5226 0 FreeSans 400 0 0 0 x3.x39.CLK
flabel locali 23393 5260 23427 5294 0 FreeSans 400 0 0 0 x3.x39.CLK
flabel locali 22657 5124 22691 5158 0 FreeSans 400 0 0 0 x3.x39.SET_B
flabel locali 21095 5056 21129 5090 0 FreeSans 400 0 0 0 x3.x39.Q
flabel locali 21095 5328 21129 5362 0 FreeSans 400 0 0 0 x3.x39.Q
flabel locali 21095 5396 21129 5430 0 FreeSans 400 0 0 0 x3.x39.Q
flabel locali 23393 5498 23427 5532 7 FreeSans 400 0 0 0 x3.x39.VPWR
flabel locali 23025 5192 23059 5226 0 FreeSans 200 0 0 0 x3.x39.D
flabel locali 23025 5260 23059 5294 0 FreeSans 200 0 0 0 x3.x39.D
flabel locali 21375 5396 21409 5430 0 FreeSans 400 0 0 0 x3.x39.Q_N
flabel locali 21375 5328 21409 5362 0 FreeSans 400 0 0 0 x3.x39.Q_N
flabel locali 21375 5056 21409 5090 0 FreeSans 400 0 0 0 x3.x39.Q_N
flabel metal1 23393 4954 23427 4988 0 FreeSans 200 0 0 0 x3.x39.VGND
flabel metal1 23393 5498 23427 5532 0 FreeSans 200 0 0 0 x3.x39.VPWR
flabel nwell 23393 5498 23427 5532 7 FreeSans 400 0 0 0 x3.x39.VPB
flabel nwell 23410 5515 23410 5515 0 FreeSans 200 0 0 0 x3.x39.VPB
flabel pwell 23393 4954 23427 4988 7 FreeSans 400 0 0 0 x3.x39.VNB
flabel pwell 23410 4971 23410 4971 0 FreeSans 200 0 0 0 x3.x39.VNB
rlabel comment 23457 4971 23457 4971 6 x3.x39.dfbbp_1
rlabel locali 21890 5118 21965 5184 1 x3.x39.SET_B
rlabel metal1 21909 5155 21967 5164 1 x3.x39.SET_B
rlabel metal1 21909 5118 21967 5127 1 x3.x39.SET_B
rlabel metal1 22645 5155 22703 5164 1 x3.x39.SET_B
rlabel metal1 21909 5127 22703 5155 1 x3.x39.SET_B
rlabel metal1 22645 5118 22703 5127 1 x3.x39.SET_B
rlabel metal1 21065 4923 23457 5019 1 x3.x39.VGND
rlabel metal1 21065 5467 23457 5563 1 x3.x39.VPWR
flabel locali 22928 5879 23003 5925 0 FreeSans 400 0 0 0 x3.x36.RESET_B
flabel locali 21095 5643 21129 5677 3 FreeSans 400 0 0 0 x3.x36.VGND
flabel locali 21095 5881 21129 5915 0 FreeSans 400 0 0 0 x3.x36.CLK
flabel locali 21095 5949 21129 5983 0 FreeSans 400 0 0 0 x3.x36.CLK
flabel locali 21831 5813 21865 5847 0 FreeSans 400 0 0 0 x3.x36.SET_B
flabel locali 23393 5745 23427 5779 0 FreeSans 400 0 0 0 x3.x36.Q
flabel locali 23393 6017 23427 6051 0 FreeSans 400 0 0 0 x3.x36.Q
flabel locali 23393 6085 23427 6119 0 FreeSans 400 0 0 0 x3.x36.Q
flabel locali 21095 6187 21129 6221 3 FreeSans 400 0 0 0 x3.x36.VPWR
flabel locali 21463 5881 21497 5915 0 FreeSans 200 0 0 0 x3.x36.D
flabel locali 21463 5949 21497 5983 0 FreeSans 200 0 0 0 x3.x36.D
flabel locali 23113 6085 23147 6119 0 FreeSans 400 0 0 0 x3.x36.Q_N
flabel locali 23113 6017 23147 6051 0 FreeSans 400 0 0 0 x3.x36.Q_N
flabel locali 23113 5745 23147 5779 0 FreeSans 400 0 0 0 x3.x36.Q_N
flabel metal1 21095 5643 21129 5677 0 FreeSans 200 0 0 0 x3.x36.VGND
flabel metal1 21095 6187 21129 6221 0 FreeSans 200 0 0 0 x3.x36.VPWR
flabel nwell 21095 6187 21129 6221 3 FreeSans 400 0 0 0 x3.x36.VPB
flabel nwell 21112 6204 21112 6204 0 FreeSans 200 0 0 0 x3.x36.VPB
flabel pwell 21095 5643 21129 5677 3 FreeSans 400 0 0 0 x3.x36.VNB
flabel pwell 21112 5660 21112 5660 0 FreeSans 200 0 0 0 x3.x36.VNB
rlabel comment 21065 5660 21065 5660 4 x3.x36.dfbbp_1
rlabel locali 22557 5807 22632 5873 1 x3.x36.SET_B
rlabel metal1 22555 5844 22613 5853 1 x3.x36.SET_B
rlabel metal1 22555 5807 22613 5816 1 x3.x36.SET_B
rlabel metal1 21819 5844 21877 5853 1 x3.x36.SET_B
rlabel metal1 21819 5816 22613 5844 1 x3.x36.SET_B
rlabel metal1 21819 5807 21877 5816 1 x3.x36.SET_B
rlabel metal1 21065 5612 23457 5708 1 x3.x36.VGND
rlabel metal1 21065 6156 23457 6252 1 x3.x36.VPWR
flabel locali 20536 5879 20611 5925 0 FreeSans 400 0 0 0 x3.x33.RESET_B
flabel locali 18703 5643 18737 5677 3 FreeSans 400 0 0 0 x3.x33.VGND
flabel locali 18703 5881 18737 5915 0 FreeSans 400 0 0 0 x3.x33.CLK
flabel locali 18703 5949 18737 5983 0 FreeSans 400 0 0 0 x3.x33.CLK
flabel locali 19439 5813 19473 5847 0 FreeSans 400 0 0 0 x3.x33.SET_B
flabel locali 21001 5745 21035 5779 0 FreeSans 400 0 0 0 x3.x33.Q
flabel locali 21001 6017 21035 6051 0 FreeSans 400 0 0 0 x3.x33.Q
flabel locali 21001 6085 21035 6119 0 FreeSans 400 0 0 0 x3.x33.Q
flabel locali 18703 6187 18737 6221 3 FreeSans 400 0 0 0 x3.x33.VPWR
flabel locali 19071 5881 19105 5915 0 FreeSans 200 0 0 0 x3.x33.D
flabel locali 19071 5949 19105 5983 0 FreeSans 200 0 0 0 x3.x33.D
flabel locali 20721 6085 20755 6119 0 FreeSans 400 0 0 0 x3.x33.Q_N
flabel locali 20721 6017 20755 6051 0 FreeSans 400 0 0 0 x3.x33.Q_N
flabel locali 20721 5745 20755 5779 0 FreeSans 400 0 0 0 x3.x33.Q_N
flabel metal1 18703 5643 18737 5677 0 FreeSans 200 0 0 0 x3.x33.VGND
flabel metal1 18703 6187 18737 6221 0 FreeSans 200 0 0 0 x3.x33.VPWR
flabel nwell 18703 6187 18737 6221 3 FreeSans 400 0 0 0 x3.x33.VPB
flabel nwell 18720 6204 18720 6204 0 FreeSans 200 0 0 0 x3.x33.VPB
flabel pwell 18703 5643 18737 5677 3 FreeSans 400 0 0 0 x3.x33.VNB
flabel pwell 18720 5660 18720 5660 0 FreeSans 200 0 0 0 x3.x33.VNB
rlabel comment 18673 5660 18673 5660 4 x3.x33.dfbbp_1
rlabel locali 20165 5807 20240 5873 1 x3.x33.SET_B
rlabel metal1 20163 5844 20221 5853 1 x3.x33.SET_B
rlabel metal1 20163 5807 20221 5816 1 x3.x33.SET_B
rlabel metal1 19427 5844 19485 5853 1 x3.x33.SET_B
rlabel metal1 19427 5816 20221 5844 1 x3.x33.SET_B
rlabel metal1 19427 5807 19485 5816 1 x3.x33.SET_B
rlabel metal1 18673 5612 21065 5708 1 x3.x33.VGND
rlabel metal1 18673 6156 21065 6252 1 x3.x33.VPWR
flabel locali 18144 5879 18219 5925 0 FreeSans 400 0 0 0 x3.x30.RESET_B
flabel locali 16311 5643 16345 5677 3 FreeSans 400 0 0 0 x3.x30.VGND
flabel locali 16311 5881 16345 5915 0 FreeSans 400 0 0 0 x3.x30.CLK
flabel locali 16311 5949 16345 5983 0 FreeSans 400 0 0 0 x3.x30.CLK
flabel locali 17047 5813 17081 5847 0 FreeSans 400 0 0 0 x3.x30.SET_B
flabel locali 18609 5745 18643 5779 0 FreeSans 400 0 0 0 x3.x30.Q
flabel locali 18609 6017 18643 6051 0 FreeSans 400 0 0 0 x3.x30.Q
flabel locali 18609 6085 18643 6119 0 FreeSans 400 0 0 0 x3.x30.Q
flabel locali 16311 6187 16345 6221 3 FreeSans 400 0 0 0 x3.x30.VPWR
flabel locali 16679 5881 16713 5915 0 FreeSans 200 0 0 0 x3.x30.D
flabel locali 16679 5949 16713 5983 0 FreeSans 200 0 0 0 x3.x30.D
flabel locali 18329 6085 18363 6119 0 FreeSans 400 0 0 0 x3.x30.Q_N
flabel locali 18329 6017 18363 6051 0 FreeSans 400 0 0 0 x3.x30.Q_N
flabel locali 18329 5745 18363 5779 0 FreeSans 400 0 0 0 x3.x30.Q_N
flabel metal1 16311 5643 16345 5677 0 FreeSans 200 0 0 0 x3.x30.VGND
flabel metal1 16311 6187 16345 6221 0 FreeSans 200 0 0 0 x3.x30.VPWR
flabel nwell 16311 6187 16345 6221 3 FreeSans 400 0 0 0 x3.x30.VPB
flabel nwell 16328 6204 16328 6204 0 FreeSans 200 0 0 0 x3.x30.VPB
flabel pwell 16311 5643 16345 5677 3 FreeSans 400 0 0 0 x3.x30.VNB
flabel pwell 16328 5660 16328 5660 0 FreeSans 200 0 0 0 x3.x30.VNB
rlabel comment 16281 5660 16281 5660 4 x3.x30.dfbbp_1
rlabel locali 17773 5807 17848 5873 1 x3.x30.SET_B
rlabel metal1 17771 5844 17829 5853 1 x3.x30.SET_B
rlabel metal1 17771 5807 17829 5816 1 x3.x30.SET_B
rlabel metal1 17035 5844 17093 5853 1 x3.x30.SET_B
rlabel metal1 17035 5816 17829 5844 1 x3.x30.SET_B
rlabel metal1 17035 5807 17093 5816 1 x3.x30.SET_B
rlabel metal1 16281 5612 18673 5708 1 x3.x30.VGND
rlabel metal1 16281 6156 18673 6252 1 x3.x30.VPWR
flabel locali 15752 5879 15827 5925 0 FreeSans 400 0 0 0 x3.x27.RESET_B
flabel locali 13919 5643 13953 5677 3 FreeSans 400 0 0 0 x3.x27.VGND
flabel locali 13919 5881 13953 5915 0 FreeSans 400 0 0 0 x3.x27.CLK
flabel locali 13919 5949 13953 5983 0 FreeSans 400 0 0 0 x3.x27.CLK
flabel locali 14655 5813 14689 5847 0 FreeSans 400 0 0 0 x3.x27.SET_B
flabel locali 16217 5745 16251 5779 0 FreeSans 400 0 0 0 x3.x27.Q
flabel locali 16217 6017 16251 6051 0 FreeSans 400 0 0 0 x3.x27.Q
flabel locali 16217 6085 16251 6119 0 FreeSans 400 0 0 0 x3.x27.Q
flabel locali 13919 6187 13953 6221 3 FreeSans 400 0 0 0 x3.x27.VPWR
flabel locali 14287 5881 14321 5915 0 FreeSans 200 0 0 0 x3.x27.D
flabel locali 14287 5949 14321 5983 0 FreeSans 200 0 0 0 x3.x27.D
flabel locali 15937 6085 15971 6119 0 FreeSans 400 0 0 0 x3.x27.Q_N
flabel locali 15937 6017 15971 6051 0 FreeSans 400 0 0 0 x3.x27.Q_N
flabel locali 15937 5745 15971 5779 0 FreeSans 400 0 0 0 x3.x27.Q_N
flabel metal1 13919 5643 13953 5677 0 FreeSans 200 0 0 0 x3.x27.VGND
flabel metal1 13919 6187 13953 6221 0 FreeSans 200 0 0 0 x3.x27.VPWR
flabel nwell 13919 6187 13953 6221 3 FreeSans 400 0 0 0 x3.x27.VPB
flabel nwell 13936 6204 13936 6204 0 FreeSans 200 0 0 0 x3.x27.VPB
flabel pwell 13919 5643 13953 5677 3 FreeSans 400 0 0 0 x3.x27.VNB
flabel pwell 13936 5660 13936 5660 0 FreeSans 200 0 0 0 x3.x27.VNB
rlabel comment 13889 5660 13889 5660 4 x3.x27.dfbbp_1
rlabel locali 15381 5807 15456 5873 1 x3.x27.SET_B
rlabel metal1 15379 5844 15437 5853 1 x3.x27.SET_B
rlabel metal1 15379 5807 15437 5816 1 x3.x27.SET_B
rlabel metal1 14643 5844 14701 5853 1 x3.x27.SET_B
rlabel metal1 14643 5816 15437 5844 1 x3.x27.SET_B
rlabel metal1 14643 5807 14701 5816 1 x3.x27.SET_B
rlabel metal1 13889 5612 16281 5708 1 x3.x27.VGND
rlabel metal1 13889 6156 16281 6252 1 x3.x27.VPWR
flabel locali 13360 5879 13435 5925 0 FreeSans 400 0 0 0 x3.x20.RESET_B
flabel locali 11527 5643 11561 5677 3 FreeSans 400 0 0 0 x3.x20.VGND
flabel locali 11527 5881 11561 5915 0 FreeSans 400 0 0 0 x3.x20.CLK
flabel locali 11527 5949 11561 5983 0 FreeSans 400 0 0 0 x3.x20.CLK
flabel locali 12263 5813 12297 5847 0 FreeSans 400 0 0 0 x3.x20.SET_B
flabel locali 13825 5745 13859 5779 0 FreeSans 400 0 0 0 x3.x20.Q
flabel locali 13825 6017 13859 6051 0 FreeSans 400 0 0 0 x3.x20.Q
flabel locali 13825 6085 13859 6119 0 FreeSans 400 0 0 0 x3.x20.Q
flabel locali 11527 6187 11561 6221 3 FreeSans 400 0 0 0 x3.x20.VPWR
flabel locali 11895 5881 11929 5915 0 FreeSans 200 0 0 0 x3.x20.D
flabel locali 11895 5949 11929 5983 0 FreeSans 200 0 0 0 x3.x20.D
flabel locali 13545 6085 13579 6119 0 FreeSans 400 0 0 0 x3.x20.Q_N
flabel locali 13545 6017 13579 6051 0 FreeSans 400 0 0 0 x3.x20.Q_N
flabel locali 13545 5745 13579 5779 0 FreeSans 400 0 0 0 x3.x20.Q_N
flabel metal1 11527 5643 11561 5677 0 FreeSans 200 0 0 0 x3.x20.VGND
flabel metal1 11527 6187 11561 6221 0 FreeSans 200 0 0 0 x3.x20.VPWR
flabel nwell 11527 6187 11561 6221 3 FreeSans 400 0 0 0 x3.x20.VPB
flabel nwell 11544 6204 11544 6204 0 FreeSans 200 0 0 0 x3.x20.VPB
flabel pwell 11527 5643 11561 5677 3 FreeSans 400 0 0 0 x3.x20.VNB
flabel pwell 11544 5660 11544 5660 0 FreeSans 200 0 0 0 x3.x20.VNB
rlabel comment 11497 5660 11497 5660 4 x3.x20.dfbbp_1
rlabel locali 12989 5807 13064 5873 1 x3.x20.SET_B
rlabel metal1 12987 5844 13045 5853 1 x3.x20.SET_B
rlabel metal1 12987 5807 13045 5816 1 x3.x20.SET_B
rlabel metal1 12251 5844 12309 5853 1 x3.x20.SET_B
rlabel metal1 12251 5816 13045 5844 1 x3.x20.SET_B
rlabel metal1 12251 5807 12309 5816 1 x3.x20.SET_B
rlabel metal1 11497 5612 13889 5708 1 x3.x20.VGND
rlabel metal1 11497 6156 13889 6252 1 x3.x20.VPWR
flabel metal1 11395 4624 11429 4658 0 FreeSans 200 0 0 0 x3.x7.VPWR
flabel metal1 11395 4080 11429 4114 0 FreeSans 200 0 0 0 x3.x7.VGND
flabel locali 11671 4318 11705 4352 0 FreeSans 200 0 0 0 x3.x7.X
flabel locali 11671 4386 11705 4420 0 FreeSans 200 0 0 0 x3.x7.X
flabel locali 11671 4250 11705 4284 0 FreeSans 200 0 0 0 x3.x7.X
flabel locali 11395 4624 11429 4658 0 FreeSans 200 0 0 0 x3.x7.VPWR
flabel locali 11395 4080 11429 4114 0 FreeSans 200 0 0 0 x3.x7.VGND
flabel locali 11395 4318 11429 4352 0 FreeSans 200 0 0 0 x3.x7.A
flabel nwell 11395 4624 11429 4658 0 FreeSans 200 0 0 0 x3.x7.VPB
flabel pwell 11395 4080 11429 4114 0 FreeSans 200 0 0 0 x3.x7.VNB
rlabel comment 11365 4097 11365 4097 4 x3.x7.buf_4
rlabel metal1 11365 4049 11917 4145 1 x3.x7.VGND
rlabel metal1 11365 4593 11917 4689 1 x3.x7.VPWR
flabel metal1 11120 4080 11154 4114 0 FreeSans 200 0 0 0 x3.x6.VGND
flabel metal1 11118 4624 11152 4658 0 FreeSans 200 0 0 0 x3.x6.VPWR
flabel locali 11118 4624 11152 4658 0 FreeSans 200 0 0 0 x3.x6.VPWR
flabel locali 11120 4080 11154 4114 0 FreeSans 200 0 0 0 x3.x6.VGND
flabel locali 11300 4182 11334 4216 0 FreeSans 200 0 0 0 x3.x6.X
flabel locali 11300 4454 11334 4488 0 FreeSans 200 0 0 0 x3.x6.X
flabel locali 11300 4522 11334 4556 0 FreeSans 200 0 0 0 x3.x6.X
flabel locali 11118 4318 11152 4352 0 FreeSans 200 0 0 0 x3.x6.A
flabel nwell 11118 4624 11152 4658 0 FreeSans 200 0 0 0 x3.x6.VPB
flabel pwell 11120 4080 11154 4114 0 FreeSans 200 0 0 0 x3.x6.VNB
rlabel comment 11089 4097 11089 4097 4 x3.x6.buf_1
rlabel metal1 11089 4049 11365 4145 1 x3.x6.VGND
rlabel metal1 11089 4593 11365 4689 1 x3.x6.VPWR
flabel metal1 11804 7060 11838 7094 0 FreeSans 200 0 0 0 x3.x5.VPWR
flabel metal1 11804 6516 11838 6550 0 FreeSans 200 0 0 0 x3.x5.VGND
flabel locali 12080 6754 12114 6788 0 FreeSans 200 0 0 0 x3.x5.X
flabel locali 12080 6822 12114 6856 0 FreeSans 200 0 0 0 x3.x5.X
flabel locali 12080 6686 12114 6720 0 FreeSans 200 0 0 0 x3.x5.X
flabel locali 11804 7060 11838 7094 0 FreeSans 200 0 0 0 x3.x5.VPWR
flabel locali 11804 6516 11838 6550 0 FreeSans 200 0 0 0 x3.x5.VGND
flabel locali 11804 6754 11838 6788 0 FreeSans 200 0 0 0 x3.x5.A
flabel nwell 11804 7060 11838 7094 0 FreeSans 200 0 0 0 x3.x5.VPB
flabel pwell 11804 6516 11838 6550 0 FreeSans 200 0 0 0 x3.x5.VNB
rlabel comment 11774 6533 11774 6533 4 x3.x5.buf_4
rlabel metal1 11774 6485 12326 6581 1 x3.x5.VGND
rlabel metal1 11774 7029 12326 7125 1 x3.x5.VPWR
flabel locali 12263 5192 12297 5226 0 FreeSans 200 0 0 0 x3.x4.A
flabel locali 12171 5192 12205 5226 0 FreeSans 200 0 0 0 x3.x4.A
flabel locali 13826 5192 13860 5226 0 FreeSans 200 0 0 0 x3.x4.X
flabel locali 13826 5260 13860 5294 0 FreeSans 200 0 0 0 x3.x4.X
flabel pwell 11895 4954 11929 4988 0 FreeSans 200 0 0 0 x3.x4.VNB
flabel nwell 11895 5498 11929 5532 0 FreeSans 200 0 0 0 x3.x4.VPB
flabel metal1 11895 4954 11929 4988 0 FreeSans 200 0 0 0 x3.x4.VGND
flabel metal1 11895 5498 11929 5532 0 FreeSans 200 0 0 0 x3.x4.VPWR
rlabel comment 11865 4971 11865 4971 4 x3.x4.buf_16
rlabel metal1 11865 4923 13889 5019 1 x3.x4.VGND
rlabel metal1 11865 5467 13889 5563 1 x3.x4.VPWR
flabel metal1 11363 5498 11397 5532 0 FreeSans 200 0 0 0 x3.x3.VPWR
flabel metal1 11363 4954 11397 4988 0 FreeSans 200 0 0 0 x3.x3.VGND
flabel locali 11639 5192 11673 5226 0 FreeSans 200 0 0 0 x3.x3.X
flabel locali 11639 5260 11673 5294 0 FreeSans 200 0 0 0 x3.x3.X
flabel locali 11639 5124 11673 5158 0 FreeSans 200 0 0 0 x3.x3.X
flabel locali 11363 5498 11397 5532 0 FreeSans 200 0 0 0 x3.x3.VPWR
flabel locali 11363 4954 11397 4988 0 FreeSans 200 0 0 0 x3.x3.VGND
flabel locali 11363 5192 11397 5226 0 FreeSans 200 0 0 0 x3.x3.A
flabel nwell 11363 5498 11397 5532 0 FreeSans 200 0 0 0 x3.x3.VPB
flabel pwell 11363 4954 11397 4988 0 FreeSans 200 0 0 0 x3.x3.VNB
rlabel comment 11333 4971 11333 4971 4 x3.x3.buf_4
rlabel metal1 11333 4923 11885 5019 1 x3.x3.VGND
rlabel metal1 11333 5467 11885 5563 1 x3.x3.VPWR
flabel metal1 11529 6516 11563 6550 0 FreeSans 200 0 0 0 x3.x2.VGND
flabel metal1 11527 7060 11561 7094 0 FreeSans 200 0 0 0 x3.x2.VPWR
flabel locali 11527 7060 11561 7094 0 FreeSans 200 0 0 0 x3.x2.VPWR
flabel locali 11529 6516 11563 6550 0 FreeSans 200 0 0 0 x3.x2.VGND
flabel locali 11709 6618 11743 6652 0 FreeSans 200 0 0 0 x3.x2.X
flabel locali 11709 6890 11743 6924 0 FreeSans 200 0 0 0 x3.x2.X
flabel locali 11709 6958 11743 6992 0 FreeSans 200 0 0 0 x3.x2.X
flabel locali 11527 6754 11561 6788 0 FreeSans 200 0 0 0 x3.x2.A
flabel nwell 11527 7060 11561 7094 0 FreeSans 200 0 0 0 x3.x2.VPB
flabel pwell 11529 6516 11563 6550 0 FreeSans 200 0 0 0 x3.x2.VNB
rlabel comment 11498 6533 11498 6533 4 x3.x2.buf_1
rlabel metal1 11498 6485 11774 6581 1 x3.x2.VGND
rlabel metal1 11498 7029 11774 7125 1 x3.x2.VPWR
flabel metal1 11088 4954 11122 4988 0 FreeSans 200 0 0 0 x3.x1.VGND
flabel metal1 11086 5498 11120 5532 0 FreeSans 200 0 0 0 x3.x1.VPWR
flabel locali 11086 5498 11120 5532 0 FreeSans 200 0 0 0 x3.x1.VPWR
flabel locali 11088 4954 11122 4988 0 FreeSans 200 0 0 0 x3.x1.VGND
flabel locali 11268 5056 11302 5090 0 FreeSans 200 0 0 0 x3.x1.X
flabel locali 11268 5328 11302 5362 0 FreeSans 200 0 0 0 x3.x1.X
flabel locali 11268 5396 11302 5430 0 FreeSans 200 0 0 0 x3.x1.X
flabel locali 11086 5192 11120 5226 0 FreeSans 200 0 0 0 x3.x1.A
flabel nwell 11086 5498 11120 5532 0 FreeSans 200 0 0 0 x3.x1.VPB
flabel pwell 11088 4954 11122 4988 0 FreeSans 200 0 0 0 x3.x1.VNB
rlabel comment 11057 4971 11057 4971 4 x3.x1.buf_1
rlabel metal1 11057 4923 11333 5019 1 x3.x1.VGND
rlabel metal1 11057 5467 11333 5563 1 x3.x1.VPWR
flabel pwell 14534 6516 14568 6550 0 FreeSans 200 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.VNB
flabel nwell 14534 7060 14568 7094 0 FreeSans 200 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.VPB
flabel metal1 14534 6516 14568 6550 0 FreeSans 200 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.VGND
flabel metal1 14534 7060 14568 7094 0 FreeSans 200 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.VPWR
flabel locali 12878 6618 12912 6652 0 FreeSans 400 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.X
flabel locali 12878 6686 12912 6720 0 FreeSans 400 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.X
flabel locali 12878 6754 12912 6788 0 FreeSans 400 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.X
flabel locali 12878 6822 12912 6856 0 FreeSans 400 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.X
flabel locali 12878 6890 12912 6924 0 FreeSans 400 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.X
flabel locali 12878 6958 12912 6992 0 FreeSans 400 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.X
flabel locali 14534 6754 14568 6788 0 FreeSans 400 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.S0
flabel locali 14534 6822 14568 6856 0 FreeSans 400 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.S0
flabel locali 14350 6686 14384 6720 0 FreeSans 400 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.A2
flabel locali 14350 6618 14384 6652 0 FreeSans 400 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.A2
flabel locali 14074 6686 14108 6720 0 FreeSans 400 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.A3
flabel locali 14074 6754 14108 6788 0 FreeSans 400 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.A3
flabel locali 13982 6754 14016 6788 0 FreeSans 400 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.S1
flabel locali 13982 6686 14016 6720 0 FreeSans 400 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.S1
flabel locali 13614 6754 13648 6788 0 FreeSans 400 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.A1
flabel locali 13614 6686 13648 6720 0 FreeSans 400 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.A1
flabel locali 13246 6686 13280 6720 0 FreeSans 400 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.A0
flabel locali 13246 6618 13280 6652 0 FreeSans 400 0 0 0 x3.sky130_fd_sc_hd__mux4_4_0.A0
rlabel comment 14598 6533 14598 6533 6 x3.sky130_fd_sc_hd__mux4_4_0.mux4_4
rlabel locali 14319 6790 14353 6822 1 x3.sky130_fd_sc_hd__mux4_4_0.S0
rlabel locali 14319 6822 14396 6856 1 x3.sky130_fd_sc_hd__mux4_4_0.S0
rlabel locali 13304 6782 13372 6862 1 x3.sky130_fd_sc_hd__mux4_4_0.S0
rlabel metal1 13326 6853 13384 6862 1 x3.sky130_fd_sc_hd__mux4_4_0.S0
rlabel metal1 13326 6816 13384 6825 1 x3.sky130_fd_sc_hd__mux4_4_0.S0
rlabel metal1 14338 6853 14396 6862 1 x3.sky130_fd_sc_hd__mux4_4_0.S0
rlabel metal1 14338 6816 14396 6825 1 x3.sky130_fd_sc_hd__mux4_4_0.S0
rlabel metal1 14522 6853 14581 6862 1 x3.sky130_fd_sc_hd__mux4_4_0.S0
rlabel metal1 13326 6825 14581 6853 1 x3.sky130_fd_sc_hd__mux4_4_0.S0
rlabel metal1 14522 6816 14581 6825 1 x3.sky130_fd_sc_hd__mux4_4_0.S0
rlabel metal1 12758 6485 14598 6581 1 x3.sky130_fd_sc_hd__mux4_4_0.VGND
rlabel metal1 12758 7029 14598 7125 1 x3.sky130_fd_sc_hd__mux4_4_0.VPWR
flabel metal1 10914 11473 10957 11531 0 FreeSans 320 0 0 0 x2.set
flabel metal1 11199 11470 11232 11528 0 FreeSans 320 0 0 0 x2.reset
flabel metal1 13473 10493 13505 10605 0 FreeSans 320 0 0 0 x2.sample_delay_offset
flabel metal1 13479 10913 13504 10941 0 FreeSans 320 0 0 0 x2.CAP_CTRL_CODE0[2]
flabel metal1 13481 10857 13506 10885 0 FreeSans 320 0 0 0 x2.CAP_CTRL_CODE0[1]
flabel metal1 13483 10801 13508 10829 0 FreeSans 320 0 0 0 x2.CAP_CTRL_CODE0[0]
flabel metal1 13484 10745 13509 10773 0 FreeSans 320 0 0 0 x2.CAP_CTRL_CODE1[2]
flabel metal1 13486 10689 13511 10717 0 FreeSans 320 0 0 0 x2.CAP_CTRL_CODE1[1]
flabel metal1 13485 10633 13510 10661 0 FreeSans 320 0 0 0 x2.CAP_CTRL_CODE1[0]
flabel metal1 13481 10437 13506 10465 0 FreeSans 320 0 0 0 x2.CAP_CTRL_CODE2[2]
flabel metal1 13484 10381 13509 10409 0 FreeSans 320 0 0 0 x2.CAP_CTRL_CODE2[1]
flabel metal1 13486 10325 13511 10353 0 FreeSans 320 0 0 0 x2.CAP_CTRL_CODE2[0]
flabel metal1 13481 10269 13506 10297 0 FreeSans 320 0 0 0 x2.CAP_CTRL_CODE3[2]
flabel metal1 13484 10213 13509 10241 0 FreeSans 320 0 0 0 x2.CAP_CTRL_CODE3[1]
flabel metal1 13484 10157 13509 10185 0 FreeSans 320 0 0 0 x2.CAP_CTRL_CODE3[0]
flabel metal1 13198 12668 13224 12702 0 FreeSans 320 0 0 0 x2.CAP_CTRL_CODE0[3]
flabel metal1 19914 12668 19940 12702 0 FreeSans 320 0 0 0 x2.CAP_CTRL_CODE1[3]
flabel metal1 26659 8407 26685 8441 0 FreeSans 320 0 0 0 x2.CAP_CTRL_CODE2[3]
flabel metal1 19956 8407 19982 8441 0 FreeSans 320 0 0 0 x2.CAP_CTRL_CODE3[3]
flabel metal4 10645 12760 13437 13747 0 FreeSans 320 0 0 0 x2.vdd
flabel metal4 10878 9481 12863 11301 0 FreeSans 320 0 0 0 x2.vss
flabel metal1 11827 7941 11873 8087 0 FreeSans 320 0 0 0 x2.sample_clk_b
flabel metal1 11826 8724 11874 8888 0 FreeSans 320 0 0 0 x2.sample_clk
flabel metal1 10869 12169 10912 12233 0 FreeSans 320 0 0 0 x2.clk
flabel locali 12771 8919 12805 8953 0 FreeSans 250 0 0 0 x2.x3.Y
flabel locali 12771 8851 12805 8885 0 FreeSans 250 0 0 0 x2.x3.Y
flabel locali 12771 8783 12805 8817 0 FreeSans 250 0 0 0 x2.x3.Y
flabel locali 12863 8783 12897 8817 0 FreeSans 250 0 0 0 x2.x3.B
flabel locali 12679 8783 12713 8817 0 FreeSans 250 0 0 0 x2.x3.A
flabel nwell 12863 8477 12897 8511 0 FreeSans 200 0 0 0 x2.x3.VPB
flabel pwell 12863 9021 12897 9055 0 FreeSans 200 0 0 0 x2.x3.VNB
flabel metal1 12863 9021 12897 9055 0 FreeSans 200 0 0 0 x2.x3.VGND
flabel metal1 12863 8477 12897 8511 0 FreeSans 200 0 0 0 x2.x3.VPWR
rlabel comment 12925 9038 12925 9038 8 x2.x3.nand2_1
rlabel metal1 12649 8990 12925 9086 5 x2.x3.VGND
rlabel metal1 12649 8446 12925 8542 5 x2.x3.VPWR
flabel locali 13003 8715 13037 8749 0 FreeSans 340 0 0 0 x2.x7.Y
flabel locali 13003 8783 13037 8817 0 FreeSans 340 0 0 0 x2.x7.Y
flabel locali 13095 8783 13129 8817 0 FreeSans 340 0 0 0 x2.x7.A
flabel metal1 13138 9021 13172 9055 0 FreeSans 200 0 0 0 x2.x7.VGND
flabel metal1 13138 8477 13172 8511 0 FreeSans 200 0 0 0 x2.x7.VPWR
rlabel comment 13201 9038 13201 9038 8 x2.x7.inv_1
rlabel metal1 12925 8990 13201 9086 5 x2.x7.VGND
rlabel metal1 12925 8446 13201 8542 5 x2.x7.VPWR
flabel pwell 13138 9021 13172 9055 0 FreeSans 200 0 0 0 x2.x7.VNB
flabel nwell 13138 8477 13172 8511 0 FreeSans 200 0 0 0 x2.x7.VPB
flabel metal1 10931 11473 10957 11531 0 FreeSans 320 0 0 0 x2.x1.set
flabel metal1 11205 11471 11228 11529 0 FreeSans 320 0 0 0 x2.x1.reset
flabel metal1 10876 12169 10912 12234 0 FreeSans 320 0 0 0 x2.x1.clk
flabel space 13214 12102 13257 12320 0 FreeSans 320 0 0 0 x2.x1.div_clk
flabel locali 12745 12184 12820 12230 0 FreeSans 400 0 0 0 x2.x1.x2.RESET_B
flabel locali 10912 12432 10946 12466 3 FreeSans 400 0 0 0 x2.x1.x2.VGND
flabel locali 10912 12194 10946 12228 0 FreeSans 400 0 0 0 x2.x1.x2.CLK
flabel locali 10912 12126 10946 12160 0 FreeSans 400 0 0 0 x2.x1.x2.CLK
flabel locali 11648 12262 11682 12296 0 FreeSans 400 0 0 0 x2.x1.x2.SET_B
flabel locali 13210 12330 13244 12364 0 FreeSans 400 0 0 0 x2.x1.x2.Q
flabel locali 13210 12058 13244 12092 0 FreeSans 400 0 0 0 x2.x1.x2.Q
flabel locali 13210 11990 13244 12024 0 FreeSans 400 0 0 0 x2.x1.x2.Q
flabel locali 10912 11888 10946 11922 3 FreeSans 400 0 0 0 x2.x1.x2.VPWR
flabel locali 11280 12194 11314 12228 0 FreeSans 200 0 0 0 x2.x1.x2.D
flabel locali 11280 12126 11314 12160 0 FreeSans 200 0 0 0 x2.x1.x2.D
flabel locali 12930 11990 12964 12024 0 FreeSans 400 0 0 0 x2.x1.x2.Q_N
flabel locali 12930 12058 12964 12092 0 FreeSans 400 0 0 0 x2.x1.x2.Q_N
flabel locali 12930 12330 12964 12364 0 FreeSans 400 0 0 0 x2.x1.x2.Q_N
flabel metal1 10912 12432 10946 12466 0 FreeSans 200 0 0 0 x2.x1.x2.VGND
flabel metal1 10912 11888 10946 11922 0 FreeSans 200 0 0 0 x2.x1.x2.VPWR
flabel nwell 10912 11888 10946 11922 3 FreeSans 400 0 0 0 x2.x1.x2.VPB
flabel nwell 10929 11905 10929 11905 0 FreeSans 200 0 0 0 x2.x1.x2.VPB
flabel pwell 10912 12432 10946 12466 3 FreeSans 400 0 0 0 x2.x1.x2.VNB
flabel pwell 10929 12449 10929 12449 0 FreeSans 200 0 0 0 x2.x1.x2.VNB
rlabel comment 10882 12449 10882 12449 2 x2.x1.x2.dfbbp_1
rlabel locali 12374 12236 12449 12302 5 x2.x1.x2.SET_B
rlabel metal1 12372 12256 12430 12265 5 x2.x1.x2.SET_B
rlabel metal1 12372 12293 12430 12302 5 x2.x1.x2.SET_B
rlabel metal1 11636 12256 11694 12265 5 x2.x1.x2.SET_B
rlabel metal1 11636 12265 12430 12293 5 x2.x1.x2.SET_B
rlabel metal1 11636 12293 11694 12302 5 x2.x1.x2.SET_B
rlabel metal1 10882 12401 13274 12497 5 x2.x1.x2.VGND
rlabel metal1 10882 11857 13274 11953 5 x2.x1.x2.VPWR
flabel locali 11322 11554 11356 11588 0 FreeSans 340 0 0 0 x2.x1.x4.Y
flabel locali 11322 11486 11356 11520 0 FreeSans 340 0 0 0 x2.x1.x4.Y
flabel locali 11230 11486 11264 11520 0 FreeSans 340 0 0 0 x2.x1.x4.A
flabel metal1 11187 11248 11221 11282 0 FreeSans 200 0 0 0 x2.x1.x4.VGND
flabel metal1 11187 11792 11221 11826 0 FreeSans 200 0 0 0 x2.x1.x4.VPWR
rlabel comment 11158 11265 11158 11265 4 x2.x1.x4.inv_1
rlabel metal1 11158 11217 11434 11313 1 x2.x1.x4.VGND
rlabel metal1 11158 11761 11434 11857 1 x2.x1.x4.VPWR
flabel pwell 11187 11248 11221 11282 0 FreeSans 200 0 0 0 x2.x1.x4.VNB
flabel nwell 11187 11792 11221 11826 0 FreeSans 200 0 0 0 x2.x1.x4.VPB
flabel locali 11046 11554 11080 11588 0 FreeSans 340 0 0 0 x2.x1.x3.Y
flabel locali 11046 11486 11080 11520 0 FreeSans 340 0 0 0 x2.x1.x3.Y
flabel locali 10954 11486 10988 11520 0 FreeSans 340 0 0 0 x2.x1.x3.A
flabel metal1 10911 11248 10945 11282 0 FreeSans 200 0 0 0 x2.x1.x3.VGND
flabel metal1 10911 11792 10945 11826 0 FreeSans 200 0 0 0 x2.x1.x3.VPWR
rlabel comment 10882 11265 10882 11265 4 x2.x1.x3.inv_1
rlabel metal1 10882 11217 11158 11313 1 x2.x1.x3.VGND
rlabel metal1 10882 11761 11158 11857 1 x2.x1.x3.VPWR
flabel pwell 10911 11248 10945 11282 0 FreeSans 200 0 0 0 x2.x1.x3.VNB
flabel nwell 10911 11792 10945 11826 0 FreeSans 200 0 0 0 x2.x1.x3.VPB
flabel metal1 13236 8780 13290 8826 0 FreeSans 320 0 0 0 x2.x2.out
flabel metal4 13318 13626 26677 13690 0 FreeSans 320 0 0 0 x2.x2.VDD
flabel metal1 13495 10493 14112 10605 0 FreeSans 320 0 0 0 x2.x2.sample_delay_offset
flabel metal1 13249 12285 13917 12332 0 FreeSans 320 0 0 0 x2.x2.in
flabel metal1 13212 12668 13350 12702 0 FreeSans 320 0 0 0 x2.x2.sample_code0[3]
flabel metal1 19921 12668 20059 12702 0 FreeSans 320 0 0 0 x2.x2.sample_code1[3]
flabel metal1 26538 8407 26676 8441 0 FreeSans 320 0 0 0 x2.x2.sample_code2[3]
flabel metal1 19829 8407 19967 8441 0 FreeSans 320 0 0 0 x2.x2.sample_code3[3]
flabel metal1 13495 10689 24894 10717 0 FreeSans 320 0 0 0 x2.x2.sample_code1[1]
flabel metal1 13495 10633 25750 10661 0 FreeSans 320 0 0 0 x2.x2.sample_code1[0]
flabel metal1 13495 10157 14196 10185 0 FreeSans 320 0 0 0 x2.x2.sample_code3[0]
flabel metal1 13495 10213 15052 10241 0 FreeSans 320 0 0 0 x2.x2.sample_code3[1]
flabel metal1 13495 10269 17478 10297 0 FreeSans 320 0 0 0 x2.x2.sample_code3[2]
flabel metal1 13495 10325 20905 10353 0 FreeSans 320 0 0 0 x2.x2.sample_code2[0]
flabel metal1 13495 10381 21761 10409 0 FreeSans 320 0 0 0 x2.x2.sample_code2[1]
flabel metal1 13495 10437 24187 10465 0 FreeSans 320 0 0 0 x2.x2.sample_code2[2]
flabel metal1 13495 10745 22468 10773 0 FreeSans 320 0 0 0 x2.x2.sample_code1[2]
flabel metal4 25767 10111 26676 11044 0 FreeSans 320 0 0 0 x2.x2.VSS
flabel metal1 13495 10913 15759 10941 0 FreeSans 320 0 0 0 x2.x2.sample_code0[2]
flabel metal1 13495 10857 18185 10885 0 FreeSans 320 0 0 0 x2.x2.sample_code0[1]
flabel metal1 13495 10801 19041 10829 0 FreeSans 320 0 0 0 x2.x2.sample_code0[0]
flabel metal1 13249 12285 13917 12332 0 FreeSans 320 0 0 0 x2.x2.x4.IN
flabel metal1 19725 12283 19907 12329 0 FreeSans 320 0 0 0 x2.x2.x4.OUT
flabel metal1 13212 12668 13350 12702 0 FreeSans 320 0 0 0 x2.x2.x4.code[3]
flabel metal1 18127 10957 18185 12134 0 FreeSans 320 0 0 0 x2.x2.x4.code[1]
flabel metal1 15701 10957 15759 12134 0 FreeSans 320 0 0 0 x2.x2.x4.code[2]
flabel metal4 13318 13027 13736 13637 0 FreeSans 320 0 0 0 x2.x2.x4.VDD
flabel metal4 13346 10980 13722 12417 0 FreeSans 320 0 0 0 x2.x2.x4.VSS
flabel metal2 13676 12083 14112 12129 0 FreeSans 320 0 0 0 x2.x2.x4.code_offset
flabel metal1 18983 10956 19042 12137 0 FreeSans 320 0 0 0 x2.x2.x4.code[0]
flabel metal1 13860 12738 13894 12772 0 FreeSans 320 0 0 0 x2.x2.x4.x8.input_stack
flabel nwell 13904 13521 13938 13581 0 FreeSans 320 0 0 0 x2.x2.x4.x8.vdd
flabel metal1 13898 12819 13944 12831 0 FreeSans 320 0 0 0 x2.x2.x4.x8.output_stack
flabel poly 13837 12081 13939 12111 0 FreeSans 320 0 0 0 x2.x2.x4.x9.input_stack
flabel metal1 13951 11028 13985 11088 0 FreeSans 320 0 0 0 x2.x2.x4.x9.vss
flabel metal1 13945 12054 13991 12066 0 FreeSans 320 0 0 0 x2.x2.x4.x9.output_stack
flabel locali 13438 12738 13472 12772 0 FreeSans 340 0 0 0 x2.x2.x4.x10.Y
flabel locali 13438 12670 13472 12704 0 FreeSans 340 0 0 0 x2.x2.x4.x10.Y
flabel locali 13346 12670 13380 12704 0 FreeSans 340 0 0 0 x2.x2.x4.x10.A
flabel metal1 13303 12432 13337 12466 0 FreeSans 200 0 0 0 x2.x2.x4.x10.VGND
flabel metal1 13303 12976 13337 13010 0 FreeSans 200 0 0 0 x2.x2.x4.x10.VPWR
rlabel comment 13274 12449 13274 12449 4 x2.x2.x4.x10.inv_1
rlabel metal1 13274 12401 13550 12497 1 x2.x2.x4.x10.VGND
rlabel metal1 13274 12945 13550 13041 1 x2.x2.x4.x10.VPWR
flabel pwell 13303 12432 13337 12466 0 FreeSans 200 0 0 0 x2.x2.x4.x10.VNB
flabel nwell 13303 12976 13337 13010 0 FreeSans 200 0 0 0 x2.x2.x4.x10.VPB
flabel locali 13536 12738 13570 12772 0 FreeSans 340 0 0 0 x2.x2.x4.x11.Y
flabel locali 13536 12670 13570 12704 0 FreeSans 340 0 0 0 x2.x2.x4.x11.Y
flabel locali 13628 12670 13662 12704 0 FreeSans 340 0 0 0 x2.x2.x4.x11.A
flabel metal1 13671 12432 13705 12466 0 FreeSans 200 0 0 0 x2.x2.x4.x11.VGND
flabel metal1 13671 12976 13705 13010 0 FreeSans 200 0 0 0 x2.x2.x4.x11.VPWR
rlabel comment 13734 12449 13734 12449 6 x2.x2.x4.x11.inv_1
rlabel metal1 13458 12401 13734 12497 1 x2.x2.x4.x11.VGND
rlabel metal1 13458 12945 13734 13041 1 x2.x2.x4.x11.VPWR
flabel pwell 13671 12432 13705 12466 0 FreeSans 200 0 0 0 x2.x2.x4.x11.VNB
flabel nwell 13671 12976 13705 13010 0 FreeSans 200 0 0 0 x2.x2.x4.x11.VPB
flabel metal1 14502 12495 14536 12529 0 FreeSans 320 0 0 0 x2.x2.x4.x6.SW
flabel nwell 13946 13557 14616 13625 0 FreeSans 320 0 0 0 x2.x2.x4.x6.VDD
flabel pdiff 14534 12364 14592 12448 0 FreeSans 320 0 0 0 x2.x2.x4.x6.delay_signal
flabel metal4 13946 13556 14047 13625 0 FreeSans 320 0 0 0 x2.x2.x4.x6.VDD
flabel via3 14047 12398 14111 12462 0 FreeSans 320 0 0 0 x2.x2.x4.x6.floating
flabel viali 14855 12094 14889 12128 0 FreeSans 320 0 0 0 x2.x2.x4.x7.SW
flabel ndiff 14887 12166 14945 12250 0 FreeSans 320 0 0 0 x2.x2.x4.x7.delay_signal
flabel metal4 14294 10989 14966 11057 0 FreeSans 320 0 0 0 x2.x2.x4.x7.VSS
flabel via3 14398 12153 14462 12217 0 FreeSans 320 0 0 0 x2.x2.x4.x7.floating
flabel viali 15587 12094 15621 12128 0 FreeSans 320 0 0 0 x2.x2.x4.x4[3].SW
flabel ndiff 15619 12166 15677 12250 0 FreeSans 320 0 0 0 x2.x2.x4.x4[3].delay_signal
flabel metal4 15026 10989 15698 11057 0 FreeSans 320 0 0 0 x2.x2.x4.x4[3].VSS
flabel via3 15130 12153 15194 12217 0 FreeSans 320 0 0 0 x2.x2.x4.x4[3].floating
flabel metal1 15360 12498 15394 12532 0 FreeSans 320 0 0 0 x2.x2.x4.x5[6].SW
flabel nwell 15280 13560 15950 13628 0 FreeSans 320 0 0 0 x2.x2.x4.x5[6].VDD
flabel pdiff 15304 12367 15362 12451 0 FreeSans 320 0 0 0 x2.x2.x4.x5[6].delay_signal
flabel metal4 15849 13559 15950 13628 0 FreeSans 320 0 0 0 x2.x2.x4.x5[6].VDD
flabel via3 15785 12401 15849 12465 0 FreeSans 320 0 0 0 x2.x2.x4.x5[6].floating
flabel metal1 15234 12498 15268 12532 0 FreeSans 320 0 0 0 x2.x2.x4.x5[7].SW
flabel nwell 14678 13560 15348 13628 0 FreeSans 320 0 0 0 x2.x2.x4.x5[7].VDD
flabel pdiff 15266 12367 15324 12451 0 FreeSans 320 0 0 0 x2.x2.x4.x5[7].delay_signal
flabel metal4 14678 13559 14779 13628 0 FreeSans 320 0 0 0 x2.x2.x4.x5[7].VDD
flabel via3 14779 12401 14843 12465 0 FreeSans 320 0 0 0 x2.x2.x4.x5[7].floating
flabel viali 15709 12094 15743 12128 0 FreeSans 320 0 0 0 x2.x2.x4.x4[2].SW
flabel ndiff 15653 12166 15711 12250 0 FreeSans 320 0 0 0 x2.x2.x4.x4[2].delay_signal
flabel metal4 15632 10989 16304 11057 0 FreeSans 320 0 0 0 x2.x2.x4.x4[2].VSS
flabel via3 16136 12153 16200 12217 0 FreeSans 320 0 0 0 x2.x2.x4.x4[2].floating
flabel metal1 16446 12498 16480 12532 0 FreeSans 320 0 0 0 x2.x2.x4.x5[5].SW
flabel nwell 15890 13560 16560 13628 0 FreeSans 320 0 0 0 x2.x2.x4.x5[5].VDD
flabel pdiff 16478 12367 16536 12451 0 FreeSans 320 0 0 0 x2.x2.x4.x5[5].delay_signal
flabel metal4 15890 13559 15991 13628 0 FreeSans 320 0 0 0 x2.x2.x4.x5[5].VDD
flabel via3 15991 12401 16055 12465 0 FreeSans 320 0 0 0 x2.x2.x4.x5[5].floating
flabel viali 16799 12094 16833 12128 0 FreeSans 320 0 0 0 x2.x2.x4.x4[1].SW
flabel ndiff 16831 12166 16889 12250 0 FreeSans 320 0 0 0 x2.x2.x4.x4[1].delay_signal
flabel metal4 16238 10989 16910 11057 0 FreeSans 320 0 0 0 x2.x2.x4.x4[1].VSS
flabel via3 16342 12153 16406 12217 0 FreeSans 320 0 0 0 x2.x2.x4.x4[1].floating
flabel metal1 16572 12498 16606 12532 0 FreeSans 320 0 0 0 x2.x2.x4.x5[4].SW
flabel nwell 16492 13560 17162 13628 0 FreeSans 320 0 0 0 x2.x2.x4.x5[4].VDD
flabel pdiff 16516 12367 16574 12451 0 FreeSans 320 0 0 0 x2.x2.x4.x5[4].delay_signal
flabel metal4 17061 13559 17162 13628 0 FreeSans 320 0 0 0 x2.x2.x4.x5[4].VDD
flabel via3 16997 12401 17061 12465 0 FreeSans 320 0 0 0 x2.x2.x4.x5[4].floating
flabel viali 16921 12094 16955 12128 0 FreeSans 320 0 0 0 x2.x2.x4.x4[0].SW
flabel ndiff 16865 12166 16923 12250 0 FreeSans 320 0 0 0 x2.x2.x4.x4[0].delay_signal
flabel metal4 16844 10989 17516 11057 0 FreeSans 320 0 0 0 x2.x2.x4.x4[0].VSS
flabel via3 17348 12153 17412 12217 0 FreeSans 320 0 0 0 x2.x2.x4.x4[0].floating
flabel metal1 17658 12498 17692 12532 0 FreeSans 320 0 0 0 x2.x2.x4.x5[3].SW
flabel nwell 17102 13560 17772 13628 0 FreeSans 320 0 0 0 x2.x2.x4.x5[3].VDD
flabel pdiff 17690 12367 17748 12451 0 FreeSans 320 0 0 0 x2.x2.x4.x5[3].delay_signal
flabel metal4 17102 13559 17203 13628 0 FreeSans 320 0 0 0 x2.x2.x4.x5[3].VDD
flabel via3 17203 12401 17267 12465 0 FreeSans 320 0 0 0 x2.x2.x4.x5[3].floating
flabel viali 18137 12094 18171 12128 0 FreeSans 320 0 0 0 x2.x2.x4.x3[1].SW
flabel ndiff 18169 12166 18227 12250 0 FreeSans 320 0 0 0 x2.x2.x4.x3[1].delay_signal
flabel metal4 17576 10989 18248 11057 0 FreeSans 320 0 0 0 x2.x2.x4.x3[1].VSS
flabel via3 17680 12153 17744 12217 0 FreeSans 320 0 0 0 x2.x2.x4.x3[1].floating
flabel metal1 17784 12498 17818 12532 0 FreeSans 320 0 0 0 x2.x2.x4.x5[2].SW
flabel nwell 17704 13560 18374 13628 0 FreeSans 320 0 0 0 x2.x2.x4.x5[2].VDD
flabel pdiff 17728 12367 17786 12451 0 FreeSans 320 0 0 0 x2.x2.x4.x5[2].delay_signal
flabel metal4 18273 13559 18374 13628 0 FreeSans 320 0 0 0 x2.x2.x4.x5[2].VDD
flabel via3 18209 12401 18273 12465 0 FreeSans 320 0 0 0 x2.x2.x4.x5[2].floating
flabel viali 18259 12094 18293 12128 0 FreeSans 320 0 0 0 x2.x2.x4.x3[0].SW
flabel ndiff 18203 12166 18261 12250 0 FreeSans 320 0 0 0 x2.x2.x4.x3[0].delay_signal
flabel metal4 18182 10989 18854 11057 0 FreeSans 320 0 0 0 x2.x2.x4.x3[0].VSS
flabel via3 18686 12153 18750 12217 0 FreeSans 320 0 0 0 x2.x2.x4.x3[0].floating
flabel metal1 18870 12498 18904 12532 0 FreeSans 320 0 0 0 x2.x2.x4.x5[1].SW
flabel nwell 18314 13560 18984 13628 0 FreeSans 320 0 0 0 x2.x2.x4.x5[1].VDD
flabel pdiff 18902 12367 18960 12451 0 FreeSans 320 0 0 0 x2.x2.x4.x5[1].delay_signal
flabel metal4 18314 13559 18415 13628 0 FreeSans 320 0 0 0 x2.x2.x4.x5[1].VDD
flabel via3 18415 12401 18479 12465 0 FreeSans 320 0 0 0 x2.x2.x4.x5[1].floating
flabel viali 18993 12094 19027 12128 0 FreeSans 320 0 0 0 x2.x2.x4.x2.SW
flabel ndiff 18937 12166 18995 12250 0 FreeSans 320 0 0 0 x2.x2.x4.x2.delay_signal
flabel metal4 18916 10989 19588 11057 0 FreeSans 320 0 0 0 x2.x2.x4.x2.VSS
flabel via3 19420 12153 19484 12217 0 FreeSans 320 0 0 0 x2.x2.x4.x2.floating
flabel metal1 18996 12498 19030 12532 0 FreeSans 320 0 0 0 x2.x2.x4.x5[0].SW
flabel nwell 18916 13560 19586 13628 0 FreeSans 320 0 0 0 x2.x2.x4.x5[0].VDD
flabel pdiff 18940 12367 18998 12451 0 FreeSans 320 0 0 0 x2.x2.x4.x5[0].delay_signal
flabel metal4 19485 13559 19586 13628 0 FreeSans 320 0 0 0 x2.x2.x4.x5[0].VDD
flabel via3 19421 12401 19485 12465 0 FreeSans 320 0 0 0 x2.x2.x4.x5[0].floating
flabel metal1 19262 8777 19930 8824 0 FreeSans 320 0 0 0 x2.x2.x3.IN
flabel metal1 13272 8780 13454 8826 0 FreeSans 320 0 0 0 x2.x2.x3.OUT
flabel metal1 19829 8407 19967 8441 0 FreeSans 320 0 0 0 x2.x2.x3.code[3]
flabel metal1 14994 8975 15052 10152 0 FreeSans 320 0 0 0 x2.x2.x3.code[1]
flabel metal1 17420 8975 17478 10152 0 FreeSans 320 0 0 0 x2.x2.x3.code[2]
flabel metal4 19443 7472 19861 8082 0 FreeSans 320 0 0 0 x2.x2.x3.VDD
flabel metal4 19457 8692 19833 10129 0 FreeSans 320 0 0 0 x2.x2.x3.VSS
flabel metal2 19067 8980 19503 9026 0 FreeSans 320 0 0 0 x2.x2.x3.code_offset
flabel metal1 14137 8972 14196 10153 0 FreeSans 320 0 0 0 x2.x2.x3.code[0]
flabel metal1 19285 8337 19319 8371 0 FreeSans 320 0 0 0 x2.x2.x3.x8.input_stack
flabel nwell 19241 7528 19275 7588 0 FreeSans 320 0 0 0 x2.x2.x3.x8.vdd
flabel metal1 19235 8278 19281 8290 0 FreeSans 320 0 0 0 x2.x2.x3.x8.output_stack
flabel poly 19240 8998 19342 9028 0 FreeSans 320 0 0 0 x2.x2.x3.x9.input_stack
flabel metal1 19194 10021 19228 10081 0 FreeSans 320 0 0 0 x2.x2.x3.x9.vss
flabel metal1 19188 9043 19234 9055 0 FreeSans 320 0 0 0 x2.x2.x3.x9.output_stack
flabel locali 19707 8337 19741 8371 0 FreeSans 340 0 0 0 x2.x2.x3.x10.Y
flabel locali 19707 8405 19741 8439 0 FreeSans 340 0 0 0 x2.x2.x3.x10.Y
flabel locali 19799 8405 19833 8439 0 FreeSans 340 0 0 0 x2.x2.x3.x10.A
flabel metal1 19842 8643 19876 8677 0 FreeSans 200 0 0 0 x2.x2.x3.x10.VGND
flabel metal1 19842 8099 19876 8133 0 FreeSans 200 0 0 0 x2.x2.x3.x10.VPWR
rlabel comment 19905 8660 19905 8660 8 x2.x2.x3.x10.inv_1
rlabel metal1 19629 8612 19905 8708 5 x2.x2.x3.x10.VGND
rlabel metal1 19629 8068 19905 8164 5 x2.x2.x3.x10.VPWR
flabel pwell 19842 8643 19876 8677 0 FreeSans 200 0 0 0 x2.x2.x3.x10.VNB
flabel nwell 19842 8099 19876 8133 0 FreeSans 200 0 0 0 x2.x2.x3.x10.VPB
flabel locali 19609 8337 19643 8371 0 FreeSans 340 0 0 0 x2.x2.x3.x11.Y
flabel locali 19609 8405 19643 8439 0 FreeSans 340 0 0 0 x2.x2.x3.x11.Y
flabel locali 19517 8405 19551 8439 0 FreeSans 340 0 0 0 x2.x2.x3.x11.A
flabel metal1 19474 8643 19508 8677 0 FreeSans 200 0 0 0 x2.x2.x3.x11.VGND
flabel metal1 19474 8099 19508 8133 0 FreeSans 200 0 0 0 x2.x2.x3.x11.VPWR
rlabel comment 19445 8660 19445 8660 2 x2.x2.x3.x11.inv_1
rlabel metal1 19445 8612 19721 8708 5 x2.x2.x3.x11.VGND
rlabel metal1 19445 8068 19721 8164 5 x2.x2.x3.x11.VPWR
flabel pwell 19474 8643 19508 8677 0 FreeSans 200 0 0 0 x2.x2.x3.x11.VNB
flabel nwell 19474 8099 19508 8133 0 FreeSans 200 0 0 0 x2.x2.x3.x11.VPB
flabel metal1 18643 8580 18677 8614 0 FreeSans 320 0 0 0 x2.x2.x3.x6.SW
flabel nwell 18563 7484 19233 7552 0 FreeSans 320 0 0 0 x2.x2.x3.x6.VDD
flabel pdiff 18587 8661 18645 8745 0 FreeSans 320 0 0 0 x2.x2.x3.x6.delay_signal
flabel metal4 19132 7484 19233 7553 0 FreeSans 320 0 0 0 x2.x2.x3.x6.VDD
flabel via3 19068 8647 19132 8711 0 FreeSans 320 0 0 0 x2.x2.x3.x6.floating
flabel viali 18290 8981 18324 9015 0 FreeSans 320 0 0 0 x2.x2.x3.x7.SW
flabel ndiff 18234 8859 18292 8943 0 FreeSans 320 0 0 0 x2.x2.x3.x7.delay_signal
flabel metal4 18213 10052 18885 10120 0 FreeSans 320 0 0 0 x2.x2.x3.x7.VSS
flabel via3 18717 8892 18781 8956 0 FreeSans 320 0 0 0 x2.x2.x3.x7.floating
flabel viali 17558 8981 17592 9015 0 FreeSans 320 0 0 0 x2.x2.x3.x4[3].SW
flabel ndiff 17502 8859 17560 8943 0 FreeSans 320 0 0 0 x2.x2.x3.x4[3].delay_signal
flabel metal4 17481 10052 18153 10120 0 FreeSans 320 0 0 0 x2.x2.x3.x4[3].VSS
flabel via3 17985 8892 18049 8956 0 FreeSans 320 0 0 0 x2.x2.x3.x4[3].floating
flabel metal1 17785 8577 17819 8611 0 FreeSans 320 0 0 0 x2.x2.x3.x5[6].SW
flabel nwell 17229 7481 17899 7549 0 FreeSans 320 0 0 0 x2.x2.x3.x5[6].VDD
flabel pdiff 17817 8658 17875 8742 0 FreeSans 320 0 0 0 x2.x2.x3.x5[6].delay_signal
flabel metal4 17229 7481 17330 7550 0 FreeSans 320 0 0 0 x2.x2.x3.x5[6].VDD
flabel via3 17330 8644 17394 8708 0 FreeSans 320 0 0 0 x2.x2.x3.x5[6].floating
flabel metal1 17911 8577 17945 8611 0 FreeSans 320 0 0 0 x2.x2.x3.x5[7].SW
flabel nwell 17831 7481 18501 7549 0 FreeSans 320 0 0 0 x2.x2.x3.x5[7].VDD
flabel pdiff 17855 8658 17913 8742 0 FreeSans 320 0 0 0 x2.x2.x3.x5[7].delay_signal
flabel metal4 18400 7481 18501 7550 0 FreeSans 320 0 0 0 x2.x2.x3.x5[7].VDD
flabel via3 18336 8644 18400 8708 0 FreeSans 320 0 0 0 x2.x2.x3.x5[7].floating
flabel viali 17436 8981 17470 9015 0 FreeSans 320 0 0 0 x2.x2.x3.x4[2].SW
flabel ndiff 17468 8859 17526 8943 0 FreeSans 320 0 0 0 x2.x2.x3.x4[2].delay_signal
flabel metal4 16875 10052 17547 10120 0 FreeSans 320 0 0 0 x2.x2.x3.x4[2].VSS
flabel via3 16979 8892 17043 8956 0 FreeSans 320 0 0 0 x2.x2.x3.x4[2].floating
flabel metal1 16699 8577 16733 8611 0 FreeSans 320 0 0 0 x2.x2.x3.x5[5].SW
flabel nwell 16619 7481 17289 7549 0 FreeSans 320 0 0 0 x2.x2.x3.x5[5].VDD
flabel pdiff 16643 8658 16701 8742 0 FreeSans 320 0 0 0 x2.x2.x3.x5[5].delay_signal
flabel metal4 17188 7481 17289 7550 0 FreeSans 320 0 0 0 x2.x2.x3.x5[5].VDD
flabel via3 17124 8644 17188 8708 0 FreeSans 320 0 0 0 x2.x2.x3.x5[5].floating
flabel viali 16346 8981 16380 9015 0 FreeSans 320 0 0 0 x2.x2.x3.x4[1].SW
flabel ndiff 16290 8859 16348 8943 0 FreeSans 320 0 0 0 x2.x2.x3.x4[1].delay_signal
flabel metal4 16269 10052 16941 10120 0 FreeSans 320 0 0 0 x2.x2.x3.x4[1].VSS
flabel via3 16773 8892 16837 8956 0 FreeSans 320 0 0 0 x2.x2.x3.x4[1].floating
flabel metal1 16573 8577 16607 8611 0 FreeSans 320 0 0 0 x2.x2.x3.x5[4].SW
flabel nwell 16017 7481 16687 7549 0 FreeSans 320 0 0 0 x2.x2.x3.x5[4].VDD
flabel pdiff 16605 8658 16663 8742 0 FreeSans 320 0 0 0 x2.x2.x3.x5[4].delay_signal
flabel metal4 16017 7481 16118 7550 0 FreeSans 320 0 0 0 x2.x2.x3.x5[4].VDD
flabel via3 16118 8644 16182 8708 0 FreeSans 320 0 0 0 x2.x2.x3.x5[4].floating
flabel viali 16224 8981 16258 9015 0 FreeSans 320 0 0 0 x2.x2.x3.x4[0].SW
flabel ndiff 16256 8859 16314 8943 0 FreeSans 320 0 0 0 x2.x2.x3.x4[0].delay_signal
flabel metal4 15663 10052 16335 10120 0 FreeSans 320 0 0 0 x2.x2.x3.x4[0].VSS
flabel via3 15767 8892 15831 8956 0 FreeSans 320 0 0 0 x2.x2.x3.x4[0].floating
flabel metal1 15487 8577 15521 8611 0 FreeSans 320 0 0 0 x2.x2.x3.x5[3].SW
flabel nwell 15407 7481 16077 7549 0 FreeSans 320 0 0 0 x2.x2.x3.x5[3].VDD
flabel pdiff 15431 8658 15489 8742 0 FreeSans 320 0 0 0 x2.x2.x3.x5[3].delay_signal
flabel metal4 15976 7481 16077 7550 0 FreeSans 320 0 0 0 x2.x2.x3.x5[3].VDD
flabel via3 15912 8644 15976 8708 0 FreeSans 320 0 0 0 x2.x2.x3.x5[3].floating
flabel viali 15008 8981 15042 9015 0 FreeSans 320 0 0 0 x2.x2.x3.x3[1].SW
flabel ndiff 14952 8859 15010 8943 0 FreeSans 320 0 0 0 x2.x2.x3.x3[1].delay_signal
flabel metal4 14931 10052 15603 10120 0 FreeSans 320 0 0 0 x2.x2.x3.x3[1].VSS
flabel via3 15435 8892 15499 8956 0 FreeSans 320 0 0 0 x2.x2.x3.x3[1].floating
flabel metal1 15361 8577 15395 8611 0 FreeSans 320 0 0 0 x2.x2.x3.x5[2].SW
flabel nwell 14805 7481 15475 7549 0 FreeSans 320 0 0 0 x2.x2.x3.x5[2].VDD
flabel pdiff 15393 8658 15451 8742 0 FreeSans 320 0 0 0 x2.x2.x3.x5[2].delay_signal
flabel metal4 14805 7481 14906 7550 0 FreeSans 320 0 0 0 x2.x2.x3.x5[2].VDD
flabel via3 14906 8644 14970 8708 0 FreeSans 320 0 0 0 x2.x2.x3.x5[2].floating
flabel viali 14886 8981 14920 9015 0 FreeSans 320 0 0 0 x2.x2.x3.x3[0].SW
flabel ndiff 14918 8859 14976 8943 0 FreeSans 320 0 0 0 x2.x2.x3.x3[0].delay_signal
flabel metal4 14325 10052 14997 10120 0 FreeSans 320 0 0 0 x2.x2.x3.x3[0].VSS
flabel via3 14429 8892 14493 8956 0 FreeSans 320 0 0 0 x2.x2.x3.x3[0].floating
flabel metal1 14275 8577 14309 8611 0 FreeSans 320 0 0 0 x2.x2.x3.x5[1].SW
flabel nwell 14195 7481 14865 7549 0 FreeSans 320 0 0 0 x2.x2.x3.x5[1].VDD
flabel pdiff 14219 8658 14277 8742 0 FreeSans 320 0 0 0 x2.x2.x3.x5[1].delay_signal
flabel metal4 14764 7481 14865 7550 0 FreeSans 320 0 0 0 x2.x2.x3.x5[1].VDD
flabel via3 14700 8644 14764 8708 0 FreeSans 320 0 0 0 x2.x2.x3.x5[1].floating
flabel viali 14152 8981 14186 9015 0 FreeSans 320 0 0 0 x2.x2.x3.x2.SW
flabel ndiff 14184 8859 14242 8943 0 FreeSans 320 0 0 0 x2.x2.x3.x2.delay_signal
flabel metal4 13591 10052 14263 10120 0 FreeSans 320 0 0 0 x2.x2.x3.x2.VSS
flabel via3 13695 8892 13759 8956 0 FreeSans 320 0 0 0 x2.x2.x3.x2.floating
flabel metal1 14149 8577 14183 8611 0 FreeSans 320 0 0 0 x2.x2.x3.x5[0].SW
flabel nwell 13593 7481 14263 7549 0 FreeSans 320 0 0 0 x2.x2.x3.x5[0].VDD
flabel pdiff 14181 8658 14239 8742 0 FreeSans 320 0 0 0 x2.x2.x3.x5[0].delay_signal
flabel metal4 13593 7481 13694 7550 0 FreeSans 320 0 0 0 x2.x2.x3.x5[0].VDD
flabel via3 13694 8644 13758 8708 0 FreeSans 320 0 0 0 x2.x2.x3.x5[0].floating
flabel metal1 25971 8777 26639 8824 0 FreeSans 320 0 0 0 x2.x2.x2.IN
flabel metal1 19981 8780 20163 8826 0 FreeSans 320 0 0 0 x2.x2.x2.OUT
flabel metal1 26538 8407 26676 8441 0 FreeSans 320 0 0 0 x2.x2.x2.code[3]
flabel metal1 21703 8975 21761 10152 0 FreeSans 320 0 0 0 x2.x2.x2.code[1]
flabel metal1 24129 8975 24187 10152 0 FreeSans 320 0 0 0 x2.x2.x2.code[2]
flabel metal4 26152 7472 26570 8082 0 FreeSans 320 0 0 0 x2.x2.x2.VDD
flabel metal4 26166 8692 26542 10129 0 FreeSans 320 0 0 0 x2.x2.x2.VSS
flabel metal2 25776 8980 26212 9026 0 FreeSans 320 0 0 0 x2.x2.x2.code_offset
flabel metal1 20846 8972 20905 10153 0 FreeSans 320 0 0 0 x2.x2.x2.code[0]
flabel metal1 25994 8337 26028 8371 0 FreeSans 320 0 0 0 x2.x2.x2.x8.input_stack
flabel nwell 25950 7528 25984 7588 0 FreeSans 320 0 0 0 x2.x2.x2.x8.vdd
flabel metal1 25944 8278 25990 8290 0 FreeSans 320 0 0 0 x2.x2.x2.x8.output_stack
flabel poly 25949 8998 26051 9028 0 FreeSans 320 0 0 0 x2.x2.x2.x9.input_stack
flabel metal1 25903 10021 25937 10081 0 FreeSans 320 0 0 0 x2.x2.x2.x9.vss
flabel metal1 25897 9043 25943 9055 0 FreeSans 320 0 0 0 x2.x2.x2.x9.output_stack
flabel locali 26416 8337 26450 8371 0 FreeSans 340 0 0 0 x2.x2.x2.x10.Y
flabel locali 26416 8405 26450 8439 0 FreeSans 340 0 0 0 x2.x2.x2.x10.Y
flabel locali 26508 8405 26542 8439 0 FreeSans 340 0 0 0 x2.x2.x2.x10.A
flabel metal1 26551 8643 26585 8677 0 FreeSans 200 0 0 0 x2.x2.x2.x10.VGND
flabel metal1 26551 8099 26585 8133 0 FreeSans 200 0 0 0 x2.x2.x2.x10.VPWR
rlabel comment 26614 8660 26614 8660 8 x2.x2.x2.x10.inv_1
rlabel metal1 26338 8612 26614 8708 5 x2.x2.x2.x10.VGND
rlabel metal1 26338 8068 26614 8164 5 x2.x2.x2.x10.VPWR
flabel pwell 26551 8643 26585 8677 0 FreeSans 200 0 0 0 x2.x2.x2.x10.VNB
flabel nwell 26551 8099 26585 8133 0 FreeSans 200 0 0 0 x2.x2.x2.x10.VPB
flabel locali 26318 8337 26352 8371 0 FreeSans 340 0 0 0 x2.x2.x2.x11.Y
flabel locali 26318 8405 26352 8439 0 FreeSans 340 0 0 0 x2.x2.x2.x11.Y
flabel locali 26226 8405 26260 8439 0 FreeSans 340 0 0 0 x2.x2.x2.x11.A
flabel metal1 26183 8643 26217 8677 0 FreeSans 200 0 0 0 x2.x2.x2.x11.VGND
flabel metal1 26183 8099 26217 8133 0 FreeSans 200 0 0 0 x2.x2.x2.x11.VPWR
rlabel comment 26154 8660 26154 8660 2 x2.x2.x2.x11.inv_1
rlabel metal1 26154 8612 26430 8708 5 x2.x2.x2.x11.VGND
rlabel metal1 26154 8068 26430 8164 5 x2.x2.x2.x11.VPWR
flabel pwell 26183 8643 26217 8677 0 FreeSans 200 0 0 0 x2.x2.x2.x11.VNB
flabel nwell 26183 8099 26217 8133 0 FreeSans 200 0 0 0 x2.x2.x2.x11.VPB
flabel metal1 25352 8580 25386 8614 0 FreeSans 320 0 0 0 x2.x2.x2.x6.SW
flabel nwell 25272 7484 25942 7552 0 FreeSans 320 0 0 0 x2.x2.x2.x6.VDD
flabel pdiff 25296 8661 25354 8745 0 FreeSans 320 0 0 0 x2.x2.x2.x6.delay_signal
flabel metal4 25841 7484 25942 7553 0 FreeSans 320 0 0 0 x2.x2.x2.x6.VDD
flabel via3 25777 8647 25841 8711 0 FreeSans 320 0 0 0 x2.x2.x2.x6.floating
flabel viali 24999 8981 25033 9015 0 FreeSans 320 0 0 0 x2.x2.x2.x7.SW
flabel ndiff 24943 8859 25001 8943 0 FreeSans 320 0 0 0 x2.x2.x2.x7.delay_signal
flabel metal4 24922 10052 25594 10120 0 FreeSans 320 0 0 0 x2.x2.x2.x7.VSS
flabel via3 25426 8892 25490 8956 0 FreeSans 320 0 0 0 x2.x2.x2.x7.floating
flabel viali 24267 8981 24301 9015 0 FreeSans 320 0 0 0 x2.x2.x2.x4[3].SW
flabel ndiff 24211 8859 24269 8943 0 FreeSans 320 0 0 0 x2.x2.x2.x4[3].delay_signal
flabel metal4 24190 10052 24862 10120 0 FreeSans 320 0 0 0 x2.x2.x2.x4[3].VSS
flabel via3 24694 8892 24758 8956 0 FreeSans 320 0 0 0 x2.x2.x2.x4[3].floating
flabel metal1 24494 8577 24528 8611 0 FreeSans 320 0 0 0 x2.x2.x2.x5[6].SW
flabel nwell 23938 7481 24608 7549 0 FreeSans 320 0 0 0 x2.x2.x2.x5[6].VDD
flabel pdiff 24526 8658 24584 8742 0 FreeSans 320 0 0 0 x2.x2.x2.x5[6].delay_signal
flabel metal4 23938 7481 24039 7550 0 FreeSans 320 0 0 0 x2.x2.x2.x5[6].VDD
flabel via3 24039 8644 24103 8708 0 FreeSans 320 0 0 0 x2.x2.x2.x5[6].floating
flabel metal1 24620 8577 24654 8611 0 FreeSans 320 0 0 0 x2.x2.x2.x5[7].SW
flabel nwell 24540 7481 25210 7549 0 FreeSans 320 0 0 0 x2.x2.x2.x5[7].VDD
flabel pdiff 24564 8658 24622 8742 0 FreeSans 320 0 0 0 x2.x2.x2.x5[7].delay_signal
flabel metal4 25109 7481 25210 7550 0 FreeSans 320 0 0 0 x2.x2.x2.x5[7].VDD
flabel via3 25045 8644 25109 8708 0 FreeSans 320 0 0 0 x2.x2.x2.x5[7].floating
flabel viali 24145 8981 24179 9015 0 FreeSans 320 0 0 0 x2.x2.x2.x4[2].SW
flabel ndiff 24177 8859 24235 8943 0 FreeSans 320 0 0 0 x2.x2.x2.x4[2].delay_signal
flabel metal4 23584 10052 24256 10120 0 FreeSans 320 0 0 0 x2.x2.x2.x4[2].VSS
flabel via3 23688 8892 23752 8956 0 FreeSans 320 0 0 0 x2.x2.x2.x4[2].floating
flabel metal1 23408 8577 23442 8611 0 FreeSans 320 0 0 0 x2.x2.x2.x5[5].SW
flabel nwell 23328 7481 23998 7549 0 FreeSans 320 0 0 0 x2.x2.x2.x5[5].VDD
flabel pdiff 23352 8658 23410 8742 0 FreeSans 320 0 0 0 x2.x2.x2.x5[5].delay_signal
flabel metal4 23897 7481 23998 7550 0 FreeSans 320 0 0 0 x2.x2.x2.x5[5].VDD
flabel via3 23833 8644 23897 8708 0 FreeSans 320 0 0 0 x2.x2.x2.x5[5].floating
flabel viali 23055 8981 23089 9015 0 FreeSans 320 0 0 0 x2.x2.x2.x4[1].SW
flabel ndiff 22999 8859 23057 8943 0 FreeSans 320 0 0 0 x2.x2.x2.x4[1].delay_signal
flabel metal4 22978 10052 23650 10120 0 FreeSans 320 0 0 0 x2.x2.x2.x4[1].VSS
flabel via3 23482 8892 23546 8956 0 FreeSans 320 0 0 0 x2.x2.x2.x4[1].floating
flabel metal1 23282 8577 23316 8611 0 FreeSans 320 0 0 0 x2.x2.x2.x5[4].SW
flabel nwell 22726 7481 23396 7549 0 FreeSans 320 0 0 0 x2.x2.x2.x5[4].VDD
flabel pdiff 23314 8658 23372 8742 0 FreeSans 320 0 0 0 x2.x2.x2.x5[4].delay_signal
flabel metal4 22726 7481 22827 7550 0 FreeSans 320 0 0 0 x2.x2.x2.x5[4].VDD
flabel via3 22827 8644 22891 8708 0 FreeSans 320 0 0 0 x2.x2.x2.x5[4].floating
flabel viali 22933 8981 22967 9015 0 FreeSans 320 0 0 0 x2.x2.x2.x4[0].SW
flabel ndiff 22965 8859 23023 8943 0 FreeSans 320 0 0 0 x2.x2.x2.x4[0].delay_signal
flabel metal4 22372 10052 23044 10120 0 FreeSans 320 0 0 0 x2.x2.x2.x4[0].VSS
flabel via3 22476 8892 22540 8956 0 FreeSans 320 0 0 0 x2.x2.x2.x4[0].floating
flabel metal1 22196 8577 22230 8611 0 FreeSans 320 0 0 0 x2.x2.x2.x5[3].SW
flabel nwell 22116 7481 22786 7549 0 FreeSans 320 0 0 0 x2.x2.x2.x5[3].VDD
flabel pdiff 22140 8658 22198 8742 0 FreeSans 320 0 0 0 x2.x2.x2.x5[3].delay_signal
flabel metal4 22685 7481 22786 7550 0 FreeSans 320 0 0 0 x2.x2.x2.x5[3].VDD
flabel via3 22621 8644 22685 8708 0 FreeSans 320 0 0 0 x2.x2.x2.x5[3].floating
flabel viali 21717 8981 21751 9015 0 FreeSans 320 0 0 0 x2.x2.x2.x3[1].SW
flabel ndiff 21661 8859 21719 8943 0 FreeSans 320 0 0 0 x2.x2.x2.x3[1].delay_signal
flabel metal4 21640 10052 22312 10120 0 FreeSans 320 0 0 0 x2.x2.x2.x3[1].VSS
flabel via3 22144 8892 22208 8956 0 FreeSans 320 0 0 0 x2.x2.x2.x3[1].floating
flabel metal1 22070 8577 22104 8611 0 FreeSans 320 0 0 0 x2.x2.x2.x5[2].SW
flabel nwell 21514 7481 22184 7549 0 FreeSans 320 0 0 0 x2.x2.x2.x5[2].VDD
flabel pdiff 22102 8658 22160 8742 0 FreeSans 320 0 0 0 x2.x2.x2.x5[2].delay_signal
flabel metal4 21514 7481 21615 7550 0 FreeSans 320 0 0 0 x2.x2.x2.x5[2].VDD
flabel via3 21615 8644 21679 8708 0 FreeSans 320 0 0 0 x2.x2.x2.x5[2].floating
flabel viali 21595 8981 21629 9015 0 FreeSans 320 0 0 0 x2.x2.x2.x3[0].SW
flabel ndiff 21627 8859 21685 8943 0 FreeSans 320 0 0 0 x2.x2.x2.x3[0].delay_signal
flabel metal4 21034 10052 21706 10120 0 FreeSans 320 0 0 0 x2.x2.x2.x3[0].VSS
flabel via3 21138 8892 21202 8956 0 FreeSans 320 0 0 0 x2.x2.x2.x3[0].floating
flabel metal1 20984 8577 21018 8611 0 FreeSans 320 0 0 0 x2.x2.x2.x5[1].SW
flabel nwell 20904 7481 21574 7549 0 FreeSans 320 0 0 0 x2.x2.x2.x5[1].VDD
flabel pdiff 20928 8658 20986 8742 0 FreeSans 320 0 0 0 x2.x2.x2.x5[1].delay_signal
flabel metal4 21473 7481 21574 7550 0 FreeSans 320 0 0 0 x2.x2.x2.x5[1].VDD
flabel via3 21409 8644 21473 8708 0 FreeSans 320 0 0 0 x2.x2.x2.x5[1].floating
flabel viali 20861 8981 20895 9015 0 FreeSans 320 0 0 0 x2.x2.x2.x2.SW
flabel ndiff 20893 8859 20951 8943 0 FreeSans 320 0 0 0 x2.x2.x2.x2.delay_signal
flabel metal4 20300 10052 20972 10120 0 FreeSans 320 0 0 0 x2.x2.x2.x2.VSS
flabel via3 20404 8892 20468 8956 0 FreeSans 320 0 0 0 x2.x2.x2.x2.floating
flabel metal1 20858 8577 20892 8611 0 FreeSans 320 0 0 0 x2.x2.x2.x5[0].SW
flabel nwell 20302 7481 20972 7549 0 FreeSans 320 0 0 0 x2.x2.x2.x5[0].VDD
flabel pdiff 20890 8658 20948 8742 0 FreeSans 320 0 0 0 x2.x2.x2.x5[0].delay_signal
flabel metal4 20302 7481 20403 7550 0 FreeSans 320 0 0 0 x2.x2.x2.x5[0].VDD
flabel via3 20403 8644 20467 8708 0 FreeSans 320 0 0 0 x2.x2.x2.x5[0].floating
flabel metal1 19958 12285 20626 12332 0 FreeSans 320 0 0 0 x2.x2.x1.IN
flabel metal1 26434 12283 26616 12329 0 FreeSans 320 0 0 0 x2.x2.x1.OUT
flabel metal1 19921 12668 20059 12702 0 FreeSans 320 0 0 0 x2.x2.x1.code[3]
flabel metal1 24836 10957 24894 12134 0 FreeSans 320 0 0 0 x2.x2.x1.code[1]
flabel metal1 22410 10957 22468 12134 0 FreeSans 320 0 0 0 x2.x2.x1.code[2]
flabel metal4 20027 13027 20445 13637 0 FreeSans 320 0 0 0 x2.x2.x1.VDD
flabel metal4 20055 10980 20431 12417 0 FreeSans 320 0 0 0 x2.x2.x1.VSS
flabel metal2 20385 12083 20821 12129 0 FreeSans 320 0 0 0 x2.x2.x1.code_offset
flabel metal1 25692 10956 25751 12137 0 FreeSans 320 0 0 0 x2.x2.x1.code[0]
flabel metal1 20569 12738 20603 12772 0 FreeSans 320 0 0 0 x2.x2.x1.x8.input_stack
flabel nwell 20613 13521 20647 13581 0 FreeSans 320 0 0 0 x2.x2.x1.x8.vdd
flabel metal1 20607 12819 20653 12831 0 FreeSans 320 0 0 0 x2.x2.x1.x8.output_stack
flabel poly 20546 12081 20648 12111 0 FreeSans 320 0 0 0 x2.x2.x1.x9.input_stack
flabel metal1 20660 11028 20694 11088 0 FreeSans 320 0 0 0 x2.x2.x1.x9.vss
flabel metal1 20654 12054 20700 12066 0 FreeSans 320 0 0 0 x2.x2.x1.x9.output_stack
flabel locali 20147 12738 20181 12772 0 FreeSans 340 0 0 0 x2.x2.x1.x10.Y
flabel locali 20147 12670 20181 12704 0 FreeSans 340 0 0 0 x2.x2.x1.x10.Y
flabel locali 20055 12670 20089 12704 0 FreeSans 340 0 0 0 x2.x2.x1.x10.A
flabel metal1 20012 12432 20046 12466 0 FreeSans 200 0 0 0 x2.x2.x1.x10.VGND
flabel metal1 20012 12976 20046 13010 0 FreeSans 200 0 0 0 x2.x2.x1.x10.VPWR
rlabel comment 19983 12449 19983 12449 4 x2.x2.x1.x10.inv_1
rlabel metal1 19983 12401 20259 12497 1 x2.x2.x1.x10.VGND
rlabel metal1 19983 12945 20259 13041 1 x2.x2.x1.x10.VPWR
flabel pwell 20012 12432 20046 12466 0 FreeSans 200 0 0 0 x2.x2.x1.x10.VNB
flabel nwell 20012 12976 20046 13010 0 FreeSans 200 0 0 0 x2.x2.x1.x10.VPB
flabel locali 20245 12738 20279 12772 0 FreeSans 340 0 0 0 x2.x2.x1.x11.Y
flabel locali 20245 12670 20279 12704 0 FreeSans 340 0 0 0 x2.x2.x1.x11.Y
flabel locali 20337 12670 20371 12704 0 FreeSans 340 0 0 0 x2.x2.x1.x11.A
flabel metal1 20380 12432 20414 12466 0 FreeSans 200 0 0 0 x2.x2.x1.x11.VGND
flabel metal1 20380 12976 20414 13010 0 FreeSans 200 0 0 0 x2.x2.x1.x11.VPWR
rlabel comment 20443 12449 20443 12449 6 x2.x2.x1.x11.inv_1
rlabel metal1 20167 12401 20443 12497 1 x2.x2.x1.x11.VGND
rlabel metal1 20167 12945 20443 13041 1 x2.x2.x1.x11.VPWR
flabel pwell 20380 12432 20414 12466 0 FreeSans 200 0 0 0 x2.x2.x1.x11.VNB
flabel nwell 20380 12976 20414 13010 0 FreeSans 200 0 0 0 x2.x2.x1.x11.VPB
flabel metal1 21211 12495 21245 12529 0 FreeSans 320 0 0 0 x2.x2.x1.x6.SW
flabel nwell 20655 13557 21325 13625 0 FreeSans 320 0 0 0 x2.x2.x1.x6.VDD
flabel pdiff 21243 12364 21301 12448 0 FreeSans 320 0 0 0 x2.x2.x1.x6.delay_signal
flabel metal4 20655 13556 20756 13625 0 FreeSans 320 0 0 0 x2.x2.x1.x6.VDD
flabel via3 20756 12398 20820 12462 0 FreeSans 320 0 0 0 x2.x2.x1.x6.floating
flabel viali 21564 12094 21598 12128 0 FreeSans 320 0 0 0 x2.x2.x1.x7.SW
flabel ndiff 21596 12166 21654 12250 0 FreeSans 320 0 0 0 x2.x2.x1.x7.delay_signal
flabel metal4 21003 10989 21675 11057 0 FreeSans 320 0 0 0 x2.x2.x1.x7.VSS
flabel via3 21107 12153 21171 12217 0 FreeSans 320 0 0 0 x2.x2.x1.x7.floating
flabel viali 22296 12094 22330 12128 0 FreeSans 320 0 0 0 x2.x2.x1.x4[3].SW
flabel ndiff 22328 12166 22386 12250 0 FreeSans 320 0 0 0 x2.x2.x1.x4[3].delay_signal
flabel metal4 21735 10989 22407 11057 0 FreeSans 320 0 0 0 x2.x2.x1.x4[3].VSS
flabel via3 21839 12153 21903 12217 0 FreeSans 320 0 0 0 x2.x2.x1.x4[3].floating
flabel metal1 22069 12498 22103 12532 0 FreeSans 320 0 0 0 x2.x2.x1.x5[6].SW
flabel nwell 21989 13560 22659 13628 0 FreeSans 320 0 0 0 x2.x2.x1.x5[6].VDD
flabel pdiff 22013 12367 22071 12451 0 FreeSans 320 0 0 0 x2.x2.x1.x5[6].delay_signal
flabel metal4 22558 13559 22659 13628 0 FreeSans 320 0 0 0 x2.x2.x1.x5[6].VDD
flabel via3 22494 12401 22558 12465 0 FreeSans 320 0 0 0 x2.x2.x1.x5[6].floating
flabel metal1 21943 12498 21977 12532 0 FreeSans 320 0 0 0 x2.x2.x1.x5[7].SW
flabel nwell 21387 13560 22057 13628 0 FreeSans 320 0 0 0 x2.x2.x1.x5[7].VDD
flabel pdiff 21975 12367 22033 12451 0 FreeSans 320 0 0 0 x2.x2.x1.x5[7].delay_signal
flabel metal4 21387 13559 21488 13628 0 FreeSans 320 0 0 0 x2.x2.x1.x5[7].VDD
flabel via3 21488 12401 21552 12465 0 FreeSans 320 0 0 0 x2.x2.x1.x5[7].floating
flabel viali 22418 12094 22452 12128 0 FreeSans 320 0 0 0 x2.x2.x1.x4[2].SW
flabel ndiff 22362 12166 22420 12250 0 FreeSans 320 0 0 0 x2.x2.x1.x4[2].delay_signal
flabel metal4 22341 10989 23013 11057 0 FreeSans 320 0 0 0 x2.x2.x1.x4[2].VSS
flabel via3 22845 12153 22909 12217 0 FreeSans 320 0 0 0 x2.x2.x1.x4[2].floating
flabel metal1 23155 12498 23189 12532 0 FreeSans 320 0 0 0 x2.x2.x1.x5[5].SW
flabel nwell 22599 13560 23269 13628 0 FreeSans 320 0 0 0 x2.x2.x1.x5[5].VDD
flabel pdiff 23187 12367 23245 12451 0 FreeSans 320 0 0 0 x2.x2.x1.x5[5].delay_signal
flabel metal4 22599 13559 22700 13628 0 FreeSans 320 0 0 0 x2.x2.x1.x5[5].VDD
flabel via3 22700 12401 22764 12465 0 FreeSans 320 0 0 0 x2.x2.x1.x5[5].floating
flabel viali 23508 12094 23542 12128 0 FreeSans 320 0 0 0 x2.x2.x1.x4[1].SW
flabel ndiff 23540 12166 23598 12250 0 FreeSans 320 0 0 0 x2.x2.x1.x4[1].delay_signal
flabel metal4 22947 10989 23619 11057 0 FreeSans 320 0 0 0 x2.x2.x1.x4[1].VSS
flabel via3 23051 12153 23115 12217 0 FreeSans 320 0 0 0 x2.x2.x1.x4[1].floating
flabel metal1 23281 12498 23315 12532 0 FreeSans 320 0 0 0 x2.x2.x1.x5[4].SW
flabel nwell 23201 13560 23871 13628 0 FreeSans 320 0 0 0 x2.x2.x1.x5[4].VDD
flabel pdiff 23225 12367 23283 12451 0 FreeSans 320 0 0 0 x2.x2.x1.x5[4].delay_signal
flabel metal4 23770 13559 23871 13628 0 FreeSans 320 0 0 0 x2.x2.x1.x5[4].VDD
flabel via3 23706 12401 23770 12465 0 FreeSans 320 0 0 0 x2.x2.x1.x5[4].floating
flabel viali 23630 12094 23664 12128 0 FreeSans 320 0 0 0 x2.x2.x1.x4[0].SW
flabel ndiff 23574 12166 23632 12250 0 FreeSans 320 0 0 0 x2.x2.x1.x4[0].delay_signal
flabel metal4 23553 10989 24225 11057 0 FreeSans 320 0 0 0 x2.x2.x1.x4[0].VSS
flabel via3 24057 12153 24121 12217 0 FreeSans 320 0 0 0 x2.x2.x1.x4[0].floating
flabel metal1 24367 12498 24401 12532 0 FreeSans 320 0 0 0 x2.x2.x1.x5[3].SW
flabel nwell 23811 13560 24481 13628 0 FreeSans 320 0 0 0 x2.x2.x1.x5[3].VDD
flabel pdiff 24399 12367 24457 12451 0 FreeSans 320 0 0 0 x2.x2.x1.x5[3].delay_signal
flabel metal4 23811 13559 23912 13628 0 FreeSans 320 0 0 0 x2.x2.x1.x5[3].VDD
flabel via3 23912 12401 23976 12465 0 FreeSans 320 0 0 0 x2.x2.x1.x5[3].floating
flabel viali 24846 12094 24880 12128 0 FreeSans 320 0 0 0 x2.x2.x1.x3[1].SW
flabel ndiff 24878 12166 24936 12250 0 FreeSans 320 0 0 0 x2.x2.x1.x3[1].delay_signal
flabel metal4 24285 10989 24957 11057 0 FreeSans 320 0 0 0 x2.x2.x1.x3[1].VSS
flabel via3 24389 12153 24453 12217 0 FreeSans 320 0 0 0 x2.x2.x1.x3[1].floating
flabel metal1 24493 12498 24527 12532 0 FreeSans 320 0 0 0 x2.x2.x1.x5[2].SW
flabel nwell 24413 13560 25083 13628 0 FreeSans 320 0 0 0 x2.x2.x1.x5[2].VDD
flabel pdiff 24437 12367 24495 12451 0 FreeSans 320 0 0 0 x2.x2.x1.x5[2].delay_signal
flabel metal4 24982 13559 25083 13628 0 FreeSans 320 0 0 0 x2.x2.x1.x5[2].VDD
flabel via3 24918 12401 24982 12465 0 FreeSans 320 0 0 0 x2.x2.x1.x5[2].floating
flabel viali 24968 12094 25002 12128 0 FreeSans 320 0 0 0 x2.x2.x1.x3[0].SW
flabel ndiff 24912 12166 24970 12250 0 FreeSans 320 0 0 0 x2.x2.x1.x3[0].delay_signal
flabel metal4 24891 10989 25563 11057 0 FreeSans 320 0 0 0 x2.x2.x1.x3[0].VSS
flabel via3 25395 12153 25459 12217 0 FreeSans 320 0 0 0 x2.x2.x1.x3[0].floating
flabel metal1 25579 12498 25613 12532 0 FreeSans 320 0 0 0 x2.x2.x1.x5[1].SW
flabel nwell 25023 13560 25693 13628 0 FreeSans 320 0 0 0 x2.x2.x1.x5[1].VDD
flabel pdiff 25611 12367 25669 12451 0 FreeSans 320 0 0 0 x2.x2.x1.x5[1].delay_signal
flabel metal4 25023 13559 25124 13628 0 FreeSans 320 0 0 0 x2.x2.x1.x5[1].VDD
flabel via3 25124 12401 25188 12465 0 FreeSans 320 0 0 0 x2.x2.x1.x5[1].floating
flabel viali 25702 12094 25736 12128 0 FreeSans 320 0 0 0 x2.x2.x1.x2.SW
flabel ndiff 25646 12166 25704 12250 0 FreeSans 320 0 0 0 x2.x2.x1.x2.delay_signal
flabel metal4 25625 10989 26297 11057 0 FreeSans 320 0 0 0 x2.x2.x1.x2.VSS
flabel via3 26129 12153 26193 12217 0 FreeSans 320 0 0 0 x2.x2.x1.x2.floating
flabel metal1 25705 12498 25739 12532 0 FreeSans 320 0 0 0 x2.x2.x1.x5[0].SW
flabel nwell 25625 13560 26295 13628 0 FreeSans 320 0 0 0 x2.x2.x1.x5[0].VDD
flabel pdiff 25649 12367 25707 12451 0 FreeSans 320 0 0 0 x2.x2.x1.x5[0].delay_signal
flabel metal4 26194 13559 26295 13628 0 FreeSans 320 0 0 0 x2.x2.x1.x5[0].VDD
flabel via3 26130 12401 26194 12465 0 FreeSans 320 0 0 0 x2.x2.x1.x5[0].floating
flabel metal2 11556 7587 11590 7616 0 FreeSans 320 0 0 0 x1.sample_clk
flabel metal2 10746 9426 10780 9459 0 FreeSans 320 0 0 0 x1.eob
flabel metal2 2737 9000 2790 11540 0 FreeSans 320 0 0 0 x1.delay_offset
flabel metal1 3038 7367 9995 7401 0 FreeSans 320 0 0 0 x1.async_clk_sar
flabel metal4 2458 10123 2570 10430 0 FreeSans 320 0 0 0 x1.vss
flabel metal4 2064 7484 2370 13066 0 FreeSans 320 0 0 0 x1.vdd
flabel metal1 2330 11810 2375 11857 0 FreeSans 320 0 0 0 x1.ready
flabel metal1 2930 10169 4871 10197 0 FreeSans 320 0 0 0 x1.async_resetb_delay_ctrl_code[2]
flabel metal1 2932 10225 7297 10253 0 FreeSans 320 0 0 0 x1.async_resetb_delay_ctrl_code[1]
flabel metal1 2928 10281 8154 10309 0 FreeSans 320 0 0 0 x1.async_resetb_delay_ctrl_code[0]
flabel metal1 2324 8419 2366 8453 0 FreeSans 320 0 0 0 x1.async_resetb_delay_ctrl_code[3]
flabel metal1 2324 12193 2356 12227 0 FreeSans 320 0 0 0 x1.async_setb_delay_ctrl_code[3]
flabel metal1 2929 10337 8154 10365 0 FreeSans 320 0 0 0 x1.async_setb_delay_ctrl_code[0]
flabel metal1 2931 10393 7297 10421 0 FreeSans 320 0 0 0 x1.async_setb_delay_ctrl_code[1]
flabel metal1 2930 10449 4871 10477 0 FreeSans 320 0 0 0 x1.async_setb_delay_ctrl_code[2]
flabel locali 9771 8786 9846 8832 0 FreeSans 400 0 0 0 x1.x27.RESET_B
flabel locali 11645 9034 11679 9068 7 FreeSans 400 0 0 0 x1.x27.VGND
flabel locali 11645 8796 11679 8830 0 FreeSans 400 0 0 0 x1.x27.CLK
flabel locali 11645 8728 11679 8762 0 FreeSans 400 0 0 0 x1.x27.CLK
flabel locali 10909 8864 10943 8898 0 FreeSans 400 0 0 0 x1.x27.SET_B
flabel locali 9347 8932 9381 8966 0 FreeSans 400 0 0 0 x1.x27.Q
flabel locali 9347 8660 9381 8694 0 FreeSans 400 0 0 0 x1.x27.Q
flabel locali 9347 8592 9381 8626 0 FreeSans 400 0 0 0 x1.x27.Q
flabel locali 11645 8490 11679 8524 7 FreeSans 400 0 0 0 x1.x27.VPWR
flabel locali 11277 8796 11311 8830 0 FreeSans 200 0 0 0 x1.x27.D
flabel locali 11277 8728 11311 8762 0 FreeSans 200 0 0 0 x1.x27.D
flabel locali 9627 8592 9661 8626 0 FreeSans 400 0 0 0 x1.x27.Q_N
flabel locali 9627 8660 9661 8694 0 FreeSans 400 0 0 0 x1.x27.Q_N
flabel locali 9627 8932 9661 8966 0 FreeSans 400 0 0 0 x1.x27.Q_N
flabel metal1 11645 9034 11679 9068 0 FreeSans 200 0 0 0 x1.x27.VGND
flabel metal1 11645 8490 11679 8524 0 FreeSans 200 0 0 0 x1.x27.VPWR
flabel nwell 11645 8490 11679 8524 7 FreeSans 400 0 0 0 x1.x27.VPB
flabel nwell 11662 8507 11662 8507 0 FreeSans 200 0 0 0 x1.x27.VPB
flabel pwell 11645 9034 11679 9068 7 FreeSans 400 0 0 0 x1.x27.VNB
flabel pwell 11662 9051 11662 9051 0 FreeSans 200 0 0 0 x1.x27.VNB
rlabel comment 11709 9051 11709 9051 8 x1.x27.dfbbp_1
rlabel locali 10142 8838 10217 8904 5 x1.x27.SET_B
rlabel metal1 10161 8858 10219 8867 5 x1.x27.SET_B
rlabel metal1 10161 8895 10219 8904 5 x1.x27.SET_B
rlabel metal1 10897 8858 10955 8867 5 x1.x27.SET_B
rlabel metal1 10161 8867 10955 8895 5 x1.x27.SET_B
rlabel metal1 10897 8895 10955 8904 5 x1.x27.SET_B
rlabel metal1 9317 9003 11709 9099 5 x1.x27.VGND
rlabel metal1 9317 8459 11709 8555 5 x1.x27.VPWR
flabel locali 9225 8728 9259 8762 0 FreeSans 340 0 0 0 x1.x10.Y
flabel locali 9225 8796 9259 8830 0 FreeSans 340 0 0 0 x1.x10.Y
flabel locali 9133 8796 9167 8830 0 FreeSans 340 0 0 0 x1.x10.A
flabel metal1 9090 9034 9124 9068 0 FreeSans 200 0 0 0 x1.x10.VGND
flabel metal1 9090 8490 9124 8524 0 FreeSans 200 0 0 0 x1.x10.VPWR
rlabel comment 9061 9051 9061 9051 2 x1.x10.inv_1
rlabel metal1 9061 9003 9337 9099 5 x1.x10.VGND
rlabel metal1 9061 8459 9337 8555 5 x1.x10.VPWR
flabel pwell 9090 9034 9124 9068 0 FreeSans 200 0 0 0 x1.x10.VNB
flabel nwell 9090 8490 9124 8524 0 FreeSans 200 0 0 0 x1.x10.VPB
flabel locali 9225 11886 9259 11920 0 FreeSans 340 0 0 0 x1.x9.Y
flabel locali 9225 11818 9259 11852 0 FreeSans 340 0 0 0 x1.x9.Y
flabel locali 9133 11818 9167 11852 0 FreeSans 340 0 0 0 x1.x9.A
flabel metal1 9090 11580 9124 11614 0 FreeSans 200 0 0 0 x1.x9.VGND
flabel metal1 9090 12124 9124 12158 0 FreeSans 200 0 0 0 x1.x9.VPWR
rlabel comment 9061 11597 9061 11597 4 x1.x9.inv_1
rlabel metal1 9061 11549 9337 11645 1 x1.x9.VGND
rlabel metal1 9061 12093 9337 12189 1 x1.x9.VPWR
flabel pwell 9090 11580 9124 11614 0 FreeSans 200 0 0 0 x1.x9.VNB
flabel nwell 9090 12124 9124 12158 0 FreeSans 200 0 0 0 x1.x9.VPB
flabel metal1 10084 7771 10118 7805 0 FreeSans 200 0 0 0 x1.x8.VGND
flabel metal1 10084 8315 10118 8349 0 FreeSans 200 0 0 0 x1.x8.VPWR
flabel locali 10728 8077 10762 8111 0 FreeSans 250 0 0 0 x1.x8.S
flabel locali 10636 8077 10670 8111 0 FreeSans 250 0 0 0 x1.x8.S
flabel locali 10544 7941 10578 7975 0 FreeSans 250 0 0 0 x1.x8.A1
flabel locali 10544 8009 10578 8043 0 FreeSans 250 0 0 0 x1.x8.A1
flabel locali 10452 8009 10486 8043 0 FreeSans 250 0 0 0 x1.x8.A0
flabel locali 10084 7873 10118 7907 0 FreeSans 250 0 0 0 x1.x8.X
flabel locali 10084 8145 10118 8179 0 FreeSans 250 0 0 0 x1.x8.X
flabel locali 10084 8213 10118 8247 0 FreeSans 250 0 0 0 x1.x8.X
flabel nwell 10128 8315 10162 8349 0 FreeSans 250 0 0 0 x1.x8.VPB
flabel pwell 10138 7771 10172 7805 0 FreeSans 250 0 0 0 x1.x8.VNB
rlabel comment 10054 7788 10054 7788 4 x1.x8.mux2_1
rlabel metal1 10054 7740 10882 7836 1 x1.x8.VGND
rlabel metal1 10054 8284 10882 8380 1 x1.x8.VPWR
flabel metal1 2361 8789 3029 8836 0 FreeSans 320 0 0 0 x1.x4.IN
flabel metal1 8837 8792 9019 8838 0 FreeSans 320 0 0 0 x1.x4.OUT
flabel metal1 2324 8419 2462 8453 0 FreeSans 320 0 0 0 x1.x4.code[3]
flabel metal1 7239 8987 7297 10164 0 FreeSans 320 0 0 0 x1.x4.code[1]
flabel metal1 4813 8987 4871 10164 0 FreeSans 320 0 0 0 x1.x4.code[2]
flabel metal4 2430 7484 2848 8094 0 FreeSans 320 0 0 0 x1.x4.VDD
flabel metal4 2458 8704 2834 10141 0 FreeSans 320 0 0 0 x1.x4.VSS
flabel metal2 2788 8992 3224 9038 0 FreeSans 320 0 0 0 x1.x4.code_offset
flabel metal1 8095 8984 8154 10165 0 FreeSans 320 0 0 0 x1.x4.code[0]
flabel metal1 2972 8349 3006 8383 0 FreeSans 320 0 0 0 x1.x4.x8.input_stack
flabel nwell 3016 7540 3050 7600 0 FreeSans 320 0 0 0 x1.x4.x8.vdd
flabel metal1 3010 8290 3056 8302 0 FreeSans 320 0 0 0 x1.x4.x8.output_stack
flabel poly 2949 9010 3051 9040 0 FreeSans 320 0 0 0 x1.x4.x9.input_stack
flabel metal1 3063 10033 3097 10093 0 FreeSans 320 0 0 0 x1.x4.x9.vss
flabel metal1 3057 9055 3103 9067 0 FreeSans 320 0 0 0 x1.x4.x9.output_stack
flabel locali 2550 8349 2584 8383 0 FreeSans 340 0 0 0 x1.x4.x10.Y
flabel locali 2550 8417 2584 8451 0 FreeSans 340 0 0 0 x1.x4.x10.Y
flabel locali 2458 8417 2492 8451 0 FreeSans 340 0 0 0 x1.x4.x10.A
flabel metal1 2415 8655 2449 8689 0 FreeSans 200 0 0 0 x1.x4.x10.VGND
flabel metal1 2415 8111 2449 8145 0 FreeSans 200 0 0 0 x1.x4.x10.VPWR
rlabel comment 2386 8672 2386 8672 2 x1.x4.x10.inv_1
rlabel metal1 2386 8624 2662 8720 5 x1.x4.x10.VGND
rlabel metal1 2386 8080 2662 8176 5 x1.x4.x10.VPWR
flabel pwell 2415 8655 2449 8689 0 FreeSans 200 0 0 0 x1.x4.x10.VNB
flabel nwell 2415 8111 2449 8145 0 FreeSans 200 0 0 0 x1.x4.x10.VPB
flabel locali 2648 8349 2682 8383 0 FreeSans 340 0 0 0 x1.x4.x11.Y
flabel locali 2648 8417 2682 8451 0 FreeSans 340 0 0 0 x1.x4.x11.Y
flabel locali 2740 8417 2774 8451 0 FreeSans 340 0 0 0 x1.x4.x11.A
flabel metal1 2783 8655 2817 8689 0 FreeSans 200 0 0 0 x1.x4.x11.VGND
flabel metal1 2783 8111 2817 8145 0 FreeSans 200 0 0 0 x1.x4.x11.VPWR
rlabel comment 2846 8672 2846 8672 8 x1.x4.x11.inv_1
rlabel metal1 2570 8624 2846 8720 5 x1.x4.x11.VGND
rlabel metal1 2570 8080 2846 8176 5 x1.x4.x11.VPWR
flabel pwell 2783 8655 2817 8689 0 FreeSans 200 0 0 0 x1.x4.x11.VNB
flabel nwell 2783 8111 2817 8145 0 FreeSans 200 0 0 0 x1.x4.x11.VPB
flabel metal1 3614 8592 3648 8626 0 FreeSans 320 0 0 0 x1.x4.x6.SW
flabel nwell 3058 7496 3728 7564 0 FreeSans 320 0 0 0 x1.x4.x6.VDD
flabel pdiff 3646 8673 3704 8757 0 FreeSans 320 0 0 0 x1.x4.x6.delay_signal
flabel metal4 3058 7496 3159 7565 0 FreeSans 320 0 0 0 x1.x4.x6.VDD
flabel via3 3159 8659 3223 8723 0 FreeSans 320 0 0 0 x1.x4.x6.floating
flabel viali 3967 8993 4001 9027 0 FreeSans 320 0 0 0 x1.x4.x7.SW
flabel ndiff 3999 8871 4057 8955 0 FreeSans 320 0 0 0 x1.x4.x7.delay_signal
flabel metal4 3406 10064 4078 10132 0 FreeSans 320 0 0 0 x1.x4.x7.VSS
flabel via3 3510 8904 3574 8968 0 FreeSans 320 0 0 0 x1.x4.x7.floating
flabel viali 4699 8993 4733 9027 0 FreeSans 320 0 0 0 x1.x4.x4[3].SW
flabel ndiff 4731 8871 4789 8955 0 FreeSans 320 0 0 0 x1.x4.x4[3].delay_signal
flabel metal4 4138 10064 4810 10132 0 FreeSans 320 0 0 0 x1.x4.x4[3].VSS
flabel via3 4242 8904 4306 8968 0 FreeSans 320 0 0 0 x1.x4.x4[3].floating
flabel metal1 4472 8589 4506 8623 0 FreeSans 320 0 0 0 x1.x4.x5[6].SW
flabel nwell 4392 7493 5062 7561 0 FreeSans 320 0 0 0 x1.x4.x5[6].VDD
flabel pdiff 4416 8670 4474 8754 0 FreeSans 320 0 0 0 x1.x4.x5[6].delay_signal
flabel metal4 4961 7493 5062 7562 0 FreeSans 320 0 0 0 x1.x4.x5[6].VDD
flabel via3 4897 8656 4961 8720 0 FreeSans 320 0 0 0 x1.x4.x5[6].floating
flabel metal1 4346 8589 4380 8623 0 FreeSans 320 0 0 0 x1.x4.x5[7].SW
flabel nwell 3790 7493 4460 7561 0 FreeSans 320 0 0 0 x1.x4.x5[7].VDD
flabel pdiff 4378 8670 4436 8754 0 FreeSans 320 0 0 0 x1.x4.x5[7].delay_signal
flabel metal4 3790 7493 3891 7562 0 FreeSans 320 0 0 0 x1.x4.x5[7].VDD
flabel via3 3891 8656 3955 8720 0 FreeSans 320 0 0 0 x1.x4.x5[7].floating
flabel viali 4821 8993 4855 9027 0 FreeSans 320 0 0 0 x1.x4.x4[2].SW
flabel ndiff 4765 8871 4823 8955 0 FreeSans 320 0 0 0 x1.x4.x4[2].delay_signal
flabel metal4 4744 10064 5416 10132 0 FreeSans 320 0 0 0 x1.x4.x4[2].VSS
flabel via3 5248 8904 5312 8968 0 FreeSans 320 0 0 0 x1.x4.x4[2].floating
flabel metal1 5558 8589 5592 8623 0 FreeSans 320 0 0 0 x1.x4.x5[5].SW
flabel nwell 5002 7493 5672 7561 0 FreeSans 320 0 0 0 x1.x4.x5[5].VDD
flabel pdiff 5590 8670 5648 8754 0 FreeSans 320 0 0 0 x1.x4.x5[5].delay_signal
flabel metal4 5002 7493 5103 7562 0 FreeSans 320 0 0 0 x1.x4.x5[5].VDD
flabel via3 5103 8656 5167 8720 0 FreeSans 320 0 0 0 x1.x4.x5[5].floating
flabel viali 5911 8993 5945 9027 0 FreeSans 320 0 0 0 x1.x4.x4[1].SW
flabel ndiff 5943 8871 6001 8955 0 FreeSans 320 0 0 0 x1.x4.x4[1].delay_signal
flabel metal4 5350 10064 6022 10132 0 FreeSans 320 0 0 0 x1.x4.x4[1].VSS
flabel via3 5454 8904 5518 8968 0 FreeSans 320 0 0 0 x1.x4.x4[1].floating
flabel metal1 5684 8589 5718 8623 0 FreeSans 320 0 0 0 x1.x4.x5[4].SW
flabel nwell 5604 7493 6274 7561 0 FreeSans 320 0 0 0 x1.x4.x5[4].VDD
flabel pdiff 5628 8670 5686 8754 0 FreeSans 320 0 0 0 x1.x4.x5[4].delay_signal
flabel metal4 6173 7493 6274 7562 0 FreeSans 320 0 0 0 x1.x4.x5[4].VDD
flabel via3 6109 8656 6173 8720 0 FreeSans 320 0 0 0 x1.x4.x5[4].floating
flabel viali 6033 8993 6067 9027 0 FreeSans 320 0 0 0 x1.x4.x4[0].SW
flabel ndiff 5977 8871 6035 8955 0 FreeSans 320 0 0 0 x1.x4.x4[0].delay_signal
flabel metal4 5956 10064 6628 10132 0 FreeSans 320 0 0 0 x1.x4.x4[0].VSS
flabel via3 6460 8904 6524 8968 0 FreeSans 320 0 0 0 x1.x4.x4[0].floating
flabel metal1 6770 8589 6804 8623 0 FreeSans 320 0 0 0 x1.x4.x5[3].SW
flabel nwell 6214 7493 6884 7561 0 FreeSans 320 0 0 0 x1.x4.x5[3].VDD
flabel pdiff 6802 8670 6860 8754 0 FreeSans 320 0 0 0 x1.x4.x5[3].delay_signal
flabel metal4 6214 7493 6315 7562 0 FreeSans 320 0 0 0 x1.x4.x5[3].VDD
flabel via3 6315 8656 6379 8720 0 FreeSans 320 0 0 0 x1.x4.x5[3].floating
flabel viali 7249 8993 7283 9027 0 FreeSans 320 0 0 0 x1.x4.x3[1].SW
flabel ndiff 7281 8871 7339 8955 0 FreeSans 320 0 0 0 x1.x4.x3[1].delay_signal
flabel metal4 6688 10064 7360 10132 0 FreeSans 320 0 0 0 x1.x4.x3[1].VSS
flabel via3 6792 8904 6856 8968 0 FreeSans 320 0 0 0 x1.x4.x3[1].floating
flabel metal1 6896 8589 6930 8623 0 FreeSans 320 0 0 0 x1.x4.x5[2].SW
flabel nwell 6816 7493 7486 7561 0 FreeSans 320 0 0 0 x1.x4.x5[2].VDD
flabel pdiff 6840 8670 6898 8754 0 FreeSans 320 0 0 0 x1.x4.x5[2].delay_signal
flabel metal4 7385 7493 7486 7562 0 FreeSans 320 0 0 0 x1.x4.x5[2].VDD
flabel via3 7321 8656 7385 8720 0 FreeSans 320 0 0 0 x1.x4.x5[2].floating
flabel viali 7371 8993 7405 9027 0 FreeSans 320 0 0 0 x1.x4.x3[0].SW
flabel ndiff 7315 8871 7373 8955 0 FreeSans 320 0 0 0 x1.x4.x3[0].delay_signal
flabel metal4 7294 10064 7966 10132 0 FreeSans 320 0 0 0 x1.x4.x3[0].VSS
flabel via3 7798 8904 7862 8968 0 FreeSans 320 0 0 0 x1.x4.x3[0].floating
flabel metal1 7982 8589 8016 8623 0 FreeSans 320 0 0 0 x1.x4.x5[1].SW
flabel nwell 7426 7493 8096 7561 0 FreeSans 320 0 0 0 x1.x4.x5[1].VDD
flabel pdiff 8014 8670 8072 8754 0 FreeSans 320 0 0 0 x1.x4.x5[1].delay_signal
flabel metal4 7426 7493 7527 7562 0 FreeSans 320 0 0 0 x1.x4.x5[1].VDD
flabel via3 7527 8656 7591 8720 0 FreeSans 320 0 0 0 x1.x4.x5[1].floating
flabel viali 8105 8993 8139 9027 0 FreeSans 320 0 0 0 x1.x4.x2.SW
flabel ndiff 8049 8871 8107 8955 0 FreeSans 320 0 0 0 x1.x4.x2.delay_signal
flabel metal4 8028 10064 8700 10132 0 FreeSans 320 0 0 0 x1.x4.x2.VSS
flabel via3 8532 8904 8596 8968 0 FreeSans 320 0 0 0 x1.x4.x2.floating
flabel metal1 8108 8589 8142 8623 0 FreeSans 320 0 0 0 x1.x4.x5[0].SW
flabel nwell 8028 7493 8698 7561 0 FreeSans 320 0 0 0 x1.x4.x5[0].VDD
flabel pdiff 8052 8670 8110 8754 0 FreeSans 320 0 0 0 x1.x4.x5[0].delay_signal
flabel metal4 8597 7493 8698 7562 0 FreeSans 320 0 0 0 x1.x4.x5[0].VDD
flabel via3 8533 8656 8597 8720 0 FreeSans 320 0 0 0 x1.x4.x5[0].floating
flabel metal1 10911 7771 10945 7805 0 FreeSans 200 0 0 0 x1.x3.VGND
flabel metal1 10911 8315 10945 8349 0 FreeSans 200 0 0 0 x1.x3.VPWR
flabel locali 11555 8077 11589 8111 0 FreeSans 250 0 0 0 x1.x3.S
flabel locali 11463 8077 11497 8111 0 FreeSans 250 0 0 0 x1.x3.S
flabel locali 11371 7941 11405 7975 0 FreeSans 250 0 0 0 x1.x3.A1
flabel locali 11371 8009 11405 8043 0 FreeSans 250 0 0 0 x1.x3.A1
flabel locali 11279 8009 11313 8043 0 FreeSans 250 0 0 0 x1.x3.A0
flabel locali 10911 7873 10945 7907 0 FreeSans 250 0 0 0 x1.x3.X
flabel locali 10911 8145 10945 8179 0 FreeSans 250 0 0 0 x1.x3.X
flabel locali 10911 8213 10945 8247 0 FreeSans 250 0 0 0 x1.x3.X
flabel nwell 10955 8315 10989 8349 0 FreeSans 250 0 0 0 x1.x3.VPB
flabel pwell 10965 7771 10999 7805 0 FreeSans 250 0 0 0 x1.x3.VNB
rlabel comment 10881 7788 10881 7788 4 x1.x3.mux2_1
rlabel metal1 10881 7740 11709 7836 1 x1.x3.VGND
rlabel metal1 10881 8284 11709 8380 1 x1.x3.VPWR
flabel metal1 2361 11810 3029 11857 0 FreeSans 320 0 0 0 x1.x2.IN
flabel metal1 8837 11808 9019 11854 0 FreeSans 320 0 0 0 x1.x2.OUT
flabel metal1 2324 12193 2462 12227 0 FreeSans 320 0 0 0 x1.x2.code[3]
flabel metal1 7239 10482 7297 11659 0 FreeSans 320 0 0 0 x1.x2.code[1]
flabel metal1 4813 10482 4871 11659 0 FreeSans 320 0 0 0 x1.x2.code[2]
flabel metal4 2430 12552 2848 13162 0 FreeSans 320 0 0 0 x1.x2.VDD
flabel metal4 2458 10505 2834 11942 0 FreeSans 320 0 0 0 x1.x2.VSS
flabel metal2 2788 11608 3224 11654 0 FreeSans 320 0 0 0 x1.x2.code_offset
flabel metal1 8095 10481 8154 11662 0 FreeSans 320 0 0 0 x1.x2.code[0]
flabel metal1 2972 12263 3006 12297 0 FreeSans 320 0 0 0 x1.x2.x8.input_stack
flabel nwell 3016 13046 3050 13106 0 FreeSans 320 0 0 0 x1.x2.x8.vdd
flabel metal1 3010 12344 3056 12356 0 FreeSans 320 0 0 0 x1.x2.x8.output_stack
flabel poly 2949 11606 3051 11636 0 FreeSans 320 0 0 0 x1.x2.x9.input_stack
flabel metal1 3063 10553 3097 10613 0 FreeSans 320 0 0 0 x1.x2.x9.vss
flabel metal1 3057 11579 3103 11591 0 FreeSans 320 0 0 0 x1.x2.x9.output_stack
flabel locali 2550 12263 2584 12297 0 FreeSans 340 0 0 0 x1.x2.x10.Y
flabel locali 2550 12195 2584 12229 0 FreeSans 340 0 0 0 x1.x2.x10.Y
flabel locali 2458 12195 2492 12229 0 FreeSans 340 0 0 0 x1.x2.x10.A
flabel metal1 2415 11957 2449 11991 0 FreeSans 200 0 0 0 x1.x2.x10.VGND
flabel metal1 2415 12501 2449 12535 0 FreeSans 200 0 0 0 x1.x2.x10.VPWR
rlabel comment 2386 11974 2386 11974 4 x1.x2.x10.inv_1
rlabel metal1 2386 11926 2662 12022 1 x1.x2.x10.VGND
rlabel metal1 2386 12470 2662 12566 1 x1.x2.x10.VPWR
flabel pwell 2415 11957 2449 11991 0 FreeSans 200 0 0 0 x1.x2.x10.VNB
flabel nwell 2415 12501 2449 12535 0 FreeSans 200 0 0 0 x1.x2.x10.VPB
flabel locali 2648 12263 2682 12297 0 FreeSans 340 0 0 0 x1.x2.x11.Y
flabel locali 2648 12195 2682 12229 0 FreeSans 340 0 0 0 x1.x2.x11.Y
flabel locali 2740 12195 2774 12229 0 FreeSans 340 0 0 0 x1.x2.x11.A
flabel metal1 2783 11957 2817 11991 0 FreeSans 200 0 0 0 x1.x2.x11.VGND
flabel metal1 2783 12501 2817 12535 0 FreeSans 200 0 0 0 x1.x2.x11.VPWR
rlabel comment 2846 11974 2846 11974 6 x1.x2.x11.inv_1
rlabel metal1 2570 11926 2846 12022 1 x1.x2.x11.VGND
rlabel metal1 2570 12470 2846 12566 1 x1.x2.x11.VPWR
flabel pwell 2783 11957 2817 11991 0 FreeSans 200 0 0 0 x1.x2.x11.VNB
flabel nwell 2783 12501 2817 12535 0 FreeSans 200 0 0 0 x1.x2.x11.VPB
flabel metal1 3614 12020 3648 12054 0 FreeSans 320 0 0 0 x1.x2.x6.SW
flabel nwell 3058 13082 3728 13150 0 FreeSans 320 0 0 0 x1.x2.x6.VDD
flabel pdiff 3646 11889 3704 11973 0 FreeSans 320 0 0 0 x1.x2.x6.delay_signal
flabel metal4 3058 13081 3159 13150 0 FreeSans 320 0 0 0 x1.x2.x6.VDD
flabel via3 3159 11923 3223 11987 0 FreeSans 320 0 0 0 x1.x2.x6.floating
flabel viali 3967 11619 4001 11653 0 FreeSans 320 0 0 0 x1.x2.x7.SW
flabel ndiff 3999 11691 4057 11775 0 FreeSans 320 0 0 0 x1.x2.x7.delay_signal
flabel metal4 3406 10514 4078 10582 0 FreeSans 320 0 0 0 x1.x2.x7.VSS
flabel via3 3510 11678 3574 11742 0 FreeSans 320 0 0 0 x1.x2.x7.floating
flabel viali 4699 11619 4733 11653 0 FreeSans 320 0 0 0 x1.x2.x4[3].SW
flabel ndiff 4731 11691 4789 11775 0 FreeSans 320 0 0 0 x1.x2.x4[3].delay_signal
flabel metal4 4138 10514 4810 10582 0 FreeSans 320 0 0 0 x1.x2.x4[3].VSS
flabel via3 4242 11678 4306 11742 0 FreeSans 320 0 0 0 x1.x2.x4[3].floating
flabel metal1 4472 12023 4506 12057 0 FreeSans 320 0 0 0 x1.x2.x5[6].SW
flabel nwell 4392 13085 5062 13153 0 FreeSans 320 0 0 0 x1.x2.x5[6].VDD
flabel pdiff 4416 11892 4474 11976 0 FreeSans 320 0 0 0 x1.x2.x5[6].delay_signal
flabel metal4 4961 13084 5062 13153 0 FreeSans 320 0 0 0 x1.x2.x5[6].VDD
flabel via3 4897 11926 4961 11990 0 FreeSans 320 0 0 0 x1.x2.x5[6].floating
flabel metal1 4346 12023 4380 12057 0 FreeSans 320 0 0 0 x1.x2.x5[7].SW
flabel nwell 3790 13085 4460 13153 0 FreeSans 320 0 0 0 x1.x2.x5[7].VDD
flabel pdiff 4378 11892 4436 11976 0 FreeSans 320 0 0 0 x1.x2.x5[7].delay_signal
flabel metal4 3790 13084 3891 13153 0 FreeSans 320 0 0 0 x1.x2.x5[7].VDD
flabel via3 3891 11926 3955 11990 0 FreeSans 320 0 0 0 x1.x2.x5[7].floating
flabel viali 4821 11619 4855 11653 0 FreeSans 320 0 0 0 x1.x2.x4[2].SW
flabel ndiff 4765 11691 4823 11775 0 FreeSans 320 0 0 0 x1.x2.x4[2].delay_signal
flabel metal4 4744 10514 5416 10582 0 FreeSans 320 0 0 0 x1.x2.x4[2].VSS
flabel via3 5248 11678 5312 11742 0 FreeSans 320 0 0 0 x1.x2.x4[2].floating
flabel metal1 5558 12023 5592 12057 0 FreeSans 320 0 0 0 x1.x2.x5[5].SW
flabel nwell 5002 13085 5672 13153 0 FreeSans 320 0 0 0 x1.x2.x5[5].VDD
flabel pdiff 5590 11892 5648 11976 0 FreeSans 320 0 0 0 x1.x2.x5[5].delay_signal
flabel metal4 5002 13084 5103 13153 0 FreeSans 320 0 0 0 x1.x2.x5[5].VDD
flabel via3 5103 11926 5167 11990 0 FreeSans 320 0 0 0 x1.x2.x5[5].floating
flabel viali 5911 11619 5945 11653 0 FreeSans 320 0 0 0 x1.x2.x4[1].SW
flabel ndiff 5943 11691 6001 11775 0 FreeSans 320 0 0 0 x1.x2.x4[1].delay_signal
flabel metal4 5350 10514 6022 10582 0 FreeSans 320 0 0 0 x1.x2.x4[1].VSS
flabel via3 5454 11678 5518 11742 0 FreeSans 320 0 0 0 x1.x2.x4[1].floating
flabel metal1 5684 12023 5718 12057 0 FreeSans 320 0 0 0 x1.x2.x5[4].SW
flabel nwell 5604 13085 6274 13153 0 FreeSans 320 0 0 0 x1.x2.x5[4].VDD
flabel pdiff 5628 11892 5686 11976 0 FreeSans 320 0 0 0 x1.x2.x5[4].delay_signal
flabel metal4 6173 13084 6274 13153 0 FreeSans 320 0 0 0 x1.x2.x5[4].VDD
flabel via3 6109 11926 6173 11990 0 FreeSans 320 0 0 0 x1.x2.x5[4].floating
flabel viali 6033 11619 6067 11653 0 FreeSans 320 0 0 0 x1.x2.x4[0].SW
flabel ndiff 5977 11691 6035 11775 0 FreeSans 320 0 0 0 x1.x2.x4[0].delay_signal
flabel metal4 5956 10514 6628 10582 0 FreeSans 320 0 0 0 x1.x2.x4[0].VSS
flabel via3 6460 11678 6524 11742 0 FreeSans 320 0 0 0 x1.x2.x4[0].floating
flabel metal1 6770 12023 6804 12057 0 FreeSans 320 0 0 0 x1.x2.x5[3].SW
flabel nwell 6214 13085 6884 13153 0 FreeSans 320 0 0 0 x1.x2.x5[3].VDD
flabel pdiff 6802 11892 6860 11976 0 FreeSans 320 0 0 0 x1.x2.x5[3].delay_signal
flabel metal4 6214 13084 6315 13153 0 FreeSans 320 0 0 0 x1.x2.x5[3].VDD
flabel via3 6315 11926 6379 11990 0 FreeSans 320 0 0 0 x1.x2.x5[3].floating
flabel viali 7249 11619 7283 11653 0 FreeSans 320 0 0 0 x1.x2.x3[1].SW
flabel ndiff 7281 11691 7339 11775 0 FreeSans 320 0 0 0 x1.x2.x3[1].delay_signal
flabel metal4 6688 10514 7360 10582 0 FreeSans 320 0 0 0 x1.x2.x3[1].VSS
flabel via3 6792 11678 6856 11742 0 FreeSans 320 0 0 0 x1.x2.x3[1].floating
flabel metal1 6896 12023 6930 12057 0 FreeSans 320 0 0 0 x1.x2.x5[2].SW
flabel nwell 6816 13085 7486 13153 0 FreeSans 320 0 0 0 x1.x2.x5[2].VDD
flabel pdiff 6840 11892 6898 11976 0 FreeSans 320 0 0 0 x1.x2.x5[2].delay_signal
flabel metal4 7385 13084 7486 13153 0 FreeSans 320 0 0 0 x1.x2.x5[2].VDD
flabel via3 7321 11926 7385 11990 0 FreeSans 320 0 0 0 x1.x2.x5[2].floating
flabel viali 7371 11619 7405 11653 0 FreeSans 320 0 0 0 x1.x2.x3[0].SW
flabel ndiff 7315 11691 7373 11775 0 FreeSans 320 0 0 0 x1.x2.x3[0].delay_signal
flabel metal4 7294 10514 7966 10582 0 FreeSans 320 0 0 0 x1.x2.x3[0].VSS
flabel via3 7798 11678 7862 11742 0 FreeSans 320 0 0 0 x1.x2.x3[0].floating
flabel metal1 7982 12023 8016 12057 0 FreeSans 320 0 0 0 x1.x2.x5[1].SW
flabel nwell 7426 13085 8096 13153 0 FreeSans 320 0 0 0 x1.x2.x5[1].VDD
flabel pdiff 8014 11892 8072 11976 0 FreeSans 320 0 0 0 x1.x2.x5[1].delay_signal
flabel metal4 7426 13084 7527 13153 0 FreeSans 320 0 0 0 x1.x2.x5[1].VDD
flabel via3 7527 11926 7591 11990 0 FreeSans 320 0 0 0 x1.x2.x5[1].floating
flabel viali 8105 11619 8139 11653 0 FreeSans 320 0 0 0 x1.x2.x2.SW
flabel ndiff 8049 11691 8107 11775 0 FreeSans 320 0 0 0 x1.x2.x2.delay_signal
flabel metal4 8028 10514 8700 10582 0 FreeSans 320 0 0 0 x1.x2.x2.VSS
flabel via3 8532 11678 8596 11742 0 FreeSans 320 0 0 0 x1.x2.x2.floating
flabel metal1 8108 12023 8142 12057 0 FreeSans 320 0 0 0 x1.x2.x5[0].SW
flabel nwell 8028 13085 8698 13153 0 FreeSans 320 0 0 0 x1.x2.x5[0].VDD
flabel pdiff 8052 11892 8110 11976 0 FreeSans 320 0 0 0 x1.x2.x5[0].delay_signal
flabel metal4 8597 13084 8698 13153 0 FreeSans 320 0 0 0 x1.x2.x5[0].VDD
flabel via3 8533 11926 8597 11990 0 FreeSans 320 0 0 0 x1.x2.x5[0].floating
<< end >>
