magic
tech sky130A
magscale 1 2
timestamp 1698578866
<< nwell >>
rect -796 -170 796 261
<< pmos >>
rect -600 -42 600 42
<< pdiff >>
rect -658 30 -600 42
rect -658 -30 -646 30
rect -612 -30 -600 30
rect -658 -42 -600 -30
rect 600 30 658 42
rect 600 -30 612 30
rect 646 -30 658 30
rect 600 -42 658 -30
<< pdiffc >>
rect -646 -30 -612 30
rect 612 -30 646 30
<< nsubdiff >>
rect -760 191 -664 225
rect 664 191 760 225
rect -760 129 -726 191
rect 726 129 760 191
rect -760 -100 -726 -66
rect 726 -100 760 -66
rect -760 -134 -664 -100
rect 664 -134 760 -100
<< nsubdiffcont >>
rect -664 191 664 225
rect -760 -66 -726 129
rect 726 -66 760 129
rect -664 -134 664 -100
<< poly >>
rect -600 123 600 139
rect -600 89 -584 123
rect 584 89 600 123
rect -600 42 600 89
rect -600 -68 600 -42
<< polycont >>
rect -584 89 584 123
<< locali >>
rect -760 191 -664 225
rect 664 191 760 225
rect -760 129 -726 191
rect 726 129 760 191
rect -600 89 -584 123
rect 584 89 600 123
rect -760 -100 -726 -66
rect -646 30 -612 46
rect -646 -100 -612 -30
rect 612 30 646 46
rect 612 -100 646 -30
rect 726 -100 760 -66
rect -760 -134 -664 -100
rect 664 -134 760 -100
<< viali >>
rect -584 89 584 123
rect -646 -30 -612 30
rect 612 -30 646 30
<< metal1 >>
rect -596 123 596 129
rect -596 89 -584 123
rect 584 89 596 123
rect -596 83 596 89
rect -652 30 -606 42
rect -652 -30 -646 30
rect -612 -30 -606 30
rect -652 -42 -606 -30
rect 606 30 652 42
rect 606 -30 612 30
rect 646 -30 652 30
rect 606 -42 652 -30
<< properties >>
string FIXED_BBOX -743 -208 743 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 6.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
