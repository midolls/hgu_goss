magic
tech sky130A
magscale 1 2
timestamp 1699171588
<< pwell >>
rect 14108 3744 14134 3776
rect 14714 3744 14740 3776
rect 15320 3744 15346 3776
rect 15926 3744 15952 3776
rect 16532 3744 16558 3776
rect 17138 3744 17164 3776
rect 17744 3744 17770 3776
rect 18350 3744 18376 3776
rect 18956 3744 18982 3776
rect 19562 3744 19588 3776
rect 20168 3744 20194 3776
rect 20774 3744 20800 3776
rect 21380 3744 21406 3776
rect 21986 3744 22012 3776
rect 22592 3744 22618 3776
rect 23198 3744 23224 3776
rect 23804 3744 23830 3776
rect 24410 3744 24436 3776
rect 25016 3744 25042 3776
rect 25622 3744 25648 3776
rect 26228 3744 26254 3776
rect 26834 3744 26860 3776
rect 27440 3744 27466 3776
rect 28046 3744 28072 3776
rect 28652 3744 28678 3776
rect 29258 3744 29284 3776
rect 29864 3744 29890 3776
rect 30470 3744 30496 3776
rect 31076 3744 31102 3776
rect 31682 3744 31708 3776
rect 32288 3744 32314 3776
rect 32894 3744 32920 3776
rect 14102 2220 14128 2252
rect 14708 2220 14734 2252
rect 15314 2220 15340 2252
rect 15920 2220 15946 2252
rect 16526 2220 16552 2252
rect 17132 2220 17158 2252
rect 17738 2220 17764 2252
rect 18344 2220 18370 2252
rect 18950 2220 18976 2252
rect 19556 2220 19582 2252
rect 20162 2220 20188 2252
rect 20768 2220 20794 2252
rect 21374 2220 21400 2252
rect 21980 2220 22006 2252
rect 22586 2220 22612 2252
rect 23192 2220 23218 2252
rect 23798 2220 23824 2252
rect 24404 2220 24430 2252
rect 25010 2220 25036 2252
rect 25616 2220 25642 2252
rect 26222 2220 26248 2252
rect 26828 2220 26854 2252
rect 27434 2220 27460 2252
rect 28040 2220 28066 2252
rect 28646 2220 28672 2252
rect 29252 2220 29278 2252
rect 29858 2220 29884 2252
rect 30464 2220 30490 2252
rect 31070 2220 31096 2252
rect 31676 2220 31702 2252
rect 32282 2220 32308 2252
rect 32888 2220 32914 2252
<< psubdiff >>
rect 22704 3266 22746 3356
<< metal3 >>
rect 13782 4190 33240 4192
rect 13782 4126 13886 4190
rect 13950 4126 13966 4190
rect 14030 4126 14046 4190
rect 14110 4126 14126 4190
rect 14190 4126 14206 4190
rect 14270 4126 14286 4190
rect 14350 4126 14492 4190
rect 14556 4126 14572 4190
rect 14636 4126 14652 4190
rect 14716 4126 14732 4190
rect 14796 4126 14812 4190
rect 14876 4126 14892 4190
rect 14956 4126 15098 4190
rect 15162 4126 15178 4190
rect 15242 4126 15258 4190
rect 15322 4126 15338 4190
rect 15402 4126 15418 4190
rect 15482 4126 15498 4190
rect 15562 4126 15704 4190
rect 15768 4126 15784 4190
rect 15848 4126 15864 4190
rect 15928 4126 15944 4190
rect 16008 4126 16024 4190
rect 16088 4126 16104 4190
rect 16168 4126 16310 4190
rect 16374 4126 16390 4190
rect 16454 4126 16470 4190
rect 16534 4126 16550 4190
rect 16614 4126 16630 4190
rect 16694 4126 16710 4190
rect 16774 4126 16916 4190
rect 16980 4126 16996 4190
rect 17060 4126 17076 4190
rect 17140 4126 17156 4190
rect 17220 4126 17236 4190
rect 17300 4126 17316 4190
rect 17380 4126 17522 4190
rect 17586 4126 17602 4190
rect 17666 4126 17682 4190
rect 17746 4126 17762 4190
rect 17826 4126 17842 4190
rect 17906 4126 17922 4190
rect 17986 4126 18128 4190
rect 18192 4126 18208 4190
rect 18272 4126 18288 4190
rect 18352 4126 18368 4190
rect 18432 4126 18448 4190
rect 18512 4126 18528 4190
rect 18592 4126 18734 4190
rect 18798 4126 18814 4190
rect 18878 4126 18894 4190
rect 18958 4126 18974 4190
rect 19038 4126 19054 4190
rect 19118 4126 19134 4190
rect 19198 4126 19340 4190
rect 19404 4126 19420 4190
rect 19484 4126 19500 4190
rect 19564 4126 19580 4190
rect 19644 4126 19660 4190
rect 19724 4126 19740 4190
rect 19804 4126 19946 4190
rect 20010 4126 20026 4190
rect 20090 4126 20106 4190
rect 20170 4126 20186 4190
rect 20250 4126 20266 4190
rect 20330 4126 20346 4190
rect 20410 4126 20552 4190
rect 20616 4126 20632 4190
rect 20696 4126 20712 4190
rect 20776 4126 20792 4190
rect 20856 4126 20872 4190
rect 20936 4126 20952 4190
rect 21016 4126 21158 4190
rect 21222 4126 21238 4190
rect 21302 4126 21318 4190
rect 21382 4126 21398 4190
rect 21462 4126 21478 4190
rect 21542 4126 21558 4190
rect 21622 4126 21764 4190
rect 21828 4126 21844 4190
rect 21908 4126 21924 4190
rect 21988 4126 22004 4190
rect 22068 4126 22084 4190
rect 22148 4126 22164 4190
rect 22228 4126 22370 4190
rect 22434 4126 22450 4190
rect 22514 4126 22530 4190
rect 22594 4126 22610 4190
rect 22674 4126 22690 4190
rect 22754 4126 22770 4190
rect 22834 4126 22976 4190
rect 23040 4126 23056 4190
rect 23120 4126 23136 4190
rect 23200 4126 23216 4190
rect 23280 4126 23296 4190
rect 23360 4126 23376 4190
rect 23440 4126 23582 4190
rect 23646 4126 23662 4190
rect 23726 4126 23742 4190
rect 23806 4126 23822 4190
rect 23886 4126 23902 4190
rect 23966 4126 23982 4190
rect 24046 4126 24188 4190
rect 24252 4126 24268 4190
rect 24332 4126 24348 4190
rect 24412 4126 24428 4190
rect 24492 4126 24508 4190
rect 24572 4126 24588 4190
rect 24652 4126 24794 4190
rect 24858 4126 24874 4190
rect 24938 4126 24954 4190
rect 25018 4126 25034 4190
rect 25098 4126 25114 4190
rect 25178 4126 25194 4190
rect 25258 4126 25400 4190
rect 25464 4126 25480 4190
rect 25544 4126 25560 4190
rect 25624 4126 25640 4190
rect 25704 4126 25720 4190
rect 25784 4126 25800 4190
rect 25864 4126 26006 4190
rect 26070 4126 26086 4190
rect 26150 4126 26166 4190
rect 26230 4126 26246 4190
rect 26310 4126 26326 4190
rect 26390 4126 26406 4190
rect 26470 4126 26612 4190
rect 26676 4126 26692 4190
rect 26756 4126 26772 4190
rect 26836 4126 26852 4190
rect 26916 4126 26932 4190
rect 26996 4126 27012 4190
rect 27076 4126 27218 4190
rect 27282 4126 27298 4190
rect 27362 4126 27378 4190
rect 27442 4126 27458 4190
rect 27522 4126 27538 4190
rect 27602 4126 27618 4190
rect 27682 4126 27824 4190
rect 27888 4126 27904 4190
rect 27968 4126 27984 4190
rect 28048 4126 28064 4190
rect 28128 4126 28144 4190
rect 28208 4126 28224 4190
rect 28288 4126 28430 4190
rect 28494 4126 28510 4190
rect 28574 4126 28590 4190
rect 28654 4126 28670 4190
rect 28734 4126 28750 4190
rect 28814 4126 28830 4190
rect 28894 4126 29036 4190
rect 29100 4126 29116 4190
rect 29180 4126 29196 4190
rect 29260 4126 29276 4190
rect 29340 4126 29356 4190
rect 29420 4126 29436 4190
rect 29500 4126 29642 4190
rect 29706 4126 29722 4190
rect 29786 4126 29802 4190
rect 29866 4126 29882 4190
rect 29946 4126 29962 4190
rect 30026 4126 30042 4190
rect 30106 4126 30248 4190
rect 30312 4126 30328 4190
rect 30392 4126 30408 4190
rect 30472 4126 30488 4190
rect 30552 4126 30568 4190
rect 30632 4126 30648 4190
rect 30712 4126 30854 4190
rect 30918 4126 30934 4190
rect 30998 4126 31014 4190
rect 31078 4126 31094 4190
rect 31158 4126 31174 4190
rect 31238 4126 31254 4190
rect 31318 4126 31460 4190
rect 31524 4126 31540 4190
rect 31604 4126 31620 4190
rect 31684 4126 31700 4190
rect 31764 4126 31780 4190
rect 31844 4126 31860 4190
rect 31924 4126 32066 4190
rect 32130 4126 32146 4190
rect 32210 4126 32226 4190
rect 32290 4126 32306 4190
rect 32370 4126 32386 4190
rect 32450 4126 32466 4190
rect 32530 4126 32672 4190
rect 32736 4126 32752 4190
rect 32816 4126 32832 4190
rect 32896 4126 32912 4190
rect 32976 4126 32992 4190
rect 33056 4126 33072 4190
rect 33136 4126 33240 4190
rect 13782 4124 33240 4126
rect 13782 3970 13848 4060
rect 13782 3906 13783 3970
rect 13847 3906 13848 3970
rect 13782 3890 13848 3906
rect 13782 3826 13783 3890
rect 13847 3826 13848 3890
rect 13782 3810 13848 3826
rect 13782 3746 13783 3810
rect 13847 3746 13848 3810
rect 13782 3730 13848 3746
rect 13782 3666 13783 3730
rect 13847 3666 13848 3730
rect 13782 3650 13848 3666
rect 13782 3586 13783 3650
rect 13847 3586 13848 3650
rect 13782 3570 13848 3586
rect 13782 3506 13783 3570
rect 13847 3506 13848 3570
rect 13782 3490 13848 3506
rect 13782 3426 13783 3490
rect 13847 3426 13848 3490
rect 13782 3410 13848 3426
rect 13782 3346 13783 3410
rect 13847 3346 13848 3410
rect 13782 3330 13848 3346
rect 13782 3266 13783 3330
rect 13847 3266 13848 3330
rect 13782 3250 13848 3266
rect 13782 3186 13783 3250
rect 13847 3186 13848 3250
rect 13782 3032 13848 3186
rect 13908 3094 13968 4124
rect 14028 3032 14088 4064
rect 14148 3094 14208 4124
rect 14268 3032 14328 4064
rect 14388 3970 14454 4060
rect 14388 3906 14389 3970
rect 14453 3906 14454 3970
rect 14388 3890 14454 3906
rect 14388 3826 14389 3890
rect 14453 3826 14454 3890
rect 14388 3810 14454 3826
rect 14388 3746 14389 3810
rect 14453 3746 14454 3810
rect 14388 3730 14454 3746
rect 14388 3666 14389 3730
rect 14453 3666 14454 3730
rect 14388 3650 14454 3666
rect 14388 3586 14389 3650
rect 14453 3586 14454 3650
rect 14388 3570 14454 3586
rect 14388 3506 14389 3570
rect 14453 3506 14454 3570
rect 14388 3490 14454 3506
rect 14388 3426 14389 3490
rect 14453 3426 14454 3490
rect 14388 3410 14454 3426
rect 14388 3346 14389 3410
rect 14453 3346 14454 3410
rect 14388 3330 14454 3346
rect 14388 3266 14389 3330
rect 14453 3266 14454 3330
rect 14388 3250 14454 3266
rect 14388 3186 14389 3250
rect 14453 3186 14454 3250
rect 14388 3032 14454 3186
rect 14514 3094 14574 4124
rect 14634 3032 14694 4064
rect 14754 3094 14814 4124
rect 14874 3032 14934 4064
rect 14994 3970 15060 4060
rect 14994 3906 14995 3970
rect 15059 3906 15060 3970
rect 14994 3890 15060 3906
rect 14994 3826 14995 3890
rect 15059 3826 15060 3890
rect 14994 3810 15060 3826
rect 14994 3746 14995 3810
rect 15059 3746 15060 3810
rect 14994 3730 15060 3746
rect 14994 3666 14995 3730
rect 15059 3666 15060 3730
rect 14994 3650 15060 3666
rect 14994 3586 14995 3650
rect 15059 3586 15060 3650
rect 14994 3570 15060 3586
rect 14994 3506 14995 3570
rect 15059 3506 15060 3570
rect 14994 3490 15060 3506
rect 14994 3426 14995 3490
rect 15059 3426 15060 3490
rect 14994 3410 15060 3426
rect 14994 3346 14995 3410
rect 15059 3346 15060 3410
rect 14994 3330 15060 3346
rect 14994 3266 14995 3330
rect 15059 3266 15060 3330
rect 14994 3250 15060 3266
rect 14994 3186 14995 3250
rect 15059 3186 15060 3250
rect 14994 3032 15060 3186
rect 15120 3094 15180 4124
rect 15240 3032 15300 4064
rect 15360 3094 15420 4124
rect 15480 3032 15540 4064
rect 15600 3970 15666 4060
rect 15600 3906 15601 3970
rect 15665 3906 15666 3970
rect 15600 3890 15666 3906
rect 15600 3826 15601 3890
rect 15665 3826 15666 3890
rect 15600 3810 15666 3826
rect 15600 3746 15601 3810
rect 15665 3746 15666 3810
rect 15600 3730 15666 3746
rect 15600 3666 15601 3730
rect 15665 3666 15666 3730
rect 15600 3650 15666 3666
rect 15600 3586 15601 3650
rect 15665 3586 15666 3650
rect 15600 3570 15666 3586
rect 15600 3506 15601 3570
rect 15665 3506 15666 3570
rect 15600 3490 15666 3506
rect 15600 3426 15601 3490
rect 15665 3426 15666 3490
rect 15600 3410 15666 3426
rect 15600 3346 15601 3410
rect 15665 3346 15666 3410
rect 15600 3330 15666 3346
rect 15600 3266 15601 3330
rect 15665 3266 15666 3330
rect 15600 3250 15666 3266
rect 15600 3186 15601 3250
rect 15665 3186 15666 3250
rect 15600 3032 15666 3186
rect 15726 3094 15786 4124
rect 15846 3032 15906 4064
rect 15966 3094 16026 4124
rect 16086 3032 16146 4064
rect 16206 3970 16272 4060
rect 16206 3906 16207 3970
rect 16271 3906 16272 3970
rect 16206 3890 16272 3906
rect 16206 3826 16207 3890
rect 16271 3826 16272 3890
rect 16206 3810 16272 3826
rect 16206 3746 16207 3810
rect 16271 3746 16272 3810
rect 16206 3730 16272 3746
rect 16206 3666 16207 3730
rect 16271 3666 16272 3730
rect 16206 3650 16272 3666
rect 16206 3586 16207 3650
rect 16271 3586 16272 3650
rect 16206 3570 16272 3586
rect 16206 3506 16207 3570
rect 16271 3506 16272 3570
rect 16206 3490 16272 3506
rect 16206 3426 16207 3490
rect 16271 3426 16272 3490
rect 16206 3410 16272 3426
rect 16206 3346 16207 3410
rect 16271 3346 16272 3410
rect 16206 3330 16272 3346
rect 16206 3266 16207 3330
rect 16271 3266 16272 3330
rect 16206 3250 16272 3266
rect 16206 3186 16207 3250
rect 16271 3186 16272 3250
rect 16206 3032 16272 3186
rect 16332 3094 16392 4124
rect 16452 3032 16512 4064
rect 16572 3094 16632 4124
rect 16692 3032 16752 4064
rect 16812 3970 16878 4060
rect 16812 3906 16813 3970
rect 16877 3906 16878 3970
rect 16812 3890 16878 3906
rect 16812 3826 16813 3890
rect 16877 3826 16878 3890
rect 16812 3810 16878 3826
rect 16812 3746 16813 3810
rect 16877 3746 16878 3810
rect 16812 3730 16878 3746
rect 16812 3666 16813 3730
rect 16877 3666 16878 3730
rect 16812 3650 16878 3666
rect 16812 3586 16813 3650
rect 16877 3586 16878 3650
rect 16812 3570 16878 3586
rect 16812 3506 16813 3570
rect 16877 3506 16878 3570
rect 16812 3490 16878 3506
rect 16812 3426 16813 3490
rect 16877 3426 16878 3490
rect 16812 3410 16878 3426
rect 16812 3346 16813 3410
rect 16877 3346 16878 3410
rect 16812 3330 16878 3346
rect 16812 3266 16813 3330
rect 16877 3266 16878 3330
rect 16812 3250 16878 3266
rect 16812 3186 16813 3250
rect 16877 3186 16878 3250
rect 16812 3032 16878 3186
rect 16938 3094 16998 4124
rect 17058 3032 17118 4064
rect 17178 3094 17238 4124
rect 17298 3032 17358 4064
rect 17418 3970 17484 4060
rect 17418 3906 17419 3970
rect 17483 3906 17484 3970
rect 17418 3890 17484 3906
rect 17418 3826 17419 3890
rect 17483 3826 17484 3890
rect 17418 3810 17484 3826
rect 17418 3746 17419 3810
rect 17483 3746 17484 3810
rect 17418 3730 17484 3746
rect 17418 3666 17419 3730
rect 17483 3666 17484 3730
rect 17418 3650 17484 3666
rect 17418 3586 17419 3650
rect 17483 3586 17484 3650
rect 17418 3570 17484 3586
rect 17418 3506 17419 3570
rect 17483 3506 17484 3570
rect 17418 3490 17484 3506
rect 17418 3426 17419 3490
rect 17483 3426 17484 3490
rect 17418 3410 17484 3426
rect 17418 3346 17419 3410
rect 17483 3346 17484 3410
rect 17418 3330 17484 3346
rect 17418 3266 17419 3330
rect 17483 3266 17484 3330
rect 17418 3250 17484 3266
rect 17418 3186 17419 3250
rect 17483 3186 17484 3250
rect 17418 3032 17484 3186
rect 17544 3094 17604 4124
rect 17664 3032 17724 4064
rect 17784 3094 17844 4124
rect 17904 3032 17964 4064
rect 18024 3970 18090 4060
rect 18024 3906 18025 3970
rect 18089 3906 18090 3970
rect 18024 3890 18090 3906
rect 18024 3826 18025 3890
rect 18089 3826 18090 3890
rect 18024 3810 18090 3826
rect 18024 3746 18025 3810
rect 18089 3746 18090 3810
rect 18024 3730 18090 3746
rect 18024 3666 18025 3730
rect 18089 3666 18090 3730
rect 18024 3650 18090 3666
rect 18024 3586 18025 3650
rect 18089 3586 18090 3650
rect 18024 3570 18090 3586
rect 18024 3506 18025 3570
rect 18089 3506 18090 3570
rect 18024 3490 18090 3506
rect 18024 3426 18025 3490
rect 18089 3426 18090 3490
rect 18024 3410 18090 3426
rect 18024 3346 18025 3410
rect 18089 3346 18090 3410
rect 18024 3330 18090 3346
rect 18024 3266 18025 3330
rect 18089 3266 18090 3330
rect 18024 3250 18090 3266
rect 18024 3186 18025 3250
rect 18089 3186 18090 3250
rect 18024 3032 18090 3186
rect 18150 3094 18210 4124
rect 18270 3032 18330 4064
rect 18390 3094 18450 4124
rect 18510 3032 18570 4064
rect 18630 3970 18696 4060
rect 18630 3906 18631 3970
rect 18695 3906 18696 3970
rect 18630 3890 18696 3906
rect 18630 3826 18631 3890
rect 18695 3826 18696 3890
rect 18630 3810 18696 3826
rect 18630 3746 18631 3810
rect 18695 3746 18696 3810
rect 18630 3730 18696 3746
rect 18630 3666 18631 3730
rect 18695 3666 18696 3730
rect 18630 3650 18696 3666
rect 18630 3586 18631 3650
rect 18695 3586 18696 3650
rect 18630 3570 18696 3586
rect 18630 3506 18631 3570
rect 18695 3506 18696 3570
rect 18630 3490 18696 3506
rect 18630 3426 18631 3490
rect 18695 3426 18696 3490
rect 18630 3410 18696 3426
rect 18630 3346 18631 3410
rect 18695 3346 18696 3410
rect 18630 3330 18696 3346
rect 18630 3266 18631 3330
rect 18695 3266 18696 3330
rect 18630 3250 18696 3266
rect 18630 3186 18631 3250
rect 18695 3186 18696 3250
rect 18630 3032 18696 3186
rect 18756 3094 18816 4124
rect 18876 3032 18936 4064
rect 18996 3094 19056 4124
rect 19116 3032 19176 4064
rect 19236 3970 19302 4060
rect 19236 3906 19237 3970
rect 19301 3906 19302 3970
rect 19236 3890 19302 3906
rect 19236 3826 19237 3890
rect 19301 3826 19302 3890
rect 19236 3810 19302 3826
rect 19236 3746 19237 3810
rect 19301 3746 19302 3810
rect 19236 3730 19302 3746
rect 19236 3666 19237 3730
rect 19301 3666 19302 3730
rect 19236 3650 19302 3666
rect 19236 3586 19237 3650
rect 19301 3586 19302 3650
rect 19236 3570 19302 3586
rect 19236 3506 19237 3570
rect 19301 3506 19302 3570
rect 19236 3490 19302 3506
rect 19236 3426 19237 3490
rect 19301 3426 19302 3490
rect 19236 3410 19302 3426
rect 19236 3346 19237 3410
rect 19301 3346 19302 3410
rect 19236 3330 19302 3346
rect 19236 3266 19237 3330
rect 19301 3266 19302 3330
rect 19236 3250 19302 3266
rect 19236 3186 19237 3250
rect 19301 3186 19302 3250
rect 19236 3032 19302 3186
rect 19362 3094 19422 4124
rect 19482 3032 19542 4064
rect 19602 3094 19662 4124
rect 19722 3032 19782 4064
rect 19842 3970 19908 4060
rect 19842 3906 19843 3970
rect 19907 3906 19908 3970
rect 19842 3890 19908 3906
rect 19842 3826 19843 3890
rect 19907 3826 19908 3890
rect 19842 3810 19908 3826
rect 19842 3746 19843 3810
rect 19907 3746 19908 3810
rect 19842 3730 19908 3746
rect 19842 3666 19843 3730
rect 19907 3666 19908 3730
rect 19842 3650 19908 3666
rect 19842 3586 19843 3650
rect 19907 3586 19908 3650
rect 19842 3570 19908 3586
rect 19842 3506 19843 3570
rect 19907 3506 19908 3570
rect 19842 3490 19908 3506
rect 19842 3426 19843 3490
rect 19907 3426 19908 3490
rect 19842 3410 19908 3426
rect 19842 3346 19843 3410
rect 19907 3346 19908 3410
rect 19842 3330 19908 3346
rect 19842 3266 19843 3330
rect 19907 3266 19908 3330
rect 19842 3250 19908 3266
rect 19842 3186 19843 3250
rect 19907 3186 19908 3250
rect 19842 3032 19908 3186
rect 19968 3094 20028 4124
rect 20088 3032 20148 4064
rect 20208 3094 20268 4124
rect 20328 3032 20388 4064
rect 20448 3970 20514 4060
rect 20448 3906 20449 3970
rect 20513 3906 20514 3970
rect 20448 3890 20514 3906
rect 20448 3826 20449 3890
rect 20513 3826 20514 3890
rect 20448 3810 20514 3826
rect 20448 3746 20449 3810
rect 20513 3746 20514 3810
rect 20448 3730 20514 3746
rect 20448 3666 20449 3730
rect 20513 3666 20514 3730
rect 20448 3650 20514 3666
rect 20448 3586 20449 3650
rect 20513 3586 20514 3650
rect 20448 3570 20514 3586
rect 20448 3506 20449 3570
rect 20513 3506 20514 3570
rect 20448 3490 20514 3506
rect 20448 3426 20449 3490
rect 20513 3426 20514 3490
rect 20448 3410 20514 3426
rect 20448 3346 20449 3410
rect 20513 3346 20514 3410
rect 20448 3330 20514 3346
rect 20448 3266 20449 3330
rect 20513 3266 20514 3330
rect 20448 3250 20514 3266
rect 20448 3186 20449 3250
rect 20513 3186 20514 3250
rect 20448 3032 20514 3186
rect 20574 3094 20634 4124
rect 20694 3032 20754 4064
rect 20814 3094 20874 4124
rect 20934 3032 20994 4064
rect 21054 3970 21120 4060
rect 21054 3906 21055 3970
rect 21119 3906 21120 3970
rect 21054 3890 21120 3906
rect 21054 3826 21055 3890
rect 21119 3826 21120 3890
rect 21054 3810 21120 3826
rect 21054 3746 21055 3810
rect 21119 3746 21120 3810
rect 21054 3730 21120 3746
rect 21054 3666 21055 3730
rect 21119 3666 21120 3730
rect 21054 3650 21120 3666
rect 21054 3586 21055 3650
rect 21119 3586 21120 3650
rect 21054 3570 21120 3586
rect 21054 3506 21055 3570
rect 21119 3506 21120 3570
rect 21054 3490 21120 3506
rect 21054 3426 21055 3490
rect 21119 3426 21120 3490
rect 21054 3410 21120 3426
rect 21054 3346 21055 3410
rect 21119 3346 21120 3410
rect 21054 3330 21120 3346
rect 21054 3266 21055 3330
rect 21119 3266 21120 3330
rect 21054 3250 21120 3266
rect 21054 3186 21055 3250
rect 21119 3186 21120 3250
rect 21054 3032 21120 3186
rect 21180 3094 21240 4124
rect 21300 3032 21360 4064
rect 21420 3094 21480 4124
rect 21540 3032 21600 4064
rect 21660 3970 21726 4060
rect 21660 3906 21661 3970
rect 21725 3906 21726 3970
rect 21660 3890 21726 3906
rect 21660 3826 21661 3890
rect 21725 3826 21726 3890
rect 21660 3810 21726 3826
rect 21660 3746 21661 3810
rect 21725 3746 21726 3810
rect 21660 3730 21726 3746
rect 21660 3666 21661 3730
rect 21725 3666 21726 3730
rect 21660 3650 21726 3666
rect 21660 3586 21661 3650
rect 21725 3586 21726 3650
rect 21660 3570 21726 3586
rect 21660 3506 21661 3570
rect 21725 3506 21726 3570
rect 21660 3490 21726 3506
rect 21660 3426 21661 3490
rect 21725 3426 21726 3490
rect 21660 3410 21726 3426
rect 21660 3346 21661 3410
rect 21725 3346 21726 3410
rect 21660 3330 21726 3346
rect 21660 3266 21661 3330
rect 21725 3266 21726 3330
rect 21660 3250 21726 3266
rect 21660 3186 21661 3250
rect 21725 3186 21726 3250
rect 21660 3032 21726 3186
rect 21786 3094 21846 4124
rect 21906 3032 21966 4064
rect 22026 3094 22086 4124
rect 22146 3032 22206 4064
rect 22266 3970 22332 4060
rect 22266 3906 22267 3970
rect 22331 3906 22332 3970
rect 22266 3890 22332 3906
rect 22266 3826 22267 3890
rect 22331 3826 22332 3890
rect 22266 3810 22332 3826
rect 22266 3746 22267 3810
rect 22331 3746 22332 3810
rect 22266 3730 22332 3746
rect 22266 3666 22267 3730
rect 22331 3666 22332 3730
rect 22266 3650 22332 3666
rect 22266 3586 22267 3650
rect 22331 3586 22332 3650
rect 22266 3570 22332 3586
rect 22266 3506 22267 3570
rect 22331 3506 22332 3570
rect 22266 3490 22332 3506
rect 22266 3426 22267 3490
rect 22331 3426 22332 3490
rect 22266 3410 22332 3426
rect 22266 3346 22267 3410
rect 22331 3346 22332 3410
rect 22266 3330 22332 3346
rect 22266 3266 22267 3330
rect 22331 3266 22332 3330
rect 22266 3250 22332 3266
rect 22266 3186 22267 3250
rect 22331 3186 22332 3250
rect 22266 3032 22332 3186
rect 22392 3094 22452 4124
rect 22512 3032 22572 4064
rect 22632 3094 22692 4124
rect 22752 3032 22812 4064
rect 22872 3970 22938 4060
rect 22872 3906 22873 3970
rect 22937 3906 22938 3970
rect 22872 3890 22938 3906
rect 22872 3826 22873 3890
rect 22937 3826 22938 3890
rect 22872 3810 22938 3826
rect 22872 3746 22873 3810
rect 22937 3746 22938 3810
rect 22872 3730 22938 3746
rect 22872 3666 22873 3730
rect 22937 3666 22938 3730
rect 22872 3650 22938 3666
rect 22872 3586 22873 3650
rect 22937 3586 22938 3650
rect 22872 3570 22938 3586
rect 22872 3506 22873 3570
rect 22937 3506 22938 3570
rect 22872 3490 22938 3506
rect 22872 3426 22873 3490
rect 22937 3426 22938 3490
rect 22872 3410 22938 3426
rect 22872 3346 22873 3410
rect 22937 3346 22938 3410
rect 22872 3330 22938 3346
rect 22872 3266 22873 3330
rect 22937 3266 22938 3330
rect 22872 3250 22938 3266
rect 22872 3186 22873 3250
rect 22937 3186 22938 3250
rect 22872 3032 22938 3186
rect 22998 3094 23058 4124
rect 23118 3032 23178 4064
rect 23238 3094 23298 4124
rect 23358 3032 23418 4064
rect 23478 3970 23544 4060
rect 23478 3906 23479 3970
rect 23543 3906 23544 3970
rect 23478 3890 23544 3906
rect 23478 3826 23479 3890
rect 23543 3826 23544 3890
rect 23478 3810 23544 3826
rect 23478 3746 23479 3810
rect 23543 3746 23544 3810
rect 23478 3730 23544 3746
rect 23478 3666 23479 3730
rect 23543 3666 23544 3730
rect 23478 3650 23544 3666
rect 23478 3586 23479 3650
rect 23543 3586 23544 3650
rect 23478 3570 23544 3586
rect 23478 3506 23479 3570
rect 23543 3506 23544 3570
rect 23478 3490 23544 3506
rect 23478 3426 23479 3490
rect 23543 3426 23544 3490
rect 23478 3410 23544 3426
rect 23478 3346 23479 3410
rect 23543 3346 23544 3410
rect 23478 3330 23544 3346
rect 23478 3266 23479 3330
rect 23543 3266 23544 3330
rect 23478 3250 23544 3266
rect 23478 3186 23479 3250
rect 23543 3186 23544 3250
rect 23478 3032 23544 3186
rect 23604 3094 23664 4124
rect 23724 3032 23784 4064
rect 23844 3094 23904 4124
rect 23964 3032 24024 4064
rect 24084 3970 24150 4060
rect 24084 3906 24085 3970
rect 24149 3906 24150 3970
rect 24084 3890 24150 3906
rect 24084 3826 24085 3890
rect 24149 3826 24150 3890
rect 24084 3810 24150 3826
rect 24084 3746 24085 3810
rect 24149 3746 24150 3810
rect 24084 3730 24150 3746
rect 24084 3666 24085 3730
rect 24149 3666 24150 3730
rect 24084 3650 24150 3666
rect 24084 3586 24085 3650
rect 24149 3586 24150 3650
rect 24084 3570 24150 3586
rect 24084 3506 24085 3570
rect 24149 3506 24150 3570
rect 24084 3490 24150 3506
rect 24084 3426 24085 3490
rect 24149 3426 24150 3490
rect 24084 3410 24150 3426
rect 24084 3346 24085 3410
rect 24149 3346 24150 3410
rect 24084 3330 24150 3346
rect 24084 3266 24085 3330
rect 24149 3266 24150 3330
rect 24084 3250 24150 3266
rect 24084 3186 24085 3250
rect 24149 3186 24150 3250
rect 24084 3032 24150 3186
rect 24210 3094 24270 4124
rect 24330 3032 24390 4064
rect 24450 3094 24510 4124
rect 24570 3032 24630 4064
rect 24690 3970 24756 4060
rect 24690 3906 24691 3970
rect 24755 3906 24756 3970
rect 24690 3890 24756 3906
rect 24690 3826 24691 3890
rect 24755 3826 24756 3890
rect 24690 3810 24756 3826
rect 24690 3746 24691 3810
rect 24755 3746 24756 3810
rect 24690 3730 24756 3746
rect 24690 3666 24691 3730
rect 24755 3666 24756 3730
rect 24690 3650 24756 3666
rect 24690 3586 24691 3650
rect 24755 3586 24756 3650
rect 24690 3570 24756 3586
rect 24690 3506 24691 3570
rect 24755 3506 24756 3570
rect 24690 3490 24756 3506
rect 24690 3426 24691 3490
rect 24755 3426 24756 3490
rect 24690 3410 24756 3426
rect 24690 3346 24691 3410
rect 24755 3346 24756 3410
rect 24690 3330 24756 3346
rect 24690 3266 24691 3330
rect 24755 3266 24756 3330
rect 24690 3250 24756 3266
rect 24690 3186 24691 3250
rect 24755 3186 24756 3250
rect 24690 3032 24756 3186
rect 24816 3094 24876 4124
rect 24936 3032 24996 4064
rect 25056 3094 25116 4124
rect 25176 3032 25236 4064
rect 25296 3970 25362 4060
rect 25296 3906 25297 3970
rect 25361 3906 25362 3970
rect 25296 3890 25362 3906
rect 25296 3826 25297 3890
rect 25361 3826 25362 3890
rect 25296 3810 25362 3826
rect 25296 3746 25297 3810
rect 25361 3746 25362 3810
rect 25296 3730 25362 3746
rect 25296 3666 25297 3730
rect 25361 3666 25362 3730
rect 25296 3650 25362 3666
rect 25296 3586 25297 3650
rect 25361 3586 25362 3650
rect 25296 3570 25362 3586
rect 25296 3506 25297 3570
rect 25361 3506 25362 3570
rect 25296 3490 25362 3506
rect 25296 3426 25297 3490
rect 25361 3426 25362 3490
rect 25296 3410 25362 3426
rect 25296 3346 25297 3410
rect 25361 3346 25362 3410
rect 25296 3330 25362 3346
rect 25296 3266 25297 3330
rect 25361 3266 25362 3330
rect 25296 3250 25362 3266
rect 25296 3186 25297 3250
rect 25361 3186 25362 3250
rect 25296 3032 25362 3186
rect 25422 3094 25482 4124
rect 25542 3032 25602 4064
rect 25662 3094 25722 4124
rect 25782 3032 25842 4064
rect 25902 3970 25968 4060
rect 25902 3906 25903 3970
rect 25967 3906 25968 3970
rect 25902 3890 25968 3906
rect 25902 3826 25903 3890
rect 25967 3826 25968 3890
rect 25902 3810 25968 3826
rect 25902 3746 25903 3810
rect 25967 3746 25968 3810
rect 25902 3730 25968 3746
rect 25902 3666 25903 3730
rect 25967 3666 25968 3730
rect 25902 3650 25968 3666
rect 25902 3586 25903 3650
rect 25967 3586 25968 3650
rect 25902 3570 25968 3586
rect 25902 3506 25903 3570
rect 25967 3506 25968 3570
rect 25902 3490 25968 3506
rect 25902 3426 25903 3490
rect 25967 3426 25968 3490
rect 25902 3410 25968 3426
rect 25902 3346 25903 3410
rect 25967 3346 25968 3410
rect 25902 3330 25968 3346
rect 25902 3266 25903 3330
rect 25967 3266 25968 3330
rect 25902 3250 25968 3266
rect 25902 3186 25903 3250
rect 25967 3186 25968 3250
rect 25902 3032 25968 3186
rect 26028 3094 26088 4124
rect 26148 3032 26208 4064
rect 26268 3094 26328 4124
rect 26388 3032 26448 4064
rect 26508 3970 26574 4060
rect 26508 3906 26509 3970
rect 26573 3906 26574 3970
rect 26508 3890 26574 3906
rect 26508 3826 26509 3890
rect 26573 3826 26574 3890
rect 26508 3810 26574 3826
rect 26508 3746 26509 3810
rect 26573 3746 26574 3810
rect 26508 3730 26574 3746
rect 26508 3666 26509 3730
rect 26573 3666 26574 3730
rect 26508 3650 26574 3666
rect 26508 3586 26509 3650
rect 26573 3586 26574 3650
rect 26508 3570 26574 3586
rect 26508 3506 26509 3570
rect 26573 3506 26574 3570
rect 26508 3490 26574 3506
rect 26508 3426 26509 3490
rect 26573 3426 26574 3490
rect 26508 3410 26574 3426
rect 26508 3346 26509 3410
rect 26573 3346 26574 3410
rect 26508 3330 26574 3346
rect 26508 3266 26509 3330
rect 26573 3266 26574 3330
rect 26508 3250 26574 3266
rect 26508 3186 26509 3250
rect 26573 3186 26574 3250
rect 26508 3032 26574 3186
rect 26634 3094 26694 4124
rect 26754 3032 26814 4064
rect 26874 3094 26934 4124
rect 26994 3032 27054 4064
rect 27114 3970 27180 4060
rect 27114 3906 27115 3970
rect 27179 3906 27180 3970
rect 27114 3890 27180 3906
rect 27114 3826 27115 3890
rect 27179 3826 27180 3890
rect 27114 3810 27180 3826
rect 27114 3746 27115 3810
rect 27179 3746 27180 3810
rect 27114 3730 27180 3746
rect 27114 3666 27115 3730
rect 27179 3666 27180 3730
rect 27114 3650 27180 3666
rect 27114 3586 27115 3650
rect 27179 3586 27180 3650
rect 27114 3570 27180 3586
rect 27114 3506 27115 3570
rect 27179 3506 27180 3570
rect 27114 3490 27180 3506
rect 27114 3426 27115 3490
rect 27179 3426 27180 3490
rect 27114 3410 27180 3426
rect 27114 3346 27115 3410
rect 27179 3346 27180 3410
rect 27114 3330 27180 3346
rect 27114 3266 27115 3330
rect 27179 3266 27180 3330
rect 27114 3250 27180 3266
rect 27114 3186 27115 3250
rect 27179 3186 27180 3250
rect 27114 3032 27180 3186
rect 27240 3094 27300 4124
rect 27360 3032 27420 4064
rect 27480 3094 27540 4124
rect 27600 3032 27660 4064
rect 27720 3970 27786 4060
rect 27720 3906 27721 3970
rect 27785 3906 27786 3970
rect 27720 3890 27786 3906
rect 27720 3826 27721 3890
rect 27785 3826 27786 3890
rect 27720 3810 27786 3826
rect 27720 3746 27721 3810
rect 27785 3746 27786 3810
rect 27720 3730 27786 3746
rect 27720 3666 27721 3730
rect 27785 3666 27786 3730
rect 27720 3650 27786 3666
rect 27720 3586 27721 3650
rect 27785 3586 27786 3650
rect 27720 3570 27786 3586
rect 27720 3506 27721 3570
rect 27785 3506 27786 3570
rect 27720 3490 27786 3506
rect 27720 3426 27721 3490
rect 27785 3426 27786 3490
rect 27720 3410 27786 3426
rect 27720 3346 27721 3410
rect 27785 3346 27786 3410
rect 27720 3330 27786 3346
rect 27720 3266 27721 3330
rect 27785 3266 27786 3330
rect 27720 3250 27786 3266
rect 27720 3186 27721 3250
rect 27785 3186 27786 3250
rect 27720 3032 27786 3186
rect 27846 3094 27906 4124
rect 27966 3032 28026 4064
rect 28086 3094 28146 4124
rect 28206 3032 28266 4064
rect 28326 3970 28392 4060
rect 28326 3906 28327 3970
rect 28391 3906 28392 3970
rect 28326 3890 28392 3906
rect 28326 3826 28327 3890
rect 28391 3826 28392 3890
rect 28326 3810 28392 3826
rect 28326 3746 28327 3810
rect 28391 3746 28392 3810
rect 28326 3730 28392 3746
rect 28326 3666 28327 3730
rect 28391 3666 28392 3730
rect 28326 3650 28392 3666
rect 28326 3586 28327 3650
rect 28391 3586 28392 3650
rect 28326 3570 28392 3586
rect 28326 3506 28327 3570
rect 28391 3506 28392 3570
rect 28326 3490 28392 3506
rect 28326 3426 28327 3490
rect 28391 3426 28392 3490
rect 28326 3410 28392 3426
rect 28326 3346 28327 3410
rect 28391 3346 28392 3410
rect 28326 3330 28392 3346
rect 28326 3266 28327 3330
rect 28391 3266 28392 3330
rect 28326 3250 28392 3266
rect 28326 3186 28327 3250
rect 28391 3186 28392 3250
rect 28326 3032 28392 3186
rect 28452 3094 28512 4124
rect 28572 3032 28632 4064
rect 28692 3094 28752 4124
rect 28812 3032 28872 4064
rect 28932 3970 28998 4060
rect 28932 3906 28933 3970
rect 28997 3906 28998 3970
rect 28932 3890 28998 3906
rect 28932 3826 28933 3890
rect 28997 3826 28998 3890
rect 28932 3810 28998 3826
rect 28932 3746 28933 3810
rect 28997 3746 28998 3810
rect 28932 3730 28998 3746
rect 28932 3666 28933 3730
rect 28997 3666 28998 3730
rect 28932 3650 28998 3666
rect 28932 3586 28933 3650
rect 28997 3586 28998 3650
rect 28932 3570 28998 3586
rect 28932 3506 28933 3570
rect 28997 3506 28998 3570
rect 28932 3490 28998 3506
rect 28932 3426 28933 3490
rect 28997 3426 28998 3490
rect 28932 3410 28998 3426
rect 28932 3346 28933 3410
rect 28997 3346 28998 3410
rect 28932 3330 28998 3346
rect 28932 3266 28933 3330
rect 28997 3266 28998 3330
rect 28932 3250 28998 3266
rect 28932 3186 28933 3250
rect 28997 3186 28998 3250
rect 28932 3032 28998 3186
rect 29058 3094 29118 4124
rect 29178 3032 29238 4064
rect 29298 3094 29358 4124
rect 29418 3032 29478 4064
rect 29538 3970 29604 4060
rect 29538 3906 29539 3970
rect 29603 3906 29604 3970
rect 29538 3890 29604 3906
rect 29538 3826 29539 3890
rect 29603 3826 29604 3890
rect 29538 3810 29604 3826
rect 29538 3746 29539 3810
rect 29603 3746 29604 3810
rect 29538 3730 29604 3746
rect 29538 3666 29539 3730
rect 29603 3666 29604 3730
rect 29538 3650 29604 3666
rect 29538 3586 29539 3650
rect 29603 3586 29604 3650
rect 29538 3570 29604 3586
rect 29538 3506 29539 3570
rect 29603 3506 29604 3570
rect 29538 3490 29604 3506
rect 29538 3426 29539 3490
rect 29603 3426 29604 3490
rect 29538 3410 29604 3426
rect 29538 3346 29539 3410
rect 29603 3346 29604 3410
rect 29538 3330 29604 3346
rect 29538 3266 29539 3330
rect 29603 3266 29604 3330
rect 29538 3250 29604 3266
rect 29538 3186 29539 3250
rect 29603 3186 29604 3250
rect 29538 3032 29604 3186
rect 29664 3094 29724 4124
rect 29784 3032 29844 4064
rect 29904 3094 29964 4124
rect 30024 3032 30084 4064
rect 30144 3970 30210 4060
rect 30144 3906 30145 3970
rect 30209 3906 30210 3970
rect 30144 3890 30210 3906
rect 30144 3826 30145 3890
rect 30209 3826 30210 3890
rect 30144 3810 30210 3826
rect 30144 3746 30145 3810
rect 30209 3746 30210 3810
rect 30144 3730 30210 3746
rect 30144 3666 30145 3730
rect 30209 3666 30210 3730
rect 30144 3650 30210 3666
rect 30144 3586 30145 3650
rect 30209 3586 30210 3650
rect 30144 3570 30210 3586
rect 30144 3506 30145 3570
rect 30209 3506 30210 3570
rect 30144 3490 30210 3506
rect 30144 3426 30145 3490
rect 30209 3426 30210 3490
rect 30144 3410 30210 3426
rect 30144 3346 30145 3410
rect 30209 3346 30210 3410
rect 30144 3330 30210 3346
rect 30144 3266 30145 3330
rect 30209 3266 30210 3330
rect 30144 3250 30210 3266
rect 30144 3186 30145 3250
rect 30209 3186 30210 3250
rect 30144 3032 30210 3186
rect 30270 3094 30330 4124
rect 30390 3032 30450 4064
rect 30510 3094 30570 4124
rect 30630 3032 30690 4064
rect 30750 3970 30816 4060
rect 30750 3906 30751 3970
rect 30815 3906 30816 3970
rect 30750 3890 30816 3906
rect 30750 3826 30751 3890
rect 30815 3826 30816 3890
rect 30750 3810 30816 3826
rect 30750 3746 30751 3810
rect 30815 3746 30816 3810
rect 30750 3730 30816 3746
rect 30750 3666 30751 3730
rect 30815 3666 30816 3730
rect 30750 3650 30816 3666
rect 30750 3586 30751 3650
rect 30815 3586 30816 3650
rect 30750 3570 30816 3586
rect 30750 3506 30751 3570
rect 30815 3506 30816 3570
rect 30750 3490 30816 3506
rect 30750 3426 30751 3490
rect 30815 3426 30816 3490
rect 30750 3410 30816 3426
rect 30750 3346 30751 3410
rect 30815 3346 30816 3410
rect 30750 3330 30816 3346
rect 30750 3266 30751 3330
rect 30815 3266 30816 3330
rect 30750 3250 30816 3266
rect 30750 3186 30751 3250
rect 30815 3186 30816 3250
rect 30750 3032 30816 3186
rect 30876 3094 30936 4124
rect 30996 3032 31056 4064
rect 31116 3094 31176 4124
rect 31236 3032 31296 4064
rect 31356 3970 31422 4060
rect 31356 3906 31357 3970
rect 31421 3906 31422 3970
rect 31356 3890 31422 3906
rect 31356 3826 31357 3890
rect 31421 3826 31422 3890
rect 31356 3810 31422 3826
rect 31356 3746 31357 3810
rect 31421 3746 31422 3810
rect 31356 3730 31422 3746
rect 31356 3666 31357 3730
rect 31421 3666 31422 3730
rect 31356 3650 31422 3666
rect 31356 3586 31357 3650
rect 31421 3586 31422 3650
rect 31356 3570 31422 3586
rect 31356 3506 31357 3570
rect 31421 3506 31422 3570
rect 31356 3490 31422 3506
rect 31356 3426 31357 3490
rect 31421 3426 31422 3490
rect 31356 3410 31422 3426
rect 31356 3346 31357 3410
rect 31421 3346 31422 3410
rect 31356 3330 31422 3346
rect 31356 3266 31357 3330
rect 31421 3266 31422 3330
rect 31356 3250 31422 3266
rect 31356 3186 31357 3250
rect 31421 3186 31422 3250
rect 31356 3032 31422 3186
rect 31482 3094 31542 4124
rect 31602 3032 31662 4064
rect 31722 3094 31782 4124
rect 31842 3032 31902 4064
rect 31962 3970 32028 4060
rect 31962 3906 31963 3970
rect 32027 3906 32028 3970
rect 31962 3890 32028 3906
rect 31962 3826 31963 3890
rect 32027 3826 32028 3890
rect 31962 3810 32028 3826
rect 31962 3746 31963 3810
rect 32027 3746 32028 3810
rect 31962 3730 32028 3746
rect 31962 3666 31963 3730
rect 32027 3666 32028 3730
rect 31962 3650 32028 3666
rect 31962 3586 31963 3650
rect 32027 3586 32028 3650
rect 31962 3570 32028 3586
rect 31962 3506 31963 3570
rect 32027 3506 32028 3570
rect 31962 3490 32028 3506
rect 31962 3426 31963 3490
rect 32027 3426 32028 3490
rect 31962 3410 32028 3426
rect 31962 3346 31963 3410
rect 32027 3346 32028 3410
rect 31962 3330 32028 3346
rect 31962 3266 31963 3330
rect 32027 3266 32028 3330
rect 31962 3250 32028 3266
rect 31962 3186 31963 3250
rect 32027 3186 32028 3250
rect 31962 3032 32028 3186
rect 32088 3094 32148 4124
rect 32208 3032 32268 4064
rect 32328 3094 32388 4124
rect 32448 3032 32508 4064
rect 32568 3970 32634 4060
rect 32568 3906 32569 3970
rect 32633 3906 32634 3970
rect 32568 3890 32634 3906
rect 32568 3826 32569 3890
rect 32633 3826 32634 3890
rect 32568 3810 32634 3826
rect 32568 3746 32569 3810
rect 32633 3746 32634 3810
rect 32568 3730 32634 3746
rect 32568 3666 32569 3730
rect 32633 3666 32634 3730
rect 32568 3650 32634 3666
rect 32568 3586 32569 3650
rect 32633 3586 32634 3650
rect 32568 3570 32634 3586
rect 32568 3506 32569 3570
rect 32633 3506 32634 3570
rect 32568 3490 32634 3506
rect 32568 3426 32569 3490
rect 32633 3426 32634 3490
rect 32568 3410 32634 3426
rect 32568 3346 32569 3410
rect 32633 3346 32634 3410
rect 32568 3330 32634 3346
rect 32568 3266 32569 3330
rect 32633 3266 32634 3330
rect 32568 3250 32634 3266
rect 32568 3186 32569 3250
rect 32633 3186 32634 3250
rect 32568 3032 32634 3186
rect 32694 3094 32754 4124
rect 32814 3032 32874 4064
rect 32934 3094 32994 4124
rect 33054 3032 33114 4064
rect 33174 3970 33240 4060
rect 33174 3906 33175 3970
rect 33239 3906 33240 3970
rect 33174 3890 33240 3906
rect 33174 3826 33175 3890
rect 33239 3826 33240 3890
rect 33174 3810 33240 3826
rect 33174 3746 33175 3810
rect 33239 3746 33240 3810
rect 33174 3730 33240 3746
rect 33174 3666 33175 3730
rect 33239 3666 33240 3730
rect 33174 3650 33240 3666
rect 33174 3586 33175 3650
rect 33239 3586 33240 3650
rect 33174 3570 33240 3586
rect 33174 3506 33175 3570
rect 33239 3506 33240 3570
rect 33174 3490 33240 3506
rect 33174 3426 33175 3490
rect 33239 3426 33240 3490
rect 33174 3410 33240 3426
rect 33174 3346 33175 3410
rect 33239 3346 33240 3410
rect 33174 3330 33240 3346
rect 33174 3266 33175 3330
rect 33239 3266 33240 3330
rect 33174 3250 33240 3266
rect 33174 3186 33175 3250
rect 33239 3186 33240 3250
rect 33174 3032 33240 3186
rect 13782 3030 33240 3032
rect 13782 2966 13886 3030
rect 13950 2966 13966 3030
rect 14030 2966 14046 3030
rect 14110 2966 14126 3030
rect 14190 2966 14206 3030
rect 14270 2966 14286 3030
rect 14350 2966 14492 3030
rect 14556 2966 14572 3030
rect 14636 2966 14652 3030
rect 14716 2966 14732 3030
rect 14796 2966 14812 3030
rect 14876 2966 14892 3030
rect 14956 2966 15098 3030
rect 15162 2966 15178 3030
rect 15242 2966 15258 3030
rect 15322 2966 15338 3030
rect 15402 2966 15418 3030
rect 15482 2966 15498 3030
rect 15562 2966 15704 3030
rect 15768 2966 15784 3030
rect 15848 2966 15864 3030
rect 15928 2966 15944 3030
rect 16008 2966 16024 3030
rect 16088 2966 16104 3030
rect 16168 2966 16310 3030
rect 16374 2966 16390 3030
rect 16454 2966 16470 3030
rect 16534 2966 16550 3030
rect 16614 2966 16630 3030
rect 16694 2966 16710 3030
rect 16774 2966 16916 3030
rect 16980 2966 16996 3030
rect 17060 2966 17076 3030
rect 17140 2966 17156 3030
rect 17220 2966 17236 3030
rect 17300 2966 17316 3030
rect 17380 2966 17522 3030
rect 17586 2966 17602 3030
rect 17666 2966 17682 3030
rect 17746 2966 17762 3030
rect 17826 2966 17842 3030
rect 17906 2966 17922 3030
rect 17986 2966 18128 3030
rect 18192 2966 18208 3030
rect 18272 2966 18288 3030
rect 18352 2966 18368 3030
rect 18432 2966 18448 3030
rect 18512 2966 18528 3030
rect 18592 2966 18734 3030
rect 18798 2966 18814 3030
rect 18878 2966 18894 3030
rect 18958 2966 18974 3030
rect 19038 2966 19054 3030
rect 19118 2966 19134 3030
rect 19198 2966 19340 3030
rect 19404 2966 19420 3030
rect 19484 2966 19500 3030
rect 19564 2966 19580 3030
rect 19644 2966 19660 3030
rect 19724 2966 19740 3030
rect 19804 2966 19946 3030
rect 20010 2966 20026 3030
rect 20090 2966 20106 3030
rect 20170 2966 20186 3030
rect 20250 2966 20266 3030
rect 20330 2966 20346 3030
rect 20410 2966 20552 3030
rect 20616 2966 20632 3030
rect 20696 2966 20712 3030
rect 20776 2966 20792 3030
rect 20856 2966 20872 3030
rect 20936 2966 20952 3030
rect 21016 2966 21158 3030
rect 21222 2966 21238 3030
rect 21302 2966 21318 3030
rect 21382 2966 21398 3030
rect 21462 2966 21478 3030
rect 21542 2966 21558 3030
rect 21622 2966 21764 3030
rect 21828 2966 21844 3030
rect 21908 2966 21924 3030
rect 21988 2966 22004 3030
rect 22068 2966 22084 3030
rect 22148 2966 22164 3030
rect 22228 2966 22370 3030
rect 22434 2966 22450 3030
rect 22514 2966 22530 3030
rect 22594 2966 22610 3030
rect 22674 2966 22690 3030
rect 22754 2966 22770 3030
rect 22834 2966 22976 3030
rect 23040 2966 23056 3030
rect 23120 2966 23136 3030
rect 23200 2966 23216 3030
rect 23280 2966 23296 3030
rect 23360 2966 23376 3030
rect 23440 2966 23582 3030
rect 23646 2966 23662 3030
rect 23726 2966 23742 3030
rect 23806 2966 23822 3030
rect 23886 2966 23902 3030
rect 23966 2966 23982 3030
rect 24046 2966 24188 3030
rect 24252 2966 24268 3030
rect 24332 2966 24348 3030
rect 24412 2966 24428 3030
rect 24492 2966 24508 3030
rect 24572 2966 24588 3030
rect 24652 2966 24794 3030
rect 24858 2966 24874 3030
rect 24938 2966 24954 3030
rect 25018 2966 25034 3030
rect 25098 2966 25114 3030
rect 25178 2966 25194 3030
rect 25258 2966 25400 3030
rect 25464 2966 25480 3030
rect 25544 2966 25560 3030
rect 25624 2966 25640 3030
rect 25704 2966 25720 3030
rect 25784 2966 25800 3030
rect 25864 2966 26006 3030
rect 26070 2966 26086 3030
rect 26150 2966 26166 3030
rect 26230 2966 26246 3030
rect 26310 2966 26326 3030
rect 26390 2966 26406 3030
rect 26470 2966 26612 3030
rect 26676 2966 26692 3030
rect 26756 2966 26772 3030
rect 26836 2966 26852 3030
rect 26916 2966 26932 3030
rect 26996 2966 27012 3030
rect 27076 2966 27218 3030
rect 27282 2966 27298 3030
rect 27362 2966 27378 3030
rect 27442 2966 27458 3030
rect 27522 2966 27538 3030
rect 27602 2966 27618 3030
rect 27682 2966 27824 3030
rect 27888 2966 27904 3030
rect 27968 2966 27984 3030
rect 28048 2966 28064 3030
rect 28128 2966 28144 3030
rect 28208 2966 28224 3030
rect 28288 2966 28430 3030
rect 28494 2966 28510 3030
rect 28574 2966 28590 3030
rect 28654 2966 28670 3030
rect 28734 2966 28750 3030
rect 28814 2966 28830 3030
rect 28894 2966 29036 3030
rect 29100 2966 29116 3030
rect 29180 2966 29196 3030
rect 29260 2966 29276 3030
rect 29340 2966 29356 3030
rect 29420 2966 29436 3030
rect 29500 2966 29642 3030
rect 29706 2966 29722 3030
rect 29786 2966 29802 3030
rect 29866 2966 29882 3030
rect 29946 2966 29962 3030
rect 30026 2966 30042 3030
rect 30106 2966 30248 3030
rect 30312 2966 30328 3030
rect 30392 2966 30408 3030
rect 30472 2966 30488 3030
rect 30552 2966 30568 3030
rect 30632 2966 30648 3030
rect 30712 2966 30854 3030
rect 30918 2966 30934 3030
rect 30998 2966 31014 3030
rect 31078 2966 31094 3030
rect 31158 2966 31174 3030
rect 31238 2966 31254 3030
rect 31318 2966 31460 3030
rect 31524 2966 31540 3030
rect 31604 2966 31620 3030
rect 31684 2966 31700 3030
rect 31764 2966 31780 3030
rect 31844 2966 31860 3030
rect 31924 2966 32066 3030
rect 32130 2966 32146 3030
rect 32210 2966 32226 3030
rect 32290 2966 32306 3030
rect 32370 2966 32386 3030
rect 32450 2966 32466 3030
rect 32530 2966 32672 3030
rect 32736 2966 32752 3030
rect 32816 2966 32832 3030
rect 32896 2966 32912 3030
rect 32976 2966 32992 3030
rect 33056 2966 33072 3030
rect 33136 2966 33240 3030
rect 13782 2964 33240 2966
rect 13782 2810 13848 2964
rect 13782 2746 13783 2810
rect 13847 2746 13848 2810
rect 13782 2730 13848 2746
rect 13782 2666 13783 2730
rect 13847 2666 13848 2730
rect 13782 2650 13848 2666
rect 13782 2586 13783 2650
rect 13847 2586 13848 2650
rect 13782 2570 13848 2586
rect 13782 2506 13783 2570
rect 13847 2506 13848 2570
rect 13782 2490 13848 2506
rect 13782 2426 13783 2490
rect 13847 2426 13848 2490
rect 13782 2410 13848 2426
rect 13782 2346 13783 2410
rect 13847 2346 13848 2410
rect 13782 2330 13848 2346
rect 13782 2266 13783 2330
rect 13847 2266 13848 2330
rect 13782 2250 13848 2266
rect 13782 2186 13783 2250
rect 13847 2186 13848 2250
rect 13782 2170 13848 2186
rect 13782 2106 13783 2170
rect 13847 2106 13848 2170
rect 13782 2090 13848 2106
rect 13782 2026 13783 2090
rect 13847 2026 13848 2090
rect 13782 1936 13848 2026
rect 13908 1932 13968 2964
rect 14028 1872 14088 2902
rect 14148 1932 14208 2964
rect 14268 1872 14328 2902
rect 14388 2810 14454 2964
rect 14388 2746 14389 2810
rect 14453 2746 14454 2810
rect 14388 2730 14454 2746
rect 14388 2666 14389 2730
rect 14453 2666 14454 2730
rect 14388 2650 14454 2666
rect 14388 2586 14389 2650
rect 14453 2586 14454 2650
rect 14388 2570 14454 2586
rect 14388 2506 14389 2570
rect 14453 2506 14454 2570
rect 14388 2490 14454 2506
rect 14388 2426 14389 2490
rect 14453 2426 14454 2490
rect 14388 2410 14454 2426
rect 14388 2346 14389 2410
rect 14453 2346 14454 2410
rect 14388 2330 14454 2346
rect 14388 2266 14389 2330
rect 14453 2266 14454 2330
rect 14388 2250 14454 2266
rect 14388 2186 14389 2250
rect 14453 2186 14454 2250
rect 14388 2170 14454 2186
rect 14388 2106 14389 2170
rect 14453 2106 14454 2170
rect 14388 2090 14454 2106
rect 14388 2026 14389 2090
rect 14453 2026 14454 2090
rect 14388 1936 14454 2026
rect 14514 1932 14574 2964
rect 14634 1872 14694 2902
rect 14754 1932 14814 2964
rect 14874 1872 14934 2902
rect 14994 2810 15060 2964
rect 14994 2746 14995 2810
rect 15059 2746 15060 2810
rect 14994 2730 15060 2746
rect 14994 2666 14995 2730
rect 15059 2666 15060 2730
rect 14994 2650 15060 2666
rect 14994 2586 14995 2650
rect 15059 2586 15060 2650
rect 14994 2570 15060 2586
rect 14994 2506 14995 2570
rect 15059 2506 15060 2570
rect 14994 2490 15060 2506
rect 14994 2426 14995 2490
rect 15059 2426 15060 2490
rect 14994 2410 15060 2426
rect 14994 2346 14995 2410
rect 15059 2346 15060 2410
rect 14994 2330 15060 2346
rect 14994 2266 14995 2330
rect 15059 2266 15060 2330
rect 14994 2250 15060 2266
rect 14994 2186 14995 2250
rect 15059 2186 15060 2250
rect 14994 2170 15060 2186
rect 14994 2106 14995 2170
rect 15059 2106 15060 2170
rect 14994 2090 15060 2106
rect 14994 2026 14995 2090
rect 15059 2026 15060 2090
rect 14994 1936 15060 2026
rect 15120 1932 15180 2964
rect 15240 1872 15300 2902
rect 15360 1932 15420 2964
rect 15480 1872 15540 2902
rect 15600 2810 15666 2964
rect 15600 2746 15601 2810
rect 15665 2746 15666 2810
rect 15600 2730 15666 2746
rect 15600 2666 15601 2730
rect 15665 2666 15666 2730
rect 15600 2650 15666 2666
rect 15600 2586 15601 2650
rect 15665 2586 15666 2650
rect 15600 2570 15666 2586
rect 15600 2506 15601 2570
rect 15665 2506 15666 2570
rect 15600 2490 15666 2506
rect 15600 2426 15601 2490
rect 15665 2426 15666 2490
rect 15600 2410 15666 2426
rect 15600 2346 15601 2410
rect 15665 2346 15666 2410
rect 15600 2330 15666 2346
rect 15600 2266 15601 2330
rect 15665 2266 15666 2330
rect 15600 2250 15666 2266
rect 15600 2186 15601 2250
rect 15665 2186 15666 2250
rect 15600 2170 15666 2186
rect 15600 2106 15601 2170
rect 15665 2106 15666 2170
rect 15600 2090 15666 2106
rect 15600 2026 15601 2090
rect 15665 2026 15666 2090
rect 15600 1936 15666 2026
rect 15726 1932 15786 2964
rect 15846 1872 15906 2902
rect 15966 1932 16026 2964
rect 16086 1872 16146 2902
rect 16206 2810 16272 2964
rect 16206 2746 16207 2810
rect 16271 2746 16272 2810
rect 16206 2730 16272 2746
rect 16206 2666 16207 2730
rect 16271 2666 16272 2730
rect 16206 2650 16272 2666
rect 16206 2586 16207 2650
rect 16271 2586 16272 2650
rect 16206 2570 16272 2586
rect 16206 2506 16207 2570
rect 16271 2506 16272 2570
rect 16206 2490 16272 2506
rect 16206 2426 16207 2490
rect 16271 2426 16272 2490
rect 16206 2410 16272 2426
rect 16206 2346 16207 2410
rect 16271 2346 16272 2410
rect 16206 2330 16272 2346
rect 16206 2266 16207 2330
rect 16271 2266 16272 2330
rect 16206 2250 16272 2266
rect 16206 2186 16207 2250
rect 16271 2186 16272 2250
rect 16206 2170 16272 2186
rect 16206 2106 16207 2170
rect 16271 2106 16272 2170
rect 16206 2090 16272 2106
rect 16206 2026 16207 2090
rect 16271 2026 16272 2090
rect 16206 1936 16272 2026
rect 16332 1932 16392 2964
rect 16452 1872 16512 2902
rect 16572 1932 16632 2964
rect 16692 1872 16752 2902
rect 16812 2810 16878 2964
rect 16812 2746 16813 2810
rect 16877 2746 16878 2810
rect 16812 2730 16878 2746
rect 16812 2666 16813 2730
rect 16877 2666 16878 2730
rect 16812 2650 16878 2666
rect 16812 2586 16813 2650
rect 16877 2586 16878 2650
rect 16812 2570 16878 2586
rect 16812 2506 16813 2570
rect 16877 2506 16878 2570
rect 16812 2490 16878 2506
rect 16812 2426 16813 2490
rect 16877 2426 16878 2490
rect 16812 2410 16878 2426
rect 16812 2346 16813 2410
rect 16877 2346 16878 2410
rect 16812 2330 16878 2346
rect 16812 2266 16813 2330
rect 16877 2266 16878 2330
rect 16812 2250 16878 2266
rect 16812 2186 16813 2250
rect 16877 2186 16878 2250
rect 16812 2170 16878 2186
rect 16812 2106 16813 2170
rect 16877 2106 16878 2170
rect 16812 2090 16878 2106
rect 16812 2026 16813 2090
rect 16877 2026 16878 2090
rect 16812 1936 16878 2026
rect 16938 1932 16998 2964
rect 17058 1872 17118 2902
rect 17178 1932 17238 2964
rect 17298 1872 17358 2902
rect 17418 2810 17484 2964
rect 17418 2746 17419 2810
rect 17483 2746 17484 2810
rect 17418 2730 17484 2746
rect 17418 2666 17419 2730
rect 17483 2666 17484 2730
rect 17418 2650 17484 2666
rect 17418 2586 17419 2650
rect 17483 2586 17484 2650
rect 17418 2570 17484 2586
rect 17418 2506 17419 2570
rect 17483 2506 17484 2570
rect 17418 2490 17484 2506
rect 17418 2426 17419 2490
rect 17483 2426 17484 2490
rect 17418 2410 17484 2426
rect 17418 2346 17419 2410
rect 17483 2346 17484 2410
rect 17418 2330 17484 2346
rect 17418 2266 17419 2330
rect 17483 2266 17484 2330
rect 17418 2250 17484 2266
rect 17418 2186 17419 2250
rect 17483 2186 17484 2250
rect 17418 2170 17484 2186
rect 17418 2106 17419 2170
rect 17483 2106 17484 2170
rect 17418 2090 17484 2106
rect 17418 2026 17419 2090
rect 17483 2026 17484 2090
rect 17418 1936 17484 2026
rect 17544 1932 17604 2964
rect 17664 1872 17724 2902
rect 17784 1932 17844 2964
rect 17904 1872 17964 2902
rect 18024 2810 18090 2964
rect 18024 2746 18025 2810
rect 18089 2746 18090 2810
rect 18024 2730 18090 2746
rect 18024 2666 18025 2730
rect 18089 2666 18090 2730
rect 18024 2650 18090 2666
rect 18024 2586 18025 2650
rect 18089 2586 18090 2650
rect 18024 2570 18090 2586
rect 18024 2506 18025 2570
rect 18089 2506 18090 2570
rect 18024 2490 18090 2506
rect 18024 2426 18025 2490
rect 18089 2426 18090 2490
rect 18024 2410 18090 2426
rect 18024 2346 18025 2410
rect 18089 2346 18090 2410
rect 18024 2330 18090 2346
rect 18024 2266 18025 2330
rect 18089 2266 18090 2330
rect 18024 2250 18090 2266
rect 18024 2186 18025 2250
rect 18089 2186 18090 2250
rect 18024 2170 18090 2186
rect 18024 2106 18025 2170
rect 18089 2106 18090 2170
rect 18024 2090 18090 2106
rect 18024 2026 18025 2090
rect 18089 2026 18090 2090
rect 18024 1936 18090 2026
rect 18150 1932 18210 2964
rect 18270 1872 18330 2902
rect 18390 1932 18450 2964
rect 18510 1872 18570 2902
rect 18630 2810 18696 2964
rect 18630 2746 18631 2810
rect 18695 2746 18696 2810
rect 18630 2730 18696 2746
rect 18630 2666 18631 2730
rect 18695 2666 18696 2730
rect 18630 2650 18696 2666
rect 18630 2586 18631 2650
rect 18695 2586 18696 2650
rect 18630 2570 18696 2586
rect 18630 2506 18631 2570
rect 18695 2506 18696 2570
rect 18630 2490 18696 2506
rect 18630 2426 18631 2490
rect 18695 2426 18696 2490
rect 18630 2410 18696 2426
rect 18630 2346 18631 2410
rect 18695 2346 18696 2410
rect 18630 2330 18696 2346
rect 18630 2266 18631 2330
rect 18695 2266 18696 2330
rect 18630 2250 18696 2266
rect 18630 2186 18631 2250
rect 18695 2186 18696 2250
rect 18630 2170 18696 2186
rect 18630 2106 18631 2170
rect 18695 2106 18696 2170
rect 18630 2090 18696 2106
rect 18630 2026 18631 2090
rect 18695 2026 18696 2090
rect 18630 1936 18696 2026
rect 18756 1932 18816 2964
rect 18876 1872 18936 2902
rect 18996 1932 19056 2964
rect 19116 1872 19176 2902
rect 19236 2810 19302 2964
rect 19236 2746 19237 2810
rect 19301 2746 19302 2810
rect 19236 2730 19302 2746
rect 19236 2666 19237 2730
rect 19301 2666 19302 2730
rect 19236 2650 19302 2666
rect 19236 2586 19237 2650
rect 19301 2586 19302 2650
rect 19236 2570 19302 2586
rect 19236 2506 19237 2570
rect 19301 2506 19302 2570
rect 19236 2490 19302 2506
rect 19236 2426 19237 2490
rect 19301 2426 19302 2490
rect 19236 2410 19302 2426
rect 19236 2346 19237 2410
rect 19301 2346 19302 2410
rect 19236 2330 19302 2346
rect 19236 2266 19237 2330
rect 19301 2266 19302 2330
rect 19236 2250 19302 2266
rect 19236 2186 19237 2250
rect 19301 2186 19302 2250
rect 19236 2170 19302 2186
rect 19236 2106 19237 2170
rect 19301 2106 19302 2170
rect 19236 2090 19302 2106
rect 19236 2026 19237 2090
rect 19301 2026 19302 2090
rect 19236 1936 19302 2026
rect 19362 1932 19422 2964
rect 19482 1872 19542 2902
rect 19602 1932 19662 2964
rect 19722 1872 19782 2902
rect 19842 2810 19908 2964
rect 19842 2746 19843 2810
rect 19907 2746 19908 2810
rect 19842 2730 19908 2746
rect 19842 2666 19843 2730
rect 19907 2666 19908 2730
rect 19842 2650 19908 2666
rect 19842 2586 19843 2650
rect 19907 2586 19908 2650
rect 19842 2570 19908 2586
rect 19842 2506 19843 2570
rect 19907 2506 19908 2570
rect 19842 2490 19908 2506
rect 19842 2426 19843 2490
rect 19907 2426 19908 2490
rect 19842 2410 19908 2426
rect 19842 2346 19843 2410
rect 19907 2346 19908 2410
rect 19842 2330 19908 2346
rect 19842 2266 19843 2330
rect 19907 2266 19908 2330
rect 19842 2250 19908 2266
rect 19842 2186 19843 2250
rect 19907 2186 19908 2250
rect 19842 2170 19908 2186
rect 19842 2106 19843 2170
rect 19907 2106 19908 2170
rect 19842 2090 19908 2106
rect 19842 2026 19843 2090
rect 19907 2026 19908 2090
rect 19842 1936 19908 2026
rect 19968 1932 20028 2964
rect 20088 1872 20148 2902
rect 20208 1932 20268 2964
rect 20328 1872 20388 2902
rect 20448 2810 20514 2964
rect 20448 2746 20449 2810
rect 20513 2746 20514 2810
rect 20448 2730 20514 2746
rect 20448 2666 20449 2730
rect 20513 2666 20514 2730
rect 20448 2650 20514 2666
rect 20448 2586 20449 2650
rect 20513 2586 20514 2650
rect 20448 2570 20514 2586
rect 20448 2506 20449 2570
rect 20513 2506 20514 2570
rect 20448 2490 20514 2506
rect 20448 2426 20449 2490
rect 20513 2426 20514 2490
rect 20448 2410 20514 2426
rect 20448 2346 20449 2410
rect 20513 2346 20514 2410
rect 20448 2330 20514 2346
rect 20448 2266 20449 2330
rect 20513 2266 20514 2330
rect 20448 2250 20514 2266
rect 20448 2186 20449 2250
rect 20513 2186 20514 2250
rect 20448 2170 20514 2186
rect 20448 2106 20449 2170
rect 20513 2106 20514 2170
rect 20448 2090 20514 2106
rect 20448 2026 20449 2090
rect 20513 2026 20514 2090
rect 20448 1936 20514 2026
rect 20574 1932 20634 2964
rect 20694 1872 20754 2902
rect 20814 1932 20874 2964
rect 20934 1872 20994 2902
rect 21054 2810 21120 2964
rect 21054 2746 21055 2810
rect 21119 2746 21120 2810
rect 21054 2730 21120 2746
rect 21054 2666 21055 2730
rect 21119 2666 21120 2730
rect 21054 2650 21120 2666
rect 21054 2586 21055 2650
rect 21119 2586 21120 2650
rect 21054 2570 21120 2586
rect 21054 2506 21055 2570
rect 21119 2506 21120 2570
rect 21054 2490 21120 2506
rect 21054 2426 21055 2490
rect 21119 2426 21120 2490
rect 21054 2410 21120 2426
rect 21054 2346 21055 2410
rect 21119 2346 21120 2410
rect 21054 2330 21120 2346
rect 21054 2266 21055 2330
rect 21119 2266 21120 2330
rect 21054 2250 21120 2266
rect 21054 2186 21055 2250
rect 21119 2186 21120 2250
rect 21054 2170 21120 2186
rect 21054 2106 21055 2170
rect 21119 2106 21120 2170
rect 21054 2090 21120 2106
rect 21054 2026 21055 2090
rect 21119 2026 21120 2090
rect 21054 1936 21120 2026
rect 21180 1932 21240 2964
rect 21300 1872 21360 2902
rect 21420 1932 21480 2964
rect 21540 1872 21600 2902
rect 21660 2810 21726 2964
rect 21660 2746 21661 2810
rect 21725 2746 21726 2810
rect 21660 2730 21726 2746
rect 21660 2666 21661 2730
rect 21725 2666 21726 2730
rect 21660 2650 21726 2666
rect 21660 2586 21661 2650
rect 21725 2586 21726 2650
rect 21660 2570 21726 2586
rect 21660 2506 21661 2570
rect 21725 2506 21726 2570
rect 21660 2490 21726 2506
rect 21660 2426 21661 2490
rect 21725 2426 21726 2490
rect 21660 2410 21726 2426
rect 21660 2346 21661 2410
rect 21725 2346 21726 2410
rect 21660 2330 21726 2346
rect 21660 2266 21661 2330
rect 21725 2266 21726 2330
rect 21660 2250 21726 2266
rect 21660 2186 21661 2250
rect 21725 2186 21726 2250
rect 21660 2170 21726 2186
rect 21660 2106 21661 2170
rect 21725 2106 21726 2170
rect 21660 2090 21726 2106
rect 21660 2026 21661 2090
rect 21725 2026 21726 2090
rect 21660 1936 21726 2026
rect 21786 1932 21846 2964
rect 21906 1872 21966 2902
rect 22026 1932 22086 2964
rect 22146 1872 22206 2902
rect 22266 2810 22332 2964
rect 22266 2746 22267 2810
rect 22331 2746 22332 2810
rect 22266 2730 22332 2746
rect 22266 2666 22267 2730
rect 22331 2666 22332 2730
rect 22266 2650 22332 2666
rect 22266 2586 22267 2650
rect 22331 2586 22332 2650
rect 22266 2570 22332 2586
rect 22266 2506 22267 2570
rect 22331 2506 22332 2570
rect 22266 2490 22332 2506
rect 22266 2426 22267 2490
rect 22331 2426 22332 2490
rect 22266 2410 22332 2426
rect 22266 2346 22267 2410
rect 22331 2346 22332 2410
rect 22266 2330 22332 2346
rect 22266 2266 22267 2330
rect 22331 2266 22332 2330
rect 22266 2250 22332 2266
rect 22266 2186 22267 2250
rect 22331 2186 22332 2250
rect 22266 2170 22332 2186
rect 22266 2106 22267 2170
rect 22331 2106 22332 2170
rect 22266 2090 22332 2106
rect 22266 2026 22267 2090
rect 22331 2026 22332 2090
rect 22266 1936 22332 2026
rect 22392 1932 22452 2964
rect 22512 1872 22572 2902
rect 22632 1932 22692 2964
rect 22752 1872 22812 2902
rect 22872 2810 22938 2964
rect 22872 2746 22873 2810
rect 22937 2746 22938 2810
rect 22872 2730 22938 2746
rect 22872 2666 22873 2730
rect 22937 2666 22938 2730
rect 22872 2650 22938 2666
rect 22872 2586 22873 2650
rect 22937 2586 22938 2650
rect 22872 2570 22938 2586
rect 22872 2506 22873 2570
rect 22937 2506 22938 2570
rect 22872 2490 22938 2506
rect 22872 2426 22873 2490
rect 22937 2426 22938 2490
rect 22872 2410 22938 2426
rect 22872 2346 22873 2410
rect 22937 2346 22938 2410
rect 22872 2330 22938 2346
rect 22872 2266 22873 2330
rect 22937 2266 22938 2330
rect 22872 2250 22938 2266
rect 22872 2186 22873 2250
rect 22937 2186 22938 2250
rect 22872 2170 22938 2186
rect 22872 2106 22873 2170
rect 22937 2106 22938 2170
rect 22872 2090 22938 2106
rect 22872 2026 22873 2090
rect 22937 2026 22938 2090
rect 22872 1936 22938 2026
rect 22998 1932 23058 2964
rect 23118 1872 23178 2902
rect 23238 1932 23298 2964
rect 23358 1872 23418 2902
rect 23478 2810 23544 2964
rect 23478 2746 23479 2810
rect 23543 2746 23544 2810
rect 23478 2730 23544 2746
rect 23478 2666 23479 2730
rect 23543 2666 23544 2730
rect 23478 2650 23544 2666
rect 23478 2586 23479 2650
rect 23543 2586 23544 2650
rect 23478 2570 23544 2586
rect 23478 2506 23479 2570
rect 23543 2506 23544 2570
rect 23478 2490 23544 2506
rect 23478 2426 23479 2490
rect 23543 2426 23544 2490
rect 23478 2410 23544 2426
rect 23478 2346 23479 2410
rect 23543 2346 23544 2410
rect 23478 2330 23544 2346
rect 23478 2266 23479 2330
rect 23543 2266 23544 2330
rect 23478 2250 23544 2266
rect 23478 2186 23479 2250
rect 23543 2186 23544 2250
rect 23478 2170 23544 2186
rect 23478 2106 23479 2170
rect 23543 2106 23544 2170
rect 23478 2090 23544 2106
rect 23478 2026 23479 2090
rect 23543 2026 23544 2090
rect 23478 1936 23544 2026
rect 23604 1932 23664 2964
rect 23724 1872 23784 2902
rect 23844 1932 23904 2964
rect 23964 1872 24024 2902
rect 24084 2810 24150 2964
rect 24084 2746 24085 2810
rect 24149 2746 24150 2810
rect 24084 2730 24150 2746
rect 24084 2666 24085 2730
rect 24149 2666 24150 2730
rect 24084 2650 24150 2666
rect 24084 2586 24085 2650
rect 24149 2586 24150 2650
rect 24084 2570 24150 2586
rect 24084 2506 24085 2570
rect 24149 2506 24150 2570
rect 24084 2490 24150 2506
rect 24084 2426 24085 2490
rect 24149 2426 24150 2490
rect 24084 2410 24150 2426
rect 24084 2346 24085 2410
rect 24149 2346 24150 2410
rect 24084 2330 24150 2346
rect 24084 2266 24085 2330
rect 24149 2266 24150 2330
rect 24084 2250 24150 2266
rect 24084 2186 24085 2250
rect 24149 2186 24150 2250
rect 24084 2170 24150 2186
rect 24084 2106 24085 2170
rect 24149 2106 24150 2170
rect 24084 2090 24150 2106
rect 24084 2026 24085 2090
rect 24149 2026 24150 2090
rect 24084 1936 24150 2026
rect 24210 1932 24270 2964
rect 24330 1872 24390 2902
rect 24450 1932 24510 2964
rect 24570 1872 24630 2902
rect 24690 2810 24756 2964
rect 24690 2746 24691 2810
rect 24755 2746 24756 2810
rect 24690 2730 24756 2746
rect 24690 2666 24691 2730
rect 24755 2666 24756 2730
rect 24690 2650 24756 2666
rect 24690 2586 24691 2650
rect 24755 2586 24756 2650
rect 24690 2570 24756 2586
rect 24690 2506 24691 2570
rect 24755 2506 24756 2570
rect 24690 2490 24756 2506
rect 24690 2426 24691 2490
rect 24755 2426 24756 2490
rect 24690 2410 24756 2426
rect 24690 2346 24691 2410
rect 24755 2346 24756 2410
rect 24690 2330 24756 2346
rect 24690 2266 24691 2330
rect 24755 2266 24756 2330
rect 24690 2250 24756 2266
rect 24690 2186 24691 2250
rect 24755 2186 24756 2250
rect 24690 2170 24756 2186
rect 24690 2106 24691 2170
rect 24755 2106 24756 2170
rect 24690 2090 24756 2106
rect 24690 2026 24691 2090
rect 24755 2026 24756 2090
rect 24690 1936 24756 2026
rect 24816 1932 24876 2964
rect 24936 1872 24996 2902
rect 25056 1932 25116 2964
rect 25176 1872 25236 2902
rect 25296 2810 25362 2964
rect 25296 2746 25297 2810
rect 25361 2746 25362 2810
rect 25296 2730 25362 2746
rect 25296 2666 25297 2730
rect 25361 2666 25362 2730
rect 25296 2650 25362 2666
rect 25296 2586 25297 2650
rect 25361 2586 25362 2650
rect 25296 2570 25362 2586
rect 25296 2506 25297 2570
rect 25361 2506 25362 2570
rect 25296 2490 25362 2506
rect 25296 2426 25297 2490
rect 25361 2426 25362 2490
rect 25296 2410 25362 2426
rect 25296 2346 25297 2410
rect 25361 2346 25362 2410
rect 25296 2330 25362 2346
rect 25296 2266 25297 2330
rect 25361 2266 25362 2330
rect 25296 2250 25362 2266
rect 25296 2186 25297 2250
rect 25361 2186 25362 2250
rect 25296 2170 25362 2186
rect 25296 2106 25297 2170
rect 25361 2106 25362 2170
rect 25296 2090 25362 2106
rect 25296 2026 25297 2090
rect 25361 2026 25362 2090
rect 25296 1936 25362 2026
rect 25422 1932 25482 2964
rect 25542 1872 25602 2902
rect 25662 1932 25722 2964
rect 25782 1872 25842 2902
rect 25902 2810 25968 2964
rect 25902 2746 25903 2810
rect 25967 2746 25968 2810
rect 25902 2730 25968 2746
rect 25902 2666 25903 2730
rect 25967 2666 25968 2730
rect 25902 2650 25968 2666
rect 25902 2586 25903 2650
rect 25967 2586 25968 2650
rect 25902 2570 25968 2586
rect 25902 2506 25903 2570
rect 25967 2506 25968 2570
rect 25902 2490 25968 2506
rect 25902 2426 25903 2490
rect 25967 2426 25968 2490
rect 25902 2410 25968 2426
rect 25902 2346 25903 2410
rect 25967 2346 25968 2410
rect 25902 2330 25968 2346
rect 25902 2266 25903 2330
rect 25967 2266 25968 2330
rect 25902 2250 25968 2266
rect 25902 2186 25903 2250
rect 25967 2186 25968 2250
rect 25902 2170 25968 2186
rect 25902 2106 25903 2170
rect 25967 2106 25968 2170
rect 25902 2090 25968 2106
rect 25902 2026 25903 2090
rect 25967 2026 25968 2090
rect 25902 1936 25968 2026
rect 26028 1932 26088 2964
rect 26148 1872 26208 2902
rect 26268 1932 26328 2964
rect 26388 1872 26448 2902
rect 26508 2810 26574 2964
rect 26508 2746 26509 2810
rect 26573 2746 26574 2810
rect 26508 2730 26574 2746
rect 26508 2666 26509 2730
rect 26573 2666 26574 2730
rect 26508 2650 26574 2666
rect 26508 2586 26509 2650
rect 26573 2586 26574 2650
rect 26508 2570 26574 2586
rect 26508 2506 26509 2570
rect 26573 2506 26574 2570
rect 26508 2490 26574 2506
rect 26508 2426 26509 2490
rect 26573 2426 26574 2490
rect 26508 2410 26574 2426
rect 26508 2346 26509 2410
rect 26573 2346 26574 2410
rect 26508 2330 26574 2346
rect 26508 2266 26509 2330
rect 26573 2266 26574 2330
rect 26508 2250 26574 2266
rect 26508 2186 26509 2250
rect 26573 2186 26574 2250
rect 26508 2170 26574 2186
rect 26508 2106 26509 2170
rect 26573 2106 26574 2170
rect 26508 2090 26574 2106
rect 26508 2026 26509 2090
rect 26573 2026 26574 2090
rect 26508 1936 26574 2026
rect 26634 1932 26694 2964
rect 26754 1872 26814 2902
rect 26874 1932 26934 2964
rect 26994 1872 27054 2902
rect 27114 2810 27180 2964
rect 27114 2746 27115 2810
rect 27179 2746 27180 2810
rect 27114 2730 27180 2746
rect 27114 2666 27115 2730
rect 27179 2666 27180 2730
rect 27114 2650 27180 2666
rect 27114 2586 27115 2650
rect 27179 2586 27180 2650
rect 27114 2570 27180 2586
rect 27114 2506 27115 2570
rect 27179 2506 27180 2570
rect 27114 2490 27180 2506
rect 27114 2426 27115 2490
rect 27179 2426 27180 2490
rect 27114 2410 27180 2426
rect 27114 2346 27115 2410
rect 27179 2346 27180 2410
rect 27114 2330 27180 2346
rect 27114 2266 27115 2330
rect 27179 2266 27180 2330
rect 27114 2250 27180 2266
rect 27114 2186 27115 2250
rect 27179 2186 27180 2250
rect 27114 2170 27180 2186
rect 27114 2106 27115 2170
rect 27179 2106 27180 2170
rect 27114 2090 27180 2106
rect 27114 2026 27115 2090
rect 27179 2026 27180 2090
rect 27114 1936 27180 2026
rect 27240 1932 27300 2964
rect 27360 1872 27420 2902
rect 27480 1932 27540 2964
rect 27600 1872 27660 2902
rect 27720 2810 27786 2964
rect 27720 2746 27721 2810
rect 27785 2746 27786 2810
rect 27720 2730 27786 2746
rect 27720 2666 27721 2730
rect 27785 2666 27786 2730
rect 27720 2650 27786 2666
rect 27720 2586 27721 2650
rect 27785 2586 27786 2650
rect 27720 2570 27786 2586
rect 27720 2506 27721 2570
rect 27785 2506 27786 2570
rect 27720 2490 27786 2506
rect 27720 2426 27721 2490
rect 27785 2426 27786 2490
rect 27720 2410 27786 2426
rect 27720 2346 27721 2410
rect 27785 2346 27786 2410
rect 27720 2330 27786 2346
rect 27720 2266 27721 2330
rect 27785 2266 27786 2330
rect 27720 2250 27786 2266
rect 27720 2186 27721 2250
rect 27785 2186 27786 2250
rect 27720 2170 27786 2186
rect 27720 2106 27721 2170
rect 27785 2106 27786 2170
rect 27720 2090 27786 2106
rect 27720 2026 27721 2090
rect 27785 2026 27786 2090
rect 27720 1936 27786 2026
rect 27846 1932 27906 2964
rect 27966 1872 28026 2902
rect 28086 1932 28146 2964
rect 28206 1872 28266 2902
rect 28326 2810 28392 2964
rect 28326 2746 28327 2810
rect 28391 2746 28392 2810
rect 28326 2730 28392 2746
rect 28326 2666 28327 2730
rect 28391 2666 28392 2730
rect 28326 2650 28392 2666
rect 28326 2586 28327 2650
rect 28391 2586 28392 2650
rect 28326 2570 28392 2586
rect 28326 2506 28327 2570
rect 28391 2506 28392 2570
rect 28326 2490 28392 2506
rect 28326 2426 28327 2490
rect 28391 2426 28392 2490
rect 28326 2410 28392 2426
rect 28326 2346 28327 2410
rect 28391 2346 28392 2410
rect 28326 2330 28392 2346
rect 28326 2266 28327 2330
rect 28391 2266 28392 2330
rect 28326 2250 28392 2266
rect 28326 2186 28327 2250
rect 28391 2186 28392 2250
rect 28326 2170 28392 2186
rect 28326 2106 28327 2170
rect 28391 2106 28392 2170
rect 28326 2090 28392 2106
rect 28326 2026 28327 2090
rect 28391 2026 28392 2090
rect 28326 1936 28392 2026
rect 28452 1932 28512 2964
rect 28572 1872 28632 2902
rect 28692 1932 28752 2964
rect 28812 1872 28872 2902
rect 28932 2810 28998 2964
rect 28932 2746 28933 2810
rect 28997 2746 28998 2810
rect 28932 2730 28998 2746
rect 28932 2666 28933 2730
rect 28997 2666 28998 2730
rect 28932 2650 28998 2666
rect 28932 2586 28933 2650
rect 28997 2586 28998 2650
rect 28932 2570 28998 2586
rect 28932 2506 28933 2570
rect 28997 2506 28998 2570
rect 28932 2490 28998 2506
rect 28932 2426 28933 2490
rect 28997 2426 28998 2490
rect 28932 2410 28998 2426
rect 28932 2346 28933 2410
rect 28997 2346 28998 2410
rect 28932 2330 28998 2346
rect 28932 2266 28933 2330
rect 28997 2266 28998 2330
rect 28932 2250 28998 2266
rect 28932 2186 28933 2250
rect 28997 2186 28998 2250
rect 28932 2170 28998 2186
rect 28932 2106 28933 2170
rect 28997 2106 28998 2170
rect 28932 2090 28998 2106
rect 28932 2026 28933 2090
rect 28997 2026 28998 2090
rect 28932 1936 28998 2026
rect 29058 1932 29118 2964
rect 29178 1872 29238 2902
rect 29298 1932 29358 2964
rect 29418 1872 29478 2902
rect 29538 2810 29604 2964
rect 29538 2746 29539 2810
rect 29603 2746 29604 2810
rect 29538 2730 29604 2746
rect 29538 2666 29539 2730
rect 29603 2666 29604 2730
rect 29538 2650 29604 2666
rect 29538 2586 29539 2650
rect 29603 2586 29604 2650
rect 29538 2570 29604 2586
rect 29538 2506 29539 2570
rect 29603 2506 29604 2570
rect 29538 2490 29604 2506
rect 29538 2426 29539 2490
rect 29603 2426 29604 2490
rect 29538 2410 29604 2426
rect 29538 2346 29539 2410
rect 29603 2346 29604 2410
rect 29538 2330 29604 2346
rect 29538 2266 29539 2330
rect 29603 2266 29604 2330
rect 29538 2250 29604 2266
rect 29538 2186 29539 2250
rect 29603 2186 29604 2250
rect 29538 2170 29604 2186
rect 29538 2106 29539 2170
rect 29603 2106 29604 2170
rect 29538 2090 29604 2106
rect 29538 2026 29539 2090
rect 29603 2026 29604 2090
rect 29538 1936 29604 2026
rect 29664 1932 29724 2964
rect 29784 1872 29844 2902
rect 29904 1932 29964 2964
rect 30024 1872 30084 2902
rect 30144 2810 30210 2964
rect 30144 2746 30145 2810
rect 30209 2746 30210 2810
rect 30144 2730 30210 2746
rect 30144 2666 30145 2730
rect 30209 2666 30210 2730
rect 30144 2650 30210 2666
rect 30144 2586 30145 2650
rect 30209 2586 30210 2650
rect 30144 2570 30210 2586
rect 30144 2506 30145 2570
rect 30209 2506 30210 2570
rect 30144 2490 30210 2506
rect 30144 2426 30145 2490
rect 30209 2426 30210 2490
rect 30144 2410 30210 2426
rect 30144 2346 30145 2410
rect 30209 2346 30210 2410
rect 30144 2330 30210 2346
rect 30144 2266 30145 2330
rect 30209 2266 30210 2330
rect 30144 2250 30210 2266
rect 30144 2186 30145 2250
rect 30209 2186 30210 2250
rect 30144 2170 30210 2186
rect 30144 2106 30145 2170
rect 30209 2106 30210 2170
rect 30144 2090 30210 2106
rect 30144 2026 30145 2090
rect 30209 2026 30210 2090
rect 30144 1936 30210 2026
rect 30270 1932 30330 2964
rect 30390 1872 30450 2902
rect 30510 1932 30570 2964
rect 30630 1872 30690 2902
rect 30750 2810 30816 2964
rect 30750 2746 30751 2810
rect 30815 2746 30816 2810
rect 30750 2730 30816 2746
rect 30750 2666 30751 2730
rect 30815 2666 30816 2730
rect 30750 2650 30816 2666
rect 30750 2586 30751 2650
rect 30815 2586 30816 2650
rect 30750 2570 30816 2586
rect 30750 2506 30751 2570
rect 30815 2506 30816 2570
rect 30750 2490 30816 2506
rect 30750 2426 30751 2490
rect 30815 2426 30816 2490
rect 30750 2410 30816 2426
rect 30750 2346 30751 2410
rect 30815 2346 30816 2410
rect 30750 2330 30816 2346
rect 30750 2266 30751 2330
rect 30815 2266 30816 2330
rect 30750 2250 30816 2266
rect 30750 2186 30751 2250
rect 30815 2186 30816 2250
rect 30750 2170 30816 2186
rect 30750 2106 30751 2170
rect 30815 2106 30816 2170
rect 30750 2090 30816 2106
rect 30750 2026 30751 2090
rect 30815 2026 30816 2090
rect 30750 1936 30816 2026
rect 30876 1932 30936 2964
rect 30996 1872 31056 2902
rect 31116 1932 31176 2964
rect 31236 1872 31296 2902
rect 31356 2810 31422 2964
rect 31356 2746 31357 2810
rect 31421 2746 31422 2810
rect 31356 2730 31422 2746
rect 31356 2666 31357 2730
rect 31421 2666 31422 2730
rect 31356 2650 31422 2666
rect 31356 2586 31357 2650
rect 31421 2586 31422 2650
rect 31356 2570 31422 2586
rect 31356 2506 31357 2570
rect 31421 2506 31422 2570
rect 31356 2490 31422 2506
rect 31356 2426 31357 2490
rect 31421 2426 31422 2490
rect 31356 2410 31422 2426
rect 31356 2346 31357 2410
rect 31421 2346 31422 2410
rect 31356 2330 31422 2346
rect 31356 2266 31357 2330
rect 31421 2266 31422 2330
rect 31356 2250 31422 2266
rect 31356 2186 31357 2250
rect 31421 2186 31422 2250
rect 31356 2170 31422 2186
rect 31356 2106 31357 2170
rect 31421 2106 31422 2170
rect 31356 2090 31422 2106
rect 31356 2026 31357 2090
rect 31421 2026 31422 2090
rect 31356 1936 31422 2026
rect 31482 1932 31542 2964
rect 31602 1872 31662 2902
rect 31722 1932 31782 2964
rect 31842 1872 31902 2902
rect 31962 2810 32028 2964
rect 31962 2746 31963 2810
rect 32027 2746 32028 2810
rect 31962 2730 32028 2746
rect 31962 2666 31963 2730
rect 32027 2666 32028 2730
rect 31962 2650 32028 2666
rect 31962 2586 31963 2650
rect 32027 2586 32028 2650
rect 31962 2570 32028 2586
rect 31962 2506 31963 2570
rect 32027 2506 32028 2570
rect 31962 2490 32028 2506
rect 31962 2426 31963 2490
rect 32027 2426 32028 2490
rect 31962 2410 32028 2426
rect 31962 2346 31963 2410
rect 32027 2346 32028 2410
rect 31962 2330 32028 2346
rect 31962 2266 31963 2330
rect 32027 2266 32028 2330
rect 31962 2250 32028 2266
rect 31962 2186 31963 2250
rect 32027 2186 32028 2250
rect 31962 2170 32028 2186
rect 31962 2106 31963 2170
rect 32027 2106 32028 2170
rect 31962 2090 32028 2106
rect 31962 2026 31963 2090
rect 32027 2026 32028 2090
rect 31962 1936 32028 2026
rect 32088 1932 32148 2964
rect 32208 1872 32268 2902
rect 32328 1932 32388 2964
rect 32448 1872 32508 2902
rect 32568 2810 32634 2964
rect 32568 2746 32569 2810
rect 32633 2746 32634 2810
rect 32568 2730 32634 2746
rect 32568 2666 32569 2730
rect 32633 2666 32634 2730
rect 32568 2650 32634 2666
rect 32568 2586 32569 2650
rect 32633 2586 32634 2650
rect 32568 2570 32634 2586
rect 32568 2506 32569 2570
rect 32633 2506 32634 2570
rect 32568 2490 32634 2506
rect 32568 2426 32569 2490
rect 32633 2426 32634 2490
rect 32568 2410 32634 2426
rect 32568 2346 32569 2410
rect 32633 2346 32634 2410
rect 32568 2330 32634 2346
rect 32568 2266 32569 2330
rect 32633 2266 32634 2330
rect 32568 2250 32634 2266
rect 32568 2186 32569 2250
rect 32633 2186 32634 2250
rect 32568 2170 32634 2186
rect 32568 2106 32569 2170
rect 32633 2106 32634 2170
rect 32568 2090 32634 2106
rect 32568 2026 32569 2090
rect 32633 2026 32634 2090
rect 32568 1936 32634 2026
rect 32694 1932 32754 2964
rect 32814 1872 32874 2902
rect 32934 1932 32994 2964
rect 33054 1872 33114 2902
rect 33174 2810 33240 2964
rect 33174 2746 33175 2810
rect 33239 2746 33240 2810
rect 33174 2730 33240 2746
rect 33174 2666 33175 2730
rect 33239 2666 33240 2730
rect 33174 2650 33240 2666
rect 33174 2586 33175 2650
rect 33239 2586 33240 2650
rect 33174 2570 33240 2586
rect 33174 2506 33175 2570
rect 33239 2506 33240 2570
rect 33174 2490 33240 2506
rect 33174 2426 33175 2490
rect 33239 2426 33240 2490
rect 33174 2410 33240 2426
rect 33174 2346 33175 2410
rect 33239 2346 33240 2410
rect 33174 2330 33240 2346
rect 33174 2266 33175 2330
rect 33239 2266 33240 2330
rect 33174 2250 33240 2266
rect 33174 2186 33175 2250
rect 33239 2186 33240 2250
rect 33174 2170 33240 2186
rect 33174 2106 33175 2170
rect 33239 2106 33240 2170
rect 33174 2090 33240 2106
rect 33174 2026 33175 2090
rect 33239 2026 33240 2090
rect 33174 1936 33240 2026
rect 13782 1870 33240 1872
rect 13782 1806 13886 1870
rect 13950 1806 13966 1870
rect 14030 1806 14046 1870
rect 14110 1806 14126 1870
rect 14190 1806 14206 1870
rect 14270 1806 14286 1870
rect 14350 1806 14492 1870
rect 14556 1806 14572 1870
rect 14636 1806 14652 1870
rect 14716 1806 14732 1870
rect 14796 1806 14812 1870
rect 14876 1806 14892 1870
rect 14956 1806 15098 1870
rect 15162 1806 15178 1870
rect 15242 1806 15258 1870
rect 15322 1806 15338 1870
rect 15402 1806 15418 1870
rect 15482 1806 15498 1870
rect 15562 1806 15704 1870
rect 15768 1806 15784 1870
rect 15848 1806 15864 1870
rect 15928 1806 15944 1870
rect 16008 1806 16024 1870
rect 16088 1806 16104 1870
rect 16168 1806 16310 1870
rect 16374 1806 16390 1870
rect 16454 1806 16470 1870
rect 16534 1806 16550 1870
rect 16614 1806 16630 1870
rect 16694 1806 16710 1870
rect 16774 1806 16916 1870
rect 16980 1806 16996 1870
rect 17060 1806 17076 1870
rect 17140 1806 17156 1870
rect 17220 1806 17236 1870
rect 17300 1806 17316 1870
rect 17380 1806 17522 1870
rect 17586 1806 17602 1870
rect 17666 1806 17682 1870
rect 17746 1806 17762 1870
rect 17826 1806 17842 1870
rect 17906 1806 17922 1870
rect 17986 1806 18128 1870
rect 18192 1806 18208 1870
rect 18272 1806 18288 1870
rect 18352 1806 18368 1870
rect 18432 1806 18448 1870
rect 18512 1806 18528 1870
rect 18592 1806 18734 1870
rect 18798 1806 18814 1870
rect 18878 1806 18894 1870
rect 18958 1806 18974 1870
rect 19038 1806 19054 1870
rect 19118 1806 19134 1870
rect 19198 1806 19340 1870
rect 19404 1806 19420 1870
rect 19484 1806 19500 1870
rect 19564 1806 19580 1870
rect 19644 1806 19660 1870
rect 19724 1806 19740 1870
rect 19804 1806 19946 1870
rect 20010 1806 20026 1870
rect 20090 1806 20106 1870
rect 20170 1806 20186 1870
rect 20250 1806 20266 1870
rect 20330 1806 20346 1870
rect 20410 1806 20552 1870
rect 20616 1806 20632 1870
rect 20696 1806 20712 1870
rect 20776 1806 20792 1870
rect 20856 1806 20872 1870
rect 20936 1806 20952 1870
rect 21016 1806 21158 1870
rect 21222 1806 21238 1870
rect 21302 1806 21318 1870
rect 21382 1806 21398 1870
rect 21462 1806 21478 1870
rect 21542 1806 21558 1870
rect 21622 1806 21764 1870
rect 21828 1806 21844 1870
rect 21908 1806 21924 1870
rect 21988 1806 22004 1870
rect 22068 1806 22084 1870
rect 22148 1806 22164 1870
rect 22228 1806 22370 1870
rect 22434 1806 22450 1870
rect 22514 1806 22530 1870
rect 22594 1806 22610 1870
rect 22674 1806 22690 1870
rect 22754 1806 22770 1870
rect 22834 1806 22976 1870
rect 23040 1806 23056 1870
rect 23120 1806 23136 1870
rect 23200 1806 23216 1870
rect 23280 1806 23296 1870
rect 23360 1806 23376 1870
rect 23440 1806 23582 1870
rect 23646 1806 23662 1870
rect 23726 1806 23742 1870
rect 23806 1806 23822 1870
rect 23886 1806 23902 1870
rect 23966 1806 23982 1870
rect 24046 1806 24188 1870
rect 24252 1806 24268 1870
rect 24332 1806 24348 1870
rect 24412 1806 24428 1870
rect 24492 1806 24508 1870
rect 24572 1806 24588 1870
rect 24652 1806 24794 1870
rect 24858 1806 24874 1870
rect 24938 1806 24954 1870
rect 25018 1806 25034 1870
rect 25098 1806 25114 1870
rect 25178 1806 25194 1870
rect 25258 1806 25400 1870
rect 25464 1806 25480 1870
rect 25544 1806 25560 1870
rect 25624 1806 25640 1870
rect 25704 1806 25720 1870
rect 25784 1806 25800 1870
rect 25864 1806 26006 1870
rect 26070 1806 26086 1870
rect 26150 1806 26166 1870
rect 26230 1806 26246 1870
rect 26310 1806 26326 1870
rect 26390 1806 26406 1870
rect 26470 1806 26612 1870
rect 26676 1806 26692 1870
rect 26756 1806 26772 1870
rect 26836 1806 26852 1870
rect 26916 1806 26932 1870
rect 26996 1806 27012 1870
rect 27076 1806 27218 1870
rect 27282 1806 27298 1870
rect 27362 1806 27378 1870
rect 27442 1806 27458 1870
rect 27522 1806 27538 1870
rect 27602 1806 27618 1870
rect 27682 1806 27824 1870
rect 27888 1806 27904 1870
rect 27968 1806 27984 1870
rect 28048 1806 28064 1870
rect 28128 1806 28144 1870
rect 28208 1806 28224 1870
rect 28288 1806 28430 1870
rect 28494 1806 28510 1870
rect 28574 1806 28590 1870
rect 28654 1806 28670 1870
rect 28734 1806 28750 1870
rect 28814 1806 28830 1870
rect 28894 1806 29036 1870
rect 29100 1806 29116 1870
rect 29180 1806 29196 1870
rect 29260 1806 29276 1870
rect 29340 1806 29356 1870
rect 29420 1806 29436 1870
rect 29500 1806 29642 1870
rect 29706 1806 29722 1870
rect 29786 1806 29802 1870
rect 29866 1806 29882 1870
rect 29946 1806 29962 1870
rect 30026 1806 30042 1870
rect 30106 1806 30248 1870
rect 30312 1806 30328 1870
rect 30392 1806 30408 1870
rect 30472 1806 30488 1870
rect 30552 1806 30568 1870
rect 30632 1806 30648 1870
rect 30712 1806 30854 1870
rect 30918 1806 30934 1870
rect 30998 1806 31014 1870
rect 31078 1806 31094 1870
rect 31158 1806 31174 1870
rect 31238 1806 31254 1870
rect 31318 1806 31460 1870
rect 31524 1806 31540 1870
rect 31604 1806 31620 1870
rect 31684 1806 31700 1870
rect 31764 1806 31780 1870
rect 31844 1806 31860 1870
rect 31924 1806 32066 1870
rect 32130 1806 32146 1870
rect 32210 1806 32226 1870
rect 32290 1806 32306 1870
rect 32370 1806 32386 1870
rect 32450 1806 32466 1870
rect 32530 1806 32672 1870
rect 32736 1806 32752 1870
rect 32816 1806 32832 1870
rect 32896 1806 32912 1870
rect 32976 1806 32992 1870
rect 33056 1806 33072 1870
rect 33136 1806 33240 1870
rect 13782 1804 33240 1806
<< via3 >>
rect 13886 4126 13950 4190
rect 13966 4126 14030 4190
rect 14046 4126 14110 4190
rect 14126 4126 14190 4190
rect 14206 4126 14270 4190
rect 14286 4126 14350 4190
rect 14492 4126 14556 4190
rect 14572 4126 14636 4190
rect 14652 4126 14716 4190
rect 14732 4126 14796 4190
rect 14812 4126 14876 4190
rect 14892 4126 14956 4190
rect 15098 4126 15162 4190
rect 15178 4126 15242 4190
rect 15258 4126 15322 4190
rect 15338 4126 15402 4190
rect 15418 4126 15482 4190
rect 15498 4126 15562 4190
rect 15704 4126 15768 4190
rect 15784 4126 15848 4190
rect 15864 4126 15928 4190
rect 15944 4126 16008 4190
rect 16024 4126 16088 4190
rect 16104 4126 16168 4190
rect 16310 4126 16374 4190
rect 16390 4126 16454 4190
rect 16470 4126 16534 4190
rect 16550 4126 16614 4190
rect 16630 4126 16694 4190
rect 16710 4126 16774 4190
rect 16916 4126 16980 4190
rect 16996 4126 17060 4190
rect 17076 4126 17140 4190
rect 17156 4126 17220 4190
rect 17236 4126 17300 4190
rect 17316 4126 17380 4190
rect 17522 4126 17586 4190
rect 17602 4126 17666 4190
rect 17682 4126 17746 4190
rect 17762 4126 17826 4190
rect 17842 4126 17906 4190
rect 17922 4126 17986 4190
rect 18128 4126 18192 4190
rect 18208 4126 18272 4190
rect 18288 4126 18352 4190
rect 18368 4126 18432 4190
rect 18448 4126 18512 4190
rect 18528 4126 18592 4190
rect 18734 4126 18798 4190
rect 18814 4126 18878 4190
rect 18894 4126 18958 4190
rect 18974 4126 19038 4190
rect 19054 4126 19118 4190
rect 19134 4126 19198 4190
rect 19340 4126 19404 4190
rect 19420 4126 19484 4190
rect 19500 4126 19564 4190
rect 19580 4126 19644 4190
rect 19660 4126 19724 4190
rect 19740 4126 19804 4190
rect 19946 4126 20010 4190
rect 20026 4126 20090 4190
rect 20106 4126 20170 4190
rect 20186 4126 20250 4190
rect 20266 4126 20330 4190
rect 20346 4126 20410 4190
rect 20552 4126 20616 4190
rect 20632 4126 20696 4190
rect 20712 4126 20776 4190
rect 20792 4126 20856 4190
rect 20872 4126 20936 4190
rect 20952 4126 21016 4190
rect 21158 4126 21222 4190
rect 21238 4126 21302 4190
rect 21318 4126 21382 4190
rect 21398 4126 21462 4190
rect 21478 4126 21542 4190
rect 21558 4126 21622 4190
rect 21764 4126 21828 4190
rect 21844 4126 21908 4190
rect 21924 4126 21988 4190
rect 22004 4126 22068 4190
rect 22084 4126 22148 4190
rect 22164 4126 22228 4190
rect 22370 4126 22434 4190
rect 22450 4126 22514 4190
rect 22530 4126 22594 4190
rect 22610 4126 22674 4190
rect 22690 4126 22754 4190
rect 22770 4126 22834 4190
rect 22976 4126 23040 4190
rect 23056 4126 23120 4190
rect 23136 4126 23200 4190
rect 23216 4126 23280 4190
rect 23296 4126 23360 4190
rect 23376 4126 23440 4190
rect 23582 4126 23646 4190
rect 23662 4126 23726 4190
rect 23742 4126 23806 4190
rect 23822 4126 23886 4190
rect 23902 4126 23966 4190
rect 23982 4126 24046 4190
rect 24188 4126 24252 4190
rect 24268 4126 24332 4190
rect 24348 4126 24412 4190
rect 24428 4126 24492 4190
rect 24508 4126 24572 4190
rect 24588 4126 24652 4190
rect 24794 4126 24858 4190
rect 24874 4126 24938 4190
rect 24954 4126 25018 4190
rect 25034 4126 25098 4190
rect 25114 4126 25178 4190
rect 25194 4126 25258 4190
rect 25400 4126 25464 4190
rect 25480 4126 25544 4190
rect 25560 4126 25624 4190
rect 25640 4126 25704 4190
rect 25720 4126 25784 4190
rect 25800 4126 25864 4190
rect 26006 4126 26070 4190
rect 26086 4126 26150 4190
rect 26166 4126 26230 4190
rect 26246 4126 26310 4190
rect 26326 4126 26390 4190
rect 26406 4126 26470 4190
rect 26612 4126 26676 4190
rect 26692 4126 26756 4190
rect 26772 4126 26836 4190
rect 26852 4126 26916 4190
rect 26932 4126 26996 4190
rect 27012 4126 27076 4190
rect 27218 4126 27282 4190
rect 27298 4126 27362 4190
rect 27378 4126 27442 4190
rect 27458 4126 27522 4190
rect 27538 4126 27602 4190
rect 27618 4126 27682 4190
rect 27824 4126 27888 4190
rect 27904 4126 27968 4190
rect 27984 4126 28048 4190
rect 28064 4126 28128 4190
rect 28144 4126 28208 4190
rect 28224 4126 28288 4190
rect 28430 4126 28494 4190
rect 28510 4126 28574 4190
rect 28590 4126 28654 4190
rect 28670 4126 28734 4190
rect 28750 4126 28814 4190
rect 28830 4126 28894 4190
rect 29036 4126 29100 4190
rect 29116 4126 29180 4190
rect 29196 4126 29260 4190
rect 29276 4126 29340 4190
rect 29356 4126 29420 4190
rect 29436 4126 29500 4190
rect 29642 4126 29706 4190
rect 29722 4126 29786 4190
rect 29802 4126 29866 4190
rect 29882 4126 29946 4190
rect 29962 4126 30026 4190
rect 30042 4126 30106 4190
rect 30248 4126 30312 4190
rect 30328 4126 30392 4190
rect 30408 4126 30472 4190
rect 30488 4126 30552 4190
rect 30568 4126 30632 4190
rect 30648 4126 30712 4190
rect 30854 4126 30918 4190
rect 30934 4126 30998 4190
rect 31014 4126 31078 4190
rect 31094 4126 31158 4190
rect 31174 4126 31238 4190
rect 31254 4126 31318 4190
rect 31460 4126 31524 4190
rect 31540 4126 31604 4190
rect 31620 4126 31684 4190
rect 31700 4126 31764 4190
rect 31780 4126 31844 4190
rect 31860 4126 31924 4190
rect 32066 4126 32130 4190
rect 32146 4126 32210 4190
rect 32226 4126 32290 4190
rect 32306 4126 32370 4190
rect 32386 4126 32450 4190
rect 32466 4126 32530 4190
rect 32672 4126 32736 4190
rect 32752 4126 32816 4190
rect 32832 4126 32896 4190
rect 32912 4126 32976 4190
rect 32992 4126 33056 4190
rect 33072 4126 33136 4190
rect 13783 3906 13847 3970
rect 13783 3826 13847 3890
rect 13783 3746 13847 3810
rect 13783 3666 13847 3730
rect 13783 3586 13847 3650
rect 13783 3506 13847 3570
rect 13783 3426 13847 3490
rect 13783 3346 13847 3410
rect 13783 3266 13847 3330
rect 13783 3186 13847 3250
rect 14389 3906 14453 3970
rect 14389 3826 14453 3890
rect 14389 3746 14453 3810
rect 14389 3666 14453 3730
rect 14389 3586 14453 3650
rect 14389 3506 14453 3570
rect 14389 3426 14453 3490
rect 14389 3346 14453 3410
rect 14389 3266 14453 3330
rect 14389 3186 14453 3250
rect 14995 3906 15059 3970
rect 14995 3826 15059 3890
rect 14995 3746 15059 3810
rect 14995 3666 15059 3730
rect 14995 3586 15059 3650
rect 14995 3506 15059 3570
rect 14995 3426 15059 3490
rect 14995 3346 15059 3410
rect 14995 3266 15059 3330
rect 14995 3186 15059 3250
rect 15601 3906 15665 3970
rect 15601 3826 15665 3890
rect 15601 3746 15665 3810
rect 15601 3666 15665 3730
rect 15601 3586 15665 3650
rect 15601 3506 15665 3570
rect 15601 3426 15665 3490
rect 15601 3346 15665 3410
rect 15601 3266 15665 3330
rect 15601 3186 15665 3250
rect 16207 3906 16271 3970
rect 16207 3826 16271 3890
rect 16207 3746 16271 3810
rect 16207 3666 16271 3730
rect 16207 3586 16271 3650
rect 16207 3506 16271 3570
rect 16207 3426 16271 3490
rect 16207 3346 16271 3410
rect 16207 3266 16271 3330
rect 16207 3186 16271 3250
rect 16813 3906 16877 3970
rect 16813 3826 16877 3890
rect 16813 3746 16877 3810
rect 16813 3666 16877 3730
rect 16813 3586 16877 3650
rect 16813 3506 16877 3570
rect 16813 3426 16877 3490
rect 16813 3346 16877 3410
rect 16813 3266 16877 3330
rect 16813 3186 16877 3250
rect 17419 3906 17483 3970
rect 17419 3826 17483 3890
rect 17419 3746 17483 3810
rect 17419 3666 17483 3730
rect 17419 3586 17483 3650
rect 17419 3506 17483 3570
rect 17419 3426 17483 3490
rect 17419 3346 17483 3410
rect 17419 3266 17483 3330
rect 17419 3186 17483 3250
rect 18025 3906 18089 3970
rect 18025 3826 18089 3890
rect 18025 3746 18089 3810
rect 18025 3666 18089 3730
rect 18025 3586 18089 3650
rect 18025 3506 18089 3570
rect 18025 3426 18089 3490
rect 18025 3346 18089 3410
rect 18025 3266 18089 3330
rect 18025 3186 18089 3250
rect 18631 3906 18695 3970
rect 18631 3826 18695 3890
rect 18631 3746 18695 3810
rect 18631 3666 18695 3730
rect 18631 3586 18695 3650
rect 18631 3506 18695 3570
rect 18631 3426 18695 3490
rect 18631 3346 18695 3410
rect 18631 3266 18695 3330
rect 18631 3186 18695 3250
rect 19237 3906 19301 3970
rect 19237 3826 19301 3890
rect 19237 3746 19301 3810
rect 19237 3666 19301 3730
rect 19237 3586 19301 3650
rect 19237 3506 19301 3570
rect 19237 3426 19301 3490
rect 19237 3346 19301 3410
rect 19237 3266 19301 3330
rect 19237 3186 19301 3250
rect 19843 3906 19907 3970
rect 19843 3826 19907 3890
rect 19843 3746 19907 3810
rect 19843 3666 19907 3730
rect 19843 3586 19907 3650
rect 19843 3506 19907 3570
rect 19843 3426 19907 3490
rect 19843 3346 19907 3410
rect 19843 3266 19907 3330
rect 19843 3186 19907 3250
rect 20449 3906 20513 3970
rect 20449 3826 20513 3890
rect 20449 3746 20513 3810
rect 20449 3666 20513 3730
rect 20449 3586 20513 3650
rect 20449 3506 20513 3570
rect 20449 3426 20513 3490
rect 20449 3346 20513 3410
rect 20449 3266 20513 3330
rect 20449 3186 20513 3250
rect 21055 3906 21119 3970
rect 21055 3826 21119 3890
rect 21055 3746 21119 3810
rect 21055 3666 21119 3730
rect 21055 3586 21119 3650
rect 21055 3506 21119 3570
rect 21055 3426 21119 3490
rect 21055 3346 21119 3410
rect 21055 3266 21119 3330
rect 21055 3186 21119 3250
rect 21661 3906 21725 3970
rect 21661 3826 21725 3890
rect 21661 3746 21725 3810
rect 21661 3666 21725 3730
rect 21661 3586 21725 3650
rect 21661 3506 21725 3570
rect 21661 3426 21725 3490
rect 21661 3346 21725 3410
rect 21661 3266 21725 3330
rect 21661 3186 21725 3250
rect 22267 3906 22331 3970
rect 22267 3826 22331 3890
rect 22267 3746 22331 3810
rect 22267 3666 22331 3730
rect 22267 3586 22331 3650
rect 22267 3506 22331 3570
rect 22267 3426 22331 3490
rect 22267 3346 22331 3410
rect 22267 3266 22331 3330
rect 22267 3186 22331 3250
rect 22873 3906 22937 3970
rect 22873 3826 22937 3890
rect 22873 3746 22937 3810
rect 22873 3666 22937 3730
rect 22873 3586 22937 3650
rect 22873 3506 22937 3570
rect 22873 3426 22937 3490
rect 22873 3346 22937 3410
rect 22873 3266 22937 3330
rect 22873 3186 22937 3250
rect 23479 3906 23543 3970
rect 23479 3826 23543 3890
rect 23479 3746 23543 3810
rect 23479 3666 23543 3730
rect 23479 3586 23543 3650
rect 23479 3506 23543 3570
rect 23479 3426 23543 3490
rect 23479 3346 23543 3410
rect 23479 3266 23543 3330
rect 23479 3186 23543 3250
rect 24085 3906 24149 3970
rect 24085 3826 24149 3890
rect 24085 3746 24149 3810
rect 24085 3666 24149 3730
rect 24085 3586 24149 3650
rect 24085 3506 24149 3570
rect 24085 3426 24149 3490
rect 24085 3346 24149 3410
rect 24085 3266 24149 3330
rect 24085 3186 24149 3250
rect 24691 3906 24755 3970
rect 24691 3826 24755 3890
rect 24691 3746 24755 3810
rect 24691 3666 24755 3730
rect 24691 3586 24755 3650
rect 24691 3506 24755 3570
rect 24691 3426 24755 3490
rect 24691 3346 24755 3410
rect 24691 3266 24755 3330
rect 24691 3186 24755 3250
rect 25297 3906 25361 3970
rect 25297 3826 25361 3890
rect 25297 3746 25361 3810
rect 25297 3666 25361 3730
rect 25297 3586 25361 3650
rect 25297 3506 25361 3570
rect 25297 3426 25361 3490
rect 25297 3346 25361 3410
rect 25297 3266 25361 3330
rect 25297 3186 25361 3250
rect 25903 3906 25967 3970
rect 25903 3826 25967 3890
rect 25903 3746 25967 3810
rect 25903 3666 25967 3730
rect 25903 3586 25967 3650
rect 25903 3506 25967 3570
rect 25903 3426 25967 3490
rect 25903 3346 25967 3410
rect 25903 3266 25967 3330
rect 25903 3186 25967 3250
rect 26509 3906 26573 3970
rect 26509 3826 26573 3890
rect 26509 3746 26573 3810
rect 26509 3666 26573 3730
rect 26509 3586 26573 3650
rect 26509 3506 26573 3570
rect 26509 3426 26573 3490
rect 26509 3346 26573 3410
rect 26509 3266 26573 3330
rect 26509 3186 26573 3250
rect 27115 3906 27179 3970
rect 27115 3826 27179 3890
rect 27115 3746 27179 3810
rect 27115 3666 27179 3730
rect 27115 3586 27179 3650
rect 27115 3506 27179 3570
rect 27115 3426 27179 3490
rect 27115 3346 27179 3410
rect 27115 3266 27179 3330
rect 27115 3186 27179 3250
rect 27721 3906 27785 3970
rect 27721 3826 27785 3890
rect 27721 3746 27785 3810
rect 27721 3666 27785 3730
rect 27721 3586 27785 3650
rect 27721 3506 27785 3570
rect 27721 3426 27785 3490
rect 27721 3346 27785 3410
rect 27721 3266 27785 3330
rect 27721 3186 27785 3250
rect 28327 3906 28391 3970
rect 28327 3826 28391 3890
rect 28327 3746 28391 3810
rect 28327 3666 28391 3730
rect 28327 3586 28391 3650
rect 28327 3506 28391 3570
rect 28327 3426 28391 3490
rect 28327 3346 28391 3410
rect 28327 3266 28391 3330
rect 28327 3186 28391 3250
rect 28933 3906 28997 3970
rect 28933 3826 28997 3890
rect 28933 3746 28997 3810
rect 28933 3666 28997 3730
rect 28933 3586 28997 3650
rect 28933 3506 28997 3570
rect 28933 3426 28997 3490
rect 28933 3346 28997 3410
rect 28933 3266 28997 3330
rect 28933 3186 28997 3250
rect 29539 3906 29603 3970
rect 29539 3826 29603 3890
rect 29539 3746 29603 3810
rect 29539 3666 29603 3730
rect 29539 3586 29603 3650
rect 29539 3506 29603 3570
rect 29539 3426 29603 3490
rect 29539 3346 29603 3410
rect 29539 3266 29603 3330
rect 29539 3186 29603 3250
rect 30145 3906 30209 3970
rect 30145 3826 30209 3890
rect 30145 3746 30209 3810
rect 30145 3666 30209 3730
rect 30145 3586 30209 3650
rect 30145 3506 30209 3570
rect 30145 3426 30209 3490
rect 30145 3346 30209 3410
rect 30145 3266 30209 3330
rect 30145 3186 30209 3250
rect 30751 3906 30815 3970
rect 30751 3826 30815 3890
rect 30751 3746 30815 3810
rect 30751 3666 30815 3730
rect 30751 3586 30815 3650
rect 30751 3506 30815 3570
rect 30751 3426 30815 3490
rect 30751 3346 30815 3410
rect 30751 3266 30815 3330
rect 30751 3186 30815 3250
rect 31357 3906 31421 3970
rect 31357 3826 31421 3890
rect 31357 3746 31421 3810
rect 31357 3666 31421 3730
rect 31357 3586 31421 3650
rect 31357 3506 31421 3570
rect 31357 3426 31421 3490
rect 31357 3346 31421 3410
rect 31357 3266 31421 3330
rect 31357 3186 31421 3250
rect 31963 3906 32027 3970
rect 31963 3826 32027 3890
rect 31963 3746 32027 3810
rect 31963 3666 32027 3730
rect 31963 3586 32027 3650
rect 31963 3506 32027 3570
rect 31963 3426 32027 3490
rect 31963 3346 32027 3410
rect 31963 3266 32027 3330
rect 31963 3186 32027 3250
rect 32569 3906 32633 3970
rect 32569 3826 32633 3890
rect 32569 3746 32633 3810
rect 32569 3666 32633 3730
rect 32569 3586 32633 3650
rect 32569 3506 32633 3570
rect 32569 3426 32633 3490
rect 32569 3346 32633 3410
rect 32569 3266 32633 3330
rect 32569 3186 32633 3250
rect 33175 3906 33239 3970
rect 33175 3826 33239 3890
rect 33175 3746 33239 3810
rect 33175 3666 33239 3730
rect 33175 3586 33239 3650
rect 33175 3506 33239 3570
rect 33175 3426 33239 3490
rect 33175 3346 33239 3410
rect 33175 3266 33239 3330
rect 33175 3186 33239 3250
rect 13886 2966 13950 3030
rect 13966 2966 14030 3030
rect 14046 2966 14110 3030
rect 14126 2966 14190 3030
rect 14206 2966 14270 3030
rect 14286 2966 14350 3030
rect 14492 2966 14556 3030
rect 14572 2966 14636 3030
rect 14652 2966 14716 3030
rect 14732 2966 14796 3030
rect 14812 2966 14876 3030
rect 14892 2966 14956 3030
rect 15098 2966 15162 3030
rect 15178 2966 15242 3030
rect 15258 2966 15322 3030
rect 15338 2966 15402 3030
rect 15418 2966 15482 3030
rect 15498 2966 15562 3030
rect 15704 2966 15768 3030
rect 15784 2966 15848 3030
rect 15864 2966 15928 3030
rect 15944 2966 16008 3030
rect 16024 2966 16088 3030
rect 16104 2966 16168 3030
rect 16310 2966 16374 3030
rect 16390 2966 16454 3030
rect 16470 2966 16534 3030
rect 16550 2966 16614 3030
rect 16630 2966 16694 3030
rect 16710 2966 16774 3030
rect 16916 2966 16980 3030
rect 16996 2966 17060 3030
rect 17076 2966 17140 3030
rect 17156 2966 17220 3030
rect 17236 2966 17300 3030
rect 17316 2966 17380 3030
rect 17522 2966 17586 3030
rect 17602 2966 17666 3030
rect 17682 2966 17746 3030
rect 17762 2966 17826 3030
rect 17842 2966 17906 3030
rect 17922 2966 17986 3030
rect 18128 2966 18192 3030
rect 18208 2966 18272 3030
rect 18288 2966 18352 3030
rect 18368 2966 18432 3030
rect 18448 2966 18512 3030
rect 18528 2966 18592 3030
rect 18734 2966 18798 3030
rect 18814 2966 18878 3030
rect 18894 2966 18958 3030
rect 18974 2966 19038 3030
rect 19054 2966 19118 3030
rect 19134 2966 19198 3030
rect 19340 2966 19404 3030
rect 19420 2966 19484 3030
rect 19500 2966 19564 3030
rect 19580 2966 19644 3030
rect 19660 2966 19724 3030
rect 19740 2966 19804 3030
rect 19946 2966 20010 3030
rect 20026 2966 20090 3030
rect 20106 2966 20170 3030
rect 20186 2966 20250 3030
rect 20266 2966 20330 3030
rect 20346 2966 20410 3030
rect 20552 2966 20616 3030
rect 20632 2966 20696 3030
rect 20712 2966 20776 3030
rect 20792 2966 20856 3030
rect 20872 2966 20936 3030
rect 20952 2966 21016 3030
rect 21158 2966 21222 3030
rect 21238 2966 21302 3030
rect 21318 2966 21382 3030
rect 21398 2966 21462 3030
rect 21478 2966 21542 3030
rect 21558 2966 21622 3030
rect 21764 2966 21828 3030
rect 21844 2966 21908 3030
rect 21924 2966 21988 3030
rect 22004 2966 22068 3030
rect 22084 2966 22148 3030
rect 22164 2966 22228 3030
rect 22370 2966 22434 3030
rect 22450 2966 22514 3030
rect 22530 2966 22594 3030
rect 22610 2966 22674 3030
rect 22690 2966 22754 3030
rect 22770 2966 22834 3030
rect 22976 2966 23040 3030
rect 23056 2966 23120 3030
rect 23136 2966 23200 3030
rect 23216 2966 23280 3030
rect 23296 2966 23360 3030
rect 23376 2966 23440 3030
rect 23582 2966 23646 3030
rect 23662 2966 23726 3030
rect 23742 2966 23806 3030
rect 23822 2966 23886 3030
rect 23902 2966 23966 3030
rect 23982 2966 24046 3030
rect 24188 2966 24252 3030
rect 24268 2966 24332 3030
rect 24348 2966 24412 3030
rect 24428 2966 24492 3030
rect 24508 2966 24572 3030
rect 24588 2966 24652 3030
rect 24794 2966 24858 3030
rect 24874 2966 24938 3030
rect 24954 2966 25018 3030
rect 25034 2966 25098 3030
rect 25114 2966 25178 3030
rect 25194 2966 25258 3030
rect 25400 2966 25464 3030
rect 25480 2966 25544 3030
rect 25560 2966 25624 3030
rect 25640 2966 25704 3030
rect 25720 2966 25784 3030
rect 25800 2966 25864 3030
rect 26006 2966 26070 3030
rect 26086 2966 26150 3030
rect 26166 2966 26230 3030
rect 26246 2966 26310 3030
rect 26326 2966 26390 3030
rect 26406 2966 26470 3030
rect 26612 2966 26676 3030
rect 26692 2966 26756 3030
rect 26772 2966 26836 3030
rect 26852 2966 26916 3030
rect 26932 2966 26996 3030
rect 27012 2966 27076 3030
rect 27218 2966 27282 3030
rect 27298 2966 27362 3030
rect 27378 2966 27442 3030
rect 27458 2966 27522 3030
rect 27538 2966 27602 3030
rect 27618 2966 27682 3030
rect 27824 2966 27888 3030
rect 27904 2966 27968 3030
rect 27984 2966 28048 3030
rect 28064 2966 28128 3030
rect 28144 2966 28208 3030
rect 28224 2966 28288 3030
rect 28430 2966 28494 3030
rect 28510 2966 28574 3030
rect 28590 2966 28654 3030
rect 28670 2966 28734 3030
rect 28750 2966 28814 3030
rect 28830 2966 28894 3030
rect 29036 2966 29100 3030
rect 29116 2966 29180 3030
rect 29196 2966 29260 3030
rect 29276 2966 29340 3030
rect 29356 2966 29420 3030
rect 29436 2966 29500 3030
rect 29642 2966 29706 3030
rect 29722 2966 29786 3030
rect 29802 2966 29866 3030
rect 29882 2966 29946 3030
rect 29962 2966 30026 3030
rect 30042 2966 30106 3030
rect 30248 2966 30312 3030
rect 30328 2966 30392 3030
rect 30408 2966 30472 3030
rect 30488 2966 30552 3030
rect 30568 2966 30632 3030
rect 30648 2966 30712 3030
rect 30854 2966 30918 3030
rect 30934 2966 30998 3030
rect 31014 2966 31078 3030
rect 31094 2966 31158 3030
rect 31174 2966 31238 3030
rect 31254 2966 31318 3030
rect 31460 2966 31524 3030
rect 31540 2966 31604 3030
rect 31620 2966 31684 3030
rect 31700 2966 31764 3030
rect 31780 2966 31844 3030
rect 31860 2966 31924 3030
rect 32066 2966 32130 3030
rect 32146 2966 32210 3030
rect 32226 2966 32290 3030
rect 32306 2966 32370 3030
rect 32386 2966 32450 3030
rect 32466 2966 32530 3030
rect 32672 2966 32736 3030
rect 32752 2966 32816 3030
rect 32832 2966 32896 3030
rect 32912 2966 32976 3030
rect 32992 2966 33056 3030
rect 33072 2966 33136 3030
rect 13783 2746 13847 2810
rect 13783 2666 13847 2730
rect 13783 2586 13847 2650
rect 13783 2506 13847 2570
rect 13783 2426 13847 2490
rect 13783 2346 13847 2410
rect 13783 2266 13847 2330
rect 13783 2186 13847 2250
rect 13783 2106 13847 2170
rect 13783 2026 13847 2090
rect 14389 2746 14453 2810
rect 14389 2666 14453 2730
rect 14389 2586 14453 2650
rect 14389 2506 14453 2570
rect 14389 2426 14453 2490
rect 14389 2346 14453 2410
rect 14389 2266 14453 2330
rect 14389 2186 14453 2250
rect 14389 2106 14453 2170
rect 14389 2026 14453 2090
rect 14995 2746 15059 2810
rect 14995 2666 15059 2730
rect 14995 2586 15059 2650
rect 14995 2506 15059 2570
rect 14995 2426 15059 2490
rect 14995 2346 15059 2410
rect 14995 2266 15059 2330
rect 14995 2186 15059 2250
rect 14995 2106 15059 2170
rect 14995 2026 15059 2090
rect 15601 2746 15665 2810
rect 15601 2666 15665 2730
rect 15601 2586 15665 2650
rect 15601 2506 15665 2570
rect 15601 2426 15665 2490
rect 15601 2346 15665 2410
rect 15601 2266 15665 2330
rect 15601 2186 15665 2250
rect 15601 2106 15665 2170
rect 15601 2026 15665 2090
rect 16207 2746 16271 2810
rect 16207 2666 16271 2730
rect 16207 2586 16271 2650
rect 16207 2506 16271 2570
rect 16207 2426 16271 2490
rect 16207 2346 16271 2410
rect 16207 2266 16271 2330
rect 16207 2186 16271 2250
rect 16207 2106 16271 2170
rect 16207 2026 16271 2090
rect 16813 2746 16877 2810
rect 16813 2666 16877 2730
rect 16813 2586 16877 2650
rect 16813 2506 16877 2570
rect 16813 2426 16877 2490
rect 16813 2346 16877 2410
rect 16813 2266 16877 2330
rect 16813 2186 16877 2250
rect 16813 2106 16877 2170
rect 16813 2026 16877 2090
rect 17419 2746 17483 2810
rect 17419 2666 17483 2730
rect 17419 2586 17483 2650
rect 17419 2506 17483 2570
rect 17419 2426 17483 2490
rect 17419 2346 17483 2410
rect 17419 2266 17483 2330
rect 17419 2186 17483 2250
rect 17419 2106 17483 2170
rect 17419 2026 17483 2090
rect 18025 2746 18089 2810
rect 18025 2666 18089 2730
rect 18025 2586 18089 2650
rect 18025 2506 18089 2570
rect 18025 2426 18089 2490
rect 18025 2346 18089 2410
rect 18025 2266 18089 2330
rect 18025 2186 18089 2250
rect 18025 2106 18089 2170
rect 18025 2026 18089 2090
rect 18631 2746 18695 2810
rect 18631 2666 18695 2730
rect 18631 2586 18695 2650
rect 18631 2506 18695 2570
rect 18631 2426 18695 2490
rect 18631 2346 18695 2410
rect 18631 2266 18695 2330
rect 18631 2186 18695 2250
rect 18631 2106 18695 2170
rect 18631 2026 18695 2090
rect 19237 2746 19301 2810
rect 19237 2666 19301 2730
rect 19237 2586 19301 2650
rect 19237 2506 19301 2570
rect 19237 2426 19301 2490
rect 19237 2346 19301 2410
rect 19237 2266 19301 2330
rect 19237 2186 19301 2250
rect 19237 2106 19301 2170
rect 19237 2026 19301 2090
rect 19843 2746 19907 2810
rect 19843 2666 19907 2730
rect 19843 2586 19907 2650
rect 19843 2506 19907 2570
rect 19843 2426 19907 2490
rect 19843 2346 19907 2410
rect 19843 2266 19907 2330
rect 19843 2186 19907 2250
rect 19843 2106 19907 2170
rect 19843 2026 19907 2090
rect 20449 2746 20513 2810
rect 20449 2666 20513 2730
rect 20449 2586 20513 2650
rect 20449 2506 20513 2570
rect 20449 2426 20513 2490
rect 20449 2346 20513 2410
rect 20449 2266 20513 2330
rect 20449 2186 20513 2250
rect 20449 2106 20513 2170
rect 20449 2026 20513 2090
rect 21055 2746 21119 2810
rect 21055 2666 21119 2730
rect 21055 2586 21119 2650
rect 21055 2506 21119 2570
rect 21055 2426 21119 2490
rect 21055 2346 21119 2410
rect 21055 2266 21119 2330
rect 21055 2186 21119 2250
rect 21055 2106 21119 2170
rect 21055 2026 21119 2090
rect 21661 2746 21725 2810
rect 21661 2666 21725 2730
rect 21661 2586 21725 2650
rect 21661 2506 21725 2570
rect 21661 2426 21725 2490
rect 21661 2346 21725 2410
rect 21661 2266 21725 2330
rect 21661 2186 21725 2250
rect 21661 2106 21725 2170
rect 21661 2026 21725 2090
rect 22267 2746 22331 2810
rect 22267 2666 22331 2730
rect 22267 2586 22331 2650
rect 22267 2506 22331 2570
rect 22267 2426 22331 2490
rect 22267 2346 22331 2410
rect 22267 2266 22331 2330
rect 22267 2186 22331 2250
rect 22267 2106 22331 2170
rect 22267 2026 22331 2090
rect 22873 2746 22937 2810
rect 22873 2666 22937 2730
rect 22873 2586 22937 2650
rect 22873 2506 22937 2570
rect 22873 2426 22937 2490
rect 22873 2346 22937 2410
rect 22873 2266 22937 2330
rect 22873 2186 22937 2250
rect 22873 2106 22937 2170
rect 22873 2026 22937 2090
rect 23479 2746 23543 2810
rect 23479 2666 23543 2730
rect 23479 2586 23543 2650
rect 23479 2506 23543 2570
rect 23479 2426 23543 2490
rect 23479 2346 23543 2410
rect 23479 2266 23543 2330
rect 23479 2186 23543 2250
rect 23479 2106 23543 2170
rect 23479 2026 23543 2090
rect 24085 2746 24149 2810
rect 24085 2666 24149 2730
rect 24085 2586 24149 2650
rect 24085 2506 24149 2570
rect 24085 2426 24149 2490
rect 24085 2346 24149 2410
rect 24085 2266 24149 2330
rect 24085 2186 24149 2250
rect 24085 2106 24149 2170
rect 24085 2026 24149 2090
rect 24691 2746 24755 2810
rect 24691 2666 24755 2730
rect 24691 2586 24755 2650
rect 24691 2506 24755 2570
rect 24691 2426 24755 2490
rect 24691 2346 24755 2410
rect 24691 2266 24755 2330
rect 24691 2186 24755 2250
rect 24691 2106 24755 2170
rect 24691 2026 24755 2090
rect 25297 2746 25361 2810
rect 25297 2666 25361 2730
rect 25297 2586 25361 2650
rect 25297 2506 25361 2570
rect 25297 2426 25361 2490
rect 25297 2346 25361 2410
rect 25297 2266 25361 2330
rect 25297 2186 25361 2250
rect 25297 2106 25361 2170
rect 25297 2026 25361 2090
rect 25903 2746 25967 2810
rect 25903 2666 25967 2730
rect 25903 2586 25967 2650
rect 25903 2506 25967 2570
rect 25903 2426 25967 2490
rect 25903 2346 25967 2410
rect 25903 2266 25967 2330
rect 25903 2186 25967 2250
rect 25903 2106 25967 2170
rect 25903 2026 25967 2090
rect 26509 2746 26573 2810
rect 26509 2666 26573 2730
rect 26509 2586 26573 2650
rect 26509 2506 26573 2570
rect 26509 2426 26573 2490
rect 26509 2346 26573 2410
rect 26509 2266 26573 2330
rect 26509 2186 26573 2250
rect 26509 2106 26573 2170
rect 26509 2026 26573 2090
rect 27115 2746 27179 2810
rect 27115 2666 27179 2730
rect 27115 2586 27179 2650
rect 27115 2506 27179 2570
rect 27115 2426 27179 2490
rect 27115 2346 27179 2410
rect 27115 2266 27179 2330
rect 27115 2186 27179 2250
rect 27115 2106 27179 2170
rect 27115 2026 27179 2090
rect 27721 2746 27785 2810
rect 27721 2666 27785 2730
rect 27721 2586 27785 2650
rect 27721 2506 27785 2570
rect 27721 2426 27785 2490
rect 27721 2346 27785 2410
rect 27721 2266 27785 2330
rect 27721 2186 27785 2250
rect 27721 2106 27785 2170
rect 27721 2026 27785 2090
rect 28327 2746 28391 2810
rect 28327 2666 28391 2730
rect 28327 2586 28391 2650
rect 28327 2506 28391 2570
rect 28327 2426 28391 2490
rect 28327 2346 28391 2410
rect 28327 2266 28391 2330
rect 28327 2186 28391 2250
rect 28327 2106 28391 2170
rect 28327 2026 28391 2090
rect 28933 2746 28997 2810
rect 28933 2666 28997 2730
rect 28933 2586 28997 2650
rect 28933 2506 28997 2570
rect 28933 2426 28997 2490
rect 28933 2346 28997 2410
rect 28933 2266 28997 2330
rect 28933 2186 28997 2250
rect 28933 2106 28997 2170
rect 28933 2026 28997 2090
rect 29539 2746 29603 2810
rect 29539 2666 29603 2730
rect 29539 2586 29603 2650
rect 29539 2506 29603 2570
rect 29539 2426 29603 2490
rect 29539 2346 29603 2410
rect 29539 2266 29603 2330
rect 29539 2186 29603 2250
rect 29539 2106 29603 2170
rect 29539 2026 29603 2090
rect 30145 2746 30209 2810
rect 30145 2666 30209 2730
rect 30145 2586 30209 2650
rect 30145 2506 30209 2570
rect 30145 2426 30209 2490
rect 30145 2346 30209 2410
rect 30145 2266 30209 2330
rect 30145 2186 30209 2250
rect 30145 2106 30209 2170
rect 30145 2026 30209 2090
rect 30751 2746 30815 2810
rect 30751 2666 30815 2730
rect 30751 2586 30815 2650
rect 30751 2506 30815 2570
rect 30751 2426 30815 2490
rect 30751 2346 30815 2410
rect 30751 2266 30815 2330
rect 30751 2186 30815 2250
rect 30751 2106 30815 2170
rect 30751 2026 30815 2090
rect 31357 2746 31421 2810
rect 31357 2666 31421 2730
rect 31357 2586 31421 2650
rect 31357 2506 31421 2570
rect 31357 2426 31421 2490
rect 31357 2346 31421 2410
rect 31357 2266 31421 2330
rect 31357 2186 31421 2250
rect 31357 2106 31421 2170
rect 31357 2026 31421 2090
rect 31963 2746 32027 2810
rect 31963 2666 32027 2730
rect 31963 2586 32027 2650
rect 31963 2506 32027 2570
rect 31963 2426 32027 2490
rect 31963 2346 32027 2410
rect 31963 2266 32027 2330
rect 31963 2186 32027 2250
rect 31963 2106 32027 2170
rect 31963 2026 32027 2090
rect 32569 2746 32633 2810
rect 32569 2666 32633 2730
rect 32569 2586 32633 2650
rect 32569 2506 32633 2570
rect 32569 2426 32633 2490
rect 32569 2346 32633 2410
rect 32569 2266 32633 2330
rect 32569 2186 32633 2250
rect 32569 2106 32633 2170
rect 32569 2026 32633 2090
rect 33175 2746 33239 2810
rect 33175 2666 33239 2730
rect 33175 2586 33239 2650
rect 33175 2506 33239 2570
rect 33175 2426 33239 2490
rect 33175 2346 33239 2410
rect 33175 2266 33239 2330
rect 33175 2186 33239 2250
rect 33175 2106 33239 2170
rect 33175 2026 33239 2090
rect 13886 1806 13950 1870
rect 13966 1806 14030 1870
rect 14046 1806 14110 1870
rect 14126 1806 14190 1870
rect 14206 1806 14270 1870
rect 14286 1806 14350 1870
rect 14492 1806 14556 1870
rect 14572 1806 14636 1870
rect 14652 1806 14716 1870
rect 14732 1806 14796 1870
rect 14812 1806 14876 1870
rect 14892 1806 14956 1870
rect 15098 1806 15162 1870
rect 15178 1806 15242 1870
rect 15258 1806 15322 1870
rect 15338 1806 15402 1870
rect 15418 1806 15482 1870
rect 15498 1806 15562 1870
rect 15704 1806 15768 1870
rect 15784 1806 15848 1870
rect 15864 1806 15928 1870
rect 15944 1806 16008 1870
rect 16024 1806 16088 1870
rect 16104 1806 16168 1870
rect 16310 1806 16374 1870
rect 16390 1806 16454 1870
rect 16470 1806 16534 1870
rect 16550 1806 16614 1870
rect 16630 1806 16694 1870
rect 16710 1806 16774 1870
rect 16916 1806 16980 1870
rect 16996 1806 17060 1870
rect 17076 1806 17140 1870
rect 17156 1806 17220 1870
rect 17236 1806 17300 1870
rect 17316 1806 17380 1870
rect 17522 1806 17586 1870
rect 17602 1806 17666 1870
rect 17682 1806 17746 1870
rect 17762 1806 17826 1870
rect 17842 1806 17906 1870
rect 17922 1806 17986 1870
rect 18128 1806 18192 1870
rect 18208 1806 18272 1870
rect 18288 1806 18352 1870
rect 18368 1806 18432 1870
rect 18448 1806 18512 1870
rect 18528 1806 18592 1870
rect 18734 1806 18798 1870
rect 18814 1806 18878 1870
rect 18894 1806 18958 1870
rect 18974 1806 19038 1870
rect 19054 1806 19118 1870
rect 19134 1806 19198 1870
rect 19340 1806 19404 1870
rect 19420 1806 19484 1870
rect 19500 1806 19564 1870
rect 19580 1806 19644 1870
rect 19660 1806 19724 1870
rect 19740 1806 19804 1870
rect 19946 1806 20010 1870
rect 20026 1806 20090 1870
rect 20106 1806 20170 1870
rect 20186 1806 20250 1870
rect 20266 1806 20330 1870
rect 20346 1806 20410 1870
rect 20552 1806 20616 1870
rect 20632 1806 20696 1870
rect 20712 1806 20776 1870
rect 20792 1806 20856 1870
rect 20872 1806 20936 1870
rect 20952 1806 21016 1870
rect 21158 1806 21222 1870
rect 21238 1806 21302 1870
rect 21318 1806 21382 1870
rect 21398 1806 21462 1870
rect 21478 1806 21542 1870
rect 21558 1806 21622 1870
rect 21764 1806 21828 1870
rect 21844 1806 21908 1870
rect 21924 1806 21988 1870
rect 22004 1806 22068 1870
rect 22084 1806 22148 1870
rect 22164 1806 22228 1870
rect 22370 1806 22434 1870
rect 22450 1806 22514 1870
rect 22530 1806 22594 1870
rect 22610 1806 22674 1870
rect 22690 1806 22754 1870
rect 22770 1806 22834 1870
rect 22976 1806 23040 1870
rect 23056 1806 23120 1870
rect 23136 1806 23200 1870
rect 23216 1806 23280 1870
rect 23296 1806 23360 1870
rect 23376 1806 23440 1870
rect 23582 1806 23646 1870
rect 23662 1806 23726 1870
rect 23742 1806 23806 1870
rect 23822 1806 23886 1870
rect 23902 1806 23966 1870
rect 23982 1806 24046 1870
rect 24188 1806 24252 1870
rect 24268 1806 24332 1870
rect 24348 1806 24412 1870
rect 24428 1806 24492 1870
rect 24508 1806 24572 1870
rect 24588 1806 24652 1870
rect 24794 1806 24858 1870
rect 24874 1806 24938 1870
rect 24954 1806 25018 1870
rect 25034 1806 25098 1870
rect 25114 1806 25178 1870
rect 25194 1806 25258 1870
rect 25400 1806 25464 1870
rect 25480 1806 25544 1870
rect 25560 1806 25624 1870
rect 25640 1806 25704 1870
rect 25720 1806 25784 1870
rect 25800 1806 25864 1870
rect 26006 1806 26070 1870
rect 26086 1806 26150 1870
rect 26166 1806 26230 1870
rect 26246 1806 26310 1870
rect 26326 1806 26390 1870
rect 26406 1806 26470 1870
rect 26612 1806 26676 1870
rect 26692 1806 26756 1870
rect 26772 1806 26836 1870
rect 26852 1806 26916 1870
rect 26932 1806 26996 1870
rect 27012 1806 27076 1870
rect 27218 1806 27282 1870
rect 27298 1806 27362 1870
rect 27378 1806 27442 1870
rect 27458 1806 27522 1870
rect 27538 1806 27602 1870
rect 27618 1806 27682 1870
rect 27824 1806 27888 1870
rect 27904 1806 27968 1870
rect 27984 1806 28048 1870
rect 28064 1806 28128 1870
rect 28144 1806 28208 1870
rect 28224 1806 28288 1870
rect 28430 1806 28494 1870
rect 28510 1806 28574 1870
rect 28590 1806 28654 1870
rect 28670 1806 28734 1870
rect 28750 1806 28814 1870
rect 28830 1806 28894 1870
rect 29036 1806 29100 1870
rect 29116 1806 29180 1870
rect 29196 1806 29260 1870
rect 29276 1806 29340 1870
rect 29356 1806 29420 1870
rect 29436 1806 29500 1870
rect 29642 1806 29706 1870
rect 29722 1806 29786 1870
rect 29802 1806 29866 1870
rect 29882 1806 29946 1870
rect 29962 1806 30026 1870
rect 30042 1806 30106 1870
rect 30248 1806 30312 1870
rect 30328 1806 30392 1870
rect 30408 1806 30472 1870
rect 30488 1806 30552 1870
rect 30568 1806 30632 1870
rect 30648 1806 30712 1870
rect 30854 1806 30918 1870
rect 30934 1806 30998 1870
rect 31014 1806 31078 1870
rect 31094 1806 31158 1870
rect 31174 1806 31238 1870
rect 31254 1806 31318 1870
rect 31460 1806 31524 1870
rect 31540 1806 31604 1870
rect 31620 1806 31684 1870
rect 31700 1806 31764 1870
rect 31780 1806 31844 1870
rect 31860 1806 31924 1870
rect 32066 1806 32130 1870
rect 32146 1806 32210 1870
rect 32226 1806 32290 1870
rect 32306 1806 32370 1870
rect 32386 1806 32450 1870
rect 32466 1806 32530 1870
rect 32672 1806 32736 1870
rect 32752 1806 32816 1870
rect 32832 1806 32896 1870
rect 32912 1806 32976 1870
rect 32992 1806 33056 1870
rect 33072 1806 33136 1870
<< metal4 >>
rect 13782 4190 33240 4192
rect 13782 4126 13886 4190
rect 13950 4126 13966 4190
rect 14030 4126 14046 4190
rect 14110 4126 14126 4190
rect 14190 4126 14206 4190
rect 14270 4126 14286 4190
rect 14350 4126 14492 4190
rect 14556 4126 14572 4190
rect 14636 4126 14652 4190
rect 14716 4126 14732 4190
rect 14796 4126 14812 4190
rect 14876 4126 14892 4190
rect 14956 4126 15098 4190
rect 15162 4126 15178 4190
rect 15242 4126 15258 4190
rect 15322 4126 15338 4190
rect 15402 4126 15418 4190
rect 15482 4126 15498 4190
rect 15562 4126 15704 4190
rect 15768 4126 15784 4190
rect 15848 4126 15864 4190
rect 15928 4126 15944 4190
rect 16008 4126 16024 4190
rect 16088 4126 16104 4190
rect 16168 4126 16310 4190
rect 16374 4126 16390 4190
rect 16454 4126 16470 4190
rect 16534 4126 16550 4190
rect 16614 4126 16630 4190
rect 16694 4126 16710 4190
rect 16774 4126 16916 4190
rect 16980 4126 16996 4190
rect 17060 4126 17076 4190
rect 17140 4126 17156 4190
rect 17220 4126 17236 4190
rect 17300 4126 17316 4190
rect 17380 4126 17522 4190
rect 17586 4126 17602 4190
rect 17666 4126 17682 4190
rect 17746 4126 17762 4190
rect 17826 4126 17842 4190
rect 17906 4126 17922 4190
rect 17986 4126 18128 4190
rect 18192 4126 18208 4190
rect 18272 4126 18288 4190
rect 18352 4126 18368 4190
rect 18432 4126 18448 4190
rect 18512 4126 18528 4190
rect 18592 4126 18734 4190
rect 18798 4126 18814 4190
rect 18878 4126 18894 4190
rect 18958 4126 18974 4190
rect 19038 4126 19054 4190
rect 19118 4126 19134 4190
rect 19198 4126 19340 4190
rect 19404 4126 19420 4190
rect 19484 4126 19500 4190
rect 19564 4126 19580 4190
rect 19644 4126 19660 4190
rect 19724 4126 19740 4190
rect 19804 4126 19946 4190
rect 20010 4126 20026 4190
rect 20090 4126 20106 4190
rect 20170 4126 20186 4190
rect 20250 4126 20266 4190
rect 20330 4126 20346 4190
rect 20410 4126 20552 4190
rect 20616 4126 20632 4190
rect 20696 4126 20712 4190
rect 20776 4126 20792 4190
rect 20856 4126 20872 4190
rect 20936 4126 20952 4190
rect 21016 4126 21158 4190
rect 21222 4126 21238 4190
rect 21302 4126 21318 4190
rect 21382 4126 21398 4190
rect 21462 4126 21478 4190
rect 21542 4126 21558 4190
rect 21622 4126 21764 4190
rect 21828 4126 21844 4190
rect 21908 4126 21924 4190
rect 21988 4126 22004 4190
rect 22068 4126 22084 4190
rect 22148 4126 22164 4190
rect 22228 4126 22370 4190
rect 22434 4126 22450 4190
rect 22514 4126 22530 4190
rect 22594 4126 22610 4190
rect 22674 4126 22690 4190
rect 22754 4126 22770 4190
rect 22834 4126 22976 4190
rect 23040 4126 23056 4190
rect 23120 4126 23136 4190
rect 23200 4126 23216 4190
rect 23280 4126 23296 4190
rect 23360 4126 23376 4190
rect 23440 4126 23582 4190
rect 23646 4126 23662 4190
rect 23726 4126 23742 4190
rect 23806 4126 23822 4190
rect 23886 4126 23902 4190
rect 23966 4126 23982 4190
rect 24046 4126 24188 4190
rect 24252 4126 24268 4190
rect 24332 4126 24348 4190
rect 24412 4126 24428 4190
rect 24492 4126 24508 4190
rect 24572 4126 24588 4190
rect 24652 4126 24794 4190
rect 24858 4126 24874 4190
rect 24938 4126 24954 4190
rect 25018 4126 25034 4190
rect 25098 4126 25114 4190
rect 25178 4126 25194 4190
rect 25258 4126 25400 4190
rect 25464 4126 25480 4190
rect 25544 4126 25560 4190
rect 25624 4126 25640 4190
rect 25704 4126 25720 4190
rect 25784 4126 25800 4190
rect 25864 4126 26006 4190
rect 26070 4126 26086 4190
rect 26150 4126 26166 4190
rect 26230 4126 26246 4190
rect 26310 4126 26326 4190
rect 26390 4126 26406 4190
rect 26470 4126 26612 4190
rect 26676 4126 26692 4190
rect 26756 4126 26772 4190
rect 26836 4126 26852 4190
rect 26916 4126 26932 4190
rect 26996 4126 27012 4190
rect 27076 4126 27218 4190
rect 27282 4126 27298 4190
rect 27362 4126 27378 4190
rect 27442 4126 27458 4190
rect 27522 4126 27538 4190
rect 27602 4126 27618 4190
rect 27682 4126 27824 4190
rect 27888 4126 27904 4190
rect 27968 4126 27984 4190
rect 28048 4126 28064 4190
rect 28128 4126 28144 4190
rect 28208 4126 28224 4190
rect 28288 4126 28430 4190
rect 28494 4126 28510 4190
rect 28574 4126 28590 4190
rect 28654 4126 28670 4190
rect 28734 4126 28750 4190
rect 28814 4126 28830 4190
rect 28894 4126 29036 4190
rect 29100 4126 29116 4190
rect 29180 4126 29196 4190
rect 29260 4126 29276 4190
rect 29340 4126 29356 4190
rect 29420 4126 29436 4190
rect 29500 4126 29642 4190
rect 29706 4126 29722 4190
rect 29786 4126 29802 4190
rect 29866 4126 29882 4190
rect 29946 4126 29962 4190
rect 30026 4126 30042 4190
rect 30106 4126 30248 4190
rect 30312 4126 30328 4190
rect 30392 4126 30408 4190
rect 30472 4126 30488 4190
rect 30552 4126 30568 4190
rect 30632 4126 30648 4190
rect 30712 4126 30854 4190
rect 30918 4126 30934 4190
rect 30998 4126 31014 4190
rect 31078 4126 31094 4190
rect 31158 4126 31174 4190
rect 31238 4126 31254 4190
rect 31318 4126 31460 4190
rect 31524 4126 31540 4190
rect 31604 4126 31620 4190
rect 31684 4126 31700 4190
rect 31764 4126 31780 4190
rect 31844 4126 31860 4190
rect 31924 4126 32066 4190
rect 32130 4126 32146 4190
rect 32210 4126 32226 4190
rect 32290 4126 32306 4190
rect 32370 4126 32386 4190
rect 32450 4126 32466 4190
rect 32530 4126 32672 4190
rect 32736 4126 32752 4190
rect 32816 4126 32832 4190
rect 32896 4126 32912 4190
rect 32976 4126 32992 4190
rect 33056 4126 33072 4190
rect 33136 4126 33240 4190
rect 13782 4124 33240 4126
rect 13782 3970 13848 4060
rect 13782 3906 13783 3970
rect 13847 3906 13848 3970
rect 13782 3890 13848 3906
rect 13782 3826 13783 3890
rect 13847 3826 13848 3890
rect 13782 3810 13848 3826
rect 13782 3746 13783 3810
rect 13847 3746 13848 3810
rect 13782 3730 13848 3746
rect 13782 3666 13783 3730
rect 13847 3666 13848 3730
rect 13782 3650 13848 3666
rect 13782 3586 13783 3650
rect 13847 3586 13848 3650
rect 13782 3570 13848 3586
rect 13782 3506 13783 3570
rect 13847 3506 13848 3570
rect 13782 3490 13848 3506
rect 13782 3426 13783 3490
rect 13847 3426 13848 3490
rect 13782 3410 13848 3426
rect 13782 3346 13783 3410
rect 13847 3346 13848 3410
rect 13782 3330 13848 3346
rect 13782 3266 13783 3330
rect 13847 3266 13848 3330
rect 13782 3250 13848 3266
rect 13782 3186 13783 3250
rect 13847 3186 13848 3250
rect 13782 3032 13848 3186
rect 13908 3032 13968 4064
rect 14028 3094 14088 4124
rect 14148 3032 14208 4064
rect 14268 3094 14328 4124
rect 14388 3970 14454 4060
rect 14388 3906 14389 3970
rect 14453 3906 14454 3970
rect 14388 3890 14454 3906
rect 14388 3826 14389 3890
rect 14453 3826 14454 3890
rect 14388 3810 14454 3826
rect 14388 3746 14389 3810
rect 14453 3746 14454 3810
rect 14388 3730 14454 3746
rect 14388 3666 14389 3730
rect 14453 3666 14454 3730
rect 14388 3650 14454 3666
rect 14388 3586 14389 3650
rect 14453 3586 14454 3650
rect 14388 3570 14454 3586
rect 14388 3506 14389 3570
rect 14453 3506 14454 3570
rect 14388 3490 14454 3506
rect 14388 3426 14389 3490
rect 14453 3426 14454 3490
rect 14388 3410 14454 3426
rect 14388 3346 14389 3410
rect 14453 3346 14454 3410
rect 14388 3330 14454 3346
rect 14388 3266 14389 3330
rect 14453 3266 14454 3330
rect 14388 3250 14454 3266
rect 14388 3186 14389 3250
rect 14453 3186 14454 3250
rect 14388 3032 14454 3186
rect 14514 3032 14574 4064
rect 14634 3094 14694 4124
rect 14754 3032 14814 4064
rect 14874 3094 14934 4124
rect 14994 3970 15060 4060
rect 14994 3906 14995 3970
rect 15059 3906 15060 3970
rect 14994 3890 15060 3906
rect 14994 3826 14995 3890
rect 15059 3826 15060 3890
rect 14994 3810 15060 3826
rect 14994 3746 14995 3810
rect 15059 3746 15060 3810
rect 14994 3730 15060 3746
rect 14994 3666 14995 3730
rect 15059 3666 15060 3730
rect 14994 3650 15060 3666
rect 14994 3586 14995 3650
rect 15059 3586 15060 3650
rect 14994 3570 15060 3586
rect 14994 3506 14995 3570
rect 15059 3506 15060 3570
rect 14994 3490 15060 3506
rect 14994 3426 14995 3490
rect 15059 3426 15060 3490
rect 14994 3410 15060 3426
rect 14994 3346 14995 3410
rect 15059 3346 15060 3410
rect 14994 3330 15060 3346
rect 14994 3266 14995 3330
rect 15059 3266 15060 3330
rect 14994 3250 15060 3266
rect 14994 3186 14995 3250
rect 15059 3186 15060 3250
rect 14994 3032 15060 3186
rect 15120 3032 15180 4064
rect 15240 3094 15300 4124
rect 15360 3032 15420 4064
rect 15480 3094 15540 4124
rect 15600 3970 15666 4060
rect 15600 3906 15601 3970
rect 15665 3906 15666 3970
rect 15600 3890 15666 3906
rect 15600 3826 15601 3890
rect 15665 3826 15666 3890
rect 15600 3810 15666 3826
rect 15600 3746 15601 3810
rect 15665 3746 15666 3810
rect 15600 3730 15666 3746
rect 15600 3666 15601 3730
rect 15665 3666 15666 3730
rect 15600 3650 15666 3666
rect 15600 3586 15601 3650
rect 15665 3586 15666 3650
rect 15600 3570 15666 3586
rect 15600 3506 15601 3570
rect 15665 3506 15666 3570
rect 15600 3490 15666 3506
rect 15600 3426 15601 3490
rect 15665 3426 15666 3490
rect 15600 3410 15666 3426
rect 15600 3346 15601 3410
rect 15665 3346 15666 3410
rect 15600 3330 15666 3346
rect 15600 3266 15601 3330
rect 15665 3266 15666 3330
rect 15600 3250 15666 3266
rect 15600 3186 15601 3250
rect 15665 3186 15666 3250
rect 15600 3032 15666 3186
rect 15726 3032 15786 4064
rect 15846 3094 15906 4124
rect 15966 3032 16026 4064
rect 16086 3094 16146 4124
rect 16206 3970 16272 4060
rect 16206 3906 16207 3970
rect 16271 3906 16272 3970
rect 16206 3890 16272 3906
rect 16206 3826 16207 3890
rect 16271 3826 16272 3890
rect 16206 3810 16272 3826
rect 16206 3746 16207 3810
rect 16271 3746 16272 3810
rect 16206 3730 16272 3746
rect 16206 3666 16207 3730
rect 16271 3666 16272 3730
rect 16206 3650 16272 3666
rect 16206 3586 16207 3650
rect 16271 3586 16272 3650
rect 16206 3570 16272 3586
rect 16206 3506 16207 3570
rect 16271 3506 16272 3570
rect 16206 3490 16272 3506
rect 16206 3426 16207 3490
rect 16271 3426 16272 3490
rect 16206 3410 16272 3426
rect 16206 3346 16207 3410
rect 16271 3346 16272 3410
rect 16206 3330 16272 3346
rect 16206 3266 16207 3330
rect 16271 3266 16272 3330
rect 16206 3250 16272 3266
rect 16206 3186 16207 3250
rect 16271 3186 16272 3250
rect 16206 3032 16272 3186
rect 16332 3032 16392 4064
rect 16452 3094 16512 4124
rect 16572 3032 16632 4064
rect 16692 3094 16752 4124
rect 16812 3970 16878 4060
rect 16812 3906 16813 3970
rect 16877 3906 16878 3970
rect 16812 3890 16878 3906
rect 16812 3826 16813 3890
rect 16877 3826 16878 3890
rect 16812 3810 16878 3826
rect 16812 3746 16813 3810
rect 16877 3746 16878 3810
rect 16812 3730 16878 3746
rect 16812 3666 16813 3730
rect 16877 3666 16878 3730
rect 16812 3650 16878 3666
rect 16812 3586 16813 3650
rect 16877 3586 16878 3650
rect 16812 3570 16878 3586
rect 16812 3506 16813 3570
rect 16877 3506 16878 3570
rect 16812 3490 16878 3506
rect 16812 3426 16813 3490
rect 16877 3426 16878 3490
rect 16812 3410 16878 3426
rect 16812 3346 16813 3410
rect 16877 3346 16878 3410
rect 16812 3330 16878 3346
rect 16812 3266 16813 3330
rect 16877 3266 16878 3330
rect 16812 3250 16878 3266
rect 16812 3186 16813 3250
rect 16877 3186 16878 3250
rect 16812 3032 16878 3186
rect 16938 3032 16998 4064
rect 17058 3094 17118 4124
rect 17178 3032 17238 4064
rect 17298 3094 17358 4124
rect 17418 3970 17484 4060
rect 17418 3906 17419 3970
rect 17483 3906 17484 3970
rect 17418 3890 17484 3906
rect 17418 3826 17419 3890
rect 17483 3826 17484 3890
rect 17418 3810 17484 3826
rect 17418 3746 17419 3810
rect 17483 3746 17484 3810
rect 17418 3730 17484 3746
rect 17418 3666 17419 3730
rect 17483 3666 17484 3730
rect 17418 3650 17484 3666
rect 17418 3586 17419 3650
rect 17483 3586 17484 3650
rect 17418 3570 17484 3586
rect 17418 3506 17419 3570
rect 17483 3506 17484 3570
rect 17418 3490 17484 3506
rect 17418 3426 17419 3490
rect 17483 3426 17484 3490
rect 17418 3410 17484 3426
rect 17418 3346 17419 3410
rect 17483 3346 17484 3410
rect 17418 3330 17484 3346
rect 17418 3266 17419 3330
rect 17483 3266 17484 3330
rect 17418 3250 17484 3266
rect 17418 3186 17419 3250
rect 17483 3186 17484 3250
rect 17418 3032 17484 3186
rect 17544 3032 17604 4064
rect 17664 3094 17724 4124
rect 17784 3032 17844 4064
rect 17904 3094 17964 4124
rect 18024 3970 18090 4060
rect 18024 3906 18025 3970
rect 18089 3906 18090 3970
rect 18024 3890 18090 3906
rect 18024 3826 18025 3890
rect 18089 3826 18090 3890
rect 18024 3810 18090 3826
rect 18024 3746 18025 3810
rect 18089 3746 18090 3810
rect 18024 3730 18090 3746
rect 18024 3666 18025 3730
rect 18089 3666 18090 3730
rect 18024 3650 18090 3666
rect 18024 3586 18025 3650
rect 18089 3586 18090 3650
rect 18024 3570 18090 3586
rect 18024 3506 18025 3570
rect 18089 3506 18090 3570
rect 18024 3490 18090 3506
rect 18024 3426 18025 3490
rect 18089 3426 18090 3490
rect 18024 3410 18090 3426
rect 18024 3346 18025 3410
rect 18089 3346 18090 3410
rect 18024 3330 18090 3346
rect 18024 3266 18025 3330
rect 18089 3266 18090 3330
rect 18024 3250 18090 3266
rect 18024 3186 18025 3250
rect 18089 3186 18090 3250
rect 18024 3032 18090 3186
rect 18150 3032 18210 4064
rect 18270 3094 18330 4124
rect 18390 3032 18450 4064
rect 18510 3094 18570 4124
rect 18630 3970 18696 4060
rect 18630 3906 18631 3970
rect 18695 3906 18696 3970
rect 18630 3890 18696 3906
rect 18630 3826 18631 3890
rect 18695 3826 18696 3890
rect 18630 3810 18696 3826
rect 18630 3746 18631 3810
rect 18695 3746 18696 3810
rect 18630 3730 18696 3746
rect 18630 3666 18631 3730
rect 18695 3666 18696 3730
rect 18630 3650 18696 3666
rect 18630 3586 18631 3650
rect 18695 3586 18696 3650
rect 18630 3570 18696 3586
rect 18630 3506 18631 3570
rect 18695 3506 18696 3570
rect 18630 3490 18696 3506
rect 18630 3426 18631 3490
rect 18695 3426 18696 3490
rect 18630 3410 18696 3426
rect 18630 3346 18631 3410
rect 18695 3346 18696 3410
rect 18630 3330 18696 3346
rect 18630 3266 18631 3330
rect 18695 3266 18696 3330
rect 18630 3250 18696 3266
rect 18630 3186 18631 3250
rect 18695 3186 18696 3250
rect 18630 3032 18696 3186
rect 18756 3032 18816 4064
rect 18876 3094 18936 4124
rect 18996 3032 19056 4064
rect 19116 3094 19176 4124
rect 19236 3970 19302 4060
rect 19236 3906 19237 3970
rect 19301 3906 19302 3970
rect 19236 3890 19302 3906
rect 19236 3826 19237 3890
rect 19301 3826 19302 3890
rect 19236 3810 19302 3826
rect 19236 3746 19237 3810
rect 19301 3746 19302 3810
rect 19236 3730 19302 3746
rect 19236 3666 19237 3730
rect 19301 3666 19302 3730
rect 19236 3650 19302 3666
rect 19236 3586 19237 3650
rect 19301 3586 19302 3650
rect 19236 3570 19302 3586
rect 19236 3506 19237 3570
rect 19301 3506 19302 3570
rect 19236 3490 19302 3506
rect 19236 3426 19237 3490
rect 19301 3426 19302 3490
rect 19236 3410 19302 3426
rect 19236 3346 19237 3410
rect 19301 3346 19302 3410
rect 19236 3330 19302 3346
rect 19236 3266 19237 3330
rect 19301 3266 19302 3330
rect 19236 3250 19302 3266
rect 19236 3186 19237 3250
rect 19301 3186 19302 3250
rect 19236 3032 19302 3186
rect 19362 3032 19422 4064
rect 19482 3094 19542 4124
rect 19602 3032 19662 4064
rect 19722 3094 19782 4124
rect 19842 3970 19908 4060
rect 19842 3906 19843 3970
rect 19907 3906 19908 3970
rect 19842 3890 19908 3906
rect 19842 3826 19843 3890
rect 19907 3826 19908 3890
rect 19842 3810 19908 3826
rect 19842 3746 19843 3810
rect 19907 3746 19908 3810
rect 19842 3730 19908 3746
rect 19842 3666 19843 3730
rect 19907 3666 19908 3730
rect 19842 3650 19908 3666
rect 19842 3586 19843 3650
rect 19907 3586 19908 3650
rect 19842 3570 19908 3586
rect 19842 3506 19843 3570
rect 19907 3506 19908 3570
rect 19842 3490 19908 3506
rect 19842 3426 19843 3490
rect 19907 3426 19908 3490
rect 19842 3410 19908 3426
rect 19842 3346 19843 3410
rect 19907 3346 19908 3410
rect 19842 3330 19908 3346
rect 19842 3266 19843 3330
rect 19907 3266 19908 3330
rect 19842 3250 19908 3266
rect 19842 3186 19843 3250
rect 19907 3186 19908 3250
rect 19842 3032 19908 3186
rect 19968 3032 20028 4064
rect 20088 3094 20148 4124
rect 20208 3032 20268 4064
rect 20328 3094 20388 4124
rect 20448 3970 20514 4060
rect 20448 3906 20449 3970
rect 20513 3906 20514 3970
rect 20448 3890 20514 3906
rect 20448 3826 20449 3890
rect 20513 3826 20514 3890
rect 20448 3810 20514 3826
rect 20448 3746 20449 3810
rect 20513 3746 20514 3810
rect 20448 3730 20514 3746
rect 20448 3666 20449 3730
rect 20513 3666 20514 3730
rect 20448 3650 20514 3666
rect 20448 3586 20449 3650
rect 20513 3586 20514 3650
rect 20448 3570 20514 3586
rect 20448 3506 20449 3570
rect 20513 3506 20514 3570
rect 20448 3490 20514 3506
rect 20448 3426 20449 3490
rect 20513 3426 20514 3490
rect 20448 3410 20514 3426
rect 20448 3346 20449 3410
rect 20513 3346 20514 3410
rect 20448 3330 20514 3346
rect 20448 3266 20449 3330
rect 20513 3266 20514 3330
rect 20448 3250 20514 3266
rect 20448 3186 20449 3250
rect 20513 3186 20514 3250
rect 20448 3032 20514 3186
rect 20574 3032 20634 4064
rect 20694 3094 20754 4124
rect 20814 3032 20874 4064
rect 20934 3094 20994 4124
rect 21054 3970 21120 4060
rect 21054 3906 21055 3970
rect 21119 3906 21120 3970
rect 21054 3890 21120 3906
rect 21054 3826 21055 3890
rect 21119 3826 21120 3890
rect 21054 3810 21120 3826
rect 21054 3746 21055 3810
rect 21119 3746 21120 3810
rect 21054 3730 21120 3746
rect 21054 3666 21055 3730
rect 21119 3666 21120 3730
rect 21054 3650 21120 3666
rect 21054 3586 21055 3650
rect 21119 3586 21120 3650
rect 21054 3570 21120 3586
rect 21054 3506 21055 3570
rect 21119 3506 21120 3570
rect 21054 3490 21120 3506
rect 21054 3426 21055 3490
rect 21119 3426 21120 3490
rect 21054 3410 21120 3426
rect 21054 3346 21055 3410
rect 21119 3346 21120 3410
rect 21054 3330 21120 3346
rect 21054 3266 21055 3330
rect 21119 3266 21120 3330
rect 21054 3250 21120 3266
rect 21054 3186 21055 3250
rect 21119 3186 21120 3250
rect 21054 3032 21120 3186
rect 21180 3032 21240 4064
rect 21300 3094 21360 4124
rect 21420 3032 21480 4064
rect 21540 3094 21600 4124
rect 21660 3970 21726 4060
rect 21660 3906 21661 3970
rect 21725 3906 21726 3970
rect 21660 3890 21726 3906
rect 21660 3826 21661 3890
rect 21725 3826 21726 3890
rect 21660 3810 21726 3826
rect 21660 3746 21661 3810
rect 21725 3746 21726 3810
rect 21660 3730 21726 3746
rect 21660 3666 21661 3730
rect 21725 3666 21726 3730
rect 21660 3650 21726 3666
rect 21660 3586 21661 3650
rect 21725 3586 21726 3650
rect 21660 3570 21726 3586
rect 21660 3506 21661 3570
rect 21725 3506 21726 3570
rect 21660 3490 21726 3506
rect 21660 3426 21661 3490
rect 21725 3426 21726 3490
rect 21660 3410 21726 3426
rect 21660 3346 21661 3410
rect 21725 3346 21726 3410
rect 21660 3330 21726 3346
rect 21660 3266 21661 3330
rect 21725 3266 21726 3330
rect 21660 3250 21726 3266
rect 21660 3186 21661 3250
rect 21725 3186 21726 3250
rect 21660 3032 21726 3186
rect 21786 3032 21846 4064
rect 21906 3094 21966 4124
rect 22026 3032 22086 4064
rect 22146 3094 22206 4124
rect 22266 3970 22332 4060
rect 22266 3906 22267 3970
rect 22331 3906 22332 3970
rect 22266 3890 22332 3906
rect 22266 3826 22267 3890
rect 22331 3826 22332 3890
rect 22266 3810 22332 3826
rect 22266 3746 22267 3810
rect 22331 3746 22332 3810
rect 22266 3730 22332 3746
rect 22266 3666 22267 3730
rect 22331 3666 22332 3730
rect 22266 3650 22332 3666
rect 22266 3586 22267 3650
rect 22331 3586 22332 3650
rect 22266 3570 22332 3586
rect 22266 3506 22267 3570
rect 22331 3506 22332 3570
rect 22266 3490 22332 3506
rect 22266 3426 22267 3490
rect 22331 3426 22332 3490
rect 22266 3410 22332 3426
rect 22266 3346 22267 3410
rect 22331 3346 22332 3410
rect 22266 3330 22332 3346
rect 22266 3266 22267 3330
rect 22331 3266 22332 3330
rect 22266 3250 22332 3266
rect 22266 3186 22267 3250
rect 22331 3186 22332 3250
rect 22266 3032 22332 3186
rect 22392 3032 22452 4064
rect 22512 3094 22572 4124
rect 22632 3032 22692 4064
rect 22752 3094 22812 4124
rect 22872 3970 22938 4060
rect 22872 3906 22873 3970
rect 22937 3906 22938 3970
rect 22872 3890 22938 3906
rect 22872 3826 22873 3890
rect 22937 3826 22938 3890
rect 22872 3810 22938 3826
rect 22872 3746 22873 3810
rect 22937 3746 22938 3810
rect 22872 3730 22938 3746
rect 22872 3666 22873 3730
rect 22937 3666 22938 3730
rect 22872 3650 22938 3666
rect 22872 3586 22873 3650
rect 22937 3586 22938 3650
rect 22872 3570 22938 3586
rect 22872 3506 22873 3570
rect 22937 3506 22938 3570
rect 22872 3490 22938 3506
rect 22872 3426 22873 3490
rect 22937 3426 22938 3490
rect 22872 3410 22938 3426
rect 22872 3346 22873 3410
rect 22937 3346 22938 3410
rect 22872 3330 22938 3346
rect 22872 3266 22873 3330
rect 22937 3266 22938 3330
rect 22872 3250 22938 3266
rect 22872 3186 22873 3250
rect 22937 3186 22938 3250
rect 22872 3032 22938 3186
rect 22998 3032 23058 4064
rect 23118 3094 23178 4124
rect 23238 3032 23298 4064
rect 23358 3094 23418 4124
rect 23478 3970 23544 4060
rect 23478 3906 23479 3970
rect 23543 3906 23544 3970
rect 23478 3890 23544 3906
rect 23478 3826 23479 3890
rect 23543 3826 23544 3890
rect 23478 3810 23544 3826
rect 23478 3746 23479 3810
rect 23543 3746 23544 3810
rect 23478 3730 23544 3746
rect 23478 3666 23479 3730
rect 23543 3666 23544 3730
rect 23478 3650 23544 3666
rect 23478 3586 23479 3650
rect 23543 3586 23544 3650
rect 23478 3570 23544 3586
rect 23478 3506 23479 3570
rect 23543 3506 23544 3570
rect 23478 3490 23544 3506
rect 23478 3426 23479 3490
rect 23543 3426 23544 3490
rect 23478 3410 23544 3426
rect 23478 3346 23479 3410
rect 23543 3346 23544 3410
rect 23478 3330 23544 3346
rect 23478 3266 23479 3330
rect 23543 3266 23544 3330
rect 23478 3250 23544 3266
rect 23478 3186 23479 3250
rect 23543 3186 23544 3250
rect 23478 3032 23544 3186
rect 23604 3032 23664 4064
rect 23724 3094 23784 4124
rect 23844 3032 23904 4064
rect 23964 3094 24024 4124
rect 24084 3970 24150 4060
rect 24084 3906 24085 3970
rect 24149 3906 24150 3970
rect 24084 3890 24150 3906
rect 24084 3826 24085 3890
rect 24149 3826 24150 3890
rect 24084 3810 24150 3826
rect 24084 3746 24085 3810
rect 24149 3746 24150 3810
rect 24084 3730 24150 3746
rect 24084 3666 24085 3730
rect 24149 3666 24150 3730
rect 24084 3650 24150 3666
rect 24084 3586 24085 3650
rect 24149 3586 24150 3650
rect 24084 3570 24150 3586
rect 24084 3506 24085 3570
rect 24149 3506 24150 3570
rect 24084 3490 24150 3506
rect 24084 3426 24085 3490
rect 24149 3426 24150 3490
rect 24084 3410 24150 3426
rect 24084 3346 24085 3410
rect 24149 3346 24150 3410
rect 24084 3330 24150 3346
rect 24084 3266 24085 3330
rect 24149 3266 24150 3330
rect 24084 3250 24150 3266
rect 24084 3186 24085 3250
rect 24149 3186 24150 3250
rect 24084 3032 24150 3186
rect 24210 3032 24270 4064
rect 24330 3094 24390 4124
rect 24450 3032 24510 4064
rect 24570 3094 24630 4124
rect 24690 3970 24756 4060
rect 24690 3906 24691 3970
rect 24755 3906 24756 3970
rect 24690 3890 24756 3906
rect 24690 3826 24691 3890
rect 24755 3826 24756 3890
rect 24690 3810 24756 3826
rect 24690 3746 24691 3810
rect 24755 3746 24756 3810
rect 24690 3730 24756 3746
rect 24690 3666 24691 3730
rect 24755 3666 24756 3730
rect 24690 3650 24756 3666
rect 24690 3586 24691 3650
rect 24755 3586 24756 3650
rect 24690 3570 24756 3586
rect 24690 3506 24691 3570
rect 24755 3506 24756 3570
rect 24690 3490 24756 3506
rect 24690 3426 24691 3490
rect 24755 3426 24756 3490
rect 24690 3410 24756 3426
rect 24690 3346 24691 3410
rect 24755 3346 24756 3410
rect 24690 3330 24756 3346
rect 24690 3266 24691 3330
rect 24755 3266 24756 3330
rect 24690 3250 24756 3266
rect 24690 3186 24691 3250
rect 24755 3186 24756 3250
rect 24690 3032 24756 3186
rect 24816 3032 24876 4064
rect 24936 3094 24996 4124
rect 25056 3032 25116 4064
rect 25176 3094 25236 4124
rect 25296 3970 25362 4060
rect 25296 3906 25297 3970
rect 25361 3906 25362 3970
rect 25296 3890 25362 3906
rect 25296 3826 25297 3890
rect 25361 3826 25362 3890
rect 25296 3810 25362 3826
rect 25296 3746 25297 3810
rect 25361 3746 25362 3810
rect 25296 3730 25362 3746
rect 25296 3666 25297 3730
rect 25361 3666 25362 3730
rect 25296 3650 25362 3666
rect 25296 3586 25297 3650
rect 25361 3586 25362 3650
rect 25296 3570 25362 3586
rect 25296 3506 25297 3570
rect 25361 3506 25362 3570
rect 25296 3490 25362 3506
rect 25296 3426 25297 3490
rect 25361 3426 25362 3490
rect 25296 3410 25362 3426
rect 25296 3346 25297 3410
rect 25361 3346 25362 3410
rect 25296 3330 25362 3346
rect 25296 3266 25297 3330
rect 25361 3266 25362 3330
rect 25296 3250 25362 3266
rect 25296 3186 25297 3250
rect 25361 3186 25362 3250
rect 25296 3032 25362 3186
rect 25422 3032 25482 4064
rect 25542 3094 25602 4124
rect 25662 3032 25722 4064
rect 25782 3094 25842 4124
rect 25902 3970 25968 4060
rect 25902 3906 25903 3970
rect 25967 3906 25968 3970
rect 25902 3890 25968 3906
rect 25902 3826 25903 3890
rect 25967 3826 25968 3890
rect 25902 3810 25968 3826
rect 25902 3746 25903 3810
rect 25967 3746 25968 3810
rect 25902 3730 25968 3746
rect 25902 3666 25903 3730
rect 25967 3666 25968 3730
rect 25902 3650 25968 3666
rect 25902 3586 25903 3650
rect 25967 3586 25968 3650
rect 25902 3570 25968 3586
rect 25902 3506 25903 3570
rect 25967 3506 25968 3570
rect 25902 3490 25968 3506
rect 25902 3426 25903 3490
rect 25967 3426 25968 3490
rect 25902 3410 25968 3426
rect 25902 3346 25903 3410
rect 25967 3346 25968 3410
rect 25902 3330 25968 3346
rect 25902 3266 25903 3330
rect 25967 3266 25968 3330
rect 25902 3250 25968 3266
rect 25902 3186 25903 3250
rect 25967 3186 25968 3250
rect 25902 3032 25968 3186
rect 26028 3032 26088 4064
rect 26148 3094 26208 4124
rect 26268 3032 26328 4064
rect 26388 3094 26448 4124
rect 26508 3970 26574 4060
rect 26508 3906 26509 3970
rect 26573 3906 26574 3970
rect 26508 3890 26574 3906
rect 26508 3826 26509 3890
rect 26573 3826 26574 3890
rect 26508 3810 26574 3826
rect 26508 3746 26509 3810
rect 26573 3746 26574 3810
rect 26508 3730 26574 3746
rect 26508 3666 26509 3730
rect 26573 3666 26574 3730
rect 26508 3650 26574 3666
rect 26508 3586 26509 3650
rect 26573 3586 26574 3650
rect 26508 3570 26574 3586
rect 26508 3506 26509 3570
rect 26573 3506 26574 3570
rect 26508 3490 26574 3506
rect 26508 3426 26509 3490
rect 26573 3426 26574 3490
rect 26508 3410 26574 3426
rect 26508 3346 26509 3410
rect 26573 3346 26574 3410
rect 26508 3330 26574 3346
rect 26508 3266 26509 3330
rect 26573 3266 26574 3330
rect 26508 3250 26574 3266
rect 26508 3186 26509 3250
rect 26573 3186 26574 3250
rect 26508 3032 26574 3186
rect 26634 3032 26694 4064
rect 26754 3094 26814 4124
rect 26874 3032 26934 4064
rect 26994 3094 27054 4124
rect 27114 3970 27180 4060
rect 27114 3906 27115 3970
rect 27179 3906 27180 3970
rect 27114 3890 27180 3906
rect 27114 3826 27115 3890
rect 27179 3826 27180 3890
rect 27114 3810 27180 3826
rect 27114 3746 27115 3810
rect 27179 3746 27180 3810
rect 27114 3730 27180 3746
rect 27114 3666 27115 3730
rect 27179 3666 27180 3730
rect 27114 3650 27180 3666
rect 27114 3586 27115 3650
rect 27179 3586 27180 3650
rect 27114 3570 27180 3586
rect 27114 3506 27115 3570
rect 27179 3506 27180 3570
rect 27114 3490 27180 3506
rect 27114 3426 27115 3490
rect 27179 3426 27180 3490
rect 27114 3410 27180 3426
rect 27114 3346 27115 3410
rect 27179 3346 27180 3410
rect 27114 3330 27180 3346
rect 27114 3266 27115 3330
rect 27179 3266 27180 3330
rect 27114 3250 27180 3266
rect 27114 3186 27115 3250
rect 27179 3186 27180 3250
rect 27114 3032 27180 3186
rect 27240 3032 27300 4064
rect 27360 3094 27420 4124
rect 27480 3032 27540 4064
rect 27600 3094 27660 4124
rect 27720 3970 27786 4060
rect 27720 3906 27721 3970
rect 27785 3906 27786 3970
rect 27720 3890 27786 3906
rect 27720 3826 27721 3890
rect 27785 3826 27786 3890
rect 27720 3810 27786 3826
rect 27720 3746 27721 3810
rect 27785 3746 27786 3810
rect 27720 3730 27786 3746
rect 27720 3666 27721 3730
rect 27785 3666 27786 3730
rect 27720 3650 27786 3666
rect 27720 3586 27721 3650
rect 27785 3586 27786 3650
rect 27720 3570 27786 3586
rect 27720 3506 27721 3570
rect 27785 3506 27786 3570
rect 27720 3490 27786 3506
rect 27720 3426 27721 3490
rect 27785 3426 27786 3490
rect 27720 3410 27786 3426
rect 27720 3346 27721 3410
rect 27785 3346 27786 3410
rect 27720 3330 27786 3346
rect 27720 3266 27721 3330
rect 27785 3266 27786 3330
rect 27720 3250 27786 3266
rect 27720 3186 27721 3250
rect 27785 3186 27786 3250
rect 27720 3032 27786 3186
rect 27846 3032 27906 4064
rect 27966 3094 28026 4124
rect 28086 3032 28146 4064
rect 28206 3094 28266 4124
rect 28326 3970 28392 4060
rect 28326 3906 28327 3970
rect 28391 3906 28392 3970
rect 28326 3890 28392 3906
rect 28326 3826 28327 3890
rect 28391 3826 28392 3890
rect 28326 3810 28392 3826
rect 28326 3746 28327 3810
rect 28391 3746 28392 3810
rect 28326 3730 28392 3746
rect 28326 3666 28327 3730
rect 28391 3666 28392 3730
rect 28326 3650 28392 3666
rect 28326 3586 28327 3650
rect 28391 3586 28392 3650
rect 28326 3570 28392 3586
rect 28326 3506 28327 3570
rect 28391 3506 28392 3570
rect 28326 3490 28392 3506
rect 28326 3426 28327 3490
rect 28391 3426 28392 3490
rect 28326 3410 28392 3426
rect 28326 3346 28327 3410
rect 28391 3346 28392 3410
rect 28326 3330 28392 3346
rect 28326 3266 28327 3330
rect 28391 3266 28392 3330
rect 28326 3250 28392 3266
rect 28326 3186 28327 3250
rect 28391 3186 28392 3250
rect 28326 3032 28392 3186
rect 28452 3032 28512 4064
rect 28572 3094 28632 4124
rect 28692 3032 28752 4064
rect 28812 3094 28872 4124
rect 28932 3970 28998 4060
rect 28932 3906 28933 3970
rect 28997 3906 28998 3970
rect 28932 3890 28998 3906
rect 28932 3826 28933 3890
rect 28997 3826 28998 3890
rect 28932 3810 28998 3826
rect 28932 3746 28933 3810
rect 28997 3746 28998 3810
rect 28932 3730 28998 3746
rect 28932 3666 28933 3730
rect 28997 3666 28998 3730
rect 28932 3650 28998 3666
rect 28932 3586 28933 3650
rect 28997 3586 28998 3650
rect 28932 3570 28998 3586
rect 28932 3506 28933 3570
rect 28997 3506 28998 3570
rect 28932 3490 28998 3506
rect 28932 3426 28933 3490
rect 28997 3426 28998 3490
rect 28932 3410 28998 3426
rect 28932 3346 28933 3410
rect 28997 3346 28998 3410
rect 28932 3330 28998 3346
rect 28932 3266 28933 3330
rect 28997 3266 28998 3330
rect 28932 3250 28998 3266
rect 28932 3186 28933 3250
rect 28997 3186 28998 3250
rect 28932 3032 28998 3186
rect 29058 3032 29118 4064
rect 29178 3094 29238 4124
rect 29298 3032 29358 4064
rect 29418 3094 29478 4124
rect 29538 3970 29604 4060
rect 29538 3906 29539 3970
rect 29603 3906 29604 3970
rect 29538 3890 29604 3906
rect 29538 3826 29539 3890
rect 29603 3826 29604 3890
rect 29538 3810 29604 3826
rect 29538 3746 29539 3810
rect 29603 3746 29604 3810
rect 29538 3730 29604 3746
rect 29538 3666 29539 3730
rect 29603 3666 29604 3730
rect 29538 3650 29604 3666
rect 29538 3586 29539 3650
rect 29603 3586 29604 3650
rect 29538 3570 29604 3586
rect 29538 3506 29539 3570
rect 29603 3506 29604 3570
rect 29538 3490 29604 3506
rect 29538 3426 29539 3490
rect 29603 3426 29604 3490
rect 29538 3410 29604 3426
rect 29538 3346 29539 3410
rect 29603 3346 29604 3410
rect 29538 3330 29604 3346
rect 29538 3266 29539 3330
rect 29603 3266 29604 3330
rect 29538 3250 29604 3266
rect 29538 3186 29539 3250
rect 29603 3186 29604 3250
rect 29538 3032 29604 3186
rect 29664 3032 29724 4064
rect 29784 3094 29844 4124
rect 29904 3032 29964 4064
rect 30024 3094 30084 4124
rect 30144 3970 30210 4060
rect 30144 3906 30145 3970
rect 30209 3906 30210 3970
rect 30144 3890 30210 3906
rect 30144 3826 30145 3890
rect 30209 3826 30210 3890
rect 30144 3810 30210 3826
rect 30144 3746 30145 3810
rect 30209 3746 30210 3810
rect 30144 3730 30210 3746
rect 30144 3666 30145 3730
rect 30209 3666 30210 3730
rect 30144 3650 30210 3666
rect 30144 3586 30145 3650
rect 30209 3586 30210 3650
rect 30144 3570 30210 3586
rect 30144 3506 30145 3570
rect 30209 3506 30210 3570
rect 30144 3490 30210 3506
rect 30144 3426 30145 3490
rect 30209 3426 30210 3490
rect 30144 3410 30210 3426
rect 30144 3346 30145 3410
rect 30209 3346 30210 3410
rect 30144 3330 30210 3346
rect 30144 3266 30145 3330
rect 30209 3266 30210 3330
rect 30144 3250 30210 3266
rect 30144 3186 30145 3250
rect 30209 3186 30210 3250
rect 30144 3032 30210 3186
rect 30270 3032 30330 4064
rect 30390 3094 30450 4124
rect 30510 3032 30570 4064
rect 30630 3094 30690 4124
rect 30750 3970 30816 4060
rect 30750 3906 30751 3970
rect 30815 3906 30816 3970
rect 30750 3890 30816 3906
rect 30750 3826 30751 3890
rect 30815 3826 30816 3890
rect 30750 3810 30816 3826
rect 30750 3746 30751 3810
rect 30815 3746 30816 3810
rect 30750 3730 30816 3746
rect 30750 3666 30751 3730
rect 30815 3666 30816 3730
rect 30750 3650 30816 3666
rect 30750 3586 30751 3650
rect 30815 3586 30816 3650
rect 30750 3570 30816 3586
rect 30750 3506 30751 3570
rect 30815 3506 30816 3570
rect 30750 3490 30816 3506
rect 30750 3426 30751 3490
rect 30815 3426 30816 3490
rect 30750 3410 30816 3426
rect 30750 3346 30751 3410
rect 30815 3346 30816 3410
rect 30750 3330 30816 3346
rect 30750 3266 30751 3330
rect 30815 3266 30816 3330
rect 30750 3250 30816 3266
rect 30750 3186 30751 3250
rect 30815 3186 30816 3250
rect 30750 3032 30816 3186
rect 30876 3032 30936 4064
rect 30996 3094 31056 4124
rect 31116 3032 31176 4064
rect 31236 3094 31296 4124
rect 31356 3970 31422 4060
rect 31356 3906 31357 3970
rect 31421 3906 31422 3970
rect 31356 3890 31422 3906
rect 31356 3826 31357 3890
rect 31421 3826 31422 3890
rect 31356 3810 31422 3826
rect 31356 3746 31357 3810
rect 31421 3746 31422 3810
rect 31356 3730 31422 3746
rect 31356 3666 31357 3730
rect 31421 3666 31422 3730
rect 31356 3650 31422 3666
rect 31356 3586 31357 3650
rect 31421 3586 31422 3650
rect 31356 3570 31422 3586
rect 31356 3506 31357 3570
rect 31421 3506 31422 3570
rect 31356 3490 31422 3506
rect 31356 3426 31357 3490
rect 31421 3426 31422 3490
rect 31356 3410 31422 3426
rect 31356 3346 31357 3410
rect 31421 3346 31422 3410
rect 31356 3330 31422 3346
rect 31356 3266 31357 3330
rect 31421 3266 31422 3330
rect 31356 3250 31422 3266
rect 31356 3186 31357 3250
rect 31421 3186 31422 3250
rect 31356 3032 31422 3186
rect 31482 3032 31542 4064
rect 31602 3094 31662 4124
rect 31722 3032 31782 4064
rect 31842 3094 31902 4124
rect 31962 3970 32028 4060
rect 31962 3906 31963 3970
rect 32027 3906 32028 3970
rect 31962 3890 32028 3906
rect 31962 3826 31963 3890
rect 32027 3826 32028 3890
rect 31962 3810 32028 3826
rect 31962 3746 31963 3810
rect 32027 3746 32028 3810
rect 31962 3730 32028 3746
rect 31962 3666 31963 3730
rect 32027 3666 32028 3730
rect 31962 3650 32028 3666
rect 31962 3586 31963 3650
rect 32027 3586 32028 3650
rect 31962 3570 32028 3586
rect 31962 3506 31963 3570
rect 32027 3506 32028 3570
rect 31962 3490 32028 3506
rect 31962 3426 31963 3490
rect 32027 3426 32028 3490
rect 31962 3410 32028 3426
rect 31962 3346 31963 3410
rect 32027 3346 32028 3410
rect 31962 3330 32028 3346
rect 31962 3266 31963 3330
rect 32027 3266 32028 3330
rect 31962 3250 32028 3266
rect 31962 3186 31963 3250
rect 32027 3186 32028 3250
rect 31962 3032 32028 3186
rect 32088 3032 32148 4064
rect 32208 3094 32268 4124
rect 32328 3032 32388 4064
rect 32448 3094 32508 4124
rect 32568 3970 32634 4060
rect 32568 3906 32569 3970
rect 32633 3906 32634 3970
rect 32568 3890 32634 3906
rect 32568 3826 32569 3890
rect 32633 3826 32634 3890
rect 32568 3810 32634 3826
rect 32568 3746 32569 3810
rect 32633 3746 32634 3810
rect 32568 3730 32634 3746
rect 32568 3666 32569 3730
rect 32633 3666 32634 3730
rect 32568 3650 32634 3666
rect 32568 3586 32569 3650
rect 32633 3586 32634 3650
rect 32568 3570 32634 3586
rect 32568 3506 32569 3570
rect 32633 3506 32634 3570
rect 32568 3490 32634 3506
rect 32568 3426 32569 3490
rect 32633 3426 32634 3490
rect 32568 3410 32634 3426
rect 32568 3346 32569 3410
rect 32633 3346 32634 3410
rect 32568 3330 32634 3346
rect 32568 3266 32569 3330
rect 32633 3266 32634 3330
rect 32568 3250 32634 3266
rect 32568 3186 32569 3250
rect 32633 3186 32634 3250
rect 32568 3032 32634 3186
rect 32694 3032 32754 4064
rect 32814 3094 32874 4124
rect 32934 3032 32994 4064
rect 33054 3094 33114 4124
rect 33174 3970 33240 4060
rect 33174 3906 33175 3970
rect 33239 3906 33240 3970
rect 33174 3890 33240 3906
rect 33174 3826 33175 3890
rect 33239 3826 33240 3890
rect 33174 3810 33240 3826
rect 33174 3746 33175 3810
rect 33239 3746 33240 3810
rect 33174 3730 33240 3746
rect 33174 3666 33175 3730
rect 33239 3666 33240 3730
rect 33174 3650 33240 3666
rect 33174 3586 33175 3650
rect 33239 3586 33240 3650
rect 33174 3570 33240 3586
rect 33174 3506 33175 3570
rect 33239 3506 33240 3570
rect 33174 3490 33240 3506
rect 33174 3426 33175 3490
rect 33239 3426 33240 3490
rect 33174 3410 33240 3426
rect 33174 3346 33175 3410
rect 33239 3346 33240 3410
rect 33174 3330 33240 3346
rect 33174 3266 33175 3330
rect 33239 3266 33240 3330
rect 33174 3250 33240 3266
rect 33174 3186 33175 3250
rect 33239 3186 33240 3250
rect 33174 3032 33240 3186
rect 13782 3030 33240 3032
rect 13782 2966 13886 3030
rect 13950 2966 13966 3030
rect 14030 2966 14046 3030
rect 14110 2966 14126 3030
rect 14190 2966 14206 3030
rect 14270 2966 14286 3030
rect 14350 2966 14492 3030
rect 14556 2966 14572 3030
rect 14636 2966 14652 3030
rect 14716 2966 14732 3030
rect 14796 2966 14812 3030
rect 14876 2966 14892 3030
rect 14956 2966 15098 3030
rect 15162 2966 15178 3030
rect 15242 2966 15258 3030
rect 15322 2966 15338 3030
rect 15402 2966 15418 3030
rect 15482 2966 15498 3030
rect 15562 2966 15704 3030
rect 15768 2966 15784 3030
rect 15848 2966 15864 3030
rect 15928 2966 15944 3030
rect 16008 2966 16024 3030
rect 16088 2966 16104 3030
rect 16168 2966 16310 3030
rect 16374 2966 16390 3030
rect 16454 2966 16470 3030
rect 16534 2966 16550 3030
rect 16614 2966 16630 3030
rect 16694 2966 16710 3030
rect 16774 2966 16916 3030
rect 16980 2966 16996 3030
rect 17060 2966 17076 3030
rect 17140 2966 17156 3030
rect 17220 2966 17236 3030
rect 17300 2966 17316 3030
rect 17380 2966 17522 3030
rect 17586 2966 17602 3030
rect 17666 2966 17682 3030
rect 17746 2966 17762 3030
rect 17826 2966 17842 3030
rect 17906 2966 17922 3030
rect 17986 2966 18128 3030
rect 18192 2966 18208 3030
rect 18272 2966 18288 3030
rect 18352 2966 18368 3030
rect 18432 2966 18448 3030
rect 18512 2966 18528 3030
rect 18592 2966 18734 3030
rect 18798 2966 18814 3030
rect 18878 2966 18894 3030
rect 18958 2966 18974 3030
rect 19038 2966 19054 3030
rect 19118 2966 19134 3030
rect 19198 2966 19340 3030
rect 19404 2966 19420 3030
rect 19484 2966 19500 3030
rect 19564 2966 19580 3030
rect 19644 2966 19660 3030
rect 19724 2966 19740 3030
rect 19804 2966 19946 3030
rect 20010 2966 20026 3030
rect 20090 2966 20106 3030
rect 20170 2966 20186 3030
rect 20250 2966 20266 3030
rect 20330 2966 20346 3030
rect 20410 2966 20552 3030
rect 20616 2966 20632 3030
rect 20696 2966 20712 3030
rect 20776 2966 20792 3030
rect 20856 2966 20872 3030
rect 20936 2966 20952 3030
rect 21016 2966 21158 3030
rect 21222 2966 21238 3030
rect 21302 2966 21318 3030
rect 21382 2966 21398 3030
rect 21462 2966 21478 3030
rect 21542 2966 21558 3030
rect 21622 2966 21764 3030
rect 21828 2966 21844 3030
rect 21908 2966 21924 3030
rect 21988 2966 22004 3030
rect 22068 2966 22084 3030
rect 22148 2966 22164 3030
rect 22228 2966 22370 3030
rect 22434 2966 22450 3030
rect 22514 2966 22530 3030
rect 22594 2966 22610 3030
rect 22674 2966 22690 3030
rect 22754 2966 22770 3030
rect 22834 2966 22976 3030
rect 23040 2966 23056 3030
rect 23120 2966 23136 3030
rect 23200 2966 23216 3030
rect 23280 2966 23296 3030
rect 23360 2966 23376 3030
rect 23440 2966 23582 3030
rect 23646 2966 23662 3030
rect 23726 2966 23742 3030
rect 23806 2966 23822 3030
rect 23886 2966 23902 3030
rect 23966 2966 23982 3030
rect 24046 2966 24188 3030
rect 24252 2966 24268 3030
rect 24332 2966 24348 3030
rect 24412 2966 24428 3030
rect 24492 2966 24508 3030
rect 24572 2966 24588 3030
rect 24652 2966 24794 3030
rect 24858 2966 24874 3030
rect 24938 2966 24954 3030
rect 25018 2966 25034 3030
rect 25098 2966 25114 3030
rect 25178 2966 25194 3030
rect 25258 2966 25400 3030
rect 25464 2966 25480 3030
rect 25544 2966 25560 3030
rect 25624 2966 25640 3030
rect 25704 2966 25720 3030
rect 25784 2966 25800 3030
rect 25864 2966 26006 3030
rect 26070 2966 26086 3030
rect 26150 2966 26166 3030
rect 26230 2966 26246 3030
rect 26310 2966 26326 3030
rect 26390 2966 26406 3030
rect 26470 2966 26612 3030
rect 26676 2966 26692 3030
rect 26756 2966 26772 3030
rect 26836 2966 26852 3030
rect 26916 2966 26932 3030
rect 26996 2966 27012 3030
rect 27076 2966 27218 3030
rect 27282 2966 27298 3030
rect 27362 2966 27378 3030
rect 27442 2966 27458 3030
rect 27522 2966 27538 3030
rect 27602 2966 27618 3030
rect 27682 2966 27824 3030
rect 27888 2966 27904 3030
rect 27968 2966 27984 3030
rect 28048 2966 28064 3030
rect 28128 2966 28144 3030
rect 28208 2966 28224 3030
rect 28288 2966 28430 3030
rect 28494 2966 28510 3030
rect 28574 2966 28590 3030
rect 28654 2966 28670 3030
rect 28734 2966 28750 3030
rect 28814 2966 28830 3030
rect 28894 2966 29036 3030
rect 29100 2966 29116 3030
rect 29180 2966 29196 3030
rect 29260 2966 29276 3030
rect 29340 2966 29356 3030
rect 29420 2966 29436 3030
rect 29500 2966 29642 3030
rect 29706 2966 29722 3030
rect 29786 2966 29802 3030
rect 29866 2966 29882 3030
rect 29946 2966 29962 3030
rect 30026 2966 30042 3030
rect 30106 2966 30248 3030
rect 30312 2966 30328 3030
rect 30392 2966 30408 3030
rect 30472 2966 30488 3030
rect 30552 2966 30568 3030
rect 30632 2966 30648 3030
rect 30712 2966 30854 3030
rect 30918 2966 30934 3030
rect 30998 2966 31014 3030
rect 31078 2966 31094 3030
rect 31158 2966 31174 3030
rect 31238 2966 31254 3030
rect 31318 2966 31460 3030
rect 31524 2966 31540 3030
rect 31604 2966 31620 3030
rect 31684 2966 31700 3030
rect 31764 2966 31780 3030
rect 31844 2966 31860 3030
rect 31924 2966 32066 3030
rect 32130 2966 32146 3030
rect 32210 2966 32226 3030
rect 32290 2966 32306 3030
rect 32370 2966 32386 3030
rect 32450 2966 32466 3030
rect 32530 2966 32672 3030
rect 32736 2966 32752 3030
rect 32816 2966 32832 3030
rect 32896 2966 32912 3030
rect 32976 2966 32992 3030
rect 33056 2966 33072 3030
rect 33136 2966 33240 3030
rect 13782 2964 33240 2966
rect 13782 2810 13848 2964
rect 13782 2746 13783 2810
rect 13847 2746 13848 2810
rect 13782 2730 13848 2746
rect 13782 2666 13783 2730
rect 13847 2666 13848 2730
rect 13782 2650 13848 2666
rect 13782 2586 13783 2650
rect 13847 2586 13848 2650
rect 13782 2570 13848 2586
rect 13782 2506 13783 2570
rect 13847 2506 13848 2570
rect 13782 2490 13848 2506
rect 13782 2426 13783 2490
rect 13847 2426 13848 2490
rect 13782 2410 13848 2426
rect 13782 2346 13783 2410
rect 13847 2346 13848 2410
rect 13782 2330 13848 2346
rect 13782 2266 13783 2330
rect 13847 2266 13848 2330
rect 13782 2250 13848 2266
rect 13782 2186 13783 2250
rect 13847 2186 13848 2250
rect 13782 2170 13848 2186
rect 13782 2106 13783 2170
rect 13847 2106 13848 2170
rect 13782 2090 13848 2106
rect 13782 2026 13783 2090
rect 13847 2026 13848 2090
rect 13782 1936 13848 2026
rect 13908 1872 13968 2902
rect 14028 1932 14088 2964
rect 14148 1872 14208 2902
rect 14268 1932 14328 2964
rect 14388 2810 14454 2964
rect 14388 2746 14389 2810
rect 14453 2746 14454 2810
rect 14388 2730 14454 2746
rect 14388 2666 14389 2730
rect 14453 2666 14454 2730
rect 14388 2650 14454 2666
rect 14388 2586 14389 2650
rect 14453 2586 14454 2650
rect 14388 2570 14454 2586
rect 14388 2506 14389 2570
rect 14453 2506 14454 2570
rect 14388 2490 14454 2506
rect 14388 2426 14389 2490
rect 14453 2426 14454 2490
rect 14388 2410 14454 2426
rect 14388 2346 14389 2410
rect 14453 2346 14454 2410
rect 14388 2330 14454 2346
rect 14388 2266 14389 2330
rect 14453 2266 14454 2330
rect 14388 2250 14454 2266
rect 14388 2186 14389 2250
rect 14453 2186 14454 2250
rect 14388 2170 14454 2186
rect 14388 2106 14389 2170
rect 14453 2106 14454 2170
rect 14388 2090 14454 2106
rect 14388 2026 14389 2090
rect 14453 2026 14454 2090
rect 14388 1936 14454 2026
rect 14514 1872 14574 2902
rect 14634 1932 14694 2964
rect 14754 1872 14814 2902
rect 14874 1932 14934 2964
rect 14994 2810 15060 2964
rect 14994 2746 14995 2810
rect 15059 2746 15060 2810
rect 14994 2730 15060 2746
rect 14994 2666 14995 2730
rect 15059 2666 15060 2730
rect 14994 2650 15060 2666
rect 14994 2586 14995 2650
rect 15059 2586 15060 2650
rect 14994 2570 15060 2586
rect 14994 2506 14995 2570
rect 15059 2506 15060 2570
rect 14994 2490 15060 2506
rect 14994 2426 14995 2490
rect 15059 2426 15060 2490
rect 14994 2410 15060 2426
rect 14994 2346 14995 2410
rect 15059 2346 15060 2410
rect 14994 2330 15060 2346
rect 14994 2266 14995 2330
rect 15059 2266 15060 2330
rect 14994 2250 15060 2266
rect 14994 2186 14995 2250
rect 15059 2186 15060 2250
rect 14994 2170 15060 2186
rect 14994 2106 14995 2170
rect 15059 2106 15060 2170
rect 14994 2090 15060 2106
rect 14994 2026 14995 2090
rect 15059 2026 15060 2090
rect 14994 1936 15060 2026
rect 15120 1872 15180 2902
rect 15240 1932 15300 2964
rect 15360 1872 15420 2902
rect 15480 1932 15540 2964
rect 15600 2810 15666 2964
rect 15600 2746 15601 2810
rect 15665 2746 15666 2810
rect 15600 2730 15666 2746
rect 15600 2666 15601 2730
rect 15665 2666 15666 2730
rect 15600 2650 15666 2666
rect 15600 2586 15601 2650
rect 15665 2586 15666 2650
rect 15600 2570 15666 2586
rect 15600 2506 15601 2570
rect 15665 2506 15666 2570
rect 15600 2490 15666 2506
rect 15600 2426 15601 2490
rect 15665 2426 15666 2490
rect 15600 2410 15666 2426
rect 15600 2346 15601 2410
rect 15665 2346 15666 2410
rect 15600 2330 15666 2346
rect 15600 2266 15601 2330
rect 15665 2266 15666 2330
rect 15600 2250 15666 2266
rect 15600 2186 15601 2250
rect 15665 2186 15666 2250
rect 15600 2170 15666 2186
rect 15600 2106 15601 2170
rect 15665 2106 15666 2170
rect 15600 2090 15666 2106
rect 15600 2026 15601 2090
rect 15665 2026 15666 2090
rect 15600 1936 15666 2026
rect 15726 1872 15786 2902
rect 15846 1932 15906 2964
rect 15966 1872 16026 2902
rect 16086 1932 16146 2964
rect 16206 2810 16272 2964
rect 16206 2746 16207 2810
rect 16271 2746 16272 2810
rect 16206 2730 16272 2746
rect 16206 2666 16207 2730
rect 16271 2666 16272 2730
rect 16206 2650 16272 2666
rect 16206 2586 16207 2650
rect 16271 2586 16272 2650
rect 16206 2570 16272 2586
rect 16206 2506 16207 2570
rect 16271 2506 16272 2570
rect 16206 2490 16272 2506
rect 16206 2426 16207 2490
rect 16271 2426 16272 2490
rect 16206 2410 16272 2426
rect 16206 2346 16207 2410
rect 16271 2346 16272 2410
rect 16206 2330 16272 2346
rect 16206 2266 16207 2330
rect 16271 2266 16272 2330
rect 16206 2250 16272 2266
rect 16206 2186 16207 2250
rect 16271 2186 16272 2250
rect 16206 2170 16272 2186
rect 16206 2106 16207 2170
rect 16271 2106 16272 2170
rect 16206 2090 16272 2106
rect 16206 2026 16207 2090
rect 16271 2026 16272 2090
rect 16206 1936 16272 2026
rect 16332 1872 16392 2902
rect 16452 1932 16512 2964
rect 16572 1872 16632 2902
rect 16692 1932 16752 2964
rect 16812 2810 16878 2964
rect 16812 2746 16813 2810
rect 16877 2746 16878 2810
rect 16812 2730 16878 2746
rect 16812 2666 16813 2730
rect 16877 2666 16878 2730
rect 16812 2650 16878 2666
rect 16812 2586 16813 2650
rect 16877 2586 16878 2650
rect 16812 2570 16878 2586
rect 16812 2506 16813 2570
rect 16877 2506 16878 2570
rect 16812 2490 16878 2506
rect 16812 2426 16813 2490
rect 16877 2426 16878 2490
rect 16812 2410 16878 2426
rect 16812 2346 16813 2410
rect 16877 2346 16878 2410
rect 16812 2330 16878 2346
rect 16812 2266 16813 2330
rect 16877 2266 16878 2330
rect 16812 2250 16878 2266
rect 16812 2186 16813 2250
rect 16877 2186 16878 2250
rect 16812 2170 16878 2186
rect 16812 2106 16813 2170
rect 16877 2106 16878 2170
rect 16812 2090 16878 2106
rect 16812 2026 16813 2090
rect 16877 2026 16878 2090
rect 16812 1936 16878 2026
rect 16938 1872 16998 2902
rect 17058 1932 17118 2964
rect 17178 1872 17238 2902
rect 17298 1932 17358 2964
rect 17418 2810 17484 2964
rect 17418 2746 17419 2810
rect 17483 2746 17484 2810
rect 17418 2730 17484 2746
rect 17418 2666 17419 2730
rect 17483 2666 17484 2730
rect 17418 2650 17484 2666
rect 17418 2586 17419 2650
rect 17483 2586 17484 2650
rect 17418 2570 17484 2586
rect 17418 2506 17419 2570
rect 17483 2506 17484 2570
rect 17418 2490 17484 2506
rect 17418 2426 17419 2490
rect 17483 2426 17484 2490
rect 17418 2410 17484 2426
rect 17418 2346 17419 2410
rect 17483 2346 17484 2410
rect 17418 2330 17484 2346
rect 17418 2266 17419 2330
rect 17483 2266 17484 2330
rect 17418 2250 17484 2266
rect 17418 2186 17419 2250
rect 17483 2186 17484 2250
rect 17418 2170 17484 2186
rect 17418 2106 17419 2170
rect 17483 2106 17484 2170
rect 17418 2090 17484 2106
rect 17418 2026 17419 2090
rect 17483 2026 17484 2090
rect 17418 1936 17484 2026
rect 17544 1872 17604 2902
rect 17664 1932 17724 2964
rect 17784 1872 17844 2902
rect 17904 1932 17964 2964
rect 18024 2810 18090 2964
rect 18024 2746 18025 2810
rect 18089 2746 18090 2810
rect 18024 2730 18090 2746
rect 18024 2666 18025 2730
rect 18089 2666 18090 2730
rect 18024 2650 18090 2666
rect 18024 2586 18025 2650
rect 18089 2586 18090 2650
rect 18024 2570 18090 2586
rect 18024 2506 18025 2570
rect 18089 2506 18090 2570
rect 18024 2490 18090 2506
rect 18024 2426 18025 2490
rect 18089 2426 18090 2490
rect 18024 2410 18090 2426
rect 18024 2346 18025 2410
rect 18089 2346 18090 2410
rect 18024 2330 18090 2346
rect 18024 2266 18025 2330
rect 18089 2266 18090 2330
rect 18024 2250 18090 2266
rect 18024 2186 18025 2250
rect 18089 2186 18090 2250
rect 18024 2170 18090 2186
rect 18024 2106 18025 2170
rect 18089 2106 18090 2170
rect 18024 2090 18090 2106
rect 18024 2026 18025 2090
rect 18089 2026 18090 2090
rect 18024 1936 18090 2026
rect 18150 1872 18210 2902
rect 18270 1932 18330 2964
rect 18390 1872 18450 2902
rect 18510 1932 18570 2964
rect 18630 2810 18696 2964
rect 18630 2746 18631 2810
rect 18695 2746 18696 2810
rect 18630 2730 18696 2746
rect 18630 2666 18631 2730
rect 18695 2666 18696 2730
rect 18630 2650 18696 2666
rect 18630 2586 18631 2650
rect 18695 2586 18696 2650
rect 18630 2570 18696 2586
rect 18630 2506 18631 2570
rect 18695 2506 18696 2570
rect 18630 2490 18696 2506
rect 18630 2426 18631 2490
rect 18695 2426 18696 2490
rect 18630 2410 18696 2426
rect 18630 2346 18631 2410
rect 18695 2346 18696 2410
rect 18630 2330 18696 2346
rect 18630 2266 18631 2330
rect 18695 2266 18696 2330
rect 18630 2250 18696 2266
rect 18630 2186 18631 2250
rect 18695 2186 18696 2250
rect 18630 2170 18696 2186
rect 18630 2106 18631 2170
rect 18695 2106 18696 2170
rect 18630 2090 18696 2106
rect 18630 2026 18631 2090
rect 18695 2026 18696 2090
rect 18630 1936 18696 2026
rect 18756 1872 18816 2902
rect 18876 1932 18936 2964
rect 18996 1872 19056 2902
rect 19116 1932 19176 2964
rect 19236 2810 19302 2964
rect 19236 2746 19237 2810
rect 19301 2746 19302 2810
rect 19236 2730 19302 2746
rect 19236 2666 19237 2730
rect 19301 2666 19302 2730
rect 19236 2650 19302 2666
rect 19236 2586 19237 2650
rect 19301 2586 19302 2650
rect 19236 2570 19302 2586
rect 19236 2506 19237 2570
rect 19301 2506 19302 2570
rect 19236 2490 19302 2506
rect 19236 2426 19237 2490
rect 19301 2426 19302 2490
rect 19236 2410 19302 2426
rect 19236 2346 19237 2410
rect 19301 2346 19302 2410
rect 19236 2330 19302 2346
rect 19236 2266 19237 2330
rect 19301 2266 19302 2330
rect 19236 2250 19302 2266
rect 19236 2186 19237 2250
rect 19301 2186 19302 2250
rect 19236 2170 19302 2186
rect 19236 2106 19237 2170
rect 19301 2106 19302 2170
rect 19236 2090 19302 2106
rect 19236 2026 19237 2090
rect 19301 2026 19302 2090
rect 19236 1936 19302 2026
rect 19362 1872 19422 2902
rect 19482 1932 19542 2964
rect 19602 1872 19662 2902
rect 19722 1932 19782 2964
rect 19842 2810 19908 2964
rect 19842 2746 19843 2810
rect 19907 2746 19908 2810
rect 19842 2730 19908 2746
rect 19842 2666 19843 2730
rect 19907 2666 19908 2730
rect 19842 2650 19908 2666
rect 19842 2586 19843 2650
rect 19907 2586 19908 2650
rect 19842 2570 19908 2586
rect 19842 2506 19843 2570
rect 19907 2506 19908 2570
rect 19842 2490 19908 2506
rect 19842 2426 19843 2490
rect 19907 2426 19908 2490
rect 19842 2410 19908 2426
rect 19842 2346 19843 2410
rect 19907 2346 19908 2410
rect 19842 2330 19908 2346
rect 19842 2266 19843 2330
rect 19907 2266 19908 2330
rect 19842 2250 19908 2266
rect 19842 2186 19843 2250
rect 19907 2186 19908 2250
rect 19842 2170 19908 2186
rect 19842 2106 19843 2170
rect 19907 2106 19908 2170
rect 19842 2090 19908 2106
rect 19842 2026 19843 2090
rect 19907 2026 19908 2090
rect 19842 1936 19908 2026
rect 19968 1872 20028 2902
rect 20088 1932 20148 2964
rect 20208 1872 20268 2902
rect 20328 1932 20388 2964
rect 20448 2810 20514 2964
rect 20448 2746 20449 2810
rect 20513 2746 20514 2810
rect 20448 2730 20514 2746
rect 20448 2666 20449 2730
rect 20513 2666 20514 2730
rect 20448 2650 20514 2666
rect 20448 2586 20449 2650
rect 20513 2586 20514 2650
rect 20448 2570 20514 2586
rect 20448 2506 20449 2570
rect 20513 2506 20514 2570
rect 20448 2490 20514 2506
rect 20448 2426 20449 2490
rect 20513 2426 20514 2490
rect 20448 2410 20514 2426
rect 20448 2346 20449 2410
rect 20513 2346 20514 2410
rect 20448 2330 20514 2346
rect 20448 2266 20449 2330
rect 20513 2266 20514 2330
rect 20448 2250 20514 2266
rect 20448 2186 20449 2250
rect 20513 2186 20514 2250
rect 20448 2170 20514 2186
rect 20448 2106 20449 2170
rect 20513 2106 20514 2170
rect 20448 2090 20514 2106
rect 20448 2026 20449 2090
rect 20513 2026 20514 2090
rect 20448 1936 20514 2026
rect 20574 1872 20634 2902
rect 20694 1932 20754 2964
rect 20814 1872 20874 2902
rect 20934 1932 20994 2964
rect 21054 2810 21120 2964
rect 21054 2746 21055 2810
rect 21119 2746 21120 2810
rect 21054 2730 21120 2746
rect 21054 2666 21055 2730
rect 21119 2666 21120 2730
rect 21054 2650 21120 2666
rect 21054 2586 21055 2650
rect 21119 2586 21120 2650
rect 21054 2570 21120 2586
rect 21054 2506 21055 2570
rect 21119 2506 21120 2570
rect 21054 2490 21120 2506
rect 21054 2426 21055 2490
rect 21119 2426 21120 2490
rect 21054 2410 21120 2426
rect 21054 2346 21055 2410
rect 21119 2346 21120 2410
rect 21054 2330 21120 2346
rect 21054 2266 21055 2330
rect 21119 2266 21120 2330
rect 21054 2250 21120 2266
rect 21054 2186 21055 2250
rect 21119 2186 21120 2250
rect 21054 2170 21120 2186
rect 21054 2106 21055 2170
rect 21119 2106 21120 2170
rect 21054 2090 21120 2106
rect 21054 2026 21055 2090
rect 21119 2026 21120 2090
rect 21054 1936 21120 2026
rect 21180 1872 21240 2902
rect 21300 1932 21360 2964
rect 21420 1872 21480 2902
rect 21540 1932 21600 2964
rect 21660 2810 21726 2964
rect 21660 2746 21661 2810
rect 21725 2746 21726 2810
rect 21660 2730 21726 2746
rect 21660 2666 21661 2730
rect 21725 2666 21726 2730
rect 21660 2650 21726 2666
rect 21660 2586 21661 2650
rect 21725 2586 21726 2650
rect 21660 2570 21726 2586
rect 21660 2506 21661 2570
rect 21725 2506 21726 2570
rect 21660 2490 21726 2506
rect 21660 2426 21661 2490
rect 21725 2426 21726 2490
rect 21660 2410 21726 2426
rect 21660 2346 21661 2410
rect 21725 2346 21726 2410
rect 21660 2330 21726 2346
rect 21660 2266 21661 2330
rect 21725 2266 21726 2330
rect 21660 2250 21726 2266
rect 21660 2186 21661 2250
rect 21725 2186 21726 2250
rect 21660 2170 21726 2186
rect 21660 2106 21661 2170
rect 21725 2106 21726 2170
rect 21660 2090 21726 2106
rect 21660 2026 21661 2090
rect 21725 2026 21726 2090
rect 21660 1936 21726 2026
rect 21786 1872 21846 2902
rect 21906 1932 21966 2964
rect 22026 1872 22086 2902
rect 22146 1932 22206 2964
rect 22266 2810 22332 2964
rect 22266 2746 22267 2810
rect 22331 2746 22332 2810
rect 22266 2730 22332 2746
rect 22266 2666 22267 2730
rect 22331 2666 22332 2730
rect 22266 2650 22332 2666
rect 22266 2586 22267 2650
rect 22331 2586 22332 2650
rect 22266 2570 22332 2586
rect 22266 2506 22267 2570
rect 22331 2506 22332 2570
rect 22266 2490 22332 2506
rect 22266 2426 22267 2490
rect 22331 2426 22332 2490
rect 22266 2410 22332 2426
rect 22266 2346 22267 2410
rect 22331 2346 22332 2410
rect 22266 2330 22332 2346
rect 22266 2266 22267 2330
rect 22331 2266 22332 2330
rect 22266 2250 22332 2266
rect 22266 2186 22267 2250
rect 22331 2186 22332 2250
rect 22266 2170 22332 2186
rect 22266 2106 22267 2170
rect 22331 2106 22332 2170
rect 22266 2090 22332 2106
rect 22266 2026 22267 2090
rect 22331 2026 22332 2090
rect 22266 1936 22332 2026
rect 22392 1872 22452 2902
rect 22512 1932 22572 2964
rect 22632 1872 22692 2902
rect 22752 1932 22812 2964
rect 22872 2810 22938 2964
rect 22872 2746 22873 2810
rect 22937 2746 22938 2810
rect 22872 2730 22938 2746
rect 22872 2666 22873 2730
rect 22937 2666 22938 2730
rect 22872 2650 22938 2666
rect 22872 2586 22873 2650
rect 22937 2586 22938 2650
rect 22872 2570 22938 2586
rect 22872 2506 22873 2570
rect 22937 2506 22938 2570
rect 22872 2490 22938 2506
rect 22872 2426 22873 2490
rect 22937 2426 22938 2490
rect 22872 2410 22938 2426
rect 22872 2346 22873 2410
rect 22937 2346 22938 2410
rect 22872 2330 22938 2346
rect 22872 2266 22873 2330
rect 22937 2266 22938 2330
rect 22872 2250 22938 2266
rect 22872 2186 22873 2250
rect 22937 2186 22938 2250
rect 22872 2170 22938 2186
rect 22872 2106 22873 2170
rect 22937 2106 22938 2170
rect 22872 2090 22938 2106
rect 22872 2026 22873 2090
rect 22937 2026 22938 2090
rect 22872 1936 22938 2026
rect 22998 1872 23058 2902
rect 23118 1932 23178 2964
rect 23238 1872 23298 2902
rect 23358 1932 23418 2964
rect 23478 2810 23544 2964
rect 23478 2746 23479 2810
rect 23543 2746 23544 2810
rect 23478 2730 23544 2746
rect 23478 2666 23479 2730
rect 23543 2666 23544 2730
rect 23478 2650 23544 2666
rect 23478 2586 23479 2650
rect 23543 2586 23544 2650
rect 23478 2570 23544 2586
rect 23478 2506 23479 2570
rect 23543 2506 23544 2570
rect 23478 2490 23544 2506
rect 23478 2426 23479 2490
rect 23543 2426 23544 2490
rect 23478 2410 23544 2426
rect 23478 2346 23479 2410
rect 23543 2346 23544 2410
rect 23478 2330 23544 2346
rect 23478 2266 23479 2330
rect 23543 2266 23544 2330
rect 23478 2250 23544 2266
rect 23478 2186 23479 2250
rect 23543 2186 23544 2250
rect 23478 2170 23544 2186
rect 23478 2106 23479 2170
rect 23543 2106 23544 2170
rect 23478 2090 23544 2106
rect 23478 2026 23479 2090
rect 23543 2026 23544 2090
rect 23478 1936 23544 2026
rect 23604 1872 23664 2902
rect 23724 1932 23784 2964
rect 23844 1872 23904 2902
rect 23964 1932 24024 2964
rect 24084 2810 24150 2964
rect 24084 2746 24085 2810
rect 24149 2746 24150 2810
rect 24084 2730 24150 2746
rect 24084 2666 24085 2730
rect 24149 2666 24150 2730
rect 24084 2650 24150 2666
rect 24084 2586 24085 2650
rect 24149 2586 24150 2650
rect 24084 2570 24150 2586
rect 24084 2506 24085 2570
rect 24149 2506 24150 2570
rect 24084 2490 24150 2506
rect 24084 2426 24085 2490
rect 24149 2426 24150 2490
rect 24084 2410 24150 2426
rect 24084 2346 24085 2410
rect 24149 2346 24150 2410
rect 24084 2330 24150 2346
rect 24084 2266 24085 2330
rect 24149 2266 24150 2330
rect 24084 2250 24150 2266
rect 24084 2186 24085 2250
rect 24149 2186 24150 2250
rect 24084 2170 24150 2186
rect 24084 2106 24085 2170
rect 24149 2106 24150 2170
rect 24084 2090 24150 2106
rect 24084 2026 24085 2090
rect 24149 2026 24150 2090
rect 24084 1936 24150 2026
rect 24210 1872 24270 2902
rect 24330 1932 24390 2964
rect 24450 1872 24510 2902
rect 24570 1932 24630 2964
rect 24690 2810 24756 2964
rect 24690 2746 24691 2810
rect 24755 2746 24756 2810
rect 24690 2730 24756 2746
rect 24690 2666 24691 2730
rect 24755 2666 24756 2730
rect 24690 2650 24756 2666
rect 24690 2586 24691 2650
rect 24755 2586 24756 2650
rect 24690 2570 24756 2586
rect 24690 2506 24691 2570
rect 24755 2506 24756 2570
rect 24690 2490 24756 2506
rect 24690 2426 24691 2490
rect 24755 2426 24756 2490
rect 24690 2410 24756 2426
rect 24690 2346 24691 2410
rect 24755 2346 24756 2410
rect 24690 2330 24756 2346
rect 24690 2266 24691 2330
rect 24755 2266 24756 2330
rect 24690 2250 24756 2266
rect 24690 2186 24691 2250
rect 24755 2186 24756 2250
rect 24690 2170 24756 2186
rect 24690 2106 24691 2170
rect 24755 2106 24756 2170
rect 24690 2090 24756 2106
rect 24690 2026 24691 2090
rect 24755 2026 24756 2090
rect 24690 1936 24756 2026
rect 24816 1872 24876 2902
rect 24936 1932 24996 2964
rect 25056 1872 25116 2902
rect 25176 1932 25236 2964
rect 25296 2810 25362 2964
rect 25296 2746 25297 2810
rect 25361 2746 25362 2810
rect 25296 2730 25362 2746
rect 25296 2666 25297 2730
rect 25361 2666 25362 2730
rect 25296 2650 25362 2666
rect 25296 2586 25297 2650
rect 25361 2586 25362 2650
rect 25296 2570 25362 2586
rect 25296 2506 25297 2570
rect 25361 2506 25362 2570
rect 25296 2490 25362 2506
rect 25296 2426 25297 2490
rect 25361 2426 25362 2490
rect 25296 2410 25362 2426
rect 25296 2346 25297 2410
rect 25361 2346 25362 2410
rect 25296 2330 25362 2346
rect 25296 2266 25297 2330
rect 25361 2266 25362 2330
rect 25296 2250 25362 2266
rect 25296 2186 25297 2250
rect 25361 2186 25362 2250
rect 25296 2170 25362 2186
rect 25296 2106 25297 2170
rect 25361 2106 25362 2170
rect 25296 2090 25362 2106
rect 25296 2026 25297 2090
rect 25361 2026 25362 2090
rect 25296 1936 25362 2026
rect 25422 1872 25482 2902
rect 25542 1932 25602 2964
rect 25662 1872 25722 2902
rect 25782 1932 25842 2964
rect 25902 2810 25968 2964
rect 25902 2746 25903 2810
rect 25967 2746 25968 2810
rect 25902 2730 25968 2746
rect 25902 2666 25903 2730
rect 25967 2666 25968 2730
rect 25902 2650 25968 2666
rect 25902 2586 25903 2650
rect 25967 2586 25968 2650
rect 25902 2570 25968 2586
rect 25902 2506 25903 2570
rect 25967 2506 25968 2570
rect 25902 2490 25968 2506
rect 25902 2426 25903 2490
rect 25967 2426 25968 2490
rect 25902 2410 25968 2426
rect 25902 2346 25903 2410
rect 25967 2346 25968 2410
rect 25902 2330 25968 2346
rect 25902 2266 25903 2330
rect 25967 2266 25968 2330
rect 25902 2250 25968 2266
rect 25902 2186 25903 2250
rect 25967 2186 25968 2250
rect 25902 2170 25968 2186
rect 25902 2106 25903 2170
rect 25967 2106 25968 2170
rect 25902 2090 25968 2106
rect 25902 2026 25903 2090
rect 25967 2026 25968 2090
rect 25902 1936 25968 2026
rect 26028 1872 26088 2902
rect 26148 1932 26208 2964
rect 26268 1872 26328 2902
rect 26388 1932 26448 2964
rect 26508 2810 26574 2964
rect 26508 2746 26509 2810
rect 26573 2746 26574 2810
rect 26508 2730 26574 2746
rect 26508 2666 26509 2730
rect 26573 2666 26574 2730
rect 26508 2650 26574 2666
rect 26508 2586 26509 2650
rect 26573 2586 26574 2650
rect 26508 2570 26574 2586
rect 26508 2506 26509 2570
rect 26573 2506 26574 2570
rect 26508 2490 26574 2506
rect 26508 2426 26509 2490
rect 26573 2426 26574 2490
rect 26508 2410 26574 2426
rect 26508 2346 26509 2410
rect 26573 2346 26574 2410
rect 26508 2330 26574 2346
rect 26508 2266 26509 2330
rect 26573 2266 26574 2330
rect 26508 2250 26574 2266
rect 26508 2186 26509 2250
rect 26573 2186 26574 2250
rect 26508 2170 26574 2186
rect 26508 2106 26509 2170
rect 26573 2106 26574 2170
rect 26508 2090 26574 2106
rect 26508 2026 26509 2090
rect 26573 2026 26574 2090
rect 26508 1936 26574 2026
rect 26634 1872 26694 2902
rect 26754 1932 26814 2964
rect 26874 1872 26934 2902
rect 26994 1932 27054 2964
rect 27114 2810 27180 2964
rect 27114 2746 27115 2810
rect 27179 2746 27180 2810
rect 27114 2730 27180 2746
rect 27114 2666 27115 2730
rect 27179 2666 27180 2730
rect 27114 2650 27180 2666
rect 27114 2586 27115 2650
rect 27179 2586 27180 2650
rect 27114 2570 27180 2586
rect 27114 2506 27115 2570
rect 27179 2506 27180 2570
rect 27114 2490 27180 2506
rect 27114 2426 27115 2490
rect 27179 2426 27180 2490
rect 27114 2410 27180 2426
rect 27114 2346 27115 2410
rect 27179 2346 27180 2410
rect 27114 2330 27180 2346
rect 27114 2266 27115 2330
rect 27179 2266 27180 2330
rect 27114 2250 27180 2266
rect 27114 2186 27115 2250
rect 27179 2186 27180 2250
rect 27114 2170 27180 2186
rect 27114 2106 27115 2170
rect 27179 2106 27180 2170
rect 27114 2090 27180 2106
rect 27114 2026 27115 2090
rect 27179 2026 27180 2090
rect 27114 1936 27180 2026
rect 27240 1872 27300 2902
rect 27360 1932 27420 2964
rect 27480 1872 27540 2902
rect 27600 1932 27660 2964
rect 27720 2810 27786 2964
rect 27720 2746 27721 2810
rect 27785 2746 27786 2810
rect 27720 2730 27786 2746
rect 27720 2666 27721 2730
rect 27785 2666 27786 2730
rect 27720 2650 27786 2666
rect 27720 2586 27721 2650
rect 27785 2586 27786 2650
rect 27720 2570 27786 2586
rect 27720 2506 27721 2570
rect 27785 2506 27786 2570
rect 27720 2490 27786 2506
rect 27720 2426 27721 2490
rect 27785 2426 27786 2490
rect 27720 2410 27786 2426
rect 27720 2346 27721 2410
rect 27785 2346 27786 2410
rect 27720 2330 27786 2346
rect 27720 2266 27721 2330
rect 27785 2266 27786 2330
rect 27720 2250 27786 2266
rect 27720 2186 27721 2250
rect 27785 2186 27786 2250
rect 27720 2170 27786 2186
rect 27720 2106 27721 2170
rect 27785 2106 27786 2170
rect 27720 2090 27786 2106
rect 27720 2026 27721 2090
rect 27785 2026 27786 2090
rect 27720 1936 27786 2026
rect 27846 1872 27906 2902
rect 27966 1932 28026 2964
rect 28086 1872 28146 2902
rect 28206 1932 28266 2964
rect 28326 2810 28392 2964
rect 28326 2746 28327 2810
rect 28391 2746 28392 2810
rect 28326 2730 28392 2746
rect 28326 2666 28327 2730
rect 28391 2666 28392 2730
rect 28326 2650 28392 2666
rect 28326 2586 28327 2650
rect 28391 2586 28392 2650
rect 28326 2570 28392 2586
rect 28326 2506 28327 2570
rect 28391 2506 28392 2570
rect 28326 2490 28392 2506
rect 28326 2426 28327 2490
rect 28391 2426 28392 2490
rect 28326 2410 28392 2426
rect 28326 2346 28327 2410
rect 28391 2346 28392 2410
rect 28326 2330 28392 2346
rect 28326 2266 28327 2330
rect 28391 2266 28392 2330
rect 28326 2250 28392 2266
rect 28326 2186 28327 2250
rect 28391 2186 28392 2250
rect 28326 2170 28392 2186
rect 28326 2106 28327 2170
rect 28391 2106 28392 2170
rect 28326 2090 28392 2106
rect 28326 2026 28327 2090
rect 28391 2026 28392 2090
rect 28326 1936 28392 2026
rect 28452 1872 28512 2902
rect 28572 1932 28632 2964
rect 28692 1872 28752 2902
rect 28812 1932 28872 2964
rect 28932 2810 28998 2964
rect 28932 2746 28933 2810
rect 28997 2746 28998 2810
rect 28932 2730 28998 2746
rect 28932 2666 28933 2730
rect 28997 2666 28998 2730
rect 28932 2650 28998 2666
rect 28932 2586 28933 2650
rect 28997 2586 28998 2650
rect 28932 2570 28998 2586
rect 28932 2506 28933 2570
rect 28997 2506 28998 2570
rect 28932 2490 28998 2506
rect 28932 2426 28933 2490
rect 28997 2426 28998 2490
rect 28932 2410 28998 2426
rect 28932 2346 28933 2410
rect 28997 2346 28998 2410
rect 28932 2330 28998 2346
rect 28932 2266 28933 2330
rect 28997 2266 28998 2330
rect 28932 2250 28998 2266
rect 28932 2186 28933 2250
rect 28997 2186 28998 2250
rect 28932 2170 28998 2186
rect 28932 2106 28933 2170
rect 28997 2106 28998 2170
rect 28932 2090 28998 2106
rect 28932 2026 28933 2090
rect 28997 2026 28998 2090
rect 28932 1936 28998 2026
rect 29058 1872 29118 2902
rect 29178 1932 29238 2964
rect 29298 1872 29358 2902
rect 29418 1932 29478 2964
rect 29538 2810 29604 2964
rect 29538 2746 29539 2810
rect 29603 2746 29604 2810
rect 29538 2730 29604 2746
rect 29538 2666 29539 2730
rect 29603 2666 29604 2730
rect 29538 2650 29604 2666
rect 29538 2586 29539 2650
rect 29603 2586 29604 2650
rect 29538 2570 29604 2586
rect 29538 2506 29539 2570
rect 29603 2506 29604 2570
rect 29538 2490 29604 2506
rect 29538 2426 29539 2490
rect 29603 2426 29604 2490
rect 29538 2410 29604 2426
rect 29538 2346 29539 2410
rect 29603 2346 29604 2410
rect 29538 2330 29604 2346
rect 29538 2266 29539 2330
rect 29603 2266 29604 2330
rect 29538 2250 29604 2266
rect 29538 2186 29539 2250
rect 29603 2186 29604 2250
rect 29538 2170 29604 2186
rect 29538 2106 29539 2170
rect 29603 2106 29604 2170
rect 29538 2090 29604 2106
rect 29538 2026 29539 2090
rect 29603 2026 29604 2090
rect 29538 1936 29604 2026
rect 29664 1872 29724 2902
rect 29784 1932 29844 2964
rect 29904 1872 29964 2902
rect 30024 1932 30084 2964
rect 30144 2810 30210 2964
rect 30144 2746 30145 2810
rect 30209 2746 30210 2810
rect 30144 2730 30210 2746
rect 30144 2666 30145 2730
rect 30209 2666 30210 2730
rect 30144 2650 30210 2666
rect 30144 2586 30145 2650
rect 30209 2586 30210 2650
rect 30144 2570 30210 2586
rect 30144 2506 30145 2570
rect 30209 2506 30210 2570
rect 30144 2490 30210 2506
rect 30144 2426 30145 2490
rect 30209 2426 30210 2490
rect 30144 2410 30210 2426
rect 30144 2346 30145 2410
rect 30209 2346 30210 2410
rect 30144 2330 30210 2346
rect 30144 2266 30145 2330
rect 30209 2266 30210 2330
rect 30144 2250 30210 2266
rect 30144 2186 30145 2250
rect 30209 2186 30210 2250
rect 30144 2170 30210 2186
rect 30144 2106 30145 2170
rect 30209 2106 30210 2170
rect 30144 2090 30210 2106
rect 30144 2026 30145 2090
rect 30209 2026 30210 2090
rect 30144 1936 30210 2026
rect 30270 1872 30330 2902
rect 30390 1932 30450 2964
rect 30510 1872 30570 2902
rect 30630 1932 30690 2964
rect 30750 2810 30816 2964
rect 30750 2746 30751 2810
rect 30815 2746 30816 2810
rect 30750 2730 30816 2746
rect 30750 2666 30751 2730
rect 30815 2666 30816 2730
rect 30750 2650 30816 2666
rect 30750 2586 30751 2650
rect 30815 2586 30816 2650
rect 30750 2570 30816 2586
rect 30750 2506 30751 2570
rect 30815 2506 30816 2570
rect 30750 2490 30816 2506
rect 30750 2426 30751 2490
rect 30815 2426 30816 2490
rect 30750 2410 30816 2426
rect 30750 2346 30751 2410
rect 30815 2346 30816 2410
rect 30750 2330 30816 2346
rect 30750 2266 30751 2330
rect 30815 2266 30816 2330
rect 30750 2250 30816 2266
rect 30750 2186 30751 2250
rect 30815 2186 30816 2250
rect 30750 2170 30816 2186
rect 30750 2106 30751 2170
rect 30815 2106 30816 2170
rect 30750 2090 30816 2106
rect 30750 2026 30751 2090
rect 30815 2026 30816 2090
rect 30750 1936 30816 2026
rect 30876 1872 30936 2902
rect 30996 1932 31056 2964
rect 31116 1872 31176 2902
rect 31236 1932 31296 2964
rect 31356 2810 31422 2964
rect 31356 2746 31357 2810
rect 31421 2746 31422 2810
rect 31356 2730 31422 2746
rect 31356 2666 31357 2730
rect 31421 2666 31422 2730
rect 31356 2650 31422 2666
rect 31356 2586 31357 2650
rect 31421 2586 31422 2650
rect 31356 2570 31422 2586
rect 31356 2506 31357 2570
rect 31421 2506 31422 2570
rect 31356 2490 31422 2506
rect 31356 2426 31357 2490
rect 31421 2426 31422 2490
rect 31356 2410 31422 2426
rect 31356 2346 31357 2410
rect 31421 2346 31422 2410
rect 31356 2330 31422 2346
rect 31356 2266 31357 2330
rect 31421 2266 31422 2330
rect 31356 2250 31422 2266
rect 31356 2186 31357 2250
rect 31421 2186 31422 2250
rect 31356 2170 31422 2186
rect 31356 2106 31357 2170
rect 31421 2106 31422 2170
rect 31356 2090 31422 2106
rect 31356 2026 31357 2090
rect 31421 2026 31422 2090
rect 31356 1936 31422 2026
rect 31482 1872 31542 2902
rect 31602 1932 31662 2964
rect 31722 1872 31782 2902
rect 31842 1932 31902 2964
rect 31962 2810 32028 2964
rect 31962 2746 31963 2810
rect 32027 2746 32028 2810
rect 31962 2730 32028 2746
rect 31962 2666 31963 2730
rect 32027 2666 32028 2730
rect 31962 2650 32028 2666
rect 31962 2586 31963 2650
rect 32027 2586 32028 2650
rect 31962 2570 32028 2586
rect 31962 2506 31963 2570
rect 32027 2506 32028 2570
rect 31962 2490 32028 2506
rect 31962 2426 31963 2490
rect 32027 2426 32028 2490
rect 31962 2410 32028 2426
rect 31962 2346 31963 2410
rect 32027 2346 32028 2410
rect 31962 2330 32028 2346
rect 31962 2266 31963 2330
rect 32027 2266 32028 2330
rect 31962 2250 32028 2266
rect 31962 2186 31963 2250
rect 32027 2186 32028 2250
rect 31962 2170 32028 2186
rect 31962 2106 31963 2170
rect 32027 2106 32028 2170
rect 31962 2090 32028 2106
rect 31962 2026 31963 2090
rect 32027 2026 32028 2090
rect 31962 1936 32028 2026
rect 32088 1872 32148 2902
rect 32208 1932 32268 2964
rect 32328 1872 32388 2902
rect 32448 1932 32508 2964
rect 32568 2810 32634 2964
rect 32568 2746 32569 2810
rect 32633 2746 32634 2810
rect 32568 2730 32634 2746
rect 32568 2666 32569 2730
rect 32633 2666 32634 2730
rect 32568 2650 32634 2666
rect 32568 2586 32569 2650
rect 32633 2586 32634 2650
rect 32568 2570 32634 2586
rect 32568 2506 32569 2570
rect 32633 2506 32634 2570
rect 32568 2490 32634 2506
rect 32568 2426 32569 2490
rect 32633 2426 32634 2490
rect 32568 2410 32634 2426
rect 32568 2346 32569 2410
rect 32633 2346 32634 2410
rect 32568 2330 32634 2346
rect 32568 2266 32569 2330
rect 32633 2266 32634 2330
rect 32568 2250 32634 2266
rect 32568 2186 32569 2250
rect 32633 2186 32634 2250
rect 32568 2170 32634 2186
rect 32568 2106 32569 2170
rect 32633 2106 32634 2170
rect 32568 2090 32634 2106
rect 32568 2026 32569 2090
rect 32633 2026 32634 2090
rect 32568 1936 32634 2026
rect 32694 1872 32754 2902
rect 32814 1932 32874 2964
rect 32934 1872 32994 2902
rect 33054 1932 33114 2964
rect 33174 2810 33240 2964
rect 33174 2746 33175 2810
rect 33239 2746 33240 2810
rect 33174 2730 33240 2746
rect 33174 2666 33175 2730
rect 33239 2666 33240 2730
rect 33174 2650 33240 2666
rect 33174 2586 33175 2650
rect 33239 2586 33240 2650
rect 33174 2570 33240 2586
rect 33174 2506 33175 2570
rect 33239 2506 33240 2570
rect 33174 2490 33240 2506
rect 33174 2426 33175 2490
rect 33239 2426 33240 2490
rect 33174 2410 33240 2426
rect 33174 2346 33175 2410
rect 33239 2346 33240 2410
rect 33174 2330 33240 2346
rect 33174 2266 33175 2330
rect 33239 2266 33240 2330
rect 33174 2250 33240 2266
rect 33174 2186 33175 2250
rect 33239 2186 33240 2250
rect 33174 2170 33240 2186
rect 33174 2106 33175 2170
rect 33239 2106 33240 2170
rect 33174 2090 33240 2106
rect 33174 2026 33175 2090
rect 33239 2026 33240 2090
rect 33174 1936 33240 2026
rect 13782 1870 33240 1872
rect 13782 1806 13886 1870
rect 13950 1806 13966 1870
rect 14030 1806 14046 1870
rect 14110 1806 14126 1870
rect 14190 1806 14206 1870
rect 14270 1806 14286 1870
rect 14350 1806 14492 1870
rect 14556 1806 14572 1870
rect 14636 1806 14652 1870
rect 14716 1806 14732 1870
rect 14796 1806 14812 1870
rect 14876 1806 14892 1870
rect 14956 1806 15098 1870
rect 15162 1806 15178 1870
rect 15242 1806 15258 1870
rect 15322 1806 15338 1870
rect 15402 1806 15418 1870
rect 15482 1806 15498 1870
rect 15562 1806 15704 1870
rect 15768 1806 15784 1870
rect 15848 1806 15864 1870
rect 15928 1806 15944 1870
rect 16008 1806 16024 1870
rect 16088 1806 16104 1870
rect 16168 1806 16310 1870
rect 16374 1806 16390 1870
rect 16454 1806 16470 1870
rect 16534 1806 16550 1870
rect 16614 1806 16630 1870
rect 16694 1806 16710 1870
rect 16774 1806 16916 1870
rect 16980 1806 16996 1870
rect 17060 1806 17076 1870
rect 17140 1806 17156 1870
rect 17220 1806 17236 1870
rect 17300 1806 17316 1870
rect 17380 1806 17522 1870
rect 17586 1806 17602 1870
rect 17666 1806 17682 1870
rect 17746 1806 17762 1870
rect 17826 1806 17842 1870
rect 17906 1806 17922 1870
rect 17986 1806 18128 1870
rect 18192 1806 18208 1870
rect 18272 1806 18288 1870
rect 18352 1806 18368 1870
rect 18432 1806 18448 1870
rect 18512 1806 18528 1870
rect 18592 1806 18734 1870
rect 18798 1806 18814 1870
rect 18878 1806 18894 1870
rect 18958 1806 18974 1870
rect 19038 1806 19054 1870
rect 19118 1806 19134 1870
rect 19198 1806 19340 1870
rect 19404 1806 19420 1870
rect 19484 1806 19500 1870
rect 19564 1806 19580 1870
rect 19644 1806 19660 1870
rect 19724 1806 19740 1870
rect 19804 1806 19946 1870
rect 20010 1806 20026 1870
rect 20090 1806 20106 1870
rect 20170 1806 20186 1870
rect 20250 1806 20266 1870
rect 20330 1806 20346 1870
rect 20410 1806 20552 1870
rect 20616 1806 20632 1870
rect 20696 1806 20712 1870
rect 20776 1806 20792 1870
rect 20856 1806 20872 1870
rect 20936 1806 20952 1870
rect 21016 1806 21158 1870
rect 21222 1806 21238 1870
rect 21302 1806 21318 1870
rect 21382 1806 21398 1870
rect 21462 1806 21478 1870
rect 21542 1806 21558 1870
rect 21622 1806 21764 1870
rect 21828 1806 21844 1870
rect 21908 1806 21924 1870
rect 21988 1806 22004 1870
rect 22068 1806 22084 1870
rect 22148 1806 22164 1870
rect 22228 1806 22370 1870
rect 22434 1806 22450 1870
rect 22514 1806 22530 1870
rect 22594 1806 22610 1870
rect 22674 1806 22690 1870
rect 22754 1806 22770 1870
rect 22834 1806 22976 1870
rect 23040 1806 23056 1870
rect 23120 1806 23136 1870
rect 23200 1806 23216 1870
rect 23280 1806 23296 1870
rect 23360 1806 23376 1870
rect 23440 1806 23582 1870
rect 23646 1806 23662 1870
rect 23726 1806 23742 1870
rect 23806 1806 23822 1870
rect 23886 1806 23902 1870
rect 23966 1806 23982 1870
rect 24046 1806 24188 1870
rect 24252 1806 24268 1870
rect 24332 1806 24348 1870
rect 24412 1806 24428 1870
rect 24492 1806 24508 1870
rect 24572 1806 24588 1870
rect 24652 1806 24794 1870
rect 24858 1806 24874 1870
rect 24938 1806 24954 1870
rect 25018 1806 25034 1870
rect 25098 1806 25114 1870
rect 25178 1806 25194 1870
rect 25258 1806 25400 1870
rect 25464 1806 25480 1870
rect 25544 1806 25560 1870
rect 25624 1806 25640 1870
rect 25704 1806 25720 1870
rect 25784 1806 25800 1870
rect 25864 1806 26006 1870
rect 26070 1806 26086 1870
rect 26150 1806 26166 1870
rect 26230 1806 26246 1870
rect 26310 1806 26326 1870
rect 26390 1806 26406 1870
rect 26470 1806 26612 1870
rect 26676 1806 26692 1870
rect 26756 1806 26772 1870
rect 26836 1806 26852 1870
rect 26916 1806 26932 1870
rect 26996 1806 27012 1870
rect 27076 1806 27218 1870
rect 27282 1806 27298 1870
rect 27362 1806 27378 1870
rect 27442 1806 27458 1870
rect 27522 1806 27538 1870
rect 27602 1806 27618 1870
rect 27682 1806 27824 1870
rect 27888 1806 27904 1870
rect 27968 1806 27984 1870
rect 28048 1806 28064 1870
rect 28128 1806 28144 1870
rect 28208 1806 28224 1870
rect 28288 1806 28430 1870
rect 28494 1806 28510 1870
rect 28574 1806 28590 1870
rect 28654 1806 28670 1870
rect 28734 1806 28750 1870
rect 28814 1806 28830 1870
rect 28894 1806 29036 1870
rect 29100 1806 29116 1870
rect 29180 1806 29196 1870
rect 29260 1806 29276 1870
rect 29340 1806 29356 1870
rect 29420 1806 29436 1870
rect 29500 1806 29642 1870
rect 29706 1806 29722 1870
rect 29786 1806 29802 1870
rect 29866 1806 29882 1870
rect 29946 1806 29962 1870
rect 30026 1806 30042 1870
rect 30106 1806 30248 1870
rect 30312 1806 30328 1870
rect 30392 1806 30408 1870
rect 30472 1806 30488 1870
rect 30552 1806 30568 1870
rect 30632 1806 30648 1870
rect 30712 1806 30854 1870
rect 30918 1806 30934 1870
rect 30998 1806 31014 1870
rect 31078 1806 31094 1870
rect 31158 1806 31174 1870
rect 31238 1806 31254 1870
rect 31318 1806 31460 1870
rect 31524 1806 31540 1870
rect 31604 1806 31620 1870
rect 31684 1806 31700 1870
rect 31764 1806 31780 1870
rect 31844 1806 31860 1870
rect 31924 1806 32066 1870
rect 32130 1806 32146 1870
rect 32210 1806 32226 1870
rect 32290 1806 32306 1870
rect 32370 1806 32386 1870
rect 32450 1806 32466 1870
rect 32530 1806 32672 1870
rect 32736 1806 32752 1870
rect 32816 1806 32832 1870
rect 32896 1806 32912 1870
rect 32976 1806 32992 1870
rect 33056 1806 33072 1870
rect 33136 1806 33240 1870
rect 13782 1804 33240 1806
<< labels >>
flabel psubdiff 22704 3266 22746 3356 0 FreeSans 320 0 0 0 SUB
port 1 nsew
flabel metal4 22520 3210 22566 3280 0 FreeSans 320 0 0 0 CTOP
port 3 nsew
flabel metal4 22638 2536 22684 2606 0 FreeSans 320 0 0 0 CTOP
port 5 nsew
flabel metal4 22760 2806 22806 2876 0 FreeSans 320 0 0 0 CBOT
port 7 nsew
flabel pwell 14102 2220 14128 2252 0 FreeSans 160 0 0 0 x1[1].SUB
flabel metal4 14044 2554 14070 2586 0 FreeSans 320 0 0 0 x1[1].CBOT
flabel metal4 14162 1964 14188 1996 0 FreeSans 320 0 0 0 x1[1].CTOP
flabel pwell 16526 2220 16552 2252 0 FreeSans 160 0 0 0 x1[9].SUB
flabel metal4 16468 2554 16494 2586 0 FreeSans 320 0 0 0 x1[9].CBOT
flabel metal4 16586 1964 16612 1996 0 FreeSans 320 0 0 0 x1[9].CTOP
flabel pwell 15920 2220 15946 2252 0 FreeSans 160 0 0 0 x1[7].SUB
flabel metal4 15862 2554 15888 2586 0 FreeSans 320 0 0 0 x1[7].CBOT
flabel metal4 15980 1964 16006 1996 0 FreeSans 320 0 0 0 x1[7].CTOP
flabel pwell 15314 2220 15340 2252 0 FreeSans 160 0 0 0 x1[5].SUB
flabel metal4 15256 2554 15282 2586 0 FreeSans 320 0 0 0 x1[5].CBOT
flabel metal4 15374 1964 15400 1996 0 FreeSans 320 0 0 0 x1[5].CTOP
flabel pwell 14708 2220 14734 2252 0 FreeSans 160 0 0 0 x1[3].SUB
flabel metal4 14650 2554 14676 2586 0 FreeSans 320 0 0 0 x1[3].CBOT
flabel metal4 14768 1964 14794 1996 0 FreeSans 320 0 0 0 x1[3].CTOP
flabel pwell 17738 2220 17764 2252 0 FreeSans 160 0 0 0 x1[13].SUB
flabel metal4 17680 2554 17706 2586 0 FreeSans 320 0 0 0 x1[13].CBOT
flabel metal4 17798 1964 17824 1996 0 FreeSans 320 0 0 0 x1[13].CTOP
flabel pwell 17132 2220 17158 2252 0 FreeSans 160 0 0 0 x1[11].SUB
flabel metal4 17074 2554 17100 2586 0 FreeSans 320 0 0 0 x1[11].CBOT
flabel metal4 17192 1964 17218 1996 0 FreeSans 320 0 0 0 x1[11].CTOP
flabel pwell 21374 2220 21400 2252 0 FreeSans 160 0 0 0 x1[25].SUB
flabel metal4 21316 2554 21342 2586 0 FreeSans 320 0 0 0 x1[25].CBOT
flabel metal4 21434 1964 21460 1996 0 FreeSans 320 0 0 0 x1[25].CTOP
flabel pwell 18950 2220 18976 2252 0 FreeSans 160 0 0 0 x1[17].SUB
flabel metal4 18892 2554 18918 2586 0 FreeSans 320 0 0 0 x1[17].CBOT
flabel metal4 19010 1964 19036 1996 0 FreeSans 320 0 0 0 x1[17].CTOP
flabel pwell 18344 2220 18370 2252 0 FreeSans 160 0 0 0 x1[15].SUB
flabel metal4 18286 2554 18312 2586 0 FreeSans 320 0 0 0 x1[15].CBOT
flabel metal4 18404 1964 18430 1996 0 FreeSans 320 0 0 0 x1[15].CTOP
flabel pwell 20768 2220 20794 2252 0 FreeSans 160 0 0 0 x1[23].SUB
flabel metal4 20710 2554 20736 2586 0 FreeSans 320 0 0 0 x1[23].CBOT
flabel metal4 20828 1964 20854 1996 0 FreeSans 320 0 0 0 x1[23].CTOP
flabel pwell 20162 2220 20188 2252 0 FreeSans 160 0 0 0 x1[21].SUB
flabel metal4 20104 2554 20130 2586 0 FreeSans 320 0 0 0 x1[21].CBOT
flabel metal4 20222 1964 20248 1996 0 FreeSans 320 0 0 0 x1[21].CTOP
flabel pwell 19556 2220 19582 2252 0 FreeSans 160 0 0 0 x1[19].SUB
flabel metal4 19498 2554 19524 2586 0 FreeSans 320 0 0 0 x1[19].CBOT
flabel metal4 19616 1964 19642 1996 0 FreeSans 320 0 0 0 x1[19].CTOP
flabel pwell 25010 2220 25036 2252 0 FreeSans 160 0 0 0 x1[37].SUB
flabel metal4 24952 2554 24978 2586 0 FreeSans 320 0 0 0 x1[37].CBOT
flabel metal4 25070 1964 25096 1996 0 FreeSans 320 0 0 0 x1[37].CTOP
flabel pwell 24404 2220 24430 2252 0 FreeSans 160 0 0 0 x1[35].SUB
flabel metal4 24346 2554 24372 2586 0 FreeSans 320 0 0 0 x1[35].CBOT
flabel metal4 24464 1964 24490 1996 0 FreeSans 320 0 0 0 x1[35].CTOP
flabel pwell 23798 2220 23824 2252 0 FreeSans 160 0 0 0 x1[33].SUB
flabel metal4 23740 2554 23766 2586 0 FreeSans 320 0 0 0 x1[33].CBOT
flabel metal4 23858 1964 23884 1996 0 FreeSans 320 0 0 0 x1[33].CTOP
flabel pwell 23192 2220 23218 2252 0 FreeSans 160 0 0 0 x1[31].SUB
flabel metal4 23134 2554 23160 2586 0 FreeSans 320 0 0 0 x1[31].CBOT
flabel metal4 23252 1964 23278 1996 0 FreeSans 320 0 0 0 x1[31].CTOP
flabel pwell 22586 2220 22612 2252 0 FreeSans 160 0 0 0 x1[29].SUB
flabel metal4 22528 2554 22554 2586 0 FreeSans 320 0 0 0 x1[29].CBOT
flabel metal4 22646 1964 22672 1996 0 FreeSans 320 0 0 0 x1[29].CTOP
flabel pwell 21980 2220 22006 2252 0 FreeSans 160 0 0 0 x1[27].SUB
flabel metal4 21922 2554 21948 2586 0 FreeSans 320 0 0 0 x1[27].CBOT
flabel metal4 22040 1964 22066 1996 0 FreeSans 320 0 0 0 x1[27].CTOP
flabel pwell 28040 2220 28066 2252 0 FreeSans 160 0 0 0 x1[47].SUB
flabel metal4 27982 2554 28008 2586 0 FreeSans 320 0 0 0 x1[47].CBOT
flabel metal4 28100 1964 28126 1996 0 FreeSans 320 0 0 0 x1[47].CTOP
flabel pwell 27434 2220 27460 2252 0 FreeSans 160 0 0 0 x1[45].SUB
flabel metal4 27376 2554 27402 2586 0 FreeSans 320 0 0 0 x1[45].CBOT
flabel metal4 27494 1964 27520 1996 0 FreeSans 320 0 0 0 x1[45].CTOP
flabel pwell 26828 2220 26854 2252 0 FreeSans 160 0 0 0 x1[43].SUB
flabel metal4 26770 2554 26796 2586 0 FreeSans 320 0 0 0 x1[43].CBOT
flabel metal4 26888 1964 26914 1996 0 FreeSans 320 0 0 0 x1[43].CTOP
flabel pwell 26222 2220 26248 2252 0 FreeSans 160 0 0 0 x1[41].SUB
flabel metal4 26164 2554 26190 2586 0 FreeSans 320 0 0 0 x1[41].CBOT
flabel metal4 26282 1964 26308 1996 0 FreeSans 320 0 0 0 x1[41].CTOP
flabel pwell 25616 2220 25642 2252 0 FreeSans 160 0 0 0 x1[39].SUB
flabel metal4 25558 2554 25584 2586 0 FreeSans 320 0 0 0 x1[39].CBOT
flabel metal4 25676 1964 25702 1996 0 FreeSans 320 0 0 0 x1[39].CTOP
flabel pwell 31676 2220 31702 2252 0 FreeSans 160 0 0 0 x1[59].SUB
flabel metal4 31618 2554 31644 2586 0 FreeSans 320 0 0 0 x1[59].CBOT
flabel metal4 31736 1964 31762 1996 0 FreeSans 320 0 0 0 x1[59].CTOP
flabel pwell 31070 2220 31096 2252 0 FreeSans 160 0 0 0 x1[57].SUB
flabel metal4 31012 2554 31038 2586 0 FreeSans 320 0 0 0 x1[57].CBOT
flabel metal4 31130 1964 31156 1996 0 FreeSans 320 0 0 0 x1[57].CTOP
flabel pwell 30464 2220 30490 2252 0 FreeSans 160 0 0 0 x1[55].SUB
flabel metal4 30406 2554 30432 2586 0 FreeSans 320 0 0 0 x1[55].CBOT
flabel metal4 30524 1964 30550 1996 0 FreeSans 320 0 0 0 x1[55].CTOP
flabel pwell 29858 2220 29884 2252 0 FreeSans 160 0 0 0 x1[53].SUB
flabel metal4 29800 2554 29826 2586 0 FreeSans 320 0 0 0 x1[53].CBOT
flabel metal4 29918 1964 29944 1996 0 FreeSans 320 0 0 0 x1[53].CTOP
flabel pwell 29252 2220 29278 2252 0 FreeSans 160 0 0 0 x1[51].SUB
flabel metal4 29194 2554 29220 2586 0 FreeSans 320 0 0 0 x1[51].CBOT
flabel metal4 29312 1964 29338 1996 0 FreeSans 320 0 0 0 x1[51].CTOP
flabel pwell 28646 2220 28672 2252 0 FreeSans 160 0 0 0 x1[49].SUB
flabel metal4 28588 2554 28614 2586 0 FreeSans 320 0 0 0 x1[49].CBOT
flabel metal4 28706 1964 28732 1996 0 FreeSans 320 0 0 0 x1[49].CTOP
flabel pwell 32888 2220 32914 2252 0 FreeSans 160 0 0 0 x1[63].SUB
flabel metal4 32830 2554 32856 2586 0 FreeSans 320 0 0 0 x1[63].CBOT
flabel metal4 32948 1964 32974 1996 0 FreeSans 320 0 0 0 x1[63].CTOP
flabel pwell 32282 2220 32308 2252 0 FreeSans 160 0 0 0 x1[61].SUB
flabel metal4 32224 2554 32250 2586 0 FreeSans 320 0 0 0 x1[61].CBOT
flabel metal4 32342 1964 32368 1996 0 FreeSans 320 0 0 0 x1[61].CTOP
flabel pwell 14108 3744 14134 3776 0 FreeSans 160 0 0 0 x1[0].SUB
flabel metal4 14166 3410 14192 3442 0 FreeSans 320 0 0 0 x1[0].CBOT
flabel metal4 14048 4000 14074 4032 0 FreeSans 320 0 0 0 x1[0].CTOP
flabel pwell 17744 3744 17770 3776 0 FreeSans 160 0 0 0 x1[12].SUB
flabel metal4 17802 3410 17828 3442 0 FreeSans 320 0 0 0 x1[12].CBOT
flabel metal4 17684 4000 17710 4032 0 FreeSans 320 0 0 0 x1[12].CTOP
flabel pwell 17138 3744 17164 3776 0 FreeSans 160 0 0 0 x1[10].SUB
flabel metal4 17196 3410 17222 3442 0 FreeSans 320 0 0 0 x1[10].CBOT
flabel metal4 17078 4000 17104 4032 0 FreeSans 320 0 0 0 x1[10].CTOP
flabel pwell 16532 3744 16558 3776 0 FreeSans 160 0 0 0 x1[8].SUB
flabel metal4 16590 3410 16616 3442 0 FreeSans 320 0 0 0 x1[8].CBOT
flabel metal4 16472 4000 16498 4032 0 FreeSans 320 0 0 0 x1[8].CTOP
flabel pwell 15926 3744 15952 3776 0 FreeSans 160 0 0 0 x1[6].SUB
flabel metal4 15984 3410 16010 3442 0 FreeSans 320 0 0 0 x1[6].CBOT
flabel metal4 15866 4000 15892 4032 0 FreeSans 320 0 0 0 x1[6].CTOP
flabel pwell 15320 3744 15346 3776 0 FreeSans 160 0 0 0 x1[4].SUB
flabel metal4 15378 3410 15404 3442 0 FreeSans 320 0 0 0 x1[4].CBOT
flabel metal4 15260 4000 15286 4032 0 FreeSans 320 0 0 0 x1[4].CTOP
flabel pwell 14714 3744 14740 3776 0 FreeSans 160 0 0 0 x1[2].SUB
flabel metal4 14772 3410 14798 3442 0 FreeSans 320 0 0 0 x1[2].CBOT
flabel metal4 14654 4000 14680 4032 0 FreeSans 320 0 0 0 x1[2].CTOP
flabel pwell 21380 3744 21406 3776 0 FreeSans 160 0 0 0 x1[24].SUB
flabel metal4 21438 3410 21464 3442 0 FreeSans 320 0 0 0 x1[24].CBOT
flabel metal4 21320 4000 21346 4032 0 FreeSans 320 0 0 0 x1[24].CTOP
flabel pwell 20774 3744 20800 3776 0 FreeSans 160 0 0 0 x1[22].SUB
flabel metal4 20832 3410 20858 3442 0 FreeSans 320 0 0 0 x1[22].CBOT
flabel metal4 20714 4000 20740 4032 0 FreeSans 320 0 0 0 x1[22].CTOP
flabel pwell 20168 3744 20194 3776 0 FreeSans 160 0 0 0 x1[20].SUB
flabel metal4 20226 3410 20252 3442 0 FreeSans 320 0 0 0 x1[20].CBOT
flabel metal4 20108 4000 20134 4032 0 FreeSans 320 0 0 0 x1[20].CTOP
flabel pwell 19562 3744 19588 3776 0 FreeSans 160 0 0 0 x1[18].SUB
flabel metal4 19620 3410 19646 3442 0 FreeSans 320 0 0 0 x1[18].CBOT
flabel metal4 19502 4000 19528 4032 0 FreeSans 320 0 0 0 x1[18].CTOP
flabel pwell 18956 3744 18982 3776 0 FreeSans 160 0 0 0 x1[16].SUB
flabel metal4 19014 3410 19040 3442 0 FreeSans 320 0 0 0 x1[16].CBOT
flabel metal4 18896 4000 18922 4032 0 FreeSans 320 0 0 0 x1[16].CTOP
flabel pwell 18350 3744 18376 3776 0 FreeSans 160 0 0 0 x1[14].SUB
flabel metal4 18408 3410 18434 3442 0 FreeSans 320 0 0 0 x1[14].CBOT
flabel metal4 18290 4000 18316 4032 0 FreeSans 320 0 0 0 x1[14].CTOP
flabel pwell 25016 3744 25042 3776 0 FreeSans 160 0 0 0 x1[36].SUB
flabel metal4 25074 3410 25100 3442 0 FreeSans 320 0 0 0 x1[36].CBOT
flabel metal4 24956 4000 24982 4032 0 FreeSans 320 0 0 0 x1[36].CTOP
flabel pwell 24410 3744 24436 3776 0 FreeSans 160 0 0 0 x1[34].SUB
flabel metal4 24468 3410 24494 3442 0 FreeSans 320 0 0 0 x1[34].CBOT
flabel metal4 24350 4000 24376 4032 0 FreeSans 320 0 0 0 x1[34].CTOP
flabel pwell 23804 3744 23830 3776 0 FreeSans 160 0 0 0 x1[32].SUB
flabel metal4 23862 3410 23888 3442 0 FreeSans 320 0 0 0 x1[32].CBOT
flabel metal4 23744 4000 23770 4032 0 FreeSans 320 0 0 0 x1[32].CTOP
flabel pwell 23198 3744 23224 3776 0 FreeSans 160 0 0 0 x1[30].SUB
flabel metal4 23256 3410 23282 3442 0 FreeSans 320 0 0 0 x1[30].CBOT
flabel metal4 23138 4000 23164 4032 0 FreeSans 320 0 0 0 x1[30].CTOP
flabel pwell 22592 3744 22618 3776 0 FreeSans 160 0 0 0 x1[28].SUB
flabel metal4 22650 3410 22676 3442 0 FreeSans 320 0 0 0 x1[28].CBOT
flabel metal4 22532 4000 22558 4032 0 FreeSans 320 0 0 0 x1[28].CTOP
flabel pwell 21986 3744 22012 3776 0 FreeSans 160 0 0 0 x1[26].SUB
flabel metal4 22044 3410 22070 3442 0 FreeSans 320 0 0 0 x1[26].CBOT
flabel metal4 21926 4000 21952 4032 0 FreeSans 320 0 0 0 x1[26].CTOP
flabel pwell 28046 3744 28072 3776 0 FreeSans 160 0 0 0 x1[46].SUB
flabel metal4 28104 3410 28130 3442 0 FreeSans 320 0 0 0 x1[46].CBOT
flabel metal4 27986 4000 28012 4032 0 FreeSans 320 0 0 0 x1[46].CTOP
flabel pwell 27440 3744 27466 3776 0 FreeSans 160 0 0 0 x1[44].SUB
flabel metal4 27498 3410 27524 3442 0 FreeSans 320 0 0 0 x1[44].CBOT
flabel metal4 27380 4000 27406 4032 0 FreeSans 320 0 0 0 x1[44].CTOP
flabel pwell 26834 3744 26860 3776 0 FreeSans 160 0 0 0 x1[42].SUB
flabel metal4 26892 3410 26918 3442 0 FreeSans 320 0 0 0 x1[42].CBOT
flabel metal4 26774 4000 26800 4032 0 FreeSans 320 0 0 0 x1[42].CTOP
flabel pwell 26228 3744 26254 3776 0 FreeSans 160 0 0 0 x1[40].SUB
flabel metal4 26286 3410 26312 3442 0 FreeSans 320 0 0 0 x1[40].CBOT
flabel metal4 26168 4000 26194 4032 0 FreeSans 320 0 0 0 x1[40].CTOP
flabel pwell 25622 3744 25648 3776 0 FreeSans 160 0 0 0 x1[38].SUB
flabel metal4 25680 3410 25706 3442 0 FreeSans 320 0 0 0 x1[38].CBOT
flabel metal4 25562 4000 25588 4032 0 FreeSans 320 0 0 0 x1[38].CTOP
flabel pwell 31682 3744 31708 3776 0 FreeSans 160 0 0 0 x1[58].SUB
flabel metal4 31740 3410 31766 3442 0 FreeSans 320 0 0 0 x1[58].CBOT
flabel metal4 31622 4000 31648 4032 0 FreeSans 320 0 0 0 x1[58].CTOP
flabel pwell 31076 3744 31102 3776 0 FreeSans 160 0 0 0 x1[56].SUB
flabel metal4 31134 3410 31160 3442 0 FreeSans 320 0 0 0 x1[56].CBOT
flabel metal4 31016 4000 31042 4032 0 FreeSans 320 0 0 0 x1[56].CTOP
flabel pwell 30470 3744 30496 3776 0 FreeSans 160 0 0 0 x1[54].SUB
flabel metal4 30528 3410 30554 3442 0 FreeSans 320 0 0 0 x1[54].CBOT
flabel metal4 30410 4000 30436 4032 0 FreeSans 320 0 0 0 x1[54].CTOP
flabel pwell 29864 3744 29890 3776 0 FreeSans 160 0 0 0 x1[52].SUB
flabel metal4 29922 3410 29948 3442 0 FreeSans 320 0 0 0 x1[52].CBOT
flabel metal4 29804 4000 29830 4032 0 FreeSans 320 0 0 0 x1[52].CTOP
flabel pwell 29258 3744 29284 3776 0 FreeSans 160 0 0 0 x1[50].SUB
flabel metal4 29316 3410 29342 3442 0 FreeSans 320 0 0 0 x1[50].CBOT
flabel metal4 29198 4000 29224 4032 0 FreeSans 320 0 0 0 x1[50].CTOP
flabel pwell 28652 3744 28678 3776 0 FreeSans 160 0 0 0 x1[48].SUB
flabel metal4 28710 3410 28736 3442 0 FreeSans 320 0 0 0 x1[48].CBOT
flabel metal4 28592 4000 28618 4032 0 FreeSans 320 0 0 0 x1[48].CTOP
flabel pwell 32894 3744 32920 3776 0 FreeSans 160 0 0 0 x1[62].SUB
flabel metal4 32952 3410 32978 3442 0 FreeSans 320 0 0 0 x1[62].CBOT
flabel metal4 32834 4000 32860 4032 0 FreeSans 320 0 0 0 x1[62].CTOP
flabel pwell 32288 3744 32314 3776 0 FreeSans 160 0 0 0 x1[60].SUB
flabel metal4 32346 3410 32372 3442 0 FreeSans 320 0 0 0 x1[60].CBOT
flabel metal4 32228 4000 32254 4032 0 FreeSans 320 0 0 0 x1[60].CTOP
<< end >>
