magic
tech sky130A
magscale 1 2
timestamp 1698286991
use hgu_inverter  x1
timestamp 1698286873
transform 1 0 53 0 1 2200
box 372 160 690 825
use hgu_inverter  x2
timestamp 1698286873
transform -1 0 1203 0 1 2200
box 372 160 690 825
<< end >>
