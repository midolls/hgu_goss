magic
tech sky130A
magscale 1 2
timestamp 1698022638
<< checkpaint >>
rect -1260 -2860 1460 1460
<< pwell >>
rect 1006 1014 1032 1046
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
<< metal3 >>
rect 686 1514 1478 1516
rect 686 1450 766 1514
rect 830 1450 846 1514
rect 910 1450 926 1514
rect 990 1450 1006 1514
rect 1070 1450 1086 1514
rect 1150 1450 1166 1514
rect 1230 1450 1246 1514
rect 1310 1450 1326 1514
rect 1390 1450 1478 1514
rect 686 1448 1478 1450
rect 686 1414 752 1448
rect 686 1350 687 1414
rect 751 1350 752 1414
rect 686 1334 752 1350
rect 686 1270 687 1334
rect 751 1270 752 1334
rect 686 1254 752 1270
rect 686 1190 687 1254
rect 751 1190 752 1254
rect 686 1174 752 1190
rect 686 1110 687 1174
rect 751 1110 752 1174
rect 686 1094 752 1110
rect 686 1030 687 1094
rect 751 1030 752 1094
rect 686 1014 752 1030
rect 686 950 687 1014
rect 751 950 752 1014
rect 686 934 752 950
rect 686 870 687 934
rect 751 870 752 934
rect 686 854 752 870
rect 686 790 687 854
rect 751 790 752 854
rect 686 724 752 790
rect 812 726 872 1448
rect 932 666 992 1388
rect 1052 726 1112 1448
rect 1172 666 1232 1388
rect 1292 726 1352 1448
rect 1412 1414 1478 1448
rect 1412 1350 1413 1414
rect 1477 1350 1478 1414
rect 1412 1334 1478 1350
rect 1412 1270 1413 1334
rect 1477 1270 1478 1334
rect 1412 1254 1478 1270
rect 1412 1190 1413 1254
rect 1477 1190 1478 1254
rect 1412 1174 1478 1190
rect 1412 1110 1413 1174
rect 1477 1110 1478 1174
rect 1412 1094 1478 1110
rect 1412 1030 1413 1094
rect 1477 1030 1478 1094
rect 1412 1014 1478 1030
rect 1412 950 1413 1014
rect 1477 950 1478 1014
rect 1412 934 1478 950
rect 1412 870 1413 934
rect 1477 870 1478 934
rect 1412 854 1478 870
rect 1412 790 1413 854
rect 1477 790 1478 854
rect 1412 724 1478 790
rect 812 664 1354 666
rect 812 600 888 664
rect 952 600 968 664
rect 1032 600 1048 664
rect 1112 600 1128 664
rect 1192 600 1208 664
rect 1272 600 1354 664
rect 812 598 1354 600
rect 862 596 1294 598
<< via3 >>
rect 766 1450 830 1514
rect 846 1450 910 1514
rect 926 1450 990 1514
rect 1006 1450 1070 1514
rect 1086 1450 1150 1514
rect 1166 1450 1230 1514
rect 1246 1450 1310 1514
rect 1326 1450 1390 1514
rect 687 1350 751 1414
rect 687 1270 751 1334
rect 687 1190 751 1254
rect 687 1110 751 1174
rect 687 1030 751 1094
rect 687 950 751 1014
rect 687 870 751 934
rect 687 790 751 854
rect 1413 1350 1477 1414
rect 1413 1270 1477 1334
rect 1413 1190 1477 1254
rect 1413 1110 1477 1174
rect 1413 1030 1477 1094
rect 1413 950 1477 1014
rect 1413 870 1477 934
rect 1413 790 1477 854
rect 888 600 952 664
rect 968 600 1032 664
rect 1048 600 1112 664
rect 1128 600 1192 664
rect 1208 600 1272 664
<< metal4 >>
rect 686 1514 1478 1516
rect 686 1450 766 1514
rect 830 1450 846 1514
rect 910 1450 926 1514
rect 990 1450 1006 1514
rect 1070 1450 1086 1514
rect 1150 1450 1166 1514
rect 1230 1450 1246 1514
rect 1310 1450 1326 1514
rect 1390 1450 1478 1514
rect 686 1448 1478 1450
rect 686 1414 752 1448
rect 686 1350 687 1414
rect 751 1350 752 1414
rect 686 1334 752 1350
rect 686 1270 687 1334
rect 751 1270 752 1334
rect 686 1254 752 1270
rect 686 1190 687 1254
rect 751 1190 752 1254
rect 686 1174 752 1190
rect 686 1110 687 1174
rect 751 1110 752 1174
rect 686 1094 752 1110
rect 686 1030 687 1094
rect 751 1030 752 1094
rect 686 1014 752 1030
rect 686 950 687 1014
rect 751 950 752 1014
rect 686 934 752 950
rect 686 870 687 934
rect 751 870 752 934
rect 686 854 752 870
rect 686 790 687 854
rect 751 790 752 854
rect 686 724 752 790
rect 812 666 872 1388
rect 932 726 992 1448
rect 1052 666 1112 1388
rect 1172 726 1232 1448
rect 1412 1414 1478 1448
rect 1292 666 1352 1388
rect 1412 1350 1413 1414
rect 1477 1350 1478 1414
rect 1412 1334 1478 1350
rect 1412 1270 1413 1334
rect 1477 1270 1478 1334
rect 1412 1254 1478 1270
rect 1412 1190 1413 1254
rect 1477 1190 1478 1254
rect 1412 1174 1478 1190
rect 1412 1110 1413 1174
rect 1477 1110 1478 1174
rect 1412 1094 1478 1110
rect 1412 1030 1413 1094
rect 1477 1030 1478 1094
rect 1412 1014 1478 1030
rect 1412 950 1413 1014
rect 1477 950 1478 1014
rect 1412 934 1478 950
rect 1412 870 1413 934
rect 1477 870 1478 934
rect 1412 854 1478 870
rect 1412 790 1413 854
rect 1477 790 1478 854
rect 1412 724 1478 790
rect 812 664 1354 666
rect 812 600 888 664
rect 952 600 968 664
rect 1032 600 1048 664
rect 1112 600 1128 664
rect 1192 600 1208 664
rect 1272 600 1354 664
rect 812 598 1354 600
rect 862 596 1294 598
use sky130_fd_pr__cap_vpp_02p4x04p6_m1m2_noshield  XC2 ../mag
timestamp 1697993263
transform 1 0 88 0 1 600
box -88 0 396 918
<< labels >>
flabel space 1006 1016 1032 1048 0 FreeSans 160 0 0 0 SUB
port 1 nsew
flabel metal4 948 1348 974 1380 0 FreeSans 320 0 0 0 C1
port 4 nsew
flabel metal4 1066 758 1092 790 0 FreeSans 320 0 0 0 C0
port 6 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 {}
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 csize=1
port 3 nsew
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 PLUS
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 MINUS
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 SUB
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 {}
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 csize=1
<< end >>
