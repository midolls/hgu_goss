* NGSPICE file created from hgu_cdac_cap_64.ext - technology: sky130A

.subckt hgu_cdac_cap_64 SUB
C0 x1[8].CTOP x1[9].CTOP 0.161p
C1 x1[9].CTOP x1[9].CBOT 0.161p
.ends

