magic
tech sky130A
magscale 1 2
timestamp 1700462216
<< nwell >>
rect -378 6072 -50 6456
rect 399 6072 855 6456
rect 1308 6072 2020 6456
rect 2841 6072 4065 6456
rect 5392 6072 7640 6456
rect 10479 6072 14775 6456
rect 20264 6072 28656 6456
rect -400 5384 -72 5768
rect 528 5384 984 5768
rect 1792 5384 2504 5768
rect 3411 5384 4635 5768
rect 7976 5384 10224 5768
rect 15134 5384 19430 5768
rect 20188 5384 28580 5768
<< pwell >>
rect 17436 3572 17468 3622
rect 17436 1084 17468 1134
<< pmoslvt >>
rect -249 6110 -179 6278
rect 528 6110 598 6278
rect 656 6110 726 6278
rect 1437 6110 1507 6278
rect 1565 6110 1635 6278
rect 1693 6110 1763 6278
rect 1821 6110 1891 6278
rect 2970 6110 3040 6278
rect 3098 6110 3168 6278
rect 3226 6110 3296 6278
rect 3354 6110 3424 6278
rect 3482 6110 3552 6278
rect 3610 6110 3680 6278
rect 3738 6110 3808 6278
rect 3866 6110 3936 6278
rect 5521 6110 5591 6278
rect 5649 6110 5719 6278
rect 5777 6110 5847 6278
rect 5905 6110 5975 6278
rect 6033 6110 6103 6278
rect 6161 6110 6231 6278
rect 6289 6110 6359 6278
rect 6417 6110 6487 6278
rect 6545 6110 6615 6278
rect 6673 6110 6743 6278
rect 6801 6110 6871 6278
rect 6929 6110 6999 6278
rect 7057 6110 7127 6278
rect 7185 6110 7255 6278
rect 7313 6110 7383 6278
rect 7441 6110 7511 6278
rect 10608 6110 10678 6278
rect 10736 6110 10806 6278
rect 10864 6110 10934 6278
rect 10992 6110 11062 6278
rect 11120 6110 11190 6278
rect 11248 6110 11318 6278
rect 11376 6110 11446 6278
rect 11504 6110 11574 6278
rect 11632 6110 11702 6278
rect 11760 6110 11830 6278
rect 11888 6110 11958 6278
rect 12016 6110 12086 6278
rect 12144 6110 12214 6278
rect 12272 6110 12342 6278
rect 12400 6110 12470 6278
rect 12528 6110 12598 6278
rect 12656 6110 12726 6278
rect 12784 6110 12854 6278
rect 12912 6110 12982 6278
rect 13040 6110 13110 6278
rect 13168 6110 13238 6278
rect 13296 6110 13366 6278
rect 13424 6110 13494 6278
rect 13552 6110 13622 6278
rect 13680 6110 13750 6278
rect 13808 6110 13878 6278
rect 13936 6110 14006 6278
rect 14064 6110 14134 6278
rect 14192 6110 14262 6278
rect 14320 6110 14390 6278
rect 14448 6110 14518 6278
rect 14576 6110 14646 6278
rect 20393 6110 20463 6278
rect 20521 6110 20591 6278
rect 20649 6110 20719 6278
rect 20777 6110 20847 6278
rect 20905 6110 20975 6278
rect 21033 6110 21103 6278
rect 21161 6110 21231 6278
rect 21289 6110 21359 6278
rect 21417 6110 21487 6278
rect 21545 6110 21615 6278
rect 21673 6110 21743 6278
rect 21801 6110 21871 6278
rect 21929 6110 21999 6278
rect 22057 6110 22127 6278
rect 22185 6110 22255 6278
rect 22313 6110 22383 6278
rect 22441 6110 22511 6278
rect 22569 6110 22639 6278
rect 22697 6110 22767 6278
rect 22825 6110 22895 6278
rect 22953 6110 23023 6278
rect 23081 6110 23151 6278
rect 23209 6110 23279 6278
rect 23337 6110 23407 6278
rect 23465 6110 23535 6278
rect 23593 6110 23663 6278
rect 23721 6110 23791 6278
rect 23849 6110 23919 6278
rect 23977 6110 24047 6278
rect 24105 6110 24175 6278
rect 24233 6110 24303 6278
rect 24361 6110 24431 6278
rect 24489 6110 24559 6278
rect 24617 6110 24687 6278
rect 24745 6110 24815 6278
rect 24873 6110 24943 6278
rect 25001 6110 25071 6278
rect 25129 6110 25199 6278
rect 25257 6110 25327 6278
rect 25385 6110 25455 6278
rect 25513 6110 25583 6278
rect 25641 6110 25711 6278
rect 25769 6110 25839 6278
rect 25897 6110 25967 6278
rect 26025 6110 26095 6278
rect 26153 6110 26223 6278
rect 26281 6110 26351 6278
rect 26409 6110 26479 6278
rect 26537 6110 26607 6278
rect 26665 6110 26735 6278
rect 26793 6110 26863 6278
rect 26921 6110 26991 6278
rect 27049 6110 27119 6278
rect 27177 6110 27247 6278
rect 27305 6110 27375 6278
rect 27433 6110 27503 6278
rect 27561 6110 27631 6278
rect 27689 6110 27759 6278
rect 27817 6110 27887 6278
rect 27945 6110 28015 6278
rect 28073 6110 28143 6278
rect 28201 6110 28271 6278
rect 28329 6110 28399 6278
rect 28457 6110 28527 6278
rect -271 5422 -201 5590
rect 657 5422 727 5590
rect 785 5422 855 5590
rect 1921 5422 1991 5590
rect 2049 5422 2119 5590
rect 2177 5422 2247 5590
rect 2305 5422 2375 5590
rect 3540 5422 3610 5590
rect 3668 5422 3738 5590
rect 3796 5422 3866 5590
rect 3924 5422 3994 5590
rect 4052 5422 4122 5590
rect 4180 5422 4250 5590
rect 4308 5422 4378 5590
rect 4436 5422 4506 5590
rect 8105 5422 8175 5590
rect 8233 5422 8303 5590
rect 8361 5422 8431 5590
rect 8489 5422 8559 5590
rect 8617 5422 8687 5590
rect 8745 5422 8815 5590
rect 8873 5422 8943 5590
rect 9001 5422 9071 5590
rect 9129 5422 9199 5590
rect 9257 5422 9327 5590
rect 9385 5422 9455 5590
rect 9513 5422 9583 5590
rect 9641 5422 9711 5590
rect 9769 5422 9839 5590
rect 9897 5422 9967 5590
rect 10025 5422 10095 5590
rect 15263 5422 15333 5590
rect 15391 5422 15461 5590
rect 15519 5422 15589 5590
rect 15647 5422 15717 5590
rect 15775 5422 15845 5590
rect 15903 5422 15973 5590
rect 16031 5422 16101 5590
rect 16159 5422 16229 5590
rect 16287 5422 16357 5590
rect 16415 5422 16485 5590
rect 16543 5422 16613 5590
rect 16671 5422 16741 5590
rect 16799 5422 16869 5590
rect 16927 5422 16997 5590
rect 17055 5422 17125 5590
rect 17183 5422 17253 5590
rect 17311 5422 17381 5590
rect 17439 5422 17509 5590
rect 17567 5422 17637 5590
rect 17695 5422 17765 5590
rect 17823 5422 17893 5590
rect 17951 5422 18021 5590
rect 18079 5422 18149 5590
rect 18207 5422 18277 5590
rect 18335 5422 18405 5590
rect 18463 5422 18533 5590
rect 18591 5422 18661 5590
rect 18719 5422 18789 5590
rect 18847 5422 18917 5590
rect 18975 5422 19045 5590
rect 19103 5422 19173 5590
rect 19231 5422 19301 5590
rect 20317 5422 20387 5590
rect 20445 5422 20515 5590
rect 20573 5422 20643 5590
rect 20701 5422 20771 5590
rect 20829 5422 20899 5590
rect 20957 5422 21027 5590
rect 21085 5422 21155 5590
rect 21213 5422 21283 5590
rect 21341 5422 21411 5590
rect 21469 5422 21539 5590
rect 21597 5422 21667 5590
rect 21725 5422 21795 5590
rect 21853 5422 21923 5590
rect 21981 5422 22051 5590
rect 22109 5422 22179 5590
rect 22237 5422 22307 5590
rect 22365 5422 22435 5590
rect 22493 5422 22563 5590
rect 22621 5422 22691 5590
rect 22749 5422 22819 5590
rect 22877 5422 22947 5590
rect 23005 5422 23075 5590
rect 23133 5422 23203 5590
rect 23261 5422 23331 5590
rect 23389 5422 23459 5590
rect 23517 5422 23587 5590
rect 23645 5422 23715 5590
rect 23773 5422 23843 5590
rect 23901 5422 23971 5590
rect 24029 5422 24099 5590
rect 24157 5422 24227 5590
rect 24285 5422 24355 5590
rect 24413 5422 24483 5590
rect 24541 5422 24611 5590
rect 24669 5422 24739 5590
rect 24797 5422 24867 5590
rect 24925 5422 24995 5590
rect 25053 5422 25123 5590
rect 25181 5422 25251 5590
rect 25309 5422 25379 5590
rect 25437 5422 25507 5590
rect 25565 5422 25635 5590
rect 25693 5422 25763 5590
rect 25821 5422 25891 5590
rect 25949 5422 26019 5590
rect 26077 5422 26147 5590
rect 26205 5422 26275 5590
rect 26333 5422 26403 5590
rect 26461 5422 26531 5590
rect 26589 5422 26659 5590
rect 26717 5422 26787 5590
rect 26845 5422 26915 5590
rect 26973 5422 27043 5590
rect 27101 5422 27171 5590
rect 27229 5422 27299 5590
rect 27357 5422 27427 5590
rect 27485 5422 27555 5590
rect 27613 5422 27683 5590
rect 27741 5422 27811 5590
rect 27869 5422 27939 5590
rect 27997 5422 28067 5590
rect 28125 5422 28195 5590
rect 28253 5422 28323 5590
rect 28381 5422 28451 5590
<< nmoslvt >>
rect -249 5894 -179 5978
rect 528 5894 598 5978
rect 656 5894 726 5978
rect 1437 5894 1507 5978
rect 1565 5894 1635 5978
rect 1693 5894 1763 5978
rect 1821 5894 1891 5978
rect 2970 5894 3040 5978
rect 3098 5894 3168 5978
rect 3226 5894 3296 5978
rect 3354 5894 3424 5978
rect 3482 5894 3552 5978
rect 3610 5894 3680 5978
rect 3738 5894 3808 5978
rect 3866 5894 3936 5978
rect 5521 5894 5591 5978
rect 5649 5894 5719 5978
rect 5777 5894 5847 5978
rect 5905 5894 5975 5978
rect 6033 5894 6103 5978
rect 6161 5894 6231 5978
rect 6289 5894 6359 5978
rect 6417 5894 6487 5978
rect 6545 5894 6615 5978
rect 6673 5894 6743 5978
rect 6801 5894 6871 5978
rect 6929 5894 6999 5978
rect 7057 5894 7127 5978
rect 7185 5894 7255 5978
rect 7313 5894 7383 5978
rect 7441 5894 7511 5978
rect 10608 5894 10678 5978
rect 10736 5894 10806 5978
rect 10864 5894 10934 5978
rect 10992 5894 11062 5978
rect 11120 5894 11190 5978
rect 11248 5894 11318 5978
rect 11376 5894 11446 5978
rect 11504 5894 11574 5978
rect 11632 5894 11702 5978
rect 11760 5894 11830 5978
rect 11888 5894 11958 5978
rect 12016 5894 12086 5978
rect 12144 5894 12214 5978
rect 12272 5894 12342 5978
rect 12400 5894 12470 5978
rect 12528 5894 12598 5978
rect 12656 5894 12726 5978
rect 12784 5894 12854 5978
rect 12912 5894 12982 5978
rect 13040 5894 13110 5978
rect 13168 5894 13238 5978
rect 13296 5894 13366 5978
rect 13424 5894 13494 5978
rect 13552 5894 13622 5978
rect 13680 5894 13750 5978
rect 13808 5894 13878 5978
rect 13936 5894 14006 5978
rect 14064 5894 14134 5978
rect 14192 5894 14262 5978
rect 14320 5894 14390 5978
rect 14448 5894 14518 5978
rect 14576 5894 14646 5978
rect 20393 5894 20463 5978
rect 20521 5894 20591 5978
rect 20649 5894 20719 5978
rect 20777 5894 20847 5978
rect 20905 5894 20975 5978
rect 21033 5894 21103 5978
rect 21161 5894 21231 5978
rect 21289 5894 21359 5978
rect 21417 5894 21487 5978
rect 21545 5894 21615 5978
rect 21673 5894 21743 5978
rect 21801 5894 21871 5978
rect 21929 5894 21999 5978
rect 22057 5894 22127 5978
rect 22185 5894 22255 5978
rect 22313 5894 22383 5978
rect 22441 5894 22511 5978
rect 22569 5894 22639 5978
rect 22697 5894 22767 5978
rect 22825 5894 22895 5978
rect 22953 5894 23023 5978
rect 23081 5894 23151 5978
rect 23209 5894 23279 5978
rect 23337 5894 23407 5978
rect 23465 5894 23535 5978
rect 23593 5894 23663 5978
rect 23721 5894 23791 5978
rect 23849 5894 23919 5978
rect 23977 5894 24047 5978
rect 24105 5894 24175 5978
rect 24233 5894 24303 5978
rect 24361 5894 24431 5978
rect 24489 5894 24559 5978
rect 24617 5894 24687 5978
rect 24745 5894 24815 5978
rect 24873 5894 24943 5978
rect 25001 5894 25071 5978
rect 25129 5894 25199 5978
rect 25257 5894 25327 5978
rect 25385 5894 25455 5978
rect 25513 5894 25583 5978
rect 25641 5894 25711 5978
rect 25769 5894 25839 5978
rect 25897 5894 25967 5978
rect 26025 5894 26095 5978
rect 26153 5894 26223 5978
rect 26281 5894 26351 5978
rect 26409 5894 26479 5978
rect 26537 5894 26607 5978
rect 26665 5894 26735 5978
rect 26793 5894 26863 5978
rect 26921 5894 26991 5978
rect 27049 5894 27119 5978
rect 27177 5894 27247 5978
rect 27305 5894 27375 5978
rect 27433 5894 27503 5978
rect 27561 5894 27631 5978
rect 27689 5894 27759 5978
rect 27817 5894 27887 5978
rect 27945 5894 28015 5978
rect 28073 5894 28143 5978
rect 28201 5894 28271 5978
rect 28329 5894 28399 5978
rect 28457 5894 28527 5978
rect -271 5206 -201 5290
rect 657 5206 727 5290
rect 785 5206 855 5290
rect 1921 5206 1991 5290
rect 2049 5206 2119 5290
rect 2177 5206 2247 5290
rect 2305 5206 2375 5290
rect 3540 5206 3610 5290
rect 3668 5206 3738 5290
rect 3796 5206 3866 5290
rect 3924 5206 3994 5290
rect 4052 5206 4122 5290
rect 4180 5206 4250 5290
rect 4308 5206 4378 5290
rect 4436 5206 4506 5290
rect 8105 5206 8175 5290
rect 8233 5206 8303 5290
rect 8361 5206 8431 5290
rect 8489 5206 8559 5290
rect 8617 5206 8687 5290
rect 8745 5206 8815 5290
rect 8873 5206 8943 5290
rect 9001 5206 9071 5290
rect 9129 5206 9199 5290
rect 9257 5206 9327 5290
rect 9385 5206 9455 5290
rect 9513 5206 9583 5290
rect 9641 5206 9711 5290
rect 9769 5206 9839 5290
rect 9897 5206 9967 5290
rect 10025 5206 10095 5290
rect 15263 5206 15333 5290
rect 15391 5206 15461 5290
rect 15519 5206 15589 5290
rect 15647 5206 15717 5290
rect 15775 5206 15845 5290
rect 15903 5206 15973 5290
rect 16031 5206 16101 5290
rect 16159 5206 16229 5290
rect 16287 5206 16357 5290
rect 16415 5206 16485 5290
rect 16543 5206 16613 5290
rect 16671 5206 16741 5290
rect 16799 5206 16869 5290
rect 16927 5206 16997 5290
rect 17055 5206 17125 5290
rect 17183 5206 17253 5290
rect 17311 5206 17381 5290
rect 17439 5206 17509 5290
rect 17567 5206 17637 5290
rect 17695 5206 17765 5290
rect 17823 5206 17893 5290
rect 17951 5206 18021 5290
rect 18079 5206 18149 5290
rect 18207 5206 18277 5290
rect 18335 5206 18405 5290
rect 18463 5206 18533 5290
rect 18591 5206 18661 5290
rect 18719 5206 18789 5290
rect 18847 5206 18917 5290
rect 18975 5206 19045 5290
rect 19103 5206 19173 5290
rect 19231 5206 19301 5290
rect 20317 5206 20387 5290
rect 20445 5206 20515 5290
rect 20573 5206 20643 5290
rect 20701 5206 20771 5290
rect 20829 5206 20899 5290
rect 20957 5206 21027 5290
rect 21085 5206 21155 5290
rect 21213 5206 21283 5290
rect 21341 5206 21411 5290
rect 21469 5206 21539 5290
rect 21597 5206 21667 5290
rect 21725 5206 21795 5290
rect 21853 5206 21923 5290
rect 21981 5206 22051 5290
rect 22109 5206 22179 5290
rect 22237 5206 22307 5290
rect 22365 5206 22435 5290
rect 22493 5206 22563 5290
rect 22621 5206 22691 5290
rect 22749 5206 22819 5290
rect 22877 5206 22947 5290
rect 23005 5206 23075 5290
rect 23133 5206 23203 5290
rect 23261 5206 23331 5290
rect 23389 5206 23459 5290
rect 23517 5206 23587 5290
rect 23645 5206 23715 5290
rect 23773 5206 23843 5290
rect 23901 5206 23971 5290
rect 24029 5206 24099 5290
rect 24157 5206 24227 5290
rect 24285 5206 24355 5290
rect 24413 5206 24483 5290
rect 24541 5206 24611 5290
rect 24669 5206 24739 5290
rect 24797 5206 24867 5290
rect 24925 5206 24995 5290
rect 25053 5206 25123 5290
rect 25181 5206 25251 5290
rect 25309 5206 25379 5290
rect 25437 5206 25507 5290
rect 25565 5206 25635 5290
rect 25693 5206 25763 5290
rect 25821 5206 25891 5290
rect 25949 5206 26019 5290
rect 26077 5206 26147 5290
rect 26205 5206 26275 5290
rect 26333 5206 26403 5290
rect 26461 5206 26531 5290
rect 26589 5206 26659 5290
rect 26717 5206 26787 5290
rect 26845 5206 26915 5290
rect 26973 5206 27043 5290
rect 27101 5206 27171 5290
rect 27229 5206 27299 5290
rect 27357 5206 27427 5290
rect 27485 5206 27555 5290
rect 27613 5206 27683 5290
rect 27741 5206 27811 5290
rect 27869 5206 27939 5290
rect 27997 5206 28067 5290
rect 28125 5206 28195 5290
rect 28253 5206 28323 5290
rect 28381 5206 28451 5290
<< ndiff >>
rect -307 5966 -249 5978
rect -307 5906 -295 5966
rect -261 5906 -249 5966
rect -307 5894 -249 5906
rect -179 5966 -121 5978
rect -179 5906 -167 5966
rect -133 5906 -121 5966
rect -179 5894 -121 5906
rect 470 5966 528 5978
rect 470 5906 482 5966
rect 516 5906 528 5966
rect 470 5894 528 5906
rect 598 5966 656 5978
rect 598 5906 610 5966
rect 644 5906 656 5966
rect 598 5894 656 5906
rect 726 5966 784 5978
rect 726 5906 738 5966
rect 772 5906 784 5966
rect 726 5894 784 5906
rect 1379 5966 1437 5978
rect 1379 5906 1391 5966
rect 1425 5906 1437 5966
rect 1379 5894 1437 5906
rect 1507 5966 1565 5978
rect 1507 5906 1519 5966
rect 1553 5906 1565 5966
rect 1507 5894 1565 5906
rect 1635 5966 1693 5978
rect 1635 5906 1647 5966
rect 1681 5906 1693 5966
rect 1635 5894 1693 5906
rect 1763 5966 1821 5978
rect 1763 5906 1775 5966
rect 1809 5906 1821 5966
rect 1763 5894 1821 5906
rect 1891 5966 1949 5978
rect 1891 5906 1903 5966
rect 1937 5906 1949 5966
rect 1891 5894 1949 5906
rect 2912 5966 2970 5978
rect 2912 5906 2924 5966
rect 2958 5906 2970 5966
rect 2912 5894 2970 5906
rect 3040 5966 3098 5978
rect 3040 5906 3052 5966
rect 3086 5906 3098 5966
rect 3040 5894 3098 5906
rect 3168 5966 3226 5978
rect 3168 5906 3180 5966
rect 3214 5906 3226 5966
rect 3168 5894 3226 5906
rect 3296 5966 3354 5978
rect 3296 5906 3308 5966
rect 3342 5906 3354 5966
rect 3296 5894 3354 5906
rect 3424 5966 3482 5978
rect 3424 5906 3436 5966
rect 3470 5906 3482 5966
rect 3424 5894 3482 5906
rect 3552 5966 3610 5978
rect 3552 5906 3564 5966
rect 3598 5906 3610 5966
rect 3552 5894 3610 5906
rect 3680 5966 3738 5978
rect 3680 5906 3692 5966
rect 3726 5906 3738 5966
rect 3680 5894 3738 5906
rect 3808 5966 3866 5978
rect 3808 5906 3820 5966
rect 3854 5906 3866 5966
rect 3808 5894 3866 5906
rect 3936 5966 3994 5978
rect 3936 5906 3948 5966
rect 3982 5906 3994 5966
rect 3936 5894 3994 5906
rect 5463 5966 5521 5978
rect 5463 5906 5475 5966
rect 5509 5906 5521 5966
rect 5463 5894 5521 5906
rect 5591 5966 5649 5978
rect 5591 5906 5603 5966
rect 5637 5906 5649 5966
rect 5591 5894 5649 5906
rect 5719 5966 5777 5978
rect 5719 5906 5731 5966
rect 5765 5906 5777 5966
rect 5719 5894 5777 5906
rect 5847 5966 5905 5978
rect 5847 5906 5859 5966
rect 5893 5906 5905 5966
rect 5847 5894 5905 5906
rect 5975 5966 6033 5978
rect 5975 5906 5987 5966
rect 6021 5906 6033 5966
rect 5975 5894 6033 5906
rect 6103 5966 6161 5978
rect 6103 5906 6115 5966
rect 6149 5906 6161 5966
rect 6103 5894 6161 5906
rect 6231 5966 6289 5978
rect 6231 5906 6243 5966
rect 6277 5906 6289 5966
rect 6231 5894 6289 5906
rect 6359 5966 6417 5978
rect 6359 5906 6371 5966
rect 6405 5906 6417 5966
rect 6359 5894 6417 5906
rect 6487 5966 6545 5978
rect 6487 5906 6499 5966
rect 6533 5906 6545 5966
rect 6487 5894 6545 5906
rect 6615 5966 6673 5978
rect 6615 5906 6627 5966
rect 6661 5906 6673 5966
rect 6615 5894 6673 5906
rect 6743 5966 6801 5978
rect 6743 5906 6755 5966
rect 6789 5906 6801 5966
rect 6743 5894 6801 5906
rect 6871 5966 6929 5978
rect 6871 5906 6883 5966
rect 6917 5906 6929 5966
rect 6871 5894 6929 5906
rect 6999 5966 7057 5978
rect 6999 5906 7011 5966
rect 7045 5906 7057 5966
rect 6999 5894 7057 5906
rect 7127 5966 7185 5978
rect 7127 5906 7139 5966
rect 7173 5906 7185 5966
rect 7127 5894 7185 5906
rect 7255 5966 7313 5978
rect 7255 5906 7267 5966
rect 7301 5906 7313 5966
rect 7255 5894 7313 5906
rect 7383 5966 7441 5978
rect 7383 5906 7395 5966
rect 7429 5906 7441 5966
rect 7383 5894 7441 5906
rect 7511 5966 7569 5978
rect 7511 5906 7523 5966
rect 7557 5906 7569 5966
rect 7511 5894 7569 5906
rect 10550 5966 10608 5978
rect 10550 5906 10562 5966
rect 10596 5906 10608 5966
rect 10550 5894 10608 5906
rect 10678 5966 10736 5978
rect 10678 5906 10690 5966
rect 10724 5906 10736 5966
rect 10678 5894 10736 5906
rect 10806 5966 10864 5978
rect 10806 5906 10818 5966
rect 10852 5906 10864 5966
rect 10806 5894 10864 5906
rect 10934 5966 10992 5978
rect 10934 5906 10946 5966
rect 10980 5906 10992 5966
rect 10934 5894 10992 5906
rect 11062 5966 11120 5978
rect 11062 5906 11074 5966
rect 11108 5906 11120 5966
rect 11062 5894 11120 5906
rect 11190 5966 11248 5978
rect 11190 5906 11202 5966
rect 11236 5906 11248 5966
rect 11190 5894 11248 5906
rect 11318 5966 11376 5978
rect 11318 5906 11330 5966
rect 11364 5906 11376 5966
rect 11318 5894 11376 5906
rect 11446 5966 11504 5978
rect 11446 5906 11458 5966
rect 11492 5906 11504 5966
rect 11446 5894 11504 5906
rect 11574 5966 11632 5978
rect 11574 5906 11586 5966
rect 11620 5906 11632 5966
rect 11574 5894 11632 5906
rect 11702 5966 11760 5978
rect 11702 5906 11714 5966
rect 11748 5906 11760 5966
rect 11702 5894 11760 5906
rect 11830 5966 11888 5978
rect 11830 5906 11842 5966
rect 11876 5906 11888 5966
rect 11830 5894 11888 5906
rect 11958 5966 12016 5978
rect 11958 5906 11970 5966
rect 12004 5906 12016 5966
rect 11958 5894 12016 5906
rect 12086 5966 12144 5978
rect 12086 5906 12098 5966
rect 12132 5906 12144 5966
rect 12086 5894 12144 5906
rect 12214 5966 12272 5978
rect 12214 5906 12226 5966
rect 12260 5906 12272 5966
rect 12214 5894 12272 5906
rect 12342 5966 12400 5978
rect 12342 5906 12354 5966
rect 12388 5906 12400 5966
rect 12342 5894 12400 5906
rect 12470 5966 12528 5978
rect 12470 5906 12482 5966
rect 12516 5906 12528 5966
rect 12470 5894 12528 5906
rect 12598 5966 12656 5978
rect 12598 5906 12610 5966
rect 12644 5906 12656 5966
rect 12598 5894 12656 5906
rect 12726 5966 12784 5978
rect 12726 5906 12738 5966
rect 12772 5906 12784 5966
rect 12726 5894 12784 5906
rect 12854 5966 12912 5978
rect 12854 5906 12866 5966
rect 12900 5906 12912 5966
rect 12854 5894 12912 5906
rect 12982 5966 13040 5978
rect 12982 5906 12994 5966
rect 13028 5906 13040 5966
rect 12982 5894 13040 5906
rect 13110 5966 13168 5978
rect 13110 5906 13122 5966
rect 13156 5906 13168 5966
rect 13110 5894 13168 5906
rect 13238 5966 13296 5978
rect 13238 5906 13250 5966
rect 13284 5906 13296 5966
rect 13238 5894 13296 5906
rect 13366 5966 13424 5978
rect 13366 5906 13378 5966
rect 13412 5906 13424 5966
rect 13366 5894 13424 5906
rect 13494 5966 13552 5978
rect 13494 5906 13506 5966
rect 13540 5906 13552 5966
rect 13494 5894 13552 5906
rect 13622 5966 13680 5978
rect 13622 5906 13634 5966
rect 13668 5906 13680 5966
rect 13622 5894 13680 5906
rect 13750 5966 13808 5978
rect 13750 5906 13762 5966
rect 13796 5906 13808 5966
rect 13750 5894 13808 5906
rect 13878 5966 13936 5978
rect 13878 5906 13890 5966
rect 13924 5906 13936 5966
rect 13878 5894 13936 5906
rect 14006 5966 14064 5978
rect 14006 5906 14018 5966
rect 14052 5906 14064 5966
rect 14006 5894 14064 5906
rect 14134 5966 14192 5978
rect 14134 5906 14146 5966
rect 14180 5906 14192 5966
rect 14134 5894 14192 5906
rect 14262 5966 14320 5978
rect 14262 5906 14274 5966
rect 14308 5906 14320 5966
rect 14262 5894 14320 5906
rect 14390 5966 14448 5978
rect 14390 5906 14402 5966
rect 14436 5906 14448 5966
rect 14390 5894 14448 5906
rect 14518 5966 14576 5978
rect 14518 5906 14530 5966
rect 14564 5906 14576 5966
rect 14518 5894 14576 5906
rect 14646 5966 14704 5978
rect 14646 5906 14658 5966
rect 14692 5906 14704 5966
rect 14646 5894 14704 5906
rect 20335 5966 20393 5978
rect 20335 5906 20347 5966
rect 20381 5906 20393 5966
rect 20335 5894 20393 5906
rect 20463 5966 20521 5978
rect 20463 5906 20475 5966
rect 20509 5906 20521 5966
rect 20463 5894 20521 5906
rect 20591 5966 20649 5978
rect 20591 5906 20603 5966
rect 20637 5906 20649 5966
rect 20591 5894 20649 5906
rect 20719 5966 20777 5978
rect 20719 5906 20731 5966
rect 20765 5906 20777 5966
rect 20719 5894 20777 5906
rect 20847 5966 20905 5978
rect 20847 5906 20859 5966
rect 20893 5906 20905 5966
rect 20847 5894 20905 5906
rect 20975 5966 21033 5978
rect 20975 5906 20987 5966
rect 21021 5906 21033 5966
rect 20975 5894 21033 5906
rect 21103 5966 21161 5978
rect 21103 5906 21115 5966
rect 21149 5906 21161 5966
rect 21103 5894 21161 5906
rect 21231 5966 21289 5978
rect 21231 5906 21243 5966
rect 21277 5906 21289 5966
rect 21231 5894 21289 5906
rect 21359 5966 21417 5978
rect 21359 5906 21371 5966
rect 21405 5906 21417 5966
rect 21359 5894 21417 5906
rect 21487 5966 21545 5978
rect 21487 5906 21499 5966
rect 21533 5906 21545 5966
rect 21487 5894 21545 5906
rect 21615 5966 21673 5978
rect 21615 5906 21627 5966
rect 21661 5906 21673 5966
rect 21615 5894 21673 5906
rect 21743 5966 21801 5978
rect 21743 5906 21755 5966
rect 21789 5906 21801 5966
rect 21743 5894 21801 5906
rect 21871 5966 21929 5978
rect 21871 5906 21883 5966
rect 21917 5906 21929 5966
rect 21871 5894 21929 5906
rect 21999 5966 22057 5978
rect 21999 5906 22011 5966
rect 22045 5906 22057 5966
rect 21999 5894 22057 5906
rect 22127 5966 22185 5978
rect 22127 5906 22139 5966
rect 22173 5906 22185 5966
rect 22127 5894 22185 5906
rect 22255 5966 22313 5978
rect 22255 5906 22267 5966
rect 22301 5906 22313 5966
rect 22255 5894 22313 5906
rect 22383 5966 22441 5978
rect 22383 5906 22395 5966
rect 22429 5906 22441 5966
rect 22383 5894 22441 5906
rect 22511 5966 22569 5978
rect 22511 5906 22523 5966
rect 22557 5906 22569 5966
rect 22511 5894 22569 5906
rect 22639 5966 22697 5978
rect 22639 5906 22651 5966
rect 22685 5906 22697 5966
rect 22639 5894 22697 5906
rect 22767 5966 22825 5978
rect 22767 5906 22779 5966
rect 22813 5906 22825 5966
rect 22767 5894 22825 5906
rect 22895 5966 22953 5978
rect 22895 5906 22907 5966
rect 22941 5906 22953 5966
rect 22895 5894 22953 5906
rect 23023 5966 23081 5978
rect 23023 5906 23035 5966
rect 23069 5906 23081 5966
rect 23023 5894 23081 5906
rect 23151 5966 23209 5978
rect 23151 5906 23163 5966
rect 23197 5906 23209 5966
rect 23151 5894 23209 5906
rect 23279 5966 23337 5978
rect 23279 5906 23291 5966
rect 23325 5906 23337 5966
rect 23279 5894 23337 5906
rect 23407 5966 23465 5978
rect 23407 5906 23419 5966
rect 23453 5906 23465 5966
rect 23407 5894 23465 5906
rect 23535 5966 23593 5978
rect 23535 5906 23547 5966
rect 23581 5906 23593 5966
rect 23535 5894 23593 5906
rect 23663 5966 23721 5978
rect 23663 5906 23675 5966
rect 23709 5906 23721 5966
rect 23663 5894 23721 5906
rect 23791 5966 23849 5978
rect 23791 5906 23803 5966
rect 23837 5906 23849 5966
rect 23791 5894 23849 5906
rect 23919 5966 23977 5978
rect 23919 5906 23931 5966
rect 23965 5906 23977 5966
rect 23919 5894 23977 5906
rect 24047 5966 24105 5978
rect 24047 5906 24059 5966
rect 24093 5906 24105 5966
rect 24047 5894 24105 5906
rect 24175 5966 24233 5978
rect 24175 5906 24187 5966
rect 24221 5906 24233 5966
rect 24175 5894 24233 5906
rect 24303 5966 24361 5978
rect 24303 5906 24315 5966
rect 24349 5906 24361 5966
rect 24303 5894 24361 5906
rect 24431 5966 24489 5978
rect 24431 5906 24443 5966
rect 24477 5906 24489 5966
rect 24431 5894 24489 5906
rect 24559 5966 24617 5978
rect 24559 5906 24571 5966
rect 24605 5906 24617 5966
rect 24559 5894 24617 5906
rect 24687 5966 24745 5978
rect 24687 5906 24699 5966
rect 24733 5906 24745 5966
rect 24687 5894 24745 5906
rect 24815 5966 24873 5978
rect 24815 5906 24827 5966
rect 24861 5906 24873 5966
rect 24815 5894 24873 5906
rect 24943 5966 25001 5978
rect 24943 5906 24955 5966
rect 24989 5906 25001 5966
rect 24943 5894 25001 5906
rect 25071 5966 25129 5978
rect 25071 5906 25083 5966
rect 25117 5906 25129 5966
rect 25071 5894 25129 5906
rect 25199 5966 25257 5978
rect 25199 5906 25211 5966
rect 25245 5906 25257 5966
rect 25199 5894 25257 5906
rect 25327 5966 25385 5978
rect 25327 5906 25339 5966
rect 25373 5906 25385 5966
rect 25327 5894 25385 5906
rect 25455 5966 25513 5978
rect 25455 5906 25467 5966
rect 25501 5906 25513 5966
rect 25455 5894 25513 5906
rect 25583 5966 25641 5978
rect 25583 5906 25595 5966
rect 25629 5906 25641 5966
rect 25583 5894 25641 5906
rect 25711 5966 25769 5978
rect 25711 5906 25723 5966
rect 25757 5906 25769 5966
rect 25711 5894 25769 5906
rect 25839 5966 25897 5978
rect 25839 5906 25851 5966
rect 25885 5906 25897 5966
rect 25839 5894 25897 5906
rect 25967 5966 26025 5978
rect 25967 5906 25979 5966
rect 26013 5906 26025 5966
rect 25967 5894 26025 5906
rect 26095 5966 26153 5978
rect 26095 5906 26107 5966
rect 26141 5906 26153 5966
rect 26095 5894 26153 5906
rect 26223 5966 26281 5978
rect 26223 5906 26235 5966
rect 26269 5906 26281 5966
rect 26223 5894 26281 5906
rect 26351 5966 26409 5978
rect 26351 5906 26363 5966
rect 26397 5906 26409 5966
rect 26351 5894 26409 5906
rect 26479 5966 26537 5978
rect 26479 5906 26491 5966
rect 26525 5906 26537 5966
rect 26479 5894 26537 5906
rect 26607 5966 26665 5978
rect 26607 5906 26619 5966
rect 26653 5906 26665 5966
rect 26607 5894 26665 5906
rect 26735 5966 26793 5978
rect 26735 5906 26747 5966
rect 26781 5906 26793 5966
rect 26735 5894 26793 5906
rect 26863 5966 26921 5978
rect 26863 5906 26875 5966
rect 26909 5906 26921 5966
rect 26863 5894 26921 5906
rect 26991 5966 27049 5978
rect 26991 5906 27003 5966
rect 27037 5906 27049 5966
rect 26991 5894 27049 5906
rect 27119 5966 27177 5978
rect 27119 5906 27131 5966
rect 27165 5906 27177 5966
rect 27119 5894 27177 5906
rect 27247 5966 27305 5978
rect 27247 5906 27259 5966
rect 27293 5906 27305 5966
rect 27247 5894 27305 5906
rect 27375 5966 27433 5978
rect 27375 5906 27387 5966
rect 27421 5906 27433 5966
rect 27375 5894 27433 5906
rect 27503 5966 27561 5978
rect 27503 5906 27515 5966
rect 27549 5906 27561 5966
rect 27503 5894 27561 5906
rect 27631 5966 27689 5978
rect 27631 5906 27643 5966
rect 27677 5906 27689 5966
rect 27631 5894 27689 5906
rect 27759 5966 27817 5978
rect 27759 5906 27771 5966
rect 27805 5906 27817 5966
rect 27759 5894 27817 5906
rect 27887 5966 27945 5978
rect 27887 5906 27899 5966
rect 27933 5906 27945 5966
rect 27887 5894 27945 5906
rect 28015 5966 28073 5978
rect 28015 5906 28027 5966
rect 28061 5906 28073 5966
rect 28015 5894 28073 5906
rect 28143 5966 28201 5978
rect 28143 5906 28155 5966
rect 28189 5906 28201 5966
rect 28143 5894 28201 5906
rect 28271 5966 28329 5978
rect 28271 5906 28283 5966
rect 28317 5906 28329 5966
rect 28271 5894 28329 5906
rect 28399 5966 28457 5978
rect 28399 5906 28411 5966
rect 28445 5906 28457 5966
rect 28399 5894 28457 5906
rect 28527 5966 28585 5978
rect 28527 5906 28539 5966
rect 28573 5906 28585 5966
rect 28527 5894 28585 5906
rect -329 5278 -271 5290
rect -329 5218 -317 5278
rect -283 5218 -271 5278
rect -329 5206 -271 5218
rect -201 5278 -143 5290
rect -201 5218 -189 5278
rect -155 5218 -143 5278
rect -201 5206 -143 5218
rect 599 5278 657 5290
rect 599 5218 611 5278
rect 645 5218 657 5278
rect 599 5206 657 5218
rect 727 5278 785 5290
rect 727 5218 739 5278
rect 773 5218 785 5278
rect 727 5206 785 5218
rect 855 5278 913 5290
rect 855 5218 867 5278
rect 901 5218 913 5278
rect 855 5206 913 5218
rect 1863 5278 1921 5290
rect 1863 5218 1875 5278
rect 1909 5218 1921 5278
rect 1863 5206 1921 5218
rect 1991 5278 2049 5290
rect 1991 5218 2003 5278
rect 2037 5218 2049 5278
rect 1991 5206 2049 5218
rect 2119 5278 2177 5290
rect 2119 5218 2131 5278
rect 2165 5218 2177 5278
rect 2119 5206 2177 5218
rect 2247 5278 2305 5290
rect 2247 5218 2259 5278
rect 2293 5218 2305 5278
rect 2247 5206 2305 5218
rect 2375 5278 2433 5290
rect 2375 5218 2387 5278
rect 2421 5218 2433 5278
rect 2375 5206 2433 5218
rect 3482 5278 3540 5290
rect 3482 5218 3494 5278
rect 3528 5218 3540 5278
rect 3482 5206 3540 5218
rect 3610 5278 3668 5290
rect 3610 5218 3622 5278
rect 3656 5218 3668 5278
rect 3610 5206 3668 5218
rect 3738 5278 3796 5290
rect 3738 5218 3750 5278
rect 3784 5218 3796 5278
rect 3738 5206 3796 5218
rect 3866 5278 3924 5290
rect 3866 5218 3878 5278
rect 3912 5218 3924 5278
rect 3866 5206 3924 5218
rect 3994 5278 4052 5290
rect 3994 5218 4006 5278
rect 4040 5218 4052 5278
rect 3994 5206 4052 5218
rect 4122 5278 4180 5290
rect 4122 5218 4134 5278
rect 4168 5218 4180 5278
rect 4122 5206 4180 5218
rect 4250 5278 4308 5290
rect 4250 5218 4262 5278
rect 4296 5218 4308 5278
rect 4250 5206 4308 5218
rect 4378 5278 4436 5290
rect 4378 5218 4390 5278
rect 4424 5218 4436 5278
rect 4378 5206 4436 5218
rect 4506 5278 4564 5290
rect 4506 5218 4518 5278
rect 4552 5218 4564 5278
rect 4506 5206 4564 5218
rect 8047 5278 8105 5290
rect 8047 5218 8059 5278
rect 8093 5218 8105 5278
rect 8047 5206 8105 5218
rect 8175 5278 8233 5290
rect 8175 5218 8187 5278
rect 8221 5218 8233 5278
rect 8175 5206 8233 5218
rect 8303 5278 8361 5290
rect 8303 5218 8315 5278
rect 8349 5218 8361 5278
rect 8303 5206 8361 5218
rect 8431 5278 8489 5290
rect 8431 5218 8443 5278
rect 8477 5218 8489 5278
rect 8431 5206 8489 5218
rect 8559 5278 8617 5290
rect 8559 5218 8571 5278
rect 8605 5218 8617 5278
rect 8559 5206 8617 5218
rect 8687 5278 8745 5290
rect 8687 5218 8699 5278
rect 8733 5218 8745 5278
rect 8687 5206 8745 5218
rect 8815 5278 8873 5290
rect 8815 5218 8827 5278
rect 8861 5218 8873 5278
rect 8815 5206 8873 5218
rect 8943 5278 9001 5290
rect 8943 5218 8955 5278
rect 8989 5218 9001 5278
rect 8943 5206 9001 5218
rect 9071 5278 9129 5290
rect 9071 5218 9083 5278
rect 9117 5218 9129 5278
rect 9071 5206 9129 5218
rect 9199 5278 9257 5290
rect 9199 5218 9211 5278
rect 9245 5218 9257 5278
rect 9199 5206 9257 5218
rect 9327 5278 9385 5290
rect 9327 5218 9339 5278
rect 9373 5218 9385 5278
rect 9327 5206 9385 5218
rect 9455 5278 9513 5290
rect 9455 5218 9467 5278
rect 9501 5218 9513 5278
rect 9455 5206 9513 5218
rect 9583 5278 9641 5290
rect 9583 5218 9595 5278
rect 9629 5218 9641 5278
rect 9583 5206 9641 5218
rect 9711 5278 9769 5290
rect 9711 5218 9723 5278
rect 9757 5218 9769 5278
rect 9711 5206 9769 5218
rect 9839 5278 9897 5290
rect 9839 5218 9851 5278
rect 9885 5218 9897 5278
rect 9839 5206 9897 5218
rect 9967 5278 10025 5290
rect 9967 5218 9979 5278
rect 10013 5218 10025 5278
rect 9967 5206 10025 5218
rect 10095 5278 10153 5290
rect 10095 5218 10107 5278
rect 10141 5218 10153 5278
rect 10095 5206 10153 5218
rect 15205 5278 15263 5290
rect 15205 5218 15217 5278
rect 15251 5218 15263 5278
rect 15205 5206 15263 5218
rect 15333 5278 15391 5290
rect 15333 5218 15345 5278
rect 15379 5218 15391 5278
rect 15333 5206 15391 5218
rect 15461 5278 15519 5290
rect 15461 5218 15473 5278
rect 15507 5218 15519 5278
rect 15461 5206 15519 5218
rect 15589 5278 15647 5290
rect 15589 5218 15601 5278
rect 15635 5218 15647 5278
rect 15589 5206 15647 5218
rect 15717 5278 15775 5290
rect 15717 5218 15729 5278
rect 15763 5218 15775 5278
rect 15717 5206 15775 5218
rect 15845 5278 15903 5290
rect 15845 5218 15857 5278
rect 15891 5218 15903 5278
rect 15845 5206 15903 5218
rect 15973 5278 16031 5290
rect 15973 5218 15985 5278
rect 16019 5218 16031 5278
rect 15973 5206 16031 5218
rect 16101 5278 16159 5290
rect 16101 5218 16113 5278
rect 16147 5218 16159 5278
rect 16101 5206 16159 5218
rect 16229 5278 16287 5290
rect 16229 5218 16241 5278
rect 16275 5218 16287 5278
rect 16229 5206 16287 5218
rect 16357 5278 16415 5290
rect 16357 5218 16369 5278
rect 16403 5218 16415 5278
rect 16357 5206 16415 5218
rect 16485 5278 16543 5290
rect 16485 5218 16497 5278
rect 16531 5218 16543 5278
rect 16485 5206 16543 5218
rect 16613 5278 16671 5290
rect 16613 5218 16625 5278
rect 16659 5218 16671 5278
rect 16613 5206 16671 5218
rect 16741 5278 16799 5290
rect 16741 5218 16753 5278
rect 16787 5218 16799 5278
rect 16741 5206 16799 5218
rect 16869 5278 16927 5290
rect 16869 5218 16881 5278
rect 16915 5218 16927 5278
rect 16869 5206 16927 5218
rect 16997 5278 17055 5290
rect 16997 5218 17009 5278
rect 17043 5218 17055 5278
rect 16997 5206 17055 5218
rect 17125 5278 17183 5290
rect 17125 5218 17137 5278
rect 17171 5218 17183 5278
rect 17125 5206 17183 5218
rect 17253 5278 17311 5290
rect 17253 5218 17265 5278
rect 17299 5218 17311 5278
rect 17253 5206 17311 5218
rect 17381 5278 17439 5290
rect 17381 5218 17393 5278
rect 17427 5218 17439 5278
rect 17381 5206 17439 5218
rect 17509 5278 17567 5290
rect 17509 5218 17521 5278
rect 17555 5218 17567 5278
rect 17509 5206 17567 5218
rect 17637 5278 17695 5290
rect 17637 5218 17649 5278
rect 17683 5218 17695 5278
rect 17637 5206 17695 5218
rect 17765 5278 17823 5290
rect 17765 5218 17777 5278
rect 17811 5218 17823 5278
rect 17765 5206 17823 5218
rect 17893 5278 17951 5290
rect 17893 5218 17905 5278
rect 17939 5218 17951 5278
rect 17893 5206 17951 5218
rect 18021 5278 18079 5290
rect 18021 5218 18033 5278
rect 18067 5218 18079 5278
rect 18021 5206 18079 5218
rect 18149 5278 18207 5290
rect 18149 5218 18161 5278
rect 18195 5218 18207 5278
rect 18149 5206 18207 5218
rect 18277 5278 18335 5290
rect 18277 5218 18289 5278
rect 18323 5218 18335 5278
rect 18277 5206 18335 5218
rect 18405 5278 18463 5290
rect 18405 5218 18417 5278
rect 18451 5218 18463 5278
rect 18405 5206 18463 5218
rect 18533 5278 18591 5290
rect 18533 5218 18545 5278
rect 18579 5218 18591 5278
rect 18533 5206 18591 5218
rect 18661 5278 18719 5290
rect 18661 5218 18673 5278
rect 18707 5218 18719 5278
rect 18661 5206 18719 5218
rect 18789 5278 18847 5290
rect 18789 5218 18801 5278
rect 18835 5218 18847 5278
rect 18789 5206 18847 5218
rect 18917 5278 18975 5290
rect 18917 5218 18929 5278
rect 18963 5218 18975 5278
rect 18917 5206 18975 5218
rect 19045 5278 19103 5290
rect 19045 5218 19057 5278
rect 19091 5218 19103 5278
rect 19045 5206 19103 5218
rect 19173 5278 19231 5290
rect 19173 5218 19185 5278
rect 19219 5218 19231 5278
rect 19173 5206 19231 5218
rect 19301 5278 19359 5290
rect 19301 5218 19313 5278
rect 19347 5218 19359 5278
rect 19301 5206 19359 5218
rect 20259 5278 20317 5290
rect 20259 5218 20271 5278
rect 20305 5218 20317 5278
rect 20259 5206 20317 5218
rect 20387 5278 20445 5290
rect 20387 5218 20399 5278
rect 20433 5218 20445 5278
rect 20387 5206 20445 5218
rect 20515 5278 20573 5290
rect 20515 5218 20527 5278
rect 20561 5218 20573 5278
rect 20515 5206 20573 5218
rect 20643 5278 20701 5290
rect 20643 5218 20655 5278
rect 20689 5218 20701 5278
rect 20643 5206 20701 5218
rect 20771 5278 20829 5290
rect 20771 5218 20783 5278
rect 20817 5218 20829 5278
rect 20771 5206 20829 5218
rect 20899 5278 20957 5290
rect 20899 5218 20911 5278
rect 20945 5218 20957 5278
rect 20899 5206 20957 5218
rect 21027 5278 21085 5290
rect 21027 5218 21039 5278
rect 21073 5218 21085 5278
rect 21027 5206 21085 5218
rect 21155 5278 21213 5290
rect 21155 5218 21167 5278
rect 21201 5218 21213 5278
rect 21155 5206 21213 5218
rect 21283 5278 21341 5290
rect 21283 5218 21295 5278
rect 21329 5218 21341 5278
rect 21283 5206 21341 5218
rect 21411 5278 21469 5290
rect 21411 5218 21423 5278
rect 21457 5218 21469 5278
rect 21411 5206 21469 5218
rect 21539 5278 21597 5290
rect 21539 5218 21551 5278
rect 21585 5218 21597 5278
rect 21539 5206 21597 5218
rect 21667 5278 21725 5290
rect 21667 5218 21679 5278
rect 21713 5218 21725 5278
rect 21667 5206 21725 5218
rect 21795 5278 21853 5290
rect 21795 5218 21807 5278
rect 21841 5218 21853 5278
rect 21795 5206 21853 5218
rect 21923 5278 21981 5290
rect 21923 5218 21935 5278
rect 21969 5218 21981 5278
rect 21923 5206 21981 5218
rect 22051 5278 22109 5290
rect 22051 5218 22063 5278
rect 22097 5218 22109 5278
rect 22051 5206 22109 5218
rect 22179 5278 22237 5290
rect 22179 5218 22191 5278
rect 22225 5218 22237 5278
rect 22179 5206 22237 5218
rect 22307 5278 22365 5290
rect 22307 5218 22319 5278
rect 22353 5218 22365 5278
rect 22307 5206 22365 5218
rect 22435 5278 22493 5290
rect 22435 5218 22447 5278
rect 22481 5218 22493 5278
rect 22435 5206 22493 5218
rect 22563 5278 22621 5290
rect 22563 5218 22575 5278
rect 22609 5218 22621 5278
rect 22563 5206 22621 5218
rect 22691 5278 22749 5290
rect 22691 5218 22703 5278
rect 22737 5218 22749 5278
rect 22691 5206 22749 5218
rect 22819 5278 22877 5290
rect 22819 5218 22831 5278
rect 22865 5218 22877 5278
rect 22819 5206 22877 5218
rect 22947 5278 23005 5290
rect 22947 5218 22959 5278
rect 22993 5218 23005 5278
rect 22947 5206 23005 5218
rect 23075 5278 23133 5290
rect 23075 5218 23087 5278
rect 23121 5218 23133 5278
rect 23075 5206 23133 5218
rect 23203 5278 23261 5290
rect 23203 5218 23215 5278
rect 23249 5218 23261 5278
rect 23203 5206 23261 5218
rect 23331 5278 23389 5290
rect 23331 5218 23343 5278
rect 23377 5218 23389 5278
rect 23331 5206 23389 5218
rect 23459 5278 23517 5290
rect 23459 5218 23471 5278
rect 23505 5218 23517 5278
rect 23459 5206 23517 5218
rect 23587 5278 23645 5290
rect 23587 5218 23599 5278
rect 23633 5218 23645 5278
rect 23587 5206 23645 5218
rect 23715 5278 23773 5290
rect 23715 5218 23727 5278
rect 23761 5218 23773 5278
rect 23715 5206 23773 5218
rect 23843 5278 23901 5290
rect 23843 5218 23855 5278
rect 23889 5218 23901 5278
rect 23843 5206 23901 5218
rect 23971 5278 24029 5290
rect 23971 5218 23983 5278
rect 24017 5218 24029 5278
rect 23971 5206 24029 5218
rect 24099 5278 24157 5290
rect 24099 5218 24111 5278
rect 24145 5218 24157 5278
rect 24099 5206 24157 5218
rect 24227 5278 24285 5290
rect 24227 5218 24239 5278
rect 24273 5218 24285 5278
rect 24227 5206 24285 5218
rect 24355 5278 24413 5290
rect 24355 5218 24367 5278
rect 24401 5218 24413 5278
rect 24355 5206 24413 5218
rect 24483 5278 24541 5290
rect 24483 5218 24495 5278
rect 24529 5218 24541 5278
rect 24483 5206 24541 5218
rect 24611 5278 24669 5290
rect 24611 5218 24623 5278
rect 24657 5218 24669 5278
rect 24611 5206 24669 5218
rect 24739 5278 24797 5290
rect 24739 5218 24751 5278
rect 24785 5218 24797 5278
rect 24739 5206 24797 5218
rect 24867 5278 24925 5290
rect 24867 5218 24879 5278
rect 24913 5218 24925 5278
rect 24867 5206 24925 5218
rect 24995 5278 25053 5290
rect 24995 5218 25007 5278
rect 25041 5218 25053 5278
rect 24995 5206 25053 5218
rect 25123 5278 25181 5290
rect 25123 5218 25135 5278
rect 25169 5218 25181 5278
rect 25123 5206 25181 5218
rect 25251 5278 25309 5290
rect 25251 5218 25263 5278
rect 25297 5218 25309 5278
rect 25251 5206 25309 5218
rect 25379 5278 25437 5290
rect 25379 5218 25391 5278
rect 25425 5218 25437 5278
rect 25379 5206 25437 5218
rect 25507 5278 25565 5290
rect 25507 5218 25519 5278
rect 25553 5218 25565 5278
rect 25507 5206 25565 5218
rect 25635 5278 25693 5290
rect 25635 5218 25647 5278
rect 25681 5218 25693 5278
rect 25635 5206 25693 5218
rect 25763 5278 25821 5290
rect 25763 5218 25775 5278
rect 25809 5218 25821 5278
rect 25763 5206 25821 5218
rect 25891 5278 25949 5290
rect 25891 5218 25903 5278
rect 25937 5218 25949 5278
rect 25891 5206 25949 5218
rect 26019 5278 26077 5290
rect 26019 5218 26031 5278
rect 26065 5218 26077 5278
rect 26019 5206 26077 5218
rect 26147 5278 26205 5290
rect 26147 5218 26159 5278
rect 26193 5218 26205 5278
rect 26147 5206 26205 5218
rect 26275 5278 26333 5290
rect 26275 5218 26287 5278
rect 26321 5218 26333 5278
rect 26275 5206 26333 5218
rect 26403 5278 26461 5290
rect 26403 5218 26415 5278
rect 26449 5218 26461 5278
rect 26403 5206 26461 5218
rect 26531 5278 26589 5290
rect 26531 5218 26543 5278
rect 26577 5218 26589 5278
rect 26531 5206 26589 5218
rect 26659 5278 26717 5290
rect 26659 5218 26671 5278
rect 26705 5218 26717 5278
rect 26659 5206 26717 5218
rect 26787 5278 26845 5290
rect 26787 5218 26799 5278
rect 26833 5218 26845 5278
rect 26787 5206 26845 5218
rect 26915 5278 26973 5290
rect 26915 5218 26927 5278
rect 26961 5218 26973 5278
rect 26915 5206 26973 5218
rect 27043 5278 27101 5290
rect 27043 5218 27055 5278
rect 27089 5218 27101 5278
rect 27043 5206 27101 5218
rect 27171 5278 27229 5290
rect 27171 5218 27183 5278
rect 27217 5218 27229 5278
rect 27171 5206 27229 5218
rect 27299 5278 27357 5290
rect 27299 5218 27311 5278
rect 27345 5218 27357 5278
rect 27299 5206 27357 5218
rect 27427 5278 27485 5290
rect 27427 5218 27439 5278
rect 27473 5218 27485 5278
rect 27427 5206 27485 5218
rect 27555 5278 27613 5290
rect 27555 5218 27567 5278
rect 27601 5218 27613 5278
rect 27555 5206 27613 5218
rect 27683 5278 27741 5290
rect 27683 5218 27695 5278
rect 27729 5218 27741 5278
rect 27683 5206 27741 5218
rect 27811 5278 27869 5290
rect 27811 5218 27823 5278
rect 27857 5218 27869 5278
rect 27811 5206 27869 5218
rect 27939 5278 27997 5290
rect 27939 5218 27951 5278
rect 27985 5218 27997 5278
rect 27939 5206 27997 5218
rect 28067 5278 28125 5290
rect 28067 5218 28079 5278
rect 28113 5218 28125 5278
rect 28067 5206 28125 5218
rect 28195 5278 28253 5290
rect 28195 5218 28207 5278
rect 28241 5218 28253 5278
rect 28195 5206 28253 5218
rect 28323 5278 28381 5290
rect 28323 5218 28335 5278
rect 28369 5218 28381 5278
rect 28323 5206 28381 5218
rect 28451 5278 28509 5290
rect 28451 5218 28463 5278
rect 28497 5218 28509 5278
rect 28451 5206 28509 5218
<< pdiff >>
rect -307 6266 -249 6278
rect -307 6122 -295 6266
rect -261 6122 -249 6266
rect -307 6110 -249 6122
rect -179 6266 -121 6278
rect -179 6122 -167 6266
rect -133 6122 -121 6266
rect -179 6110 -121 6122
rect 470 6266 528 6278
rect 470 6122 482 6266
rect 516 6122 528 6266
rect 470 6110 528 6122
rect 598 6266 656 6278
rect 598 6122 610 6266
rect 644 6122 656 6266
rect 598 6110 656 6122
rect 726 6266 784 6278
rect 726 6122 738 6266
rect 772 6122 784 6266
rect 726 6110 784 6122
rect 1379 6266 1437 6278
rect 1379 6122 1391 6266
rect 1425 6122 1437 6266
rect 1379 6110 1437 6122
rect 1507 6266 1565 6278
rect 1507 6122 1519 6266
rect 1553 6122 1565 6266
rect 1507 6110 1565 6122
rect 1635 6266 1693 6278
rect 1635 6122 1647 6266
rect 1681 6122 1693 6266
rect 1635 6110 1693 6122
rect 1763 6266 1821 6278
rect 1763 6122 1775 6266
rect 1809 6122 1821 6266
rect 1763 6110 1821 6122
rect 1891 6266 1949 6278
rect 1891 6122 1903 6266
rect 1937 6122 1949 6266
rect 1891 6110 1949 6122
rect 2912 6266 2970 6278
rect 2912 6122 2924 6266
rect 2958 6122 2970 6266
rect 2912 6110 2970 6122
rect 3040 6266 3098 6278
rect 3040 6122 3052 6266
rect 3086 6122 3098 6266
rect 3040 6110 3098 6122
rect 3168 6266 3226 6278
rect 3168 6122 3180 6266
rect 3214 6122 3226 6266
rect 3168 6110 3226 6122
rect 3296 6266 3354 6278
rect 3296 6122 3308 6266
rect 3342 6122 3354 6266
rect 3296 6110 3354 6122
rect 3424 6266 3482 6278
rect 3424 6122 3436 6266
rect 3470 6122 3482 6266
rect 3424 6110 3482 6122
rect 3552 6266 3610 6278
rect 3552 6122 3564 6266
rect 3598 6122 3610 6266
rect 3552 6110 3610 6122
rect 3680 6266 3738 6278
rect 3680 6122 3692 6266
rect 3726 6122 3738 6266
rect 3680 6110 3738 6122
rect 3808 6266 3866 6278
rect 3808 6122 3820 6266
rect 3854 6122 3866 6266
rect 3808 6110 3866 6122
rect 3936 6266 3994 6278
rect 3936 6122 3948 6266
rect 3982 6122 3994 6266
rect 3936 6110 3994 6122
rect 5463 6266 5521 6278
rect 5463 6122 5475 6266
rect 5509 6122 5521 6266
rect 5463 6110 5521 6122
rect 5591 6266 5649 6278
rect 5591 6122 5603 6266
rect 5637 6122 5649 6266
rect 5591 6110 5649 6122
rect 5719 6266 5777 6278
rect 5719 6122 5731 6266
rect 5765 6122 5777 6266
rect 5719 6110 5777 6122
rect 5847 6266 5905 6278
rect 5847 6122 5859 6266
rect 5893 6122 5905 6266
rect 5847 6110 5905 6122
rect 5975 6266 6033 6278
rect 5975 6122 5987 6266
rect 6021 6122 6033 6266
rect 5975 6110 6033 6122
rect 6103 6266 6161 6278
rect 6103 6122 6115 6266
rect 6149 6122 6161 6266
rect 6103 6110 6161 6122
rect 6231 6266 6289 6278
rect 6231 6122 6243 6266
rect 6277 6122 6289 6266
rect 6231 6110 6289 6122
rect 6359 6266 6417 6278
rect 6359 6122 6371 6266
rect 6405 6122 6417 6266
rect 6359 6110 6417 6122
rect 6487 6266 6545 6278
rect 6487 6122 6499 6266
rect 6533 6122 6545 6266
rect 6487 6110 6545 6122
rect 6615 6266 6673 6278
rect 6615 6122 6627 6266
rect 6661 6122 6673 6266
rect 6615 6110 6673 6122
rect 6743 6266 6801 6278
rect 6743 6122 6755 6266
rect 6789 6122 6801 6266
rect 6743 6110 6801 6122
rect 6871 6266 6929 6278
rect 6871 6122 6883 6266
rect 6917 6122 6929 6266
rect 6871 6110 6929 6122
rect 6999 6266 7057 6278
rect 6999 6122 7011 6266
rect 7045 6122 7057 6266
rect 6999 6110 7057 6122
rect 7127 6266 7185 6278
rect 7127 6122 7139 6266
rect 7173 6122 7185 6266
rect 7127 6110 7185 6122
rect 7255 6266 7313 6278
rect 7255 6122 7267 6266
rect 7301 6122 7313 6266
rect 7255 6110 7313 6122
rect 7383 6266 7441 6278
rect 7383 6122 7395 6266
rect 7429 6122 7441 6266
rect 7383 6110 7441 6122
rect 7511 6266 7569 6278
rect 7511 6122 7523 6266
rect 7557 6122 7569 6266
rect 7511 6110 7569 6122
rect 10550 6266 10608 6278
rect 10550 6122 10562 6266
rect 10596 6122 10608 6266
rect 10550 6110 10608 6122
rect 10678 6266 10736 6278
rect 10678 6122 10690 6266
rect 10724 6122 10736 6266
rect 10678 6110 10736 6122
rect 10806 6266 10864 6278
rect 10806 6122 10818 6266
rect 10852 6122 10864 6266
rect 10806 6110 10864 6122
rect 10934 6266 10992 6278
rect 10934 6122 10946 6266
rect 10980 6122 10992 6266
rect 10934 6110 10992 6122
rect 11062 6266 11120 6278
rect 11062 6122 11074 6266
rect 11108 6122 11120 6266
rect 11062 6110 11120 6122
rect 11190 6266 11248 6278
rect 11190 6122 11202 6266
rect 11236 6122 11248 6266
rect 11190 6110 11248 6122
rect 11318 6266 11376 6278
rect 11318 6122 11330 6266
rect 11364 6122 11376 6266
rect 11318 6110 11376 6122
rect 11446 6266 11504 6278
rect 11446 6122 11458 6266
rect 11492 6122 11504 6266
rect 11446 6110 11504 6122
rect 11574 6266 11632 6278
rect 11574 6122 11586 6266
rect 11620 6122 11632 6266
rect 11574 6110 11632 6122
rect 11702 6266 11760 6278
rect 11702 6122 11714 6266
rect 11748 6122 11760 6266
rect 11702 6110 11760 6122
rect 11830 6266 11888 6278
rect 11830 6122 11842 6266
rect 11876 6122 11888 6266
rect 11830 6110 11888 6122
rect 11958 6266 12016 6278
rect 11958 6122 11970 6266
rect 12004 6122 12016 6266
rect 11958 6110 12016 6122
rect 12086 6266 12144 6278
rect 12086 6122 12098 6266
rect 12132 6122 12144 6266
rect 12086 6110 12144 6122
rect 12214 6266 12272 6278
rect 12214 6122 12226 6266
rect 12260 6122 12272 6266
rect 12214 6110 12272 6122
rect 12342 6266 12400 6278
rect 12342 6122 12354 6266
rect 12388 6122 12400 6266
rect 12342 6110 12400 6122
rect 12470 6266 12528 6278
rect 12470 6122 12482 6266
rect 12516 6122 12528 6266
rect 12470 6110 12528 6122
rect 12598 6266 12656 6278
rect 12598 6122 12610 6266
rect 12644 6122 12656 6266
rect 12598 6110 12656 6122
rect 12726 6266 12784 6278
rect 12726 6122 12738 6266
rect 12772 6122 12784 6266
rect 12726 6110 12784 6122
rect 12854 6266 12912 6278
rect 12854 6122 12866 6266
rect 12900 6122 12912 6266
rect 12854 6110 12912 6122
rect 12982 6266 13040 6278
rect 12982 6122 12994 6266
rect 13028 6122 13040 6266
rect 12982 6110 13040 6122
rect 13110 6266 13168 6278
rect 13110 6122 13122 6266
rect 13156 6122 13168 6266
rect 13110 6110 13168 6122
rect 13238 6266 13296 6278
rect 13238 6122 13250 6266
rect 13284 6122 13296 6266
rect 13238 6110 13296 6122
rect 13366 6266 13424 6278
rect 13366 6122 13378 6266
rect 13412 6122 13424 6266
rect 13366 6110 13424 6122
rect 13494 6266 13552 6278
rect 13494 6122 13506 6266
rect 13540 6122 13552 6266
rect 13494 6110 13552 6122
rect 13622 6266 13680 6278
rect 13622 6122 13634 6266
rect 13668 6122 13680 6266
rect 13622 6110 13680 6122
rect 13750 6266 13808 6278
rect 13750 6122 13762 6266
rect 13796 6122 13808 6266
rect 13750 6110 13808 6122
rect 13878 6266 13936 6278
rect 13878 6122 13890 6266
rect 13924 6122 13936 6266
rect 13878 6110 13936 6122
rect 14006 6266 14064 6278
rect 14006 6122 14018 6266
rect 14052 6122 14064 6266
rect 14006 6110 14064 6122
rect 14134 6266 14192 6278
rect 14134 6122 14146 6266
rect 14180 6122 14192 6266
rect 14134 6110 14192 6122
rect 14262 6266 14320 6278
rect 14262 6122 14274 6266
rect 14308 6122 14320 6266
rect 14262 6110 14320 6122
rect 14390 6266 14448 6278
rect 14390 6122 14402 6266
rect 14436 6122 14448 6266
rect 14390 6110 14448 6122
rect 14518 6266 14576 6278
rect 14518 6122 14530 6266
rect 14564 6122 14576 6266
rect 14518 6110 14576 6122
rect 14646 6266 14704 6278
rect 14646 6122 14658 6266
rect 14692 6122 14704 6266
rect 14646 6110 14704 6122
rect 20335 6266 20393 6278
rect 20335 6122 20347 6266
rect 20381 6122 20393 6266
rect 20335 6110 20393 6122
rect 20463 6266 20521 6278
rect 20463 6122 20475 6266
rect 20509 6122 20521 6266
rect 20463 6110 20521 6122
rect 20591 6266 20649 6278
rect 20591 6122 20603 6266
rect 20637 6122 20649 6266
rect 20591 6110 20649 6122
rect 20719 6266 20777 6278
rect 20719 6122 20731 6266
rect 20765 6122 20777 6266
rect 20719 6110 20777 6122
rect 20847 6266 20905 6278
rect 20847 6122 20859 6266
rect 20893 6122 20905 6266
rect 20847 6110 20905 6122
rect 20975 6266 21033 6278
rect 20975 6122 20987 6266
rect 21021 6122 21033 6266
rect 20975 6110 21033 6122
rect 21103 6266 21161 6278
rect 21103 6122 21115 6266
rect 21149 6122 21161 6266
rect 21103 6110 21161 6122
rect 21231 6266 21289 6278
rect 21231 6122 21243 6266
rect 21277 6122 21289 6266
rect 21231 6110 21289 6122
rect 21359 6266 21417 6278
rect 21359 6122 21371 6266
rect 21405 6122 21417 6266
rect 21359 6110 21417 6122
rect 21487 6266 21545 6278
rect 21487 6122 21499 6266
rect 21533 6122 21545 6266
rect 21487 6110 21545 6122
rect 21615 6266 21673 6278
rect 21615 6122 21627 6266
rect 21661 6122 21673 6266
rect 21615 6110 21673 6122
rect 21743 6266 21801 6278
rect 21743 6122 21755 6266
rect 21789 6122 21801 6266
rect 21743 6110 21801 6122
rect 21871 6266 21929 6278
rect 21871 6122 21883 6266
rect 21917 6122 21929 6266
rect 21871 6110 21929 6122
rect 21999 6266 22057 6278
rect 21999 6122 22011 6266
rect 22045 6122 22057 6266
rect 21999 6110 22057 6122
rect 22127 6266 22185 6278
rect 22127 6122 22139 6266
rect 22173 6122 22185 6266
rect 22127 6110 22185 6122
rect 22255 6266 22313 6278
rect 22255 6122 22267 6266
rect 22301 6122 22313 6266
rect 22255 6110 22313 6122
rect 22383 6266 22441 6278
rect 22383 6122 22395 6266
rect 22429 6122 22441 6266
rect 22383 6110 22441 6122
rect 22511 6266 22569 6278
rect 22511 6122 22523 6266
rect 22557 6122 22569 6266
rect 22511 6110 22569 6122
rect 22639 6266 22697 6278
rect 22639 6122 22651 6266
rect 22685 6122 22697 6266
rect 22639 6110 22697 6122
rect 22767 6266 22825 6278
rect 22767 6122 22779 6266
rect 22813 6122 22825 6266
rect 22767 6110 22825 6122
rect 22895 6266 22953 6278
rect 22895 6122 22907 6266
rect 22941 6122 22953 6266
rect 22895 6110 22953 6122
rect 23023 6266 23081 6278
rect 23023 6122 23035 6266
rect 23069 6122 23081 6266
rect 23023 6110 23081 6122
rect 23151 6266 23209 6278
rect 23151 6122 23163 6266
rect 23197 6122 23209 6266
rect 23151 6110 23209 6122
rect 23279 6266 23337 6278
rect 23279 6122 23291 6266
rect 23325 6122 23337 6266
rect 23279 6110 23337 6122
rect 23407 6266 23465 6278
rect 23407 6122 23419 6266
rect 23453 6122 23465 6266
rect 23407 6110 23465 6122
rect 23535 6266 23593 6278
rect 23535 6122 23547 6266
rect 23581 6122 23593 6266
rect 23535 6110 23593 6122
rect 23663 6266 23721 6278
rect 23663 6122 23675 6266
rect 23709 6122 23721 6266
rect 23663 6110 23721 6122
rect 23791 6266 23849 6278
rect 23791 6122 23803 6266
rect 23837 6122 23849 6266
rect 23791 6110 23849 6122
rect 23919 6266 23977 6278
rect 23919 6122 23931 6266
rect 23965 6122 23977 6266
rect 23919 6110 23977 6122
rect 24047 6266 24105 6278
rect 24047 6122 24059 6266
rect 24093 6122 24105 6266
rect 24047 6110 24105 6122
rect 24175 6266 24233 6278
rect 24175 6122 24187 6266
rect 24221 6122 24233 6266
rect 24175 6110 24233 6122
rect 24303 6266 24361 6278
rect 24303 6122 24315 6266
rect 24349 6122 24361 6266
rect 24303 6110 24361 6122
rect 24431 6266 24489 6278
rect 24431 6122 24443 6266
rect 24477 6122 24489 6266
rect 24431 6110 24489 6122
rect 24559 6266 24617 6278
rect 24559 6122 24571 6266
rect 24605 6122 24617 6266
rect 24559 6110 24617 6122
rect 24687 6266 24745 6278
rect 24687 6122 24699 6266
rect 24733 6122 24745 6266
rect 24687 6110 24745 6122
rect 24815 6266 24873 6278
rect 24815 6122 24827 6266
rect 24861 6122 24873 6266
rect 24815 6110 24873 6122
rect 24943 6266 25001 6278
rect 24943 6122 24955 6266
rect 24989 6122 25001 6266
rect 24943 6110 25001 6122
rect 25071 6266 25129 6278
rect 25071 6122 25083 6266
rect 25117 6122 25129 6266
rect 25071 6110 25129 6122
rect 25199 6266 25257 6278
rect 25199 6122 25211 6266
rect 25245 6122 25257 6266
rect 25199 6110 25257 6122
rect 25327 6266 25385 6278
rect 25327 6122 25339 6266
rect 25373 6122 25385 6266
rect 25327 6110 25385 6122
rect 25455 6266 25513 6278
rect 25455 6122 25467 6266
rect 25501 6122 25513 6266
rect 25455 6110 25513 6122
rect 25583 6266 25641 6278
rect 25583 6122 25595 6266
rect 25629 6122 25641 6266
rect 25583 6110 25641 6122
rect 25711 6266 25769 6278
rect 25711 6122 25723 6266
rect 25757 6122 25769 6266
rect 25711 6110 25769 6122
rect 25839 6266 25897 6278
rect 25839 6122 25851 6266
rect 25885 6122 25897 6266
rect 25839 6110 25897 6122
rect 25967 6266 26025 6278
rect 25967 6122 25979 6266
rect 26013 6122 26025 6266
rect 25967 6110 26025 6122
rect 26095 6266 26153 6278
rect 26095 6122 26107 6266
rect 26141 6122 26153 6266
rect 26095 6110 26153 6122
rect 26223 6266 26281 6278
rect 26223 6122 26235 6266
rect 26269 6122 26281 6266
rect 26223 6110 26281 6122
rect 26351 6266 26409 6278
rect 26351 6122 26363 6266
rect 26397 6122 26409 6266
rect 26351 6110 26409 6122
rect 26479 6266 26537 6278
rect 26479 6122 26491 6266
rect 26525 6122 26537 6266
rect 26479 6110 26537 6122
rect 26607 6266 26665 6278
rect 26607 6122 26619 6266
rect 26653 6122 26665 6266
rect 26607 6110 26665 6122
rect 26735 6266 26793 6278
rect 26735 6122 26747 6266
rect 26781 6122 26793 6266
rect 26735 6110 26793 6122
rect 26863 6266 26921 6278
rect 26863 6122 26875 6266
rect 26909 6122 26921 6266
rect 26863 6110 26921 6122
rect 26991 6266 27049 6278
rect 26991 6122 27003 6266
rect 27037 6122 27049 6266
rect 26991 6110 27049 6122
rect 27119 6266 27177 6278
rect 27119 6122 27131 6266
rect 27165 6122 27177 6266
rect 27119 6110 27177 6122
rect 27247 6266 27305 6278
rect 27247 6122 27259 6266
rect 27293 6122 27305 6266
rect 27247 6110 27305 6122
rect 27375 6266 27433 6278
rect 27375 6122 27387 6266
rect 27421 6122 27433 6266
rect 27375 6110 27433 6122
rect 27503 6266 27561 6278
rect 27503 6122 27515 6266
rect 27549 6122 27561 6266
rect 27503 6110 27561 6122
rect 27631 6266 27689 6278
rect 27631 6122 27643 6266
rect 27677 6122 27689 6266
rect 27631 6110 27689 6122
rect 27759 6266 27817 6278
rect 27759 6122 27771 6266
rect 27805 6122 27817 6266
rect 27759 6110 27817 6122
rect 27887 6266 27945 6278
rect 27887 6122 27899 6266
rect 27933 6122 27945 6266
rect 27887 6110 27945 6122
rect 28015 6266 28073 6278
rect 28015 6122 28027 6266
rect 28061 6122 28073 6266
rect 28015 6110 28073 6122
rect 28143 6266 28201 6278
rect 28143 6122 28155 6266
rect 28189 6122 28201 6266
rect 28143 6110 28201 6122
rect 28271 6266 28329 6278
rect 28271 6122 28283 6266
rect 28317 6122 28329 6266
rect 28271 6110 28329 6122
rect 28399 6266 28457 6278
rect 28399 6122 28411 6266
rect 28445 6122 28457 6266
rect 28399 6110 28457 6122
rect 28527 6266 28585 6278
rect 28527 6122 28539 6266
rect 28573 6122 28585 6266
rect 28527 6110 28585 6122
rect -329 5578 -271 5590
rect -329 5434 -317 5578
rect -283 5434 -271 5578
rect -329 5422 -271 5434
rect -201 5578 -143 5590
rect -201 5434 -189 5578
rect -155 5434 -143 5578
rect -201 5422 -143 5434
rect 599 5578 657 5590
rect 599 5434 611 5578
rect 645 5434 657 5578
rect 599 5422 657 5434
rect 727 5578 785 5590
rect 727 5434 739 5578
rect 773 5434 785 5578
rect 727 5422 785 5434
rect 855 5578 913 5590
rect 855 5434 867 5578
rect 901 5434 913 5578
rect 855 5422 913 5434
rect 1863 5578 1921 5590
rect 1863 5434 1875 5578
rect 1909 5434 1921 5578
rect 1863 5422 1921 5434
rect 1991 5578 2049 5590
rect 1991 5434 2003 5578
rect 2037 5434 2049 5578
rect 1991 5422 2049 5434
rect 2119 5578 2177 5590
rect 2119 5434 2131 5578
rect 2165 5434 2177 5578
rect 2119 5422 2177 5434
rect 2247 5578 2305 5590
rect 2247 5434 2259 5578
rect 2293 5434 2305 5578
rect 2247 5422 2305 5434
rect 2375 5578 2433 5590
rect 2375 5434 2387 5578
rect 2421 5434 2433 5578
rect 2375 5422 2433 5434
rect 3482 5578 3540 5590
rect 3482 5434 3494 5578
rect 3528 5434 3540 5578
rect 3482 5422 3540 5434
rect 3610 5578 3668 5590
rect 3610 5434 3622 5578
rect 3656 5434 3668 5578
rect 3610 5422 3668 5434
rect 3738 5578 3796 5590
rect 3738 5434 3750 5578
rect 3784 5434 3796 5578
rect 3738 5422 3796 5434
rect 3866 5578 3924 5590
rect 3866 5434 3878 5578
rect 3912 5434 3924 5578
rect 3866 5422 3924 5434
rect 3994 5578 4052 5590
rect 3994 5434 4006 5578
rect 4040 5434 4052 5578
rect 3994 5422 4052 5434
rect 4122 5578 4180 5590
rect 4122 5434 4134 5578
rect 4168 5434 4180 5578
rect 4122 5422 4180 5434
rect 4250 5578 4308 5590
rect 4250 5434 4262 5578
rect 4296 5434 4308 5578
rect 4250 5422 4308 5434
rect 4378 5578 4436 5590
rect 4378 5434 4390 5578
rect 4424 5434 4436 5578
rect 4378 5422 4436 5434
rect 4506 5578 4564 5590
rect 4506 5434 4518 5578
rect 4552 5434 4564 5578
rect 4506 5422 4564 5434
rect 8047 5578 8105 5590
rect 8047 5434 8059 5578
rect 8093 5434 8105 5578
rect 8047 5422 8105 5434
rect 8175 5578 8233 5590
rect 8175 5434 8187 5578
rect 8221 5434 8233 5578
rect 8175 5422 8233 5434
rect 8303 5578 8361 5590
rect 8303 5434 8315 5578
rect 8349 5434 8361 5578
rect 8303 5422 8361 5434
rect 8431 5578 8489 5590
rect 8431 5434 8443 5578
rect 8477 5434 8489 5578
rect 8431 5422 8489 5434
rect 8559 5578 8617 5590
rect 8559 5434 8571 5578
rect 8605 5434 8617 5578
rect 8559 5422 8617 5434
rect 8687 5578 8745 5590
rect 8687 5434 8699 5578
rect 8733 5434 8745 5578
rect 8687 5422 8745 5434
rect 8815 5578 8873 5590
rect 8815 5434 8827 5578
rect 8861 5434 8873 5578
rect 8815 5422 8873 5434
rect 8943 5578 9001 5590
rect 8943 5434 8955 5578
rect 8989 5434 9001 5578
rect 8943 5422 9001 5434
rect 9071 5578 9129 5590
rect 9071 5434 9083 5578
rect 9117 5434 9129 5578
rect 9071 5422 9129 5434
rect 9199 5578 9257 5590
rect 9199 5434 9211 5578
rect 9245 5434 9257 5578
rect 9199 5422 9257 5434
rect 9327 5578 9385 5590
rect 9327 5434 9339 5578
rect 9373 5434 9385 5578
rect 9327 5422 9385 5434
rect 9455 5578 9513 5590
rect 9455 5434 9467 5578
rect 9501 5434 9513 5578
rect 9455 5422 9513 5434
rect 9583 5578 9641 5590
rect 9583 5434 9595 5578
rect 9629 5434 9641 5578
rect 9583 5422 9641 5434
rect 9711 5578 9769 5590
rect 9711 5434 9723 5578
rect 9757 5434 9769 5578
rect 9711 5422 9769 5434
rect 9839 5578 9897 5590
rect 9839 5434 9851 5578
rect 9885 5434 9897 5578
rect 9839 5422 9897 5434
rect 9967 5578 10025 5590
rect 9967 5434 9979 5578
rect 10013 5434 10025 5578
rect 9967 5422 10025 5434
rect 10095 5578 10153 5590
rect 10095 5434 10107 5578
rect 10141 5434 10153 5578
rect 10095 5422 10153 5434
rect 15205 5578 15263 5590
rect 15205 5434 15217 5578
rect 15251 5434 15263 5578
rect 15205 5422 15263 5434
rect 15333 5578 15391 5590
rect 15333 5434 15345 5578
rect 15379 5434 15391 5578
rect 15333 5422 15391 5434
rect 15461 5578 15519 5590
rect 15461 5434 15473 5578
rect 15507 5434 15519 5578
rect 15461 5422 15519 5434
rect 15589 5578 15647 5590
rect 15589 5434 15601 5578
rect 15635 5434 15647 5578
rect 15589 5422 15647 5434
rect 15717 5578 15775 5590
rect 15717 5434 15729 5578
rect 15763 5434 15775 5578
rect 15717 5422 15775 5434
rect 15845 5578 15903 5590
rect 15845 5434 15857 5578
rect 15891 5434 15903 5578
rect 15845 5422 15903 5434
rect 15973 5578 16031 5590
rect 15973 5434 15985 5578
rect 16019 5434 16031 5578
rect 15973 5422 16031 5434
rect 16101 5578 16159 5590
rect 16101 5434 16113 5578
rect 16147 5434 16159 5578
rect 16101 5422 16159 5434
rect 16229 5578 16287 5590
rect 16229 5434 16241 5578
rect 16275 5434 16287 5578
rect 16229 5422 16287 5434
rect 16357 5578 16415 5590
rect 16357 5434 16369 5578
rect 16403 5434 16415 5578
rect 16357 5422 16415 5434
rect 16485 5578 16543 5590
rect 16485 5434 16497 5578
rect 16531 5434 16543 5578
rect 16485 5422 16543 5434
rect 16613 5578 16671 5590
rect 16613 5434 16625 5578
rect 16659 5434 16671 5578
rect 16613 5422 16671 5434
rect 16741 5578 16799 5590
rect 16741 5434 16753 5578
rect 16787 5434 16799 5578
rect 16741 5422 16799 5434
rect 16869 5578 16927 5590
rect 16869 5434 16881 5578
rect 16915 5434 16927 5578
rect 16869 5422 16927 5434
rect 16997 5578 17055 5590
rect 16997 5434 17009 5578
rect 17043 5434 17055 5578
rect 16997 5422 17055 5434
rect 17125 5578 17183 5590
rect 17125 5434 17137 5578
rect 17171 5434 17183 5578
rect 17125 5422 17183 5434
rect 17253 5578 17311 5590
rect 17253 5434 17265 5578
rect 17299 5434 17311 5578
rect 17253 5422 17311 5434
rect 17381 5578 17439 5590
rect 17381 5434 17393 5578
rect 17427 5434 17439 5578
rect 17381 5422 17439 5434
rect 17509 5578 17567 5590
rect 17509 5434 17521 5578
rect 17555 5434 17567 5578
rect 17509 5422 17567 5434
rect 17637 5578 17695 5590
rect 17637 5434 17649 5578
rect 17683 5434 17695 5578
rect 17637 5422 17695 5434
rect 17765 5578 17823 5590
rect 17765 5434 17777 5578
rect 17811 5434 17823 5578
rect 17765 5422 17823 5434
rect 17893 5578 17951 5590
rect 17893 5434 17905 5578
rect 17939 5434 17951 5578
rect 17893 5422 17951 5434
rect 18021 5578 18079 5590
rect 18021 5434 18033 5578
rect 18067 5434 18079 5578
rect 18021 5422 18079 5434
rect 18149 5578 18207 5590
rect 18149 5434 18161 5578
rect 18195 5434 18207 5578
rect 18149 5422 18207 5434
rect 18277 5578 18335 5590
rect 18277 5434 18289 5578
rect 18323 5434 18335 5578
rect 18277 5422 18335 5434
rect 18405 5578 18463 5590
rect 18405 5434 18417 5578
rect 18451 5434 18463 5578
rect 18405 5422 18463 5434
rect 18533 5578 18591 5590
rect 18533 5434 18545 5578
rect 18579 5434 18591 5578
rect 18533 5422 18591 5434
rect 18661 5578 18719 5590
rect 18661 5434 18673 5578
rect 18707 5434 18719 5578
rect 18661 5422 18719 5434
rect 18789 5578 18847 5590
rect 18789 5434 18801 5578
rect 18835 5434 18847 5578
rect 18789 5422 18847 5434
rect 18917 5578 18975 5590
rect 18917 5434 18929 5578
rect 18963 5434 18975 5578
rect 18917 5422 18975 5434
rect 19045 5578 19103 5590
rect 19045 5434 19057 5578
rect 19091 5434 19103 5578
rect 19045 5422 19103 5434
rect 19173 5578 19231 5590
rect 19173 5434 19185 5578
rect 19219 5434 19231 5578
rect 19173 5422 19231 5434
rect 19301 5578 19359 5590
rect 19301 5434 19313 5578
rect 19347 5434 19359 5578
rect 19301 5422 19359 5434
rect 20259 5578 20317 5590
rect 20259 5434 20271 5578
rect 20305 5434 20317 5578
rect 20259 5422 20317 5434
rect 20387 5578 20445 5590
rect 20387 5434 20399 5578
rect 20433 5434 20445 5578
rect 20387 5422 20445 5434
rect 20515 5578 20573 5590
rect 20515 5434 20527 5578
rect 20561 5434 20573 5578
rect 20515 5422 20573 5434
rect 20643 5578 20701 5590
rect 20643 5434 20655 5578
rect 20689 5434 20701 5578
rect 20643 5422 20701 5434
rect 20771 5578 20829 5590
rect 20771 5434 20783 5578
rect 20817 5434 20829 5578
rect 20771 5422 20829 5434
rect 20899 5578 20957 5590
rect 20899 5434 20911 5578
rect 20945 5434 20957 5578
rect 20899 5422 20957 5434
rect 21027 5578 21085 5590
rect 21027 5434 21039 5578
rect 21073 5434 21085 5578
rect 21027 5422 21085 5434
rect 21155 5578 21213 5590
rect 21155 5434 21167 5578
rect 21201 5434 21213 5578
rect 21155 5422 21213 5434
rect 21283 5578 21341 5590
rect 21283 5434 21295 5578
rect 21329 5434 21341 5578
rect 21283 5422 21341 5434
rect 21411 5578 21469 5590
rect 21411 5434 21423 5578
rect 21457 5434 21469 5578
rect 21411 5422 21469 5434
rect 21539 5578 21597 5590
rect 21539 5434 21551 5578
rect 21585 5434 21597 5578
rect 21539 5422 21597 5434
rect 21667 5578 21725 5590
rect 21667 5434 21679 5578
rect 21713 5434 21725 5578
rect 21667 5422 21725 5434
rect 21795 5578 21853 5590
rect 21795 5434 21807 5578
rect 21841 5434 21853 5578
rect 21795 5422 21853 5434
rect 21923 5578 21981 5590
rect 21923 5434 21935 5578
rect 21969 5434 21981 5578
rect 21923 5422 21981 5434
rect 22051 5578 22109 5590
rect 22051 5434 22063 5578
rect 22097 5434 22109 5578
rect 22051 5422 22109 5434
rect 22179 5578 22237 5590
rect 22179 5434 22191 5578
rect 22225 5434 22237 5578
rect 22179 5422 22237 5434
rect 22307 5578 22365 5590
rect 22307 5434 22319 5578
rect 22353 5434 22365 5578
rect 22307 5422 22365 5434
rect 22435 5578 22493 5590
rect 22435 5434 22447 5578
rect 22481 5434 22493 5578
rect 22435 5422 22493 5434
rect 22563 5578 22621 5590
rect 22563 5434 22575 5578
rect 22609 5434 22621 5578
rect 22563 5422 22621 5434
rect 22691 5578 22749 5590
rect 22691 5434 22703 5578
rect 22737 5434 22749 5578
rect 22691 5422 22749 5434
rect 22819 5578 22877 5590
rect 22819 5434 22831 5578
rect 22865 5434 22877 5578
rect 22819 5422 22877 5434
rect 22947 5578 23005 5590
rect 22947 5434 22959 5578
rect 22993 5434 23005 5578
rect 22947 5422 23005 5434
rect 23075 5578 23133 5590
rect 23075 5434 23087 5578
rect 23121 5434 23133 5578
rect 23075 5422 23133 5434
rect 23203 5578 23261 5590
rect 23203 5434 23215 5578
rect 23249 5434 23261 5578
rect 23203 5422 23261 5434
rect 23331 5578 23389 5590
rect 23331 5434 23343 5578
rect 23377 5434 23389 5578
rect 23331 5422 23389 5434
rect 23459 5578 23517 5590
rect 23459 5434 23471 5578
rect 23505 5434 23517 5578
rect 23459 5422 23517 5434
rect 23587 5578 23645 5590
rect 23587 5434 23599 5578
rect 23633 5434 23645 5578
rect 23587 5422 23645 5434
rect 23715 5578 23773 5590
rect 23715 5434 23727 5578
rect 23761 5434 23773 5578
rect 23715 5422 23773 5434
rect 23843 5578 23901 5590
rect 23843 5434 23855 5578
rect 23889 5434 23901 5578
rect 23843 5422 23901 5434
rect 23971 5578 24029 5590
rect 23971 5434 23983 5578
rect 24017 5434 24029 5578
rect 23971 5422 24029 5434
rect 24099 5578 24157 5590
rect 24099 5434 24111 5578
rect 24145 5434 24157 5578
rect 24099 5422 24157 5434
rect 24227 5578 24285 5590
rect 24227 5434 24239 5578
rect 24273 5434 24285 5578
rect 24227 5422 24285 5434
rect 24355 5578 24413 5590
rect 24355 5434 24367 5578
rect 24401 5434 24413 5578
rect 24355 5422 24413 5434
rect 24483 5578 24541 5590
rect 24483 5434 24495 5578
rect 24529 5434 24541 5578
rect 24483 5422 24541 5434
rect 24611 5578 24669 5590
rect 24611 5434 24623 5578
rect 24657 5434 24669 5578
rect 24611 5422 24669 5434
rect 24739 5578 24797 5590
rect 24739 5434 24751 5578
rect 24785 5434 24797 5578
rect 24739 5422 24797 5434
rect 24867 5578 24925 5590
rect 24867 5434 24879 5578
rect 24913 5434 24925 5578
rect 24867 5422 24925 5434
rect 24995 5578 25053 5590
rect 24995 5434 25007 5578
rect 25041 5434 25053 5578
rect 24995 5422 25053 5434
rect 25123 5578 25181 5590
rect 25123 5434 25135 5578
rect 25169 5434 25181 5578
rect 25123 5422 25181 5434
rect 25251 5578 25309 5590
rect 25251 5434 25263 5578
rect 25297 5434 25309 5578
rect 25251 5422 25309 5434
rect 25379 5578 25437 5590
rect 25379 5434 25391 5578
rect 25425 5434 25437 5578
rect 25379 5422 25437 5434
rect 25507 5578 25565 5590
rect 25507 5434 25519 5578
rect 25553 5434 25565 5578
rect 25507 5422 25565 5434
rect 25635 5578 25693 5590
rect 25635 5434 25647 5578
rect 25681 5434 25693 5578
rect 25635 5422 25693 5434
rect 25763 5578 25821 5590
rect 25763 5434 25775 5578
rect 25809 5434 25821 5578
rect 25763 5422 25821 5434
rect 25891 5578 25949 5590
rect 25891 5434 25903 5578
rect 25937 5434 25949 5578
rect 25891 5422 25949 5434
rect 26019 5578 26077 5590
rect 26019 5434 26031 5578
rect 26065 5434 26077 5578
rect 26019 5422 26077 5434
rect 26147 5578 26205 5590
rect 26147 5434 26159 5578
rect 26193 5434 26205 5578
rect 26147 5422 26205 5434
rect 26275 5578 26333 5590
rect 26275 5434 26287 5578
rect 26321 5434 26333 5578
rect 26275 5422 26333 5434
rect 26403 5578 26461 5590
rect 26403 5434 26415 5578
rect 26449 5434 26461 5578
rect 26403 5422 26461 5434
rect 26531 5578 26589 5590
rect 26531 5434 26543 5578
rect 26577 5434 26589 5578
rect 26531 5422 26589 5434
rect 26659 5578 26717 5590
rect 26659 5434 26671 5578
rect 26705 5434 26717 5578
rect 26659 5422 26717 5434
rect 26787 5578 26845 5590
rect 26787 5434 26799 5578
rect 26833 5434 26845 5578
rect 26787 5422 26845 5434
rect 26915 5578 26973 5590
rect 26915 5434 26927 5578
rect 26961 5434 26973 5578
rect 26915 5422 26973 5434
rect 27043 5578 27101 5590
rect 27043 5434 27055 5578
rect 27089 5434 27101 5578
rect 27043 5422 27101 5434
rect 27171 5578 27229 5590
rect 27171 5434 27183 5578
rect 27217 5434 27229 5578
rect 27171 5422 27229 5434
rect 27299 5578 27357 5590
rect 27299 5434 27311 5578
rect 27345 5434 27357 5578
rect 27299 5422 27357 5434
rect 27427 5578 27485 5590
rect 27427 5434 27439 5578
rect 27473 5434 27485 5578
rect 27427 5422 27485 5434
rect 27555 5578 27613 5590
rect 27555 5434 27567 5578
rect 27601 5434 27613 5578
rect 27555 5422 27613 5434
rect 27683 5578 27741 5590
rect 27683 5434 27695 5578
rect 27729 5434 27741 5578
rect 27683 5422 27741 5434
rect 27811 5578 27869 5590
rect 27811 5434 27823 5578
rect 27857 5434 27869 5578
rect 27811 5422 27869 5434
rect 27939 5578 27997 5590
rect 27939 5434 27951 5578
rect 27985 5434 27997 5578
rect 27939 5422 27997 5434
rect 28067 5578 28125 5590
rect 28067 5434 28079 5578
rect 28113 5434 28125 5578
rect 28067 5422 28125 5434
rect 28195 5578 28253 5590
rect 28195 5434 28207 5578
rect 28241 5434 28253 5578
rect 28195 5422 28253 5434
rect 28323 5578 28381 5590
rect 28323 5434 28335 5578
rect 28369 5434 28381 5578
rect 28323 5422 28381 5434
rect 28451 5578 28509 5590
rect 28451 5434 28463 5578
rect 28497 5434 28509 5578
rect 28451 5422 28509 5434
<< ndiffc >>
rect -295 5906 -261 5966
rect -167 5906 -133 5966
rect 482 5906 516 5966
rect 610 5906 644 5966
rect 738 5906 772 5966
rect 1391 5906 1425 5966
rect 1519 5906 1553 5966
rect 1647 5906 1681 5966
rect 1775 5906 1809 5966
rect 1903 5906 1937 5966
rect 2924 5906 2958 5966
rect 3052 5906 3086 5966
rect 3180 5906 3214 5966
rect 3308 5906 3342 5966
rect 3436 5906 3470 5966
rect 3564 5906 3598 5966
rect 3692 5906 3726 5966
rect 3820 5906 3854 5966
rect 3948 5906 3982 5966
rect 5475 5906 5509 5966
rect 5603 5906 5637 5966
rect 5731 5906 5765 5966
rect 5859 5906 5893 5966
rect 5987 5906 6021 5966
rect 6115 5906 6149 5966
rect 6243 5906 6277 5966
rect 6371 5906 6405 5966
rect 6499 5906 6533 5966
rect 6627 5906 6661 5966
rect 6755 5906 6789 5966
rect 6883 5906 6917 5966
rect 7011 5906 7045 5966
rect 7139 5906 7173 5966
rect 7267 5906 7301 5966
rect 7395 5906 7429 5966
rect 7523 5906 7557 5966
rect 10562 5906 10596 5966
rect 10690 5906 10724 5966
rect 10818 5906 10852 5966
rect 10946 5906 10980 5966
rect 11074 5906 11108 5966
rect 11202 5906 11236 5966
rect 11330 5906 11364 5966
rect 11458 5906 11492 5966
rect 11586 5906 11620 5966
rect 11714 5906 11748 5966
rect 11842 5906 11876 5966
rect 11970 5906 12004 5966
rect 12098 5906 12132 5966
rect 12226 5906 12260 5966
rect 12354 5906 12388 5966
rect 12482 5906 12516 5966
rect 12610 5906 12644 5966
rect 12738 5906 12772 5966
rect 12866 5906 12900 5966
rect 12994 5906 13028 5966
rect 13122 5906 13156 5966
rect 13250 5906 13284 5966
rect 13378 5906 13412 5966
rect 13506 5906 13540 5966
rect 13634 5906 13668 5966
rect 13762 5906 13796 5966
rect 13890 5906 13924 5966
rect 14018 5906 14052 5966
rect 14146 5906 14180 5966
rect 14274 5906 14308 5966
rect 14402 5906 14436 5966
rect 14530 5906 14564 5966
rect 14658 5906 14692 5966
rect 20347 5906 20381 5966
rect 20475 5906 20509 5966
rect 20603 5906 20637 5966
rect 20731 5906 20765 5966
rect 20859 5906 20893 5966
rect 20987 5906 21021 5966
rect 21115 5906 21149 5966
rect 21243 5906 21277 5966
rect 21371 5906 21405 5966
rect 21499 5906 21533 5966
rect 21627 5906 21661 5966
rect 21755 5906 21789 5966
rect 21883 5906 21917 5966
rect 22011 5906 22045 5966
rect 22139 5906 22173 5966
rect 22267 5906 22301 5966
rect 22395 5906 22429 5966
rect 22523 5906 22557 5966
rect 22651 5906 22685 5966
rect 22779 5906 22813 5966
rect 22907 5906 22941 5966
rect 23035 5906 23069 5966
rect 23163 5906 23197 5966
rect 23291 5906 23325 5966
rect 23419 5906 23453 5966
rect 23547 5906 23581 5966
rect 23675 5906 23709 5966
rect 23803 5906 23837 5966
rect 23931 5906 23965 5966
rect 24059 5906 24093 5966
rect 24187 5906 24221 5966
rect 24315 5906 24349 5966
rect 24443 5906 24477 5966
rect 24571 5906 24605 5966
rect 24699 5906 24733 5966
rect 24827 5906 24861 5966
rect 24955 5906 24989 5966
rect 25083 5906 25117 5966
rect 25211 5906 25245 5966
rect 25339 5906 25373 5966
rect 25467 5906 25501 5966
rect 25595 5906 25629 5966
rect 25723 5906 25757 5966
rect 25851 5906 25885 5966
rect 25979 5906 26013 5966
rect 26107 5906 26141 5966
rect 26235 5906 26269 5966
rect 26363 5906 26397 5966
rect 26491 5906 26525 5966
rect 26619 5906 26653 5966
rect 26747 5906 26781 5966
rect 26875 5906 26909 5966
rect 27003 5906 27037 5966
rect 27131 5906 27165 5966
rect 27259 5906 27293 5966
rect 27387 5906 27421 5966
rect 27515 5906 27549 5966
rect 27643 5906 27677 5966
rect 27771 5906 27805 5966
rect 27899 5906 27933 5966
rect 28027 5906 28061 5966
rect 28155 5906 28189 5966
rect 28283 5906 28317 5966
rect 28411 5906 28445 5966
rect 28539 5906 28573 5966
rect -317 5218 -283 5278
rect -189 5218 -155 5278
rect 611 5218 645 5278
rect 739 5218 773 5278
rect 867 5218 901 5278
rect 1875 5218 1909 5278
rect 2003 5218 2037 5278
rect 2131 5218 2165 5278
rect 2259 5218 2293 5278
rect 2387 5218 2421 5278
rect 3494 5218 3528 5278
rect 3622 5218 3656 5278
rect 3750 5218 3784 5278
rect 3878 5218 3912 5278
rect 4006 5218 4040 5278
rect 4134 5218 4168 5278
rect 4262 5218 4296 5278
rect 4390 5218 4424 5278
rect 4518 5218 4552 5278
rect 8059 5218 8093 5278
rect 8187 5218 8221 5278
rect 8315 5218 8349 5278
rect 8443 5218 8477 5278
rect 8571 5218 8605 5278
rect 8699 5218 8733 5278
rect 8827 5218 8861 5278
rect 8955 5218 8989 5278
rect 9083 5218 9117 5278
rect 9211 5218 9245 5278
rect 9339 5218 9373 5278
rect 9467 5218 9501 5278
rect 9595 5218 9629 5278
rect 9723 5218 9757 5278
rect 9851 5218 9885 5278
rect 9979 5218 10013 5278
rect 10107 5218 10141 5278
rect 15217 5218 15251 5278
rect 15345 5218 15379 5278
rect 15473 5218 15507 5278
rect 15601 5218 15635 5278
rect 15729 5218 15763 5278
rect 15857 5218 15891 5278
rect 15985 5218 16019 5278
rect 16113 5218 16147 5278
rect 16241 5218 16275 5278
rect 16369 5218 16403 5278
rect 16497 5218 16531 5278
rect 16625 5218 16659 5278
rect 16753 5218 16787 5278
rect 16881 5218 16915 5278
rect 17009 5218 17043 5278
rect 17137 5218 17171 5278
rect 17265 5218 17299 5278
rect 17393 5218 17427 5278
rect 17521 5218 17555 5278
rect 17649 5218 17683 5278
rect 17777 5218 17811 5278
rect 17905 5218 17939 5278
rect 18033 5218 18067 5278
rect 18161 5218 18195 5278
rect 18289 5218 18323 5278
rect 18417 5218 18451 5278
rect 18545 5218 18579 5278
rect 18673 5218 18707 5278
rect 18801 5218 18835 5278
rect 18929 5218 18963 5278
rect 19057 5218 19091 5278
rect 19185 5218 19219 5278
rect 19313 5218 19347 5278
rect 20271 5218 20305 5278
rect 20399 5218 20433 5278
rect 20527 5218 20561 5278
rect 20655 5218 20689 5278
rect 20783 5218 20817 5278
rect 20911 5218 20945 5278
rect 21039 5218 21073 5278
rect 21167 5218 21201 5278
rect 21295 5218 21329 5278
rect 21423 5218 21457 5278
rect 21551 5218 21585 5278
rect 21679 5218 21713 5278
rect 21807 5218 21841 5278
rect 21935 5218 21969 5278
rect 22063 5218 22097 5278
rect 22191 5218 22225 5278
rect 22319 5218 22353 5278
rect 22447 5218 22481 5278
rect 22575 5218 22609 5278
rect 22703 5218 22737 5278
rect 22831 5218 22865 5278
rect 22959 5218 22993 5278
rect 23087 5218 23121 5278
rect 23215 5218 23249 5278
rect 23343 5218 23377 5278
rect 23471 5218 23505 5278
rect 23599 5218 23633 5278
rect 23727 5218 23761 5278
rect 23855 5218 23889 5278
rect 23983 5218 24017 5278
rect 24111 5218 24145 5278
rect 24239 5218 24273 5278
rect 24367 5218 24401 5278
rect 24495 5218 24529 5278
rect 24623 5218 24657 5278
rect 24751 5218 24785 5278
rect 24879 5218 24913 5278
rect 25007 5218 25041 5278
rect 25135 5218 25169 5278
rect 25263 5218 25297 5278
rect 25391 5218 25425 5278
rect 25519 5218 25553 5278
rect 25647 5218 25681 5278
rect 25775 5218 25809 5278
rect 25903 5218 25937 5278
rect 26031 5218 26065 5278
rect 26159 5218 26193 5278
rect 26287 5218 26321 5278
rect 26415 5218 26449 5278
rect 26543 5218 26577 5278
rect 26671 5218 26705 5278
rect 26799 5218 26833 5278
rect 26927 5218 26961 5278
rect 27055 5218 27089 5278
rect 27183 5218 27217 5278
rect 27311 5218 27345 5278
rect 27439 5218 27473 5278
rect 27567 5218 27601 5278
rect 27695 5218 27729 5278
rect 27823 5218 27857 5278
rect 27951 5218 27985 5278
rect 28079 5218 28113 5278
rect 28207 5218 28241 5278
rect 28335 5218 28369 5278
rect 28463 5218 28497 5278
<< pdiffc >>
rect -295 6122 -261 6266
rect -167 6122 -133 6266
rect 482 6122 516 6266
rect 610 6122 644 6266
rect 738 6122 772 6266
rect 1391 6122 1425 6266
rect 1519 6122 1553 6266
rect 1647 6122 1681 6266
rect 1775 6122 1809 6266
rect 1903 6122 1937 6266
rect 2924 6122 2958 6266
rect 3052 6122 3086 6266
rect 3180 6122 3214 6266
rect 3308 6122 3342 6266
rect 3436 6122 3470 6266
rect 3564 6122 3598 6266
rect 3692 6122 3726 6266
rect 3820 6122 3854 6266
rect 3948 6122 3982 6266
rect 5475 6122 5509 6266
rect 5603 6122 5637 6266
rect 5731 6122 5765 6266
rect 5859 6122 5893 6266
rect 5987 6122 6021 6266
rect 6115 6122 6149 6266
rect 6243 6122 6277 6266
rect 6371 6122 6405 6266
rect 6499 6122 6533 6266
rect 6627 6122 6661 6266
rect 6755 6122 6789 6266
rect 6883 6122 6917 6266
rect 7011 6122 7045 6266
rect 7139 6122 7173 6266
rect 7267 6122 7301 6266
rect 7395 6122 7429 6266
rect 7523 6122 7557 6266
rect 10562 6122 10596 6266
rect 10690 6122 10724 6266
rect 10818 6122 10852 6266
rect 10946 6122 10980 6266
rect 11074 6122 11108 6266
rect 11202 6122 11236 6266
rect 11330 6122 11364 6266
rect 11458 6122 11492 6266
rect 11586 6122 11620 6266
rect 11714 6122 11748 6266
rect 11842 6122 11876 6266
rect 11970 6122 12004 6266
rect 12098 6122 12132 6266
rect 12226 6122 12260 6266
rect 12354 6122 12388 6266
rect 12482 6122 12516 6266
rect 12610 6122 12644 6266
rect 12738 6122 12772 6266
rect 12866 6122 12900 6266
rect 12994 6122 13028 6266
rect 13122 6122 13156 6266
rect 13250 6122 13284 6266
rect 13378 6122 13412 6266
rect 13506 6122 13540 6266
rect 13634 6122 13668 6266
rect 13762 6122 13796 6266
rect 13890 6122 13924 6266
rect 14018 6122 14052 6266
rect 14146 6122 14180 6266
rect 14274 6122 14308 6266
rect 14402 6122 14436 6266
rect 14530 6122 14564 6266
rect 14658 6122 14692 6266
rect 20347 6122 20381 6266
rect 20475 6122 20509 6266
rect 20603 6122 20637 6266
rect 20731 6122 20765 6266
rect 20859 6122 20893 6266
rect 20987 6122 21021 6266
rect 21115 6122 21149 6266
rect 21243 6122 21277 6266
rect 21371 6122 21405 6266
rect 21499 6122 21533 6266
rect 21627 6122 21661 6266
rect 21755 6122 21789 6266
rect 21883 6122 21917 6266
rect 22011 6122 22045 6266
rect 22139 6122 22173 6266
rect 22267 6122 22301 6266
rect 22395 6122 22429 6266
rect 22523 6122 22557 6266
rect 22651 6122 22685 6266
rect 22779 6122 22813 6266
rect 22907 6122 22941 6266
rect 23035 6122 23069 6266
rect 23163 6122 23197 6266
rect 23291 6122 23325 6266
rect 23419 6122 23453 6266
rect 23547 6122 23581 6266
rect 23675 6122 23709 6266
rect 23803 6122 23837 6266
rect 23931 6122 23965 6266
rect 24059 6122 24093 6266
rect 24187 6122 24221 6266
rect 24315 6122 24349 6266
rect 24443 6122 24477 6266
rect 24571 6122 24605 6266
rect 24699 6122 24733 6266
rect 24827 6122 24861 6266
rect 24955 6122 24989 6266
rect 25083 6122 25117 6266
rect 25211 6122 25245 6266
rect 25339 6122 25373 6266
rect 25467 6122 25501 6266
rect 25595 6122 25629 6266
rect 25723 6122 25757 6266
rect 25851 6122 25885 6266
rect 25979 6122 26013 6266
rect 26107 6122 26141 6266
rect 26235 6122 26269 6266
rect 26363 6122 26397 6266
rect 26491 6122 26525 6266
rect 26619 6122 26653 6266
rect 26747 6122 26781 6266
rect 26875 6122 26909 6266
rect 27003 6122 27037 6266
rect 27131 6122 27165 6266
rect 27259 6122 27293 6266
rect 27387 6122 27421 6266
rect 27515 6122 27549 6266
rect 27643 6122 27677 6266
rect 27771 6122 27805 6266
rect 27899 6122 27933 6266
rect 28027 6122 28061 6266
rect 28155 6122 28189 6266
rect 28283 6122 28317 6266
rect 28411 6122 28445 6266
rect 28539 6122 28573 6266
rect -317 5434 -283 5578
rect -189 5434 -155 5578
rect 611 5434 645 5578
rect 739 5434 773 5578
rect 867 5434 901 5578
rect 1875 5434 1909 5578
rect 2003 5434 2037 5578
rect 2131 5434 2165 5578
rect 2259 5434 2293 5578
rect 2387 5434 2421 5578
rect 3494 5434 3528 5578
rect 3622 5434 3656 5578
rect 3750 5434 3784 5578
rect 3878 5434 3912 5578
rect 4006 5434 4040 5578
rect 4134 5434 4168 5578
rect 4262 5434 4296 5578
rect 4390 5434 4424 5578
rect 4518 5434 4552 5578
rect 8059 5434 8093 5578
rect 8187 5434 8221 5578
rect 8315 5434 8349 5578
rect 8443 5434 8477 5578
rect 8571 5434 8605 5578
rect 8699 5434 8733 5578
rect 8827 5434 8861 5578
rect 8955 5434 8989 5578
rect 9083 5434 9117 5578
rect 9211 5434 9245 5578
rect 9339 5434 9373 5578
rect 9467 5434 9501 5578
rect 9595 5434 9629 5578
rect 9723 5434 9757 5578
rect 9851 5434 9885 5578
rect 9979 5434 10013 5578
rect 10107 5434 10141 5578
rect 15217 5434 15251 5578
rect 15345 5434 15379 5578
rect 15473 5434 15507 5578
rect 15601 5434 15635 5578
rect 15729 5434 15763 5578
rect 15857 5434 15891 5578
rect 15985 5434 16019 5578
rect 16113 5434 16147 5578
rect 16241 5434 16275 5578
rect 16369 5434 16403 5578
rect 16497 5434 16531 5578
rect 16625 5434 16659 5578
rect 16753 5434 16787 5578
rect 16881 5434 16915 5578
rect 17009 5434 17043 5578
rect 17137 5434 17171 5578
rect 17265 5434 17299 5578
rect 17393 5434 17427 5578
rect 17521 5434 17555 5578
rect 17649 5434 17683 5578
rect 17777 5434 17811 5578
rect 17905 5434 17939 5578
rect 18033 5434 18067 5578
rect 18161 5434 18195 5578
rect 18289 5434 18323 5578
rect 18417 5434 18451 5578
rect 18545 5434 18579 5578
rect 18673 5434 18707 5578
rect 18801 5434 18835 5578
rect 18929 5434 18963 5578
rect 19057 5434 19091 5578
rect 19185 5434 19219 5578
rect 19313 5434 19347 5578
rect 20271 5434 20305 5578
rect 20399 5434 20433 5578
rect 20527 5434 20561 5578
rect 20655 5434 20689 5578
rect 20783 5434 20817 5578
rect 20911 5434 20945 5578
rect 21039 5434 21073 5578
rect 21167 5434 21201 5578
rect 21295 5434 21329 5578
rect 21423 5434 21457 5578
rect 21551 5434 21585 5578
rect 21679 5434 21713 5578
rect 21807 5434 21841 5578
rect 21935 5434 21969 5578
rect 22063 5434 22097 5578
rect 22191 5434 22225 5578
rect 22319 5434 22353 5578
rect 22447 5434 22481 5578
rect 22575 5434 22609 5578
rect 22703 5434 22737 5578
rect 22831 5434 22865 5578
rect 22959 5434 22993 5578
rect 23087 5434 23121 5578
rect 23215 5434 23249 5578
rect 23343 5434 23377 5578
rect 23471 5434 23505 5578
rect 23599 5434 23633 5578
rect 23727 5434 23761 5578
rect 23855 5434 23889 5578
rect 23983 5434 24017 5578
rect 24111 5434 24145 5578
rect 24239 5434 24273 5578
rect 24367 5434 24401 5578
rect 24495 5434 24529 5578
rect 24623 5434 24657 5578
rect 24751 5434 24785 5578
rect 24879 5434 24913 5578
rect 25007 5434 25041 5578
rect 25135 5434 25169 5578
rect 25263 5434 25297 5578
rect 25391 5434 25425 5578
rect 25519 5434 25553 5578
rect 25647 5434 25681 5578
rect 25775 5434 25809 5578
rect 25903 5434 25937 5578
rect 26031 5434 26065 5578
rect 26159 5434 26193 5578
rect 26287 5434 26321 5578
rect 26415 5434 26449 5578
rect 26543 5434 26577 5578
rect 26671 5434 26705 5578
rect 26799 5434 26833 5578
rect 26927 5434 26961 5578
rect 27055 5434 27089 5578
rect 27183 5434 27217 5578
rect 27311 5434 27345 5578
rect 27439 5434 27473 5578
rect 27567 5434 27601 5578
rect 27695 5434 27729 5578
rect 27823 5434 27857 5578
rect 27951 5434 27985 5578
rect 28079 5434 28113 5578
rect 28207 5434 28241 5578
rect 28335 5434 28369 5578
rect 28463 5434 28497 5578
<< psubdiff >>
rect -341 5836 7603 5840
rect -341 5798 -297 5836
rect -259 5798 -169 5836
rect -131 5798 480 5836
rect 518 5798 608 5836
rect 646 5798 736 5836
rect 774 5798 1389 5836
rect 1427 5798 1517 5836
rect 1555 5798 1645 5836
rect 1683 5798 1773 5836
rect 1811 5798 1901 5836
rect 1939 5798 2922 5836
rect 2960 5798 3050 5836
rect 3088 5798 3178 5836
rect 3216 5798 3306 5836
rect 3344 5798 3434 5836
rect 3472 5798 3562 5836
rect 3600 5798 3690 5836
rect 3728 5798 3818 5836
rect 3856 5798 3946 5836
rect 3984 5798 5473 5836
rect 5511 5798 5601 5836
rect 5639 5798 5729 5836
rect 5767 5798 5857 5836
rect 5895 5798 5985 5836
rect 6023 5798 6113 5836
rect 6151 5798 6241 5836
rect 6279 5798 6369 5836
rect 6407 5798 6497 5836
rect 6535 5798 6625 5836
rect 6663 5798 6753 5836
rect 6791 5798 6881 5836
rect 6919 5798 7009 5836
rect 7047 5798 7137 5836
rect 7175 5798 7265 5836
rect 7303 5798 7393 5836
rect 7431 5798 7521 5836
rect 7559 5798 7603 5836
rect -341 5794 7603 5798
rect 10516 5836 28619 5840
rect 10516 5798 10560 5836
rect 10598 5798 10688 5836
rect 10726 5798 10816 5836
rect 10854 5798 10944 5836
rect 10982 5798 11072 5836
rect 11110 5798 11200 5836
rect 11238 5798 11328 5836
rect 11366 5798 11456 5836
rect 11494 5798 11584 5836
rect 11622 5798 11712 5836
rect 11750 5798 11840 5836
rect 11878 5798 11968 5836
rect 12006 5798 12096 5836
rect 12134 5798 12224 5836
rect 12262 5798 12352 5836
rect 12390 5798 12480 5836
rect 12518 5798 12608 5836
rect 12646 5798 12736 5836
rect 12774 5798 12864 5836
rect 12902 5798 12992 5836
rect 13030 5798 13120 5836
rect 13158 5798 13248 5836
rect 13286 5798 13376 5836
rect 13414 5798 13504 5836
rect 13542 5798 13632 5836
rect 13670 5798 13760 5836
rect 13798 5798 13888 5836
rect 13926 5798 14016 5836
rect 14054 5798 14144 5836
rect 14182 5798 14272 5836
rect 14310 5798 14400 5836
rect 14438 5798 14528 5836
rect 14566 5798 14656 5836
rect 14694 5798 20345 5836
rect 20383 5798 20473 5836
rect 20511 5798 20601 5836
rect 20639 5798 20729 5836
rect 20767 5798 20857 5836
rect 20895 5798 20985 5836
rect 21023 5798 21113 5836
rect 21151 5798 21241 5836
rect 21279 5798 21369 5836
rect 21407 5798 21497 5836
rect 21535 5798 21625 5836
rect 21663 5798 21753 5836
rect 21791 5798 21881 5836
rect 21919 5798 22009 5836
rect 22047 5798 22137 5836
rect 22175 5798 22265 5836
rect 22303 5798 22393 5836
rect 22431 5798 22521 5836
rect 22559 5798 22649 5836
rect 22687 5798 22777 5836
rect 22815 5798 22905 5836
rect 22943 5798 23033 5836
rect 23071 5798 23161 5836
rect 23199 5798 23289 5836
rect 23327 5798 23417 5836
rect 23455 5798 23545 5836
rect 23583 5798 23673 5836
rect 23711 5798 23801 5836
rect 23839 5798 23929 5836
rect 23967 5798 24057 5836
rect 24095 5798 24185 5836
rect 24223 5798 24313 5836
rect 24351 5798 24441 5836
rect 24479 5798 24569 5836
rect 24607 5798 24697 5836
rect 24735 5798 24825 5836
rect 24863 5798 24953 5836
rect 24991 5798 25081 5836
rect 25119 5798 25209 5836
rect 25247 5798 25337 5836
rect 25375 5798 25465 5836
rect 25503 5798 25593 5836
rect 25631 5798 25721 5836
rect 25759 5798 25849 5836
rect 25887 5798 25977 5836
rect 26015 5798 26105 5836
rect 26143 5798 26233 5836
rect 26271 5798 26361 5836
rect 26399 5798 26489 5836
rect 26527 5798 26617 5836
rect 26655 5798 26745 5836
rect 26783 5798 26873 5836
rect 26911 5798 27001 5836
rect 27039 5798 27129 5836
rect 27167 5798 27257 5836
rect 27295 5798 27385 5836
rect 27423 5798 27513 5836
rect 27551 5798 27641 5836
rect 27679 5798 27769 5836
rect 27807 5798 27897 5836
rect 27935 5798 28025 5836
rect 28063 5798 28153 5836
rect 28191 5798 28281 5836
rect 28319 5798 28409 5836
rect 28447 5798 28537 5836
rect 28575 5798 28619 5836
rect 10516 5794 28619 5798
rect -363 5148 947 5152
rect -363 5110 -319 5148
rect -281 5110 -191 5148
rect -153 5110 609 5148
rect 647 5110 737 5148
rect 775 5110 865 5148
rect 903 5110 947 5148
rect -363 5106 947 5110
rect 1829 5148 2467 5152
rect 1829 5110 1873 5148
rect 1911 5110 2001 5148
rect 2039 5110 2129 5148
rect 2167 5110 2257 5148
rect 2295 5110 2385 5148
rect 2423 5110 2467 5148
rect 1829 5106 2467 5110
rect 3448 5148 28543 5152
rect 3448 5110 3492 5148
rect 3530 5110 3620 5148
rect 3658 5110 3748 5148
rect 3786 5110 3876 5148
rect 3914 5110 4004 5148
rect 4042 5110 4132 5148
rect 4170 5110 4260 5148
rect 4298 5110 4388 5148
rect 4426 5110 4516 5148
rect 4554 5110 8057 5148
rect 8095 5110 8185 5148
rect 8223 5110 8313 5148
rect 8351 5110 8441 5148
rect 8479 5110 8569 5148
rect 8607 5110 8697 5148
rect 8735 5110 8825 5148
rect 8863 5110 8953 5148
rect 8991 5110 9081 5148
rect 9119 5110 9209 5148
rect 9247 5110 9337 5148
rect 9375 5110 9465 5148
rect 9503 5110 9593 5148
rect 9631 5110 9721 5148
rect 9759 5110 9849 5148
rect 9887 5110 9977 5148
rect 10015 5110 10105 5148
rect 10143 5110 15215 5148
rect 15253 5110 15343 5148
rect 15381 5110 15471 5148
rect 15509 5110 15599 5148
rect 15637 5110 15727 5148
rect 15765 5110 15855 5148
rect 15893 5110 15983 5148
rect 16021 5110 16111 5148
rect 16149 5110 16239 5148
rect 16277 5110 16367 5148
rect 16405 5110 16495 5148
rect 16533 5110 16623 5148
rect 16661 5110 16751 5148
rect 16789 5110 16879 5148
rect 16917 5110 17007 5148
rect 17045 5110 17135 5148
rect 17173 5110 17263 5148
rect 17301 5110 17391 5148
rect 17429 5110 17519 5148
rect 17557 5110 17647 5148
rect 17685 5110 17775 5148
rect 17813 5110 17903 5148
rect 17941 5110 18031 5148
rect 18069 5110 18159 5148
rect 18197 5110 18287 5148
rect 18325 5110 18415 5148
rect 18453 5110 18543 5148
rect 18581 5110 18671 5148
rect 18709 5110 18799 5148
rect 18837 5110 18927 5148
rect 18965 5110 19055 5148
rect 19093 5110 19183 5148
rect 19221 5110 19311 5148
rect 19349 5110 20269 5148
rect 20307 5110 20397 5148
rect 20435 5110 20525 5148
rect 20563 5110 20653 5148
rect 20691 5110 20781 5148
rect 20819 5110 20909 5148
rect 20947 5110 21037 5148
rect 21075 5110 21165 5148
rect 21203 5110 21293 5148
rect 21331 5110 21421 5148
rect 21459 5110 21549 5148
rect 21587 5110 21677 5148
rect 21715 5110 21805 5148
rect 21843 5110 21933 5148
rect 21971 5110 22061 5148
rect 22099 5110 22189 5148
rect 22227 5110 22317 5148
rect 22355 5110 22445 5148
rect 22483 5110 22573 5148
rect 22611 5110 22701 5148
rect 22739 5110 22829 5148
rect 22867 5110 22957 5148
rect 22995 5110 23085 5148
rect 23123 5110 23213 5148
rect 23251 5110 23341 5148
rect 23379 5110 23469 5148
rect 23507 5110 23597 5148
rect 23635 5110 23725 5148
rect 23763 5110 23853 5148
rect 23891 5110 23981 5148
rect 24019 5110 24109 5148
rect 24147 5110 24237 5148
rect 24275 5110 24365 5148
rect 24403 5110 24493 5148
rect 24531 5110 24621 5148
rect 24659 5110 24749 5148
rect 24787 5110 24877 5148
rect 24915 5110 25005 5148
rect 25043 5110 25133 5148
rect 25171 5110 25261 5148
rect 25299 5110 25389 5148
rect 25427 5110 25517 5148
rect 25555 5110 25645 5148
rect 25683 5110 25773 5148
rect 25811 5110 25901 5148
rect 25939 5110 26029 5148
rect 26067 5110 26157 5148
rect 26195 5110 26285 5148
rect 26323 5110 26413 5148
rect 26451 5110 26541 5148
rect 26579 5110 26669 5148
rect 26707 5110 26797 5148
rect 26835 5110 26925 5148
rect 26963 5110 27053 5148
rect 27091 5110 27181 5148
rect 27219 5110 27309 5148
rect 27347 5110 27437 5148
rect 27475 5110 27565 5148
rect 27603 5110 27693 5148
rect 27731 5110 27821 5148
rect 27859 5110 27949 5148
rect 27987 5110 28077 5148
rect 28115 5110 28205 5148
rect 28243 5110 28333 5148
rect 28371 5110 28461 5148
rect 28499 5110 28543 5148
rect 3448 5106 28543 5110
rect 675 4600 713 4678
rect 1587 4600 1625 4678
rect 2193 4600 2231 4678
rect 3121 4600 3159 4678
rect 3727 4600 3765 4678
rect 4333 4600 4371 4678
rect 4939 4600 4977 4678
rect 5672 4600 5710 4678
rect 6278 4600 6316 4678
rect 6884 4600 6922 4678
rect 7490 4600 7528 4678
rect 8096 4600 8134 4678
rect 8702 4600 8740 4678
rect 9308 4600 9346 4678
rect 9914 4600 9952 4678
rect 10646 4600 10684 4678
rect 11252 4600 11290 4678
rect 11858 4600 11896 4678
rect 12464 4600 12502 4678
rect 13070 4600 13108 4678
rect 13676 4600 13714 4678
rect 14282 4600 14320 4678
rect 14888 4600 14926 4678
rect 15494 4600 15532 4678
rect 16100 4600 16138 4678
rect 16706 4600 16744 4678
rect 17312 4600 17350 4678
rect 17918 4600 17956 4678
rect 18524 4600 18562 4678
rect 19130 4600 19168 4678
rect 19736 4600 19774 4678
rect 20468 4600 20506 4678
rect 21074 4600 21112 4678
rect 21680 4600 21718 4678
rect 22286 4600 22324 4678
rect 22892 4600 22930 4678
rect 23498 4600 23536 4678
rect 24104 4600 24142 4678
rect 24710 4600 24748 4678
rect 25316 4600 25354 4678
rect 25922 4600 25960 4678
rect 26528 4600 26566 4678
rect 27134 4600 27172 4678
rect 27740 4600 27778 4678
rect 28346 4600 28384 4678
rect 28952 4600 28990 4678
rect 29558 4600 29596 4678
rect 30164 4600 30202 4678
rect 30770 4600 30808 4678
rect 31376 4600 31414 4678
rect 31982 4600 32020 4678
rect 32588 4600 32626 4678
rect 33194 4600 33232 4678
rect 33800 4600 33838 4678
rect 34406 4600 34444 4678
rect 35012 4600 35050 4678
rect 35618 4600 35656 4678
rect 36224 4600 36262 4678
rect 36830 4600 36868 4678
rect 37436 4600 37474 4678
rect 38042 4600 38080 4678
rect 38648 4600 38686 4678
rect 39254 4600 39292 4678
rect -145 4282 -107 4360
rect 7850 3958 7894 4040
rect 669 3615 717 3729
rect 2069 3708 2109 3818
rect 4207 3754 4251 3854
rect 14766 3754 14810 3846
rect 29070 3542 29112 3632
rect -139 3440 -101 3518
rect 669 3122 707 3200
rect 1581 3122 1619 3200
rect 2187 3122 2225 3200
rect 3115 3122 3153 3200
rect 3721 3122 3759 3200
rect 4327 3122 4365 3200
rect 4933 3122 4971 3200
rect 5666 3122 5704 3200
rect 6272 3122 6310 3200
rect 6878 3122 6916 3200
rect 7484 3122 7522 3200
rect 8090 3122 8128 3200
rect 8696 3122 8734 3200
rect 9302 3122 9340 3200
rect 9908 3122 9946 3200
rect 10640 3122 10678 3200
rect 11246 3122 11284 3200
rect 11852 3122 11890 3200
rect 12458 3122 12496 3200
rect 13064 3122 13102 3200
rect 13670 3122 13708 3200
rect 14276 3122 14314 3200
rect 14882 3122 14920 3200
rect 15488 3122 15526 3200
rect 16094 3122 16132 3200
rect 16700 3122 16738 3200
rect 17306 3122 17344 3200
rect 17912 3122 17950 3200
rect 18518 3122 18556 3200
rect 19124 3122 19162 3200
rect 19730 3122 19768 3200
rect 20462 3122 20500 3200
rect 21068 3122 21106 3200
rect 21674 3122 21712 3200
rect 22280 3122 22318 3200
rect 22886 3122 22924 3200
rect 23492 3122 23530 3200
rect 24098 3122 24136 3200
rect 24704 3122 24742 3200
rect 25310 3122 25348 3200
rect 25916 3122 25954 3200
rect 26522 3122 26560 3200
rect 27128 3122 27166 3200
rect 27734 3122 27772 3200
rect 28340 3122 28378 3200
rect 28946 3122 28984 3200
rect 29552 3122 29590 3200
rect 30158 3122 30196 3200
rect 30764 3122 30802 3200
rect 31370 3122 31408 3200
rect 31976 3122 32014 3200
rect 32582 3122 32620 3200
rect 33188 3122 33226 3200
rect 33794 3122 33832 3200
rect 34400 3122 34438 3200
rect 35006 3122 35044 3200
rect 35612 3122 35650 3200
rect 36218 3122 36256 3200
rect 36824 3122 36862 3200
rect 37430 3122 37468 3200
rect 38036 3122 38074 3200
rect 38642 3122 38680 3200
rect 39248 3122 39286 3200
rect 675 2112 713 2190
rect 1587 2112 1625 2190
rect 2193 2112 2231 2190
rect 3121 2112 3159 2190
rect 3727 2112 3765 2190
rect 4333 2112 4371 2190
rect 4939 2112 4977 2190
rect 5672 2112 5710 2190
rect 6278 2112 6316 2190
rect 6884 2112 6922 2190
rect 7490 2112 7528 2190
rect 8096 2112 8134 2190
rect 8702 2112 8740 2190
rect 9308 2112 9346 2190
rect 9914 2112 9952 2190
rect 10646 2112 10684 2190
rect 11252 2112 11290 2190
rect 11858 2112 11896 2190
rect 12464 2112 12502 2190
rect 13070 2112 13108 2190
rect 13676 2112 13714 2190
rect 14282 2112 14320 2190
rect 14888 2112 14926 2190
rect 15494 2112 15532 2190
rect 16100 2112 16138 2190
rect 16706 2112 16744 2190
rect 17312 2112 17350 2190
rect 17918 2112 17956 2190
rect 18524 2112 18562 2190
rect 19130 2112 19168 2190
rect 19736 2112 19774 2190
rect 20468 2112 20506 2190
rect 21074 2112 21112 2190
rect 21680 2112 21718 2190
rect 22286 2112 22324 2190
rect 22892 2112 22930 2190
rect 23498 2112 23536 2190
rect 24104 2112 24142 2190
rect 24710 2112 24748 2190
rect 25316 2112 25354 2190
rect 25922 2112 25960 2190
rect 26528 2112 26566 2190
rect 27134 2112 27172 2190
rect 27740 2112 27778 2190
rect 28346 2112 28384 2190
rect 28952 2112 28990 2190
rect 29558 2112 29596 2190
rect 30164 2112 30202 2190
rect 30770 2112 30808 2190
rect 31376 2112 31414 2190
rect 31982 2112 32020 2190
rect 32588 2112 32626 2190
rect 33194 2112 33232 2190
rect 33800 2112 33838 2190
rect 34406 2112 34444 2190
rect 35012 2112 35050 2190
rect 35618 2112 35656 2190
rect 36224 2112 36262 2190
rect 36830 2112 36868 2190
rect 37436 2112 37474 2190
rect 38042 2112 38080 2190
rect 38648 2112 38686 2190
rect 39254 2112 39292 2190
rect -145 1794 -107 1872
rect 7850 1470 7894 1552
rect 669 1127 717 1241
rect 2069 1220 2109 1330
rect 4207 1266 4251 1366
rect 14766 1266 14810 1358
rect 29070 1054 29112 1144
rect -139 952 -101 1030
rect 669 634 707 712
rect 1581 634 1619 712
rect 2187 634 2225 712
rect 3115 634 3153 712
rect 3721 634 3759 712
rect 4327 634 4365 712
rect 4933 634 4971 712
rect 5666 634 5704 712
rect 6272 634 6310 712
rect 6878 634 6916 712
rect 7484 634 7522 712
rect 8090 634 8128 712
rect 8696 634 8734 712
rect 9302 634 9340 712
rect 9908 634 9946 712
rect 10640 634 10678 712
rect 11246 634 11284 712
rect 11852 634 11890 712
rect 12458 634 12496 712
rect 13064 634 13102 712
rect 13670 634 13708 712
rect 14276 634 14314 712
rect 14882 634 14920 712
rect 15488 634 15526 712
rect 16094 634 16132 712
rect 16700 634 16738 712
rect 17306 634 17344 712
rect 17912 634 17950 712
rect 18518 634 18556 712
rect 19124 634 19162 712
rect 19730 634 19768 712
rect 20462 634 20500 712
rect 21068 634 21106 712
rect 21674 634 21712 712
rect 22280 634 22318 712
rect 22886 634 22924 712
rect 23492 634 23530 712
rect 24098 634 24136 712
rect 24704 634 24742 712
rect 25310 634 25348 712
rect 25916 634 25954 712
rect 26522 634 26560 712
rect 27128 634 27166 712
rect 27734 634 27772 712
rect 28340 634 28378 712
rect 28946 634 28984 712
rect 29552 634 29590 712
rect 30158 634 30196 712
rect 30764 634 30802 712
rect 31370 634 31408 712
rect 31976 634 32014 712
rect 32582 634 32620 712
rect 33188 634 33226 712
rect 33794 634 33832 712
rect 34400 634 34438 712
rect 35006 634 35044 712
rect 35612 634 35650 712
rect 36218 634 36256 712
rect 36824 634 36862 712
rect 37430 634 37468 712
rect 38036 634 38074 712
rect 38642 634 38680 712
rect 39248 634 39286 712
<< nsubdiff >>
rect -341 6416 -87 6420
rect -341 6378 -297 6416
rect -259 6378 -169 6416
rect -131 6378 -87 6416
rect -341 6374 -87 6378
rect 436 6416 818 6420
rect 436 6378 480 6416
rect 518 6378 608 6416
rect 646 6378 736 6416
rect 774 6378 818 6416
rect 436 6374 818 6378
rect 1345 6416 1983 6420
rect 1345 6378 1389 6416
rect 1427 6378 1517 6416
rect 1555 6378 1645 6416
rect 1683 6378 1773 6416
rect 1811 6378 1901 6416
rect 1939 6378 1983 6416
rect 1345 6374 1983 6378
rect 2878 6416 4028 6420
rect 2878 6378 2922 6416
rect 2960 6378 3050 6416
rect 3088 6378 3178 6416
rect 3216 6378 3306 6416
rect 3344 6378 3434 6416
rect 3472 6378 3562 6416
rect 3600 6378 3690 6416
rect 3728 6378 3818 6416
rect 3856 6378 3946 6416
rect 3984 6378 4028 6416
rect 2878 6374 4028 6378
rect 5429 6416 7603 6420
rect 5429 6378 5473 6416
rect 5511 6378 5601 6416
rect 5639 6378 5729 6416
rect 5767 6378 5857 6416
rect 5895 6378 5985 6416
rect 6023 6378 6113 6416
rect 6151 6378 6241 6416
rect 6279 6378 6369 6416
rect 6407 6378 6497 6416
rect 6535 6378 6625 6416
rect 6663 6378 6753 6416
rect 6791 6378 6881 6416
rect 6919 6378 7009 6416
rect 7047 6378 7137 6416
rect 7175 6378 7265 6416
rect 7303 6378 7393 6416
rect 7431 6378 7521 6416
rect 7559 6378 7603 6416
rect 5429 6374 7603 6378
rect 10516 6416 14738 6420
rect 10516 6378 10560 6416
rect 10598 6378 10688 6416
rect 10726 6378 10816 6416
rect 10854 6378 10944 6416
rect 10982 6378 11072 6416
rect 11110 6378 11200 6416
rect 11238 6378 11328 6416
rect 11366 6378 11456 6416
rect 11494 6378 11584 6416
rect 11622 6378 11712 6416
rect 11750 6378 11840 6416
rect 11878 6378 11968 6416
rect 12006 6378 12096 6416
rect 12134 6378 12224 6416
rect 12262 6378 12352 6416
rect 12390 6378 12480 6416
rect 12518 6378 12608 6416
rect 12646 6378 12736 6416
rect 12774 6378 12864 6416
rect 12902 6378 12992 6416
rect 13030 6378 13120 6416
rect 13158 6378 13248 6416
rect 13286 6378 13376 6416
rect 13414 6378 13504 6416
rect 13542 6378 13632 6416
rect 13670 6378 13760 6416
rect 13798 6378 13888 6416
rect 13926 6378 14016 6416
rect 14054 6378 14144 6416
rect 14182 6378 14272 6416
rect 14310 6378 14400 6416
rect 14438 6378 14528 6416
rect 14566 6378 14656 6416
rect 14694 6378 14738 6416
rect 10516 6374 14738 6378
rect 20301 6416 28619 6420
rect 20301 6378 20345 6416
rect 20383 6378 20473 6416
rect 20511 6378 20601 6416
rect 20639 6378 20729 6416
rect 20767 6378 20857 6416
rect 20895 6378 20985 6416
rect 21023 6378 21113 6416
rect 21151 6378 21241 6416
rect 21279 6378 21369 6416
rect 21407 6378 21497 6416
rect 21535 6378 21625 6416
rect 21663 6378 21753 6416
rect 21791 6378 21881 6416
rect 21919 6378 22009 6416
rect 22047 6378 22137 6416
rect 22175 6378 22265 6416
rect 22303 6378 22393 6416
rect 22431 6378 22521 6416
rect 22559 6378 22649 6416
rect 22687 6378 22777 6416
rect 22815 6378 22905 6416
rect 22943 6378 23033 6416
rect 23071 6378 23161 6416
rect 23199 6378 23289 6416
rect 23327 6378 23417 6416
rect 23455 6378 23545 6416
rect 23583 6378 23673 6416
rect 23711 6378 23801 6416
rect 23839 6378 23929 6416
rect 23967 6378 24057 6416
rect 24095 6378 24185 6416
rect 24223 6378 24313 6416
rect 24351 6378 24441 6416
rect 24479 6378 24569 6416
rect 24607 6378 24697 6416
rect 24735 6378 24825 6416
rect 24863 6378 24953 6416
rect 24991 6378 25081 6416
rect 25119 6378 25209 6416
rect 25247 6378 25337 6416
rect 25375 6378 25465 6416
rect 25503 6378 25593 6416
rect 25631 6378 25721 6416
rect 25759 6378 25849 6416
rect 25887 6378 25977 6416
rect 26015 6378 26105 6416
rect 26143 6378 26233 6416
rect 26271 6378 26361 6416
rect 26399 6378 26489 6416
rect 26527 6378 26617 6416
rect 26655 6378 26745 6416
rect 26783 6378 26873 6416
rect 26911 6378 27001 6416
rect 27039 6378 27129 6416
rect 27167 6378 27257 6416
rect 27295 6378 27385 6416
rect 27423 6378 27513 6416
rect 27551 6378 27641 6416
rect 27679 6378 27769 6416
rect 27807 6378 27897 6416
rect 27935 6378 28025 6416
rect 28063 6378 28153 6416
rect 28191 6378 28281 6416
rect 28319 6378 28409 6416
rect 28447 6378 28537 6416
rect 28575 6378 28619 6416
rect 20301 6374 28619 6378
rect -363 5728 -109 5732
rect -363 5690 -319 5728
rect -281 5690 -191 5728
rect -153 5690 -109 5728
rect -363 5686 -109 5690
rect 565 5728 947 5732
rect 565 5690 609 5728
rect 647 5690 737 5728
rect 775 5690 865 5728
rect 903 5690 947 5728
rect 565 5686 947 5690
rect 1829 5728 2467 5732
rect 1829 5690 1873 5728
rect 1911 5690 2001 5728
rect 2039 5690 2129 5728
rect 2167 5690 2257 5728
rect 2295 5690 2385 5728
rect 2423 5690 2467 5728
rect 1829 5686 2467 5690
rect 3448 5728 4598 5732
rect 3448 5690 3492 5728
rect 3530 5690 3620 5728
rect 3658 5690 3748 5728
rect 3786 5690 3876 5728
rect 3914 5690 4004 5728
rect 4042 5690 4132 5728
rect 4170 5690 4260 5728
rect 4298 5690 4388 5728
rect 4426 5690 4516 5728
rect 4554 5690 4598 5728
rect 3448 5686 4598 5690
rect 8013 5728 10187 5732
rect 8013 5690 8057 5728
rect 8095 5690 8185 5728
rect 8223 5690 8313 5728
rect 8351 5690 8441 5728
rect 8479 5690 8569 5728
rect 8607 5690 8697 5728
rect 8735 5690 8825 5728
rect 8863 5690 8953 5728
rect 8991 5690 9081 5728
rect 9119 5690 9209 5728
rect 9247 5690 9337 5728
rect 9375 5690 9465 5728
rect 9503 5690 9593 5728
rect 9631 5690 9721 5728
rect 9759 5690 9849 5728
rect 9887 5690 9977 5728
rect 10015 5690 10105 5728
rect 10143 5690 10187 5728
rect 8013 5686 10187 5690
rect 15171 5728 19393 5732
rect 15171 5690 15215 5728
rect 15253 5690 15343 5728
rect 15381 5690 15471 5728
rect 15509 5690 15599 5728
rect 15637 5690 15727 5728
rect 15765 5690 15855 5728
rect 15893 5690 15983 5728
rect 16021 5690 16111 5728
rect 16149 5690 16239 5728
rect 16277 5690 16367 5728
rect 16405 5690 16495 5728
rect 16533 5690 16623 5728
rect 16661 5690 16751 5728
rect 16789 5690 16879 5728
rect 16917 5690 17007 5728
rect 17045 5690 17135 5728
rect 17173 5690 17263 5728
rect 17301 5690 17391 5728
rect 17429 5690 17519 5728
rect 17557 5690 17647 5728
rect 17685 5690 17775 5728
rect 17813 5690 17903 5728
rect 17941 5690 18031 5728
rect 18069 5690 18159 5728
rect 18197 5690 18287 5728
rect 18325 5690 18415 5728
rect 18453 5690 18543 5728
rect 18581 5690 18671 5728
rect 18709 5690 18799 5728
rect 18837 5690 18927 5728
rect 18965 5690 19055 5728
rect 19093 5690 19183 5728
rect 19221 5690 19311 5728
rect 19349 5690 19393 5728
rect 15171 5686 19393 5690
rect 20225 5728 28543 5732
rect 20225 5690 20269 5728
rect 20307 5690 20397 5728
rect 20435 5690 20525 5728
rect 20563 5690 20653 5728
rect 20691 5690 20781 5728
rect 20819 5690 20909 5728
rect 20947 5690 21037 5728
rect 21075 5690 21165 5728
rect 21203 5690 21293 5728
rect 21331 5690 21421 5728
rect 21459 5690 21549 5728
rect 21587 5690 21677 5728
rect 21715 5690 21805 5728
rect 21843 5690 21933 5728
rect 21971 5690 22061 5728
rect 22099 5690 22189 5728
rect 22227 5690 22317 5728
rect 22355 5690 22445 5728
rect 22483 5690 22573 5728
rect 22611 5690 22701 5728
rect 22739 5690 22829 5728
rect 22867 5690 22957 5728
rect 22995 5690 23085 5728
rect 23123 5690 23213 5728
rect 23251 5690 23341 5728
rect 23379 5690 23469 5728
rect 23507 5690 23597 5728
rect 23635 5690 23725 5728
rect 23763 5690 23853 5728
rect 23891 5690 23981 5728
rect 24019 5690 24109 5728
rect 24147 5690 24237 5728
rect 24275 5690 24365 5728
rect 24403 5690 24493 5728
rect 24531 5690 24621 5728
rect 24659 5690 24749 5728
rect 24787 5690 24877 5728
rect 24915 5690 25005 5728
rect 25043 5690 25133 5728
rect 25171 5690 25261 5728
rect 25299 5690 25389 5728
rect 25427 5690 25517 5728
rect 25555 5690 25645 5728
rect 25683 5690 25773 5728
rect 25811 5690 25901 5728
rect 25939 5690 26029 5728
rect 26067 5690 26157 5728
rect 26195 5690 26285 5728
rect 26323 5690 26413 5728
rect 26451 5690 26541 5728
rect 26579 5690 26669 5728
rect 26707 5690 26797 5728
rect 26835 5690 26925 5728
rect 26963 5690 27053 5728
rect 27091 5690 27181 5728
rect 27219 5690 27309 5728
rect 27347 5690 27437 5728
rect 27475 5690 27565 5728
rect 27603 5690 27693 5728
rect 27731 5690 27821 5728
rect 27859 5690 27949 5728
rect 27987 5690 28077 5728
rect 28115 5690 28205 5728
rect 28243 5690 28333 5728
rect 28371 5690 28461 5728
rect 28499 5690 28543 5728
rect 20225 5686 28543 5690
<< psubdiffcont >>
rect -297 5798 -259 5836
rect -169 5798 -131 5836
rect 480 5798 518 5836
rect 608 5798 646 5836
rect 736 5798 774 5836
rect 1389 5798 1427 5836
rect 1517 5798 1555 5836
rect 1645 5798 1683 5836
rect 1773 5798 1811 5836
rect 1901 5798 1939 5836
rect 2922 5798 2960 5836
rect 3050 5798 3088 5836
rect 3178 5798 3216 5836
rect 3306 5798 3344 5836
rect 3434 5798 3472 5836
rect 3562 5798 3600 5836
rect 3690 5798 3728 5836
rect 3818 5798 3856 5836
rect 3946 5798 3984 5836
rect 5473 5798 5511 5836
rect 5601 5798 5639 5836
rect 5729 5798 5767 5836
rect 5857 5798 5895 5836
rect 5985 5798 6023 5836
rect 6113 5798 6151 5836
rect 6241 5798 6279 5836
rect 6369 5798 6407 5836
rect 6497 5798 6535 5836
rect 6625 5798 6663 5836
rect 6753 5798 6791 5836
rect 6881 5798 6919 5836
rect 7009 5798 7047 5836
rect 7137 5798 7175 5836
rect 7265 5798 7303 5836
rect 7393 5798 7431 5836
rect 7521 5798 7559 5836
rect 10560 5798 10598 5836
rect 10688 5798 10726 5836
rect 10816 5798 10854 5836
rect 10944 5798 10982 5836
rect 11072 5798 11110 5836
rect 11200 5798 11238 5836
rect 11328 5798 11366 5836
rect 11456 5798 11494 5836
rect 11584 5798 11622 5836
rect 11712 5798 11750 5836
rect 11840 5798 11878 5836
rect 11968 5798 12006 5836
rect 12096 5798 12134 5836
rect 12224 5798 12262 5836
rect 12352 5798 12390 5836
rect 12480 5798 12518 5836
rect 12608 5798 12646 5836
rect 12736 5798 12774 5836
rect 12864 5798 12902 5836
rect 12992 5798 13030 5836
rect 13120 5798 13158 5836
rect 13248 5798 13286 5836
rect 13376 5798 13414 5836
rect 13504 5798 13542 5836
rect 13632 5798 13670 5836
rect 13760 5798 13798 5836
rect 13888 5798 13926 5836
rect 14016 5798 14054 5836
rect 14144 5798 14182 5836
rect 14272 5798 14310 5836
rect 14400 5798 14438 5836
rect 14528 5798 14566 5836
rect 14656 5798 14694 5836
rect 20345 5798 20383 5836
rect 20473 5798 20511 5836
rect 20601 5798 20639 5836
rect 20729 5798 20767 5836
rect 20857 5798 20895 5836
rect 20985 5798 21023 5836
rect 21113 5798 21151 5836
rect 21241 5798 21279 5836
rect 21369 5798 21407 5836
rect 21497 5798 21535 5836
rect 21625 5798 21663 5836
rect 21753 5798 21791 5836
rect 21881 5798 21919 5836
rect 22009 5798 22047 5836
rect 22137 5798 22175 5836
rect 22265 5798 22303 5836
rect 22393 5798 22431 5836
rect 22521 5798 22559 5836
rect 22649 5798 22687 5836
rect 22777 5798 22815 5836
rect 22905 5798 22943 5836
rect 23033 5798 23071 5836
rect 23161 5798 23199 5836
rect 23289 5798 23327 5836
rect 23417 5798 23455 5836
rect 23545 5798 23583 5836
rect 23673 5798 23711 5836
rect 23801 5798 23839 5836
rect 23929 5798 23967 5836
rect 24057 5798 24095 5836
rect 24185 5798 24223 5836
rect 24313 5798 24351 5836
rect 24441 5798 24479 5836
rect 24569 5798 24607 5836
rect 24697 5798 24735 5836
rect 24825 5798 24863 5836
rect 24953 5798 24991 5836
rect 25081 5798 25119 5836
rect 25209 5798 25247 5836
rect 25337 5798 25375 5836
rect 25465 5798 25503 5836
rect 25593 5798 25631 5836
rect 25721 5798 25759 5836
rect 25849 5798 25887 5836
rect 25977 5798 26015 5836
rect 26105 5798 26143 5836
rect 26233 5798 26271 5836
rect 26361 5798 26399 5836
rect 26489 5798 26527 5836
rect 26617 5798 26655 5836
rect 26745 5798 26783 5836
rect 26873 5798 26911 5836
rect 27001 5798 27039 5836
rect 27129 5798 27167 5836
rect 27257 5798 27295 5836
rect 27385 5798 27423 5836
rect 27513 5798 27551 5836
rect 27641 5798 27679 5836
rect 27769 5798 27807 5836
rect 27897 5798 27935 5836
rect 28025 5798 28063 5836
rect 28153 5798 28191 5836
rect 28281 5798 28319 5836
rect 28409 5798 28447 5836
rect 28537 5798 28575 5836
rect -319 5110 -281 5148
rect -191 5110 -153 5148
rect 609 5110 647 5148
rect 737 5110 775 5148
rect 865 5110 903 5148
rect 1873 5110 1911 5148
rect 2001 5110 2039 5148
rect 2129 5110 2167 5148
rect 2257 5110 2295 5148
rect 2385 5110 2423 5148
rect 3492 5110 3530 5148
rect 3620 5110 3658 5148
rect 3748 5110 3786 5148
rect 3876 5110 3914 5148
rect 4004 5110 4042 5148
rect 4132 5110 4170 5148
rect 4260 5110 4298 5148
rect 4388 5110 4426 5148
rect 4516 5110 4554 5148
rect 8057 5110 8095 5148
rect 8185 5110 8223 5148
rect 8313 5110 8351 5148
rect 8441 5110 8479 5148
rect 8569 5110 8607 5148
rect 8697 5110 8735 5148
rect 8825 5110 8863 5148
rect 8953 5110 8991 5148
rect 9081 5110 9119 5148
rect 9209 5110 9247 5148
rect 9337 5110 9375 5148
rect 9465 5110 9503 5148
rect 9593 5110 9631 5148
rect 9721 5110 9759 5148
rect 9849 5110 9887 5148
rect 9977 5110 10015 5148
rect 10105 5110 10143 5148
rect 15215 5110 15253 5148
rect 15343 5110 15381 5148
rect 15471 5110 15509 5148
rect 15599 5110 15637 5148
rect 15727 5110 15765 5148
rect 15855 5110 15893 5148
rect 15983 5110 16021 5148
rect 16111 5110 16149 5148
rect 16239 5110 16277 5148
rect 16367 5110 16405 5148
rect 16495 5110 16533 5148
rect 16623 5110 16661 5148
rect 16751 5110 16789 5148
rect 16879 5110 16917 5148
rect 17007 5110 17045 5148
rect 17135 5110 17173 5148
rect 17263 5110 17301 5148
rect 17391 5110 17429 5148
rect 17519 5110 17557 5148
rect 17647 5110 17685 5148
rect 17775 5110 17813 5148
rect 17903 5110 17941 5148
rect 18031 5110 18069 5148
rect 18159 5110 18197 5148
rect 18287 5110 18325 5148
rect 18415 5110 18453 5148
rect 18543 5110 18581 5148
rect 18671 5110 18709 5148
rect 18799 5110 18837 5148
rect 18927 5110 18965 5148
rect 19055 5110 19093 5148
rect 19183 5110 19221 5148
rect 19311 5110 19349 5148
rect 20269 5110 20307 5148
rect 20397 5110 20435 5148
rect 20525 5110 20563 5148
rect 20653 5110 20691 5148
rect 20781 5110 20819 5148
rect 20909 5110 20947 5148
rect 21037 5110 21075 5148
rect 21165 5110 21203 5148
rect 21293 5110 21331 5148
rect 21421 5110 21459 5148
rect 21549 5110 21587 5148
rect 21677 5110 21715 5148
rect 21805 5110 21843 5148
rect 21933 5110 21971 5148
rect 22061 5110 22099 5148
rect 22189 5110 22227 5148
rect 22317 5110 22355 5148
rect 22445 5110 22483 5148
rect 22573 5110 22611 5148
rect 22701 5110 22739 5148
rect 22829 5110 22867 5148
rect 22957 5110 22995 5148
rect 23085 5110 23123 5148
rect 23213 5110 23251 5148
rect 23341 5110 23379 5148
rect 23469 5110 23507 5148
rect 23597 5110 23635 5148
rect 23725 5110 23763 5148
rect 23853 5110 23891 5148
rect 23981 5110 24019 5148
rect 24109 5110 24147 5148
rect 24237 5110 24275 5148
rect 24365 5110 24403 5148
rect 24493 5110 24531 5148
rect 24621 5110 24659 5148
rect 24749 5110 24787 5148
rect 24877 5110 24915 5148
rect 25005 5110 25043 5148
rect 25133 5110 25171 5148
rect 25261 5110 25299 5148
rect 25389 5110 25427 5148
rect 25517 5110 25555 5148
rect 25645 5110 25683 5148
rect 25773 5110 25811 5148
rect 25901 5110 25939 5148
rect 26029 5110 26067 5148
rect 26157 5110 26195 5148
rect 26285 5110 26323 5148
rect 26413 5110 26451 5148
rect 26541 5110 26579 5148
rect 26669 5110 26707 5148
rect 26797 5110 26835 5148
rect 26925 5110 26963 5148
rect 27053 5110 27091 5148
rect 27181 5110 27219 5148
rect 27309 5110 27347 5148
rect 27437 5110 27475 5148
rect 27565 5110 27603 5148
rect 27693 5110 27731 5148
rect 27821 5110 27859 5148
rect 27949 5110 27987 5148
rect 28077 5110 28115 5148
rect 28205 5110 28243 5148
rect 28333 5110 28371 5148
rect 28461 5110 28499 5148
<< nsubdiffcont >>
rect -297 6378 -259 6416
rect -169 6378 -131 6416
rect 480 6378 518 6416
rect 608 6378 646 6416
rect 736 6378 774 6416
rect 1389 6378 1427 6416
rect 1517 6378 1555 6416
rect 1645 6378 1683 6416
rect 1773 6378 1811 6416
rect 1901 6378 1939 6416
rect 2922 6378 2960 6416
rect 3050 6378 3088 6416
rect 3178 6378 3216 6416
rect 3306 6378 3344 6416
rect 3434 6378 3472 6416
rect 3562 6378 3600 6416
rect 3690 6378 3728 6416
rect 3818 6378 3856 6416
rect 3946 6378 3984 6416
rect 5473 6378 5511 6416
rect 5601 6378 5639 6416
rect 5729 6378 5767 6416
rect 5857 6378 5895 6416
rect 5985 6378 6023 6416
rect 6113 6378 6151 6416
rect 6241 6378 6279 6416
rect 6369 6378 6407 6416
rect 6497 6378 6535 6416
rect 6625 6378 6663 6416
rect 6753 6378 6791 6416
rect 6881 6378 6919 6416
rect 7009 6378 7047 6416
rect 7137 6378 7175 6416
rect 7265 6378 7303 6416
rect 7393 6378 7431 6416
rect 7521 6378 7559 6416
rect 10560 6378 10598 6416
rect 10688 6378 10726 6416
rect 10816 6378 10854 6416
rect 10944 6378 10982 6416
rect 11072 6378 11110 6416
rect 11200 6378 11238 6416
rect 11328 6378 11366 6416
rect 11456 6378 11494 6416
rect 11584 6378 11622 6416
rect 11712 6378 11750 6416
rect 11840 6378 11878 6416
rect 11968 6378 12006 6416
rect 12096 6378 12134 6416
rect 12224 6378 12262 6416
rect 12352 6378 12390 6416
rect 12480 6378 12518 6416
rect 12608 6378 12646 6416
rect 12736 6378 12774 6416
rect 12864 6378 12902 6416
rect 12992 6378 13030 6416
rect 13120 6378 13158 6416
rect 13248 6378 13286 6416
rect 13376 6378 13414 6416
rect 13504 6378 13542 6416
rect 13632 6378 13670 6416
rect 13760 6378 13798 6416
rect 13888 6378 13926 6416
rect 14016 6378 14054 6416
rect 14144 6378 14182 6416
rect 14272 6378 14310 6416
rect 14400 6378 14438 6416
rect 14528 6378 14566 6416
rect 14656 6378 14694 6416
rect 20345 6378 20383 6416
rect 20473 6378 20511 6416
rect 20601 6378 20639 6416
rect 20729 6378 20767 6416
rect 20857 6378 20895 6416
rect 20985 6378 21023 6416
rect 21113 6378 21151 6416
rect 21241 6378 21279 6416
rect 21369 6378 21407 6416
rect 21497 6378 21535 6416
rect 21625 6378 21663 6416
rect 21753 6378 21791 6416
rect 21881 6378 21919 6416
rect 22009 6378 22047 6416
rect 22137 6378 22175 6416
rect 22265 6378 22303 6416
rect 22393 6378 22431 6416
rect 22521 6378 22559 6416
rect 22649 6378 22687 6416
rect 22777 6378 22815 6416
rect 22905 6378 22943 6416
rect 23033 6378 23071 6416
rect 23161 6378 23199 6416
rect 23289 6378 23327 6416
rect 23417 6378 23455 6416
rect 23545 6378 23583 6416
rect 23673 6378 23711 6416
rect 23801 6378 23839 6416
rect 23929 6378 23967 6416
rect 24057 6378 24095 6416
rect 24185 6378 24223 6416
rect 24313 6378 24351 6416
rect 24441 6378 24479 6416
rect 24569 6378 24607 6416
rect 24697 6378 24735 6416
rect 24825 6378 24863 6416
rect 24953 6378 24991 6416
rect 25081 6378 25119 6416
rect 25209 6378 25247 6416
rect 25337 6378 25375 6416
rect 25465 6378 25503 6416
rect 25593 6378 25631 6416
rect 25721 6378 25759 6416
rect 25849 6378 25887 6416
rect 25977 6378 26015 6416
rect 26105 6378 26143 6416
rect 26233 6378 26271 6416
rect 26361 6378 26399 6416
rect 26489 6378 26527 6416
rect 26617 6378 26655 6416
rect 26745 6378 26783 6416
rect 26873 6378 26911 6416
rect 27001 6378 27039 6416
rect 27129 6378 27167 6416
rect 27257 6378 27295 6416
rect 27385 6378 27423 6416
rect 27513 6378 27551 6416
rect 27641 6378 27679 6416
rect 27769 6378 27807 6416
rect 27897 6378 27935 6416
rect 28025 6378 28063 6416
rect 28153 6378 28191 6416
rect 28281 6378 28319 6416
rect 28409 6378 28447 6416
rect 28537 6378 28575 6416
rect -319 5690 -281 5728
rect -191 5690 -153 5728
rect 609 5690 647 5728
rect 737 5690 775 5728
rect 865 5690 903 5728
rect 1873 5690 1911 5728
rect 2001 5690 2039 5728
rect 2129 5690 2167 5728
rect 2257 5690 2295 5728
rect 2385 5690 2423 5728
rect 3492 5690 3530 5728
rect 3620 5690 3658 5728
rect 3748 5690 3786 5728
rect 3876 5690 3914 5728
rect 4004 5690 4042 5728
rect 4132 5690 4170 5728
rect 4260 5690 4298 5728
rect 4388 5690 4426 5728
rect 4516 5690 4554 5728
rect 8057 5690 8095 5728
rect 8185 5690 8223 5728
rect 8313 5690 8351 5728
rect 8441 5690 8479 5728
rect 8569 5690 8607 5728
rect 8697 5690 8735 5728
rect 8825 5690 8863 5728
rect 8953 5690 8991 5728
rect 9081 5690 9119 5728
rect 9209 5690 9247 5728
rect 9337 5690 9375 5728
rect 9465 5690 9503 5728
rect 9593 5690 9631 5728
rect 9721 5690 9759 5728
rect 9849 5690 9887 5728
rect 9977 5690 10015 5728
rect 10105 5690 10143 5728
rect 15215 5690 15253 5728
rect 15343 5690 15381 5728
rect 15471 5690 15509 5728
rect 15599 5690 15637 5728
rect 15727 5690 15765 5728
rect 15855 5690 15893 5728
rect 15983 5690 16021 5728
rect 16111 5690 16149 5728
rect 16239 5690 16277 5728
rect 16367 5690 16405 5728
rect 16495 5690 16533 5728
rect 16623 5690 16661 5728
rect 16751 5690 16789 5728
rect 16879 5690 16917 5728
rect 17007 5690 17045 5728
rect 17135 5690 17173 5728
rect 17263 5690 17301 5728
rect 17391 5690 17429 5728
rect 17519 5690 17557 5728
rect 17647 5690 17685 5728
rect 17775 5690 17813 5728
rect 17903 5690 17941 5728
rect 18031 5690 18069 5728
rect 18159 5690 18197 5728
rect 18287 5690 18325 5728
rect 18415 5690 18453 5728
rect 18543 5690 18581 5728
rect 18671 5690 18709 5728
rect 18799 5690 18837 5728
rect 18927 5690 18965 5728
rect 19055 5690 19093 5728
rect 19183 5690 19221 5728
rect 19311 5690 19349 5728
rect 20269 5690 20307 5728
rect 20397 5690 20435 5728
rect 20525 5690 20563 5728
rect 20653 5690 20691 5728
rect 20781 5690 20819 5728
rect 20909 5690 20947 5728
rect 21037 5690 21075 5728
rect 21165 5690 21203 5728
rect 21293 5690 21331 5728
rect 21421 5690 21459 5728
rect 21549 5690 21587 5728
rect 21677 5690 21715 5728
rect 21805 5690 21843 5728
rect 21933 5690 21971 5728
rect 22061 5690 22099 5728
rect 22189 5690 22227 5728
rect 22317 5690 22355 5728
rect 22445 5690 22483 5728
rect 22573 5690 22611 5728
rect 22701 5690 22739 5728
rect 22829 5690 22867 5728
rect 22957 5690 22995 5728
rect 23085 5690 23123 5728
rect 23213 5690 23251 5728
rect 23341 5690 23379 5728
rect 23469 5690 23507 5728
rect 23597 5690 23635 5728
rect 23725 5690 23763 5728
rect 23853 5690 23891 5728
rect 23981 5690 24019 5728
rect 24109 5690 24147 5728
rect 24237 5690 24275 5728
rect 24365 5690 24403 5728
rect 24493 5690 24531 5728
rect 24621 5690 24659 5728
rect 24749 5690 24787 5728
rect 24877 5690 24915 5728
rect 25005 5690 25043 5728
rect 25133 5690 25171 5728
rect 25261 5690 25299 5728
rect 25389 5690 25427 5728
rect 25517 5690 25555 5728
rect 25645 5690 25683 5728
rect 25773 5690 25811 5728
rect 25901 5690 25939 5728
rect 26029 5690 26067 5728
rect 26157 5690 26195 5728
rect 26285 5690 26323 5728
rect 26413 5690 26451 5728
rect 26541 5690 26579 5728
rect 26669 5690 26707 5728
rect 26797 5690 26835 5728
rect 26925 5690 26963 5728
rect 27053 5690 27091 5728
rect 27181 5690 27219 5728
rect 27309 5690 27347 5728
rect 27437 5690 27475 5728
rect 27565 5690 27603 5728
rect 27693 5690 27731 5728
rect 27821 5690 27859 5728
rect 27949 5690 27987 5728
rect 28077 5690 28115 5728
rect 28205 5690 28243 5728
rect 28333 5690 28371 5728
rect 28461 5690 28499 5728
<< poly >>
rect -249 6278 -179 6309
rect 528 6278 598 6309
rect 656 6278 726 6309
rect 1437 6278 1507 6309
rect 1565 6278 1635 6309
rect 1693 6278 1763 6309
rect 1821 6278 1891 6309
rect 2970 6278 3040 6309
rect 3098 6278 3168 6309
rect 3226 6278 3296 6309
rect 3354 6278 3424 6309
rect 3482 6278 3552 6309
rect 3610 6278 3680 6309
rect 3738 6278 3808 6309
rect 3866 6278 3936 6309
rect 5521 6278 5591 6309
rect 5649 6278 5719 6309
rect 5777 6278 5847 6309
rect 5905 6278 5975 6309
rect 6033 6278 6103 6309
rect 6161 6278 6231 6309
rect 6289 6278 6359 6309
rect 6417 6278 6487 6309
rect 6545 6278 6615 6309
rect 6673 6278 6743 6309
rect 6801 6278 6871 6309
rect 6929 6278 6999 6309
rect 7057 6278 7127 6309
rect 7185 6278 7255 6309
rect 7313 6278 7383 6309
rect 7441 6278 7511 6309
rect 10608 6278 10678 6309
rect 10736 6278 10806 6309
rect 10864 6278 10934 6309
rect 10992 6278 11062 6309
rect 11120 6278 11190 6309
rect 11248 6278 11318 6309
rect 11376 6278 11446 6309
rect 11504 6278 11574 6309
rect 11632 6278 11702 6309
rect 11760 6278 11830 6309
rect 11888 6278 11958 6309
rect 12016 6278 12086 6309
rect 12144 6278 12214 6309
rect 12272 6278 12342 6309
rect 12400 6278 12470 6309
rect 12528 6278 12598 6309
rect 12656 6278 12726 6309
rect 12784 6278 12854 6309
rect 12912 6278 12982 6309
rect 13040 6278 13110 6309
rect 13168 6278 13238 6309
rect 13296 6278 13366 6309
rect 13424 6278 13494 6309
rect 13552 6278 13622 6309
rect 13680 6278 13750 6309
rect 13808 6278 13878 6309
rect 13936 6278 14006 6309
rect 14064 6278 14134 6309
rect 14192 6278 14262 6309
rect 14320 6278 14390 6309
rect 14448 6278 14518 6309
rect 14576 6278 14646 6309
rect 20393 6278 20463 6309
rect 20521 6278 20591 6309
rect 20649 6278 20719 6309
rect 20777 6278 20847 6309
rect 20905 6278 20975 6309
rect 21033 6278 21103 6309
rect 21161 6278 21231 6309
rect 21289 6278 21359 6309
rect 21417 6278 21487 6309
rect 21545 6278 21615 6309
rect 21673 6278 21743 6309
rect 21801 6278 21871 6309
rect 21929 6278 21999 6309
rect 22057 6278 22127 6309
rect 22185 6278 22255 6309
rect 22313 6278 22383 6309
rect 22441 6278 22511 6309
rect 22569 6278 22639 6309
rect 22697 6278 22767 6309
rect 22825 6278 22895 6309
rect 22953 6278 23023 6309
rect 23081 6278 23151 6309
rect 23209 6278 23279 6309
rect 23337 6278 23407 6309
rect 23465 6278 23535 6309
rect 23593 6278 23663 6309
rect 23721 6278 23791 6309
rect 23849 6278 23919 6309
rect 23977 6278 24047 6309
rect 24105 6278 24175 6309
rect 24233 6278 24303 6309
rect 24361 6278 24431 6309
rect 24489 6278 24559 6309
rect 24617 6278 24687 6309
rect 24745 6278 24815 6309
rect 24873 6278 24943 6309
rect 25001 6278 25071 6309
rect 25129 6278 25199 6309
rect 25257 6278 25327 6309
rect 25385 6278 25455 6309
rect 25513 6278 25583 6309
rect 25641 6278 25711 6309
rect 25769 6278 25839 6309
rect 25897 6278 25967 6309
rect 26025 6278 26095 6309
rect 26153 6278 26223 6309
rect 26281 6278 26351 6309
rect 26409 6278 26479 6309
rect 26537 6278 26607 6309
rect 26665 6278 26735 6309
rect 26793 6278 26863 6309
rect 26921 6278 26991 6309
rect 27049 6278 27119 6309
rect 27177 6278 27247 6309
rect 27305 6278 27375 6309
rect 27433 6278 27503 6309
rect 27561 6278 27631 6309
rect 27689 6278 27759 6309
rect 27817 6278 27887 6309
rect 27945 6278 28015 6309
rect 28073 6278 28143 6309
rect 28201 6278 28271 6309
rect 28329 6278 28399 6309
rect 28457 6278 28527 6309
rect -249 5978 -179 6110
rect 528 6093 598 6110
rect 656 6093 726 6110
rect 528 6023 726 6093
rect 528 5978 598 6023
rect 656 5978 726 6023
rect 1437 6093 1507 6110
rect 1565 6093 1635 6110
rect 1693 6093 1763 6110
rect 1821 6093 1891 6110
rect 1437 6023 1891 6093
rect 1437 5978 1507 6023
rect 1565 5978 1635 6023
rect 1693 5978 1763 6023
rect 1821 5978 1891 6023
rect 2970 6093 3040 6110
rect 3098 6093 3168 6110
rect 3226 6093 3296 6110
rect 3354 6093 3424 6110
rect 3482 6093 3552 6110
rect 3610 6093 3680 6110
rect 3738 6093 3808 6110
rect 3866 6093 3936 6110
rect 2970 6023 3936 6093
rect 2970 5978 3040 6023
rect 3098 5978 3168 6023
rect 3226 5978 3296 6023
rect 3354 5978 3424 6023
rect 3482 5978 3552 6023
rect 3610 5978 3680 6023
rect 3738 5978 3808 6023
rect 3866 5978 3936 6023
rect 5521 6093 5591 6110
rect 5649 6093 5719 6110
rect 5777 6093 5847 6110
rect 5905 6093 5975 6110
rect 6033 6093 6103 6110
rect 6161 6093 6231 6110
rect 6289 6093 6359 6110
rect 6417 6093 6487 6110
rect 6545 6093 6615 6110
rect 6673 6093 6743 6110
rect 6801 6093 6871 6110
rect 6929 6093 6999 6110
rect 7057 6093 7127 6110
rect 7185 6093 7255 6110
rect 7313 6093 7383 6110
rect 7441 6093 7511 6110
rect 5521 6023 7511 6093
rect 5521 5978 5591 6023
rect 5649 5978 5719 6023
rect 5777 5978 5847 6023
rect 5905 5978 5975 6023
rect 6033 5978 6103 6023
rect 6161 5978 6231 6023
rect 6289 5978 6359 6023
rect 6417 5978 6487 6023
rect 6545 5978 6615 6023
rect 6673 5978 6743 6023
rect 6801 5978 6871 6023
rect 6929 5978 6999 6023
rect 7057 5978 7127 6023
rect 7185 5978 7255 6023
rect 7313 5978 7383 6023
rect 7441 5978 7511 6023
rect 10608 6093 10678 6110
rect 10736 6093 10806 6110
rect 10864 6093 10934 6110
rect 10992 6093 11062 6110
rect 11120 6093 11190 6110
rect 11248 6093 11318 6110
rect 11376 6093 11446 6110
rect 11504 6093 11574 6110
rect 11632 6093 11702 6110
rect 11760 6093 11830 6110
rect 11888 6093 11958 6110
rect 12016 6093 12086 6110
rect 12144 6093 12214 6110
rect 12272 6093 12342 6110
rect 12400 6093 12470 6110
rect 12528 6093 12598 6110
rect 12656 6093 12726 6110
rect 12784 6093 12854 6110
rect 12912 6093 12982 6110
rect 13040 6093 13110 6110
rect 13168 6093 13238 6110
rect 13296 6093 13366 6110
rect 13424 6093 13494 6110
rect 13552 6093 13622 6110
rect 13680 6093 13750 6110
rect 13808 6093 13878 6110
rect 13936 6093 14006 6110
rect 14064 6093 14134 6110
rect 14192 6093 14262 6110
rect 14320 6093 14390 6110
rect 14448 6093 14518 6110
rect 14576 6093 14646 6110
rect 10608 6023 14646 6093
rect 10608 5978 10678 6023
rect 10736 5978 10806 6023
rect 10864 5978 10934 6023
rect 10992 5978 11062 6023
rect 11120 5978 11190 6023
rect 11248 5978 11318 6023
rect 11376 5978 11446 6023
rect 11504 5978 11574 6023
rect 11632 5978 11702 6023
rect 11760 5978 11830 6023
rect 11888 5978 11958 6023
rect 12016 5978 12086 6023
rect 12144 5978 12214 6023
rect 12272 5978 12342 6023
rect 12400 5978 12470 6023
rect 12528 5978 12598 6023
rect 12656 5978 12726 6023
rect 12784 5978 12854 6023
rect 12912 5978 12982 6023
rect 13040 5978 13110 6023
rect 13168 5978 13238 6023
rect 13296 5978 13366 6023
rect 13424 5978 13494 6023
rect 13552 5978 13622 6023
rect 13680 5978 13750 6023
rect 13808 5978 13878 6023
rect 13936 5978 14006 6023
rect 14064 5978 14134 6023
rect 14192 5978 14262 6023
rect 14320 5978 14390 6023
rect 14448 5978 14518 6023
rect 14576 5978 14646 6023
rect 20393 6093 20463 6110
rect 20521 6093 20591 6110
rect 20649 6093 20719 6110
rect 20777 6093 20847 6110
rect 20905 6093 20975 6110
rect 21033 6093 21103 6110
rect 21161 6093 21231 6110
rect 21289 6093 21359 6110
rect 21417 6093 21487 6110
rect 21545 6093 21615 6110
rect 21673 6093 21743 6110
rect 21801 6093 21871 6110
rect 21929 6093 21999 6110
rect 22057 6093 22127 6110
rect 22185 6093 22255 6110
rect 22313 6093 22383 6110
rect 22441 6093 22511 6110
rect 22569 6093 22639 6110
rect 22697 6093 22767 6110
rect 22825 6093 22895 6110
rect 22953 6093 23023 6110
rect 23081 6093 23151 6110
rect 23209 6093 23279 6110
rect 23337 6093 23407 6110
rect 23465 6093 23535 6110
rect 23593 6093 23663 6110
rect 23721 6093 23791 6110
rect 23849 6093 23919 6110
rect 23977 6093 24047 6110
rect 24105 6093 24175 6110
rect 24233 6093 24303 6110
rect 24361 6093 24431 6110
rect 24489 6093 24559 6110
rect 24617 6093 24687 6110
rect 24745 6093 24815 6110
rect 24873 6093 24943 6110
rect 25001 6093 25071 6110
rect 25129 6093 25199 6110
rect 25257 6093 25327 6110
rect 25385 6093 25455 6110
rect 25513 6093 25583 6110
rect 25641 6093 25711 6110
rect 25769 6093 25839 6110
rect 25897 6093 25967 6110
rect 26025 6093 26095 6110
rect 26153 6093 26223 6110
rect 26281 6093 26351 6110
rect 26409 6093 26479 6110
rect 26537 6093 26607 6110
rect 26665 6093 26735 6110
rect 26793 6093 26863 6110
rect 26921 6093 26991 6110
rect 27049 6093 27119 6110
rect 27177 6093 27247 6110
rect 27305 6093 27375 6110
rect 27433 6093 27503 6110
rect 27561 6093 27631 6110
rect 27689 6093 27759 6110
rect 27817 6093 27887 6110
rect 27945 6093 28015 6110
rect 28073 6093 28143 6110
rect 28201 6093 28271 6110
rect 28329 6093 28399 6110
rect 28457 6093 28527 6110
rect 20393 6023 28527 6093
rect 20393 5978 20463 6023
rect 20521 5978 20591 6023
rect 20649 5978 20719 6023
rect 20777 5978 20847 6023
rect 20905 5978 20975 6023
rect 21033 5978 21103 6023
rect 21161 5978 21231 6023
rect 21289 5978 21359 6023
rect 21417 5978 21487 6023
rect 21545 5978 21615 6023
rect 21673 5978 21743 6023
rect 21801 5978 21871 6023
rect 21929 5978 21999 6023
rect 22057 5978 22127 6023
rect 22185 5978 22255 6023
rect 22313 5978 22383 6023
rect 22441 5978 22511 6023
rect 22569 5978 22639 6023
rect 22697 5978 22767 6023
rect 22825 5978 22895 6023
rect 22953 5978 23023 6023
rect 23081 5978 23151 6023
rect 23209 5978 23279 6023
rect 23337 5978 23407 6023
rect 23465 5978 23535 6023
rect 23593 5978 23663 6023
rect 23721 5978 23791 6023
rect 23849 5978 23919 6023
rect 23977 5978 24047 6023
rect 24105 5978 24175 6023
rect 24233 5978 24303 6023
rect 24361 5978 24431 6023
rect 24489 5978 24559 6023
rect 24617 5978 24687 6023
rect 24745 5978 24815 6023
rect 24873 5978 24943 6023
rect 25001 5978 25071 6023
rect 25129 5978 25199 6023
rect 25257 5978 25327 6023
rect 25385 5978 25455 6023
rect 25513 5978 25583 6023
rect 25641 5978 25711 6023
rect 25769 5978 25839 6023
rect 25897 5978 25967 6023
rect 26025 5978 26095 6023
rect 26153 5978 26223 6023
rect 26281 5978 26351 6023
rect 26409 5978 26479 6023
rect 26537 5978 26607 6023
rect 26665 5978 26735 6023
rect 26793 5978 26863 6023
rect 26921 5978 26991 6023
rect 27049 5978 27119 6023
rect 27177 5978 27247 6023
rect 27305 5978 27375 6023
rect 27433 5978 27503 6023
rect 27561 5978 27631 6023
rect 27689 5978 27759 6023
rect 27817 5978 27887 6023
rect 27945 5978 28015 6023
rect 28073 5978 28143 6023
rect 28201 5978 28271 6023
rect 28329 5978 28399 6023
rect 28457 5978 28527 6023
rect -249 5868 -179 5894
rect 528 5868 598 5894
rect 656 5868 726 5894
rect 1437 5868 1507 5894
rect 1565 5868 1635 5894
rect 1693 5868 1763 5894
rect 1821 5868 1891 5894
rect 2970 5868 3040 5894
rect 3098 5868 3168 5894
rect 3226 5868 3296 5894
rect 3354 5868 3424 5894
rect 3482 5868 3552 5894
rect 3610 5868 3680 5894
rect 3738 5868 3808 5894
rect 3866 5868 3936 5894
rect 5521 5868 5591 5894
rect 5649 5868 5719 5894
rect 5777 5868 5847 5894
rect 5905 5868 5975 5894
rect 6033 5868 6103 5894
rect 6161 5868 6231 5894
rect 6289 5868 6359 5894
rect 6417 5868 6487 5894
rect 6545 5868 6615 5894
rect 6673 5868 6743 5894
rect 6801 5868 6871 5894
rect 6929 5868 6999 5894
rect 7057 5868 7127 5894
rect 7185 5868 7255 5894
rect 7313 5868 7383 5894
rect 7441 5868 7511 5894
rect 10608 5868 10678 5894
rect 10736 5868 10806 5894
rect 10864 5868 10934 5894
rect 10992 5868 11062 5894
rect 11120 5868 11190 5894
rect 11248 5868 11318 5894
rect 11376 5868 11446 5894
rect 11504 5868 11574 5894
rect 11632 5868 11702 5894
rect 11760 5868 11830 5894
rect 11888 5868 11958 5894
rect 12016 5868 12086 5894
rect 12144 5868 12214 5894
rect 12272 5868 12342 5894
rect 12400 5868 12470 5894
rect 12528 5868 12598 5894
rect 12656 5868 12726 5894
rect 12784 5868 12854 5894
rect 12912 5868 12982 5894
rect 13040 5868 13110 5894
rect 13168 5868 13238 5894
rect 13296 5868 13366 5894
rect 13424 5868 13494 5894
rect 13552 5868 13622 5894
rect 13680 5868 13750 5894
rect 13808 5868 13878 5894
rect 13936 5868 14006 5894
rect 14064 5868 14134 5894
rect 14192 5868 14262 5894
rect 14320 5868 14390 5894
rect 14448 5868 14518 5894
rect 14576 5868 14646 5894
rect 20393 5868 20463 5894
rect 20521 5868 20591 5894
rect 20649 5868 20719 5894
rect 20777 5868 20847 5894
rect 20905 5868 20975 5894
rect 21033 5868 21103 5894
rect 21161 5868 21231 5894
rect 21289 5868 21359 5894
rect 21417 5868 21487 5894
rect 21545 5868 21615 5894
rect 21673 5868 21743 5894
rect 21801 5868 21871 5894
rect 21929 5868 21999 5894
rect 22057 5868 22127 5894
rect 22185 5868 22255 5894
rect 22313 5868 22383 5894
rect 22441 5868 22511 5894
rect 22569 5868 22639 5894
rect 22697 5868 22767 5894
rect 22825 5868 22895 5894
rect 22953 5868 23023 5894
rect 23081 5868 23151 5894
rect 23209 5868 23279 5894
rect 23337 5868 23407 5894
rect 23465 5868 23535 5894
rect 23593 5868 23663 5894
rect 23721 5868 23791 5894
rect 23849 5868 23919 5894
rect 23977 5868 24047 5894
rect 24105 5868 24175 5894
rect 24233 5868 24303 5894
rect 24361 5868 24431 5894
rect 24489 5868 24559 5894
rect 24617 5868 24687 5894
rect 24745 5868 24815 5894
rect 24873 5868 24943 5894
rect 25001 5868 25071 5894
rect 25129 5868 25199 5894
rect 25257 5868 25327 5894
rect 25385 5868 25455 5894
rect 25513 5868 25583 5894
rect 25641 5868 25711 5894
rect 25769 5868 25839 5894
rect 25897 5868 25967 5894
rect 26025 5868 26095 5894
rect 26153 5868 26223 5894
rect 26281 5868 26351 5894
rect 26409 5868 26479 5894
rect 26537 5868 26607 5894
rect 26665 5868 26735 5894
rect 26793 5868 26863 5894
rect 26921 5868 26991 5894
rect 27049 5868 27119 5894
rect 27177 5868 27247 5894
rect 27305 5868 27375 5894
rect 27433 5868 27503 5894
rect 27561 5868 27631 5894
rect 27689 5868 27759 5894
rect 27817 5868 27887 5894
rect 27945 5868 28015 5894
rect 28073 5868 28143 5894
rect 28201 5868 28271 5894
rect 28329 5868 28399 5894
rect 28457 5868 28527 5894
rect -271 5590 -201 5621
rect 657 5590 727 5621
rect 785 5590 855 5621
rect 1921 5590 1991 5621
rect 2049 5590 2119 5621
rect 2177 5590 2247 5621
rect 2305 5590 2375 5621
rect 3540 5590 3610 5621
rect 3668 5590 3738 5621
rect 3796 5590 3866 5621
rect 3924 5590 3994 5621
rect 4052 5590 4122 5621
rect 4180 5590 4250 5621
rect 4308 5590 4378 5621
rect 4436 5590 4506 5621
rect 8105 5590 8175 5621
rect 8233 5590 8303 5621
rect 8361 5590 8431 5621
rect 8489 5590 8559 5621
rect 8617 5590 8687 5621
rect 8745 5590 8815 5621
rect 8873 5590 8943 5621
rect 9001 5590 9071 5621
rect 9129 5590 9199 5621
rect 9257 5590 9327 5621
rect 9385 5590 9455 5621
rect 9513 5590 9583 5621
rect 9641 5590 9711 5621
rect 9769 5590 9839 5621
rect 9897 5590 9967 5621
rect 10025 5590 10095 5621
rect 15263 5590 15333 5621
rect 15391 5590 15461 5621
rect 15519 5590 15589 5621
rect 15647 5590 15717 5621
rect 15775 5590 15845 5621
rect 15903 5590 15973 5621
rect 16031 5590 16101 5621
rect 16159 5590 16229 5621
rect 16287 5590 16357 5621
rect 16415 5590 16485 5621
rect 16543 5590 16613 5621
rect 16671 5590 16741 5621
rect 16799 5590 16869 5621
rect 16927 5590 16997 5621
rect 17055 5590 17125 5621
rect 17183 5590 17253 5621
rect 17311 5590 17381 5621
rect 17439 5590 17509 5621
rect 17567 5590 17637 5621
rect 17695 5590 17765 5621
rect 17823 5590 17893 5621
rect 17951 5590 18021 5621
rect 18079 5590 18149 5621
rect 18207 5590 18277 5621
rect 18335 5590 18405 5621
rect 18463 5590 18533 5621
rect 18591 5590 18661 5621
rect 18719 5590 18789 5621
rect 18847 5590 18917 5621
rect 18975 5590 19045 5621
rect 19103 5590 19173 5621
rect 19231 5590 19301 5621
rect 20317 5590 20387 5621
rect 20445 5590 20515 5621
rect 20573 5590 20643 5621
rect 20701 5590 20771 5621
rect 20829 5590 20899 5621
rect 20957 5590 21027 5621
rect 21085 5590 21155 5621
rect 21213 5590 21283 5621
rect 21341 5590 21411 5621
rect 21469 5590 21539 5621
rect 21597 5590 21667 5621
rect 21725 5590 21795 5621
rect 21853 5590 21923 5621
rect 21981 5590 22051 5621
rect 22109 5590 22179 5621
rect 22237 5590 22307 5621
rect 22365 5590 22435 5621
rect 22493 5590 22563 5621
rect 22621 5590 22691 5621
rect 22749 5590 22819 5621
rect 22877 5590 22947 5621
rect 23005 5590 23075 5621
rect 23133 5590 23203 5621
rect 23261 5590 23331 5621
rect 23389 5590 23459 5621
rect 23517 5590 23587 5621
rect 23645 5590 23715 5621
rect 23773 5590 23843 5621
rect 23901 5590 23971 5621
rect 24029 5590 24099 5621
rect 24157 5590 24227 5621
rect 24285 5590 24355 5621
rect 24413 5590 24483 5621
rect 24541 5590 24611 5621
rect 24669 5590 24739 5621
rect 24797 5590 24867 5621
rect 24925 5590 24995 5621
rect 25053 5590 25123 5621
rect 25181 5590 25251 5621
rect 25309 5590 25379 5621
rect 25437 5590 25507 5621
rect 25565 5590 25635 5621
rect 25693 5590 25763 5621
rect 25821 5590 25891 5621
rect 25949 5590 26019 5621
rect 26077 5590 26147 5621
rect 26205 5590 26275 5621
rect 26333 5590 26403 5621
rect 26461 5590 26531 5621
rect 26589 5590 26659 5621
rect 26717 5590 26787 5621
rect 26845 5590 26915 5621
rect 26973 5590 27043 5621
rect 27101 5590 27171 5621
rect 27229 5590 27299 5621
rect 27357 5590 27427 5621
rect 27485 5590 27555 5621
rect 27613 5590 27683 5621
rect 27741 5590 27811 5621
rect 27869 5590 27939 5621
rect 27997 5590 28067 5621
rect 28125 5590 28195 5621
rect 28253 5590 28323 5621
rect 28381 5590 28451 5621
rect -271 5290 -201 5422
rect 657 5405 727 5422
rect 785 5405 855 5422
rect 657 5335 855 5405
rect 657 5290 727 5335
rect 785 5290 855 5335
rect 1921 5405 1991 5422
rect 2049 5405 2119 5422
rect 2177 5405 2247 5422
rect 2305 5405 2375 5422
rect 1921 5335 2375 5405
rect 1921 5290 1991 5335
rect 2049 5290 2119 5335
rect 2177 5290 2247 5335
rect 2305 5290 2375 5335
rect 3540 5405 3610 5422
rect 3668 5405 3738 5422
rect 3796 5405 3866 5422
rect 3924 5405 3994 5422
rect 4052 5405 4122 5422
rect 4180 5405 4250 5422
rect 4308 5405 4378 5422
rect 4436 5405 4506 5422
rect 3540 5335 4506 5405
rect 3540 5290 3610 5335
rect 3668 5290 3738 5335
rect 3796 5290 3866 5335
rect 3924 5290 3994 5335
rect 4052 5290 4122 5335
rect 4180 5290 4250 5335
rect 4308 5290 4378 5335
rect 4436 5290 4506 5335
rect 8105 5405 8175 5422
rect 8233 5405 8303 5422
rect 8361 5405 8431 5422
rect 8489 5405 8559 5422
rect 8617 5405 8687 5422
rect 8745 5405 8815 5422
rect 8873 5405 8943 5422
rect 9001 5405 9071 5422
rect 9129 5405 9199 5422
rect 9257 5405 9327 5422
rect 9385 5405 9455 5422
rect 9513 5405 9583 5422
rect 9641 5405 9711 5422
rect 9769 5405 9839 5422
rect 9897 5405 9967 5422
rect 10025 5405 10095 5422
rect 8105 5335 10095 5405
rect 8105 5290 8175 5335
rect 8233 5290 8303 5335
rect 8361 5290 8431 5335
rect 8489 5290 8559 5335
rect 8617 5290 8687 5335
rect 8745 5290 8815 5335
rect 8873 5290 8943 5335
rect 9001 5290 9071 5335
rect 9129 5290 9199 5335
rect 9257 5290 9327 5335
rect 9385 5290 9455 5335
rect 9513 5290 9583 5335
rect 9641 5290 9711 5335
rect 9769 5290 9839 5335
rect 9897 5290 9967 5335
rect 10025 5290 10095 5335
rect 15263 5405 15333 5422
rect 15391 5405 15461 5422
rect 15519 5405 15589 5422
rect 15647 5405 15717 5422
rect 15775 5405 15845 5422
rect 15903 5405 15973 5422
rect 16031 5405 16101 5422
rect 16159 5405 16229 5422
rect 16287 5405 16357 5422
rect 16415 5405 16485 5422
rect 16543 5405 16613 5422
rect 16671 5405 16741 5422
rect 16799 5405 16869 5422
rect 16927 5405 16997 5422
rect 17055 5405 17125 5422
rect 17183 5405 17253 5422
rect 17311 5405 17381 5422
rect 17439 5405 17509 5422
rect 17567 5405 17637 5422
rect 17695 5405 17765 5422
rect 17823 5405 17893 5422
rect 17951 5405 18021 5422
rect 18079 5405 18149 5422
rect 18207 5405 18277 5422
rect 18335 5405 18405 5422
rect 18463 5405 18533 5422
rect 18591 5405 18661 5422
rect 18719 5405 18789 5422
rect 18847 5405 18917 5422
rect 18975 5405 19045 5422
rect 19103 5405 19173 5422
rect 19231 5405 19301 5422
rect 15263 5335 19301 5405
rect 15263 5290 15333 5335
rect 15391 5290 15461 5335
rect 15519 5290 15589 5335
rect 15647 5290 15717 5335
rect 15775 5290 15845 5335
rect 15903 5290 15973 5335
rect 16031 5290 16101 5335
rect 16159 5290 16229 5335
rect 16287 5290 16357 5335
rect 16415 5290 16485 5335
rect 16543 5290 16613 5335
rect 16671 5290 16741 5335
rect 16799 5290 16869 5335
rect 16927 5290 16997 5335
rect 17055 5290 17125 5335
rect 17183 5290 17253 5335
rect 17311 5290 17381 5335
rect 17439 5290 17509 5335
rect 17567 5290 17637 5335
rect 17695 5290 17765 5335
rect 17823 5290 17893 5335
rect 17951 5290 18021 5335
rect 18079 5290 18149 5335
rect 18207 5290 18277 5335
rect 18335 5290 18405 5335
rect 18463 5290 18533 5335
rect 18591 5290 18661 5335
rect 18719 5290 18789 5335
rect 18847 5290 18917 5335
rect 18975 5290 19045 5335
rect 19103 5290 19173 5335
rect 19231 5290 19301 5335
rect 20317 5405 20387 5422
rect 20445 5405 20515 5422
rect 20573 5405 20643 5422
rect 20701 5405 20771 5422
rect 20829 5405 20899 5422
rect 20957 5405 21027 5422
rect 21085 5405 21155 5422
rect 21213 5405 21283 5422
rect 21341 5405 21411 5422
rect 21469 5405 21539 5422
rect 21597 5405 21667 5422
rect 21725 5405 21795 5422
rect 21853 5405 21923 5422
rect 21981 5405 22051 5422
rect 22109 5405 22179 5422
rect 22237 5405 22307 5422
rect 22365 5405 22435 5422
rect 22493 5405 22563 5422
rect 22621 5405 22691 5422
rect 22749 5405 22819 5422
rect 22877 5405 22947 5422
rect 23005 5405 23075 5422
rect 23133 5405 23203 5422
rect 23261 5405 23331 5422
rect 23389 5405 23459 5422
rect 23517 5405 23587 5422
rect 23645 5405 23715 5422
rect 23773 5405 23843 5422
rect 23901 5405 23971 5422
rect 24029 5405 24099 5422
rect 24157 5405 24227 5422
rect 24285 5405 24355 5422
rect 24413 5405 24483 5422
rect 24541 5405 24611 5422
rect 24669 5405 24739 5422
rect 24797 5405 24867 5422
rect 24925 5405 24995 5422
rect 25053 5405 25123 5422
rect 25181 5405 25251 5422
rect 25309 5405 25379 5422
rect 25437 5405 25507 5422
rect 25565 5405 25635 5422
rect 25693 5405 25763 5422
rect 25821 5405 25891 5422
rect 25949 5405 26019 5422
rect 26077 5405 26147 5422
rect 26205 5405 26275 5422
rect 26333 5405 26403 5422
rect 26461 5405 26531 5422
rect 26589 5405 26659 5422
rect 26717 5405 26787 5422
rect 26845 5405 26915 5422
rect 26973 5405 27043 5422
rect 27101 5405 27171 5422
rect 27229 5405 27299 5422
rect 27357 5405 27427 5422
rect 27485 5405 27555 5422
rect 27613 5405 27683 5422
rect 27741 5405 27811 5422
rect 27869 5405 27939 5422
rect 27997 5405 28067 5422
rect 28125 5405 28195 5422
rect 28253 5405 28323 5422
rect 28381 5405 28451 5422
rect 20317 5335 28451 5405
rect 20317 5290 20387 5335
rect 20445 5290 20515 5335
rect 20573 5290 20643 5335
rect 20701 5290 20771 5335
rect 20829 5290 20899 5335
rect 20957 5290 21027 5335
rect 21085 5290 21155 5335
rect 21213 5290 21283 5335
rect 21341 5290 21411 5335
rect 21469 5290 21539 5335
rect 21597 5290 21667 5335
rect 21725 5290 21795 5335
rect 21853 5290 21923 5335
rect 21981 5290 22051 5335
rect 22109 5290 22179 5335
rect 22237 5290 22307 5335
rect 22365 5290 22435 5335
rect 22493 5290 22563 5335
rect 22621 5290 22691 5335
rect 22749 5290 22819 5335
rect 22877 5290 22947 5335
rect 23005 5290 23075 5335
rect 23133 5290 23203 5335
rect 23261 5290 23331 5335
rect 23389 5290 23459 5335
rect 23517 5290 23587 5335
rect 23645 5290 23715 5335
rect 23773 5290 23843 5335
rect 23901 5290 23971 5335
rect 24029 5290 24099 5335
rect 24157 5290 24227 5335
rect 24285 5290 24355 5335
rect 24413 5290 24483 5335
rect 24541 5290 24611 5335
rect 24669 5290 24739 5335
rect 24797 5290 24867 5335
rect 24925 5290 24995 5335
rect 25053 5290 25123 5335
rect 25181 5290 25251 5335
rect 25309 5290 25379 5335
rect 25437 5290 25507 5335
rect 25565 5290 25635 5335
rect 25693 5290 25763 5335
rect 25821 5290 25891 5335
rect 25949 5290 26019 5335
rect 26077 5290 26147 5335
rect 26205 5290 26275 5335
rect 26333 5290 26403 5335
rect 26461 5290 26531 5335
rect 26589 5290 26659 5335
rect 26717 5290 26787 5335
rect 26845 5290 26915 5335
rect 26973 5290 27043 5335
rect 27101 5290 27171 5335
rect 27229 5290 27299 5335
rect 27357 5290 27427 5335
rect 27485 5290 27555 5335
rect 27613 5290 27683 5335
rect 27741 5290 27811 5335
rect 27869 5290 27939 5335
rect 27997 5290 28067 5335
rect 28125 5290 28195 5335
rect 28253 5290 28323 5335
rect 28381 5290 28451 5335
rect -271 5180 -201 5206
rect 657 5180 727 5206
rect 785 5180 855 5206
rect 1921 5180 1991 5206
rect 2049 5180 2119 5206
rect 2177 5180 2247 5206
rect 2305 5180 2375 5206
rect 3540 5180 3610 5206
rect 3668 5180 3738 5206
rect 3796 5180 3866 5206
rect 3924 5180 3994 5206
rect 4052 5180 4122 5206
rect 4180 5180 4250 5206
rect 4308 5180 4378 5206
rect 4436 5180 4506 5206
rect 8105 5180 8175 5206
rect 8233 5180 8303 5206
rect 8361 5180 8431 5206
rect 8489 5180 8559 5206
rect 8617 5180 8687 5206
rect 8745 5180 8815 5206
rect 8873 5180 8943 5206
rect 9001 5180 9071 5206
rect 9129 5180 9199 5206
rect 9257 5180 9327 5206
rect 9385 5180 9455 5206
rect 9513 5180 9583 5206
rect 9641 5180 9711 5206
rect 9769 5180 9839 5206
rect 9897 5180 9967 5206
rect 10025 5180 10095 5206
rect 15263 5180 15333 5206
rect 15391 5180 15461 5206
rect 15519 5180 15589 5206
rect 15647 5180 15717 5206
rect 15775 5180 15845 5206
rect 15903 5180 15973 5206
rect 16031 5180 16101 5206
rect 16159 5180 16229 5206
rect 16287 5180 16357 5206
rect 16415 5180 16485 5206
rect 16543 5180 16613 5206
rect 16671 5180 16741 5206
rect 16799 5180 16869 5206
rect 16927 5180 16997 5206
rect 17055 5180 17125 5206
rect 17183 5180 17253 5206
rect 17311 5180 17381 5206
rect 17439 5180 17509 5206
rect 17567 5180 17637 5206
rect 17695 5180 17765 5206
rect 17823 5180 17893 5206
rect 17951 5180 18021 5206
rect 18079 5180 18149 5206
rect 18207 5180 18277 5206
rect 18335 5180 18405 5206
rect 18463 5180 18533 5206
rect 18591 5180 18661 5206
rect 18719 5180 18789 5206
rect 18847 5180 18917 5206
rect 18975 5180 19045 5206
rect 19103 5180 19173 5206
rect 19231 5180 19301 5206
rect 20317 5180 20387 5206
rect 20445 5180 20515 5206
rect 20573 5180 20643 5206
rect 20701 5180 20771 5206
rect 20829 5180 20899 5206
rect 20957 5180 21027 5206
rect 21085 5180 21155 5206
rect 21213 5180 21283 5206
rect 21341 5180 21411 5206
rect 21469 5180 21539 5206
rect 21597 5180 21667 5206
rect 21725 5180 21795 5206
rect 21853 5180 21923 5206
rect 21981 5180 22051 5206
rect 22109 5180 22179 5206
rect 22237 5180 22307 5206
rect 22365 5180 22435 5206
rect 22493 5180 22563 5206
rect 22621 5180 22691 5206
rect 22749 5180 22819 5206
rect 22877 5180 22947 5206
rect 23005 5180 23075 5206
rect 23133 5180 23203 5206
rect 23261 5180 23331 5206
rect 23389 5180 23459 5206
rect 23517 5180 23587 5206
rect 23645 5180 23715 5206
rect 23773 5180 23843 5206
rect 23901 5180 23971 5206
rect 24029 5180 24099 5206
rect 24157 5180 24227 5206
rect 24285 5180 24355 5206
rect 24413 5180 24483 5206
rect 24541 5180 24611 5206
rect 24669 5180 24739 5206
rect 24797 5180 24867 5206
rect 24925 5180 24995 5206
rect 25053 5180 25123 5206
rect 25181 5180 25251 5206
rect 25309 5180 25379 5206
rect 25437 5180 25507 5206
rect 25565 5180 25635 5206
rect 25693 5180 25763 5206
rect 25821 5180 25891 5206
rect 25949 5180 26019 5206
rect 26077 5180 26147 5206
rect 26205 5180 26275 5206
rect 26333 5180 26403 5206
rect 26461 5180 26531 5206
rect 26589 5180 26659 5206
rect 26717 5180 26787 5206
rect 26845 5180 26915 5206
rect 26973 5180 27043 5206
rect 27101 5180 27171 5206
rect 27229 5180 27299 5206
rect 27357 5180 27427 5206
rect 27485 5180 27555 5206
rect 27613 5180 27683 5206
rect 27741 5180 27811 5206
rect 27869 5180 27939 5206
rect 27997 5180 28067 5206
rect 28125 5180 28195 5206
rect 28253 5180 28323 5206
rect 28381 5180 28451 5206
<< locali >>
rect -341 6416 28619 6420
rect -341 6378 -297 6416
rect -259 6378 -169 6416
rect -131 6378 480 6416
rect 518 6378 608 6416
rect 646 6378 736 6416
rect 774 6378 1389 6416
rect 1427 6378 1517 6416
rect 1555 6378 1645 6416
rect 1683 6378 1773 6416
rect 1811 6378 1901 6416
rect 1939 6378 2922 6416
rect 2960 6378 3050 6416
rect 3088 6378 3178 6416
rect 3216 6378 3306 6416
rect 3344 6378 3434 6416
rect 3472 6378 3562 6416
rect 3600 6378 3690 6416
rect 3728 6378 3818 6416
rect 3856 6378 3946 6416
rect 3984 6378 5473 6416
rect 5511 6378 5601 6416
rect 5639 6378 5729 6416
rect 5767 6378 5857 6416
rect 5895 6378 5985 6416
rect 6023 6378 6113 6416
rect 6151 6378 6241 6416
rect 6279 6378 6369 6416
rect 6407 6378 6497 6416
rect 6535 6378 6625 6416
rect 6663 6378 6753 6416
rect 6791 6378 6881 6416
rect 6919 6378 7009 6416
rect 7047 6378 7137 6416
rect 7175 6378 7265 6416
rect 7303 6378 7393 6416
rect 7431 6378 7521 6416
rect 7559 6378 10560 6416
rect 10598 6378 10688 6416
rect 10726 6378 10816 6416
rect 10854 6378 10944 6416
rect 10982 6378 11072 6416
rect 11110 6378 11200 6416
rect 11238 6378 11328 6416
rect 11366 6378 11456 6416
rect 11494 6378 11584 6416
rect 11622 6378 11712 6416
rect 11750 6378 11840 6416
rect 11878 6378 11968 6416
rect 12006 6378 12096 6416
rect 12134 6378 12224 6416
rect 12262 6378 12352 6416
rect 12390 6378 12480 6416
rect 12518 6378 12608 6416
rect 12646 6378 12736 6416
rect 12774 6378 12864 6416
rect 12902 6378 12992 6416
rect 13030 6378 13120 6416
rect 13158 6378 13248 6416
rect 13286 6378 13376 6416
rect 13414 6378 13504 6416
rect 13542 6378 13632 6416
rect 13670 6378 13760 6416
rect 13798 6378 13888 6416
rect 13926 6378 14016 6416
rect 14054 6378 14144 6416
rect 14182 6378 14272 6416
rect 14310 6378 14400 6416
rect 14438 6378 14528 6416
rect 14566 6378 14656 6416
rect 14694 6378 20345 6416
rect 20383 6378 20473 6416
rect 20511 6378 20601 6416
rect 20639 6378 20729 6416
rect 20767 6378 20857 6416
rect 20895 6378 20985 6416
rect 21023 6378 21113 6416
rect 21151 6378 21241 6416
rect 21279 6378 21369 6416
rect 21407 6378 21497 6416
rect 21535 6378 21625 6416
rect 21663 6378 21753 6416
rect 21791 6378 21881 6416
rect 21919 6378 22009 6416
rect 22047 6378 22137 6416
rect 22175 6378 22265 6416
rect 22303 6378 22393 6416
rect 22431 6378 22521 6416
rect 22559 6378 22649 6416
rect 22687 6378 22777 6416
rect 22815 6378 22905 6416
rect 22943 6378 23033 6416
rect 23071 6378 23161 6416
rect 23199 6378 23289 6416
rect 23327 6378 23417 6416
rect 23455 6378 23545 6416
rect 23583 6378 23673 6416
rect 23711 6378 23801 6416
rect 23839 6378 23929 6416
rect 23967 6378 24057 6416
rect 24095 6378 24185 6416
rect 24223 6378 24313 6416
rect 24351 6378 24441 6416
rect 24479 6378 24569 6416
rect 24607 6378 24697 6416
rect 24735 6378 24825 6416
rect 24863 6378 24953 6416
rect 24991 6378 25081 6416
rect 25119 6378 25209 6416
rect 25247 6378 25337 6416
rect 25375 6378 25465 6416
rect 25503 6378 25593 6416
rect 25631 6378 25721 6416
rect 25759 6378 25849 6416
rect 25887 6378 25977 6416
rect 26015 6378 26105 6416
rect 26143 6378 26233 6416
rect 26271 6378 26361 6416
rect 26399 6378 26489 6416
rect 26527 6378 26617 6416
rect 26655 6378 26745 6416
rect 26783 6378 26873 6416
rect 26911 6378 27001 6416
rect 27039 6378 27129 6416
rect 27167 6378 27257 6416
rect 27295 6378 27385 6416
rect 27423 6378 27513 6416
rect 27551 6378 27641 6416
rect 27679 6378 27769 6416
rect 27807 6378 27897 6416
rect 27935 6378 28025 6416
rect 28063 6378 28153 6416
rect 28191 6378 28281 6416
rect 28319 6378 28409 6416
rect 28447 6378 28537 6416
rect 28575 6378 28619 6416
rect -341 6374 28619 6378
rect -295 6266 -261 6282
rect -295 6106 -261 6122
rect -167 6266 -133 6282
rect -167 6106 -133 6122
rect 482 6266 516 6282
rect 482 6106 516 6122
rect 610 6266 644 6282
rect 610 6106 644 6122
rect 738 6266 772 6282
rect 738 6106 772 6122
rect 1391 6266 1425 6282
rect 1391 6106 1425 6122
rect 1519 6266 1553 6282
rect 1519 6106 1553 6122
rect 1647 6266 1681 6282
rect 1647 6106 1681 6122
rect 1775 6266 1809 6282
rect 1775 6106 1809 6122
rect 1903 6266 1937 6282
rect 1903 6106 1937 6122
rect 2924 6266 2958 6282
rect 2924 6106 2958 6122
rect 3052 6266 3086 6282
rect 3052 6106 3086 6122
rect 3180 6266 3214 6282
rect 3180 6106 3214 6122
rect 3308 6266 3342 6282
rect 3308 6106 3342 6122
rect 3436 6266 3470 6282
rect 3436 6106 3470 6122
rect 3564 6266 3598 6282
rect 3564 6106 3598 6122
rect 3692 6266 3726 6282
rect 3692 6106 3726 6122
rect 3820 6266 3854 6282
rect 3820 6106 3854 6122
rect 3948 6266 3982 6282
rect 3948 6106 3982 6122
rect 5475 6266 5509 6282
rect 5475 6106 5509 6122
rect 5603 6266 5637 6282
rect 5603 6106 5637 6122
rect 5731 6266 5765 6282
rect 5731 6106 5765 6122
rect 5859 6266 5893 6282
rect 5859 6106 5893 6122
rect 5987 6266 6021 6282
rect 5987 6106 6021 6122
rect 6115 6266 6149 6282
rect 6115 6106 6149 6122
rect 6243 6266 6277 6282
rect 6243 6106 6277 6122
rect 6371 6266 6405 6282
rect 6371 6106 6405 6122
rect 6499 6266 6533 6282
rect 6499 6106 6533 6122
rect 6627 6266 6661 6282
rect 6627 6106 6661 6122
rect 6755 6266 6789 6282
rect 6755 6106 6789 6122
rect 6883 6266 6917 6282
rect 6883 6106 6917 6122
rect 7011 6266 7045 6282
rect 7011 6106 7045 6122
rect 7139 6266 7173 6282
rect 7139 6106 7173 6122
rect 7267 6266 7301 6282
rect 7267 6106 7301 6122
rect 7395 6266 7429 6282
rect 7395 6106 7429 6122
rect 7523 6266 7557 6282
rect 7523 6106 7557 6122
rect 10562 6266 10596 6282
rect 10562 6106 10596 6122
rect 10690 6266 10724 6282
rect 10690 6106 10724 6122
rect 10818 6266 10852 6282
rect 10818 6106 10852 6122
rect 10946 6266 10980 6282
rect 10946 6106 10980 6122
rect 11074 6266 11108 6282
rect 11074 6106 11108 6122
rect 11202 6266 11236 6282
rect 11202 6106 11236 6122
rect 11330 6266 11364 6282
rect 11330 6106 11364 6122
rect 11458 6266 11492 6282
rect 11458 6106 11492 6122
rect 11586 6266 11620 6282
rect 11586 6106 11620 6122
rect 11714 6266 11748 6282
rect 11714 6106 11748 6122
rect 11842 6266 11876 6282
rect 11842 6106 11876 6122
rect 11970 6266 12004 6282
rect 11970 6106 12004 6122
rect 12098 6266 12132 6282
rect 12098 6106 12132 6122
rect 12226 6266 12260 6282
rect 12226 6106 12260 6122
rect 12354 6266 12388 6282
rect 12354 6106 12388 6122
rect 12482 6266 12516 6282
rect 12482 6106 12516 6122
rect 12610 6266 12644 6282
rect 12610 6106 12644 6122
rect 12738 6266 12772 6282
rect 12738 6106 12772 6122
rect 12866 6266 12900 6282
rect 12866 6106 12900 6122
rect 12994 6266 13028 6282
rect 12994 6106 13028 6122
rect 13122 6266 13156 6282
rect 13122 6106 13156 6122
rect 13250 6266 13284 6282
rect 13250 6106 13284 6122
rect 13378 6266 13412 6282
rect 13378 6106 13412 6122
rect 13506 6266 13540 6282
rect 13506 6106 13540 6122
rect 13634 6266 13668 6282
rect 13634 6106 13668 6122
rect 13762 6266 13796 6282
rect 13762 6106 13796 6122
rect 13890 6266 13924 6282
rect 13890 6106 13924 6122
rect 14018 6266 14052 6282
rect 14018 6106 14052 6122
rect 14146 6266 14180 6282
rect 14146 6106 14180 6122
rect 14274 6266 14308 6282
rect 14274 6106 14308 6122
rect 14402 6266 14436 6282
rect 14402 6106 14436 6122
rect 14530 6266 14564 6282
rect 14530 6106 14564 6122
rect 14658 6266 14692 6282
rect 14658 6106 14692 6122
rect 20347 6266 20381 6282
rect 20347 6106 20381 6122
rect 20475 6266 20509 6282
rect 20475 6106 20509 6122
rect 20603 6266 20637 6282
rect 20603 6106 20637 6122
rect 20731 6266 20765 6282
rect 20731 6106 20765 6122
rect 20859 6266 20893 6282
rect 20859 6106 20893 6122
rect 20987 6266 21021 6282
rect 20987 6106 21021 6122
rect 21115 6266 21149 6282
rect 21115 6106 21149 6122
rect 21243 6266 21277 6282
rect 21243 6106 21277 6122
rect 21371 6266 21405 6282
rect 21371 6106 21405 6122
rect 21499 6266 21533 6282
rect 21499 6106 21533 6122
rect 21627 6266 21661 6282
rect 21627 6106 21661 6122
rect 21755 6266 21789 6282
rect 21755 6106 21789 6122
rect 21883 6266 21917 6282
rect 21883 6106 21917 6122
rect 22011 6266 22045 6282
rect 22011 6106 22045 6122
rect 22139 6266 22173 6282
rect 22139 6106 22173 6122
rect 22267 6266 22301 6282
rect 22267 6106 22301 6122
rect 22395 6266 22429 6282
rect 22395 6106 22429 6122
rect 22523 6266 22557 6282
rect 22523 6106 22557 6122
rect 22651 6266 22685 6282
rect 22651 6106 22685 6122
rect 22779 6266 22813 6282
rect 22779 6106 22813 6122
rect 22907 6266 22941 6282
rect 22907 6106 22941 6122
rect 23035 6266 23069 6282
rect 23035 6106 23069 6122
rect 23163 6266 23197 6282
rect 23163 6106 23197 6122
rect 23291 6266 23325 6282
rect 23291 6106 23325 6122
rect 23419 6266 23453 6282
rect 23419 6106 23453 6122
rect 23547 6266 23581 6282
rect 23547 6106 23581 6122
rect 23675 6266 23709 6282
rect 23675 6106 23709 6122
rect 23803 6266 23837 6282
rect 23803 6106 23837 6122
rect 23931 6266 23965 6282
rect 23931 6106 23965 6122
rect 24059 6266 24093 6282
rect 24059 6106 24093 6122
rect 24187 6266 24221 6282
rect 24187 6106 24221 6122
rect 24315 6266 24349 6282
rect 24315 6106 24349 6122
rect 24443 6266 24477 6282
rect 24443 6106 24477 6122
rect 24571 6266 24605 6282
rect 24571 6106 24605 6122
rect 24699 6266 24733 6282
rect 24699 6106 24733 6122
rect 24827 6266 24861 6282
rect 24827 6106 24861 6122
rect 24955 6266 24989 6282
rect 24955 6106 24989 6122
rect 25083 6266 25117 6282
rect 25083 6106 25117 6122
rect 25211 6266 25245 6282
rect 25211 6106 25245 6122
rect 25339 6266 25373 6282
rect 25339 6106 25373 6122
rect 25467 6266 25501 6282
rect 25467 6106 25501 6122
rect 25595 6266 25629 6282
rect 25595 6106 25629 6122
rect 25723 6266 25757 6282
rect 25723 6106 25757 6122
rect 25851 6266 25885 6282
rect 25851 6106 25885 6122
rect 25979 6266 26013 6282
rect 25979 6106 26013 6122
rect 26107 6266 26141 6282
rect 26107 6106 26141 6122
rect 26235 6266 26269 6282
rect 26235 6106 26269 6122
rect 26363 6266 26397 6282
rect 26363 6106 26397 6122
rect 26491 6266 26525 6282
rect 26491 6106 26525 6122
rect 26619 6266 26653 6282
rect 26619 6106 26653 6122
rect 26747 6266 26781 6282
rect 26747 6106 26781 6122
rect 26875 6266 26909 6282
rect 26875 6106 26909 6122
rect 27003 6266 27037 6282
rect 27003 6106 27037 6122
rect 27131 6266 27165 6282
rect 27131 6106 27165 6122
rect 27259 6266 27293 6282
rect 27259 6106 27293 6122
rect 27387 6266 27421 6282
rect 27387 6106 27421 6122
rect 27515 6266 27549 6282
rect 27515 6106 27549 6122
rect 27643 6266 27677 6282
rect 27643 6106 27677 6122
rect 27771 6266 27805 6282
rect 27771 6106 27805 6122
rect 27899 6266 27933 6282
rect 27899 6106 27933 6122
rect 28027 6266 28061 6282
rect 28027 6106 28061 6122
rect 28155 6266 28189 6282
rect 28155 6106 28189 6122
rect 28283 6266 28317 6282
rect 28283 6106 28317 6122
rect 28411 6266 28445 6282
rect 28411 6106 28445 6122
rect 28539 6266 28573 6282
rect 28539 6106 28573 6122
rect -295 5966 -261 5982
rect -295 5890 -261 5906
rect -167 5966 -133 5982
rect -167 5890 -133 5906
rect 482 5966 516 5982
rect 482 5890 516 5906
rect 610 5966 644 5982
rect 610 5890 644 5906
rect 738 5966 772 5982
rect 738 5890 772 5906
rect 1391 5966 1425 5982
rect 1391 5890 1425 5906
rect 1519 5966 1553 5982
rect 1519 5890 1553 5906
rect 1647 5966 1681 5982
rect 1647 5890 1681 5906
rect 1775 5966 1809 5982
rect 1775 5890 1809 5906
rect 1903 5966 1937 5982
rect 1903 5890 1937 5906
rect 2924 5966 2958 5982
rect 2924 5890 2958 5906
rect 3052 5966 3086 5982
rect 3052 5890 3086 5906
rect 3180 5966 3214 5982
rect 3180 5890 3214 5906
rect 3308 5966 3342 5982
rect 3308 5890 3342 5906
rect 3436 5966 3470 5982
rect 3436 5890 3470 5906
rect 3564 5966 3598 5982
rect 3564 5890 3598 5906
rect 3692 5966 3726 5982
rect 3692 5890 3726 5906
rect 3820 5966 3854 5982
rect 3820 5890 3854 5906
rect 3948 5966 3982 5982
rect 3948 5890 3982 5906
rect 5475 5966 5509 5982
rect 5475 5890 5509 5906
rect 5603 5966 5637 5982
rect 5603 5890 5637 5906
rect 5731 5966 5765 5982
rect 5731 5890 5765 5906
rect 5859 5966 5893 5982
rect 5859 5890 5893 5906
rect 5987 5966 6021 5982
rect 5987 5890 6021 5906
rect 6115 5966 6149 5982
rect 6115 5890 6149 5906
rect 6243 5966 6277 5982
rect 6243 5890 6277 5906
rect 6371 5966 6405 5982
rect 6371 5890 6405 5906
rect 6499 5966 6533 5982
rect 6499 5890 6533 5906
rect 6627 5966 6661 5982
rect 6627 5890 6661 5906
rect 6755 5966 6789 5982
rect 6755 5890 6789 5906
rect 6883 5966 6917 5982
rect 6883 5890 6917 5906
rect 7011 5966 7045 5982
rect 7011 5890 7045 5906
rect 7139 5966 7173 5982
rect 7139 5890 7173 5906
rect 7267 5966 7301 5982
rect 7267 5890 7301 5906
rect 7395 5966 7429 5982
rect 7395 5890 7429 5906
rect 7523 5966 7557 5982
rect 7523 5890 7557 5906
rect 10562 5966 10596 5982
rect 10562 5890 10596 5906
rect 10690 5966 10724 5982
rect 10690 5890 10724 5906
rect 10818 5966 10852 5982
rect 10818 5890 10852 5906
rect 10946 5966 10980 5982
rect 10946 5890 10980 5906
rect 11074 5966 11108 5982
rect 11074 5890 11108 5906
rect 11202 5966 11236 5982
rect 11202 5890 11236 5906
rect 11330 5966 11364 5982
rect 11330 5890 11364 5906
rect 11458 5966 11492 5982
rect 11458 5890 11492 5906
rect 11586 5966 11620 5982
rect 11586 5890 11620 5906
rect 11714 5966 11748 5982
rect 11714 5890 11748 5906
rect 11842 5966 11876 5982
rect 11842 5890 11876 5906
rect 11970 5966 12004 5982
rect 11970 5890 12004 5906
rect 12098 5966 12132 5982
rect 12098 5890 12132 5906
rect 12226 5966 12260 5982
rect 12226 5890 12260 5906
rect 12354 5966 12388 5982
rect 12354 5890 12388 5906
rect 12482 5966 12516 5982
rect 12482 5890 12516 5906
rect 12610 5966 12644 5982
rect 12610 5890 12644 5906
rect 12738 5966 12772 5982
rect 12738 5890 12772 5906
rect 12866 5966 12900 5982
rect 12866 5890 12900 5906
rect 12994 5966 13028 5982
rect 12994 5890 13028 5906
rect 13122 5966 13156 5982
rect 13122 5890 13156 5906
rect 13250 5966 13284 5982
rect 13250 5890 13284 5906
rect 13378 5966 13412 5982
rect 13378 5890 13412 5906
rect 13506 5966 13540 5982
rect 13506 5890 13540 5906
rect 13634 5966 13668 5982
rect 13634 5890 13668 5906
rect 13762 5966 13796 5982
rect 13762 5890 13796 5906
rect 13890 5966 13924 5982
rect 13890 5890 13924 5906
rect 14018 5966 14052 5982
rect 14018 5890 14052 5906
rect 14146 5966 14180 5982
rect 14146 5890 14180 5906
rect 14274 5966 14308 5982
rect 14274 5890 14308 5906
rect 14402 5966 14436 5982
rect 14402 5890 14436 5906
rect 14530 5966 14564 5982
rect 14530 5890 14564 5906
rect 14658 5966 14692 5982
rect 14658 5890 14692 5906
rect 20347 5966 20381 5982
rect 20347 5890 20381 5906
rect 20475 5966 20509 5982
rect 20475 5890 20509 5906
rect 20603 5966 20637 5982
rect 20603 5890 20637 5906
rect 20731 5966 20765 5982
rect 20731 5890 20765 5906
rect 20859 5966 20893 5982
rect 20859 5890 20893 5906
rect 20987 5966 21021 5982
rect 20987 5890 21021 5906
rect 21115 5966 21149 5982
rect 21115 5890 21149 5906
rect 21243 5966 21277 5982
rect 21243 5890 21277 5906
rect 21371 5966 21405 5982
rect 21371 5890 21405 5906
rect 21499 5966 21533 5982
rect 21499 5890 21533 5906
rect 21627 5966 21661 5982
rect 21627 5890 21661 5906
rect 21755 5966 21789 5982
rect 21755 5890 21789 5906
rect 21883 5966 21917 5982
rect 21883 5890 21917 5906
rect 22011 5966 22045 5982
rect 22011 5890 22045 5906
rect 22139 5966 22173 5982
rect 22139 5890 22173 5906
rect 22267 5966 22301 5982
rect 22267 5890 22301 5906
rect 22395 5966 22429 5982
rect 22395 5890 22429 5906
rect 22523 5966 22557 5982
rect 22523 5890 22557 5906
rect 22651 5966 22685 5982
rect 22651 5890 22685 5906
rect 22779 5966 22813 5982
rect 22779 5890 22813 5906
rect 22907 5966 22941 5982
rect 22907 5890 22941 5906
rect 23035 5966 23069 5982
rect 23035 5890 23069 5906
rect 23163 5966 23197 5982
rect 23163 5890 23197 5906
rect 23291 5966 23325 5982
rect 23291 5890 23325 5906
rect 23419 5966 23453 5982
rect 23419 5890 23453 5906
rect 23547 5966 23581 5982
rect 23547 5890 23581 5906
rect 23675 5966 23709 5982
rect 23675 5890 23709 5906
rect 23803 5966 23837 5982
rect 23803 5890 23837 5906
rect 23931 5966 23965 5982
rect 23931 5890 23965 5906
rect 24059 5966 24093 5982
rect 24059 5890 24093 5906
rect 24187 5966 24221 5982
rect 24187 5890 24221 5906
rect 24315 5966 24349 5982
rect 24315 5890 24349 5906
rect 24443 5966 24477 5982
rect 24443 5890 24477 5906
rect 24571 5966 24605 5982
rect 24571 5890 24605 5906
rect 24699 5966 24733 5982
rect 24699 5890 24733 5906
rect 24827 5966 24861 5982
rect 24827 5890 24861 5906
rect 24955 5966 24989 5982
rect 24955 5890 24989 5906
rect 25083 5966 25117 5982
rect 25083 5890 25117 5906
rect 25211 5966 25245 5982
rect 25211 5890 25245 5906
rect 25339 5966 25373 5982
rect 25339 5890 25373 5906
rect 25467 5966 25501 5982
rect 25467 5890 25501 5906
rect 25595 5966 25629 5982
rect 25595 5890 25629 5906
rect 25723 5966 25757 5982
rect 25723 5890 25757 5906
rect 25851 5966 25885 5982
rect 25851 5890 25885 5906
rect 25979 5966 26013 5982
rect 25979 5890 26013 5906
rect 26107 5966 26141 5982
rect 26107 5890 26141 5906
rect 26235 5966 26269 5982
rect 26235 5890 26269 5906
rect 26363 5966 26397 5982
rect 26363 5890 26397 5906
rect 26491 5966 26525 5982
rect 26491 5890 26525 5906
rect 26619 5966 26653 5982
rect 26619 5890 26653 5906
rect 26747 5966 26781 5982
rect 26747 5890 26781 5906
rect 26875 5966 26909 5982
rect 26875 5890 26909 5906
rect 27003 5966 27037 5982
rect 27003 5890 27037 5906
rect 27131 5966 27165 5982
rect 27131 5890 27165 5906
rect 27259 5966 27293 5982
rect 27259 5890 27293 5906
rect 27387 5966 27421 5982
rect 27387 5890 27421 5906
rect 27515 5966 27549 5982
rect 27515 5890 27549 5906
rect 27643 5966 27677 5982
rect 27643 5890 27677 5906
rect 27771 5966 27805 5982
rect 27771 5890 27805 5906
rect 27899 5966 27933 5982
rect 27899 5890 27933 5906
rect 28027 5966 28061 5982
rect 28027 5890 28061 5906
rect 28155 5966 28189 5982
rect 28155 5890 28189 5906
rect 28283 5966 28317 5982
rect 28283 5890 28317 5906
rect 28411 5966 28445 5982
rect 28411 5890 28445 5906
rect 28539 5966 28573 5982
rect 28539 5890 28573 5906
rect -341 5836 28619 5840
rect -341 5798 -297 5836
rect -259 5798 -169 5836
rect -131 5798 480 5836
rect 518 5798 608 5836
rect 646 5798 736 5836
rect 774 5798 1389 5836
rect 1427 5798 1517 5836
rect 1555 5798 1645 5836
rect 1683 5798 1773 5836
rect 1811 5798 1901 5836
rect 1939 5798 2922 5836
rect 2960 5798 3050 5836
rect 3088 5798 3178 5836
rect 3216 5798 3306 5836
rect 3344 5798 3434 5836
rect 3472 5798 3562 5836
rect 3600 5798 3690 5836
rect 3728 5798 3818 5836
rect 3856 5798 3946 5836
rect 3984 5798 5473 5836
rect 5511 5798 5601 5836
rect 5639 5798 5729 5836
rect 5767 5798 5857 5836
rect 5895 5798 5985 5836
rect 6023 5798 6113 5836
rect 6151 5798 6241 5836
rect 6279 5798 6369 5836
rect 6407 5798 6497 5836
rect 6535 5798 6625 5836
rect 6663 5798 6753 5836
rect 6791 5798 6881 5836
rect 6919 5798 7009 5836
rect 7047 5798 7137 5836
rect 7175 5798 7265 5836
rect 7303 5798 7393 5836
rect 7431 5798 7521 5836
rect 7559 5798 10560 5836
rect 10598 5798 10688 5836
rect 10726 5798 10816 5836
rect 10854 5798 10944 5836
rect 10982 5798 11072 5836
rect 11110 5798 11200 5836
rect 11238 5798 11328 5836
rect 11366 5798 11456 5836
rect 11494 5798 11584 5836
rect 11622 5798 11712 5836
rect 11750 5798 11840 5836
rect 11878 5798 11968 5836
rect 12006 5798 12096 5836
rect 12134 5798 12224 5836
rect 12262 5798 12352 5836
rect 12390 5798 12480 5836
rect 12518 5798 12608 5836
rect 12646 5798 12736 5836
rect 12774 5798 12864 5836
rect 12902 5798 12992 5836
rect 13030 5798 13120 5836
rect 13158 5798 13248 5836
rect 13286 5798 13376 5836
rect 13414 5798 13504 5836
rect 13542 5798 13632 5836
rect 13670 5798 13760 5836
rect 13798 5798 13888 5836
rect 13926 5798 14016 5836
rect 14054 5798 14144 5836
rect 14182 5798 14272 5836
rect 14310 5798 14400 5836
rect 14438 5798 14528 5836
rect 14566 5798 14656 5836
rect 14694 5798 20345 5836
rect 20383 5798 20473 5836
rect 20511 5798 20601 5836
rect 20639 5798 20729 5836
rect 20767 5798 20857 5836
rect 20895 5798 20985 5836
rect 21023 5798 21113 5836
rect 21151 5798 21241 5836
rect 21279 5798 21369 5836
rect 21407 5798 21497 5836
rect 21535 5798 21625 5836
rect 21663 5798 21753 5836
rect 21791 5798 21881 5836
rect 21919 5798 22009 5836
rect 22047 5798 22137 5836
rect 22175 5798 22265 5836
rect 22303 5798 22393 5836
rect 22431 5798 22521 5836
rect 22559 5798 22649 5836
rect 22687 5798 22777 5836
rect 22815 5798 22905 5836
rect 22943 5798 23033 5836
rect 23071 5798 23161 5836
rect 23199 5798 23289 5836
rect 23327 5798 23417 5836
rect 23455 5798 23545 5836
rect 23583 5798 23673 5836
rect 23711 5798 23801 5836
rect 23839 5798 23929 5836
rect 23967 5798 24057 5836
rect 24095 5798 24185 5836
rect 24223 5798 24313 5836
rect 24351 5798 24441 5836
rect 24479 5798 24569 5836
rect 24607 5798 24697 5836
rect 24735 5798 24825 5836
rect 24863 5798 24953 5836
rect 24991 5798 25081 5836
rect 25119 5798 25209 5836
rect 25247 5798 25337 5836
rect 25375 5798 25465 5836
rect 25503 5798 25593 5836
rect 25631 5798 25721 5836
rect 25759 5798 25849 5836
rect 25887 5798 25977 5836
rect 26015 5798 26105 5836
rect 26143 5798 26233 5836
rect 26271 5798 26361 5836
rect 26399 5798 26489 5836
rect 26527 5798 26617 5836
rect 26655 5798 26745 5836
rect 26783 5798 26873 5836
rect 26911 5798 27001 5836
rect 27039 5798 27129 5836
rect 27167 5798 27257 5836
rect 27295 5798 27385 5836
rect 27423 5798 27513 5836
rect 27551 5798 27641 5836
rect 27679 5798 27769 5836
rect 27807 5798 27897 5836
rect 27935 5798 28025 5836
rect 28063 5798 28153 5836
rect 28191 5798 28281 5836
rect 28319 5798 28409 5836
rect 28447 5798 28537 5836
rect 28575 5798 28619 5836
rect -341 5794 28619 5798
rect -363 5728 28543 5732
rect -363 5690 -319 5728
rect -281 5690 -191 5728
rect -153 5690 609 5728
rect 647 5690 737 5728
rect 775 5690 865 5728
rect 903 5690 1873 5728
rect 1911 5690 2001 5728
rect 2039 5690 2129 5728
rect 2167 5690 2257 5728
rect 2295 5690 2385 5728
rect 2423 5690 3492 5728
rect 3530 5690 3620 5728
rect 3658 5690 3748 5728
rect 3786 5690 3876 5728
rect 3914 5690 4004 5728
rect 4042 5690 4132 5728
rect 4170 5690 4260 5728
rect 4298 5690 4388 5728
rect 4426 5690 4516 5728
rect 4554 5690 8057 5728
rect 8095 5690 8185 5728
rect 8223 5690 8313 5728
rect 8351 5690 8441 5728
rect 8479 5690 8569 5728
rect 8607 5690 8697 5728
rect 8735 5690 8825 5728
rect 8863 5690 8953 5728
rect 8991 5690 9081 5728
rect 9119 5690 9209 5728
rect 9247 5690 9337 5728
rect 9375 5690 9465 5728
rect 9503 5690 9593 5728
rect 9631 5690 9721 5728
rect 9759 5690 9849 5728
rect 9887 5690 9977 5728
rect 10015 5690 10105 5728
rect 10143 5690 15215 5728
rect 15253 5690 15343 5728
rect 15381 5690 15471 5728
rect 15509 5690 15599 5728
rect 15637 5690 15727 5728
rect 15765 5690 15855 5728
rect 15893 5690 15983 5728
rect 16021 5690 16111 5728
rect 16149 5690 16239 5728
rect 16277 5690 16367 5728
rect 16405 5690 16495 5728
rect 16533 5690 16623 5728
rect 16661 5690 16751 5728
rect 16789 5690 16879 5728
rect 16917 5690 17007 5728
rect 17045 5690 17135 5728
rect 17173 5690 17263 5728
rect 17301 5690 17391 5728
rect 17429 5690 17519 5728
rect 17557 5690 17647 5728
rect 17685 5690 17775 5728
rect 17813 5690 17903 5728
rect 17941 5690 18031 5728
rect 18069 5690 18159 5728
rect 18197 5690 18287 5728
rect 18325 5690 18415 5728
rect 18453 5690 18543 5728
rect 18581 5690 18671 5728
rect 18709 5690 18799 5728
rect 18837 5690 18927 5728
rect 18965 5690 19055 5728
rect 19093 5690 19183 5728
rect 19221 5690 19311 5728
rect 19349 5690 20269 5728
rect 20307 5690 20397 5728
rect 20435 5690 20525 5728
rect 20563 5690 20653 5728
rect 20691 5690 20781 5728
rect 20819 5690 20909 5728
rect 20947 5690 21037 5728
rect 21075 5690 21165 5728
rect 21203 5690 21293 5728
rect 21331 5690 21421 5728
rect 21459 5690 21549 5728
rect 21587 5690 21677 5728
rect 21715 5690 21805 5728
rect 21843 5690 21933 5728
rect 21971 5690 22061 5728
rect 22099 5690 22189 5728
rect 22227 5690 22317 5728
rect 22355 5690 22445 5728
rect 22483 5690 22573 5728
rect 22611 5690 22701 5728
rect 22739 5690 22829 5728
rect 22867 5690 22957 5728
rect 22995 5690 23085 5728
rect 23123 5690 23213 5728
rect 23251 5690 23341 5728
rect 23379 5690 23469 5728
rect 23507 5690 23597 5728
rect 23635 5690 23725 5728
rect 23763 5690 23853 5728
rect 23891 5690 23981 5728
rect 24019 5690 24109 5728
rect 24147 5690 24237 5728
rect 24275 5690 24365 5728
rect 24403 5690 24493 5728
rect 24531 5690 24621 5728
rect 24659 5690 24749 5728
rect 24787 5690 24877 5728
rect 24915 5690 25005 5728
rect 25043 5690 25133 5728
rect 25171 5690 25261 5728
rect 25299 5690 25389 5728
rect 25427 5690 25517 5728
rect 25555 5690 25645 5728
rect 25683 5690 25773 5728
rect 25811 5690 25901 5728
rect 25939 5690 26029 5728
rect 26067 5690 26157 5728
rect 26195 5690 26285 5728
rect 26323 5690 26413 5728
rect 26451 5690 26541 5728
rect 26579 5690 26669 5728
rect 26707 5690 26797 5728
rect 26835 5690 26925 5728
rect 26963 5690 27053 5728
rect 27091 5690 27181 5728
rect 27219 5690 27309 5728
rect 27347 5690 27437 5728
rect 27475 5690 27565 5728
rect 27603 5690 27693 5728
rect 27731 5690 27821 5728
rect 27859 5690 27949 5728
rect 27987 5690 28077 5728
rect 28115 5690 28205 5728
rect 28243 5690 28333 5728
rect 28371 5690 28461 5728
rect 28499 5690 28543 5728
rect -363 5686 28543 5690
rect -317 5578 -283 5594
rect -317 5418 -283 5434
rect -189 5578 -155 5594
rect -189 5418 -155 5434
rect 611 5578 645 5594
rect 611 5418 645 5434
rect 739 5578 773 5594
rect 739 5418 773 5434
rect 867 5578 901 5594
rect 867 5418 901 5434
rect 1875 5578 1909 5594
rect 1875 5418 1909 5434
rect 2003 5578 2037 5594
rect 2003 5418 2037 5434
rect 2131 5578 2165 5594
rect 2131 5418 2165 5434
rect 2259 5578 2293 5594
rect 2259 5418 2293 5434
rect 2387 5578 2421 5594
rect 2387 5418 2421 5434
rect 3494 5578 3528 5594
rect 3494 5418 3528 5434
rect 3622 5578 3656 5594
rect 3622 5418 3656 5434
rect 3750 5578 3784 5594
rect 3750 5418 3784 5434
rect 3878 5578 3912 5594
rect 3878 5418 3912 5434
rect 4006 5578 4040 5594
rect 4006 5418 4040 5434
rect 4134 5578 4168 5594
rect 4134 5418 4168 5434
rect 4262 5578 4296 5594
rect 4262 5418 4296 5434
rect 4390 5578 4424 5594
rect 4390 5418 4424 5434
rect 4518 5578 4552 5594
rect 4518 5418 4552 5434
rect 8059 5578 8093 5594
rect 8059 5418 8093 5434
rect 8187 5578 8221 5594
rect 8187 5418 8221 5434
rect 8315 5578 8349 5594
rect 8315 5418 8349 5434
rect 8443 5578 8477 5594
rect 8443 5418 8477 5434
rect 8571 5578 8605 5594
rect 8571 5418 8605 5434
rect 8699 5578 8733 5594
rect 8699 5418 8733 5434
rect 8827 5578 8861 5594
rect 8827 5418 8861 5434
rect 8955 5578 8989 5594
rect 8955 5418 8989 5434
rect 9083 5578 9117 5594
rect 9083 5418 9117 5434
rect 9211 5578 9245 5594
rect 9211 5418 9245 5434
rect 9339 5578 9373 5594
rect 9339 5418 9373 5434
rect 9467 5578 9501 5594
rect 9467 5418 9501 5434
rect 9595 5578 9629 5594
rect 9595 5418 9629 5434
rect 9723 5578 9757 5594
rect 9723 5418 9757 5434
rect 9851 5578 9885 5594
rect 9851 5418 9885 5434
rect 9979 5578 10013 5594
rect 9979 5418 10013 5434
rect 10107 5578 10141 5594
rect 10107 5418 10141 5434
rect 15217 5578 15251 5594
rect 15217 5418 15251 5434
rect 15345 5578 15379 5594
rect 15345 5418 15379 5434
rect 15473 5578 15507 5594
rect 15473 5418 15507 5434
rect 15601 5578 15635 5594
rect 15601 5418 15635 5434
rect 15729 5578 15763 5594
rect 15729 5418 15763 5434
rect 15857 5578 15891 5594
rect 15857 5418 15891 5434
rect 15985 5578 16019 5594
rect 15985 5418 16019 5434
rect 16113 5578 16147 5594
rect 16113 5418 16147 5434
rect 16241 5578 16275 5594
rect 16241 5418 16275 5434
rect 16369 5578 16403 5594
rect 16369 5418 16403 5434
rect 16497 5578 16531 5594
rect 16497 5418 16531 5434
rect 16625 5578 16659 5594
rect 16625 5418 16659 5434
rect 16753 5578 16787 5594
rect 16753 5418 16787 5434
rect 16881 5578 16915 5594
rect 16881 5418 16915 5434
rect 17009 5578 17043 5594
rect 17009 5418 17043 5434
rect 17137 5578 17171 5594
rect 17137 5418 17171 5434
rect 17265 5578 17299 5594
rect 17265 5418 17299 5434
rect 17393 5578 17427 5594
rect 17393 5418 17427 5434
rect 17521 5578 17555 5594
rect 17521 5418 17555 5434
rect 17649 5578 17683 5594
rect 17649 5418 17683 5434
rect 17777 5578 17811 5594
rect 17777 5418 17811 5434
rect 17905 5578 17939 5594
rect 17905 5418 17939 5434
rect 18033 5578 18067 5594
rect 18033 5418 18067 5434
rect 18161 5578 18195 5594
rect 18161 5418 18195 5434
rect 18289 5578 18323 5594
rect 18289 5418 18323 5434
rect 18417 5578 18451 5594
rect 18417 5418 18451 5434
rect 18545 5578 18579 5594
rect 18545 5418 18579 5434
rect 18673 5578 18707 5594
rect 18673 5418 18707 5434
rect 18801 5578 18835 5594
rect 18801 5418 18835 5434
rect 18929 5578 18963 5594
rect 18929 5418 18963 5434
rect 19057 5578 19091 5594
rect 19057 5418 19091 5434
rect 19185 5578 19219 5594
rect 19185 5418 19219 5434
rect 19313 5578 19347 5594
rect 19313 5418 19347 5434
rect 20271 5578 20305 5594
rect 20271 5418 20305 5434
rect 20399 5578 20433 5594
rect 20399 5418 20433 5434
rect 20527 5578 20561 5594
rect 20527 5418 20561 5434
rect 20655 5578 20689 5594
rect 20655 5418 20689 5434
rect 20783 5578 20817 5594
rect 20783 5418 20817 5434
rect 20911 5578 20945 5594
rect 20911 5418 20945 5434
rect 21039 5578 21073 5594
rect 21039 5418 21073 5434
rect 21167 5578 21201 5594
rect 21167 5418 21201 5434
rect 21295 5578 21329 5594
rect 21295 5418 21329 5434
rect 21423 5578 21457 5594
rect 21423 5418 21457 5434
rect 21551 5578 21585 5594
rect 21551 5418 21585 5434
rect 21679 5578 21713 5594
rect 21679 5418 21713 5434
rect 21807 5578 21841 5594
rect 21807 5418 21841 5434
rect 21935 5578 21969 5594
rect 21935 5418 21969 5434
rect 22063 5578 22097 5594
rect 22063 5418 22097 5434
rect 22191 5578 22225 5594
rect 22191 5418 22225 5434
rect 22319 5578 22353 5594
rect 22319 5418 22353 5434
rect 22447 5578 22481 5594
rect 22447 5418 22481 5434
rect 22575 5578 22609 5594
rect 22575 5418 22609 5434
rect 22703 5578 22737 5594
rect 22703 5418 22737 5434
rect 22831 5578 22865 5594
rect 22831 5418 22865 5434
rect 22959 5578 22993 5594
rect 22959 5418 22993 5434
rect 23087 5578 23121 5594
rect 23087 5418 23121 5434
rect 23215 5578 23249 5594
rect 23215 5418 23249 5434
rect 23343 5578 23377 5594
rect 23343 5418 23377 5434
rect 23471 5578 23505 5594
rect 23471 5418 23505 5434
rect 23599 5578 23633 5594
rect 23599 5418 23633 5434
rect 23727 5578 23761 5594
rect 23727 5418 23761 5434
rect 23855 5578 23889 5594
rect 23855 5418 23889 5434
rect 23983 5578 24017 5594
rect 23983 5418 24017 5434
rect 24111 5578 24145 5594
rect 24111 5418 24145 5434
rect 24239 5578 24273 5594
rect 24239 5418 24273 5434
rect 24367 5578 24401 5594
rect 24367 5418 24401 5434
rect 24495 5578 24529 5594
rect 24495 5418 24529 5434
rect 24623 5578 24657 5594
rect 24623 5418 24657 5434
rect 24751 5578 24785 5594
rect 24751 5418 24785 5434
rect 24879 5578 24913 5594
rect 24879 5418 24913 5434
rect 25007 5578 25041 5594
rect 25007 5418 25041 5434
rect 25135 5578 25169 5594
rect 25135 5418 25169 5434
rect 25263 5578 25297 5594
rect 25263 5418 25297 5434
rect 25391 5578 25425 5594
rect 25391 5418 25425 5434
rect 25519 5578 25553 5594
rect 25519 5418 25553 5434
rect 25647 5578 25681 5594
rect 25647 5418 25681 5434
rect 25775 5578 25809 5594
rect 25775 5418 25809 5434
rect 25903 5578 25937 5594
rect 25903 5418 25937 5434
rect 26031 5578 26065 5594
rect 26031 5418 26065 5434
rect 26159 5578 26193 5594
rect 26159 5418 26193 5434
rect 26287 5578 26321 5594
rect 26287 5418 26321 5434
rect 26415 5578 26449 5594
rect 26415 5418 26449 5434
rect 26543 5578 26577 5594
rect 26543 5418 26577 5434
rect 26671 5578 26705 5594
rect 26671 5418 26705 5434
rect 26799 5578 26833 5594
rect 26799 5418 26833 5434
rect 26927 5578 26961 5594
rect 26927 5418 26961 5434
rect 27055 5578 27089 5594
rect 27055 5418 27089 5434
rect 27183 5578 27217 5594
rect 27183 5418 27217 5434
rect 27311 5578 27345 5594
rect 27311 5418 27345 5434
rect 27439 5578 27473 5594
rect 27439 5418 27473 5434
rect 27567 5578 27601 5594
rect 27567 5418 27601 5434
rect 27695 5578 27729 5594
rect 27695 5418 27729 5434
rect 27823 5578 27857 5594
rect 27823 5418 27857 5434
rect 27951 5578 27985 5594
rect 27951 5418 27985 5434
rect 28079 5578 28113 5594
rect 28079 5418 28113 5434
rect 28207 5578 28241 5594
rect 28207 5418 28241 5434
rect 28335 5578 28369 5594
rect 28335 5418 28369 5434
rect 28463 5578 28497 5594
rect 28463 5418 28497 5434
rect -317 5278 -283 5294
rect -317 5202 -283 5218
rect -189 5278 -155 5294
rect -189 5202 -155 5218
rect 611 5278 645 5294
rect 611 5202 645 5218
rect 739 5278 773 5294
rect 739 5202 773 5218
rect 867 5278 901 5294
rect 867 5202 901 5218
rect 1875 5278 1909 5294
rect 1875 5202 1909 5218
rect 2003 5278 2037 5294
rect 2003 5202 2037 5218
rect 2131 5278 2165 5294
rect 2131 5202 2165 5218
rect 2259 5278 2293 5294
rect 2259 5202 2293 5218
rect 2387 5278 2421 5294
rect 2387 5202 2421 5218
rect 3494 5278 3528 5294
rect 3494 5202 3528 5218
rect 3622 5278 3656 5294
rect 3622 5202 3656 5218
rect 3750 5278 3784 5294
rect 3750 5202 3784 5218
rect 3878 5278 3912 5294
rect 3878 5202 3912 5218
rect 4006 5278 4040 5294
rect 4006 5202 4040 5218
rect 4134 5278 4168 5294
rect 4134 5202 4168 5218
rect 4262 5278 4296 5294
rect 4262 5202 4296 5218
rect 4390 5278 4424 5294
rect 4390 5202 4424 5218
rect 4518 5278 4552 5294
rect 4518 5202 4552 5218
rect 8059 5278 8093 5294
rect 8059 5202 8093 5218
rect 8187 5278 8221 5294
rect 8187 5202 8221 5218
rect 8315 5278 8349 5294
rect 8315 5202 8349 5218
rect 8443 5278 8477 5294
rect 8443 5202 8477 5218
rect 8571 5278 8605 5294
rect 8571 5202 8605 5218
rect 8699 5278 8733 5294
rect 8699 5202 8733 5218
rect 8827 5278 8861 5294
rect 8827 5202 8861 5218
rect 8955 5278 8989 5294
rect 8955 5202 8989 5218
rect 9083 5278 9117 5294
rect 9083 5202 9117 5218
rect 9211 5278 9245 5294
rect 9211 5202 9245 5218
rect 9339 5278 9373 5294
rect 9339 5202 9373 5218
rect 9467 5278 9501 5294
rect 9467 5202 9501 5218
rect 9595 5278 9629 5294
rect 9595 5202 9629 5218
rect 9723 5278 9757 5294
rect 9723 5202 9757 5218
rect 9851 5278 9885 5294
rect 9851 5202 9885 5218
rect 9979 5278 10013 5294
rect 9979 5202 10013 5218
rect 10107 5278 10141 5294
rect 10107 5202 10141 5218
rect 15217 5278 15251 5294
rect 15217 5202 15251 5218
rect 15345 5278 15379 5294
rect 15345 5202 15379 5218
rect 15473 5278 15507 5294
rect 15473 5202 15507 5218
rect 15601 5278 15635 5294
rect 15601 5202 15635 5218
rect 15729 5278 15763 5294
rect 15729 5202 15763 5218
rect 15857 5278 15891 5294
rect 15857 5202 15891 5218
rect 15985 5278 16019 5294
rect 15985 5202 16019 5218
rect 16113 5278 16147 5294
rect 16113 5202 16147 5218
rect 16241 5278 16275 5294
rect 16241 5202 16275 5218
rect 16369 5278 16403 5294
rect 16369 5202 16403 5218
rect 16497 5278 16531 5294
rect 16497 5202 16531 5218
rect 16625 5278 16659 5294
rect 16625 5202 16659 5218
rect 16753 5278 16787 5294
rect 16753 5202 16787 5218
rect 16881 5278 16915 5294
rect 16881 5202 16915 5218
rect 17009 5278 17043 5294
rect 17009 5202 17043 5218
rect 17137 5278 17171 5294
rect 17137 5202 17171 5218
rect 17265 5278 17299 5294
rect 17265 5202 17299 5218
rect 17393 5278 17427 5294
rect 17393 5202 17427 5218
rect 17521 5278 17555 5294
rect 17521 5202 17555 5218
rect 17649 5278 17683 5294
rect 17649 5202 17683 5218
rect 17777 5278 17811 5294
rect 17777 5202 17811 5218
rect 17905 5278 17939 5294
rect 17905 5202 17939 5218
rect 18033 5278 18067 5294
rect 18033 5202 18067 5218
rect 18161 5278 18195 5294
rect 18161 5202 18195 5218
rect 18289 5278 18323 5294
rect 18289 5202 18323 5218
rect 18417 5278 18451 5294
rect 18417 5202 18451 5218
rect 18545 5278 18579 5294
rect 18545 5202 18579 5218
rect 18673 5278 18707 5294
rect 18673 5202 18707 5218
rect 18801 5278 18835 5294
rect 18801 5202 18835 5218
rect 18929 5278 18963 5294
rect 18929 5202 18963 5218
rect 19057 5278 19091 5294
rect 19057 5202 19091 5218
rect 19185 5278 19219 5294
rect 19185 5202 19219 5218
rect 19313 5278 19347 5294
rect 19313 5202 19347 5218
rect 20271 5278 20305 5294
rect 20271 5202 20305 5218
rect 20399 5278 20433 5294
rect 20399 5202 20433 5218
rect 20527 5278 20561 5294
rect 20527 5202 20561 5218
rect 20655 5278 20689 5294
rect 20655 5202 20689 5218
rect 20783 5278 20817 5294
rect 20783 5202 20817 5218
rect 20911 5278 20945 5294
rect 20911 5202 20945 5218
rect 21039 5278 21073 5294
rect 21039 5202 21073 5218
rect 21167 5278 21201 5294
rect 21167 5202 21201 5218
rect 21295 5278 21329 5294
rect 21295 5202 21329 5218
rect 21423 5278 21457 5294
rect 21423 5202 21457 5218
rect 21551 5278 21585 5294
rect 21551 5202 21585 5218
rect 21679 5278 21713 5294
rect 21679 5202 21713 5218
rect 21807 5278 21841 5294
rect 21807 5202 21841 5218
rect 21935 5278 21969 5294
rect 21935 5202 21969 5218
rect 22063 5278 22097 5294
rect 22063 5202 22097 5218
rect 22191 5278 22225 5294
rect 22191 5202 22225 5218
rect 22319 5278 22353 5294
rect 22319 5202 22353 5218
rect 22447 5278 22481 5294
rect 22447 5202 22481 5218
rect 22575 5278 22609 5294
rect 22575 5202 22609 5218
rect 22703 5278 22737 5294
rect 22703 5202 22737 5218
rect 22831 5278 22865 5294
rect 22831 5202 22865 5218
rect 22959 5278 22993 5294
rect 22959 5202 22993 5218
rect 23087 5278 23121 5294
rect 23087 5202 23121 5218
rect 23215 5278 23249 5294
rect 23215 5202 23249 5218
rect 23343 5278 23377 5294
rect 23343 5202 23377 5218
rect 23471 5278 23505 5294
rect 23471 5202 23505 5218
rect 23599 5278 23633 5294
rect 23599 5202 23633 5218
rect 23727 5278 23761 5294
rect 23727 5202 23761 5218
rect 23855 5278 23889 5294
rect 23855 5202 23889 5218
rect 23983 5278 24017 5294
rect 23983 5202 24017 5218
rect 24111 5278 24145 5294
rect 24111 5202 24145 5218
rect 24239 5278 24273 5294
rect 24239 5202 24273 5218
rect 24367 5278 24401 5294
rect 24367 5202 24401 5218
rect 24495 5278 24529 5294
rect 24495 5202 24529 5218
rect 24623 5278 24657 5294
rect 24623 5202 24657 5218
rect 24751 5278 24785 5294
rect 24751 5202 24785 5218
rect 24879 5278 24913 5294
rect 24879 5202 24913 5218
rect 25007 5278 25041 5294
rect 25007 5202 25041 5218
rect 25135 5278 25169 5294
rect 25135 5202 25169 5218
rect 25263 5278 25297 5294
rect 25263 5202 25297 5218
rect 25391 5278 25425 5294
rect 25391 5202 25425 5218
rect 25519 5278 25553 5294
rect 25519 5202 25553 5218
rect 25647 5278 25681 5294
rect 25647 5202 25681 5218
rect 25775 5278 25809 5294
rect 25775 5202 25809 5218
rect 25903 5278 25937 5294
rect 25903 5202 25937 5218
rect 26031 5278 26065 5294
rect 26031 5202 26065 5218
rect 26159 5278 26193 5294
rect 26159 5202 26193 5218
rect 26287 5278 26321 5294
rect 26287 5202 26321 5218
rect 26415 5278 26449 5294
rect 26415 5202 26449 5218
rect 26543 5278 26577 5294
rect 26543 5202 26577 5218
rect 26671 5278 26705 5294
rect 26671 5202 26705 5218
rect 26799 5278 26833 5294
rect 26799 5202 26833 5218
rect 26927 5278 26961 5294
rect 26927 5202 26961 5218
rect 27055 5278 27089 5294
rect 27055 5202 27089 5218
rect 27183 5278 27217 5294
rect 27183 5202 27217 5218
rect 27311 5278 27345 5294
rect 27311 5202 27345 5218
rect 27439 5278 27473 5294
rect 27439 5202 27473 5218
rect 27567 5278 27601 5294
rect 27567 5202 27601 5218
rect 27695 5278 27729 5294
rect 27695 5202 27729 5218
rect 27823 5278 27857 5294
rect 27823 5202 27857 5218
rect 27951 5278 27985 5294
rect 27951 5202 27985 5218
rect 28079 5278 28113 5294
rect 28079 5202 28113 5218
rect 28207 5278 28241 5294
rect 28207 5202 28241 5218
rect 28335 5278 28369 5294
rect 28335 5202 28369 5218
rect 28463 5278 28497 5294
rect 28463 5202 28497 5218
rect -363 5148 28543 5152
rect -363 5110 -319 5148
rect -281 5110 -191 5148
rect -153 5110 609 5148
rect 647 5110 737 5148
rect 775 5110 865 5148
rect 903 5110 1873 5148
rect 1911 5110 2001 5148
rect 2039 5110 2129 5148
rect 2167 5110 2257 5148
rect 2295 5110 2385 5148
rect 2423 5110 3492 5148
rect 3530 5110 3620 5148
rect 3658 5110 3748 5148
rect 3786 5110 3876 5148
rect 3914 5110 4004 5148
rect 4042 5110 4132 5148
rect 4170 5110 4260 5148
rect 4298 5110 4388 5148
rect 4426 5110 4516 5148
rect 4554 5110 8057 5148
rect 8095 5110 8185 5148
rect 8223 5110 8313 5148
rect 8351 5110 8441 5148
rect 8479 5110 8569 5148
rect 8607 5110 8697 5148
rect 8735 5110 8825 5148
rect 8863 5110 8953 5148
rect 8991 5110 9081 5148
rect 9119 5110 9209 5148
rect 9247 5110 9337 5148
rect 9375 5110 9465 5148
rect 9503 5110 9593 5148
rect 9631 5110 9721 5148
rect 9759 5110 9849 5148
rect 9887 5110 9977 5148
rect 10015 5110 10105 5148
rect 10143 5110 15215 5148
rect 15253 5110 15343 5148
rect 15381 5110 15471 5148
rect 15509 5110 15599 5148
rect 15637 5110 15727 5148
rect 15765 5110 15855 5148
rect 15893 5110 15983 5148
rect 16021 5110 16111 5148
rect 16149 5110 16239 5148
rect 16277 5110 16367 5148
rect 16405 5110 16495 5148
rect 16533 5110 16623 5148
rect 16661 5110 16751 5148
rect 16789 5110 16879 5148
rect 16917 5110 17007 5148
rect 17045 5110 17135 5148
rect 17173 5110 17263 5148
rect 17301 5110 17391 5148
rect 17429 5110 17519 5148
rect 17557 5110 17647 5148
rect 17685 5110 17775 5148
rect 17813 5110 17903 5148
rect 17941 5110 18031 5148
rect 18069 5110 18159 5148
rect 18197 5110 18287 5148
rect 18325 5110 18415 5148
rect 18453 5110 18543 5148
rect 18581 5110 18671 5148
rect 18709 5110 18799 5148
rect 18837 5110 18927 5148
rect 18965 5110 19055 5148
rect 19093 5110 19183 5148
rect 19221 5110 19311 5148
rect 19349 5110 20269 5148
rect 20307 5110 20397 5148
rect 20435 5110 20525 5148
rect 20563 5110 20653 5148
rect 20691 5110 20781 5148
rect 20819 5110 20909 5148
rect 20947 5110 21037 5148
rect 21075 5110 21165 5148
rect 21203 5110 21293 5148
rect 21331 5110 21421 5148
rect 21459 5110 21549 5148
rect 21587 5110 21677 5148
rect 21715 5110 21805 5148
rect 21843 5110 21933 5148
rect 21971 5110 22061 5148
rect 22099 5110 22189 5148
rect 22227 5110 22317 5148
rect 22355 5110 22445 5148
rect 22483 5110 22573 5148
rect 22611 5110 22701 5148
rect 22739 5110 22829 5148
rect 22867 5110 22957 5148
rect 22995 5110 23085 5148
rect 23123 5110 23213 5148
rect 23251 5110 23341 5148
rect 23379 5110 23469 5148
rect 23507 5110 23597 5148
rect 23635 5110 23725 5148
rect 23763 5110 23853 5148
rect 23891 5110 23981 5148
rect 24019 5110 24109 5148
rect 24147 5110 24237 5148
rect 24275 5110 24365 5148
rect 24403 5110 24493 5148
rect 24531 5110 24621 5148
rect 24659 5110 24749 5148
rect 24787 5110 24877 5148
rect 24915 5110 25005 5148
rect 25043 5110 25133 5148
rect 25171 5110 25261 5148
rect 25299 5110 25389 5148
rect 25427 5110 25517 5148
rect 25555 5110 25645 5148
rect 25683 5110 25773 5148
rect 25811 5110 25901 5148
rect 25939 5110 26029 5148
rect 26067 5110 26157 5148
rect 26195 5110 26285 5148
rect 26323 5110 26413 5148
rect 26451 5110 26541 5148
rect 26579 5110 26669 5148
rect 26707 5110 26797 5148
rect 26835 5110 26925 5148
rect 26963 5110 27053 5148
rect 27091 5110 27181 5148
rect 27219 5110 27309 5148
rect 27347 5110 27437 5148
rect 27475 5110 27565 5148
rect 27603 5110 27693 5148
rect 27731 5110 27821 5148
rect 27859 5110 27949 5148
rect 27987 5110 28077 5148
rect 28115 5110 28205 5148
rect 28243 5110 28333 5148
rect 28371 5110 28461 5148
rect 28499 5110 28543 5148
rect -363 5106 28543 5110
<< viali >>
rect -297 6378 -259 6416
rect -169 6378 -131 6416
rect 480 6378 518 6416
rect 608 6378 646 6416
rect 736 6378 774 6416
rect 1389 6378 1427 6416
rect 1517 6378 1555 6416
rect 1645 6378 1683 6416
rect 1773 6378 1811 6416
rect 1901 6378 1939 6416
rect 2922 6378 2960 6416
rect 3050 6378 3088 6416
rect 3178 6378 3216 6416
rect 3306 6378 3344 6416
rect 3434 6378 3472 6416
rect 3562 6378 3600 6416
rect 3690 6378 3728 6416
rect 3818 6378 3856 6416
rect 3946 6378 3984 6416
rect 5473 6378 5511 6416
rect 5601 6378 5639 6416
rect 5729 6378 5767 6416
rect 5857 6378 5895 6416
rect 5985 6378 6023 6416
rect 6113 6378 6151 6416
rect 6241 6378 6279 6416
rect 6369 6378 6407 6416
rect 6497 6378 6535 6416
rect 6625 6378 6663 6416
rect 6753 6378 6791 6416
rect 6881 6378 6919 6416
rect 7009 6378 7047 6416
rect 7137 6378 7175 6416
rect 7265 6378 7303 6416
rect 7393 6378 7431 6416
rect 7521 6378 7559 6416
rect 10560 6378 10598 6416
rect 10688 6378 10726 6416
rect 10816 6378 10854 6416
rect 10944 6378 10982 6416
rect 11072 6378 11110 6416
rect 11200 6378 11238 6416
rect 11328 6378 11366 6416
rect 11456 6378 11494 6416
rect 11584 6378 11622 6416
rect 11712 6378 11750 6416
rect 11840 6378 11878 6416
rect 11968 6378 12006 6416
rect 12096 6378 12134 6416
rect 12224 6378 12262 6416
rect 12352 6378 12390 6416
rect 12480 6378 12518 6416
rect 12608 6378 12646 6416
rect 12736 6378 12774 6416
rect 12864 6378 12902 6416
rect 12992 6378 13030 6416
rect 13120 6378 13158 6416
rect 13248 6378 13286 6416
rect 13376 6378 13414 6416
rect 13504 6378 13542 6416
rect 13632 6378 13670 6416
rect 13760 6378 13798 6416
rect 13888 6378 13926 6416
rect 14016 6378 14054 6416
rect 14144 6378 14182 6416
rect 14272 6378 14310 6416
rect 14400 6378 14438 6416
rect 14528 6378 14566 6416
rect 14656 6378 14694 6416
rect 20345 6378 20383 6416
rect 20473 6378 20511 6416
rect 20601 6378 20639 6416
rect 20729 6378 20767 6416
rect 20857 6378 20895 6416
rect 20985 6378 21023 6416
rect 21113 6378 21151 6416
rect 21241 6378 21279 6416
rect 21369 6378 21407 6416
rect 21497 6378 21535 6416
rect 21625 6378 21663 6416
rect 21753 6378 21791 6416
rect 21881 6378 21919 6416
rect 22009 6378 22047 6416
rect 22137 6378 22175 6416
rect 22265 6378 22303 6416
rect 22393 6378 22431 6416
rect 22521 6378 22559 6416
rect 22649 6378 22687 6416
rect 22777 6378 22815 6416
rect 22905 6378 22943 6416
rect 23033 6378 23071 6416
rect 23161 6378 23199 6416
rect 23289 6378 23327 6416
rect 23417 6378 23455 6416
rect 23545 6378 23583 6416
rect 23673 6378 23711 6416
rect 23801 6378 23839 6416
rect 23929 6378 23967 6416
rect 24057 6378 24095 6416
rect 24185 6378 24223 6416
rect 24313 6378 24351 6416
rect 24441 6378 24479 6416
rect 24569 6378 24607 6416
rect 24697 6378 24735 6416
rect 24825 6378 24863 6416
rect 24953 6378 24991 6416
rect 25081 6378 25119 6416
rect 25209 6378 25247 6416
rect 25337 6378 25375 6416
rect 25465 6378 25503 6416
rect 25593 6378 25631 6416
rect 25721 6378 25759 6416
rect 25849 6378 25887 6416
rect 25977 6378 26015 6416
rect 26105 6378 26143 6416
rect 26233 6378 26271 6416
rect 26361 6378 26399 6416
rect 26489 6378 26527 6416
rect 26617 6378 26655 6416
rect 26745 6378 26783 6416
rect 26873 6378 26911 6416
rect 27001 6378 27039 6416
rect 27129 6378 27167 6416
rect 27257 6378 27295 6416
rect 27385 6378 27423 6416
rect 27513 6378 27551 6416
rect 27641 6378 27679 6416
rect 27769 6378 27807 6416
rect 27897 6378 27935 6416
rect 28025 6378 28063 6416
rect 28153 6378 28191 6416
rect 28281 6378 28319 6416
rect 28409 6378 28447 6416
rect 28537 6378 28575 6416
rect -295 6122 -261 6266
rect -167 6122 -133 6266
rect 482 6122 516 6266
rect 610 6122 644 6266
rect 738 6122 772 6266
rect 1391 6122 1425 6266
rect 1519 6122 1553 6266
rect 1647 6122 1681 6266
rect 1775 6122 1809 6266
rect 1903 6122 1937 6266
rect 2924 6122 2958 6266
rect 3052 6122 3086 6266
rect 3180 6122 3214 6266
rect 3308 6122 3342 6266
rect 3436 6122 3470 6266
rect 3564 6122 3598 6266
rect 3692 6122 3726 6266
rect 3820 6122 3854 6266
rect 3948 6122 3982 6266
rect 5475 6122 5509 6266
rect 5603 6122 5637 6266
rect 5731 6122 5765 6266
rect 5859 6122 5893 6266
rect 5987 6122 6021 6266
rect 6115 6122 6149 6266
rect 6243 6122 6277 6266
rect 6371 6122 6405 6266
rect 6499 6122 6533 6266
rect 6627 6122 6661 6266
rect 6755 6122 6789 6266
rect 6883 6122 6917 6266
rect 7011 6122 7045 6266
rect 7139 6122 7173 6266
rect 7267 6122 7301 6266
rect 7395 6122 7429 6266
rect 7523 6122 7557 6266
rect 10562 6122 10596 6266
rect 10690 6122 10724 6266
rect 10818 6122 10852 6266
rect 10946 6122 10980 6266
rect 11074 6122 11108 6266
rect 11202 6122 11236 6266
rect 11330 6122 11364 6266
rect 11458 6122 11492 6266
rect 11586 6122 11620 6266
rect 11714 6122 11748 6266
rect 11842 6122 11876 6266
rect 11970 6122 12004 6266
rect 12098 6122 12132 6266
rect 12226 6122 12260 6266
rect 12354 6122 12388 6266
rect 12482 6122 12516 6266
rect 12610 6122 12644 6266
rect 12738 6122 12772 6266
rect 12866 6122 12900 6266
rect 12994 6122 13028 6266
rect 13122 6122 13156 6266
rect 13250 6122 13284 6266
rect 13378 6122 13412 6266
rect 13506 6122 13540 6266
rect 13634 6122 13668 6266
rect 13762 6122 13796 6266
rect 13890 6122 13924 6266
rect 14018 6122 14052 6266
rect 14146 6122 14180 6266
rect 14274 6122 14308 6266
rect 14402 6122 14436 6266
rect 14530 6122 14564 6266
rect 14658 6122 14692 6266
rect 20347 6122 20381 6266
rect 20475 6122 20509 6266
rect 20603 6122 20637 6266
rect 20731 6122 20765 6266
rect 20859 6122 20893 6266
rect 20987 6122 21021 6266
rect 21115 6122 21149 6266
rect 21243 6122 21277 6266
rect 21371 6122 21405 6266
rect 21499 6122 21533 6266
rect 21627 6122 21661 6266
rect 21755 6122 21789 6266
rect 21883 6122 21917 6266
rect 22011 6122 22045 6266
rect 22139 6122 22173 6266
rect 22267 6122 22301 6266
rect 22395 6122 22429 6266
rect 22523 6122 22557 6266
rect 22651 6122 22685 6266
rect 22779 6122 22813 6266
rect 22907 6122 22941 6266
rect 23035 6122 23069 6266
rect 23163 6122 23197 6266
rect 23291 6122 23325 6266
rect 23419 6122 23453 6266
rect 23547 6122 23581 6266
rect 23675 6122 23709 6266
rect 23803 6122 23837 6266
rect 23931 6122 23965 6266
rect 24059 6122 24093 6266
rect 24187 6122 24221 6266
rect 24315 6122 24349 6266
rect 24443 6122 24477 6266
rect 24571 6122 24605 6266
rect 24699 6122 24733 6266
rect 24827 6122 24861 6266
rect 24955 6122 24989 6266
rect 25083 6122 25117 6266
rect 25211 6122 25245 6266
rect 25339 6122 25373 6266
rect 25467 6122 25501 6266
rect 25595 6122 25629 6266
rect 25723 6122 25757 6266
rect 25851 6122 25885 6266
rect 25979 6122 26013 6266
rect 26107 6122 26141 6266
rect 26235 6122 26269 6266
rect 26363 6122 26397 6266
rect 26491 6122 26525 6266
rect 26619 6122 26653 6266
rect 26747 6122 26781 6266
rect 26875 6122 26909 6266
rect 27003 6122 27037 6266
rect 27131 6122 27165 6266
rect 27259 6122 27293 6266
rect 27387 6122 27421 6266
rect 27515 6122 27549 6266
rect 27643 6122 27677 6266
rect 27771 6122 27805 6266
rect 27899 6122 27933 6266
rect 28027 6122 28061 6266
rect 28155 6122 28189 6266
rect 28283 6122 28317 6266
rect 28411 6122 28445 6266
rect 28539 6122 28573 6266
rect -295 5906 -261 5966
rect -167 5906 -133 5966
rect 482 5906 516 5966
rect 610 5906 644 5966
rect 738 5906 772 5966
rect 1391 5906 1425 5966
rect 1519 5906 1553 5966
rect 1647 5906 1681 5966
rect 1775 5906 1809 5966
rect 1903 5906 1937 5966
rect 2924 5906 2958 5966
rect 3052 5906 3086 5966
rect 3180 5906 3214 5966
rect 3308 5906 3342 5966
rect 3436 5906 3470 5966
rect 3564 5906 3598 5966
rect 3692 5906 3726 5966
rect 3820 5906 3854 5966
rect 3948 5906 3982 5966
rect 5475 5906 5509 5966
rect 5603 5906 5637 5966
rect 5731 5906 5765 5966
rect 5859 5906 5893 5966
rect 5987 5906 6021 5966
rect 6115 5906 6149 5966
rect 6243 5906 6277 5966
rect 6371 5906 6405 5966
rect 6499 5906 6533 5966
rect 6627 5906 6661 5966
rect 6755 5906 6789 5966
rect 6883 5906 6917 5966
rect 7011 5906 7045 5966
rect 7139 5906 7173 5966
rect 7267 5906 7301 5966
rect 7395 5906 7429 5966
rect 7523 5906 7557 5966
rect 10562 5906 10596 5966
rect 10690 5906 10724 5966
rect 10818 5906 10852 5966
rect 10946 5906 10980 5966
rect 11074 5906 11108 5966
rect 11202 5906 11236 5966
rect 11330 5906 11364 5966
rect 11458 5906 11492 5966
rect 11586 5906 11620 5966
rect 11714 5906 11748 5966
rect 11842 5906 11876 5966
rect 11970 5906 12004 5966
rect 12098 5906 12132 5966
rect 12226 5906 12260 5966
rect 12354 5906 12388 5966
rect 12482 5906 12516 5966
rect 12610 5906 12644 5966
rect 12738 5906 12772 5966
rect 12866 5906 12900 5966
rect 12994 5906 13028 5966
rect 13122 5906 13156 5966
rect 13250 5906 13284 5966
rect 13378 5906 13412 5966
rect 13506 5906 13540 5966
rect 13634 5906 13668 5966
rect 13762 5906 13796 5966
rect 13890 5906 13924 5966
rect 14018 5906 14052 5966
rect 14146 5906 14180 5966
rect 14274 5906 14308 5966
rect 14402 5906 14436 5966
rect 14530 5906 14564 5966
rect 14658 5906 14692 5966
rect 20347 5906 20381 5966
rect 20475 5906 20509 5966
rect 20603 5906 20637 5966
rect 20731 5906 20765 5966
rect 20859 5906 20893 5966
rect 20987 5906 21021 5966
rect 21115 5906 21149 5966
rect 21243 5906 21277 5966
rect 21371 5906 21405 5966
rect 21499 5906 21533 5966
rect 21627 5906 21661 5966
rect 21755 5906 21789 5966
rect 21883 5906 21917 5966
rect 22011 5906 22045 5966
rect 22139 5906 22173 5966
rect 22267 5906 22301 5966
rect 22395 5906 22429 5966
rect 22523 5906 22557 5966
rect 22651 5906 22685 5966
rect 22779 5906 22813 5966
rect 22907 5906 22941 5966
rect 23035 5906 23069 5966
rect 23163 5906 23197 5966
rect 23291 5906 23325 5966
rect 23419 5906 23453 5966
rect 23547 5906 23581 5966
rect 23675 5906 23709 5966
rect 23803 5906 23837 5966
rect 23931 5906 23965 5966
rect 24059 5906 24093 5966
rect 24187 5906 24221 5966
rect 24315 5906 24349 5966
rect 24443 5906 24477 5966
rect 24571 5906 24605 5966
rect 24699 5906 24733 5966
rect 24827 5906 24861 5966
rect 24955 5906 24989 5966
rect 25083 5906 25117 5966
rect 25211 5906 25245 5966
rect 25339 5906 25373 5966
rect 25467 5906 25501 5966
rect 25595 5906 25629 5966
rect 25723 5906 25757 5966
rect 25851 5906 25885 5966
rect 25979 5906 26013 5966
rect 26107 5906 26141 5966
rect 26235 5906 26269 5966
rect 26363 5906 26397 5966
rect 26491 5906 26525 5966
rect 26619 5906 26653 5966
rect 26747 5906 26781 5966
rect 26875 5906 26909 5966
rect 27003 5906 27037 5966
rect 27131 5906 27165 5966
rect 27259 5906 27293 5966
rect 27387 5906 27421 5966
rect 27515 5906 27549 5966
rect 27643 5906 27677 5966
rect 27771 5906 27805 5966
rect 27899 5906 27933 5966
rect 28027 5906 28061 5966
rect 28155 5906 28189 5966
rect 28283 5906 28317 5966
rect 28411 5906 28445 5966
rect 28539 5906 28573 5966
rect -297 5798 -259 5836
rect -169 5798 -131 5836
rect 480 5798 518 5836
rect 608 5798 646 5836
rect 736 5798 774 5836
rect 1389 5798 1427 5836
rect 1517 5798 1555 5836
rect 1645 5798 1683 5836
rect 1773 5798 1811 5836
rect 1901 5798 1939 5836
rect 2922 5798 2960 5836
rect 3050 5798 3088 5836
rect 3178 5798 3216 5836
rect 3306 5798 3344 5836
rect 3434 5798 3472 5836
rect 3562 5798 3600 5836
rect 3690 5798 3728 5836
rect 3818 5798 3856 5836
rect 3946 5798 3984 5836
rect 5473 5798 5511 5836
rect 5601 5798 5639 5836
rect 5729 5798 5767 5836
rect 5857 5798 5895 5836
rect 5985 5798 6023 5836
rect 6113 5798 6151 5836
rect 6241 5798 6279 5836
rect 6369 5798 6407 5836
rect 6497 5798 6535 5836
rect 6625 5798 6663 5836
rect 6753 5798 6791 5836
rect 6881 5798 6919 5836
rect 7009 5798 7047 5836
rect 7137 5798 7175 5836
rect 7265 5798 7303 5836
rect 7393 5798 7431 5836
rect 7521 5798 7559 5836
rect 10560 5798 10598 5836
rect 10688 5798 10726 5836
rect 10816 5798 10854 5836
rect 10944 5798 10982 5836
rect 11072 5798 11110 5836
rect 11200 5798 11238 5836
rect 11328 5798 11366 5836
rect 11456 5798 11494 5836
rect 11584 5798 11622 5836
rect 11712 5798 11750 5836
rect 11840 5798 11878 5836
rect 11968 5798 12006 5836
rect 12096 5798 12134 5836
rect 12224 5798 12262 5836
rect 12352 5798 12390 5836
rect 12480 5798 12518 5836
rect 12608 5798 12646 5836
rect 12736 5798 12774 5836
rect 12864 5798 12902 5836
rect 12992 5798 13030 5836
rect 13120 5798 13158 5836
rect 13248 5798 13286 5836
rect 13376 5798 13414 5836
rect 13504 5798 13542 5836
rect 13632 5798 13670 5836
rect 13760 5798 13798 5836
rect 13888 5798 13926 5836
rect 14016 5798 14054 5836
rect 14144 5798 14182 5836
rect 14272 5798 14310 5836
rect 14400 5798 14438 5836
rect 14528 5798 14566 5836
rect 14656 5798 14694 5836
rect 20345 5798 20383 5836
rect 20473 5798 20511 5836
rect 20601 5798 20639 5836
rect 20729 5798 20767 5836
rect 20857 5798 20895 5836
rect 20985 5798 21023 5836
rect 21113 5798 21151 5836
rect 21241 5798 21279 5836
rect 21369 5798 21407 5836
rect 21497 5798 21535 5836
rect 21625 5798 21663 5836
rect 21753 5798 21791 5836
rect 21881 5798 21919 5836
rect 22009 5798 22047 5836
rect 22137 5798 22175 5836
rect 22265 5798 22303 5836
rect 22393 5798 22431 5836
rect 22521 5798 22559 5836
rect 22649 5798 22687 5836
rect 22777 5798 22815 5836
rect 22905 5798 22943 5836
rect 23033 5798 23071 5836
rect 23161 5798 23199 5836
rect 23289 5798 23327 5836
rect 23417 5798 23455 5836
rect 23545 5798 23583 5836
rect 23673 5798 23711 5836
rect 23801 5798 23839 5836
rect 23929 5798 23967 5836
rect 24057 5798 24095 5836
rect 24185 5798 24223 5836
rect 24313 5798 24351 5836
rect 24441 5798 24479 5836
rect 24569 5798 24607 5836
rect 24697 5798 24735 5836
rect 24825 5798 24863 5836
rect 24953 5798 24991 5836
rect 25081 5798 25119 5836
rect 25209 5798 25247 5836
rect 25337 5798 25375 5836
rect 25465 5798 25503 5836
rect 25593 5798 25631 5836
rect 25721 5798 25759 5836
rect 25849 5798 25887 5836
rect 25977 5798 26015 5836
rect 26105 5798 26143 5836
rect 26233 5798 26271 5836
rect 26361 5798 26399 5836
rect 26489 5798 26527 5836
rect 26617 5798 26655 5836
rect 26745 5798 26783 5836
rect 26873 5798 26911 5836
rect 27001 5798 27039 5836
rect 27129 5798 27167 5836
rect 27257 5798 27295 5836
rect 27385 5798 27423 5836
rect 27513 5798 27551 5836
rect 27641 5798 27679 5836
rect 27769 5798 27807 5836
rect 27897 5798 27935 5836
rect 28025 5798 28063 5836
rect 28153 5798 28191 5836
rect 28281 5798 28319 5836
rect 28409 5798 28447 5836
rect 28537 5798 28575 5836
rect -319 5690 -281 5728
rect -191 5690 -153 5728
rect 609 5690 647 5728
rect 737 5690 775 5728
rect 865 5690 903 5728
rect 1873 5690 1911 5728
rect 2001 5690 2039 5728
rect 2129 5690 2167 5728
rect 2257 5690 2295 5728
rect 2385 5690 2423 5728
rect 3492 5690 3530 5728
rect 3620 5690 3658 5728
rect 3748 5690 3786 5728
rect 3876 5690 3914 5728
rect 4004 5690 4042 5728
rect 4132 5690 4170 5728
rect 4260 5690 4298 5728
rect 4388 5690 4426 5728
rect 4516 5690 4554 5728
rect 8057 5690 8095 5728
rect 8185 5690 8223 5728
rect 8313 5690 8351 5728
rect 8441 5690 8479 5728
rect 8569 5690 8607 5728
rect 8697 5690 8735 5728
rect 8825 5690 8863 5728
rect 8953 5690 8991 5728
rect 9081 5690 9119 5728
rect 9209 5690 9247 5728
rect 9337 5690 9375 5728
rect 9465 5690 9503 5728
rect 9593 5690 9631 5728
rect 9721 5690 9759 5728
rect 9849 5690 9887 5728
rect 9977 5690 10015 5728
rect 10105 5690 10143 5728
rect 15215 5690 15253 5728
rect 15343 5690 15381 5728
rect 15471 5690 15509 5728
rect 15599 5690 15637 5728
rect 15727 5690 15765 5728
rect 15855 5690 15893 5728
rect 15983 5690 16021 5728
rect 16111 5690 16149 5728
rect 16239 5690 16277 5728
rect 16367 5690 16405 5728
rect 16495 5690 16533 5728
rect 16623 5690 16661 5728
rect 16751 5690 16789 5728
rect 16879 5690 16917 5728
rect 17007 5690 17045 5728
rect 17135 5690 17173 5728
rect 17263 5690 17301 5728
rect 17391 5690 17429 5728
rect 17519 5690 17557 5728
rect 17647 5690 17685 5728
rect 17775 5690 17813 5728
rect 17903 5690 17941 5728
rect 18031 5690 18069 5728
rect 18159 5690 18197 5728
rect 18287 5690 18325 5728
rect 18415 5690 18453 5728
rect 18543 5690 18581 5728
rect 18671 5690 18709 5728
rect 18799 5690 18837 5728
rect 18927 5690 18965 5728
rect 19055 5690 19093 5728
rect 19183 5690 19221 5728
rect 19311 5690 19349 5728
rect 20269 5690 20307 5728
rect 20397 5690 20435 5728
rect 20525 5690 20563 5728
rect 20653 5690 20691 5728
rect 20781 5690 20819 5728
rect 20909 5690 20947 5728
rect 21037 5690 21075 5728
rect 21165 5690 21203 5728
rect 21293 5690 21331 5728
rect 21421 5690 21459 5728
rect 21549 5690 21587 5728
rect 21677 5690 21715 5728
rect 21805 5690 21843 5728
rect 21933 5690 21971 5728
rect 22061 5690 22099 5728
rect 22189 5690 22227 5728
rect 22317 5690 22355 5728
rect 22445 5690 22483 5728
rect 22573 5690 22611 5728
rect 22701 5690 22739 5728
rect 22829 5690 22867 5728
rect 22957 5690 22995 5728
rect 23085 5690 23123 5728
rect 23213 5690 23251 5728
rect 23341 5690 23379 5728
rect 23469 5690 23507 5728
rect 23597 5690 23635 5728
rect 23725 5690 23763 5728
rect 23853 5690 23891 5728
rect 23981 5690 24019 5728
rect 24109 5690 24147 5728
rect 24237 5690 24275 5728
rect 24365 5690 24403 5728
rect 24493 5690 24531 5728
rect 24621 5690 24659 5728
rect 24749 5690 24787 5728
rect 24877 5690 24915 5728
rect 25005 5690 25043 5728
rect 25133 5690 25171 5728
rect 25261 5690 25299 5728
rect 25389 5690 25427 5728
rect 25517 5690 25555 5728
rect 25645 5690 25683 5728
rect 25773 5690 25811 5728
rect 25901 5690 25939 5728
rect 26029 5690 26067 5728
rect 26157 5690 26195 5728
rect 26285 5690 26323 5728
rect 26413 5690 26451 5728
rect 26541 5690 26579 5728
rect 26669 5690 26707 5728
rect 26797 5690 26835 5728
rect 26925 5690 26963 5728
rect 27053 5690 27091 5728
rect 27181 5690 27219 5728
rect 27309 5690 27347 5728
rect 27437 5690 27475 5728
rect 27565 5690 27603 5728
rect 27693 5690 27731 5728
rect 27821 5690 27859 5728
rect 27949 5690 27987 5728
rect 28077 5690 28115 5728
rect 28205 5690 28243 5728
rect 28333 5690 28371 5728
rect 28461 5690 28499 5728
rect -317 5434 -283 5578
rect -189 5434 -155 5578
rect 611 5434 645 5578
rect 739 5434 773 5578
rect 867 5434 901 5578
rect 1875 5434 1909 5578
rect 2003 5434 2037 5578
rect 2131 5434 2165 5578
rect 2259 5434 2293 5578
rect 2387 5434 2421 5578
rect 3494 5434 3528 5578
rect 3622 5434 3656 5578
rect 3750 5434 3784 5578
rect 3878 5434 3912 5578
rect 4006 5434 4040 5578
rect 4134 5434 4168 5578
rect 4262 5434 4296 5578
rect 4390 5434 4424 5578
rect 4518 5434 4552 5578
rect 8059 5434 8093 5578
rect 8187 5434 8221 5578
rect 8315 5434 8349 5578
rect 8443 5434 8477 5578
rect 8571 5434 8605 5578
rect 8699 5434 8733 5578
rect 8827 5434 8861 5578
rect 8955 5434 8989 5578
rect 9083 5434 9117 5578
rect 9211 5434 9245 5578
rect 9339 5434 9373 5578
rect 9467 5434 9501 5578
rect 9595 5434 9629 5578
rect 9723 5434 9757 5578
rect 9851 5434 9885 5578
rect 9979 5434 10013 5578
rect 10107 5434 10141 5578
rect 15217 5434 15251 5578
rect 15345 5434 15379 5578
rect 15473 5434 15507 5578
rect 15601 5434 15635 5578
rect 15729 5434 15763 5578
rect 15857 5434 15891 5578
rect 15985 5434 16019 5578
rect 16113 5434 16147 5578
rect 16241 5434 16275 5578
rect 16369 5434 16403 5578
rect 16497 5434 16531 5578
rect 16625 5434 16659 5578
rect 16753 5434 16787 5578
rect 16881 5434 16915 5578
rect 17009 5434 17043 5578
rect 17137 5434 17171 5578
rect 17265 5434 17299 5578
rect 17393 5434 17427 5578
rect 17521 5434 17555 5578
rect 17649 5434 17683 5578
rect 17777 5434 17811 5578
rect 17905 5434 17939 5578
rect 18033 5434 18067 5578
rect 18161 5434 18195 5578
rect 18289 5434 18323 5578
rect 18417 5434 18451 5578
rect 18545 5434 18579 5578
rect 18673 5434 18707 5578
rect 18801 5434 18835 5578
rect 18929 5434 18963 5578
rect 19057 5434 19091 5578
rect 19185 5434 19219 5578
rect 19313 5434 19347 5578
rect 20271 5434 20305 5578
rect 20399 5434 20433 5578
rect 20527 5434 20561 5578
rect 20655 5434 20689 5578
rect 20783 5434 20817 5578
rect 20911 5434 20945 5578
rect 21039 5434 21073 5578
rect 21167 5434 21201 5578
rect 21295 5434 21329 5578
rect 21423 5434 21457 5578
rect 21551 5434 21585 5578
rect 21679 5434 21713 5578
rect 21807 5434 21841 5578
rect 21935 5434 21969 5578
rect 22063 5434 22097 5578
rect 22191 5434 22225 5578
rect 22319 5434 22353 5578
rect 22447 5434 22481 5578
rect 22575 5434 22609 5578
rect 22703 5434 22737 5578
rect 22831 5434 22865 5578
rect 22959 5434 22993 5578
rect 23087 5434 23121 5578
rect 23215 5434 23249 5578
rect 23343 5434 23377 5578
rect 23471 5434 23505 5578
rect 23599 5434 23633 5578
rect 23727 5434 23761 5578
rect 23855 5434 23889 5578
rect 23983 5434 24017 5578
rect 24111 5434 24145 5578
rect 24239 5434 24273 5578
rect 24367 5434 24401 5578
rect 24495 5434 24529 5578
rect 24623 5434 24657 5578
rect 24751 5434 24785 5578
rect 24879 5434 24913 5578
rect 25007 5434 25041 5578
rect 25135 5434 25169 5578
rect 25263 5434 25297 5578
rect 25391 5434 25425 5578
rect 25519 5434 25553 5578
rect 25647 5434 25681 5578
rect 25775 5434 25809 5578
rect 25903 5434 25937 5578
rect 26031 5434 26065 5578
rect 26159 5434 26193 5578
rect 26287 5434 26321 5578
rect 26415 5434 26449 5578
rect 26543 5434 26577 5578
rect 26671 5434 26705 5578
rect 26799 5434 26833 5578
rect 26927 5434 26961 5578
rect 27055 5434 27089 5578
rect 27183 5434 27217 5578
rect 27311 5434 27345 5578
rect 27439 5434 27473 5578
rect 27567 5434 27601 5578
rect 27695 5434 27729 5578
rect 27823 5434 27857 5578
rect 27951 5434 27985 5578
rect 28079 5434 28113 5578
rect 28207 5434 28241 5578
rect 28335 5434 28369 5578
rect 28463 5434 28497 5578
rect -317 5218 -283 5278
rect -189 5218 -155 5278
rect 611 5218 645 5278
rect 739 5218 773 5278
rect 867 5218 901 5278
rect 1875 5218 1909 5278
rect 2003 5218 2037 5278
rect 2131 5218 2165 5278
rect 2259 5218 2293 5278
rect 2387 5218 2421 5278
rect 3494 5218 3528 5278
rect 3622 5218 3656 5278
rect 3750 5218 3784 5278
rect 3878 5218 3912 5278
rect 4006 5218 4040 5278
rect 4134 5218 4168 5278
rect 4262 5218 4296 5278
rect 4390 5218 4424 5278
rect 4518 5218 4552 5278
rect 8059 5218 8093 5278
rect 8187 5218 8221 5278
rect 8315 5218 8349 5278
rect 8443 5218 8477 5278
rect 8571 5218 8605 5278
rect 8699 5218 8733 5278
rect 8827 5218 8861 5278
rect 8955 5218 8989 5278
rect 9083 5218 9117 5278
rect 9211 5218 9245 5278
rect 9339 5218 9373 5278
rect 9467 5218 9501 5278
rect 9595 5218 9629 5278
rect 9723 5218 9757 5278
rect 9851 5218 9885 5278
rect 9979 5218 10013 5278
rect 10107 5218 10141 5278
rect 15217 5218 15251 5278
rect 15345 5218 15379 5278
rect 15473 5218 15507 5278
rect 15601 5218 15635 5278
rect 15729 5218 15763 5278
rect 15857 5218 15891 5278
rect 15985 5218 16019 5278
rect 16113 5218 16147 5278
rect 16241 5218 16275 5278
rect 16369 5218 16403 5278
rect 16497 5218 16531 5278
rect 16625 5218 16659 5278
rect 16753 5218 16787 5278
rect 16881 5218 16915 5278
rect 17009 5218 17043 5278
rect 17137 5218 17171 5278
rect 17265 5218 17299 5278
rect 17393 5218 17427 5278
rect 17521 5218 17555 5278
rect 17649 5218 17683 5278
rect 17777 5218 17811 5278
rect 17905 5218 17939 5278
rect 18033 5218 18067 5278
rect 18161 5218 18195 5278
rect 18289 5218 18323 5278
rect 18417 5218 18451 5278
rect 18545 5218 18579 5278
rect 18673 5218 18707 5278
rect 18801 5218 18835 5278
rect 18929 5218 18963 5278
rect 19057 5218 19091 5278
rect 19185 5218 19219 5278
rect 19313 5218 19347 5278
rect 20271 5218 20305 5278
rect 20399 5218 20433 5278
rect 20527 5218 20561 5278
rect 20655 5218 20689 5278
rect 20783 5218 20817 5278
rect 20911 5218 20945 5278
rect 21039 5218 21073 5278
rect 21167 5218 21201 5278
rect 21295 5218 21329 5278
rect 21423 5218 21457 5278
rect 21551 5218 21585 5278
rect 21679 5218 21713 5278
rect 21807 5218 21841 5278
rect 21935 5218 21969 5278
rect 22063 5218 22097 5278
rect 22191 5218 22225 5278
rect 22319 5218 22353 5278
rect 22447 5218 22481 5278
rect 22575 5218 22609 5278
rect 22703 5218 22737 5278
rect 22831 5218 22865 5278
rect 22959 5218 22993 5278
rect 23087 5218 23121 5278
rect 23215 5218 23249 5278
rect 23343 5218 23377 5278
rect 23471 5218 23505 5278
rect 23599 5218 23633 5278
rect 23727 5218 23761 5278
rect 23855 5218 23889 5278
rect 23983 5218 24017 5278
rect 24111 5218 24145 5278
rect 24239 5218 24273 5278
rect 24367 5218 24401 5278
rect 24495 5218 24529 5278
rect 24623 5218 24657 5278
rect 24751 5218 24785 5278
rect 24879 5218 24913 5278
rect 25007 5218 25041 5278
rect 25135 5218 25169 5278
rect 25263 5218 25297 5278
rect 25391 5218 25425 5278
rect 25519 5218 25553 5278
rect 25647 5218 25681 5278
rect 25775 5218 25809 5278
rect 25903 5218 25937 5278
rect 26031 5218 26065 5278
rect 26159 5218 26193 5278
rect 26287 5218 26321 5278
rect 26415 5218 26449 5278
rect 26543 5218 26577 5278
rect 26671 5218 26705 5278
rect 26799 5218 26833 5278
rect 26927 5218 26961 5278
rect 27055 5218 27089 5278
rect 27183 5218 27217 5278
rect 27311 5218 27345 5278
rect 27439 5218 27473 5278
rect 27567 5218 27601 5278
rect 27695 5218 27729 5278
rect 27823 5218 27857 5278
rect 27951 5218 27985 5278
rect 28079 5218 28113 5278
rect 28207 5218 28241 5278
rect 28335 5218 28369 5278
rect 28463 5218 28497 5278
rect -319 5110 -281 5148
rect -191 5110 -153 5148
rect 609 5110 647 5148
rect 737 5110 775 5148
rect 865 5110 903 5148
rect 1873 5110 1911 5148
rect 2001 5110 2039 5148
rect 2129 5110 2167 5148
rect 2257 5110 2295 5148
rect 2385 5110 2423 5148
rect 3492 5110 3530 5148
rect 3620 5110 3658 5148
rect 3748 5110 3786 5148
rect 3876 5110 3914 5148
rect 4004 5110 4042 5148
rect 4132 5110 4170 5148
rect 4260 5110 4298 5148
rect 4388 5110 4426 5148
rect 4516 5110 4554 5148
rect 8057 5110 8095 5148
rect 8185 5110 8223 5148
rect 8313 5110 8351 5148
rect 8441 5110 8479 5148
rect 8569 5110 8607 5148
rect 8697 5110 8735 5148
rect 8825 5110 8863 5148
rect 8953 5110 8991 5148
rect 9081 5110 9119 5148
rect 9209 5110 9247 5148
rect 9337 5110 9375 5148
rect 9465 5110 9503 5148
rect 9593 5110 9631 5148
rect 9721 5110 9759 5148
rect 9849 5110 9887 5148
rect 9977 5110 10015 5148
rect 10105 5110 10143 5148
rect 15215 5110 15253 5148
rect 15343 5110 15381 5148
rect 15471 5110 15509 5148
rect 15599 5110 15637 5148
rect 15727 5110 15765 5148
rect 15855 5110 15893 5148
rect 15983 5110 16021 5148
rect 16111 5110 16149 5148
rect 16239 5110 16277 5148
rect 16367 5110 16405 5148
rect 16495 5110 16533 5148
rect 16623 5110 16661 5148
rect 16751 5110 16789 5148
rect 16879 5110 16917 5148
rect 17007 5110 17045 5148
rect 17135 5110 17173 5148
rect 17263 5110 17301 5148
rect 17391 5110 17429 5148
rect 17519 5110 17557 5148
rect 17647 5110 17685 5148
rect 17775 5110 17813 5148
rect 17903 5110 17941 5148
rect 18031 5110 18069 5148
rect 18159 5110 18197 5148
rect 18287 5110 18325 5148
rect 18415 5110 18453 5148
rect 18543 5110 18581 5148
rect 18671 5110 18709 5148
rect 18799 5110 18837 5148
rect 18927 5110 18965 5148
rect 19055 5110 19093 5148
rect 19183 5110 19221 5148
rect 19311 5110 19349 5148
rect 20269 5110 20307 5148
rect 20397 5110 20435 5148
rect 20525 5110 20563 5148
rect 20653 5110 20691 5148
rect 20781 5110 20819 5148
rect 20909 5110 20947 5148
rect 21037 5110 21075 5148
rect 21165 5110 21203 5148
rect 21293 5110 21331 5148
rect 21421 5110 21459 5148
rect 21549 5110 21587 5148
rect 21677 5110 21715 5148
rect 21805 5110 21843 5148
rect 21933 5110 21971 5148
rect 22061 5110 22099 5148
rect 22189 5110 22227 5148
rect 22317 5110 22355 5148
rect 22445 5110 22483 5148
rect 22573 5110 22611 5148
rect 22701 5110 22739 5148
rect 22829 5110 22867 5148
rect 22957 5110 22995 5148
rect 23085 5110 23123 5148
rect 23213 5110 23251 5148
rect 23341 5110 23379 5148
rect 23469 5110 23507 5148
rect 23597 5110 23635 5148
rect 23725 5110 23763 5148
rect 23853 5110 23891 5148
rect 23981 5110 24019 5148
rect 24109 5110 24147 5148
rect 24237 5110 24275 5148
rect 24365 5110 24403 5148
rect 24493 5110 24531 5148
rect 24621 5110 24659 5148
rect 24749 5110 24787 5148
rect 24877 5110 24915 5148
rect 25005 5110 25043 5148
rect 25133 5110 25171 5148
rect 25261 5110 25299 5148
rect 25389 5110 25427 5148
rect 25517 5110 25555 5148
rect 25645 5110 25683 5148
rect 25773 5110 25811 5148
rect 25901 5110 25939 5148
rect 26029 5110 26067 5148
rect 26157 5110 26195 5148
rect 26285 5110 26323 5148
rect 26413 5110 26451 5148
rect 26541 5110 26579 5148
rect 26669 5110 26707 5148
rect 26797 5110 26835 5148
rect 26925 5110 26963 5148
rect 27053 5110 27091 5148
rect 27181 5110 27219 5148
rect 27309 5110 27347 5148
rect 27437 5110 27475 5148
rect 27565 5110 27603 5148
rect 27693 5110 27731 5148
rect 27821 5110 27859 5148
rect 27949 5110 27987 5148
rect 28077 5110 28115 5148
rect 28205 5110 28243 5148
rect 28333 5110 28371 5148
rect 28461 5110 28499 5148
<< metal1 >>
rect 29502 6422 29566 6426
rect -341 6420 29566 6422
rect -341 6416 29508 6420
rect -341 6378 -297 6416
rect -259 6378 -169 6416
rect -131 6378 480 6416
rect 518 6378 608 6416
rect 646 6378 736 6416
rect 774 6378 1389 6416
rect 1427 6378 1517 6416
rect 1555 6378 1645 6416
rect 1683 6378 1773 6416
rect 1811 6378 1901 6416
rect 1939 6378 2922 6416
rect 2960 6378 3050 6416
rect 3088 6378 3178 6416
rect 3216 6378 3306 6416
rect 3344 6378 3434 6416
rect 3472 6378 3562 6416
rect 3600 6378 3690 6416
rect 3728 6378 3818 6416
rect 3856 6378 3946 6416
rect 3984 6378 5473 6416
rect 5511 6378 5601 6416
rect 5639 6378 5729 6416
rect 5767 6378 5857 6416
rect 5895 6378 5985 6416
rect 6023 6378 6113 6416
rect 6151 6378 6241 6416
rect 6279 6378 6369 6416
rect 6407 6378 6497 6416
rect 6535 6378 6625 6416
rect 6663 6378 6753 6416
rect 6791 6378 6881 6416
rect 6919 6378 7009 6416
rect 7047 6378 7137 6416
rect 7175 6378 7265 6416
rect 7303 6378 7393 6416
rect 7431 6378 7521 6416
rect 7559 6378 10560 6416
rect 10598 6378 10688 6416
rect 10726 6378 10816 6416
rect 10854 6378 10944 6416
rect 10982 6378 11072 6416
rect 11110 6378 11200 6416
rect 11238 6378 11328 6416
rect 11366 6378 11456 6416
rect 11494 6378 11584 6416
rect 11622 6378 11712 6416
rect 11750 6378 11840 6416
rect 11878 6378 11968 6416
rect 12006 6378 12096 6416
rect 12134 6378 12224 6416
rect 12262 6378 12352 6416
rect 12390 6378 12480 6416
rect 12518 6378 12608 6416
rect 12646 6378 12736 6416
rect 12774 6378 12864 6416
rect 12902 6378 12992 6416
rect 13030 6378 13120 6416
rect 13158 6378 13248 6416
rect 13286 6378 13376 6416
rect 13414 6378 13504 6416
rect 13542 6378 13632 6416
rect 13670 6378 13760 6416
rect 13798 6378 13888 6416
rect 13926 6378 14016 6416
rect 14054 6378 14144 6416
rect 14182 6378 14272 6416
rect 14310 6378 14400 6416
rect 14438 6378 14528 6416
rect 14566 6378 14656 6416
rect 14694 6378 20345 6416
rect 20383 6378 20473 6416
rect 20511 6378 20601 6416
rect 20639 6378 20729 6416
rect 20767 6378 20857 6416
rect 20895 6378 20985 6416
rect 21023 6378 21113 6416
rect 21151 6378 21241 6416
rect 21279 6378 21369 6416
rect 21407 6378 21497 6416
rect 21535 6378 21625 6416
rect 21663 6378 21753 6416
rect 21791 6378 21881 6416
rect 21919 6378 22009 6416
rect 22047 6378 22137 6416
rect 22175 6378 22265 6416
rect 22303 6378 22393 6416
rect 22431 6378 22521 6416
rect 22559 6378 22649 6416
rect 22687 6378 22777 6416
rect 22815 6378 22905 6416
rect 22943 6378 23033 6416
rect 23071 6378 23161 6416
rect 23199 6378 23289 6416
rect 23327 6378 23417 6416
rect 23455 6378 23545 6416
rect 23583 6378 23673 6416
rect 23711 6378 23801 6416
rect 23839 6378 23929 6416
rect 23967 6378 24057 6416
rect 24095 6378 24185 6416
rect 24223 6378 24313 6416
rect 24351 6378 24441 6416
rect 24479 6378 24569 6416
rect 24607 6378 24697 6416
rect 24735 6378 24825 6416
rect 24863 6378 24953 6416
rect 24991 6378 25081 6416
rect 25119 6378 25209 6416
rect 25247 6378 25337 6416
rect 25375 6378 25465 6416
rect 25503 6378 25593 6416
rect 25631 6378 25721 6416
rect 25759 6378 25849 6416
rect 25887 6378 25977 6416
rect 26015 6378 26105 6416
rect 26143 6378 26233 6416
rect 26271 6378 26361 6416
rect 26399 6378 26489 6416
rect 26527 6378 26617 6416
rect 26655 6378 26745 6416
rect 26783 6378 26873 6416
rect 26911 6378 27001 6416
rect 27039 6378 27129 6416
rect 27167 6378 27257 6416
rect 27295 6378 27385 6416
rect 27423 6378 27513 6416
rect 27551 6378 27641 6416
rect 27679 6378 27769 6416
rect 27807 6378 27897 6416
rect 27935 6378 28025 6416
rect 28063 6378 28153 6416
rect 28191 6378 28281 6416
rect 28319 6378 28409 6416
rect 28447 6378 28537 6416
rect 28575 6378 29508 6416
rect -341 6372 29508 6378
rect 29502 6368 29508 6372
rect 29560 6368 29566 6420
rect 29502 6362 29566 6368
rect -341 6337 28783 6343
rect -341 6311 28725 6337
rect -295 6278 -261 6311
rect 482 6278 516 6311
rect 738 6278 772 6311
rect 1391 6278 1425 6311
rect 1647 6278 1681 6311
rect 1903 6278 1937 6311
rect 2924 6278 2958 6311
rect 3180 6278 3214 6311
rect 3436 6278 3470 6311
rect 3692 6278 3726 6311
rect 3948 6278 3982 6311
rect 5475 6278 5509 6311
rect 5731 6278 5765 6311
rect 5987 6278 6021 6311
rect 6243 6278 6277 6311
rect 6499 6278 6533 6311
rect 6755 6278 6789 6311
rect 7011 6278 7045 6311
rect 7267 6278 7301 6311
rect 7523 6278 7557 6311
rect 10562 6278 10596 6311
rect 10818 6278 10852 6311
rect 11074 6278 11108 6311
rect 11330 6278 11364 6311
rect 11586 6278 11620 6311
rect 11842 6278 11876 6311
rect 12098 6278 12132 6311
rect 12354 6278 12388 6311
rect 12610 6278 12644 6311
rect 12866 6278 12900 6311
rect 13122 6278 13156 6311
rect 13378 6278 13412 6311
rect 13634 6278 13668 6311
rect 13890 6278 13924 6311
rect 14146 6278 14180 6311
rect 14402 6278 14436 6311
rect 14658 6278 14692 6311
rect 20347 6278 20381 6311
rect 20603 6278 20637 6311
rect 20859 6278 20893 6311
rect 21115 6278 21149 6311
rect 21371 6278 21405 6311
rect 21627 6278 21661 6311
rect 21883 6278 21917 6311
rect 22139 6278 22173 6311
rect 22395 6278 22429 6311
rect 22651 6278 22685 6311
rect 22907 6278 22941 6311
rect 23163 6278 23197 6311
rect 23419 6278 23453 6311
rect 23675 6278 23709 6311
rect 23931 6278 23965 6311
rect 24187 6278 24221 6311
rect 24443 6278 24477 6311
rect 24699 6278 24733 6311
rect 24955 6278 24989 6311
rect 25211 6278 25245 6311
rect 25467 6278 25501 6311
rect 25723 6278 25757 6311
rect 25979 6278 26013 6311
rect 26235 6278 26269 6311
rect 26491 6278 26525 6311
rect 26747 6278 26781 6311
rect 27003 6278 27037 6311
rect 27259 6278 27293 6311
rect 27515 6278 27549 6311
rect 27771 6278 27805 6311
rect 28027 6278 28061 6311
rect 28283 6278 28317 6311
rect 28539 6278 28573 6311
rect 28719 6285 28725 6311
rect 28777 6285 28783 6337
rect 28719 6279 28783 6285
rect -301 6266 -255 6278
rect -301 6122 -295 6266
rect -261 6122 -255 6266
rect -301 6110 -255 6122
rect -173 6266 -127 6278
rect -173 6122 -167 6266
rect -133 6122 -127 6266
rect -173 6110 -127 6122
rect 476 6266 522 6278
rect 476 6122 482 6266
rect 516 6122 522 6266
rect 476 6110 522 6122
rect 604 6266 650 6278
rect 604 6122 610 6266
rect 644 6122 650 6266
rect 604 6110 650 6122
rect 732 6266 778 6278
rect 732 6122 738 6266
rect 772 6122 778 6266
rect 732 6110 778 6122
rect 1385 6266 1431 6278
rect 1385 6122 1391 6266
rect 1425 6122 1431 6266
rect 1385 6110 1431 6122
rect 1513 6266 1559 6278
rect 1513 6122 1519 6266
rect 1553 6122 1559 6266
rect 1513 6110 1559 6122
rect 1641 6266 1687 6278
rect 1641 6122 1647 6266
rect 1681 6122 1687 6266
rect 1641 6110 1687 6122
rect 1769 6266 1815 6278
rect 1769 6122 1775 6266
rect 1809 6122 1815 6266
rect 1769 6110 1815 6122
rect 1897 6266 1943 6278
rect 1897 6122 1903 6266
rect 1937 6122 1943 6266
rect 1897 6110 1943 6122
rect 2918 6266 2964 6278
rect 2918 6122 2924 6266
rect 2958 6122 2964 6266
rect 2918 6110 2964 6122
rect 3046 6266 3092 6278
rect 3046 6122 3052 6266
rect 3086 6122 3092 6266
rect 3046 6110 3092 6122
rect 3174 6266 3220 6278
rect 3174 6122 3180 6266
rect 3214 6122 3220 6266
rect 3174 6110 3220 6122
rect 3302 6266 3348 6278
rect 3302 6122 3308 6266
rect 3342 6122 3348 6266
rect 3302 6110 3348 6122
rect 3430 6266 3476 6278
rect 3430 6122 3436 6266
rect 3470 6122 3476 6266
rect 3430 6110 3476 6122
rect 3558 6266 3604 6278
rect 3558 6122 3564 6266
rect 3598 6122 3604 6266
rect 3558 6110 3604 6122
rect 3686 6266 3732 6278
rect 3686 6122 3692 6266
rect 3726 6122 3732 6266
rect 3686 6110 3732 6122
rect 3814 6266 3860 6278
rect 3814 6122 3820 6266
rect 3854 6122 3860 6266
rect 3814 6110 3860 6122
rect 3942 6266 3988 6278
rect 3942 6122 3948 6266
rect 3982 6122 3988 6266
rect 3942 6110 3988 6122
rect 5469 6266 5515 6278
rect 5469 6122 5475 6266
rect 5509 6122 5515 6266
rect 5469 6110 5515 6122
rect 5597 6266 5643 6278
rect 5597 6122 5603 6266
rect 5637 6122 5643 6266
rect 5597 6110 5643 6122
rect 5725 6266 5771 6278
rect 5725 6122 5731 6266
rect 5765 6122 5771 6266
rect 5725 6110 5771 6122
rect 5853 6266 5899 6278
rect 5853 6122 5859 6266
rect 5893 6122 5899 6266
rect 5853 6110 5899 6122
rect 5981 6266 6027 6278
rect 5981 6122 5987 6266
rect 6021 6122 6027 6266
rect 5981 6110 6027 6122
rect 6109 6266 6155 6278
rect 6109 6122 6115 6266
rect 6149 6122 6155 6266
rect 6109 6110 6155 6122
rect 6237 6266 6283 6278
rect 6237 6122 6243 6266
rect 6277 6122 6283 6266
rect 6237 6110 6283 6122
rect 6365 6266 6411 6278
rect 6365 6122 6371 6266
rect 6405 6122 6411 6266
rect 6365 6110 6411 6122
rect 6493 6266 6539 6278
rect 6493 6122 6499 6266
rect 6533 6122 6539 6266
rect 6493 6110 6539 6122
rect 6621 6266 6667 6278
rect 6621 6122 6627 6266
rect 6661 6122 6667 6266
rect 6621 6110 6667 6122
rect 6749 6266 6795 6278
rect 6749 6122 6755 6266
rect 6789 6122 6795 6266
rect 6749 6110 6795 6122
rect 6877 6266 6923 6278
rect 6877 6122 6883 6266
rect 6917 6122 6923 6266
rect 6877 6110 6923 6122
rect 7005 6266 7051 6278
rect 7005 6122 7011 6266
rect 7045 6122 7051 6266
rect 7005 6110 7051 6122
rect 7133 6266 7179 6278
rect 7133 6122 7139 6266
rect 7173 6122 7179 6266
rect 7133 6110 7179 6122
rect 7261 6266 7307 6278
rect 7261 6122 7267 6266
rect 7301 6122 7307 6266
rect 7261 6110 7307 6122
rect 7389 6266 7435 6278
rect 7389 6122 7395 6266
rect 7429 6122 7435 6266
rect 7389 6110 7435 6122
rect 7517 6266 7563 6278
rect 7517 6122 7523 6266
rect 7557 6122 7563 6266
rect 7517 6110 7563 6122
rect 10556 6266 10602 6278
rect 10556 6122 10562 6266
rect 10596 6122 10602 6266
rect 10556 6110 10602 6122
rect 10684 6266 10730 6278
rect 10684 6122 10690 6266
rect 10724 6122 10730 6266
rect 10684 6110 10730 6122
rect 10812 6266 10858 6278
rect 10812 6122 10818 6266
rect 10852 6122 10858 6266
rect 10812 6110 10858 6122
rect 10940 6266 10986 6278
rect 10940 6122 10946 6266
rect 10980 6122 10986 6266
rect 10940 6110 10986 6122
rect 11068 6266 11114 6278
rect 11068 6122 11074 6266
rect 11108 6122 11114 6266
rect 11068 6110 11114 6122
rect 11196 6266 11242 6278
rect 11196 6122 11202 6266
rect 11236 6122 11242 6266
rect 11196 6110 11242 6122
rect 11324 6266 11370 6278
rect 11324 6122 11330 6266
rect 11364 6122 11370 6266
rect 11324 6110 11370 6122
rect 11452 6266 11498 6278
rect 11452 6122 11458 6266
rect 11492 6122 11498 6266
rect 11452 6110 11498 6122
rect 11580 6266 11626 6278
rect 11580 6122 11586 6266
rect 11620 6122 11626 6266
rect 11580 6110 11626 6122
rect 11708 6266 11754 6278
rect 11708 6122 11714 6266
rect 11748 6122 11754 6266
rect 11708 6110 11754 6122
rect 11836 6266 11882 6278
rect 11836 6122 11842 6266
rect 11876 6122 11882 6266
rect 11836 6110 11882 6122
rect 11964 6266 12010 6278
rect 11964 6122 11970 6266
rect 12004 6122 12010 6266
rect 11964 6110 12010 6122
rect 12092 6266 12138 6278
rect 12092 6122 12098 6266
rect 12132 6122 12138 6266
rect 12092 6110 12138 6122
rect 12220 6266 12266 6278
rect 12220 6122 12226 6266
rect 12260 6122 12266 6266
rect 12220 6110 12266 6122
rect 12348 6266 12394 6278
rect 12348 6122 12354 6266
rect 12388 6122 12394 6266
rect 12348 6110 12394 6122
rect 12476 6266 12522 6278
rect 12476 6122 12482 6266
rect 12516 6122 12522 6266
rect 12476 6110 12522 6122
rect 12604 6266 12650 6278
rect 12604 6122 12610 6266
rect 12644 6122 12650 6266
rect 12604 6110 12650 6122
rect 12732 6266 12778 6278
rect 12732 6122 12738 6266
rect 12772 6122 12778 6266
rect 12732 6110 12778 6122
rect 12860 6266 12906 6278
rect 12860 6122 12866 6266
rect 12900 6122 12906 6266
rect 12860 6110 12906 6122
rect 12988 6266 13034 6278
rect 12988 6122 12994 6266
rect 13028 6122 13034 6266
rect 12988 6110 13034 6122
rect 13116 6266 13162 6278
rect 13116 6122 13122 6266
rect 13156 6122 13162 6266
rect 13116 6110 13162 6122
rect 13244 6266 13290 6278
rect 13244 6122 13250 6266
rect 13284 6122 13290 6266
rect 13244 6110 13290 6122
rect 13372 6266 13418 6278
rect 13372 6122 13378 6266
rect 13412 6122 13418 6266
rect 13372 6110 13418 6122
rect 13500 6266 13546 6278
rect 13500 6122 13506 6266
rect 13540 6122 13546 6266
rect 13500 6110 13546 6122
rect 13628 6266 13674 6278
rect 13628 6122 13634 6266
rect 13668 6122 13674 6266
rect 13628 6110 13674 6122
rect 13756 6266 13802 6278
rect 13756 6122 13762 6266
rect 13796 6122 13802 6266
rect 13756 6110 13802 6122
rect 13884 6266 13930 6278
rect 13884 6122 13890 6266
rect 13924 6122 13930 6266
rect 13884 6110 13930 6122
rect 14012 6266 14058 6278
rect 14012 6122 14018 6266
rect 14052 6122 14058 6266
rect 14012 6110 14058 6122
rect 14140 6266 14186 6278
rect 14140 6122 14146 6266
rect 14180 6122 14186 6266
rect 14140 6110 14186 6122
rect 14268 6266 14314 6278
rect 14268 6122 14274 6266
rect 14308 6122 14314 6266
rect 14268 6110 14314 6122
rect 14396 6266 14442 6278
rect 14396 6122 14402 6266
rect 14436 6122 14442 6266
rect 14396 6110 14442 6122
rect 14524 6266 14570 6278
rect 14524 6122 14530 6266
rect 14564 6122 14570 6266
rect 14524 6110 14570 6122
rect 14652 6266 14698 6278
rect 14652 6122 14658 6266
rect 14692 6122 14698 6266
rect 14652 6110 14698 6122
rect 20341 6266 20387 6278
rect 20341 6122 20347 6266
rect 20381 6122 20387 6266
rect 20341 6110 20387 6122
rect 20469 6266 20515 6278
rect 20469 6122 20475 6266
rect 20509 6122 20515 6266
rect 20469 6110 20515 6122
rect 20597 6266 20643 6278
rect 20597 6122 20603 6266
rect 20637 6122 20643 6266
rect 20597 6110 20643 6122
rect 20725 6266 20771 6278
rect 20725 6122 20731 6266
rect 20765 6122 20771 6266
rect 20725 6110 20771 6122
rect 20853 6266 20899 6278
rect 20853 6122 20859 6266
rect 20893 6122 20899 6266
rect 20853 6110 20899 6122
rect 20981 6266 21027 6278
rect 20981 6122 20987 6266
rect 21021 6122 21027 6266
rect 20981 6110 21027 6122
rect 21109 6266 21155 6278
rect 21109 6122 21115 6266
rect 21149 6122 21155 6266
rect 21109 6110 21155 6122
rect 21237 6266 21283 6278
rect 21237 6122 21243 6266
rect 21277 6122 21283 6266
rect 21237 6110 21283 6122
rect 21365 6266 21411 6278
rect 21365 6122 21371 6266
rect 21405 6122 21411 6266
rect 21365 6110 21411 6122
rect 21493 6266 21539 6278
rect 21493 6122 21499 6266
rect 21533 6122 21539 6266
rect 21493 6110 21539 6122
rect 21621 6266 21667 6278
rect 21621 6122 21627 6266
rect 21661 6122 21667 6266
rect 21621 6110 21667 6122
rect 21749 6266 21795 6278
rect 21749 6122 21755 6266
rect 21789 6122 21795 6266
rect 21749 6110 21795 6122
rect 21877 6266 21923 6278
rect 21877 6122 21883 6266
rect 21917 6122 21923 6266
rect 21877 6110 21923 6122
rect 22005 6266 22051 6278
rect 22005 6122 22011 6266
rect 22045 6122 22051 6266
rect 22005 6110 22051 6122
rect 22133 6266 22179 6278
rect 22133 6122 22139 6266
rect 22173 6122 22179 6266
rect 22133 6110 22179 6122
rect 22261 6266 22307 6278
rect 22261 6122 22267 6266
rect 22301 6122 22307 6266
rect 22261 6110 22307 6122
rect 22389 6266 22435 6278
rect 22389 6122 22395 6266
rect 22429 6122 22435 6266
rect 22389 6110 22435 6122
rect 22517 6266 22563 6278
rect 22517 6122 22523 6266
rect 22557 6122 22563 6266
rect 22517 6110 22563 6122
rect 22645 6266 22691 6278
rect 22645 6122 22651 6266
rect 22685 6122 22691 6266
rect 22645 6110 22691 6122
rect 22773 6266 22819 6278
rect 22773 6122 22779 6266
rect 22813 6122 22819 6266
rect 22773 6110 22819 6122
rect 22901 6266 22947 6278
rect 22901 6122 22907 6266
rect 22941 6122 22947 6266
rect 22901 6110 22947 6122
rect 23029 6266 23075 6278
rect 23029 6122 23035 6266
rect 23069 6122 23075 6266
rect 23029 6110 23075 6122
rect 23157 6266 23203 6278
rect 23157 6122 23163 6266
rect 23197 6122 23203 6266
rect 23157 6110 23203 6122
rect 23285 6266 23331 6278
rect 23285 6122 23291 6266
rect 23325 6122 23331 6266
rect 23285 6110 23331 6122
rect 23413 6266 23459 6278
rect 23413 6122 23419 6266
rect 23453 6122 23459 6266
rect 23413 6110 23459 6122
rect 23541 6266 23587 6278
rect 23541 6122 23547 6266
rect 23581 6122 23587 6266
rect 23541 6110 23587 6122
rect 23669 6266 23715 6278
rect 23669 6122 23675 6266
rect 23709 6122 23715 6266
rect 23669 6110 23715 6122
rect 23797 6266 23843 6278
rect 23797 6122 23803 6266
rect 23837 6122 23843 6266
rect 23797 6110 23843 6122
rect 23925 6266 23971 6278
rect 23925 6122 23931 6266
rect 23965 6122 23971 6266
rect 23925 6110 23971 6122
rect 24053 6266 24099 6278
rect 24053 6122 24059 6266
rect 24093 6122 24099 6266
rect 24053 6110 24099 6122
rect 24181 6266 24227 6278
rect 24181 6122 24187 6266
rect 24221 6122 24227 6266
rect 24181 6110 24227 6122
rect 24309 6266 24355 6278
rect 24309 6122 24315 6266
rect 24349 6122 24355 6266
rect 24309 6110 24355 6122
rect 24437 6266 24483 6278
rect 24437 6122 24443 6266
rect 24477 6122 24483 6266
rect 24437 6110 24483 6122
rect 24565 6266 24611 6278
rect 24565 6122 24571 6266
rect 24605 6122 24611 6266
rect 24565 6110 24611 6122
rect 24693 6266 24739 6278
rect 24693 6122 24699 6266
rect 24733 6122 24739 6266
rect 24693 6110 24739 6122
rect 24821 6266 24867 6278
rect 24821 6122 24827 6266
rect 24861 6122 24867 6266
rect 24821 6110 24867 6122
rect 24949 6266 24995 6278
rect 24949 6122 24955 6266
rect 24989 6122 24995 6266
rect 24949 6110 24995 6122
rect 25077 6266 25123 6278
rect 25077 6122 25083 6266
rect 25117 6122 25123 6266
rect 25077 6110 25123 6122
rect 25205 6266 25251 6278
rect 25205 6122 25211 6266
rect 25245 6122 25251 6266
rect 25205 6110 25251 6122
rect 25333 6266 25379 6278
rect 25333 6122 25339 6266
rect 25373 6122 25379 6266
rect 25333 6110 25379 6122
rect 25461 6266 25507 6278
rect 25461 6122 25467 6266
rect 25501 6122 25507 6266
rect 25461 6110 25507 6122
rect 25589 6266 25635 6278
rect 25589 6122 25595 6266
rect 25629 6122 25635 6266
rect 25589 6110 25635 6122
rect 25717 6266 25763 6278
rect 25717 6122 25723 6266
rect 25757 6122 25763 6266
rect 25717 6110 25763 6122
rect 25845 6266 25891 6278
rect 25845 6122 25851 6266
rect 25885 6122 25891 6266
rect 25845 6110 25891 6122
rect 25973 6266 26019 6278
rect 25973 6122 25979 6266
rect 26013 6122 26019 6266
rect 25973 6110 26019 6122
rect 26101 6266 26147 6278
rect 26101 6122 26107 6266
rect 26141 6122 26147 6266
rect 26101 6110 26147 6122
rect 26229 6266 26275 6278
rect 26229 6122 26235 6266
rect 26269 6122 26275 6266
rect 26229 6110 26275 6122
rect 26357 6266 26403 6278
rect 26357 6122 26363 6266
rect 26397 6122 26403 6266
rect 26357 6110 26403 6122
rect 26485 6266 26531 6278
rect 26485 6122 26491 6266
rect 26525 6122 26531 6266
rect 26485 6110 26531 6122
rect 26613 6266 26659 6278
rect 26613 6122 26619 6266
rect 26653 6122 26659 6266
rect 26613 6110 26659 6122
rect 26741 6266 26787 6278
rect 26741 6122 26747 6266
rect 26781 6122 26787 6266
rect 26741 6110 26787 6122
rect 26869 6266 26915 6278
rect 26869 6122 26875 6266
rect 26909 6122 26915 6266
rect 26869 6110 26915 6122
rect 26997 6266 27043 6278
rect 26997 6122 27003 6266
rect 27037 6122 27043 6266
rect 26997 6110 27043 6122
rect 27125 6266 27171 6278
rect 27125 6122 27131 6266
rect 27165 6122 27171 6266
rect 27125 6110 27171 6122
rect 27253 6266 27299 6278
rect 27253 6122 27259 6266
rect 27293 6122 27299 6266
rect 27253 6110 27299 6122
rect 27381 6266 27427 6278
rect 27381 6122 27387 6266
rect 27421 6122 27427 6266
rect 27381 6110 27427 6122
rect 27509 6266 27555 6278
rect 27509 6122 27515 6266
rect 27549 6122 27555 6266
rect 27509 6110 27555 6122
rect 27637 6266 27683 6278
rect 27637 6122 27643 6266
rect 27677 6122 27683 6266
rect 27637 6110 27683 6122
rect 27765 6266 27811 6278
rect 27765 6122 27771 6266
rect 27805 6122 27811 6266
rect 27765 6110 27811 6122
rect 27893 6266 27939 6278
rect 27893 6122 27899 6266
rect 27933 6122 27939 6266
rect 27893 6110 27939 6122
rect 28021 6266 28067 6278
rect 28021 6122 28027 6266
rect 28061 6122 28067 6266
rect 28021 6110 28067 6122
rect 28149 6266 28195 6278
rect 28149 6122 28155 6266
rect 28189 6122 28195 6266
rect 28149 6110 28195 6122
rect 28277 6266 28323 6278
rect 28277 6122 28283 6266
rect 28317 6122 28323 6266
rect 28277 6110 28323 6122
rect 28405 6266 28451 6278
rect 28405 6122 28411 6266
rect 28445 6122 28451 6266
rect 28405 6110 28451 6122
rect 28533 6266 28579 6278
rect 28533 6122 28539 6266
rect 28573 6122 28579 6266
rect 28533 6110 28579 6122
rect -167 6073 -133 6110
rect -95 6083 -31 6089
rect -95 6073 -89 6083
rect -167 6040 -89 6073
rect -167 5978 -133 6040
rect -95 6031 -89 6040
rect -37 6031 -31 6083
rect -95 6025 -31 6031
rect 357 6061 421 6067
rect 357 6009 363 6061
rect 415 6053 421 6061
rect 610 6053 644 6110
rect 415 6017 644 6053
rect 415 6009 421 6017
rect 357 6003 421 6009
rect 610 5978 644 6017
rect 1268 6061 1332 6067
rect 1268 6009 1274 6061
rect 1326 6050 1332 6061
rect 1519 6050 1553 6110
rect 1326 6036 1553 6050
rect 1775 6036 1809 6110
rect 1326 6019 1809 6036
rect 1326 6009 1332 6019
rect 1268 6003 1332 6009
rect 1519 6007 1809 6019
rect 1519 5978 1553 6007
rect 1775 5978 1809 6007
rect 2803 6049 2867 6055
rect 2803 5997 2809 6049
rect 2861 6038 2867 6049
rect 3052 6038 3086 6110
rect 2861 6036 3086 6038
rect 3308 6036 3342 6110
rect 3564 6036 3598 6110
rect 3820 6036 3854 6110
rect 2861 6009 3854 6036
rect 2861 5997 2867 6009
rect 2803 5991 2867 5997
rect 3052 6007 3854 6009
rect 3052 5978 3086 6007
rect 3308 5978 3342 6007
rect 3564 5978 3598 6007
rect 3820 5978 3854 6007
rect 5353 6047 5417 6053
rect 5353 5995 5359 6047
rect 5411 6036 5417 6047
rect 5603 6036 5637 6110
rect 5859 6036 5893 6110
rect 6115 6036 6149 6110
rect 6371 6036 6405 6110
rect 6627 6036 6661 6110
rect 6883 6036 6917 6110
rect 7139 6036 7173 6110
rect 7395 6036 7429 6110
rect 5411 6007 7429 6036
rect 5411 5995 5417 6007
rect 5353 5989 5417 5995
rect 5603 5978 5637 6007
rect 5859 5978 5893 6007
rect 6115 5978 6149 6007
rect 6371 5978 6405 6007
rect 6627 5978 6661 6007
rect 6883 5978 6917 6007
rect 7139 5978 7173 6007
rect 7395 5978 7429 6007
rect 10326 6047 10390 6053
rect 10326 5995 10332 6047
rect 10384 6036 10390 6047
rect 10690 6036 10724 6110
rect 10946 6036 10980 6110
rect 11202 6036 11236 6110
rect 11458 6036 11492 6110
rect 11714 6036 11748 6110
rect 11970 6036 12004 6110
rect 12226 6036 12260 6110
rect 12482 6036 12516 6110
rect 12738 6036 12772 6110
rect 12994 6036 13028 6110
rect 13250 6036 13284 6110
rect 13506 6036 13540 6110
rect 13762 6036 13796 6110
rect 14018 6036 14052 6110
rect 14274 6036 14308 6110
rect 14530 6036 14564 6110
rect 10384 6007 14564 6036
rect 10384 6006 10724 6007
rect 10384 5995 10390 6006
rect 10326 5989 10390 5995
rect 10690 5978 10724 6006
rect 10946 5978 10980 6007
rect 11202 5978 11236 6007
rect 11458 5978 11492 6007
rect 11714 5978 11748 6007
rect 11970 5978 12004 6007
rect 12226 5978 12260 6007
rect 12482 5978 12516 6007
rect 12738 5978 12772 6007
rect 12994 5978 13028 6007
rect 13250 5978 13284 6007
rect 13506 5978 13540 6007
rect 13762 5978 13796 6007
rect 14018 5978 14052 6007
rect 14274 5978 14308 6007
rect 14530 5978 14564 6007
rect 20475 6036 20509 6110
rect 20731 6036 20765 6110
rect 20987 6036 21021 6110
rect 21243 6036 21277 6110
rect 21499 6036 21533 6110
rect 21755 6036 21789 6110
rect 22011 6036 22045 6110
rect 22267 6036 22301 6110
rect 22523 6036 22557 6110
rect 22779 6036 22813 6110
rect 23035 6036 23069 6110
rect 23291 6036 23325 6110
rect 23547 6036 23581 6110
rect 23803 6036 23837 6110
rect 24059 6036 24093 6110
rect 24315 6036 24349 6110
rect 24571 6036 24605 6110
rect 24827 6036 24861 6110
rect 25083 6036 25117 6110
rect 25339 6036 25373 6110
rect 25595 6036 25629 6110
rect 25851 6036 25885 6110
rect 26107 6036 26141 6110
rect 26363 6036 26397 6110
rect 26619 6036 26653 6110
rect 26875 6036 26909 6110
rect 27131 6036 27165 6110
rect 27387 6036 27421 6110
rect 27643 6036 27677 6110
rect 27899 6036 27933 6110
rect 28155 6036 28189 6110
rect 28411 6036 28445 6110
rect 28631 6047 28695 6053
rect 28631 6036 28637 6047
rect 20475 6007 28637 6036
rect 20475 5978 20509 6007
rect 20731 5978 20765 6007
rect 20987 5978 21021 6007
rect 21243 5978 21277 6007
rect 21499 5978 21533 6007
rect 21755 5978 21789 6007
rect 22011 5978 22045 6007
rect 22267 5978 22301 6007
rect 22523 5978 22557 6007
rect 22779 5978 22813 6007
rect 23035 5978 23069 6007
rect 23291 5978 23325 6007
rect 23547 5978 23581 6007
rect 23803 5978 23837 6007
rect 24059 5978 24093 6007
rect 24315 5978 24349 6007
rect 24571 5978 24605 6007
rect 24827 5978 24861 6007
rect 25083 5978 25117 6007
rect 25339 5978 25373 6007
rect 25595 5978 25629 6007
rect 25851 5978 25885 6007
rect 26107 5978 26141 6007
rect 26363 5978 26397 6007
rect 26619 5978 26653 6007
rect 26875 5978 26909 6007
rect 27131 5978 27165 6007
rect 27387 5978 27421 6007
rect 27643 5978 27677 6007
rect 27899 5978 27933 6007
rect 28155 5978 28189 6007
rect 28411 5978 28445 6007
rect 28631 5995 28637 6007
rect 28689 5995 28695 6047
rect 28631 5989 28695 5995
rect -301 5966 -255 5978
rect -301 5906 -295 5966
rect -261 5906 -255 5966
rect -301 5894 -255 5906
rect -173 5966 -127 5978
rect -173 5906 -167 5966
rect -133 5906 -127 5966
rect -173 5894 -127 5906
rect 476 5966 522 5978
rect 476 5906 482 5966
rect 516 5906 522 5966
rect 476 5894 522 5906
rect 604 5966 650 5978
rect 604 5906 610 5966
rect 644 5906 650 5966
rect 604 5894 650 5906
rect 732 5966 778 5978
rect 732 5906 738 5966
rect 772 5906 778 5966
rect 732 5894 778 5906
rect 1385 5966 1431 5978
rect 1385 5906 1391 5966
rect 1425 5906 1431 5966
rect 1385 5894 1431 5906
rect 1513 5966 1559 5978
rect 1513 5906 1519 5966
rect 1553 5906 1559 5966
rect 1513 5894 1559 5906
rect 1641 5966 1687 5978
rect 1641 5906 1647 5966
rect 1681 5906 1687 5966
rect 1641 5894 1687 5906
rect 1769 5966 1815 5978
rect 1769 5906 1775 5966
rect 1809 5906 1815 5966
rect 1769 5894 1815 5906
rect 1897 5966 1943 5978
rect 1897 5906 1903 5966
rect 1937 5906 1943 5966
rect 1897 5894 1943 5906
rect 2918 5966 2964 5978
rect 2918 5906 2924 5966
rect 2958 5906 2964 5966
rect 2918 5894 2964 5906
rect 3046 5966 3092 5978
rect 3046 5906 3052 5966
rect 3086 5906 3092 5966
rect 3046 5894 3092 5906
rect 3174 5966 3220 5978
rect 3174 5906 3180 5966
rect 3214 5906 3220 5966
rect 3174 5894 3220 5906
rect 3302 5966 3348 5978
rect 3302 5906 3308 5966
rect 3342 5906 3348 5966
rect 3302 5894 3348 5906
rect 3430 5966 3476 5978
rect 3430 5906 3436 5966
rect 3470 5906 3476 5966
rect 3430 5894 3476 5906
rect 3558 5966 3604 5978
rect 3558 5906 3564 5966
rect 3598 5906 3604 5966
rect 3558 5894 3604 5906
rect 3686 5966 3732 5978
rect 3686 5906 3692 5966
rect 3726 5906 3732 5966
rect 3686 5894 3732 5906
rect 3814 5966 3860 5978
rect 3814 5906 3820 5966
rect 3854 5906 3860 5966
rect 3814 5894 3860 5906
rect 3942 5966 3988 5978
rect 3942 5906 3948 5966
rect 3982 5906 3988 5966
rect 3942 5894 3988 5906
rect 5469 5966 5515 5978
rect 5469 5906 5475 5966
rect 5509 5906 5515 5966
rect 5469 5894 5515 5906
rect 5597 5966 5643 5978
rect 5597 5906 5603 5966
rect 5637 5906 5643 5966
rect 5597 5894 5643 5906
rect 5725 5966 5771 5978
rect 5725 5906 5731 5966
rect 5765 5906 5771 5966
rect 5725 5894 5771 5906
rect 5853 5966 5899 5978
rect 5853 5906 5859 5966
rect 5893 5906 5899 5966
rect 5853 5894 5899 5906
rect 5981 5966 6027 5978
rect 5981 5906 5987 5966
rect 6021 5906 6027 5966
rect 5981 5894 6027 5906
rect 6109 5966 6155 5978
rect 6109 5906 6115 5966
rect 6149 5906 6155 5966
rect 6109 5894 6155 5906
rect 6237 5966 6283 5978
rect 6237 5906 6243 5966
rect 6277 5906 6283 5966
rect 6237 5894 6283 5906
rect 6365 5966 6411 5978
rect 6365 5906 6371 5966
rect 6405 5906 6411 5966
rect 6365 5894 6411 5906
rect 6493 5966 6539 5978
rect 6493 5906 6499 5966
rect 6533 5906 6539 5966
rect 6493 5894 6539 5906
rect 6621 5966 6667 5978
rect 6621 5906 6627 5966
rect 6661 5906 6667 5966
rect 6621 5894 6667 5906
rect 6749 5966 6795 5978
rect 6749 5906 6755 5966
rect 6789 5906 6795 5966
rect 6749 5894 6795 5906
rect 6877 5966 6923 5978
rect 6877 5906 6883 5966
rect 6917 5906 6923 5966
rect 6877 5894 6923 5906
rect 7005 5966 7051 5978
rect 7005 5906 7011 5966
rect 7045 5906 7051 5966
rect 7005 5894 7051 5906
rect 7133 5966 7179 5978
rect 7133 5906 7139 5966
rect 7173 5906 7179 5966
rect 7133 5894 7179 5906
rect 7261 5966 7307 5978
rect 7261 5906 7267 5966
rect 7301 5906 7307 5966
rect 7261 5894 7307 5906
rect 7389 5966 7435 5978
rect 7389 5906 7395 5966
rect 7429 5906 7435 5966
rect 7389 5894 7435 5906
rect 7517 5966 7563 5978
rect 7517 5906 7523 5966
rect 7557 5906 7563 5966
rect 7517 5894 7563 5906
rect 10556 5966 10602 5978
rect 10556 5906 10562 5966
rect 10596 5906 10602 5966
rect 10556 5894 10602 5906
rect 10684 5966 10730 5978
rect 10684 5906 10690 5966
rect 10724 5906 10730 5966
rect 10684 5894 10730 5906
rect 10812 5966 10858 5978
rect 10812 5906 10818 5966
rect 10852 5906 10858 5966
rect 10812 5894 10858 5906
rect 10940 5966 10986 5978
rect 10940 5906 10946 5966
rect 10980 5906 10986 5966
rect 10940 5894 10986 5906
rect 11068 5966 11114 5978
rect 11068 5906 11074 5966
rect 11108 5906 11114 5966
rect 11068 5894 11114 5906
rect 11196 5966 11242 5978
rect 11196 5906 11202 5966
rect 11236 5906 11242 5966
rect 11196 5894 11242 5906
rect 11324 5966 11370 5978
rect 11324 5906 11330 5966
rect 11364 5906 11370 5966
rect 11324 5894 11370 5906
rect 11452 5966 11498 5978
rect 11452 5906 11458 5966
rect 11492 5906 11498 5966
rect 11452 5894 11498 5906
rect 11580 5966 11626 5978
rect 11580 5906 11586 5966
rect 11620 5906 11626 5966
rect 11580 5894 11626 5906
rect 11708 5966 11754 5978
rect 11708 5906 11714 5966
rect 11748 5906 11754 5966
rect 11708 5894 11754 5906
rect 11836 5966 11882 5978
rect 11836 5906 11842 5966
rect 11876 5906 11882 5966
rect 11836 5894 11882 5906
rect 11964 5966 12010 5978
rect 11964 5906 11970 5966
rect 12004 5906 12010 5966
rect 11964 5894 12010 5906
rect 12092 5966 12138 5978
rect 12092 5906 12098 5966
rect 12132 5906 12138 5966
rect 12092 5894 12138 5906
rect 12220 5966 12266 5978
rect 12220 5906 12226 5966
rect 12260 5906 12266 5966
rect 12220 5894 12266 5906
rect 12348 5966 12394 5978
rect 12348 5906 12354 5966
rect 12388 5906 12394 5966
rect 12348 5894 12394 5906
rect 12476 5966 12522 5978
rect 12476 5906 12482 5966
rect 12516 5906 12522 5966
rect 12476 5894 12522 5906
rect 12604 5966 12650 5978
rect 12604 5906 12610 5966
rect 12644 5906 12650 5966
rect 12604 5894 12650 5906
rect 12732 5966 12778 5978
rect 12732 5906 12738 5966
rect 12772 5906 12778 5966
rect 12732 5894 12778 5906
rect 12860 5966 12906 5978
rect 12860 5906 12866 5966
rect 12900 5906 12906 5966
rect 12860 5894 12906 5906
rect 12988 5966 13034 5978
rect 12988 5906 12994 5966
rect 13028 5906 13034 5966
rect 12988 5894 13034 5906
rect 13116 5966 13162 5978
rect 13116 5906 13122 5966
rect 13156 5906 13162 5966
rect 13116 5894 13162 5906
rect 13244 5966 13290 5978
rect 13244 5906 13250 5966
rect 13284 5906 13290 5966
rect 13244 5894 13290 5906
rect 13372 5966 13418 5978
rect 13372 5906 13378 5966
rect 13412 5906 13418 5966
rect 13372 5894 13418 5906
rect 13500 5966 13546 5978
rect 13500 5906 13506 5966
rect 13540 5906 13546 5966
rect 13500 5894 13546 5906
rect 13628 5966 13674 5978
rect 13628 5906 13634 5966
rect 13668 5906 13674 5966
rect 13628 5894 13674 5906
rect 13756 5966 13802 5978
rect 13756 5906 13762 5966
rect 13796 5906 13802 5966
rect 13756 5894 13802 5906
rect 13884 5966 13930 5978
rect 13884 5906 13890 5966
rect 13924 5906 13930 5966
rect 13884 5894 13930 5906
rect 14012 5966 14058 5978
rect 14012 5906 14018 5966
rect 14052 5906 14058 5966
rect 14012 5894 14058 5906
rect 14140 5966 14186 5978
rect 14140 5906 14146 5966
rect 14180 5906 14186 5966
rect 14140 5894 14186 5906
rect 14268 5966 14314 5978
rect 14268 5906 14274 5966
rect 14308 5906 14314 5966
rect 14268 5894 14314 5906
rect 14396 5966 14442 5978
rect 14396 5906 14402 5966
rect 14436 5906 14442 5966
rect 14396 5894 14442 5906
rect 14524 5966 14570 5978
rect 14524 5906 14530 5966
rect 14564 5906 14570 5966
rect 14524 5894 14570 5906
rect 14652 5966 14698 5978
rect 14652 5906 14658 5966
rect 14692 5906 14698 5966
rect 14652 5894 14698 5906
rect 20341 5966 20387 5978
rect 20341 5906 20347 5966
rect 20381 5906 20387 5966
rect 20341 5894 20387 5906
rect 20469 5966 20515 5978
rect 20469 5906 20475 5966
rect 20509 5906 20515 5966
rect 20469 5894 20515 5906
rect 20597 5966 20643 5978
rect 20597 5906 20603 5966
rect 20637 5906 20643 5966
rect 20597 5894 20643 5906
rect 20725 5966 20771 5978
rect 20725 5906 20731 5966
rect 20765 5906 20771 5966
rect 20725 5894 20771 5906
rect 20853 5966 20899 5978
rect 20853 5906 20859 5966
rect 20893 5906 20899 5966
rect 20853 5894 20899 5906
rect 20981 5966 21027 5978
rect 20981 5906 20987 5966
rect 21021 5906 21027 5966
rect 20981 5894 21027 5906
rect 21109 5966 21155 5978
rect 21109 5906 21115 5966
rect 21149 5906 21155 5966
rect 21109 5894 21155 5906
rect 21237 5966 21283 5978
rect 21237 5906 21243 5966
rect 21277 5906 21283 5966
rect 21237 5894 21283 5906
rect 21365 5966 21411 5978
rect 21365 5906 21371 5966
rect 21405 5906 21411 5966
rect 21365 5894 21411 5906
rect 21493 5966 21539 5978
rect 21493 5906 21499 5966
rect 21533 5906 21539 5966
rect 21493 5894 21539 5906
rect 21621 5966 21667 5978
rect 21621 5906 21627 5966
rect 21661 5906 21667 5966
rect 21621 5894 21667 5906
rect 21749 5966 21795 5978
rect 21749 5906 21755 5966
rect 21789 5906 21795 5966
rect 21749 5894 21795 5906
rect 21877 5966 21923 5978
rect 21877 5906 21883 5966
rect 21917 5906 21923 5966
rect 21877 5894 21923 5906
rect 22005 5966 22051 5978
rect 22005 5906 22011 5966
rect 22045 5906 22051 5966
rect 22005 5894 22051 5906
rect 22133 5966 22179 5978
rect 22133 5906 22139 5966
rect 22173 5906 22179 5966
rect 22133 5894 22179 5906
rect 22261 5966 22307 5978
rect 22261 5906 22267 5966
rect 22301 5906 22307 5966
rect 22261 5894 22307 5906
rect 22389 5966 22435 5978
rect 22389 5906 22395 5966
rect 22429 5906 22435 5966
rect 22389 5894 22435 5906
rect 22517 5966 22563 5978
rect 22517 5906 22523 5966
rect 22557 5906 22563 5966
rect 22517 5894 22563 5906
rect 22645 5966 22691 5978
rect 22645 5906 22651 5966
rect 22685 5906 22691 5966
rect 22645 5894 22691 5906
rect 22773 5966 22819 5978
rect 22773 5906 22779 5966
rect 22813 5906 22819 5966
rect 22773 5894 22819 5906
rect 22901 5966 22947 5978
rect 22901 5906 22907 5966
rect 22941 5906 22947 5966
rect 22901 5894 22947 5906
rect 23029 5966 23075 5978
rect 23029 5906 23035 5966
rect 23069 5906 23075 5966
rect 23029 5894 23075 5906
rect 23157 5966 23203 5978
rect 23157 5906 23163 5966
rect 23197 5906 23203 5966
rect 23157 5894 23203 5906
rect 23285 5966 23331 5978
rect 23285 5906 23291 5966
rect 23325 5906 23331 5966
rect 23285 5894 23331 5906
rect 23413 5966 23459 5978
rect 23413 5906 23419 5966
rect 23453 5906 23459 5966
rect 23413 5894 23459 5906
rect 23541 5966 23587 5978
rect 23541 5906 23547 5966
rect 23581 5906 23587 5966
rect 23541 5894 23587 5906
rect 23669 5966 23715 5978
rect 23669 5906 23675 5966
rect 23709 5906 23715 5966
rect 23669 5894 23715 5906
rect 23797 5966 23843 5978
rect 23797 5906 23803 5966
rect 23837 5906 23843 5966
rect 23797 5894 23843 5906
rect 23925 5966 23971 5978
rect 23925 5906 23931 5966
rect 23965 5906 23971 5966
rect 23925 5894 23971 5906
rect 24053 5966 24099 5978
rect 24053 5906 24059 5966
rect 24093 5906 24099 5966
rect 24053 5894 24099 5906
rect 24181 5966 24227 5978
rect 24181 5906 24187 5966
rect 24221 5906 24227 5966
rect 24181 5894 24227 5906
rect 24309 5966 24355 5978
rect 24309 5906 24315 5966
rect 24349 5906 24355 5966
rect 24309 5894 24355 5906
rect 24437 5966 24483 5978
rect 24437 5906 24443 5966
rect 24477 5906 24483 5966
rect 24437 5894 24483 5906
rect 24565 5966 24611 5978
rect 24565 5906 24571 5966
rect 24605 5906 24611 5966
rect 24565 5894 24611 5906
rect 24693 5966 24739 5978
rect 24693 5906 24699 5966
rect 24733 5906 24739 5966
rect 24693 5894 24739 5906
rect 24821 5966 24867 5978
rect 24821 5906 24827 5966
rect 24861 5906 24867 5966
rect 24821 5894 24867 5906
rect 24949 5966 24995 5978
rect 24949 5906 24955 5966
rect 24989 5906 24995 5966
rect 24949 5894 24995 5906
rect 25077 5966 25123 5978
rect 25077 5906 25083 5966
rect 25117 5906 25123 5966
rect 25077 5894 25123 5906
rect 25205 5966 25251 5978
rect 25205 5906 25211 5966
rect 25245 5906 25251 5966
rect 25205 5894 25251 5906
rect 25333 5966 25379 5978
rect 25333 5906 25339 5966
rect 25373 5906 25379 5966
rect 25333 5894 25379 5906
rect 25461 5966 25507 5978
rect 25461 5906 25467 5966
rect 25501 5906 25507 5966
rect 25461 5894 25507 5906
rect 25589 5966 25635 5978
rect 25589 5906 25595 5966
rect 25629 5906 25635 5966
rect 25589 5894 25635 5906
rect 25717 5966 25763 5978
rect 25717 5906 25723 5966
rect 25757 5906 25763 5966
rect 25717 5894 25763 5906
rect 25845 5966 25891 5978
rect 25845 5906 25851 5966
rect 25885 5906 25891 5966
rect 25845 5894 25891 5906
rect 25973 5966 26019 5978
rect 25973 5906 25979 5966
rect 26013 5906 26019 5966
rect 25973 5894 26019 5906
rect 26101 5966 26147 5978
rect 26101 5906 26107 5966
rect 26141 5906 26147 5966
rect 26101 5894 26147 5906
rect 26229 5966 26275 5978
rect 26229 5906 26235 5966
rect 26269 5906 26275 5966
rect 26229 5894 26275 5906
rect 26357 5966 26403 5978
rect 26357 5906 26363 5966
rect 26397 5906 26403 5966
rect 26357 5894 26403 5906
rect 26485 5966 26531 5978
rect 26485 5906 26491 5966
rect 26525 5906 26531 5966
rect 26485 5894 26531 5906
rect 26613 5966 26659 5978
rect 26613 5906 26619 5966
rect 26653 5906 26659 5966
rect 26613 5894 26659 5906
rect 26741 5966 26787 5978
rect 26741 5906 26747 5966
rect 26781 5906 26787 5966
rect 26741 5894 26787 5906
rect 26869 5966 26915 5978
rect 26869 5906 26875 5966
rect 26909 5906 26915 5966
rect 26869 5894 26915 5906
rect 26997 5966 27043 5978
rect 26997 5906 27003 5966
rect 27037 5906 27043 5966
rect 26997 5894 27043 5906
rect 27125 5966 27171 5978
rect 27125 5906 27131 5966
rect 27165 5906 27171 5966
rect 27125 5894 27171 5906
rect 27253 5966 27299 5978
rect 27253 5906 27259 5966
rect 27293 5906 27299 5966
rect 27253 5894 27299 5906
rect 27381 5966 27427 5978
rect 27381 5906 27387 5966
rect 27421 5906 27427 5966
rect 27381 5894 27427 5906
rect 27509 5966 27555 5978
rect 27509 5906 27515 5966
rect 27549 5906 27555 5966
rect 27509 5894 27555 5906
rect 27637 5966 27683 5978
rect 27637 5906 27643 5966
rect 27677 5906 27683 5966
rect 27637 5894 27683 5906
rect 27765 5966 27811 5978
rect 27765 5906 27771 5966
rect 27805 5906 27811 5966
rect 27765 5894 27811 5906
rect 27893 5966 27939 5978
rect 27893 5906 27899 5966
rect 27933 5906 27939 5966
rect 27893 5894 27939 5906
rect 28021 5966 28067 5978
rect 28021 5906 28027 5966
rect 28061 5906 28067 5966
rect 28021 5894 28067 5906
rect 28149 5966 28195 5978
rect 28149 5906 28155 5966
rect 28189 5906 28195 5966
rect 28149 5894 28195 5906
rect 28277 5966 28323 5978
rect 28277 5906 28283 5966
rect 28317 5906 28323 5966
rect 28277 5894 28323 5906
rect 28405 5966 28451 5978
rect 28405 5906 28411 5966
rect 28445 5906 28451 5966
rect 28405 5894 28451 5906
rect 28533 5966 28579 5978
rect 28533 5906 28539 5966
rect 28573 5906 28579 5966
rect 28533 5894 28579 5906
rect -295 5842 -261 5894
rect 482 5842 516 5894
rect 738 5842 772 5894
rect 1391 5842 1425 5894
rect 1647 5842 1681 5894
rect 1903 5842 1937 5894
rect 2924 5842 2958 5894
rect 3180 5842 3214 5894
rect 3436 5842 3470 5894
rect 3692 5842 3726 5894
rect 3948 5842 3982 5894
rect 5475 5842 5509 5894
rect 5731 5842 5765 5894
rect 5987 5842 6021 5894
rect 6243 5842 6277 5894
rect 6499 5842 6533 5894
rect 6755 5842 6789 5894
rect 7011 5842 7045 5894
rect 7267 5842 7301 5894
rect 7523 5842 7557 5894
rect 10562 5842 10596 5894
rect 10818 5842 10852 5894
rect 11074 5842 11108 5894
rect 11330 5842 11364 5894
rect 11586 5842 11620 5894
rect 11842 5842 11876 5894
rect 12098 5842 12132 5894
rect 12354 5842 12388 5894
rect 12610 5842 12644 5894
rect 12866 5842 12900 5894
rect 13122 5842 13156 5894
rect 13378 5842 13412 5894
rect 13634 5842 13668 5894
rect 13890 5842 13924 5894
rect 14146 5842 14180 5894
rect 14402 5842 14436 5894
rect 14658 5842 14692 5894
rect 20347 5842 20381 5894
rect 20603 5842 20637 5894
rect 20859 5842 20893 5894
rect 21115 5842 21149 5894
rect 21371 5842 21405 5894
rect 21627 5842 21661 5894
rect 21883 5842 21917 5894
rect 22139 5842 22173 5894
rect 22395 5842 22429 5894
rect 22651 5842 22685 5894
rect 22907 5842 22941 5894
rect 23163 5842 23197 5894
rect 23419 5842 23453 5894
rect 23675 5842 23709 5894
rect 23931 5842 23965 5894
rect 24187 5842 24221 5894
rect 24443 5842 24477 5894
rect 24699 5842 24733 5894
rect 24955 5842 24989 5894
rect 25211 5842 25245 5894
rect 25467 5842 25501 5894
rect 25723 5842 25757 5894
rect 25979 5842 26013 5894
rect 26235 5842 26269 5894
rect 26491 5842 26525 5894
rect 26747 5842 26781 5894
rect 27003 5842 27037 5894
rect 27259 5842 27293 5894
rect 27515 5842 27549 5894
rect 27771 5842 27805 5894
rect 28027 5842 28061 5894
rect 28283 5842 28317 5894
rect 28539 5842 28573 5894
rect 28824 5843 28888 5849
rect 28824 5842 28830 5843
rect -341 5836 28830 5842
rect -341 5798 -297 5836
rect -259 5798 -169 5836
rect -131 5798 480 5836
rect 518 5798 608 5836
rect 646 5798 736 5836
rect 774 5798 1389 5836
rect 1427 5798 1517 5836
rect 1555 5798 1645 5836
rect 1683 5798 1773 5836
rect 1811 5798 1901 5836
rect 1939 5798 2922 5836
rect 2960 5798 3050 5836
rect 3088 5798 3178 5836
rect 3216 5798 3306 5836
rect 3344 5798 3434 5836
rect 3472 5798 3562 5836
rect 3600 5798 3690 5836
rect 3728 5798 3818 5836
rect 3856 5798 3946 5836
rect 3984 5798 5473 5836
rect 5511 5798 5601 5836
rect 5639 5798 5729 5836
rect 5767 5798 5857 5836
rect 5895 5798 5985 5836
rect 6023 5798 6113 5836
rect 6151 5798 6241 5836
rect 6279 5798 6369 5836
rect 6407 5798 6497 5836
rect 6535 5798 6625 5836
rect 6663 5798 6753 5836
rect 6791 5798 6881 5836
rect 6919 5798 7009 5836
rect 7047 5798 7137 5836
rect 7175 5798 7265 5836
rect 7303 5798 7393 5836
rect 7431 5798 7521 5836
rect 7559 5798 10560 5836
rect 10598 5798 10688 5836
rect 10726 5798 10816 5836
rect 10854 5798 10944 5836
rect 10982 5798 11072 5836
rect 11110 5798 11200 5836
rect 11238 5798 11328 5836
rect 11366 5798 11456 5836
rect 11494 5798 11584 5836
rect 11622 5798 11712 5836
rect 11750 5798 11840 5836
rect 11878 5798 11968 5836
rect 12006 5798 12096 5836
rect 12134 5798 12224 5836
rect 12262 5798 12352 5836
rect 12390 5798 12480 5836
rect 12518 5798 12608 5836
rect 12646 5798 12736 5836
rect 12774 5798 12864 5836
rect 12902 5798 12992 5836
rect 13030 5798 13120 5836
rect 13158 5798 13248 5836
rect 13286 5798 13376 5836
rect 13414 5798 13504 5836
rect 13542 5798 13632 5836
rect 13670 5798 13760 5836
rect 13798 5798 13888 5836
rect 13926 5798 14016 5836
rect 14054 5798 14144 5836
rect 14182 5798 14272 5836
rect 14310 5798 14400 5836
rect 14438 5798 14528 5836
rect 14566 5798 14656 5836
rect 14694 5798 20345 5836
rect 20383 5798 20473 5836
rect 20511 5798 20601 5836
rect 20639 5798 20729 5836
rect 20767 5798 20857 5836
rect 20895 5798 20985 5836
rect 21023 5798 21113 5836
rect 21151 5798 21241 5836
rect 21279 5798 21369 5836
rect 21407 5798 21497 5836
rect 21535 5798 21625 5836
rect 21663 5798 21753 5836
rect 21791 5798 21881 5836
rect 21919 5798 22009 5836
rect 22047 5798 22137 5836
rect 22175 5798 22265 5836
rect 22303 5798 22393 5836
rect 22431 5798 22521 5836
rect 22559 5798 22649 5836
rect 22687 5798 22777 5836
rect 22815 5798 22905 5836
rect 22943 5798 23033 5836
rect 23071 5798 23161 5836
rect 23199 5798 23289 5836
rect 23327 5798 23417 5836
rect 23455 5798 23545 5836
rect 23583 5798 23673 5836
rect 23711 5798 23801 5836
rect 23839 5798 23929 5836
rect 23967 5798 24057 5836
rect 24095 5798 24185 5836
rect 24223 5798 24313 5836
rect 24351 5798 24441 5836
rect 24479 5798 24569 5836
rect 24607 5798 24697 5836
rect 24735 5798 24825 5836
rect 24863 5798 24953 5836
rect 24991 5798 25081 5836
rect 25119 5798 25209 5836
rect 25247 5798 25337 5836
rect 25375 5798 25465 5836
rect 25503 5798 25593 5836
rect 25631 5798 25721 5836
rect 25759 5798 25849 5836
rect 25887 5798 25977 5836
rect 26015 5798 26105 5836
rect 26143 5798 26233 5836
rect 26271 5798 26361 5836
rect 26399 5798 26489 5836
rect 26527 5798 26617 5836
rect 26655 5798 26745 5836
rect 26783 5798 26873 5836
rect 26911 5798 27001 5836
rect 27039 5798 27129 5836
rect 27167 5798 27257 5836
rect 27295 5798 27385 5836
rect 27423 5798 27513 5836
rect 27551 5798 27641 5836
rect 27679 5798 27769 5836
rect 27807 5798 27897 5836
rect 27935 5798 28025 5836
rect 28063 5798 28153 5836
rect 28191 5798 28281 5836
rect 28319 5798 28409 5836
rect 28447 5798 28537 5836
rect 28575 5798 28830 5836
rect -341 5792 28830 5798
rect 28824 5791 28830 5792
rect 28882 5791 28888 5843
rect 28824 5785 28888 5791
rect 29504 5736 29568 5742
rect 29504 5734 29510 5736
rect -363 5728 29510 5734
rect -363 5690 -319 5728
rect -281 5690 -191 5728
rect -153 5690 609 5728
rect 647 5690 737 5728
rect 775 5690 865 5728
rect 903 5690 1873 5728
rect 1911 5690 2001 5728
rect 2039 5690 2129 5728
rect 2167 5690 2257 5728
rect 2295 5690 2385 5728
rect 2423 5690 3492 5728
rect 3530 5690 3620 5728
rect 3658 5690 3748 5728
rect 3786 5690 3876 5728
rect 3914 5690 4004 5728
rect 4042 5690 4132 5728
rect 4170 5690 4260 5728
rect 4298 5690 4388 5728
rect 4426 5690 4516 5728
rect 4554 5690 8057 5728
rect 8095 5690 8185 5728
rect 8223 5690 8313 5728
rect 8351 5690 8441 5728
rect 8479 5690 8569 5728
rect 8607 5690 8697 5728
rect 8735 5690 8825 5728
rect 8863 5690 8953 5728
rect 8991 5690 9081 5728
rect 9119 5690 9209 5728
rect 9247 5690 9337 5728
rect 9375 5690 9465 5728
rect 9503 5690 9593 5728
rect 9631 5690 9721 5728
rect 9759 5690 9849 5728
rect 9887 5690 9977 5728
rect 10015 5690 10105 5728
rect 10143 5690 15215 5728
rect 15253 5690 15343 5728
rect 15381 5690 15471 5728
rect 15509 5690 15599 5728
rect 15637 5690 15727 5728
rect 15765 5690 15855 5728
rect 15893 5690 15983 5728
rect 16021 5690 16111 5728
rect 16149 5690 16239 5728
rect 16277 5690 16367 5728
rect 16405 5690 16495 5728
rect 16533 5690 16623 5728
rect 16661 5690 16751 5728
rect 16789 5690 16879 5728
rect 16917 5690 17007 5728
rect 17045 5690 17135 5728
rect 17173 5690 17263 5728
rect 17301 5690 17391 5728
rect 17429 5690 17519 5728
rect 17557 5690 17647 5728
rect 17685 5690 17775 5728
rect 17813 5690 17903 5728
rect 17941 5690 18031 5728
rect 18069 5690 18159 5728
rect 18197 5690 18287 5728
rect 18325 5690 18415 5728
rect 18453 5690 18543 5728
rect 18581 5690 18671 5728
rect 18709 5690 18799 5728
rect 18837 5690 18927 5728
rect 18965 5690 19055 5728
rect 19093 5690 19183 5728
rect 19221 5690 19311 5728
rect 19349 5690 20269 5728
rect 20307 5690 20397 5728
rect 20435 5690 20525 5728
rect 20563 5690 20653 5728
rect 20691 5690 20781 5728
rect 20819 5690 20909 5728
rect 20947 5690 21037 5728
rect 21075 5690 21165 5728
rect 21203 5690 21293 5728
rect 21331 5690 21421 5728
rect 21459 5690 21549 5728
rect 21587 5690 21677 5728
rect 21715 5690 21805 5728
rect 21843 5690 21933 5728
rect 21971 5690 22061 5728
rect 22099 5690 22189 5728
rect 22227 5690 22317 5728
rect 22355 5690 22445 5728
rect 22483 5690 22573 5728
rect 22611 5690 22701 5728
rect 22739 5690 22829 5728
rect 22867 5690 22957 5728
rect 22995 5690 23085 5728
rect 23123 5690 23213 5728
rect 23251 5690 23341 5728
rect 23379 5690 23469 5728
rect 23507 5690 23597 5728
rect 23635 5690 23725 5728
rect 23763 5690 23853 5728
rect 23891 5690 23981 5728
rect 24019 5690 24109 5728
rect 24147 5690 24237 5728
rect 24275 5690 24365 5728
rect 24403 5690 24493 5728
rect 24531 5690 24621 5728
rect 24659 5690 24749 5728
rect 24787 5690 24877 5728
rect 24915 5690 25005 5728
rect 25043 5690 25133 5728
rect 25171 5690 25261 5728
rect 25299 5690 25389 5728
rect 25427 5690 25517 5728
rect 25555 5690 25645 5728
rect 25683 5690 25773 5728
rect 25811 5690 25901 5728
rect 25939 5690 26029 5728
rect 26067 5690 26157 5728
rect 26195 5690 26285 5728
rect 26323 5690 26413 5728
rect 26451 5690 26541 5728
rect 26579 5690 26669 5728
rect 26707 5690 26797 5728
rect 26835 5690 26925 5728
rect 26963 5690 27053 5728
rect 27091 5690 27181 5728
rect 27219 5690 27309 5728
rect 27347 5690 27437 5728
rect 27475 5690 27565 5728
rect 27603 5690 27693 5728
rect 27731 5690 27821 5728
rect 27859 5690 27949 5728
rect 27987 5690 28077 5728
rect 28115 5690 28205 5728
rect 28243 5690 28333 5728
rect 28371 5690 28461 5728
rect 28499 5690 29510 5728
rect -363 5684 29510 5690
rect 29562 5684 29568 5736
rect 29504 5678 29568 5684
rect -363 5649 28783 5655
rect -363 5623 28725 5649
rect -317 5590 -283 5623
rect 611 5590 645 5623
rect 867 5590 901 5623
rect 1875 5590 1909 5623
rect 2131 5590 2165 5623
rect 2387 5590 2421 5623
rect 3494 5590 3528 5623
rect 3750 5590 3784 5623
rect 4006 5590 4040 5623
rect 4262 5590 4296 5623
rect 4518 5590 4552 5623
rect 8059 5590 8093 5623
rect 8315 5590 8349 5623
rect 8571 5590 8605 5623
rect 8827 5590 8861 5623
rect 9083 5590 9117 5623
rect 9339 5590 9373 5623
rect 9595 5590 9629 5623
rect 9851 5590 9885 5623
rect 10107 5590 10141 5623
rect 15217 5590 15251 5623
rect 15473 5590 15507 5623
rect 15729 5590 15763 5623
rect 15985 5590 16019 5623
rect 16241 5590 16275 5623
rect 16497 5590 16531 5623
rect 16753 5590 16787 5623
rect 17009 5590 17043 5623
rect 17265 5590 17299 5623
rect 17521 5590 17555 5623
rect 17777 5590 17811 5623
rect 18033 5590 18067 5623
rect 18289 5590 18323 5623
rect 18545 5590 18579 5623
rect 18801 5590 18835 5623
rect 19057 5590 19091 5623
rect 19313 5590 19347 5623
rect 20271 5590 20305 5623
rect 20527 5590 20561 5623
rect 20783 5590 20817 5623
rect 21039 5590 21073 5623
rect 21295 5590 21329 5623
rect 21551 5590 21585 5623
rect 21807 5590 21841 5623
rect 22063 5590 22097 5623
rect 22319 5590 22353 5623
rect 22575 5590 22609 5623
rect 22831 5590 22865 5623
rect 23087 5590 23121 5623
rect 23343 5590 23377 5623
rect 23599 5590 23633 5623
rect 23855 5590 23889 5623
rect 24111 5590 24145 5623
rect 24367 5590 24401 5623
rect 24623 5590 24657 5623
rect 24879 5590 24913 5623
rect 25135 5590 25169 5623
rect 25391 5590 25425 5623
rect 25647 5590 25681 5623
rect 25903 5590 25937 5623
rect 26159 5590 26193 5623
rect 26415 5590 26449 5623
rect 26671 5590 26705 5623
rect 26927 5590 26961 5623
rect 27183 5590 27217 5623
rect 27439 5590 27473 5623
rect 27695 5590 27729 5623
rect 27951 5590 27985 5623
rect 28207 5590 28241 5623
rect 28463 5590 28497 5623
rect 28719 5597 28725 5623
rect 28777 5597 28783 5649
rect 28719 5591 28783 5597
rect -323 5578 -277 5590
rect -323 5434 -317 5578
rect -283 5434 -277 5578
rect -323 5422 -277 5434
rect -195 5578 -149 5590
rect -195 5434 -189 5578
rect -155 5434 -149 5578
rect -195 5422 -149 5434
rect 605 5578 651 5590
rect 605 5434 611 5578
rect 645 5434 651 5578
rect 605 5422 651 5434
rect 733 5578 779 5590
rect 733 5434 739 5578
rect 773 5434 779 5578
rect 733 5422 779 5434
rect 861 5578 907 5590
rect 861 5434 867 5578
rect 901 5434 907 5578
rect 861 5422 907 5434
rect 1869 5578 1915 5590
rect 1869 5434 1875 5578
rect 1909 5434 1915 5578
rect 1869 5422 1915 5434
rect 1997 5578 2043 5590
rect 1997 5434 2003 5578
rect 2037 5434 2043 5578
rect 1997 5422 2043 5434
rect 2125 5578 2171 5590
rect 2125 5434 2131 5578
rect 2165 5434 2171 5578
rect 2125 5422 2171 5434
rect 2253 5578 2299 5590
rect 2253 5434 2259 5578
rect 2293 5434 2299 5578
rect 2253 5422 2299 5434
rect 2381 5578 2427 5590
rect 2381 5434 2387 5578
rect 2421 5434 2427 5578
rect 2381 5422 2427 5434
rect 3488 5578 3534 5590
rect 3488 5434 3494 5578
rect 3528 5434 3534 5578
rect 3488 5422 3534 5434
rect 3616 5578 3662 5590
rect 3616 5434 3622 5578
rect 3656 5434 3662 5578
rect 3616 5422 3662 5434
rect 3744 5578 3790 5590
rect 3744 5434 3750 5578
rect 3784 5434 3790 5578
rect 3744 5422 3790 5434
rect 3872 5578 3918 5590
rect 3872 5434 3878 5578
rect 3912 5434 3918 5578
rect 3872 5422 3918 5434
rect 4000 5578 4046 5590
rect 4000 5434 4006 5578
rect 4040 5434 4046 5578
rect 4000 5422 4046 5434
rect 4128 5578 4174 5590
rect 4128 5434 4134 5578
rect 4168 5434 4174 5578
rect 4128 5422 4174 5434
rect 4256 5578 4302 5590
rect 4256 5434 4262 5578
rect 4296 5434 4302 5578
rect 4256 5422 4302 5434
rect 4384 5578 4430 5590
rect 4384 5434 4390 5578
rect 4424 5434 4430 5578
rect 4384 5422 4430 5434
rect 4512 5578 4558 5590
rect 4512 5434 4518 5578
rect 4552 5434 4558 5578
rect 4512 5422 4558 5434
rect 8053 5578 8099 5590
rect 8053 5434 8059 5578
rect 8093 5434 8099 5578
rect 8053 5422 8099 5434
rect 8181 5578 8227 5590
rect 8181 5434 8187 5578
rect 8221 5434 8227 5578
rect 8181 5422 8227 5434
rect 8309 5578 8355 5590
rect 8309 5434 8315 5578
rect 8349 5434 8355 5578
rect 8309 5422 8355 5434
rect 8437 5578 8483 5590
rect 8437 5434 8443 5578
rect 8477 5434 8483 5578
rect 8437 5422 8483 5434
rect 8565 5578 8611 5590
rect 8565 5434 8571 5578
rect 8605 5434 8611 5578
rect 8565 5422 8611 5434
rect 8693 5578 8739 5590
rect 8693 5434 8699 5578
rect 8733 5434 8739 5578
rect 8693 5422 8739 5434
rect 8821 5578 8867 5590
rect 8821 5434 8827 5578
rect 8861 5434 8867 5578
rect 8821 5422 8867 5434
rect 8949 5578 8995 5590
rect 8949 5434 8955 5578
rect 8989 5434 8995 5578
rect 8949 5422 8995 5434
rect 9077 5578 9123 5590
rect 9077 5434 9083 5578
rect 9117 5434 9123 5578
rect 9077 5422 9123 5434
rect 9205 5578 9251 5590
rect 9205 5434 9211 5578
rect 9245 5434 9251 5578
rect 9205 5422 9251 5434
rect 9333 5578 9379 5590
rect 9333 5434 9339 5578
rect 9373 5434 9379 5578
rect 9333 5422 9379 5434
rect 9461 5578 9507 5590
rect 9461 5434 9467 5578
rect 9501 5434 9507 5578
rect 9461 5422 9507 5434
rect 9589 5578 9635 5590
rect 9589 5434 9595 5578
rect 9629 5434 9635 5578
rect 9589 5422 9635 5434
rect 9717 5578 9763 5590
rect 9717 5434 9723 5578
rect 9757 5434 9763 5578
rect 9717 5422 9763 5434
rect 9845 5578 9891 5590
rect 9845 5434 9851 5578
rect 9885 5434 9891 5578
rect 9845 5422 9891 5434
rect 9973 5578 10019 5590
rect 9973 5434 9979 5578
rect 10013 5434 10019 5578
rect 9973 5422 10019 5434
rect 10101 5578 10147 5590
rect 10101 5434 10107 5578
rect 10141 5434 10147 5578
rect 10101 5422 10147 5434
rect 15211 5578 15257 5590
rect 15211 5434 15217 5578
rect 15251 5434 15257 5578
rect 15211 5422 15257 5434
rect 15339 5578 15385 5590
rect 15339 5434 15345 5578
rect 15379 5434 15385 5578
rect 15339 5422 15385 5434
rect 15467 5578 15513 5590
rect 15467 5434 15473 5578
rect 15507 5434 15513 5578
rect 15467 5422 15513 5434
rect 15595 5578 15641 5590
rect 15595 5434 15601 5578
rect 15635 5434 15641 5578
rect 15595 5422 15641 5434
rect 15723 5578 15769 5590
rect 15723 5434 15729 5578
rect 15763 5434 15769 5578
rect 15723 5422 15769 5434
rect 15851 5578 15897 5590
rect 15851 5434 15857 5578
rect 15891 5434 15897 5578
rect 15851 5422 15897 5434
rect 15979 5578 16025 5590
rect 15979 5434 15985 5578
rect 16019 5434 16025 5578
rect 15979 5422 16025 5434
rect 16107 5578 16153 5590
rect 16107 5434 16113 5578
rect 16147 5434 16153 5578
rect 16107 5422 16153 5434
rect 16235 5578 16281 5590
rect 16235 5434 16241 5578
rect 16275 5434 16281 5578
rect 16235 5422 16281 5434
rect 16363 5578 16409 5590
rect 16363 5434 16369 5578
rect 16403 5434 16409 5578
rect 16363 5422 16409 5434
rect 16491 5578 16537 5590
rect 16491 5434 16497 5578
rect 16531 5434 16537 5578
rect 16491 5422 16537 5434
rect 16619 5578 16665 5590
rect 16619 5434 16625 5578
rect 16659 5434 16665 5578
rect 16619 5422 16665 5434
rect 16747 5578 16793 5590
rect 16747 5434 16753 5578
rect 16787 5434 16793 5578
rect 16747 5422 16793 5434
rect 16875 5578 16921 5590
rect 16875 5434 16881 5578
rect 16915 5434 16921 5578
rect 16875 5422 16921 5434
rect 17003 5578 17049 5590
rect 17003 5434 17009 5578
rect 17043 5434 17049 5578
rect 17003 5422 17049 5434
rect 17131 5578 17177 5590
rect 17131 5434 17137 5578
rect 17171 5434 17177 5578
rect 17131 5422 17177 5434
rect 17259 5578 17305 5590
rect 17259 5434 17265 5578
rect 17299 5434 17305 5578
rect 17259 5422 17305 5434
rect 17387 5578 17433 5590
rect 17387 5434 17393 5578
rect 17427 5434 17433 5578
rect 17387 5422 17433 5434
rect 17515 5578 17561 5590
rect 17515 5434 17521 5578
rect 17555 5434 17561 5578
rect 17515 5422 17561 5434
rect 17643 5578 17689 5590
rect 17643 5434 17649 5578
rect 17683 5434 17689 5578
rect 17643 5422 17689 5434
rect 17771 5578 17817 5590
rect 17771 5434 17777 5578
rect 17811 5434 17817 5578
rect 17771 5422 17817 5434
rect 17899 5578 17945 5590
rect 17899 5434 17905 5578
rect 17939 5434 17945 5578
rect 17899 5422 17945 5434
rect 18027 5578 18073 5590
rect 18027 5434 18033 5578
rect 18067 5434 18073 5578
rect 18027 5422 18073 5434
rect 18155 5578 18201 5590
rect 18155 5434 18161 5578
rect 18195 5434 18201 5578
rect 18155 5422 18201 5434
rect 18283 5578 18329 5590
rect 18283 5434 18289 5578
rect 18323 5434 18329 5578
rect 18283 5422 18329 5434
rect 18411 5578 18457 5590
rect 18411 5434 18417 5578
rect 18451 5434 18457 5578
rect 18411 5422 18457 5434
rect 18539 5578 18585 5590
rect 18539 5434 18545 5578
rect 18579 5434 18585 5578
rect 18539 5422 18585 5434
rect 18667 5578 18713 5590
rect 18667 5434 18673 5578
rect 18707 5434 18713 5578
rect 18667 5422 18713 5434
rect 18795 5578 18841 5590
rect 18795 5434 18801 5578
rect 18835 5434 18841 5578
rect 18795 5422 18841 5434
rect 18923 5578 18969 5590
rect 18923 5434 18929 5578
rect 18963 5434 18969 5578
rect 18923 5422 18969 5434
rect 19051 5578 19097 5590
rect 19051 5434 19057 5578
rect 19091 5434 19097 5578
rect 19051 5422 19097 5434
rect 19179 5578 19225 5590
rect 19179 5434 19185 5578
rect 19219 5434 19225 5578
rect 19179 5422 19225 5434
rect 19307 5578 19353 5590
rect 19307 5434 19313 5578
rect 19347 5434 19353 5578
rect 19307 5422 19353 5434
rect 20265 5578 20311 5590
rect 20265 5434 20271 5578
rect 20305 5434 20311 5578
rect 20265 5422 20311 5434
rect 20393 5578 20439 5590
rect 20393 5434 20399 5578
rect 20433 5434 20439 5578
rect 20393 5422 20439 5434
rect 20521 5578 20567 5590
rect 20521 5434 20527 5578
rect 20561 5434 20567 5578
rect 20521 5422 20567 5434
rect 20649 5578 20695 5590
rect 20649 5434 20655 5578
rect 20689 5434 20695 5578
rect 20649 5422 20695 5434
rect 20777 5578 20823 5590
rect 20777 5434 20783 5578
rect 20817 5434 20823 5578
rect 20777 5422 20823 5434
rect 20905 5578 20951 5590
rect 20905 5434 20911 5578
rect 20945 5434 20951 5578
rect 20905 5422 20951 5434
rect 21033 5578 21079 5590
rect 21033 5434 21039 5578
rect 21073 5434 21079 5578
rect 21033 5422 21079 5434
rect 21161 5578 21207 5590
rect 21161 5434 21167 5578
rect 21201 5434 21207 5578
rect 21161 5422 21207 5434
rect 21289 5578 21335 5590
rect 21289 5434 21295 5578
rect 21329 5434 21335 5578
rect 21289 5422 21335 5434
rect 21417 5578 21463 5590
rect 21417 5434 21423 5578
rect 21457 5434 21463 5578
rect 21417 5422 21463 5434
rect 21545 5578 21591 5590
rect 21545 5434 21551 5578
rect 21585 5434 21591 5578
rect 21545 5422 21591 5434
rect 21673 5578 21719 5590
rect 21673 5434 21679 5578
rect 21713 5434 21719 5578
rect 21673 5422 21719 5434
rect 21801 5578 21847 5590
rect 21801 5434 21807 5578
rect 21841 5434 21847 5578
rect 21801 5422 21847 5434
rect 21929 5578 21975 5590
rect 21929 5434 21935 5578
rect 21969 5434 21975 5578
rect 21929 5422 21975 5434
rect 22057 5578 22103 5590
rect 22057 5434 22063 5578
rect 22097 5434 22103 5578
rect 22057 5422 22103 5434
rect 22185 5578 22231 5590
rect 22185 5434 22191 5578
rect 22225 5434 22231 5578
rect 22185 5422 22231 5434
rect 22313 5578 22359 5590
rect 22313 5434 22319 5578
rect 22353 5434 22359 5578
rect 22313 5422 22359 5434
rect 22441 5578 22487 5590
rect 22441 5434 22447 5578
rect 22481 5434 22487 5578
rect 22441 5422 22487 5434
rect 22569 5578 22615 5590
rect 22569 5434 22575 5578
rect 22609 5434 22615 5578
rect 22569 5422 22615 5434
rect 22697 5578 22743 5590
rect 22697 5434 22703 5578
rect 22737 5434 22743 5578
rect 22697 5422 22743 5434
rect 22825 5578 22871 5590
rect 22825 5434 22831 5578
rect 22865 5434 22871 5578
rect 22825 5422 22871 5434
rect 22953 5578 22999 5590
rect 22953 5434 22959 5578
rect 22993 5434 22999 5578
rect 22953 5422 22999 5434
rect 23081 5578 23127 5590
rect 23081 5434 23087 5578
rect 23121 5434 23127 5578
rect 23081 5422 23127 5434
rect 23209 5578 23255 5590
rect 23209 5434 23215 5578
rect 23249 5434 23255 5578
rect 23209 5422 23255 5434
rect 23337 5578 23383 5590
rect 23337 5434 23343 5578
rect 23377 5434 23383 5578
rect 23337 5422 23383 5434
rect 23465 5578 23511 5590
rect 23465 5434 23471 5578
rect 23505 5434 23511 5578
rect 23465 5422 23511 5434
rect 23593 5578 23639 5590
rect 23593 5434 23599 5578
rect 23633 5434 23639 5578
rect 23593 5422 23639 5434
rect 23721 5578 23767 5590
rect 23721 5434 23727 5578
rect 23761 5434 23767 5578
rect 23721 5422 23767 5434
rect 23849 5578 23895 5590
rect 23849 5434 23855 5578
rect 23889 5434 23895 5578
rect 23849 5422 23895 5434
rect 23977 5578 24023 5590
rect 23977 5434 23983 5578
rect 24017 5434 24023 5578
rect 23977 5422 24023 5434
rect 24105 5578 24151 5590
rect 24105 5434 24111 5578
rect 24145 5434 24151 5578
rect 24105 5422 24151 5434
rect 24233 5578 24279 5590
rect 24233 5434 24239 5578
rect 24273 5434 24279 5578
rect 24233 5422 24279 5434
rect 24361 5578 24407 5590
rect 24361 5434 24367 5578
rect 24401 5434 24407 5578
rect 24361 5422 24407 5434
rect 24489 5578 24535 5590
rect 24489 5434 24495 5578
rect 24529 5434 24535 5578
rect 24489 5422 24535 5434
rect 24617 5578 24663 5590
rect 24617 5434 24623 5578
rect 24657 5434 24663 5578
rect 24617 5422 24663 5434
rect 24745 5578 24791 5590
rect 24745 5434 24751 5578
rect 24785 5434 24791 5578
rect 24745 5422 24791 5434
rect 24873 5578 24919 5590
rect 24873 5434 24879 5578
rect 24913 5434 24919 5578
rect 24873 5422 24919 5434
rect 25001 5578 25047 5590
rect 25001 5434 25007 5578
rect 25041 5434 25047 5578
rect 25001 5422 25047 5434
rect 25129 5578 25175 5590
rect 25129 5434 25135 5578
rect 25169 5434 25175 5578
rect 25129 5422 25175 5434
rect 25257 5578 25303 5590
rect 25257 5434 25263 5578
rect 25297 5434 25303 5578
rect 25257 5422 25303 5434
rect 25385 5578 25431 5590
rect 25385 5434 25391 5578
rect 25425 5434 25431 5578
rect 25385 5422 25431 5434
rect 25513 5578 25559 5590
rect 25513 5434 25519 5578
rect 25553 5434 25559 5578
rect 25513 5422 25559 5434
rect 25641 5578 25687 5590
rect 25641 5434 25647 5578
rect 25681 5434 25687 5578
rect 25641 5422 25687 5434
rect 25769 5578 25815 5590
rect 25769 5434 25775 5578
rect 25809 5434 25815 5578
rect 25769 5422 25815 5434
rect 25897 5578 25943 5590
rect 25897 5434 25903 5578
rect 25937 5434 25943 5578
rect 25897 5422 25943 5434
rect 26025 5578 26071 5590
rect 26025 5434 26031 5578
rect 26065 5434 26071 5578
rect 26025 5422 26071 5434
rect 26153 5578 26199 5590
rect 26153 5434 26159 5578
rect 26193 5434 26199 5578
rect 26153 5422 26199 5434
rect 26281 5578 26327 5590
rect 26281 5434 26287 5578
rect 26321 5434 26327 5578
rect 26281 5422 26327 5434
rect 26409 5578 26455 5590
rect 26409 5434 26415 5578
rect 26449 5434 26455 5578
rect 26409 5422 26455 5434
rect 26537 5578 26583 5590
rect 26537 5434 26543 5578
rect 26577 5434 26583 5578
rect 26537 5422 26583 5434
rect 26665 5578 26711 5590
rect 26665 5434 26671 5578
rect 26705 5434 26711 5578
rect 26665 5422 26711 5434
rect 26793 5578 26839 5590
rect 26793 5434 26799 5578
rect 26833 5434 26839 5578
rect 26793 5422 26839 5434
rect 26921 5578 26967 5590
rect 26921 5434 26927 5578
rect 26961 5434 26967 5578
rect 26921 5422 26967 5434
rect 27049 5578 27095 5590
rect 27049 5434 27055 5578
rect 27089 5434 27095 5578
rect 27049 5422 27095 5434
rect 27177 5578 27223 5590
rect 27177 5434 27183 5578
rect 27217 5434 27223 5578
rect 27177 5422 27223 5434
rect 27305 5578 27351 5590
rect 27305 5434 27311 5578
rect 27345 5434 27351 5578
rect 27305 5422 27351 5434
rect 27433 5578 27479 5590
rect 27433 5434 27439 5578
rect 27473 5434 27479 5578
rect 27433 5422 27479 5434
rect 27561 5578 27607 5590
rect 27561 5434 27567 5578
rect 27601 5434 27607 5578
rect 27561 5422 27607 5434
rect 27689 5578 27735 5590
rect 27689 5434 27695 5578
rect 27729 5434 27735 5578
rect 27689 5422 27735 5434
rect 27817 5578 27863 5590
rect 27817 5434 27823 5578
rect 27857 5434 27863 5578
rect 27817 5422 27863 5434
rect 27945 5578 27991 5590
rect 27945 5434 27951 5578
rect 27985 5434 27991 5578
rect 27945 5422 27991 5434
rect 28073 5578 28119 5590
rect 28073 5434 28079 5578
rect 28113 5434 28119 5578
rect 28073 5422 28119 5434
rect 28201 5578 28247 5590
rect 28201 5434 28207 5578
rect 28241 5434 28247 5578
rect 28201 5422 28247 5434
rect 28329 5578 28375 5590
rect 28329 5434 28335 5578
rect 28369 5434 28375 5578
rect 28329 5422 28375 5434
rect 28457 5578 28503 5590
rect 28457 5434 28463 5578
rect 28497 5434 28503 5578
rect 28457 5422 28503 5434
rect -189 5356 -155 5422
rect 739 5394 773 5422
rect 962 5401 1026 5407
rect 962 5394 968 5401
rect -95 5363 -31 5369
rect -95 5356 -89 5363
rect -189 5322 -89 5356
rect -189 5290 -155 5322
rect -95 5311 -89 5322
rect -37 5311 -31 5363
rect -95 5305 -31 5311
rect 739 5358 968 5394
rect 739 5290 773 5358
rect 962 5349 968 5358
rect 1020 5349 1026 5401
rect 962 5343 1026 5349
rect 2003 5348 2037 5422
rect 2259 5354 2293 5422
rect 2480 5364 2544 5370
rect 2480 5354 2486 5364
rect 2259 5348 2486 5354
rect 2003 5323 2486 5348
rect 2003 5319 2293 5323
rect 2003 5290 2037 5319
rect 2259 5290 2293 5319
rect 2480 5312 2486 5323
rect 2538 5312 2544 5364
rect 2480 5306 2544 5312
rect 3622 5348 3656 5422
rect 3878 5348 3912 5422
rect 4134 5348 4168 5422
rect 4390 5348 4424 5422
rect 4620 5359 4684 5365
rect 4620 5348 4626 5359
rect 3622 5319 4626 5348
rect 3622 5290 3656 5319
rect 3878 5290 3912 5319
rect 4134 5290 4168 5319
rect 4390 5290 4424 5319
rect 4620 5307 4626 5319
rect 4678 5307 4684 5359
rect 4620 5301 4684 5307
rect 8187 5348 8221 5422
rect 8443 5348 8477 5422
rect 8699 5348 8733 5422
rect 8955 5348 8989 5422
rect 9211 5348 9245 5422
rect 9467 5348 9501 5422
rect 9723 5348 9757 5422
rect 9979 5353 10013 5422
rect 10200 5362 10264 5368
rect 10200 5353 10206 5362
rect 9979 5348 10206 5353
rect 8187 5324 10206 5348
rect 8187 5319 10013 5324
rect 8187 5290 8221 5319
rect 8443 5290 8477 5319
rect 8699 5290 8733 5319
rect 8955 5290 8989 5319
rect 9211 5290 9245 5319
rect 9467 5290 9501 5319
rect 9723 5290 9757 5319
rect 9979 5290 10013 5319
rect 10200 5310 10206 5324
rect 10258 5310 10264 5362
rect 10200 5304 10264 5310
rect 15345 5348 15379 5422
rect 15601 5348 15635 5422
rect 15857 5348 15891 5422
rect 16113 5348 16147 5422
rect 16369 5348 16403 5422
rect 16625 5348 16659 5422
rect 16881 5348 16915 5422
rect 17137 5348 17171 5422
rect 17393 5348 17427 5422
rect 17649 5348 17683 5422
rect 17905 5348 17939 5422
rect 18161 5348 18195 5422
rect 18417 5348 18451 5422
rect 18673 5348 18707 5422
rect 18929 5348 18963 5422
rect 19185 5348 19219 5422
rect 15345 5347 19219 5348
rect 19416 5358 19480 5364
rect 19416 5347 19422 5358
rect 15345 5319 19422 5347
rect 15345 5290 15379 5319
rect 15601 5290 15635 5319
rect 15857 5290 15891 5319
rect 16113 5290 16147 5319
rect 16369 5290 16403 5319
rect 16625 5290 16659 5319
rect 16881 5290 16915 5319
rect 17137 5290 17171 5319
rect 17393 5290 17427 5319
rect 17649 5290 17683 5319
rect 17905 5290 17939 5319
rect 18161 5290 18195 5319
rect 18417 5290 18451 5319
rect 18673 5290 18707 5319
rect 18929 5290 18963 5319
rect 19185 5318 19422 5319
rect 19185 5290 19219 5318
rect 19416 5306 19422 5318
rect 19474 5306 19480 5358
rect 19416 5300 19480 5306
rect 20149 5358 20213 5364
rect 20149 5306 20155 5358
rect 20207 5348 20213 5358
rect 20399 5348 20433 5422
rect 20655 5348 20689 5422
rect 20911 5348 20945 5422
rect 21167 5348 21201 5422
rect 21423 5348 21457 5422
rect 21679 5348 21713 5422
rect 21935 5348 21969 5422
rect 22191 5348 22225 5422
rect 22447 5348 22481 5422
rect 22703 5348 22737 5422
rect 22959 5348 22993 5422
rect 23215 5348 23249 5422
rect 23471 5348 23505 5422
rect 23727 5348 23761 5422
rect 23983 5348 24017 5422
rect 24239 5348 24273 5422
rect 24495 5348 24529 5422
rect 24751 5348 24785 5422
rect 25007 5348 25041 5422
rect 25263 5348 25297 5422
rect 25519 5348 25553 5422
rect 25775 5348 25809 5422
rect 26031 5348 26065 5422
rect 26287 5348 26321 5422
rect 26543 5348 26577 5422
rect 26799 5348 26833 5422
rect 27055 5348 27089 5422
rect 27311 5348 27345 5422
rect 27567 5348 27601 5422
rect 27823 5348 27857 5422
rect 28079 5348 28113 5422
rect 28335 5348 28369 5422
rect 20207 5319 28369 5348
rect 20207 5306 20213 5319
rect 20149 5300 20213 5306
rect 20399 5290 20433 5319
rect 20655 5290 20689 5319
rect 20911 5290 20945 5319
rect 21167 5290 21201 5319
rect 21423 5290 21457 5319
rect 21679 5290 21713 5319
rect 21935 5290 21969 5319
rect 22191 5290 22225 5319
rect 22447 5290 22481 5319
rect 22703 5290 22737 5319
rect 22959 5290 22993 5319
rect 23215 5290 23249 5319
rect 23471 5290 23505 5319
rect 23727 5290 23761 5319
rect 23983 5290 24017 5319
rect 24239 5290 24273 5319
rect 24495 5290 24529 5319
rect 24751 5290 24785 5319
rect 25007 5290 25041 5319
rect 25263 5290 25297 5319
rect 25519 5290 25553 5319
rect 25775 5290 25809 5319
rect 26031 5290 26065 5319
rect 26287 5290 26321 5319
rect 26543 5290 26577 5319
rect 26799 5290 26833 5319
rect 27055 5290 27089 5319
rect 27311 5290 27345 5319
rect 27567 5290 27601 5319
rect 27823 5290 27857 5319
rect 28079 5290 28113 5319
rect 28335 5290 28369 5319
rect -323 5278 -277 5290
rect -323 5218 -317 5278
rect -283 5218 -277 5278
rect -323 5206 -277 5218
rect -195 5278 -149 5290
rect -195 5218 -189 5278
rect -155 5218 -149 5278
rect -195 5206 -149 5218
rect 605 5278 651 5290
rect 605 5218 611 5278
rect 645 5218 651 5278
rect 605 5206 651 5218
rect 733 5278 779 5290
rect 733 5218 739 5278
rect 773 5218 779 5278
rect 733 5206 779 5218
rect 861 5278 907 5290
rect 861 5218 867 5278
rect 901 5218 907 5278
rect 861 5206 907 5218
rect 1869 5278 1915 5290
rect 1869 5218 1875 5278
rect 1909 5218 1915 5278
rect 1869 5206 1915 5218
rect 1997 5278 2043 5290
rect 1997 5218 2003 5278
rect 2037 5218 2043 5278
rect 1997 5206 2043 5218
rect 2125 5278 2171 5290
rect 2125 5218 2131 5278
rect 2165 5218 2171 5278
rect 2125 5206 2171 5218
rect 2253 5278 2299 5290
rect 2253 5218 2259 5278
rect 2293 5218 2299 5278
rect 2253 5206 2299 5218
rect 2381 5278 2427 5290
rect 2381 5218 2387 5278
rect 2421 5218 2427 5278
rect 2381 5206 2427 5218
rect 3488 5278 3534 5290
rect 3488 5218 3494 5278
rect 3528 5218 3534 5278
rect 3488 5206 3534 5218
rect 3616 5278 3662 5290
rect 3616 5218 3622 5278
rect 3656 5218 3662 5278
rect 3616 5206 3662 5218
rect 3744 5278 3790 5290
rect 3744 5218 3750 5278
rect 3784 5218 3790 5278
rect 3744 5206 3790 5218
rect 3872 5278 3918 5290
rect 3872 5218 3878 5278
rect 3912 5218 3918 5278
rect 3872 5206 3918 5218
rect 4000 5278 4046 5290
rect 4000 5218 4006 5278
rect 4040 5218 4046 5278
rect 4000 5206 4046 5218
rect 4128 5278 4174 5290
rect 4128 5218 4134 5278
rect 4168 5218 4174 5278
rect 4128 5206 4174 5218
rect 4256 5278 4302 5290
rect 4256 5218 4262 5278
rect 4296 5218 4302 5278
rect 4256 5206 4302 5218
rect 4384 5278 4430 5290
rect 4384 5218 4390 5278
rect 4424 5218 4430 5278
rect 4384 5206 4430 5218
rect 4512 5278 4558 5290
rect 4512 5218 4518 5278
rect 4552 5218 4558 5278
rect 4512 5206 4558 5218
rect 8053 5278 8099 5290
rect 8053 5218 8059 5278
rect 8093 5218 8099 5278
rect 8053 5206 8099 5218
rect 8181 5278 8227 5290
rect 8181 5218 8187 5278
rect 8221 5218 8227 5278
rect 8181 5206 8227 5218
rect 8309 5278 8355 5290
rect 8309 5218 8315 5278
rect 8349 5218 8355 5278
rect 8309 5206 8355 5218
rect 8437 5278 8483 5290
rect 8437 5218 8443 5278
rect 8477 5218 8483 5278
rect 8437 5206 8483 5218
rect 8565 5278 8611 5290
rect 8565 5218 8571 5278
rect 8605 5218 8611 5278
rect 8565 5206 8611 5218
rect 8693 5278 8739 5290
rect 8693 5218 8699 5278
rect 8733 5218 8739 5278
rect 8693 5206 8739 5218
rect 8821 5278 8867 5290
rect 8821 5218 8827 5278
rect 8861 5218 8867 5278
rect 8821 5206 8867 5218
rect 8949 5278 8995 5290
rect 8949 5218 8955 5278
rect 8989 5218 8995 5278
rect 8949 5206 8995 5218
rect 9077 5278 9123 5290
rect 9077 5218 9083 5278
rect 9117 5218 9123 5278
rect 9077 5206 9123 5218
rect 9205 5278 9251 5290
rect 9205 5218 9211 5278
rect 9245 5218 9251 5278
rect 9205 5206 9251 5218
rect 9333 5278 9379 5290
rect 9333 5218 9339 5278
rect 9373 5218 9379 5278
rect 9333 5206 9379 5218
rect 9461 5278 9507 5290
rect 9461 5218 9467 5278
rect 9501 5218 9507 5278
rect 9461 5206 9507 5218
rect 9589 5278 9635 5290
rect 9589 5218 9595 5278
rect 9629 5218 9635 5278
rect 9589 5206 9635 5218
rect 9717 5278 9763 5290
rect 9717 5218 9723 5278
rect 9757 5218 9763 5278
rect 9717 5206 9763 5218
rect 9845 5278 9891 5290
rect 9845 5218 9851 5278
rect 9885 5218 9891 5278
rect 9845 5206 9891 5218
rect 9973 5278 10019 5290
rect 9973 5218 9979 5278
rect 10013 5218 10019 5278
rect 9973 5206 10019 5218
rect 10101 5278 10147 5290
rect 10101 5218 10107 5278
rect 10141 5218 10147 5278
rect 10101 5206 10147 5218
rect 15211 5278 15257 5290
rect 15211 5218 15217 5278
rect 15251 5218 15257 5278
rect 15211 5206 15257 5218
rect 15339 5278 15385 5290
rect 15339 5218 15345 5278
rect 15379 5218 15385 5278
rect 15339 5206 15385 5218
rect 15467 5278 15513 5290
rect 15467 5218 15473 5278
rect 15507 5218 15513 5278
rect 15467 5206 15513 5218
rect 15595 5278 15641 5290
rect 15595 5218 15601 5278
rect 15635 5218 15641 5278
rect 15595 5206 15641 5218
rect 15723 5278 15769 5290
rect 15723 5218 15729 5278
rect 15763 5218 15769 5278
rect 15723 5206 15769 5218
rect 15851 5278 15897 5290
rect 15851 5218 15857 5278
rect 15891 5218 15897 5278
rect 15851 5206 15897 5218
rect 15979 5278 16025 5290
rect 15979 5218 15985 5278
rect 16019 5218 16025 5278
rect 15979 5206 16025 5218
rect 16107 5278 16153 5290
rect 16107 5218 16113 5278
rect 16147 5218 16153 5278
rect 16107 5206 16153 5218
rect 16235 5278 16281 5290
rect 16235 5218 16241 5278
rect 16275 5218 16281 5278
rect 16235 5206 16281 5218
rect 16363 5278 16409 5290
rect 16363 5218 16369 5278
rect 16403 5218 16409 5278
rect 16363 5206 16409 5218
rect 16491 5278 16537 5290
rect 16491 5218 16497 5278
rect 16531 5218 16537 5278
rect 16491 5206 16537 5218
rect 16619 5278 16665 5290
rect 16619 5218 16625 5278
rect 16659 5218 16665 5278
rect 16619 5206 16665 5218
rect 16747 5278 16793 5290
rect 16747 5218 16753 5278
rect 16787 5218 16793 5278
rect 16747 5206 16793 5218
rect 16875 5278 16921 5290
rect 16875 5218 16881 5278
rect 16915 5218 16921 5278
rect 16875 5206 16921 5218
rect 17003 5278 17049 5290
rect 17003 5218 17009 5278
rect 17043 5218 17049 5278
rect 17003 5206 17049 5218
rect 17131 5278 17177 5290
rect 17131 5218 17137 5278
rect 17171 5218 17177 5278
rect 17131 5206 17177 5218
rect 17259 5278 17305 5290
rect 17259 5218 17265 5278
rect 17299 5218 17305 5278
rect 17259 5206 17305 5218
rect 17387 5278 17433 5290
rect 17387 5218 17393 5278
rect 17427 5218 17433 5278
rect 17387 5206 17433 5218
rect 17515 5278 17561 5290
rect 17515 5218 17521 5278
rect 17555 5218 17561 5278
rect 17515 5206 17561 5218
rect 17643 5278 17689 5290
rect 17643 5218 17649 5278
rect 17683 5218 17689 5278
rect 17643 5206 17689 5218
rect 17771 5278 17817 5290
rect 17771 5218 17777 5278
rect 17811 5218 17817 5278
rect 17771 5206 17817 5218
rect 17899 5278 17945 5290
rect 17899 5218 17905 5278
rect 17939 5218 17945 5278
rect 17899 5206 17945 5218
rect 18027 5278 18073 5290
rect 18027 5218 18033 5278
rect 18067 5218 18073 5278
rect 18027 5206 18073 5218
rect 18155 5278 18201 5290
rect 18155 5218 18161 5278
rect 18195 5218 18201 5278
rect 18155 5206 18201 5218
rect 18283 5278 18329 5290
rect 18283 5218 18289 5278
rect 18323 5218 18329 5278
rect 18283 5206 18329 5218
rect 18411 5278 18457 5290
rect 18411 5218 18417 5278
rect 18451 5218 18457 5278
rect 18411 5206 18457 5218
rect 18539 5278 18585 5290
rect 18539 5218 18545 5278
rect 18579 5218 18585 5278
rect 18539 5206 18585 5218
rect 18667 5278 18713 5290
rect 18667 5218 18673 5278
rect 18707 5218 18713 5278
rect 18667 5206 18713 5218
rect 18795 5278 18841 5290
rect 18795 5218 18801 5278
rect 18835 5218 18841 5278
rect 18795 5206 18841 5218
rect 18923 5278 18969 5290
rect 18923 5218 18929 5278
rect 18963 5218 18969 5278
rect 18923 5206 18969 5218
rect 19051 5278 19097 5290
rect 19051 5218 19057 5278
rect 19091 5218 19097 5278
rect 19051 5206 19097 5218
rect 19179 5278 19225 5290
rect 19179 5218 19185 5278
rect 19219 5218 19225 5278
rect 19179 5206 19225 5218
rect 19307 5278 19353 5290
rect 19307 5218 19313 5278
rect 19347 5218 19353 5278
rect 19307 5206 19353 5218
rect 20265 5278 20311 5290
rect 20265 5218 20271 5278
rect 20305 5218 20311 5278
rect 20265 5206 20311 5218
rect 20393 5278 20439 5290
rect 20393 5218 20399 5278
rect 20433 5218 20439 5278
rect 20393 5206 20439 5218
rect 20521 5278 20567 5290
rect 20521 5218 20527 5278
rect 20561 5218 20567 5278
rect 20521 5206 20567 5218
rect 20649 5278 20695 5290
rect 20649 5218 20655 5278
rect 20689 5218 20695 5278
rect 20649 5206 20695 5218
rect 20777 5278 20823 5290
rect 20777 5218 20783 5278
rect 20817 5218 20823 5278
rect 20777 5206 20823 5218
rect 20905 5278 20951 5290
rect 20905 5218 20911 5278
rect 20945 5218 20951 5278
rect 20905 5206 20951 5218
rect 21033 5278 21079 5290
rect 21033 5218 21039 5278
rect 21073 5218 21079 5278
rect 21033 5206 21079 5218
rect 21161 5278 21207 5290
rect 21161 5218 21167 5278
rect 21201 5218 21207 5278
rect 21161 5206 21207 5218
rect 21289 5278 21335 5290
rect 21289 5218 21295 5278
rect 21329 5218 21335 5278
rect 21289 5206 21335 5218
rect 21417 5278 21463 5290
rect 21417 5218 21423 5278
rect 21457 5218 21463 5278
rect 21417 5206 21463 5218
rect 21545 5278 21591 5290
rect 21545 5218 21551 5278
rect 21585 5218 21591 5278
rect 21545 5206 21591 5218
rect 21673 5278 21719 5290
rect 21673 5218 21679 5278
rect 21713 5218 21719 5278
rect 21673 5206 21719 5218
rect 21801 5278 21847 5290
rect 21801 5218 21807 5278
rect 21841 5218 21847 5278
rect 21801 5206 21847 5218
rect 21929 5278 21975 5290
rect 21929 5218 21935 5278
rect 21969 5218 21975 5278
rect 21929 5206 21975 5218
rect 22057 5278 22103 5290
rect 22057 5218 22063 5278
rect 22097 5218 22103 5278
rect 22057 5206 22103 5218
rect 22185 5278 22231 5290
rect 22185 5218 22191 5278
rect 22225 5218 22231 5278
rect 22185 5206 22231 5218
rect 22313 5278 22359 5290
rect 22313 5218 22319 5278
rect 22353 5218 22359 5278
rect 22313 5206 22359 5218
rect 22441 5278 22487 5290
rect 22441 5218 22447 5278
rect 22481 5218 22487 5278
rect 22441 5206 22487 5218
rect 22569 5278 22615 5290
rect 22569 5218 22575 5278
rect 22609 5218 22615 5278
rect 22569 5206 22615 5218
rect 22697 5278 22743 5290
rect 22697 5218 22703 5278
rect 22737 5218 22743 5278
rect 22697 5206 22743 5218
rect 22825 5278 22871 5290
rect 22825 5218 22831 5278
rect 22865 5218 22871 5278
rect 22825 5206 22871 5218
rect 22953 5278 22999 5290
rect 22953 5218 22959 5278
rect 22993 5218 22999 5278
rect 22953 5206 22999 5218
rect 23081 5278 23127 5290
rect 23081 5218 23087 5278
rect 23121 5218 23127 5278
rect 23081 5206 23127 5218
rect 23209 5278 23255 5290
rect 23209 5218 23215 5278
rect 23249 5218 23255 5278
rect 23209 5206 23255 5218
rect 23337 5278 23383 5290
rect 23337 5218 23343 5278
rect 23377 5218 23383 5278
rect 23337 5206 23383 5218
rect 23465 5278 23511 5290
rect 23465 5218 23471 5278
rect 23505 5218 23511 5278
rect 23465 5206 23511 5218
rect 23593 5278 23639 5290
rect 23593 5218 23599 5278
rect 23633 5218 23639 5278
rect 23593 5206 23639 5218
rect 23721 5278 23767 5290
rect 23721 5218 23727 5278
rect 23761 5218 23767 5278
rect 23721 5206 23767 5218
rect 23849 5278 23895 5290
rect 23849 5218 23855 5278
rect 23889 5218 23895 5278
rect 23849 5206 23895 5218
rect 23977 5278 24023 5290
rect 23977 5218 23983 5278
rect 24017 5218 24023 5278
rect 23977 5206 24023 5218
rect 24105 5278 24151 5290
rect 24105 5218 24111 5278
rect 24145 5218 24151 5278
rect 24105 5206 24151 5218
rect 24233 5278 24279 5290
rect 24233 5218 24239 5278
rect 24273 5218 24279 5278
rect 24233 5206 24279 5218
rect 24361 5278 24407 5290
rect 24361 5218 24367 5278
rect 24401 5218 24407 5278
rect 24361 5206 24407 5218
rect 24489 5278 24535 5290
rect 24489 5218 24495 5278
rect 24529 5218 24535 5278
rect 24489 5206 24535 5218
rect 24617 5278 24663 5290
rect 24617 5218 24623 5278
rect 24657 5218 24663 5278
rect 24617 5206 24663 5218
rect 24745 5278 24791 5290
rect 24745 5218 24751 5278
rect 24785 5218 24791 5278
rect 24745 5206 24791 5218
rect 24873 5278 24919 5290
rect 24873 5218 24879 5278
rect 24913 5218 24919 5278
rect 24873 5206 24919 5218
rect 25001 5278 25047 5290
rect 25001 5218 25007 5278
rect 25041 5218 25047 5278
rect 25001 5206 25047 5218
rect 25129 5278 25175 5290
rect 25129 5218 25135 5278
rect 25169 5218 25175 5278
rect 25129 5206 25175 5218
rect 25257 5278 25303 5290
rect 25257 5218 25263 5278
rect 25297 5218 25303 5278
rect 25257 5206 25303 5218
rect 25385 5278 25431 5290
rect 25385 5218 25391 5278
rect 25425 5218 25431 5278
rect 25385 5206 25431 5218
rect 25513 5278 25559 5290
rect 25513 5218 25519 5278
rect 25553 5218 25559 5278
rect 25513 5206 25559 5218
rect 25641 5278 25687 5290
rect 25641 5218 25647 5278
rect 25681 5218 25687 5278
rect 25641 5206 25687 5218
rect 25769 5278 25815 5290
rect 25769 5218 25775 5278
rect 25809 5218 25815 5278
rect 25769 5206 25815 5218
rect 25897 5278 25943 5290
rect 25897 5218 25903 5278
rect 25937 5218 25943 5278
rect 25897 5206 25943 5218
rect 26025 5278 26071 5290
rect 26025 5218 26031 5278
rect 26065 5218 26071 5278
rect 26025 5206 26071 5218
rect 26153 5278 26199 5290
rect 26153 5218 26159 5278
rect 26193 5218 26199 5278
rect 26153 5206 26199 5218
rect 26281 5278 26327 5290
rect 26281 5218 26287 5278
rect 26321 5218 26327 5278
rect 26281 5206 26327 5218
rect 26409 5278 26455 5290
rect 26409 5218 26415 5278
rect 26449 5218 26455 5278
rect 26409 5206 26455 5218
rect 26537 5278 26583 5290
rect 26537 5218 26543 5278
rect 26577 5218 26583 5278
rect 26537 5206 26583 5218
rect 26665 5278 26711 5290
rect 26665 5218 26671 5278
rect 26705 5218 26711 5278
rect 26665 5206 26711 5218
rect 26793 5278 26839 5290
rect 26793 5218 26799 5278
rect 26833 5218 26839 5278
rect 26793 5206 26839 5218
rect 26921 5278 26967 5290
rect 26921 5218 26927 5278
rect 26961 5218 26967 5278
rect 26921 5206 26967 5218
rect 27049 5278 27095 5290
rect 27049 5218 27055 5278
rect 27089 5218 27095 5278
rect 27049 5206 27095 5218
rect 27177 5278 27223 5290
rect 27177 5218 27183 5278
rect 27217 5218 27223 5278
rect 27177 5206 27223 5218
rect 27305 5278 27351 5290
rect 27305 5218 27311 5278
rect 27345 5218 27351 5278
rect 27305 5206 27351 5218
rect 27433 5278 27479 5290
rect 27433 5218 27439 5278
rect 27473 5218 27479 5278
rect 27433 5206 27479 5218
rect 27561 5278 27607 5290
rect 27561 5218 27567 5278
rect 27601 5218 27607 5278
rect 27561 5206 27607 5218
rect 27689 5278 27735 5290
rect 27689 5218 27695 5278
rect 27729 5218 27735 5278
rect 27689 5206 27735 5218
rect 27817 5278 27863 5290
rect 27817 5218 27823 5278
rect 27857 5218 27863 5278
rect 27817 5206 27863 5218
rect 27945 5278 27991 5290
rect 27945 5218 27951 5278
rect 27985 5218 27991 5278
rect 27945 5206 27991 5218
rect 28073 5278 28119 5290
rect 28073 5218 28079 5278
rect 28113 5218 28119 5278
rect 28073 5206 28119 5218
rect 28201 5278 28247 5290
rect 28201 5218 28207 5278
rect 28241 5218 28247 5278
rect 28201 5206 28247 5218
rect 28329 5278 28375 5290
rect 28329 5218 28335 5278
rect 28369 5218 28375 5278
rect 28329 5206 28375 5218
rect 28457 5278 28503 5290
rect 28457 5218 28463 5278
rect 28497 5218 28503 5278
rect 28457 5206 28503 5218
rect -317 5154 -283 5206
rect 611 5154 645 5206
rect 867 5154 901 5206
rect 1875 5154 1909 5206
rect 2131 5154 2165 5206
rect 2387 5154 2421 5206
rect 3494 5154 3528 5206
rect 3750 5154 3784 5206
rect 4006 5154 4040 5206
rect 4262 5154 4296 5206
rect 4518 5154 4552 5206
rect 8059 5154 8093 5206
rect 8315 5154 8349 5206
rect 8571 5154 8605 5206
rect 8827 5154 8861 5206
rect 9083 5154 9117 5206
rect 9339 5154 9373 5206
rect 9595 5154 9629 5206
rect 9851 5154 9885 5206
rect 10107 5154 10141 5206
rect 15217 5154 15251 5206
rect 15473 5154 15507 5206
rect 15729 5154 15763 5206
rect 15985 5154 16019 5206
rect 16241 5154 16275 5206
rect 16497 5154 16531 5206
rect 16753 5154 16787 5206
rect 17009 5154 17043 5206
rect 17265 5154 17299 5206
rect 17521 5154 17555 5206
rect 17777 5154 17811 5206
rect 18033 5154 18067 5206
rect 18289 5154 18323 5206
rect 18545 5154 18579 5206
rect 18801 5154 18835 5206
rect 19057 5154 19091 5206
rect 19313 5154 19347 5206
rect 20271 5154 20305 5206
rect 20527 5154 20561 5206
rect 20783 5154 20817 5206
rect 21039 5154 21073 5206
rect 21295 5154 21329 5206
rect 21551 5154 21585 5206
rect 21807 5154 21841 5206
rect 22063 5154 22097 5206
rect 22319 5154 22353 5206
rect 22575 5154 22609 5206
rect 22831 5154 22865 5206
rect 23087 5154 23121 5206
rect 23343 5154 23377 5206
rect 23599 5154 23633 5206
rect 23855 5154 23889 5206
rect 24111 5154 24145 5206
rect 24367 5154 24401 5206
rect 24623 5154 24657 5206
rect 24879 5154 24913 5206
rect 25135 5154 25169 5206
rect 25391 5154 25425 5206
rect 25647 5154 25681 5206
rect 25903 5154 25937 5206
rect 26159 5154 26193 5206
rect 26415 5154 26449 5206
rect 26671 5154 26705 5206
rect 26927 5154 26961 5206
rect 27183 5154 27217 5206
rect 27439 5154 27473 5206
rect 27695 5154 27729 5206
rect 27951 5154 27985 5206
rect 28207 5154 28241 5206
rect 28463 5154 28497 5206
rect 28825 5158 28889 5164
rect 28825 5154 28831 5158
rect -363 5148 28831 5154
rect -363 5110 -319 5148
rect -281 5110 -191 5148
rect -153 5110 609 5148
rect 647 5110 737 5148
rect 775 5110 865 5148
rect 903 5110 1873 5148
rect 1911 5110 2001 5148
rect 2039 5110 2129 5148
rect 2167 5110 2257 5148
rect 2295 5110 2385 5148
rect 2423 5110 3492 5148
rect 3530 5110 3620 5148
rect 3658 5110 3748 5148
rect 3786 5110 3876 5148
rect 3914 5110 4004 5148
rect 4042 5110 4132 5148
rect 4170 5110 4260 5148
rect 4298 5110 4388 5148
rect 4426 5110 4516 5148
rect 4554 5110 8057 5148
rect 8095 5110 8185 5148
rect 8223 5110 8313 5148
rect 8351 5110 8441 5148
rect 8479 5110 8569 5148
rect 8607 5110 8697 5148
rect 8735 5110 8825 5148
rect 8863 5110 8953 5148
rect 8991 5110 9081 5148
rect 9119 5110 9209 5148
rect 9247 5110 9337 5148
rect 9375 5110 9465 5148
rect 9503 5110 9593 5148
rect 9631 5110 9721 5148
rect 9759 5110 9849 5148
rect 9887 5110 9977 5148
rect 10015 5110 10105 5148
rect 10143 5110 15215 5148
rect 15253 5110 15343 5148
rect 15381 5110 15471 5148
rect 15509 5110 15599 5148
rect 15637 5110 15727 5148
rect 15765 5110 15855 5148
rect 15893 5110 15983 5148
rect 16021 5110 16111 5148
rect 16149 5110 16239 5148
rect 16277 5110 16367 5148
rect 16405 5110 16495 5148
rect 16533 5110 16623 5148
rect 16661 5110 16751 5148
rect 16789 5110 16879 5148
rect 16917 5110 17007 5148
rect 17045 5110 17135 5148
rect 17173 5110 17263 5148
rect 17301 5110 17391 5148
rect 17429 5110 17519 5148
rect 17557 5110 17647 5148
rect 17685 5110 17775 5148
rect 17813 5110 17903 5148
rect 17941 5110 18031 5148
rect 18069 5110 18159 5148
rect 18197 5110 18287 5148
rect 18325 5110 18415 5148
rect 18453 5110 18543 5148
rect 18581 5110 18671 5148
rect 18709 5110 18799 5148
rect 18837 5110 18927 5148
rect 18965 5110 19055 5148
rect 19093 5110 19183 5148
rect 19221 5110 19311 5148
rect 19349 5110 20269 5148
rect 20307 5110 20397 5148
rect 20435 5110 20525 5148
rect 20563 5110 20653 5148
rect 20691 5110 20781 5148
rect 20819 5110 20909 5148
rect 20947 5110 21037 5148
rect 21075 5110 21165 5148
rect 21203 5110 21293 5148
rect 21331 5110 21421 5148
rect 21459 5110 21549 5148
rect 21587 5110 21677 5148
rect 21715 5110 21805 5148
rect 21843 5110 21933 5148
rect 21971 5110 22061 5148
rect 22099 5110 22189 5148
rect 22227 5110 22317 5148
rect 22355 5110 22445 5148
rect 22483 5110 22573 5148
rect 22611 5110 22701 5148
rect 22739 5110 22829 5148
rect 22867 5110 22957 5148
rect 22995 5110 23085 5148
rect 23123 5110 23213 5148
rect 23251 5110 23341 5148
rect 23379 5110 23469 5148
rect 23507 5110 23597 5148
rect 23635 5110 23725 5148
rect 23763 5110 23853 5148
rect 23891 5110 23981 5148
rect 24019 5110 24109 5148
rect 24147 5110 24237 5148
rect 24275 5110 24365 5148
rect 24403 5110 24493 5148
rect 24531 5110 24621 5148
rect 24659 5110 24749 5148
rect 24787 5110 24877 5148
rect 24915 5110 25005 5148
rect 25043 5110 25133 5148
rect 25171 5110 25261 5148
rect 25299 5110 25389 5148
rect 25427 5110 25517 5148
rect 25555 5110 25645 5148
rect 25683 5110 25773 5148
rect 25811 5110 25901 5148
rect 25939 5110 26029 5148
rect 26067 5110 26157 5148
rect 26195 5110 26285 5148
rect 26323 5110 26413 5148
rect 26451 5110 26541 5148
rect 26579 5110 26669 5148
rect 26707 5110 26797 5148
rect 26835 5110 26925 5148
rect 26963 5110 27053 5148
rect 27091 5110 27181 5148
rect 27219 5110 27309 5148
rect 27347 5110 27437 5148
rect 27475 5110 27565 5148
rect 27603 5110 27693 5148
rect 27731 5110 27821 5148
rect 27859 5110 27949 5148
rect 27987 5110 28077 5148
rect 28115 5110 28205 5148
rect 28243 5110 28333 5148
rect 28371 5110 28461 5148
rect 28499 5110 28831 5148
rect -363 5106 28831 5110
rect 28883 5106 28889 5158
rect -363 5104 28889 5106
rect 28825 5100 28889 5104
rect 150 4070 210 4078
rect 150 4018 154 4070
rect 206 4018 210 4070
rect 150 4007 210 4018
rect 162 3998 196 4007
rect 10327 3271 10391 3282
rect 10327 3219 10332 3271
rect 10384 3219 10391 3271
rect 10327 3208 10391 3219
rect 10341 3204 10375 3208
rect 28633 3177 28697 3183
rect 5352 3163 5418 3174
rect 1270 3143 1330 3149
rect 1270 3091 1274 3143
rect 1326 3091 1330 3143
rect 1270 3082 1330 3091
rect 2804 3131 2864 3137
rect 358 3074 418 3080
rect 358 3022 362 3074
rect 414 3022 418 3074
rect 1282 3071 1316 3082
rect 2804 3079 2808 3131
rect 2860 3079 2864 3131
rect 5352 3111 5358 3163
rect 5410 3111 5418 3163
rect 28633 3125 28639 3177
rect 28691 3125 28697 3177
rect 28633 3119 28697 3125
rect 28647 3114 28681 3119
rect 5352 3100 5418 3111
rect 5367 3096 5401 3100
rect 2804 3070 2864 3079
rect 2816 3059 2850 3070
rect 358 3013 418 3022
rect 370 3002 404 3013
rect -93 2598 -33 2604
rect -93 2546 -89 2598
rect -37 2546 -33 2598
rect -93 2540 -33 2546
rect -81 2526 -47 2540
rect 964 2459 1024 2465
rect 964 2407 968 2459
rect 1020 2407 1024 2459
rect 964 2398 1024 2407
rect 2482 2459 2542 2465
rect 2482 2407 2486 2459
rect 2538 2407 2542 2459
rect 2482 2398 2542 2407
rect 4620 2449 4684 2455
rect 976 2387 1010 2398
rect 2494 2387 2528 2398
rect 4620 2397 4626 2449
rect 4678 2397 4684 2449
rect 4620 2391 4684 2397
rect 10200 2451 10266 2462
rect 10200 2399 10206 2451
rect 10258 2399 10266 2451
rect 19417 2459 19481 2465
rect 19417 2407 19423 2459
rect 19475 2407 19481 2459
rect 19417 2401 19481 2407
rect 20149 2460 20213 2466
rect 20149 2408 20155 2460
rect 20207 2408 20213 2460
rect 20149 2402 20213 2408
rect 4634 2377 4668 2391
rect 10200 2388 10266 2399
rect 19431 2396 19465 2401
rect 20163 2397 20197 2402
rect 10215 2379 10249 2388
<< via1 >>
rect 29508 6368 29560 6420
rect 28725 6285 28777 6337
rect -89 6031 -37 6083
rect 363 6009 415 6061
rect 1274 6009 1326 6061
rect 2809 5997 2861 6049
rect 5359 5995 5411 6047
rect 10332 5995 10384 6047
rect 28637 5995 28689 6047
rect 28830 5791 28882 5843
rect 29510 5684 29562 5736
rect 28725 5597 28777 5649
rect -89 5311 -37 5363
rect 968 5349 1020 5401
rect 2486 5312 2538 5364
rect 4626 5307 4678 5359
rect 10206 5310 10258 5362
rect 19422 5306 19474 5358
rect 20155 5306 20207 5358
rect 28831 5106 28883 5158
rect 154 4018 206 4070
rect 10332 3219 10384 3271
rect 1274 3091 1326 3143
rect 362 3022 414 3074
rect 2808 3079 2860 3131
rect 5358 3111 5410 3163
rect 28639 3125 28691 3177
rect -89 2546 -37 2598
rect 968 2407 1020 2459
rect 2486 2407 2538 2459
rect 4626 2397 4678 2449
rect 10206 2399 10258 2451
rect 19423 2407 19475 2459
rect 20155 2408 20207 2460
<< metal2 >>
rect 29502 6420 29566 6426
rect 29502 6368 29508 6420
rect 29560 6368 29566 6420
rect 29502 6362 29566 6368
rect 28719 6337 28783 6343
rect 28719 6285 28725 6337
rect 28777 6285 28783 6337
rect 81 6248 196 6281
rect 28719 6279 28783 6285
rect -95 6083 -31 6089
rect -95 6031 -89 6083
rect -37 6073 -31 6083
rect 81 6073 114 6248
rect -37 6040 114 6073
rect -37 6031 -31 6040
rect -95 6025 -31 6031
rect -95 5363 -31 5369
rect -95 5311 -89 5363
rect -37 5311 -31 5363
rect -95 5305 -31 5311
rect -80 2609 -47 5305
rect 163 4081 196 6248
rect 357 6061 421 6067
rect 357 6009 363 6061
rect 415 6009 421 6061
rect 357 6003 421 6009
rect 1268 6061 1332 6067
rect 1268 6009 1274 6061
rect 1326 6009 1332 6061
rect 28734 6058 28768 6279
rect 29518 6060 29552 6362
rect 29753 6061 29828 6063
rect 29749 6060 29828 6061
rect 28946 6058 29021 6060
rect 1268 6003 1332 6009
rect 2803 6049 2867 6055
rect 150 4072 210 4081
rect 150 4016 152 4072
rect 208 4016 210 4072
rect 150 4007 210 4016
rect 371 3085 405 6003
rect 962 5401 1026 5407
rect 962 5349 968 5401
rect 1020 5349 1026 5401
rect 962 5343 1026 5349
rect 358 3076 418 3085
rect 358 3020 360 3076
rect 416 3020 418 3076
rect 358 3011 418 3020
rect -93 2600 -33 2609
rect -93 2544 -91 2600
rect -35 2544 -33 2600
rect -93 2535 -33 2544
rect 977 2470 1011 5343
rect 1283 3154 1317 6003
rect 2803 5997 2809 6049
rect 2861 5997 2867 6049
rect 2803 5991 2867 5997
rect 5353 6047 5417 6053
rect 5353 5995 5359 6047
rect 5411 5995 5417 6047
rect 2480 5364 2544 5370
rect 2480 5312 2486 5364
rect 2538 5312 2544 5364
rect 2480 5306 2544 5312
rect 1270 3145 1330 3154
rect 1270 3089 1272 3145
rect 1328 3089 1330 3145
rect 1270 3080 1330 3089
rect 2495 2470 2529 5306
rect 2817 3142 2850 5991
rect 5353 5989 5417 5995
rect 10326 6047 10390 6053
rect 10326 5995 10332 6047
rect 10384 5995 10390 6047
rect 10326 5989 10390 5995
rect 28631 6047 28695 6053
rect 28631 5995 28637 6047
rect 28689 5995 28695 6047
rect 28631 5989 28695 5995
rect 28734 6051 29021 6058
rect 28734 5995 28955 6051
rect 29011 5995 29021 6051
rect 4620 5359 4684 5365
rect 4620 5307 4626 5359
rect 4678 5307 4684 5359
rect 4620 5301 4684 5307
rect 2804 3133 2864 3142
rect 2804 3077 2806 3133
rect 2862 3077 2864 3133
rect 2804 3068 2864 3077
rect 964 2461 1024 2470
rect 964 2405 966 2461
rect 1022 2405 1024 2461
rect 964 2396 1024 2405
rect 2482 2461 2542 2470
rect 2482 2405 2484 2461
rect 2540 2405 2542 2461
rect 4635 2460 4669 5301
rect 5367 3174 5401 5989
rect 10200 5362 10264 5368
rect 10200 5310 10206 5362
rect 10258 5310 10264 5362
rect 10200 5304 10264 5310
rect 5352 3165 5418 3174
rect 5352 3109 5357 3165
rect 5413 3109 5418 3165
rect 5352 3100 5418 3109
rect 10215 2462 10249 5304
rect 10341 3282 10375 5989
rect 19416 5358 19480 5364
rect 19416 5306 19422 5358
rect 19474 5306 19480 5358
rect 19416 5300 19480 5306
rect 20149 5358 20213 5364
rect 20149 5306 20155 5358
rect 20207 5306 20213 5358
rect 20149 5300 20213 5306
rect 10327 3273 10391 3282
rect 10327 3217 10331 3273
rect 10387 3217 10391 3273
rect 10327 3208 10391 3217
rect 19431 2470 19465 5300
rect 20163 2471 20197 5300
rect 28647 3188 28681 5989
rect 28734 5988 29021 5995
rect 28734 5655 28768 5988
rect 28946 5986 29021 5988
rect 29518 6054 29828 6060
rect 29518 5998 29762 6054
rect 29818 5998 29828 6054
rect 29518 5992 29828 5998
rect 28824 5843 28888 5849
rect 28824 5791 28830 5843
rect 28882 5791 28888 5843
rect 28824 5785 28888 5791
rect 28719 5649 28783 5655
rect 28719 5597 28725 5649
rect 28777 5597 28783 5649
rect 28719 5591 28783 5597
rect 28839 5429 28873 5785
rect 29518 5742 29552 5992
rect 29749 5991 29828 5992
rect 29753 5989 29828 5991
rect 29504 5736 29568 5742
rect 29504 5684 29510 5736
rect 29562 5684 29568 5736
rect 29504 5678 29568 5684
rect 28839 5425 28874 5429
rect 29142 5426 29217 5428
rect 29138 5425 29217 5426
rect 28839 5419 29217 5425
rect 28839 5363 29151 5419
rect 29207 5363 29217 5419
rect 28839 5357 29217 5363
rect 28839 5352 28874 5357
rect 29138 5356 29217 5357
rect 29142 5354 29217 5356
rect 28839 5164 28873 5352
rect 28825 5158 28889 5164
rect 28825 5106 28831 5158
rect 28883 5106 28889 5158
rect 28825 5100 28889 5106
rect 28633 3179 28697 3188
rect 28633 3123 28637 3179
rect 28693 3123 28697 3179
rect 28633 3114 28697 3123
rect 2482 2396 2542 2405
rect 4620 2451 4684 2460
rect 4620 2395 4624 2451
rect 4680 2395 4684 2451
rect 4620 2386 4684 2395
rect 10200 2453 10266 2462
rect 10200 2397 10205 2453
rect 10261 2397 10266 2453
rect 10200 2388 10266 2397
rect 19417 2461 19481 2470
rect 19417 2405 19421 2461
rect 19477 2405 19481 2461
rect 19417 2396 19481 2405
rect 20149 2462 20213 2471
rect 20149 2406 20153 2462
rect 20209 2406 20213 2462
rect 20149 2397 20213 2406
<< via2 >>
rect 152 4070 208 4072
rect 152 4018 154 4070
rect 154 4018 206 4070
rect 206 4018 208 4070
rect 152 4016 208 4018
rect 360 3074 416 3076
rect 360 3022 362 3074
rect 362 3022 414 3074
rect 414 3022 416 3074
rect 360 3020 416 3022
rect -91 2598 -35 2600
rect -91 2546 -89 2598
rect -89 2546 -37 2598
rect -37 2546 -35 2598
rect -91 2544 -35 2546
rect 1272 3143 1328 3145
rect 1272 3091 1274 3143
rect 1274 3091 1326 3143
rect 1326 3091 1328 3143
rect 1272 3089 1328 3091
rect 28955 5995 29011 6051
rect 2806 3131 2862 3133
rect 2806 3079 2808 3131
rect 2808 3079 2860 3131
rect 2860 3079 2862 3131
rect 2806 3077 2862 3079
rect 966 2459 1022 2461
rect 966 2407 968 2459
rect 968 2407 1020 2459
rect 1020 2407 1022 2459
rect 966 2405 1022 2407
rect 2484 2459 2540 2461
rect 2484 2407 2486 2459
rect 2486 2407 2538 2459
rect 2538 2407 2540 2459
rect 2484 2405 2540 2407
rect 5357 3163 5413 3165
rect 5357 3111 5358 3163
rect 5358 3111 5410 3163
rect 5410 3111 5413 3163
rect 5357 3109 5413 3111
rect 10331 3271 10387 3273
rect 10331 3219 10332 3271
rect 10332 3219 10384 3271
rect 10384 3219 10387 3271
rect 10331 3217 10387 3219
rect 29762 5998 29818 6054
rect 29151 5363 29207 5419
rect 28637 3177 28693 3179
rect 28637 3125 28639 3177
rect 28639 3125 28691 3177
rect 28691 3125 28693 3177
rect 28637 3123 28693 3125
rect 4624 2449 4680 2451
rect 4624 2397 4626 2449
rect 4626 2397 4678 2449
rect 4678 2397 4680 2449
rect 4624 2395 4680 2397
rect 10205 2451 10261 2453
rect 10205 2399 10206 2451
rect 10206 2399 10258 2451
rect 10258 2399 10261 2451
rect 10205 2397 10261 2399
rect 19421 2459 19477 2461
rect 19421 2407 19423 2459
rect 19423 2407 19475 2459
rect 19475 2407 19477 2459
rect 19421 2405 19477 2407
rect 20153 2460 20209 2462
rect 20153 2408 20155 2460
rect 20155 2408 20207 2460
rect 20207 2408 20209 2460
rect 20153 2406 20209 2408
<< metal3 >>
rect 28942 6055 29039 6075
rect 28942 5991 28951 6055
rect 29015 5991 29039 6055
rect 28942 5971 29039 5991
rect 29749 6058 29846 6078
rect 29749 5994 29758 6058
rect 29822 5994 29846 6058
rect 29749 5974 29846 5994
rect 29138 5423 29235 5443
rect 29138 5359 29147 5423
rect 29211 5359 29235 5423
rect 29138 5339 29235 5359
rect -459 5092 213 5094
rect -459 5028 -355 5092
rect -291 5028 -275 5092
rect -211 5028 -195 5092
rect -131 5028 -115 5092
rect -51 5028 -35 5092
rect 29 5028 45 5092
rect 109 5028 213 5092
rect -459 5026 213 5028
rect 355 5092 1027 5094
rect 355 5028 459 5092
rect 523 5028 539 5092
rect 603 5028 619 5092
rect 683 5028 699 5092
rect 763 5028 779 5092
rect 843 5028 859 5092
rect 923 5028 1027 5092
rect 355 5026 1027 5028
rect 1267 5092 2545 5094
rect 1267 5028 1371 5092
rect 1435 5028 1451 5092
rect 1515 5028 1531 5092
rect 1595 5028 1611 5092
rect 1675 5028 1691 5092
rect 1755 5028 1771 5092
rect 1835 5028 1977 5092
rect 2041 5028 2057 5092
rect 2121 5028 2137 5092
rect 2201 5028 2217 5092
rect 2281 5028 2297 5092
rect 2361 5028 2377 5092
rect 2441 5028 2545 5092
rect 1267 5026 2545 5028
rect 2801 5092 5291 5094
rect 2801 5028 2905 5092
rect 2969 5028 2985 5092
rect 3049 5028 3065 5092
rect 3129 5028 3145 5092
rect 3209 5028 3225 5092
rect 3289 5028 3305 5092
rect 3369 5028 3511 5092
rect 3575 5028 3591 5092
rect 3655 5028 3671 5092
rect 3735 5028 3751 5092
rect 3815 5028 3831 5092
rect 3895 5028 3911 5092
rect 3975 5028 4117 5092
rect 4181 5028 4197 5092
rect 4261 5028 4277 5092
rect 4341 5028 4357 5092
rect 4421 5028 4437 5092
rect 4501 5028 4517 5092
rect 4581 5028 4723 5092
rect 4787 5028 4803 5092
rect 4867 5028 4883 5092
rect 4947 5028 4963 5092
rect 5027 5028 5043 5092
rect 5107 5028 5123 5092
rect 5187 5028 5291 5092
rect 2801 5026 5291 5028
rect 5352 5092 10266 5094
rect 5352 5028 5456 5092
rect 5520 5028 5536 5092
rect 5600 5028 5616 5092
rect 5680 5028 5696 5092
rect 5760 5028 5776 5092
rect 5840 5028 5856 5092
rect 5920 5028 6062 5092
rect 6126 5028 6142 5092
rect 6206 5028 6222 5092
rect 6286 5028 6302 5092
rect 6366 5028 6382 5092
rect 6446 5028 6462 5092
rect 6526 5028 6668 5092
rect 6732 5028 6748 5092
rect 6812 5028 6828 5092
rect 6892 5028 6908 5092
rect 6972 5028 6988 5092
rect 7052 5028 7068 5092
rect 7132 5028 7274 5092
rect 7338 5028 7354 5092
rect 7418 5028 7434 5092
rect 7498 5028 7514 5092
rect 7578 5028 7594 5092
rect 7658 5028 7674 5092
rect 7738 5028 7880 5092
rect 7944 5028 7960 5092
rect 8024 5028 8040 5092
rect 8104 5028 8120 5092
rect 8184 5028 8200 5092
rect 8264 5028 8280 5092
rect 8344 5028 8486 5092
rect 8550 5028 8566 5092
rect 8630 5028 8646 5092
rect 8710 5028 8726 5092
rect 8790 5028 8806 5092
rect 8870 5028 8886 5092
rect 8950 5028 9092 5092
rect 9156 5028 9172 5092
rect 9236 5028 9252 5092
rect 9316 5028 9332 5092
rect 9396 5028 9412 5092
rect 9476 5028 9492 5092
rect 9556 5028 9698 5092
rect 9762 5028 9778 5092
rect 9842 5028 9858 5092
rect 9922 5028 9938 5092
rect 10002 5028 10018 5092
rect 10082 5028 10098 5092
rect 10162 5028 10266 5092
rect 5352 5026 10266 5028
rect 10326 5092 20088 5094
rect 10326 5028 10430 5092
rect 10494 5028 10510 5092
rect 10574 5028 10590 5092
rect 10654 5028 10670 5092
rect 10734 5028 10750 5092
rect 10814 5028 10830 5092
rect 10894 5028 11036 5092
rect 11100 5028 11116 5092
rect 11180 5028 11196 5092
rect 11260 5028 11276 5092
rect 11340 5028 11356 5092
rect 11420 5028 11436 5092
rect 11500 5028 11642 5092
rect 11706 5028 11722 5092
rect 11786 5028 11802 5092
rect 11866 5028 11882 5092
rect 11946 5028 11962 5092
rect 12026 5028 12042 5092
rect 12106 5028 12248 5092
rect 12312 5028 12328 5092
rect 12392 5028 12408 5092
rect 12472 5028 12488 5092
rect 12552 5028 12568 5092
rect 12632 5028 12648 5092
rect 12712 5028 12854 5092
rect 12918 5028 12934 5092
rect 12998 5028 13014 5092
rect 13078 5028 13094 5092
rect 13158 5028 13174 5092
rect 13238 5028 13254 5092
rect 13318 5028 13460 5092
rect 13524 5028 13540 5092
rect 13604 5028 13620 5092
rect 13684 5028 13700 5092
rect 13764 5028 13780 5092
rect 13844 5028 13860 5092
rect 13924 5028 14066 5092
rect 14130 5028 14146 5092
rect 14210 5028 14226 5092
rect 14290 5028 14306 5092
rect 14370 5028 14386 5092
rect 14450 5028 14466 5092
rect 14530 5028 14672 5092
rect 14736 5028 14752 5092
rect 14816 5028 14832 5092
rect 14896 5028 14912 5092
rect 14976 5028 14992 5092
rect 15056 5028 15072 5092
rect 15136 5028 15278 5092
rect 15342 5028 15358 5092
rect 15422 5028 15438 5092
rect 15502 5028 15518 5092
rect 15582 5028 15598 5092
rect 15662 5028 15678 5092
rect 15742 5028 15884 5092
rect 15948 5028 15964 5092
rect 16028 5028 16044 5092
rect 16108 5028 16124 5092
rect 16188 5028 16204 5092
rect 16268 5028 16284 5092
rect 16348 5028 16490 5092
rect 16554 5028 16570 5092
rect 16634 5028 16650 5092
rect 16714 5028 16730 5092
rect 16794 5028 16810 5092
rect 16874 5028 16890 5092
rect 16954 5028 17096 5092
rect 17160 5028 17176 5092
rect 17240 5028 17256 5092
rect 17320 5028 17336 5092
rect 17400 5028 17416 5092
rect 17480 5028 17496 5092
rect 17560 5028 17702 5092
rect 17766 5028 17782 5092
rect 17846 5028 17862 5092
rect 17926 5028 17942 5092
rect 18006 5028 18022 5092
rect 18086 5028 18102 5092
rect 18166 5028 18308 5092
rect 18372 5028 18388 5092
rect 18452 5028 18468 5092
rect 18532 5028 18548 5092
rect 18612 5028 18628 5092
rect 18692 5028 18708 5092
rect 18772 5028 18914 5092
rect 18978 5028 18994 5092
rect 19058 5028 19074 5092
rect 19138 5028 19154 5092
rect 19218 5028 19234 5092
rect 19298 5028 19314 5092
rect 19378 5028 19520 5092
rect 19584 5028 19600 5092
rect 19664 5028 19680 5092
rect 19744 5028 19760 5092
rect 19824 5028 19840 5092
rect 19904 5028 19920 5092
rect 19984 5028 20088 5092
rect 10326 5026 20088 5028
rect 20148 5092 39606 5094
rect 20148 5028 20252 5092
rect 20316 5028 20332 5092
rect 20396 5028 20412 5092
rect 20476 5028 20492 5092
rect 20556 5028 20572 5092
rect 20636 5028 20652 5092
rect 20716 5028 20858 5092
rect 20922 5028 20938 5092
rect 21002 5028 21018 5092
rect 21082 5028 21098 5092
rect 21162 5028 21178 5092
rect 21242 5028 21258 5092
rect 21322 5028 21464 5092
rect 21528 5028 21544 5092
rect 21608 5028 21624 5092
rect 21688 5028 21704 5092
rect 21768 5028 21784 5092
rect 21848 5028 21864 5092
rect 21928 5028 22070 5092
rect 22134 5028 22150 5092
rect 22214 5028 22230 5092
rect 22294 5028 22310 5092
rect 22374 5028 22390 5092
rect 22454 5028 22470 5092
rect 22534 5028 22676 5092
rect 22740 5028 22756 5092
rect 22820 5028 22836 5092
rect 22900 5028 22916 5092
rect 22980 5028 22996 5092
rect 23060 5028 23076 5092
rect 23140 5028 23282 5092
rect 23346 5028 23362 5092
rect 23426 5028 23442 5092
rect 23506 5028 23522 5092
rect 23586 5028 23602 5092
rect 23666 5028 23682 5092
rect 23746 5028 23888 5092
rect 23952 5028 23968 5092
rect 24032 5028 24048 5092
rect 24112 5028 24128 5092
rect 24192 5028 24208 5092
rect 24272 5028 24288 5092
rect 24352 5028 24494 5092
rect 24558 5028 24574 5092
rect 24638 5028 24654 5092
rect 24718 5028 24734 5092
rect 24798 5028 24814 5092
rect 24878 5028 24894 5092
rect 24958 5028 25100 5092
rect 25164 5028 25180 5092
rect 25244 5028 25260 5092
rect 25324 5028 25340 5092
rect 25404 5028 25420 5092
rect 25484 5028 25500 5092
rect 25564 5028 25706 5092
rect 25770 5028 25786 5092
rect 25850 5028 25866 5092
rect 25930 5028 25946 5092
rect 26010 5028 26026 5092
rect 26090 5028 26106 5092
rect 26170 5028 26312 5092
rect 26376 5028 26392 5092
rect 26456 5028 26472 5092
rect 26536 5028 26552 5092
rect 26616 5028 26632 5092
rect 26696 5028 26712 5092
rect 26776 5028 26918 5092
rect 26982 5028 26998 5092
rect 27062 5028 27078 5092
rect 27142 5028 27158 5092
rect 27222 5028 27238 5092
rect 27302 5028 27318 5092
rect 27382 5028 27524 5092
rect 27588 5028 27604 5092
rect 27668 5028 27684 5092
rect 27748 5028 27764 5092
rect 27828 5028 27844 5092
rect 27908 5028 27924 5092
rect 27988 5028 28130 5092
rect 28194 5028 28210 5092
rect 28274 5028 28290 5092
rect 28354 5028 28370 5092
rect 28434 5028 28450 5092
rect 28514 5028 28530 5092
rect 28594 5028 28736 5092
rect 28800 5028 28816 5092
rect 28880 5028 28896 5092
rect 28960 5028 28976 5092
rect 29040 5028 29056 5092
rect 29120 5028 29136 5092
rect 29200 5028 29342 5092
rect 29406 5028 29422 5092
rect 29486 5028 29502 5092
rect 29566 5028 29582 5092
rect 29646 5028 29662 5092
rect 29726 5028 29742 5092
rect 29806 5028 29948 5092
rect 30012 5028 30028 5092
rect 30092 5028 30108 5092
rect 30172 5028 30188 5092
rect 30252 5028 30268 5092
rect 30332 5028 30348 5092
rect 30412 5028 30554 5092
rect 30618 5028 30634 5092
rect 30698 5028 30714 5092
rect 30778 5028 30794 5092
rect 30858 5028 30874 5092
rect 30938 5028 30954 5092
rect 31018 5028 31160 5092
rect 31224 5028 31240 5092
rect 31304 5028 31320 5092
rect 31384 5028 31400 5092
rect 31464 5028 31480 5092
rect 31544 5028 31560 5092
rect 31624 5028 31766 5092
rect 31830 5028 31846 5092
rect 31910 5028 31926 5092
rect 31990 5028 32006 5092
rect 32070 5028 32086 5092
rect 32150 5028 32166 5092
rect 32230 5028 32372 5092
rect 32436 5028 32452 5092
rect 32516 5028 32532 5092
rect 32596 5028 32612 5092
rect 32676 5028 32692 5092
rect 32756 5028 32772 5092
rect 32836 5028 32978 5092
rect 33042 5028 33058 5092
rect 33122 5028 33138 5092
rect 33202 5028 33218 5092
rect 33282 5028 33298 5092
rect 33362 5028 33378 5092
rect 33442 5028 33584 5092
rect 33648 5028 33664 5092
rect 33728 5028 33744 5092
rect 33808 5028 33824 5092
rect 33888 5028 33904 5092
rect 33968 5028 33984 5092
rect 34048 5028 34190 5092
rect 34254 5028 34270 5092
rect 34334 5028 34350 5092
rect 34414 5028 34430 5092
rect 34494 5028 34510 5092
rect 34574 5028 34590 5092
rect 34654 5028 34796 5092
rect 34860 5028 34876 5092
rect 34940 5028 34956 5092
rect 35020 5028 35036 5092
rect 35100 5028 35116 5092
rect 35180 5028 35196 5092
rect 35260 5028 35402 5092
rect 35466 5028 35482 5092
rect 35546 5028 35562 5092
rect 35626 5028 35642 5092
rect 35706 5028 35722 5092
rect 35786 5028 35802 5092
rect 35866 5028 36008 5092
rect 36072 5028 36088 5092
rect 36152 5028 36168 5092
rect 36232 5028 36248 5092
rect 36312 5028 36328 5092
rect 36392 5028 36408 5092
rect 36472 5028 36614 5092
rect 36678 5028 36694 5092
rect 36758 5028 36774 5092
rect 36838 5028 36854 5092
rect 36918 5028 36934 5092
rect 36998 5028 37014 5092
rect 37078 5028 37220 5092
rect 37284 5028 37300 5092
rect 37364 5028 37380 5092
rect 37444 5028 37460 5092
rect 37524 5028 37540 5092
rect 37604 5028 37620 5092
rect 37684 5028 37826 5092
rect 37890 5028 37906 5092
rect 37970 5028 37986 5092
rect 38050 5028 38066 5092
rect 38130 5028 38146 5092
rect 38210 5028 38226 5092
rect 38290 5028 38432 5092
rect 38496 5028 38512 5092
rect 38576 5028 38592 5092
rect 38656 5028 38672 5092
rect 38736 5028 38752 5092
rect 38816 5028 38832 5092
rect 38896 5028 39038 5092
rect 39102 5028 39118 5092
rect 39182 5028 39198 5092
rect 39262 5028 39278 5092
rect 39342 5028 39358 5092
rect 39422 5028 39438 5092
rect 39502 5028 39606 5092
rect 20148 5026 39606 5028
rect -459 4872 -393 5026
rect -459 4808 -458 4872
rect -394 4808 -393 4872
rect -459 4792 -393 4808
rect -459 4728 -458 4792
rect -394 4728 -393 4792
rect -459 4712 -393 4728
rect -459 4648 -458 4712
rect -394 4648 -393 4712
rect -459 4632 -393 4648
rect -459 4568 -458 4632
rect -394 4568 -393 4632
rect -459 4552 -393 4568
rect -459 4488 -458 4552
rect -394 4488 -393 4552
rect -459 4472 -393 4488
rect -459 4408 -458 4472
rect -394 4408 -393 4472
rect -459 4392 -393 4408
rect -459 4328 -458 4392
rect -394 4328 -393 4392
rect -459 4312 -393 4328
rect -459 4248 -458 4312
rect -394 4248 -393 4312
rect -459 4232 -393 4248
rect -459 4168 -458 4232
rect -394 4168 -393 4232
rect -459 4152 -393 4168
rect -459 4088 -458 4152
rect -394 4088 -393 4152
rect -459 3998 -393 4088
rect -333 3934 -273 4964
rect -213 3994 -153 5026
rect -93 3934 -33 4964
rect 27 3994 87 5026
rect 147 4872 213 5026
rect 147 4808 148 4872
rect 212 4808 213 4872
rect 147 4792 213 4808
rect 147 4728 148 4792
rect 212 4728 213 4792
rect 147 4712 213 4728
rect 147 4648 148 4712
rect 212 4648 213 4712
rect 147 4632 213 4648
rect 147 4568 148 4632
rect 212 4568 213 4632
rect 147 4552 213 4568
rect 147 4488 148 4552
rect 212 4488 213 4552
rect 147 4472 213 4488
rect 147 4408 148 4472
rect 212 4408 213 4472
rect 147 4392 213 4408
rect 147 4328 148 4392
rect 212 4328 213 4392
rect 147 4312 213 4328
rect 147 4248 148 4312
rect 212 4248 213 4312
rect 147 4232 213 4248
rect 147 4168 148 4232
rect 212 4168 213 4232
rect 147 4152 213 4168
rect 147 4088 148 4152
rect 212 4088 213 4152
rect 147 4072 213 4088
rect 147 4016 152 4072
rect 208 4016 213 4072
rect 147 3998 213 4016
rect 355 4872 421 4962
rect 355 4808 356 4872
rect 420 4808 421 4872
rect 355 4792 421 4808
rect 355 4728 356 4792
rect 420 4728 421 4792
rect 355 4712 421 4728
rect 355 4648 356 4712
rect 420 4648 421 4712
rect 355 4632 421 4648
rect 355 4568 356 4632
rect 420 4568 421 4632
rect 355 4552 421 4568
rect 355 4488 356 4552
rect 420 4488 421 4552
rect 355 4472 421 4488
rect 355 4408 356 4472
rect 420 4408 421 4472
rect 355 4392 421 4408
rect 355 4328 356 4392
rect 420 4328 421 4392
rect 355 4312 421 4328
rect 355 4248 356 4312
rect 420 4248 421 4312
rect 355 4232 421 4248
rect 355 4168 356 4232
rect 420 4168 421 4232
rect 355 4152 421 4168
rect 355 4088 356 4152
rect 420 4088 421 4152
rect 355 3934 421 4088
rect 481 3934 541 4966
rect 601 3996 661 5026
rect 721 3934 781 4966
rect 841 3996 901 5026
rect 961 4872 1027 4962
rect 961 4808 962 4872
rect 1026 4808 1027 4872
rect 961 4792 1027 4808
rect 961 4728 962 4792
rect 1026 4728 1027 4792
rect 961 4712 1027 4728
rect 961 4648 962 4712
rect 1026 4648 1027 4712
rect 961 4632 1027 4648
rect 961 4568 962 4632
rect 1026 4568 1027 4632
rect 961 4552 1027 4568
rect 961 4488 962 4552
rect 1026 4488 1027 4552
rect 961 4472 1027 4488
rect 961 4408 962 4472
rect 1026 4408 1027 4472
rect 961 4392 1027 4408
rect 961 4328 962 4392
rect 1026 4328 1027 4392
rect 961 4312 1027 4328
rect 961 4248 962 4312
rect 1026 4248 1027 4312
rect 961 4232 1027 4248
rect 961 4168 962 4232
rect 1026 4168 1027 4232
rect 961 4152 1027 4168
rect 961 4088 962 4152
rect 1026 4088 1027 4152
rect 961 3934 1027 4088
rect -459 3932 213 3934
rect -459 3868 -355 3932
rect -291 3868 -275 3932
rect -211 3868 -195 3932
rect -131 3868 -115 3932
rect -51 3868 -35 3932
rect 29 3868 45 3932
rect 109 3868 213 3932
rect -459 3866 213 3868
rect 355 3932 1027 3934
rect 355 3868 459 3932
rect 523 3868 539 3932
rect 603 3868 619 3932
rect 683 3868 699 3932
rect 763 3868 779 3932
rect 843 3868 859 3932
rect 923 3868 1027 3932
rect 355 3866 1027 3868
rect -459 3712 -393 3802
rect -459 3648 -458 3712
rect -394 3648 -393 3712
rect -459 3632 -393 3648
rect -459 3568 -458 3632
rect -394 3568 -393 3632
rect -459 3552 -393 3568
rect -459 3488 -458 3552
rect -394 3488 -393 3552
rect -459 3472 -393 3488
rect -459 3408 -458 3472
rect -394 3408 -393 3472
rect -459 3392 -393 3408
rect -459 3328 -458 3392
rect -394 3328 -393 3392
rect -459 3312 -393 3328
rect -459 3248 -458 3312
rect -394 3248 -393 3312
rect -459 3232 -393 3248
rect -459 3168 -458 3232
rect -394 3168 -393 3232
rect -459 3152 -393 3168
rect -459 3088 -458 3152
rect -394 3088 -393 3152
rect -459 3072 -393 3088
rect -459 3008 -458 3072
rect -394 3008 -393 3072
rect -459 2992 -393 3008
rect -459 2928 -458 2992
rect -394 2928 -393 2992
rect -459 2774 -393 2928
rect -333 2774 -273 3806
rect -213 2836 -153 3866
rect -93 2774 -33 3806
rect 27 2836 87 3866
rect 147 3712 213 3802
rect 147 3648 148 3712
rect 212 3648 213 3712
rect 147 3632 213 3648
rect 147 3568 148 3632
rect 212 3568 213 3632
rect 147 3552 213 3568
rect 147 3488 148 3552
rect 212 3488 213 3552
rect 147 3472 213 3488
rect 147 3408 148 3472
rect 212 3408 213 3472
rect 147 3392 213 3408
rect 147 3328 148 3392
rect 212 3328 213 3392
rect 147 3312 213 3328
rect 147 3248 148 3312
rect 212 3248 213 3312
rect 147 3232 213 3248
rect 147 3168 148 3232
rect 212 3168 213 3232
rect 147 3152 213 3168
rect 147 3088 148 3152
rect 212 3088 213 3152
rect 147 3072 213 3088
rect 147 3008 148 3072
rect 212 3008 213 3072
rect 147 2992 213 3008
rect 147 2928 148 2992
rect 212 2928 213 2992
rect 147 2774 213 2928
rect 355 3712 421 3866
rect 355 3648 356 3712
rect 420 3648 421 3712
rect 355 3632 421 3648
rect 355 3568 356 3632
rect 420 3568 421 3632
rect 355 3552 421 3568
rect 355 3488 356 3552
rect 420 3488 421 3552
rect 355 3472 421 3488
rect 355 3408 356 3472
rect 420 3408 421 3472
rect 355 3392 421 3408
rect 355 3328 356 3392
rect 420 3328 421 3392
rect 355 3312 421 3328
rect 355 3248 356 3312
rect 420 3248 421 3312
rect 355 3232 421 3248
rect 355 3168 356 3232
rect 420 3168 421 3232
rect 355 3152 421 3168
rect 355 3088 356 3152
rect 420 3088 421 3152
rect 355 3076 421 3088
rect 355 3072 360 3076
rect 416 3072 421 3076
rect 355 3008 356 3072
rect 420 3008 421 3072
rect 355 2992 421 3008
rect 355 2928 356 2992
rect 420 2928 421 2992
rect 355 2838 421 2928
rect 481 2774 541 3804
rect 601 2834 661 3866
rect 721 2774 781 3804
rect 841 2834 901 3866
rect 961 3712 1027 3866
rect 961 3648 962 3712
rect 1026 3648 1027 3712
rect 961 3632 1027 3648
rect 961 3568 962 3632
rect 1026 3568 1027 3632
rect 961 3552 1027 3568
rect 961 3488 962 3552
rect 1026 3488 1027 3552
rect 961 3472 1027 3488
rect 961 3408 962 3472
rect 1026 3408 1027 3472
rect 961 3392 1027 3408
rect 961 3328 962 3392
rect 1026 3328 1027 3392
rect 961 3312 1027 3328
rect 961 3248 962 3312
rect 1026 3248 1027 3312
rect 961 3232 1027 3248
rect 961 3168 962 3232
rect 1026 3168 1027 3232
rect 961 3152 1027 3168
rect 961 3088 962 3152
rect 1026 3088 1027 3152
rect 961 3072 1027 3088
rect 961 3008 962 3072
rect 1026 3008 1027 3072
rect 961 2992 1027 3008
rect 961 2928 962 2992
rect 1026 2928 1027 2992
rect 961 2838 1027 2928
rect 1267 4872 1333 4962
rect 1267 4808 1268 4872
rect 1332 4808 1333 4872
rect 1267 4792 1333 4808
rect 1267 4728 1268 4792
rect 1332 4728 1333 4792
rect 1267 4712 1333 4728
rect 1267 4648 1268 4712
rect 1332 4648 1333 4712
rect 1267 4632 1333 4648
rect 1267 4568 1268 4632
rect 1332 4568 1333 4632
rect 1267 4552 1333 4568
rect 1267 4488 1268 4552
rect 1332 4488 1333 4552
rect 1267 4472 1333 4488
rect 1267 4408 1268 4472
rect 1332 4408 1333 4472
rect 1267 4392 1333 4408
rect 1267 4328 1268 4392
rect 1332 4328 1333 4392
rect 1267 4312 1333 4328
rect 1267 4248 1268 4312
rect 1332 4248 1333 4312
rect 1267 4232 1333 4248
rect 1267 4168 1268 4232
rect 1332 4168 1333 4232
rect 1267 4152 1333 4168
rect 1267 4088 1268 4152
rect 1332 4088 1333 4152
rect 1267 3934 1333 4088
rect 1393 3934 1453 4966
rect 1513 3996 1573 5026
rect 1633 3934 1693 4966
rect 1753 3996 1813 5026
rect 1873 4872 1939 4962
rect 1873 4808 1874 4872
rect 1938 4808 1939 4872
rect 1873 4792 1939 4808
rect 1873 4728 1874 4792
rect 1938 4728 1939 4792
rect 1873 4712 1939 4728
rect 1873 4648 1874 4712
rect 1938 4648 1939 4712
rect 1873 4632 1939 4648
rect 1873 4568 1874 4632
rect 1938 4568 1939 4632
rect 1873 4552 1939 4568
rect 1873 4488 1874 4552
rect 1938 4488 1939 4552
rect 1873 4472 1939 4488
rect 1873 4408 1874 4472
rect 1938 4408 1939 4472
rect 1873 4392 1939 4408
rect 1873 4328 1874 4392
rect 1938 4328 1939 4392
rect 1873 4312 1939 4328
rect 1873 4248 1874 4312
rect 1938 4248 1939 4312
rect 1873 4232 1939 4248
rect 1873 4168 1874 4232
rect 1938 4168 1939 4232
rect 1873 4152 1939 4168
rect 1873 4088 1874 4152
rect 1938 4088 1939 4152
rect 1873 3934 1939 4088
rect 1999 3934 2059 4966
rect 2119 3996 2179 5026
rect 2239 3934 2299 4966
rect 2359 3996 2419 5026
rect 2479 4872 2545 4962
rect 2479 4808 2480 4872
rect 2544 4808 2545 4872
rect 2479 4792 2545 4808
rect 2479 4728 2480 4792
rect 2544 4728 2545 4792
rect 2479 4712 2545 4728
rect 2479 4648 2480 4712
rect 2544 4648 2545 4712
rect 2479 4632 2545 4648
rect 2479 4568 2480 4632
rect 2544 4568 2545 4632
rect 2479 4552 2545 4568
rect 2479 4488 2480 4552
rect 2544 4488 2545 4552
rect 2479 4472 2545 4488
rect 2479 4408 2480 4472
rect 2544 4408 2545 4472
rect 2479 4392 2545 4408
rect 2479 4328 2480 4392
rect 2544 4328 2545 4392
rect 2479 4312 2545 4328
rect 2479 4248 2480 4312
rect 2544 4248 2545 4312
rect 2479 4232 2545 4248
rect 2479 4168 2480 4232
rect 2544 4168 2545 4232
rect 2479 4152 2545 4168
rect 2479 4088 2480 4152
rect 2544 4088 2545 4152
rect 2479 3934 2545 4088
rect 1267 3932 2545 3934
rect 1267 3868 1371 3932
rect 1435 3868 1451 3932
rect 1515 3868 1531 3932
rect 1595 3868 1611 3932
rect 1675 3868 1691 3932
rect 1755 3868 1771 3932
rect 1835 3868 1977 3932
rect 2041 3868 2057 3932
rect 2121 3868 2137 3932
rect 2201 3868 2217 3932
rect 2281 3868 2297 3932
rect 2361 3868 2377 3932
rect 2441 3868 2545 3932
rect 1267 3866 2545 3868
rect 1267 3712 1333 3866
rect 1267 3648 1268 3712
rect 1332 3648 1333 3712
rect 1267 3632 1333 3648
rect 1267 3568 1268 3632
rect 1332 3568 1333 3632
rect 1267 3552 1333 3568
rect 1267 3488 1268 3552
rect 1332 3488 1333 3552
rect 1267 3472 1333 3488
rect 1267 3408 1268 3472
rect 1332 3408 1333 3472
rect 1267 3392 1333 3408
rect 1267 3328 1268 3392
rect 1332 3328 1333 3392
rect 1267 3312 1333 3328
rect 1267 3248 1268 3312
rect 1332 3248 1333 3312
rect 1267 3232 1333 3248
rect 1267 3168 1268 3232
rect 1332 3168 1333 3232
rect 1267 3152 1333 3168
rect 1267 3088 1268 3152
rect 1332 3088 1333 3152
rect 1267 3072 1333 3088
rect 1267 3008 1268 3072
rect 1332 3008 1333 3072
rect 1267 2992 1333 3008
rect 1267 2928 1268 2992
rect 1332 2928 1333 2992
rect 1267 2838 1333 2928
rect 1393 2774 1453 3804
rect 1513 2834 1573 3866
rect 1633 2774 1693 3804
rect 1753 2834 1813 3866
rect 1873 3712 1939 3866
rect 1873 3648 1874 3712
rect 1938 3648 1939 3712
rect 1873 3632 1939 3648
rect 1873 3568 1874 3632
rect 1938 3568 1939 3632
rect 1873 3552 1939 3568
rect 1873 3488 1874 3552
rect 1938 3488 1939 3552
rect 1873 3472 1939 3488
rect 1873 3408 1874 3472
rect 1938 3408 1939 3472
rect 1873 3392 1939 3408
rect 1873 3328 1874 3392
rect 1938 3328 1939 3392
rect 1873 3312 1939 3328
rect 1873 3248 1874 3312
rect 1938 3248 1939 3312
rect 1873 3232 1939 3248
rect 1873 3168 1874 3232
rect 1938 3168 1939 3232
rect 1873 3152 1939 3168
rect 1873 3088 1874 3152
rect 1938 3088 1939 3152
rect 1873 3072 1939 3088
rect 1873 3008 1874 3072
rect 1938 3008 1939 3072
rect 1873 2992 1939 3008
rect 1873 2928 1874 2992
rect 1938 2928 1939 2992
rect 1873 2838 1939 2928
rect 1999 2774 2059 3804
rect 2119 2834 2179 3866
rect 2239 2774 2299 3804
rect 2359 2834 2419 3866
rect 2479 3712 2545 3866
rect 2479 3648 2480 3712
rect 2544 3648 2545 3712
rect 2479 3632 2545 3648
rect 2479 3568 2480 3632
rect 2544 3568 2545 3632
rect 2479 3552 2545 3568
rect 2479 3488 2480 3552
rect 2544 3488 2545 3552
rect 2479 3472 2545 3488
rect 2479 3408 2480 3472
rect 2544 3408 2545 3472
rect 2479 3392 2545 3408
rect 2479 3328 2480 3392
rect 2544 3328 2545 3392
rect 2479 3312 2545 3328
rect 2479 3248 2480 3312
rect 2544 3248 2545 3312
rect 2479 3232 2545 3248
rect 2479 3168 2480 3232
rect 2544 3168 2545 3232
rect 2479 3152 2545 3168
rect 2479 3088 2480 3152
rect 2544 3088 2545 3152
rect 2479 3072 2545 3088
rect 2479 3008 2480 3072
rect 2544 3008 2545 3072
rect 2479 2992 2545 3008
rect 2479 2928 2480 2992
rect 2544 2928 2545 2992
rect 2479 2838 2545 2928
rect 2801 4872 2867 4962
rect 2801 4808 2802 4872
rect 2866 4808 2867 4872
rect 2801 4792 2867 4808
rect 2801 4728 2802 4792
rect 2866 4728 2867 4792
rect 2801 4712 2867 4728
rect 2801 4648 2802 4712
rect 2866 4648 2867 4712
rect 2801 4632 2867 4648
rect 2801 4568 2802 4632
rect 2866 4568 2867 4632
rect 2801 4552 2867 4568
rect 2801 4488 2802 4552
rect 2866 4488 2867 4552
rect 2801 4472 2867 4488
rect 2801 4408 2802 4472
rect 2866 4408 2867 4472
rect 2801 4392 2867 4408
rect 2801 4328 2802 4392
rect 2866 4328 2867 4392
rect 2801 4312 2867 4328
rect 2801 4248 2802 4312
rect 2866 4248 2867 4312
rect 2801 4232 2867 4248
rect 2801 4168 2802 4232
rect 2866 4168 2867 4232
rect 2801 4152 2867 4168
rect 2801 4088 2802 4152
rect 2866 4088 2867 4152
rect 2801 3934 2867 4088
rect 2927 3934 2987 4966
rect 3047 3996 3107 5026
rect 3167 3934 3227 4966
rect 3287 3996 3347 5026
rect 3407 4872 3473 4962
rect 3407 4808 3408 4872
rect 3472 4808 3473 4872
rect 3407 4792 3473 4808
rect 3407 4728 3408 4792
rect 3472 4728 3473 4792
rect 3407 4712 3473 4728
rect 3407 4648 3408 4712
rect 3472 4648 3473 4712
rect 3407 4632 3473 4648
rect 3407 4568 3408 4632
rect 3472 4568 3473 4632
rect 3407 4552 3473 4568
rect 3407 4488 3408 4552
rect 3472 4488 3473 4552
rect 3407 4472 3473 4488
rect 3407 4408 3408 4472
rect 3472 4408 3473 4472
rect 3407 4392 3473 4408
rect 3407 4328 3408 4392
rect 3472 4328 3473 4392
rect 3407 4312 3473 4328
rect 3407 4248 3408 4312
rect 3472 4248 3473 4312
rect 3407 4232 3473 4248
rect 3407 4168 3408 4232
rect 3472 4168 3473 4232
rect 3407 4152 3473 4168
rect 3407 4088 3408 4152
rect 3472 4088 3473 4152
rect 3407 3934 3473 4088
rect 3533 3934 3593 4966
rect 3653 3996 3713 5026
rect 3773 3934 3833 4966
rect 3893 3996 3953 5026
rect 4013 4872 4079 4962
rect 4013 4808 4014 4872
rect 4078 4808 4079 4872
rect 4013 4792 4079 4808
rect 4013 4728 4014 4792
rect 4078 4728 4079 4792
rect 4013 4712 4079 4728
rect 4013 4648 4014 4712
rect 4078 4648 4079 4712
rect 4013 4632 4079 4648
rect 4013 4568 4014 4632
rect 4078 4568 4079 4632
rect 4013 4552 4079 4568
rect 4013 4488 4014 4552
rect 4078 4488 4079 4552
rect 4013 4472 4079 4488
rect 4013 4408 4014 4472
rect 4078 4408 4079 4472
rect 4013 4392 4079 4408
rect 4013 4328 4014 4392
rect 4078 4328 4079 4392
rect 4013 4312 4079 4328
rect 4013 4248 4014 4312
rect 4078 4248 4079 4312
rect 4013 4232 4079 4248
rect 4013 4168 4014 4232
rect 4078 4168 4079 4232
rect 4013 4152 4079 4168
rect 4013 4088 4014 4152
rect 4078 4088 4079 4152
rect 4013 3934 4079 4088
rect 4139 3934 4199 4966
rect 4259 3996 4319 5026
rect 4379 3934 4439 4966
rect 4499 3996 4559 5026
rect 4619 4872 4685 4962
rect 4619 4808 4620 4872
rect 4684 4808 4685 4872
rect 4619 4792 4685 4808
rect 4619 4728 4620 4792
rect 4684 4728 4685 4792
rect 4619 4712 4685 4728
rect 4619 4648 4620 4712
rect 4684 4648 4685 4712
rect 4619 4632 4685 4648
rect 4619 4568 4620 4632
rect 4684 4568 4685 4632
rect 4619 4552 4685 4568
rect 4619 4488 4620 4552
rect 4684 4488 4685 4552
rect 4619 4472 4685 4488
rect 4619 4408 4620 4472
rect 4684 4408 4685 4472
rect 4619 4392 4685 4408
rect 4619 4328 4620 4392
rect 4684 4328 4685 4392
rect 4619 4312 4685 4328
rect 4619 4248 4620 4312
rect 4684 4248 4685 4312
rect 4619 4232 4685 4248
rect 4619 4168 4620 4232
rect 4684 4168 4685 4232
rect 4619 4152 4685 4168
rect 4619 4088 4620 4152
rect 4684 4088 4685 4152
rect 4619 3934 4685 4088
rect 4745 3934 4805 4966
rect 4865 3996 4925 5026
rect 4985 3934 5045 4966
rect 5105 3996 5165 5026
rect 5225 4872 5291 4962
rect 5225 4808 5226 4872
rect 5290 4808 5291 4872
rect 5225 4792 5291 4808
rect 5225 4728 5226 4792
rect 5290 4728 5291 4792
rect 5225 4712 5291 4728
rect 5225 4648 5226 4712
rect 5290 4648 5291 4712
rect 5225 4632 5291 4648
rect 5225 4568 5226 4632
rect 5290 4568 5291 4632
rect 5225 4552 5291 4568
rect 5225 4488 5226 4552
rect 5290 4488 5291 4552
rect 5225 4472 5291 4488
rect 5225 4408 5226 4472
rect 5290 4408 5291 4472
rect 5225 4392 5291 4408
rect 5225 4328 5226 4392
rect 5290 4328 5291 4392
rect 5225 4312 5291 4328
rect 5225 4248 5226 4312
rect 5290 4248 5291 4312
rect 5225 4232 5291 4248
rect 5225 4168 5226 4232
rect 5290 4168 5291 4232
rect 5225 4152 5291 4168
rect 5225 4088 5226 4152
rect 5290 4088 5291 4152
rect 5225 3934 5291 4088
rect 2801 3932 5291 3934
rect 2801 3868 2905 3932
rect 2969 3868 2985 3932
rect 3049 3868 3065 3932
rect 3129 3868 3145 3932
rect 3209 3868 3225 3932
rect 3289 3868 3305 3932
rect 3369 3868 3511 3932
rect 3575 3868 3591 3932
rect 3655 3868 3671 3932
rect 3735 3868 3751 3932
rect 3815 3868 3831 3932
rect 3895 3868 3911 3932
rect 3975 3868 4117 3932
rect 4181 3868 4197 3932
rect 4261 3868 4277 3932
rect 4341 3868 4357 3932
rect 4421 3868 4437 3932
rect 4501 3868 4517 3932
rect 4581 3868 4723 3932
rect 4787 3868 4803 3932
rect 4867 3868 4883 3932
rect 4947 3868 4963 3932
rect 5027 3868 5043 3932
rect 5107 3868 5123 3932
rect 5187 3868 5291 3932
rect 2801 3866 5291 3868
rect 2801 3712 2867 3866
rect 2801 3648 2802 3712
rect 2866 3648 2867 3712
rect 2801 3632 2867 3648
rect 2801 3568 2802 3632
rect 2866 3568 2867 3632
rect 2801 3552 2867 3568
rect 2801 3488 2802 3552
rect 2866 3488 2867 3552
rect 2801 3472 2867 3488
rect 2801 3408 2802 3472
rect 2866 3408 2867 3472
rect 2801 3392 2867 3408
rect 2801 3328 2802 3392
rect 2866 3328 2867 3392
rect 2801 3312 2867 3328
rect 2801 3248 2802 3312
rect 2866 3248 2867 3312
rect 2801 3232 2867 3248
rect 2801 3168 2802 3232
rect 2866 3168 2867 3232
rect 2801 3152 2867 3168
rect 2801 3088 2802 3152
rect 2866 3088 2867 3152
rect 2801 3077 2806 3088
rect 2862 3077 2867 3088
rect 2801 3072 2867 3077
rect 2801 3008 2802 3072
rect 2866 3008 2867 3072
rect 2801 2992 2867 3008
rect 2801 2928 2802 2992
rect 2866 2928 2867 2992
rect 2801 2838 2867 2928
rect 2927 2774 2987 3804
rect 3047 2834 3107 3866
rect 3167 2774 3227 3804
rect 3287 2834 3347 3866
rect 3407 3712 3473 3866
rect 3407 3648 3408 3712
rect 3472 3648 3473 3712
rect 3407 3632 3473 3648
rect 3407 3568 3408 3632
rect 3472 3568 3473 3632
rect 3407 3552 3473 3568
rect 3407 3488 3408 3552
rect 3472 3488 3473 3552
rect 3407 3472 3473 3488
rect 3407 3408 3408 3472
rect 3472 3408 3473 3472
rect 3407 3392 3473 3408
rect 3407 3328 3408 3392
rect 3472 3328 3473 3392
rect 3407 3312 3473 3328
rect 3407 3248 3408 3312
rect 3472 3248 3473 3312
rect 3407 3232 3473 3248
rect 3407 3168 3408 3232
rect 3472 3168 3473 3232
rect 3407 3152 3473 3168
rect 3407 3088 3408 3152
rect 3472 3088 3473 3152
rect 3407 3072 3473 3088
rect 3407 3008 3408 3072
rect 3472 3008 3473 3072
rect 3407 2992 3473 3008
rect 3407 2928 3408 2992
rect 3472 2928 3473 2992
rect 3407 2838 3473 2928
rect 3533 2774 3593 3804
rect 3653 2834 3713 3866
rect 3773 2774 3833 3804
rect 3893 2834 3953 3866
rect 4013 3712 4079 3866
rect 4013 3648 4014 3712
rect 4078 3648 4079 3712
rect 4013 3632 4079 3648
rect 4013 3568 4014 3632
rect 4078 3568 4079 3632
rect 4013 3552 4079 3568
rect 4013 3488 4014 3552
rect 4078 3488 4079 3552
rect 4013 3472 4079 3488
rect 4013 3408 4014 3472
rect 4078 3408 4079 3472
rect 4013 3392 4079 3408
rect 4013 3328 4014 3392
rect 4078 3328 4079 3392
rect 4013 3312 4079 3328
rect 4013 3248 4014 3312
rect 4078 3248 4079 3312
rect 4013 3232 4079 3248
rect 4013 3168 4014 3232
rect 4078 3168 4079 3232
rect 4013 3152 4079 3168
rect 4013 3088 4014 3152
rect 4078 3088 4079 3152
rect 4013 3072 4079 3088
rect 4013 3008 4014 3072
rect 4078 3008 4079 3072
rect 4013 2992 4079 3008
rect 4013 2928 4014 2992
rect 4078 2928 4079 2992
rect 4013 2838 4079 2928
rect 4139 2774 4199 3804
rect 4259 2834 4319 3866
rect 4379 2774 4439 3804
rect 4499 2834 4559 3866
rect 4619 3712 4685 3866
rect 4619 3648 4620 3712
rect 4684 3648 4685 3712
rect 4619 3632 4685 3648
rect 4619 3568 4620 3632
rect 4684 3568 4685 3632
rect 4619 3552 4685 3568
rect 4619 3488 4620 3552
rect 4684 3488 4685 3552
rect 4619 3472 4685 3488
rect 4619 3408 4620 3472
rect 4684 3408 4685 3472
rect 4619 3392 4685 3408
rect 4619 3328 4620 3392
rect 4684 3328 4685 3392
rect 4619 3312 4685 3328
rect 4619 3248 4620 3312
rect 4684 3248 4685 3312
rect 4619 3232 4685 3248
rect 4619 3168 4620 3232
rect 4684 3168 4685 3232
rect 4619 3152 4685 3168
rect 4619 3088 4620 3152
rect 4684 3088 4685 3152
rect 4619 3072 4685 3088
rect 4619 3008 4620 3072
rect 4684 3008 4685 3072
rect 4619 2992 4685 3008
rect 4619 2928 4620 2992
rect 4684 2928 4685 2992
rect 4619 2838 4685 2928
rect 4745 2774 4805 3804
rect 4865 2834 4925 3866
rect 4985 2774 5045 3804
rect 5105 2834 5165 3866
rect 5225 3712 5291 3866
rect 5225 3648 5226 3712
rect 5290 3648 5291 3712
rect 5225 3632 5291 3648
rect 5225 3568 5226 3632
rect 5290 3568 5291 3632
rect 5225 3552 5291 3568
rect 5225 3488 5226 3552
rect 5290 3488 5291 3552
rect 5225 3472 5291 3488
rect 5225 3408 5226 3472
rect 5290 3408 5291 3472
rect 5225 3392 5291 3408
rect 5225 3328 5226 3392
rect 5290 3328 5291 3392
rect 5225 3312 5291 3328
rect 5225 3248 5226 3312
rect 5290 3248 5291 3312
rect 5225 3232 5291 3248
rect 5225 3168 5226 3232
rect 5290 3168 5291 3232
rect 5225 3152 5291 3168
rect 5225 3088 5226 3152
rect 5290 3088 5291 3152
rect 5225 3072 5291 3088
rect 5225 3008 5226 3072
rect 5290 3008 5291 3072
rect 5225 2992 5291 3008
rect 5225 2928 5226 2992
rect 5290 2928 5291 2992
rect 5225 2838 5291 2928
rect 5352 4872 5418 4962
rect 5352 4808 5353 4872
rect 5417 4808 5418 4872
rect 5352 4792 5418 4808
rect 5352 4728 5353 4792
rect 5417 4728 5418 4792
rect 5352 4712 5418 4728
rect 5352 4648 5353 4712
rect 5417 4648 5418 4712
rect 5352 4632 5418 4648
rect 5352 4568 5353 4632
rect 5417 4568 5418 4632
rect 5352 4552 5418 4568
rect 5352 4488 5353 4552
rect 5417 4488 5418 4552
rect 5352 4472 5418 4488
rect 5352 4408 5353 4472
rect 5417 4408 5418 4472
rect 5352 4392 5418 4408
rect 5352 4328 5353 4392
rect 5417 4328 5418 4392
rect 5352 4312 5418 4328
rect 5352 4248 5353 4312
rect 5417 4248 5418 4312
rect 5352 4232 5418 4248
rect 5352 4168 5353 4232
rect 5417 4168 5418 4232
rect 5352 4152 5418 4168
rect 5352 4088 5353 4152
rect 5417 4088 5418 4152
rect 5352 3934 5418 4088
rect 5478 3934 5538 4966
rect 5598 3996 5658 5026
rect 5718 3934 5778 4966
rect 5838 3996 5898 5026
rect 5958 4872 6024 4962
rect 5958 4808 5959 4872
rect 6023 4808 6024 4872
rect 5958 4792 6024 4808
rect 5958 4728 5959 4792
rect 6023 4728 6024 4792
rect 5958 4712 6024 4728
rect 5958 4648 5959 4712
rect 6023 4648 6024 4712
rect 5958 4632 6024 4648
rect 5958 4568 5959 4632
rect 6023 4568 6024 4632
rect 5958 4552 6024 4568
rect 5958 4488 5959 4552
rect 6023 4488 6024 4552
rect 5958 4472 6024 4488
rect 5958 4408 5959 4472
rect 6023 4408 6024 4472
rect 5958 4392 6024 4408
rect 5958 4328 5959 4392
rect 6023 4328 6024 4392
rect 5958 4312 6024 4328
rect 5958 4248 5959 4312
rect 6023 4248 6024 4312
rect 5958 4232 6024 4248
rect 5958 4168 5959 4232
rect 6023 4168 6024 4232
rect 5958 4152 6024 4168
rect 5958 4088 5959 4152
rect 6023 4088 6024 4152
rect 5958 3934 6024 4088
rect 6084 3934 6144 4966
rect 6204 3996 6264 5026
rect 6324 3934 6384 4966
rect 6444 3996 6504 5026
rect 6564 4872 6630 4962
rect 6564 4808 6565 4872
rect 6629 4808 6630 4872
rect 6564 4792 6630 4808
rect 6564 4728 6565 4792
rect 6629 4728 6630 4792
rect 6564 4712 6630 4728
rect 6564 4648 6565 4712
rect 6629 4648 6630 4712
rect 6564 4632 6630 4648
rect 6564 4568 6565 4632
rect 6629 4568 6630 4632
rect 6564 4552 6630 4568
rect 6564 4488 6565 4552
rect 6629 4488 6630 4552
rect 6564 4472 6630 4488
rect 6564 4408 6565 4472
rect 6629 4408 6630 4472
rect 6564 4392 6630 4408
rect 6564 4328 6565 4392
rect 6629 4328 6630 4392
rect 6564 4312 6630 4328
rect 6564 4248 6565 4312
rect 6629 4248 6630 4312
rect 6564 4232 6630 4248
rect 6564 4168 6565 4232
rect 6629 4168 6630 4232
rect 6564 4152 6630 4168
rect 6564 4088 6565 4152
rect 6629 4088 6630 4152
rect 6564 3934 6630 4088
rect 6690 3934 6750 4966
rect 6810 3996 6870 5026
rect 6930 3934 6990 4966
rect 7050 3996 7110 5026
rect 7170 4872 7236 4962
rect 7170 4808 7171 4872
rect 7235 4808 7236 4872
rect 7170 4792 7236 4808
rect 7170 4728 7171 4792
rect 7235 4728 7236 4792
rect 7170 4712 7236 4728
rect 7170 4648 7171 4712
rect 7235 4648 7236 4712
rect 7170 4632 7236 4648
rect 7170 4568 7171 4632
rect 7235 4568 7236 4632
rect 7170 4552 7236 4568
rect 7170 4488 7171 4552
rect 7235 4488 7236 4552
rect 7170 4472 7236 4488
rect 7170 4408 7171 4472
rect 7235 4408 7236 4472
rect 7170 4392 7236 4408
rect 7170 4328 7171 4392
rect 7235 4328 7236 4392
rect 7170 4312 7236 4328
rect 7170 4248 7171 4312
rect 7235 4248 7236 4312
rect 7170 4232 7236 4248
rect 7170 4168 7171 4232
rect 7235 4168 7236 4232
rect 7170 4152 7236 4168
rect 7170 4088 7171 4152
rect 7235 4088 7236 4152
rect 7170 3934 7236 4088
rect 7296 3934 7356 4966
rect 7416 3996 7476 5026
rect 7536 3934 7596 4966
rect 7656 3996 7716 5026
rect 7776 4872 7842 4962
rect 7776 4808 7777 4872
rect 7841 4808 7842 4872
rect 7776 4792 7842 4808
rect 7776 4728 7777 4792
rect 7841 4728 7842 4792
rect 7776 4712 7842 4728
rect 7776 4648 7777 4712
rect 7841 4648 7842 4712
rect 7776 4632 7842 4648
rect 7776 4568 7777 4632
rect 7841 4568 7842 4632
rect 7776 4552 7842 4568
rect 7776 4488 7777 4552
rect 7841 4488 7842 4552
rect 7776 4472 7842 4488
rect 7776 4408 7777 4472
rect 7841 4408 7842 4472
rect 7776 4392 7842 4408
rect 7776 4328 7777 4392
rect 7841 4328 7842 4392
rect 7776 4312 7842 4328
rect 7776 4248 7777 4312
rect 7841 4248 7842 4312
rect 7776 4232 7842 4248
rect 7776 4168 7777 4232
rect 7841 4168 7842 4232
rect 7776 4152 7842 4168
rect 7776 4088 7777 4152
rect 7841 4088 7842 4152
rect 7776 3934 7842 4088
rect 7902 3934 7962 4966
rect 8022 3996 8082 5026
rect 8142 3934 8202 4966
rect 8262 3996 8322 5026
rect 8382 4872 8448 4962
rect 8382 4808 8383 4872
rect 8447 4808 8448 4872
rect 8382 4792 8448 4808
rect 8382 4728 8383 4792
rect 8447 4728 8448 4792
rect 8382 4712 8448 4728
rect 8382 4648 8383 4712
rect 8447 4648 8448 4712
rect 8382 4632 8448 4648
rect 8382 4568 8383 4632
rect 8447 4568 8448 4632
rect 8382 4552 8448 4568
rect 8382 4488 8383 4552
rect 8447 4488 8448 4552
rect 8382 4472 8448 4488
rect 8382 4408 8383 4472
rect 8447 4408 8448 4472
rect 8382 4392 8448 4408
rect 8382 4328 8383 4392
rect 8447 4328 8448 4392
rect 8382 4312 8448 4328
rect 8382 4248 8383 4312
rect 8447 4248 8448 4312
rect 8382 4232 8448 4248
rect 8382 4168 8383 4232
rect 8447 4168 8448 4232
rect 8382 4152 8448 4168
rect 8382 4088 8383 4152
rect 8447 4088 8448 4152
rect 8382 3934 8448 4088
rect 8508 3934 8568 4966
rect 8628 3996 8688 5026
rect 8748 3934 8808 4966
rect 8868 3996 8928 5026
rect 8988 4872 9054 4962
rect 8988 4808 8989 4872
rect 9053 4808 9054 4872
rect 8988 4792 9054 4808
rect 8988 4728 8989 4792
rect 9053 4728 9054 4792
rect 8988 4712 9054 4728
rect 8988 4648 8989 4712
rect 9053 4648 9054 4712
rect 8988 4632 9054 4648
rect 8988 4568 8989 4632
rect 9053 4568 9054 4632
rect 8988 4552 9054 4568
rect 8988 4488 8989 4552
rect 9053 4488 9054 4552
rect 8988 4472 9054 4488
rect 8988 4408 8989 4472
rect 9053 4408 9054 4472
rect 8988 4392 9054 4408
rect 8988 4328 8989 4392
rect 9053 4328 9054 4392
rect 8988 4312 9054 4328
rect 8988 4248 8989 4312
rect 9053 4248 9054 4312
rect 8988 4232 9054 4248
rect 8988 4168 8989 4232
rect 9053 4168 9054 4232
rect 8988 4152 9054 4168
rect 8988 4088 8989 4152
rect 9053 4088 9054 4152
rect 8988 3934 9054 4088
rect 9114 3934 9174 4966
rect 9234 3996 9294 5026
rect 9354 3934 9414 4966
rect 9474 3996 9534 5026
rect 9594 4872 9660 4962
rect 9594 4808 9595 4872
rect 9659 4808 9660 4872
rect 9594 4792 9660 4808
rect 9594 4728 9595 4792
rect 9659 4728 9660 4792
rect 9594 4712 9660 4728
rect 9594 4648 9595 4712
rect 9659 4648 9660 4712
rect 9594 4632 9660 4648
rect 9594 4568 9595 4632
rect 9659 4568 9660 4632
rect 9594 4552 9660 4568
rect 9594 4488 9595 4552
rect 9659 4488 9660 4552
rect 9594 4472 9660 4488
rect 9594 4408 9595 4472
rect 9659 4408 9660 4472
rect 9594 4392 9660 4408
rect 9594 4328 9595 4392
rect 9659 4328 9660 4392
rect 9594 4312 9660 4328
rect 9594 4248 9595 4312
rect 9659 4248 9660 4312
rect 9594 4232 9660 4248
rect 9594 4168 9595 4232
rect 9659 4168 9660 4232
rect 9594 4152 9660 4168
rect 9594 4088 9595 4152
rect 9659 4088 9660 4152
rect 9594 3934 9660 4088
rect 9720 3934 9780 4966
rect 9840 3996 9900 5026
rect 9960 3934 10020 4966
rect 10080 3996 10140 5026
rect 10200 4872 10266 4962
rect 10200 4808 10201 4872
rect 10265 4808 10266 4872
rect 10200 4792 10266 4808
rect 10200 4728 10201 4792
rect 10265 4728 10266 4792
rect 10200 4712 10266 4728
rect 10200 4648 10201 4712
rect 10265 4648 10266 4712
rect 10200 4632 10266 4648
rect 10200 4568 10201 4632
rect 10265 4568 10266 4632
rect 10200 4552 10266 4568
rect 10200 4488 10201 4552
rect 10265 4488 10266 4552
rect 10200 4472 10266 4488
rect 10200 4408 10201 4472
rect 10265 4408 10266 4472
rect 10200 4392 10266 4408
rect 10200 4328 10201 4392
rect 10265 4328 10266 4392
rect 10200 4312 10266 4328
rect 10200 4248 10201 4312
rect 10265 4248 10266 4312
rect 10200 4232 10266 4248
rect 10200 4168 10201 4232
rect 10265 4168 10266 4232
rect 10200 4152 10266 4168
rect 10200 4088 10201 4152
rect 10265 4088 10266 4152
rect 10200 3934 10266 4088
rect 5352 3932 10266 3934
rect 5352 3868 5456 3932
rect 5520 3868 5536 3932
rect 5600 3868 5616 3932
rect 5680 3868 5696 3932
rect 5760 3868 5776 3932
rect 5840 3868 5856 3932
rect 5920 3868 6062 3932
rect 6126 3868 6142 3932
rect 6206 3868 6222 3932
rect 6286 3868 6302 3932
rect 6366 3868 6382 3932
rect 6446 3868 6462 3932
rect 6526 3868 6668 3932
rect 6732 3868 6748 3932
rect 6812 3868 6828 3932
rect 6892 3868 6908 3932
rect 6972 3868 6988 3932
rect 7052 3868 7068 3932
rect 7132 3868 7274 3932
rect 7338 3868 7354 3932
rect 7418 3868 7434 3932
rect 7498 3868 7514 3932
rect 7578 3868 7594 3932
rect 7658 3868 7674 3932
rect 7738 3868 7880 3932
rect 7944 3868 7960 3932
rect 8024 3868 8040 3932
rect 8104 3868 8120 3932
rect 8184 3868 8200 3932
rect 8264 3868 8280 3932
rect 8344 3868 8486 3932
rect 8550 3868 8566 3932
rect 8630 3868 8646 3932
rect 8710 3868 8726 3932
rect 8790 3868 8806 3932
rect 8870 3868 8886 3932
rect 8950 3868 9092 3932
rect 9156 3868 9172 3932
rect 9236 3868 9252 3932
rect 9316 3868 9332 3932
rect 9396 3868 9412 3932
rect 9476 3868 9492 3932
rect 9556 3868 9698 3932
rect 9762 3868 9778 3932
rect 9842 3868 9858 3932
rect 9922 3868 9938 3932
rect 10002 3868 10018 3932
rect 10082 3868 10098 3932
rect 10162 3868 10266 3932
rect 5352 3866 10266 3868
rect 5352 3712 5418 3866
rect 5352 3648 5353 3712
rect 5417 3648 5418 3712
rect 5352 3632 5418 3648
rect 5352 3568 5353 3632
rect 5417 3568 5418 3632
rect 5352 3552 5418 3568
rect 5352 3488 5353 3552
rect 5417 3488 5418 3552
rect 5352 3472 5418 3488
rect 5352 3408 5353 3472
rect 5417 3408 5418 3472
rect 5352 3392 5418 3408
rect 5352 3328 5353 3392
rect 5417 3328 5418 3392
rect 5352 3312 5418 3328
rect 5352 3248 5353 3312
rect 5417 3248 5418 3312
rect 5352 3232 5418 3248
rect 5352 3168 5353 3232
rect 5417 3168 5418 3232
rect 5352 3165 5418 3168
rect 5352 3152 5357 3165
rect 5413 3152 5418 3165
rect 5352 3088 5353 3152
rect 5417 3088 5418 3152
rect 5352 3072 5418 3088
rect 5352 3008 5353 3072
rect 5417 3008 5418 3072
rect 5352 2992 5418 3008
rect 5352 2928 5353 2992
rect 5417 2928 5418 2992
rect 5352 2838 5418 2928
rect 5478 2774 5538 3804
rect 5598 2834 5658 3866
rect 5718 2774 5778 3804
rect 5838 2834 5898 3866
rect 5958 3712 6024 3866
rect 5958 3648 5959 3712
rect 6023 3648 6024 3712
rect 5958 3632 6024 3648
rect 5958 3568 5959 3632
rect 6023 3568 6024 3632
rect 5958 3552 6024 3568
rect 5958 3488 5959 3552
rect 6023 3488 6024 3552
rect 5958 3472 6024 3488
rect 5958 3408 5959 3472
rect 6023 3408 6024 3472
rect 5958 3392 6024 3408
rect 5958 3328 5959 3392
rect 6023 3328 6024 3392
rect 5958 3312 6024 3328
rect 5958 3248 5959 3312
rect 6023 3248 6024 3312
rect 5958 3232 6024 3248
rect 5958 3168 5959 3232
rect 6023 3168 6024 3232
rect 5958 3152 6024 3168
rect 5958 3088 5959 3152
rect 6023 3088 6024 3152
rect 5958 3072 6024 3088
rect 5958 3008 5959 3072
rect 6023 3008 6024 3072
rect 5958 2992 6024 3008
rect 5958 2928 5959 2992
rect 6023 2928 6024 2992
rect 5958 2838 6024 2928
rect 6084 2774 6144 3804
rect 6204 2834 6264 3866
rect 6324 2774 6384 3804
rect 6444 2834 6504 3866
rect 6564 3712 6630 3866
rect 6564 3648 6565 3712
rect 6629 3648 6630 3712
rect 6564 3632 6630 3648
rect 6564 3568 6565 3632
rect 6629 3568 6630 3632
rect 6564 3552 6630 3568
rect 6564 3488 6565 3552
rect 6629 3488 6630 3552
rect 6564 3472 6630 3488
rect 6564 3408 6565 3472
rect 6629 3408 6630 3472
rect 6564 3392 6630 3408
rect 6564 3328 6565 3392
rect 6629 3328 6630 3392
rect 6564 3312 6630 3328
rect 6564 3248 6565 3312
rect 6629 3248 6630 3312
rect 6564 3232 6630 3248
rect 6564 3168 6565 3232
rect 6629 3168 6630 3232
rect 6564 3152 6630 3168
rect 6564 3088 6565 3152
rect 6629 3088 6630 3152
rect 6564 3072 6630 3088
rect 6564 3008 6565 3072
rect 6629 3008 6630 3072
rect 6564 2992 6630 3008
rect 6564 2928 6565 2992
rect 6629 2928 6630 2992
rect 6564 2838 6630 2928
rect 6690 2774 6750 3804
rect 6810 2834 6870 3866
rect 6930 2774 6990 3804
rect 7050 2834 7110 3866
rect 7170 3712 7236 3866
rect 7170 3648 7171 3712
rect 7235 3648 7236 3712
rect 7170 3632 7236 3648
rect 7170 3568 7171 3632
rect 7235 3568 7236 3632
rect 7170 3552 7236 3568
rect 7170 3488 7171 3552
rect 7235 3488 7236 3552
rect 7170 3472 7236 3488
rect 7170 3408 7171 3472
rect 7235 3408 7236 3472
rect 7170 3392 7236 3408
rect 7170 3328 7171 3392
rect 7235 3328 7236 3392
rect 7170 3312 7236 3328
rect 7170 3248 7171 3312
rect 7235 3248 7236 3312
rect 7170 3232 7236 3248
rect 7170 3168 7171 3232
rect 7235 3168 7236 3232
rect 7170 3152 7236 3168
rect 7170 3088 7171 3152
rect 7235 3088 7236 3152
rect 7170 3072 7236 3088
rect 7170 3008 7171 3072
rect 7235 3008 7236 3072
rect 7170 2992 7236 3008
rect 7170 2928 7171 2992
rect 7235 2928 7236 2992
rect 7170 2838 7236 2928
rect 7296 2774 7356 3804
rect 7416 2834 7476 3866
rect 7536 2774 7596 3804
rect 7656 2834 7716 3866
rect 7776 3712 7842 3866
rect 7776 3648 7777 3712
rect 7841 3648 7842 3712
rect 7776 3632 7842 3648
rect 7776 3568 7777 3632
rect 7841 3568 7842 3632
rect 7776 3552 7842 3568
rect 7776 3488 7777 3552
rect 7841 3488 7842 3552
rect 7776 3472 7842 3488
rect 7776 3408 7777 3472
rect 7841 3408 7842 3472
rect 7776 3392 7842 3408
rect 7776 3328 7777 3392
rect 7841 3328 7842 3392
rect 7776 3312 7842 3328
rect 7776 3248 7777 3312
rect 7841 3248 7842 3312
rect 7776 3232 7842 3248
rect 7776 3168 7777 3232
rect 7841 3168 7842 3232
rect 7776 3152 7842 3168
rect 7776 3088 7777 3152
rect 7841 3088 7842 3152
rect 7776 3072 7842 3088
rect 7776 3008 7777 3072
rect 7841 3008 7842 3072
rect 7776 2992 7842 3008
rect 7776 2928 7777 2992
rect 7841 2928 7842 2992
rect 7776 2838 7842 2928
rect 7902 2774 7962 3804
rect 8022 2834 8082 3866
rect 8142 2774 8202 3804
rect 8262 2834 8322 3866
rect 8382 3712 8448 3866
rect 8382 3648 8383 3712
rect 8447 3648 8448 3712
rect 8382 3632 8448 3648
rect 8382 3568 8383 3632
rect 8447 3568 8448 3632
rect 8382 3552 8448 3568
rect 8382 3488 8383 3552
rect 8447 3488 8448 3552
rect 8382 3472 8448 3488
rect 8382 3408 8383 3472
rect 8447 3408 8448 3472
rect 8382 3392 8448 3408
rect 8382 3328 8383 3392
rect 8447 3328 8448 3392
rect 8382 3312 8448 3328
rect 8382 3248 8383 3312
rect 8447 3248 8448 3312
rect 8382 3232 8448 3248
rect 8382 3168 8383 3232
rect 8447 3168 8448 3232
rect 8382 3152 8448 3168
rect 8382 3088 8383 3152
rect 8447 3088 8448 3152
rect 8382 3072 8448 3088
rect 8382 3008 8383 3072
rect 8447 3008 8448 3072
rect 8382 2992 8448 3008
rect 8382 2928 8383 2992
rect 8447 2928 8448 2992
rect 8382 2838 8448 2928
rect 8508 2774 8568 3804
rect 8628 2834 8688 3866
rect 8748 2774 8808 3804
rect 8868 2834 8928 3866
rect 8988 3712 9054 3866
rect 8988 3648 8989 3712
rect 9053 3648 9054 3712
rect 8988 3632 9054 3648
rect 8988 3568 8989 3632
rect 9053 3568 9054 3632
rect 8988 3552 9054 3568
rect 8988 3488 8989 3552
rect 9053 3488 9054 3552
rect 8988 3472 9054 3488
rect 8988 3408 8989 3472
rect 9053 3408 9054 3472
rect 8988 3392 9054 3408
rect 8988 3328 8989 3392
rect 9053 3328 9054 3392
rect 8988 3312 9054 3328
rect 8988 3248 8989 3312
rect 9053 3248 9054 3312
rect 8988 3232 9054 3248
rect 8988 3168 8989 3232
rect 9053 3168 9054 3232
rect 8988 3152 9054 3168
rect 8988 3088 8989 3152
rect 9053 3088 9054 3152
rect 8988 3072 9054 3088
rect 8988 3008 8989 3072
rect 9053 3008 9054 3072
rect 8988 2992 9054 3008
rect 8988 2928 8989 2992
rect 9053 2928 9054 2992
rect 8988 2838 9054 2928
rect 9114 2774 9174 3804
rect 9234 2834 9294 3866
rect 9354 2774 9414 3804
rect 9474 2834 9534 3866
rect 9594 3712 9660 3866
rect 9594 3648 9595 3712
rect 9659 3648 9660 3712
rect 9594 3632 9660 3648
rect 9594 3568 9595 3632
rect 9659 3568 9660 3632
rect 9594 3552 9660 3568
rect 9594 3488 9595 3552
rect 9659 3488 9660 3552
rect 9594 3472 9660 3488
rect 9594 3408 9595 3472
rect 9659 3408 9660 3472
rect 9594 3392 9660 3408
rect 9594 3328 9595 3392
rect 9659 3328 9660 3392
rect 9594 3312 9660 3328
rect 9594 3248 9595 3312
rect 9659 3248 9660 3312
rect 9594 3232 9660 3248
rect 9594 3168 9595 3232
rect 9659 3168 9660 3232
rect 9594 3152 9660 3168
rect 9594 3088 9595 3152
rect 9659 3088 9660 3152
rect 9594 3072 9660 3088
rect 9594 3008 9595 3072
rect 9659 3008 9660 3072
rect 9594 2992 9660 3008
rect 9594 2928 9595 2992
rect 9659 2928 9660 2992
rect 9594 2838 9660 2928
rect 9720 2774 9780 3804
rect 9840 2834 9900 3866
rect 9960 2774 10020 3804
rect 10080 2834 10140 3866
rect 10200 3712 10266 3866
rect 10200 3648 10201 3712
rect 10265 3648 10266 3712
rect 10200 3632 10266 3648
rect 10200 3568 10201 3632
rect 10265 3568 10266 3632
rect 10200 3552 10266 3568
rect 10200 3488 10201 3552
rect 10265 3488 10266 3552
rect 10200 3472 10266 3488
rect 10200 3408 10201 3472
rect 10265 3408 10266 3472
rect 10200 3392 10266 3408
rect 10200 3328 10201 3392
rect 10265 3328 10266 3392
rect 10200 3312 10266 3328
rect 10200 3248 10201 3312
rect 10265 3248 10266 3312
rect 10200 3232 10266 3248
rect 10200 3168 10201 3232
rect 10265 3168 10266 3232
rect 10200 3152 10266 3168
rect 10200 3088 10201 3152
rect 10265 3088 10266 3152
rect 10200 3072 10266 3088
rect 10200 3008 10201 3072
rect 10265 3008 10266 3072
rect 10200 2992 10266 3008
rect 10200 2928 10201 2992
rect 10265 2928 10266 2992
rect 10200 2838 10266 2928
rect 10326 4872 10392 4962
rect 10326 4808 10327 4872
rect 10391 4808 10392 4872
rect 10326 4792 10392 4808
rect 10326 4728 10327 4792
rect 10391 4728 10392 4792
rect 10326 4712 10392 4728
rect 10326 4648 10327 4712
rect 10391 4648 10392 4712
rect 10326 4632 10392 4648
rect 10326 4568 10327 4632
rect 10391 4568 10392 4632
rect 10326 4552 10392 4568
rect 10326 4488 10327 4552
rect 10391 4488 10392 4552
rect 10326 4472 10392 4488
rect 10326 4408 10327 4472
rect 10391 4408 10392 4472
rect 10326 4392 10392 4408
rect 10326 4328 10327 4392
rect 10391 4328 10392 4392
rect 10326 4312 10392 4328
rect 10326 4248 10327 4312
rect 10391 4248 10392 4312
rect 10326 4232 10392 4248
rect 10326 4168 10327 4232
rect 10391 4168 10392 4232
rect 10326 4152 10392 4168
rect 10326 4088 10327 4152
rect 10391 4088 10392 4152
rect 10326 3934 10392 4088
rect 10452 3934 10512 4966
rect 10572 3996 10632 5026
rect 10692 3934 10752 4966
rect 10812 3996 10872 5026
rect 10932 4872 10998 4962
rect 10932 4808 10933 4872
rect 10997 4808 10998 4872
rect 10932 4792 10998 4808
rect 10932 4728 10933 4792
rect 10997 4728 10998 4792
rect 10932 4712 10998 4728
rect 10932 4648 10933 4712
rect 10997 4648 10998 4712
rect 10932 4632 10998 4648
rect 10932 4568 10933 4632
rect 10997 4568 10998 4632
rect 10932 4552 10998 4568
rect 10932 4488 10933 4552
rect 10997 4488 10998 4552
rect 10932 4472 10998 4488
rect 10932 4408 10933 4472
rect 10997 4408 10998 4472
rect 10932 4392 10998 4408
rect 10932 4328 10933 4392
rect 10997 4328 10998 4392
rect 10932 4312 10998 4328
rect 10932 4248 10933 4312
rect 10997 4248 10998 4312
rect 10932 4232 10998 4248
rect 10932 4168 10933 4232
rect 10997 4168 10998 4232
rect 10932 4152 10998 4168
rect 10932 4088 10933 4152
rect 10997 4088 10998 4152
rect 10932 3934 10998 4088
rect 11058 3934 11118 4966
rect 11178 3996 11238 5026
rect 11298 3934 11358 4966
rect 11418 3996 11478 5026
rect 11538 4872 11604 4962
rect 11538 4808 11539 4872
rect 11603 4808 11604 4872
rect 11538 4792 11604 4808
rect 11538 4728 11539 4792
rect 11603 4728 11604 4792
rect 11538 4712 11604 4728
rect 11538 4648 11539 4712
rect 11603 4648 11604 4712
rect 11538 4632 11604 4648
rect 11538 4568 11539 4632
rect 11603 4568 11604 4632
rect 11538 4552 11604 4568
rect 11538 4488 11539 4552
rect 11603 4488 11604 4552
rect 11538 4472 11604 4488
rect 11538 4408 11539 4472
rect 11603 4408 11604 4472
rect 11538 4392 11604 4408
rect 11538 4328 11539 4392
rect 11603 4328 11604 4392
rect 11538 4312 11604 4328
rect 11538 4248 11539 4312
rect 11603 4248 11604 4312
rect 11538 4232 11604 4248
rect 11538 4168 11539 4232
rect 11603 4168 11604 4232
rect 11538 4152 11604 4168
rect 11538 4088 11539 4152
rect 11603 4088 11604 4152
rect 11538 3934 11604 4088
rect 11664 3934 11724 4966
rect 11784 3996 11844 5026
rect 11904 3934 11964 4966
rect 12024 3996 12084 5026
rect 12144 4872 12210 4962
rect 12144 4808 12145 4872
rect 12209 4808 12210 4872
rect 12144 4792 12210 4808
rect 12144 4728 12145 4792
rect 12209 4728 12210 4792
rect 12144 4712 12210 4728
rect 12144 4648 12145 4712
rect 12209 4648 12210 4712
rect 12144 4632 12210 4648
rect 12144 4568 12145 4632
rect 12209 4568 12210 4632
rect 12144 4552 12210 4568
rect 12144 4488 12145 4552
rect 12209 4488 12210 4552
rect 12144 4472 12210 4488
rect 12144 4408 12145 4472
rect 12209 4408 12210 4472
rect 12144 4392 12210 4408
rect 12144 4328 12145 4392
rect 12209 4328 12210 4392
rect 12144 4312 12210 4328
rect 12144 4248 12145 4312
rect 12209 4248 12210 4312
rect 12144 4232 12210 4248
rect 12144 4168 12145 4232
rect 12209 4168 12210 4232
rect 12144 4152 12210 4168
rect 12144 4088 12145 4152
rect 12209 4088 12210 4152
rect 12144 3934 12210 4088
rect 12270 3934 12330 4966
rect 12390 3996 12450 5026
rect 12510 3934 12570 4966
rect 12630 3996 12690 5026
rect 12750 4872 12816 4962
rect 12750 4808 12751 4872
rect 12815 4808 12816 4872
rect 12750 4792 12816 4808
rect 12750 4728 12751 4792
rect 12815 4728 12816 4792
rect 12750 4712 12816 4728
rect 12750 4648 12751 4712
rect 12815 4648 12816 4712
rect 12750 4632 12816 4648
rect 12750 4568 12751 4632
rect 12815 4568 12816 4632
rect 12750 4552 12816 4568
rect 12750 4488 12751 4552
rect 12815 4488 12816 4552
rect 12750 4472 12816 4488
rect 12750 4408 12751 4472
rect 12815 4408 12816 4472
rect 12750 4392 12816 4408
rect 12750 4328 12751 4392
rect 12815 4328 12816 4392
rect 12750 4312 12816 4328
rect 12750 4248 12751 4312
rect 12815 4248 12816 4312
rect 12750 4232 12816 4248
rect 12750 4168 12751 4232
rect 12815 4168 12816 4232
rect 12750 4152 12816 4168
rect 12750 4088 12751 4152
rect 12815 4088 12816 4152
rect 12750 3934 12816 4088
rect 12876 3934 12936 4966
rect 12996 3996 13056 5026
rect 13116 3934 13176 4966
rect 13236 3996 13296 5026
rect 13356 4872 13422 4962
rect 13356 4808 13357 4872
rect 13421 4808 13422 4872
rect 13356 4792 13422 4808
rect 13356 4728 13357 4792
rect 13421 4728 13422 4792
rect 13356 4712 13422 4728
rect 13356 4648 13357 4712
rect 13421 4648 13422 4712
rect 13356 4632 13422 4648
rect 13356 4568 13357 4632
rect 13421 4568 13422 4632
rect 13356 4552 13422 4568
rect 13356 4488 13357 4552
rect 13421 4488 13422 4552
rect 13356 4472 13422 4488
rect 13356 4408 13357 4472
rect 13421 4408 13422 4472
rect 13356 4392 13422 4408
rect 13356 4328 13357 4392
rect 13421 4328 13422 4392
rect 13356 4312 13422 4328
rect 13356 4248 13357 4312
rect 13421 4248 13422 4312
rect 13356 4232 13422 4248
rect 13356 4168 13357 4232
rect 13421 4168 13422 4232
rect 13356 4152 13422 4168
rect 13356 4088 13357 4152
rect 13421 4088 13422 4152
rect 13356 3934 13422 4088
rect 13482 3934 13542 4966
rect 13602 3996 13662 5026
rect 13722 3934 13782 4966
rect 13842 3996 13902 5026
rect 13962 4872 14028 4962
rect 13962 4808 13963 4872
rect 14027 4808 14028 4872
rect 13962 4792 14028 4808
rect 13962 4728 13963 4792
rect 14027 4728 14028 4792
rect 13962 4712 14028 4728
rect 13962 4648 13963 4712
rect 14027 4648 14028 4712
rect 13962 4632 14028 4648
rect 13962 4568 13963 4632
rect 14027 4568 14028 4632
rect 13962 4552 14028 4568
rect 13962 4488 13963 4552
rect 14027 4488 14028 4552
rect 13962 4472 14028 4488
rect 13962 4408 13963 4472
rect 14027 4408 14028 4472
rect 13962 4392 14028 4408
rect 13962 4328 13963 4392
rect 14027 4328 14028 4392
rect 13962 4312 14028 4328
rect 13962 4248 13963 4312
rect 14027 4248 14028 4312
rect 13962 4232 14028 4248
rect 13962 4168 13963 4232
rect 14027 4168 14028 4232
rect 13962 4152 14028 4168
rect 13962 4088 13963 4152
rect 14027 4088 14028 4152
rect 13962 3934 14028 4088
rect 14088 3934 14148 4966
rect 14208 3996 14268 5026
rect 14328 3934 14388 4966
rect 14448 3996 14508 5026
rect 14568 4872 14634 4962
rect 14568 4808 14569 4872
rect 14633 4808 14634 4872
rect 14568 4792 14634 4808
rect 14568 4728 14569 4792
rect 14633 4728 14634 4792
rect 14568 4712 14634 4728
rect 14568 4648 14569 4712
rect 14633 4648 14634 4712
rect 14568 4632 14634 4648
rect 14568 4568 14569 4632
rect 14633 4568 14634 4632
rect 14568 4552 14634 4568
rect 14568 4488 14569 4552
rect 14633 4488 14634 4552
rect 14568 4472 14634 4488
rect 14568 4408 14569 4472
rect 14633 4408 14634 4472
rect 14568 4392 14634 4408
rect 14568 4328 14569 4392
rect 14633 4328 14634 4392
rect 14568 4312 14634 4328
rect 14568 4248 14569 4312
rect 14633 4248 14634 4312
rect 14568 4232 14634 4248
rect 14568 4168 14569 4232
rect 14633 4168 14634 4232
rect 14568 4152 14634 4168
rect 14568 4088 14569 4152
rect 14633 4088 14634 4152
rect 14568 3934 14634 4088
rect 14694 3934 14754 4966
rect 14814 3996 14874 5026
rect 14934 3934 14994 4966
rect 15054 3996 15114 5026
rect 15174 4872 15240 4962
rect 15174 4808 15175 4872
rect 15239 4808 15240 4872
rect 15174 4792 15240 4808
rect 15174 4728 15175 4792
rect 15239 4728 15240 4792
rect 15174 4712 15240 4728
rect 15174 4648 15175 4712
rect 15239 4648 15240 4712
rect 15174 4632 15240 4648
rect 15174 4568 15175 4632
rect 15239 4568 15240 4632
rect 15174 4552 15240 4568
rect 15174 4488 15175 4552
rect 15239 4488 15240 4552
rect 15174 4472 15240 4488
rect 15174 4408 15175 4472
rect 15239 4408 15240 4472
rect 15174 4392 15240 4408
rect 15174 4328 15175 4392
rect 15239 4328 15240 4392
rect 15174 4312 15240 4328
rect 15174 4248 15175 4312
rect 15239 4248 15240 4312
rect 15174 4232 15240 4248
rect 15174 4168 15175 4232
rect 15239 4168 15240 4232
rect 15174 4152 15240 4168
rect 15174 4088 15175 4152
rect 15239 4088 15240 4152
rect 15174 3934 15240 4088
rect 15300 3934 15360 4966
rect 15420 3996 15480 5026
rect 15540 3934 15600 4966
rect 15660 3996 15720 5026
rect 15780 4872 15846 4962
rect 15780 4808 15781 4872
rect 15845 4808 15846 4872
rect 15780 4792 15846 4808
rect 15780 4728 15781 4792
rect 15845 4728 15846 4792
rect 15780 4712 15846 4728
rect 15780 4648 15781 4712
rect 15845 4648 15846 4712
rect 15780 4632 15846 4648
rect 15780 4568 15781 4632
rect 15845 4568 15846 4632
rect 15780 4552 15846 4568
rect 15780 4488 15781 4552
rect 15845 4488 15846 4552
rect 15780 4472 15846 4488
rect 15780 4408 15781 4472
rect 15845 4408 15846 4472
rect 15780 4392 15846 4408
rect 15780 4328 15781 4392
rect 15845 4328 15846 4392
rect 15780 4312 15846 4328
rect 15780 4248 15781 4312
rect 15845 4248 15846 4312
rect 15780 4232 15846 4248
rect 15780 4168 15781 4232
rect 15845 4168 15846 4232
rect 15780 4152 15846 4168
rect 15780 4088 15781 4152
rect 15845 4088 15846 4152
rect 15780 3934 15846 4088
rect 15906 3934 15966 4966
rect 16026 3996 16086 5026
rect 16146 3934 16206 4966
rect 16266 3996 16326 5026
rect 16386 4872 16452 4962
rect 16386 4808 16387 4872
rect 16451 4808 16452 4872
rect 16386 4792 16452 4808
rect 16386 4728 16387 4792
rect 16451 4728 16452 4792
rect 16386 4712 16452 4728
rect 16386 4648 16387 4712
rect 16451 4648 16452 4712
rect 16386 4632 16452 4648
rect 16386 4568 16387 4632
rect 16451 4568 16452 4632
rect 16386 4552 16452 4568
rect 16386 4488 16387 4552
rect 16451 4488 16452 4552
rect 16386 4472 16452 4488
rect 16386 4408 16387 4472
rect 16451 4408 16452 4472
rect 16386 4392 16452 4408
rect 16386 4328 16387 4392
rect 16451 4328 16452 4392
rect 16386 4312 16452 4328
rect 16386 4248 16387 4312
rect 16451 4248 16452 4312
rect 16386 4232 16452 4248
rect 16386 4168 16387 4232
rect 16451 4168 16452 4232
rect 16386 4152 16452 4168
rect 16386 4088 16387 4152
rect 16451 4088 16452 4152
rect 16386 3934 16452 4088
rect 16512 3934 16572 4966
rect 16632 3996 16692 5026
rect 16752 3934 16812 4966
rect 16872 3996 16932 5026
rect 16992 4872 17058 4962
rect 16992 4808 16993 4872
rect 17057 4808 17058 4872
rect 16992 4792 17058 4808
rect 16992 4728 16993 4792
rect 17057 4728 17058 4792
rect 16992 4712 17058 4728
rect 16992 4648 16993 4712
rect 17057 4648 17058 4712
rect 16992 4632 17058 4648
rect 16992 4568 16993 4632
rect 17057 4568 17058 4632
rect 16992 4552 17058 4568
rect 16992 4488 16993 4552
rect 17057 4488 17058 4552
rect 16992 4472 17058 4488
rect 16992 4408 16993 4472
rect 17057 4408 17058 4472
rect 16992 4392 17058 4408
rect 16992 4328 16993 4392
rect 17057 4328 17058 4392
rect 16992 4312 17058 4328
rect 16992 4248 16993 4312
rect 17057 4248 17058 4312
rect 16992 4232 17058 4248
rect 16992 4168 16993 4232
rect 17057 4168 17058 4232
rect 16992 4152 17058 4168
rect 16992 4088 16993 4152
rect 17057 4088 17058 4152
rect 16992 3934 17058 4088
rect 17118 3934 17178 4966
rect 17238 3996 17298 5026
rect 17358 3934 17418 4966
rect 17478 3996 17538 5026
rect 17598 4872 17664 4962
rect 17598 4808 17599 4872
rect 17663 4808 17664 4872
rect 17598 4792 17664 4808
rect 17598 4728 17599 4792
rect 17663 4728 17664 4792
rect 17598 4712 17664 4728
rect 17598 4648 17599 4712
rect 17663 4648 17664 4712
rect 17598 4632 17664 4648
rect 17598 4568 17599 4632
rect 17663 4568 17664 4632
rect 17598 4552 17664 4568
rect 17598 4488 17599 4552
rect 17663 4488 17664 4552
rect 17598 4472 17664 4488
rect 17598 4408 17599 4472
rect 17663 4408 17664 4472
rect 17598 4392 17664 4408
rect 17598 4328 17599 4392
rect 17663 4328 17664 4392
rect 17598 4312 17664 4328
rect 17598 4248 17599 4312
rect 17663 4248 17664 4312
rect 17598 4232 17664 4248
rect 17598 4168 17599 4232
rect 17663 4168 17664 4232
rect 17598 4152 17664 4168
rect 17598 4088 17599 4152
rect 17663 4088 17664 4152
rect 17598 3934 17664 4088
rect 17724 3934 17784 4966
rect 17844 3996 17904 5026
rect 17964 3934 18024 4966
rect 18084 3996 18144 5026
rect 18204 4872 18270 4962
rect 18204 4808 18205 4872
rect 18269 4808 18270 4872
rect 18204 4792 18270 4808
rect 18204 4728 18205 4792
rect 18269 4728 18270 4792
rect 18204 4712 18270 4728
rect 18204 4648 18205 4712
rect 18269 4648 18270 4712
rect 18204 4632 18270 4648
rect 18204 4568 18205 4632
rect 18269 4568 18270 4632
rect 18204 4552 18270 4568
rect 18204 4488 18205 4552
rect 18269 4488 18270 4552
rect 18204 4472 18270 4488
rect 18204 4408 18205 4472
rect 18269 4408 18270 4472
rect 18204 4392 18270 4408
rect 18204 4328 18205 4392
rect 18269 4328 18270 4392
rect 18204 4312 18270 4328
rect 18204 4248 18205 4312
rect 18269 4248 18270 4312
rect 18204 4232 18270 4248
rect 18204 4168 18205 4232
rect 18269 4168 18270 4232
rect 18204 4152 18270 4168
rect 18204 4088 18205 4152
rect 18269 4088 18270 4152
rect 18204 3934 18270 4088
rect 18330 3934 18390 4966
rect 18450 3996 18510 5026
rect 18570 3934 18630 4966
rect 18690 3996 18750 5026
rect 18810 4872 18876 4962
rect 18810 4808 18811 4872
rect 18875 4808 18876 4872
rect 18810 4792 18876 4808
rect 18810 4728 18811 4792
rect 18875 4728 18876 4792
rect 18810 4712 18876 4728
rect 18810 4648 18811 4712
rect 18875 4648 18876 4712
rect 18810 4632 18876 4648
rect 18810 4568 18811 4632
rect 18875 4568 18876 4632
rect 18810 4552 18876 4568
rect 18810 4488 18811 4552
rect 18875 4488 18876 4552
rect 18810 4472 18876 4488
rect 18810 4408 18811 4472
rect 18875 4408 18876 4472
rect 18810 4392 18876 4408
rect 18810 4328 18811 4392
rect 18875 4328 18876 4392
rect 18810 4312 18876 4328
rect 18810 4248 18811 4312
rect 18875 4248 18876 4312
rect 18810 4232 18876 4248
rect 18810 4168 18811 4232
rect 18875 4168 18876 4232
rect 18810 4152 18876 4168
rect 18810 4088 18811 4152
rect 18875 4088 18876 4152
rect 18810 3934 18876 4088
rect 18936 3934 18996 4966
rect 19056 3996 19116 5026
rect 19176 3934 19236 4966
rect 19296 3996 19356 5026
rect 19416 4872 19482 4962
rect 19416 4808 19417 4872
rect 19481 4808 19482 4872
rect 19416 4792 19482 4808
rect 19416 4728 19417 4792
rect 19481 4728 19482 4792
rect 19416 4712 19482 4728
rect 19416 4648 19417 4712
rect 19481 4648 19482 4712
rect 19416 4632 19482 4648
rect 19416 4568 19417 4632
rect 19481 4568 19482 4632
rect 19416 4552 19482 4568
rect 19416 4488 19417 4552
rect 19481 4488 19482 4552
rect 19416 4472 19482 4488
rect 19416 4408 19417 4472
rect 19481 4408 19482 4472
rect 19416 4392 19482 4408
rect 19416 4328 19417 4392
rect 19481 4328 19482 4392
rect 19416 4312 19482 4328
rect 19416 4248 19417 4312
rect 19481 4248 19482 4312
rect 19416 4232 19482 4248
rect 19416 4168 19417 4232
rect 19481 4168 19482 4232
rect 19416 4152 19482 4168
rect 19416 4088 19417 4152
rect 19481 4088 19482 4152
rect 19416 3934 19482 4088
rect 19542 3934 19602 4966
rect 19662 3996 19722 5026
rect 19782 3934 19842 4966
rect 19902 3996 19962 5026
rect 20022 4872 20088 4962
rect 20022 4808 20023 4872
rect 20087 4808 20088 4872
rect 20022 4792 20088 4808
rect 20022 4728 20023 4792
rect 20087 4728 20088 4792
rect 20022 4712 20088 4728
rect 20022 4648 20023 4712
rect 20087 4648 20088 4712
rect 20022 4632 20088 4648
rect 20022 4568 20023 4632
rect 20087 4568 20088 4632
rect 20022 4552 20088 4568
rect 20022 4488 20023 4552
rect 20087 4488 20088 4552
rect 20022 4472 20088 4488
rect 20022 4408 20023 4472
rect 20087 4408 20088 4472
rect 20022 4392 20088 4408
rect 20022 4328 20023 4392
rect 20087 4328 20088 4392
rect 20022 4312 20088 4328
rect 20022 4248 20023 4312
rect 20087 4248 20088 4312
rect 20022 4232 20088 4248
rect 20022 4168 20023 4232
rect 20087 4168 20088 4232
rect 20022 4152 20088 4168
rect 20022 4088 20023 4152
rect 20087 4088 20088 4152
rect 20022 3934 20088 4088
rect 10326 3932 20088 3934
rect 10326 3868 10430 3932
rect 10494 3868 10510 3932
rect 10574 3868 10590 3932
rect 10654 3868 10670 3932
rect 10734 3868 10750 3932
rect 10814 3868 10830 3932
rect 10894 3868 11036 3932
rect 11100 3868 11116 3932
rect 11180 3868 11196 3932
rect 11260 3868 11276 3932
rect 11340 3868 11356 3932
rect 11420 3868 11436 3932
rect 11500 3868 11642 3932
rect 11706 3868 11722 3932
rect 11786 3868 11802 3932
rect 11866 3868 11882 3932
rect 11946 3868 11962 3932
rect 12026 3868 12042 3932
rect 12106 3868 12248 3932
rect 12312 3868 12328 3932
rect 12392 3868 12408 3932
rect 12472 3868 12488 3932
rect 12552 3868 12568 3932
rect 12632 3868 12648 3932
rect 12712 3868 12854 3932
rect 12918 3868 12934 3932
rect 12998 3868 13014 3932
rect 13078 3868 13094 3932
rect 13158 3868 13174 3932
rect 13238 3868 13254 3932
rect 13318 3868 13460 3932
rect 13524 3868 13540 3932
rect 13604 3868 13620 3932
rect 13684 3868 13700 3932
rect 13764 3868 13780 3932
rect 13844 3868 13860 3932
rect 13924 3868 14066 3932
rect 14130 3868 14146 3932
rect 14210 3868 14226 3932
rect 14290 3868 14306 3932
rect 14370 3868 14386 3932
rect 14450 3868 14466 3932
rect 14530 3868 14672 3932
rect 14736 3868 14752 3932
rect 14816 3868 14832 3932
rect 14896 3868 14912 3932
rect 14976 3868 14992 3932
rect 15056 3868 15072 3932
rect 15136 3868 15278 3932
rect 15342 3868 15358 3932
rect 15422 3868 15438 3932
rect 15502 3868 15518 3932
rect 15582 3868 15598 3932
rect 15662 3868 15678 3932
rect 15742 3868 15884 3932
rect 15948 3868 15964 3932
rect 16028 3868 16044 3932
rect 16108 3868 16124 3932
rect 16188 3868 16204 3932
rect 16268 3868 16284 3932
rect 16348 3868 16490 3932
rect 16554 3868 16570 3932
rect 16634 3868 16650 3932
rect 16714 3868 16730 3932
rect 16794 3868 16810 3932
rect 16874 3868 16890 3932
rect 16954 3868 17096 3932
rect 17160 3868 17176 3932
rect 17240 3868 17256 3932
rect 17320 3868 17336 3932
rect 17400 3868 17416 3932
rect 17480 3868 17496 3932
rect 17560 3868 17702 3932
rect 17766 3868 17782 3932
rect 17846 3868 17862 3932
rect 17926 3868 17942 3932
rect 18006 3868 18022 3932
rect 18086 3868 18102 3932
rect 18166 3868 18308 3932
rect 18372 3868 18388 3932
rect 18452 3868 18468 3932
rect 18532 3868 18548 3932
rect 18612 3868 18628 3932
rect 18692 3868 18708 3932
rect 18772 3868 18914 3932
rect 18978 3868 18994 3932
rect 19058 3868 19074 3932
rect 19138 3868 19154 3932
rect 19218 3868 19234 3932
rect 19298 3868 19314 3932
rect 19378 3868 19520 3932
rect 19584 3868 19600 3932
rect 19664 3868 19680 3932
rect 19744 3868 19760 3932
rect 19824 3868 19840 3932
rect 19904 3868 19920 3932
rect 19984 3868 20088 3932
rect 10326 3866 20088 3868
rect 10326 3712 10392 3866
rect 10326 3648 10327 3712
rect 10391 3648 10392 3712
rect 10326 3632 10392 3648
rect 10326 3568 10327 3632
rect 10391 3568 10392 3632
rect 10326 3552 10392 3568
rect 10326 3488 10327 3552
rect 10391 3488 10392 3552
rect 10326 3472 10392 3488
rect 10326 3408 10327 3472
rect 10391 3408 10392 3472
rect 10326 3392 10392 3408
rect 10326 3328 10327 3392
rect 10391 3328 10392 3392
rect 10326 3312 10392 3328
rect 10326 3248 10327 3312
rect 10391 3248 10392 3312
rect 10326 3232 10331 3248
rect 10387 3232 10392 3248
rect 10326 3168 10327 3232
rect 10391 3168 10392 3232
rect 10326 3152 10392 3168
rect 10326 3088 10327 3152
rect 10391 3088 10392 3152
rect 10326 3072 10392 3088
rect 10326 3008 10327 3072
rect 10391 3008 10392 3072
rect 10326 2992 10392 3008
rect 10326 2928 10327 2992
rect 10391 2928 10392 2992
rect 10326 2838 10392 2928
rect 10452 2774 10512 3804
rect 10572 2834 10632 3866
rect 10692 2774 10752 3804
rect 10812 2834 10872 3866
rect 10932 3712 10998 3866
rect 10932 3648 10933 3712
rect 10997 3648 10998 3712
rect 10932 3632 10998 3648
rect 10932 3568 10933 3632
rect 10997 3568 10998 3632
rect 10932 3552 10998 3568
rect 10932 3488 10933 3552
rect 10997 3488 10998 3552
rect 10932 3472 10998 3488
rect 10932 3408 10933 3472
rect 10997 3408 10998 3472
rect 10932 3392 10998 3408
rect 10932 3328 10933 3392
rect 10997 3328 10998 3392
rect 10932 3312 10998 3328
rect 10932 3248 10933 3312
rect 10997 3248 10998 3312
rect 10932 3232 10998 3248
rect 10932 3168 10933 3232
rect 10997 3168 10998 3232
rect 10932 3152 10998 3168
rect 10932 3088 10933 3152
rect 10997 3088 10998 3152
rect 10932 3072 10998 3088
rect 10932 3008 10933 3072
rect 10997 3008 10998 3072
rect 10932 2992 10998 3008
rect 10932 2928 10933 2992
rect 10997 2928 10998 2992
rect 10932 2838 10998 2928
rect 11058 2774 11118 3804
rect 11178 2834 11238 3866
rect 11298 2774 11358 3804
rect 11418 2834 11478 3866
rect 11538 3712 11604 3866
rect 11538 3648 11539 3712
rect 11603 3648 11604 3712
rect 11538 3632 11604 3648
rect 11538 3568 11539 3632
rect 11603 3568 11604 3632
rect 11538 3552 11604 3568
rect 11538 3488 11539 3552
rect 11603 3488 11604 3552
rect 11538 3472 11604 3488
rect 11538 3408 11539 3472
rect 11603 3408 11604 3472
rect 11538 3392 11604 3408
rect 11538 3328 11539 3392
rect 11603 3328 11604 3392
rect 11538 3312 11604 3328
rect 11538 3248 11539 3312
rect 11603 3248 11604 3312
rect 11538 3232 11604 3248
rect 11538 3168 11539 3232
rect 11603 3168 11604 3232
rect 11538 3152 11604 3168
rect 11538 3088 11539 3152
rect 11603 3088 11604 3152
rect 11538 3072 11604 3088
rect 11538 3008 11539 3072
rect 11603 3008 11604 3072
rect 11538 2992 11604 3008
rect 11538 2928 11539 2992
rect 11603 2928 11604 2992
rect 11538 2838 11604 2928
rect 11664 2774 11724 3804
rect 11784 2834 11844 3866
rect 11904 2774 11964 3804
rect 12024 2834 12084 3866
rect 12144 3712 12210 3866
rect 12144 3648 12145 3712
rect 12209 3648 12210 3712
rect 12144 3632 12210 3648
rect 12144 3568 12145 3632
rect 12209 3568 12210 3632
rect 12144 3552 12210 3568
rect 12144 3488 12145 3552
rect 12209 3488 12210 3552
rect 12144 3472 12210 3488
rect 12144 3408 12145 3472
rect 12209 3408 12210 3472
rect 12144 3392 12210 3408
rect 12144 3328 12145 3392
rect 12209 3328 12210 3392
rect 12144 3312 12210 3328
rect 12144 3248 12145 3312
rect 12209 3248 12210 3312
rect 12144 3232 12210 3248
rect 12144 3168 12145 3232
rect 12209 3168 12210 3232
rect 12144 3152 12210 3168
rect 12144 3088 12145 3152
rect 12209 3088 12210 3152
rect 12144 3072 12210 3088
rect 12144 3008 12145 3072
rect 12209 3008 12210 3072
rect 12144 2992 12210 3008
rect 12144 2928 12145 2992
rect 12209 2928 12210 2992
rect 12144 2838 12210 2928
rect 12270 2774 12330 3804
rect 12390 2834 12450 3866
rect 12510 2774 12570 3804
rect 12630 2834 12690 3866
rect 12750 3712 12816 3866
rect 12750 3648 12751 3712
rect 12815 3648 12816 3712
rect 12750 3632 12816 3648
rect 12750 3568 12751 3632
rect 12815 3568 12816 3632
rect 12750 3552 12816 3568
rect 12750 3488 12751 3552
rect 12815 3488 12816 3552
rect 12750 3472 12816 3488
rect 12750 3408 12751 3472
rect 12815 3408 12816 3472
rect 12750 3392 12816 3408
rect 12750 3328 12751 3392
rect 12815 3328 12816 3392
rect 12750 3312 12816 3328
rect 12750 3248 12751 3312
rect 12815 3248 12816 3312
rect 12750 3232 12816 3248
rect 12750 3168 12751 3232
rect 12815 3168 12816 3232
rect 12750 3152 12816 3168
rect 12750 3088 12751 3152
rect 12815 3088 12816 3152
rect 12750 3072 12816 3088
rect 12750 3008 12751 3072
rect 12815 3008 12816 3072
rect 12750 2992 12816 3008
rect 12750 2928 12751 2992
rect 12815 2928 12816 2992
rect 12750 2838 12816 2928
rect 12876 2774 12936 3804
rect 12996 2834 13056 3866
rect 13116 2774 13176 3804
rect 13236 2834 13296 3866
rect 13356 3712 13422 3866
rect 13356 3648 13357 3712
rect 13421 3648 13422 3712
rect 13356 3632 13422 3648
rect 13356 3568 13357 3632
rect 13421 3568 13422 3632
rect 13356 3552 13422 3568
rect 13356 3488 13357 3552
rect 13421 3488 13422 3552
rect 13356 3472 13422 3488
rect 13356 3408 13357 3472
rect 13421 3408 13422 3472
rect 13356 3392 13422 3408
rect 13356 3328 13357 3392
rect 13421 3328 13422 3392
rect 13356 3312 13422 3328
rect 13356 3248 13357 3312
rect 13421 3248 13422 3312
rect 13356 3232 13422 3248
rect 13356 3168 13357 3232
rect 13421 3168 13422 3232
rect 13356 3152 13422 3168
rect 13356 3088 13357 3152
rect 13421 3088 13422 3152
rect 13356 3072 13422 3088
rect 13356 3008 13357 3072
rect 13421 3008 13422 3072
rect 13356 2992 13422 3008
rect 13356 2928 13357 2992
rect 13421 2928 13422 2992
rect 13356 2838 13422 2928
rect 13482 2774 13542 3804
rect 13602 2834 13662 3866
rect 13722 2774 13782 3804
rect 13842 2834 13902 3866
rect 13962 3712 14028 3866
rect 13962 3648 13963 3712
rect 14027 3648 14028 3712
rect 13962 3632 14028 3648
rect 13962 3568 13963 3632
rect 14027 3568 14028 3632
rect 13962 3552 14028 3568
rect 13962 3488 13963 3552
rect 14027 3488 14028 3552
rect 13962 3472 14028 3488
rect 13962 3408 13963 3472
rect 14027 3408 14028 3472
rect 13962 3392 14028 3408
rect 13962 3328 13963 3392
rect 14027 3328 14028 3392
rect 13962 3312 14028 3328
rect 13962 3248 13963 3312
rect 14027 3248 14028 3312
rect 13962 3232 14028 3248
rect 13962 3168 13963 3232
rect 14027 3168 14028 3232
rect 13962 3152 14028 3168
rect 13962 3088 13963 3152
rect 14027 3088 14028 3152
rect 13962 3072 14028 3088
rect 13962 3008 13963 3072
rect 14027 3008 14028 3072
rect 13962 2992 14028 3008
rect 13962 2928 13963 2992
rect 14027 2928 14028 2992
rect 13962 2838 14028 2928
rect 14088 2774 14148 3804
rect 14208 2834 14268 3866
rect 14328 2774 14388 3804
rect 14448 2834 14508 3866
rect 14568 3712 14634 3866
rect 14568 3648 14569 3712
rect 14633 3648 14634 3712
rect 14568 3632 14634 3648
rect 14568 3568 14569 3632
rect 14633 3568 14634 3632
rect 14568 3552 14634 3568
rect 14568 3488 14569 3552
rect 14633 3488 14634 3552
rect 14568 3472 14634 3488
rect 14568 3408 14569 3472
rect 14633 3408 14634 3472
rect 14568 3392 14634 3408
rect 14568 3328 14569 3392
rect 14633 3328 14634 3392
rect 14568 3312 14634 3328
rect 14568 3248 14569 3312
rect 14633 3248 14634 3312
rect 14568 3232 14634 3248
rect 14568 3168 14569 3232
rect 14633 3168 14634 3232
rect 14568 3152 14634 3168
rect 14568 3088 14569 3152
rect 14633 3088 14634 3152
rect 14568 3072 14634 3088
rect 14568 3008 14569 3072
rect 14633 3008 14634 3072
rect 14568 2992 14634 3008
rect 14568 2928 14569 2992
rect 14633 2928 14634 2992
rect 14568 2838 14634 2928
rect 14694 2774 14754 3804
rect 14814 2834 14874 3866
rect 14934 2774 14994 3804
rect 15054 2834 15114 3866
rect 15174 3712 15240 3866
rect 15174 3648 15175 3712
rect 15239 3648 15240 3712
rect 15174 3632 15240 3648
rect 15174 3568 15175 3632
rect 15239 3568 15240 3632
rect 15174 3552 15240 3568
rect 15174 3488 15175 3552
rect 15239 3488 15240 3552
rect 15174 3472 15240 3488
rect 15174 3408 15175 3472
rect 15239 3408 15240 3472
rect 15174 3392 15240 3408
rect 15174 3328 15175 3392
rect 15239 3328 15240 3392
rect 15174 3312 15240 3328
rect 15174 3248 15175 3312
rect 15239 3248 15240 3312
rect 15174 3232 15240 3248
rect 15174 3168 15175 3232
rect 15239 3168 15240 3232
rect 15174 3152 15240 3168
rect 15174 3088 15175 3152
rect 15239 3088 15240 3152
rect 15174 3072 15240 3088
rect 15174 3008 15175 3072
rect 15239 3008 15240 3072
rect 15174 2992 15240 3008
rect 15174 2928 15175 2992
rect 15239 2928 15240 2992
rect 15174 2838 15240 2928
rect 15300 2774 15360 3804
rect 15420 2834 15480 3866
rect 15540 2774 15600 3804
rect 15660 2834 15720 3866
rect 15780 3712 15846 3866
rect 15780 3648 15781 3712
rect 15845 3648 15846 3712
rect 15780 3632 15846 3648
rect 15780 3568 15781 3632
rect 15845 3568 15846 3632
rect 15780 3552 15846 3568
rect 15780 3488 15781 3552
rect 15845 3488 15846 3552
rect 15780 3472 15846 3488
rect 15780 3408 15781 3472
rect 15845 3408 15846 3472
rect 15780 3392 15846 3408
rect 15780 3328 15781 3392
rect 15845 3328 15846 3392
rect 15780 3312 15846 3328
rect 15780 3248 15781 3312
rect 15845 3248 15846 3312
rect 15780 3232 15846 3248
rect 15780 3168 15781 3232
rect 15845 3168 15846 3232
rect 15780 3152 15846 3168
rect 15780 3088 15781 3152
rect 15845 3088 15846 3152
rect 15780 3072 15846 3088
rect 15780 3008 15781 3072
rect 15845 3008 15846 3072
rect 15780 2992 15846 3008
rect 15780 2928 15781 2992
rect 15845 2928 15846 2992
rect 15780 2838 15846 2928
rect 15906 2774 15966 3804
rect 16026 2834 16086 3866
rect 16146 2774 16206 3804
rect 16266 2834 16326 3866
rect 16386 3712 16452 3866
rect 16386 3648 16387 3712
rect 16451 3648 16452 3712
rect 16386 3632 16452 3648
rect 16386 3568 16387 3632
rect 16451 3568 16452 3632
rect 16386 3552 16452 3568
rect 16386 3488 16387 3552
rect 16451 3488 16452 3552
rect 16386 3472 16452 3488
rect 16386 3408 16387 3472
rect 16451 3408 16452 3472
rect 16386 3392 16452 3408
rect 16386 3328 16387 3392
rect 16451 3328 16452 3392
rect 16386 3312 16452 3328
rect 16386 3248 16387 3312
rect 16451 3248 16452 3312
rect 16386 3232 16452 3248
rect 16386 3168 16387 3232
rect 16451 3168 16452 3232
rect 16386 3152 16452 3168
rect 16386 3088 16387 3152
rect 16451 3088 16452 3152
rect 16386 3072 16452 3088
rect 16386 3008 16387 3072
rect 16451 3008 16452 3072
rect 16386 2992 16452 3008
rect 16386 2928 16387 2992
rect 16451 2928 16452 2992
rect 16386 2838 16452 2928
rect 16512 2774 16572 3804
rect 16632 2834 16692 3866
rect 16752 2774 16812 3804
rect 16872 2834 16932 3866
rect 16992 3712 17058 3866
rect 16992 3648 16993 3712
rect 17057 3648 17058 3712
rect 16992 3632 17058 3648
rect 16992 3568 16993 3632
rect 17057 3568 17058 3632
rect 16992 3552 17058 3568
rect 16992 3488 16993 3552
rect 17057 3488 17058 3552
rect 16992 3472 17058 3488
rect 16992 3408 16993 3472
rect 17057 3408 17058 3472
rect 16992 3392 17058 3408
rect 16992 3328 16993 3392
rect 17057 3328 17058 3392
rect 16992 3312 17058 3328
rect 16992 3248 16993 3312
rect 17057 3248 17058 3312
rect 16992 3232 17058 3248
rect 16992 3168 16993 3232
rect 17057 3168 17058 3232
rect 16992 3152 17058 3168
rect 16992 3088 16993 3152
rect 17057 3088 17058 3152
rect 16992 3072 17058 3088
rect 16992 3008 16993 3072
rect 17057 3008 17058 3072
rect 16992 2992 17058 3008
rect 16992 2928 16993 2992
rect 17057 2928 17058 2992
rect 16992 2838 17058 2928
rect 17118 2774 17178 3804
rect 17238 2834 17298 3866
rect 17358 2774 17418 3804
rect 17478 2834 17538 3866
rect 17598 3712 17664 3866
rect 17598 3648 17599 3712
rect 17663 3648 17664 3712
rect 17598 3632 17664 3648
rect 17598 3568 17599 3632
rect 17663 3568 17664 3632
rect 17598 3552 17664 3568
rect 17598 3488 17599 3552
rect 17663 3488 17664 3552
rect 17598 3472 17664 3488
rect 17598 3408 17599 3472
rect 17663 3408 17664 3472
rect 17598 3392 17664 3408
rect 17598 3328 17599 3392
rect 17663 3328 17664 3392
rect 17598 3312 17664 3328
rect 17598 3248 17599 3312
rect 17663 3248 17664 3312
rect 17598 3232 17664 3248
rect 17598 3168 17599 3232
rect 17663 3168 17664 3232
rect 17598 3152 17664 3168
rect 17598 3088 17599 3152
rect 17663 3088 17664 3152
rect 17598 3072 17664 3088
rect 17598 3008 17599 3072
rect 17663 3008 17664 3072
rect 17598 2992 17664 3008
rect 17598 2928 17599 2992
rect 17663 2928 17664 2992
rect 17598 2838 17664 2928
rect 17724 2774 17784 3804
rect 17844 2834 17904 3866
rect 17964 2774 18024 3804
rect 18084 2834 18144 3866
rect 18204 3712 18270 3866
rect 18204 3648 18205 3712
rect 18269 3648 18270 3712
rect 18204 3632 18270 3648
rect 18204 3568 18205 3632
rect 18269 3568 18270 3632
rect 18204 3552 18270 3568
rect 18204 3488 18205 3552
rect 18269 3488 18270 3552
rect 18204 3472 18270 3488
rect 18204 3408 18205 3472
rect 18269 3408 18270 3472
rect 18204 3392 18270 3408
rect 18204 3328 18205 3392
rect 18269 3328 18270 3392
rect 18204 3312 18270 3328
rect 18204 3248 18205 3312
rect 18269 3248 18270 3312
rect 18204 3232 18270 3248
rect 18204 3168 18205 3232
rect 18269 3168 18270 3232
rect 18204 3152 18270 3168
rect 18204 3088 18205 3152
rect 18269 3088 18270 3152
rect 18204 3072 18270 3088
rect 18204 3008 18205 3072
rect 18269 3008 18270 3072
rect 18204 2992 18270 3008
rect 18204 2928 18205 2992
rect 18269 2928 18270 2992
rect 18204 2838 18270 2928
rect 18330 2774 18390 3804
rect 18450 2834 18510 3866
rect 18570 2774 18630 3804
rect 18690 2834 18750 3866
rect 18810 3712 18876 3866
rect 18810 3648 18811 3712
rect 18875 3648 18876 3712
rect 18810 3632 18876 3648
rect 18810 3568 18811 3632
rect 18875 3568 18876 3632
rect 18810 3552 18876 3568
rect 18810 3488 18811 3552
rect 18875 3488 18876 3552
rect 18810 3472 18876 3488
rect 18810 3408 18811 3472
rect 18875 3408 18876 3472
rect 18810 3392 18876 3408
rect 18810 3328 18811 3392
rect 18875 3328 18876 3392
rect 18810 3312 18876 3328
rect 18810 3248 18811 3312
rect 18875 3248 18876 3312
rect 18810 3232 18876 3248
rect 18810 3168 18811 3232
rect 18875 3168 18876 3232
rect 18810 3152 18876 3168
rect 18810 3088 18811 3152
rect 18875 3088 18876 3152
rect 18810 3072 18876 3088
rect 18810 3008 18811 3072
rect 18875 3008 18876 3072
rect 18810 2992 18876 3008
rect 18810 2928 18811 2992
rect 18875 2928 18876 2992
rect 18810 2838 18876 2928
rect 18936 2774 18996 3804
rect 19056 2834 19116 3866
rect 19176 2774 19236 3804
rect 19296 2834 19356 3866
rect 19416 3712 19482 3866
rect 19416 3648 19417 3712
rect 19481 3648 19482 3712
rect 19416 3632 19482 3648
rect 19416 3568 19417 3632
rect 19481 3568 19482 3632
rect 19416 3552 19482 3568
rect 19416 3488 19417 3552
rect 19481 3488 19482 3552
rect 19416 3472 19482 3488
rect 19416 3408 19417 3472
rect 19481 3408 19482 3472
rect 19416 3392 19482 3408
rect 19416 3328 19417 3392
rect 19481 3328 19482 3392
rect 19416 3312 19482 3328
rect 19416 3248 19417 3312
rect 19481 3248 19482 3312
rect 19416 3232 19482 3248
rect 19416 3168 19417 3232
rect 19481 3168 19482 3232
rect 19416 3152 19482 3168
rect 19416 3088 19417 3152
rect 19481 3088 19482 3152
rect 19416 3072 19482 3088
rect 19416 3008 19417 3072
rect 19481 3008 19482 3072
rect 19416 2992 19482 3008
rect 19416 2928 19417 2992
rect 19481 2928 19482 2992
rect 19416 2838 19482 2928
rect 19542 2774 19602 3804
rect 19662 2834 19722 3866
rect 19782 2774 19842 3804
rect 19902 2834 19962 3866
rect 20022 3712 20088 3866
rect 20022 3648 20023 3712
rect 20087 3648 20088 3712
rect 20022 3632 20088 3648
rect 20022 3568 20023 3632
rect 20087 3568 20088 3632
rect 20022 3552 20088 3568
rect 20022 3488 20023 3552
rect 20087 3488 20088 3552
rect 20022 3472 20088 3488
rect 20022 3408 20023 3472
rect 20087 3408 20088 3472
rect 20022 3392 20088 3408
rect 20022 3328 20023 3392
rect 20087 3328 20088 3392
rect 20022 3312 20088 3328
rect 20022 3248 20023 3312
rect 20087 3248 20088 3312
rect 20022 3232 20088 3248
rect 20022 3168 20023 3232
rect 20087 3168 20088 3232
rect 20022 3152 20088 3168
rect 20022 3088 20023 3152
rect 20087 3088 20088 3152
rect 20022 3072 20088 3088
rect 20022 3008 20023 3072
rect 20087 3008 20088 3072
rect 20022 2992 20088 3008
rect 20022 2928 20023 2992
rect 20087 2928 20088 2992
rect 20022 2838 20088 2928
rect 20148 4872 20214 4962
rect 20148 4808 20149 4872
rect 20213 4808 20214 4872
rect 20148 4792 20214 4808
rect 20148 4728 20149 4792
rect 20213 4728 20214 4792
rect 20148 4712 20214 4728
rect 20148 4648 20149 4712
rect 20213 4648 20214 4712
rect 20148 4632 20214 4648
rect 20148 4568 20149 4632
rect 20213 4568 20214 4632
rect 20148 4552 20214 4568
rect 20148 4488 20149 4552
rect 20213 4488 20214 4552
rect 20148 4472 20214 4488
rect 20148 4408 20149 4472
rect 20213 4408 20214 4472
rect 20148 4392 20214 4408
rect 20148 4328 20149 4392
rect 20213 4328 20214 4392
rect 20148 4312 20214 4328
rect 20148 4248 20149 4312
rect 20213 4248 20214 4312
rect 20148 4232 20214 4248
rect 20148 4168 20149 4232
rect 20213 4168 20214 4232
rect 20148 4152 20214 4168
rect 20148 4088 20149 4152
rect 20213 4088 20214 4152
rect 20148 3934 20214 4088
rect 20274 3934 20334 4966
rect 20394 3996 20454 5026
rect 20514 3934 20574 4966
rect 20634 3996 20694 5026
rect 20754 4872 20820 4962
rect 20754 4808 20755 4872
rect 20819 4808 20820 4872
rect 20754 4792 20820 4808
rect 20754 4728 20755 4792
rect 20819 4728 20820 4792
rect 20754 4712 20820 4728
rect 20754 4648 20755 4712
rect 20819 4648 20820 4712
rect 20754 4632 20820 4648
rect 20754 4568 20755 4632
rect 20819 4568 20820 4632
rect 20754 4552 20820 4568
rect 20754 4488 20755 4552
rect 20819 4488 20820 4552
rect 20754 4472 20820 4488
rect 20754 4408 20755 4472
rect 20819 4408 20820 4472
rect 20754 4392 20820 4408
rect 20754 4328 20755 4392
rect 20819 4328 20820 4392
rect 20754 4312 20820 4328
rect 20754 4248 20755 4312
rect 20819 4248 20820 4312
rect 20754 4232 20820 4248
rect 20754 4168 20755 4232
rect 20819 4168 20820 4232
rect 20754 4152 20820 4168
rect 20754 4088 20755 4152
rect 20819 4088 20820 4152
rect 20754 3934 20820 4088
rect 20880 3934 20940 4966
rect 21000 3996 21060 5026
rect 21120 3934 21180 4966
rect 21240 3996 21300 5026
rect 21360 4872 21426 4962
rect 21360 4808 21361 4872
rect 21425 4808 21426 4872
rect 21360 4792 21426 4808
rect 21360 4728 21361 4792
rect 21425 4728 21426 4792
rect 21360 4712 21426 4728
rect 21360 4648 21361 4712
rect 21425 4648 21426 4712
rect 21360 4632 21426 4648
rect 21360 4568 21361 4632
rect 21425 4568 21426 4632
rect 21360 4552 21426 4568
rect 21360 4488 21361 4552
rect 21425 4488 21426 4552
rect 21360 4472 21426 4488
rect 21360 4408 21361 4472
rect 21425 4408 21426 4472
rect 21360 4392 21426 4408
rect 21360 4328 21361 4392
rect 21425 4328 21426 4392
rect 21360 4312 21426 4328
rect 21360 4248 21361 4312
rect 21425 4248 21426 4312
rect 21360 4232 21426 4248
rect 21360 4168 21361 4232
rect 21425 4168 21426 4232
rect 21360 4152 21426 4168
rect 21360 4088 21361 4152
rect 21425 4088 21426 4152
rect 21360 3934 21426 4088
rect 21486 3934 21546 4966
rect 21606 3996 21666 5026
rect 21726 3934 21786 4966
rect 21846 3996 21906 5026
rect 21966 4872 22032 4962
rect 21966 4808 21967 4872
rect 22031 4808 22032 4872
rect 21966 4792 22032 4808
rect 21966 4728 21967 4792
rect 22031 4728 22032 4792
rect 21966 4712 22032 4728
rect 21966 4648 21967 4712
rect 22031 4648 22032 4712
rect 21966 4632 22032 4648
rect 21966 4568 21967 4632
rect 22031 4568 22032 4632
rect 21966 4552 22032 4568
rect 21966 4488 21967 4552
rect 22031 4488 22032 4552
rect 21966 4472 22032 4488
rect 21966 4408 21967 4472
rect 22031 4408 22032 4472
rect 21966 4392 22032 4408
rect 21966 4328 21967 4392
rect 22031 4328 22032 4392
rect 21966 4312 22032 4328
rect 21966 4248 21967 4312
rect 22031 4248 22032 4312
rect 21966 4232 22032 4248
rect 21966 4168 21967 4232
rect 22031 4168 22032 4232
rect 21966 4152 22032 4168
rect 21966 4088 21967 4152
rect 22031 4088 22032 4152
rect 21966 3934 22032 4088
rect 22092 3934 22152 4966
rect 22212 3996 22272 5026
rect 22332 3934 22392 4966
rect 22452 3996 22512 5026
rect 22572 4872 22638 4962
rect 22572 4808 22573 4872
rect 22637 4808 22638 4872
rect 22572 4792 22638 4808
rect 22572 4728 22573 4792
rect 22637 4728 22638 4792
rect 22572 4712 22638 4728
rect 22572 4648 22573 4712
rect 22637 4648 22638 4712
rect 22572 4632 22638 4648
rect 22572 4568 22573 4632
rect 22637 4568 22638 4632
rect 22572 4552 22638 4568
rect 22572 4488 22573 4552
rect 22637 4488 22638 4552
rect 22572 4472 22638 4488
rect 22572 4408 22573 4472
rect 22637 4408 22638 4472
rect 22572 4392 22638 4408
rect 22572 4328 22573 4392
rect 22637 4328 22638 4392
rect 22572 4312 22638 4328
rect 22572 4248 22573 4312
rect 22637 4248 22638 4312
rect 22572 4232 22638 4248
rect 22572 4168 22573 4232
rect 22637 4168 22638 4232
rect 22572 4152 22638 4168
rect 22572 4088 22573 4152
rect 22637 4088 22638 4152
rect 22572 3934 22638 4088
rect 22698 3934 22758 4966
rect 22818 3996 22878 5026
rect 22938 3934 22998 4966
rect 23058 3996 23118 5026
rect 23178 4872 23244 4962
rect 23178 4808 23179 4872
rect 23243 4808 23244 4872
rect 23178 4792 23244 4808
rect 23178 4728 23179 4792
rect 23243 4728 23244 4792
rect 23178 4712 23244 4728
rect 23178 4648 23179 4712
rect 23243 4648 23244 4712
rect 23178 4632 23244 4648
rect 23178 4568 23179 4632
rect 23243 4568 23244 4632
rect 23178 4552 23244 4568
rect 23178 4488 23179 4552
rect 23243 4488 23244 4552
rect 23178 4472 23244 4488
rect 23178 4408 23179 4472
rect 23243 4408 23244 4472
rect 23178 4392 23244 4408
rect 23178 4328 23179 4392
rect 23243 4328 23244 4392
rect 23178 4312 23244 4328
rect 23178 4248 23179 4312
rect 23243 4248 23244 4312
rect 23178 4232 23244 4248
rect 23178 4168 23179 4232
rect 23243 4168 23244 4232
rect 23178 4152 23244 4168
rect 23178 4088 23179 4152
rect 23243 4088 23244 4152
rect 23178 3934 23244 4088
rect 23304 3934 23364 4966
rect 23424 3996 23484 5026
rect 23544 3934 23604 4966
rect 23664 3996 23724 5026
rect 23784 4872 23850 4962
rect 23784 4808 23785 4872
rect 23849 4808 23850 4872
rect 23784 4792 23850 4808
rect 23784 4728 23785 4792
rect 23849 4728 23850 4792
rect 23784 4712 23850 4728
rect 23784 4648 23785 4712
rect 23849 4648 23850 4712
rect 23784 4632 23850 4648
rect 23784 4568 23785 4632
rect 23849 4568 23850 4632
rect 23784 4552 23850 4568
rect 23784 4488 23785 4552
rect 23849 4488 23850 4552
rect 23784 4472 23850 4488
rect 23784 4408 23785 4472
rect 23849 4408 23850 4472
rect 23784 4392 23850 4408
rect 23784 4328 23785 4392
rect 23849 4328 23850 4392
rect 23784 4312 23850 4328
rect 23784 4248 23785 4312
rect 23849 4248 23850 4312
rect 23784 4232 23850 4248
rect 23784 4168 23785 4232
rect 23849 4168 23850 4232
rect 23784 4152 23850 4168
rect 23784 4088 23785 4152
rect 23849 4088 23850 4152
rect 23784 3934 23850 4088
rect 23910 3934 23970 4966
rect 24030 3996 24090 5026
rect 24150 3934 24210 4966
rect 24270 3996 24330 5026
rect 24390 4872 24456 4962
rect 24390 4808 24391 4872
rect 24455 4808 24456 4872
rect 24390 4792 24456 4808
rect 24390 4728 24391 4792
rect 24455 4728 24456 4792
rect 24390 4712 24456 4728
rect 24390 4648 24391 4712
rect 24455 4648 24456 4712
rect 24390 4632 24456 4648
rect 24390 4568 24391 4632
rect 24455 4568 24456 4632
rect 24390 4552 24456 4568
rect 24390 4488 24391 4552
rect 24455 4488 24456 4552
rect 24390 4472 24456 4488
rect 24390 4408 24391 4472
rect 24455 4408 24456 4472
rect 24390 4392 24456 4408
rect 24390 4328 24391 4392
rect 24455 4328 24456 4392
rect 24390 4312 24456 4328
rect 24390 4248 24391 4312
rect 24455 4248 24456 4312
rect 24390 4232 24456 4248
rect 24390 4168 24391 4232
rect 24455 4168 24456 4232
rect 24390 4152 24456 4168
rect 24390 4088 24391 4152
rect 24455 4088 24456 4152
rect 24390 3934 24456 4088
rect 24516 3934 24576 4966
rect 24636 3996 24696 5026
rect 24756 3934 24816 4966
rect 24876 3996 24936 5026
rect 24996 4872 25062 4962
rect 24996 4808 24997 4872
rect 25061 4808 25062 4872
rect 24996 4792 25062 4808
rect 24996 4728 24997 4792
rect 25061 4728 25062 4792
rect 24996 4712 25062 4728
rect 24996 4648 24997 4712
rect 25061 4648 25062 4712
rect 24996 4632 25062 4648
rect 24996 4568 24997 4632
rect 25061 4568 25062 4632
rect 24996 4552 25062 4568
rect 24996 4488 24997 4552
rect 25061 4488 25062 4552
rect 24996 4472 25062 4488
rect 24996 4408 24997 4472
rect 25061 4408 25062 4472
rect 24996 4392 25062 4408
rect 24996 4328 24997 4392
rect 25061 4328 25062 4392
rect 24996 4312 25062 4328
rect 24996 4248 24997 4312
rect 25061 4248 25062 4312
rect 24996 4232 25062 4248
rect 24996 4168 24997 4232
rect 25061 4168 25062 4232
rect 24996 4152 25062 4168
rect 24996 4088 24997 4152
rect 25061 4088 25062 4152
rect 24996 3934 25062 4088
rect 25122 3934 25182 4966
rect 25242 3996 25302 5026
rect 25362 3934 25422 4966
rect 25482 3996 25542 5026
rect 25602 4872 25668 4962
rect 25602 4808 25603 4872
rect 25667 4808 25668 4872
rect 25602 4792 25668 4808
rect 25602 4728 25603 4792
rect 25667 4728 25668 4792
rect 25602 4712 25668 4728
rect 25602 4648 25603 4712
rect 25667 4648 25668 4712
rect 25602 4632 25668 4648
rect 25602 4568 25603 4632
rect 25667 4568 25668 4632
rect 25602 4552 25668 4568
rect 25602 4488 25603 4552
rect 25667 4488 25668 4552
rect 25602 4472 25668 4488
rect 25602 4408 25603 4472
rect 25667 4408 25668 4472
rect 25602 4392 25668 4408
rect 25602 4328 25603 4392
rect 25667 4328 25668 4392
rect 25602 4312 25668 4328
rect 25602 4248 25603 4312
rect 25667 4248 25668 4312
rect 25602 4232 25668 4248
rect 25602 4168 25603 4232
rect 25667 4168 25668 4232
rect 25602 4152 25668 4168
rect 25602 4088 25603 4152
rect 25667 4088 25668 4152
rect 25602 3934 25668 4088
rect 25728 3934 25788 4966
rect 25848 3996 25908 5026
rect 25968 3934 26028 4966
rect 26088 3996 26148 5026
rect 26208 4872 26274 4962
rect 26208 4808 26209 4872
rect 26273 4808 26274 4872
rect 26208 4792 26274 4808
rect 26208 4728 26209 4792
rect 26273 4728 26274 4792
rect 26208 4712 26274 4728
rect 26208 4648 26209 4712
rect 26273 4648 26274 4712
rect 26208 4632 26274 4648
rect 26208 4568 26209 4632
rect 26273 4568 26274 4632
rect 26208 4552 26274 4568
rect 26208 4488 26209 4552
rect 26273 4488 26274 4552
rect 26208 4472 26274 4488
rect 26208 4408 26209 4472
rect 26273 4408 26274 4472
rect 26208 4392 26274 4408
rect 26208 4328 26209 4392
rect 26273 4328 26274 4392
rect 26208 4312 26274 4328
rect 26208 4248 26209 4312
rect 26273 4248 26274 4312
rect 26208 4232 26274 4248
rect 26208 4168 26209 4232
rect 26273 4168 26274 4232
rect 26208 4152 26274 4168
rect 26208 4088 26209 4152
rect 26273 4088 26274 4152
rect 26208 3934 26274 4088
rect 26334 3934 26394 4966
rect 26454 3996 26514 5026
rect 26574 3934 26634 4966
rect 26694 3996 26754 5026
rect 26814 4872 26880 4962
rect 26814 4808 26815 4872
rect 26879 4808 26880 4872
rect 26814 4792 26880 4808
rect 26814 4728 26815 4792
rect 26879 4728 26880 4792
rect 26814 4712 26880 4728
rect 26814 4648 26815 4712
rect 26879 4648 26880 4712
rect 26814 4632 26880 4648
rect 26814 4568 26815 4632
rect 26879 4568 26880 4632
rect 26814 4552 26880 4568
rect 26814 4488 26815 4552
rect 26879 4488 26880 4552
rect 26814 4472 26880 4488
rect 26814 4408 26815 4472
rect 26879 4408 26880 4472
rect 26814 4392 26880 4408
rect 26814 4328 26815 4392
rect 26879 4328 26880 4392
rect 26814 4312 26880 4328
rect 26814 4248 26815 4312
rect 26879 4248 26880 4312
rect 26814 4232 26880 4248
rect 26814 4168 26815 4232
rect 26879 4168 26880 4232
rect 26814 4152 26880 4168
rect 26814 4088 26815 4152
rect 26879 4088 26880 4152
rect 26814 3934 26880 4088
rect 26940 3934 27000 4966
rect 27060 3996 27120 5026
rect 27180 3934 27240 4966
rect 27300 3996 27360 5026
rect 27420 4872 27486 4962
rect 27420 4808 27421 4872
rect 27485 4808 27486 4872
rect 27420 4792 27486 4808
rect 27420 4728 27421 4792
rect 27485 4728 27486 4792
rect 27420 4712 27486 4728
rect 27420 4648 27421 4712
rect 27485 4648 27486 4712
rect 27420 4632 27486 4648
rect 27420 4568 27421 4632
rect 27485 4568 27486 4632
rect 27420 4552 27486 4568
rect 27420 4488 27421 4552
rect 27485 4488 27486 4552
rect 27420 4472 27486 4488
rect 27420 4408 27421 4472
rect 27485 4408 27486 4472
rect 27420 4392 27486 4408
rect 27420 4328 27421 4392
rect 27485 4328 27486 4392
rect 27420 4312 27486 4328
rect 27420 4248 27421 4312
rect 27485 4248 27486 4312
rect 27420 4232 27486 4248
rect 27420 4168 27421 4232
rect 27485 4168 27486 4232
rect 27420 4152 27486 4168
rect 27420 4088 27421 4152
rect 27485 4088 27486 4152
rect 27420 3934 27486 4088
rect 27546 3934 27606 4966
rect 27666 3996 27726 5026
rect 27786 3934 27846 4966
rect 27906 3996 27966 5026
rect 28026 4872 28092 4962
rect 28026 4808 28027 4872
rect 28091 4808 28092 4872
rect 28026 4792 28092 4808
rect 28026 4728 28027 4792
rect 28091 4728 28092 4792
rect 28026 4712 28092 4728
rect 28026 4648 28027 4712
rect 28091 4648 28092 4712
rect 28026 4632 28092 4648
rect 28026 4568 28027 4632
rect 28091 4568 28092 4632
rect 28026 4552 28092 4568
rect 28026 4488 28027 4552
rect 28091 4488 28092 4552
rect 28026 4472 28092 4488
rect 28026 4408 28027 4472
rect 28091 4408 28092 4472
rect 28026 4392 28092 4408
rect 28026 4328 28027 4392
rect 28091 4328 28092 4392
rect 28026 4312 28092 4328
rect 28026 4248 28027 4312
rect 28091 4248 28092 4312
rect 28026 4232 28092 4248
rect 28026 4168 28027 4232
rect 28091 4168 28092 4232
rect 28026 4152 28092 4168
rect 28026 4088 28027 4152
rect 28091 4088 28092 4152
rect 28026 3934 28092 4088
rect 28152 3934 28212 4966
rect 28272 3996 28332 5026
rect 28392 3934 28452 4966
rect 28512 3996 28572 5026
rect 28632 4872 28698 4962
rect 28632 4808 28633 4872
rect 28697 4808 28698 4872
rect 28632 4792 28698 4808
rect 28632 4728 28633 4792
rect 28697 4728 28698 4792
rect 28632 4712 28698 4728
rect 28632 4648 28633 4712
rect 28697 4648 28698 4712
rect 28632 4632 28698 4648
rect 28632 4568 28633 4632
rect 28697 4568 28698 4632
rect 28632 4552 28698 4568
rect 28632 4488 28633 4552
rect 28697 4488 28698 4552
rect 28632 4472 28698 4488
rect 28632 4408 28633 4472
rect 28697 4408 28698 4472
rect 28632 4392 28698 4408
rect 28632 4328 28633 4392
rect 28697 4328 28698 4392
rect 28632 4312 28698 4328
rect 28632 4248 28633 4312
rect 28697 4248 28698 4312
rect 28632 4232 28698 4248
rect 28632 4168 28633 4232
rect 28697 4168 28698 4232
rect 28632 4152 28698 4168
rect 28632 4088 28633 4152
rect 28697 4088 28698 4152
rect 28632 3934 28698 4088
rect 28758 3934 28818 4966
rect 28878 3996 28938 5026
rect 28998 3934 29058 4966
rect 29118 3996 29178 5026
rect 29238 4872 29304 4962
rect 29238 4808 29239 4872
rect 29303 4808 29304 4872
rect 29238 4792 29304 4808
rect 29238 4728 29239 4792
rect 29303 4728 29304 4792
rect 29238 4712 29304 4728
rect 29238 4648 29239 4712
rect 29303 4648 29304 4712
rect 29238 4632 29304 4648
rect 29238 4568 29239 4632
rect 29303 4568 29304 4632
rect 29238 4552 29304 4568
rect 29238 4488 29239 4552
rect 29303 4488 29304 4552
rect 29238 4472 29304 4488
rect 29238 4408 29239 4472
rect 29303 4408 29304 4472
rect 29238 4392 29304 4408
rect 29238 4328 29239 4392
rect 29303 4328 29304 4392
rect 29238 4312 29304 4328
rect 29238 4248 29239 4312
rect 29303 4248 29304 4312
rect 29238 4232 29304 4248
rect 29238 4168 29239 4232
rect 29303 4168 29304 4232
rect 29238 4152 29304 4168
rect 29238 4088 29239 4152
rect 29303 4088 29304 4152
rect 29238 3934 29304 4088
rect 29364 3934 29424 4966
rect 29484 3996 29544 5026
rect 29604 3934 29664 4966
rect 29724 3996 29784 5026
rect 29844 4872 29910 4962
rect 29844 4808 29845 4872
rect 29909 4808 29910 4872
rect 29844 4792 29910 4808
rect 29844 4728 29845 4792
rect 29909 4728 29910 4792
rect 29844 4712 29910 4728
rect 29844 4648 29845 4712
rect 29909 4648 29910 4712
rect 29844 4632 29910 4648
rect 29844 4568 29845 4632
rect 29909 4568 29910 4632
rect 29844 4552 29910 4568
rect 29844 4488 29845 4552
rect 29909 4488 29910 4552
rect 29844 4472 29910 4488
rect 29844 4408 29845 4472
rect 29909 4408 29910 4472
rect 29844 4392 29910 4408
rect 29844 4328 29845 4392
rect 29909 4328 29910 4392
rect 29844 4312 29910 4328
rect 29844 4248 29845 4312
rect 29909 4248 29910 4312
rect 29844 4232 29910 4248
rect 29844 4168 29845 4232
rect 29909 4168 29910 4232
rect 29844 4152 29910 4168
rect 29844 4088 29845 4152
rect 29909 4088 29910 4152
rect 29844 3934 29910 4088
rect 29970 3934 30030 4966
rect 30090 3996 30150 5026
rect 30210 3934 30270 4966
rect 30330 3996 30390 5026
rect 30450 4872 30516 4962
rect 30450 4808 30451 4872
rect 30515 4808 30516 4872
rect 30450 4792 30516 4808
rect 30450 4728 30451 4792
rect 30515 4728 30516 4792
rect 30450 4712 30516 4728
rect 30450 4648 30451 4712
rect 30515 4648 30516 4712
rect 30450 4632 30516 4648
rect 30450 4568 30451 4632
rect 30515 4568 30516 4632
rect 30450 4552 30516 4568
rect 30450 4488 30451 4552
rect 30515 4488 30516 4552
rect 30450 4472 30516 4488
rect 30450 4408 30451 4472
rect 30515 4408 30516 4472
rect 30450 4392 30516 4408
rect 30450 4328 30451 4392
rect 30515 4328 30516 4392
rect 30450 4312 30516 4328
rect 30450 4248 30451 4312
rect 30515 4248 30516 4312
rect 30450 4232 30516 4248
rect 30450 4168 30451 4232
rect 30515 4168 30516 4232
rect 30450 4152 30516 4168
rect 30450 4088 30451 4152
rect 30515 4088 30516 4152
rect 30450 3934 30516 4088
rect 30576 3934 30636 4966
rect 30696 3996 30756 5026
rect 30816 3934 30876 4966
rect 30936 3996 30996 5026
rect 31056 4872 31122 4962
rect 31056 4808 31057 4872
rect 31121 4808 31122 4872
rect 31056 4792 31122 4808
rect 31056 4728 31057 4792
rect 31121 4728 31122 4792
rect 31056 4712 31122 4728
rect 31056 4648 31057 4712
rect 31121 4648 31122 4712
rect 31056 4632 31122 4648
rect 31056 4568 31057 4632
rect 31121 4568 31122 4632
rect 31056 4552 31122 4568
rect 31056 4488 31057 4552
rect 31121 4488 31122 4552
rect 31056 4472 31122 4488
rect 31056 4408 31057 4472
rect 31121 4408 31122 4472
rect 31056 4392 31122 4408
rect 31056 4328 31057 4392
rect 31121 4328 31122 4392
rect 31056 4312 31122 4328
rect 31056 4248 31057 4312
rect 31121 4248 31122 4312
rect 31056 4232 31122 4248
rect 31056 4168 31057 4232
rect 31121 4168 31122 4232
rect 31056 4152 31122 4168
rect 31056 4088 31057 4152
rect 31121 4088 31122 4152
rect 31056 3934 31122 4088
rect 31182 3934 31242 4966
rect 31302 3996 31362 5026
rect 31422 3934 31482 4966
rect 31542 3996 31602 5026
rect 31662 4872 31728 4962
rect 31662 4808 31663 4872
rect 31727 4808 31728 4872
rect 31662 4792 31728 4808
rect 31662 4728 31663 4792
rect 31727 4728 31728 4792
rect 31662 4712 31728 4728
rect 31662 4648 31663 4712
rect 31727 4648 31728 4712
rect 31662 4632 31728 4648
rect 31662 4568 31663 4632
rect 31727 4568 31728 4632
rect 31662 4552 31728 4568
rect 31662 4488 31663 4552
rect 31727 4488 31728 4552
rect 31662 4472 31728 4488
rect 31662 4408 31663 4472
rect 31727 4408 31728 4472
rect 31662 4392 31728 4408
rect 31662 4328 31663 4392
rect 31727 4328 31728 4392
rect 31662 4312 31728 4328
rect 31662 4248 31663 4312
rect 31727 4248 31728 4312
rect 31662 4232 31728 4248
rect 31662 4168 31663 4232
rect 31727 4168 31728 4232
rect 31662 4152 31728 4168
rect 31662 4088 31663 4152
rect 31727 4088 31728 4152
rect 31662 3934 31728 4088
rect 31788 3934 31848 4966
rect 31908 3996 31968 5026
rect 32028 3934 32088 4966
rect 32148 3996 32208 5026
rect 32268 4872 32334 4962
rect 32268 4808 32269 4872
rect 32333 4808 32334 4872
rect 32268 4792 32334 4808
rect 32268 4728 32269 4792
rect 32333 4728 32334 4792
rect 32268 4712 32334 4728
rect 32268 4648 32269 4712
rect 32333 4648 32334 4712
rect 32268 4632 32334 4648
rect 32268 4568 32269 4632
rect 32333 4568 32334 4632
rect 32268 4552 32334 4568
rect 32268 4488 32269 4552
rect 32333 4488 32334 4552
rect 32268 4472 32334 4488
rect 32268 4408 32269 4472
rect 32333 4408 32334 4472
rect 32268 4392 32334 4408
rect 32268 4328 32269 4392
rect 32333 4328 32334 4392
rect 32268 4312 32334 4328
rect 32268 4248 32269 4312
rect 32333 4248 32334 4312
rect 32268 4232 32334 4248
rect 32268 4168 32269 4232
rect 32333 4168 32334 4232
rect 32268 4152 32334 4168
rect 32268 4088 32269 4152
rect 32333 4088 32334 4152
rect 32268 3934 32334 4088
rect 32394 3934 32454 4966
rect 32514 3996 32574 5026
rect 32634 3934 32694 4966
rect 32754 3996 32814 5026
rect 32874 4872 32940 4962
rect 32874 4808 32875 4872
rect 32939 4808 32940 4872
rect 32874 4792 32940 4808
rect 32874 4728 32875 4792
rect 32939 4728 32940 4792
rect 32874 4712 32940 4728
rect 32874 4648 32875 4712
rect 32939 4648 32940 4712
rect 32874 4632 32940 4648
rect 32874 4568 32875 4632
rect 32939 4568 32940 4632
rect 32874 4552 32940 4568
rect 32874 4488 32875 4552
rect 32939 4488 32940 4552
rect 32874 4472 32940 4488
rect 32874 4408 32875 4472
rect 32939 4408 32940 4472
rect 32874 4392 32940 4408
rect 32874 4328 32875 4392
rect 32939 4328 32940 4392
rect 32874 4312 32940 4328
rect 32874 4248 32875 4312
rect 32939 4248 32940 4312
rect 32874 4232 32940 4248
rect 32874 4168 32875 4232
rect 32939 4168 32940 4232
rect 32874 4152 32940 4168
rect 32874 4088 32875 4152
rect 32939 4088 32940 4152
rect 32874 3934 32940 4088
rect 33000 3934 33060 4966
rect 33120 3996 33180 5026
rect 33240 3934 33300 4966
rect 33360 3996 33420 5026
rect 33480 4872 33546 4962
rect 33480 4808 33481 4872
rect 33545 4808 33546 4872
rect 33480 4792 33546 4808
rect 33480 4728 33481 4792
rect 33545 4728 33546 4792
rect 33480 4712 33546 4728
rect 33480 4648 33481 4712
rect 33545 4648 33546 4712
rect 33480 4632 33546 4648
rect 33480 4568 33481 4632
rect 33545 4568 33546 4632
rect 33480 4552 33546 4568
rect 33480 4488 33481 4552
rect 33545 4488 33546 4552
rect 33480 4472 33546 4488
rect 33480 4408 33481 4472
rect 33545 4408 33546 4472
rect 33480 4392 33546 4408
rect 33480 4328 33481 4392
rect 33545 4328 33546 4392
rect 33480 4312 33546 4328
rect 33480 4248 33481 4312
rect 33545 4248 33546 4312
rect 33480 4232 33546 4248
rect 33480 4168 33481 4232
rect 33545 4168 33546 4232
rect 33480 4152 33546 4168
rect 33480 4088 33481 4152
rect 33545 4088 33546 4152
rect 33480 3934 33546 4088
rect 33606 3934 33666 4966
rect 33726 3996 33786 5026
rect 33846 3934 33906 4966
rect 33966 3996 34026 5026
rect 34086 4872 34152 4962
rect 34086 4808 34087 4872
rect 34151 4808 34152 4872
rect 34086 4792 34152 4808
rect 34086 4728 34087 4792
rect 34151 4728 34152 4792
rect 34086 4712 34152 4728
rect 34086 4648 34087 4712
rect 34151 4648 34152 4712
rect 34086 4632 34152 4648
rect 34086 4568 34087 4632
rect 34151 4568 34152 4632
rect 34086 4552 34152 4568
rect 34086 4488 34087 4552
rect 34151 4488 34152 4552
rect 34086 4472 34152 4488
rect 34086 4408 34087 4472
rect 34151 4408 34152 4472
rect 34086 4392 34152 4408
rect 34086 4328 34087 4392
rect 34151 4328 34152 4392
rect 34086 4312 34152 4328
rect 34086 4248 34087 4312
rect 34151 4248 34152 4312
rect 34086 4232 34152 4248
rect 34086 4168 34087 4232
rect 34151 4168 34152 4232
rect 34086 4152 34152 4168
rect 34086 4088 34087 4152
rect 34151 4088 34152 4152
rect 34086 3934 34152 4088
rect 34212 3934 34272 4966
rect 34332 3996 34392 5026
rect 34452 3934 34512 4966
rect 34572 3996 34632 5026
rect 34692 4872 34758 4962
rect 34692 4808 34693 4872
rect 34757 4808 34758 4872
rect 34692 4792 34758 4808
rect 34692 4728 34693 4792
rect 34757 4728 34758 4792
rect 34692 4712 34758 4728
rect 34692 4648 34693 4712
rect 34757 4648 34758 4712
rect 34692 4632 34758 4648
rect 34692 4568 34693 4632
rect 34757 4568 34758 4632
rect 34692 4552 34758 4568
rect 34692 4488 34693 4552
rect 34757 4488 34758 4552
rect 34692 4472 34758 4488
rect 34692 4408 34693 4472
rect 34757 4408 34758 4472
rect 34692 4392 34758 4408
rect 34692 4328 34693 4392
rect 34757 4328 34758 4392
rect 34692 4312 34758 4328
rect 34692 4248 34693 4312
rect 34757 4248 34758 4312
rect 34692 4232 34758 4248
rect 34692 4168 34693 4232
rect 34757 4168 34758 4232
rect 34692 4152 34758 4168
rect 34692 4088 34693 4152
rect 34757 4088 34758 4152
rect 34692 3934 34758 4088
rect 34818 3934 34878 4966
rect 34938 3996 34998 5026
rect 35058 3934 35118 4966
rect 35178 3996 35238 5026
rect 35298 4872 35364 4962
rect 35298 4808 35299 4872
rect 35363 4808 35364 4872
rect 35298 4792 35364 4808
rect 35298 4728 35299 4792
rect 35363 4728 35364 4792
rect 35298 4712 35364 4728
rect 35298 4648 35299 4712
rect 35363 4648 35364 4712
rect 35298 4632 35364 4648
rect 35298 4568 35299 4632
rect 35363 4568 35364 4632
rect 35298 4552 35364 4568
rect 35298 4488 35299 4552
rect 35363 4488 35364 4552
rect 35298 4472 35364 4488
rect 35298 4408 35299 4472
rect 35363 4408 35364 4472
rect 35298 4392 35364 4408
rect 35298 4328 35299 4392
rect 35363 4328 35364 4392
rect 35298 4312 35364 4328
rect 35298 4248 35299 4312
rect 35363 4248 35364 4312
rect 35298 4232 35364 4248
rect 35298 4168 35299 4232
rect 35363 4168 35364 4232
rect 35298 4152 35364 4168
rect 35298 4088 35299 4152
rect 35363 4088 35364 4152
rect 35298 3934 35364 4088
rect 35424 3934 35484 4966
rect 35544 3996 35604 5026
rect 35664 3934 35724 4966
rect 35784 3996 35844 5026
rect 35904 4872 35970 4962
rect 35904 4808 35905 4872
rect 35969 4808 35970 4872
rect 35904 4792 35970 4808
rect 35904 4728 35905 4792
rect 35969 4728 35970 4792
rect 35904 4712 35970 4728
rect 35904 4648 35905 4712
rect 35969 4648 35970 4712
rect 35904 4632 35970 4648
rect 35904 4568 35905 4632
rect 35969 4568 35970 4632
rect 35904 4552 35970 4568
rect 35904 4488 35905 4552
rect 35969 4488 35970 4552
rect 35904 4472 35970 4488
rect 35904 4408 35905 4472
rect 35969 4408 35970 4472
rect 35904 4392 35970 4408
rect 35904 4328 35905 4392
rect 35969 4328 35970 4392
rect 35904 4312 35970 4328
rect 35904 4248 35905 4312
rect 35969 4248 35970 4312
rect 35904 4232 35970 4248
rect 35904 4168 35905 4232
rect 35969 4168 35970 4232
rect 35904 4152 35970 4168
rect 35904 4088 35905 4152
rect 35969 4088 35970 4152
rect 35904 3934 35970 4088
rect 36030 3934 36090 4966
rect 36150 3996 36210 5026
rect 36270 3934 36330 4966
rect 36390 3996 36450 5026
rect 36510 4872 36576 4962
rect 36510 4808 36511 4872
rect 36575 4808 36576 4872
rect 36510 4792 36576 4808
rect 36510 4728 36511 4792
rect 36575 4728 36576 4792
rect 36510 4712 36576 4728
rect 36510 4648 36511 4712
rect 36575 4648 36576 4712
rect 36510 4632 36576 4648
rect 36510 4568 36511 4632
rect 36575 4568 36576 4632
rect 36510 4552 36576 4568
rect 36510 4488 36511 4552
rect 36575 4488 36576 4552
rect 36510 4472 36576 4488
rect 36510 4408 36511 4472
rect 36575 4408 36576 4472
rect 36510 4392 36576 4408
rect 36510 4328 36511 4392
rect 36575 4328 36576 4392
rect 36510 4312 36576 4328
rect 36510 4248 36511 4312
rect 36575 4248 36576 4312
rect 36510 4232 36576 4248
rect 36510 4168 36511 4232
rect 36575 4168 36576 4232
rect 36510 4152 36576 4168
rect 36510 4088 36511 4152
rect 36575 4088 36576 4152
rect 36510 3934 36576 4088
rect 36636 3934 36696 4966
rect 36756 3996 36816 5026
rect 36876 3934 36936 4966
rect 36996 3996 37056 5026
rect 37116 4872 37182 4962
rect 37116 4808 37117 4872
rect 37181 4808 37182 4872
rect 37116 4792 37182 4808
rect 37116 4728 37117 4792
rect 37181 4728 37182 4792
rect 37116 4712 37182 4728
rect 37116 4648 37117 4712
rect 37181 4648 37182 4712
rect 37116 4632 37182 4648
rect 37116 4568 37117 4632
rect 37181 4568 37182 4632
rect 37116 4552 37182 4568
rect 37116 4488 37117 4552
rect 37181 4488 37182 4552
rect 37116 4472 37182 4488
rect 37116 4408 37117 4472
rect 37181 4408 37182 4472
rect 37116 4392 37182 4408
rect 37116 4328 37117 4392
rect 37181 4328 37182 4392
rect 37116 4312 37182 4328
rect 37116 4248 37117 4312
rect 37181 4248 37182 4312
rect 37116 4232 37182 4248
rect 37116 4168 37117 4232
rect 37181 4168 37182 4232
rect 37116 4152 37182 4168
rect 37116 4088 37117 4152
rect 37181 4088 37182 4152
rect 37116 3934 37182 4088
rect 37242 3934 37302 4966
rect 37362 3996 37422 5026
rect 37482 3934 37542 4966
rect 37602 3996 37662 5026
rect 37722 4872 37788 4962
rect 37722 4808 37723 4872
rect 37787 4808 37788 4872
rect 37722 4792 37788 4808
rect 37722 4728 37723 4792
rect 37787 4728 37788 4792
rect 37722 4712 37788 4728
rect 37722 4648 37723 4712
rect 37787 4648 37788 4712
rect 37722 4632 37788 4648
rect 37722 4568 37723 4632
rect 37787 4568 37788 4632
rect 37722 4552 37788 4568
rect 37722 4488 37723 4552
rect 37787 4488 37788 4552
rect 37722 4472 37788 4488
rect 37722 4408 37723 4472
rect 37787 4408 37788 4472
rect 37722 4392 37788 4408
rect 37722 4328 37723 4392
rect 37787 4328 37788 4392
rect 37722 4312 37788 4328
rect 37722 4248 37723 4312
rect 37787 4248 37788 4312
rect 37722 4232 37788 4248
rect 37722 4168 37723 4232
rect 37787 4168 37788 4232
rect 37722 4152 37788 4168
rect 37722 4088 37723 4152
rect 37787 4088 37788 4152
rect 37722 3934 37788 4088
rect 37848 3934 37908 4966
rect 37968 3996 38028 5026
rect 38088 3934 38148 4966
rect 38208 3996 38268 5026
rect 38328 4872 38394 4962
rect 38328 4808 38329 4872
rect 38393 4808 38394 4872
rect 38328 4792 38394 4808
rect 38328 4728 38329 4792
rect 38393 4728 38394 4792
rect 38328 4712 38394 4728
rect 38328 4648 38329 4712
rect 38393 4648 38394 4712
rect 38328 4632 38394 4648
rect 38328 4568 38329 4632
rect 38393 4568 38394 4632
rect 38328 4552 38394 4568
rect 38328 4488 38329 4552
rect 38393 4488 38394 4552
rect 38328 4472 38394 4488
rect 38328 4408 38329 4472
rect 38393 4408 38394 4472
rect 38328 4392 38394 4408
rect 38328 4328 38329 4392
rect 38393 4328 38394 4392
rect 38328 4312 38394 4328
rect 38328 4248 38329 4312
rect 38393 4248 38394 4312
rect 38328 4232 38394 4248
rect 38328 4168 38329 4232
rect 38393 4168 38394 4232
rect 38328 4152 38394 4168
rect 38328 4088 38329 4152
rect 38393 4088 38394 4152
rect 38328 3934 38394 4088
rect 38454 3934 38514 4966
rect 38574 3996 38634 5026
rect 38694 3934 38754 4966
rect 38814 3996 38874 5026
rect 38934 4872 39000 4962
rect 38934 4808 38935 4872
rect 38999 4808 39000 4872
rect 38934 4792 39000 4808
rect 38934 4728 38935 4792
rect 38999 4728 39000 4792
rect 38934 4712 39000 4728
rect 38934 4648 38935 4712
rect 38999 4648 39000 4712
rect 38934 4632 39000 4648
rect 38934 4568 38935 4632
rect 38999 4568 39000 4632
rect 38934 4552 39000 4568
rect 38934 4488 38935 4552
rect 38999 4488 39000 4552
rect 38934 4472 39000 4488
rect 38934 4408 38935 4472
rect 38999 4408 39000 4472
rect 38934 4392 39000 4408
rect 38934 4328 38935 4392
rect 38999 4328 39000 4392
rect 38934 4312 39000 4328
rect 38934 4248 38935 4312
rect 38999 4248 39000 4312
rect 38934 4232 39000 4248
rect 38934 4168 38935 4232
rect 38999 4168 39000 4232
rect 38934 4152 39000 4168
rect 38934 4088 38935 4152
rect 38999 4088 39000 4152
rect 38934 3934 39000 4088
rect 39060 3934 39120 4966
rect 39180 3996 39240 5026
rect 39300 3934 39360 4966
rect 39420 3996 39480 5026
rect 39540 4872 39606 4962
rect 39540 4808 39541 4872
rect 39605 4808 39606 4872
rect 39540 4792 39606 4808
rect 39540 4728 39541 4792
rect 39605 4728 39606 4792
rect 39540 4712 39606 4728
rect 39540 4648 39541 4712
rect 39605 4648 39606 4712
rect 39540 4632 39606 4648
rect 39540 4568 39541 4632
rect 39605 4568 39606 4632
rect 39540 4552 39606 4568
rect 39540 4488 39541 4552
rect 39605 4488 39606 4552
rect 39540 4472 39606 4488
rect 39540 4408 39541 4472
rect 39605 4408 39606 4472
rect 39540 4392 39606 4408
rect 39540 4328 39541 4392
rect 39605 4328 39606 4392
rect 39540 4312 39606 4328
rect 39540 4248 39541 4312
rect 39605 4248 39606 4312
rect 39540 4232 39606 4248
rect 39540 4168 39541 4232
rect 39605 4168 39606 4232
rect 39540 4152 39606 4168
rect 39540 4088 39541 4152
rect 39605 4088 39606 4152
rect 39540 3934 39606 4088
rect 20148 3932 39606 3934
rect 20148 3868 20252 3932
rect 20316 3868 20332 3932
rect 20396 3868 20412 3932
rect 20476 3868 20492 3932
rect 20556 3868 20572 3932
rect 20636 3868 20652 3932
rect 20716 3868 20858 3932
rect 20922 3868 20938 3932
rect 21002 3868 21018 3932
rect 21082 3868 21098 3932
rect 21162 3868 21178 3932
rect 21242 3868 21258 3932
rect 21322 3868 21464 3932
rect 21528 3868 21544 3932
rect 21608 3868 21624 3932
rect 21688 3868 21704 3932
rect 21768 3868 21784 3932
rect 21848 3868 21864 3932
rect 21928 3868 22070 3932
rect 22134 3868 22150 3932
rect 22214 3868 22230 3932
rect 22294 3868 22310 3932
rect 22374 3868 22390 3932
rect 22454 3868 22470 3932
rect 22534 3868 22676 3932
rect 22740 3868 22756 3932
rect 22820 3868 22836 3932
rect 22900 3868 22916 3932
rect 22980 3868 22996 3932
rect 23060 3868 23076 3932
rect 23140 3868 23282 3932
rect 23346 3868 23362 3932
rect 23426 3868 23442 3932
rect 23506 3868 23522 3932
rect 23586 3868 23602 3932
rect 23666 3868 23682 3932
rect 23746 3868 23888 3932
rect 23952 3868 23968 3932
rect 24032 3868 24048 3932
rect 24112 3868 24128 3932
rect 24192 3868 24208 3932
rect 24272 3868 24288 3932
rect 24352 3868 24494 3932
rect 24558 3868 24574 3932
rect 24638 3868 24654 3932
rect 24718 3868 24734 3932
rect 24798 3868 24814 3932
rect 24878 3868 24894 3932
rect 24958 3868 25100 3932
rect 25164 3868 25180 3932
rect 25244 3868 25260 3932
rect 25324 3868 25340 3932
rect 25404 3868 25420 3932
rect 25484 3868 25500 3932
rect 25564 3868 25706 3932
rect 25770 3868 25786 3932
rect 25850 3868 25866 3932
rect 25930 3868 25946 3932
rect 26010 3868 26026 3932
rect 26090 3868 26106 3932
rect 26170 3868 26312 3932
rect 26376 3868 26392 3932
rect 26456 3868 26472 3932
rect 26536 3868 26552 3932
rect 26616 3868 26632 3932
rect 26696 3868 26712 3932
rect 26776 3868 26918 3932
rect 26982 3868 26998 3932
rect 27062 3868 27078 3932
rect 27142 3868 27158 3932
rect 27222 3868 27238 3932
rect 27302 3868 27318 3932
rect 27382 3868 27524 3932
rect 27588 3868 27604 3932
rect 27668 3868 27684 3932
rect 27748 3868 27764 3932
rect 27828 3868 27844 3932
rect 27908 3868 27924 3932
rect 27988 3868 28130 3932
rect 28194 3868 28210 3932
rect 28274 3868 28290 3932
rect 28354 3868 28370 3932
rect 28434 3868 28450 3932
rect 28514 3868 28530 3932
rect 28594 3868 28736 3932
rect 28800 3868 28816 3932
rect 28880 3868 28896 3932
rect 28960 3868 28976 3932
rect 29040 3868 29056 3932
rect 29120 3868 29136 3932
rect 29200 3868 29342 3932
rect 29406 3868 29422 3932
rect 29486 3868 29502 3932
rect 29566 3868 29582 3932
rect 29646 3868 29662 3932
rect 29726 3868 29742 3932
rect 29806 3868 29948 3932
rect 30012 3868 30028 3932
rect 30092 3868 30108 3932
rect 30172 3868 30188 3932
rect 30252 3868 30268 3932
rect 30332 3868 30348 3932
rect 30412 3868 30554 3932
rect 30618 3868 30634 3932
rect 30698 3868 30714 3932
rect 30778 3868 30794 3932
rect 30858 3868 30874 3932
rect 30938 3868 30954 3932
rect 31018 3868 31160 3932
rect 31224 3868 31240 3932
rect 31304 3868 31320 3932
rect 31384 3868 31400 3932
rect 31464 3868 31480 3932
rect 31544 3868 31560 3932
rect 31624 3868 31766 3932
rect 31830 3868 31846 3932
rect 31910 3868 31926 3932
rect 31990 3868 32006 3932
rect 32070 3868 32086 3932
rect 32150 3868 32166 3932
rect 32230 3868 32372 3932
rect 32436 3868 32452 3932
rect 32516 3868 32532 3932
rect 32596 3868 32612 3932
rect 32676 3868 32692 3932
rect 32756 3868 32772 3932
rect 32836 3868 32978 3932
rect 33042 3868 33058 3932
rect 33122 3868 33138 3932
rect 33202 3868 33218 3932
rect 33282 3868 33298 3932
rect 33362 3868 33378 3932
rect 33442 3868 33584 3932
rect 33648 3868 33664 3932
rect 33728 3868 33744 3932
rect 33808 3868 33824 3932
rect 33888 3868 33904 3932
rect 33968 3868 33984 3932
rect 34048 3868 34190 3932
rect 34254 3868 34270 3932
rect 34334 3868 34350 3932
rect 34414 3868 34430 3932
rect 34494 3868 34510 3932
rect 34574 3868 34590 3932
rect 34654 3868 34796 3932
rect 34860 3868 34876 3932
rect 34940 3868 34956 3932
rect 35020 3868 35036 3932
rect 35100 3868 35116 3932
rect 35180 3868 35196 3932
rect 35260 3868 35402 3932
rect 35466 3868 35482 3932
rect 35546 3868 35562 3932
rect 35626 3868 35642 3932
rect 35706 3868 35722 3932
rect 35786 3868 35802 3932
rect 35866 3868 36008 3932
rect 36072 3868 36088 3932
rect 36152 3868 36168 3932
rect 36232 3868 36248 3932
rect 36312 3868 36328 3932
rect 36392 3868 36408 3932
rect 36472 3868 36614 3932
rect 36678 3868 36694 3932
rect 36758 3868 36774 3932
rect 36838 3868 36854 3932
rect 36918 3868 36934 3932
rect 36998 3868 37014 3932
rect 37078 3868 37220 3932
rect 37284 3868 37300 3932
rect 37364 3868 37380 3932
rect 37444 3868 37460 3932
rect 37524 3868 37540 3932
rect 37604 3868 37620 3932
rect 37684 3868 37826 3932
rect 37890 3868 37906 3932
rect 37970 3868 37986 3932
rect 38050 3868 38066 3932
rect 38130 3868 38146 3932
rect 38210 3868 38226 3932
rect 38290 3868 38432 3932
rect 38496 3868 38512 3932
rect 38576 3868 38592 3932
rect 38656 3868 38672 3932
rect 38736 3868 38752 3932
rect 38816 3868 38832 3932
rect 38896 3868 39038 3932
rect 39102 3868 39118 3932
rect 39182 3868 39198 3932
rect 39262 3868 39278 3932
rect 39342 3868 39358 3932
rect 39422 3868 39438 3932
rect 39502 3868 39606 3932
rect 20148 3866 39606 3868
rect 20148 3712 20214 3866
rect 20148 3648 20149 3712
rect 20213 3648 20214 3712
rect 20148 3632 20214 3648
rect 20148 3568 20149 3632
rect 20213 3568 20214 3632
rect 20148 3552 20214 3568
rect 20148 3488 20149 3552
rect 20213 3488 20214 3552
rect 20148 3472 20214 3488
rect 20148 3408 20149 3472
rect 20213 3408 20214 3472
rect 20148 3392 20214 3408
rect 20148 3328 20149 3392
rect 20213 3328 20214 3392
rect 20148 3312 20214 3328
rect 20148 3248 20149 3312
rect 20213 3248 20214 3312
rect 20148 3232 20214 3248
rect 20148 3168 20149 3232
rect 20213 3168 20214 3232
rect 20148 3152 20214 3168
rect 20148 3088 20149 3152
rect 20213 3088 20214 3152
rect 20148 3072 20214 3088
rect 20148 3008 20149 3072
rect 20213 3008 20214 3072
rect 20148 2992 20214 3008
rect 20148 2928 20149 2992
rect 20213 2928 20214 2992
rect 20148 2838 20214 2928
rect 20274 2774 20334 3804
rect 20394 2834 20454 3866
rect 20514 2774 20574 3804
rect 20634 2834 20694 3866
rect 20754 3712 20820 3866
rect 20754 3648 20755 3712
rect 20819 3648 20820 3712
rect 20754 3632 20820 3648
rect 20754 3568 20755 3632
rect 20819 3568 20820 3632
rect 20754 3552 20820 3568
rect 20754 3488 20755 3552
rect 20819 3488 20820 3552
rect 20754 3472 20820 3488
rect 20754 3408 20755 3472
rect 20819 3408 20820 3472
rect 20754 3392 20820 3408
rect 20754 3328 20755 3392
rect 20819 3328 20820 3392
rect 20754 3312 20820 3328
rect 20754 3248 20755 3312
rect 20819 3248 20820 3312
rect 20754 3232 20820 3248
rect 20754 3168 20755 3232
rect 20819 3168 20820 3232
rect 20754 3152 20820 3168
rect 20754 3088 20755 3152
rect 20819 3088 20820 3152
rect 20754 3072 20820 3088
rect 20754 3008 20755 3072
rect 20819 3008 20820 3072
rect 20754 2992 20820 3008
rect 20754 2928 20755 2992
rect 20819 2928 20820 2992
rect 20754 2838 20820 2928
rect 20880 2774 20940 3804
rect 21000 2834 21060 3866
rect 21120 2774 21180 3804
rect 21240 2834 21300 3866
rect 21360 3712 21426 3866
rect 21360 3648 21361 3712
rect 21425 3648 21426 3712
rect 21360 3632 21426 3648
rect 21360 3568 21361 3632
rect 21425 3568 21426 3632
rect 21360 3552 21426 3568
rect 21360 3488 21361 3552
rect 21425 3488 21426 3552
rect 21360 3472 21426 3488
rect 21360 3408 21361 3472
rect 21425 3408 21426 3472
rect 21360 3392 21426 3408
rect 21360 3328 21361 3392
rect 21425 3328 21426 3392
rect 21360 3312 21426 3328
rect 21360 3248 21361 3312
rect 21425 3248 21426 3312
rect 21360 3232 21426 3248
rect 21360 3168 21361 3232
rect 21425 3168 21426 3232
rect 21360 3152 21426 3168
rect 21360 3088 21361 3152
rect 21425 3088 21426 3152
rect 21360 3072 21426 3088
rect 21360 3008 21361 3072
rect 21425 3008 21426 3072
rect 21360 2992 21426 3008
rect 21360 2928 21361 2992
rect 21425 2928 21426 2992
rect 21360 2838 21426 2928
rect 21486 2774 21546 3804
rect 21606 2834 21666 3866
rect 21726 2774 21786 3804
rect 21846 2834 21906 3866
rect 21966 3712 22032 3866
rect 21966 3648 21967 3712
rect 22031 3648 22032 3712
rect 21966 3632 22032 3648
rect 21966 3568 21967 3632
rect 22031 3568 22032 3632
rect 21966 3552 22032 3568
rect 21966 3488 21967 3552
rect 22031 3488 22032 3552
rect 21966 3472 22032 3488
rect 21966 3408 21967 3472
rect 22031 3408 22032 3472
rect 21966 3392 22032 3408
rect 21966 3328 21967 3392
rect 22031 3328 22032 3392
rect 21966 3312 22032 3328
rect 21966 3248 21967 3312
rect 22031 3248 22032 3312
rect 21966 3232 22032 3248
rect 21966 3168 21967 3232
rect 22031 3168 22032 3232
rect 21966 3152 22032 3168
rect 21966 3088 21967 3152
rect 22031 3088 22032 3152
rect 21966 3072 22032 3088
rect 21966 3008 21967 3072
rect 22031 3008 22032 3072
rect 21966 2992 22032 3008
rect 21966 2928 21967 2992
rect 22031 2928 22032 2992
rect 21966 2838 22032 2928
rect 22092 2774 22152 3804
rect 22212 2834 22272 3866
rect 22332 2774 22392 3804
rect 22452 2834 22512 3866
rect 22572 3712 22638 3866
rect 22572 3648 22573 3712
rect 22637 3648 22638 3712
rect 22572 3632 22638 3648
rect 22572 3568 22573 3632
rect 22637 3568 22638 3632
rect 22572 3552 22638 3568
rect 22572 3488 22573 3552
rect 22637 3488 22638 3552
rect 22572 3472 22638 3488
rect 22572 3408 22573 3472
rect 22637 3408 22638 3472
rect 22572 3392 22638 3408
rect 22572 3328 22573 3392
rect 22637 3328 22638 3392
rect 22572 3312 22638 3328
rect 22572 3248 22573 3312
rect 22637 3248 22638 3312
rect 22572 3232 22638 3248
rect 22572 3168 22573 3232
rect 22637 3168 22638 3232
rect 22572 3152 22638 3168
rect 22572 3088 22573 3152
rect 22637 3088 22638 3152
rect 22572 3072 22638 3088
rect 22572 3008 22573 3072
rect 22637 3008 22638 3072
rect 22572 2992 22638 3008
rect 22572 2928 22573 2992
rect 22637 2928 22638 2992
rect 22572 2838 22638 2928
rect 22698 2774 22758 3804
rect 22818 2834 22878 3866
rect 22938 2774 22998 3804
rect 23058 2834 23118 3866
rect 23178 3712 23244 3866
rect 23178 3648 23179 3712
rect 23243 3648 23244 3712
rect 23178 3632 23244 3648
rect 23178 3568 23179 3632
rect 23243 3568 23244 3632
rect 23178 3552 23244 3568
rect 23178 3488 23179 3552
rect 23243 3488 23244 3552
rect 23178 3472 23244 3488
rect 23178 3408 23179 3472
rect 23243 3408 23244 3472
rect 23178 3392 23244 3408
rect 23178 3328 23179 3392
rect 23243 3328 23244 3392
rect 23178 3312 23244 3328
rect 23178 3248 23179 3312
rect 23243 3248 23244 3312
rect 23178 3232 23244 3248
rect 23178 3168 23179 3232
rect 23243 3168 23244 3232
rect 23178 3152 23244 3168
rect 23178 3088 23179 3152
rect 23243 3088 23244 3152
rect 23178 3072 23244 3088
rect 23178 3008 23179 3072
rect 23243 3008 23244 3072
rect 23178 2992 23244 3008
rect 23178 2928 23179 2992
rect 23243 2928 23244 2992
rect 23178 2838 23244 2928
rect 23304 2774 23364 3804
rect 23424 2834 23484 3866
rect 23544 2774 23604 3804
rect 23664 2834 23724 3866
rect 23784 3712 23850 3866
rect 23784 3648 23785 3712
rect 23849 3648 23850 3712
rect 23784 3632 23850 3648
rect 23784 3568 23785 3632
rect 23849 3568 23850 3632
rect 23784 3552 23850 3568
rect 23784 3488 23785 3552
rect 23849 3488 23850 3552
rect 23784 3472 23850 3488
rect 23784 3408 23785 3472
rect 23849 3408 23850 3472
rect 23784 3392 23850 3408
rect 23784 3328 23785 3392
rect 23849 3328 23850 3392
rect 23784 3312 23850 3328
rect 23784 3248 23785 3312
rect 23849 3248 23850 3312
rect 23784 3232 23850 3248
rect 23784 3168 23785 3232
rect 23849 3168 23850 3232
rect 23784 3152 23850 3168
rect 23784 3088 23785 3152
rect 23849 3088 23850 3152
rect 23784 3072 23850 3088
rect 23784 3008 23785 3072
rect 23849 3008 23850 3072
rect 23784 2992 23850 3008
rect 23784 2928 23785 2992
rect 23849 2928 23850 2992
rect 23784 2838 23850 2928
rect 23910 2774 23970 3804
rect 24030 2834 24090 3866
rect 24150 2774 24210 3804
rect 24270 2834 24330 3866
rect 24390 3712 24456 3866
rect 24390 3648 24391 3712
rect 24455 3648 24456 3712
rect 24390 3632 24456 3648
rect 24390 3568 24391 3632
rect 24455 3568 24456 3632
rect 24390 3552 24456 3568
rect 24390 3488 24391 3552
rect 24455 3488 24456 3552
rect 24390 3472 24456 3488
rect 24390 3408 24391 3472
rect 24455 3408 24456 3472
rect 24390 3392 24456 3408
rect 24390 3328 24391 3392
rect 24455 3328 24456 3392
rect 24390 3312 24456 3328
rect 24390 3248 24391 3312
rect 24455 3248 24456 3312
rect 24390 3232 24456 3248
rect 24390 3168 24391 3232
rect 24455 3168 24456 3232
rect 24390 3152 24456 3168
rect 24390 3088 24391 3152
rect 24455 3088 24456 3152
rect 24390 3072 24456 3088
rect 24390 3008 24391 3072
rect 24455 3008 24456 3072
rect 24390 2992 24456 3008
rect 24390 2928 24391 2992
rect 24455 2928 24456 2992
rect 24390 2838 24456 2928
rect 24516 2774 24576 3804
rect 24636 2834 24696 3866
rect 24756 2774 24816 3804
rect 24876 2834 24936 3866
rect 24996 3712 25062 3866
rect 24996 3648 24997 3712
rect 25061 3648 25062 3712
rect 24996 3632 25062 3648
rect 24996 3568 24997 3632
rect 25061 3568 25062 3632
rect 24996 3552 25062 3568
rect 24996 3488 24997 3552
rect 25061 3488 25062 3552
rect 24996 3472 25062 3488
rect 24996 3408 24997 3472
rect 25061 3408 25062 3472
rect 24996 3392 25062 3408
rect 24996 3328 24997 3392
rect 25061 3328 25062 3392
rect 24996 3312 25062 3328
rect 24996 3248 24997 3312
rect 25061 3248 25062 3312
rect 24996 3232 25062 3248
rect 24996 3168 24997 3232
rect 25061 3168 25062 3232
rect 24996 3152 25062 3168
rect 24996 3088 24997 3152
rect 25061 3088 25062 3152
rect 24996 3072 25062 3088
rect 24996 3008 24997 3072
rect 25061 3008 25062 3072
rect 24996 2992 25062 3008
rect 24996 2928 24997 2992
rect 25061 2928 25062 2992
rect 24996 2838 25062 2928
rect 25122 2774 25182 3804
rect 25242 2834 25302 3866
rect 25362 2774 25422 3804
rect 25482 2834 25542 3866
rect 25602 3712 25668 3866
rect 25602 3648 25603 3712
rect 25667 3648 25668 3712
rect 25602 3632 25668 3648
rect 25602 3568 25603 3632
rect 25667 3568 25668 3632
rect 25602 3552 25668 3568
rect 25602 3488 25603 3552
rect 25667 3488 25668 3552
rect 25602 3472 25668 3488
rect 25602 3408 25603 3472
rect 25667 3408 25668 3472
rect 25602 3392 25668 3408
rect 25602 3328 25603 3392
rect 25667 3328 25668 3392
rect 25602 3312 25668 3328
rect 25602 3248 25603 3312
rect 25667 3248 25668 3312
rect 25602 3232 25668 3248
rect 25602 3168 25603 3232
rect 25667 3168 25668 3232
rect 25602 3152 25668 3168
rect 25602 3088 25603 3152
rect 25667 3088 25668 3152
rect 25602 3072 25668 3088
rect 25602 3008 25603 3072
rect 25667 3008 25668 3072
rect 25602 2992 25668 3008
rect 25602 2928 25603 2992
rect 25667 2928 25668 2992
rect 25602 2838 25668 2928
rect 25728 2774 25788 3804
rect 25848 2834 25908 3866
rect 25968 2774 26028 3804
rect 26088 2834 26148 3866
rect 26208 3712 26274 3866
rect 26208 3648 26209 3712
rect 26273 3648 26274 3712
rect 26208 3632 26274 3648
rect 26208 3568 26209 3632
rect 26273 3568 26274 3632
rect 26208 3552 26274 3568
rect 26208 3488 26209 3552
rect 26273 3488 26274 3552
rect 26208 3472 26274 3488
rect 26208 3408 26209 3472
rect 26273 3408 26274 3472
rect 26208 3392 26274 3408
rect 26208 3328 26209 3392
rect 26273 3328 26274 3392
rect 26208 3312 26274 3328
rect 26208 3248 26209 3312
rect 26273 3248 26274 3312
rect 26208 3232 26274 3248
rect 26208 3168 26209 3232
rect 26273 3168 26274 3232
rect 26208 3152 26274 3168
rect 26208 3088 26209 3152
rect 26273 3088 26274 3152
rect 26208 3072 26274 3088
rect 26208 3008 26209 3072
rect 26273 3008 26274 3072
rect 26208 2992 26274 3008
rect 26208 2928 26209 2992
rect 26273 2928 26274 2992
rect 26208 2838 26274 2928
rect 26334 2774 26394 3804
rect 26454 2834 26514 3866
rect 26574 2774 26634 3804
rect 26694 2834 26754 3866
rect 26814 3712 26880 3866
rect 26814 3648 26815 3712
rect 26879 3648 26880 3712
rect 26814 3632 26880 3648
rect 26814 3568 26815 3632
rect 26879 3568 26880 3632
rect 26814 3552 26880 3568
rect 26814 3488 26815 3552
rect 26879 3488 26880 3552
rect 26814 3472 26880 3488
rect 26814 3408 26815 3472
rect 26879 3408 26880 3472
rect 26814 3392 26880 3408
rect 26814 3328 26815 3392
rect 26879 3328 26880 3392
rect 26814 3312 26880 3328
rect 26814 3248 26815 3312
rect 26879 3248 26880 3312
rect 26814 3232 26880 3248
rect 26814 3168 26815 3232
rect 26879 3168 26880 3232
rect 26814 3152 26880 3168
rect 26814 3088 26815 3152
rect 26879 3088 26880 3152
rect 26814 3072 26880 3088
rect 26814 3008 26815 3072
rect 26879 3008 26880 3072
rect 26814 2992 26880 3008
rect 26814 2928 26815 2992
rect 26879 2928 26880 2992
rect 26814 2838 26880 2928
rect 26940 2774 27000 3804
rect 27060 2834 27120 3866
rect 27180 2774 27240 3804
rect 27300 2834 27360 3866
rect 27420 3712 27486 3866
rect 27420 3648 27421 3712
rect 27485 3648 27486 3712
rect 27420 3632 27486 3648
rect 27420 3568 27421 3632
rect 27485 3568 27486 3632
rect 27420 3552 27486 3568
rect 27420 3488 27421 3552
rect 27485 3488 27486 3552
rect 27420 3472 27486 3488
rect 27420 3408 27421 3472
rect 27485 3408 27486 3472
rect 27420 3392 27486 3408
rect 27420 3328 27421 3392
rect 27485 3328 27486 3392
rect 27420 3312 27486 3328
rect 27420 3248 27421 3312
rect 27485 3248 27486 3312
rect 27420 3232 27486 3248
rect 27420 3168 27421 3232
rect 27485 3168 27486 3232
rect 27420 3152 27486 3168
rect 27420 3088 27421 3152
rect 27485 3088 27486 3152
rect 27420 3072 27486 3088
rect 27420 3008 27421 3072
rect 27485 3008 27486 3072
rect 27420 2992 27486 3008
rect 27420 2928 27421 2992
rect 27485 2928 27486 2992
rect 27420 2838 27486 2928
rect 27546 2774 27606 3804
rect 27666 2834 27726 3866
rect 27786 2774 27846 3804
rect 27906 2834 27966 3866
rect 28026 3712 28092 3866
rect 28026 3648 28027 3712
rect 28091 3648 28092 3712
rect 28026 3632 28092 3648
rect 28026 3568 28027 3632
rect 28091 3568 28092 3632
rect 28026 3552 28092 3568
rect 28026 3488 28027 3552
rect 28091 3488 28092 3552
rect 28026 3472 28092 3488
rect 28026 3408 28027 3472
rect 28091 3408 28092 3472
rect 28026 3392 28092 3408
rect 28026 3328 28027 3392
rect 28091 3328 28092 3392
rect 28026 3312 28092 3328
rect 28026 3248 28027 3312
rect 28091 3248 28092 3312
rect 28026 3232 28092 3248
rect 28026 3168 28027 3232
rect 28091 3168 28092 3232
rect 28026 3152 28092 3168
rect 28026 3088 28027 3152
rect 28091 3088 28092 3152
rect 28026 3072 28092 3088
rect 28026 3008 28027 3072
rect 28091 3008 28092 3072
rect 28026 2992 28092 3008
rect 28026 2928 28027 2992
rect 28091 2928 28092 2992
rect 28026 2838 28092 2928
rect 28152 2774 28212 3804
rect 28272 2834 28332 3866
rect 28392 2774 28452 3804
rect 28512 2834 28572 3866
rect 28632 3712 28698 3866
rect 28632 3648 28633 3712
rect 28697 3648 28698 3712
rect 28632 3632 28698 3648
rect 28632 3568 28633 3632
rect 28697 3568 28698 3632
rect 28632 3552 28698 3568
rect 28632 3488 28633 3552
rect 28697 3488 28698 3552
rect 28632 3472 28698 3488
rect 28632 3408 28633 3472
rect 28697 3408 28698 3472
rect 28632 3392 28698 3408
rect 28632 3328 28633 3392
rect 28697 3328 28698 3392
rect 28632 3312 28698 3328
rect 28632 3248 28633 3312
rect 28697 3248 28698 3312
rect 28632 3232 28698 3248
rect 28632 3168 28633 3232
rect 28697 3168 28698 3232
rect 28632 3152 28637 3168
rect 28693 3152 28698 3168
rect 28632 3088 28633 3152
rect 28697 3088 28698 3152
rect 28632 3072 28698 3088
rect 28632 3008 28633 3072
rect 28697 3008 28698 3072
rect 28632 2992 28698 3008
rect 28632 2928 28633 2992
rect 28697 2928 28698 2992
rect 28632 2838 28698 2928
rect 28758 2774 28818 3804
rect 28878 2834 28938 3866
rect 28998 2774 29058 3804
rect 29118 2834 29178 3866
rect 29238 3712 29304 3866
rect 29238 3648 29239 3712
rect 29303 3648 29304 3712
rect 29238 3632 29304 3648
rect 29238 3568 29239 3632
rect 29303 3568 29304 3632
rect 29238 3552 29304 3568
rect 29238 3488 29239 3552
rect 29303 3488 29304 3552
rect 29238 3472 29304 3488
rect 29238 3408 29239 3472
rect 29303 3408 29304 3472
rect 29238 3392 29304 3408
rect 29238 3328 29239 3392
rect 29303 3328 29304 3392
rect 29238 3312 29304 3328
rect 29238 3248 29239 3312
rect 29303 3248 29304 3312
rect 29238 3232 29304 3248
rect 29238 3168 29239 3232
rect 29303 3168 29304 3232
rect 29238 3152 29304 3168
rect 29238 3088 29239 3152
rect 29303 3088 29304 3152
rect 29238 3072 29304 3088
rect 29238 3008 29239 3072
rect 29303 3008 29304 3072
rect 29238 2992 29304 3008
rect 29238 2928 29239 2992
rect 29303 2928 29304 2992
rect 29238 2838 29304 2928
rect 29364 2774 29424 3804
rect 29484 2834 29544 3866
rect 29604 2774 29664 3804
rect 29724 2834 29784 3866
rect 29844 3712 29910 3866
rect 29844 3648 29845 3712
rect 29909 3648 29910 3712
rect 29844 3632 29910 3648
rect 29844 3568 29845 3632
rect 29909 3568 29910 3632
rect 29844 3552 29910 3568
rect 29844 3488 29845 3552
rect 29909 3488 29910 3552
rect 29844 3472 29910 3488
rect 29844 3408 29845 3472
rect 29909 3408 29910 3472
rect 29844 3392 29910 3408
rect 29844 3328 29845 3392
rect 29909 3328 29910 3392
rect 29844 3312 29910 3328
rect 29844 3248 29845 3312
rect 29909 3248 29910 3312
rect 29844 3232 29910 3248
rect 29844 3168 29845 3232
rect 29909 3168 29910 3232
rect 29844 3152 29910 3168
rect 29844 3088 29845 3152
rect 29909 3088 29910 3152
rect 29844 3072 29910 3088
rect 29844 3008 29845 3072
rect 29909 3008 29910 3072
rect 29844 2992 29910 3008
rect 29844 2928 29845 2992
rect 29909 2928 29910 2992
rect 29844 2838 29910 2928
rect 29970 2774 30030 3804
rect 30090 2834 30150 3866
rect 30210 2774 30270 3804
rect 30330 2834 30390 3866
rect 30450 3712 30516 3866
rect 30450 3648 30451 3712
rect 30515 3648 30516 3712
rect 30450 3632 30516 3648
rect 30450 3568 30451 3632
rect 30515 3568 30516 3632
rect 30450 3552 30516 3568
rect 30450 3488 30451 3552
rect 30515 3488 30516 3552
rect 30450 3472 30516 3488
rect 30450 3408 30451 3472
rect 30515 3408 30516 3472
rect 30450 3392 30516 3408
rect 30450 3328 30451 3392
rect 30515 3328 30516 3392
rect 30450 3312 30516 3328
rect 30450 3248 30451 3312
rect 30515 3248 30516 3312
rect 30450 3232 30516 3248
rect 30450 3168 30451 3232
rect 30515 3168 30516 3232
rect 30450 3152 30516 3168
rect 30450 3088 30451 3152
rect 30515 3088 30516 3152
rect 30450 3072 30516 3088
rect 30450 3008 30451 3072
rect 30515 3008 30516 3072
rect 30450 2992 30516 3008
rect 30450 2928 30451 2992
rect 30515 2928 30516 2992
rect 30450 2838 30516 2928
rect 30576 2774 30636 3804
rect 30696 2834 30756 3866
rect 30816 2774 30876 3804
rect 30936 2834 30996 3866
rect 31056 3712 31122 3866
rect 31056 3648 31057 3712
rect 31121 3648 31122 3712
rect 31056 3632 31122 3648
rect 31056 3568 31057 3632
rect 31121 3568 31122 3632
rect 31056 3552 31122 3568
rect 31056 3488 31057 3552
rect 31121 3488 31122 3552
rect 31056 3472 31122 3488
rect 31056 3408 31057 3472
rect 31121 3408 31122 3472
rect 31056 3392 31122 3408
rect 31056 3328 31057 3392
rect 31121 3328 31122 3392
rect 31056 3312 31122 3328
rect 31056 3248 31057 3312
rect 31121 3248 31122 3312
rect 31056 3232 31122 3248
rect 31056 3168 31057 3232
rect 31121 3168 31122 3232
rect 31056 3152 31122 3168
rect 31056 3088 31057 3152
rect 31121 3088 31122 3152
rect 31056 3072 31122 3088
rect 31056 3008 31057 3072
rect 31121 3008 31122 3072
rect 31056 2992 31122 3008
rect 31056 2928 31057 2992
rect 31121 2928 31122 2992
rect 31056 2838 31122 2928
rect 31182 2774 31242 3804
rect 31302 2834 31362 3866
rect 31422 2774 31482 3804
rect 31542 2834 31602 3866
rect 31662 3712 31728 3866
rect 31662 3648 31663 3712
rect 31727 3648 31728 3712
rect 31662 3632 31728 3648
rect 31662 3568 31663 3632
rect 31727 3568 31728 3632
rect 31662 3552 31728 3568
rect 31662 3488 31663 3552
rect 31727 3488 31728 3552
rect 31662 3472 31728 3488
rect 31662 3408 31663 3472
rect 31727 3408 31728 3472
rect 31662 3392 31728 3408
rect 31662 3328 31663 3392
rect 31727 3328 31728 3392
rect 31662 3312 31728 3328
rect 31662 3248 31663 3312
rect 31727 3248 31728 3312
rect 31662 3232 31728 3248
rect 31662 3168 31663 3232
rect 31727 3168 31728 3232
rect 31662 3152 31728 3168
rect 31662 3088 31663 3152
rect 31727 3088 31728 3152
rect 31662 3072 31728 3088
rect 31662 3008 31663 3072
rect 31727 3008 31728 3072
rect 31662 2992 31728 3008
rect 31662 2928 31663 2992
rect 31727 2928 31728 2992
rect 31662 2838 31728 2928
rect 31788 2774 31848 3804
rect 31908 2834 31968 3866
rect 32028 2774 32088 3804
rect 32148 2834 32208 3866
rect 32268 3712 32334 3866
rect 32268 3648 32269 3712
rect 32333 3648 32334 3712
rect 32268 3632 32334 3648
rect 32268 3568 32269 3632
rect 32333 3568 32334 3632
rect 32268 3552 32334 3568
rect 32268 3488 32269 3552
rect 32333 3488 32334 3552
rect 32268 3472 32334 3488
rect 32268 3408 32269 3472
rect 32333 3408 32334 3472
rect 32268 3392 32334 3408
rect 32268 3328 32269 3392
rect 32333 3328 32334 3392
rect 32268 3312 32334 3328
rect 32268 3248 32269 3312
rect 32333 3248 32334 3312
rect 32268 3232 32334 3248
rect 32268 3168 32269 3232
rect 32333 3168 32334 3232
rect 32268 3152 32334 3168
rect 32268 3088 32269 3152
rect 32333 3088 32334 3152
rect 32268 3072 32334 3088
rect 32268 3008 32269 3072
rect 32333 3008 32334 3072
rect 32268 2992 32334 3008
rect 32268 2928 32269 2992
rect 32333 2928 32334 2992
rect 32268 2838 32334 2928
rect 32394 2774 32454 3804
rect 32514 2834 32574 3866
rect 32634 2774 32694 3804
rect 32754 2834 32814 3866
rect 32874 3712 32940 3866
rect 32874 3648 32875 3712
rect 32939 3648 32940 3712
rect 32874 3632 32940 3648
rect 32874 3568 32875 3632
rect 32939 3568 32940 3632
rect 32874 3552 32940 3568
rect 32874 3488 32875 3552
rect 32939 3488 32940 3552
rect 32874 3472 32940 3488
rect 32874 3408 32875 3472
rect 32939 3408 32940 3472
rect 32874 3392 32940 3408
rect 32874 3328 32875 3392
rect 32939 3328 32940 3392
rect 32874 3312 32940 3328
rect 32874 3248 32875 3312
rect 32939 3248 32940 3312
rect 32874 3232 32940 3248
rect 32874 3168 32875 3232
rect 32939 3168 32940 3232
rect 32874 3152 32940 3168
rect 32874 3088 32875 3152
rect 32939 3088 32940 3152
rect 32874 3072 32940 3088
rect 32874 3008 32875 3072
rect 32939 3008 32940 3072
rect 32874 2992 32940 3008
rect 32874 2928 32875 2992
rect 32939 2928 32940 2992
rect 32874 2838 32940 2928
rect 33000 2774 33060 3804
rect 33120 2834 33180 3866
rect 33240 2774 33300 3804
rect 33360 2834 33420 3866
rect 33480 3712 33546 3866
rect 33480 3648 33481 3712
rect 33545 3648 33546 3712
rect 33480 3632 33546 3648
rect 33480 3568 33481 3632
rect 33545 3568 33546 3632
rect 33480 3552 33546 3568
rect 33480 3488 33481 3552
rect 33545 3488 33546 3552
rect 33480 3472 33546 3488
rect 33480 3408 33481 3472
rect 33545 3408 33546 3472
rect 33480 3392 33546 3408
rect 33480 3328 33481 3392
rect 33545 3328 33546 3392
rect 33480 3312 33546 3328
rect 33480 3248 33481 3312
rect 33545 3248 33546 3312
rect 33480 3232 33546 3248
rect 33480 3168 33481 3232
rect 33545 3168 33546 3232
rect 33480 3152 33546 3168
rect 33480 3088 33481 3152
rect 33545 3088 33546 3152
rect 33480 3072 33546 3088
rect 33480 3008 33481 3072
rect 33545 3008 33546 3072
rect 33480 2992 33546 3008
rect 33480 2928 33481 2992
rect 33545 2928 33546 2992
rect 33480 2838 33546 2928
rect 33606 2774 33666 3804
rect 33726 2834 33786 3866
rect 33846 2774 33906 3804
rect 33966 2834 34026 3866
rect 34086 3712 34152 3866
rect 34086 3648 34087 3712
rect 34151 3648 34152 3712
rect 34086 3632 34152 3648
rect 34086 3568 34087 3632
rect 34151 3568 34152 3632
rect 34086 3552 34152 3568
rect 34086 3488 34087 3552
rect 34151 3488 34152 3552
rect 34086 3472 34152 3488
rect 34086 3408 34087 3472
rect 34151 3408 34152 3472
rect 34086 3392 34152 3408
rect 34086 3328 34087 3392
rect 34151 3328 34152 3392
rect 34086 3312 34152 3328
rect 34086 3248 34087 3312
rect 34151 3248 34152 3312
rect 34086 3232 34152 3248
rect 34086 3168 34087 3232
rect 34151 3168 34152 3232
rect 34086 3152 34152 3168
rect 34086 3088 34087 3152
rect 34151 3088 34152 3152
rect 34086 3072 34152 3088
rect 34086 3008 34087 3072
rect 34151 3008 34152 3072
rect 34086 2992 34152 3008
rect 34086 2928 34087 2992
rect 34151 2928 34152 2992
rect 34086 2838 34152 2928
rect 34212 2774 34272 3804
rect 34332 2834 34392 3866
rect 34452 2774 34512 3804
rect 34572 2834 34632 3866
rect 34692 3712 34758 3866
rect 34692 3648 34693 3712
rect 34757 3648 34758 3712
rect 34692 3632 34758 3648
rect 34692 3568 34693 3632
rect 34757 3568 34758 3632
rect 34692 3552 34758 3568
rect 34692 3488 34693 3552
rect 34757 3488 34758 3552
rect 34692 3472 34758 3488
rect 34692 3408 34693 3472
rect 34757 3408 34758 3472
rect 34692 3392 34758 3408
rect 34692 3328 34693 3392
rect 34757 3328 34758 3392
rect 34692 3312 34758 3328
rect 34692 3248 34693 3312
rect 34757 3248 34758 3312
rect 34692 3232 34758 3248
rect 34692 3168 34693 3232
rect 34757 3168 34758 3232
rect 34692 3152 34758 3168
rect 34692 3088 34693 3152
rect 34757 3088 34758 3152
rect 34692 3072 34758 3088
rect 34692 3008 34693 3072
rect 34757 3008 34758 3072
rect 34692 2992 34758 3008
rect 34692 2928 34693 2992
rect 34757 2928 34758 2992
rect 34692 2838 34758 2928
rect 34818 2774 34878 3804
rect 34938 2834 34998 3866
rect 35058 2774 35118 3804
rect 35178 2834 35238 3866
rect 35298 3712 35364 3866
rect 35298 3648 35299 3712
rect 35363 3648 35364 3712
rect 35298 3632 35364 3648
rect 35298 3568 35299 3632
rect 35363 3568 35364 3632
rect 35298 3552 35364 3568
rect 35298 3488 35299 3552
rect 35363 3488 35364 3552
rect 35298 3472 35364 3488
rect 35298 3408 35299 3472
rect 35363 3408 35364 3472
rect 35298 3392 35364 3408
rect 35298 3328 35299 3392
rect 35363 3328 35364 3392
rect 35298 3312 35364 3328
rect 35298 3248 35299 3312
rect 35363 3248 35364 3312
rect 35298 3232 35364 3248
rect 35298 3168 35299 3232
rect 35363 3168 35364 3232
rect 35298 3152 35364 3168
rect 35298 3088 35299 3152
rect 35363 3088 35364 3152
rect 35298 3072 35364 3088
rect 35298 3008 35299 3072
rect 35363 3008 35364 3072
rect 35298 2992 35364 3008
rect 35298 2928 35299 2992
rect 35363 2928 35364 2992
rect 35298 2838 35364 2928
rect 35424 2774 35484 3804
rect 35544 2834 35604 3866
rect 35664 2774 35724 3804
rect 35784 2834 35844 3866
rect 35904 3712 35970 3866
rect 35904 3648 35905 3712
rect 35969 3648 35970 3712
rect 35904 3632 35970 3648
rect 35904 3568 35905 3632
rect 35969 3568 35970 3632
rect 35904 3552 35970 3568
rect 35904 3488 35905 3552
rect 35969 3488 35970 3552
rect 35904 3472 35970 3488
rect 35904 3408 35905 3472
rect 35969 3408 35970 3472
rect 35904 3392 35970 3408
rect 35904 3328 35905 3392
rect 35969 3328 35970 3392
rect 35904 3312 35970 3328
rect 35904 3248 35905 3312
rect 35969 3248 35970 3312
rect 35904 3232 35970 3248
rect 35904 3168 35905 3232
rect 35969 3168 35970 3232
rect 35904 3152 35970 3168
rect 35904 3088 35905 3152
rect 35969 3088 35970 3152
rect 35904 3072 35970 3088
rect 35904 3008 35905 3072
rect 35969 3008 35970 3072
rect 35904 2992 35970 3008
rect 35904 2928 35905 2992
rect 35969 2928 35970 2992
rect 35904 2838 35970 2928
rect 36030 2774 36090 3804
rect 36150 2834 36210 3866
rect 36270 2774 36330 3804
rect 36390 2834 36450 3866
rect 36510 3712 36576 3866
rect 36510 3648 36511 3712
rect 36575 3648 36576 3712
rect 36510 3632 36576 3648
rect 36510 3568 36511 3632
rect 36575 3568 36576 3632
rect 36510 3552 36576 3568
rect 36510 3488 36511 3552
rect 36575 3488 36576 3552
rect 36510 3472 36576 3488
rect 36510 3408 36511 3472
rect 36575 3408 36576 3472
rect 36510 3392 36576 3408
rect 36510 3328 36511 3392
rect 36575 3328 36576 3392
rect 36510 3312 36576 3328
rect 36510 3248 36511 3312
rect 36575 3248 36576 3312
rect 36510 3232 36576 3248
rect 36510 3168 36511 3232
rect 36575 3168 36576 3232
rect 36510 3152 36576 3168
rect 36510 3088 36511 3152
rect 36575 3088 36576 3152
rect 36510 3072 36576 3088
rect 36510 3008 36511 3072
rect 36575 3008 36576 3072
rect 36510 2992 36576 3008
rect 36510 2928 36511 2992
rect 36575 2928 36576 2992
rect 36510 2838 36576 2928
rect 36636 2774 36696 3804
rect 36756 2834 36816 3866
rect 36876 2774 36936 3804
rect 36996 2834 37056 3866
rect 37116 3712 37182 3866
rect 37116 3648 37117 3712
rect 37181 3648 37182 3712
rect 37116 3632 37182 3648
rect 37116 3568 37117 3632
rect 37181 3568 37182 3632
rect 37116 3552 37182 3568
rect 37116 3488 37117 3552
rect 37181 3488 37182 3552
rect 37116 3472 37182 3488
rect 37116 3408 37117 3472
rect 37181 3408 37182 3472
rect 37116 3392 37182 3408
rect 37116 3328 37117 3392
rect 37181 3328 37182 3392
rect 37116 3312 37182 3328
rect 37116 3248 37117 3312
rect 37181 3248 37182 3312
rect 37116 3232 37182 3248
rect 37116 3168 37117 3232
rect 37181 3168 37182 3232
rect 37116 3152 37182 3168
rect 37116 3088 37117 3152
rect 37181 3088 37182 3152
rect 37116 3072 37182 3088
rect 37116 3008 37117 3072
rect 37181 3008 37182 3072
rect 37116 2992 37182 3008
rect 37116 2928 37117 2992
rect 37181 2928 37182 2992
rect 37116 2838 37182 2928
rect 37242 2774 37302 3804
rect 37362 2834 37422 3866
rect 37482 2774 37542 3804
rect 37602 2834 37662 3866
rect 37722 3712 37788 3866
rect 37722 3648 37723 3712
rect 37787 3648 37788 3712
rect 37722 3632 37788 3648
rect 37722 3568 37723 3632
rect 37787 3568 37788 3632
rect 37722 3552 37788 3568
rect 37722 3488 37723 3552
rect 37787 3488 37788 3552
rect 37722 3472 37788 3488
rect 37722 3408 37723 3472
rect 37787 3408 37788 3472
rect 37722 3392 37788 3408
rect 37722 3328 37723 3392
rect 37787 3328 37788 3392
rect 37722 3312 37788 3328
rect 37722 3248 37723 3312
rect 37787 3248 37788 3312
rect 37722 3232 37788 3248
rect 37722 3168 37723 3232
rect 37787 3168 37788 3232
rect 37722 3152 37788 3168
rect 37722 3088 37723 3152
rect 37787 3088 37788 3152
rect 37722 3072 37788 3088
rect 37722 3008 37723 3072
rect 37787 3008 37788 3072
rect 37722 2992 37788 3008
rect 37722 2928 37723 2992
rect 37787 2928 37788 2992
rect 37722 2838 37788 2928
rect 37848 2774 37908 3804
rect 37968 2834 38028 3866
rect 38088 2774 38148 3804
rect 38208 2834 38268 3866
rect 38328 3712 38394 3866
rect 38328 3648 38329 3712
rect 38393 3648 38394 3712
rect 38328 3632 38394 3648
rect 38328 3568 38329 3632
rect 38393 3568 38394 3632
rect 38328 3552 38394 3568
rect 38328 3488 38329 3552
rect 38393 3488 38394 3552
rect 38328 3472 38394 3488
rect 38328 3408 38329 3472
rect 38393 3408 38394 3472
rect 38328 3392 38394 3408
rect 38328 3328 38329 3392
rect 38393 3328 38394 3392
rect 38328 3312 38394 3328
rect 38328 3248 38329 3312
rect 38393 3248 38394 3312
rect 38328 3232 38394 3248
rect 38328 3168 38329 3232
rect 38393 3168 38394 3232
rect 38328 3152 38394 3168
rect 38328 3088 38329 3152
rect 38393 3088 38394 3152
rect 38328 3072 38394 3088
rect 38328 3008 38329 3072
rect 38393 3008 38394 3072
rect 38328 2992 38394 3008
rect 38328 2928 38329 2992
rect 38393 2928 38394 2992
rect 38328 2838 38394 2928
rect 38454 2774 38514 3804
rect 38574 2834 38634 3866
rect 38694 2774 38754 3804
rect 38814 2834 38874 3866
rect 38934 3712 39000 3866
rect 38934 3648 38935 3712
rect 38999 3648 39000 3712
rect 38934 3632 39000 3648
rect 38934 3568 38935 3632
rect 38999 3568 39000 3632
rect 38934 3552 39000 3568
rect 38934 3488 38935 3552
rect 38999 3488 39000 3552
rect 38934 3472 39000 3488
rect 38934 3408 38935 3472
rect 38999 3408 39000 3472
rect 38934 3392 39000 3408
rect 38934 3328 38935 3392
rect 38999 3328 39000 3392
rect 38934 3312 39000 3328
rect 38934 3248 38935 3312
rect 38999 3248 39000 3312
rect 38934 3232 39000 3248
rect 38934 3168 38935 3232
rect 38999 3168 39000 3232
rect 38934 3152 39000 3168
rect 38934 3088 38935 3152
rect 38999 3088 39000 3152
rect 38934 3072 39000 3088
rect 38934 3008 38935 3072
rect 38999 3008 39000 3072
rect 38934 2992 39000 3008
rect 38934 2928 38935 2992
rect 38999 2928 39000 2992
rect 38934 2838 39000 2928
rect 39060 2774 39120 3804
rect 39180 2834 39240 3866
rect 39300 2774 39360 3804
rect 39420 2834 39480 3866
rect 39540 3712 39606 3866
rect 39540 3648 39541 3712
rect 39605 3648 39606 3712
rect 39540 3632 39606 3648
rect 39540 3568 39541 3632
rect 39605 3568 39606 3632
rect 39540 3552 39606 3568
rect 39540 3488 39541 3552
rect 39605 3488 39606 3552
rect 39540 3472 39606 3488
rect 39540 3408 39541 3472
rect 39605 3408 39606 3472
rect 39540 3392 39606 3408
rect 39540 3328 39541 3392
rect 39605 3328 39606 3392
rect 39540 3312 39606 3328
rect 39540 3248 39541 3312
rect 39605 3248 39606 3312
rect 39540 3232 39606 3248
rect 39540 3168 39541 3232
rect 39605 3168 39606 3232
rect 39540 3152 39606 3168
rect 39540 3088 39541 3152
rect 39605 3088 39606 3152
rect 39540 3072 39606 3088
rect 39540 3008 39541 3072
rect 39605 3008 39606 3072
rect 39540 2992 39606 3008
rect 39540 2928 39541 2992
rect 39605 2928 39606 2992
rect 39540 2838 39606 2928
rect -459 2772 213 2774
rect -459 2708 -355 2772
rect -291 2708 -275 2772
rect -211 2708 -195 2772
rect -131 2708 -115 2772
rect -51 2708 -35 2772
rect 29 2708 45 2772
rect 109 2708 213 2772
rect -459 2706 213 2708
rect 355 2772 1027 2774
rect 355 2708 459 2772
rect 523 2708 539 2772
rect 603 2708 619 2772
rect 683 2708 699 2772
rect 763 2708 779 2772
rect 843 2708 859 2772
rect 923 2708 1027 2772
rect 355 2706 1027 2708
rect 1267 2772 2545 2774
rect 1267 2708 1371 2772
rect 1435 2708 1451 2772
rect 1515 2708 1531 2772
rect 1595 2708 1611 2772
rect 1675 2708 1691 2772
rect 1755 2708 1771 2772
rect 1835 2708 1977 2772
rect 2041 2708 2057 2772
rect 2121 2708 2137 2772
rect 2201 2708 2217 2772
rect 2281 2708 2297 2772
rect 2361 2708 2377 2772
rect 2441 2708 2545 2772
rect 1267 2706 2545 2708
rect 2801 2772 5291 2774
rect 2801 2708 2905 2772
rect 2969 2708 2985 2772
rect 3049 2708 3065 2772
rect 3129 2708 3145 2772
rect 3209 2708 3225 2772
rect 3289 2708 3305 2772
rect 3369 2708 3511 2772
rect 3575 2708 3591 2772
rect 3655 2708 3671 2772
rect 3735 2708 3751 2772
rect 3815 2708 3831 2772
rect 3895 2708 3911 2772
rect 3975 2708 4117 2772
rect 4181 2708 4197 2772
rect 4261 2708 4277 2772
rect 4341 2708 4357 2772
rect 4421 2708 4437 2772
rect 4501 2708 4517 2772
rect 4581 2708 4723 2772
rect 4787 2708 4803 2772
rect 4867 2708 4883 2772
rect 4947 2708 4963 2772
rect 5027 2708 5043 2772
rect 5107 2708 5123 2772
rect 5187 2708 5291 2772
rect 2801 2706 5291 2708
rect 5352 2772 10266 2774
rect 5352 2708 5456 2772
rect 5520 2708 5536 2772
rect 5600 2708 5616 2772
rect 5680 2708 5696 2772
rect 5760 2708 5776 2772
rect 5840 2708 5856 2772
rect 5920 2708 6062 2772
rect 6126 2708 6142 2772
rect 6206 2708 6222 2772
rect 6286 2708 6302 2772
rect 6366 2708 6382 2772
rect 6446 2708 6462 2772
rect 6526 2708 6668 2772
rect 6732 2708 6748 2772
rect 6812 2708 6828 2772
rect 6892 2708 6908 2772
rect 6972 2708 6988 2772
rect 7052 2708 7068 2772
rect 7132 2708 7274 2772
rect 7338 2708 7354 2772
rect 7418 2708 7434 2772
rect 7498 2708 7514 2772
rect 7578 2708 7594 2772
rect 7658 2708 7674 2772
rect 7738 2708 7880 2772
rect 7944 2708 7960 2772
rect 8024 2708 8040 2772
rect 8104 2708 8120 2772
rect 8184 2708 8200 2772
rect 8264 2708 8280 2772
rect 8344 2708 8486 2772
rect 8550 2708 8566 2772
rect 8630 2708 8646 2772
rect 8710 2708 8726 2772
rect 8790 2708 8806 2772
rect 8870 2708 8886 2772
rect 8950 2708 9092 2772
rect 9156 2708 9172 2772
rect 9236 2708 9252 2772
rect 9316 2708 9332 2772
rect 9396 2708 9412 2772
rect 9476 2708 9492 2772
rect 9556 2708 9698 2772
rect 9762 2708 9778 2772
rect 9842 2708 9858 2772
rect 9922 2708 9938 2772
rect 10002 2708 10018 2772
rect 10082 2708 10098 2772
rect 10162 2708 10266 2772
rect 5352 2706 10266 2708
rect 10326 2772 20088 2774
rect 10326 2708 10430 2772
rect 10494 2708 10510 2772
rect 10574 2708 10590 2772
rect 10654 2708 10670 2772
rect 10734 2708 10750 2772
rect 10814 2708 10830 2772
rect 10894 2708 11036 2772
rect 11100 2708 11116 2772
rect 11180 2708 11196 2772
rect 11260 2708 11276 2772
rect 11340 2708 11356 2772
rect 11420 2708 11436 2772
rect 11500 2708 11642 2772
rect 11706 2708 11722 2772
rect 11786 2708 11802 2772
rect 11866 2708 11882 2772
rect 11946 2708 11962 2772
rect 12026 2708 12042 2772
rect 12106 2708 12248 2772
rect 12312 2708 12328 2772
rect 12392 2708 12408 2772
rect 12472 2708 12488 2772
rect 12552 2708 12568 2772
rect 12632 2708 12648 2772
rect 12712 2708 12854 2772
rect 12918 2708 12934 2772
rect 12998 2708 13014 2772
rect 13078 2708 13094 2772
rect 13158 2708 13174 2772
rect 13238 2708 13254 2772
rect 13318 2708 13460 2772
rect 13524 2708 13540 2772
rect 13604 2708 13620 2772
rect 13684 2708 13700 2772
rect 13764 2708 13780 2772
rect 13844 2708 13860 2772
rect 13924 2708 14066 2772
rect 14130 2708 14146 2772
rect 14210 2708 14226 2772
rect 14290 2708 14306 2772
rect 14370 2708 14386 2772
rect 14450 2708 14466 2772
rect 14530 2708 14672 2772
rect 14736 2708 14752 2772
rect 14816 2708 14832 2772
rect 14896 2708 14912 2772
rect 14976 2708 14992 2772
rect 15056 2708 15072 2772
rect 15136 2708 15278 2772
rect 15342 2708 15358 2772
rect 15422 2708 15438 2772
rect 15502 2708 15518 2772
rect 15582 2708 15598 2772
rect 15662 2708 15678 2772
rect 15742 2708 15884 2772
rect 15948 2708 15964 2772
rect 16028 2708 16044 2772
rect 16108 2708 16124 2772
rect 16188 2708 16204 2772
rect 16268 2708 16284 2772
rect 16348 2708 16490 2772
rect 16554 2708 16570 2772
rect 16634 2708 16650 2772
rect 16714 2708 16730 2772
rect 16794 2708 16810 2772
rect 16874 2708 16890 2772
rect 16954 2708 17096 2772
rect 17160 2708 17176 2772
rect 17240 2708 17256 2772
rect 17320 2708 17336 2772
rect 17400 2708 17416 2772
rect 17480 2708 17496 2772
rect 17560 2708 17702 2772
rect 17766 2708 17782 2772
rect 17846 2708 17862 2772
rect 17926 2708 17942 2772
rect 18006 2708 18022 2772
rect 18086 2708 18102 2772
rect 18166 2708 18308 2772
rect 18372 2708 18388 2772
rect 18452 2708 18468 2772
rect 18532 2708 18548 2772
rect 18612 2708 18628 2772
rect 18692 2708 18708 2772
rect 18772 2708 18914 2772
rect 18978 2708 18994 2772
rect 19058 2708 19074 2772
rect 19138 2708 19154 2772
rect 19218 2708 19234 2772
rect 19298 2708 19314 2772
rect 19378 2708 19520 2772
rect 19584 2708 19600 2772
rect 19664 2708 19680 2772
rect 19744 2708 19760 2772
rect 19824 2708 19840 2772
rect 19904 2708 19920 2772
rect 19984 2708 20088 2772
rect 10326 2706 20088 2708
rect 20148 2772 39606 2774
rect 20148 2708 20252 2772
rect 20316 2708 20332 2772
rect 20396 2708 20412 2772
rect 20476 2708 20492 2772
rect 20556 2708 20572 2772
rect 20636 2708 20652 2772
rect 20716 2708 20858 2772
rect 20922 2708 20938 2772
rect 21002 2708 21018 2772
rect 21082 2708 21098 2772
rect 21162 2708 21178 2772
rect 21242 2708 21258 2772
rect 21322 2708 21464 2772
rect 21528 2708 21544 2772
rect 21608 2708 21624 2772
rect 21688 2708 21704 2772
rect 21768 2708 21784 2772
rect 21848 2708 21864 2772
rect 21928 2708 22070 2772
rect 22134 2708 22150 2772
rect 22214 2708 22230 2772
rect 22294 2708 22310 2772
rect 22374 2708 22390 2772
rect 22454 2708 22470 2772
rect 22534 2708 22676 2772
rect 22740 2708 22756 2772
rect 22820 2708 22836 2772
rect 22900 2708 22916 2772
rect 22980 2708 22996 2772
rect 23060 2708 23076 2772
rect 23140 2708 23282 2772
rect 23346 2708 23362 2772
rect 23426 2708 23442 2772
rect 23506 2708 23522 2772
rect 23586 2708 23602 2772
rect 23666 2708 23682 2772
rect 23746 2708 23888 2772
rect 23952 2708 23968 2772
rect 24032 2708 24048 2772
rect 24112 2708 24128 2772
rect 24192 2708 24208 2772
rect 24272 2708 24288 2772
rect 24352 2708 24494 2772
rect 24558 2708 24574 2772
rect 24638 2708 24654 2772
rect 24718 2708 24734 2772
rect 24798 2708 24814 2772
rect 24878 2708 24894 2772
rect 24958 2708 25100 2772
rect 25164 2708 25180 2772
rect 25244 2708 25260 2772
rect 25324 2708 25340 2772
rect 25404 2708 25420 2772
rect 25484 2708 25500 2772
rect 25564 2708 25706 2772
rect 25770 2708 25786 2772
rect 25850 2708 25866 2772
rect 25930 2708 25946 2772
rect 26010 2708 26026 2772
rect 26090 2708 26106 2772
rect 26170 2708 26312 2772
rect 26376 2708 26392 2772
rect 26456 2708 26472 2772
rect 26536 2708 26552 2772
rect 26616 2708 26632 2772
rect 26696 2708 26712 2772
rect 26776 2708 26918 2772
rect 26982 2708 26998 2772
rect 27062 2708 27078 2772
rect 27142 2708 27158 2772
rect 27222 2708 27238 2772
rect 27302 2708 27318 2772
rect 27382 2708 27524 2772
rect 27588 2708 27604 2772
rect 27668 2708 27684 2772
rect 27748 2708 27764 2772
rect 27828 2708 27844 2772
rect 27908 2708 27924 2772
rect 27988 2708 28130 2772
rect 28194 2708 28210 2772
rect 28274 2708 28290 2772
rect 28354 2708 28370 2772
rect 28434 2708 28450 2772
rect 28514 2708 28530 2772
rect 28594 2708 28736 2772
rect 28800 2708 28816 2772
rect 28880 2708 28896 2772
rect 28960 2708 28976 2772
rect 29040 2708 29056 2772
rect 29120 2708 29136 2772
rect 29200 2708 29342 2772
rect 29406 2708 29422 2772
rect 29486 2708 29502 2772
rect 29566 2708 29582 2772
rect 29646 2708 29662 2772
rect 29726 2708 29742 2772
rect 29806 2708 29948 2772
rect 30012 2708 30028 2772
rect 30092 2708 30108 2772
rect 30172 2708 30188 2772
rect 30252 2708 30268 2772
rect 30332 2708 30348 2772
rect 30412 2708 30554 2772
rect 30618 2708 30634 2772
rect 30698 2708 30714 2772
rect 30778 2708 30794 2772
rect 30858 2708 30874 2772
rect 30938 2708 30954 2772
rect 31018 2708 31160 2772
rect 31224 2708 31240 2772
rect 31304 2708 31320 2772
rect 31384 2708 31400 2772
rect 31464 2708 31480 2772
rect 31544 2708 31560 2772
rect 31624 2708 31766 2772
rect 31830 2708 31846 2772
rect 31910 2708 31926 2772
rect 31990 2708 32006 2772
rect 32070 2708 32086 2772
rect 32150 2708 32166 2772
rect 32230 2708 32372 2772
rect 32436 2708 32452 2772
rect 32516 2708 32532 2772
rect 32596 2708 32612 2772
rect 32676 2708 32692 2772
rect 32756 2708 32772 2772
rect 32836 2708 32978 2772
rect 33042 2708 33058 2772
rect 33122 2708 33138 2772
rect 33202 2708 33218 2772
rect 33282 2708 33298 2772
rect 33362 2708 33378 2772
rect 33442 2708 33584 2772
rect 33648 2708 33664 2772
rect 33728 2708 33744 2772
rect 33808 2708 33824 2772
rect 33888 2708 33904 2772
rect 33968 2708 33984 2772
rect 34048 2708 34190 2772
rect 34254 2708 34270 2772
rect 34334 2708 34350 2772
rect 34414 2708 34430 2772
rect 34494 2708 34510 2772
rect 34574 2708 34590 2772
rect 34654 2708 34796 2772
rect 34860 2708 34876 2772
rect 34940 2708 34956 2772
rect 35020 2708 35036 2772
rect 35100 2708 35116 2772
rect 35180 2708 35196 2772
rect 35260 2708 35402 2772
rect 35466 2708 35482 2772
rect 35546 2708 35562 2772
rect 35626 2708 35642 2772
rect 35706 2708 35722 2772
rect 35786 2708 35802 2772
rect 35866 2708 36008 2772
rect 36072 2708 36088 2772
rect 36152 2708 36168 2772
rect 36232 2708 36248 2772
rect 36312 2708 36328 2772
rect 36392 2708 36408 2772
rect 36472 2708 36614 2772
rect 36678 2708 36694 2772
rect 36758 2708 36774 2772
rect 36838 2708 36854 2772
rect 36918 2708 36934 2772
rect 36998 2708 37014 2772
rect 37078 2708 37220 2772
rect 37284 2708 37300 2772
rect 37364 2708 37380 2772
rect 37444 2708 37460 2772
rect 37524 2708 37540 2772
rect 37604 2708 37620 2772
rect 37684 2708 37826 2772
rect 37890 2708 37906 2772
rect 37970 2708 37986 2772
rect 38050 2708 38066 2772
rect 38130 2708 38146 2772
rect 38210 2708 38226 2772
rect 38290 2708 38432 2772
rect 38496 2708 38512 2772
rect 38576 2708 38592 2772
rect 38656 2708 38672 2772
rect 38736 2708 38752 2772
rect 38816 2708 38832 2772
rect 38896 2708 39038 2772
rect 39102 2708 39118 2772
rect 39182 2708 39198 2772
rect 39262 2708 39278 2772
rect 39342 2708 39358 2772
rect 39422 2708 39438 2772
rect 39502 2708 39606 2772
rect 20148 2706 39606 2708
rect -93 2606 -33 2615
rect -459 2604 213 2606
rect -459 2540 -355 2604
rect -291 2540 -275 2604
rect -211 2540 -195 2604
rect -131 2540 -115 2604
rect -51 2600 -35 2604
rect -51 2540 -35 2544
rect 29 2540 45 2604
rect 109 2540 213 2604
rect -459 2538 213 2540
rect 355 2604 1027 2606
rect 355 2540 459 2604
rect 523 2540 539 2604
rect 603 2540 619 2604
rect 683 2540 699 2604
rect 763 2540 779 2604
rect 843 2540 859 2604
rect 923 2540 1027 2604
rect 355 2538 1027 2540
rect 1267 2604 2545 2606
rect 1267 2540 1371 2604
rect 1435 2540 1451 2604
rect 1515 2540 1531 2604
rect 1595 2540 1611 2604
rect 1675 2540 1691 2604
rect 1755 2540 1771 2604
rect 1835 2540 1977 2604
rect 2041 2540 2057 2604
rect 2121 2540 2137 2604
rect 2201 2540 2217 2604
rect 2281 2540 2297 2604
rect 2361 2540 2377 2604
rect 2441 2540 2545 2604
rect 1267 2538 2545 2540
rect 2801 2604 5291 2606
rect 2801 2540 2905 2604
rect 2969 2540 2985 2604
rect 3049 2540 3065 2604
rect 3129 2540 3145 2604
rect 3209 2540 3225 2604
rect 3289 2540 3305 2604
rect 3369 2540 3511 2604
rect 3575 2540 3591 2604
rect 3655 2540 3671 2604
rect 3735 2540 3751 2604
rect 3815 2540 3831 2604
rect 3895 2540 3911 2604
rect 3975 2540 4117 2604
rect 4181 2540 4197 2604
rect 4261 2540 4277 2604
rect 4341 2540 4357 2604
rect 4421 2540 4437 2604
rect 4501 2540 4517 2604
rect 4581 2540 4723 2604
rect 4787 2540 4803 2604
rect 4867 2540 4883 2604
rect 4947 2540 4963 2604
rect 5027 2540 5043 2604
rect 5107 2540 5123 2604
rect 5187 2540 5291 2604
rect 2801 2538 5291 2540
rect 5352 2604 10266 2606
rect 5352 2540 5456 2604
rect 5520 2540 5536 2604
rect 5600 2540 5616 2604
rect 5680 2540 5696 2604
rect 5760 2540 5776 2604
rect 5840 2540 5856 2604
rect 5920 2540 6062 2604
rect 6126 2540 6142 2604
rect 6206 2540 6222 2604
rect 6286 2540 6302 2604
rect 6366 2540 6382 2604
rect 6446 2540 6462 2604
rect 6526 2540 6668 2604
rect 6732 2540 6748 2604
rect 6812 2540 6828 2604
rect 6892 2540 6908 2604
rect 6972 2540 6988 2604
rect 7052 2540 7068 2604
rect 7132 2540 7274 2604
rect 7338 2540 7354 2604
rect 7418 2540 7434 2604
rect 7498 2540 7514 2604
rect 7578 2540 7594 2604
rect 7658 2540 7674 2604
rect 7738 2540 7880 2604
rect 7944 2540 7960 2604
rect 8024 2540 8040 2604
rect 8104 2540 8120 2604
rect 8184 2540 8200 2604
rect 8264 2540 8280 2604
rect 8344 2540 8486 2604
rect 8550 2540 8566 2604
rect 8630 2540 8646 2604
rect 8710 2540 8726 2604
rect 8790 2540 8806 2604
rect 8870 2540 8886 2604
rect 8950 2540 9092 2604
rect 9156 2540 9172 2604
rect 9236 2540 9252 2604
rect 9316 2540 9332 2604
rect 9396 2540 9412 2604
rect 9476 2540 9492 2604
rect 9556 2540 9698 2604
rect 9762 2540 9778 2604
rect 9842 2540 9858 2604
rect 9922 2540 9938 2604
rect 10002 2540 10018 2604
rect 10082 2540 10098 2604
rect 10162 2540 10266 2604
rect 5352 2538 10266 2540
rect 10326 2604 20088 2606
rect 10326 2540 10430 2604
rect 10494 2540 10510 2604
rect 10574 2540 10590 2604
rect 10654 2540 10670 2604
rect 10734 2540 10750 2604
rect 10814 2540 10830 2604
rect 10894 2540 11036 2604
rect 11100 2540 11116 2604
rect 11180 2540 11196 2604
rect 11260 2540 11276 2604
rect 11340 2540 11356 2604
rect 11420 2540 11436 2604
rect 11500 2540 11642 2604
rect 11706 2540 11722 2604
rect 11786 2540 11802 2604
rect 11866 2540 11882 2604
rect 11946 2540 11962 2604
rect 12026 2540 12042 2604
rect 12106 2540 12248 2604
rect 12312 2540 12328 2604
rect 12392 2540 12408 2604
rect 12472 2540 12488 2604
rect 12552 2540 12568 2604
rect 12632 2540 12648 2604
rect 12712 2540 12854 2604
rect 12918 2540 12934 2604
rect 12998 2540 13014 2604
rect 13078 2540 13094 2604
rect 13158 2540 13174 2604
rect 13238 2540 13254 2604
rect 13318 2540 13460 2604
rect 13524 2540 13540 2604
rect 13604 2540 13620 2604
rect 13684 2540 13700 2604
rect 13764 2540 13780 2604
rect 13844 2540 13860 2604
rect 13924 2540 14066 2604
rect 14130 2540 14146 2604
rect 14210 2540 14226 2604
rect 14290 2540 14306 2604
rect 14370 2540 14386 2604
rect 14450 2540 14466 2604
rect 14530 2540 14672 2604
rect 14736 2540 14752 2604
rect 14816 2540 14832 2604
rect 14896 2540 14912 2604
rect 14976 2540 14992 2604
rect 15056 2540 15072 2604
rect 15136 2540 15278 2604
rect 15342 2540 15358 2604
rect 15422 2540 15438 2604
rect 15502 2540 15518 2604
rect 15582 2540 15598 2604
rect 15662 2540 15678 2604
rect 15742 2540 15884 2604
rect 15948 2540 15964 2604
rect 16028 2540 16044 2604
rect 16108 2540 16124 2604
rect 16188 2540 16204 2604
rect 16268 2540 16284 2604
rect 16348 2540 16490 2604
rect 16554 2540 16570 2604
rect 16634 2540 16650 2604
rect 16714 2540 16730 2604
rect 16794 2540 16810 2604
rect 16874 2540 16890 2604
rect 16954 2540 17096 2604
rect 17160 2540 17176 2604
rect 17240 2540 17256 2604
rect 17320 2540 17336 2604
rect 17400 2540 17416 2604
rect 17480 2540 17496 2604
rect 17560 2540 17702 2604
rect 17766 2540 17782 2604
rect 17846 2540 17862 2604
rect 17926 2540 17942 2604
rect 18006 2540 18022 2604
rect 18086 2540 18102 2604
rect 18166 2540 18308 2604
rect 18372 2540 18388 2604
rect 18452 2540 18468 2604
rect 18532 2540 18548 2604
rect 18612 2540 18628 2604
rect 18692 2540 18708 2604
rect 18772 2540 18914 2604
rect 18978 2540 18994 2604
rect 19058 2540 19074 2604
rect 19138 2540 19154 2604
rect 19218 2540 19234 2604
rect 19298 2540 19314 2604
rect 19378 2540 19520 2604
rect 19584 2540 19600 2604
rect 19664 2540 19680 2604
rect 19744 2540 19760 2604
rect 19824 2540 19840 2604
rect 19904 2540 19920 2604
rect 19984 2540 20088 2604
rect 10326 2538 20088 2540
rect 20148 2604 39606 2606
rect 20148 2540 20252 2604
rect 20316 2540 20332 2604
rect 20396 2540 20412 2604
rect 20476 2540 20492 2604
rect 20556 2540 20572 2604
rect 20636 2540 20652 2604
rect 20716 2540 20858 2604
rect 20922 2540 20938 2604
rect 21002 2540 21018 2604
rect 21082 2540 21098 2604
rect 21162 2540 21178 2604
rect 21242 2540 21258 2604
rect 21322 2540 21464 2604
rect 21528 2540 21544 2604
rect 21608 2540 21624 2604
rect 21688 2540 21704 2604
rect 21768 2540 21784 2604
rect 21848 2540 21864 2604
rect 21928 2540 22070 2604
rect 22134 2540 22150 2604
rect 22214 2540 22230 2604
rect 22294 2540 22310 2604
rect 22374 2540 22390 2604
rect 22454 2540 22470 2604
rect 22534 2540 22676 2604
rect 22740 2540 22756 2604
rect 22820 2540 22836 2604
rect 22900 2540 22916 2604
rect 22980 2540 22996 2604
rect 23060 2540 23076 2604
rect 23140 2540 23282 2604
rect 23346 2540 23362 2604
rect 23426 2540 23442 2604
rect 23506 2540 23522 2604
rect 23586 2540 23602 2604
rect 23666 2540 23682 2604
rect 23746 2540 23888 2604
rect 23952 2540 23968 2604
rect 24032 2540 24048 2604
rect 24112 2540 24128 2604
rect 24192 2540 24208 2604
rect 24272 2540 24288 2604
rect 24352 2540 24494 2604
rect 24558 2540 24574 2604
rect 24638 2540 24654 2604
rect 24718 2540 24734 2604
rect 24798 2540 24814 2604
rect 24878 2540 24894 2604
rect 24958 2540 25100 2604
rect 25164 2540 25180 2604
rect 25244 2540 25260 2604
rect 25324 2540 25340 2604
rect 25404 2540 25420 2604
rect 25484 2540 25500 2604
rect 25564 2540 25706 2604
rect 25770 2540 25786 2604
rect 25850 2540 25866 2604
rect 25930 2540 25946 2604
rect 26010 2540 26026 2604
rect 26090 2540 26106 2604
rect 26170 2540 26312 2604
rect 26376 2540 26392 2604
rect 26456 2540 26472 2604
rect 26536 2540 26552 2604
rect 26616 2540 26632 2604
rect 26696 2540 26712 2604
rect 26776 2540 26918 2604
rect 26982 2540 26998 2604
rect 27062 2540 27078 2604
rect 27142 2540 27158 2604
rect 27222 2540 27238 2604
rect 27302 2540 27318 2604
rect 27382 2540 27524 2604
rect 27588 2540 27604 2604
rect 27668 2540 27684 2604
rect 27748 2540 27764 2604
rect 27828 2540 27844 2604
rect 27908 2540 27924 2604
rect 27988 2540 28130 2604
rect 28194 2540 28210 2604
rect 28274 2540 28290 2604
rect 28354 2540 28370 2604
rect 28434 2540 28450 2604
rect 28514 2540 28530 2604
rect 28594 2540 28736 2604
rect 28800 2540 28816 2604
rect 28880 2540 28896 2604
rect 28960 2540 28976 2604
rect 29040 2540 29056 2604
rect 29120 2540 29136 2604
rect 29200 2540 29342 2604
rect 29406 2540 29422 2604
rect 29486 2540 29502 2604
rect 29566 2540 29582 2604
rect 29646 2540 29662 2604
rect 29726 2540 29742 2604
rect 29806 2540 29948 2604
rect 30012 2540 30028 2604
rect 30092 2540 30108 2604
rect 30172 2540 30188 2604
rect 30252 2540 30268 2604
rect 30332 2540 30348 2604
rect 30412 2540 30554 2604
rect 30618 2540 30634 2604
rect 30698 2540 30714 2604
rect 30778 2540 30794 2604
rect 30858 2540 30874 2604
rect 30938 2540 30954 2604
rect 31018 2540 31160 2604
rect 31224 2540 31240 2604
rect 31304 2540 31320 2604
rect 31384 2540 31400 2604
rect 31464 2540 31480 2604
rect 31544 2540 31560 2604
rect 31624 2540 31766 2604
rect 31830 2540 31846 2604
rect 31910 2540 31926 2604
rect 31990 2540 32006 2604
rect 32070 2540 32086 2604
rect 32150 2540 32166 2604
rect 32230 2540 32372 2604
rect 32436 2540 32452 2604
rect 32516 2540 32532 2604
rect 32596 2540 32612 2604
rect 32676 2540 32692 2604
rect 32756 2540 32772 2604
rect 32836 2540 32978 2604
rect 33042 2540 33058 2604
rect 33122 2540 33138 2604
rect 33202 2540 33218 2604
rect 33282 2540 33298 2604
rect 33362 2540 33378 2604
rect 33442 2540 33584 2604
rect 33648 2540 33664 2604
rect 33728 2540 33744 2604
rect 33808 2540 33824 2604
rect 33888 2540 33904 2604
rect 33968 2540 33984 2604
rect 34048 2540 34190 2604
rect 34254 2540 34270 2604
rect 34334 2540 34350 2604
rect 34414 2540 34430 2604
rect 34494 2540 34510 2604
rect 34574 2540 34590 2604
rect 34654 2540 34796 2604
rect 34860 2540 34876 2604
rect 34940 2540 34956 2604
rect 35020 2540 35036 2604
rect 35100 2540 35116 2604
rect 35180 2540 35196 2604
rect 35260 2540 35402 2604
rect 35466 2540 35482 2604
rect 35546 2540 35562 2604
rect 35626 2540 35642 2604
rect 35706 2540 35722 2604
rect 35786 2540 35802 2604
rect 35866 2540 36008 2604
rect 36072 2540 36088 2604
rect 36152 2540 36168 2604
rect 36232 2540 36248 2604
rect 36312 2540 36328 2604
rect 36392 2540 36408 2604
rect 36472 2540 36614 2604
rect 36678 2540 36694 2604
rect 36758 2540 36774 2604
rect 36838 2540 36854 2604
rect 36918 2540 36934 2604
rect 36998 2540 37014 2604
rect 37078 2540 37220 2604
rect 37284 2540 37300 2604
rect 37364 2540 37380 2604
rect 37444 2540 37460 2604
rect 37524 2540 37540 2604
rect 37604 2540 37620 2604
rect 37684 2540 37826 2604
rect 37890 2540 37906 2604
rect 37970 2540 37986 2604
rect 38050 2540 38066 2604
rect 38130 2540 38146 2604
rect 38210 2540 38226 2604
rect 38290 2540 38432 2604
rect 38496 2540 38512 2604
rect 38576 2540 38592 2604
rect 38656 2540 38672 2604
rect 38736 2540 38752 2604
rect 38816 2540 38832 2604
rect 38896 2540 39038 2604
rect 39102 2540 39118 2604
rect 39182 2540 39198 2604
rect 39262 2540 39278 2604
rect 39342 2540 39358 2604
rect 39422 2540 39438 2604
rect 39502 2540 39606 2604
rect 20148 2538 39606 2540
rect -459 2384 -393 2538
rect -459 2320 -458 2384
rect -394 2320 -393 2384
rect -459 2304 -393 2320
rect -459 2240 -458 2304
rect -394 2240 -393 2304
rect -459 2224 -393 2240
rect -459 2160 -458 2224
rect -394 2160 -393 2224
rect -459 2144 -393 2160
rect -459 2080 -458 2144
rect -394 2080 -393 2144
rect -459 2064 -393 2080
rect -459 2000 -458 2064
rect -394 2000 -393 2064
rect -459 1984 -393 2000
rect -459 1920 -458 1984
rect -394 1920 -393 1984
rect -459 1904 -393 1920
rect -459 1840 -458 1904
rect -394 1840 -393 1904
rect -459 1824 -393 1840
rect -459 1760 -458 1824
rect -394 1760 -393 1824
rect -459 1744 -393 1760
rect -459 1680 -458 1744
rect -394 1680 -393 1744
rect -459 1664 -393 1680
rect -459 1600 -458 1664
rect -394 1600 -393 1664
rect -459 1510 -393 1600
rect -333 1446 -273 2476
rect -213 1506 -153 2538
rect -93 1446 -33 2476
rect 27 1506 87 2538
rect 147 2384 213 2538
rect 147 2320 148 2384
rect 212 2320 213 2384
rect 147 2304 213 2320
rect 147 2240 148 2304
rect 212 2240 213 2304
rect 147 2224 213 2240
rect 147 2160 148 2224
rect 212 2160 213 2224
rect 147 2144 213 2160
rect 147 2080 148 2144
rect 212 2080 213 2144
rect 147 2064 213 2080
rect 147 2000 148 2064
rect 212 2000 213 2064
rect 147 1984 213 2000
rect 147 1920 148 1984
rect 212 1920 213 1984
rect 147 1904 213 1920
rect 147 1840 148 1904
rect 212 1840 213 1904
rect 147 1824 213 1840
rect 147 1760 148 1824
rect 212 1760 213 1824
rect 147 1744 213 1760
rect 147 1680 148 1744
rect 212 1680 213 1744
rect 147 1664 213 1680
rect 147 1600 148 1664
rect 212 1600 213 1664
rect 147 1510 213 1600
rect 355 2384 421 2474
rect 355 2320 356 2384
rect 420 2320 421 2384
rect 355 2304 421 2320
rect 355 2240 356 2304
rect 420 2240 421 2304
rect 355 2224 421 2240
rect 355 2160 356 2224
rect 420 2160 421 2224
rect 355 2144 421 2160
rect 355 2080 356 2144
rect 420 2080 421 2144
rect 355 2064 421 2080
rect 355 2000 356 2064
rect 420 2000 421 2064
rect 355 1984 421 2000
rect 355 1920 356 1984
rect 420 1920 421 1984
rect 355 1904 421 1920
rect 355 1840 356 1904
rect 420 1840 421 1904
rect 355 1824 421 1840
rect 355 1760 356 1824
rect 420 1760 421 1824
rect 355 1744 421 1760
rect 355 1680 356 1744
rect 420 1680 421 1744
rect 355 1664 421 1680
rect 355 1600 356 1664
rect 420 1600 421 1664
rect 355 1446 421 1600
rect 481 1446 541 2478
rect 601 1508 661 2538
rect 721 1446 781 2478
rect 841 1508 901 2538
rect 964 2474 1024 2476
rect 961 2465 1027 2474
rect 961 2401 962 2465
rect 1026 2401 1027 2465
rect 961 2384 1027 2401
rect 961 2320 962 2384
rect 1026 2320 1027 2384
rect 961 2304 1027 2320
rect 961 2240 962 2304
rect 1026 2240 1027 2304
rect 961 2224 1027 2240
rect 961 2160 962 2224
rect 1026 2160 1027 2224
rect 961 2144 1027 2160
rect 961 2080 962 2144
rect 1026 2080 1027 2144
rect 961 2064 1027 2080
rect 961 2000 962 2064
rect 1026 2000 1027 2064
rect 961 1984 1027 2000
rect 961 1920 962 1984
rect 1026 1920 1027 1984
rect 961 1904 1027 1920
rect 961 1840 962 1904
rect 1026 1840 1027 1904
rect 961 1824 1027 1840
rect 961 1760 962 1824
rect 1026 1760 1027 1824
rect 961 1744 1027 1760
rect 961 1680 962 1744
rect 1026 1680 1027 1744
rect 961 1664 1027 1680
rect 961 1600 962 1664
rect 1026 1600 1027 1664
rect 961 1446 1027 1600
rect -459 1444 213 1446
rect -459 1380 -355 1444
rect -291 1380 -275 1444
rect -211 1380 -195 1444
rect -131 1380 -115 1444
rect -51 1380 -35 1444
rect 29 1380 45 1444
rect 109 1380 213 1444
rect -459 1378 213 1380
rect 355 1444 1027 1446
rect 355 1380 459 1444
rect 523 1380 539 1444
rect 603 1380 619 1444
rect 683 1380 699 1444
rect 763 1380 779 1444
rect 843 1380 859 1444
rect 923 1380 1027 1444
rect 355 1378 1027 1380
rect -459 1224 -393 1314
rect -459 1160 -458 1224
rect -394 1160 -393 1224
rect -459 1144 -393 1160
rect -459 1080 -458 1144
rect -394 1080 -393 1144
rect -459 1064 -393 1080
rect -459 1000 -458 1064
rect -394 1000 -393 1064
rect -459 984 -393 1000
rect -459 920 -458 984
rect -394 920 -393 984
rect -459 904 -393 920
rect -459 840 -458 904
rect -394 840 -393 904
rect -459 824 -393 840
rect -459 760 -458 824
rect -394 760 -393 824
rect -459 744 -393 760
rect -459 680 -458 744
rect -394 680 -393 744
rect -459 664 -393 680
rect -459 600 -458 664
rect -394 600 -393 664
rect -459 584 -393 600
rect -459 520 -458 584
rect -394 520 -393 584
rect -459 504 -393 520
rect -459 440 -458 504
rect -394 440 -393 504
rect -459 286 -393 440
rect -333 286 -273 1318
rect -213 348 -153 1378
rect -93 286 -33 1318
rect 27 348 87 1378
rect 147 1224 213 1314
rect 147 1160 148 1224
rect 212 1160 213 1224
rect 147 1144 213 1160
rect 147 1080 148 1144
rect 212 1080 213 1144
rect 147 1064 213 1080
rect 147 1000 148 1064
rect 212 1000 213 1064
rect 147 984 213 1000
rect 147 920 148 984
rect 212 920 213 984
rect 147 904 213 920
rect 147 840 148 904
rect 212 840 213 904
rect 147 824 213 840
rect 147 760 148 824
rect 212 760 213 824
rect 147 744 213 760
rect 147 680 148 744
rect 212 680 213 744
rect 147 664 213 680
rect 147 600 148 664
rect 212 600 213 664
rect 147 584 213 600
rect 147 520 148 584
rect 212 520 213 584
rect 147 504 213 520
rect 147 440 148 504
rect 212 440 213 504
rect 147 286 213 440
rect 355 1224 421 1378
rect 355 1160 356 1224
rect 420 1160 421 1224
rect 355 1144 421 1160
rect 355 1080 356 1144
rect 420 1080 421 1144
rect 355 1064 421 1080
rect 355 1000 356 1064
rect 420 1000 421 1064
rect 355 984 421 1000
rect 355 920 356 984
rect 420 920 421 984
rect 355 904 421 920
rect 355 840 356 904
rect 420 840 421 904
rect 355 824 421 840
rect 355 760 356 824
rect 420 760 421 824
rect 355 744 421 760
rect 355 680 356 744
rect 420 680 421 744
rect 355 664 421 680
rect 355 600 356 664
rect 420 600 421 664
rect 355 584 421 600
rect 355 520 356 584
rect 420 520 421 584
rect 355 504 421 520
rect 355 440 356 504
rect 420 440 421 504
rect 355 350 421 440
rect 481 286 541 1316
rect 601 346 661 1378
rect 721 286 781 1316
rect 841 346 901 1378
rect 961 1224 1027 1378
rect 961 1160 962 1224
rect 1026 1160 1027 1224
rect 961 1144 1027 1160
rect 961 1080 962 1144
rect 1026 1080 1027 1144
rect 961 1064 1027 1080
rect 961 1000 962 1064
rect 1026 1000 1027 1064
rect 961 984 1027 1000
rect 961 920 962 984
rect 1026 920 1027 984
rect 961 904 1027 920
rect 961 840 962 904
rect 1026 840 1027 904
rect 961 824 1027 840
rect 961 760 962 824
rect 1026 760 1027 824
rect 961 744 1027 760
rect 961 680 962 744
rect 1026 680 1027 744
rect 961 664 1027 680
rect 961 600 962 664
rect 1026 600 1027 664
rect 961 584 1027 600
rect 961 520 962 584
rect 1026 520 1027 584
rect 961 504 1027 520
rect 961 440 962 504
rect 1026 440 1027 504
rect 961 350 1027 440
rect 1267 2384 1333 2474
rect 1267 2320 1268 2384
rect 1332 2320 1333 2384
rect 1267 2304 1333 2320
rect 1267 2240 1268 2304
rect 1332 2240 1333 2304
rect 1267 2224 1333 2240
rect 1267 2160 1268 2224
rect 1332 2160 1333 2224
rect 1267 2144 1333 2160
rect 1267 2080 1268 2144
rect 1332 2080 1333 2144
rect 1267 2064 1333 2080
rect 1267 2000 1268 2064
rect 1332 2000 1333 2064
rect 1267 1984 1333 2000
rect 1267 1920 1268 1984
rect 1332 1920 1333 1984
rect 1267 1904 1333 1920
rect 1267 1840 1268 1904
rect 1332 1840 1333 1904
rect 1267 1824 1333 1840
rect 1267 1760 1268 1824
rect 1332 1760 1333 1824
rect 1267 1744 1333 1760
rect 1267 1680 1268 1744
rect 1332 1680 1333 1744
rect 1267 1664 1333 1680
rect 1267 1600 1268 1664
rect 1332 1600 1333 1664
rect 1267 1446 1333 1600
rect 1393 1446 1453 2478
rect 1513 1508 1573 2538
rect 1633 1446 1693 2478
rect 1753 1508 1813 2538
rect 1873 2384 1939 2474
rect 1873 2320 1874 2384
rect 1938 2320 1939 2384
rect 1873 2304 1939 2320
rect 1873 2240 1874 2304
rect 1938 2240 1939 2304
rect 1873 2224 1939 2240
rect 1873 2160 1874 2224
rect 1938 2160 1939 2224
rect 1873 2144 1939 2160
rect 1873 2080 1874 2144
rect 1938 2080 1939 2144
rect 1873 2064 1939 2080
rect 1873 2000 1874 2064
rect 1938 2000 1939 2064
rect 1873 1984 1939 2000
rect 1873 1920 1874 1984
rect 1938 1920 1939 1984
rect 1873 1904 1939 1920
rect 1873 1840 1874 1904
rect 1938 1840 1939 1904
rect 1873 1824 1939 1840
rect 1873 1760 1874 1824
rect 1938 1760 1939 1824
rect 1873 1744 1939 1760
rect 1873 1680 1874 1744
rect 1938 1680 1939 1744
rect 1873 1664 1939 1680
rect 1873 1600 1874 1664
rect 1938 1600 1939 1664
rect 1873 1446 1939 1600
rect 1999 1446 2059 2478
rect 2119 1508 2179 2538
rect 2239 1446 2299 2478
rect 2359 1508 2419 2538
rect 2482 2474 2542 2476
rect 2479 2465 2545 2474
rect 2479 2401 2480 2465
rect 2544 2401 2545 2465
rect 2479 2384 2545 2401
rect 2479 2320 2480 2384
rect 2544 2320 2545 2384
rect 2479 2304 2545 2320
rect 2479 2240 2480 2304
rect 2544 2240 2545 2304
rect 2479 2224 2545 2240
rect 2479 2160 2480 2224
rect 2544 2160 2545 2224
rect 2479 2144 2545 2160
rect 2479 2080 2480 2144
rect 2544 2080 2545 2144
rect 2479 2064 2545 2080
rect 2479 2000 2480 2064
rect 2544 2000 2545 2064
rect 2479 1984 2545 2000
rect 2479 1920 2480 1984
rect 2544 1920 2545 1984
rect 2479 1904 2545 1920
rect 2479 1840 2480 1904
rect 2544 1840 2545 1904
rect 2479 1824 2545 1840
rect 2479 1760 2480 1824
rect 2544 1760 2545 1824
rect 2479 1744 2545 1760
rect 2479 1680 2480 1744
rect 2544 1680 2545 1744
rect 2479 1664 2545 1680
rect 2479 1600 2480 1664
rect 2544 1600 2545 1664
rect 2479 1446 2545 1600
rect 1267 1444 2545 1446
rect 1267 1380 1371 1444
rect 1435 1380 1451 1444
rect 1515 1380 1531 1444
rect 1595 1380 1611 1444
rect 1675 1380 1691 1444
rect 1755 1380 1771 1444
rect 1835 1380 1977 1444
rect 2041 1380 2057 1444
rect 2121 1380 2137 1444
rect 2201 1380 2217 1444
rect 2281 1380 2297 1444
rect 2361 1380 2377 1444
rect 2441 1380 2545 1444
rect 1267 1378 2545 1380
rect 1267 1224 1333 1378
rect 1267 1160 1268 1224
rect 1332 1160 1333 1224
rect 1267 1144 1333 1160
rect 1267 1080 1268 1144
rect 1332 1080 1333 1144
rect 1267 1064 1333 1080
rect 1267 1000 1268 1064
rect 1332 1000 1333 1064
rect 1267 984 1333 1000
rect 1267 920 1268 984
rect 1332 920 1333 984
rect 1267 904 1333 920
rect 1267 840 1268 904
rect 1332 840 1333 904
rect 1267 824 1333 840
rect 1267 760 1268 824
rect 1332 760 1333 824
rect 1267 744 1333 760
rect 1267 680 1268 744
rect 1332 680 1333 744
rect 1267 664 1333 680
rect 1267 600 1268 664
rect 1332 600 1333 664
rect 1267 584 1333 600
rect 1267 520 1268 584
rect 1332 520 1333 584
rect 1267 504 1333 520
rect 1267 440 1268 504
rect 1332 440 1333 504
rect 1267 350 1333 440
rect 1393 286 1453 1316
rect 1513 346 1573 1378
rect 1633 286 1693 1316
rect 1753 346 1813 1378
rect 1873 1224 1939 1378
rect 1873 1160 1874 1224
rect 1938 1160 1939 1224
rect 1873 1144 1939 1160
rect 1873 1080 1874 1144
rect 1938 1080 1939 1144
rect 1873 1064 1939 1080
rect 1873 1000 1874 1064
rect 1938 1000 1939 1064
rect 1873 984 1939 1000
rect 1873 920 1874 984
rect 1938 920 1939 984
rect 1873 904 1939 920
rect 1873 840 1874 904
rect 1938 840 1939 904
rect 1873 824 1939 840
rect 1873 760 1874 824
rect 1938 760 1939 824
rect 1873 744 1939 760
rect 1873 680 1874 744
rect 1938 680 1939 744
rect 1873 664 1939 680
rect 1873 600 1874 664
rect 1938 600 1939 664
rect 1873 584 1939 600
rect 1873 520 1874 584
rect 1938 520 1939 584
rect 1873 504 1939 520
rect 1873 440 1874 504
rect 1938 440 1939 504
rect 1873 350 1939 440
rect 1999 286 2059 1316
rect 2119 346 2179 1378
rect 2239 286 2299 1316
rect 2359 346 2419 1378
rect 2479 1224 2545 1378
rect 2479 1160 2480 1224
rect 2544 1160 2545 1224
rect 2479 1144 2545 1160
rect 2479 1080 2480 1144
rect 2544 1080 2545 1144
rect 2479 1064 2545 1080
rect 2479 1000 2480 1064
rect 2544 1000 2545 1064
rect 2479 984 2545 1000
rect 2479 920 2480 984
rect 2544 920 2545 984
rect 2479 904 2545 920
rect 2479 840 2480 904
rect 2544 840 2545 904
rect 2479 824 2545 840
rect 2479 760 2480 824
rect 2544 760 2545 824
rect 2479 744 2545 760
rect 2479 680 2480 744
rect 2544 680 2545 744
rect 2479 664 2545 680
rect 2479 600 2480 664
rect 2544 600 2545 664
rect 2479 584 2545 600
rect 2479 520 2480 584
rect 2544 520 2545 584
rect 2479 504 2545 520
rect 2479 440 2480 504
rect 2544 440 2545 504
rect 2479 350 2545 440
rect 2801 2384 2867 2474
rect 2801 2320 2802 2384
rect 2866 2320 2867 2384
rect 2801 2304 2867 2320
rect 2801 2240 2802 2304
rect 2866 2240 2867 2304
rect 2801 2224 2867 2240
rect 2801 2160 2802 2224
rect 2866 2160 2867 2224
rect 2801 2144 2867 2160
rect 2801 2080 2802 2144
rect 2866 2080 2867 2144
rect 2801 2064 2867 2080
rect 2801 2000 2802 2064
rect 2866 2000 2867 2064
rect 2801 1984 2867 2000
rect 2801 1920 2802 1984
rect 2866 1920 2867 1984
rect 2801 1904 2867 1920
rect 2801 1840 2802 1904
rect 2866 1840 2867 1904
rect 2801 1824 2867 1840
rect 2801 1760 2802 1824
rect 2866 1760 2867 1824
rect 2801 1744 2867 1760
rect 2801 1680 2802 1744
rect 2866 1680 2867 1744
rect 2801 1664 2867 1680
rect 2801 1600 2802 1664
rect 2866 1600 2867 1664
rect 2801 1446 2867 1600
rect 2927 1446 2987 2478
rect 3047 1508 3107 2538
rect 3167 1446 3227 2478
rect 3287 1508 3347 2538
rect 3407 2384 3473 2474
rect 3407 2320 3408 2384
rect 3472 2320 3473 2384
rect 3407 2304 3473 2320
rect 3407 2240 3408 2304
rect 3472 2240 3473 2304
rect 3407 2224 3473 2240
rect 3407 2160 3408 2224
rect 3472 2160 3473 2224
rect 3407 2144 3473 2160
rect 3407 2080 3408 2144
rect 3472 2080 3473 2144
rect 3407 2064 3473 2080
rect 3407 2000 3408 2064
rect 3472 2000 3473 2064
rect 3407 1984 3473 2000
rect 3407 1920 3408 1984
rect 3472 1920 3473 1984
rect 3407 1904 3473 1920
rect 3407 1840 3408 1904
rect 3472 1840 3473 1904
rect 3407 1824 3473 1840
rect 3407 1760 3408 1824
rect 3472 1760 3473 1824
rect 3407 1744 3473 1760
rect 3407 1680 3408 1744
rect 3472 1680 3473 1744
rect 3407 1664 3473 1680
rect 3407 1600 3408 1664
rect 3472 1600 3473 1664
rect 3407 1446 3473 1600
rect 3533 1446 3593 2478
rect 3653 1508 3713 2538
rect 3773 1446 3833 2478
rect 3893 1508 3953 2538
rect 4013 2384 4079 2474
rect 4013 2320 4014 2384
rect 4078 2320 4079 2384
rect 4013 2304 4079 2320
rect 4013 2240 4014 2304
rect 4078 2240 4079 2304
rect 4013 2224 4079 2240
rect 4013 2160 4014 2224
rect 4078 2160 4079 2224
rect 4013 2144 4079 2160
rect 4013 2080 4014 2144
rect 4078 2080 4079 2144
rect 4013 2064 4079 2080
rect 4013 2000 4014 2064
rect 4078 2000 4079 2064
rect 4013 1984 4079 2000
rect 4013 1920 4014 1984
rect 4078 1920 4079 1984
rect 4013 1904 4079 1920
rect 4013 1840 4014 1904
rect 4078 1840 4079 1904
rect 4013 1824 4079 1840
rect 4013 1760 4014 1824
rect 4078 1760 4079 1824
rect 4013 1744 4079 1760
rect 4013 1680 4014 1744
rect 4078 1680 4079 1744
rect 4013 1664 4079 1680
rect 4013 1600 4014 1664
rect 4078 1600 4079 1664
rect 4013 1446 4079 1600
rect 4139 1446 4199 2478
rect 4259 1508 4319 2538
rect 4379 1446 4439 2478
rect 4499 1508 4559 2538
rect 4619 2451 4685 2474
rect 4619 2395 4624 2451
rect 4680 2395 4685 2451
rect 4619 2384 4685 2395
rect 4619 2320 4620 2384
rect 4684 2320 4685 2384
rect 4619 2304 4685 2320
rect 4619 2240 4620 2304
rect 4684 2240 4685 2304
rect 4619 2224 4685 2240
rect 4619 2160 4620 2224
rect 4684 2160 4685 2224
rect 4619 2144 4685 2160
rect 4619 2080 4620 2144
rect 4684 2080 4685 2144
rect 4619 2064 4685 2080
rect 4619 2000 4620 2064
rect 4684 2000 4685 2064
rect 4619 1984 4685 2000
rect 4619 1920 4620 1984
rect 4684 1920 4685 1984
rect 4619 1904 4685 1920
rect 4619 1840 4620 1904
rect 4684 1840 4685 1904
rect 4619 1824 4685 1840
rect 4619 1760 4620 1824
rect 4684 1760 4685 1824
rect 4619 1744 4685 1760
rect 4619 1680 4620 1744
rect 4684 1680 4685 1744
rect 4619 1664 4685 1680
rect 4619 1600 4620 1664
rect 4684 1600 4685 1664
rect 4619 1446 4685 1600
rect 4745 1446 4805 2478
rect 4865 1508 4925 2538
rect 4985 1446 5045 2478
rect 5105 1508 5165 2538
rect 5225 2384 5291 2474
rect 5225 2320 5226 2384
rect 5290 2320 5291 2384
rect 5225 2304 5291 2320
rect 5225 2240 5226 2304
rect 5290 2240 5291 2304
rect 5225 2224 5291 2240
rect 5225 2160 5226 2224
rect 5290 2160 5291 2224
rect 5225 2144 5291 2160
rect 5225 2080 5226 2144
rect 5290 2080 5291 2144
rect 5225 2064 5291 2080
rect 5225 2000 5226 2064
rect 5290 2000 5291 2064
rect 5225 1984 5291 2000
rect 5225 1920 5226 1984
rect 5290 1920 5291 1984
rect 5225 1904 5291 1920
rect 5225 1840 5226 1904
rect 5290 1840 5291 1904
rect 5225 1824 5291 1840
rect 5225 1760 5226 1824
rect 5290 1760 5291 1824
rect 5225 1744 5291 1760
rect 5225 1680 5226 1744
rect 5290 1680 5291 1744
rect 5225 1664 5291 1680
rect 5225 1600 5226 1664
rect 5290 1600 5291 1664
rect 5225 1446 5291 1600
rect 2801 1444 5291 1446
rect 2801 1380 2905 1444
rect 2969 1380 2985 1444
rect 3049 1380 3065 1444
rect 3129 1380 3145 1444
rect 3209 1380 3225 1444
rect 3289 1380 3305 1444
rect 3369 1380 3511 1444
rect 3575 1380 3591 1444
rect 3655 1380 3671 1444
rect 3735 1380 3751 1444
rect 3815 1380 3831 1444
rect 3895 1380 3911 1444
rect 3975 1380 4117 1444
rect 4181 1380 4197 1444
rect 4261 1380 4277 1444
rect 4341 1380 4357 1444
rect 4421 1380 4437 1444
rect 4501 1380 4517 1444
rect 4581 1380 4723 1444
rect 4787 1380 4803 1444
rect 4867 1380 4883 1444
rect 4947 1380 4963 1444
rect 5027 1380 5043 1444
rect 5107 1380 5123 1444
rect 5187 1380 5291 1444
rect 2801 1378 5291 1380
rect 2801 1224 2867 1378
rect 2801 1160 2802 1224
rect 2866 1160 2867 1224
rect 2801 1144 2867 1160
rect 2801 1080 2802 1144
rect 2866 1080 2867 1144
rect 2801 1064 2867 1080
rect 2801 1000 2802 1064
rect 2866 1000 2867 1064
rect 2801 984 2867 1000
rect 2801 920 2802 984
rect 2866 920 2867 984
rect 2801 904 2867 920
rect 2801 840 2802 904
rect 2866 840 2867 904
rect 2801 824 2867 840
rect 2801 760 2802 824
rect 2866 760 2867 824
rect 2801 744 2867 760
rect 2801 680 2802 744
rect 2866 680 2867 744
rect 2801 664 2867 680
rect 2801 600 2802 664
rect 2866 600 2867 664
rect 2801 584 2867 600
rect 2801 520 2802 584
rect 2866 520 2867 584
rect 2801 504 2867 520
rect 2801 440 2802 504
rect 2866 440 2867 504
rect 2801 350 2867 440
rect 2927 286 2987 1316
rect 3047 346 3107 1378
rect 3167 286 3227 1316
rect 3287 346 3347 1378
rect 3407 1224 3473 1378
rect 3407 1160 3408 1224
rect 3472 1160 3473 1224
rect 3407 1144 3473 1160
rect 3407 1080 3408 1144
rect 3472 1080 3473 1144
rect 3407 1064 3473 1080
rect 3407 1000 3408 1064
rect 3472 1000 3473 1064
rect 3407 984 3473 1000
rect 3407 920 3408 984
rect 3472 920 3473 984
rect 3407 904 3473 920
rect 3407 840 3408 904
rect 3472 840 3473 904
rect 3407 824 3473 840
rect 3407 760 3408 824
rect 3472 760 3473 824
rect 3407 744 3473 760
rect 3407 680 3408 744
rect 3472 680 3473 744
rect 3407 664 3473 680
rect 3407 600 3408 664
rect 3472 600 3473 664
rect 3407 584 3473 600
rect 3407 520 3408 584
rect 3472 520 3473 584
rect 3407 504 3473 520
rect 3407 440 3408 504
rect 3472 440 3473 504
rect 3407 350 3473 440
rect 3533 286 3593 1316
rect 3653 346 3713 1378
rect 3773 286 3833 1316
rect 3893 346 3953 1378
rect 4013 1224 4079 1378
rect 4013 1160 4014 1224
rect 4078 1160 4079 1224
rect 4013 1144 4079 1160
rect 4013 1080 4014 1144
rect 4078 1080 4079 1144
rect 4013 1064 4079 1080
rect 4013 1000 4014 1064
rect 4078 1000 4079 1064
rect 4013 984 4079 1000
rect 4013 920 4014 984
rect 4078 920 4079 984
rect 4013 904 4079 920
rect 4013 840 4014 904
rect 4078 840 4079 904
rect 4013 824 4079 840
rect 4013 760 4014 824
rect 4078 760 4079 824
rect 4013 744 4079 760
rect 4013 680 4014 744
rect 4078 680 4079 744
rect 4013 664 4079 680
rect 4013 600 4014 664
rect 4078 600 4079 664
rect 4013 584 4079 600
rect 4013 520 4014 584
rect 4078 520 4079 584
rect 4013 504 4079 520
rect 4013 440 4014 504
rect 4078 440 4079 504
rect 4013 350 4079 440
rect 4139 286 4199 1316
rect 4259 346 4319 1378
rect 4379 286 4439 1316
rect 4499 346 4559 1378
rect 4619 1224 4685 1378
rect 4619 1160 4620 1224
rect 4684 1160 4685 1224
rect 4619 1144 4685 1160
rect 4619 1080 4620 1144
rect 4684 1080 4685 1144
rect 4619 1064 4685 1080
rect 4619 1000 4620 1064
rect 4684 1000 4685 1064
rect 4619 984 4685 1000
rect 4619 920 4620 984
rect 4684 920 4685 984
rect 4619 904 4685 920
rect 4619 840 4620 904
rect 4684 840 4685 904
rect 4619 824 4685 840
rect 4619 760 4620 824
rect 4684 760 4685 824
rect 4619 744 4685 760
rect 4619 680 4620 744
rect 4684 680 4685 744
rect 4619 664 4685 680
rect 4619 600 4620 664
rect 4684 600 4685 664
rect 4619 584 4685 600
rect 4619 520 4620 584
rect 4684 520 4685 584
rect 4619 504 4685 520
rect 4619 440 4620 504
rect 4684 440 4685 504
rect 4619 350 4685 440
rect 4745 286 4805 1316
rect 4865 346 4925 1378
rect 4985 286 5045 1316
rect 5105 346 5165 1378
rect 5225 1224 5291 1378
rect 5225 1160 5226 1224
rect 5290 1160 5291 1224
rect 5225 1144 5291 1160
rect 5225 1080 5226 1144
rect 5290 1080 5291 1144
rect 5225 1064 5291 1080
rect 5225 1000 5226 1064
rect 5290 1000 5291 1064
rect 5225 984 5291 1000
rect 5225 920 5226 984
rect 5290 920 5291 984
rect 5225 904 5291 920
rect 5225 840 5226 904
rect 5290 840 5291 904
rect 5225 824 5291 840
rect 5225 760 5226 824
rect 5290 760 5291 824
rect 5225 744 5291 760
rect 5225 680 5226 744
rect 5290 680 5291 744
rect 5225 664 5291 680
rect 5225 600 5226 664
rect 5290 600 5291 664
rect 5225 584 5291 600
rect 5225 520 5226 584
rect 5290 520 5291 584
rect 5225 504 5291 520
rect 5225 440 5226 504
rect 5290 440 5291 504
rect 5225 350 5291 440
rect 5352 2384 5418 2474
rect 5352 2320 5353 2384
rect 5417 2320 5418 2384
rect 5352 2304 5418 2320
rect 5352 2240 5353 2304
rect 5417 2240 5418 2304
rect 5352 2224 5418 2240
rect 5352 2160 5353 2224
rect 5417 2160 5418 2224
rect 5352 2144 5418 2160
rect 5352 2080 5353 2144
rect 5417 2080 5418 2144
rect 5352 2064 5418 2080
rect 5352 2000 5353 2064
rect 5417 2000 5418 2064
rect 5352 1984 5418 2000
rect 5352 1920 5353 1984
rect 5417 1920 5418 1984
rect 5352 1904 5418 1920
rect 5352 1840 5353 1904
rect 5417 1840 5418 1904
rect 5352 1824 5418 1840
rect 5352 1760 5353 1824
rect 5417 1760 5418 1824
rect 5352 1744 5418 1760
rect 5352 1680 5353 1744
rect 5417 1680 5418 1744
rect 5352 1664 5418 1680
rect 5352 1600 5353 1664
rect 5417 1600 5418 1664
rect 5352 1446 5418 1600
rect 5478 1446 5538 2478
rect 5598 1508 5658 2538
rect 5718 1446 5778 2478
rect 5838 1508 5898 2538
rect 5958 2384 6024 2474
rect 5958 2320 5959 2384
rect 6023 2320 6024 2384
rect 5958 2304 6024 2320
rect 5958 2240 5959 2304
rect 6023 2240 6024 2304
rect 5958 2224 6024 2240
rect 5958 2160 5959 2224
rect 6023 2160 6024 2224
rect 5958 2144 6024 2160
rect 5958 2080 5959 2144
rect 6023 2080 6024 2144
rect 5958 2064 6024 2080
rect 5958 2000 5959 2064
rect 6023 2000 6024 2064
rect 5958 1984 6024 2000
rect 5958 1920 5959 1984
rect 6023 1920 6024 1984
rect 5958 1904 6024 1920
rect 5958 1840 5959 1904
rect 6023 1840 6024 1904
rect 5958 1824 6024 1840
rect 5958 1760 5959 1824
rect 6023 1760 6024 1824
rect 5958 1744 6024 1760
rect 5958 1680 5959 1744
rect 6023 1680 6024 1744
rect 5958 1664 6024 1680
rect 5958 1600 5959 1664
rect 6023 1600 6024 1664
rect 5958 1446 6024 1600
rect 6084 1446 6144 2478
rect 6204 1508 6264 2538
rect 6324 1446 6384 2478
rect 6444 1508 6504 2538
rect 6564 2384 6630 2474
rect 6564 2320 6565 2384
rect 6629 2320 6630 2384
rect 6564 2304 6630 2320
rect 6564 2240 6565 2304
rect 6629 2240 6630 2304
rect 6564 2224 6630 2240
rect 6564 2160 6565 2224
rect 6629 2160 6630 2224
rect 6564 2144 6630 2160
rect 6564 2080 6565 2144
rect 6629 2080 6630 2144
rect 6564 2064 6630 2080
rect 6564 2000 6565 2064
rect 6629 2000 6630 2064
rect 6564 1984 6630 2000
rect 6564 1920 6565 1984
rect 6629 1920 6630 1984
rect 6564 1904 6630 1920
rect 6564 1840 6565 1904
rect 6629 1840 6630 1904
rect 6564 1824 6630 1840
rect 6564 1760 6565 1824
rect 6629 1760 6630 1824
rect 6564 1744 6630 1760
rect 6564 1680 6565 1744
rect 6629 1680 6630 1744
rect 6564 1664 6630 1680
rect 6564 1600 6565 1664
rect 6629 1600 6630 1664
rect 6564 1446 6630 1600
rect 6690 1446 6750 2478
rect 6810 1508 6870 2538
rect 6930 1446 6990 2478
rect 7050 1508 7110 2538
rect 7170 2384 7236 2474
rect 7170 2320 7171 2384
rect 7235 2320 7236 2384
rect 7170 2304 7236 2320
rect 7170 2240 7171 2304
rect 7235 2240 7236 2304
rect 7170 2224 7236 2240
rect 7170 2160 7171 2224
rect 7235 2160 7236 2224
rect 7170 2144 7236 2160
rect 7170 2080 7171 2144
rect 7235 2080 7236 2144
rect 7170 2064 7236 2080
rect 7170 2000 7171 2064
rect 7235 2000 7236 2064
rect 7170 1984 7236 2000
rect 7170 1920 7171 1984
rect 7235 1920 7236 1984
rect 7170 1904 7236 1920
rect 7170 1840 7171 1904
rect 7235 1840 7236 1904
rect 7170 1824 7236 1840
rect 7170 1760 7171 1824
rect 7235 1760 7236 1824
rect 7170 1744 7236 1760
rect 7170 1680 7171 1744
rect 7235 1680 7236 1744
rect 7170 1664 7236 1680
rect 7170 1600 7171 1664
rect 7235 1600 7236 1664
rect 7170 1446 7236 1600
rect 7296 1446 7356 2478
rect 7416 1508 7476 2538
rect 7536 1446 7596 2478
rect 7656 1508 7716 2538
rect 7776 2384 7842 2474
rect 7776 2320 7777 2384
rect 7841 2320 7842 2384
rect 7776 2304 7842 2320
rect 7776 2240 7777 2304
rect 7841 2240 7842 2304
rect 7776 2224 7842 2240
rect 7776 2160 7777 2224
rect 7841 2160 7842 2224
rect 7776 2144 7842 2160
rect 7776 2080 7777 2144
rect 7841 2080 7842 2144
rect 7776 2064 7842 2080
rect 7776 2000 7777 2064
rect 7841 2000 7842 2064
rect 7776 1984 7842 2000
rect 7776 1920 7777 1984
rect 7841 1920 7842 1984
rect 7776 1904 7842 1920
rect 7776 1840 7777 1904
rect 7841 1840 7842 1904
rect 7776 1824 7842 1840
rect 7776 1760 7777 1824
rect 7841 1760 7842 1824
rect 7776 1744 7842 1760
rect 7776 1680 7777 1744
rect 7841 1680 7842 1744
rect 7776 1664 7842 1680
rect 7776 1600 7777 1664
rect 7841 1600 7842 1664
rect 7776 1446 7842 1600
rect 7902 1446 7962 2478
rect 8022 1508 8082 2538
rect 8142 1446 8202 2478
rect 8262 1508 8322 2538
rect 8382 2384 8448 2474
rect 8382 2320 8383 2384
rect 8447 2320 8448 2384
rect 8382 2304 8448 2320
rect 8382 2240 8383 2304
rect 8447 2240 8448 2304
rect 8382 2224 8448 2240
rect 8382 2160 8383 2224
rect 8447 2160 8448 2224
rect 8382 2144 8448 2160
rect 8382 2080 8383 2144
rect 8447 2080 8448 2144
rect 8382 2064 8448 2080
rect 8382 2000 8383 2064
rect 8447 2000 8448 2064
rect 8382 1984 8448 2000
rect 8382 1920 8383 1984
rect 8447 1920 8448 1984
rect 8382 1904 8448 1920
rect 8382 1840 8383 1904
rect 8447 1840 8448 1904
rect 8382 1824 8448 1840
rect 8382 1760 8383 1824
rect 8447 1760 8448 1824
rect 8382 1744 8448 1760
rect 8382 1680 8383 1744
rect 8447 1680 8448 1744
rect 8382 1664 8448 1680
rect 8382 1600 8383 1664
rect 8447 1600 8448 1664
rect 8382 1446 8448 1600
rect 8508 1446 8568 2478
rect 8628 1508 8688 2538
rect 8748 1446 8808 2478
rect 8868 1508 8928 2538
rect 8988 2384 9054 2474
rect 8988 2320 8989 2384
rect 9053 2320 9054 2384
rect 8988 2304 9054 2320
rect 8988 2240 8989 2304
rect 9053 2240 9054 2304
rect 8988 2224 9054 2240
rect 8988 2160 8989 2224
rect 9053 2160 9054 2224
rect 8988 2144 9054 2160
rect 8988 2080 8989 2144
rect 9053 2080 9054 2144
rect 8988 2064 9054 2080
rect 8988 2000 8989 2064
rect 9053 2000 9054 2064
rect 8988 1984 9054 2000
rect 8988 1920 8989 1984
rect 9053 1920 9054 1984
rect 8988 1904 9054 1920
rect 8988 1840 8989 1904
rect 9053 1840 9054 1904
rect 8988 1824 9054 1840
rect 8988 1760 8989 1824
rect 9053 1760 9054 1824
rect 8988 1744 9054 1760
rect 8988 1680 8989 1744
rect 9053 1680 9054 1744
rect 8988 1664 9054 1680
rect 8988 1600 8989 1664
rect 9053 1600 9054 1664
rect 8988 1446 9054 1600
rect 9114 1446 9174 2478
rect 9234 1508 9294 2538
rect 9354 1446 9414 2478
rect 9474 1508 9534 2538
rect 9594 2384 9660 2474
rect 9594 2320 9595 2384
rect 9659 2320 9660 2384
rect 9594 2304 9660 2320
rect 9594 2240 9595 2304
rect 9659 2240 9660 2304
rect 9594 2224 9660 2240
rect 9594 2160 9595 2224
rect 9659 2160 9660 2224
rect 9594 2144 9660 2160
rect 9594 2080 9595 2144
rect 9659 2080 9660 2144
rect 9594 2064 9660 2080
rect 9594 2000 9595 2064
rect 9659 2000 9660 2064
rect 9594 1984 9660 2000
rect 9594 1920 9595 1984
rect 9659 1920 9660 1984
rect 9594 1904 9660 1920
rect 9594 1840 9595 1904
rect 9659 1840 9660 1904
rect 9594 1824 9660 1840
rect 9594 1760 9595 1824
rect 9659 1760 9660 1824
rect 9594 1744 9660 1760
rect 9594 1680 9595 1744
rect 9659 1680 9660 1744
rect 9594 1664 9660 1680
rect 9594 1600 9595 1664
rect 9659 1600 9660 1664
rect 9594 1446 9660 1600
rect 9720 1446 9780 2478
rect 9840 1508 9900 2538
rect 9960 1446 10020 2478
rect 10080 1508 10140 2538
rect 10200 2453 10266 2474
rect 10200 2397 10205 2453
rect 10261 2397 10266 2453
rect 10200 2384 10266 2397
rect 10200 2320 10201 2384
rect 10265 2320 10266 2384
rect 10200 2304 10266 2320
rect 10200 2240 10201 2304
rect 10265 2240 10266 2304
rect 10200 2224 10266 2240
rect 10200 2160 10201 2224
rect 10265 2160 10266 2224
rect 10200 2144 10266 2160
rect 10200 2080 10201 2144
rect 10265 2080 10266 2144
rect 10200 2064 10266 2080
rect 10200 2000 10201 2064
rect 10265 2000 10266 2064
rect 10200 1984 10266 2000
rect 10200 1920 10201 1984
rect 10265 1920 10266 1984
rect 10200 1904 10266 1920
rect 10200 1840 10201 1904
rect 10265 1840 10266 1904
rect 10200 1824 10266 1840
rect 10200 1760 10201 1824
rect 10265 1760 10266 1824
rect 10200 1744 10266 1760
rect 10200 1680 10201 1744
rect 10265 1680 10266 1744
rect 10200 1664 10266 1680
rect 10200 1600 10201 1664
rect 10265 1600 10266 1664
rect 10200 1446 10266 1600
rect 5352 1444 10266 1446
rect 5352 1380 5456 1444
rect 5520 1380 5536 1444
rect 5600 1380 5616 1444
rect 5680 1380 5696 1444
rect 5760 1380 5776 1444
rect 5840 1380 5856 1444
rect 5920 1380 6062 1444
rect 6126 1380 6142 1444
rect 6206 1380 6222 1444
rect 6286 1380 6302 1444
rect 6366 1380 6382 1444
rect 6446 1380 6462 1444
rect 6526 1380 6668 1444
rect 6732 1380 6748 1444
rect 6812 1380 6828 1444
rect 6892 1380 6908 1444
rect 6972 1380 6988 1444
rect 7052 1380 7068 1444
rect 7132 1380 7274 1444
rect 7338 1380 7354 1444
rect 7418 1380 7434 1444
rect 7498 1380 7514 1444
rect 7578 1380 7594 1444
rect 7658 1380 7674 1444
rect 7738 1380 7880 1444
rect 7944 1380 7960 1444
rect 8024 1380 8040 1444
rect 8104 1380 8120 1444
rect 8184 1380 8200 1444
rect 8264 1380 8280 1444
rect 8344 1380 8486 1444
rect 8550 1380 8566 1444
rect 8630 1380 8646 1444
rect 8710 1380 8726 1444
rect 8790 1380 8806 1444
rect 8870 1380 8886 1444
rect 8950 1380 9092 1444
rect 9156 1380 9172 1444
rect 9236 1380 9252 1444
rect 9316 1380 9332 1444
rect 9396 1380 9412 1444
rect 9476 1380 9492 1444
rect 9556 1380 9698 1444
rect 9762 1380 9778 1444
rect 9842 1380 9858 1444
rect 9922 1380 9938 1444
rect 10002 1380 10018 1444
rect 10082 1380 10098 1444
rect 10162 1380 10266 1444
rect 5352 1378 10266 1380
rect 5352 1224 5418 1378
rect 5352 1160 5353 1224
rect 5417 1160 5418 1224
rect 5352 1144 5418 1160
rect 5352 1080 5353 1144
rect 5417 1080 5418 1144
rect 5352 1064 5418 1080
rect 5352 1000 5353 1064
rect 5417 1000 5418 1064
rect 5352 984 5418 1000
rect 5352 920 5353 984
rect 5417 920 5418 984
rect 5352 904 5418 920
rect 5352 840 5353 904
rect 5417 840 5418 904
rect 5352 824 5418 840
rect 5352 760 5353 824
rect 5417 760 5418 824
rect 5352 744 5418 760
rect 5352 680 5353 744
rect 5417 680 5418 744
rect 5352 664 5418 680
rect 5352 600 5353 664
rect 5417 600 5418 664
rect 5352 584 5418 600
rect 5352 520 5353 584
rect 5417 520 5418 584
rect 5352 504 5418 520
rect 5352 440 5353 504
rect 5417 440 5418 504
rect 5352 350 5418 440
rect 5478 286 5538 1316
rect 5598 346 5658 1378
rect 5718 286 5778 1316
rect 5838 346 5898 1378
rect 5958 1224 6024 1378
rect 5958 1160 5959 1224
rect 6023 1160 6024 1224
rect 5958 1144 6024 1160
rect 5958 1080 5959 1144
rect 6023 1080 6024 1144
rect 5958 1064 6024 1080
rect 5958 1000 5959 1064
rect 6023 1000 6024 1064
rect 5958 984 6024 1000
rect 5958 920 5959 984
rect 6023 920 6024 984
rect 5958 904 6024 920
rect 5958 840 5959 904
rect 6023 840 6024 904
rect 5958 824 6024 840
rect 5958 760 5959 824
rect 6023 760 6024 824
rect 5958 744 6024 760
rect 5958 680 5959 744
rect 6023 680 6024 744
rect 5958 664 6024 680
rect 5958 600 5959 664
rect 6023 600 6024 664
rect 5958 584 6024 600
rect 5958 520 5959 584
rect 6023 520 6024 584
rect 5958 504 6024 520
rect 5958 440 5959 504
rect 6023 440 6024 504
rect 5958 350 6024 440
rect 6084 286 6144 1316
rect 6204 346 6264 1378
rect 6324 286 6384 1316
rect 6444 346 6504 1378
rect 6564 1224 6630 1378
rect 6564 1160 6565 1224
rect 6629 1160 6630 1224
rect 6564 1144 6630 1160
rect 6564 1080 6565 1144
rect 6629 1080 6630 1144
rect 6564 1064 6630 1080
rect 6564 1000 6565 1064
rect 6629 1000 6630 1064
rect 6564 984 6630 1000
rect 6564 920 6565 984
rect 6629 920 6630 984
rect 6564 904 6630 920
rect 6564 840 6565 904
rect 6629 840 6630 904
rect 6564 824 6630 840
rect 6564 760 6565 824
rect 6629 760 6630 824
rect 6564 744 6630 760
rect 6564 680 6565 744
rect 6629 680 6630 744
rect 6564 664 6630 680
rect 6564 600 6565 664
rect 6629 600 6630 664
rect 6564 584 6630 600
rect 6564 520 6565 584
rect 6629 520 6630 584
rect 6564 504 6630 520
rect 6564 440 6565 504
rect 6629 440 6630 504
rect 6564 350 6630 440
rect 6690 286 6750 1316
rect 6810 346 6870 1378
rect 6930 286 6990 1316
rect 7050 346 7110 1378
rect 7170 1224 7236 1378
rect 7170 1160 7171 1224
rect 7235 1160 7236 1224
rect 7170 1144 7236 1160
rect 7170 1080 7171 1144
rect 7235 1080 7236 1144
rect 7170 1064 7236 1080
rect 7170 1000 7171 1064
rect 7235 1000 7236 1064
rect 7170 984 7236 1000
rect 7170 920 7171 984
rect 7235 920 7236 984
rect 7170 904 7236 920
rect 7170 840 7171 904
rect 7235 840 7236 904
rect 7170 824 7236 840
rect 7170 760 7171 824
rect 7235 760 7236 824
rect 7170 744 7236 760
rect 7170 680 7171 744
rect 7235 680 7236 744
rect 7170 664 7236 680
rect 7170 600 7171 664
rect 7235 600 7236 664
rect 7170 584 7236 600
rect 7170 520 7171 584
rect 7235 520 7236 584
rect 7170 504 7236 520
rect 7170 440 7171 504
rect 7235 440 7236 504
rect 7170 350 7236 440
rect 7296 286 7356 1316
rect 7416 346 7476 1378
rect 7536 286 7596 1316
rect 7656 346 7716 1378
rect 7776 1224 7842 1378
rect 7776 1160 7777 1224
rect 7841 1160 7842 1224
rect 7776 1144 7842 1160
rect 7776 1080 7777 1144
rect 7841 1080 7842 1144
rect 7776 1064 7842 1080
rect 7776 1000 7777 1064
rect 7841 1000 7842 1064
rect 7776 984 7842 1000
rect 7776 920 7777 984
rect 7841 920 7842 984
rect 7776 904 7842 920
rect 7776 840 7777 904
rect 7841 840 7842 904
rect 7776 824 7842 840
rect 7776 760 7777 824
rect 7841 760 7842 824
rect 7776 744 7842 760
rect 7776 680 7777 744
rect 7841 680 7842 744
rect 7776 664 7842 680
rect 7776 600 7777 664
rect 7841 600 7842 664
rect 7776 584 7842 600
rect 7776 520 7777 584
rect 7841 520 7842 584
rect 7776 504 7842 520
rect 7776 440 7777 504
rect 7841 440 7842 504
rect 7776 350 7842 440
rect 7902 286 7962 1316
rect 8022 346 8082 1378
rect 8142 286 8202 1316
rect 8262 346 8322 1378
rect 8382 1224 8448 1378
rect 8382 1160 8383 1224
rect 8447 1160 8448 1224
rect 8382 1144 8448 1160
rect 8382 1080 8383 1144
rect 8447 1080 8448 1144
rect 8382 1064 8448 1080
rect 8382 1000 8383 1064
rect 8447 1000 8448 1064
rect 8382 984 8448 1000
rect 8382 920 8383 984
rect 8447 920 8448 984
rect 8382 904 8448 920
rect 8382 840 8383 904
rect 8447 840 8448 904
rect 8382 824 8448 840
rect 8382 760 8383 824
rect 8447 760 8448 824
rect 8382 744 8448 760
rect 8382 680 8383 744
rect 8447 680 8448 744
rect 8382 664 8448 680
rect 8382 600 8383 664
rect 8447 600 8448 664
rect 8382 584 8448 600
rect 8382 520 8383 584
rect 8447 520 8448 584
rect 8382 504 8448 520
rect 8382 440 8383 504
rect 8447 440 8448 504
rect 8382 350 8448 440
rect 8508 286 8568 1316
rect 8628 346 8688 1378
rect 8748 286 8808 1316
rect 8868 346 8928 1378
rect 8988 1224 9054 1378
rect 8988 1160 8989 1224
rect 9053 1160 9054 1224
rect 8988 1144 9054 1160
rect 8988 1080 8989 1144
rect 9053 1080 9054 1144
rect 8988 1064 9054 1080
rect 8988 1000 8989 1064
rect 9053 1000 9054 1064
rect 8988 984 9054 1000
rect 8988 920 8989 984
rect 9053 920 9054 984
rect 8988 904 9054 920
rect 8988 840 8989 904
rect 9053 840 9054 904
rect 8988 824 9054 840
rect 8988 760 8989 824
rect 9053 760 9054 824
rect 8988 744 9054 760
rect 8988 680 8989 744
rect 9053 680 9054 744
rect 8988 664 9054 680
rect 8988 600 8989 664
rect 9053 600 9054 664
rect 8988 584 9054 600
rect 8988 520 8989 584
rect 9053 520 9054 584
rect 8988 504 9054 520
rect 8988 440 8989 504
rect 9053 440 9054 504
rect 8988 350 9054 440
rect 9114 286 9174 1316
rect 9234 346 9294 1378
rect 9354 286 9414 1316
rect 9474 346 9534 1378
rect 9594 1224 9660 1378
rect 9594 1160 9595 1224
rect 9659 1160 9660 1224
rect 9594 1144 9660 1160
rect 9594 1080 9595 1144
rect 9659 1080 9660 1144
rect 9594 1064 9660 1080
rect 9594 1000 9595 1064
rect 9659 1000 9660 1064
rect 9594 984 9660 1000
rect 9594 920 9595 984
rect 9659 920 9660 984
rect 9594 904 9660 920
rect 9594 840 9595 904
rect 9659 840 9660 904
rect 9594 824 9660 840
rect 9594 760 9595 824
rect 9659 760 9660 824
rect 9594 744 9660 760
rect 9594 680 9595 744
rect 9659 680 9660 744
rect 9594 664 9660 680
rect 9594 600 9595 664
rect 9659 600 9660 664
rect 9594 584 9660 600
rect 9594 520 9595 584
rect 9659 520 9660 584
rect 9594 504 9660 520
rect 9594 440 9595 504
rect 9659 440 9660 504
rect 9594 350 9660 440
rect 9720 286 9780 1316
rect 9840 346 9900 1378
rect 9960 286 10020 1316
rect 10080 346 10140 1378
rect 10200 1224 10266 1378
rect 10200 1160 10201 1224
rect 10265 1160 10266 1224
rect 10200 1144 10266 1160
rect 10200 1080 10201 1144
rect 10265 1080 10266 1144
rect 10200 1064 10266 1080
rect 10200 1000 10201 1064
rect 10265 1000 10266 1064
rect 10200 984 10266 1000
rect 10200 920 10201 984
rect 10265 920 10266 984
rect 10200 904 10266 920
rect 10200 840 10201 904
rect 10265 840 10266 904
rect 10200 824 10266 840
rect 10200 760 10201 824
rect 10265 760 10266 824
rect 10200 744 10266 760
rect 10200 680 10201 744
rect 10265 680 10266 744
rect 10200 664 10266 680
rect 10200 600 10201 664
rect 10265 600 10266 664
rect 10200 584 10266 600
rect 10200 520 10201 584
rect 10265 520 10266 584
rect 10200 504 10266 520
rect 10200 440 10201 504
rect 10265 440 10266 504
rect 10200 350 10266 440
rect 10326 2384 10392 2474
rect 10326 2320 10327 2384
rect 10391 2320 10392 2384
rect 10326 2304 10392 2320
rect 10326 2240 10327 2304
rect 10391 2240 10392 2304
rect 10326 2224 10392 2240
rect 10326 2160 10327 2224
rect 10391 2160 10392 2224
rect 10326 2144 10392 2160
rect 10326 2080 10327 2144
rect 10391 2080 10392 2144
rect 10326 2064 10392 2080
rect 10326 2000 10327 2064
rect 10391 2000 10392 2064
rect 10326 1984 10392 2000
rect 10326 1920 10327 1984
rect 10391 1920 10392 1984
rect 10326 1904 10392 1920
rect 10326 1840 10327 1904
rect 10391 1840 10392 1904
rect 10326 1824 10392 1840
rect 10326 1760 10327 1824
rect 10391 1760 10392 1824
rect 10326 1744 10392 1760
rect 10326 1680 10327 1744
rect 10391 1680 10392 1744
rect 10326 1664 10392 1680
rect 10326 1600 10327 1664
rect 10391 1600 10392 1664
rect 10326 1446 10392 1600
rect 10452 1446 10512 2478
rect 10572 1508 10632 2538
rect 10692 1446 10752 2478
rect 10812 1508 10872 2538
rect 10932 2384 10998 2474
rect 10932 2320 10933 2384
rect 10997 2320 10998 2384
rect 10932 2304 10998 2320
rect 10932 2240 10933 2304
rect 10997 2240 10998 2304
rect 10932 2224 10998 2240
rect 10932 2160 10933 2224
rect 10997 2160 10998 2224
rect 10932 2144 10998 2160
rect 10932 2080 10933 2144
rect 10997 2080 10998 2144
rect 10932 2064 10998 2080
rect 10932 2000 10933 2064
rect 10997 2000 10998 2064
rect 10932 1984 10998 2000
rect 10932 1920 10933 1984
rect 10997 1920 10998 1984
rect 10932 1904 10998 1920
rect 10932 1840 10933 1904
rect 10997 1840 10998 1904
rect 10932 1824 10998 1840
rect 10932 1760 10933 1824
rect 10997 1760 10998 1824
rect 10932 1744 10998 1760
rect 10932 1680 10933 1744
rect 10997 1680 10998 1744
rect 10932 1664 10998 1680
rect 10932 1600 10933 1664
rect 10997 1600 10998 1664
rect 10932 1446 10998 1600
rect 11058 1446 11118 2478
rect 11178 1508 11238 2538
rect 11298 1446 11358 2478
rect 11418 1508 11478 2538
rect 11538 2384 11604 2474
rect 11538 2320 11539 2384
rect 11603 2320 11604 2384
rect 11538 2304 11604 2320
rect 11538 2240 11539 2304
rect 11603 2240 11604 2304
rect 11538 2224 11604 2240
rect 11538 2160 11539 2224
rect 11603 2160 11604 2224
rect 11538 2144 11604 2160
rect 11538 2080 11539 2144
rect 11603 2080 11604 2144
rect 11538 2064 11604 2080
rect 11538 2000 11539 2064
rect 11603 2000 11604 2064
rect 11538 1984 11604 2000
rect 11538 1920 11539 1984
rect 11603 1920 11604 1984
rect 11538 1904 11604 1920
rect 11538 1840 11539 1904
rect 11603 1840 11604 1904
rect 11538 1824 11604 1840
rect 11538 1760 11539 1824
rect 11603 1760 11604 1824
rect 11538 1744 11604 1760
rect 11538 1680 11539 1744
rect 11603 1680 11604 1744
rect 11538 1664 11604 1680
rect 11538 1600 11539 1664
rect 11603 1600 11604 1664
rect 11538 1446 11604 1600
rect 11664 1446 11724 2478
rect 11784 1508 11844 2538
rect 11904 1446 11964 2478
rect 12024 1508 12084 2538
rect 12144 2384 12210 2474
rect 12144 2320 12145 2384
rect 12209 2320 12210 2384
rect 12144 2304 12210 2320
rect 12144 2240 12145 2304
rect 12209 2240 12210 2304
rect 12144 2224 12210 2240
rect 12144 2160 12145 2224
rect 12209 2160 12210 2224
rect 12144 2144 12210 2160
rect 12144 2080 12145 2144
rect 12209 2080 12210 2144
rect 12144 2064 12210 2080
rect 12144 2000 12145 2064
rect 12209 2000 12210 2064
rect 12144 1984 12210 2000
rect 12144 1920 12145 1984
rect 12209 1920 12210 1984
rect 12144 1904 12210 1920
rect 12144 1840 12145 1904
rect 12209 1840 12210 1904
rect 12144 1824 12210 1840
rect 12144 1760 12145 1824
rect 12209 1760 12210 1824
rect 12144 1744 12210 1760
rect 12144 1680 12145 1744
rect 12209 1680 12210 1744
rect 12144 1664 12210 1680
rect 12144 1600 12145 1664
rect 12209 1600 12210 1664
rect 12144 1446 12210 1600
rect 12270 1446 12330 2478
rect 12390 1508 12450 2538
rect 12510 1446 12570 2478
rect 12630 1508 12690 2538
rect 12750 2384 12816 2474
rect 12750 2320 12751 2384
rect 12815 2320 12816 2384
rect 12750 2304 12816 2320
rect 12750 2240 12751 2304
rect 12815 2240 12816 2304
rect 12750 2224 12816 2240
rect 12750 2160 12751 2224
rect 12815 2160 12816 2224
rect 12750 2144 12816 2160
rect 12750 2080 12751 2144
rect 12815 2080 12816 2144
rect 12750 2064 12816 2080
rect 12750 2000 12751 2064
rect 12815 2000 12816 2064
rect 12750 1984 12816 2000
rect 12750 1920 12751 1984
rect 12815 1920 12816 1984
rect 12750 1904 12816 1920
rect 12750 1840 12751 1904
rect 12815 1840 12816 1904
rect 12750 1824 12816 1840
rect 12750 1760 12751 1824
rect 12815 1760 12816 1824
rect 12750 1744 12816 1760
rect 12750 1680 12751 1744
rect 12815 1680 12816 1744
rect 12750 1664 12816 1680
rect 12750 1600 12751 1664
rect 12815 1600 12816 1664
rect 12750 1446 12816 1600
rect 12876 1446 12936 2478
rect 12996 1508 13056 2538
rect 13116 1446 13176 2478
rect 13236 1508 13296 2538
rect 13356 2384 13422 2474
rect 13356 2320 13357 2384
rect 13421 2320 13422 2384
rect 13356 2304 13422 2320
rect 13356 2240 13357 2304
rect 13421 2240 13422 2304
rect 13356 2224 13422 2240
rect 13356 2160 13357 2224
rect 13421 2160 13422 2224
rect 13356 2144 13422 2160
rect 13356 2080 13357 2144
rect 13421 2080 13422 2144
rect 13356 2064 13422 2080
rect 13356 2000 13357 2064
rect 13421 2000 13422 2064
rect 13356 1984 13422 2000
rect 13356 1920 13357 1984
rect 13421 1920 13422 1984
rect 13356 1904 13422 1920
rect 13356 1840 13357 1904
rect 13421 1840 13422 1904
rect 13356 1824 13422 1840
rect 13356 1760 13357 1824
rect 13421 1760 13422 1824
rect 13356 1744 13422 1760
rect 13356 1680 13357 1744
rect 13421 1680 13422 1744
rect 13356 1664 13422 1680
rect 13356 1600 13357 1664
rect 13421 1600 13422 1664
rect 13356 1446 13422 1600
rect 13482 1446 13542 2478
rect 13602 1508 13662 2538
rect 13722 1446 13782 2478
rect 13842 1508 13902 2538
rect 13962 2384 14028 2474
rect 13962 2320 13963 2384
rect 14027 2320 14028 2384
rect 13962 2304 14028 2320
rect 13962 2240 13963 2304
rect 14027 2240 14028 2304
rect 13962 2224 14028 2240
rect 13962 2160 13963 2224
rect 14027 2160 14028 2224
rect 13962 2144 14028 2160
rect 13962 2080 13963 2144
rect 14027 2080 14028 2144
rect 13962 2064 14028 2080
rect 13962 2000 13963 2064
rect 14027 2000 14028 2064
rect 13962 1984 14028 2000
rect 13962 1920 13963 1984
rect 14027 1920 14028 1984
rect 13962 1904 14028 1920
rect 13962 1840 13963 1904
rect 14027 1840 14028 1904
rect 13962 1824 14028 1840
rect 13962 1760 13963 1824
rect 14027 1760 14028 1824
rect 13962 1744 14028 1760
rect 13962 1680 13963 1744
rect 14027 1680 14028 1744
rect 13962 1664 14028 1680
rect 13962 1600 13963 1664
rect 14027 1600 14028 1664
rect 13962 1446 14028 1600
rect 14088 1446 14148 2478
rect 14208 1508 14268 2538
rect 14328 1446 14388 2478
rect 14448 1508 14508 2538
rect 14568 2384 14634 2474
rect 14568 2320 14569 2384
rect 14633 2320 14634 2384
rect 14568 2304 14634 2320
rect 14568 2240 14569 2304
rect 14633 2240 14634 2304
rect 14568 2224 14634 2240
rect 14568 2160 14569 2224
rect 14633 2160 14634 2224
rect 14568 2144 14634 2160
rect 14568 2080 14569 2144
rect 14633 2080 14634 2144
rect 14568 2064 14634 2080
rect 14568 2000 14569 2064
rect 14633 2000 14634 2064
rect 14568 1984 14634 2000
rect 14568 1920 14569 1984
rect 14633 1920 14634 1984
rect 14568 1904 14634 1920
rect 14568 1840 14569 1904
rect 14633 1840 14634 1904
rect 14568 1824 14634 1840
rect 14568 1760 14569 1824
rect 14633 1760 14634 1824
rect 14568 1744 14634 1760
rect 14568 1680 14569 1744
rect 14633 1680 14634 1744
rect 14568 1664 14634 1680
rect 14568 1600 14569 1664
rect 14633 1600 14634 1664
rect 14568 1446 14634 1600
rect 14694 1446 14754 2478
rect 14814 1508 14874 2538
rect 14934 1446 14994 2478
rect 15054 1508 15114 2538
rect 15174 2384 15240 2474
rect 15174 2320 15175 2384
rect 15239 2320 15240 2384
rect 15174 2304 15240 2320
rect 15174 2240 15175 2304
rect 15239 2240 15240 2304
rect 15174 2224 15240 2240
rect 15174 2160 15175 2224
rect 15239 2160 15240 2224
rect 15174 2144 15240 2160
rect 15174 2080 15175 2144
rect 15239 2080 15240 2144
rect 15174 2064 15240 2080
rect 15174 2000 15175 2064
rect 15239 2000 15240 2064
rect 15174 1984 15240 2000
rect 15174 1920 15175 1984
rect 15239 1920 15240 1984
rect 15174 1904 15240 1920
rect 15174 1840 15175 1904
rect 15239 1840 15240 1904
rect 15174 1824 15240 1840
rect 15174 1760 15175 1824
rect 15239 1760 15240 1824
rect 15174 1744 15240 1760
rect 15174 1680 15175 1744
rect 15239 1680 15240 1744
rect 15174 1664 15240 1680
rect 15174 1600 15175 1664
rect 15239 1600 15240 1664
rect 15174 1446 15240 1600
rect 15300 1446 15360 2478
rect 15420 1508 15480 2538
rect 15540 1446 15600 2478
rect 15660 1508 15720 2538
rect 15780 2384 15846 2474
rect 15780 2320 15781 2384
rect 15845 2320 15846 2384
rect 15780 2304 15846 2320
rect 15780 2240 15781 2304
rect 15845 2240 15846 2304
rect 15780 2224 15846 2240
rect 15780 2160 15781 2224
rect 15845 2160 15846 2224
rect 15780 2144 15846 2160
rect 15780 2080 15781 2144
rect 15845 2080 15846 2144
rect 15780 2064 15846 2080
rect 15780 2000 15781 2064
rect 15845 2000 15846 2064
rect 15780 1984 15846 2000
rect 15780 1920 15781 1984
rect 15845 1920 15846 1984
rect 15780 1904 15846 1920
rect 15780 1840 15781 1904
rect 15845 1840 15846 1904
rect 15780 1824 15846 1840
rect 15780 1760 15781 1824
rect 15845 1760 15846 1824
rect 15780 1744 15846 1760
rect 15780 1680 15781 1744
rect 15845 1680 15846 1744
rect 15780 1664 15846 1680
rect 15780 1600 15781 1664
rect 15845 1600 15846 1664
rect 15780 1446 15846 1600
rect 15906 1446 15966 2478
rect 16026 1508 16086 2538
rect 16146 1446 16206 2478
rect 16266 1508 16326 2538
rect 16386 2384 16452 2474
rect 16386 2320 16387 2384
rect 16451 2320 16452 2384
rect 16386 2304 16452 2320
rect 16386 2240 16387 2304
rect 16451 2240 16452 2304
rect 16386 2224 16452 2240
rect 16386 2160 16387 2224
rect 16451 2160 16452 2224
rect 16386 2144 16452 2160
rect 16386 2080 16387 2144
rect 16451 2080 16452 2144
rect 16386 2064 16452 2080
rect 16386 2000 16387 2064
rect 16451 2000 16452 2064
rect 16386 1984 16452 2000
rect 16386 1920 16387 1984
rect 16451 1920 16452 1984
rect 16386 1904 16452 1920
rect 16386 1840 16387 1904
rect 16451 1840 16452 1904
rect 16386 1824 16452 1840
rect 16386 1760 16387 1824
rect 16451 1760 16452 1824
rect 16386 1744 16452 1760
rect 16386 1680 16387 1744
rect 16451 1680 16452 1744
rect 16386 1664 16452 1680
rect 16386 1600 16387 1664
rect 16451 1600 16452 1664
rect 16386 1446 16452 1600
rect 16512 1446 16572 2478
rect 16632 1508 16692 2538
rect 16752 1446 16812 2478
rect 16872 1508 16932 2538
rect 16992 2384 17058 2474
rect 16992 2320 16993 2384
rect 17057 2320 17058 2384
rect 16992 2304 17058 2320
rect 16992 2240 16993 2304
rect 17057 2240 17058 2304
rect 16992 2224 17058 2240
rect 16992 2160 16993 2224
rect 17057 2160 17058 2224
rect 16992 2144 17058 2160
rect 16992 2080 16993 2144
rect 17057 2080 17058 2144
rect 16992 2064 17058 2080
rect 16992 2000 16993 2064
rect 17057 2000 17058 2064
rect 16992 1984 17058 2000
rect 16992 1920 16993 1984
rect 17057 1920 17058 1984
rect 16992 1904 17058 1920
rect 16992 1840 16993 1904
rect 17057 1840 17058 1904
rect 16992 1824 17058 1840
rect 16992 1760 16993 1824
rect 17057 1760 17058 1824
rect 16992 1744 17058 1760
rect 16992 1680 16993 1744
rect 17057 1680 17058 1744
rect 16992 1664 17058 1680
rect 16992 1600 16993 1664
rect 17057 1600 17058 1664
rect 16992 1446 17058 1600
rect 17118 1446 17178 2478
rect 17238 1508 17298 2538
rect 17358 1446 17418 2478
rect 17478 1508 17538 2538
rect 17598 2384 17664 2474
rect 17598 2320 17599 2384
rect 17663 2320 17664 2384
rect 17598 2304 17664 2320
rect 17598 2240 17599 2304
rect 17663 2240 17664 2304
rect 17598 2224 17664 2240
rect 17598 2160 17599 2224
rect 17663 2160 17664 2224
rect 17598 2144 17664 2160
rect 17598 2080 17599 2144
rect 17663 2080 17664 2144
rect 17598 2064 17664 2080
rect 17598 2000 17599 2064
rect 17663 2000 17664 2064
rect 17598 1984 17664 2000
rect 17598 1920 17599 1984
rect 17663 1920 17664 1984
rect 17598 1904 17664 1920
rect 17598 1840 17599 1904
rect 17663 1840 17664 1904
rect 17598 1824 17664 1840
rect 17598 1760 17599 1824
rect 17663 1760 17664 1824
rect 17598 1744 17664 1760
rect 17598 1680 17599 1744
rect 17663 1680 17664 1744
rect 17598 1664 17664 1680
rect 17598 1600 17599 1664
rect 17663 1600 17664 1664
rect 17598 1446 17664 1600
rect 17724 1446 17784 2478
rect 17844 1508 17904 2538
rect 17964 1446 18024 2478
rect 18084 1508 18144 2538
rect 18204 2384 18270 2474
rect 18204 2320 18205 2384
rect 18269 2320 18270 2384
rect 18204 2304 18270 2320
rect 18204 2240 18205 2304
rect 18269 2240 18270 2304
rect 18204 2224 18270 2240
rect 18204 2160 18205 2224
rect 18269 2160 18270 2224
rect 18204 2144 18270 2160
rect 18204 2080 18205 2144
rect 18269 2080 18270 2144
rect 18204 2064 18270 2080
rect 18204 2000 18205 2064
rect 18269 2000 18270 2064
rect 18204 1984 18270 2000
rect 18204 1920 18205 1984
rect 18269 1920 18270 1984
rect 18204 1904 18270 1920
rect 18204 1840 18205 1904
rect 18269 1840 18270 1904
rect 18204 1824 18270 1840
rect 18204 1760 18205 1824
rect 18269 1760 18270 1824
rect 18204 1744 18270 1760
rect 18204 1680 18205 1744
rect 18269 1680 18270 1744
rect 18204 1664 18270 1680
rect 18204 1600 18205 1664
rect 18269 1600 18270 1664
rect 18204 1446 18270 1600
rect 18330 1446 18390 2478
rect 18450 1508 18510 2538
rect 18570 1446 18630 2478
rect 18690 1508 18750 2538
rect 18810 2384 18876 2474
rect 18810 2320 18811 2384
rect 18875 2320 18876 2384
rect 18810 2304 18876 2320
rect 18810 2240 18811 2304
rect 18875 2240 18876 2304
rect 18810 2224 18876 2240
rect 18810 2160 18811 2224
rect 18875 2160 18876 2224
rect 18810 2144 18876 2160
rect 18810 2080 18811 2144
rect 18875 2080 18876 2144
rect 18810 2064 18876 2080
rect 18810 2000 18811 2064
rect 18875 2000 18876 2064
rect 18810 1984 18876 2000
rect 18810 1920 18811 1984
rect 18875 1920 18876 1984
rect 18810 1904 18876 1920
rect 18810 1840 18811 1904
rect 18875 1840 18876 1904
rect 18810 1824 18876 1840
rect 18810 1760 18811 1824
rect 18875 1760 18876 1824
rect 18810 1744 18876 1760
rect 18810 1680 18811 1744
rect 18875 1680 18876 1744
rect 18810 1664 18876 1680
rect 18810 1600 18811 1664
rect 18875 1600 18876 1664
rect 18810 1446 18876 1600
rect 18936 1446 18996 2478
rect 19056 1508 19116 2538
rect 19176 1446 19236 2478
rect 19296 1508 19356 2538
rect 19416 2461 19482 2474
rect 19416 2405 19421 2461
rect 19477 2405 19482 2461
rect 19416 2384 19482 2405
rect 19416 2320 19417 2384
rect 19481 2320 19482 2384
rect 19416 2304 19482 2320
rect 19416 2240 19417 2304
rect 19481 2240 19482 2304
rect 19416 2224 19482 2240
rect 19416 2160 19417 2224
rect 19481 2160 19482 2224
rect 19416 2144 19482 2160
rect 19416 2080 19417 2144
rect 19481 2080 19482 2144
rect 19416 2064 19482 2080
rect 19416 2000 19417 2064
rect 19481 2000 19482 2064
rect 19416 1984 19482 2000
rect 19416 1920 19417 1984
rect 19481 1920 19482 1984
rect 19416 1904 19482 1920
rect 19416 1840 19417 1904
rect 19481 1840 19482 1904
rect 19416 1824 19482 1840
rect 19416 1760 19417 1824
rect 19481 1760 19482 1824
rect 19416 1744 19482 1760
rect 19416 1680 19417 1744
rect 19481 1680 19482 1744
rect 19416 1664 19482 1680
rect 19416 1600 19417 1664
rect 19481 1600 19482 1664
rect 19416 1446 19482 1600
rect 19542 1446 19602 2478
rect 19662 1508 19722 2538
rect 19782 1446 19842 2478
rect 19902 1508 19962 2538
rect 20022 2384 20088 2474
rect 20022 2320 20023 2384
rect 20087 2320 20088 2384
rect 20022 2304 20088 2320
rect 20022 2240 20023 2304
rect 20087 2240 20088 2304
rect 20022 2224 20088 2240
rect 20022 2160 20023 2224
rect 20087 2160 20088 2224
rect 20022 2144 20088 2160
rect 20022 2080 20023 2144
rect 20087 2080 20088 2144
rect 20022 2064 20088 2080
rect 20022 2000 20023 2064
rect 20087 2000 20088 2064
rect 20022 1984 20088 2000
rect 20022 1920 20023 1984
rect 20087 1920 20088 1984
rect 20022 1904 20088 1920
rect 20022 1840 20023 1904
rect 20087 1840 20088 1904
rect 20022 1824 20088 1840
rect 20022 1760 20023 1824
rect 20087 1760 20088 1824
rect 20022 1744 20088 1760
rect 20022 1680 20023 1744
rect 20087 1680 20088 1744
rect 20022 1664 20088 1680
rect 20022 1600 20023 1664
rect 20087 1600 20088 1664
rect 20022 1446 20088 1600
rect 10326 1444 20088 1446
rect 10326 1380 10430 1444
rect 10494 1380 10510 1444
rect 10574 1380 10590 1444
rect 10654 1380 10670 1444
rect 10734 1380 10750 1444
rect 10814 1380 10830 1444
rect 10894 1380 11036 1444
rect 11100 1380 11116 1444
rect 11180 1380 11196 1444
rect 11260 1380 11276 1444
rect 11340 1380 11356 1444
rect 11420 1380 11436 1444
rect 11500 1380 11642 1444
rect 11706 1380 11722 1444
rect 11786 1380 11802 1444
rect 11866 1380 11882 1444
rect 11946 1380 11962 1444
rect 12026 1380 12042 1444
rect 12106 1380 12248 1444
rect 12312 1380 12328 1444
rect 12392 1380 12408 1444
rect 12472 1380 12488 1444
rect 12552 1380 12568 1444
rect 12632 1380 12648 1444
rect 12712 1380 12854 1444
rect 12918 1380 12934 1444
rect 12998 1380 13014 1444
rect 13078 1380 13094 1444
rect 13158 1380 13174 1444
rect 13238 1380 13254 1444
rect 13318 1380 13460 1444
rect 13524 1380 13540 1444
rect 13604 1380 13620 1444
rect 13684 1380 13700 1444
rect 13764 1380 13780 1444
rect 13844 1380 13860 1444
rect 13924 1380 14066 1444
rect 14130 1380 14146 1444
rect 14210 1380 14226 1444
rect 14290 1380 14306 1444
rect 14370 1380 14386 1444
rect 14450 1380 14466 1444
rect 14530 1380 14672 1444
rect 14736 1380 14752 1444
rect 14816 1380 14832 1444
rect 14896 1380 14912 1444
rect 14976 1380 14992 1444
rect 15056 1380 15072 1444
rect 15136 1380 15278 1444
rect 15342 1380 15358 1444
rect 15422 1380 15438 1444
rect 15502 1380 15518 1444
rect 15582 1380 15598 1444
rect 15662 1380 15678 1444
rect 15742 1380 15884 1444
rect 15948 1380 15964 1444
rect 16028 1380 16044 1444
rect 16108 1380 16124 1444
rect 16188 1380 16204 1444
rect 16268 1380 16284 1444
rect 16348 1380 16490 1444
rect 16554 1380 16570 1444
rect 16634 1380 16650 1444
rect 16714 1380 16730 1444
rect 16794 1380 16810 1444
rect 16874 1380 16890 1444
rect 16954 1380 17096 1444
rect 17160 1380 17176 1444
rect 17240 1380 17256 1444
rect 17320 1380 17336 1444
rect 17400 1380 17416 1444
rect 17480 1380 17496 1444
rect 17560 1380 17702 1444
rect 17766 1380 17782 1444
rect 17846 1380 17862 1444
rect 17926 1380 17942 1444
rect 18006 1380 18022 1444
rect 18086 1380 18102 1444
rect 18166 1380 18308 1444
rect 18372 1380 18388 1444
rect 18452 1380 18468 1444
rect 18532 1380 18548 1444
rect 18612 1380 18628 1444
rect 18692 1380 18708 1444
rect 18772 1380 18914 1444
rect 18978 1380 18994 1444
rect 19058 1380 19074 1444
rect 19138 1380 19154 1444
rect 19218 1380 19234 1444
rect 19298 1380 19314 1444
rect 19378 1380 19520 1444
rect 19584 1380 19600 1444
rect 19664 1380 19680 1444
rect 19744 1380 19760 1444
rect 19824 1380 19840 1444
rect 19904 1380 19920 1444
rect 19984 1380 20088 1444
rect 10326 1378 20088 1380
rect 10326 1224 10392 1378
rect 10326 1160 10327 1224
rect 10391 1160 10392 1224
rect 10326 1144 10392 1160
rect 10326 1080 10327 1144
rect 10391 1080 10392 1144
rect 10326 1064 10392 1080
rect 10326 1000 10327 1064
rect 10391 1000 10392 1064
rect 10326 984 10392 1000
rect 10326 920 10327 984
rect 10391 920 10392 984
rect 10326 904 10392 920
rect 10326 840 10327 904
rect 10391 840 10392 904
rect 10326 824 10392 840
rect 10326 760 10327 824
rect 10391 760 10392 824
rect 10326 744 10392 760
rect 10326 680 10327 744
rect 10391 680 10392 744
rect 10326 664 10392 680
rect 10326 600 10327 664
rect 10391 600 10392 664
rect 10326 584 10392 600
rect 10326 520 10327 584
rect 10391 520 10392 584
rect 10326 504 10392 520
rect 10326 440 10327 504
rect 10391 440 10392 504
rect 10326 350 10392 440
rect 10452 286 10512 1316
rect 10572 346 10632 1378
rect 10692 286 10752 1316
rect 10812 346 10872 1378
rect 10932 1224 10998 1378
rect 10932 1160 10933 1224
rect 10997 1160 10998 1224
rect 10932 1144 10998 1160
rect 10932 1080 10933 1144
rect 10997 1080 10998 1144
rect 10932 1064 10998 1080
rect 10932 1000 10933 1064
rect 10997 1000 10998 1064
rect 10932 984 10998 1000
rect 10932 920 10933 984
rect 10997 920 10998 984
rect 10932 904 10998 920
rect 10932 840 10933 904
rect 10997 840 10998 904
rect 10932 824 10998 840
rect 10932 760 10933 824
rect 10997 760 10998 824
rect 10932 744 10998 760
rect 10932 680 10933 744
rect 10997 680 10998 744
rect 10932 664 10998 680
rect 10932 600 10933 664
rect 10997 600 10998 664
rect 10932 584 10998 600
rect 10932 520 10933 584
rect 10997 520 10998 584
rect 10932 504 10998 520
rect 10932 440 10933 504
rect 10997 440 10998 504
rect 10932 350 10998 440
rect 11058 286 11118 1316
rect 11178 346 11238 1378
rect 11298 286 11358 1316
rect 11418 346 11478 1378
rect 11538 1224 11604 1378
rect 11538 1160 11539 1224
rect 11603 1160 11604 1224
rect 11538 1144 11604 1160
rect 11538 1080 11539 1144
rect 11603 1080 11604 1144
rect 11538 1064 11604 1080
rect 11538 1000 11539 1064
rect 11603 1000 11604 1064
rect 11538 984 11604 1000
rect 11538 920 11539 984
rect 11603 920 11604 984
rect 11538 904 11604 920
rect 11538 840 11539 904
rect 11603 840 11604 904
rect 11538 824 11604 840
rect 11538 760 11539 824
rect 11603 760 11604 824
rect 11538 744 11604 760
rect 11538 680 11539 744
rect 11603 680 11604 744
rect 11538 664 11604 680
rect 11538 600 11539 664
rect 11603 600 11604 664
rect 11538 584 11604 600
rect 11538 520 11539 584
rect 11603 520 11604 584
rect 11538 504 11604 520
rect 11538 440 11539 504
rect 11603 440 11604 504
rect 11538 350 11604 440
rect 11664 286 11724 1316
rect 11784 346 11844 1378
rect 11904 286 11964 1316
rect 12024 346 12084 1378
rect 12144 1224 12210 1378
rect 12144 1160 12145 1224
rect 12209 1160 12210 1224
rect 12144 1144 12210 1160
rect 12144 1080 12145 1144
rect 12209 1080 12210 1144
rect 12144 1064 12210 1080
rect 12144 1000 12145 1064
rect 12209 1000 12210 1064
rect 12144 984 12210 1000
rect 12144 920 12145 984
rect 12209 920 12210 984
rect 12144 904 12210 920
rect 12144 840 12145 904
rect 12209 840 12210 904
rect 12144 824 12210 840
rect 12144 760 12145 824
rect 12209 760 12210 824
rect 12144 744 12210 760
rect 12144 680 12145 744
rect 12209 680 12210 744
rect 12144 664 12210 680
rect 12144 600 12145 664
rect 12209 600 12210 664
rect 12144 584 12210 600
rect 12144 520 12145 584
rect 12209 520 12210 584
rect 12144 504 12210 520
rect 12144 440 12145 504
rect 12209 440 12210 504
rect 12144 350 12210 440
rect 12270 286 12330 1316
rect 12390 346 12450 1378
rect 12510 286 12570 1316
rect 12630 346 12690 1378
rect 12750 1224 12816 1378
rect 12750 1160 12751 1224
rect 12815 1160 12816 1224
rect 12750 1144 12816 1160
rect 12750 1080 12751 1144
rect 12815 1080 12816 1144
rect 12750 1064 12816 1080
rect 12750 1000 12751 1064
rect 12815 1000 12816 1064
rect 12750 984 12816 1000
rect 12750 920 12751 984
rect 12815 920 12816 984
rect 12750 904 12816 920
rect 12750 840 12751 904
rect 12815 840 12816 904
rect 12750 824 12816 840
rect 12750 760 12751 824
rect 12815 760 12816 824
rect 12750 744 12816 760
rect 12750 680 12751 744
rect 12815 680 12816 744
rect 12750 664 12816 680
rect 12750 600 12751 664
rect 12815 600 12816 664
rect 12750 584 12816 600
rect 12750 520 12751 584
rect 12815 520 12816 584
rect 12750 504 12816 520
rect 12750 440 12751 504
rect 12815 440 12816 504
rect 12750 350 12816 440
rect 12876 286 12936 1316
rect 12996 346 13056 1378
rect 13116 286 13176 1316
rect 13236 346 13296 1378
rect 13356 1224 13422 1378
rect 13356 1160 13357 1224
rect 13421 1160 13422 1224
rect 13356 1144 13422 1160
rect 13356 1080 13357 1144
rect 13421 1080 13422 1144
rect 13356 1064 13422 1080
rect 13356 1000 13357 1064
rect 13421 1000 13422 1064
rect 13356 984 13422 1000
rect 13356 920 13357 984
rect 13421 920 13422 984
rect 13356 904 13422 920
rect 13356 840 13357 904
rect 13421 840 13422 904
rect 13356 824 13422 840
rect 13356 760 13357 824
rect 13421 760 13422 824
rect 13356 744 13422 760
rect 13356 680 13357 744
rect 13421 680 13422 744
rect 13356 664 13422 680
rect 13356 600 13357 664
rect 13421 600 13422 664
rect 13356 584 13422 600
rect 13356 520 13357 584
rect 13421 520 13422 584
rect 13356 504 13422 520
rect 13356 440 13357 504
rect 13421 440 13422 504
rect 13356 350 13422 440
rect 13482 286 13542 1316
rect 13602 346 13662 1378
rect 13722 286 13782 1316
rect 13842 346 13902 1378
rect 13962 1224 14028 1378
rect 13962 1160 13963 1224
rect 14027 1160 14028 1224
rect 13962 1144 14028 1160
rect 13962 1080 13963 1144
rect 14027 1080 14028 1144
rect 13962 1064 14028 1080
rect 13962 1000 13963 1064
rect 14027 1000 14028 1064
rect 13962 984 14028 1000
rect 13962 920 13963 984
rect 14027 920 14028 984
rect 13962 904 14028 920
rect 13962 840 13963 904
rect 14027 840 14028 904
rect 13962 824 14028 840
rect 13962 760 13963 824
rect 14027 760 14028 824
rect 13962 744 14028 760
rect 13962 680 13963 744
rect 14027 680 14028 744
rect 13962 664 14028 680
rect 13962 600 13963 664
rect 14027 600 14028 664
rect 13962 584 14028 600
rect 13962 520 13963 584
rect 14027 520 14028 584
rect 13962 504 14028 520
rect 13962 440 13963 504
rect 14027 440 14028 504
rect 13962 350 14028 440
rect 14088 286 14148 1316
rect 14208 346 14268 1378
rect 14328 286 14388 1316
rect 14448 346 14508 1378
rect 14568 1224 14634 1378
rect 14568 1160 14569 1224
rect 14633 1160 14634 1224
rect 14568 1144 14634 1160
rect 14568 1080 14569 1144
rect 14633 1080 14634 1144
rect 14568 1064 14634 1080
rect 14568 1000 14569 1064
rect 14633 1000 14634 1064
rect 14568 984 14634 1000
rect 14568 920 14569 984
rect 14633 920 14634 984
rect 14568 904 14634 920
rect 14568 840 14569 904
rect 14633 840 14634 904
rect 14568 824 14634 840
rect 14568 760 14569 824
rect 14633 760 14634 824
rect 14568 744 14634 760
rect 14568 680 14569 744
rect 14633 680 14634 744
rect 14568 664 14634 680
rect 14568 600 14569 664
rect 14633 600 14634 664
rect 14568 584 14634 600
rect 14568 520 14569 584
rect 14633 520 14634 584
rect 14568 504 14634 520
rect 14568 440 14569 504
rect 14633 440 14634 504
rect 14568 350 14634 440
rect 14694 286 14754 1316
rect 14814 346 14874 1378
rect 14934 286 14994 1316
rect 15054 346 15114 1378
rect 15174 1224 15240 1378
rect 15174 1160 15175 1224
rect 15239 1160 15240 1224
rect 15174 1144 15240 1160
rect 15174 1080 15175 1144
rect 15239 1080 15240 1144
rect 15174 1064 15240 1080
rect 15174 1000 15175 1064
rect 15239 1000 15240 1064
rect 15174 984 15240 1000
rect 15174 920 15175 984
rect 15239 920 15240 984
rect 15174 904 15240 920
rect 15174 840 15175 904
rect 15239 840 15240 904
rect 15174 824 15240 840
rect 15174 760 15175 824
rect 15239 760 15240 824
rect 15174 744 15240 760
rect 15174 680 15175 744
rect 15239 680 15240 744
rect 15174 664 15240 680
rect 15174 600 15175 664
rect 15239 600 15240 664
rect 15174 584 15240 600
rect 15174 520 15175 584
rect 15239 520 15240 584
rect 15174 504 15240 520
rect 15174 440 15175 504
rect 15239 440 15240 504
rect 15174 350 15240 440
rect 15300 286 15360 1316
rect 15420 346 15480 1378
rect 15540 286 15600 1316
rect 15660 346 15720 1378
rect 15780 1224 15846 1378
rect 15780 1160 15781 1224
rect 15845 1160 15846 1224
rect 15780 1144 15846 1160
rect 15780 1080 15781 1144
rect 15845 1080 15846 1144
rect 15780 1064 15846 1080
rect 15780 1000 15781 1064
rect 15845 1000 15846 1064
rect 15780 984 15846 1000
rect 15780 920 15781 984
rect 15845 920 15846 984
rect 15780 904 15846 920
rect 15780 840 15781 904
rect 15845 840 15846 904
rect 15780 824 15846 840
rect 15780 760 15781 824
rect 15845 760 15846 824
rect 15780 744 15846 760
rect 15780 680 15781 744
rect 15845 680 15846 744
rect 15780 664 15846 680
rect 15780 600 15781 664
rect 15845 600 15846 664
rect 15780 584 15846 600
rect 15780 520 15781 584
rect 15845 520 15846 584
rect 15780 504 15846 520
rect 15780 440 15781 504
rect 15845 440 15846 504
rect 15780 350 15846 440
rect 15906 286 15966 1316
rect 16026 346 16086 1378
rect 16146 286 16206 1316
rect 16266 346 16326 1378
rect 16386 1224 16452 1378
rect 16386 1160 16387 1224
rect 16451 1160 16452 1224
rect 16386 1144 16452 1160
rect 16386 1080 16387 1144
rect 16451 1080 16452 1144
rect 16386 1064 16452 1080
rect 16386 1000 16387 1064
rect 16451 1000 16452 1064
rect 16386 984 16452 1000
rect 16386 920 16387 984
rect 16451 920 16452 984
rect 16386 904 16452 920
rect 16386 840 16387 904
rect 16451 840 16452 904
rect 16386 824 16452 840
rect 16386 760 16387 824
rect 16451 760 16452 824
rect 16386 744 16452 760
rect 16386 680 16387 744
rect 16451 680 16452 744
rect 16386 664 16452 680
rect 16386 600 16387 664
rect 16451 600 16452 664
rect 16386 584 16452 600
rect 16386 520 16387 584
rect 16451 520 16452 584
rect 16386 504 16452 520
rect 16386 440 16387 504
rect 16451 440 16452 504
rect 16386 350 16452 440
rect 16512 286 16572 1316
rect 16632 346 16692 1378
rect 16752 286 16812 1316
rect 16872 346 16932 1378
rect 16992 1224 17058 1378
rect 16992 1160 16993 1224
rect 17057 1160 17058 1224
rect 16992 1144 17058 1160
rect 16992 1080 16993 1144
rect 17057 1080 17058 1144
rect 16992 1064 17058 1080
rect 16992 1000 16993 1064
rect 17057 1000 17058 1064
rect 16992 984 17058 1000
rect 16992 920 16993 984
rect 17057 920 17058 984
rect 16992 904 17058 920
rect 16992 840 16993 904
rect 17057 840 17058 904
rect 16992 824 17058 840
rect 16992 760 16993 824
rect 17057 760 17058 824
rect 16992 744 17058 760
rect 16992 680 16993 744
rect 17057 680 17058 744
rect 16992 664 17058 680
rect 16992 600 16993 664
rect 17057 600 17058 664
rect 16992 584 17058 600
rect 16992 520 16993 584
rect 17057 520 17058 584
rect 16992 504 17058 520
rect 16992 440 16993 504
rect 17057 440 17058 504
rect 16992 350 17058 440
rect 17118 286 17178 1316
rect 17238 346 17298 1378
rect 17358 286 17418 1316
rect 17478 346 17538 1378
rect 17598 1224 17664 1378
rect 17598 1160 17599 1224
rect 17663 1160 17664 1224
rect 17598 1144 17664 1160
rect 17598 1080 17599 1144
rect 17663 1080 17664 1144
rect 17598 1064 17664 1080
rect 17598 1000 17599 1064
rect 17663 1000 17664 1064
rect 17598 984 17664 1000
rect 17598 920 17599 984
rect 17663 920 17664 984
rect 17598 904 17664 920
rect 17598 840 17599 904
rect 17663 840 17664 904
rect 17598 824 17664 840
rect 17598 760 17599 824
rect 17663 760 17664 824
rect 17598 744 17664 760
rect 17598 680 17599 744
rect 17663 680 17664 744
rect 17598 664 17664 680
rect 17598 600 17599 664
rect 17663 600 17664 664
rect 17598 584 17664 600
rect 17598 520 17599 584
rect 17663 520 17664 584
rect 17598 504 17664 520
rect 17598 440 17599 504
rect 17663 440 17664 504
rect 17598 350 17664 440
rect 17724 286 17784 1316
rect 17844 346 17904 1378
rect 17964 286 18024 1316
rect 18084 346 18144 1378
rect 18204 1224 18270 1378
rect 18204 1160 18205 1224
rect 18269 1160 18270 1224
rect 18204 1144 18270 1160
rect 18204 1080 18205 1144
rect 18269 1080 18270 1144
rect 18204 1064 18270 1080
rect 18204 1000 18205 1064
rect 18269 1000 18270 1064
rect 18204 984 18270 1000
rect 18204 920 18205 984
rect 18269 920 18270 984
rect 18204 904 18270 920
rect 18204 840 18205 904
rect 18269 840 18270 904
rect 18204 824 18270 840
rect 18204 760 18205 824
rect 18269 760 18270 824
rect 18204 744 18270 760
rect 18204 680 18205 744
rect 18269 680 18270 744
rect 18204 664 18270 680
rect 18204 600 18205 664
rect 18269 600 18270 664
rect 18204 584 18270 600
rect 18204 520 18205 584
rect 18269 520 18270 584
rect 18204 504 18270 520
rect 18204 440 18205 504
rect 18269 440 18270 504
rect 18204 350 18270 440
rect 18330 286 18390 1316
rect 18450 346 18510 1378
rect 18570 286 18630 1316
rect 18690 346 18750 1378
rect 18810 1224 18876 1378
rect 18810 1160 18811 1224
rect 18875 1160 18876 1224
rect 18810 1144 18876 1160
rect 18810 1080 18811 1144
rect 18875 1080 18876 1144
rect 18810 1064 18876 1080
rect 18810 1000 18811 1064
rect 18875 1000 18876 1064
rect 18810 984 18876 1000
rect 18810 920 18811 984
rect 18875 920 18876 984
rect 18810 904 18876 920
rect 18810 840 18811 904
rect 18875 840 18876 904
rect 18810 824 18876 840
rect 18810 760 18811 824
rect 18875 760 18876 824
rect 18810 744 18876 760
rect 18810 680 18811 744
rect 18875 680 18876 744
rect 18810 664 18876 680
rect 18810 600 18811 664
rect 18875 600 18876 664
rect 18810 584 18876 600
rect 18810 520 18811 584
rect 18875 520 18876 584
rect 18810 504 18876 520
rect 18810 440 18811 504
rect 18875 440 18876 504
rect 18810 350 18876 440
rect 18936 286 18996 1316
rect 19056 346 19116 1378
rect 19176 286 19236 1316
rect 19296 346 19356 1378
rect 19416 1224 19482 1378
rect 19416 1160 19417 1224
rect 19481 1160 19482 1224
rect 19416 1144 19482 1160
rect 19416 1080 19417 1144
rect 19481 1080 19482 1144
rect 19416 1064 19482 1080
rect 19416 1000 19417 1064
rect 19481 1000 19482 1064
rect 19416 984 19482 1000
rect 19416 920 19417 984
rect 19481 920 19482 984
rect 19416 904 19482 920
rect 19416 840 19417 904
rect 19481 840 19482 904
rect 19416 824 19482 840
rect 19416 760 19417 824
rect 19481 760 19482 824
rect 19416 744 19482 760
rect 19416 680 19417 744
rect 19481 680 19482 744
rect 19416 664 19482 680
rect 19416 600 19417 664
rect 19481 600 19482 664
rect 19416 584 19482 600
rect 19416 520 19417 584
rect 19481 520 19482 584
rect 19416 504 19482 520
rect 19416 440 19417 504
rect 19481 440 19482 504
rect 19416 350 19482 440
rect 19542 286 19602 1316
rect 19662 346 19722 1378
rect 19782 286 19842 1316
rect 19902 346 19962 1378
rect 20022 1224 20088 1378
rect 20022 1160 20023 1224
rect 20087 1160 20088 1224
rect 20022 1144 20088 1160
rect 20022 1080 20023 1144
rect 20087 1080 20088 1144
rect 20022 1064 20088 1080
rect 20022 1000 20023 1064
rect 20087 1000 20088 1064
rect 20022 984 20088 1000
rect 20022 920 20023 984
rect 20087 920 20088 984
rect 20022 904 20088 920
rect 20022 840 20023 904
rect 20087 840 20088 904
rect 20022 824 20088 840
rect 20022 760 20023 824
rect 20087 760 20088 824
rect 20022 744 20088 760
rect 20022 680 20023 744
rect 20087 680 20088 744
rect 20022 664 20088 680
rect 20022 600 20023 664
rect 20087 600 20088 664
rect 20022 584 20088 600
rect 20022 520 20023 584
rect 20087 520 20088 584
rect 20022 504 20088 520
rect 20022 440 20023 504
rect 20087 440 20088 504
rect 20022 350 20088 440
rect 20148 2462 20214 2474
rect 20148 2406 20153 2462
rect 20209 2406 20214 2462
rect 20148 2384 20214 2406
rect 20148 2320 20149 2384
rect 20213 2320 20214 2384
rect 20148 2304 20214 2320
rect 20148 2240 20149 2304
rect 20213 2240 20214 2304
rect 20148 2224 20214 2240
rect 20148 2160 20149 2224
rect 20213 2160 20214 2224
rect 20148 2144 20214 2160
rect 20148 2080 20149 2144
rect 20213 2080 20214 2144
rect 20148 2064 20214 2080
rect 20148 2000 20149 2064
rect 20213 2000 20214 2064
rect 20148 1984 20214 2000
rect 20148 1920 20149 1984
rect 20213 1920 20214 1984
rect 20148 1904 20214 1920
rect 20148 1840 20149 1904
rect 20213 1840 20214 1904
rect 20148 1824 20214 1840
rect 20148 1760 20149 1824
rect 20213 1760 20214 1824
rect 20148 1744 20214 1760
rect 20148 1680 20149 1744
rect 20213 1680 20214 1744
rect 20148 1664 20214 1680
rect 20148 1600 20149 1664
rect 20213 1600 20214 1664
rect 20148 1446 20214 1600
rect 20274 1446 20334 2478
rect 20394 1508 20454 2538
rect 20514 1446 20574 2478
rect 20634 1508 20694 2538
rect 20754 2384 20820 2474
rect 20754 2320 20755 2384
rect 20819 2320 20820 2384
rect 20754 2304 20820 2320
rect 20754 2240 20755 2304
rect 20819 2240 20820 2304
rect 20754 2224 20820 2240
rect 20754 2160 20755 2224
rect 20819 2160 20820 2224
rect 20754 2144 20820 2160
rect 20754 2080 20755 2144
rect 20819 2080 20820 2144
rect 20754 2064 20820 2080
rect 20754 2000 20755 2064
rect 20819 2000 20820 2064
rect 20754 1984 20820 2000
rect 20754 1920 20755 1984
rect 20819 1920 20820 1984
rect 20754 1904 20820 1920
rect 20754 1840 20755 1904
rect 20819 1840 20820 1904
rect 20754 1824 20820 1840
rect 20754 1760 20755 1824
rect 20819 1760 20820 1824
rect 20754 1744 20820 1760
rect 20754 1680 20755 1744
rect 20819 1680 20820 1744
rect 20754 1664 20820 1680
rect 20754 1600 20755 1664
rect 20819 1600 20820 1664
rect 20754 1446 20820 1600
rect 20880 1446 20940 2478
rect 21000 1508 21060 2538
rect 21120 1446 21180 2478
rect 21240 1508 21300 2538
rect 21360 2384 21426 2474
rect 21360 2320 21361 2384
rect 21425 2320 21426 2384
rect 21360 2304 21426 2320
rect 21360 2240 21361 2304
rect 21425 2240 21426 2304
rect 21360 2224 21426 2240
rect 21360 2160 21361 2224
rect 21425 2160 21426 2224
rect 21360 2144 21426 2160
rect 21360 2080 21361 2144
rect 21425 2080 21426 2144
rect 21360 2064 21426 2080
rect 21360 2000 21361 2064
rect 21425 2000 21426 2064
rect 21360 1984 21426 2000
rect 21360 1920 21361 1984
rect 21425 1920 21426 1984
rect 21360 1904 21426 1920
rect 21360 1840 21361 1904
rect 21425 1840 21426 1904
rect 21360 1824 21426 1840
rect 21360 1760 21361 1824
rect 21425 1760 21426 1824
rect 21360 1744 21426 1760
rect 21360 1680 21361 1744
rect 21425 1680 21426 1744
rect 21360 1664 21426 1680
rect 21360 1600 21361 1664
rect 21425 1600 21426 1664
rect 21360 1446 21426 1600
rect 21486 1446 21546 2478
rect 21606 1508 21666 2538
rect 21726 1446 21786 2478
rect 21846 1508 21906 2538
rect 21966 2384 22032 2474
rect 21966 2320 21967 2384
rect 22031 2320 22032 2384
rect 21966 2304 22032 2320
rect 21966 2240 21967 2304
rect 22031 2240 22032 2304
rect 21966 2224 22032 2240
rect 21966 2160 21967 2224
rect 22031 2160 22032 2224
rect 21966 2144 22032 2160
rect 21966 2080 21967 2144
rect 22031 2080 22032 2144
rect 21966 2064 22032 2080
rect 21966 2000 21967 2064
rect 22031 2000 22032 2064
rect 21966 1984 22032 2000
rect 21966 1920 21967 1984
rect 22031 1920 22032 1984
rect 21966 1904 22032 1920
rect 21966 1840 21967 1904
rect 22031 1840 22032 1904
rect 21966 1824 22032 1840
rect 21966 1760 21967 1824
rect 22031 1760 22032 1824
rect 21966 1744 22032 1760
rect 21966 1680 21967 1744
rect 22031 1680 22032 1744
rect 21966 1664 22032 1680
rect 21966 1600 21967 1664
rect 22031 1600 22032 1664
rect 21966 1446 22032 1600
rect 22092 1446 22152 2478
rect 22212 1508 22272 2538
rect 22332 1446 22392 2478
rect 22452 1508 22512 2538
rect 22572 2384 22638 2474
rect 22572 2320 22573 2384
rect 22637 2320 22638 2384
rect 22572 2304 22638 2320
rect 22572 2240 22573 2304
rect 22637 2240 22638 2304
rect 22572 2224 22638 2240
rect 22572 2160 22573 2224
rect 22637 2160 22638 2224
rect 22572 2144 22638 2160
rect 22572 2080 22573 2144
rect 22637 2080 22638 2144
rect 22572 2064 22638 2080
rect 22572 2000 22573 2064
rect 22637 2000 22638 2064
rect 22572 1984 22638 2000
rect 22572 1920 22573 1984
rect 22637 1920 22638 1984
rect 22572 1904 22638 1920
rect 22572 1840 22573 1904
rect 22637 1840 22638 1904
rect 22572 1824 22638 1840
rect 22572 1760 22573 1824
rect 22637 1760 22638 1824
rect 22572 1744 22638 1760
rect 22572 1680 22573 1744
rect 22637 1680 22638 1744
rect 22572 1664 22638 1680
rect 22572 1600 22573 1664
rect 22637 1600 22638 1664
rect 22572 1446 22638 1600
rect 22698 1446 22758 2478
rect 22818 1508 22878 2538
rect 22938 1446 22998 2478
rect 23058 1508 23118 2538
rect 23178 2384 23244 2474
rect 23178 2320 23179 2384
rect 23243 2320 23244 2384
rect 23178 2304 23244 2320
rect 23178 2240 23179 2304
rect 23243 2240 23244 2304
rect 23178 2224 23244 2240
rect 23178 2160 23179 2224
rect 23243 2160 23244 2224
rect 23178 2144 23244 2160
rect 23178 2080 23179 2144
rect 23243 2080 23244 2144
rect 23178 2064 23244 2080
rect 23178 2000 23179 2064
rect 23243 2000 23244 2064
rect 23178 1984 23244 2000
rect 23178 1920 23179 1984
rect 23243 1920 23244 1984
rect 23178 1904 23244 1920
rect 23178 1840 23179 1904
rect 23243 1840 23244 1904
rect 23178 1824 23244 1840
rect 23178 1760 23179 1824
rect 23243 1760 23244 1824
rect 23178 1744 23244 1760
rect 23178 1680 23179 1744
rect 23243 1680 23244 1744
rect 23178 1664 23244 1680
rect 23178 1600 23179 1664
rect 23243 1600 23244 1664
rect 23178 1446 23244 1600
rect 23304 1446 23364 2478
rect 23424 1508 23484 2538
rect 23544 1446 23604 2478
rect 23664 1508 23724 2538
rect 23784 2384 23850 2474
rect 23784 2320 23785 2384
rect 23849 2320 23850 2384
rect 23784 2304 23850 2320
rect 23784 2240 23785 2304
rect 23849 2240 23850 2304
rect 23784 2224 23850 2240
rect 23784 2160 23785 2224
rect 23849 2160 23850 2224
rect 23784 2144 23850 2160
rect 23784 2080 23785 2144
rect 23849 2080 23850 2144
rect 23784 2064 23850 2080
rect 23784 2000 23785 2064
rect 23849 2000 23850 2064
rect 23784 1984 23850 2000
rect 23784 1920 23785 1984
rect 23849 1920 23850 1984
rect 23784 1904 23850 1920
rect 23784 1840 23785 1904
rect 23849 1840 23850 1904
rect 23784 1824 23850 1840
rect 23784 1760 23785 1824
rect 23849 1760 23850 1824
rect 23784 1744 23850 1760
rect 23784 1680 23785 1744
rect 23849 1680 23850 1744
rect 23784 1664 23850 1680
rect 23784 1600 23785 1664
rect 23849 1600 23850 1664
rect 23784 1446 23850 1600
rect 23910 1446 23970 2478
rect 24030 1508 24090 2538
rect 24150 1446 24210 2478
rect 24270 1508 24330 2538
rect 24390 2384 24456 2474
rect 24390 2320 24391 2384
rect 24455 2320 24456 2384
rect 24390 2304 24456 2320
rect 24390 2240 24391 2304
rect 24455 2240 24456 2304
rect 24390 2224 24456 2240
rect 24390 2160 24391 2224
rect 24455 2160 24456 2224
rect 24390 2144 24456 2160
rect 24390 2080 24391 2144
rect 24455 2080 24456 2144
rect 24390 2064 24456 2080
rect 24390 2000 24391 2064
rect 24455 2000 24456 2064
rect 24390 1984 24456 2000
rect 24390 1920 24391 1984
rect 24455 1920 24456 1984
rect 24390 1904 24456 1920
rect 24390 1840 24391 1904
rect 24455 1840 24456 1904
rect 24390 1824 24456 1840
rect 24390 1760 24391 1824
rect 24455 1760 24456 1824
rect 24390 1744 24456 1760
rect 24390 1680 24391 1744
rect 24455 1680 24456 1744
rect 24390 1664 24456 1680
rect 24390 1600 24391 1664
rect 24455 1600 24456 1664
rect 24390 1446 24456 1600
rect 24516 1446 24576 2478
rect 24636 1508 24696 2538
rect 24756 1446 24816 2478
rect 24876 1508 24936 2538
rect 24996 2384 25062 2474
rect 24996 2320 24997 2384
rect 25061 2320 25062 2384
rect 24996 2304 25062 2320
rect 24996 2240 24997 2304
rect 25061 2240 25062 2304
rect 24996 2224 25062 2240
rect 24996 2160 24997 2224
rect 25061 2160 25062 2224
rect 24996 2144 25062 2160
rect 24996 2080 24997 2144
rect 25061 2080 25062 2144
rect 24996 2064 25062 2080
rect 24996 2000 24997 2064
rect 25061 2000 25062 2064
rect 24996 1984 25062 2000
rect 24996 1920 24997 1984
rect 25061 1920 25062 1984
rect 24996 1904 25062 1920
rect 24996 1840 24997 1904
rect 25061 1840 25062 1904
rect 24996 1824 25062 1840
rect 24996 1760 24997 1824
rect 25061 1760 25062 1824
rect 24996 1744 25062 1760
rect 24996 1680 24997 1744
rect 25061 1680 25062 1744
rect 24996 1664 25062 1680
rect 24996 1600 24997 1664
rect 25061 1600 25062 1664
rect 24996 1446 25062 1600
rect 25122 1446 25182 2478
rect 25242 1508 25302 2538
rect 25362 1446 25422 2478
rect 25482 1508 25542 2538
rect 25602 2384 25668 2474
rect 25602 2320 25603 2384
rect 25667 2320 25668 2384
rect 25602 2304 25668 2320
rect 25602 2240 25603 2304
rect 25667 2240 25668 2304
rect 25602 2224 25668 2240
rect 25602 2160 25603 2224
rect 25667 2160 25668 2224
rect 25602 2144 25668 2160
rect 25602 2080 25603 2144
rect 25667 2080 25668 2144
rect 25602 2064 25668 2080
rect 25602 2000 25603 2064
rect 25667 2000 25668 2064
rect 25602 1984 25668 2000
rect 25602 1920 25603 1984
rect 25667 1920 25668 1984
rect 25602 1904 25668 1920
rect 25602 1840 25603 1904
rect 25667 1840 25668 1904
rect 25602 1824 25668 1840
rect 25602 1760 25603 1824
rect 25667 1760 25668 1824
rect 25602 1744 25668 1760
rect 25602 1680 25603 1744
rect 25667 1680 25668 1744
rect 25602 1664 25668 1680
rect 25602 1600 25603 1664
rect 25667 1600 25668 1664
rect 25602 1446 25668 1600
rect 25728 1446 25788 2478
rect 25848 1508 25908 2538
rect 25968 1446 26028 2478
rect 26088 1508 26148 2538
rect 26208 2384 26274 2474
rect 26208 2320 26209 2384
rect 26273 2320 26274 2384
rect 26208 2304 26274 2320
rect 26208 2240 26209 2304
rect 26273 2240 26274 2304
rect 26208 2224 26274 2240
rect 26208 2160 26209 2224
rect 26273 2160 26274 2224
rect 26208 2144 26274 2160
rect 26208 2080 26209 2144
rect 26273 2080 26274 2144
rect 26208 2064 26274 2080
rect 26208 2000 26209 2064
rect 26273 2000 26274 2064
rect 26208 1984 26274 2000
rect 26208 1920 26209 1984
rect 26273 1920 26274 1984
rect 26208 1904 26274 1920
rect 26208 1840 26209 1904
rect 26273 1840 26274 1904
rect 26208 1824 26274 1840
rect 26208 1760 26209 1824
rect 26273 1760 26274 1824
rect 26208 1744 26274 1760
rect 26208 1680 26209 1744
rect 26273 1680 26274 1744
rect 26208 1664 26274 1680
rect 26208 1600 26209 1664
rect 26273 1600 26274 1664
rect 26208 1446 26274 1600
rect 26334 1446 26394 2478
rect 26454 1508 26514 2538
rect 26574 1446 26634 2478
rect 26694 1508 26754 2538
rect 26814 2384 26880 2474
rect 26814 2320 26815 2384
rect 26879 2320 26880 2384
rect 26814 2304 26880 2320
rect 26814 2240 26815 2304
rect 26879 2240 26880 2304
rect 26814 2224 26880 2240
rect 26814 2160 26815 2224
rect 26879 2160 26880 2224
rect 26814 2144 26880 2160
rect 26814 2080 26815 2144
rect 26879 2080 26880 2144
rect 26814 2064 26880 2080
rect 26814 2000 26815 2064
rect 26879 2000 26880 2064
rect 26814 1984 26880 2000
rect 26814 1920 26815 1984
rect 26879 1920 26880 1984
rect 26814 1904 26880 1920
rect 26814 1840 26815 1904
rect 26879 1840 26880 1904
rect 26814 1824 26880 1840
rect 26814 1760 26815 1824
rect 26879 1760 26880 1824
rect 26814 1744 26880 1760
rect 26814 1680 26815 1744
rect 26879 1680 26880 1744
rect 26814 1664 26880 1680
rect 26814 1600 26815 1664
rect 26879 1600 26880 1664
rect 26814 1446 26880 1600
rect 26940 1446 27000 2478
rect 27060 1508 27120 2538
rect 27180 1446 27240 2478
rect 27300 1508 27360 2538
rect 27420 2384 27486 2474
rect 27420 2320 27421 2384
rect 27485 2320 27486 2384
rect 27420 2304 27486 2320
rect 27420 2240 27421 2304
rect 27485 2240 27486 2304
rect 27420 2224 27486 2240
rect 27420 2160 27421 2224
rect 27485 2160 27486 2224
rect 27420 2144 27486 2160
rect 27420 2080 27421 2144
rect 27485 2080 27486 2144
rect 27420 2064 27486 2080
rect 27420 2000 27421 2064
rect 27485 2000 27486 2064
rect 27420 1984 27486 2000
rect 27420 1920 27421 1984
rect 27485 1920 27486 1984
rect 27420 1904 27486 1920
rect 27420 1840 27421 1904
rect 27485 1840 27486 1904
rect 27420 1824 27486 1840
rect 27420 1760 27421 1824
rect 27485 1760 27486 1824
rect 27420 1744 27486 1760
rect 27420 1680 27421 1744
rect 27485 1680 27486 1744
rect 27420 1664 27486 1680
rect 27420 1600 27421 1664
rect 27485 1600 27486 1664
rect 27420 1446 27486 1600
rect 27546 1446 27606 2478
rect 27666 1508 27726 2538
rect 27786 1446 27846 2478
rect 27906 1508 27966 2538
rect 28026 2384 28092 2474
rect 28026 2320 28027 2384
rect 28091 2320 28092 2384
rect 28026 2304 28092 2320
rect 28026 2240 28027 2304
rect 28091 2240 28092 2304
rect 28026 2224 28092 2240
rect 28026 2160 28027 2224
rect 28091 2160 28092 2224
rect 28026 2144 28092 2160
rect 28026 2080 28027 2144
rect 28091 2080 28092 2144
rect 28026 2064 28092 2080
rect 28026 2000 28027 2064
rect 28091 2000 28092 2064
rect 28026 1984 28092 2000
rect 28026 1920 28027 1984
rect 28091 1920 28092 1984
rect 28026 1904 28092 1920
rect 28026 1840 28027 1904
rect 28091 1840 28092 1904
rect 28026 1824 28092 1840
rect 28026 1760 28027 1824
rect 28091 1760 28092 1824
rect 28026 1744 28092 1760
rect 28026 1680 28027 1744
rect 28091 1680 28092 1744
rect 28026 1664 28092 1680
rect 28026 1600 28027 1664
rect 28091 1600 28092 1664
rect 28026 1446 28092 1600
rect 28152 1446 28212 2478
rect 28272 1508 28332 2538
rect 28392 1446 28452 2478
rect 28512 1508 28572 2538
rect 28632 2384 28698 2474
rect 28632 2320 28633 2384
rect 28697 2320 28698 2384
rect 28632 2304 28698 2320
rect 28632 2240 28633 2304
rect 28697 2240 28698 2304
rect 28632 2224 28698 2240
rect 28632 2160 28633 2224
rect 28697 2160 28698 2224
rect 28632 2144 28698 2160
rect 28632 2080 28633 2144
rect 28697 2080 28698 2144
rect 28632 2064 28698 2080
rect 28632 2000 28633 2064
rect 28697 2000 28698 2064
rect 28632 1984 28698 2000
rect 28632 1920 28633 1984
rect 28697 1920 28698 1984
rect 28632 1904 28698 1920
rect 28632 1840 28633 1904
rect 28697 1840 28698 1904
rect 28632 1824 28698 1840
rect 28632 1760 28633 1824
rect 28697 1760 28698 1824
rect 28632 1744 28698 1760
rect 28632 1680 28633 1744
rect 28697 1680 28698 1744
rect 28632 1664 28698 1680
rect 28632 1600 28633 1664
rect 28697 1600 28698 1664
rect 28632 1446 28698 1600
rect 28758 1446 28818 2478
rect 28878 1508 28938 2538
rect 28998 1446 29058 2478
rect 29118 1508 29178 2538
rect 29238 2384 29304 2474
rect 29238 2320 29239 2384
rect 29303 2320 29304 2384
rect 29238 2304 29304 2320
rect 29238 2240 29239 2304
rect 29303 2240 29304 2304
rect 29238 2224 29304 2240
rect 29238 2160 29239 2224
rect 29303 2160 29304 2224
rect 29238 2144 29304 2160
rect 29238 2080 29239 2144
rect 29303 2080 29304 2144
rect 29238 2064 29304 2080
rect 29238 2000 29239 2064
rect 29303 2000 29304 2064
rect 29238 1984 29304 2000
rect 29238 1920 29239 1984
rect 29303 1920 29304 1984
rect 29238 1904 29304 1920
rect 29238 1840 29239 1904
rect 29303 1840 29304 1904
rect 29238 1824 29304 1840
rect 29238 1760 29239 1824
rect 29303 1760 29304 1824
rect 29238 1744 29304 1760
rect 29238 1680 29239 1744
rect 29303 1680 29304 1744
rect 29238 1664 29304 1680
rect 29238 1600 29239 1664
rect 29303 1600 29304 1664
rect 29238 1446 29304 1600
rect 29364 1446 29424 2478
rect 29484 1508 29544 2538
rect 29604 1446 29664 2478
rect 29724 1508 29784 2538
rect 29844 2384 29910 2474
rect 29844 2320 29845 2384
rect 29909 2320 29910 2384
rect 29844 2304 29910 2320
rect 29844 2240 29845 2304
rect 29909 2240 29910 2304
rect 29844 2224 29910 2240
rect 29844 2160 29845 2224
rect 29909 2160 29910 2224
rect 29844 2144 29910 2160
rect 29844 2080 29845 2144
rect 29909 2080 29910 2144
rect 29844 2064 29910 2080
rect 29844 2000 29845 2064
rect 29909 2000 29910 2064
rect 29844 1984 29910 2000
rect 29844 1920 29845 1984
rect 29909 1920 29910 1984
rect 29844 1904 29910 1920
rect 29844 1840 29845 1904
rect 29909 1840 29910 1904
rect 29844 1824 29910 1840
rect 29844 1760 29845 1824
rect 29909 1760 29910 1824
rect 29844 1744 29910 1760
rect 29844 1680 29845 1744
rect 29909 1680 29910 1744
rect 29844 1664 29910 1680
rect 29844 1600 29845 1664
rect 29909 1600 29910 1664
rect 29844 1446 29910 1600
rect 29970 1446 30030 2478
rect 30090 1508 30150 2538
rect 30210 1446 30270 2478
rect 30330 1508 30390 2538
rect 30450 2384 30516 2474
rect 30450 2320 30451 2384
rect 30515 2320 30516 2384
rect 30450 2304 30516 2320
rect 30450 2240 30451 2304
rect 30515 2240 30516 2304
rect 30450 2224 30516 2240
rect 30450 2160 30451 2224
rect 30515 2160 30516 2224
rect 30450 2144 30516 2160
rect 30450 2080 30451 2144
rect 30515 2080 30516 2144
rect 30450 2064 30516 2080
rect 30450 2000 30451 2064
rect 30515 2000 30516 2064
rect 30450 1984 30516 2000
rect 30450 1920 30451 1984
rect 30515 1920 30516 1984
rect 30450 1904 30516 1920
rect 30450 1840 30451 1904
rect 30515 1840 30516 1904
rect 30450 1824 30516 1840
rect 30450 1760 30451 1824
rect 30515 1760 30516 1824
rect 30450 1744 30516 1760
rect 30450 1680 30451 1744
rect 30515 1680 30516 1744
rect 30450 1664 30516 1680
rect 30450 1600 30451 1664
rect 30515 1600 30516 1664
rect 30450 1446 30516 1600
rect 30576 1446 30636 2478
rect 30696 1508 30756 2538
rect 30816 1446 30876 2478
rect 30936 1508 30996 2538
rect 31056 2384 31122 2474
rect 31056 2320 31057 2384
rect 31121 2320 31122 2384
rect 31056 2304 31122 2320
rect 31056 2240 31057 2304
rect 31121 2240 31122 2304
rect 31056 2224 31122 2240
rect 31056 2160 31057 2224
rect 31121 2160 31122 2224
rect 31056 2144 31122 2160
rect 31056 2080 31057 2144
rect 31121 2080 31122 2144
rect 31056 2064 31122 2080
rect 31056 2000 31057 2064
rect 31121 2000 31122 2064
rect 31056 1984 31122 2000
rect 31056 1920 31057 1984
rect 31121 1920 31122 1984
rect 31056 1904 31122 1920
rect 31056 1840 31057 1904
rect 31121 1840 31122 1904
rect 31056 1824 31122 1840
rect 31056 1760 31057 1824
rect 31121 1760 31122 1824
rect 31056 1744 31122 1760
rect 31056 1680 31057 1744
rect 31121 1680 31122 1744
rect 31056 1664 31122 1680
rect 31056 1600 31057 1664
rect 31121 1600 31122 1664
rect 31056 1446 31122 1600
rect 31182 1446 31242 2478
rect 31302 1508 31362 2538
rect 31422 1446 31482 2478
rect 31542 1508 31602 2538
rect 31662 2384 31728 2474
rect 31662 2320 31663 2384
rect 31727 2320 31728 2384
rect 31662 2304 31728 2320
rect 31662 2240 31663 2304
rect 31727 2240 31728 2304
rect 31662 2224 31728 2240
rect 31662 2160 31663 2224
rect 31727 2160 31728 2224
rect 31662 2144 31728 2160
rect 31662 2080 31663 2144
rect 31727 2080 31728 2144
rect 31662 2064 31728 2080
rect 31662 2000 31663 2064
rect 31727 2000 31728 2064
rect 31662 1984 31728 2000
rect 31662 1920 31663 1984
rect 31727 1920 31728 1984
rect 31662 1904 31728 1920
rect 31662 1840 31663 1904
rect 31727 1840 31728 1904
rect 31662 1824 31728 1840
rect 31662 1760 31663 1824
rect 31727 1760 31728 1824
rect 31662 1744 31728 1760
rect 31662 1680 31663 1744
rect 31727 1680 31728 1744
rect 31662 1664 31728 1680
rect 31662 1600 31663 1664
rect 31727 1600 31728 1664
rect 31662 1446 31728 1600
rect 31788 1446 31848 2478
rect 31908 1508 31968 2538
rect 32028 1446 32088 2478
rect 32148 1508 32208 2538
rect 32268 2384 32334 2474
rect 32268 2320 32269 2384
rect 32333 2320 32334 2384
rect 32268 2304 32334 2320
rect 32268 2240 32269 2304
rect 32333 2240 32334 2304
rect 32268 2224 32334 2240
rect 32268 2160 32269 2224
rect 32333 2160 32334 2224
rect 32268 2144 32334 2160
rect 32268 2080 32269 2144
rect 32333 2080 32334 2144
rect 32268 2064 32334 2080
rect 32268 2000 32269 2064
rect 32333 2000 32334 2064
rect 32268 1984 32334 2000
rect 32268 1920 32269 1984
rect 32333 1920 32334 1984
rect 32268 1904 32334 1920
rect 32268 1840 32269 1904
rect 32333 1840 32334 1904
rect 32268 1824 32334 1840
rect 32268 1760 32269 1824
rect 32333 1760 32334 1824
rect 32268 1744 32334 1760
rect 32268 1680 32269 1744
rect 32333 1680 32334 1744
rect 32268 1664 32334 1680
rect 32268 1600 32269 1664
rect 32333 1600 32334 1664
rect 32268 1446 32334 1600
rect 32394 1446 32454 2478
rect 32514 1508 32574 2538
rect 32634 1446 32694 2478
rect 32754 1508 32814 2538
rect 32874 2384 32940 2474
rect 32874 2320 32875 2384
rect 32939 2320 32940 2384
rect 32874 2304 32940 2320
rect 32874 2240 32875 2304
rect 32939 2240 32940 2304
rect 32874 2224 32940 2240
rect 32874 2160 32875 2224
rect 32939 2160 32940 2224
rect 32874 2144 32940 2160
rect 32874 2080 32875 2144
rect 32939 2080 32940 2144
rect 32874 2064 32940 2080
rect 32874 2000 32875 2064
rect 32939 2000 32940 2064
rect 32874 1984 32940 2000
rect 32874 1920 32875 1984
rect 32939 1920 32940 1984
rect 32874 1904 32940 1920
rect 32874 1840 32875 1904
rect 32939 1840 32940 1904
rect 32874 1824 32940 1840
rect 32874 1760 32875 1824
rect 32939 1760 32940 1824
rect 32874 1744 32940 1760
rect 32874 1680 32875 1744
rect 32939 1680 32940 1744
rect 32874 1664 32940 1680
rect 32874 1600 32875 1664
rect 32939 1600 32940 1664
rect 32874 1446 32940 1600
rect 33000 1446 33060 2478
rect 33120 1508 33180 2538
rect 33240 1446 33300 2478
rect 33360 1508 33420 2538
rect 33480 2384 33546 2474
rect 33480 2320 33481 2384
rect 33545 2320 33546 2384
rect 33480 2304 33546 2320
rect 33480 2240 33481 2304
rect 33545 2240 33546 2304
rect 33480 2224 33546 2240
rect 33480 2160 33481 2224
rect 33545 2160 33546 2224
rect 33480 2144 33546 2160
rect 33480 2080 33481 2144
rect 33545 2080 33546 2144
rect 33480 2064 33546 2080
rect 33480 2000 33481 2064
rect 33545 2000 33546 2064
rect 33480 1984 33546 2000
rect 33480 1920 33481 1984
rect 33545 1920 33546 1984
rect 33480 1904 33546 1920
rect 33480 1840 33481 1904
rect 33545 1840 33546 1904
rect 33480 1824 33546 1840
rect 33480 1760 33481 1824
rect 33545 1760 33546 1824
rect 33480 1744 33546 1760
rect 33480 1680 33481 1744
rect 33545 1680 33546 1744
rect 33480 1664 33546 1680
rect 33480 1600 33481 1664
rect 33545 1600 33546 1664
rect 33480 1446 33546 1600
rect 33606 1446 33666 2478
rect 33726 1508 33786 2538
rect 33846 1446 33906 2478
rect 33966 1508 34026 2538
rect 34086 2384 34152 2474
rect 34086 2320 34087 2384
rect 34151 2320 34152 2384
rect 34086 2304 34152 2320
rect 34086 2240 34087 2304
rect 34151 2240 34152 2304
rect 34086 2224 34152 2240
rect 34086 2160 34087 2224
rect 34151 2160 34152 2224
rect 34086 2144 34152 2160
rect 34086 2080 34087 2144
rect 34151 2080 34152 2144
rect 34086 2064 34152 2080
rect 34086 2000 34087 2064
rect 34151 2000 34152 2064
rect 34086 1984 34152 2000
rect 34086 1920 34087 1984
rect 34151 1920 34152 1984
rect 34086 1904 34152 1920
rect 34086 1840 34087 1904
rect 34151 1840 34152 1904
rect 34086 1824 34152 1840
rect 34086 1760 34087 1824
rect 34151 1760 34152 1824
rect 34086 1744 34152 1760
rect 34086 1680 34087 1744
rect 34151 1680 34152 1744
rect 34086 1664 34152 1680
rect 34086 1600 34087 1664
rect 34151 1600 34152 1664
rect 34086 1446 34152 1600
rect 34212 1446 34272 2478
rect 34332 1508 34392 2538
rect 34452 1446 34512 2478
rect 34572 1508 34632 2538
rect 34692 2384 34758 2474
rect 34692 2320 34693 2384
rect 34757 2320 34758 2384
rect 34692 2304 34758 2320
rect 34692 2240 34693 2304
rect 34757 2240 34758 2304
rect 34692 2224 34758 2240
rect 34692 2160 34693 2224
rect 34757 2160 34758 2224
rect 34692 2144 34758 2160
rect 34692 2080 34693 2144
rect 34757 2080 34758 2144
rect 34692 2064 34758 2080
rect 34692 2000 34693 2064
rect 34757 2000 34758 2064
rect 34692 1984 34758 2000
rect 34692 1920 34693 1984
rect 34757 1920 34758 1984
rect 34692 1904 34758 1920
rect 34692 1840 34693 1904
rect 34757 1840 34758 1904
rect 34692 1824 34758 1840
rect 34692 1760 34693 1824
rect 34757 1760 34758 1824
rect 34692 1744 34758 1760
rect 34692 1680 34693 1744
rect 34757 1680 34758 1744
rect 34692 1664 34758 1680
rect 34692 1600 34693 1664
rect 34757 1600 34758 1664
rect 34692 1446 34758 1600
rect 34818 1446 34878 2478
rect 34938 1508 34998 2538
rect 35058 1446 35118 2478
rect 35178 1508 35238 2538
rect 35298 2384 35364 2474
rect 35298 2320 35299 2384
rect 35363 2320 35364 2384
rect 35298 2304 35364 2320
rect 35298 2240 35299 2304
rect 35363 2240 35364 2304
rect 35298 2224 35364 2240
rect 35298 2160 35299 2224
rect 35363 2160 35364 2224
rect 35298 2144 35364 2160
rect 35298 2080 35299 2144
rect 35363 2080 35364 2144
rect 35298 2064 35364 2080
rect 35298 2000 35299 2064
rect 35363 2000 35364 2064
rect 35298 1984 35364 2000
rect 35298 1920 35299 1984
rect 35363 1920 35364 1984
rect 35298 1904 35364 1920
rect 35298 1840 35299 1904
rect 35363 1840 35364 1904
rect 35298 1824 35364 1840
rect 35298 1760 35299 1824
rect 35363 1760 35364 1824
rect 35298 1744 35364 1760
rect 35298 1680 35299 1744
rect 35363 1680 35364 1744
rect 35298 1664 35364 1680
rect 35298 1600 35299 1664
rect 35363 1600 35364 1664
rect 35298 1446 35364 1600
rect 35424 1446 35484 2478
rect 35544 1508 35604 2538
rect 35664 1446 35724 2478
rect 35784 1508 35844 2538
rect 35904 2384 35970 2474
rect 35904 2320 35905 2384
rect 35969 2320 35970 2384
rect 35904 2304 35970 2320
rect 35904 2240 35905 2304
rect 35969 2240 35970 2304
rect 35904 2224 35970 2240
rect 35904 2160 35905 2224
rect 35969 2160 35970 2224
rect 35904 2144 35970 2160
rect 35904 2080 35905 2144
rect 35969 2080 35970 2144
rect 35904 2064 35970 2080
rect 35904 2000 35905 2064
rect 35969 2000 35970 2064
rect 35904 1984 35970 2000
rect 35904 1920 35905 1984
rect 35969 1920 35970 1984
rect 35904 1904 35970 1920
rect 35904 1840 35905 1904
rect 35969 1840 35970 1904
rect 35904 1824 35970 1840
rect 35904 1760 35905 1824
rect 35969 1760 35970 1824
rect 35904 1744 35970 1760
rect 35904 1680 35905 1744
rect 35969 1680 35970 1744
rect 35904 1664 35970 1680
rect 35904 1600 35905 1664
rect 35969 1600 35970 1664
rect 35904 1446 35970 1600
rect 36030 1446 36090 2478
rect 36150 1508 36210 2538
rect 36270 1446 36330 2478
rect 36390 1508 36450 2538
rect 36510 2384 36576 2474
rect 36510 2320 36511 2384
rect 36575 2320 36576 2384
rect 36510 2304 36576 2320
rect 36510 2240 36511 2304
rect 36575 2240 36576 2304
rect 36510 2224 36576 2240
rect 36510 2160 36511 2224
rect 36575 2160 36576 2224
rect 36510 2144 36576 2160
rect 36510 2080 36511 2144
rect 36575 2080 36576 2144
rect 36510 2064 36576 2080
rect 36510 2000 36511 2064
rect 36575 2000 36576 2064
rect 36510 1984 36576 2000
rect 36510 1920 36511 1984
rect 36575 1920 36576 1984
rect 36510 1904 36576 1920
rect 36510 1840 36511 1904
rect 36575 1840 36576 1904
rect 36510 1824 36576 1840
rect 36510 1760 36511 1824
rect 36575 1760 36576 1824
rect 36510 1744 36576 1760
rect 36510 1680 36511 1744
rect 36575 1680 36576 1744
rect 36510 1664 36576 1680
rect 36510 1600 36511 1664
rect 36575 1600 36576 1664
rect 36510 1446 36576 1600
rect 36636 1446 36696 2478
rect 36756 1508 36816 2538
rect 36876 1446 36936 2478
rect 36996 1508 37056 2538
rect 37116 2384 37182 2474
rect 37116 2320 37117 2384
rect 37181 2320 37182 2384
rect 37116 2304 37182 2320
rect 37116 2240 37117 2304
rect 37181 2240 37182 2304
rect 37116 2224 37182 2240
rect 37116 2160 37117 2224
rect 37181 2160 37182 2224
rect 37116 2144 37182 2160
rect 37116 2080 37117 2144
rect 37181 2080 37182 2144
rect 37116 2064 37182 2080
rect 37116 2000 37117 2064
rect 37181 2000 37182 2064
rect 37116 1984 37182 2000
rect 37116 1920 37117 1984
rect 37181 1920 37182 1984
rect 37116 1904 37182 1920
rect 37116 1840 37117 1904
rect 37181 1840 37182 1904
rect 37116 1824 37182 1840
rect 37116 1760 37117 1824
rect 37181 1760 37182 1824
rect 37116 1744 37182 1760
rect 37116 1680 37117 1744
rect 37181 1680 37182 1744
rect 37116 1664 37182 1680
rect 37116 1600 37117 1664
rect 37181 1600 37182 1664
rect 37116 1446 37182 1600
rect 37242 1446 37302 2478
rect 37362 1508 37422 2538
rect 37482 1446 37542 2478
rect 37602 1508 37662 2538
rect 37722 2384 37788 2474
rect 37722 2320 37723 2384
rect 37787 2320 37788 2384
rect 37722 2304 37788 2320
rect 37722 2240 37723 2304
rect 37787 2240 37788 2304
rect 37722 2224 37788 2240
rect 37722 2160 37723 2224
rect 37787 2160 37788 2224
rect 37722 2144 37788 2160
rect 37722 2080 37723 2144
rect 37787 2080 37788 2144
rect 37722 2064 37788 2080
rect 37722 2000 37723 2064
rect 37787 2000 37788 2064
rect 37722 1984 37788 2000
rect 37722 1920 37723 1984
rect 37787 1920 37788 1984
rect 37722 1904 37788 1920
rect 37722 1840 37723 1904
rect 37787 1840 37788 1904
rect 37722 1824 37788 1840
rect 37722 1760 37723 1824
rect 37787 1760 37788 1824
rect 37722 1744 37788 1760
rect 37722 1680 37723 1744
rect 37787 1680 37788 1744
rect 37722 1664 37788 1680
rect 37722 1600 37723 1664
rect 37787 1600 37788 1664
rect 37722 1446 37788 1600
rect 37848 1446 37908 2478
rect 37968 1508 38028 2538
rect 38088 1446 38148 2478
rect 38208 1508 38268 2538
rect 38328 2384 38394 2474
rect 38328 2320 38329 2384
rect 38393 2320 38394 2384
rect 38328 2304 38394 2320
rect 38328 2240 38329 2304
rect 38393 2240 38394 2304
rect 38328 2224 38394 2240
rect 38328 2160 38329 2224
rect 38393 2160 38394 2224
rect 38328 2144 38394 2160
rect 38328 2080 38329 2144
rect 38393 2080 38394 2144
rect 38328 2064 38394 2080
rect 38328 2000 38329 2064
rect 38393 2000 38394 2064
rect 38328 1984 38394 2000
rect 38328 1920 38329 1984
rect 38393 1920 38394 1984
rect 38328 1904 38394 1920
rect 38328 1840 38329 1904
rect 38393 1840 38394 1904
rect 38328 1824 38394 1840
rect 38328 1760 38329 1824
rect 38393 1760 38394 1824
rect 38328 1744 38394 1760
rect 38328 1680 38329 1744
rect 38393 1680 38394 1744
rect 38328 1664 38394 1680
rect 38328 1600 38329 1664
rect 38393 1600 38394 1664
rect 38328 1446 38394 1600
rect 38454 1446 38514 2478
rect 38574 1508 38634 2538
rect 38694 1446 38754 2478
rect 38814 1508 38874 2538
rect 38934 2384 39000 2474
rect 38934 2320 38935 2384
rect 38999 2320 39000 2384
rect 38934 2304 39000 2320
rect 38934 2240 38935 2304
rect 38999 2240 39000 2304
rect 38934 2224 39000 2240
rect 38934 2160 38935 2224
rect 38999 2160 39000 2224
rect 38934 2144 39000 2160
rect 38934 2080 38935 2144
rect 38999 2080 39000 2144
rect 38934 2064 39000 2080
rect 38934 2000 38935 2064
rect 38999 2000 39000 2064
rect 38934 1984 39000 2000
rect 38934 1920 38935 1984
rect 38999 1920 39000 1984
rect 38934 1904 39000 1920
rect 38934 1840 38935 1904
rect 38999 1840 39000 1904
rect 38934 1824 39000 1840
rect 38934 1760 38935 1824
rect 38999 1760 39000 1824
rect 38934 1744 39000 1760
rect 38934 1680 38935 1744
rect 38999 1680 39000 1744
rect 38934 1664 39000 1680
rect 38934 1600 38935 1664
rect 38999 1600 39000 1664
rect 38934 1446 39000 1600
rect 39060 1446 39120 2478
rect 39180 1508 39240 2538
rect 39300 1446 39360 2478
rect 39420 1508 39480 2538
rect 39540 2384 39606 2474
rect 39540 2320 39541 2384
rect 39605 2320 39606 2384
rect 39540 2304 39606 2320
rect 39540 2240 39541 2304
rect 39605 2240 39606 2304
rect 39540 2224 39606 2240
rect 39540 2160 39541 2224
rect 39605 2160 39606 2224
rect 39540 2144 39606 2160
rect 39540 2080 39541 2144
rect 39605 2080 39606 2144
rect 39540 2064 39606 2080
rect 39540 2000 39541 2064
rect 39605 2000 39606 2064
rect 39540 1984 39606 2000
rect 39540 1920 39541 1984
rect 39605 1920 39606 1984
rect 39540 1904 39606 1920
rect 39540 1840 39541 1904
rect 39605 1840 39606 1904
rect 39540 1824 39606 1840
rect 39540 1760 39541 1824
rect 39605 1760 39606 1824
rect 39540 1744 39606 1760
rect 39540 1680 39541 1744
rect 39605 1680 39606 1744
rect 39540 1664 39606 1680
rect 39540 1600 39541 1664
rect 39605 1600 39606 1664
rect 39540 1446 39606 1600
rect 20148 1444 39606 1446
rect 20148 1380 20252 1444
rect 20316 1380 20332 1444
rect 20396 1380 20412 1444
rect 20476 1380 20492 1444
rect 20556 1380 20572 1444
rect 20636 1380 20652 1444
rect 20716 1380 20858 1444
rect 20922 1380 20938 1444
rect 21002 1380 21018 1444
rect 21082 1380 21098 1444
rect 21162 1380 21178 1444
rect 21242 1380 21258 1444
rect 21322 1380 21464 1444
rect 21528 1380 21544 1444
rect 21608 1380 21624 1444
rect 21688 1380 21704 1444
rect 21768 1380 21784 1444
rect 21848 1380 21864 1444
rect 21928 1380 22070 1444
rect 22134 1380 22150 1444
rect 22214 1380 22230 1444
rect 22294 1380 22310 1444
rect 22374 1380 22390 1444
rect 22454 1380 22470 1444
rect 22534 1380 22676 1444
rect 22740 1380 22756 1444
rect 22820 1380 22836 1444
rect 22900 1380 22916 1444
rect 22980 1380 22996 1444
rect 23060 1380 23076 1444
rect 23140 1380 23282 1444
rect 23346 1380 23362 1444
rect 23426 1380 23442 1444
rect 23506 1380 23522 1444
rect 23586 1380 23602 1444
rect 23666 1380 23682 1444
rect 23746 1380 23888 1444
rect 23952 1380 23968 1444
rect 24032 1380 24048 1444
rect 24112 1380 24128 1444
rect 24192 1380 24208 1444
rect 24272 1380 24288 1444
rect 24352 1380 24494 1444
rect 24558 1380 24574 1444
rect 24638 1380 24654 1444
rect 24718 1380 24734 1444
rect 24798 1380 24814 1444
rect 24878 1380 24894 1444
rect 24958 1380 25100 1444
rect 25164 1380 25180 1444
rect 25244 1380 25260 1444
rect 25324 1380 25340 1444
rect 25404 1380 25420 1444
rect 25484 1380 25500 1444
rect 25564 1380 25706 1444
rect 25770 1380 25786 1444
rect 25850 1380 25866 1444
rect 25930 1380 25946 1444
rect 26010 1380 26026 1444
rect 26090 1380 26106 1444
rect 26170 1380 26312 1444
rect 26376 1380 26392 1444
rect 26456 1380 26472 1444
rect 26536 1380 26552 1444
rect 26616 1380 26632 1444
rect 26696 1380 26712 1444
rect 26776 1380 26918 1444
rect 26982 1380 26998 1444
rect 27062 1380 27078 1444
rect 27142 1380 27158 1444
rect 27222 1380 27238 1444
rect 27302 1380 27318 1444
rect 27382 1380 27524 1444
rect 27588 1380 27604 1444
rect 27668 1380 27684 1444
rect 27748 1380 27764 1444
rect 27828 1380 27844 1444
rect 27908 1380 27924 1444
rect 27988 1380 28130 1444
rect 28194 1380 28210 1444
rect 28274 1380 28290 1444
rect 28354 1380 28370 1444
rect 28434 1380 28450 1444
rect 28514 1380 28530 1444
rect 28594 1380 28736 1444
rect 28800 1380 28816 1444
rect 28880 1380 28896 1444
rect 28960 1380 28976 1444
rect 29040 1380 29056 1444
rect 29120 1380 29136 1444
rect 29200 1380 29342 1444
rect 29406 1380 29422 1444
rect 29486 1380 29502 1444
rect 29566 1380 29582 1444
rect 29646 1380 29662 1444
rect 29726 1380 29742 1444
rect 29806 1380 29948 1444
rect 30012 1380 30028 1444
rect 30092 1380 30108 1444
rect 30172 1380 30188 1444
rect 30252 1380 30268 1444
rect 30332 1380 30348 1444
rect 30412 1380 30554 1444
rect 30618 1380 30634 1444
rect 30698 1380 30714 1444
rect 30778 1380 30794 1444
rect 30858 1380 30874 1444
rect 30938 1380 30954 1444
rect 31018 1380 31160 1444
rect 31224 1380 31240 1444
rect 31304 1380 31320 1444
rect 31384 1380 31400 1444
rect 31464 1380 31480 1444
rect 31544 1380 31560 1444
rect 31624 1380 31766 1444
rect 31830 1380 31846 1444
rect 31910 1380 31926 1444
rect 31990 1380 32006 1444
rect 32070 1380 32086 1444
rect 32150 1380 32166 1444
rect 32230 1380 32372 1444
rect 32436 1380 32452 1444
rect 32516 1380 32532 1444
rect 32596 1380 32612 1444
rect 32676 1380 32692 1444
rect 32756 1380 32772 1444
rect 32836 1380 32978 1444
rect 33042 1380 33058 1444
rect 33122 1380 33138 1444
rect 33202 1380 33218 1444
rect 33282 1380 33298 1444
rect 33362 1380 33378 1444
rect 33442 1380 33584 1444
rect 33648 1380 33664 1444
rect 33728 1380 33744 1444
rect 33808 1380 33824 1444
rect 33888 1380 33904 1444
rect 33968 1380 33984 1444
rect 34048 1380 34190 1444
rect 34254 1380 34270 1444
rect 34334 1380 34350 1444
rect 34414 1380 34430 1444
rect 34494 1380 34510 1444
rect 34574 1380 34590 1444
rect 34654 1380 34796 1444
rect 34860 1380 34876 1444
rect 34940 1380 34956 1444
rect 35020 1380 35036 1444
rect 35100 1380 35116 1444
rect 35180 1380 35196 1444
rect 35260 1380 35402 1444
rect 35466 1380 35482 1444
rect 35546 1380 35562 1444
rect 35626 1380 35642 1444
rect 35706 1380 35722 1444
rect 35786 1380 35802 1444
rect 35866 1380 36008 1444
rect 36072 1380 36088 1444
rect 36152 1380 36168 1444
rect 36232 1380 36248 1444
rect 36312 1380 36328 1444
rect 36392 1380 36408 1444
rect 36472 1380 36614 1444
rect 36678 1380 36694 1444
rect 36758 1380 36774 1444
rect 36838 1380 36854 1444
rect 36918 1380 36934 1444
rect 36998 1380 37014 1444
rect 37078 1380 37220 1444
rect 37284 1380 37300 1444
rect 37364 1380 37380 1444
rect 37444 1380 37460 1444
rect 37524 1380 37540 1444
rect 37604 1380 37620 1444
rect 37684 1380 37826 1444
rect 37890 1380 37906 1444
rect 37970 1380 37986 1444
rect 38050 1380 38066 1444
rect 38130 1380 38146 1444
rect 38210 1380 38226 1444
rect 38290 1380 38432 1444
rect 38496 1380 38512 1444
rect 38576 1380 38592 1444
rect 38656 1380 38672 1444
rect 38736 1380 38752 1444
rect 38816 1380 38832 1444
rect 38896 1380 39038 1444
rect 39102 1380 39118 1444
rect 39182 1380 39198 1444
rect 39262 1380 39278 1444
rect 39342 1380 39358 1444
rect 39422 1380 39438 1444
rect 39502 1380 39606 1444
rect 20148 1378 39606 1380
rect 20148 1224 20214 1378
rect 20148 1160 20149 1224
rect 20213 1160 20214 1224
rect 20148 1144 20214 1160
rect 20148 1080 20149 1144
rect 20213 1080 20214 1144
rect 20148 1064 20214 1080
rect 20148 1000 20149 1064
rect 20213 1000 20214 1064
rect 20148 984 20214 1000
rect 20148 920 20149 984
rect 20213 920 20214 984
rect 20148 904 20214 920
rect 20148 840 20149 904
rect 20213 840 20214 904
rect 20148 824 20214 840
rect 20148 760 20149 824
rect 20213 760 20214 824
rect 20148 744 20214 760
rect 20148 680 20149 744
rect 20213 680 20214 744
rect 20148 664 20214 680
rect 20148 600 20149 664
rect 20213 600 20214 664
rect 20148 584 20214 600
rect 20148 520 20149 584
rect 20213 520 20214 584
rect 20148 504 20214 520
rect 20148 440 20149 504
rect 20213 440 20214 504
rect 20148 350 20214 440
rect 20274 286 20334 1316
rect 20394 346 20454 1378
rect 20514 286 20574 1316
rect 20634 346 20694 1378
rect 20754 1224 20820 1378
rect 20754 1160 20755 1224
rect 20819 1160 20820 1224
rect 20754 1144 20820 1160
rect 20754 1080 20755 1144
rect 20819 1080 20820 1144
rect 20754 1064 20820 1080
rect 20754 1000 20755 1064
rect 20819 1000 20820 1064
rect 20754 984 20820 1000
rect 20754 920 20755 984
rect 20819 920 20820 984
rect 20754 904 20820 920
rect 20754 840 20755 904
rect 20819 840 20820 904
rect 20754 824 20820 840
rect 20754 760 20755 824
rect 20819 760 20820 824
rect 20754 744 20820 760
rect 20754 680 20755 744
rect 20819 680 20820 744
rect 20754 664 20820 680
rect 20754 600 20755 664
rect 20819 600 20820 664
rect 20754 584 20820 600
rect 20754 520 20755 584
rect 20819 520 20820 584
rect 20754 504 20820 520
rect 20754 440 20755 504
rect 20819 440 20820 504
rect 20754 350 20820 440
rect 20880 286 20940 1316
rect 21000 346 21060 1378
rect 21120 286 21180 1316
rect 21240 346 21300 1378
rect 21360 1224 21426 1378
rect 21360 1160 21361 1224
rect 21425 1160 21426 1224
rect 21360 1144 21426 1160
rect 21360 1080 21361 1144
rect 21425 1080 21426 1144
rect 21360 1064 21426 1080
rect 21360 1000 21361 1064
rect 21425 1000 21426 1064
rect 21360 984 21426 1000
rect 21360 920 21361 984
rect 21425 920 21426 984
rect 21360 904 21426 920
rect 21360 840 21361 904
rect 21425 840 21426 904
rect 21360 824 21426 840
rect 21360 760 21361 824
rect 21425 760 21426 824
rect 21360 744 21426 760
rect 21360 680 21361 744
rect 21425 680 21426 744
rect 21360 664 21426 680
rect 21360 600 21361 664
rect 21425 600 21426 664
rect 21360 584 21426 600
rect 21360 520 21361 584
rect 21425 520 21426 584
rect 21360 504 21426 520
rect 21360 440 21361 504
rect 21425 440 21426 504
rect 21360 350 21426 440
rect 21486 286 21546 1316
rect 21606 346 21666 1378
rect 21726 286 21786 1316
rect 21846 346 21906 1378
rect 21966 1224 22032 1378
rect 21966 1160 21967 1224
rect 22031 1160 22032 1224
rect 21966 1144 22032 1160
rect 21966 1080 21967 1144
rect 22031 1080 22032 1144
rect 21966 1064 22032 1080
rect 21966 1000 21967 1064
rect 22031 1000 22032 1064
rect 21966 984 22032 1000
rect 21966 920 21967 984
rect 22031 920 22032 984
rect 21966 904 22032 920
rect 21966 840 21967 904
rect 22031 840 22032 904
rect 21966 824 22032 840
rect 21966 760 21967 824
rect 22031 760 22032 824
rect 21966 744 22032 760
rect 21966 680 21967 744
rect 22031 680 22032 744
rect 21966 664 22032 680
rect 21966 600 21967 664
rect 22031 600 22032 664
rect 21966 584 22032 600
rect 21966 520 21967 584
rect 22031 520 22032 584
rect 21966 504 22032 520
rect 21966 440 21967 504
rect 22031 440 22032 504
rect 21966 350 22032 440
rect 22092 286 22152 1316
rect 22212 346 22272 1378
rect 22332 286 22392 1316
rect 22452 346 22512 1378
rect 22572 1224 22638 1378
rect 22572 1160 22573 1224
rect 22637 1160 22638 1224
rect 22572 1144 22638 1160
rect 22572 1080 22573 1144
rect 22637 1080 22638 1144
rect 22572 1064 22638 1080
rect 22572 1000 22573 1064
rect 22637 1000 22638 1064
rect 22572 984 22638 1000
rect 22572 920 22573 984
rect 22637 920 22638 984
rect 22572 904 22638 920
rect 22572 840 22573 904
rect 22637 840 22638 904
rect 22572 824 22638 840
rect 22572 760 22573 824
rect 22637 760 22638 824
rect 22572 744 22638 760
rect 22572 680 22573 744
rect 22637 680 22638 744
rect 22572 664 22638 680
rect 22572 600 22573 664
rect 22637 600 22638 664
rect 22572 584 22638 600
rect 22572 520 22573 584
rect 22637 520 22638 584
rect 22572 504 22638 520
rect 22572 440 22573 504
rect 22637 440 22638 504
rect 22572 350 22638 440
rect 22698 286 22758 1316
rect 22818 346 22878 1378
rect 22938 286 22998 1316
rect 23058 346 23118 1378
rect 23178 1224 23244 1378
rect 23178 1160 23179 1224
rect 23243 1160 23244 1224
rect 23178 1144 23244 1160
rect 23178 1080 23179 1144
rect 23243 1080 23244 1144
rect 23178 1064 23244 1080
rect 23178 1000 23179 1064
rect 23243 1000 23244 1064
rect 23178 984 23244 1000
rect 23178 920 23179 984
rect 23243 920 23244 984
rect 23178 904 23244 920
rect 23178 840 23179 904
rect 23243 840 23244 904
rect 23178 824 23244 840
rect 23178 760 23179 824
rect 23243 760 23244 824
rect 23178 744 23244 760
rect 23178 680 23179 744
rect 23243 680 23244 744
rect 23178 664 23244 680
rect 23178 600 23179 664
rect 23243 600 23244 664
rect 23178 584 23244 600
rect 23178 520 23179 584
rect 23243 520 23244 584
rect 23178 504 23244 520
rect 23178 440 23179 504
rect 23243 440 23244 504
rect 23178 350 23244 440
rect 23304 286 23364 1316
rect 23424 346 23484 1378
rect 23544 286 23604 1316
rect 23664 346 23724 1378
rect 23784 1224 23850 1378
rect 23784 1160 23785 1224
rect 23849 1160 23850 1224
rect 23784 1144 23850 1160
rect 23784 1080 23785 1144
rect 23849 1080 23850 1144
rect 23784 1064 23850 1080
rect 23784 1000 23785 1064
rect 23849 1000 23850 1064
rect 23784 984 23850 1000
rect 23784 920 23785 984
rect 23849 920 23850 984
rect 23784 904 23850 920
rect 23784 840 23785 904
rect 23849 840 23850 904
rect 23784 824 23850 840
rect 23784 760 23785 824
rect 23849 760 23850 824
rect 23784 744 23850 760
rect 23784 680 23785 744
rect 23849 680 23850 744
rect 23784 664 23850 680
rect 23784 600 23785 664
rect 23849 600 23850 664
rect 23784 584 23850 600
rect 23784 520 23785 584
rect 23849 520 23850 584
rect 23784 504 23850 520
rect 23784 440 23785 504
rect 23849 440 23850 504
rect 23784 350 23850 440
rect 23910 286 23970 1316
rect 24030 346 24090 1378
rect 24150 286 24210 1316
rect 24270 346 24330 1378
rect 24390 1224 24456 1378
rect 24390 1160 24391 1224
rect 24455 1160 24456 1224
rect 24390 1144 24456 1160
rect 24390 1080 24391 1144
rect 24455 1080 24456 1144
rect 24390 1064 24456 1080
rect 24390 1000 24391 1064
rect 24455 1000 24456 1064
rect 24390 984 24456 1000
rect 24390 920 24391 984
rect 24455 920 24456 984
rect 24390 904 24456 920
rect 24390 840 24391 904
rect 24455 840 24456 904
rect 24390 824 24456 840
rect 24390 760 24391 824
rect 24455 760 24456 824
rect 24390 744 24456 760
rect 24390 680 24391 744
rect 24455 680 24456 744
rect 24390 664 24456 680
rect 24390 600 24391 664
rect 24455 600 24456 664
rect 24390 584 24456 600
rect 24390 520 24391 584
rect 24455 520 24456 584
rect 24390 504 24456 520
rect 24390 440 24391 504
rect 24455 440 24456 504
rect 24390 350 24456 440
rect 24516 286 24576 1316
rect 24636 346 24696 1378
rect 24756 286 24816 1316
rect 24876 346 24936 1378
rect 24996 1224 25062 1378
rect 24996 1160 24997 1224
rect 25061 1160 25062 1224
rect 24996 1144 25062 1160
rect 24996 1080 24997 1144
rect 25061 1080 25062 1144
rect 24996 1064 25062 1080
rect 24996 1000 24997 1064
rect 25061 1000 25062 1064
rect 24996 984 25062 1000
rect 24996 920 24997 984
rect 25061 920 25062 984
rect 24996 904 25062 920
rect 24996 840 24997 904
rect 25061 840 25062 904
rect 24996 824 25062 840
rect 24996 760 24997 824
rect 25061 760 25062 824
rect 24996 744 25062 760
rect 24996 680 24997 744
rect 25061 680 25062 744
rect 24996 664 25062 680
rect 24996 600 24997 664
rect 25061 600 25062 664
rect 24996 584 25062 600
rect 24996 520 24997 584
rect 25061 520 25062 584
rect 24996 504 25062 520
rect 24996 440 24997 504
rect 25061 440 25062 504
rect 24996 350 25062 440
rect 25122 286 25182 1316
rect 25242 346 25302 1378
rect 25362 286 25422 1316
rect 25482 346 25542 1378
rect 25602 1224 25668 1378
rect 25602 1160 25603 1224
rect 25667 1160 25668 1224
rect 25602 1144 25668 1160
rect 25602 1080 25603 1144
rect 25667 1080 25668 1144
rect 25602 1064 25668 1080
rect 25602 1000 25603 1064
rect 25667 1000 25668 1064
rect 25602 984 25668 1000
rect 25602 920 25603 984
rect 25667 920 25668 984
rect 25602 904 25668 920
rect 25602 840 25603 904
rect 25667 840 25668 904
rect 25602 824 25668 840
rect 25602 760 25603 824
rect 25667 760 25668 824
rect 25602 744 25668 760
rect 25602 680 25603 744
rect 25667 680 25668 744
rect 25602 664 25668 680
rect 25602 600 25603 664
rect 25667 600 25668 664
rect 25602 584 25668 600
rect 25602 520 25603 584
rect 25667 520 25668 584
rect 25602 504 25668 520
rect 25602 440 25603 504
rect 25667 440 25668 504
rect 25602 350 25668 440
rect 25728 286 25788 1316
rect 25848 346 25908 1378
rect 25968 286 26028 1316
rect 26088 346 26148 1378
rect 26208 1224 26274 1378
rect 26208 1160 26209 1224
rect 26273 1160 26274 1224
rect 26208 1144 26274 1160
rect 26208 1080 26209 1144
rect 26273 1080 26274 1144
rect 26208 1064 26274 1080
rect 26208 1000 26209 1064
rect 26273 1000 26274 1064
rect 26208 984 26274 1000
rect 26208 920 26209 984
rect 26273 920 26274 984
rect 26208 904 26274 920
rect 26208 840 26209 904
rect 26273 840 26274 904
rect 26208 824 26274 840
rect 26208 760 26209 824
rect 26273 760 26274 824
rect 26208 744 26274 760
rect 26208 680 26209 744
rect 26273 680 26274 744
rect 26208 664 26274 680
rect 26208 600 26209 664
rect 26273 600 26274 664
rect 26208 584 26274 600
rect 26208 520 26209 584
rect 26273 520 26274 584
rect 26208 504 26274 520
rect 26208 440 26209 504
rect 26273 440 26274 504
rect 26208 350 26274 440
rect 26334 286 26394 1316
rect 26454 346 26514 1378
rect 26574 286 26634 1316
rect 26694 346 26754 1378
rect 26814 1224 26880 1378
rect 26814 1160 26815 1224
rect 26879 1160 26880 1224
rect 26814 1144 26880 1160
rect 26814 1080 26815 1144
rect 26879 1080 26880 1144
rect 26814 1064 26880 1080
rect 26814 1000 26815 1064
rect 26879 1000 26880 1064
rect 26814 984 26880 1000
rect 26814 920 26815 984
rect 26879 920 26880 984
rect 26814 904 26880 920
rect 26814 840 26815 904
rect 26879 840 26880 904
rect 26814 824 26880 840
rect 26814 760 26815 824
rect 26879 760 26880 824
rect 26814 744 26880 760
rect 26814 680 26815 744
rect 26879 680 26880 744
rect 26814 664 26880 680
rect 26814 600 26815 664
rect 26879 600 26880 664
rect 26814 584 26880 600
rect 26814 520 26815 584
rect 26879 520 26880 584
rect 26814 504 26880 520
rect 26814 440 26815 504
rect 26879 440 26880 504
rect 26814 350 26880 440
rect 26940 286 27000 1316
rect 27060 346 27120 1378
rect 27180 286 27240 1316
rect 27300 346 27360 1378
rect 27420 1224 27486 1378
rect 27420 1160 27421 1224
rect 27485 1160 27486 1224
rect 27420 1144 27486 1160
rect 27420 1080 27421 1144
rect 27485 1080 27486 1144
rect 27420 1064 27486 1080
rect 27420 1000 27421 1064
rect 27485 1000 27486 1064
rect 27420 984 27486 1000
rect 27420 920 27421 984
rect 27485 920 27486 984
rect 27420 904 27486 920
rect 27420 840 27421 904
rect 27485 840 27486 904
rect 27420 824 27486 840
rect 27420 760 27421 824
rect 27485 760 27486 824
rect 27420 744 27486 760
rect 27420 680 27421 744
rect 27485 680 27486 744
rect 27420 664 27486 680
rect 27420 600 27421 664
rect 27485 600 27486 664
rect 27420 584 27486 600
rect 27420 520 27421 584
rect 27485 520 27486 584
rect 27420 504 27486 520
rect 27420 440 27421 504
rect 27485 440 27486 504
rect 27420 350 27486 440
rect 27546 286 27606 1316
rect 27666 346 27726 1378
rect 27786 286 27846 1316
rect 27906 346 27966 1378
rect 28026 1224 28092 1378
rect 28026 1160 28027 1224
rect 28091 1160 28092 1224
rect 28026 1144 28092 1160
rect 28026 1080 28027 1144
rect 28091 1080 28092 1144
rect 28026 1064 28092 1080
rect 28026 1000 28027 1064
rect 28091 1000 28092 1064
rect 28026 984 28092 1000
rect 28026 920 28027 984
rect 28091 920 28092 984
rect 28026 904 28092 920
rect 28026 840 28027 904
rect 28091 840 28092 904
rect 28026 824 28092 840
rect 28026 760 28027 824
rect 28091 760 28092 824
rect 28026 744 28092 760
rect 28026 680 28027 744
rect 28091 680 28092 744
rect 28026 664 28092 680
rect 28026 600 28027 664
rect 28091 600 28092 664
rect 28026 584 28092 600
rect 28026 520 28027 584
rect 28091 520 28092 584
rect 28026 504 28092 520
rect 28026 440 28027 504
rect 28091 440 28092 504
rect 28026 350 28092 440
rect 28152 286 28212 1316
rect 28272 346 28332 1378
rect 28392 286 28452 1316
rect 28512 346 28572 1378
rect 28632 1224 28698 1378
rect 28632 1160 28633 1224
rect 28697 1160 28698 1224
rect 28632 1144 28698 1160
rect 28632 1080 28633 1144
rect 28697 1080 28698 1144
rect 28632 1064 28698 1080
rect 28632 1000 28633 1064
rect 28697 1000 28698 1064
rect 28632 984 28698 1000
rect 28632 920 28633 984
rect 28697 920 28698 984
rect 28632 904 28698 920
rect 28632 840 28633 904
rect 28697 840 28698 904
rect 28632 824 28698 840
rect 28632 760 28633 824
rect 28697 760 28698 824
rect 28632 744 28698 760
rect 28632 680 28633 744
rect 28697 680 28698 744
rect 28632 664 28698 680
rect 28632 600 28633 664
rect 28697 600 28698 664
rect 28632 584 28698 600
rect 28632 520 28633 584
rect 28697 520 28698 584
rect 28632 504 28698 520
rect 28632 440 28633 504
rect 28697 440 28698 504
rect 28632 350 28698 440
rect 28758 286 28818 1316
rect 28878 346 28938 1378
rect 28998 286 29058 1316
rect 29118 346 29178 1378
rect 29238 1224 29304 1378
rect 29238 1160 29239 1224
rect 29303 1160 29304 1224
rect 29238 1144 29304 1160
rect 29238 1080 29239 1144
rect 29303 1080 29304 1144
rect 29238 1064 29304 1080
rect 29238 1000 29239 1064
rect 29303 1000 29304 1064
rect 29238 984 29304 1000
rect 29238 920 29239 984
rect 29303 920 29304 984
rect 29238 904 29304 920
rect 29238 840 29239 904
rect 29303 840 29304 904
rect 29238 824 29304 840
rect 29238 760 29239 824
rect 29303 760 29304 824
rect 29238 744 29304 760
rect 29238 680 29239 744
rect 29303 680 29304 744
rect 29238 664 29304 680
rect 29238 600 29239 664
rect 29303 600 29304 664
rect 29238 584 29304 600
rect 29238 520 29239 584
rect 29303 520 29304 584
rect 29238 504 29304 520
rect 29238 440 29239 504
rect 29303 440 29304 504
rect 29238 350 29304 440
rect 29364 286 29424 1316
rect 29484 346 29544 1378
rect 29604 286 29664 1316
rect 29724 346 29784 1378
rect 29844 1224 29910 1378
rect 29844 1160 29845 1224
rect 29909 1160 29910 1224
rect 29844 1144 29910 1160
rect 29844 1080 29845 1144
rect 29909 1080 29910 1144
rect 29844 1064 29910 1080
rect 29844 1000 29845 1064
rect 29909 1000 29910 1064
rect 29844 984 29910 1000
rect 29844 920 29845 984
rect 29909 920 29910 984
rect 29844 904 29910 920
rect 29844 840 29845 904
rect 29909 840 29910 904
rect 29844 824 29910 840
rect 29844 760 29845 824
rect 29909 760 29910 824
rect 29844 744 29910 760
rect 29844 680 29845 744
rect 29909 680 29910 744
rect 29844 664 29910 680
rect 29844 600 29845 664
rect 29909 600 29910 664
rect 29844 584 29910 600
rect 29844 520 29845 584
rect 29909 520 29910 584
rect 29844 504 29910 520
rect 29844 440 29845 504
rect 29909 440 29910 504
rect 29844 350 29910 440
rect 29970 286 30030 1316
rect 30090 346 30150 1378
rect 30210 286 30270 1316
rect 30330 346 30390 1378
rect 30450 1224 30516 1378
rect 30450 1160 30451 1224
rect 30515 1160 30516 1224
rect 30450 1144 30516 1160
rect 30450 1080 30451 1144
rect 30515 1080 30516 1144
rect 30450 1064 30516 1080
rect 30450 1000 30451 1064
rect 30515 1000 30516 1064
rect 30450 984 30516 1000
rect 30450 920 30451 984
rect 30515 920 30516 984
rect 30450 904 30516 920
rect 30450 840 30451 904
rect 30515 840 30516 904
rect 30450 824 30516 840
rect 30450 760 30451 824
rect 30515 760 30516 824
rect 30450 744 30516 760
rect 30450 680 30451 744
rect 30515 680 30516 744
rect 30450 664 30516 680
rect 30450 600 30451 664
rect 30515 600 30516 664
rect 30450 584 30516 600
rect 30450 520 30451 584
rect 30515 520 30516 584
rect 30450 504 30516 520
rect 30450 440 30451 504
rect 30515 440 30516 504
rect 30450 350 30516 440
rect 30576 286 30636 1316
rect 30696 346 30756 1378
rect 30816 286 30876 1316
rect 30936 346 30996 1378
rect 31056 1224 31122 1378
rect 31056 1160 31057 1224
rect 31121 1160 31122 1224
rect 31056 1144 31122 1160
rect 31056 1080 31057 1144
rect 31121 1080 31122 1144
rect 31056 1064 31122 1080
rect 31056 1000 31057 1064
rect 31121 1000 31122 1064
rect 31056 984 31122 1000
rect 31056 920 31057 984
rect 31121 920 31122 984
rect 31056 904 31122 920
rect 31056 840 31057 904
rect 31121 840 31122 904
rect 31056 824 31122 840
rect 31056 760 31057 824
rect 31121 760 31122 824
rect 31056 744 31122 760
rect 31056 680 31057 744
rect 31121 680 31122 744
rect 31056 664 31122 680
rect 31056 600 31057 664
rect 31121 600 31122 664
rect 31056 584 31122 600
rect 31056 520 31057 584
rect 31121 520 31122 584
rect 31056 504 31122 520
rect 31056 440 31057 504
rect 31121 440 31122 504
rect 31056 350 31122 440
rect 31182 286 31242 1316
rect 31302 346 31362 1378
rect 31422 286 31482 1316
rect 31542 346 31602 1378
rect 31662 1224 31728 1378
rect 31662 1160 31663 1224
rect 31727 1160 31728 1224
rect 31662 1144 31728 1160
rect 31662 1080 31663 1144
rect 31727 1080 31728 1144
rect 31662 1064 31728 1080
rect 31662 1000 31663 1064
rect 31727 1000 31728 1064
rect 31662 984 31728 1000
rect 31662 920 31663 984
rect 31727 920 31728 984
rect 31662 904 31728 920
rect 31662 840 31663 904
rect 31727 840 31728 904
rect 31662 824 31728 840
rect 31662 760 31663 824
rect 31727 760 31728 824
rect 31662 744 31728 760
rect 31662 680 31663 744
rect 31727 680 31728 744
rect 31662 664 31728 680
rect 31662 600 31663 664
rect 31727 600 31728 664
rect 31662 584 31728 600
rect 31662 520 31663 584
rect 31727 520 31728 584
rect 31662 504 31728 520
rect 31662 440 31663 504
rect 31727 440 31728 504
rect 31662 350 31728 440
rect 31788 286 31848 1316
rect 31908 346 31968 1378
rect 32028 286 32088 1316
rect 32148 346 32208 1378
rect 32268 1224 32334 1378
rect 32268 1160 32269 1224
rect 32333 1160 32334 1224
rect 32268 1144 32334 1160
rect 32268 1080 32269 1144
rect 32333 1080 32334 1144
rect 32268 1064 32334 1080
rect 32268 1000 32269 1064
rect 32333 1000 32334 1064
rect 32268 984 32334 1000
rect 32268 920 32269 984
rect 32333 920 32334 984
rect 32268 904 32334 920
rect 32268 840 32269 904
rect 32333 840 32334 904
rect 32268 824 32334 840
rect 32268 760 32269 824
rect 32333 760 32334 824
rect 32268 744 32334 760
rect 32268 680 32269 744
rect 32333 680 32334 744
rect 32268 664 32334 680
rect 32268 600 32269 664
rect 32333 600 32334 664
rect 32268 584 32334 600
rect 32268 520 32269 584
rect 32333 520 32334 584
rect 32268 504 32334 520
rect 32268 440 32269 504
rect 32333 440 32334 504
rect 32268 350 32334 440
rect 32394 286 32454 1316
rect 32514 346 32574 1378
rect 32634 286 32694 1316
rect 32754 346 32814 1378
rect 32874 1224 32940 1378
rect 32874 1160 32875 1224
rect 32939 1160 32940 1224
rect 32874 1144 32940 1160
rect 32874 1080 32875 1144
rect 32939 1080 32940 1144
rect 32874 1064 32940 1080
rect 32874 1000 32875 1064
rect 32939 1000 32940 1064
rect 32874 984 32940 1000
rect 32874 920 32875 984
rect 32939 920 32940 984
rect 32874 904 32940 920
rect 32874 840 32875 904
rect 32939 840 32940 904
rect 32874 824 32940 840
rect 32874 760 32875 824
rect 32939 760 32940 824
rect 32874 744 32940 760
rect 32874 680 32875 744
rect 32939 680 32940 744
rect 32874 664 32940 680
rect 32874 600 32875 664
rect 32939 600 32940 664
rect 32874 584 32940 600
rect 32874 520 32875 584
rect 32939 520 32940 584
rect 32874 504 32940 520
rect 32874 440 32875 504
rect 32939 440 32940 504
rect 32874 350 32940 440
rect 33000 286 33060 1316
rect 33120 346 33180 1378
rect 33240 286 33300 1316
rect 33360 346 33420 1378
rect 33480 1224 33546 1378
rect 33480 1160 33481 1224
rect 33545 1160 33546 1224
rect 33480 1144 33546 1160
rect 33480 1080 33481 1144
rect 33545 1080 33546 1144
rect 33480 1064 33546 1080
rect 33480 1000 33481 1064
rect 33545 1000 33546 1064
rect 33480 984 33546 1000
rect 33480 920 33481 984
rect 33545 920 33546 984
rect 33480 904 33546 920
rect 33480 840 33481 904
rect 33545 840 33546 904
rect 33480 824 33546 840
rect 33480 760 33481 824
rect 33545 760 33546 824
rect 33480 744 33546 760
rect 33480 680 33481 744
rect 33545 680 33546 744
rect 33480 664 33546 680
rect 33480 600 33481 664
rect 33545 600 33546 664
rect 33480 584 33546 600
rect 33480 520 33481 584
rect 33545 520 33546 584
rect 33480 504 33546 520
rect 33480 440 33481 504
rect 33545 440 33546 504
rect 33480 350 33546 440
rect 33606 286 33666 1316
rect 33726 346 33786 1378
rect 33846 286 33906 1316
rect 33966 346 34026 1378
rect 34086 1224 34152 1378
rect 34086 1160 34087 1224
rect 34151 1160 34152 1224
rect 34086 1144 34152 1160
rect 34086 1080 34087 1144
rect 34151 1080 34152 1144
rect 34086 1064 34152 1080
rect 34086 1000 34087 1064
rect 34151 1000 34152 1064
rect 34086 984 34152 1000
rect 34086 920 34087 984
rect 34151 920 34152 984
rect 34086 904 34152 920
rect 34086 840 34087 904
rect 34151 840 34152 904
rect 34086 824 34152 840
rect 34086 760 34087 824
rect 34151 760 34152 824
rect 34086 744 34152 760
rect 34086 680 34087 744
rect 34151 680 34152 744
rect 34086 664 34152 680
rect 34086 600 34087 664
rect 34151 600 34152 664
rect 34086 584 34152 600
rect 34086 520 34087 584
rect 34151 520 34152 584
rect 34086 504 34152 520
rect 34086 440 34087 504
rect 34151 440 34152 504
rect 34086 350 34152 440
rect 34212 286 34272 1316
rect 34332 346 34392 1378
rect 34452 286 34512 1316
rect 34572 346 34632 1378
rect 34692 1224 34758 1378
rect 34692 1160 34693 1224
rect 34757 1160 34758 1224
rect 34692 1144 34758 1160
rect 34692 1080 34693 1144
rect 34757 1080 34758 1144
rect 34692 1064 34758 1080
rect 34692 1000 34693 1064
rect 34757 1000 34758 1064
rect 34692 984 34758 1000
rect 34692 920 34693 984
rect 34757 920 34758 984
rect 34692 904 34758 920
rect 34692 840 34693 904
rect 34757 840 34758 904
rect 34692 824 34758 840
rect 34692 760 34693 824
rect 34757 760 34758 824
rect 34692 744 34758 760
rect 34692 680 34693 744
rect 34757 680 34758 744
rect 34692 664 34758 680
rect 34692 600 34693 664
rect 34757 600 34758 664
rect 34692 584 34758 600
rect 34692 520 34693 584
rect 34757 520 34758 584
rect 34692 504 34758 520
rect 34692 440 34693 504
rect 34757 440 34758 504
rect 34692 350 34758 440
rect 34818 286 34878 1316
rect 34938 346 34998 1378
rect 35058 286 35118 1316
rect 35178 346 35238 1378
rect 35298 1224 35364 1378
rect 35298 1160 35299 1224
rect 35363 1160 35364 1224
rect 35298 1144 35364 1160
rect 35298 1080 35299 1144
rect 35363 1080 35364 1144
rect 35298 1064 35364 1080
rect 35298 1000 35299 1064
rect 35363 1000 35364 1064
rect 35298 984 35364 1000
rect 35298 920 35299 984
rect 35363 920 35364 984
rect 35298 904 35364 920
rect 35298 840 35299 904
rect 35363 840 35364 904
rect 35298 824 35364 840
rect 35298 760 35299 824
rect 35363 760 35364 824
rect 35298 744 35364 760
rect 35298 680 35299 744
rect 35363 680 35364 744
rect 35298 664 35364 680
rect 35298 600 35299 664
rect 35363 600 35364 664
rect 35298 584 35364 600
rect 35298 520 35299 584
rect 35363 520 35364 584
rect 35298 504 35364 520
rect 35298 440 35299 504
rect 35363 440 35364 504
rect 35298 350 35364 440
rect 35424 286 35484 1316
rect 35544 346 35604 1378
rect 35664 286 35724 1316
rect 35784 346 35844 1378
rect 35904 1224 35970 1378
rect 35904 1160 35905 1224
rect 35969 1160 35970 1224
rect 35904 1144 35970 1160
rect 35904 1080 35905 1144
rect 35969 1080 35970 1144
rect 35904 1064 35970 1080
rect 35904 1000 35905 1064
rect 35969 1000 35970 1064
rect 35904 984 35970 1000
rect 35904 920 35905 984
rect 35969 920 35970 984
rect 35904 904 35970 920
rect 35904 840 35905 904
rect 35969 840 35970 904
rect 35904 824 35970 840
rect 35904 760 35905 824
rect 35969 760 35970 824
rect 35904 744 35970 760
rect 35904 680 35905 744
rect 35969 680 35970 744
rect 35904 664 35970 680
rect 35904 600 35905 664
rect 35969 600 35970 664
rect 35904 584 35970 600
rect 35904 520 35905 584
rect 35969 520 35970 584
rect 35904 504 35970 520
rect 35904 440 35905 504
rect 35969 440 35970 504
rect 35904 350 35970 440
rect 36030 286 36090 1316
rect 36150 346 36210 1378
rect 36270 286 36330 1316
rect 36390 346 36450 1378
rect 36510 1224 36576 1378
rect 36510 1160 36511 1224
rect 36575 1160 36576 1224
rect 36510 1144 36576 1160
rect 36510 1080 36511 1144
rect 36575 1080 36576 1144
rect 36510 1064 36576 1080
rect 36510 1000 36511 1064
rect 36575 1000 36576 1064
rect 36510 984 36576 1000
rect 36510 920 36511 984
rect 36575 920 36576 984
rect 36510 904 36576 920
rect 36510 840 36511 904
rect 36575 840 36576 904
rect 36510 824 36576 840
rect 36510 760 36511 824
rect 36575 760 36576 824
rect 36510 744 36576 760
rect 36510 680 36511 744
rect 36575 680 36576 744
rect 36510 664 36576 680
rect 36510 600 36511 664
rect 36575 600 36576 664
rect 36510 584 36576 600
rect 36510 520 36511 584
rect 36575 520 36576 584
rect 36510 504 36576 520
rect 36510 440 36511 504
rect 36575 440 36576 504
rect 36510 350 36576 440
rect 36636 286 36696 1316
rect 36756 346 36816 1378
rect 36876 286 36936 1316
rect 36996 346 37056 1378
rect 37116 1224 37182 1378
rect 37116 1160 37117 1224
rect 37181 1160 37182 1224
rect 37116 1144 37182 1160
rect 37116 1080 37117 1144
rect 37181 1080 37182 1144
rect 37116 1064 37182 1080
rect 37116 1000 37117 1064
rect 37181 1000 37182 1064
rect 37116 984 37182 1000
rect 37116 920 37117 984
rect 37181 920 37182 984
rect 37116 904 37182 920
rect 37116 840 37117 904
rect 37181 840 37182 904
rect 37116 824 37182 840
rect 37116 760 37117 824
rect 37181 760 37182 824
rect 37116 744 37182 760
rect 37116 680 37117 744
rect 37181 680 37182 744
rect 37116 664 37182 680
rect 37116 600 37117 664
rect 37181 600 37182 664
rect 37116 584 37182 600
rect 37116 520 37117 584
rect 37181 520 37182 584
rect 37116 504 37182 520
rect 37116 440 37117 504
rect 37181 440 37182 504
rect 37116 350 37182 440
rect 37242 286 37302 1316
rect 37362 346 37422 1378
rect 37482 286 37542 1316
rect 37602 346 37662 1378
rect 37722 1224 37788 1378
rect 37722 1160 37723 1224
rect 37787 1160 37788 1224
rect 37722 1144 37788 1160
rect 37722 1080 37723 1144
rect 37787 1080 37788 1144
rect 37722 1064 37788 1080
rect 37722 1000 37723 1064
rect 37787 1000 37788 1064
rect 37722 984 37788 1000
rect 37722 920 37723 984
rect 37787 920 37788 984
rect 37722 904 37788 920
rect 37722 840 37723 904
rect 37787 840 37788 904
rect 37722 824 37788 840
rect 37722 760 37723 824
rect 37787 760 37788 824
rect 37722 744 37788 760
rect 37722 680 37723 744
rect 37787 680 37788 744
rect 37722 664 37788 680
rect 37722 600 37723 664
rect 37787 600 37788 664
rect 37722 584 37788 600
rect 37722 520 37723 584
rect 37787 520 37788 584
rect 37722 504 37788 520
rect 37722 440 37723 504
rect 37787 440 37788 504
rect 37722 350 37788 440
rect 37848 286 37908 1316
rect 37968 346 38028 1378
rect 38088 286 38148 1316
rect 38208 346 38268 1378
rect 38328 1224 38394 1378
rect 38328 1160 38329 1224
rect 38393 1160 38394 1224
rect 38328 1144 38394 1160
rect 38328 1080 38329 1144
rect 38393 1080 38394 1144
rect 38328 1064 38394 1080
rect 38328 1000 38329 1064
rect 38393 1000 38394 1064
rect 38328 984 38394 1000
rect 38328 920 38329 984
rect 38393 920 38394 984
rect 38328 904 38394 920
rect 38328 840 38329 904
rect 38393 840 38394 904
rect 38328 824 38394 840
rect 38328 760 38329 824
rect 38393 760 38394 824
rect 38328 744 38394 760
rect 38328 680 38329 744
rect 38393 680 38394 744
rect 38328 664 38394 680
rect 38328 600 38329 664
rect 38393 600 38394 664
rect 38328 584 38394 600
rect 38328 520 38329 584
rect 38393 520 38394 584
rect 38328 504 38394 520
rect 38328 440 38329 504
rect 38393 440 38394 504
rect 38328 350 38394 440
rect 38454 286 38514 1316
rect 38574 346 38634 1378
rect 38694 286 38754 1316
rect 38814 346 38874 1378
rect 38934 1224 39000 1378
rect 38934 1160 38935 1224
rect 38999 1160 39000 1224
rect 38934 1144 39000 1160
rect 38934 1080 38935 1144
rect 38999 1080 39000 1144
rect 38934 1064 39000 1080
rect 38934 1000 38935 1064
rect 38999 1000 39000 1064
rect 38934 984 39000 1000
rect 38934 920 38935 984
rect 38999 920 39000 984
rect 38934 904 39000 920
rect 38934 840 38935 904
rect 38999 840 39000 904
rect 38934 824 39000 840
rect 38934 760 38935 824
rect 38999 760 39000 824
rect 38934 744 39000 760
rect 38934 680 38935 744
rect 38999 680 39000 744
rect 38934 664 39000 680
rect 38934 600 38935 664
rect 38999 600 39000 664
rect 38934 584 39000 600
rect 38934 520 38935 584
rect 38999 520 39000 584
rect 38934 504 39000 520
rect 38934 440 38935 504
rect 38999 440 39000 504
rect 38934 350 39000 440
rect 39060 286 39120 1316
rect 39180 346 39240 1378
rect 39300 286 39360 1316
rect 39420 346 39480 1378
rect 39540 1224 39606 1378
rect 39540 1160 39541 1224
rect 39605 1160 39606 1224
rect 39540 1144 39606 1160
rect 39540 1080 39541 1144
rect 39605 1080 39606 1144
rect 39540 1064 39606 1080
rect 39540 1000 39541 1064
rect 39605 1000 39606 1064
rect 39540 984 39606 1000
rect 39540 920 39541 984
rect 39605 920 39606 984
rect 39540 904 39606 920
rect 39540 840 39541 904
rect 39605 840 39606 904
rect 39540 824 39606 840
rect 39540 760 39541 824
rect 39605 760 39606 824
rect 39540 744 39606 760
rect 39540 680 39541 744
rect 39605 680 39606 744
rect 39540 664 39606 680
rect 39540 600 39541 664
rect 39605 600 39606 664
rect 39540 584 39606 600
rect 39540 520 39541 584
rect 39605 520 39606 584
rect 39540 504 39606 520
rect 39540 440 39541 504
rect 39605 440 39606 504
rect 39540 350 39606 440
rect -459 284 213 286
rect -459 220 -355 284
rect -291 220 -275 284
rect -211 220 -195 284
rect -131 220 -115 284
rect -51 220 -35 284
rect 29 220 45 284
rect 109 220 213 284
rect -459 218 213 220
rect 355 284 1027 286
rect 355 220 459 284
rect 523 220 539 284
rect 603 220 619 284
rect 683 220 699 284
rect 763 220 779 284
rect 843 220 859 284
rect 923 220 1027 284
rect 355 218 1027 220
rect 1267 284 2545 286
rect 1267 220 1371 284
rect 1435 220 1451 284
rect 1515 220 1531 284
rect 1595 220 1611 284
rect 1675 220 1691 284
rect 1755 220 1771 284
rect 1835 220 1977 284
rect 2041 220 2057 284
rect 2121 220 2137 284
rect 2201 220 2217 284
rect 2281 220 2297 284
rect 2361 220 2377 284
rect 2441 220 2545 284
rect 1267 218 2545 220
rect 2801 284 5291 286
rect 2801 220 2905 284
rect 2969 220 2985 284
rect 3049 220 3065 284
rect 3129 220 3145 284
rect 3209 220 3225 284
rect 3289 220 3305 284
rect 3369 220 3511 284
rect 3575 220 3591 284
rect 3655 220 3671 284
rect 3735 220 3751 284
rect 3815 220 3831 284
rect 3895 220 3911 284
rect 3975 220 4117 284
rect 4181 220 4197 284
rect 4261 220 4277 284
rect 4341 220 4357 284
rect 4421 220 4437 284
rect 4501 220 4517 284
rect 4581 220 4723 284
rect 4787 220 4803 284
rect 4867 220 4883 284
rect 4947 220 4963 284
rect 5027 220 5043 284
rect 5107 220 5123 284
rect 5187 220 5291 284
rect 2801 218 5291 220
rect 5352 284 10266 286
rect 5352 220 5456 284
rect 5520 220 5536 284
rect 5600 220 5616 284
rect 5680 220 5696 284
rect 5760 220 5776 284
rect 5840 220 5856 284
rect 5920 220 6062 284
rect 6126 220 6142 284
rect 6206 220 6222 284
rect 6286 220 6302 284
rect 6366 220 6382 284
rect 6446 220 6462 284
rect 6526 220 6668 284
rect 6732 220 6748 284
rect 6812 220 6828 284
rect 6892 220 6908 284
rect 6972 220 6988 284
rect 7052 220 7068 284
rect 7132 220 7274 284
rect 7338 220 7354 284
rect 7418 220 7434 284
rect 7498 220 7514 284
rect 7578 220 7594 284
rect 7658 220 7674 284
rect 7738 220 7880 284
rect 7944 220 7960 284
rect 8024 220 8040 284
rect 8104 220 8120 284
rect 8184 220 8200 284
rect 8264 220 8280 284
rect 8344 220 8486 284
rect 8550 220 8566 284
rect 8630 220 8646 284
rect 8710 220 8726 284
rect 8790 220 8806 284
rect 8870 220 8886 284
rect 8950 220 9092 284
rect 9156 220 9172 284
rect 9236 220 9252 284
rect 9316 220 9332 284
rect 9396 220 9412 284
rect 9476 220 9492 284
rect 9556 220 9698 284
rect 9762 220 9778 284
rect 9842 220 9858 284
rect 9922 220 9938 284
rect 10002 220 10018 284
rect 10082 220 10098 284
rect 10162 220 10266 284
rect 5352 218 10266 220
rect 10326 284 20088 286
rect 10326 220 10430 284
rect 10494 220 10510 284
rect 10574 220 10590 284
rect 10654 220 10670 284
rect 10734 220 10750 284
rect 10814 220 10830 284
rect 10894 220 11036 284
rect 11100 220 11116 284
rect 11180 220 11196 284
rect 11260 220 11276 284
rect 11340 220 11356 284
rect 11420 220 11436 284
rect 11500 220 11642 284
rect 11706 220 11722 284
rect 11786 220 11802 284
rect 11866 220 11882 284
rect 11946 220 11962 284
rect 12026 220 12042 284
rect 12106 220 12248 284
rect 12312 220 12328 284
rect 12392 220 12408 284
rect 12472 220 12488 284
rect 12552 220 12568 284
rect 12632 220 12648 284
rect 12712 220 12854 284
rect 12918 220 12934 284
rect 12998 220 13014 284
rect 13078 220 13094 284
rect 13158 220 13174 284
rect 13238 220 13254 284
rect 13318 220 13460 284
rect 13524 220 13540 284
rect 13604 220 13620 284
rect 13684 220 13700 284
rect 13764 220 13780 284
rect 13844 220 13860 284
rect 13924 220 14066 284
rect 14130 220 14146 284
rect 14210 220 14226 284
rect 14290 220 14306 284
rect 14370 220 14386 284
rect 14450 220 14466 284
rect 14530 220 14672 284
rect 14736 220 14752 284
rect 14816 220 14832 284
rect 14896 220 14912 284
rect 14976 220 14992 284
rect 15056 220 15072 284
rect 15136 220 15278 284
rect 15342 220 15358 284
rect 15422 220 15438 284
rect 15502 220 15518 284
rect 15582 220 15598 284
rect 15662 220 15678 284
rect 15742 220 15884 284
rect 15948 220 15964 284
rect 16028 220 16044 284
rect 16108 220 16124 284
rect 16188 220 16204 284
rect 16268 220 16284 284
rect 16348 220 16490 284
rect 16554 220 16570 284
rect 16634 220 16650 284
rect 16714 220 16730 284
rect 16794 220 16810 284
rect 16874 220 16890 284
rect 16954 220 17096 284
rect 17160 220 17176 284
rect 17240 220 17256 284
rect 17320 220 17336 284
rect 17400 220 17416 284
rect 17480 220 17496 284
rect 17560 220 17702 284
rect 17766 220 17782 284
rect 17846 220 17862 284
rect 17926 220 17942 284
rect 18006 220 18022 284
rect 18086 220 18102 284
rect 18166 220 18308 284
rect 18372 220 18388 284
rect 18452 220 18468 284
rect 18532 220 18548 284
rect 18612 220 18628 284
rect 18692 220 18708 284
rect 18772 220 18914 284
rect 18978 220 18994 284
rect 19058 220 19074 284
rect 19138 220 19154 284
rect 19218 220 19234 284
rect 19298 220 19314 284
rect 19378 220 19520 284
rect 19584 220 19600 284
rect 19664 220 19680 284
rect 19744 220 19760 284
rect 19824 220 19840 284
rect 19904 220 19920 284
rect 19984 220 20088 284
rect 10326 218 20088 220
rect 20148 284 39606 286
rect 20148 220 20252 284
rect 20316 220 20332 284
rect 20396 220 20412 284
rect 20476 220 20492 284
rect 20556 220 20572 284
rect 20636 220 20652 284
rect 20716 220 20858 284
rect 20922 220 20938 284
rect 21002 220 21018 284
rect 21082 220 21098 284
rect 21162 220 21178 284
rect 21242 220 21258 284
rect 21322 220 21464 284
rect 21528 220 21544 284
rect 21608 220 21624 284
rect 21688 220 21704 284
rect 21768 220 21784 284
rect 21848 220 21864 284
rect 21928 220 22070 284
rect 22134 220 22150 284
rect 22214 220 22230 284
rect 22294 220 22310 284
rect 22374 220 22390 284
rect 22454 220 22470 284
rect 22534 220 22676 284
rect 22740 220 22756 284
rect 22820 220 22836 284
rect 22900 220 22916 284
rect 22980 220 22996 284
rect 23060 220 23076 284
rect 23140 220 23282 284
rect 23346 220 23362 284
rect 23426 220 23442 284
rect 23506 220 23522 284
rect 23586 220 23602 284
rect 23666 220 23682 284
rect 23746 220 23888 284
rect 23952 220 23968 284
rect 24032 220 24048 284
rect 24112 220 24128 284
rect 24192 220 24208 284
rect 24272 220 24288 284
rect 24352 220 24494 284
rect 24558 220 24574 284
rect 24638 220 24654 284
rect 24718 220 24734 284
rect 24798 220 24814 284
rect 24878 220 24894 284
rect 24958 220 25100 284
rect 25164 220 25180 284
rect 25244 220 25260 284
rect 25324 220 25340 284
rect 25404 220 25420 284
rect 25484 220 25500 284
rect 25564 220 25706 284
rect 25770 220 25786 284
rect 25850 220 25866 284
rect 25930 220 25946 284
rect 26010 220 26026 284
rect 26090 220 26106 284
rect 26170 220 26312 284
rect 26376 220 26392 284
rect 26456 220 26472 284
rect 26536 220 26552 284
rect 26616 220 26632 284
rect 26696 220 26712 284
rect 26776 220 26918 284
rect 26982 220 26998 284
rect 27062 220 27078 284
rect 27142 220 27158 284
rect 27222 220 27238 284
rect 27302 220 27318 284
rect 27382 220 27524 284
rect 27588 220 27604 284
rect 27668 220 27684 284
rect 27748 220 27764 284
rect 27828 220 27844 284
rect 27908 220 27924 284
rect 27988 220 28130 284
rect 28194 220 28210 284
rect 28274 220 28290 284
rect 28354 220 28370 284
rect 28434 220 28450 284
rect 28514 220 28530 284
rect 28594 220 28736 284
rect 28800 220 28816 284
rect 28880 220 28896 284
rect 28960 220 28976 284
rect 29040 220 29056 284
rect 29120 220 29136 284
rect 29200 220 29342 284
rect 29406 220 29422 284
rect 29486 220 29502 284
rect 29566 220 29582 284
rect 29646 220 29662 284
rect 29726 220 29742 284
rect 29806 220 29948 284
rect 30012 220 30028 284
rect 30092 220 30108 284
rect 30172 220 30188 284
rect 30252 220 30268 284
rect 30332 220 30348 284
rect 30412 220 30554 284
rect 30618 220 30634 284
rect 30698 220 30714 284
rect 30778 220 30794 284
rect 30858 220 30874 284
rect 30938 220 30954 284
rect 31018 220 31160 284
rect 31224 220 31240 284
rect 31304 220 31320 284
rect 31384 220 31400 284
rect 31464 220 31480 284
rect 31544 220 31560 284
rect 31624 220 31766 284
rect 31830 220 31846 284
rect 31910 220 31926 284
rect 31990 220 32006 284
rect 32070 220 32086 284
rect 32150 220 32166 284
rect 32230 220 32372 284
rect 32436 220 32452 284
rect 32516 220 32532 284
rect 32596 220 32612 284
rect 32676 220 32692 284
rect 32756 220 32772 284
rect 32836 220 32978 284
rect 33042 220 33058 284
rect 33122 220 33138 284
rect 33202 220 33218 284
rect 33282 220 33298 284
rect 33362 220 33378 284
rect 33442 220 33584 284
rect 33648 220 33664 284
rect 33728 220 33744 284
rect 33808 220 33824 284
rect 33888 220 33904 284
rect 33968 220 33984 284
rect 34048 220 34190 284
rect 34254 220 34270 284
rect 34334 220 34350 284
rect 34414 220 34430 284
rect 34494 220 34510 284
rect 34574 220 34590 284
rect 34654 220 34796 284
rect 34860 220 34876 284
rect 34940 220 34956 284
rect 35020 220 35036 284
rect 35100 220 35116 284
rect 35180 220 35196 284
rect 35260 220 35402 284
rect 35466 220 35482 284
rect 35546 220 35562 284
rect 35626 220 35642 284
rect 35706 220 35722 284
rect 35786 220 35802 284
rect 35866 220 36008 284
rect 36072 220 36088 284
rect 36152 220 36168 284
rect 36232 220 36248 284
rect 36312 220 36328 284
rect 36392 220 36408 284
rect 36472 220 36614 284
rect 36678 220 36694 284
rect 36758 220 36774 284
rect 36838 220 36854 284
rect 36918 220 36934 284
rect 36998 220 37014 284
rect 37078 220 37220 284
rect 37284 220 37300 284
rect 37364 220 37380 284
rect 37444 220 37460 284
rect 37524 220 37540 284
rect 37604 220 37620 284
rect 37684 220 37826 284
rect 37890 220 37906 284
rect 37970 220 37986 284
rect 38050 220 38066 284
rect 38130 220 38146 284
rect 38210 220 38226 284
rect 38290 220 38432 284
rect 38496 220 38512 284
rect 38576 220 38592 284
rect 38656 220 38672 284
rect 38736 220 38752 284
rect 38816 220 38832 284
rect 38896 220 39038 284
rect 39102 220 39118 284
rect 39182 220 39198 284
rect 39262 220 39278 284
rect 39342 220 39358 284
rect 39422 220 39438 284
rect 39502 220 39606 284
rect 20148 218 39606 220
<< via3 >>
rect 28951 6051 29015 6055
rect 28951 5995 28955 6051
rect 28955 5995 29011 6051
rect 29011 5995 29015 6051
rect 28951 5991 29015 5995
rect 29758 6054 29822 6058
rect 29758 5998 29762 6054
rect 29762 5998 29818 6054
rect 29818 5998 29822 6054
rect 29758 5994 29822 5998
rect 29147 5419 29211 5423
rect 29147 5363 29151 5419
rect 29151 5363 29207 5419
rect 29207 5363 29211 5419
rect 29147 5359 29211 5363
rect -355 5028 -291 5092
rect -275 5028 -211 5092
rect -195 5028 -131 5092
rect -115 5028 -51 5092
rect -35 5028 29 5092
rect 45 5028 109 5092
rect 459 5028 523 5092
rect 539 5028 603 5092
rect 619 5028 683 5092
rect 699 5028 763 5092
rect 779 5028 843 5092
rect 859 5028 923 5092
rect 1371 5028 1435 5092
rect 1451 5028 1515 5092
rect 1531 5028 1595 5092
rect 1611 5028 1675 5092
rect 1691 5028 1755 5092
rect 1771 5028 1835 5092
rect 1977 5028 2041 5092
rect 2057 5028 2121 5092
rect 2137 5028 2201 5092
rect 2217 5028 2281 5092
rect 2297 5028 2361 5092
rect 2377 5028 2441 5092
rect 2905 5028 2969 5092
rect 2985 5028 3049 5092
rect 3065 5028 3129 5092
rect 3145 5028 3209 5092
rect 3225 5028 3289 5092
rect 3305 5028 3369 5092
rect 3511 5028 3575 5092
rect 3591 5028 3655 5092
rect 3671 5028 3735 5092
rect 3751 5028 3815 5092
rect 3831 5028 3895 5092
rect 3911 5028 3975 5092
rect 4117 5028 4181 5092
rect 4197 5028 4261 5092
rect 4277 5028 4341 5092
rect 4357 5028 4421 5092
rect 4437 5028 4501 5092
rect 4517 5028 4581 5092
rect 4723 5028 4787 5092
rect 4803 5028 4867 5092
rect 4883 5028 4947 5092
rect 4963 5028 5027 5092
rect 5043 5028 5107 5092
rect 5123 5028 5187 5092
rect 5456 5028 5520 5092
rect 5536 5028 5600 5092
rect 5616 5028 5680 5092
rect 5696 5028 5760 5092
rect 5776 5028 5840 5092
rect 5856 5028 5920 5092
rect 6062 5028 6126 5092
rect 6142 5028 6206 5092
rect 6222 5028 6286 5092
rect 6302 5028 6366 5092
rect 6382 5028 6446 5092
rect 6462 5028 6526 5092
rect 6668 5028 6732 5092
rect 6748 5028 6812 5092
rect 6828 5028 6892 5092
rect 6908 5028 6972 5092
rect 6988 5028 7052 5092
rect 7068 5028 7132 5092
rect 7274 5028 7338 5092
rect 7354 5028 7418 5092
rect 7434 5028 7498 5092
rect 7514 5028 7578 5092
rect 7594 5028 7658 5092
rect 7674 5028 7738 5092
rect 7880 5028 7944 5092
rect 7960 5028 8024 5092
rect 8040 5028 8104 5092
rect 8120 5028 8184 5092
rect 8200 5028 8264 5092
rect 8280 5028 8344 5092
rect 8486 5028 8550 5092
rect 8566 5028 8630 5092
rect 8646 5028 8710 5092
rect 8726 5028 8790 5092
rect 8806 5028 8870 5092
rect 8886 5028 8950 5092
rect 9092 5028 9156 5092
rect 9172 5028 9236 5092
rect 9252 5028 9316 5092
rect 9332 5028 9396 5092
rect 9412 5028 9476 5092
rect 9492 5028 9556 5092
rect 9698 5028 9762 5092
rect 9778 5028 9842 5092
rect 9858 5028 9922 5092
rect 9938 5028 10002 5092
rect 10018 5028 10082 5092
rect 10098 5028 10162 5092
rect 10430 5028 10494 5092
rect 10510 5028 10574 5092
rect 10590 5028 10654 5092
rect 10670 5028 10734 5092
rect 10750 5028 10814 5092
rect 10830 5028 10894 5092
rect 11036 5028 11100 5092
rect 11116 5028 11180 5092
rect 11196 5028 11260 5092
rect 11276 5028 11340 5092
rect 11356 5028 11420 5092
rect 11436 5028 11500 5092
rect 11642 5028 11706 5092
rect 11722 5028 11786 5092
rect 11802 5028 11866 5092
rect 11882 5028 11946 5092
rect 11962 5028 12026 5092
rect 12042 5028 12106 5092
rect 12248 5028 12312 5092
rect 12328 5028 12392 5092
rect 12408 5028 12472 5092
rect 12488 5028 12552 5092
rect 12568 5028 12632 5092
rect 12648 5028 12712 5092
rect 12854 5028 12918 5092
rect 12934 5028 12998 5092
rect 13014 5028 13078 5092
rect 13094 5028 13158 5092
rect 13174 5028 13238 5092
rect 13254 5028 13318 5092
rect 13460 5028 13524 5092
rect 13540 5028 13604 5092
rect 13620 5028 13684 5092
rect 13700 5028 13764 5092
rect 13780 5028 13844 5092
rect 13860 5028 13924 5092
rect 14066 5028 14130 5092
rect 14146 5028 14210 5092
rect 14226 5028 14290 5092
rect 14306 5028 14370 5092
rect 14386 5028 14450 5092
rect 14466 5028 14530 5092
rect 14672 5028 14736 5092
rect 14752 5028 14816 5092
rect 14832 5028 14896 5092
rect 14912 5028 14976 5092
rect 14992 5028 15056 5092
rect 15072 5028 15136 5092
rect 15278 5028 15342 5092
rect 15358 5028 15422 5092
rect 15438 5028 15502 5092
rect 15518 5028 15582 5092
rect 15598 5028 15662 5092
rect 15678 5028 15742 5092
rect 15884 5028 15948 5092
rect 15964 5028 16028 5092
rect 16044 5028 16108 5092
rect 16124 5028 16188 5092
rect 16204 5028 16268 5092
rect 16284 5028 16348 5092
rect 16490 5028 16554 5092
rect 16570 5028 16634 5092
rect 16650 5028 16714 5092
rect 16730 5028 16794 5092
rect 16810 5028 16874 5092
rect 16890 5028 16954 5092
rect 17096 5028 17160 5092
rect 17176 5028 17240 5092
rect 17256 5028 17320 5092
rect 17336 5028 17400 5092
rect 17416 5028 17480 5092
rect 17496 5028 17560 5092
rect 17702 5028 17766 5092
rect 17782 5028 17846 5092
rect 17862 5028 17926 5092
rect 17942 5028 18006 5092
rect 18022 5028 18086 5092
rect 18102 5028 18166 5092
rect 18308 5028 18372 5092
rect 18388 5028 18452 5092
rect 18468 5028 18532 5092
rect 18548 5028 18612 5092
rect 18628 5028 18692 5092
rect 18708 5028 18772 5092
rect 18914 5028 18978 5092
rect 18994 5028 19058 5092
rect 19074 5028 19138 5092
rect 19154 5028 19218 5092
rect 19234 5028 19298 5092
rect 19314 5028 19378 5092
rect 19520 5028 19584 5092
rect 19600 5028 19664 5092
rect 19680 5028 19744 5092
rect 19760 5028 19824 5092
rect 19840 5028 19904 5092
rect 19920 5028 19984 5092
rect 20252 5028 20316 5092
rect 20332 5028 20396 5092
rect 20412 5028 20476 5092
rect 20492 5028 20556 5092
rect 20572 5028 20636 5092
rect 20652 5028 20716 5092
rect 20858 5028 20922 5092
rect 20938 5028 21002 5092
rect 21018 5028 21082 5092
rect 21098 5028 21162 5092
rect 21178 5028 21242 5092
rect 21258 5028 21322 5092
rect 21464 5028 21528 5092
rect 21544 5028 21608 5092
rect 21624 5028 21688 5092
rect 21704 5028 21768 5092
rect 21784 5028 21848 5092
rect 21864 5028 21928 5092
rect 22070 5028 22134 5092
rect 22150 5028 22214 5092
rect 22230 5028 22294 5092
rect 22310 5028 22374 5092
rect 22390 5028 22454 5092
rect 22470 5028 22534 5092
rect 22676 5028 22740 5092
rect 22756 5028 22820 5092
rect 22836 5028 22900 5092
rect 22916 5028 22980 5092
rect 22996 5028 23060 5092
rect 23076 5028 23140 5092
rect 23282 5028 23346 5092
rect 23362 5028 23426 5092
rect 23442 5028 23506 5092
rect 23522 5028 23586 5092
rect 23602 5028 23666 5092
rect 23682 5028 23746 5092
rect 23888 5028 23952 5092
rect 23968 5028 24032 5092
rect 24048 5028 24112 5092
rect 24128 5028 24192 5092
rect 24208 5028 24272 5092
rect 24288 5028 24352 5092
rect 24494 5028 24558 5092
rect 24574 5028 24638 5092
rect 24654 5028 24718 5092
rect 24734 5028 24798 5092
rect 24814 5028 24878 5092
rect 24894 5028 24958 5092
rect 25100 5028 25164 5092
rect 25180 5028 25244 5092
rect 25260 5028 25324 5092
rect 25340 5028 25404 5092
rect 25420 5028 25484 5092
rect 25500 5028 25564 5092
rect 25706 5028 25770 5092
rect 25786 5028 25850 5092
rect 25866 5028 25930 5092
rect 25946 5028 26010 5092
rect 26026 5028 26090 5092
rect 26106 5028 26170 5092
rect 26312 5028 26376 5092
rect 26392 5028 26456 5092
rect 26472 5028 26536 5092
rect 26552 5028 26616 5092
rect 26632 5028 26696 5092
rect 26712 5028 26776 5092
rect 26918 5028 26982 5092
rect 26998 5028 27062 5092
rect 27078 5028 27142 5092
rect 27158 5028 27222 5092
rect 27238 5028 27302 5092
rect 27318 5028 27382 5092
rect 27524 5028 27588 5092
rect 27604 5028 27668 5092
rect 27684 5028 27748 5092
rect 27764 5028 27828 5092
rect 27844 5028 27908 5092
rect 27924 5028 27988 5092
rect 28130 5028 28194 5092
rect 28210 5028 28274 5092
rect 28290 5028 28354 5092
rect 28370 5028 28434 5092
rect 28450 5028 28514 5092
rect 28530 5028 28594 5092
rect 28736 5028 28800 5092
rect 28816 5028 28880 5092
rect 28896 5028 28960 5092
rect 28976 5028 29040 5092
rect 29056 5028 29120 5092
rect 29136 5028 29200 5092
rect 29342 5028 29406 5092
rect 29422 5028 29486 5092
rect 29502 5028 29566 5092
rect 29582 5028 29646 5092
rect 29662 5028 29726 5092
rect 29742 5028 29806 5092
rect 29948 5028 30012 5092
rect 30028 5028 30092 5092
rect 30108 5028 30172 5092
rect 30188 5028 30252 5092
rect 30268 5028 30332 5092
rect 30348 5028 30412 5092
rect 30554 5028 30618 5092
rect 30634 5028 30698 5092
rect 30714 5028 30778 5092
rect 30794 5028 30858 5092
rect 30874 5028 30938 5092
rect 30954 5028 31018 5092
rect 31160 5028 31224 5092
rect 31240 5028 31304 5092
rect 31320 5028 31384 5092
rect 31400 5028 31464 5092
rect 31480 5028 31544 5092
rect 31560 5028 31624 5092
rect 31766 5028 31830 5092
rect 31846 5028 31910 5092
rect 31926 5028 31990 5092
rect 32006 5028 32070 5092
rect 32086 5028 32150 5092
rect 32166 5028 32230 5092
rect 32372 5028 32436 5092
rect 32452 5028 32516 5092
rect 32532 5028 32596 5092
rect 32612 5028 32676 5092
rect 32692 5028 32756 5092
rect 32772 5028 32836 5092
rect 32978 5028 33042 5092
rect 33058 5028 33122 5092
rect 33138 5028 33202 5092
rect 33218 5028 33282 5092
rect 33298 5028 33362 5092
rect 33378 5028 33442 5092
rect 33584 5028 33648 5092
rect 33664 5028 33728 5092
rect 33744 5028 33808 5092
rect 33824 5028 33888 5092
rect 33904 5028 33968 5092
rect 33984 5028 34048 5092
rect 34190 5028 34254 5092
rect 34270 5028 34334 5092
rect 34350 5028 34414 5092
rect 34430 5028 34494 5092
rect 34510 5028 34574 5092
rect 34590 5028 34654 5092
rect 34796 5028 34860 5092
rect 34876 5028 34940 5092
rect 34956 5028 35020 5092
rect 35036 5028 35100 5092
rect 35116 5028 35180 5092
rect 35196 5028 35260 5092
rect 35402 5028 35466 5092
rect 35482 5028 35546 5092
rect 35562 5028 35626 5092
rect 35642 5028 35706 5092
rect 35722 5028 35786 5092
rect 35802 5028 35866 5092
rect 36008 5028 36072 5092
rect 36088 5028 36152 5092
rect 36168 5028 36232 5092
rect 36248 5028 36312 5092
rect 36328 5028 36392 5092
rect 36408 5028 36472 5092
rect 36614 5028 36678 5092
rect 36694 5028 36758 5092
rect 36774 5028 36838 5092
rect 36854 5028 36918 5092
rect 36934 5028 36998 5092
rect 37014 5028 37078 5092
rect 37220 5028 37284 5092
rect 37300 5028 37364 5092
rect 37380 5028 37444 5092
rect 37460 5028 37524 5092
rect 37540 5028 37604 5092
rect 37620 5028 37684 5092
rect 37826 5028 37890 5092
rect 37906 5028 37970 5092
rect 37986 5028 38050 5092
rect 38066 5028 38130 5092
rect 38146 5028 38210 5092
rect 38226 5028 38290 5092
rect 38432 5028 38496 5092
rect 38512 5028 38576 5092
rect 38592 5028 38656 5092
rect 38672 5028 38736 5092
rect 38752 5028 38816 5092
rect 38832 5028 38896 5092
rect 39038 5028 39102 5092
rect 39118 5028 39182 5092
rect 39198 5028 39262 5092
rect 39278 5028 39342 5092
rect 39358 5028 39422 5092
rect 39438 5028 39502 5092
rect -458 4808 -394 4872
rect -458 4728 -394 4792
rect -458 4648 -394 4712
rect -458 4568 -394 4632
rect -458 4488 -394 4552
rect -458 4408 -394 4472
rect -458 4328 -394 4392
rect -458 4248 -394 4312
rect -458 4168 -394 4232
rect -458 4088 -394 4152
rect 148 4808 212 4872
rect 148 4728 212 4792
rect 148 4648 212 4712
rect 148 4568 212 4632
rect 148 4488 212 4552
rect 148 4408 212 4472
rect 148 4328 212 4392
rect 148 4248 212 4312
rect 148 4168 212 4232
rect 148 4088 212 4152
rect 356 4808 420 4872
rect 356 4728 420 4792
rect 356 4648 420 4712
rect 356 4568 420 4632
rect 356 4488 420 4552
rect 356 4408 420 4472
rect 356 4328 420 4392
rect 356 4248 420 4312
rect 356 4168 420 4232
rect 356 4088 420 4152
rect 962 4808 1026 4872
rect 962 4728 1026 4792
rect 962 4648 1026 4712
rect 962 4568 1026 4632
rect 962 4488 1026 4552
rect 962 4408 1026 4472
rect 962 4328 1026 4392
rect 962 4248 1026 4312
rect 962 4168 1026 4232
rect 962 4088 1026 4152
rect -355 3868 -291 3932
rect -275 3868 -211 3932
rect -195 3868 -131 3932
rect -115 3868 -51 3932
rect -35 3868 29 3932
rect 45 3868 109 3932
rect 459 3868 523 3932
rect 539 3868 603 3932
rect 619 3868 683 3932
rect 699 3868 763 3932
rect 779 3868 843 3932
rect 859 3868 923 3932
rect -458 3648 -394 3712
rect -458 3568 -394 3632
rect -458 3488 -394 3552
rect -458 3408 -394 3472
rect -458 3328 -394 3392
rect -458 3248 -394 3312
rect -458 3168 -394 3232
rect -458 3088 -394 3152
rect -458 3008 -394 3072
rect -458 2928 -394 2992
rect 148 3648 212 3712
rect 148 3568 212 3632
rect 148 3488 212 3552
rect 148 3408 212 3472
rect 148 3328 212 3392
rect 148 3248 212 3312
rect 148 3168 212 3232
rect 148 3088 212 3152
rect 148 3008 212 3072
rect 148 2928 212 2992
rect 356 3648 420 3712
rect 356 3568 420 3632
rect 356 3488 420 3552
rect 356 3408 420 3472
rect 356 3328 420 3392
rect 356 3248 420 3312
rect 356 3168 420 3232
rect 356 3088 420 3152
rect 356 3020 360 3072
rect 360 3020 416 3072
rect 416 3020 420 3072
rect 356 3008 420 3020
rect 356 2928 420 2992
rect 962 3648 1026 3712
rect 962 3568 1026 3632
rect 962 3488 1026 3552
rect 962 3408 1026 3472
rect 962 3328 1026 3392
rect 962 3248 1026 3312
rect 962 3168 1026 3232
rect 962 3088 1026 3152
rect 962 3008 1026 3072
rect 962 2928 1026 2992
rect 1268 4808 1332 4872
rect 1268 4728 1332 4792
rect 1268 4648 1332 4712
rect 1268 4568 1332 4632
rect 1268 4488 1332 4552
rect 1268 4408 1332 4472
rect 1268 4328 1332 4392
rect 1268 4248 1332 4312
rect 1268 4168 1332 4232
rect 1268 4088 1332 4152
rect 1874 4808 1938 4872
rect 1874 4728 1938 4792
rect 1874 4648 1938 4712
rect 1874 4568 1938 4632
rect 1874 4488 1938 4552
rect 1874 4408 1938 4472
rect 1874 4328 1938 4392
rect 1874 4248 1938 4312
rect 1874 4168 1938 4232
rect 1874 4088 1938 4152
rect 2480 4808 2544 4872
rect 2480 4728 2544 4792
rect 2480 4648 2544 4712
rect 2480 4568 2544 4632
rect 2480 4488 2544 4552
rect 2480 4408 2544 4472
rect 2480 4328 2544 4392
rect 2480 4248 2544 4312
rect 2480 4168 2544 4232
rect 2480 4088 2544 4152
rect 1371 3868 1435 3932
rect 1451 3868 1515 3932
rect 1531 3868 1595 3932
rect 1611 3868 1675 3932
rect 1691 3868 1755 3932
rect 1771 3868 1835 3932
rect 1977 3868 2041 3932
rect 2057 3868 2121 3932
rect 2137 3868 2201 3932
rect 2217 3868 2281 3932
rect 2297 3868 2361 3932
rect 2377 3868 2441 3932
rect 1268 3648 1332 3712
rect 1268 3568 1332 3632
rect 1268 3488 1332 3552
rect 1268 3408 1332 3472
rect 1268 3328 1332 3392
rect 1268 3248 1332 3312
rect 1268 3168 1332 3232
rect 1268 3145 1332 3152
rect 1268 3089 1272 3145
rect 1272 3089 1328 3145
rect 1328 3089 1332 3145
rect 1268 3088 1332 3089
rect 1268 3008 1332 3072
rect 1268 2928 1332 2992
rect 1874 3648 1938 3712
rect 1874 3568 1938 3632
rect 1874 3488 1938 3552
rect 1874 3408 1938 3472
rect 1874 3328 1938 3392
rect 1874 3248 1938 3312
rect 1874 3168 1938 3232
rect 1874 3088 1938 3152
rect 1874 3008 1938 3072
rect 1874 2928 1938 2992
rect 2480 3648 2544 3712
rect 2480 3568 2544 3632
rect 2480 3488 2544 3552
rect 2480 3408 2544 3472
rect 2480 3328 2544 3392
rect 2480 3248 2544 3312
rect 2480 3168 2544 3232
rect 2480 3088 2544 3152
rect 2480 3008 2544 3072
rect 2480 2928 2544 2992
rect 2802 4808 2866 4872
rect 2802 4728 2866 4792
rect 2802 4648 2866 4712
rect 2802 4568 2866 4632
rect 2802 4488 2866 4552
rect 2802 4408 2866 4472
rect 2802 4328 2866 4392
rect 2802 4248 2866 4312
rect 2802 4168 2866 4232
rect 2802 4088 2866 4152
rect 3408 4808 3472 4872
rect 3408 4728 3472 4792
rect 3408 4648 3472 4712
rect 3408 4568 3472 4632
rect 3408 4488 3472 4552
rect 3408 4408 3472 4472
rect 3408 4328 3472 4392
rect 3408 4248 3472 4312
rect 3408 4168 3472 4232
rect 3408 4088 3472 4152
rect 4014 4808 4078 4872
rect 4014 4728 4078 4792
rect 4014 4648 4078 4712
rect 4014 4568 4078 4632
rect 4014 4488 4078 4552
rect 4014 4408 4078 4472
rect 4014 4328 4078 4392
rect 4014 4248 4078 4312
rect 4014 4168 4078 4232
rect 4014 4088 4078 4152
rect 4620 4808 4684 4872
rect 4620 4728 4684 4792
rect 4620 4648 4684 4712
rect 4620 4568 4684 4632
rect 4620 4488 4684 4552
rect 4620 4408 4684 4472
rect 4620 4328 4684 4392
rect 4620 4248 4684 4312
rect 4620 4168 4684 4232
rect 4620 4088 4684 4152
rect 5226 4808 5290 4872
rect 5226 4728 5290 4792
rect 5226 4648 5290 4712
rect 5226 4568 5290 4632
rect 5226 4488 5290 4552
rect 5226 4408 5290 4472
rect 5226 4328 5290 4392
rect 5226 4248 5290 4312
rect 5226 4168 5290 4232
rect 5226 4088 5290 4152
rect 2905 3868 2969 3932
rect 2985 3868 3049 3932
rect 3065 3868 3129 3932
rect 3145 3868 3209 3932
rect 3225 3868 3289 3932
rect 3305 3868 3369 3932
rect 3511 3868 3575 3932
rect 3591 3868 3655 3932
rect 3671 3868 3735 3932
rect 3751 3868 3815 3932
rect 3831 3868 3895 3932
rect 3911 3868 3975 3932
rect 4117 3868 4181 3932
rect 4197 3868 4261 3932
rect 4277 3868 4341 3932
rect 4357 3868 4421 3932
rect 4437 3868 4501 3932
rect 4517 3868 4581 3932
rect 4723 3868 4787 3932
rect 4803 3868 4867 3932
rect 4883 3868 4947 3932
rect 4963 3868 5027 3932
rect 5043 3868 5107 3932
rect 5123 3868 5187 3932
rect 2802 3648 2866 3712
rect 2802 3568 2866 3632
rect 2802 3488 2866 3552
rect 2802 3408 2866 3472
rect 2802 3328 2866 3392
rect 2802 3248 2866 3312
rect 2802 3168 2866 3232
rect 2802 3133 2866 3152
rect 2802 3088 2806 3133
rect 2806 3088 2862 3133
rect 2862 3088 2866 3133
rect 2802 3008 2866 3072
rect 2802 2928 2866 2992
rect 3408 3648 3472 3712
rect 3408 3568 3472 3632
rect 3408 3488 3472 3552
rect 3408 3408 3472 3472
rect 3408 3328 3472 3392
rect 3408 3248 3472 3312
rect 3408 3168 3472 3232
rect 3408 3088 3472 3152
rect 3408 3008 3472 3072
rect 3408 2928 3472 2992
rect 4014 3648 4078 3712
rect 4014 3568 4078 3632
rect 4014 3488 4078 3552
rect 4014 3408 4078 3472
rect 4014 3328 4078 3392
rect 4014 3248 4078 3312
rect 4014 3168 4078 3232
rect 4014 3088 4078 3152
rect 4014 3008 4078 3072
rect 4014 2928 4078 2992
rect 4620 3648 4684 3712
rect 4620 3568 4684 3632
rect 4620 3488 4684 3552
rect 4620 3408 4684 3472
rect 4620 3328 4684 3392
rect 4620 3248 4684 3312
rect 4620 3168 4684 3232
rect 4620 3088 4684 3152
rect 4620 3008 4684 3072
rect 4620 2928 4684 2992
rect 5226 3648 5290 3712
rect 5226 3568 5290 3632
rect 5226 3488 5290 3552
rect 5226 3408 5290 3472
rect 5226 3328 5290 3392
rect 5226 3248 5290 3312
rect 5226 3168 5290 3232
rect 5226 3088 5290 3152
rect 5226 3008 5290 3072
rect 5226 2928 5290 2992
rect 5353 4808 5417 4872
rect 5353 4728 5417 4792
rect 5353 4648 5417 4712
rect 5353 4568 5417 4632
rect 5353 4488 5417 4552
rect 5353 4408 5417 4472
rect 5353 4328 5417 4392
rect 5353 4248 5417 4312
rect 5353 4168 5417 4232
rect 5353 4088 5417 4152
rect 5959 4808 6023 4872
rect 5959 4728 6023 4792
rect 5959 4648 6023 4712
rect 5959 4568 6023 4632
rect 5959 4488 6023 4552
rect 5959 4408 6023 4472
rect 5959 4328 6023 4392
rect 5959 4248 6023 4312
rect 5959 4168 6023 4232
rect 5959 4088 6023 4152
rect 6565 4808 6629 4872
rect 6565 4728 6629 4792
rect 6565 4648 6629 4712
rect 6565 4568 6629 4632
rect 6565 4488 6629 4552
rect 6565 4408 6629 4472
rect 6565 4328 6629 4392
rect 6565 4248 6629 4312
rect 6565 4168 6629 4232
rect 6565 4088 6629 4152
rect 7171 4808 7235 4872
rect 7171 4728 7235 4792
rect 7171 4648 7235 4712
rect 7171 4568 7235 4632
rect 7171 4488 7235 4552
rect 7171 4408 7235 4472
rect 7171 4328 7235 4392
rect 7171 4248 7235 4312
rect 7171 4168 7235 4232
rect 7171 4088 7235 4152
rect 7777 4808 7841 4872
rect 7777 4728 7841 4792
rect 7777 4648 7841 4712
rect 7777 4568 7841 4632
rect 7777 4488 7841 4552
rect 7777 4408 7841 4472
rect 7777 4328 7841 4392
rect 7777 4248 7841 4312
rect 7777 4168 7841 4232
rect 7777 4088 7841 4152
rect 8383 4808 8447 4872
rect 8383 4728 8447 4792
rect 8383 4648 8447 4712
rect 8383 4568 8447 4632
rect 8383 4488 8447 4552
rect 8383 4408 8447 4472
rect 8383 4328 8447 4392
rect 8383 4248 8447 4312
rect 8383 4168 8447 4232
rect 8383 4088 8447 4152
rect 8989 4808 9053 4872
rect 8989 4728 9053 4792
rect 8989 4648 9053 4712
rect 8989 4568 9053 4632
rect 8989 4488 9053 4552
rect 8989 4408 9053 4472
rect 8989 4328 9053 4392
rect 8989 4248 9053 4312
rect 8989 4168 9053 4232
rect 8989 4088 9053 4152
rect 9595 4808 9659 4872
rect 9595 4728 9659 4792
rect 9595 4648 9659 4712
rect 9595 4568 9659 4632
rect 9595 4488 9659 4552
rect 9595 4408 9659 4472
rect 9595 4328 9659 4392
rect 9595 4248 9659 4312
rect 9595 4168 9659 4232
rect 9595 4088 9659 4152
rect 10201 4808 10265 4872
rect 10201 4728 10265 4792
rect 10201 4648 10265 4712
rect 10201 4568 10265 4632
rect 10201 4488 10265 4552
rect 10201 4408 10265 4472
rect 10201 4328 10265 4392
rect 10201 4248 10265 4312
rect 10201 4168 10265 4232
rect 10201 4088 10265 4152
rect 5456 3868 5520 3932
rect 5536 3868 5600 3932
rect 5616 3868 5680 3932
rect 5696 3868 5760 3932
rect 5776 3868 5840 3932
rect 5856 3868 5920 3932
rect 6062 3868 6126 3932
rect 6142 3868 6206 3932
rect 6222 3868 6286 3932
rect 6302 3868 6366 3932
rect 6382 3868 6446 3932
rect 6462 3868 6526 3932
rect 6668 3868 6732 3932
rect 6748 3868 6812 3932
rect 6828 3868 6892 3932
rect 6908 3868 6972 3932
rect 6988 3868 7052 3932
rect 7068 3868 7132 3932
rect 7274 3868 7338 3932
rect 7354 3868 7418 3932
rect 7434 3868 7498 3932
rect 7514 3868 7578 3932
rect 7594 3868 7658 3932
rect 7674 3868 7738 3932
rect 7880 3868 7944 3932
rect 7960 3868 8024 3932
rect 8040 3868 8104 3932
rect 8120 3868 8184 3932
rect 8200 3868 8264 3932
rect 8280 3868 8344 3932
rect 8486 3868 8550 3932
rect 8566 3868 8630 3932
rect 8646 3868 8710 3932
rect 8726 3868 8790 3932
rect 8806 3868 8870 3932
rect 8886 3868 8950 3932
rect 9092 3868 9156 3932
rect 9172 3868 9236 3932
rect 9252 3868 9316 3932
rect 9332 3868 9396 3932
rect 9412 3868 9476 3932
rect 9492 3868 9556 3932
rect 9698 3868 9762 3932
rect 9778 3868 9842 3932
rect 9858 3868 9922 3932
rect 9938 3868 10002 3932
rect 10018 3868 10082 3932
rect 10098 3868 10162 3932
rect 5353 3648 5417 3712
rect 5353 3568 5417 3632
rect 5353 3488 5417 3552
rect 5353 3408 5417 3472
rect 5353 3328 5417 3392
rect 5353 3248 5417 3312
rect 5353 3168 5417 3232
rect 5353 3109 5357 3152
rect 5357 3109 5413 3152
rect 5413 3109 5417 3152
rect 5353 3088 5417 3109
rect 5353 3008 5417 3072
rect 5353 2928 5417 2992
rect 5959 3648 6023 3712
rect 5959 3568 6023 3632
rect 5959 3488 6023 3552
rect 5959 3408 6023 3472
rect 5959 3328 6023 3392
rect 5959 3248 6023 3312
rect 5959 3168 6023 3232
rect 5959 3088 6023 3152
rect 5959 3008 6023 3072
rect 5959 2928 6023 2992
rect 6565 3648 6629 3712
rect 6565 3568 6629 3632
rect 6565 3488 6629 3552
rect 6565 3408 6629 3472
rect 6565 3328 6629 3392
rect 6565 3248 6629 3312
rect 6565 3168 6629 3232
rect 6565 3088 6629 3152
rect 6565 3008 6629 3072
rect 6565 2928 6629 2992
rect 7171 3648 7235 3712
rect 7171 3568 7235 3632
rect 7171 3488 7235 3552
rect 7171 3408 7235 3472
rect 7171 3328 7235 3392
rect 7171 3248 7235 3312
rect 7171 3168 7235 3232
rect 7171 3088 7235 3152
rect 7171 3008 7235 3072
rect 7171 2928 7235 2992
rect 7777 3648 7841 3712
rect 7777 3568 7841 3632
rect 7777 3488 7841 3552
rect 7777 3408 7841 3472
rect 7777 3328 7841 3392
rect 7777 3248 7841 3312
rect 7777 3168 7841 3232
rect 7777 3088 7841 3152
rect 7777 3008 7841 3072
rect 7777 2928 7841 2992
rect 8383 3648 8447 3712
rect 8383 3568 8447 3632
rect 8383 3488 8447 3552
rect 8383 3408 8447 3472
rect 8383 3328 8447 3392
rect 8383 3248 8447 3312
rect 8383 3168 8447 3232
rect 8383 3088 8447 3152
rect 8383 3008 8447 3072
rect 8383 2928 8447 2992
rect 8989 3648 9053 3712
rect 8989 3568 9053 3632
rect 8989 3488 9053 3552
rect 8989 3408 9053 3472
rect 8989 3328 9053 3392
rect 8989 3248 9053 3312
rect 8989 3168 9053 3232
rect 8989 3088 9053 3152
rect 8989 3008 9053 3072
rect 8989 2928 9053 2992
rect 9595 3648 9659 3712
rect 9595 3568 9659 3632
rect 9595 3488 9659 3552
rect 9595 3408 9659 3472
rect 9595 3328 9659 3392
rect 9595 3248 9659 3312
rect 9595 3168 9659 3232
rect 9595 3088 9659 3152
rect 9595 3008 9659 3072
rect 9595 2928 9659 2992
rect 10201 3648 10265 3712
rect 10201 3568 10265 3632
rect 10201 3488 10265 3552
rect 10201 3408 10265 3472
rect 10201 3328 10265 3392
rect 10201 3248 10265 3312
rect 10201 3168 10265 3232
rect 10201 3088 10265 3152
rect 10201 3008 10265 3072
rect 10201 2928 10265 2992
rect 10327 4808 10391 4872
rect 10327 4728 10391 4792
rect 10327 4648 10391 4712
rect 10327 4568 10391 4632
rect 10327 4488 10391 4552
rect 10327 4408 10391 4472
rect 10327 4328 10391 4392
rect 10327 4248 10391 4312
rect 10327 4168 10391 4232
rect 10327 4088 10391 4152
rect 10933 4808 10997 4872
rect 10933 4728 10997 4792
rect 10933 4648 10997 4712
rect 10933 4568 10997 4632
rect 10933 4488 10997 4552
rect 10933 4408 10997 4472
rect 10933 4328 10997 4392
rect 10933 4248 10997 4312
rect 10933 4168 10997 4232
rect 10933 4088 10997 4152
rect 11539 4808 11603 4872
rect 11539 4728 11603 4792
rect 11539 4648 11603 4712
rect 11539 4568 11603 4632
rect 11539 4488 11603 4552
rect 11539 4408 11603 4472
rect 11539 4328 11603 4392
rect 11539 4248 11603 4312
rect 11539 4168 11603 4232
rect 11539 4088 11603 4152
rect 12145 4808 12209 4872
rect 12145 4728 12209 4792
rect 12145 4648 12209 4712
rect 12145 4568 12209 4632
rect 12145 4488 12209 4552
rect 12145 4408 12209 4472
rect 12145 4328 12209 4392
rect 12145 4248 12209 4312
rect 12145 4168 12209 4232
rect 12145 4088 12209 4152
rect 12751 4808 12815 4872
rect 12751 4728 12815 4792
rect 12751 4648 12815 4712
rect 12751 4568 12815 4632
rect 12751 4488 12815 4552
rect 12751 4408 12815 4472
rect 12751 4328 12815 4392
rect 12751 4248 12815 4312
rect 12751 4168 12815 4232
rect 12751 4088 12815 4152
rect 13357 4808 13421 4872
rect 13357 4728 13421 4792
rect 13357 4648 13421 4712
rect 13357 4568 13421 4632
rect 13357 4488 13421 4552
rect 13357 4408 13421 4472
rect 13357 4328 13421 4392
rect 13357 4248 13421 4312
rect 13357 4168 13421 4232
rect 13357 4088 13421 4152
rect 13963 4808 14027 4872
rect 13963 4728 14027 4792
rect 13963 4648 14027 4712
rect 13963 4568 14027 4632
rect 13963 4488 14027 4552
rect 13963 4408 14027 4472
rect 13963 4328 14027 4392
rect 13963 4248 14027 4312
rect 13963 4168 14027 4232
rect 13963 4088 14027 4152
rect 14569 4808 14633 4872
rect 14569 4728 14633 4792
rect 14569 4648 14633 4712
rect 14569 4568 14633 4632
rect 14569 4488 14633 4552
rect 14569 4408 14633 4472
rect 14569 4328 14633 4392
rect 14569 4248 14633 4312
rect 14569 4168 14633 4232
rect 14569 4088 14633 4152
rect 15175 4808 15239 4872
rect 15175 4728 15239 4792
rect 15175 4648 15239 4712
rect 15175 4568 15239 4632
rect 15175 4488 15239 4552
rect 15175 4408 15239 4472
rect 15175 4328 15239 4392
rect 15175 4248 15239 4312
rect 15175 4168 15239 4232
rect 15175 4088 15239 4152
rect 15781 4808 15845 4872
rect 15781 4728 15845 4792
rect 15781 4648 15845 4712
rect 15781 4568 15845 4632
rect 15781 4488 15845 4552
rect 15781 4408 15845 4472
rect 15781 4328 15845 4392
rect 15781 4248 15845 4312
rect 15781 4168 15845 4232
rect 15781 4088 15845 4152
rect 16387 4808 16451 4872
rect 16387 4728 16451 4792
rect 16387 4648 16451 4712
rect 16387 4568 16451 4632
rect 16387 4488 16451 4552
rect 16387 4408 16451 4472
rect 16387 4328 16451 4392
rect 16387 4248 16451 4312
rect 16387 4168 16451 4232
rect 16387 4088 16451 4152
rect 16993 4808 17057 4872
rect 16993 4728 17057 4792
rect 16993 4648 17057 4712
rect 16993 4568 17057 4632
rect 16993 4488 17057 4552
rect 16993 4408 17057 4472
rect 16993 4328 17057 4392
rect 16993 4248 17057 4312
rect 16993 4168 17057 4232
rect 16993 4088 17057 4152
rect 17599 4808 17663 4872
rect 17599 4728 17663 4792
rect 17599 4648 17663 4712
rect 17599 4568 17663 4632
rect 17599 4488 17663 4552
rect 17599 4408 17663 4472
rect 17599 4328 17663 4392
rect 17599 4248 17663 4312
rect 17599 4168 17663 4232
rect 17599 4088 17663 4152
rect 18205 4808 18269 4872
rect 18205 4728 18269 4792
rect 18205 4648 18269 4712
rect 18205 4568 18269 4632
rect 18205 4488 18269 4552
rect 18205 4408 18269 4472
rect 18205 4328 18269 4392
rect 18205 4248 18269 4312
rect 18205 4168 18269 4232
rect 18205 4088 18269 4152
rect 18811 4808 18875 4872
rect 18811 4728 18875 4792
rect 18811 4648 18875 4712
rect 18811 4568 18875 4632
rect 18811 4488 18875 4552
rect 18811 4408 18875 4472
rect 18811 4328 18875 4392
rect 18811 4248 18875 4312
rect 18811 4168 18875 4232
rect 18811 4088 18875 4152
rect 19417 4808 19481 4872
rect 19417 4728 19481 4792
rect 19417 4648 19481 4712
rect 19417 4568 19481 4632
rect 19417 4488 19481 4552
rect 19417 4408 19481 4472
rect 19417 4328 19481 4392
rect 19417 4248 19481 4312
rect 19417 4168 19481 4232
rect 19417 4088 19481 4152
rect 20023 4808 20087 4872
rect 20023 4728 20087 4792
rect 20023 4648 20087 4712
rect 20023 4568 20087 4632
rect 20023 4488 20087 4552
rect 20023 4408 20087 4472
rect 20023 4328 20087 4392
rect 20023 4248 20087 4312
rect 20023 4168 20087 4232
rect 20023 4088 20087 4152
rect 10430 3868 10494 3932
rect 10510 3868 10574 3932
rect 10590 3868 10654 3932
rect 10670 3868 10734 3932
rect 10750 3868 10814 3932
rect 10830 3868 10894 3932
rect 11036 3868 11100 3932
rect 11116 3868 11180 3932
rect 11196 3868 11260 3932
rect 11276 3868 11340 3932
rect 11356 3868 11420 3932
rect 11436 3868 11500 3932
rect 11642 3868 11706 3932
rect 11722 3868 11786 3932
rect 11802 3868 11866 3932
rect 11882 3868 11946 3932
rect 11962 3868 12026 3932
rect 12042 3868 12106 3932
rect 12248 3868 12312 3932
rect 12328 3868 12392 3932
rect 12408 3868 12472 3932
rect 12488 3868 12552 3932
rect 12568 3868 12632 3932
rect 12648 3868 12712 3932
rect 12854 3868 12918 3932
rect 12934 3868 12998 3932
rect 13014 3868 13078 3932
rect 13094 3868 13158 3932
rect 13174 3868 13238 3932
rect 13254 3868 13318 3932
rect 13460 3868 13524 3932
rect 13540 3868 13604 3932
rect 13620 3868 13684 3932
rect 13700 3868 13764 3932
rect 13780 3868 13844 3932
rect 13860 3868 13924 3932
rect 14066 3868 14130 3932
rect 14146 3868 14210 3932
rect 14226 3868 14290 3932
rect 14306 3868 14370 3932
rect 14386 3868 14450 3932
rect 14466 3868 14530 3932
rect 14672 3868 14736 3932
rect 14752 3868 14816 3932
rect 14832 3868 14896 3932
rect 14912 3868 14976 3932
rect 14992 3868 15056 3932
rect 15072 3868 15136 3932
rect 15278 3868 15342 3932
rect 15358 3868 15422 3932
rect 15438 3868 15502 3932
rect 15518 3868 15582 3932
rect 15598 3868 15662 3932
rect 15678 3868 15742 3932
rect 15884 3868 15948 3932
rect 15964 3868 16028 3932
rect 16044 3868 16108 3932
rect 16124 3868 16188 3932
rect 16204 3868 16268 3932
rect 16284 3868 16348 3932
rect 16490 3868 16554 3932
rect 16570 3868 16634 3932
rect 16650 3868 16714 3932
rect 16730 3868 16794 3932
rect 16810 3868 16874 3932
rect 16890 3868 16954 3932
rect 17096 3868 17160 3932
rect 17176 3868 17240 3932
rect 17256 3868 17320 3932
rect 17336 3868 17400 3932
rect 17416 3868 17480 3932
rect 17496 3868 17560 3932
rect 17702 3868 17766 3932
rect 17782 3868 17846 3932
rect 17862 3868 17926 3932
rect 17942 3868 18006 3932
rect 18022 3868 18086 3932
rect 18102 3868 18166 3932
rect 18308 3868 18372 3932
rect 18388 3868 18452 3932
rect 18468 3868 18532 3932
rect 18548 3868 18612 3932
rect 18628 3868 18692 3932
rect 18708 3868 18772 3932
rect 18914 3868 18978 3932
rect 18994 3868 19058 3932
rect 19074 3868 19138 3932
rect 19154 3868 19218 3932
rect 19234 3868 19298 3932
rect 19314 3868 19378 3932
rect 19520 3868 19584 3932
rect 19600 3868 19664 3932
rect 19680 3868 19744 3932
rect 19760 3868 19824 3932
rect 19840 3868 19904 3932
rect 19920 3868 19984 3932
rect 10327 3648 10391 3712
rect 10327 3568 10391 3632
rect 10327 3488 10391 3552
rect 10327 3408 10391 3472
rect 10327 3328 10391 3392
rect 10327 3273 10391 3312
rect 10327 3248 10331 3273
rect 10331 3248 10387 3273
rect 10387 3248 10391 3273
rect 10327 3217 10331 3232
rect 10331 3217 10387 3232
rect 10387 3217 10391 3232
rect 10327 3168 10391 3217
rect 10327 3088 10391 3152
rect 10327 3008 10391 3072
rect 10327 2928 10391 2992
rect 10933 3648 10997 3712
rect 10933 3568 10997 3632
rect 10933 3488 10997 3552
rect 10933 3408 10997 3472
rect 10933 3328 10997 3392
rect 10933 3248 10997 3312
rect 10933 3168 10997 3232
rect 10933 3088 10997 3152
rect 10933 3008 10997 3072
rect 10933 2928 10997 2992
rect 11539 3648 11603 3712
rect 11539 3568 11603 3632
rect 11539 3488 11603 3552
rect 11539 3408 11603 3472
rect 11539 3328 11603 3392
rect 11539 3248 11603 3312
rect 11539 3168 11603 3232
rect 11539 3088 11603 3152
rect 11539 3008 11603 3072
rect 11539 2928 11603 2992
rect 12145 3648 12209 3712
rect 12145 3568 12209 3632
rect 12145 3488 12209 3552
rect 12145 3408 12209 3472
rect 12145 3328 12209 3392
rect 12145 3248 12209 3312
rect 12145 3168 12209 3232
rect 12145 3088 12209 3152
rect 12145 3008 12209 3072
rect 12145 2928 12209 2992
rect 12751 3648 12815 3712
rect 12751 3568 12815 3632
rect 12751 3488 12815 3552
rect 12751 3408 12815 3472
rect 12751 3328 12815 3392
rect 12751 3248 12815 3312
rect 12751 3168 12815 3232
rect 12751 3088 12815 3152
rect 12751 3008 12815 3072
rect 12751 2928 12815 2992
rect 13357 3648 13421 3712
rect 13357 3568 13421 3632
rect 13357 3488 13421 3552
rect 13357 3408 13421 3472
rect 13357 3328 13421 3392
rect 13357 3248 13421 3312
rect 13357 3168 13421 3232
rect 13357 3088 13421 3152
rect 13357 3008 13421 3072
rect 13357 2928 13421 2992
rect 13963 3648 14027 3712
rect 13963 3568 14027 3632
rect 13963 3488 14027 3552
rect 13963 3408 14027 3472
rect 13963 3328 14027 3392
rect 13963 3248 14027 3312
rect 13963 3168 14027 3232
rect 13963 3088 14027 3152
rect 13963 3008 14027 3072
rect 13963 2928 14027 2992
rect 14569 3648 14633 3712
rect 14569 3568 14633 3632
rect 14569 3488 14633 3552
rect 14569 3408 14633 3472
rect 14569 3328 14633 3392
rect 14569 3248 14633 3312
rect 14569 3168 14633 3232
rect 14569 3088 14633 3152
rect 14569 3008 14633 3072
rect 14569 2928 14633 2992
rect 15175 3648 15239 3712
rect 15175 3568 15239 3632
rect 15175 3488 15239 3552
rect 15175 3408 15239 3472
rect 15175 3328 15239 3392
rect 15175 3248 15239 3312
rect 15175 3168 15239 3232
rect 15175 3088 15239 3152
rect 15175 3008 15239 3072
rect 15175 2928 15239 2992
rect 15781 3648 15845 3712
rect 15781 3568 15845 3632
rect 15781 3488 15845 3552
rect 15781 3408 15845 3472
rect 15781 3328 15845 3392
rect 15781 3248 15845 3312
rect 15781 3168 15845 3232
rect 15781 3088 15845 3152
rect 15781 3008 15845 3072
rect 15781 2928 15845 2992
rect 16387 3648 16451 3712
rect 16387 3568 16451 3632
rect 16387 3488 16451 3552
rect 16387 3408 16451 3472
rect 16387 3328 16451 3392
rect 16387 3248 16451 3312
rect 16387 3168 16451 3232
rect 16387 3088 16451 3152
rect 16387 3008 16451 3072
rect 16387 2928 16451 2992
rect 16993 3648 17057 3712
rect 16993 3568 17057 3632
rect 16993 3488 17057 3552
rect 16993 3408 17057 3472
rect 16993 3328 17057 3392
rect 16993 3248 17057 3312
rect 16993 3168 17057 3232
rect 16993 3088 17057 3152
rect 16993 3008 17057 3072
rect 16993 2928 17057 2992
rect 17599 3648 17663 3712
rect 17599 3568 17663 3632
rect 17599 3488 17663 3552
rect 17599 3408 17663 3472
rect 17599 3328 17663 3392
rect 17599 3248 17663 3312
rect 17599 3168 17663 3232
rect 17599 3088 17663 3152
rect 17599 3008 17663 3072
rect 17599 2928 17663 2992
rect 18205 3648 18269 3712
rect 18205 3568 18269 3632
rect 18205 3488 18269 3552
rect 18205 3408 18269 3472
rect 18205 3328 18269 3392
rect 18205 3248 18269 3312
rect 18205 3168 18269 3232
rect 18205 3088 18269 3152
rect 18205 3008 18269 3072
rect 18205 2928 18269 2992
rect 18811 3648 18875 3712
rect 18811 3568 18875 3632
rect 18811 3488 18875 3552
rect 18811 3408 18875 3472
rect 18811 3328 18875 3392
rect 18811 3248 18875 3312
rect 18811 3168 18875 3232
rect 18811 3088 18875 3152
rect 18811 3008 18875 3072
rect 18811 2928 18875 2992
rect 19417 3648 19481 3712
rect 19417 3568 19481 3632
rect 19417 3488 19481 3552
rect 19417 3408 19481 3472
rect 19417 3328 19481 3392
rect 19417 3248 19481 3312
rect 19417 3168 19481 3232
rect 19417 3088 19481 3152
rect 19417 3008 19481 3072
rect 19417 2928 19481 2992
rect 20023 3648 20087 3712
rect 20023 3568 20087 3632
rect 20023 3488 20087 3552
rect 20023 3408 20087 3472
rect 20023 3328 20087 3392
rect 20023 3248 20087 3312
rect 20023 3168 20087 3232
rect 20023 3088 20087 3152
rect 20023 3008 20087 3072
rect 20023 2928 20087 2992
rect 20149 4808 20213 4872
rect 20149 4728 20213 4792
rect 20149 4648 20213 4712
rect 20149 4568 20213 4632
rect 20149 4488 20213 4552
rect 20149 4408 20213 4472
rect 20149 4328 20213 4392
rect 20149 4248 20213 4312
rect 20149 4168 20213 4232
rect 20149 4088 20213 4152
rect 20755 4808 20819 4872
rect 20755 4728 20819 4792
rect 20755 4648 20819 4712
rect 20755 4568 20819 4632
rect 20755 4488 20819 4552
rect 20755 4408 20819 4472
rect 20755 4328 20819 4392
rect 20755 4248 20819 4312
rect 20755 4168 20819 4232
rect 20755 4088 20819 4152
rect 21361 4808 21425 4872
rect 21361 4728 21425 4792
rect 21361 4648 21425 4712
rect 21361 4568 21425 4632
rect 21361 4488 21425 4552
rect 21361 4408 21425 4472
rect 21361 4328 21425 4392
rect 21361 4248 21425 4312
rect 21361 4168 21425 4232
rect 21361 4088 21425 4152
rect 21967 4808 22031 4872
rect 21967 4728 22031 4792
rect 21967 4648 22031 4712
rect 21967 4568 22031 4632
rect 21967 4488 22031 4552
rect 21967 4408 22031 4472
rect 21967 4328 22031 4392
rect 21967 4248 22031 4312
rect 21967 4168 22031 4232
rect 21967 4088 22031 4152
rect 22573 4808 22637 4872
rect 22573 4728 22637 4792
rect 22573 4648 22637 4712
rect 22573 4568 22637 4632
rect 22573 4488 22637 4552
rect 22573 4408 22637 4472
rect 22573 4328 22637 4392
rect 22573 4248 22637 4312
rect 22573 4168 22637 4232
rect 22573 4088 22637 4152
rect 23179 4808 23243 4872
rect 23179 4728 23243 4792
rect 23179 4648 23243 4712
rect 23179 4568 23243 4632
rect 23179 4488 23243 4552
rect 23179 4408 23243 4472
rect 23179 4328 23243 4392
rect 23179 4248 23243 4312
rect 23179 4168 23243 4232
rect 23179 4088 23243 4152
rect 23785 4808 23849 4872
rect 23785 4728 23849 4792
rect 23785 4648 23849 4712
rect 23785 4568 23849 4632
rect 23785 4488 23849 4552
rect 23785 4408 23849 4472
rect 23785 4328 23849 4392
rect 23785 4248 23849 4312
rect 23785 4168 23849 4232
rect 23785 4088 23849 4152
rect 24391 4808 24455 4872
rect 24391 4728 24455 4792
rect 24391 4648 24455 4712
rect 24391 4568 24455 4632
rect 24391 4488 24455 4552
rect 24391 4408 24455 4472
rect 24391 4328 24455 4392
rect 24391 4248 24455 4312
rect 24391 4168 24455 4232
rect 24391 4088 24455 4152
rect 24997 4808 25061 4872
rect 24997 4728 25061 4792
rect 24997 4648 25061 4712
rect 24997 4568 25061 4632
rect 24997 4488 25061 4552
rect 24997 4408 25061 4472
rect 24997 4328 25061 4392
rect 24997 4248 25061 4312
rect 24997 4168 25061 4232
rect 24997 4088 25061 4152
rect 25603 4808 25667 4872
rect 25603 4728 25667 4792
rect 25603 4648 25667 4712
rect 25603 4568 25667 4632
rect 25603 4488 25667 4552
rect 25603 4408 25667 4472
rect 25603 4328 25667 4392
rect 25603 4248 25667 4312
rect 25603 4168 25667 4232
rect 25603 4088 25667 4152
rect 26209 4808 26273 4872
rect 26209 4728 26273 4792
rect 26209 4648 26273 4712
rect 26209 4568 26273 4632
rect 26209 4488 26273 4552
rect 26209 4408 26273 4472
rect 26209 4328 26273 4392
rect 26209 4248 26273 4312
rect 26209 4168 26273 4232
rect 26209 4088 26273 4152
rect 26815 4808 26879 4872
rect 26815 4728 26879 4792
rect 26815 4648 26879 4712
rect 26815 4568 26879 4632
rect 26815 4488 26879 4552
rect 26815 4408 26879 4472
rect 26815 4328 26879 4392
rect 26815 4248 26879 4312
rect 26815 4168 26879 4232
rect 26815 4088 26879 4152
rect 27421 4808 27485 4872
rect 27421 4728 27485 4792
rect 27421 4648 27485 4712
rect 27421 4568 27485 4632
rect 27421 4488 27485 4552
rect 27421 4408 27485 4472
rect 27421 4328 27485 4392
rect 27421 4248 27485 4312
rect 27421 4168 27485 4232
rect 27421 4088 27485 4152
rect 28027 4808 28091 4872
rect 28027 4728 28091 4792
rect 28027 4648 28091 4712
rect 28027 4568 28091 4632
rect 28027 4488 28091 4552
rect 28027 4408 28091 4472
rect 28027 4328 28091 4392
rect 28027 4248 28091 4312
rect 28027 4168 28091 4232
rect 28027 4088 28091 4152
rect 28633 4808 28697 4872
rect 28633 4728 28697 4792
rect 28633 4648 28697 4712
rect 28633 4568 28697 4632
rect 28633 4488 28697 4552
rect 28633 4408 28697 4472
rect 28633 4328 28697 4392
rect 28633 4248 28697 4312
rect 28633 4168 28697 4232
rect 28633 4088 28697 4152
rect 29239 4808 29303 4872
rect 29239 4728 29303 4792
rect 29239 4648 29303 4712
rect 29239 4568 29303 4632
rect 29239 4488 29303 4552
rect 29239 4408 29303 4472
rect 29239 4328 29303 4392
rect 29239 4248 29303 4312
rect 29239 4168 29303 4232
rect 29239 4088 29303 4152
rect 29845 4808 29909 4872
rect 29845 4728 29909 4792
rect 29845 4648 29909 4712
rect 29845 4568 29909 4632
rect 29845 4488 29909 4552
rect 29845 4408 29909 4472
rect 29845 4328 29909 4392
rect 29845 4248 29909 4312
rect 29845 4168 29909 4232
rect 29845 4088 29909 4152
rect 30451 4808 30515 4872
rect 30451 4728 30515 4792
rect 30451 4648 30515 4712
rect 30451 4568 30515 4632
rect 30451 4488 30515 4552
rect 30451 4408 30515 4472
rect 30451 4328 30515 4392
rect 30451 4248 30515 4312
rect 30451 4168 30515 4232
rect 30451 4088 30515 4152
rect 31057 4808 31121 4872
rect 31057 4728 31121 4792
rect 31057 4648 31121 4712
rect 31057 4568 31121 4632
rect 31057 4488 31121 4552
rect 31057 4408 31121 4472
rect 31057 4328 31121 4392
rect 31057 4248 31121 4312
rect 31057 4168 31121 4232
rect 31057 4088 31121 4152
rect 31663 4808 31727 4872
rect 31663 4728 31727 4792
rect 31663 4648 31727 4712
rect 31663 4568 31727 4632
rect 31663 4488 31727 4552
rect 31663 4408 31727 4472
rect 31663 4328 31727 4392
rect 31663 4248 31727 4312
rect 31663 4168 31727 4232
rect 31663 4088 31727 4152
rect 32269 4808 32333 4872
rect 32269 4728 32333 4792
rect 32269 4648 32333 4712
rect 32269 4568 32333 4632
rect 32269 4488 32333 4552
rect 32269 4408 32333 4472
rect 32269 4328 32333 4392
rect 32269 4248 32333 4312
rect 32269 4168 32333 4232
rect 32269 4088 32333 4152
rect 32875 4808 32939 4872
rect 32875 4728 32939 4792
rect 32875 4648 32939 4712
rect 32875 4568 32939 4632
rect 32875 4488 32939 4552
rect 32875 4408 32939 4472
rect 32875 4328 32939 4392
rect 32875 4248 32939 4312
rect 32875 4168 32939 4232
rect 32875 4088 32939 4152
rect 33481 4808 33545 4872
rect 33481 4728 33545 4792
rect 33481 4648 33545 4712
rect 33481 4568 33545 4632
rect 33481 4488 33545 4552
rect 33481 4408 33545 4472
rect 33481 4328 33545 4392
rect 33481 4248 33545 4312
rect 33481 4168 33545 4232
rect 33481 4088 33545 4152
rect 34087 4808 34151 4872
rect 34087 4728 34151 4792
rect 34087 4648 34151 4712
rect 34087 4568 34151 4632
rect 34087 4488 34151 4552
rect 34087 4408 34151 4472
rect 34087 4328 34151 4392
rect 34087 4248 34151 4312
rect 34087 4168 34151 4232
rect 34087 4088 34151 4152
rect 34693 4808 34757 4872
rect 34693 4728 34757 4792
rect 34693 4648 34757 4712
rect 34693 4568 34757 4632
rect 34693 4488 34757 4552
rect 34693 4408 34757 4472
rect 34693 4328 34757 4392
rect 34693 4248 34757 4312
rect 34693 4168 34757 4232
rect 34693 4088 34757 4152
rect 35299 4808 35363 4872
rect 35299 4728 35363 4792
rect 35299 4648 35363 4712
rect 35299 4568 35363 4632
rect 35299 4488 35363 4552
rect 35299 4408 35363 4472
rect 35299 4328 35363 4392
rect 35299 4248 35363 4312
rect 35299 4168 35363 4232
rect 35299 4088 35363 4152
rect 35905 4808 35969 4872
rect 35905 4728 35969 4792
rect 35905 4648 35969 4712
rect 35905 4568 35969 4632
rect 35905 4488 35969 4552
rect 35905 4408 35969 4472
rect 35905 4328 35969 4392
rect 35905 4248 35969 4312
rect 35905 4168 35969 4232
rect 35905 4088 35969 4152
rect 36511 4808 36575 4872
rect 36511 4728 36575 4792
rect 36511 4648 36575 4712
rect 36511 4568 36575 4632
rect 36511 4488 36575 4552
rect 36511 4408 36575 4472
rect 36511 4328 36575 4392
rect 36511 4248 36575 4312
rect 36511 4168 36575 4232
rect 36511 4088 36575 4152
rect 37117 4808 37181 4872
rect 37117 4728 37181 4792
rect 37117 4648 37181 4712
rect 37117 4568 37181 4632
rect 37117 4488 37181 4552
rect 37117 4408 37181 4472
rect 37117 4328 37181 4392
rect 37117 4248 37181 4312
rect 37117 4168 37181 4232
rect 37117 4088 37181 4152
rect 37723 4808 37787 4872
rect 37723 4728 37787 4792
rect 37723 4648 37787 4712
rect 37723 4568 37787 4632
rect 37723 4488 37787 4552
rect 37723 4408 37787 4472
rect 37723 4328 37787 4392
rect 37723 4248 37787 4312
rect 37723 4168 37787 4232
rect 37723 4088 37787 4152
rect 38329 4808 38393 4872
rect 38329 4728 38393 4792
rect 38329 4648 38393 4712
rect 38329 4568 38393 4632
rect 38329 4488 38393 4552
rect 38329 4408 38393 4472
rect 38329 4328 38393 4392
rect 38329 4248 38393 4312
rect 38329 4168 38393 4232
rect 38329 4088 38393 4152
rect 38935 4808 38999 4872
rect 38935 4728 38999 4792
rect 38935 4648 38999 4712
rect 38935 4568 38999 4632
rect 38935 4488 38999 4552
rect 38935 4408 38999 4472
rect 38935 4328 38999 4392
rect 38935 4248 38999 4312
rect 38935 4168 38999 4232
rect 38935 4088 38999 4152
rect 39541 4808 39605 4872
rect 39541 4728 39605 4792
rect 39541 4648 39605 4712
rect 39541 4568 39605 4632
rect 39541 4488 39605 4552
rect 39541 4408 39605 4472
rect 39541 4328 39605 4392
rect 39541 4248 39605 4312
rect 39541 4168 39605 4232
rect 39541 4088 39605 4152
rect 20252 3868 20316 3932
rect 20332 3868 20396 3932
rect 20412 3868 20476 3932
rect 20492 3868 20556 3932
rect 20572 3868 20636 3932
rect 20652 3868 20716 3932
rect 20858 3868 20922 3932
rect 20938 3868 21002 3932
rect 21018 3868 21082 3932
rect 21098 3868 21162 3932
rect 21178 3868 21242 3932
rect 21258 3868 21322 3932
rect 21464 3868 21528 3932
rect 21544 3868 21608 3932
rect 21624 3868 21688 3932
rect 21704 3868 21768 3932
rect 21784 3868 21848 3932
rect 21864 3868 21928 3932
rect 22070 3868 22134 3932
rect 22150 3868 22214 3932
rect 22230 3868 22294 3932
rect 22310 3868 22374 3932
rect 22390 3868 22454 3932
rect 22470 3868 22534 3932
rect 22676 3868 22740 3932
rect 22756 3868 22820 3932
rect 22836 3868 22900 3932
rect 22916 3868 22980 3932
rect 22996 3868 23060 3932
rect 23076 3868 23140 3932
rect 23282 3868 23346 3932
rect 23362 3868 23426 3932
rect 23442 3868 23506 3932
rect 23522 3868 23586 3932
rect 23602 3868 23666 3932
rect 23682 3868 23746 3932
rect 23888 3868 23952 3932
rect 23968 3868 24032 3932
rect 24048 3868 24112 3932
rect 24128 3868 24192 3932
rect 24208 3868 24272 3932
rect 24288 3868 24352 3932
rect 24494 3868 24558 3932
rect 24574 3868 24638 3932
rect 24654 3868 24718 3932
rect 24734 3868 24798 3932
rect 24814 3868 24878 3932
rect 24894 3868 24958 3932
rect 25100 3868 25164 3932
rect 25180 3868 25244 3932
rect 25260 3868 25324 3932
rect 25340 3868 25404 3932
rect 25420 3868 25484 3932
rect 25500 3868 25564 3932
rect 25706 3868 25770 3932
rect 25786 3868 25850 3932
rect 25866 3868 25930 3932
rect 25946 3868 26010 3932
rect 26026 3868 26090 3932
rect 26106 3868 26170 3932
rect 26312 3868 26376 3932
rect 26392 3868 26456 3932
rect 26472 3868 26536 3932
rect 26552 3868 26616 3932
rect 26632 3868 26696 3932
rect 26712 3868 26776 3932
rect 26918 3868 26982 3932
rect 26998 3868 27062 3932
rect 27078 3868 27142 3932
rect 27158 3868 27222 3932
rect 27238 3868 27302 3932
rect 27318 3868 27382 3932
rect 27524 3868 27588 3932
rect 27604 3868 27668 3932
rect 27684 3868 27748 3932
rect 27764 3868 27828 3932
rect 27844 3868 27908 3932
rect 27924 3868 27988 3932
rect 28130 3868 28194 3932
rect 28210 3868 28274 3932
rect 28290 3868 28354 3932
rect 28370 3868 28434 3932
rect 28450 3868 28514 3932
rect 28530 3868 28594 3932
rect 28736 3868 28800 3932
rect 28816 3868 28880 3932
rect 28896 3868 28960 3932
rect 28976 3868 29040 3932
rect 29056 3868 29120 3932
rect 29136 3868 29200 3932
rect 29342 3868 29406 3932
rect 29422 3868 29486 3932
rect 29502 3868 29566 3932
rect 29582 3868 29646 3932
rect 29662 3868 29726 3932
rect 29742 3868 29806 3932
rect 29948 3868 30012 3932
rect 30028 3868 30092 3932
rect 30108 3868 30172 3932
rect 30188 3868 30252 3932
rect 30268 3868 30332 3932
rect 30348 3868 30412 3932
rect 30554 3868 30618 3932
rect 30634 3868 30698 3932
rect 30714 3868 30778 3932
rect 30794 3868 30858 3932
rect 30874 3868 30938 3932
rect 30954 3868 31018 3932
rect 31160 3868 31224 3932
rect 31240 3868 31304 3932
rect 31320 3868 31384 3932
rect 31400 3868 31464 3932
rect 31480 3868 31544 3932
rect 31560 3868 31624 3932
rect 31766 3868 31830 3932
rect 31846 3868 31910 3932
rect 31926 3868 31990 3932
rect 32006 3868 32070 3932
rect 32086 3868 32150 3932
rect 32166 3868 32230 3932
rect 32372 3868 32436 3932
rect 32452 3868 32516 3932
rect 32532 3868 32596 3932
rect 32612 3868 32676 3932
rect 32692 3868 32756 3932
rect 32772 3868 32836 3932
rect 32978 3868 33042 3932
rect 33058 3868 33122 3932
rect 33138 3868 33202 3932
rect 33218 3868 33282 3932
rect 33298 3868 33362 3932
rect 33378 3868 33442 3932
rect 33584 3868 33648 3932
rect 33664 3868 33728 3932
rect 33744 3868 33808 3932
rect 33824 3868 33888 3932
rect 33904 3868 33968 3932
rect 33984 3868 34048 3932
rect 34190 3868 34254 3932
rect 34270 3868 34334 3932
rect 34350 3868 34414 3932
rect 34430 3868 34494 3932
rect 34510 3868 34574 3932
rect 34590 3868 34654 3932
rect 34796 3868 34860 3932
rect 34876 3868 34940 3932
rect 34956 3868 35020 3932
rect 35036 3868 35100 3932
rect 35116 3868 35180 3932
rect 35196 3868 35260 3932
rect 35402 3868 35466 3932
rect 35482 3868 35546 3932
rect 35562 3868 35626 3932
rect 35642 3868 35706 3932
rect 35722 3868 35786 3932
rect 35802 3868 35866 3932
rect 36008 3868 36072 3932
rect 36088 3868 36152 3932
rect 36168 3868 36232 3932
rect 36248 3868 36312 3932
rect 36328 3868 36392 3932
rect 36408 3868 36472 3932
rect 36614 3868 36678 3932
rect 36694 3868 36758 3932
rect 36774 3868 36838 3932
rect 36854 3868 36918 3932
rect 36934 3868 36998 3932
rect 37014 3868 37078 3932
rect 37220 3868 37284 3932
rect 37300 3868 37364 3932
rect 37380 3868 37444 3932
rect 37460 3868 37524 3932
rect 37540 3868 37604 3932
rect 37620 3868 37684 3932
rect 37826 3868 37890 3932
rect 37906 3868 37970 3932
rect 37986 3868 38050 3932
rect 38066 3868 38130 3932
rect 38146 3868 38210 3932
rect 38226 3868 38290 3932
rect 38432 3868 38496 3932
rect 38512 3868 38576 3932
rect 38592 3868 38656 3932
rect 38672 3868 38736 3932
rect 38752 3868 38816 3932
rect 38832 3868 38896 3932
rect 39038 3868 39102 3932
rect 39118 3868 39182 3932
rect 39198 3868 39262 3932
rect 39278 3868 39342 3932
rect 39358 3868 39422 3932
rect 39438 3868 39502 3932
rect 20149 3648 20213 3712
rect 20149 3568 20213 3632
rect 20149 3488 20213 3552
rect 20149 3408 20213 3472
rect 20149 3328 20213 3392
rect 20149 3248 20213 3312
rect 20149 3168 20213 3232
rect 20149 3088 20213 3152
rect 20149 3008 20213 3072
rect 20149 2928 20213 2992
rect 20755 3648 20819 3712
rect 20755 3568 20819 3632
rect 20755 3488 20819 3552
rect 20755 3408 20819 3472
rect 20755 3328 20819 3392
rect 20755 3248 20819 3312
rect 20755 3168 20819 3232
rect 20755 3088 20819 3152
rect 20755 3008 20819 3072
rect 20755 2928 20819 2992
rect 21361 3648 21425 3712
rect 21361 3568 21425 3632
rect 21361 3488 21425 3552
rect 21361 3408 21425 3472
rect 21361 3328 21425 3392
rect 21361 3248 21425 3312
rect 21361 3168 21425 3232
rect 21361 3088 21425 3152
rect 21361 3008 21425 3072
rect 21361 2928 21425 2992
rect 21967 3648 22031 3712
rect 21967 3568 22031 3632
rect 21967 3488 22031 3552
rect 21967 3408 22031 3472
rect 21967 3328 22031 3392
rect 21967 3248 22031 3312
rect 21967 3168 22031 3232
rect 21967 3088 22031 3152
rect 21967 3008 22031 3072
rect 21967 2928 22031 2992
rect 22573 3648 22637 3712
rect 22573 3568 22637 3632
rect 22573 3488 22637 3552
rect 22573 3408 22637 3472
rect 22573 3328 22637 3392
rect 22573 3248 22637 3312
rect 22573 3168 22637 3232
rect 22573 3088 22637 3152
rect 22573 3008 22637 3072
rect 22573 2928 22637 2992
rect 23179 3648 23243 3712
rect 23179 3568 23243 3632
rect 23179 3488 23243 3552
rect 23179 3408 23243 3472
rect 23179 3328 23243 3392
rect 23179 3248 23243 3312
rect 23179 3168 23243 3232
rect 23179 3088 23243 3152
rect 23179 3008 23243 3072
rect 23179 2928 23243 2992
rect 23785 3648 23849 3712
rect 23785 3568 23849 3632
rect 23785 3488 23849 3552
rect 23785 3408 23849 3472
rect 23785 3328 23849 3392
rect 23785 3248 23849 3312
rect 23785 3168 23849 3232
rect 23785 3088 23849 3152
rect 23785 3008 23849 3072
rect 23785 2928 23849 2992
rect 24391 3648 24455 3712
rect 24391 3568 24455 3632
rect 24391 3488 24455 3552
rect 24391 3408 24455 3472
rect 24391 3328 24455 3392
rect 24391 3248 24455 3312
rect 24391 3168 24455 3232
rect 24391 3088 24455 3152
rect 24391 3008 24455 3072
rect 24391 2928 24455 2992
rect 24997 3648 25061 3712
rect 24997 3568 25061 3632
rect 24997 3488 25061 3552
rect 24997 3408 25061 3472
rect 24997 3328 25061 3392
rect 24997 3248 25061 3312
rect 24997 3168 25061 3232
rect 24997 3088 25061 3152
rect 24997 3008 25061 3072
rect 24997 2928 25061 2992
rect 25603 3648 25667 3712
rect 25603 3568 25667 3632
rect 25603 3488 25667 3552
rect 25603 3408 25667 3472
rect 25603 3328 25667 3392
rect 25603 3248 25667 3312
rect 25603 3168 25667 3232
rect 25603 3088 25667 3152
rect 25603 3008 25667 3072
rect 25603 2928 25667 2992
rect 26209 3648 26273 3712
rect 26209 3568 26273 3632
rect 26209 3488 26273 3552
rect 26209 3408 26273 3472
rect 26209 3328 26273 3392
rect 26209 3248 26273 3312
rect 26209 3168 26273 3232
rect 26209 3088 26273 3152
rect 26209 3008 26273 3072
rect 26209 2928 26273 2992
rect 26815 3648 26879 3712
rect 26815 3568 26879 3632
rect 26815 3488 26879 3552
rect 26815 3408 26879 3472
rect 26815 3328 26879 3392
rect 26815 3248 26879 3312
rect 26815 3168 26879 3232
rect 26815 3088 26879 3152
rect 26815 3008 26879 3072
rect 26815 2928 26879 2992
rect 27421 3648 27485 3712
rect 27421 3568 27485 3632
rect 27421 3488 27485 3552
rect 27421 3408 27485 3472
rect 27421 3328 27485 3392
rect 27421 3248 27485 3312
rect 27421 3168 27485 3232
rect 27421 3088 27485 3152
rect 27421 3008 27485 3072
rect 27421 2928 27485 2992
rect 28027 3648 28091 3712
rect 28027 3568 28091 3632
rect 28027 3488 28091 3552
rect 28027 3408 28091 3472
rect 28027 3328 28091 3392
rect 28027 3248 28091 3312
rect 28027 3168 28091 3232
rect 28027 3088 28091 3152
rect 28027 3008 28091 3072
rect 28027 2928 28091 2992
rect 28633 3648 28697 3712
rect 28633 3568 28697 3632
rect 28633 3488 28697 3552
rect 28633 3408 28697 3472
rect 28633 3328 28697 3392
rect 28633 3248 28697 3312
rect 28633 3179 28697 3232
rect 28633 3168 28637 3179
rect 28637 3168 28693 3179
rect 28693 3168 28697 3179
rect 28633 3123 28637 3152
rect 28637 3123 28693 3152
rect 28693 3123 28697 3152
rect 28633 3088 28697 3123
rect 28633 3008 28697 3072
rect 28633 2928 28697 2992
rect 29239 3648 29303 3712
rect 29239 3568 29303 3632
rect 29239 3488 29303 3552
rect 29239 3408 29303 3472
rect 29239 3328 29303 3392
rect 29239 3248 29303 3312
rect 29239 3168 29303 3232
rect 29239 3088 29303 3152
rect 29239 3008 29303 3072
rect 29239 2928 29303 2992
rect 29845 3648 29909 3712
rect 29845 3568 29909 3632
rect 29845 3488 29909 3552
rect 29845 3408 29909 3472
rect 29845 3328 29909 3392
rect 29845 3248 29909 3312
rect 29845 3168 29909 3232
rect 29845 3088 29909 3152
rect 29845 3008 29909 3072
rect 29845 2928 29909 2992
rect 30451 3648 30515 3712
rect 30451 3568 30515 3632
rect 30451 3488 30515 3552
rect 30451 3408 30515 3472
rect 30451 3328 30515 3392
rect 30451 3248 30515 3312
rect 30451 3168 30515 3232
rect 30451 3088 30515 3152
rect 30451 3008 30515 3072
rect 30451 2928 30515 2992
rect 31057 3648 31121 3712
rect 31057 3568 31121 3632
rect 31057 3488 31121 3552
rect 31057 3408 31121 3472
rect 31057 3328 31121 3392
rect 31057 3248 31121 3312
rect 31057 3168 31121 3232
rect 31057 3088 31121 3152
rect 31057 3008 31121 3072
rect 31057 2928 31121 2992
rect 31663 3648 31727 3712
rect 31663 3568 31727 3632
rect 31663 3488 31727 3552
rect 31663 3408 31727 3472
rect 31663 3328 31727 3392
rect 31663 3248 31727 3312
rect 31663 3168 31727 3232
rect 31663 3088 31727 3152
rect 31663 3008 31727 3072
rect 31663 2928 31727 2992
rect 32269 3648 32333 3712
rect 32269 3568 32333 3632
rect 32269 3488 32333 3552
rect 32269 3408 32333 3472
rect 32269 3328 32333 3392
rect 32269 3248 32333 3312
rect 32269 3168 32333 3232
rect 32269 3088 32333 3152
rect 32269 3008 32333 3072
rect 32269 2928 32333 2992
rect 32875 3648 32939 3712
rect 32875 3568 32939 3632
rect 32875 3488 32939 3552
rect 32875 3408 32939 3472
rect 32875 3328 32939 3392
rect 32875 3248 32939 3312
rect 32875 3168 32939 3232
rect 32875 3088 32939 3152
rect 32875 3008 32939 3072
rect 32875 2928 32939 2992
rect 33481 3648 33545 3712
rect 33481 3568 33545 3632
rect 33481 3488 33545 3552
rect 33481 3408 33545 3472
rect 33481 3328 33545 3392
rect 33481 3248 33545 3312
rect 33481 3168 33545 3232
rect 33481 3088 33545 3152
rect 33481 3008 33545 3072
rect 33481 2928 33545 2992
rect 34087 3648 34151 3712
rect 34087 3568 34151 3632
rect 34087 3488 34151 3552
rect 34087 3408 34151 3472
rect 34087 3328 34151 3392
rect 34087 3248 34151 3312
rect 34087 3168 34151 3232
rect 34087 3088 34151 3152
rect 34087 3008 34151 3072
rect 34087 2928 34151 2992
rect 34693 3648 34757 3712
rect 34693 3568 34757 3632
rect 34693 3488 34757 3552
rect 34693 3408 34757 3472
rect 34693 3328 34757 3392
rect 34693 3248 34757 3312
rect 34693 3168 34757 3232
rect 34693 3088 34757 3152
rect 34693 3008 34757 3072
rect 34693 2928 34757 2992
rect 35299 3648 35363 3712
rect 35299 3568 35363 3632
rect 35299 3488 35363 3552
rect 35299 3408 35363 3472
rect 35299 3328 35363 3392
rect 35299 3248 35363 3312
rect 35299 3168 35363 3232
rect 35299 3088 35363 3152
rect 35299 3008 35363 3072
rect 35299 2928 35363 2992
rect 35905 3648 35969 3712
rect 35905 3568 35969 3632
rect 35905 3488 35969 3552
rect 35905 3408 35969 3472
rect 35905 3328 35969 3392
rect 35905 3248 35969 3312
rect 35905 3168 35969 3232
rect 35905 3088 35969 3152
rect 35905 3008 35969 3072
rect 35905 2928 35969 2992
rect 36511 3648 36575 3712
rect 36511 3568 36575 3632
rect 36511 3488 36575 3552
rect 36511 3408 36575 3472
rect 36511 3328 36575 3392
rect 36511 3248 36575 3312
rect 36511 3168 36575 3232
rect 36511 3088 36575 3152
rect 36511 3008 36575 3072
rect 36511 2928 36575 2992
rect 37117 3648 37181 3712
rect 37117 3568 37181 3632
rect 37117 3488 37181 3552
rect 37117 3408 37181 3472
rect 37117 3328 37181 3392
rect 37117 3248 37181 3312
rect 37117 3168 37181 3232
rect 37117 3088 37181 3152
rect 37117 3008 37181 3072
rect 37117 2928 37181 2992
rect 37723 3648 37787 3712
rect 37723 3568 37787 3632
rect 37723 3488 37787 3552
rect 37723 3408 37787 3472
rect 37723 3328 37787 3392
rect 37723 3248 37787 3312
rect 37723 3168 37787 3232
rect 37723 3088 37787 3152
rect 37723 3008 37787 3072
rect 37723 2928 37787 2992
rect 38329 3648 38393 3712
rect 38329 3568 38393 3632
rect 38329 3488 38393 3552
rect 38329 3408 38393 3472
rect 38329 3328 38393 3392
rect 38329 3248 38393 3312
rect 38329 3168 38393 3232
rect 38329 3088 38393 3152
rect 38329 3008 38393 3072
rect 38329 2928 38393 2992
rect 38935 3648 38999 3712
rect 38935 3568 38999 3632
rect 38935 3488 38999 3552
rect 38935 3408 38999 3472
rect 38935 3328 38999 3392
rect 38935 3248 38999 3312
rect 38935 3168 38999 3232
rect 38935 3088 38999 3152
rect 38935 3008 38999 3072
rect 38935 2928 38999 2992
rect 39541 3648 39605 3712
rect 39541 3568 39605 3632
rect 39541 3488 39605 3552
rect 39541 3408 39605 3472
rect 39541 3328 39605 3392
rect 39541 3248 39605 3312
rect 39541 3168 39605 3232
rect 39541 3088 39605 3152
rect 39541 3008 39605 3072
rect 39541 2928 39605 2992
rect -355 2708 -291 2772
rect -275 2708 -211 2772
rect -195 2708 -131 2772
rect -115 2708 -51 2772
rect -35 2708 29 2772
rect 45 2708 109 2772
rect 459 2708 523 2772
rect 539 2708 603 2772
rect 619 2708 683 2772
rect 699 2708 763 2772
rect 779 2708 843 2772
rect 859 2708 923 2772
rect 1371 2708 1435 2772
rect 1451 2708 1515 2772
rect 1531 2708 1595 2772
rect 1611 2708 1675 2772
rect 1691 2708 1755 2772
rect 1771 2708 1835 2772
rect 1977 2708 2041 2772
rect 2057 2708 2121 2772
rect 2137 2708 2201 2772
rect 2217 2708 2281 2772
rect 2297 2708 2361 2772
rect 2377 2708 2441 2772
rect 2905 2708 2969 2772
rect 2985 2708 3049 2772
rect 3065 2708 3129 2772
rect 3145 2708 3209 2772
rect 3225 2708 3289 2772
rect 3305 2708 3369 2772
rect 3511 2708 3575 2772
rect 3591 2708 3655 2772
rect 3671 2708 3735 2772
rect 3751 2708 3815 2772
rect 3831 2708 3895 2772
rect 3911 2708 3975 2772
rect 4117 2708 4181 2772
rect 4197 2708 4261 2772
rect 4277 2708 4341 2772
rect 4357 2708 4421 2772
rect 4437 2708 4501 2772
rect 4517 2708 4581 2772
rect 4723 2708 4787 2772
rect 4803 2708 4867 2772
rect 4883 2708 4947 2772
rect 4963 2708 5027 2772
rect 5043 2708 5107 2772
rect 5123 2708 5187 2772
rect 5456 2708 5520 2772
rect 5536 2708 5600 2772
rect 5616 2708 5680 2772
rect 5696 2708 5760 2772
rect 5776 2708 5840 2772
rect 5856 2708 5920 2772
rect 6062 2708 6126 2772
rect 6142 2708 6206 2772
rect 6222 2708 6286 2772
rect 6302 2708 6366 2772
rect 6382 2708 6446 2772
rect 6462 2708 6526 2772
rect 6668 2708 6732 2772
rect 6748 2708 6812 2772
rect 6828 2708 6892 2772
rect 6908 2708 6972 2772
rect 6988 2708 7052 2772
rect 7068 2708 7132 2772
rect 7274 2708 7338 2772
rect 7354 2708 7418 2772
rect 7434 2708 7498 2772
rect 7514 2708 7578 2772
rect 7594 2708 7658 2772
rect 7674 2708 7738 2772
rect 7880 2708 7944 2772
rect 7960 2708 8024 2772
rect 8040 2708 8104 2772
rect 8120 2708 8184 2772
rect 8200 2708 8264 2772
rect 8280 2708 8344 2772
rect 8486 2708 8550 2772
rect 8566 2708 8630 2772
rect 8646 2708 8710 2772
rect 8726 2708 8790 2772
rect 8806 2708 8870 2772
rect 8886 2708 8950 2772
rect 9092 2708 9156 2772
rect 9172 2708 9236 2772
rect 9252 2708 9316 2772
rect 9332 2708 9396 2772
rect 9412 2708 9476 2772
rect 9492 2708 9556 2772
rect 9698 2708 9762 2772
rect 9778 2708 9842 2772
rect 9858 2708 9922 2772
rect 9938 2708 10002 2772
rect 10018 2708 10082 2772
rect 10098 2708 10162 2772
rect 10430 2708 10494 2772
rect 10510 2708 10574 2772
rect 10590 2708 10654 2772
rect 10670 2708 10734 2772
rect 10750 2708 10814 2772
rect 10830 2708 10894 2772
rect 11036 2708 11100 2772
rect 11116 2708 11180 2772
rect 11196 2708 11260 2772
rect 11276 2708 11340 2772
rect 11356 2708 11420 2772
rect 11436 2708 11500 2772
rect 11642 2708 11706 2772
rect 11722 2708 11786 2772
rect 11802 2708 11866 2772
rect 11882 2708 11946 2772
rect 11962 2708 12026 2772
rect 12042 2708 12106 2772
rect 12248 2708 12312 2772
rect 12328 2708 12392 2772
rect 12408 2708 12472 2772
rect 12488 2708 12552 2772
rect 12568 2708 12632 2772
rect 12648 2708 12712 2772
rect 12854 2708 12918 2772
rect 12934 2708 12998 2772
rect 13014 2708 13078 2772
rect 13094 2708 13158 2772
rect 13174 2708 13238 2772
rect 13254 2708 13318 2772
rect 13460 2708 13524 2772
rect 13540 2708 13604 2772
rect 13620 2708 13684 2772
rect 13700 2708 13764 2772
rect 13780 2708 13844 2772
rect 13860 2708 13924 2772
rect 14066 2708 14130 2772
rect 14146 2708 14210 2772
rect 14226 2708 14290 2772
rect 14306 2708 14370 2772
rect 14386 2708 14450 2772
rect 14466 2708 14530 2772
rect 14672 2708 14736 2772
rect 14752 2708 14816 2772
rect 14832 2708 14896 2772
rect 14912 2708 14976 2772
rect 14992 2708 15056 2772
rect 15072 2708 15136 2772
rect 15278 2708 15342 2772
rect 15358 2708 15422 2772
rect 15438 2708 15502 2772
rect 15518 2708 15582 2772
rect 15598 2708 15662 2772
rect 15678 2708 15742 2772
rect 15884 2708 15948 2772
rect 15964 2708 16028 2772
rect 16044 2708 16108 2772
rect 16124 2708 16188 2772
rect 16204 2708 16268 2772
rect 16284 2708 16348 2772
rect 16490 2708 16554 2772
rect 16570 2708 16634 2772
rect 16650 2708 16714 2772
rect 16730 2708 16794 2772
rect 16810 2708 16874 2772
rect 16890 2708 16954 2772
rect 17096 2708 17160 2772
rect 17176 2708 17240 2772
rect 17256 2708 17320 2772
rect 17336 2708 17400 2772
rect 17416 2708 17480 2772
rect 17496 2708 17560 2772
rect 17702 2708 17766 2772
rect 17782 2708 17846 2772
rect 17862 2708 17926 2772
rect 17942 2708 18006 2772
rect 18022 2708 18086 2772
rect 18102 2708 18166 2772
rect 18308 2708 18372 2772
rect 18388 2708 18452 2772
rect 18468 2708 18532 2772
rect 18548 2708 18612 2772
rect 18628 2708 18692 2772
rect 18708 2708 18772 2772
rect 18914 2708 18978 2772
rect 18994 2708 19058 2772
rect 19074 2708 19138 2772
rect 19154 2708 19218 2772
rect 19234 2708 19298 2772
rect 19314 2708 19378 2772
rect 19520 2708 19584 2772
rect 19600 2708 19664 2772
rect 19680 2708 19744 2772
rect 19760 2708 19824 2772
rect 19840 2708 19904 2772
rect 19920 2708 19984 2772
rect 20252 2708 20316 2772
rect 20332 2708 20396 2772
rect 20412 2708 20476 2772
rect 20492 2708 20556 2772
rect 20572 2708 20636 2772
rect 20652 2708 20716 2772
rect 20858 2708 20922 2772
rect 20938 2708 21002 2772
rect 21018 2708 21082 2772
rect 21098 2708 21162 2772
rect 21178 2708 21242 2772
rect 21258 2708 21322 2772
rect 21464 2708 21528 2772
rect 21544 2708 21608 2772
rect 21624 2708 21688 2772
rect 21704 2708 21768 2772
rect 21784 2708 21848 2772
rect 21864 2708 21928 2772
rect 22070 2708 22134 2772
rect 22150 2708 22214 2772
rect 22230 2708 22294 2772
rect 22310 2708 22374 2772
rect 22390 2708 22454 2772
rect 22470 2708 22534 2772
rect 22676 2708 22740 2772
rect 22756 2708 22820 2772
rect 22836 2708 22900 2772
rect 22916 2708 22980 2772
rect 22996 2708 23060 2772
rect 23076 2708 23140 2772
rect 23282 2708 23346 2772
rect 23362 2708 23426 2772
rect 23442 2708 23506 2772
rect 23522 2708 23586 2772
rect 23602 2708 23666 2772
rect 23682 2708 23746 2772
rect 23888 2708 23952 2772
rect 23968 2708 24032 2772
rect 24048 2708 24112 2772
rect 24128 2708 24192 2772
rect 24208 2708 24272 2772
rect 24288 2708 24352 2772
rect 24494 2708 24558 2772
rect 24574 2708 24638 2772
rect 24654 2708 24718 2772
rect 24734 2708 24798 2772
rect 24814 2708 24878 2772
rect 24894 2708 24958 2772
rect 25100 2708 25164 2772
rect 25180 2708 25244 2772
rect 25260 2708 25324 2772
rect 25340 2708 25404 2772
rect 25420 2708 25484 2772
rect 25500 2708 25564 2772
rect 25706 2708 25770 2772
rect 25786 2708 25850 2772
rect 25866 2708 25930 2772
rect 25946 2708 26010 2772
rect 26026 2708 26090 2772
rect 26106 2708 26170 2772
rect 26312 2708 26376 2772
rect 26392 2708 26456 2772
rect 26472 2708 26536 2772
rect 26552 2708 26616 2772
rect 26632 2708 26696 2772
rect 26712 2708 26776 2772
rect 26918 2708 26982 2772
rect 26998 2708 27062 2772
rect 27078 2708 27142 2772
rect 27158 2708 27222 2772
rect 27238 2708 27302 2772
rect 27318 2708 27382 2772
rect 27524 2708 27588 2772
rect 27604 2708 27668 2772
rect 27684 2708 27748 2772
rect 27764 2708 27828 2772
rect 27844 2708 27908 2772
rect 27924 2708 27988 2772
rect 28130 2708 28194 2772
rect 28210 2708 28274 2772
rect 28290 2708 28354 2772
rect 28370 2708 28434 2772
rect 28450 2708 28514 2772
rect 28530 2708 28594 2772
rect 28736 2708 28800 2772
rect 28816 2708 28880 2772
rect 28896 2708 28960 2772
rect 28976 2708 29040 2772
rect 29056 2708 29120 2772
rect 29136 2708 29200 2772
rect 29342 2708 29406 2772
rect 29422 2708 29486 2772
rect 29502 2708 29566 2772
rect 29582 2708 29646 2772
rect 29662 2708 29726 2772
rect 29742 2708 29806 2772
rect 29948 2708 30012 2772
rect 30028 2708 30092 2772
rect 30108 2708 30172 2772
rect 30188 2708 30252 2772
rect 30268 2708 30332 2772
rect 30348 2708 30412 2772
rect 30554 2708 30618 2772
rect 30634 2708 30698 2772
rect 30714 2708 30778 2772
rect 30794 2708 30858 2772
rect 30874 2708 30938 2772
rect 30954 2708 31018 2772
rect 31160 2708 31224 2772
rect 31240 2708 31304 2772
rect 31320 2708 31384 2772
rect 31400 2708 31464 2772
rect 31480 2708 31544 2772
rect 31560 2708 31624 2772
rect 31766 2708 31830 2772
rect 31846 2708 31910 2772
rect 31926 2708 31990 2772
rect 32006 2708 32070 2772
rect 32086 2708 32150 2772
rect 32166 2708 32230 2772
rect 32372 2708 32436 2772
rect 32452 2708 32516 2772
rect 32532 2708 32596 2772
rect 32612 2708 32676 2772
rect 32692 2708 32756 2772
rect 32772 2708 32836 2772
rect 32978 2708 33042 2772
rect 33058 2708 33122 2772
rect 33138 2708 33202 2772
rect 33218 2708 33282 2772
rect 33298 2708 33362 2772
rect 33378 2708 33442 2772
rect 33584 2708 33648 2772
rect 33664 2708 33728 2772
rect 33744 2708 33808 2772
rect 33824 2708 33888 2772
rect 33904 2708 33968 2772
rect 33984 2708 34048 2772
rect 34190 2708 34254 2772
rect 34270 2708 34334 2772
rect 34350 2708 34414 2772
rect 34430 2708 34494 2772
rect 34510 2708 34574 2772
rect 34590 2708 34654 2772
rect 34796 2708 34860 2772
rect 34876 2708 34940 2772
rect 34956 2708 35020 2772
rect 35036 2708 35100 2772
rect 35116 2708 35180 2772
rect 35196 2708 35260 2772
rect 35402 2708 35466 2772
rect 35482 2708 35546 2772
rect 35562 2708 35626 2772
rect 35642 2708 35706 2772
rect 35722 2708 35786 2772
rect 35802 2708 35866 2772
rect 36008 2708 36072 2772
rect 36088 2708 36152 2772
rect 36168 2708 36232 2772
rect 36248 2708 36312 2772
rect 36328 2708 36392 2772
rect 36408 2708 36472 2772
rect 36614 2708 36678 2772
rect 36694 2708 36758 2772
rect 36774 2708 36838 2772
rect 36854 2708 36918 2772
rect 36934 2708 36998 2772
rect 37014 2708 37078 2772
rect 37220 2708 37284 2772
rect 37300 2708 37364 2772
rect 37380 2708 37444 2772
rect 37460 2708 37524 2772
rect 37540 2708 37604 2772
rect 37620 2708 37684 2772
rect 37826 2708 37890 2772
rect 37906 2708 37970 2772
rect 37986 2708 38050 2772
rect 38066 2708 38130 2772
rect 38146 2708 38210 2772
rect 38226 2708 38290 2772
rect 38432 2708 38496 2772
rect 38512 2708 38576 2772
rect 38592 2708 38656 2772
rect 38672 2708 38736 2772
rect 38752 2708 38816 2772
rect 38832 2708 38896 2772
rect 39038 2708 39102 2772
rect 39118 2708 39182 2772
rect 39198 2708 39262 2772
rect 39278 2708 39342 2772
rect 39358 2708 39422 2772
rect 39438 2708 39502 2772
rect -355 2540 -291 2604
rect -275 2540 -211 2604
rect -195 2540 -131 2604
rect -115 2600 -51 2604
rect -115 2544 -91 2600
rect -91 2544 -51 2600
rect -115 2540 -51 2544
rect -35 2540 29 2604
rect 45 2540 109 2604
rect 459 2540 523 2604
rect 539 2540 603 2604
rect 619 2540 683 2604
rect 699 2540 763 2604
rect 779 2540 843 2604
rect 859 2540 923 2604
rect 1371 2540 1435 2604
rect 1451 2540 1515 2604
rect 1531 2540 1595 2604
rect 1611 2540 1675 2604
rect 1691 2540 1755 2604
rect 1771 2540 1835 2604
rect 1977 2540 2041 2604
rect 2057 2540 2121 2604
rect 2137 2540 2201 2604
rect 2217 2540 2281 2604
rect 2297 2540 2361 2604
rect 2377 2540 2441 2604
rect 2905 2540 2969 2604
rect 2985 2540 3049 2604
rect 3065 2540 3129 2604
rect 3145 2540 3209 2604
rect 3225 2540 3289 2604
rect 3305 2540 3369 2604
rect 3511 2540 3575 2604
rect 3591 2540 3655 2604
rect 3671 2540 3735 2604
rect 3751 2540 3815 2604
rect 3831 2540 3895 2604
rect 3911 2540 3975 2604
rect 4117 2540 4181 2604
rect 4197 2540 4261 2604
rect 4277 2540 4341 2604
rect 4357 2540 4421 2604
rect 4437 2540 4501 2604
rect 4517 2540 4581 2604
rect 4723 2540 4787 2604
rect 4803 2540 4867 2604
rect 4883 2540 4947 2604
rect 4963 2540 5027 2604
rect 5043 2540 5107 2604
rect 5123 2540 5187 2604
rect 5456 2540 5520 2604
rect 5536 2540 5600 2604
rect 5616 2540 5680 2604
rect 5696 2540 5760 2604
rect 5776 2540 5840 2604
rect 5856 2540 5920 2604
rect 6062 2540 6126 2604
rect 6142 2540 6206 2604
rect 6222 2540 6286 2604
rect 6302 2540 6366 2604
rect 6382 2540 6446 2604
rect 6462 2540 6526 2604
rect 6668 2540 6732 2604
rect 6748 2540 6812 2604
rect 6828 2540 6892 2604
rect 6908 2540 6972 2604
rect 6988 2540 7052 2604
rect 7068 2540 7132 2604
rect 7274 2540 7338 2604
rect 7354 2540 7418 2604
rect 7434 2540 7498 2604
rect 7514 2540 7578 2604
rect 7594 2540 7658 2604
rect 7674 2540 7738 2604
rect 7880 2540 7944 2604
rect 7960 2540 8024 2604
rect 8040 2540 8104 2604
rect 8120 2540 8184 2604
rect 8200 2540 8264 2604
rect 8280 2540 8344 2604
rect 8486 2540 8550 2604
rect 8566 2540 8630 2604
rect 8646 2540 8710 2604
rect 8726 2540 8790 2604
rect 8806 2540 8870 2604
rect 8886 2540 8950 2604
rect 9092 2540 9156 2604
rect 9172 2540 9236 2604
rect 9252 2540 9316 2604
rect 9332 2540 9396 2604
rect 9412 2540 9476 2604
rect 9492 2540 9556 2604
rect 9698 2540 9762 2604
rect 9778 2540 9842 2604
rect 9858 2540 9922 2604
rect 9938 2540 10002 2604
rect 10018 2540 10082 2604
rect 10098 2540 10162 2604
rect 10430 2540 10494 2604
rect 10510 2540 10574 2604
rect 10590 2540 10654 2604
rect 10670 2540 10734 2604
rect 10750 2540 10814 2604
rect 10830 2540 10894 2604
rect 11036 2540 11100 2604
rect 11116 2540 11180 2604
rect 11196 2540 11260 2604
rect 11276 2540 11340 2604
rect 11356 2540 11420 2604
rect 11436 2540 11500 2604
rect 11642 2540 11706 2604
rect 11722 2540 11786 2604
rect 11802 2540 11866 2604
rect 11882 2540 11946 2604
rect 11962 2540 12026 2604
rect 12042 2540 12106 2604
rect 12248 2540 12312 2604
rect 12328 2540 12392 2604
rect 12408 2540 12472 2604
rect 12488 2540 12552 2604
rect 12568 2540 12632 2604
rect 12648 2540 12712 2604
rect 12854 2540 12918 2604
rect 12934 2540 12998 2604
rect 13014 2540 13078 2604
rect 13094 2540 13158 2604
rect 13174 2540 13238 2604
rect 13254 2540 13318 2604
rect 13460 2540 13524 2604
rect 13540 2540 13604 2604
rect 13620 2540 13684 2604
rect 13700 2540 13764 2604
rect 13780 2540 13844 2604
rect 13860 2540 13924 2604
rect 14066 2540 14130 2604
rect 14146 2540 14210 2604
rect 14226 2540 14290 2604
rect 14306 2540 14370 2604
rect 14386 2540 14450 2604
rect 14466 2540 14530 2604
rect 14672 2540 14736 2604
rect 14752 2540 14816 2604
rect 14832 2540 14896 2604
rect 14912 2540 14976 2604
rect 14992 2540 15056 2604
rect 15072 2540 15136 2604
rect 15278 2540 15342 2604
rect 15358 2540 15422 2604
rect 15438 2540 15502 2604
rect 15518 2540 15582 2604
rect 15598 2540 15662 2604
rect 15678 2540 15742 2604
rect 15884 2540 15948 2604
rect 15964 2540 16028 2604
rect 16044 2540 16108 2604
rect 16124 2540 16188 2604
rect 16204 2540 16268 2604
rect 16284 2540 16348 2604
rect 16490 2540 16554 2604
rect 16570 2540 16634 2604
rect 16650 2540 16714 2604
rect 16730 2540 16794 2604
rect 16810 2540 16874 2604
rect 16890 2540 16954 2604
rect 17096 2540 17160 2604
rect 17176 2540 17240 2604
rect 17256 2540 17320 2604
rect 17336 2540 17400 2604
rect 17416 2540 17480 2604
rect 17496 2540 17560 2604
rect 17702 2540 17766 2604
rect 17782 2540 17846 2604
rect 17862 2540 17926 2604
rect 17942 2540 18006 2604
rect 18022 2540 18086 2604
rect 18102 2540 18166 2604
rect 18308 2540 18372 2604
rect 18388 2540 18452 2604
rect 18468 2540 18532 2604
rect 18548 2540 18612 2604
rect 18628 2540 18692 2604
rect 18708 2540 18772 2604
rect 18914 2540 18978 2604
rect 18994 2540 19058 2604
rect 19074 2540 19138 2604
rect 19154 2540 19218 2604
rect 19234 2540 19298 2604
rect 19314 2540 19378 2604
rect 19520 2540 19584 2604
rect 19600 2540 19664 2604
rect 19680 2540 19744 2604
rect 19760 2540 19824 2604
rect 19840 2540 19904 2604
rect 19920 2540 19984 2604
rect 20252 2540 20316 2604
rect 20332 2540 20396 2604
rect 20412 2540 20476 2604
rect 20492 2540 20556 2604
rect 20572 2540 20636 2604
rect 20652 2540 20716 2604
rect 20858 2540 20922 2604
rect 20938 2540 21002 2604
rect 21018 2540 21082 2604
rect 21098 2540 21162 2604
rect 21178 2540 21242 2604
rect 21258 2540 21322 2604
rect 21464 2540 21528 2604
rect 21544 2540 21608 2604
rect 21624 2540 21688 2604
rect 21704 2540 21768 2604
rect 21784 2540 21848 2604
rect 21864 2540 21928 2604
rect 22070 2540 22134 2604
rect 22150 2540 22214 2604
rect 22230 2540 22294 2604
rect 22310 2540 22374 2604
rect 22390 2540 22454 2604
rect 22470 2540 22534 2604
rect 22676 2540 22740 2604
rect 22756 2540 22820 2604
rect 22836 2540 22900 2604
rect 22916 2540 22980 2604
rect 22996 2540 23060 2604
rect 23076 2540 23140 2604
rect 23282 2540 23346 2604
rect 23362 2540 23426 2604
rect 23442 2540 23506 2604
rect 23522 2540 23586 2604
rect 23602 2540 23666 2604
rect 23682 2540 23746 2604
rect 23888 2540 23952 2604
rect 23968 2540 24032 2604
rect 24048 2540 24112 2604
rect 24128 2540 24192 2604
rect 24208 2540 24272 2604
rect 24288 2540 24352 2604
rect 24494 2540 24558 2604
rect 24574 2540 24638 2604
rect 24654 2540 24718 2604
rect 24734 2540 24798 2604
rect 24814 2540 24878 2604
rect 24894 2540 24958 2604
rect 25100 2540 25164 2604
rect 25180 2540 25244 2604
rect 25260 2540 25324 2604
rect 25340 2540 25404 2604
rect 25420 2540 25484 2604
rect 25500 2540 25564 2604
rect 25706 2540 25770 2604
rect 25786 2540 25850 2604
rect 25866 2540 25930 2604
rect 25946 2540 26010 2604
rect 26026 2540 26090 2604
rect 26106 2540 26170 2604
rect 26312 2540 26376 2604
rect 26392 2540 26456 2604
rect 26472 2540 26536 2604
rect 26552 2540 26616 2604
rect 26632 2540 26696 2604
rect 26712 2540 26776 2604
rect 26918 2540 26982 2604
rect 26998 2540 27062 2604
rect 27078 2540 27142 2604
rect 27158 2540 27222 2604
rect 27238 2540 27302 2604
rect 27318 2540 27382 2604
rect 27524 2540 27588 2604
rect 27604 2540 27668 2604
rect 27684 2540 27748 2604
rect 27764 2540 27828 2604
rect 27844 2540 27908 2604
rect 27924 2540 27988 2604
rect 28130 2540 28194 2604
rect 28210 2540 28274 2604
rect 28290 2540 28354 2604
rect 28370 2540 28434 2604
rect 28450 2540 28514 2604
rect 28530 2540 28594 2604
rect 28736 2540 28800 2604
rect 28816 2540 28880 2604
rect 28896 2540 28960 2604
rect 28976 2540 29040 2604
rect 29056 2540 29120 2604
rect 29136 2540 29200 2604
rect 29342 2540 29406 2604
rect 29422 2540 29486 2604
rect 29502 2540 29566 2604
rect 29582 2540 29646 2604
rect 29662 2540 29726 2604
rect 29742 2540 29806 2604
rect 29948 2540 30012 2604
rect 30028 2540 30092 2604
rect 30108 2540 30172 2604
rect 30188 2540 30252 2604
rect 30268 2540 30332 2604
rect 30348 2540 30412 2604
rect 30554 2540 30618 2604
rect 30634 2540 30698 2604
rect 30714 2540 30778 2604
rect 30794 2540 30858 2604
rect 30874 2540 30938 2604
rect 30954 2540 31018 2604
rect 31160 2540 31224 2604
rect 31240 2540 31304 2604
rect 31320 2540 31384 2604
rect 31400 2540 31464 2604
rect 31480 2540 31544 2604
rect 31560 2540 31624 2604
rect 31766 2540 31830 2604
rect 31846 2540 31910 2604
rect 31926 2540 31990 2604
rect 32006 2540 32070 2604
rect 32086 2540 32150 2604
rect 32166 2540 32230 2604
rect 32372 2540 32436 2604
rect 32452 2540 32516 2604
rect 32532 2540 32596 2604
rect 32612 2540 32676 2604
rect 32692 2540 32756 2604
rect 32772 2540 32836 2604
rect 32978 2540 33042 2604
rect 33058 2540 33122 2604
rect 33138 2540 33202 2604
rect 33218 2540 33282 2604
rect 33298 2540 33362 2604
rect 33378 2540 33442 2604
rect 33584 2540 33648 2604
rect 33664 2540 33728 2604
rect 33744 2540 33808 2604
rect 33824 2540 33888 2604
rect 33904 2540 33968 2604
rect 33984 2540 34048 2604
rect 34190 2540 34254 2604
rect 34270 2540 34334 2604
rect 34350 2540 34414 2604
rect 34430 2540 34494 2604
rect 34510 2540 34574 2604
rect 34590 2540 34654 2604
rect 34796 2540 34860 2604
rect 34876 2540 34940 2604
rect 34956 2540 35020 2604
rect 35036 2540 35100 2604
rect 35116 2540 35180 2604
rect 35196 2540 35260 2604
rect 35402 2540 35466 2604
rect 35482 2540 35546 2604
rect 35562 2540 35626 2604
rect 35642 2540 35706 2604
rect 35722 2540 35786 2604
rect 35802 2540 35866 2604
rect 36008 2540 36072 2604
rect 36088 2540 36152 2604
rect 36168 2540 36232 2604
rect 36248 2540 36312 2604
rect 36328 2540 36392 2604
rect 36408 2540 36472 2604
rect 36614 2540 36678 2604
rect 36694 2540 36758 2604
rect 36774 2540 36838 2604
rect 36854 2540 36918 2604
rect 36934 2540 36998 2604
rect 37014 2540 37078 2604
rect 37220 2540 37284 2604
rect 37300 2540 37364 2604
rect 37380 2540 37444 2604
rect 37460 2540 37524 2604
rect 37540 2540 37604 2604
rect 37620 2540 37684 2604
rect 37826 2540 37890 2604
rect 37906 2540 37970 2604
rect 37986 2540 38050 2604
rect 38066 2540 38130 2604
rect 38146 2540 38210 2604
rect 38226 2540 38290 2604
rect 38432 2540 38496 2604
rect 38512 2540 38576 2604
rect 38592 2540 38656 2604
rect 38672 2540 38736 2604
rect 38752 2540 38816 2604
rect 38832 2540 38896 2604
rect 39038 2540 39102 2604
rect 39118 2540 39182 2604
rect 39198 2540 39262 2604
rect 39278 2540 39342 2604
rect 39358 2540 39422 2604
rect 39438 2540 39502 2604
rect -458 2320 -394 2384
rect -458 2240 -394 2304
rect -458 2160 -394 2224
rect -458 2080 -394 2144
rect -458 2000 -394 2064
rect -458 1920 -394 1984
rect -458 1840 -394 1904
rect -458 1760 -394 1824
rect -458 1680 -394 1744
rect -458 1600 -394 1664
rect 148 2320 212 2384
rect 148 2240 212 2304
rect 148 2160 212 2224
rect 148 2080 212 2144
rect 148 2000 212 2064
rect 148 1920 212 1984
rect 148 1840 212 1904
rect 148 1760 212 1824
rect 148 1680 212 1744
rect 148 1600 212 1664
rect 356 2320 420 2384
rect 356 2240 420 2304
rect 356 2160 420 2224
rect 356 2080 420 2144
rect 356 2000 420 2064
rect 356 1920 420 1984
rect 356 1840 420 1904
rect 356 1760 420 1824
rect 356 1680 420 1744
rect 356 1600 420 1664
rect 962 2461 1026 2465
rect 962 2405 966 2461
rect 966 2405 1022 2461
rect 1022 2405 1026 2461
rect 962 2401 1026 2405
rect 962 2320 1026 2384
rect 962 2240 1026 2304
rect 962 2160 1026 2224
rect 962 2080 1026 2144
rect 962 2000 1026 2064
rect 962 1920 1026 1984
rect 962 1840 1026 1904
rect 962 1760 1026 1824
rect 962 1680 1026 1744
rect 962 1600 1026 1664
rect -355 1380 -291 1444
rect -275 1380 -211 1444
rect -195 1380 -131 1444
rect -115 1380 -51 1444
rect -35 1380 29 1444
rect 45 1380 109 1444
rect 459 1380 523 1444
rect 539 1380 603 1444
rect 619 1380 683 1444
rect 699 1380 763 1444
rect 779 1380 843 1444
rect 859 1380 923 1444
rect -458 1160 -394 1224
rect -458 1080 -394 1144
rect -458 1000 -394 1064
rect -458 920 -394 984
rect -458 840 -394 904
rect -458 760 -394 824
rect -458 680 -394 744
rect -458 600 -394 664
rect -458 520 -394 584
rect -458 440 -394 504
rect 148 1160 212 1224
rect 148 1080 212 1144
rect 148 1000 212 1064
rect 148 920 212 984
rect 148 840 212 904
rect 148 760 212 824
rect 148 680 212 744
rect 148 600 212 664
rect 148 520 212 584
rect 148 440 212 504
rect 356 1160 420 1224
rect 356 1080 420 1144
rect 356 1000 420 1064
rect 356 920 420 984
rect 356 840 420 904
rect 356 760 420 824
rect 356 680 420 744
rect 356 600 420 664
rect 356 520 420 584
rect 356 440 420 504
rect 962 1160 1026 1224
rect 962 1080 1026 1144
rect 962 1000 1026 1064
rect 962 920 1026 984
rect 962 840 1026 904
rect 962 760 1026 824
rect 962 680 1026 744
rect 962 600 1026 664
rect 962 520 1026 584
rect 962 440 1026 504
rect 1268 2320 1332 2384
rect 1268 2240 1332 2304
rect 1268 2160 1332 2224
rect 1268 2080 1332 2144
rect 1268 2000 1332 2064
rect 1268 1920 1332 1984
rect 1268 1840 1332 1904
rect 1268 1760 1332 1824
rect 1268 1680 1332 1744
rect 1268 1600 1332 1664
rect 1874 2320 1938 2384
rect 1874 2240 1938 2304
rect 1874 2160 1938 2224
rect 1874 2080 1938 2144
rect 1874 2000 1938 2064
rect 1874 1920 1938 1984
rect 1874 1840 1938 1904
rect 1874 1760 1938 1824
rect 1874 1680 1938 1744
rect 1874 1600 1938 1664
rect 2480 2461 2544 2465
rect 2480 2405 2484 2461
rect 2484 2405 2540 2461
rect 2540 2405 2544 2461
rect 2480 2401 2544 2405
rect 2480 2320 2544 2384
rect 2480 2240 2544 2304
rect 2480 2160 2544 2224
rect 2480 2080 2544 2144
rect 2480 2000 2544 2064
rect 2480 1920 2544 1984
rect 2480 1840 2544 1904
rect 2480 1760 2544 1824
rect 2480 1680 2544 1744
rect 2480 1600 2544 1664
rect 1371 1380 1435 1444
rect 1451 1380 1515 1444
rect 1531 1380 1595 1444
rect 1611 1380 1675 1444
rect 1691 1380 1755 1444
rect 1771 1380 1835 1444
rect 1977 1380 2041 1444
rect 2057 1380 2121 1444
rect 2137 1380 2201 1444
rect 2217 1380 2281 1444
rect 2297 1380 2361 1444
rect 2377 1380 2441 1444
rect 1268 1160 1332 1224
rect 1268 1080 1332 1144
rect 1268 1000 1332 1064
rect 1268 920 1332 984
rect 1268 840 1332 904
rect 1268 760 1332 824
rect 1268 680 1332 744
rect 1268 600 1332 664
rect 1268 520 1332 584
rect 1268 440 1332 504
rect 1874 1160 1938 1224
rect 1874 1080 1938 1144
rect 1874 1000 1938 1064
rect 1874 920 1938 984
rect 1874 840 1938 904
rect 1874 760 1938 824
rect 1874 680 1938 744
rect 1874 600 1938 664
rect 1874 520 1938 584
rect 1874 440 1938 504
rect 2480 1160 2544 1224
rect 2480 1080 2544 1144
rect 2480 1000 2544 1064
rect 2480 920 2544 984
rect 2480 840 2544 904
rect 2480 760 2544 824
rect 2480 680 2544 744
rect 2480 600 2544 664
rect 2480 520 2544 584
rect 2480 440 2544 504
rect 2802 2320 2866 2384
rect 2802 2240 2866 2304
rect 2802 2160 2866 2224
rect 2802 2080 2866 2144
rect 2802 2000 2866 2064
rect 2802 1920 2866 1984
rect 2802 1840 2866 1904
rect 2802 1760 2866 1824
rect 2802 1680 2866 1744
rect 2802 1600 2866 1664
rect 3408 2320 3472 2384
rect 3408 2240 3472 2304
rect 3408 2160 3472 2224
rect 3408 2080 3472 2144
rect 3408 2000 3472 2064
rect 3408 1920 3472 1984
rect 3408 1840 3472 1904
rect 3408 1760 3472 1824
rect 3408 1680 3472 1744
rect 3408 1600 3472 1664
rect 4014 2320 4078 2384
rect 4014 2240 4078 2304
rect 4014 2160 4078 2224
rect 4014 2080 4078 2144
rect 4014 2000 4078 2064
rect 4014 1920 4078 1984
rect 4014 1840 4078 1904
rect 4014 1760 4078 1824
rect 4014 1680 4078 1744
rect 4014 1600 4078 1664
rect 4620 2320 4684 2384
rect 4620 2240 4684 2304
rect 4620 2160 4684 2224
rect 4620 2080 4684 2144
rect 4620 2000 4684 2064
rect 4620 1920 4684 1984
rect 4620 1840 4684 1904
rect 4620 1760 4684 1824
rect 4620 1680 4684 1744
rect 4620 1600 4684 1664
rect 5226 2320 5290 2384
rect 5226 2240 5290 2304
rect 5226 2160 5290 2224
rect 5226 2080 5290 2144
rect 5226 2000 5290 2064
rect 5226 1920 5290 1984
rect 5226 1840 5290 1904
rect 5226 1760 5290 1824
rect 5226 1680 5290 1744
rect 5226 1600 5290 1664
rect 2905 1380 2969 1444
rect 2985 1380 3049 1444
rect 3065 1380 3129 1444
rect 3145 1380 3209 1444
rect 3225 1380 3289 1444
rect 3305 1380 3369 1444
rect 3511 1380 3575 1444
rect 3591 1380 3655 1444
rect 3671 1380 3735 1444
rect 3751 1380 3815 1444
rect 3831 1380 3895 1444
rect 3911 1380 3975 1444
rect 4117 1380 4181 1444
rect 4197 1380 4261 1444
rect 4277 1380 4341 1444
rect 4357 1380 4421 1444
rect 4437 1380 4501 1444
rect 4517 1380 4581 1444
rect 4723 1380 4787 1444
rect 4803 1380 4867 1444
rect 4883 1380 4947 1444
rect 4963 1380 5027 1444
rect 5043 1380 5107 1444
rect 5123 1380 5187 1444
rect 2802 1160 2866 1224
rect 2802 1080 2866 1144
rect 2802 1000 2866 1064
rect 2802 920 2866 984
rect 2802 840 2866 904
rect 2802 760 2866 824
rect 2802 680 2866 744
rect 2802 600 2866 664
rect 2802 520 2866 584
rect 2802 440 2866 504
rect 3408 1160 3472 1224
rect 3408 1080 3472 1144
rect 3408 1000 3472 1064
rect 3408 920 3472 984
rect 3408 840 3472 904
rect 3408 760 3472 824
rect 3408 680 3472 744
rect 3408 600 3472 664
rect 3408 520 3472 584
rect 3408 440 3472 504
rect 4014 1160 4078 1224
rect 4014 1080 4078 1144
rect 4014 1000 4078 1064
rect 4014 920 4078 984
rect 4014 840 4078 904
rect 4014 760 4078 824
rect 4014 680 4078 744
rect 4014 600 4078 664
rect 4014 520 4078 584
rect 4014 440 4078 504
rect 4620 1160 4684 1224
rect 4620 1080 4684 1144
rect 4620 1000 4684 1064
rect 4620 920 4684 984
rect 4620 840 4684 904
rect 4620 760 4684 824
rect 4620 680 4684 744
rect 4620 600 4684 664
rect 4620 520 4684 584
rect 4620 440 4684 504
rect 5226 1160 5290 1224
rect 5226 1080 5290 1144
rect 5226 1000 5290 1064
rect 5226 920 5290 984
rect 5226 840 5290 904
rect 5226 760 5290 824
rect 5226 680 5290 744
rect 5226 600 5290 664
rect 5226 520 5290 584
rect 5226 440 5290 504
rect 5353 2320 5417 2384
rect 5353 2240 5417 2304
rect 5353 2160 5417 2224
rect 5353 2080 5417 2144
rect 5353 2000 5417 2064
rect 5353 1920 5417 1984
rect 5353 1840 5417 1904
rect 5353 1760 5417 1824
rect 5353 1680 5417 1744
rect 5353 1600 5417 1664
rect 5959 2320 6023 2384
rect 5959 2240 6023 2304
rect 5959 2160 6023 2224
rect 5959 2080 6023 2144
rect 5959 2000 6023 2064
rect 5959 1920 6023 1984
rect 5959 1840 6023 1904
rect 5959 1760 6023 1824
rect 5959 1680 6023 1744
rect 5959 1600 6023 1664
rect 6565 2320 6629 2384
rect 6565 2240 6629 2304
rect 6565 2160 6629 2224
rect 6565 2080 6629 2144
rect 6565 2000 6629 2064
rect 6565 1920 6629 1984
rect 6565 1840 6629 1904
rect 6565 1760 6629 1824
rect 6565 1680 6629 1744
rect 6565 1600 6629 1664
rect 7171 2320 7235 2384
rect 7171 2240 7235 2304
rect 7171 2160 7235 2224
rect 7171 2080 7235 2144
rect 7171 2000 7235 2064
rect 7171 1920 7235 1984
rect 7171 1840 7235 1904
rect 7171 1760 7235 1824
rect 7171 1680 7235 1744
rect 7171 1600 7235 1664
rect 7777 2320 7841 2384
rect 7777 2240 7841 2304
rect 7777 2160 7841 2224
rect 7777 2080 7841 2144
rect 7777 2000 7841 2064
rect 7777 1920 7841 1984
rect 7777 1840 7841 1904
rect 7777 1760 7841 1824
rect 7777 1680 7841 1744
rect 7777 1600 7841 1664
rect 8383 2320 8447 2384
rect 8383 2240 8447 2304
rect 8383 2160 8447 2224
rect 8383 2080 8447 2144
rect 8383 2000 8447 2064
rect 8383 1920 8447 1984
rect 8383 1840 8447 1904
rect 8383 1760 8447 1824
rect 8383 1680 8447 1744
rect 8383 1600 8447 1664
rect 8989 2320 9053 2384
rect 8989 2240 9053 2304
rect 8989 2160 9053 2224
rect 8989 2080 9053 2144
rect 8989 2000 9053 2064
rect 8989 1920 9053 1984
rect 8989 1840 9053 1904
rect 8989 1760 9053 1824
rect 8989 1680 9053 1744
rect 8989 1600 9053 1664
rect 9595 2320 9659 2384
rect 9595 2240 9659 2304
rect 9595 2160 9659 2224
rect 9595 2080 9659 2144
rect 9595 2000 9659 2064
rect 9595 1920 9659 1984
rect 9595 1840 9659 1904
rect 9595 1760 9659 1824
rect 9595 1680 9659 1744
rect 9595 1600 9659 1664
rect 10201 2320 10265 2384
rect 10201 2240 10265 2304
rect 10201 2160 10265 2224
rect 10201 2080 10265 2144
rect 10201 2000 10265 2064
rect 10201 1920 10265 1984
rect 10201 1840 10265 1904
rect 10201 1760 10265 1824
rect 10201 1680 10265 1744
rect 10201 1600 10265 1664
rect 5456 1380 5520 1444
rect 5536 1380 5600 1444
rect 5616 1380 5680 1444
rect 5696 1380 5760 1444
rect 5776 1380 5840 1444
rect 5856 1380 5920 1444
rect 6062 1380 6126 1444
rect 6142 1380 6206 1444
rect 6222 1380 6286 1444
rect 6302 1380 6366 1444
rect 6382 1380 6446 1444
rect 6462 1380 6526 1444
rect 6668 1380 6732 1444
rect 6748 1380 6812 1444
rect 6828 1380 6892 1444
rect 6908 1380 6972 1444
rect 6988 1380 7052 1444
rect 7068 1380 7132 1444
rect 7274 1380 7338 1444
rect 7354 1380 7418 1444
rect 7434 1380 7498 1444
rect 7514 1380 7578 1444
rect 7594 1380 7658 1444
rect 7674 1380 7738 1444
rect 7880 1380 7944 1444
rect 7960 1380 8024 1444
rect 8040 1380 8104 1444
rect 8120 1380 8184 1444
rect 8200 1380 8264 1444
rect 8280 1380 8344 1444
rect 8486 1380 8550 1444
rect 8566 1380 8630 1444
rect 8646 1380 8710 1444
rect 8726 1380 8790 1444
rect 8806 1380 8870 1444
rect 8886 1380 8950 1444
rect 9092 1380 9156 1444
rect 9172 1380 9236 1444
rect 9252 1380 9316 1444
rect 9332 1380 9396 1444
rect 9412 1380 9476 1444
rect 9492 1380 9556 1444
rect 9698 1380 9762 1444
rect 9778 1380 9842 1444
rect 9858 1380 9922 1444
rect 9938 1380 10002 1444
rect 10018 1380 10082 1444
rect 10098 1380 10162 1444
rect 5353 1160 5417 1224
rect 5353 1080 5417 1144
rect 5353 1000 5417 1064
rect 5353 920 5417 984
rect 5353 840 5417 904
rect 5353 760 5417 824
rect 5353 680 5417 744
rect 5353 600 5417 664
rect 5353 520 5417 584
rect 5353 440 5417 504
rect 5959 1160 6023 1224
rect 5959 1080 6023 1144
rect 5959 1000 6023 1064
rect 5959 920 6023 984
rect 5959 840 6023 904
rect 5959 760 6023 824
rect 5959 680 6023 744
rect 5959 600 6023 664
rect 5959 520 6023 584
rect 5959 440 6023 504
rect 6565 1160 6629 1224
rect 6565 1080 6629 1144
rect 6565 1000 6629 1064
rect 6565 920 6629 984
rect 6565 840 6629 904
rect 6565 760 6629 824
rect 6565 680 6629 744
rect 6565 600 6629 664
rect 6565 520 6629 584
rect 6565 440 6629 504
rect 7171 1160 7235 1224
rect 7171 1080 7235 1144
rect 7171 1000 7235 1064
rect 7171 920 7235 984
rect 7171 840 7235 904
rect 7171 760 7235 824
rect 7171 680 7235 744
rect 7171 600 7235 664
rect 7171 520 7235 584
rect 7171 440 7235 504
rect 7777 1160 7841 1224
rect 7777 1080 7841 1144
rect 7777 1000 7841 1064
rect 7777 920 7841 984
rect 7777 840 7841 904
rect 7777 760 7841 824
rect 7777 680 7841 744
rect 7777 600 7841 664
rect 7777 520 7841 584
rect 7777 440 7841 504
rect 8383 1160 8447 1224
rect 8383 1080 8447 1144
rect 8383 1000 8447 1064
rect 8383 920 8447 984
rect 8383 840 8447 904
rect 8383 760 8447 824
rect 8383 680 8447 744
rect 8383 600 8447 664
rect 8383 520 8447 584
rect 8383 440 8447 504
rect 8989 1160 9053 1224
rect 8989 1080 9053 1144
rect 8989 1000 9053 1064
rect 8989 920 9053 984
rect 8989 840 9053 904
rect 8989 760 9053 824
rect 8989 680 9053 744
rect 8989 600 9053 664
rect 8989 520 9053 584
rect 8989 440 9053 504
rect 9595 1160 9659 1224
rect 9595 1080 9659 1144
rect 9595 1000 9659 1064
rect 9595 920 9659 984
rect 9595 840 9659 904
rect 9595 760 9659 824
rect 9595 680 9659 744
rect 9595 600 9659 664
rect 9595 520 9659 584
rect 9595 440 9659 504
rect 10201 1160 10265 1224
rect 10201 1080 10265 1144
rect 10201 1000 10265 1064
rect 10201 920 10265 984
rect 10201 840 10265 904
rect 10201 760 10265 824
rect 10201 680 10265 744
rect 10201 600 10265 664
rect 10201 520 10265 584
rect 10201 440 10265 504
rect 10327 2320 10391 2384
rect 10327 2240 10391 2304
rect 10327 2160 10391 2224
rect 10327 2080 10391 2144
rect 10327 2000 10391 2064
rect 10327 1920 10391 1984
rect 10327 1840 10391 1904
rect 10327 1760 10391 1824
rect 10327 1680 10391 1744
rect 10327 1600 10391 1664
rect 10933 2320 10997 2384
rect 10933 2240 10997 2304
rect 10933 2160 10997 2224
rect 10933 2080 10997 2144
rect 10933 2000 10997 2064
rect 10933 1920 10997 1984
rect 10933 1840 10997 1904
rect 10933 1760 10997 1824
rect 10933 1680 10997 1744
rect 10933 1600 10997 1664
rect 11539 2320 11603 2384
rect 11539 2240 11603 2304
rect 11539 2160 11603 2224
rect 11539 2080 11603 2144
rect 11539 2000 11603 2064
rect 11539 1920 11603 1984
rect 11539 1840 11603 1904
rect 11539 1760 11603 1824
rect 11539 1680 11603 1744
rect 11539 1600 11603 1664
rect 12145 2320 12209 2384
rect 12145 2240 12209 2304
rect 12145 2160 12209 2224
rect 12145 2080 12209 2144
rect 12145 2000 12209 2064
rect 12145 1920 12209 1984
rect 12145 1840 12209 1904
rect 12145 1760 12209 1824
rect 12145 1680 12209 1744
rect 12145 1600 12209 1664
rect 12751 2320 12815 2384
rect 12751 2240 12815 2304
rect 12751 2160 12815 2224
rect 12751 2080 12815 2144
rect 12751 2000 12815 2064
rect 12751 1920 12815 1984
rect 12751 1840 12815 1904
rect 12751 1760 12815 1824
rect 12751 1680 12815 1744
rect 12751 1600 12815 1664
rect 13357 2320 13421 2384
rect 13357 2240 13421 2304
rect 13357 2160 13421 2224
rect 13357 2080 13421 2144
rect 13357 2000 13421 2064
rect 13357 1920 13421 1984
rect 13357 1840 13421 1904
rect 13357 1760 13421 1824
rect 13357 1680 13421 1744
rect 13357 1600 13421 1664
rect 13963 2320 14027 2384
rect 13963 2240 14027 2304
rect 13963 2160 14027 2224
rect 13963 2080 14027 2144
rect 13963 2000 14027 2064
rect 13963 1920 14027 1984
rect 13963 1840 14027 1904
rect 13963 1760 14027 1824
rect 13963 1680 14027 1744
rect 13963 1600 14027 1664
rect 14569 2320 14633 2384
rect 14569 2240 14633 2304
rect 14569 2160 14633 2224
rect 14569 2080 14633 2144
rect 14569 2000 14633 2064
rect 14569 1920 14633 1984
rect 14569 1840 14633 1904
rect 14569 1760 14633 1824
rect 14569 1680 14633 1744
rect 14569 1600 14633 1664
rect 15175 2320 15239 2384
rect 15175 2240 15239 2304
rect 15175 2160 15239 2224
rect 15175 2080 15239 2144
rect 15175 2000 15239 2064
rect 15175 1920 15239 1984
rect 15175 1840 15239 1904
rect 15175 1760 15239 1824
rect 15175 1680 15239 1744
rect 15175 1600 15239 1664
rect 15781 2320 15845 2384
rect 15781 2240 15845 2304
rect 15781 2160 15845 2224
rect 15781 2080 15845 2144
rect 15781 2000 15845 2064
rect 15781 1920 15845 1984
rect 15781 1840 15845 1904
rect 15781 1760 15845 1824
rect 15781 1680 15845 1744
rect 15781 1600 15845 1664
rect 16387 2320 16451 2384
rect 16387 2240 16451 2304
rect 16387 2160 16451 2224
rect 16387 2080 16451 2144
rect 16387 2000 16451 2064
rect 16387 1920 16451 1984
rect 16387 1840 16451 1904
rect 16387 1760 16451 1824
rect 16387 1680 16451 1744
rect 16387 1600 16451 1664
rect 16993 2320 17057 2384
rect 16993 2240 17057 2304
rect 16993 2160 17057 2224
rect 16993 2080 17057 2144
rect 16993 2000 17057 2064
rect 16993 1920 17057 1984
rect 16993 1840 17057 1904
rect 16993 1760 17057 1824
rect 16993 1680 17057 1744
rect 16993 1600 17057 1664
rect 17599 2320 17663 2384
rect 17599 2240 17663 2304
rect 17599 2160 17663 2224
rect 17599 2080 17663 2144
rect 17599 2000 17663 2064
rect 17599 1920 17663 1984
rect 17599 1840 17663 1904
rect 17599 1760 17663 1824
rect 17599 1680 17663 1744
rect 17599 1600 17663 1664
rect 18205 2320 18269 2384
rect 18205 2240 18269 2304
rect 18205 2160 18269 2224
rect 18205 2080 18269 2144
rect 18205 2000 18269 2064
rect 18205 1920 18269 1984
rect 18205 1840 18269 1904
rect 18205 1760 18269 1824
rect 18205 1680 18269 1744
rect 18205 1600 18269 1664
rect 18811 2320 18875 2384
rect 18811 2240 18875 2304
rect 18811 2160 18875 2224
rect 18811 2080 18875 2144
rect 18811 2000 18875 2064
rect 18811 1920 18875 1984
rect 18811 1840 18875 1904
rect 18811 1760 18875 1824
rect 18811 1680 18875 1744
rect 18811 1600 18875 1664
rect 19417 2320 19481 2384
rect 19417 2240 19481 2304
rect 19417 2160 19481 2224
rect 19417 2080 19481 2144
rect 19417 2000 19481 2064
rect 19417 1920 19481 1984
rect 19417 1840 19481 1904
rect 19417 1760 19481 1824
rect 19417 1680 19481 1744
rect 19417 1600 19481 1664
rect 20023 2320 20087 2384
rect 20023 2240 20087 2304
rect 20023 2160 20087 2224
rect 20023 2080 20087 2144
rect 20023 2000 20087 2064
rect 20023 1920 20087 1984
rect 20023 1840 20087 1904
rect 20023 1760 20087 1824
rect 20023 1680 20087 1744
rect 20023 1600 20087 1664
rect 10430 1380 10494 1444
rect 10510 1380 10574 1444
rect 10590 1380 10654 1444
rect 10670 1380 10734 1444
rect 10750 1380 10814 1444
rect 10830 1380 10894 1444
rect 11036 1380 11100 1444
rect 11116 1380 11180 1444
rect 11196 1380 11260 1444
rect 11276 1380 11340 1444
rect 11356 1380 11420 1444
rect 11436 1380 11500 1444
rect 11642 1380 11706 1444
rect 11722 1380 11786 1444
rect 11802 1380 11866 1444
rect 11882 1380 11946 1444
rect 11962 1380 12026 1444
rect 12042 1380 12106 1444
rect 12248 1380 12312 1444
rect 12328 1380 12392 1444
rect 12408 1380 12472 1444
rect 12488 1380 12552 1444
rect 12568 1380 12632 1444
rect 12648 1380 12712 1444
rect 12854 1380 12918 1444
rect 12934 1380 12998 1444
rect 13014 1380 13078 1444
rect 13094 1380 13158 1444
rect 13174 1380 13238 1444
rect 13254 1380 13318 1444
rect 13460 1380 13524 1444
rect 13540 1380 13604 1444
rect 13620 1380 13684 1444
rect 13700 1380 13764 1444
rect 13780 1380 13844 1444
rect 13860 1380 13924 1444
rect 14066 1380 14130 1444
rect 14146 1380 14210 1444
rect 14226 1380 14290 1444
rect 14306 1380 14370 1444
rect 14386 1380 14450 1444
rect 14466 1380 14530 1444
rect 14672 1380 14736 1444
rect 14752 1380 14816 1444
rect 14832 1380 14896 1444
rect 14912 1380 14976 1444
rect 14992 1380 15056 1444
rect 15072 1380 15136 1444
rect 15278 1380 15342 1444
rect 15358 1380 15422 1444
rect 15438 1380 15502 1444
rect 15518 1380 15582 1444
rect 15598 1380 15662 1444
rect 15678 1380 15742 1444
rect 15884 1380 15948 1444
rect 15964 1380 16028 1444
rect 16044 1380 16108 1444
rect 16124 1380 16188 1444
rect 16204 1380 16268 1444
rect 16284 1380 16348 1444
rect 16490 1380 16554 1444
rect 16570 1380 16634 1444
rect 16650 1380 16714 1444
rect 16730 1380 16794 1444
rect 16810 1380 16874 1444
rect 16890 1380 16954 1444
rect 17096 1380 17160 1444
rect 17176 1380 17240 1444
rect 17256 1380 17320 1444
rect 17336 1380 17400 1444
rect 17416 1380 17480 1444
rect 17496 1380 17560 1444
rect 17702 1380 17766 1444
rect 17782 1380 17846 1444
rect 17862 1380 17926 1444
rect 17942 1380 18006 1444
rect 18022 1380 18086 1444
rect 18102 1380 18166 1444
rect 18308 1380 18372 1444
rect 18388 1380 18452 1444
rect 18468 1380 18532 1444
rect 18548 1380 18612 1444
rect 18628 1380 18692 1444
rect 18708 1380 18772 1444
rect 18914 1380 18978 1444
rect 18994 1380 19058 1444
rect 19074 1380 19138 1444
rect 19154 1380 19218 1444
rect 19234 1380 19298 1444
rect 19314 1380 19378 1444
rect 19520 1380 19584 1444
rect 19600 1380 19664 1444
rect 19680 1380 19744 1444
rect 19760 1380 19824 1444
rect 19840 1380 19904 1444
rect 19920 1380 19984 1444
rect 10327 1160 10391 1224
rect 10327 1080 10391 1144
rect 10327 1000 10391 1064
rect 10327 920 10391 984
rect 10327 840 10391 904
rect 10327 760 10391 824
rect 10327 680 10391 744
rect 10327 600 10391 664
rect 10327 520 10391 584
rect 10327 440 10391 504
rect 10933 1160 10997 1224
rect 10933 1080 10997 1144
rect 10933 1000 10997 1064
rect 10933 920 10997 984
rect 10933 840 10997 904
rect 10933 760 10997 824
rect 10933 680 10997 744
rect 10933 600 10997 664
rect 10933 520 10997 584
rect 10933 440 10997 504
rect 11539 1160 11603 1224
rect 11539 1080 11603 1144
rect 11539 1000 11603 1064
rect 11539 920 11603 984
rect 11539 840 11603 904
rect 11539 760 11603 824
rect 11539 680 11603 744
rect 11539 600 11603 664
rect 11539 520 11603 584
rect 11539 440 11603 504
rect 12145 1160 12209 1224
rect 12145 1080 12209 1144
rect 12145 1000 12209 1064
rect 12145 920 12209 984
rect 12145 840 12209 904
rect 12145 760 12209 824
rect 12145 680 12209 744
rect 12145 600 12209 664
rect 12145 520 12209 584
rect 12145 440 12209 504
rect 12751 1160 12815 1224
rect 12751 1080 12815 1144
rect 12751 1000 12815 1064
rect 12751 920 12815 984
rect 12751 840 12815 904
rect 12751 760 12815 824
rect 12751 680 12815 744
rect 12751 600 12815 664
rect 12751 520 12815 584
rect 12751 440 12815 504
rect 13357 1160 13421 1224
rect 13357 1080 13421 1144
rect 13357 1000 13421 1064
rect 13357 920 13421 984
rect 13357 840 13421 904
rect 13357 760 13421 824
rect 13357 680 13421 744
rect 13357 600 13421 664
rect 13357 520 13421 584
rect 13357 440 13421 504
rect 13963 1160 14027 1224
rect 13963 1080 14027 1144
rect 13963 1000 14027 1064
rect 13963 920 14027 984
rect 13963 840 14027 904
rect 13963 760 14027 824
rect 13963 680 14027 744
rect 13963 600 14027 664
rect 13963 520 14027 584
rect 13963 440 14027 504
rect 14569 1160 14633 1224
rect 14569 1080 14633 1144
rect 14569 1000 14633 1064
rect 14569 920 14633 984
rect 14569 840 14633 904
rect 14569 760 14633 824
rect 14569 680 14633 744
rect 14569 600 14633 664
rect 14569 520 14633 584
rect 14569 440 14633 504
rect 15175 1160 15239 1224
rect 15175 1080 15239 1144
rect 15175 1000 15239 1064
rect 15175 920 15239 984
rect 15175 840 15239 904
rect 15175 760 15239 824
rect 15175 680 15239 744
rect 15175 600 15239 664
rect 15175 520 15239 584
rect 15175 440 15239 504
rect 15781 1160 15845 1224
rect 15781 1080 15845 1144
rect 15781 1000 15845 1064
rect 15781 920 15845 984
rect 15781 840 15845 904
rect 15781 760 15845 824
rect 15781 680 15845 744
rect 15781 600 15845 664
rect 15781 520 15845 584
rect 15781 440 15845 504
rect 16387 1160 16451 1224
rect 16387 1080 16451 1144
rect 16387 1000 16451 1064
rect 16387 920 16451 984
rect 16387 840 16451 904
rect 16387 760 16451 824
rect 16387 680 16451 744
rect 16387 600 16451 664
rect 16387 520 16451 584
rect 16387 440 16451 504
rect 16993 1160 17057 1224
rect 16993 1080 17057 1144
rect 16993 1000 17057 1064
rect 16993 920 17057 984
rect 16993 840 17057 904
rect 16993 760 17057 824
rect 16993 680 17057 744
rect 16993 600 17057 664
rect 16993 520 17057 584
rect 16993 440 17057 504
rect 17599 1160 17663 1224
rect 17599 1080 17663 1144
rect 17599 1000 17663 1064
rect 17599 920 17663 984
rect 17599 840 17663 904
rect 17599 760 17663 824
rect 17599 680 17663 744
rect 17599 600 17663 664
rect 17599 520 17663 584
rect 17599 440 17663 504
rect 18205 1160 18269 1224
rect 18205 1080 18269 1144
rect 18205 1000 18269 1064
rect 18205 920 18269 984
rect 18205 840 18269 904
rect 18205 760 18269 824
rect 18205 680 18269 744
rect 18205 600 18269 664
rect 18205 520 18269 584
rect 18205 440 18269 504
rect 18811 1160 18875 1224
rect 18811 1080 18875 1144
rect 18811 1000 18875 1064
rect 18811 920 18875 984
rect 18811 840 18875 904
rect 18811 760 18875 824
rect 18811 680 18875 744
rect 18811 600 18875 664
rect 18811 520 18875 584
rect 18811 440 18875 504
rect 19417 1160 19481 1224
rect 19417 1080 19481 1144
rect 19417 1000 19481 1064
rect 19417 920 19481 984
rect 19417 840 19481 904
rect 19417 760 19481 824
rect 19417 680 19481 744
rect 19417 600 19481 664
rect 19417 520 19481 584
rect 19417 440 19481 504
rect 20023 1160 20087 1224
rect 20023 1080 20087 1144
rect 20023 1000 20087 1064
rect 20023 920 20087 984
rect 20023 840 20087 904
rect 20023 760 20087 824
rect 20023 680 20087 744
rect 20023 600 20087 664
rect 20023 520 20087 584
rect 20023 440 20087 504
rect 20149 2320 20213 2384
rect 20149 2240 20213 2304
rect 20149 2160 20213 2224
rect 20149 2080 20213 2144
rect 20149 2000 20213 2064
rect 20149 1920 20213 1984
rect 20149 1840 20213 1904
rect 20149 1760 20213 1824
rect 20149 1680 20213 1744
rect 20149 1600 20213 1664
rect 20755 2320 20819 2384
rect 20755 2240 20819 2304
rect 20755 2160 20819 2224
rect 20755 2080 20819 2144
rect 20755 2000 20819 2064
rect 20755 1920 20819 1984
rect 20755 1840 20819 1904
rect 20755 1760 20819 1824
rect 20755 1680 20819 1744
rect 20755 1600 20819 1664
rect 21361 2320 21425 2384
rect 21361 2240 21425 2304
rect 21361 2160 21425 2224
rect 21361 2080 21425 2144
rect 21361 2000 21425 2064
rect 21361 1920 21425 1984
rect 21361 1840 21425 1904
rect 21361 1760 21425 1824
rect 21361 1680 21425 1744
rect 21361 1600 21425 1664
rect 21967 2320 22031 2384
rect 21967 2240 22031 2304
rect 21967 2160 22031 2224
rect 21967 2080 22031 2144
rect 21967 2000 22031 2064
rect 21967 1920 22031 1984
rect 21967 1840 22031 1904
rect 21967 1760 22031 1824
rect 21967 1680 22031 1744
rect 21967 1600 22031 1664
rect 22573 2320 22637 2384
rect 22573 2240 22637 2304
rect 22573 2160 22637 2224
rect 22573 2080 22637 2144
rect 22573 2000 22637 2064
rect 22573 1920 22637 1984
rect 22573 1840 22637 1904
rect 22573 1760 22637 1824
rect 22573 1680 22637 1744
rect 22573 1600 22637 1664
rect 23179 2320 23243 2384
rect 23179 2240 23243 2304
rect 23179 2160 23243 2224
rect 23179 2080 23243 2144
rect 23179 2000 23243 2064
rect 23179 1920 23243 1984
rect 23179 1840 23243 1904
rect 23179 1760 23243 1824
rect 23179 1680 23243 1744
rect 23179 1600 23243 1664
rect 23785 2320 23849 2384
rect 23785 2240 23849 2304
rect 23785 2160 23849 2224
rect 23785 2080 23849 2144
rect 23785 2000 23849 2064
rect 23785 1920 23849 1984
rect 23785 1840 23849 1904
rect 23785 1760 23849 1824
rect 23785 1680 23849 1744
rect 23785 1600 23849 1664
rect 24391 2320 24455 2384
rect 24391 2240 24455 2304
rect 24391 2160 24455 2224
rect 24391 2080 24455 2144
rect 24391 2000 24455 2064
rect 24391 1920 24455 1984
rect 24391 1840 24455 1904
rect 24391 1760 24455 1824
rect 24391 1680 24455 1744
rect 24391 1600 24455 1664
rect 24997 2320 25061 2384
rect 24997 2240 25061 2304
rect 24997 2160 25061 2224
rect 24997 2080 25061 2144
rect 24997 2000 25061 2064
rect 24997 1920 25061 1984
rect 24997 1840 25061 1904
rect 24997 1760 25061 1824
rect 24997 1680 25061 1744
rect 24997 1600 25061 1664
rect 25603 2320 25667 2384
rect 25603 2240 25667 2304
rect 25603 2160 25667 2224
rect 25603 2080 25667 2144
rect 25603 2000 25667 2064
rect 25603 1920 25667 1984
rect 25603 1840 25667 1904
rect 25603 1760 25667 1824
rect 25603 1680 25667 1744
rect 25603 1600 25667 1664
rect 26209 2320 26273 2384
rect 26209 2240 26273 2304
rect 26209 2160 26273 2224
rect 26209 2080 26273 2144
rect 26209 2000 26273 2064
rect 26209 1920 26273 1984
rect 26209 1840 26273 1904
rect 26209 1760 26273 1824
rect 26209 1680 26273 1744
rect 26209 1600 26273 1664
rect 26815 2320 26879 2384
rect 26815 2240 26879 2304
rect 26815 2160 26879 2224
rect 26815 2080 26879 2144
rect 26815 2000 26879 2064
rect 26815 1920 26879 1984
rect 26815 1840 26879 1904
rect 26815 1760 26879 1824
rect 26815 1680 26879 1744
rect 26815 1600 26879 1664
rect 27421 2320 27485 2384
rect 27421 2240 27485 2304
rect 27421 2160 27485 2224
rect 27421 2080 27485 2144
rect 27421 2000 27485 2064
rect 27421 1920 27485 1984
rect 27421 1840 27485 1904
rect 27421 1760 27485 1824
rect 27421 1680 27485 1744
rect 27421 1600 27485 1664
rect 28027 2320 28091 2384
rect 28027 2240 28091 2304
rect 28027 2160 28091 2224
rect 28027 2080 28091 2144
rect 28027 2000 28091 2064
rect 28027 1920 28091 1984
rect 28027 1840 28091 1904
rect 28027 1760 28091 1824
rect 28027 1680 28091 1744
rect 28027 1600 28091 1664
rect 28633 2320 28697 2384
rect 28633 2240 28697 2304
rect 28633 2160 28697 2224
rect 28633 2080 28697 2144
rect 28633 2000 28697 2064
rect 28633 1920 28697 1984
rect 28633 1840 28697 1904
rect 28633 1760 28697 1824
rect 28633 1680 28697 1744
rect 28633 1600 28697 1664
rect 29239 2320 29303 2384
rect 29239 2240 29303 2304
rect 29239 2160 29303 2224
rect 29239 2080 29303 2144
rect 29239 2000 29303 2064
rect 29239 1920 29303 1984
rect 29239 1840 29303 1904
rect 29239 1760 29303 1824
rect 29239 1680 29303 1744
rect 29239 1600 29303 1664
rect 29845 2320 29909 2384
rect 29845 2240 29909 2304
rect 29845 2160 29909 2224
rect 29845 2080 29909 2144
rect 29845 2000 29909 2064
rect 29845 1920 29909 1984
rect 29845 1840 29909 1904
rect 29845 1760 29909 1824
rect 29845 1680 29909 1744
rect 29845 1600 29909 1664
rect 30451 2320 30515 2384
rect 30451 2240 30515 2304
rect 30451 2160 30515 2224
rect 30451 2080 30515 2144
rect 30451 2000 30515 2064
rect 30451 1920 30515 1984
rect 30451 1840 30515 1904
rect 30451 1760 30515 1824
rect 30451 1680 30515 1744
rect 30451 1600 30515 1664
rect 31057 2320 31121 2384
rect 31057 2240 31121 2304
rect 31057 2160 31121 2224
rect 31057 2080 31121 2144
rect 31057 2000 31121 2064
rect 31057 1920 31121 1984
rect 31057 1840 31121 1904
rect 31057 1760 31121 1824
rect 31057 1680 31121 1744
rect 31057 1600 31121 1664
rect 31663 2320 31727 2384
rect 31663 2240 31727 2304
rect 31663 2160 31727 2224
rect 31663 2080 31727 2144
rect 31663 2000 31727 2064
rect 31663 1920 31727 1984
rect 31663 1840 31727 1904
rect 31663 1760 31727 1824
rect 31663 1680 31727 1744
rect 31663 1600 31727 1664
rect 32269 2320 32333 2384
rect 32269 2240 32333 2304
rect 32269 2160 32333 2224
rect 32269 2080 32333 2144
rect 32269 2000 32333 2064
rect 32269 1920 32333 1984
rect 32269 1840 32333 1904
rect 32269 1760 32333 1824
rect 32269 1680 32333 1744
rect 32269 1600 32333 1664
rect 32875 2320 32939 2384
rect 32875 2240 32939 2304
rect 32875 2160 32939 2224
rect 32875 2080 32939 2144
rect 32875 2000 32939 2064
rect 32875 1920 32939 1984
rect 32875 1840 32939 1904
rect 32875 1760 32939 1824
rect 32875 1680 32939 1744
rect 32875 1600 32939 1664
rect 33481 2320 33545 2384
rect 33481 2240 33545 2304
rect 33481 2160 33545 2224
rect 33481 2080 33545 2144
rect 33481 2000 33545 2064
rect 33481 1920 33545 1984
rect 33481 1840 33545 1904
rect 33481 1760 33545 1824
rect 33481 1680 33545 1744
rect 33481 1600 33545 1664
rect 34087 2320 34151 2384
rect 34087 2240 34151 2304
rect 34087 2160 34151 2224
rect 34087 2080 34151 2144
rect 34087 2000 34151 2064
rect 34087 1920 34151 1984
rect 34087 1840 34151 1904
rect 34087 1760 34151 1824
rect 34087 1680 34151 1744
rect 34087 1600 34151 1664
rect 34693 2320 34757 2384
rect 34693 2240 34757 2304
rect 34693 2160 34757 2224
rect 34693 2080 34757 2144
rect 34693 2000 34757 2064
rect 34693 1920 34757 1984
rect 34693 1840 34757 1904
rect 34693 1760 34757 1824
rect 34693 1680 34757 1744
rect 34693 1600 34757 1664
rect 35299 2320 35363 2384
rect 35299 2240 35363 2304
rect 35299 2160 35363 2224
rect 35299 2080 35363 2144
rect 35299 2000 35363 2064
rect 35299 1920 35363 1984
rect 35299 1840 35363 1904
rect 35299 1760 35363 1824
rect 35299 1680 35363 1744
rect 35299 1600 35363 1664
rect 35905 2320 35969 2384
rect 35905 2240 35969 2304
rect 35905 2160 35969 2224
rect 35905 2080 35969 2144
rect 35905 2000 35969 2064
rect 35905 1920 35969 1984
rect 35905 1840 35969 1904
rect 35905 1760 35969 1824
rect 35905 1680 35969 1744
rect 35905 1600 35969 1664
rect 36511 2320 36575 2384
rect 36511 2240 36575 2304
rect 36511 2160 36575 2224
rect 36511 2080 36575 2144
rect 36511 2000 36575 2064
rect 36511 1920 36575 1984
rect 36511 1840 36575 1904
rect 36511 1760 36575 1824
rect 36511 1680 36575 1744
rect 36511 1600 36575 1664
rect 37117 2320 37181 2384
rect 37117 2240 37181 2304
rect 37117 2160 37181 2224
rect 37117 2080 37181 2144
rect 37117 2000 37181 2064
rect 37117 1920 37181 1984
rect 37117 1840 37181 1904
rect 37117 1760 37181 1824
rect 37117 1680 37181 1744
rect 37117 1600 37181 1664
rect 37723 2320 37787 2384
rect 37723 2240 37787 2304
rect 37723 2160 37787 2224
rect 37723 2080 37787 2144
rect 37723 2000 37787 2064
rect 37723 1920 37787 1984
rect 37723 1840 37787 1904
rect 37723 1760 37787 1824
rect 37723 1680 37787 1744
rect 37723 1600 37787 1664
rect 38329 2320 38393 2384
rect 38329 2240 38393 2304
rect 38329 2160 38393 2224
rect 38329 2080 38393 2144
rect 38329 2000 38393 2064
rect 38329 1920 38393 1984
rect 38329 1840 38393 1904
rect 38329 1760 38393 1824
rect 38329 1680 38393 1744
rect 38329 1600 38393 1664
rect 38935 2320 38999 2384
rect 38935 2240 38999 2304
rect 38935 2160 38999 2224
rect 38935 2080 38999 2144
rect 38935 2000 38999 2064
rect 38935 1920 38999 1984
rect 38935 1840 38999 1904
rect 38935 1760 38999 1824
rect 38935 1680 38999 1744
rect 38935 1600 38999 1664
rect 39541 2320 39605 2384
rect 39541 2240 39605 2304
rect 39541 2160 39605 2224
rect 39541 2080 39605 2144
rect 39541 2000 39605 2064
rect 39541 1920 39605 1984
rect 39541 1840 39605 1904
rect 39541 1760 39605 1824
rect 39541 1680 39605 1744
rect 39541 1600 39605 1664
rect 20252 1380 20316 1444
rect 20332 1380 20396 1444
rect 20412 1380 20476 1444
rect 20492 1380 20556 1444
rect 20572 1380 20636 1444
rect 20652 1380 20716 1444
rect 20858 1380 20922 1444
rect 20938 1380 21002 1444
rect 21018 1380 21082 1444
rect 21098 1380 21162 1444
rect 21178 1380 21242 1444
rect 21258 1380 21322 1444
rect 21464 1380 21528 1444
rect 21544 1380 21608 1444
rect 21624 1380 21688 1444
rect 21704 1380 21768 1444
rect 21784 1380 21848 1444
rect 21864 1380 21928 1444
rect 22070 1380 22134 1444
rect 22150 1380 22214 1444
rect 22230 1380 22294 1444
rect 22310 1380 22374 1444
rect 22390 1380 22454 1444
rect 22470 1380 22534 1444
rect 22676 1380 22740 1444
rect 22756 1380 22820 1444
rect 22836 1380 22900 1444
rect 22916 1380 22980 1444
rect 22996 1380 23060 1444
rect 23076 1380 23140 1444
rect 23282 1380 23346 1444
rect 23362 1380 23426 1444
rect 23442 1380 23506 1444
rect 23522 1380 23586 1444
rect 23602 1380 23666 1444
rect 23682 1380 23746 1444
rect 23888 1380 23952 1444
rect 23968 1380 24032 1444
rect 24048 1380 24112 1444
rect 24128 1380 24192 1444
rect 24208 1380 24272 1444
rect 24288 1380 24352 1444
rect 24494 1380 24558 1444
rect 24574 1380 24638 1444
rect 24654 1380 24718 1444
rect 24734 1380 24798 1444
rect 24814 1380 24878 1444
rect 24894 1380 24958 1444
rect 25100 1380 25164 1444
rect 25180 1380 25244 1444
rect 25260 1380 25324 1444
rect 25340 1380 25404 1444
rect 25420 1380 25484 1444
rect 25500 1380 25564 1444
rect 25706 1380 25770 1444
rect 25786 1380 25850 1444
rect 25866 1380 25930 1444
rect 25946 1380 26010 1444
rect 26026 1380 26090 1444
rect 26106 1380 26170 1444
rect 26312 1380 26376 1444
rect 26392 1380 26456 1444
rect 26472 1380 26536 1444
rect 26552 1380 26616 1444
rect 26632 1380 26696 1444
rect 26712 1380 26776 1444
rect 26918 1380 26982 1444
rect 26998 1380 27062 1444
rect 27078 1380 27142 1444
rect 27158 1380 27222 1444
rect 27238 1380 27302 1444
rect 27318 1380 27382 1444
rect 27524 1380 27588 1444
rect 27604 1380 27668 1444
rect 27684 1380 27748 1444
rect 27764 1380 27828 1444
rect 27844 1380 27908 1444
rect 27924 1380 27988 1444
rect 28130 1380 28194 1444
rect 28210 1380 28274 1444
rect 28290 1380 28354 1444
rect 28370 1380 28434 1444
rect 28450 1380 28514 1444
rect 28530 1380 28594 1444
rect 28736 1380 28800 1444
rect 28816 1380 28880 1444
rect 28896 1380 28960 1444
rect 28976 1380 29040 1444
rect 29056 1380 29120 1444
rect 29136 1380 29200 1444
rect 29342 1380 29406 1444
rect 29422 1380 29486 1444
rect 29502 1380 29566 1444
rect 29582 1380 29646 1444
rect 29662 1380 29726 1444
rect 29742 1380 29806 1444
rect 29948 1380 30012 1444
rect 30028 1380 30092 1444
rect 30108 1380 30172 1444
rect 30188 1380 30252 1444
rect 30268 1380 30332 1444
rect 30348 1380 30412 1444
rect 30554 1380 30618 1444
rect 30634 1380 30698 1444
rect 30714 1380 30778 1444
rect 30794 1380 30858 1444
rect 30874 1380 30938 1444
rect 30954 1380 31018 1444
rect 31160 1380 31224 1444
rect 31240 1380 31304 1444
rect 31320 1380 31384 1444
rect 31400 1380 31464 1444
rect 31480 1380 31544 1444
rect 31560 1380 31624 1444
rect 31766 1380 31830 1444
rect 31846 1380 31910 1444
rect 31926 1380 31990 1444
rect 32006 1380 32070 1444
rect 32086 1380 32150 1444
rect 32166 1380 32230 1444
rect 32372 1380 32436 1444
rect 32452 1380 32516 1444
rect 32532 1380 32596 1444
rect 32612 1380 32676 1444
rect 32692 1380 32756 1444
rect 32772 1380 32836 1444
rect 32978 1380 33042 1444
rect 33058 1380 33122 1444
rect 33138 1380 33202 1444
rect 33218 1380 33282 1444
rect 33298 1380 33362 1444
rect 33378 1380 33442 1444
rect 33584 1380 33648 1444
rect 33664 1380 33728 1444
rect 33744 1380 33808 1444
rect 33824 1380 33888 1444
rect 33904 1380 33968 1444
rect 33984 1380 34048 1444
rect 34190 1380 34254 1444
rect 34270 1380 34334 1444
rect 34350 1380 34414 1444
rect 34430 1380 34494 1444
rect 34510 1380 34574 1444
rect 34590 1380 34654 1444
rect 34796 1380 34860 1444
rect 34876 1380 34940 1444
rect 34956 1380 35020 1444
rect 35036 1380 35100 1444
rect 35116 1380 35180 1444
rect 35196 1380 35260 1444
rect 35402 1380 35466 1444
rect 35482 1380 35546 1444
rect 35562 1380 35626 1444
rect 35642 1380 35706 1444
rect 35722 1380 35786 1444
rect 35802 1380 35866 1444
rect 36008 1380 36072 1444
rect 36088 1380 36152 1444
rect 36168 1380 36232 1444
rect 36248 1380 36312 1444
rect 36328 1380 36392 1444
rect 36408 1380 36472 1444
rect 36614 1380 36678 1444
rect 36694 1380 36758 1444
rect 36774 1380 36838 1444
rect 36854 1380 36918 1444
rect 36934 1380 36998 1444
rect 37014 1380 37078 1444
rect 37220 1380 37284 1444
rect 37300 1380 37364 1444
rect 37380 1380 37444 1444
rect 37460 1380 37524 1444
rect 37540 1380 37604 1444
rect 37620 1380 37684 1444
rect 37826 1380 37890 1444
rect 37906 1380 37970 1444
rect 37986 1380 38050 1444
rect 38066 1380 38130 1444
rect 38146 1380 38210 1444
rect 38226 1380 38290 1444
rect 38432 1380 38496 1444
rect 38512 1380 38576 1444
rect 38592 1380 38656 1444
rect 38672 1380 38736 1444
rect 38752 1380 38816 1444
rect 38832 1380 38896 1444
rect 39038 1380 39102 1444
rect 39118 1380 39182 1444
rect 39198 1380 39262 1444
rect 39278 1380 39342 1444
rect 39358 1380 39422 1444
rect 39438 1380 39502 1444
rect 20149 1160 20213 1224
rect 20149 1080 20213 1144
rect 20149 1000 20213 1064
rect 20149 920 20213 984
rect 20149 840 20213 904
rect 20149 760 20213 824
rect 20149 680 20213 744
rect 20149 600 20213 664
rect 20149 520 20213 584
rect 20149 440 20213 504
rect 20755 1160 20819 1224
rect 20755 1080 20819 1144
rect 20755 1000 20819 1064
rect 20755 920 20819 984
rect 20755 840 20819 904
rect 20755 760 20819 824
rect 20755 680 20819 744
rect 20755 600 20819 664
rect 20755 520 20819 584
rect 20755 440 20819 504
rect 21361 1160 21425 1224
rect 21361 1080 21425 1144
rect 21361 1000 21425 1064
rect 21361 920 21425 984
rect 21361 840 21425 904
rect 21361 760 21425 824
rect 21361 680 21425 744
rect 21361 600 21425 664
rect 21361 520 21425 584
rect 21361 440 21425 504
rect 21967 1160 22031 1224
rect 21967 1080 22031 1144
rect 21967 1000 22031 1064
rect 21967 920 22031 984
rect 21967 840 22031 904
rect 21967 760 22031 824
rect 21967 680 22031 744
rect 21967 600 22031 664
rect 21967 520 22031 584
rect 21967 440 22031 504
rect 22573 1160 22637 1224
rect 22573 1080 22637 1144
rect 22573 1000 22637 1064
rect 22573 920 22637 984
rect 22573 840 22637 904
rect 22573 760 22637 824
rect 22573 680 22637 744
rect 22573 600 22637 664
rect 22573 520 22637 584
rect 22573 440 22637 504
rect 23179 1160 23243 1224
rect 23179 1080 23243 1144
rect 23179 1000 23243 1064
rect 23179 920 23243 984
rect 23179 840 23243 904
rect 23179 760 23243 824
rect 23179 680 23243 744
rect 23179 600 23243 664
rect 23179 520 23243 584
rect 23179 440 23243 504
rect 23785 1160 23849 1224
rect 23785 1080 23849 1144
rect 23785 1000 23849 1064
rect 23785 920 23849 984
rect 23785 840 23849 904
rect 23785 760 23849 824
rect 23785 680 23849 744
rect 23785 600 23849 664
rect 23785 520 23849 584
rect 23785 440 23849 504
rect 24391 1160 24455 1224
rect 24391 1080 24455 1144
rect 24391 1000 24455 1064
rect 24391 920 24455 984
rect 24391 840 24455 904
rect 24391 760 24455 824
rect 24391 680 24455 744
rect 24391 600 24455 664
rect 24391 520 24455 584
rect 24391 440 24455 504
rect 24997 1160 25061 1224
rect 24997 1080 25061 1144
rect 24997 1000 25061 1064
rect 24997 920 25061 984
rect 24997 840 25061 904
rect 24997 760 25061 824
rect 24997 680 25061 744
rect 24997 600 25061 664
rect 24997 520 25061 584
rect 24997 440 25061 504
rect 25603 1160 25667 1224
rect 25603 1080 25667 1144
rect 25603 1000 25667 1064
rect 25603 920 25667 984
rect 25603 840 25667 904
rect 25603 760 25667 824
rect 25603 680 25667 744
rect 25603 600 25667 664
rect 25603 520 25667 584
rect 25603 440 25667 504
rect 26209 1160 26273 1224
rect 26209 1080 26273 1144
rect 26209 1000 26273 1064
rect 26209 920 26273 984
rect 26209 840 26273 904
rect 26209 760 26273 824
rect 26209 680 26273 744
rect 26209 600 26273 664
rect 26209 520 26273 584
rect 26209 440 26273 504
rect 26815 1160 26879 1224
rect 26815 1080 26879 1144
rect 26815 1000 26879 1064
rect 26815 920 26879 984
rect 26815 840 26879 904
rect 26815 760 26879 824
rect 26815 680 26879 744
rect 26815 600 26879 664
rect 26815 520 26879 584
rect 26815 440 26879 504
rect 27421 1160 27485 1224
rect 27421 1080 27485 1144
rect 27421 1000 27485 1064
rect 27421 920 27485 984
rect 27421 840 27485 904
rect 27421 760 27485 824
rect 27421 680 27485 744
rect 27421 600 27485 664
rect 27421 520 27485 584
rect 27421 440 27485 504
rect 28027 1160 28091 1224
rect 28027 1080 28091 1144
rect 28027 1000 28091 1064
rect 28027 920 28091 984
rect 28027 840 28091 904
rect 28027 760 28091 824
rect 28027 680 28091 744
rect 28027 600 28091 664
rect 28027 520 28091 584
rect 28027 440 28091 504
rect 28633 1160 28697 1224
rect 28633 1080 28697 1144
rect 28633 1000 28697 1064
rect 28633 920 28697 984
rect 28633 840 28697 904
rect 28633 760 28697 824
rect 28633 680 28697 744
rect 28633 600 28697 664
rect 28633 520 28697 584
rect 28633 440 28697 504
rect 29239 1160 29303 1224
rect 29239 1080 29303 1144
rect 29239 1000 29303 1064
rect 29239 920 29303 984
rect 29239 840 29303 904
rect 29239 760 29303 824
rect 29239 680 29303 744
rect 29239 600 29303 664
rect 29239 520 29303 584
rect 29239 440 29303 504
rect 29845 1160 29909 1224
rect 29845 1080 29909 1144
rect 29845 1000 29909 1064
rect 29845 920 29909 984
rect 29845 840 29909 904
rect 29845 760 29909 824
rect 29845 680 29909 744
rect 29845 600 29909 664
rect 29845 520 29909 584
rect 29845 440 29909 504
rect 30451 1160 30515 1224
rect 30451 1080 30515 1144
rect 30451 1000 30515 1064
rect 30451 920 30515 984
rect 30451 840 30515 904
rect 30451 760 30515 824
rect 30451 680 30515 744
rect 30451 600 30515 664
rect 30451 520 30515 584
rect 30451 440 30515 504
rect 31057 1160 31121 1224
rect 31057 1080 31121 1144
rect 31057 1000 31121 1064
rect 31057 920 31121 984
rect 31057 840 31121 904
rect 31057 760 31121 824
rect 31057 680 31121 744
rect 31057 600 31121 664
rect 31057 520 31121 584
rect 31057 440 31121 504
rect 31663 1160 31727 1224
rect 31663 1080 31727 1144
rect 31663 1000 31727 1064
rect 31663 920 31727 984
rect 31663 840 31727 904
rect 31663 760 31727 824
rect 31663 680 31727 744
rect 31663 600 31727 664
rect 31663 520 31727 584
rect 31663 440 31727 504
rect 32269 1160 32333 1224
rect 32269 1080 32333 1144
rect 32269 1000 32333 1064
rect 32269 920 32333 984
rect 32269 840 32333 904
rect 32269 760 32333 824
rect 32269 680 32333 744
rect 32269 600 32333 664
rect 32269 520 32333 584
rect 32269 440 32333 504
rect 32875 1160 32939 1224
rect 32875 1080 32939 1144
rect 32875 1000 32939 1064
rect 32875 920 32939 984
rect 32875 840 32939 904
rect 32875 760 32939 824
rect 32875 680 32939 744
rect 32875 600 32939 664
rect 32875 520 32939 584
rect 32875 440 32939 504
rect 33481 1160 33545 1224
rect 33481 1080 33545 1144
rect 33481 1000 33545 1064
rect 33481 920 33545 984
rect 33481 840 33545 904
rect 33481 760 33545 824
rect 33481 680 33545 744
rect 33481 600 33545 664
rect 33481 520 33545 584
rect 33481 440 33545 504
rect 34087 1160 34151 1224
rect 34087 1080 34151 1144
rect 34087 1000 34151 1064
rect 34087 920 34151 984
rect 34087 840 34151 904
rect 34087 760 34151 824
rect 34087 680 34151 744
rect 34087 600 34151 664
rect 34087 520 34151 584
rect 34087 440 34151 504
rect 34693 1160 34757 1224
rect 34693 1080 34757 1144
rect 34693 1000 34757 1064
rect 34693 920 34757 984
rect 34693 840 34757 904
rect 34693 760 34757 824
rect 34693 680 34757 744
rect 34693 600 34757 664
rect 34693 520 34757 584
rect 34693 440 34757 504
rect 35299 1160 35363 1224
rect 35299 1080 35363 1144
rect 35299 1000 35363 1064
rect 35299 920 35363 984
rect 35299 840 35363 904
rect 35299 760 35363 824
rect 35299 680 35363 744
rect 35299 600 35363 664
rect 35299 520 35363 584
rect 35299 440 35363 504
rect 35905 1160 35969 1224
rect 35905 1080 35969 1144
rect 35905 1000 35969 1064
rect 35905 920 35969 984
rect 35905 840 35969 904
rect 35905 760 35969 824
rect 35905 680 35969 744
rect 35905 600 35969 664
rect 35905 520 35969 584
rect 35905 440 35969 504
rect 36511 1160 36575 1224
rect 36511 1080 36575 1144
rect 36511 1000 36575 1064
rect 36511 920 36575 984
rect 36511 840 36575 904
rect 36511 760 36575 824
rect 36511 680 36575 744
rect 36511 600 36575 664
rect 36511 520 36575 584
rect 36511 440 36575 504
rect 37117 1160 37181 1224
rect 37117 1080 37181 1144
rect 37117 1000 37181 1064
rect 37117 920 37181 984
rect 37117 840 37181 904
rect 37117 760 37181 824
rect 37117 680 37181 744
rect 37117 600 37181 664
rect 37117 520 37181 584
rect 37117 440 37181 504
rect 37723 1160 37787 1224
rect 37723 1080 37787 1144
rect 37723 1000 37787 1064
rect 37723 920 37787 984
rect 37723 840 37787 904
rect 37723 760 37787 824
rect 37723 680 37787 744
rect 37723 600 37787 664
rect 37723 520 37787 584
rect 37723 440 37787 504
rect 38329 1160 38393 1224
rect 38329 1080 38393 1144
rect 38329 1000 38393 1064
rect 38329 920 38393 984
rect 38329 840 38393 904
rect 38329 760 38393 824
rect 38329 680 38393 744
rect 38329 600 38393 664
rect 38329 520 38393 584
rect 38329 440 38393 504
rect 38935 1160 38999 1224
rect 38935 1080 38999 1144
rect 38935 1000 38999 1064
rect 38935 920 38999 984
rect 38935 840 38999 904
rect 38935 760 38999 824
rect 38935 680 38999 744
rect 38935 600 38999 664
rect 38935 520 38999 584
rect 38935 440 38999 504
rect 39541 1160 39605 1224
rect 39541 1080 39605 1144
rect 39541 1000 39605 1064
rect 39541 920 39605 984
rect 39541 840 39605 904
rect 39541 760 39605 824
rect 39541 680 39605 744
rect 39541 600 39605 664
rect 39541 520 39605 584
rect 39541 440 39605 504
rect -355 220 -291 284
rect -275 220 -211 284
rect -195 220 -131 284
rect -115 220 -51 284
rect -35 220 29 284
rect 45 220 109 284
rect 459 220 523 284
rect 539 220 603 284
rect 619 220 683 284
rect 699 220 763 284
rect 779 220 843 284
rect 859 220 923 284
rect 1371 220 1435 284
rect 1451 220 1515 284
rect 1531 220 1595 284
rect 1611 220 1675 284
rect 1691 220 1755 284
rect 1771 220 1835 284
rect 1977 220 2041 284
rect 2057 220 2121 284
rect 2137 220 2201 284
rect 2217 220 2281 284
rect 2297 220 2361 284
rect 2377 220 2441 284
rect 2905 220 2969 284
rect 2985 220 3049 284
rect 3065 220 3129 284
rect 3145 220 3209 284
rect 3225 220 3289 284
rect 3305 220 3369 284
rect 3511 220 3575 284
rect 3591 220 3655 284
rect 3671 220 3735 284
rect 3751 220 3815 284
rect 3831 220 3895 284
rect 3911 220 3975 284
rect 4117 220 4181 284
rect 4197 220 4261 284
rect 4277 220 4341 284
rect 4357 220 4421 284
rect 4437 220 4501 284
rect 4517 220 4581 284
rect 4723 220 4787 284
rect 4803 220 4867 284
rect 4883 220 4947 284
rect 4963 220 5027 284
rect 5043 220 5107 284
rect 5123 220 5187 284
rect 5456 220 5520 284
rect 5536 220 5600 284
rect 5616 220 5680 284
rect 5696 220 5760 284
rect 5776 220 5840 284
rect 5856 220 5920 284
rect 6062 220 6126 284
rect 6142 220 6206 284
rect 6222 220 6286 284
rect 6302 220 6366 284
rect 6382 220 6446 284
rect 6462 220 6526 284
rect 6668 220 6732 284
rect 6748 220 6812 284
rect 6828 220 6892 284
rect 6908 220 6972 284
rect 6988 220 7052 284
rect 7068 220 7132 284
rect 7274 220 7338 284
rect 7354 220 7418 284
rect 7434 220 7498 284
rect 7514 220 7578 284
rect 7594 220 7658 284
rect 7674 220 7738 284
rect 7880 220 7944 284
rect 7960 220 8024 284
rect 8040 220 8104 284
rect 8120 220 8184 284
rect 8200 220 8264 284
rect 8280 220 8344 284
rect 8486 220 8550 284
rect 8566 220 8630 284
rect 8646 220 8710 284
rect 8726 220 8790 284
rect 8806 220 8870 284
rect 8886 220 8950 284
rect 9092 220 9156 284
rect 9172 220 9236 284
rect 9252 220 9316 284
rect 9332 220 9396 284
rect 9412 220 9476 284
rect 9492 220 9556 284
rect 9698 220 9762 284
rect 9778 220 9842 284
rect 9858 220 9922 284
rect 9938 220 10002 284
rect 10018 220 10082 284
rect 10098 220 10162 284
rect 10430 220 10494 284
rect 10510 220 10574 284
rect 10590 220 10654 284
rect 10670 220 10734 284
rect 10750 220 10814 284
rect 10830 220 10894 284
rect 11036 220 11100 284
rect 11116 220 11180 284
rect 11196 220 11260 284
rect 11276 220 11340 284
rect 11356 220 11420 284
rect 11436 220 11500 284
rect 11642 220 11706 284
rect 11722 220 11786 284
rect 11802 220 11866 284
rect 11882 220 11946 284
rect 11962 220 12026 284
rect 12042 220 12106 284
rect 12248 220 12312 284
rect 12328 220 12392 284
rect 12408 220 12472 284
rect 12488 220 12552 284
rect 12568 220 12632 284
rect 12648 220 12712 284
rect 12854 220 12918 284
rect 12934 220 12998 284
rect 13014 220 13078 284
rect 13094 220 13158 284
rect 13174 220 13238 284
rect 13254 220 13318 284
rect 13460 220 13524 284
rect 13540 220 13604 284
rect 13620 220 13684 284
rect 13700 220 13764 284
rect 13780 220 13844 284
rect 13860 220 13924 284
rect 14066 220 14130 284
rect 14146 220 14210 284
rect 14226 220 14290 284
rect 14306 220 14370 284
rect 14386 220 14450 284
rect 14466 220 14530 284
rect 14672 220 14736 284
rect 14752 220 14816 284
rect 14832 220 14896 284
rect 14912 220 14976 284
rect 14992 220 15056 284
rect 15072 220 15136 284
rect 15278 220 15342 284
rect 15358 220 15422 284
rect 15438 220 15502 284
rect 15518 220 15582 284
rect 15598 220 15662 284
rect 15678 220 15742 284
rect 15884 220 15948 284
rect 15964 220 16028 284
rect 16044 220 16108 284
rect 16124 220 16188 284
rect 16204 220 16268 284
rect 16284 220 16348 284
rect 16490 220 16554 284
rect 16570 220 16634 284
rect 16650 220 16714 284
rect 16730 220 16794 284
rect 16810 220 16874 284
rect 16890 220 16954 284
rect 17096 220 17160 284
rect 17176 220 17240 284
rect 17256 220 17320 284
rect 17336 220 17400 284
rect 17416 220 17480 284
rect 17496 220 17560 284
rect 17702 220 17766 284
rect 17782 220 17846 284
rect 17862 220 17926 284
rect 17942 220 18006 284
rect 18022 220 18086 284
rect 18102 220 18166 284
rect 18308 220 18372 284
rect 18388 220 18452 284
rect 18468 220 18532 284
rect 18548 220 18612 284
rect 18628 220 18692 284
rect 18708 220 18772 284
rect 18914 220 18978 284
rect 18994 220 19058 284
rect 19074 220 19138 284
rect 19154 220 19218 284
rect 19234 220 19298 284
rect 19314 220 19378 284
rect 19520 220 19584 284
rect 19600 220 19664 284
rect 19680 220 19744 284
rect 19760 220 19824 284
rect 19840 220 19904 284
rect 19920 220 19984 284
rect 20252 220 20316 284
rect 20332 220 20396 284
rect 20412 220 20476 284
rect 20492 220 20556 284
rect 20572 220 20636 284
rect 20652 220 20716 284
rect 20858 220 20922 284
rect 20938 220 21002 284
rect 21018 220 21082 284
rect 21098 220 21162 284
rect 21178 220 21242 284
rect 21258 220 21322 284
rect 21464 220 21528 284
rect 21544 220 21608 284
rect 21624 220 21688 284
rect 21704 220 21768 284
rect 21784 220 21848 284
rect 21864 220 21928 284
rect 22070 220 22134 284
rect 22150 220 22214 284
rect 22230 220 22294 284
rect 22310 220 22374 284
rect 22390 220 22454 284
rect 22470 220 22534 284
rect 22676 220 22740 284
rect 22756 220 22820 284
rect 22836 220 22900 284
rect 22916 220 22980 284
rect 22996 220 23060 284
rect 23076 220 23140 284
rect 23282 220 23346 284
rect 23362 220 23426 284
rect 23442 220 23506 284
rect 23522 220 23586 284
rect 23602 220 23666 284
rect 23682 220 23746 284
rect 23888 220 23952 284
rect 23968 220 24032 284
rect 24048 220 24112 284
rect 24128 220 24192 284
rect 24208 220 24272 284
rect 24288 220 24352 284
rect 24494 220 24558 284
rect 24574 220 24638 284
rect 24654 220 24718 284
rect 24734 220 24798 284
rect 24814 220 24878 284
rect 24894 220 24958 284
rect 25100 220 25164 284
rect 25180 220 25244 284
rect 25260 220 25324 284
rect 25340 220 25404 284
rect 25420 220 25484 284
rect 25500 220 25564 284
rect 25706 220 25770 284
rect 25786 220 25850 284
rect 25866 220 25930 284
rect 25946 220 26010 284
rect 26026 220 26090 284
rect 26106 220 26170 284
rect 26312 220 26376 284
rect 26392 220 26456 284
rect 26472 220 26536 284
rect 26552 220 26616 284
rect 26632 220 26696 284
rect 26712 220 26776 284
rect 26918 220 26982 284
rect 26998 220 27062 284
rect 27078 220 27142 284
rect 27158 220 27222 284
rect 27238 220 27302 284
rect 27318 220 27382 284
rect 27524 220 27588 284
rect 27604 220 27668 284
rect 27684 220 27748 284
rect 27764 220 27828 284
rect 27844 220 27908 284
rect 27924 220 27988 284
rect 28130 220 28194 284
rect 28210 220 28274 284
rect 28290 220 28354 284
rect 28370 220 28434 284
rect 28450 220 28514 284
rect 28530 220 28594 284
rect 28736 220 28800 284
rect 28816 220 28880 284
rect 28896 220 28960 284
rect 28976 220 29040 284
rect 29056 220 29120 284
rect 29136 220 29200 284
rect 29342 220 29406 284
rect 29422 220 29486 284
rect 29502 220 29566 284
rect 29582 220 29646 284
rect 29662 220 29726 284
rect 29742 220 29806 284
rect 29948 220 30012 284
rect 30028 220 30092 284
rect 30108 220 30172 284
rect 30188 220 30252 284
rect 30268 220 30332 284
rect 30348 220 30412 284
rect 30554 220 30618 284
rect 30634 220 30698 284
rect 30714 220 30778 284
rect 30794 220 30858 284
rect 30874 220 30938 284
rect 30954 220 31018 284
rect 31160 220 31224 284
rect 31240 220 31304 284
rect 31320 220 31384 284
rect 31400 220 31464 284
rect 31480 220 31544 284
rect 31560 220 31624 284
rect 31766 220 31830 284
rect 31846 220 31910 284
rect 31926 220 31990 284
rect 32006 220 32070 284
rect 32086 220 32150 284
rect 32166 220 32230 284
rect 32372 220 32436 284
rect 32452 220 32516 284
rect 32532 220 32596 284
rect 32612 220 32676 284
rect 32692 220 32756 284
rect 32772 220 32836 284
rect 32978 220 33042 284
rect 33058 220 33122 284
rect 33138 220 33202 284
rect 33218 220 33282 284
rect 33298 220 33362 284
rect 33378 220 33442 284
rect 33584 220 33648 284
rect 33664 220 33728 284
rect 33744 220 33808 284
rect 33824 220 33888 284
rect 33904 220 33968 284
rect 33984 220 34048 284
rect 34190 220 34254 284
rect 34270 220 34334 284
rect 34350 220 34414 284
rect 34430 220 34494 284
rect 34510 220 34574 284
rect 34590 220 34654 284
rect 34796 220 34860 284
rect 34876 220 34940 284
rect 34956 220 35020 284
rect 35036 220 35100 284
rect 35116 220 35180 284
rect 35196 220 35260 284
rect 35402 220 35466 284
rect 35482 220 35546 284
rect 35562 220 35626 284
rect 35642 220 35706 284
rect 35722 220 35786 284
rect 35802 220 35866 284
rect 36008 220 36072 284
rect 36088 220 36152 284
rect 36168 220 36232 284
rect 36248 220 36312 284
rect 36328 220 36392 284
rect 36408 220 36472 284
rect 36614 220 36678 284
rect 36694 220 36758 284
rect 36774 220 36838 284
rect 36854 220 36918 284
rect 36934 220 36998 284
rect 37014 220 37078 284
rect 37220 220 37284 284
rect 37300 220 37364 284
rect 37380 220 37444 284
rect 37460 220 37524 284
rect 37540 220 37604 284
rect 37620 220 37684 284
rect 37826 220 37890 284
rect 37906 220 37970 284
rect 37986 220 38050 284
rect 38066 220 38130 284
rect 38146 220 38210 284
rect 38226 220 38290 284
rect 38432 220 38496 284
rect 38512 220 38576 284
rect 38592 220 38656 284
rect 38672 220 38736 284
rect 38752 220 38816 284
rect 38832 220 38896 284
rect 39038 220 39102 284
rect 39118 220 39182 284
rect 39198 220 39262 284
rect 39278 220 39342 284
rect 39358 220 39422 284
rect 39438 220 39502 284
<< metal4 >>
rect 29171 6320 29404 6321
rect 28942 6055 29404 6320
rect 28942 5991 28951 6055
rect 29015 5991 29404 6055
rect 28942 5756 29404 5991
rect 29171 5755 29404 5756
rect 29745 6058 30233 6365
rect 29745 5994 29758 6058
rect 29822 5994 30233 6058
rect 29745 5731 30233 5994
rect 29133 5423 29572 5639
rect 29133 5359 29147 5423
rect 29211 5359 29572 5423
rect -459 5092 213 5094
rect -459 5028 -355 5092
rect -291 5028 -275 5092
rect -211 5028 -195 5092
rect -131 5028 -115 5092
rect -51 5028 -35 5092
rect 29 5028 45 5092
rect 109 5028 213 5092
rect -459 5026 213 5028
rect 524 5092 1027 5094
rect 524 5028 539 5092
rect 603 5028 619 5092
rect 683 5028 699 5092
rect 763 5028 779 5092
rect 843 5028 859 5092
rect 923 5028 1027 5092
rect 524 5026 1027 5028
rect 1267 5092 1717 5094
rect 1954 5092 2545 5094
rect 1267 5028 1371 5092
rect 1435 5028 1451 5092
rect 1515 5028 1531 5092
rect 1595 5028 1611 5092
rect 1675 5028 1691 5092
rect 1954 5028 1977 5092
rect 2041 5028 2057 5092
rect 2121 5028 2137 5092
rect 2201 5028 2217 5092
rect 2281 5028 2297 5092
rect 2361 5028 2377 5092
rect 2441 5028 2545 5092
rect 1267 5026 1717 5028
rect 1954 5026 2545 5028
rect 2801 5092 3301 5094
rect 3538 5092 5291 5094
rect 2801 5028 2905 5092
rect 2969 5028 2985 5092
rect 3049 5028 3065 5092
rect 3129 5028 3145 5092
rect 3209 5028 3225 5092
rect 3289 5028 3301 5092
rect 3575 5028 3591 5092
rect 3655 5028 3671 5092
rect 3735 5028 3751 5092
rect 3815 5028 3831 5092
rect 3895 5028 3911 5092
rect 3975 5028 4117 5092
rect 4181 5028 4197 5092
rect 4261 5028 4277 5092
rect 4341 5028 4357 5092
rect 4421 5028 4437 5092
rect 4501 5028 4517 5092
rect 4581 5028 4723 5092
rect 4787 5028 4803 5092
rect 4867 5028 4883 5092
rect 4947 5028 4963 5092
rect 5027 5028 5043 5092
rect 5107 5028 5123 5092
rect 5187 5028 5291 5092
rect 2801 5026 3301 5028
rect 3538 5026 5291 5028
rect 5352 5026 5394 5094
rect 5631 5092 10266 5094
rect 5680 5028 5696 5092
rect 5760 5028 5776 5092
rect 5840 5028 5856 5092
rect 5920 5028 6062 5092
rect 6126 5028 6142 5092
rect 6206 5028 6222 5092
rect 6286 5028 6302 5092
rect 6366 5028 6382 5092
rect 6446 5028 6462 5092
rect 6526 5028 6668 5092
rect 6732 5028 6748 5092
rect 6812 5028 6828 5092
rect 6892 5028 6908 5092
rect 6972 5028 6988 5092
rect 7052 5028 7068 5092
rect 7132 5028 7274 5092
rect 7338 5028 7354 5092
rect 7418 5028 7434 5092
rect 7498 5028 7514 5092
rect 7578 5028 7594 5092
rect 7658 5028 7674 5092
rect 7738 5028 7880 5092
rect 7944 5028 7960 5092
rect 8024 5028 8040 5092
rect 8104 5028 8120 5092
rect 8184 5028 8200 5092
rect 8264 5028 8280 5092
rect 8344 5028 8486 5092
rect 8550 5028 8566 5092
rect 8630 5028 8646 5092
rect 8710 5028 8726 5092
rect 8790 5028 8806 5092
rect 8870 5028 8886 5092
rect 8950 5028 9092 5092
rect 9156 5028 9172 5092
rect 9236 5028 9252 5092
rect 9316 5028 9332 5092
rect 9396 5028 9412 5092
rect 9476 5028 9492 5092
rect 9556 5028 9698 5092
rect 9762 5028 9778 5092
rect 9842 5028 9858 5092
rect 9922 5028 9938 5092
rect 10002 5028 10018 5092
rect 10082 5028 10098 5092
rect 10162 5028 10266 5092
rect 5631 5026 10266 5028
rect 10326 5026 10368 5094
rect 29133 5154 29572 5359
rect 10605 5092 20088 5094
rect 10654 5028 10670 5092
rect 10734 5028 10750 5092
rect 10814 5028 10830 5092
rect 10894 5028 11036 5092
rect 11100 5028 11116 5092
rect 11180 5028 11196 5092
rect 11260 5028 11276 5092
rect 11340 5028 11356 5092
rect 11420 5028 11436 5092
rect 11500 5028 11642 5092
rect 11706 5028 11722 5092
rect 11786 5028 11802 5092
rect 11866 5028 11882 5092
rect 11946 5028 11962 5092
rect 12026 5028 12042 5092
rect 12106 5028 12248 5092
rect 12312 5028 12328 5092
rect 12392 5028 12408 5092
rect 12472 5028 12488 5092
rect 12552 5028 12568 5092
rect 12632 5028 12648 5092
rect 12712 5028 12854 5092
rect 12918 5028 12934 5092
rect 12998 5028 13014 5092
rect 13078 5028 13094 5092
rect 13158 5028 13174 5092
rect 13238 5028 13254 5092
rect 13318 5028 13460 5092
rect 13524 5028 13540 5092
rect 13604 5028 13620 5092
rect 13684 5028 13700 5092
rect 13764 5028 13780 5092
rect 13844 5028 13860 5092
rect 13924 5028 14066 5092
rect 14130 5028 14146 5092
rect 14210 5028 14226 5092
rect 14290 5028 14306 5092
rect 14370 5028 14386 5092
rect 14450 5028 14466 5092
rect 14530 5028 14672 5092
rect 14736 5028 14752 5092
rect 14816 5028 14832 5092
rect 14896 5028 14912 5092
rect 14976 5028 14992 5092
rect 15056 5028 15072 5092
rect 15136 5028 15278 5092
rect 15342 5028 15358 5092
rect 15422 5028 15438 5092
rect 15502 5028 15518 5092
rect 15582 5028 15598 5092
rect 15662 5028 15678 5092
rect 15742 5028 15884 5092
rect 15948 5028 15964 5092
rect 16028 5028 16044 5092
rect 16108 5028 16124 5092
rect 16188 5028 16204 5092
rect 16268 5028 16284 5092
rect 16348 5028 16490 5092
rect 16554 5028 16570 5092
rect 16634 5028 16650 5092
rect 16714 5028 16730 5092
rect 16794 5028 16810 5092
rect 16874 5028 16890 5092
rect 16954 5028 17096 5092
rect 17160 5028 17176 5092
rect 17240 5028 17256 5092
rect 17320 5028 17336 5092
rect 17400 5028 17416 5092
rect 17480 5028 17496 5092
rect 17560 5028 17702 5092
rect 17766 5028 17782 5092
rect 17846 5028 17862 5092
rect 17926 5028 17942 5092
rect 18006 5028 18022 5092
rect 18086 5028 18102 5092
rect 18166 5028 18308 5092
rect 18372 5028 18388 5092
rect 18452 5028 18468 5092
rect 18532 5028 18548 5092
rect 18612 5028 18628 5092
rect 18692 5028 18708 5092
rect 18772 5028 18914 5092
rect 18978 5028 18994 5092
rect 19058 5028 19074 5092
rect 19138 5028 19154 5092
rect 19218 5028 19234 5092
rect 19298 5028 19314 5092
rect 19378 5028 19520 5092
rect 19584 5028 19600 5092
rect 19664 5028 19680 5092
rect 19744 5028 19760 5092
rect 19824 5028 19840 5092
rect 19904 5028 19920 5092
rect 19984 5028 20088 5092
rect 10605 5026 20088 5028
rect 20148 5092 39298 5094
rect 20148 5028 20252 5092
rect 20316 5028 20332 5092
rect 20396 5028 20412 5092
rect 20476 5028 20492 5092
rect 20556 5028 20572 5092
rect 20636 5028 20652 5092
rect 20716 5028 20858 5092
rect 20922 5028 20938 5092
rect 21002 5028 21018 5092
rect 21082 5028 21098 5092
rect 21162 5028 21178 5092
rect 21242 5028 21258 5092
rect 21322 5028 21464 5092
rect 21528 5028 21544 5092
rect 21608 5028 21624 5092
rect 21688 5028 21704 5092
rect 21768 5028 21784 5092
rect 21848 5028 21864 5092
rect 21928 5028 22070 5092
rect 22134 5028 22150 5092
rect 22214 5028 22230 5092
rect 22294 5028 22310 5092
rect 22374 5028 22390 5092
rect 22454 5028 22470 5092
rect 22534 5028 22676 5092
rect 22740 5028 22756 5092
rect 22820 5028 22836 5092
rect 22900 5028 22916 5092
rect 22980 5028 22996 5092
rect 23060 5028 23076 5092
rect 23140 5028 23282 5092
rect 23346 5028 23362 5092
rect 23426 5028 23442 5092
rect 23506 5028 23522 5092
rect 23586 5028 23602 5092
rect 23666 5028 23682 5092
rect 23746 5028 23888 5092
rect 23952 5028 23968 5092
rect 24032 5028 24048 5092
rect 24112 5028 24128 5092
rect 24192 5028 24208 5092
rect 24272 5028 24288 5092
rect 24352 5028 24494 5092
rect 24558 5028 24574 5092
rect 24638 5028 24654 5092
rect 24718 5028 24734 5092
rect 24798 5028 24814 5092
rect 24878 5028 24894 5092
rect 24958 5028 25100 5092
rect 25164 5028 25180 5092
rect 25244 5028 25260 5092
rect 25324 5028 25340 5092
rect 25404 5028 25420 5092
rect 25484 5028 25500 5092
rect 25564 5028 25706 5092
rect 25770 5028 25786 5092
rect 25850 5028 25866 5092
rect 25930 5028 25946 5092
rect 26010 5028 26026 5092
rect 26090 5028 26106 5092
rect 26170 5028 26312 5092
rect 26376 5028 26392 5092
rect 26456 5028 26472 5092
rect 26536 5028 26552 5092
rect 26616 5028 26632 5092
rect 26696 5028 26712 5092
rect 26776 5028 26918 5092
rect 26982 5028 26998 5092
rect 27062 5028 27078 5092
rect 27142 5028 27158 5092
rect 27222 5028 27238 5092
rect 27302 5028 27318 5092
rect 27382 5028 27524 5092
rect 27588 5028 27604 5092
rect 27668 5028 27684 5092
rect 27748 5028 27764 5092
rect 27828 5028 27844 5092
rect 27908 5028 27924 5092
rect 27988 5028 28130 5092
rect 28194 5028 28210 5092
rect 28274 5028 28290 5092
rect 28354 5028 28370 5092
rect 28434 5028 28450 5092
rect 28514 5028 28530 5092
rect 28594 5028 28736 5092
rect 28800 5028 28816 5092
rect 28880 5028 28896 5092
rect 28960 5028 28976 5092
rect 29040 5028 29056 5092
rect 29120 5028 29136 5092
rect 29200 5028 29342 5092
rect 29406 5028 29422 5092
rect 29486 5028 29502 5092
rect 29566 5028 29582 5092
rect 29646 5028 29662 5092
rect 29726 5028 29742 5092
rect 29806 5028 29948 5092
rect 30012 5028 30028 5092
rect 30092 5028 30108 5092
rect 30172 5028 30188 5092
rect 30252 5028 30268 5092
rect 30332 5028 30348 5092
rect 30412 5028 30554 5092
rect 30618 5028 30634 5092
rect 30698 5028 30714 5092
rect 30778 5028 30794 5092
rect 30858 5028 30874 5092
rect 30938 5028 30954 5092
rect 31018 5028 31160 5092
rect 31224 5028 31240 5092
rect 31304 5028 31320 5092
rect 31384 5028 31400 5092
rect 31464 5028 31480 5092
rect 31544 5028 31560 5092
rect 31624 5028 31766 5092
rect 31830 5028 31846 5092
rect 31910 5028 31926 5092
rect 31990 5028 32006 5092
rect 32070 5028 32086 5092
rect 32150 5028 32166 5092
rect 32230 5028 32372 5092
rect 32436 5028 32452 5092
rect 32516 5028 32532 5092
rect 32596 5028 32612 5092
rect 32676 5028 32692 5092
rect 32756 5028 32772 5092
rect 32836 5028 32978 5092
rect 33042 5028 33058 5092
rect 33122 5028 33138 5092
rect 33202 5028 33218 5092
rect 33282 5028 33298 5092
rect 33362 5028 33378 5092
rect 33442 5028 33584 5092
rect 33648 5028 33664 5092
rect 33728 5028 33744 5092
rect 33808 5028 33824 5092
rect 33888 5028 33904 5092
rect 33968 5028 33984 5092
rect 34048 5028 34190 5092
rect 34254 5028 34270 5092
rect 34334 5028 34350 5092
rect 34414 5028 34430 5092
rect 34494 5028 34510 5092
rect 34574 5028 34590 5092
rect 34654 5028 34796 5092
rect 34860 5028 34876 5092
rect 34940 5028 34956 5092
rect 35020 5028 35036 5092
rect 35100 5028 35116 5092
rect 35180 5028 35196 5092
rect 35260 5028 35402 5092
rect 35466 5028 35482 5092
rect 35546 5028 35562 5092
rect 35626 5028 35642 5092
rect 35706 5028 35722 5092
rect 35786 5028 35802 5092
rect 35866 5028 36008 5092
rect 36072 5028 36088 5092
rect 36152 5028 36168 5092
rect 36232 5028 36248 5092
rect 36312 5028 36328 5092
rect 36392 5028 36408 5092
rect 36472 5028 36614 5092
rect 36678 5028 36694 5092
rect 36758 5028 36774 5092
rect 36838 5028 36854 5092
rect 36918 5028 36934 5092
rect 36998 5028 37014 5092
rect 37078 5028 37220 5092
rect 37284 5028 37300 5092
rect 37364 5028 37380 5092
rect 37444 5028 37460 5092
rect 37524 5028 37540 5092
rect 37604 5028 37620 5092
rect 37684 5028 37826 5092
rect 37890 5028 37906 5092
rect 37970 5028 37986 5092
rect 38050 5028 38066 5092
rect 38130 5028 38146 5092
rect 38210 5028 38226 5092
rect 38290 5028 38432 5092
rect 38496 5028 38512 5092
rect 38576 5028 38592 5092
rect 38656 5028 38672 5092
rect 38736 5028 38752 5092
rect 38816 5028 38832 5092
rect 38896 5028 39038 5092
rect 39102 5028 39118 5092
rect 39182 5028 39198 5092
rect 39262 5028 39278 5092
rect 20148 5026 39298 5028
rect 39534 5026 39606 5094
rect -459 4872 -393 5026
rect -459 4808 -458 4872
rect -394 4808 -393 4872
rect -459 4792 -393 4808
rect -459 4728 -458 4792
rect -394 4728 -393 4792
rect -459 4712 -393 4728
rect -459 4648 -458 4712
rect -394 4648 -393 4712
rect -459 4632 -393 4648
rect -459 4568 -458 4632
rect -394 4568 -393 4632
rect -459 4552 -393 4568
rect -459 4488 -458 4552
rect -394 4488 -393 4552
rect -459 4472 -393 4488
rect -459 4408 -458 4472
rect -394 4408 -393 4472
rect -459 4392 -393 4408
rect -459 4328 -458 4392
rect -394 4328 -393 4392
rect -459 4312 -393 4328
rect -459 4248 -458 4312
rect -394 4248 -393 4312
rect -459 4232 -393 4248
rect -459 4168 -458 4232
rect -394 4168 -393 4232
rect -459 4152 -393 4168
rect -459 4088 -458 4152
rect -394 4088 -393 4152
rect -459 3998 -393 4088
rect -333 3994 -273 5026
rect -213 3934 -153 4964
rect -93 3994 -33 5026
rect 27 3934 87 4964
rect 147 4872 213 5026
rect 147 4808 148 4872
rect 212 4808 213 4872
rect 147 4792 213 4808
rect 147 4728 148 4792
rect 212 4728 213 4792
rect 147 4712 213 4728
rect 147 4648 148 4712
rect 212 4648 213 4712
rect 147 4632 213 4648
rect 147 4568 148 4632
rect 212 4568 213 4632
rect 147 4552 213 4568
rect 147 4488 148 4552
rect 212 4488 213 4552
rect 147 4472 213 4488
rect 147 4408 148 4472
rect 212 4408 213 4472
rect 147 4392 213 4408
rect 147 4328 148 4392
rect 212 4328 213 4392
rect 147 4312 213 4328
rect 147 4248 148 4312
rect 212 4248 213 4312
rect 147 4232 213 4248
rect 147 4168 148 4232
rect 212 4168 213 4232
rect 147 4152 213 4168
rect 147 4088 148 4152
rect 212 4088 213 4152
rect 147 3998 213 4088
rect 355 4872 421 4962
rect 355 4808 356 4872
rect 420 4808 421 4872
rect 355 4792 421 4808
rect 355 4728 356 4792
rect 420 4728 421 4792
rect 355 4712 421 4728
rect 355 4648 356 4712
rect 420 4648 421 4712
rect 355 4632 421 4648
rect 355 4568 356 4632
rect 420 4568 421 4632
rect 355 4552 421 4568
rect 355 4488 356 4552
rect 420 4488 421 4552
rect 355 4472 421 4488
rect 355 4408 356 4472
rect 420 4408 421 4472
rect 355 4392 421 4408
rect 355 4328 356 4392
rect 420 4328 421 4392
rect 355 4312 421 4328
rect 355 4248 356 4312
rect 420 4248 421 4312
rect 355 4232 421 4248
rect 355 4168 356 4232
rect 420 4168 421 4232
rect 355 4152 421 4168
rect 355 4088 356 4152
rect 420 4088 421 4152
rect 150 3994 210 3998
rect 355 3934 421 4088
rect 481 3996 541 5026
rect 601 3934 661 4966
rect 721 3996 781 5026
rect 841 3934 901 4966
rect 961 4872 1027 4962
rect 961 4808 962 4872
rect 1026 4808 1027 4872
rect 961 4792 1027 4808
rect 961 4728 962 4792
rect 1026 4728 1027 4792
rect 961 4712 1027 4728
rect 961 4648 962 4712
rect 1026 4648 1027 4712
rect 961 4632 1027 4648
rect 961 4568 962 4632
rect 1026 4568 1027 4632
rect 961 4552 1027 4568
rect 961 4488 962 4552
rect 1026 4488 1027 4552
rect 961 4472 1027 4488
rect 961 4408 962 4472
rect 1026 4408 1027 4472
rect 961 4392 1027 4408
rect 961 4328 962 4392
rect 1026 4328 1027 4392
rect 961 4312 1027 4328
rect 961 4248 962 4312
rect 1026 4248 1027 4312
rect 961 4232 1027 4248
rect 961 4168 962 4232
rect 1026 4168 1027 4232
rect 961 4152 1027 4168
rect 961 4088 962 4152
rect 1026 4088 1027 4152
rect 961 3934 1027 4088
rect -459 3932 213 3934
rect -459 3868 -355 3932
rect -291 3868 -275 3932
rect -211 3868 -195 3932
rect -131 3868 -115 3932
rect -51 3868 -35 3932
rect 29 3868 45 3932
rect 109 3868 213 3932
rect -459 3866 213 3868
rect 355 3932 1027 3934
rect 355 3868 459 3932
rect 523 3868 539 3932
rect 603 3868 619 3932
rect 683 3868 699 3932
rect 763 3868 779 3932
rect 843 3868 859 3932
rect 923 3868 1027 3932
rect 355 3866 1027 3868
rect -459 3712 -393 3802
rect -459 3648 -458 3712
rect -394 3648 -393 3712
rect -459 3632 -393 3648
rect -459 3568 -458 3632
rect -394 3568 -393 3632
rect -459 3552 -393 3568
rect -459 3488 -458 3552
rect -394 3488 -393 3552
rect -459 3472 -393 3488
rect -459 3408 -458 3472
rect -394 3408 -393 3472
rect -459 3392 -393 3408
rect -459 3328 -458 3392
rect -394 3328 -393 3392
rect -459 3312 -393 3328
rect -459 3248 -458 3312
rect -394 3248 -393 3312
rect -459 3232 -393 3248
rect -459 3168 -458 3232
rect -394 3168 -393 3232
rect -459 3152 -393 3168
rect -459 3088 -458 3152
rect -394 3088 -393 3152
rect -459 3072 -393 3088
rect -459 3008 -458 3072
rect -394 3008 -393 3072
rect -459 2992 -393 3008
rect -459 2928 -458 2992
rect -394 2928 -393 2992
rect -459 2774 -393 2928
rect -333 2836 -273 3866
rect -213 2774 -153 3806
rect -93 2836 -33 3866
rect 27 2774 87 3806
rect 147 3712 213 3802
rect 147 3648 148 3712
rect 212 3648 213 3712
rect 147 3632 213 3648
rect 147 3568 148 3632
rect 212 3568 213 3632
rect 147 3552 213 3568
rect 147 3488 148 3552
rect 212 3488 213 3552
rect 147 3472 213 3488
rect 147 3408 148 3472
rect 212 3408 213 3472
rect 147 3392 213 3408
rect 147 3328 148 3392
rect 212 3328 213 3392
rect 147 3312 213 3328
rect 147 3248 148 3312
rect 212 3248 213 3312
rect 147 3232 213 3248
rect 147 3168 148 3232
rect 212 3168 213 3232
rect 147 3152 213 3168
rect 147 3088 148 3152
rect 212 3088 213 3152
rect 147 3072 213 3088
rect 147 3008 148 3072
rect 212 3008 213 3072
rect 147 2992 213 3008
rect 147 2928 148 2992
rect 212 2928 213 2992
rect 147 2774 213 2928
rect 355 3712 421 3866
rect 355 3648 356 3712
rect 420 3648 421 3712
rect 355 3632 421 3648
rect 355 3568 356 3632
rect 420 3568 421 3632
rect 355 3552 421 3568
rect 355 3488 356 3552
rect 420 3488 421 3552
rect 355 3472 421 3488
rect 355 3408 356 3472
rect 420 3408 421 3472
rect 355 3392 421 3408
rect 355 3328 356 3392
rect 420 3328 421 3392
rect 355 3312 421 3328
rect 355 3248 356 3312
rect 420 3248 421 3312
rect 355 3232 421 3248
rect 355 3168 356 3232
rect 420 3168 421 3232
rect 355 3152 421 3168
rect 355 3088 356 3152
rect 420 3088 421 3152
rect 355 3072 421 3088
rect 355 3008 356 3072
rect 420 3008 421 3072
rect 355 2992 421 3008
rect 355 2928 356 2992
rect 420 2928 421 2992
rect 355 2838 421 2928
rect 481 2834 541 3866
rect 601 2774 661 3804
rect 721 2834 781 3866
rect 841 2774 901 3804
rect 961 3712 1027 3866
rect 961 3648 962 3712
rect 1026 3648 1027 3712
rect 961 3632 1027 3648
rect 961 3568 962 3632
rect 1026 3568 1027 3632
rect 961 3552 1027 3568
rect 961 3488 962 3552
rect 1026 3488 1027 3552
rect 961 3472 1027 3488
rect 961 3408 962 3472
rect 1026 3408 1027 3472
rect 961 3392 1027 3408
rect 961 3328 962 3392
rect 1026 3328 1027 3392
rect 961 3312 1027 3328
rect 961 3248 962 3312
rect 1026 3248 1027 3312
rect 961 3232 1027 3248
rect 961 3168 962 3232
rect 1026 3168 1027 3232
rect 961 3152 1027 3168
rect 961 3088 962 3152
rect 1026 3088 1027 3152
rect 961 3072 1027 3088
rect 961 3008 962 3072
rect 1026 3008 1027 3072
rect 961 2992 1027 3008
rect 961 2928 962 2992
rect 1026 2928 1027 2992
rect 961 2838 1027 2928
rect 1267 4872 1333 4962
rect 1267 4808 1268 4872
rect 1332 4808 1333 4872
rect 1267 4792 1333 4808
rect 1267 4728 1268 4792
rect 1332 4728 1333 4792
rect 1267 4712 1333 4728
rect 1267 4648 1268 4712
rect 1332 4648 1333 4712
rect 1267 4632 1333 4648
rect 1267 4568 1268 4632
rect 1332 4568 1333 4632
rect 1267 4552 1333 4568
rect 1267 4488 1268 4552
rect 1332 4488 1333 4552
rect 1267 4472 1333 4488
rect 1267 4408 1268 4472
rect 1332 4408 1333 4472
rect 1267 4392 1333 4408
rect 1267 4328 1268 4392
rect 1332 4328 1333 4392
rect 1267 4312 1333 4328
rect 1267 4248 1268 4312
rect 1332 4248 1333 4312
rect 1267 4232 1333 4248
rect 1267 4168 1268 4232
rect 1332 4168 1333 4232
rect 1267 4152 1333 4168
rect 1267 4088 1268 4152
rect 1332 4088 1333 4152
rect 1267 3934 1333 4088
rect 1393 3996 1453 5026
rect 1513 3934 1573 4966
rect 1633 3996 1693 5026
rect 1753 3934 1813 4966
rect 1873 4872 1939 4962
rect 1873 4808 1874 4872
rect 1938 4808 1939 4872
rect 1873 4792 1939 4808
rect 1873 4728 1874 4792
rect 1938 4728 1939 4792
rect 1873 4712 1939 4728
rect 1873 4648 1874 4712
rect 1938 4648 1939 4712
rect 1873 4632 1939 4648
rect 1873 4568 1874 4632
rect 1938 4568 1939 4632
rect 1873 4552 1939 4568
rect 1873 4488 1874 4552
rect 1938 4488 1939 4552
rect 1873 4472 1939 4488
rect 1873 4408 1874 4472
rect 1938 4408 1939 4472
rect 1873 4392 1939 4408
rect 1873 4328 1874 4392
rect 1938 4328 1939 4392
rect 1873 4312 1939 4328
rect 1873 4248 1874 4312
rect 1938 4248 1939 4312
rect 1873 4232 1939 4248
rect 1873 4168 1874 4232
rect 1938 4168 1939 4232
rect 1873 4152 1939 4168
rect 1873 4088 1874 4152
rect 1938 4088 1939 4152
rect 1873 3934 1939 4088
rect 1999 3996 2059 5026
rect 2119 3934 2179 4966
rect 2239 3996 2299 5026
rect 2359 3934 2419 4966
rect 2479 4872 2545 4962
rect 2479 4808 2480 4872
rect 2544 4808 2545 4872
rect 2479 4792 2545 4808
rect 2479 4728 2480 4792
rect 2544 4728 2545 4792
rect 2479 4712 2545 4728
rect 2479 4648 2480 4712
rect 2544 4648 2545 4712
rect 2479 4632 2545 4648
rect 2479 4568 2480 4632
rect 2544 4568 2545 4632
rect 2479 4552 2545 4568
rect 2479 4488 2480 4552
rect 2544 4488 2545 4552
rect 2479 4472 2545 4488
rect 2479 4408 2480 4472
rect 2544 4408 2545 4472
rect 2479 4392 2545 4408
rect 2479 4328 2480 4392
rect 2544 4328 2545 4392
rect 2479 4312 2545 4328
rect 2479 4248 2480 4312
rect 2544 4248 2545 4312
rect 2479 4232 2545 4248
rect 2479 4168 2480 4232
rect 2544 4168 2545 4232
rect 2479 4152 2545 4168
rect 2479 4088 2480 4152
rect 2544 4088 2545 4152
rect 2479 3934 2545 4088
rect 1267 3932 2545 3934
rect 1267 3868 1371 3932
rect 1435 3868 1451 3932
rect 1515 3868 1531 3932
rect 1595 3868 1611 3932
rect 1675 3868 1691 3932
rect 1755 3868 1771 3932
rect 1835 3868 1977 3932
rect 2041 3868 2057 3932
rect 2121 3868 2137 3932
rect 2201 3868 2217 3932
rect 2281 3868 2297 3932
rect 2361 3868 2377 3932
rect 2441 3868 2545 3932
rect 1267 3866 2545 3868
rect 1267 3712 1333 3866
rect 1267 3648 1268 3712
rect 1332 3648 1333 3712
rect 1267 3632 1333 3648
rect 1267 3568 1268 3632
rect 1332 3568 1333 3632
rect 1267 3552 1333 3568
rect 1267 3488 1268 3552
rect 1332 3488 1333 3552
rect 1267 3472 1333 3488
rect 1267 3408 1268 3472
rect 1332 3408 1333 3472
rect 1267 3392 1333 3408
rect 1267 3328 1268 3392
rect 1332 3328 1333 3392
rect 1267 3312 1333 3328
rect 1267 3248 1268 3312
rect 1332 3248 1333 3312
rect 1267 3232 1333 3248
rect 1267 3168 1268 3232
rect 1332 3168 1333 3232
rect 1267 3152 1333 3168
rect 1267 3088 1268 3152
rect 1332 3088 1333 3152
rect 1267 3072 1333 3088
rect 1267 3008 1268 3072
rect 1332 3008 1333 3072
rect 1267 2992 1333 3008
rect 1267 2928 1268 2992
rect 1332 2928 1333 2992
rect 1267 2838 1333 2928
rect 1393 2834 1453 3866
rect 1513 2774 1573 3804
rect 1633 2834 1693 3866
rect 1753 2774 1813 3804
rect 1873 3712 1939 3866
rect 1873 3648 1874 3712
rect 1938 3648 1939 3712
rect 1873 3632 1939 3648
rect 1873 3568 1874 3632
rect 1938 3568 1939 3632
rect 1873 3552 1939 3568
rect 1873 3488 1874 3552
rect 1938 3488 1939 3552
rect 1873 3472 1939 3488
rect 1873 3408 1874 3472
rect 1938 3408 1939 3472
rect 1873 3392 1939 3408
rect 1873 3328 1874 3392
rect 1938 3328 1939 3392
rect 1873 3312 1939 3328
rect 1873 3248 1874 3312
rect 1938 3248 1939 3312
rect 1873 3232 1939 3248
rect 1873 3168 1874 3232
rect 1938 3168 1939 3232
rect 1873 3152 1939 3168
rect 1873 3088 1874 3152
rect 1938 3088 1939 3152
rect 1873 3072 1939 3088
rect 1873 3008 1874 3072
rect 1938 3008 1939 3072
rect 1873 2992 1939 3008
rect 1873 2928 1874 2992
rect 1938 2928 1939 2992
rect 1873 2838 1939 2928
rect 1999 2834 2059 3866
rect 2119 2774 2179 3804
rect 2239 2834 2299 3866
rect 2359 2774 2419 3804
rect 2479 3712 2545 3866
rect 2479 3648 2480 3712
rect 2544 3648 2545 3712
rect 2479 3632 2545 3648
rect 2479 3568 2480 3632
rect 2544 3568 2545 3632
rect 2479 3552 2545 3568
rect 2479 3488 2480 3552
rect 2544 3488 2545 3552
rect 2479 3472 2545 3488
rect 2479 3408 2480 3472
rect 2544 3408 2545 3472
rect 2479 3392 2545 3408
rect 2479 3328 2480 3392
rect 2544 3328 2545 3392
rect 2479 3312 2545 3328
rect 2479 3248 2480 3312
rect 2544 3248 2545 3312
rect 2479 3232 2545 3248
rect 2479 3168 2480 3232
rect 2544 3168 2545 3232
rect 2479 3152 2545 3168
rect 2479 3088 2480 3152
rect 2544 3088 2545 3152
rect 2479 3072 2545 3088
rect 2479 3008 2480 3072
rect 2544 3008 2545 3072
rect 2479 2992 2545 3008
rect 2479 2928 2480 2992
rect 2544 2928 2545 2992
rect 2479 2838 2545 2928
rect 2801 4872 2867 4962
rect 2801 4808 2802 4872
rect 2866 4808 2867 4872
rect 2801 4792 2867 4808
rect 2801 4728 2802 4792
rect 2866 4728 2867 4792
rect 2801 4712 2867 4728
rect 2801 4648 2802 4712
rect 2866 4648 2867 4712
rect 2801 4632 2867 4648
rect 2801 4568 2802 4632
rect 2866 4568 2867 4632
rect 2801 4552 2867 4568
rect 2801 4488 2802 4552
rect 2866 4488 2867 4552
rect 2801 4472 2867 4488
rect 2801 4408 2802 4472
rect 2866 4408 2867 4472
rect 2801 4392 2867 4408
rect 2801 4328 2802 4392
rect 2866 4328 2867 4392
rect 2801 4312 2867 4328
rect 2801 4248 2802 4312
rect 2866 4248 2867 4312
rect 2801 4232 2867 4248
rect 2801 4168 2802 4232
rect 2866 4168 2867 4232
rect 2801 4152 2867 4168
rect 2801 4088 2802 4152
rect 2866 4088 2867 4152
rect 2801 3934 2867 4088
rect 2927 3996 2987 5026
rect 3047 3934 3107 4966
rect 3167 3996 3227 5026
rect 3287 3934 3347 4966
rect 3407 4872 3473 4962
rect 3407 4808 3408 4872
rect 3472 4808 3473 4872
rect 3407 4792 3473 4808
rect 3407 4728 3408 4792
rect 3472 4728 3473 4792
rect 3407 4712 3473 4728
rect 3407 4648 3408 4712
rect 3472 4648 3473 4712
rect 3407 4632 3473 4648
rect 3407 4568 3408 4632
rect 3472 4568 3473 4632
rect 3407 4552 3473 4568
rect 3407 4488 3408 4552
rect 3472 4488 3473 4552
rect 3407 4472 3473 4488
rect 3407 4408 3408 4472
rect 3472 4408 3473 4472
rect 3407 4392 3473 4408
rect 3407 4328 3408 4392
rect 3472 4328 3473 4392
rect 3407 4312 3473 4328
rect 3407 4248 3408 4312
rect 3472 4248 3473 4312
rect 3407 4232 3473 4248
rect 3407 4168 3408 4232
rect 3472 4168 3473 4232
rect 3407 4152 3473 4168
rect 3407 4088 3408 4152
rect 3472 4088 3473 4152
rect 3407 3934 3473 4088
rect 3533 3996 3593 5026
rect 3653 3934 3713 4966
rect 3773 3996 3833 5026
rect 3893 3934 3953 4966
rect 4013 4872 4079 4962
rect 4013 4808 4014 4872
rect 4078 4808 4079 4872
rect 4013 4792 4079 4808
rect 4013 4728 4014 4792
rect 4078 4728 4079 4792
rect 4013 4712 4079 4728
rect 4013 4648 4014 4712
rect 4078 4648 4079 4712
rect 4013 4632 4079 4648
rect 4013 4568 4014 4632
rect 4078 4568 4079 4632
rect 4013 4552 4079 4568
rect 4013 4488 4014 4552
rect 4078 4488 4079 4552
rect 4013 4472 4079 4488
rect 4013 4408 4014 4472
rect 4078 4408 4079 4472
rect 4013 4392 4079 4408
rect 4013 4328 4014 4392
rect 4078 4328 4079 4392
rect 4013 4312 4079 4328
rect 4013 4248 4014 4312
rect 4078 4248 4079 4312
rect 4013 4232 4079 4248
rect 4013 4168 4014 4232
rect 4078 4168 4079 4232
rect 4013 4152 4079 4168
rect 4013 4088 4014 4152
rect 4078 4088 4079 4152
rect 4013 3934 4079 4088
rect 4139 3996 4199 5026
rect 4259 3934 4319 4966
rect 4379 3996 4439 5026
rect 4499 3934 4559 4966
rect 4619 4872 4685 4962
rect 4619 4808 4620 4872
rect 4684 4808 4685 4872
rect 4619 4792 4685 4808
rect 4619 4728 4620 4792
rect 4684 4728 4685 4792
rect 4619 4712 4685 4728
rect 4619 4648 4620 4712
rect 4684 4648 4685 4712
rect 4619 4632 4685 4648
rect 4619 4568 4620 4632
rect 4684 4568 4685 4632
rect 4619 4552 4685 4568
rect 4619 4488 4620 4552
rect 4684 4488 4685 4552
rect 4619 4472 4685 4488
rect 4619 4408 4620 4472
rect 4684 4408 4685 4472
rect 4619 4392 4685 4408
rect 4619 4328 4620 4392
rect 4684 4328 4685 4392
rect 4619 4312 4685 4328
rect 4619 4248 4620 4312
rect 4684 4248 4685 4312
rect 4619 4232 4685 4248
rect 4619 4168 4620 4232
rect 4684 4168 4685 4232
rect 4619 4152 4685 4168
rect 4619 4088 4620 4152
rect 4684 4088 4685 4152
rect 4619 3934 4685 4088
rect 4745 3996 4805 5026
rect 4865 3934 4925 4966
rect 4985 3996 5045 5026
rect 5105 3934 5165 4966
rect 5225 4872 5291 4962
rect 5225 4808 5226 4872
rect 5290 4808 5291 4872
rect 5225 4792 5291 4808
rect 5225 4728 5226 4792
rect 5290 4728 5291 4792
rect 5225 4712 5291 4728
rect 5225 4648 5226 4712
rect 5290 4648 5291 4712
rect 5225 4632 5291 4648
rect 5225 4568 5226 4632
rect 5290 4568 5291 4632
rect 5225 4552 5291 4568
rect 5225 4488 5226 4552
rect 5290 4488 5291 4552
rect 5225 4472 5291 4488
rect 5225 4408 5226 4472
rect 5290 4408 5291 4472
rect 5225 4392 5291 4408
rect 5225 4328 5226 4392
rect 5290 4328 5291 4392
rect 5225 4312 5291 4328
rect 5225 4248 5226 4312
rect 5290 4248 5291 4312
rect 5225 4232 5291 4248
rect 5225 4168 5226 4232
rect 5290 4168 5291 4232
rect 5225 4152 5291 4168
rect 5225 4088 5226 4152
rect 5290 4088 5291 4152
rect 5225 3934 5291 4088
rect 2801 3932 5291 3934
rect 2801 3868 2905 3932
rect 2969 3868 2985 3932
rect 3049 3868 3065 3932
rect 3129 3868 3145 3932
rect 3209 3868 3225 3932
rect 3289 3868 3305 3932
rect 3369 3868 3511 3932
rect 3575 3868 3591 3932
rect 3655 3868 3671 3932
rect 3735 3868 3751 3932
rect 3815 3868 3831 3932
rect 3895 3868 3911 3932
rect 3975 3868 4117 3932
rect 4181 3868 4197 3932
rect 4261 3868 4277 3932
rect 4341 3868 4357 3932
rect 4421 3868 4437 3932
rect 4501 3868 4517 3932
rect 4581 3868 4723 3932
rect 4787 3868 4803 3932
rect 4867 3868 4883 3932
rect 4947 3868 4963 3932
rect 5027 3868 5043 3932
rect 5107 3868 5123 3932
rect 5187 3868 5291 3932
rect 2801 3866 5291 3868
rect 2801 3712 2867 3866
rect 2801 3648 2802 3712
rect 2866 3648 2867 3712
rect 2801 3632 2867 3648
rect 2801 3568 2802 3632
rect 2866 3568 2867 3632
rect 2801 3552 2867 3568
rect 2801 3488 2802 3552
rect 2866 3488 2867 3552
rect 2801 3472 2867 3488
rect 2801 3408 2802 3472
rect 2866 3408 2867 3472
rect 2801 3392 2867 3408
rect 2801 3328 2802 3392
rect 2866 3328 2867 3392
rect 2801 3312 2867 3328
rect 2801 3248 2802 3312
rect 2866 3248 2867 3312
rect 2801 3232 2867 3248
rect 2801 3168 2802 3232
rect 2866 3168 2867 3232
rect 2801 3152 2867 3168
rect 2801 3088 2802 3152
rect 2866 3088 2867 3152
rect 2801 3072 2867 3088
rect 2801 3008 2802 3072
rect 2866 3008 2867 3072
rect 2801 2992 2867 3008
rect 2801 2928 2802 2992
rect 2866 2928 2867 2992
rect 2801 2838 2867 2928
rect 2927 2834 2987 3866
rect 3047 2774 3107 3804
rect 3167 2834 3227 3866
rect 3287 2774 3347 3804
rect 3407 3712 3473 3866
rect 3407 3648 3408 3712
rect 3472 3648 3473 3712
rect 3407 3632 3473 3648
rect 3407 3568 3408 3632
rect 3472 3568 3473 3632
rect 3407 3552 3473 3568
rect 3407 3488 3408 3552
rect 3472 3488 3473 3552
rect 3407 3472 3473 3488
rect 3407 3408 3408 3472
rect 3472 3408 3473 3472
rect 3407 3392 3473 3408
rect 3407 3328 3408 3392
rect 3472 3328 3473 3392
rect 3407 3312 3473 3328
rect 3407 3248 3408 3312
rect 3472 3248 3473 3312
rect 3407 3232 3473 3248
rect 3407 3168 3408 3232
rect 3472 3168 3473 3232
rect 3407 3152 3473 3168
rect 3407 3088 3408 3152
rect 3472 3088 3473 3152
rect 3407 3072 3473 3088
rect 3407 3008 3408 3072
rect 3472 3008 3473 3072
rect 3407 2992 3473 3008
rect 3407 2928 3408 2992
rect 3472 2928 3473 2992
rect 3407 2838 3473 2928
rect 3533 2834 3593 3866
rect 3653 2774 3713 3804
rect 3773 2834 3833 3866
rect 3893 2774 3953 3804
rect 4013 3712 4079 3866
rect 4013 3648 4014 3712
rect 4078 3648 4079 3712
rect 4013 3632 4079 3648
rect 4013 3568 4014 3632
rect 4078 3568 4079 3632
rect 4013 3552 4079 3568
rect 4013 3488 4014 3552
rect 4078 3488 4079 3552
rect 4013 3472 4079 3488
rect 4013 3408 4014 3472
rect 4078 3408 4079 3472
rect 4013 3392 4079 3408
rect 4013 3328 4014 3392
rect 4078 3328 4079 3392
rect 4013 3312 4079 3328
rect 4013 3248 4014 3312
rect 4078 3248 4079 3312
rect 4013 3232 4079 3248
rect 4013 3168 4014 3232
rect 4078 3168 4079 3232
rect 4013 3152 4079 3168
rect 4013 3088 4014 3152
rect 4078 3088 4079 3152
rect 4013 3072 4079 3088
rect 4013 3008 4014 3072
rect 4078 3008 4079 3072
rect 4013 2992 4079 3008
rect 4013 2928 4014 2992
rect 4078 2928 4079 2992
rect 4013 2838 4079 2928
rect 4139 2834 4199 3866
rect 4259 2774 4319 3804
rect 4379 2834 4439 3866
rect 4499 2774 4559 3804
rect 4619 3712 4685 3866
rect 4619 3648 4620 3712
rect 4684 3648 4685 3712
rect 4619 3632 4685 3648
rect 4619 3568 4620 3632
rect 4684 3568 4685 3632
rect 4619 3552 4685 3568
rect 4619 3488 4620 3552
rect 4684 3488 4685 3552
rect 4619 3472 4685 3488
rect 4619 3408 4620 3472
rect 4684 3408 4685 3472
rect 4619 3392 4685 3408
rect 4619 3328 4620 3392
rect 4684 3328 4685 3392
rect 4619 3312 4685 3328
rect 4619 3248 4620 3312
rect 4684 3248 4685 3312
rect 4619 3232 4685 3248
rect 4619 3168 4620 3232
rect 4684 3168 4685 3232
rect 4619 3152 4685 3168
rect 4619 3088 4620 3152
rect 4684 3088 4685 3152
rect 4619 3072 4685 3088
rect 4619 3008 4620 3072
rect 4684 3008 4685 3072
rect 4619 2992 4685 3008
rect 4619 2928 4620 2992
rect 4684 2928 4685 2992
rect 4619 2838 4685 2928
rect 4745 2834 4805 3866
rect 4865 2774 4925 3804
rect 4985 2834 5045 3866
rect 5105 2774 5165 3804
rect 5225 3712 5291 3866
rect 5225 3648 5226 3712
rect 5290 3648 5291 3712
rect 5225 3632 5291 3648
rect 5225 3568 5226 3632
rect 5290 3568 5291 3632
rect 5225 3552 5291 3568
rect 5225 3488 5226 3552
rect 5290 3488 5291 3552
rect 5225 3472 5291 3488
rect 5225 3408 5226 3472
rect 5290 3408 5291 3472
rect 5225 3392 5291 3408
rect 5225 3328 5226 3392
rect 5290 3328 5291 3392
rect 5225 3312 5291 3328
rect 5225 3248 5226 3312
rect 5290 3248 5291 3312
rect 5225 3232 5291 3248
rect 5225 3168 5226 3232
rect 5290 3168 5291 3232
rect 5225 3152 5291 3168
rect 5225 3088 5226 3152
rect 5290 3088 5291 3152
rect 5225 3072 5291 3088
rect 5225 3008 5226 3072
rect 5290 3008 5291 3072
rect 5225 2992 5291 3008
rect 5225 2928 5226 2992
rect 5290 2928 5291 2992
rect 5225 2838 5291 2928
rect 5352 4872 5418 4962
rect 5352 4808 5353 4872
rect 5417 4808 5418 4872
rect 5352 4792 5418 4808
rect 5352 4728 5353 4792
rect 5417 4728 5418 4792
rect 5352 4712 5418 4728
rect 5352 4648 5353 4712
rect 5417 4648 5418 4712
rect 5352 4632 5418 4648
rect 5352 4568 5353 4632
rect 5417 4568 5418 4632
rect 5352 4552 5418 4568
rect 5352 4488 5353 4552
rect 5417 4488 5418 4552
rect 5352 4472 5418 4488
rect 5352 4408 5353 4472
rect 5417 4408 5418 4472
rect 5352 4392 5418 4408
rect 5352 4328 5353 4392
rect 5417 4328 5418 4392
rect 5352 4312 5418 4328
rect 5352 4248 5353 4312
rect 5417 4248 5418 4312
rect 5352 4232 5418 4248
rect 5352 4168 5353 4232
rect 5417 4168 5418 4232
rect 5352 4152 5418 4168
rect 5352 4088 5353 4152
rect 5417 4088 5418 4152
rect 5352 3934 5418 4088
rect 5478 3996 5538 5026
rect 5598 3934 5658 4966
rect 5718 3996 5778 5026
rect 5838 3934 5898 4966
rect 5958 4872 6024 4962
rect 5958 4808 5959 4872
rect 6023 4808 6024 4872
rect 5958 4792 6024 4808
rect 5958 4728 5959 4792
rect 6023 4728 6024 4792
rect 5958 4712 6024 4728
rect 5958 4648 5959 4712
rect 6023 4648 6024 4712
rect 5958 4632 6024 4648
rect 5958 4568 5959 4632
rect 6023 4568 6024 4632
rect 5958 4552 6024 4568
rect 5958 4488 5959 4552
rect 6023 4488 6024 4552
rect 5958 4472 6024 4488
rect 5958 4408 5959 4472
rect 6023 4408 6024 4472
rect 5958 4392 6024 4408
rect 5958 4328 5959 4392
rect 6023 4328 6024 4392
rect 5958 4312 6024 4328
rect 5958 4248 5959 4312
rect 6023 4248 6024 4312
rect 5958 4232 6024 4248
rect 5958 4168 5959 4232
rect 6023 4168 6024 4232
rect 5958 4152 6024 4168
rect 5958 4088 5959 4152
rect 6023 4088 6024 4152
rect 5958 3934 6024 4088
rect 6084 3996 6144 5026
rect 6204 3934 6264 4966
rect 6324 3996 6384 5026
rect 6444 3934 6504 4966
rect 6564 4872 6630 4962
rect 6564 4808 6565 4872
rect 6629 4808 6630 4872
rect 6564 4792 6630 4808
rect 6564 4728 6565 4792
rect 6629 4728 6630 4792
rect 6564 4712 6630 4728
rect 6564 4648 6565 4712
rect 6629 4648 6630 4712
rect 6564 4632 6630 4648
rect 6564 4568 6565 4632
rect 6629 4568 6630 4632
rect 6564 4552 6630 4568
rect 6564 4488 6565 4552
rect 6629 4488 6630 4552
rect 6564 4472 6630 4488
rect 6564 4408 6565 4472
rect 6629 4408 6630 4472
rect 6564 4392 6630 4408
rect 6564 4328 6565 4392
rect 6629 4328 6630 4392
rect 6564 4312 6630 4328
rect 6564 4248 6565 4312
rect 6629 4248 6630 4312
rect 6564 4232 6630 4248
rect 6564 4168 6565 4232
rect 6629 4168 6630 4232
rect 6564 4152 6630 4168
rect 6564 4088 6565 4152
rect 6629 4088 6630 4152
rect 6564 3934 6630 4088
rect 6690 3996 6750 5026
rect 6810 3934 6870 4966
rect 6930 3996 6990 5026
rect 7050 3934 7110 4966
rect 7170 4872 7236 4962
rect 7170 4808 7171 4872
rect 7235 4808 7236 4872
rect 7170 4792 7236 4808
rect 7170 4728 7171 4792
rect 7235 4728 7236 4792
rect 7170 4712 7236 4728
rect 7170 4648 7171 4712
rect 7235 4648 7236 4712
rect 7170 4632 7236 4648
rect 7170 4568 7171 4632
rect 7235 4568 7236 4632
rect 7170 4552 7236 4568
rect 7170 4488 7171 4552
rect 7235 4488 7236 4552
rect 7170 4472 7236 4488
rect 7170 4408 7171 4472
rect 7235 4408 7236 4472
rect 7170 4392 7236 4408
rect 7170 4328 7171 4392
rect 7235 4328 7236 4392
rect 7170 4312 7236 4328
rect 7170 4248 7171 4312
rect 7235 4248 7236 4312
rect 7170 4232 7236 4248
rect 7170 4168 7171 4232
rect 7235 4168 7236 4232
rect 7170 4152 7236 4168
rect 7170 4088 7171 4152
rect 7235 4088 7236 4152
rect 7170 3934 7236 4088
rect 7296 3996 7356 5026
rect 7416 3934 7476 4966
rect 7536 3996 7596 5026
rect 7656 3934 7716 4966
rect 7776 4872 7842 4962
rect 7776 4808 7777 4872
rect 7841 4808 7842 4872
rect 7776 4792 7842 4808
rect 7776 4728 7777 4792
rect 7841 4728 7842 4792
rect 7776 4712 7842 4728
rect 7776 4648 7777 4712
rect 7841 4648 7842 4712
rect 7776 4632 7842 4648
rect 7776 4568 7777 4632
rect 7841 4568 7842 4632
rect 7776 4552 7842 4568
rect 7776 4488 7777 4552
rect 7841 4488 7842 4552
rect 7776 4472 7842 4488
rect 7776 4408 7777 4472
rect 7841 4408 7842 4472
rect 7776 4392 7842 4408
rect 7776 4328 7777 4392
rect 7841 4328 7842 4392
rect 7776 4312 7842 4328
rect 7776 4248 7777 4312
rect 7841 4248 7842 4312
rect 7776 4232 7842 4248
rect 7776 4168 7777 4232
rect 7841 4168 7842 4232
rect 7776 4152 7842 4168
rect 7776 4088 7777 4152
rect 7841 4088 7842 4152
rect 7776 3934 7842 4088
rect 7902 3996 7962 5026
rect 8022 3934 8082 4966
rect 8142 3996 8202 5026
rect 8262 3934 8322 4966
rect 8382 4872 8448 4962
rect 8382 4808 8383 4872
rect 8447 4808 8448 4872
rect 8382 4792 8448 4808
rect 8382 4728 8383 4792
rect 8447 4728 8448 4792
rect 8382 4712 8448 4728
rect 8382 4648 8383 4712
rect 8447 4648 8448 4712
rect 8382 4632 8448 4648
rect 8382 4568 8383 4632
rect 8447 4568 8448 4632
rect 8382 4552 8448 4568
rect 8382 4488 8383 4552
rect 8447 4488 8448 4552
rect 8382 4472 8448 4488
rect 8382 4408 8383 4472
rect 8447 4408 8448 4472
rect 8382 4392 8448 4408
rect 8382 4328 8383 4392
rect 8447 4328 8448 4392
rect 8382 4312 8448 4328
rect 8382 4248 8383 4312
rect 8447 4248 8448 4312
rect 8382 4232 8448 4248
rect 8382 4168 8383 4232
rect 8447 4168 8448 4232
rect 8382 4152 8448 4168
rect 8382 4088 8383 4152
rect 8447 4088 8448 4152
rect 8382 3934 8448 4088
rect 8508 3996 8568 5026
rect 8628 3934 8688 4966
rect 8748 3996 8808 5026
rect 8868 3934 8928 4966
rect 8988 4872 9054 4962
rect 8988 4808 8989 4872
rect 9053 4808 9054 4872
rect 8988 4792 9054 4808
rect 8988 4728 8989 4792
rect 9053 4728 9054 4792
rect 8988 4712 9054 4728
rect 8988 4648 8989 4712
rect 9053 4648 9054 4712
rect 8988 4632 9054 4648
rect 8988 4568 8989 4632
rect 9053 4568 9054 4632
rect 8988 4552 9054 4568
rect 8988 4488 8989 4552
rect 9053 4488 9054 4552
rect 8988 4472 9054 4488
rect 8988 4408 8989 4472
rect 9053 4408 9054 4472
rect 8988 4392 9054 4408
rect 8988 4328 8989 4392
rect 9053 4328 9054 4392
rect 8988 4312 9054 4328
rect 8988 4248 8989 4312
rect 9053 4248 9054 4312
rect 8988 4232 9054 4248
rect 8988 4168 8989 4232
rect 9053 4168 9054 4232
rect 8988 4152 9054 4168
rect 8988 4088 8989 4152
rect 9053 4088 9054 4152
rect 8988 3934 9054 4088
rect 9114 3996 9174 5026
rect 9234 3934 9294 4966
rect 9354 3996 9414 5026
rect 9474 3934 9534 4966
rect 9594 4872 9660 4962
rect 9594 4808 9595 4872
rect 9659 4808 9660 4872
rect 9594 4792 9660 4808
rect 9594 4728 9595 4792
rect 9659 4728 9660 4792
rect 9594 4712 9660 4728
rect 9594 4648 9595 4712
rect 9659 4648 9660 4712
rect 9594 4632 9660 4648
rect 9594 4568 9595 4632
rect 9659 4568 9660 4632
rect 9594 4552 9660 4568
rect 9594 4488 9595 4552
rect 9659 4488 9660 4552
rect 9594 4472 9660 4488
rect 9594 4408 9595 4472
rect 9659 4408 9660 4472
rect 9594 4392 9660 4408
rect 9594 4328 9595 4392
rect 9659 4328 9660 4392
rect 9594 4312 9660 4328
rect 9594 4248 9595 4312
rect 9659 4248 9660 4312
rect 9594 4232 9660 4248
rect 9594 4168 9595 4232
rect 9659 4168 9660 4232
rect 9594 4152 9660 4168
rect 9594 4088 9595 4152
rect 9659 4088 9660 4152
rect 9594 3934 9660 4088
rect 9720 3996 9780 5026
rect 9840 3934 9900 4966
rect 9960 3996 10020 5026
rect 10080 3934 10140 4966
rect 10200 4872 10266 4962
rect 10200 4808 10201 4872
rect 10265 4808 10266 4872
rect 10200 4792 10266 4808
rect 10200 4728 10201 4792
rect 10265 4728 10266 4792
rect 10200 4712 10266 4728
rect 10200 4648 10201 4712
rect 10265 4648 10266 4712
rect 10200 4632 10266 4648
rect 10200 4568 10201 4632
rect 10265 4568 10266 4632
rect 10200 4552 10266 4568
rect 10200 4488 10201 4552
rect 10265 4488 10266 4552
rect 10200 4472 10266 4488
rect 10200 4408 10201 4472
rect 10265 4408 10266 4472
rect 10200 4392 10266 4408
rect 10200 4328 10201 4392
rect 10265 4328 10266 4392
rect 10200 4312 10266 4328
rect 10200 4248 10201 4312
rect 10265 4248 10266 4312
rect 10200 4232 10266 4248
rect 10200 4168 10201 4232
rect 10265 4168 10266 4232
rect 10200 4152 10266 4168
rect 10200 4088 10201 4152
rect 10265 4088 10266 4152
rect 10200 3934 10266 4088
rect 5352 3932 10266 3934
rect 5352 3868 5456 3932
rect 5520 3868 5536 3932
rect 5600 3868 5616 3932
rect 5680 3868 5696 3932
rect 5760 3868 5776 3932
rect 5840 3868 5856 3932
rect 5920 3868 6062 3932
rect 6126 3868 6142 3932
rect 6206 3868 6222 3932
rect 6286 3868 6302 3932
rect 6366 3868 6382 3932
rect 6446 3868 6462 3932
rect 6526 3868 6668 3932
rect 6732 3868 6748 3932
rect 6812 3868 6828 3932
rect 6892 3868 6908 3932
rect 6972 3868 6988 3932
rect 7052 3868 7068 3932
rect 7132 3868 7274 3932
rect 7338 3868 7354 3932
rect 7418 3868 7434 3932
rect 7498 3868 7514 3932
rect 7578 3868 7594 3932
rect 7658 3868 7674 3932
rect 7738 3868 7880 3932
rect 7944 3868 7960 3932
rect 8024 3868 8040 3932
rect 8104 3868 8120 3932
rect 8184 3868 8200 3932
rect 8264 3868 8280 3932
rect 8344 3868 8486 3932
rect 8550 3868 8566 3932
rect 8630 3868 8646 3932
rect 8710 3868 8726 3932
rect 8790 3868 8806 3932
rect 8870 3868 8886 3932
rect 8950 3868 9092 3932
rect 9156 3868 9172 3932
rect 9236 3868 9252 3932
rect 9316 3868 9332 3932
rect 9396 3868 9412 3932
rect 9476 3868 9492 3932
rect 9556 3868 9698 3932
rect 9762 3868 9778 3932
rect 9842 3868 9858 3932
rect 9922 3868 9938 3932
rect 10002 3868 10018 3932
rect 10082 3868 10098 3932
rect 10162 3868 10266 3932
rect 5352 3866 10266 3868
rect 5352 3712 5418 3866
rect 5352 3648 5353 3712
rect 5417 3648 5418 3712
rect 5352 3632 5418 3648
rect 5352 3568 5353 3632
rect 5417 3568 5418 3632
rect 5352 3552 5418 3568
rect 5352 3488 5353 3552
rect 5417 3488 5418 3552
rect 5352 3472 5418 3488
rect 5352 3408 5353 3472
rect 5417 3408 5418 3472
rect 5352 3392 5418 3408
rect 5352 3328 5353 3392
rect 5417 3328 5418 3392
rect 5352 3312 5418 3328
rect 5352 3248 5353 3312
rect 5417 3248 5418 3312
rect 5352 3232 5418 3248
rect 5352 3168 5353 3232
rect 5417 3168 5418 3232
rect 5352 3152 5418 3168
rect 5352 3088 5353 3152
rect 5417 3088 5418 3152
rect 5352 3072 5418 3088
rect 5352 3008 5353 3072
rect 5417 3008 5418 3072
rect 5352 2992 5418 3008
rect 5352 2928 5353 2992
rect 5417 2928 5418 2992
rect 5352 2838 5418 2928
rect 5478 2834 5538 3866
rect 5598 2774 5658 3804
rect 5718 2834 5778 3866
rect 5838 2774 5898 3804
rect 5958 3712 6024 3866
rect 5958 3648 5959 3712
rect 6023 3648 6024 3712
rect 5958 3632 6024 3648
rect 5958 3568 5959 3632
rect 6023 3568 6024 3632
rect 5958 3552 6024 3568
rect 5958 3488 5959 3552
rect 6023 3488 6024 3552
rect 5958 3472 6024 3488
rect 5958 3408 5959 3472
rect 6023 3408 6024 3472
rect 5958 3392 6024 3408
rect 5958 3328 5959 3392
rect 6023 3328 6024 3392
rect 5958 3312 6024 3328
rect 5958 3248 5959 3312
rect 6023 3248 6024 3312
rect 5958 3232 6024 3248
rect 5958 3168 5959 3232
rect 6023 3168 6024 3232
rect 5958 3152 6024 3168
rect 5958 3088 5959 3152
rect 6023 3088 6024 3152
rect 5958 3072 6024 3088
rect 5958 3008 5959 3072
rect 6023 3008 6024 3072
rect 5958 2992 6024 3008
rect 5958 2928 5959 2992
rect 6023 2928 6024 2992
rect 5958 2838 6024 2928
rect 6084 2834 6144 3866
rect 6204 2774 6264 3804
rect 6324 2834 6384 3866
rect 6444 2774 6504 3804
rect 6564 3712 6630 3866
rect 6564 3648 6565 3712
rect 6629 3648 6630 3712
rect 6564 3632 6630 3648
rect 6564 3568 6565 3632
rect 6629 3568 6630 3632
rect 6564 3552 6630 3568
rect 6564 3488 6565 3552
rect 6629 3488 6630 3552
rect 6564 3472 6630 3488
rect 6564 3408 6565 3472
rect 6629 3408 6630 3472
rect 6564 3392 6630 3408
rect 6564 3328 6565 3392
rect 6629 3328 6630 3392
rect 6564 3312 6630 3328
rect 6564 3248 6565 3312
rect 6629 3248 6630 3312
rect 6564 3232 6630 3248
rect 6564 3168 6565 3232
rect 6629 3168 6630 3232
rect 6564 3152 6630 3168
rect 6564 3088 6565 3152
rect 6629 3088 6630 3152
rect 6564 3072 6630 3088
rect 6564 3008 6565 3072
rect 6629 3008 6630 3072
rect 6564 2992 6630 3008
rect 6564 2928 6565 2992
rect 6629 2928 6630 2992
rect 6564 2838 6630 2928
rect 6690 2834 6750 3866
rect 6810 2774 6870 3804
rect 6930 2834 6990 3866
rect 7050 2774 7110 3804
rect 7170 3712 7236 3866
rect 7170 3648 7171 3712
rect 7235 3648 7236 3712
rect 7170 3632 7236 3648
rect 7170 3568 7171 3632
rect 7235 3568 7236 3632
rect 7170 3552 7236 3568
rect 7170 3488 7171 3552
rect 7235 3488 7236 3552
rect 7170 3472 7236 3488
rect 7170 3408 7171 3472
rect 7235 3408 7236 3472
rect 7170 3392 7236 3408
rect 7170 3328 7171 3392
rect 7235 3328 7236 3392
rect 7170 3312 7236 3328
rect 7170 3248 7171 3312
rect 7235 3248 7236 3312
rect 7170 3232 7236 3248
rect 7170 3168 7171 3232
rect 7235 3168 7236 3232
rect 7170 3152 7236 3168
rect 7170 3088 7171 3152
rect 7235 3088 7236 3152
rect 7170 3072 7236 3088
rect 7170 3008 7171 3072
rect 7235 3008 7236 3072
rect 7170 2992 7236 3008
rect 7170 2928 7171 2992
rect 7235 2928 7236 2992
rect 7170 2838 7236 2928
rect 7296 2834 7356 3866
rect 7416 2774 7476 3804
rect 7536 2834 7596 3866
rect 7656 2774 7716 3804
rect 7776 3712 7842 3866
rect 7776 3648 7777 3712
rect 7841 3648 7842 3712
rect 7776 3632 7842 3648
rect 7776 3568 7777 3632
rect 7841 3568 7842 3632
rect 7776 3552 7842 3568
rect 7776 3488 7777 3552
rect 7841 3488 7842 3552
rect 7776 3472 7842 3488
rect 7776 3408 7777 3472
rect 7841 3408 7842 3472
rect 7776 3392 7842 3408
rect 7776 3328 7777 3392
rect 7841 3328 7842 3392
rect 7776 3312 7842 3328
rect 7776 3248 7777 3312
rect 7841 3248 7842 3312
rect 7776 3232 7842 3248
rect 7776 3168 7777 3232
rect 7841 3168 7842 3232
rect 7776 3152 7842 3168
rect 7776 3088 7777 3152
rect 7841 3088 7842 3152
rect 7776 3072 7842 3088
rect 7776 3008 7777 3072
rect 7841 3008 7842 3072
rect 7776 2992 7842 3008
rect 7776 2928 7777 2992
rect 7841 2928 7842 2992
rect 7776 2838 7842 2928
rect 7902 2834 7962 3866
rect 8022 2774 8082 3804
rect 8142 2834 8202 3866
rect 8262 2774 8322 3804
rect 8382 3712 8448 3866
rect 8382 3648 8383 3712
rect 8447 3648 8448 3712
rect 8382 3632 8448 3648
rect 8382 3568 8383 3632
rect 8447 3568 8448 3632
rect 8382 3552 8448 3568
rect 8382 3488 8383 3552
rect 8447 3488 8448 3552
rect 8382 3472 8448 3488
rect 8382 3408 8383 3472
rect 8447 3408 8448 3472
rect 8382 3392 8448 3408
rect 8382 3328 8383 3392
rect 8447 3328 8448 3392
rect 8382 3312 8448 3328
rect 8382 3248 8383 3312
rect 8447 3248 8448 3312
rect 8382 3232 8448 3248
rect 8382 3168 8383 3232
rect 8447 3168 8448 3232
rect 8382 3152 8448 3168
rect 8382 3088 8383 3152
rect 8447 3088 8448 3152
rect 8382 3072 8448 3088
rect 8382 3008 8383 3072
rect 8447 3008 8448 3072
rect 8382 2992 8448 3008
rect 8382 2928 8383 2992
rect 8447 2928 8448 2992
rect 8382 2838 8448 2928
rect 8508 2834 8568 3866
rect 8628 2774 8688 3804
rect 8748 2834 8808 3866
rect 8868 2774 8928 3804
rect 8988 3712 9054 3866
rect 8988 3648 8989 3712
rect 9053 3648 9054 3712
rect 8988 3632 9054 3648
rect 8988 3568 8989 3632
rect 9053 3568 9054 3632
rect 8988 3552 9054 3568
rect 8988 3488 8989 3552
rect 9053 3488 9054 3552
rect 8988 3472 9054 3488
rect 8988 3408 8989 3472
rect 9053 3408 9054 3472
rect 8988 3392 9054 3408
rect 8988 3328 8989 3392
rect 9053 3328 9054 3392
rect 8988 3312 9054 3328
rect 8988 3248 8989 3312
rect 9053 3248 9054 3312
rect 8988 3232 9054 3248
rect 8988 3168 8989 3232
rect 9053 3168 9054 3232
rect 8988 3152 9054 3168
rect 8988 3088 8989 3152
rect 9053 3088 9054 3152
rect 8988 3072 9054 3088
rect 8988 3008 8989 3072
rect 9053 3008 9054 3072
rect 8988 2992 9054 3008
rect 8988 2928 8989 2992
rect 9053 2928 9054 2992
rect 8988 2838 9054 2928
rect 9114 2834 9174 3866
rect 9234 2774 9294 3804
rect 9354 2834 9414 3866
rect 9474 2774 9534 3804
rect 9594 3712 9660 3866
rect 9594 3648 9595 3712
rect 9659 3648 9660 3712
rect 9594 3632 9660 3648
rect 9594 3568 9595 3632
rect 9659 3568 9660 3632
rect 9594 3552 9660 3568
rect 9594 3488 9595 3552
rect 9659 3488 9660 3552
rect 9594 3472 9660 3488
rect 9594 3408 9595 3472
rect 9659 3408 9660 3472
rect 9594 3392 9660 3408
rect 9594 3328 9595 3392
rect 9659 3328 9660 3392
rect 9594 3312 9660 3328
rect 9594 3248 9595 3312
rect 9659 3248 9660 3312
rect 9594 3232 9660 3248
rect 9594 3168 9595 3232
rect 9659 3168 9660 3232
rect 9594 3152 9660 3168
rect 9594 3088 9595 3152
rect 9659 3088 9660 3152
rect 9594 3072 9660 3088
rect 9594 3008 9595 3072
rect 9659 3008 9660 3072
rect 9594 2992 9660 3008
rect 9594 2928 9595 2992
rect 9659 2928 9660 2992
rect 9594 2838 9660 2928
rect 9720 2834 9780 3866
rect 9840 2774 9900 3804
rect 9960 2834 10020 3866
rect 10080 2774 10140 3804
rect 10200 3712 10266 3866
rect 10200 3648 10201 3712
rect 10265 3648 10266 3712
rect 10200 3632 10266 3648
rect 10200 3568 10201 3632
rect 10265 3568 10266 3632
rect 10200 3552 10266 3568
rect 10200 3488 10201 3552
rect 10265 3488 10266 3552
rect 10200 3472 10266 3488
rect 10200 3408 10201 3472
rect 10265 3408 10266 3472
rect 10200 3392 10266 3408
rect 10200 3328 10201 3392
rect 10265 3328 10266 3392
rect 10200 3312 10266 3328
rect 10200 3248 10201 3312
rect 10265 3248 10266 3312
rect 10200 3232 10266 3248
rect 10200 3168 10201 3232
rect 10265 3168 10266 3232
rect 10200 3152 10266 3168
rect 10200 3088 10201 3152
rect 10265 3088 10266 3152
rect 10200 3072 10266 3088
rect 10200 3008 10201 3072
rect 10265 3008 10266 3072
rect 10200 2992 10266 3008
rect 10200 2928 10201 2992
rect 10265 2928 10266 2992
rect 10200 2838 10266 2928
rect 10326 4872 10392 4962
rect 10326 4808 10327 4872
rect 10391 4808 10392 4872
rect 10326 4792 10392 4808
rect 10326 4728 10327 4792
rect 10391 4728 10392 4792
rect 10326 4712 10392 4728
rect 10326 4648 10327 4712
rect 10391 4648 10392 4712
rect 10326 4632 10392 4648
rect 10326 4568 10327 4632
rect 10391 4568 10392 4632
rect 10326 4552 10392 4568
rect 10326 4488 10327 4552
rect 10391 4488 10392 4552
rect 10326 4472 10392 4488
rect 10326 4408 10327 4472
rect 10391 4408 10392 4472
rect 10326 4392 10392 4408
rect 10326 4328 10327 4392
rect 10391 4328 10392 4392
rect 10326 4312 10392 4328
rect 10326 4248 10327 4312
rect 10391 4248 10392 4312
rect 10326 4232 10392 4248
rect 10326 4168 10327 4232
rect 10391 4168 10392 4232
rect 10326 4152 10392 4168
rect 10326 4088 10327 4152
rect 10391 4088 10392 4152
rect 10326 3934 10392 4088
rect 10452 3996 10512 5026
rect 10572 3934 10632 4966
rect 10692 3996 10752 5026
rect 10812 3934 10872 4966
rect 10932 4872 10998 4962
rect 10932 4808 10933 4872
rect 10997 4808 10998 4872
rect 10932 4792 10998 4808
rect 10932 4728 10933 4792
rect 10997 4728 10998 4792
rect 10932 4712 10998 4728
rect 10932 4648 10933 4712
rect 10997 4648 10998 4712
rect 10932 4632 10998 4648
rect 10932 4568 10933 4632
rect 10997 4568 10998 4632
rect 10932 4552 10998 4568
rect 10932 4488 10933 4552
rect 10997 4488 10998 4552
rect 10932 4472 10998 4488
rect 10932 4408 10933 4472
rect 10997 4408 10998 4472
rect 10932 4392 10998 4408
rect 10932 4328 10933 4392
rect 10997 4328 10998 4392
rect 10932 4312 10998 4328
rect 10932 4248 10933 4312
rect 10997 4248 10998 4312
rect 10932 4232 10998 4248
rect 10932 4168 10933 4232
rect 10997 4168 10998 4232
rect 10932 4152 10998 4168
rect 10932 4088 10933 4152
rect 10997 4088 10998 4152
rect 10932 3934 10998 4088
rect 11058 3996 11118 5026
rect 11178 3934 11238 4966
rect 11298 3996 11358 5026
rect 11418 3934 11478 4966
rect 11538 4872 11604 4962
rect 11538 4808 11539 4872
rect 11603 4808 11604 4872
rect 11538 4792 11604 4808
rect 11538 4728 11539 4792
rect 11603 4728 11604 4792
rect 11538 4712 11604 4728
rect 11538 4648 11539 4712
rect 11603 4648 11604 4712
rect 11538 4632 11604 4648
rect 11538 4568 11539 4632
rect 11603 4568 11604 4632
rect 11538 4552 11604 4568
rect 11538 4488 11539 4552
rect 11603 4488 11604 4552
rect 11538 4472 11604 4488
rect 11538 4408 11539 4472
rect 11603 4408 11604 4472
rect 11538 4392 11604 4408
rect 11538 4328 11539 4392
rect 11603 4328 11604 4392
rect 11538 4312 11604 4328
rect 11538 4248 11539 4312
rect 11603 4248 11604 4312
rect 11538 4232 11604 4248
rect 11538 4168 11539 4232
rect 11603 4168 11604 4232
rect 11538 4152 11604 4168
rect 11538 4088 11539 4152
rect 11603 4088 11604 4152
rect 11538 3934 11604 4088
rect 11664 3996 11724 5026
rect 11784 3934 11844 4966
rect 11904 3996 11964 5026
rect 12024 3934 12084 4966
rect 12144 4872 12210 4962
rect 12144 4808 12145 4872
rect 12209 4808 12210 4872
rect 12144 4792 12210 4808
rect 12144 4728 12145 4792
rect 12209 4728 12210 4792
rect 12144 4712 12210 4728
rect 12144 4648 12145 4712
rect 12209 4648 12210 4712
rect 12144 4632 12210 4648
rect 12144 4568 12145 4632
rect 12209 4568 12210 4632
rect 12144 4552 12210 4568
rect 12144 4488 12145 4552
rect 12209 4488 12210 4552
rect 12144 4472 12210 4488
rect 12144 4408 12145 4472
rect 12209 4408 12210 4472
rect 12144 4392 12210 4408
rect 12144 4328 12145 4392
rect 12209 4328 12210 4392
rect 12144 4312 12210 4328
rect 12144 4248 12145 4312
rect 12209 4248 12210 4312
rect 12144 4232 12210 4248
rect 12144 4168 12145 4232
rect 12209 4168 12210 4232
rect 12144 4152 12210 4168
rect 12144 4088 12145 4152
rect 12209 4088 12210 4152
rect 12144 3934 12210 4088
rect 12270 3996 12330 5026
rect 12390 3934 12450 4966
rect 12510 3996 12570 5026
rect 12630 3934 12690 4966
rect 12750 4872 12816 4962
rect 12750 4808 12751 4872
rect 12815 4808 12816 4872
rect 12750 4792 12816 4808
rect 12750 4728 12751 4792
rect 12815 4728 12816 4792
rect 12750 4712 12816 4728
rect 12750 4648 12751 4712
rect 12815 4648 12816 4712
rect 12750 4632 12816 4648
rect 12750 4568 12751 4632
rect 12815 4568 12816 4632
rect 12750 4552 12816 4568
rect 12750 4488 12751 4552
rect 12815 4488 12816 4552
rect 12750 4472 12816 4488
rect 12750 4408 12751 4472
rect 12815 4408 12816 4472
rect 12750 4392 12816 4408
rect 12750 4328 12751 4392
rect 12815 4328 12816 4392
rect 12750 4312 12816 4328
rect 12750 4248 12751 4312
rect 12815 4248 12816 4312
rect 12750 4232 12816 4248
rect 12750 4168 12751 4232
rect 12815 4168 12816 4232
rect 12750 4152 12816 4168
rect 12750 4088 12751 4152
rect 12815 4088 12816 4152
rect 12750 3934 12816 4088
rect 12876 3996 12936 5026
rect 12996 3934 13056 4966
rect 13116 3996 13176 5026
rect 13236 3934 13296 4966
rect 13356 4872 13422 4962
rect 13356 4808 13357 4872
rect 13421 4808 13422 4872
rect 13356 4792 13422 4808
rect 13356 4728 13357 4792
rect 13421 4728 13422 4792
rect 13356 4712 13422 4728
rect 13356 4648 13357 4712
rect 13421 4648 13422 4712
rect 13356 4632 13422 4648
rect 13356 4568 13357 4632
rect 13421 4568 13422 4632
rect 13356 4552 13422 4568
rect 13356 4488 13357 4552
rect 13421 4488 13422 4552
rect 13356 4472 13422 4488
rect 13356 4408 13357 4472
rect 13421 4408 13422 4472
rect 13356 4392 13422 4408
rect 13356 4328 13357 4392
rect 13421 4328 13422 4392
rect 13356 4312 13422 4328
rect 13356 4248 13357 4312
rect 13421 4248 13422 4312
rect 13356 4232 13422 4248
rect 13356 4168 13357 4232
rect 13421 4168 13422 4232
rect 13356 4152 13422 4168
rect 13356 4088 13357 4152
rect 13421 4088 13422 4152
rect 13356 3934 13422 4088
rect 13482 3996 13542 5026
rect 13602 3934 13662 4966
rect 13722 3996 13782 5026
rect 13842 3934 13902 4966
rect 13962 4872 14028 4962
rect 13962 4808 13963 4872
rect 14027 4808 14028 4872
rect 13962 4792 14028 4808
rect 13962 4728 13963 4792
rect 14027 4728 14028 4792
rect 13962 4712 14028 4728
rect 13962 4648 13963 4712
rect 14027 4648 14028 4712
rect 13962 4632 14028 4648
rect 13962 4568 13963 4632
rect 14027 4568 14028 4632
rect 13962 4552 14028 4568
rect 13962 4488 13963 4552
rect 14027 4488 14028 4552
rect 13962 4472 14028 4488
rect 13962 4408 13963 4472
rect 14027 4408 14028 4472
rect 13962 4392 14028 4408
rect 13962 4328 13963 4392
rect 14027 4328 14028 4392
rect 13962 4312 14028 4328
rect 13962 4248 13963 4312
rect 14027 4248 14028 4312
rect 13962 4232 14028 4248
rect 13962 4168 13963 4232
rect 14027 4168 14028 4232
rect 13962 4152 14028 4168
rect 13962 4088 13963 4152
rect 14027 4088 14028 4152
rect 13962 3934 14028 4088
rect 14088 3996 14148 5026
rect 14208 3934 14268 4966
rect 14328 3996 14388 5026
rect 14448 3934 14508 4966
rect 14568 4872 14634 4962
rect 14568 4808 14569 4872
rect 14633 4808 14634 4872
rect 14568 4792 14634 4808
rect 14568 4728 14569 4792
rect 14633 4728 14634 4792
rect 14568 4712 14634 4728
rect 14568 4648 14569 4712
rect 14633 4648 14634 4712
rect 14568 4632 14634 4648
rect 14568 4568 14569 4632
rect 14633 4568 14634 4632
rect 14568 4552 14634 4568
rect 14568 4488 14569 4552
rect 14633 4488 14634 4552
rect 14568 4472 14634 4488
rect 14568 4408 14569 4472
rect 14633 4408 14634 4472
rect 14568 4392 14634 4408
rect 14568 4328 14569 4392
rect 14633 4328 14634 4392
rect 14568 4312 14634 4328
rect 14568 4248 14569 4312
rect 14633 4248 14634 4312
rect 14568 4232 14634 4248
rect 14568 4168 14569 4232
rect 14633 4168 14634 4232
rect 14568 4152 14634 4168
rect 14568 4088 14569 4152
rect 14633 4088 14634 4152
rect 14568 3934 14634 4088
rect 14694 3996 14754 5026
rect 14814 3934 14874 4966
rect 14934 3996 14994 5026
rect 15054 3934 15114 4966
rect 15174 4872 15240 4962
rect 15174 4808 15175 4872
rect 15239 4808 15240 4872
rect 15174 4792 15240 4808
rect 15174 4728 15175 4792
rect 15239 4728 15240 4792
rect 15174 4712 15240 4728
rect 15174 4648 15175 4712
rect 15239 4648 15240 4712
rect 15174 4632 15240 4648
rect 15174 4568 15175 4632
rect 15239 4568 15240 4632
rect 15174 4552 15240 4568
rect 15174 4488 15175 4552
rect 15239 4488 15240 4552
rect 15174 4472 15240 4488
rect 15174 4408 15175 4472
rect 15239 4408 15240 4472
rect 15174 4392 15240 4408
rect 15174 4328 15175 4392
rect 15239 4328 15240 4392
rect 15174 4312 15240 4328
rect 15174 4248 15175 4312
rect 15239 4248 15240 4312
rect 15174 4232 15240 4248
rect 15174 4168 15175 4232
rect 15239 4168 15240 4232
rect 15174 4152 15240 4168
rect 15174 4088 15175 4152
rect 15239 4088 15240 4152
rect 15174 3934 15240 4088
rect 15300 3996 15360 5026
rect 15420 3934 15480 4966
rect 15540 3996 15600 5026
rect 15660 3934 15720 4966
rect 15780 4872 15846 4962
rect 15780 4808 15781 4872
rect 15845 4808 15846 4872
rect 15780 4792 15846 4808
rect 15780 4728 15781 4792
rect 15845 4728 15846 4792
rect 15780 4712 15846 4728
rect 15780 4648 15781 4712
rect 15845 4648 15846 4712
rect 15780 4632 15846 4648
rect 15780 4568 15781 4632
rect 15845 4568 15846 4632
rect 15780 4552 15846 4568
rect 15780 4488 15781 4552
rect 15845 4488 15846 4552
rect 15780 4472 15846 4488
rect 15780 4408 15781 4472
rect 15845 4408 15846 4472
rect 15780 4392 15846 4408
rect 15780 4328 15781 4392
rect 15845 4328 15846 4392
rect 15780 4312 15846 4328
rect 15780 4248 15781 4312
rect 15845 4248 15846 4312
rect 15780 4232 15846 4248
rect 15780 4168 15781 4232
rect 15845 4168 15846 4232
rect 15780 4152 15846 4168
rect 15780 4088 15781 4152
rect 15845 4088 15846 4152
rect 15780 3934 15846 4088
rect 15906 3996 15966 5026
rect 16026 3934 16086 4966
rect 16146 3996 16206 5026
rect 16266 3934 16326 4966
rect 16386 4872 16452 4962
rect 16386 4808 16387 4872
rect 16451 4808 16452 4872
rect 16386 4792 16452 4808
rect 16386 4728 16387 4792
rect 16451 4728 16452 4792
rect 16386 4712 16452 4728
rect 16386 4648 16387 4712
rect 16451 4648 16452 4712
rect 16386 4632 16452 4648
rect 16386 4568 16387 4632
rect 16451 4568 16452 4632
rect 16386 4552 16452 4568
rect 16386 4488 16387 4552
rect 16451 4488 16452 4552
rect 16386 4472 16452 4488
rect 16386 4408 16387 4472
rect 16451 4408 16452 4472
rect 16386 4392 16452 4408
rect 16386 4328 16387 4392
rect 16451 4328 16452 4392
rect 16386 4312 16452 4328
rect 16386 4248 16387 4312
rect 16451 4248 16452 4312
rect 16386 4232 16452 4248
rect 16386 4168 16387 4232
rect 16451 4168 16452 4232
rect 16386 4152 16452 4168
rect 16386 4088 16387 4152
rect 16451 4088 16452 4152
rect 16386 3934 16452 4088
rect 16512 3996 16572 5026
rect 16632 3934 16692 4966
rect 16752 3996 16812 5026
rect 16872 3934 16932 4966
rect 16992 4872 17058 4962
rect 16992 4808 16993 4872
rect 17057 4808 17058 4872
rect 16992 4792 17058 4808
rect 16992 4728 16993 4792
rect 17057 4728 17058 4792
rect 16992 4712 17058 4728
rect 16992 4648 16993 4712
rect 17057 4648 17058 4712
rect 16992 4632 17058 4648
rect 16992 4568 16993 4632
rect 17057 4568 17058 4632
rect 16992 4552 17058 4568
rect 16992 4488 16993 4552
rect 17057 4488 17058 4552
rect 16992 4472 17058 4488
rect 16992 4408 16993 4472
rect 17057 4408 17058 4472
rect 16992 4392 17058 4408
rect 16992 4328 16993 4392
rect 17057 4328 17058 4392
rect 16992 4312 17058 4328
rect 16992 4248 16993 4312
rect 17057 4248 17058 4312
rect 16992 4232 17058 4248
rect 16992 4168 16993 4232
rect 17057 4168 17058 4232
rect 16992 4152 17058 4168
rect 16992 4088 16993 4152
rect 17057 4088 17058 4152
rect 16992 3934 17058 4088
rect 17118 3996 17178 5026
rect 17238 3934 17298 4966
rect 17358 3996 17418 5026
rect 17478 3934 17538 4966
rect 17598 4872 17664 4962
rect 17598 4808 17599 4872
rect 17663 4808 17664 4872
rect 17598 4792 17664 4808
rect 17598 4728 17599 4792
rect 17663 4728 17664 4792
rect 17598 4712 17664 4728
rect 17598 4648 17599 4712
rect 17663 4648 17664 4712
rect 17598 4632 17664 4648
rect 17598 4568 17599 4632
rect 17663 4568 17664 4632
rect 17598 4552 17664 4568
rect 17598 4488 17599 4552
rect 17663 4488 17664 4552
rect 17598 4472 17664 4488
rect 17598 4408 17599 4472
rect 17663 4408 17664 4472
rect 17598 4392 17664 4408
rect 17598 4328 17599 4392
rect 17663 4328 17664 4392
rect 17598 4312 17664 4328
rect 17598 4248 17599 4312
rect 17663 4248 17664 4312
rect 17598 4232 17664 4248
rect 17598 4168 17599 4232
rect 17663 4168 17664 4232
rect 17598 4152 17664 4168
rect 17598 4088 17599 4152
rect 17663 4088 17664 4152
rect 17598 3934 17664 4088
rect 17724 3996 17784 5026
rect 17844 3934 17904 4966
rect 17964 3996 18024 5026
rect 18084 3934 18144 4966
rect 18204 4872 18270 4962
rect 18204 4808 18205 4872
rect 18269 4808 18270 4872
rect 18204 4792 18270 4808
rect 18204 4728 18205 4792
rect 18269 4728 18270 4792
rect 18204 4712 18270 4728
rect 18204 4648 18205 4712
rect 18269 4648 18270 4712
rect 18204 4632 18270 4648
rect 18204 4568 18205 4632
rect 18269 4568 18270 4632
rect 18204 4552 18270 4568
rect 18204 4488 18205 4552
rect 18269 4488 18270 4552
rect 18204 4472 18270 4488
rect 18204 4408 18205 4472
rect 18269 4408 18270 4472
rect 18204 4392 18270 4408
rect 18204 4328 18205 4392
rect 18269 4328 18270 4392
rect 18204 4312 18270 4328
rect 18204 4248 18205 4312
rect 18269 4248 18270 4312
rect 18204 4232 18270 4248
rect 18204 4168 18205 4232
rect 18269 4168 18270 4232
rect 18204 4152 18270 4168
rect 18204 4088 18205 4152
rect 18269 4088 18270 4152
rect 18204 3934 18270 4088
rect 18330 3996 18390 5026
rect 18450 3934 18510 4966
rect 18570 3996 18630 5026
rect 18690 3934 18750 4966
rect 18810 4872 18876 4962
rect 18810 4808 18811 4872
rect 18875 4808 18876 4872
rect 18810 4792 18876 4808
rect 18810 4728 18811 4792
rect 18875 4728 18876 4792
rect 18810 4712 18876 4728
rect 18810 4648 18811 4712
rect 18875 4648 18876 4712
rect 18810 4632 18876 4648
rect 18810 4568 18811 4632
rect 18875 4568 18876 4632
rect 18810 4552 18876 4568
rect 18810 4488 18811 4552
rect 18875 4488 18876 4552
rect 18810 4472 18876 4488
rect 18810 4408 18811 4472
rect 18875 4408 18876 4472
rect 18810 4392 18876 4408
rect 18810 4328 18811 4392
rect 18875 4328 18876 4392
rect 18810 4312 18876 4328
rect 18810 4248 18811 4312
rect 18875 4248 18876 4312
rect 18810 4232 18876 4248
rect 18810 4168 18811 4232
rect 18875 4168 18876 4232
rect 18810 4152 18876 4168
rect 18810 4088 18811 4152
rect 18875 4088 18876 4152
rect 18810 3934 18876 4088
rect 18936 3996 18996 5026
rect 19056 3934 19116 4966
rect 19176 3996 19236 5026
rect 19296 3934 19356 4966
rect 19416 4872 19482 4962
rect 19416 4808 19417 4872
rect 19481 4808 19482 4872
rect 19416 4792 19482 4808
rect 19416 4728 19417 4792
rect 19481 4728 19482 4792
rect 19416 4712 19482 4728
rect 19416 4648 19417 4712
rect 19481 4648 19482 4712
rect 19416 4632 19482 4648
rect 19416 4568 19417 4632
rect 19481 4568 19482 4632
rect 19416 4552 19482 4568
rect 19416 4488 19417 4552
rect 19481 4488 19482 4552
rect 19416 4472 19482 4488
rect 19416 4408 19417 4472
rect 19481 4408 19482 4472
rect 19416 4392 19482 4408
rect 19416 4328 19417 4392
rect 19481 4328 19482 4392
rect 19416 4312 19482 4328
rect 19416 4248 19417 4312
rect 19481 4248 19482 4312
rect 19416 4232 19482 4248
rect 19416 4168 19417 4232
rect 19481 4168 19482 4232
rect 19416 4152 19482 4168
rect 19416 4088 19417 4152
rect 19481 4088 19482 4152
rect 19416 3934 19482 4088
rect 19542 3996 19602 5026
rect 19662 3934 19722 4966
rect 19782 3996 19842 5026
rect 19902 3934 19962 4966
rect 20022 4872 20088 4962
rect 20022 4808 20023 4872
rect 20087 4808 20088 4872
rect 20022 4792 20088 4808
rect 20022 4728 20023 4792
rect 20087 4728 20088 4792
rect 20022 4712 20088 4728
rect 20022 4648 20023 4712
rect 20087 4648 20088 4712
rect 20022 4632 20088 4648
rect 20022 4568 20023 4632
rect 20087 4568 20088 4632
rect 20022 4552 20088 4568
rect 20022 4488 20023 4552
rect 20087 4488 20088 4552
rect 20022 4472 20088 4488
rect 20022 4408 20023 4472
rect 20087 4408 20088 4472
rect 20022 4392 20088 4408
rect 20022 4328 20023 4392
rect 20087 4328 20088 4392
rect 20022 4312 20088 4328
rect 20022 4248 20023 4312
rect 20087 4248 20088 4312
rect 20022 4232 20088 4248
rect 20022 4168 20023 4232
rect 20087 4168 20088 4232
rect 20022 4152 20088 4168
rect 20022 4088 20023 4152
rect 20087 4088 20088 4152
rect 20022 3934 20088 4088
rect 10326 3932 20088 3934
rect 10326 3868 10430 3932
rect 10494 3868 10510 3932
rect 10574 3868 10590 3932
rect 10654 3868 10670 3932
rect 10734 3868 10750 3932
rect 10814 3868 10830 3932
rect 10894 3868 11036 3932
rect 11100 3868 11116 3932
rect 11180 3868 11196 3932
rect 11260 3868 11276 3932
rect 11340 3868 11356 3932
rect 11420 3868 11436 3932
rect 11500 3868 11642 3932
rect 11706 3868 11722 3932
rect 11786 3868 11802 3932
rect 11866 3868 11882 3932
rect 11946 3868 11962 3932
rect 12026 3868 12042 3932
rect 12106 3868 12248 3932
rect 12312 3868 12328 3932
rect 12392 3868 12408 3932
rect 12472 3868 12488 3932
rect 12552 3868 12568 3932
rect 12632 3868 12648 3932
rect 12712 3868 12854 3932
rect 12918 3868 12934 3932
rect 12998 3868 13014 3932
rect 13078 3868 13094 3932
rect 13158 3868 13174 3932
rect 13238 3868 13254 3932
rect 13318 3868 13460 3932
rect 13524 3868 13540 3932
rect 13604 3868 13620 3932
rect 13684 3868 13700 3932
rect 13764 3868 13780 3932
rect 13844 3868 13860 3932
rect 13924 3868 14066 3932
rect 14130 3868 14146 3932
rect 14210 3868 14226 3932
rect 14290 3868 14306 3932
rect 14370 3868 14386 3932
rect 14450 3868 14466 3932
rect 14530 3868 14672 3932
rect 14736 3868 14752 3932
rect 14816 3868 14832 3932
rect 14896 3868 14912 3932
rect 14976 3868 14992 3932
rect 15056 3868 15072 3932
rect 15136 3868 15278 3932
rect 15342 3868 15358 3932
rect 15422 3868 15438 3932
rect 15502 3868 15518 3932
rect 15582 3868 15598 3932
rect 15662 3868 15678 3932
rect 15742 3868 15884 3932
rect 15948 3868 15964 3932
rect 16028 3868 16044 3932
rect 16108 3868 16124 3932
rect 16188 3868 16204 3932
rect 16268 3868 16284 3932
rect 16348 3868 16490 3932
rect 16554 3868 16570 3932
rect 16634 3868 16650 3932
rect 16714 3868 16730 3932
rect 16794 3868 16810 3932
rect 16874 3868 16890 3932
rect 16954 3868 17096 3932
rect 17160 3868 17176 3932
rect 17240 3868 17256 3932
rect 17320 3868 17336 3932
rect 17400 3868 17416 3932
rect 17480 3868 17496 3932
rect 17560 3868 17702 3932
rect 17766 3868 17782 3932
rect 17846 3868 17862 3932
rect 17926 3868 17942 3932
rect 18006 3868 18022 3932
rect 18086 3868 18102 3932
rect 18166 3868 18308 3932
rect 18372 3868 18388 3932
rect 18452 3868 18468 3932
rect 18532 3868 18548 3932
rect 18612 3868 18628 3932
rect 18692 3868 18708 3932
rect 18772 3868 18914 3932
rect 18978 3868 18994 3932
rect 19058 3868 19074 3932
rect 19138 3868 19154 3932
rect 19218 3868 19234 3932
rect 19298 3868 19314 3932
rect 19378 3868 19520 3932
rect 19584 3868 19600 3932
rect 19664 3868 19680 3932
rect 19744 3868 19760 3932
rect 19824 3868 19840 3932
rect 19904 3868 19920 3932
rect 19984 3868 20088 3932
rect 10326 3866 20088 3868
rect 10326 3712 10392 3866
rect 10326 3648 10327 3712
rect 10391 3648 10392 3712
rect 10326 3632 10392 3648
rect 10326 3568 10327 3632
rect 10391 3568 10392 3632
rect 10326 3552 10392 3568
rect 10326 3488 10327 3552
rect 10391 3488 10392 3552
rect 10326 3472 10392 3488
rect 10326 3408 10327 3472
rect 10391 3408 10392 3472
rect 10326 3392 10392 3408
rect 10326 3328 10327 3392
rect 10391 3328 10392 3392
rect 10326 3312 10392 3328
rect 10326 3248 10327 3312
rect 10391 3248 10392 3312
rect 10326 3232 10392 3248
rect 10326 3168 10327 3232
rect 10391 3168 10392 3232
rect 10326 3152 10392 3168
rect 10326 3088 10327 3152
rect 10391 3088 10392 3152
rect 10326 3072 10392 3088
rect 10326 3008 10327 3072
rect 10391 3008 10392 3072
rect 10326 2992 10392 3008
rect 10326 2928 10327 2992
rect 10391 2928 10392 2992
rect 10326 2838 10392 2928
rect 10452 2834 10512 3866
rect 10572 2774 10632 3804
rect 10692 2834 10752 3866
rect 10812 2774 10872 3804
rect 10932 3712 10998 3866
rect 10932 3648 10933 3712
rect 10997 3648 10998 3712
rect 10932 3632 10998 3648
rect 10932 3568 10933 3632
rect 10997 3568 10998 3632
rect 10932 3552 10998 3568
rect 10932 3488 10933 3552
rect 10997 3488 10998 3552
rect 10932 3472 10998 3488
rect 10932 3408 10933 3472
rect 10997 3408 10998 3472
rect 10932 3392 10998 3408
rect 10932 3328 10933 3392
rect 10997 3328 10998 3392
rect 10932 3312 10998 3328
rect 10932 3248 10933 3312
rect 10997 3248 10998 3312
rect 10932 3232 10998 3248
rect 10932 3168 10933 3232
rect 10997 3168 10998 3232
rect 10932 3152 10998 3168
rect 10932 3088 10933 3152
rect 10997 3088 10998 3152
rect 10932 3072 10998 3088
rect 10932 3008 10933 3072
rect 10997 3008 10998 3072
rect 10932 2992 10998 3008
rect 10932 2928 10933 2992
rect 10997 2928 10998 2992
rect 10932 2838 10998 2928
rect 11058 2834 11118 3866
rect 11178 2774 11238 3804
rect 11298 2834 11358 3866
rect 11418 2774 11478 3804
rect 11538 3712 11604 3866
rect 11538 3648 11539 3712
rect 11603 3648 11604 3712
rect 11538 3632 11604 3648
rect 11538 3568 11539 3632
rect 11603 3568 11604 3632
rect 11538 3552 11604 3568
rect 11538 3488 11539 3552
rect 11603 3488 11604 3552
rect 11538 3472 11604 3488
rect 11538 3408 11539 3472
rect 11603 3408 11604 3472
rect 11538 3392 11604 3408
rect 11538 3328 11539 3392
rect 11603 3328 11604 3392
rect 11538 3312 11604 3328
rect 11538 3248 11539 3312
rect 11603 3248 11604 3312
rect 11538 3232 11604 3248
rect 11538 3168 11539 3232
rect 11603 3168 11604 3232
rect 11538 3152 11604 3168
rect 11538 3088 11539 3152
rect 11603 3088 11604 3152
rect 11538 3072 11604 3088
rect 11538 3008 11539 3072
rect 11603 3008 11604 3072
rect 11538 2992 11604 3008
rect 11538 2928 11539 2992
rect 11603 2928 11604 2992
rect 11538 2838 11604 2928
rect 11664 2834 11724 3866
rect 11784 2774 11844 3804
rect 11904 2834 11964 3866
rect 12024 2774 12084 3804
rect 12144 3712 12210 3866
rect 12144 3648 12145 3712
rect 12209 3648 12210 3712
rect 12144 3632 12210 3648
rect 12144 3568 12145 3632
rect 12209 3568 12210 3632
rect 12144 3552 12210 3568
rect 12144 3488 12145 3552
rect 12209 3488 12210 3552
rect 12144 3472 12210 3488
rect 12144 3408 12145 3472
rect 12209 3408 12210 3472
rect 12144 3392 12210 3408
rect 12144 3328 12145 3392
rect 12209 3328 12210 3392
rect 12144 3312 12210 3328
rect 12144 3248 12145 3312
rect 12209 3248 12210 3312
rect 12144 3232 12210 3248
rect 12144 3168 12145 3232
rect 12209 3168 12210 3232
rect 12144 3152 12210 3168
rect 12144 3088 12145 3152
rect 12209 3088 12210 3152
rect 12144 3072 12210 3088
rect 12144 3008 12145 3072
rect 12209 3008 12210 3072
rect 12144 2992 12210 3008
rect 12144 2928 12145 2992
rect 12209 2928 12210 2992
rect 12144 2838 12210 2928
rect 12270 2834 12330 3866
rect 12390 2774 12450 3804
rect 12510 2834 12570 3866
rect 12630 2774 12690 3804
rect 12750 3712 12816 3866
rect 12750 3648 12751 3712
rect 12815 3648 12816 3712
rect 12750 3632 12816 3648
rect 12750 3568 12751 3632
rect 12815 3568 12816 3632
rect 12750 3552 12816 3568
rect 12750 3488 12751 3552
rect 12815 3488 12816 3552
rect 12750 3472 12816 3488
rect 12750 3408 12751 3472
rect 12815 3408 12816 3472
rect 12750 3392 12816 3408
rect 12750 3328 12751 3392
rect 12815 3328 12816 3392
rect 12750 3312 12816 3328
rect 12750 3248 12751 3312
rect 12815 3248 12816 3312
rect 12750 3232 12816 3248
rect 12750 3168 12751 3232
rect 12815 3168 12816 3232
rect 12750 3152 12816 3168
rect 12750 3088 12751 3152
rect 12815 3088 12816 3152
rect 12750 3072 12816 3088
rect 12750 3008 12751 3072
rect 12815 3008 12816 3072
rect 12750 2992 12816 3008
rect 12750 2928 12751 2992
rect 12815 2928 12816 2992
rect 12750 2838 12816 2928
rect 12876 2834 12936 3866
rect 12996 2774 13056 3804
rect 13116 2834 13176 3866
rect 13236 2774 13296 3804
rect 13356 3712 13422 3866
rect 13356 3648 13357 3712
rect 13421 3648 13422 3712
rect 13356 3632 13422 3648
rect 13356 3568 13357 3632
rect 13421 3568 13422 3632
rect 13356 3552 13422 3568
rect 13356 3488 13357 3552
rect 13421 3488 13422 3552
rect 13356 3472 13422 3488
rect 13356 3408 13357 3472
rect 13421 3408 13422 3472
rect 13356 3392 13422 3408
rect 13356 3328 13357 3392
rect 13421 3328 13422 3392
rect 13356 3312 13422 3328
rect 13356 3248 13357 3312
rect 13421 3248 13422 3312
rect 13356 3232 13422 3248
rect 13356 3168 13357 3232
rect 13421 3168 13422 3232
rect 13356 3152 13422 3168
rect 13356 3088 13357 3152
rect 13421 3088 13422 3152
rect 13356 3072 13422 3088
rect 13356 3008 13357 3072
rect 13421 3008 13422 3072
rect 13356 2992 13422 3008
rect 13356 2928 13357 2992
rect 13421 2928 13422 2992
rect 13356 2838 13422 2928
rect 13482 2834 13542 3866
rect 13602 2774 13662 3804
rect 13722 2834 13782 3866
rect 13842 2774 13902 3804
rect 13962 3712 14028 3866
rect 13962 3648 13963 3712
rect 14027 3648 14028 3712
rect 13962 3632 14028 3648
rect 13962 3568 13963 3632
rect 14027 3568 14028 3632
rect 13962 3552 14028 3568
rect 13962 3488 13963 3552
rect 14027 3488 14028 3552
rect 13962 3472 14028 3488
rect 13962 3408 13963 3472
rect 14027 3408 14028 3472
rect 13962 3392 14028 3408
rect 13962 3328 13963 3392
rect 14027 3328 14028 3392
rect 13962 3312 14028 3328
rect 13962 3248 13963 3312
rect 14027 3248 14028 3312
rect 13962 3232 14028 3248
rect 13962 3168 13963 3232
rect 14027 3168 14028 3232
rect 13962 3152 14028 3168
rect 13962 3088 13963 3152
rect 14027 3088 14028 3152
rect 13962 3072 14028 3088
rect 13962 3008 13963 3072
rect 14027 3008 14028 3072
rect 13962 2992 14028 3008
rect 13962 2928 13963 2992
rect 14027 2928 14028 2992
rect 13962 2838 14028 2928
rect 14088 2834 14148 3866
rect 14208 2774 14268 3804
rect 14328 2834 14388 3866
rect 14448 2774 14508 3804
rect 14568 3712 14634 3866
rect 14568 3648 14569 3712
rect 14633 3648 14634 3712
rect 14568 3632 14634 3648
rect 14568 3568 14569 3632
rect 14633 3568 14634 3632
rect 14568 3552 14634 3568
rect 14568 3488 14569 3552
rect 14633 3488 14634 3552
rect 14568 3472 14634 3488
rect 14568 3408 14569 3472
rect 14633 3408 14634 3472
rect 14568 3392 14634 3408
rect 14568 3328 14569 3392
rect 14633 3328 14634 3392
rect 14568 3312 14634 3328
rect 14568 3248 14569 3312
rect 14633 3248 14634 3312
rect 14568 3232 14634 3248
rect 14568 3168 14569 3232
rect 14633 3168 14634 3232
rect 14568 3152 14634 3168
rect 14568 3088 14569 3152
rect 14633 3088 14634 3152
rect 14568 3072 14634 3088
rect 14568 3008 14569 3072
rect 14633 3008 14634 3072
rect 14568 2992 14634 3008
rect 14568 2928 14569 2992
rect 14633 2928 14634 2992
rect 14568 2838 14634 2928
rect 14694 2834 14754 3866
rect 14814 2774 14874 3804
rect 14934 2834 14994 3866
rect 15054 2774 15114 3804
rect 15174 3712 15240 3866
rect 15174 3648 15175 3712
rect 15239 3648 15240 3712
rect 15174 3632 15240 3648
rect 15174 3568 15175 3632
rect 15239 3568 15240 3632
rect 15174 3552 15240 3568
rect 15174 3488 15175 3552
rect 15239 3488 15240 3552
rect 15174 3472 15240 3488
rect 15174 3408 15175 3472
rect 15239 3408 15240 3472
rect 15174 3392 15240 3408
rect 15174 3328 15175 3392
rect 15239 3328 15240 3392
rect 15174 3312 15240 3328
rect 15174 3248 15175 3312
rect 15239 3248 15240 3312
rect 15174 3232 15240 3248
rect 15174 3168 15175 3232
rect 15239 3168 15240 3232
rect 15174 3152 15240 3168
rect 15174 3088 15175 3152
rect 15239 3088 15240 3152
rect 15174 3072 15240 3088
rect 15174 3008 15175 3072
rect 15239 3008 15240 3072
rect 15174 2992 15240 3008
rect 15174 2928 15175 2992
rect 15239 2928 15240 2992
rect 15174 2838 15240 2928
rect 15300 2834 15360 3866
rect 15420 2774 15480 3804
rect 15540 2834 15600 3866
rect 15660 2774 15720 3804
rect 15780 3712 15846 3866
rect 15780 3648 15781 3712
rect 15845 3648 15846 3712
rect 15780 3632 15846 3648
rect 15780 3568 15781 3632
rect 15845 3568 15846 3632
rect 15780 3552 15846 3568
rect 15780 3488 15781 3552
rect 15845 3488 15846 3552
rect 15780 3472 15846 3488
rect 15780 3408 15781 3472
rect 15845 3408 15846 3472
rect 15780 3392 15846 3408
rect 15780 3328 15781 3392
rect 15845 3328 15846 3392
rect 15780 3312 15846 3328
rect 15780 3248 15781 3312
rect 15845 3248 15846 3312
rect 15780 3232 15846 3248
rect 15780 3168 15781 3232
rect 15845 3168 15846 3232
rect 15780 3152 15846 3168
rect 15780 3088 15781 3152
rect 15845 3088 15846 3152
rect 15780 3072 15846 3088
rect 15780 3008 15781 3072
rect 15845 3008 15846 3072
rect 15780 2992 15846 3008
rect 15780 2928 15781 2992
rect 15845 2928 15846 2992
rect 15780 2838 15846 2928
rect 15906 2834 15966 3866
rect 16026 2774 16086 3804
rect 16146 2834 16206 3866
rect 16266 2774 16326 3804
rect 16386 3712 16452 3866
rect 16386 3648 16387 3712
rect 16451 3648 16452 3712
rect 16386 3632 16452 3648
rect 16386 3568 16387 3632
rect 16451 3568 16452 3632
rect 16386 3552 16452 3568
rect 16386 3488 16387 3552
rect 16451 3488 16452 3552
rect 16386 3472 16452 3488
rect 16386 3408 16387 3472
rect 16451 3408 16452 3472
rect 16386 3392 16452 3408
rect 16386 3328 16387 3392
rect 16451 3328 16452 3392
rect 16386 3312 16452 3328
rect 16386 3248 16387 3312
rect 16451 3248 16452 3312
rect 16386 3232 16452 3248
rect 16386 3168 16387 3232
rect 16451 3168 16452 3232
rect 16386 3152 16452 3168
rect 16386 3088 16387 3152
rect 16451 3088 16452 3152
rect 16386 3072 16452 3088
rect 16386 3008 16387 3072
rect 16451 3008 16452 3072
rect 16386 2992 16452 3008
rect 16386 2928 16387 2992
rect 16451 2928 16452 2992
rect 16386 2838 16452 2928
rect 16512 2834 16572 3866
rect 16632 2774 16692 3804
rect 16752 2834 16812 3866
rect 16872 2774 16932 3804
rect 16992 3712 17058 3866
rect 16992 3648 16993 3712
rect 17057 3648 17058 3712
rect 16992 3632 17058 3648
rect 16992 3568 16993 3632
rect 17057 3568 17058 3632
rect 16992 3552 17058 3568
rect 16992 3488 16993 3552
rect 17057 3488 17058 3552
rect 16992 3472 17058 3488
rect 16992 3408 16993 3472
rect 17057 3408 17058 3472
rect 16992 3392 17058 3408
rect 16992 3328 16993 3392
rect 17057 3328 17058 3392
rect 16992 3312 17058 3328
rect 16992 3248 16993 3312
rect 17057 3248 17058 3312
rect 16992 3232 17058 3248
rect 16992 3168 16993 3232
rect 17057 3168 17058 3232
rect 16992 3152 17058 3168
rect 16992 3088 16993 3152
rect 17057 3088 17058 3152
rect 16992 3072 17058 3088
rect 16992 3008 16993 3072
rect 17057 3008 17058 3072
rect 16992 2992 17058 3008
rect 16992 2928 16993 2992
rect 17057 2928 17058 2992
rect 16992 2838 17058 2928
rect 17118 2834 17178 3866
rect 17238 2774 17298 3804
rect 17358 2834 17418 3866
rect 17478 2774 17538 3804
rect 17598 3712 17664 3866
rect 17598 3648 17599 3712
rect 17663 3648 17664 3712
rect 17598 3632 17664 3648
rect 17598 3568 17599 3632
rect 17663 3568 17664 3632
rect 17598 3552 17664 3568
rect 17598 3488 17599 3552
rect 17663 3488 17664 3552
rect 17598 3472 17664 3488
rect 17598 3408 17599 3472
rect 17663 3408 17664 3472
rect 17598 3392 17664 3408
rect 17598 3328 17599 3392
rect 17663 3328 17664 3392
rect 17598 3312 17664 3328
rect 17598 3248 17599 3312
rect 17663 3248 17664 3312
rect 17598 3232 17664 3248
rect 17598 3168 17599 3232
rect 17663 3168 17664 3232
rect 17598 3152 17664 3168
rect 17598 3088 17599 3152
rect 17663 3088 17664 3152
rect 17598 3072 17664 3088
rect 17598 3008 17599 3072
rect 17663 3008 17664 3072
rect 17598 2992 17664 3008
rect 17598 2928 17599 2992
rect 17663 2928 17664 2992
rect 17598 2838 17664 2928
rect 17724 2834 17784 3866
rect 17844 2774 17904 3804
rect 17964 2834 18024 3866
rect 18084 2774 18144 3804
rect 18204 3712 18270 3866
rect 18204 3648 18205 3712
rect 18269 3648 18270 3712
rect 18204 3632 18270 3648
rect 18204 3568 18205 3632
rect 18269 3568 18270 3632
rect 18204 3552 18270 3568
rect 18204 3488 18205 3552
rect 18269 3488 18270 3552
rect 18204 3472 18270 3488
rect 18204 3408 18205 3472
rect 18269 3408 18270 3472
rect 18204 3392 18270 3408
rect 18204 3328 18205 3392
rect 18269 3328 18270 3392
rect 18204 3312 18270 3328
rect 18204 3248 18205 3312
rect 18269 3248 18270 3312
rect 18204 3232 18270 3248
rect 18204 3168 18205 3232
rect 18269 3168 18270 3232
rect 18204 3152 18270 3168
rect 18204 3088 18205 3152
rect 18269 3088 18270 3152
rect 18204 3072 18270 3088
rect 18204 3008 18205 3072
rect 18269 3008 18270 3072
rect 18204 2992 18270 3008
rect 18204 2928 18205 2992
rect 18269 2928 18270 2992
rect 18204 2838 18270 2928
rect 18330 2834 18390 3866
rect 18450 2774 18510 3804
rect 18570 2834 18630 3866
rect 18690 2774 18750 3804
rect 18810 3712 18876 3866
rect 18810 3648 18811 3712
rect 18875 3648 18876 3712
rect 18810 3632 18876 3648
rect 18810 3568 18811 3632
rect 18875 3568 18876 3632
rect 18810 3552 18876 3568
rect 18810 3488 18811 3552
rect 18875 3488 18876 3552
rect 18810 3472 18876 3488
rect 18810 3408 18811 3472
rect 18875 3408 18876 3472
rect 18810 3392 18876 3408
rect 18810 3328 18811 3392
rect 18875 3328 18876 3392
rect 18810 3312 18876 3328
rect 18810 3248 18811 3312
rect 18875 3248 18876 3312
rect 18810 3232 18876 3248
rect 18810 3168 18811 3232
rect 18875 3168 18876 3232
rect 18810 3152 18876 3168
rect 18810 3088 18811 3152
rect 18875 3088 18876 3152
rect 18810 3072 18876 3088
rect 18810 3008 18811 3072
rect 18875 3008 18876 3072
rect 18810 2992 18876 3008
rect 18810 2928 18811 2992
rect 18875 2928 18876 2992
rect 18810 2838 18876 2928
rect 18936 2834 18996 3866
rect 19056 2774 19116 3804
rect 19176 2834 19236 3866
rect 19296 2774 19356 3804
rect 19416 3712 19482 3866
rect 19416 3648 19417 3712
rect 19481 3648 19482 3712
rect 19416 3632 19482 3648
rect 19416 3568 19417 3632
rect 19481 3568 19482 3632
rect 19416 3552 19482 3568
rect 19416 3488 19417 3552
rect 19481 3488 19482 3552
rect 19416 3472 19482 3488
rect 19416 3408 19417 3472
rect 19481 3408 19482 3472
rect 19416 3392 19482 3408
rect 19416 3328 19417 3392
rect 19481 3328 19482 3392
rect 19416 3312 19482 3328
rect 19416 3248 19417 3312
rect 19481 3248 19482 3312
rect 19416 3232 19482 3248
rect 19416 3168 19417 3232
rect 19481 3168 19482 3232
rect 19416 3152 19482 3168
rect 19416 3088 19417 3152
rect 19481 3088 19482 3152
rect 19416 3072 19482 3088
rect 19416 3008 19417 3072
rect 19481 3008 19482 3072
rect 19416 2992 19482 3008
rect 19416 2928 19417 2992
rect 19481 2928 19482 2992
rect 19416 2838 19482 2928
rect 19542 2834 19602 3866
rect 19662 2774 19722 3804
rect 19782 2834 19842 3866
rect 19902 2774 19962 3804
rect 20022 3712 20088 3866
rect 20022 3648 20023 3712
rect 20087 3648 20088 3712
rect 20022 3632 20088 3648
rect 20022 3568 20023 3632
rect 20087 3568 20088 3632
rect 20022 3552 20088 3568
rect 20022 3488 20023 3552
rect 20087 3488 20088 3552
rect 20022 3472 20088 3488
rect 20022 3408 20023 3472
rect 20087 3408 20088 3472
rect 20022 3392 20088 3408
rect 20022 3328 20023 3392
rect 20087 3328 20088 3392
rect 20022 3312 20088 3328
rect 20022 3248 20023 3312
rect 20087 3248 20088 3312
rect 20022 3232 20088 3248
rect 20022 3168 20023 3232
rect 20087 3168 20088 3232
rect 20022 3152 20088 3168
rect 20022 3088 20023 3152
rect 20087 3088 20088 3152
rect 20022 3072 20088 3088
rect 20022 3008 20023 3072
rect 20087 3008 20088 3072
rect 20022 2992 20088 3008
rect 20022 2928 20023 2992
rect 20087 2928 20088 2992
rect 20022 2838 20088 2928
rect 20148 4872 20214 4962
rect 20148 4808 20149 4872
rect 20213 4808 20214 4872
rect 20148 4792 20214 4808
rect 20148 4728 20149 4792
rect 20213 4728 20214 4792
rect 20148 4712 20214 4728
rect 20148 4648 20149 4712
rect 20213 4648 20214 4712
rect 20148 4632 20214 4648
rect 20148 4568 20149 4632
rect 20213 4568 20214 4632
rect 20148 4552 20214 4568
rect 20148 4488 20149 4552
rect 20213 4488 20214 4552
rect 20148 4472 20214 4488
rect 20148 4408 20149 4472
rect 20213 4408 20214 4472
rect 20148 4392 20214 4408
rect 20148 4328 20149 4392
rect 20213 4328 20214 4392
rect 20148 4312 20214 4328
rect 20148 4248 20149 4312
rect 20213 4248 20214 4312
rect 20148 4232 20214 4248
rect 20148 4168 20149 4232
rect 20213 4168 20214 4232
rect 20148 4152 20214 4168
rect 20148 4088 20149 4152
rect 20213 4088 20214 4152
rect 20148 3934 20214 4088
rect 20274 3996 20334 5026
rect 20394 3934 20454 4966
rect 20514 3996 20574 5026
rect 20634 3934 20694 4966
rect 20754 4872 20820 4962
rect 20754 4808 20755 4872
rect 20819 4808 20820 4872
rect 20754 4792 20820 4808
rect 20754 4728 20755 4792
rect 20819 4728 20820 4792
rect 20754 4712 20820 4728
rect 20754 4648 20755 4712
rect 20819 4648 20820 4712
rect 20754 4632 20820 4648
rect 20754 4568 20755 4632
rect 20819 4568 20820 4632
rect 20754 4552 20820 4568
rect 20754 4488 20755 4552
rect 20819 4488 20820 4552
rect 20754 4472 20820 4488
rect 20754 4408 20755 4472
rect 20819 4408 20820 4472
rect 20754 4392 20820 4408
rect 20754 4328 20755 4392
rect 20819 4328 20820 4392
rect 20754 4312 20820 4328
rect 20754 4248 20755 4312
rect 20819 4248 20820 4312
rect 20754 4232 20820 4248
rect 20754 4168 20755 4232
rect 20819 4168 20820 4232
rect 20754 4152 20820 4168
rect 20754 4088 20755 4152
rect 20819 4088 20820 4152
rect 20754 3934 20820 4088
rect 20880 3996 20940 5026
rect 21000 3934 21060 4966
rect 21120 3996 21180 5026
rect 21240 3934 21300 4966
rect 21360 4872 21426 4962
rect 21360 4808 21361 4872
rect 21425 4808 21426 4872
rect 21360 4792 21426 4808
rect 21360 4728 21361 4792
rect 21425 4728 21426 4792
rect 21360 4712 21426 4728
rect 21360 4648 21361 4712
rect 21425 4648 21426 4712
rect 21360 4632 21426 4648
rect 21360 4568 21361 4632
rect 21425 4568 21426 4632
rect 21360 4552 21426 4568
rect 21360 4488 21361 4552
rect 21425 4488 21426 4552
rect 21360 4472 21426 4488
rect 21360 4408 21361 4472
rect 21425 4408 21426 4472
rect 21360 4392 21426 4408
rect 21360 4328 21361 4392
rect 21425 4328 21426 4392
rect 21360 4312 21426 4328
rect 21360 4248 21361 4312
rect 21425 4248 21426 4312
rect 21360 4232 21426 4248
rect 21360 4168 21361 4232
rect 21425 4168 21426 4232
rect 21360 4152 21426 4168
rect 21360 4088 21361 4152
rect 21425 4088 21426 4152
rect 21360 3934 21426 4088
rect 21486 3996 21546 5026
rect 21606 3934 21666 4966
rect 21726 3996 21786 5026
rect 21846 3934 21906 4966
rect 21966 4872 22032 4962
rect 21966 4808 21967 4872
rect 22031 4808 22032 4872
rect 21966 4792 22032 4808
rect 21966 4728 21967 4792
rect 22031 4728 22032 4792
rect 21966 4712 22032 4728
rect 21966 4648 21967 4712
rect 22031 4648 22032 4712
rect 21966 4632 22032 4648
rect 21966 4568 21967 4632
rect 22031 4568 22032 4632
rect 21966 4552 22032 4568
rect 21966 4488 21967 4552
rect 22031 4488 22032 4552
rect 21966 4472 22032 4488
rect 21966 4408 21967 4472
rect 22031 4408 22032 4472
rect 21966 4392 22032 4408
rect 21966 4328 21967 4392
rect 22031 4328 22032 4392
rect 21966 4312 22032 4328
rect 21966 4248 21967 4312
rect 22031 4248 22032 4312
rect 21966 4232 22032 4248
rect 21966 4168 21967 4232
rect 22031 4168 22032 4232
rect 21966 4152 22032 4168
rect 21966 4088 21967 4152
rect 22031 4088 22032 4152
rect 21966 3934 22032 4088
rect 22092 3996 22152 5026
rect 22212 3934 22272 4966
rect 22332 3996 22392 5026
rect 22452 3934 22512 4966
rect 22572 4872 22638 4962
rect 22572 4808 22573 4872
rect 22637 4808 22638 4872
rect 22572 4792 22638 4808
rect 22572 4728 22573 4792
rect 22637 4728 22638 4792
rect 22572 4712 22638 4728
rect 22572 4648 22573 4712
rect 22637 4648 22638 4712
rect 22572 4632 22638 4648
rect 22572 4568 22573 4632
rect 22637 4568 22638 4632
rect 22572 4552 22638 4568
rect 22572 4488 22573 4552
rect 22637 4488 22638 4552
rect 22572 4472 22638 4488
rect 22572 4408 22573 4472
rect 22637 4408 22638 4472
rect 22572 4392 22638 4408
rect 22572 4328 22573 4392
rect 22637 4328 22638 4392
rect 22572 4312 22638 4328
rect 22572 4248 22573 4312
rect 22637 4248 22638 4312
rect 22572 4232 22638 4248
rect 22572 4168 22573 4232
rect 22637 4168 22638 4232
rect 22572 4152 22638 4168
rect 22572 4088 22573 4152
rect 22637 4088 22638 4152
rect 22572 3934 22638 4088
rect 22698 3996 22758 5026
rect 22818 3934 22878 4966
rect 22938 3996 22998 5026
rect 23058 3934 23118 4966
rect 23178 4872 23244 4962
rect 23178 4808 23179 4872
rect 23243 4808 23244 4872
rect 23178 4792 23244 4808
rect 23178 4728 23179 4792
rect 23243 4728 23244 4792
rect 23178 4712 23244 4728
rect 23178 4648 23179 4712
rect 23243 4648 23244 4712
rect 23178 4632 23244 4648
rect 23178 4568 23179 4632
rect 23243 4568 23244 4632
rect 23178 4552 23244 4568
rect 23178 4488 23179 4552
rect 23243 4488 23244 4552
rect 23178 4472 23244 4488
rect 23178 4408 23179 4472
rect 23243 4408 23244 4472
rect 23178 4392 23244 4408
rect 23178 4328 23179 4392
rect 23243 4328 23244 4392
rect 23178 4312 23244 4328
rect 23178 4248 23179 4312
rect 23243 4248 23244 4312
rect 23178 4232 23244 4248
rect 23178 4168 23179 4232
rect 23243 4168 23244 4232
rect 23178 4152 23244 4168
rect 23178 4088 23179 4152
rect 23243 4088 23244 4152
rect 23178 3934 23244 4088
rect 23304 3996 23364 5026
rect 23424 3934 23484 4966
rect 23544 3996 23604 5026
rect 23664 3934 23724 4966
rect 23784 4872 23850 4962
rect 23784 4808 23785 4872
rect 23849 4808 23850 4872
rect 23784 4792 23850 4808
rect 23784 4728 23785 4792
rect 23849 4728 23850 4792
rect 23784 4712 23850 4728
rect 23784 4648 23785 4712
rect 23849 4648 23850 4712
rect 23784 4632 23850 4648
rect 23784 4568 23785 4632
rect 23849 4568 23850 4632
rect 23784 4552 23850 4568
rect 23784 4488 23785 4552
rect 23849 4488 23850 4552
rect 23784 4472 23850 4488
rect 23784 4408 23785 4472
rect 23849 4408 23850 4472
rect 23784 4392 23850 4408
rect 23784 4328 23785 4392
rect 23849 4328 23850 4392
rect 23784 4312 23850 4328
rect 23784 4248 23785 4312
rect 23849 4248 23850 4312
rect 23784 4232 23850 4248
rect 23784 4168 23785 4232
rect 23849 4168 23850 4232
rect 23784 4152 23850 4168
rect 23784 4088 23785 4152
rect 23849 4088 23850 4152
rect 23784 3934 23850 4088
rect 23910 3996 23970 5026
rect 24030 3934 24090 4966
rect 24150 3996 24210 5026
rect 24270 3934 24330 4966
rect 24390 4872 24456 4962
rect 24390 4808 24391 4872
rect 24455 4808 24456 4872
rect 24390 4792 24456 4808
rect 24390 4728 24391 4792
rect 24455 4728 24456 4792
rect 24390 4712 24456 4728
rect 24390 4648 24391 4712
rect 24455 4648 24456 4712
rect 24390 4632 24456 4648
rect 24390 4568 24391 4632
rect 24455 4568 24456 4632
rect 24390 4552 24456 4568
rect 24390 4488 24391 4552
rect 24455 4488 24456 4552
rect 24390 4472 24456 4488
rect 24390 4408 24391 4472
rect 24455 4408 24456 4472
rect 24390 4392 24456 4408
rect 24390 4328 24391 4392
rect 24455 4328 24456 4392
rect 24390 4312 24456 4328
rect 24390 4248 24391 4312
rect 24455 4248 24456 4312
rect 24390 4232 24456 4248
rect 24390 4168 24391 4232
rect 24455 4168 24456 4232
rect 24390 4152 24456 4168
rect 24390 4088 24391 4152
rect 24455 4088 24456 4152
rect 24390 3934 24456 4088
rect 24516 3996 24576 5026
rect 24636 3934 24696 4966
rect 24756 3996 24816 5026
rect 24876 3934 24936 4966
rect 24996 4872 25062 4962
rect 24996 4808 24997 4872
rect 25061 4808 25062 4872
rect 24996 4792 25062 4808
rect 24996 4728 24997 4792
rect 25061 4728 25062 4792
rect 24996 4712 25062 4728
rect 24996 4648 24997 4712
rect 25061 4648 25062 4712
rect 24996 4632 25062 4648
rect 24996 4568 24997 4632
rect 25061 4568 25062 4632
rect 24996 4552 25062 4568
rect 24996 4488 24997 4552
rect 25061 4488 25062 4552
rect 24996 4472 25062 4488
rect 24996 4408 24997 4472
rect 25061 4408 25062 4472
rect 24996 4392 25062 4408
rect 24996 4328 24997 4392
rect 25061 4328 25062 4392
rect 24996 4312 25062 4328
rect 24996 4248 24997 4312
rect 25061 4248 25062 4312
rect 24996 4232 25062 4248
rect 24996 4168 24997 4232
rect 25061 4168 25062 4232
rect 24996 4152 25062 4168
rect 24996 4088 24997 4152
rect 25061 4088 25062 4152
rect 24996 3934 25062 4088
rect 25122 3996 25182 5026
rect 25242 3934 25302 4966
rect 25362 3996 25422 5026
rect 25482 3934 25542 4966
rect 25602 4872 25668 4962
rect 25602 4808 25603 4872
rect 25667 4808 25668 4872
rect 25602 4792 25668 4808
rect 25602 4728 25603 4792
rect 25667 4728 25668 4792
rect 25602 4712 25668 4728
rect 25602 4648 25603 4712
rect 25667 4648 25668 4712
rect 25602 4632 25668 4648
rect 25602 4568 25603 4632
rect 25667 4568 25668 4632
rect 25602 4552 25668 4568
rect 25602 4488 25603 4552
rect 25667 4488 25668 4552
rect 25602 4472 25668 4488
rect 25602 4408 25603 4472
rect 25667 4408 25668 4472
rect 25602 4392 25668 4408
rect 25602 4328 25603 4392
rect 25667 4328 25668 4392
rect 25602 4312 25668 4328
rect 25602 4248 25603 4312
rect 25667 4248 25668 4312
rect 25602 4232 25668 4248
rect 25602 4168 25603 4232
rect 25667 4168 25668 4232
rect 25602 4152 25668 4168
rect 25602 4088 25603 4152
rect 25667 4088 25668 4152
rect 25602 3934 25668 4088
rect 25728 3996 25788 5026
rect 25848 3934 25908 4966
rect 25968 3996 26028 5026
rect 26088 3934 26148 4966
rect 26208 4872 26274 4962
rect 26208 4808 26209 4872
rect 26273 4808 26274 4872
rect 26208 4792 26274 4808
rect 26208 4728 26209 4792
rect 26273 4728 26274 4792
rect 26208 4712 26274 4728
rect 26208 4648 26209 4712
rect 26273 4648 26274 4712
rect 26208 4632 26274 4648
rect 26208 4568 26209 4632
rect 26273 4568 26274 4632
rect 26208 4552 26274 4568
rect 26208 4488 26209 4552
rect 26273 4488 26274 4552
rect 26208 4472 26274 4488
rect 26208 4408 26209 4472
rect 26273 4408 26274 4472
rect 26208 4392 26274 4408
rect 26208 4328 26209 4392
rect 26273 4328 26274 4392
rect 26208 4312 26274 4328
rect 26208 4248 26209 4312
rect 26273 4248 26274 4312
rect 26208 4232 26274 4248
rect 26208 4168 26209 4232
rect 26273 4168 26274 4232
rect 26208 4152 26274 4168
rect 26208 4088 26209 4152
rect 26273 4088 26274 4152
rect 26208 3934 26274 4088
rect 26334 3996 26394 5026
rect 26454 3934 26514 4966
rect 26574 3996 26634 5026
rect 26694 3934 26754 4966
rect 26814 4872 26880 4962
rect 26814 4808 26815 4872
rect 26879 4808 26880 4872
rect 26814 4792 26880 4808
rect 26814 4728 26815 4792
rect 26879 4728 26880 4792
rect 26814 4712 26880 4728
rect 26814 4648 26815 4712
rect 26879 4648 26880 4712
rect 26814 4632 26880 4648
rect 26814 4568 26815 4632
rect 26879 4568 26880 4632
rect 26814 4552 26880 4568
rect 26814 4488 26815 4552
rect 26879 4488 26880 4552
rect 26814 4472 26880 4488
rect 26814 4408 26815 4472
rect 26879 4408 26880 4472
rect 26814 4392 26880 4408
rect 26814 4328 26815 4392
rect 26879 4328 26880 4392
rect 26814 4312 26880 4328
rect 26814 4248 26815 4312
rect 26879 4248 26880 4312
rect 26814 4232 26880 4248
rect 26814 4168 26815 4232
rect 26879 4168 26880 4232
rect 26814 4152 26880 4168
rect 26814 4088 26815 4152
rect 26879 4088 26880 4152
rect 26814 3934 26880 4088
rect 26940 3996 27000 5026
rect 27060 3934 27120 4966
rect 27180 3996 27240 5026
rect 27300 3934 27360 4966
rect 27420 4872 27486 4962
rect 27420 4808 27421 4872
rect 27485 4808 27486 4872
rect 27420 4792 27486 4808
rect 27420 4728 27421 4792
rect 27485 4728 27486 4792
rect 27420 4712 27486 4728
rect 27420 4648 27421 4712
rect 27485 4648 27486 4712
rect 27420 4632 27486 4648
rect 27420 4568 27421 4632
rect 27485 4568 27486 4632
rect 27420 4552 27486 4568
rect 27420 4488 27421 4552
rect 27485 4488 27486 4552
rect 27420 4472 27486 4488
rect 27420 4408 27421 4472
rect 27485 4408 27486 4472
rect 27420 4392 27486 4408
rect 27420 4328 27421 4392
rect 27485 4328 27486 4392
rect 27420 4312 27486 4328
rect 27420 4248 27421 4312
rect 27485 4248 27486 4312
rect 27420 4232 27486 4248
rect 27420 4168 27421 4232
rect 27485 4168 27486 4232
rect 27420 4152 27486 4168
rect 27420 4088 27421 4152
rect 27485 4088 27486 4152
rect 27420 3934 27486 4088
rect 27546 3996 27606 5026
rect 27666 3934 27726 4966
rect 27786 3996 27846 5026
rect 27906 3934 27966 4966
rect 28026 4872 28092 4962
rect 28026 4808 28027 4872
rect 28091 4808 28092 4872
rect 28026 4792 28092 4808
rect 28026 4728 28027 4792
rect 28091 4728 28092 4792
rect 28026 4712 28092 4728
rect 28026 4648 28027 4712
rect 28091 4648 28092 4712
rect 28026 4632 28092 4648
rect 28026 4568 28027 4632
rect 28091 4568 28092 4632
rect 28026 4552 28092 4568
rect 28026 4488 28027 4552
rect 28091 4488 28092 4552
rect 28026 4472 28092 4488
rect 28026 4408 28027 4472
rect 28091 4408 28092 4472
rect 28026 4392 28092 4408
rect 28026 4328 28027 4392
rect 28091 4328 28092 4392
rect 28026 4312 28092 4328
rect 28026 4248 28027 4312
rect 28091 4248 28092 4312
rect 28026 4232 28092 4248
rect 28026 4168 28027 4232
rect 28091 4168 28092 4232
rect 28026 4152 28092 4168
rect 28026 4088 28027 4152
rect 28091 4088 28092 4152
rect 28026 3934 28092 4088
rect 28152 3996 28212 5026
rect 28272 3934 28332 4966
rect 28392 3996 28452 5026
rect 28512 3934 28572 4966
rect 28632 4872 28698 4962
rect 28632 4808 28633 4872
rect 28697 4808 28698 4872
rect 28632 4792 28698 4808
rect 28632 4728 28633 4792
rect 28697 4728 28698 4792
rect 28632 4712 28698 4728
rect 28632 4648 28633 4712
rect 28697 4648 28698 4712
rect 28632 4632 28698 4648
rect 28632 4568 28633 4632
rect 28697 4568 28698 4632
rect 28632 4552 28698 4568
rect 28632 4488 28633 4552
rect 28697 4488 28698 4552
rect 28632 4472 28698 4488
rect 28632 4408 28633 4472
rect 28697 4408 28698 4472
rect 28632 4392 28698 4408
rect 28632 4328 28633 4392
rect 28697 4328 28698 4392
rect 28632 4312 28698 4328
rect 28632 4248 28633 4312
rect 28697 4248 28698 4312
rect 28632 4232 28698 4248
rect 28632 4168 28633 4232
rect 28697 4168 28698 4232
rect 28632 4152 28698 4168
rect 28632 4088 28633 4152
rect 28697 4088 28698 4152
rect 28632 3934 28698 4088
rect 28758 3996 28818 5026
rect 28878 3934 28938 4966
rect 28998 3996 29058 5026
rect 29118 3934 29178 4966
rect 29238 4872 29304 4962
rect 29238 4808 29239 4872
rect 29303 4808 29304 4872
rect 29238 4792 29304 4808
rect 29238 4728 29239 4792
rect 29303 4728 29304 4792
rect 29238 4712 29304 4728
rect 29238 4648 29239 4712
rect 29303 4648 29304 4712
rect 29238 4632 29304 4648
rect 29238 4568 29239 4632
rect 29303 4568 29304 4632
rect 29238 4552 29304 4568
rect 29238 4488 29239 4552
rect 29303 4488 29304 4552
rect 29238 4472 29304 4488
rect 29238 4408 29239 4472
rect 29303 4408 29304 4472
rect 29238 4392 29304 4408
rect 29238 4328 29239 4392
rect 29303 4328 29304 4392
rect 29238 4312 29304 4328
rect 29238 4248 29239 4312
rect 29303 4248 29304 4312
rect 29238 4232 29304 4248
rect 29238 4168 29239 4232
rect 29303 4168 29304 4232
rect 29238 4152 29304 4168
rect 29238 4088 29239 4152
rect 29303 4088 29304 4152
rect 29238 3934 29304 4088
rect 29364 3996 29424 5026
rect 29484 3934 29544 4966
rect 29604 3996 29664 5026
rect 29724 3934 29784 4966
rect 29844 4872 29910 4962
rect 29844 4808 29845 4872
rect 29909 4808 29910 4872
rect 29844 4792 29910 4808
rect 29844 4728 29845 4792
rect 29909 4728 29910 4792
rect 29844 4712 29910 4728
rect 29844 4648 29845 4712
rect 29909 4648 29910 4712
rect 29844 4632 29910 4648
rect 29844 4568 29845 4632
rect 29909 4568 29910 4632
rect 29844 4552 29910 4568
rect 29844 4488 29845 4552
rect 29909 4488 29910 4552
rect 29844 4472 29910 4488
rect 29844 4408 29845 4472
rect 29909 4408 29910 4472
rect 29844 4392 29910 4408
rect 29844 4328 29845 4392
rect 29909 4328 29910 4392
rect 29844 4312 29910 4328
rect 29844 4248 29845 4312
rect 29909 4248 29910 4312
rect 29844 4232 29910 4248
rect 29844 4168 29845 4232
rect 29909 4168 29910 4232
rect 29844 4152 29910 4168
rect 29844 4088 29845 4152
rect 29909 4088 29910 4152
rect 29844 3934 29910 4088
rect 29970 3996 30030 5026
rect 30090 3934 30150 4966
rect 30210 3996 30270 5026
rect 30330 3934 30390 4966
rect 30450 4872 30516 4962
rect 30450 4808 30451 4872
rect 30515 4808 30516 4872
rect 30450 4792 30516 4808
rect 30450 4728 30451 4792
rect 30515 4728 30516 4792
rect 30450 4712 30516 4728
rect 30450 4648 30451 4712
rect 30515 4648 30516 4712
rect 30450 4632 30516 4648
rect 30450 4568 30451 4632
rect 30515 4568 30516 4632
rect 30450 4552 30516 4568
rect 30450 4488 30451 4552
rect 30515 4488 30516 4552
rect 30450 4472 30516 4488
rect 30450 4408 30451 4472
rect 30515 4408 30516 4472
rect 30450 4392 30516 4408
rect 30450 4328 30451 4392
rect 30515 4328 30516 4392
rect 30450 4312 30516 4328
rect 30450 4248 30451 4312
rect 30515 4248 30516 4312
rect 30450 4232 30516 4248
rect 30450 4168 30451 4232
rect 30515 4168 30516 4232
rect 30450 4152 30516 4168
rect 30450 4088 30451 4152
rect 30515 4088 30516 4152
rect 30450 3934 30516 4088
rect 30576 3996 30636 5026
rect 30696 3934 30756 4966
rect 30816 3996 30876 5026
rect 30936 3934 30996 4966
rect 31056 4872 31122 4962
rect 31056 4808 31057 4872
rect 31121 4808 31122 4872
rect 31056 4792 31122 4808
rect 31056 4728 31057 4792
rect 31121 4728 31122 4792
rect 31056 4712 31122 4728
rect 31056 4648 31057 4712
rect 31121 4648 31122 4712
rect 31056 4632 31122 4648
rect 31056 4568 31057 4632
rect 31121 4568 31122 4632
rect 31056 4552 31122 4568
rect 31056 4488 31057 4552
rect 31121 4488 31122 4552
rect 31056 4472 31122 4488
rect 31056 4408 31057 4472
rect 31121 4408 31122 4472
rect 31056 4392 31122 4408
rect 31056 4328 31057 4392
rect 31121 4328 31122 4392
rect 31056 4312 31122 4328
rect 31056 4248 31057 4312
rect 31121 4248 31122 4312
rect 31056 4232 31122 4248
rect 31056 4168 31057 4232
rect 31121 4168 31122 4232
rect 31056 4152 31122 4168
rect 31056 4088 31057 4152
rect 31121 4088 31122 4152
rect 31056 3934 31122 4088
rect 31182 3996 31242 5026
rect 31302 3934 31362 4966
rect 31422 3996 31482 5026
rect 31542 3934 31602 4966
rect 31662 4872 31728 4962
rect 31662 4808 31663 4872
rect 31727 4808 31728 4872
rect 31662 4792 31728 4808
rect 31662 4728 31663 4792
rect 31727 4728 31728 4792
rect 31662 4712 31728 4728
rect 31662 4648 31663 4712
rect 31727 4648 31728 4712
rect 31662 4632 31728 4648
rect 31662 4568 31663 4632
rect 31727 4568 31728 4632
rect 31662 4552 31728 4568
rect 31662 4488 31663 4552
rect 31727 4488 31728 4552
rect 31662 4472 31728 4488
rect 31662 4408 31663 4472
rect 31727 4408 31728 4472
rect 31662 4392 31728 4408
rect 31662 4328 31663 4392
rect 31727 4328 31728 4392
rect 31662 4312 31728 4328
rect 31662 4248 31663 4312
rect 31727 4248 31728 4312
rect 31662 4232 31728 4248
rect 31662 4168 31663 4232
rect 31727 4168 31728 4232
rect 31662 4152 31728 4168
rect 31662 4088 31663 4152
rect 31727 4088 31728 4152
rect 31662 3934 31728 4088
rect 31788 3996 31848 5026
rect 31908 3934 31968 4966
rect 32028 3996 32088 5026
rect 32148 3934 32208 4966
rect 32268 4872 32334 4962
rect 32268 4808 32269 4872
rect 32333 4808 32334 4872
rect 32268 4792 32334 4808
rect 32268 4728 32269 4792
rect 32333 4728 32334 4792
rect 32268 4712 32334 4728
rect 32268 4648 32269 4712
rect 32333 4648 32334 4712
rect 32268 4632 32334 4648
rect 32268 4568 32269 4632
rect 32333 4568 32334 4632
rect 32268 4552 32334 4568
rect 32268 4488 32269 4552
rect 32333 4488 32334 4552
rect 32268 4472 32334 4488
rect 32268 4408 32269 4472
rect 32333 4408 32334 4472
rect 32268 4392 32334 4408
rect 32268 4328 32269 4392
rect 32333 4328 32334 4392
rect 32268 4312 32334 4328
rect 32268 4248 32269 4312
rect 32333 4248 32334 4312
rect 32268 4232 32334 4248
rect 32268 4168 32269 4232
rect 32333 4168 32334 4232
rect 32268 4152 32334 4168
rect 32268 4088 32269 4152
rect 32333 4088 32334 4152
rect 32268 3934 32334 4088
rect 32394 3996 32454 5026
rect 32514 3934 32574 4966
rect 32634 3996 32694 5026
rect 32754 3934 32814 4966
rect 32874 4872 32940 4962
rect 32874 4808 32875 4872
rect 32939 4808 32940 4872
rect 32874 4792 32940 4808
rect 32874 4728 32875 4792
rect 32939 4728 32940 4792
rect 32874 4712 32940 4728
rect 32874 4648 32875 4712
rect 32939 4648 32940 4712
rect 32874 4632 32940 4648
rect 32874 4568 32875 4632
rect 32939 4568 32940 4632
rect 32874 4552 32940 4568
rect 32874 4488 32875 4552
rect 32939 4488 32940 4552
rect 32874 4472 32940 4488
rect 32874 4408 32875 4472
rect 32939 4408 32940 4472
rect 32874 4392 32940 4408
rect 32874 4328 32875 4392
rect 32939 4328 32940 4392
rect 32874 4312 32940 4328
rect 32874 4248 32875 4312
rect 32939 4248 32940 4312
rect 32874 4232 32940 4248
rect 32874 4168 32875 4232
rect 32939 4168 32940 4232
rect 32874 4152 32940 4168
rect 32874 4088 32875 4152
rect 32939 4088 32940 4152
rect 32874 3934 32940 4088
rect 33000 3996 33060 5026
rect 33120 3934 33180 4966
rect 33240 3996 33300 5026
rect 33360 3934 33420 4966
rect 33480 4872 33546 4962
rect 33480 4808 33481 4872
rect 33545 4808 33546 4872
rect 33480 4792 33546 4808
rect 33480 4728 33481 4792
rect 33545 4728 33546 4792
rect 33480 4712 33546 4728
rect 33480 4648 33481 4712
rect 33545 4648 33546 4712
rect 33480 4632 33546 4648
rect 33480 4568 33481 4632
rect 33545 4568 33546 4632
rect 33480 4552 33546 4568
rect 33480 4488 33481 4552
rect 33545 4488 33546 4552
rect 33480 4472 33546 4488
rect 33480 4408 33481 4472
rect 33545 4408 33546 4472
rect 33480 4392 33546 4408
rect 33480 4328 33481 4392
rect 33545 4328 33546 4392
rect 33480 4312 33546 4328
rect 33480 4248 33481 4312
rect 33545 4248 33546 4312
rect 33480 4232 33546 4248
rect 33480 4168 33481 4232
rect 33545 4168 33546 4232
rect 33480 4152 33546 4168
rect 33480 4088 33481 4152
rect 33545 4088 33546 4152
rect 33480 3934 33546 4088
rect 33606 3996 33666 5026
rect 33726 3934 33786 4966
rect 33846 3996 33906 5026
rect 33966 3934 34026 4966
rect 34086 4872 34152 4962
rect 34086 4808 34087 4872
rect 34151 4808 34152 4872
rect 34086 4792 34152 4808
rect 34086 4728 34087 4792
rect 34151 4728 34152 4792
rect 34086 4712 34152 4728
rect 34086 4648 34087 4712
rect 34151 4648 34152 4712
rect 34086 4632 34152 4648
rect 34086 4568 34087 4632
rect 34151 4568 34152 4632
rect 34086 4552 34152 4568
rect 34086 4488 34087 4552
rect 34151 4488 34152 4552
rect 34086 4472 34152 4488
rect 34086 4408 34087 4472
rect 34151 4408 34152 4472
rect 34086 4392 34152 4408
rect 34086 4328 34087 4392
rect 34151 4328 34152 4392
rect 34086 4312 34152 4328
rect 34086 4248 34087 4312
rect 34151 4248 34152 4312
rect 34086 4232 34152 4248
rect 34086 4168 34087 4232
rect 34151 4168 34152 4232
rect 34086 4152 34152 4168
rect 34086 4088 34087 4152
rect 34151 4088 34152 4152
rect 34086 3934 34152 4088
rect 34212 3996 34272 5026
rect 34332 3934 34392 4966
rect 34452 3996 34512 5026
rect 34572 3934 34632 4966
rect 34692 4872 34758 4962
rect 34692 4808 34693 4872
rect 34757 4808 34758 4872
rect 34692 4792 34758 4808
rect 34692 4728 34693 4792
rect 34757 4728 34758 4792
rect 34692 4712 34758 4728
rect 34692 4648 34693 4712
rect 34757 4648 34758 4712
rect 34692 4632 34758 4648
rect 34692 4568 34693 4632
rect 34757 4568 34758 4632
rect 34692 4552 34758 4568
rect 34692 4488 34693 4552
rect 34757 4488 34758 4552
rect 34692 4472 34758 4488
rect 34692 4408 34693 4472
rect 34757 4408 34758 4472
rect 34692 4392 34758 4408
rect 34692 4328 34693 4392
rect 34757 4328 34758 4392
rect 34692 4312 34758 4328
rect 34692 4248 34693 4312
rect 34757 4248 34758 4312
rect 34692 4232 34758 4248
rect 34692 4168 34693 4232
rect 34757 4168 34758 4232
rect 34692 4152 34758 4168
rect 34692 4088 34693 4152
rect 34757 4088 34758 4152
rect 34692 3934 34758 4088
rect 34818 3996 34878 5026
rect 34938 3934 34998 4966
rect 35058 3996 35118 5026
rect 35178 3934 35238 4966
rect 35298 4872 35364 4962
rect 35298 4808 35299 4872
rect 35363 4808 35364 4872
rect 35298 4792 35364 4808
rect 35298 4728 35299 4792
rect 35363 4728 35364 4792
rect 35298 4712 35364 4728
rect 35298 4648 35299 4712
rect 35363 4648 35364 4712
rect 35298 4632 35364 4648
rect 35298 4568 35299 4632
rect 35363 4568 35364 4632
rect 35298 4552 35364 4568
rect 35298 4488 35299 4552
rect 35363 4488 35364 4552
rect 35298 4472 35364 4488
rect 35298 4408 35299 4472
rect 35363 4408 35364 4472
rect 35298 4392 35364 4408
rect 35298 4328 35299 4392
rect 35363 4328 35364 4392
rect 35298 4312 35364 4328
rect 35298 4248 35299 4312
rect 35363 4248 35364 4312
rect 35298 4232 35364 4248
rect 35298 4168 35299 4232
rect 35363 4168 35364 4232
rect 35298 4152 35364 4168
rect 35298 4088 35299 4152
rect 35363 4088 35364 4152
rect 35298 3934 35364 4088
rect 35424 3996 35484 5026
rect 35544 3934 35604 4966
rect 35664 3996 35724 5026
rect 35784 3934 35844 4966
rect 35904 4872 35970 4962
rect 35904 4808 35905 4872
rect 35969 4808 35970 4872
rect 35904 4792 35970 4808
rect 35904 4728 35905 4792
rect 35969 4728 35970 4792
rect 35904 4712 35970 4728
rect 35904 4648 35905 4712
rect 35969 4648 35970 4712
rect 35904 4632 35970 4648
rect 35904 4568 35905 4632
rect 35969 4568 35970 4632
rect 35904 4552 35970 4568
rect 35904 4488 35905 4552
rect 35969 4488 35970 4552
rect 35904 4472 35970 4488
rect 35904 4408 35905 4472
rect 35969 4408 35970 4472
rect 35904 4392 35970 4408
rect 35904 4328 35905 4392
rect 35969 4328 35970 4392
rect 35904 4312 35970 4328
rect 35904 4248 35905 4312
rect 35969 4248 35970 4312
rect 35904 4232 35970 4248
rect 35904 4168 35905 4232
rect 35969 4168 35970 4232
rect 35904 4152 35970 4168
rect 35904 4088 35905 4152
rect 35969 4088 35970 4152
rect 35904 3934 35970 4088
rect 36030 3996 36090 5026
rect 36150 3934 36210 4966
rect 36270 3996 36330 5026
rect 36390 3934 36450 4966
rect 36510 4872 36576 4962
rect 36510 4808 36511 4872
rect 36575 4808 36576 4872
rect 36510 4792 36576 4808
rect 36510 4728 36511 4792
rect 36575 4728 36576 4792
rect 36510 4712 36576 4728
rect 36510 4648 36511 4712
rect 36575 4648 36576 4712
rect 36510 4632 36576 4648
rect 36510 4568 36511 4632
rect 36575 4568 36576 4632
rect 36510 4552 36576 4568
rect 36510 4488 36511 4552
rect 36575 4488 36576 4552
rect 36510 4472 36576 4488
rect 36510 4408 36511 4472
rect 36575 4408 36576 4472
rect 36510 4392 36576 4408
rect 36510 4328 36511 4392
rect 36575 4328 36576 4392
rect 36510 4312 36576 4328
rect 36510 4248 36511 4312
rect 36575 4248 36576 4312
rect 36510 4232 36576 4248
rect 36510 4168 36511 4232
rect 36575 4168 36576 4232
rect 36510 4152 36576 4168
rect 36510 4088 36511 4152
rect 36575 4088 36576 4152
rect 36510 3934 36576 4088
rect 36636 3996 36696 5026
rect 36756 3934 36816 4966
rect 36876 3996 36936 5026
rect 36996 3934 37056 4966
rect 37116 4872 37182 4962
rect 37116 4808 37117 4872
rect 37181 4808 37182 4872
rect 37116 4792 37182 4808
rect 37116 4728 37117 4792
rect 37181 4728 37182 4792
rect 37116 4712 37182 4728
rect 37116 4648 37117 4712
rect 37181 4648 37182 4712
rect 37116 4632 37182 4648
rect 37116 4568 37117 4632
rect 37181 4568 37182 4632
rect 37116 4552 37182 4568
rect 37116 4488 37117 4552
rect 37181 4488 37182 4552
rect 37116 4472 37182 4488
rect 37116 4408 37117 4472
rect 37181 4408 37182 4472
rect 37116 4392 37182 4408
rect 37116 4328 37117 4392
rect 37181 4328 37182 4392
rect 37116 4312 37182 4328
rect 37116 4248 37117 4312
rect 37181 4248 37182 4312
rect 37116 4232 37182 4248
rect 37116 4168 37117 4232
rect 37181 4168 37182 4232
rect 37116 4152 37182 4168
rect 37116 4088 37117 4152
rect 37181 4088 37182 4152
rect 37116 3934 37182 4088
rect 37242 3996 37302 5026
rect 37362 3934 37422 4966
rect 37482 3996 37542 5026
rect 37602 3934 37662 4966
rect 37722 4872 37788 4962
rect 37722 4808 37723 4872
rect 37787 4808 37788 4872
rect 37722 4792 37788 4808
rect 37722 4728 37723 4792
rect 37787 4728 37788 4792
rect 37722 4712 37788 4728
rect 37722 4648 37723 4712
rect 37787 4648 37788 4712
rect 37722 4632 37788 4648
rect 37722 4568 37723 4632
rect 37787 4568 37788 4632
rect 37722 4552 37788 4568
rect 37722 4488 37723 4552
rect 37787 4488 37788 4552
rect 37722 4472 37788 4488
rect 37722 4408 37723 4472
rect 37787 4408 37788 4472
rect 37722 4392 37788 4408
rect 37722 4328 37723 4392
rect 37787 4328 37788 4392
rect 37722 4312 37788 4328
rect 37722 4248 37723 4312
rect 37787 4248 37788 4312
rect 37722 4232 37788 4248
rect 37722 4168 37723 4232
rect 37787 4168 37788 4232
rect 37722 4152 37788 4168
rect 37722 4088 37723 4152
rect 37787 4088 37788 4152
rect 37722 3934 37788 4088
rect 37848 3996 37908 5026
rect 37968 3934 38028 4966
rect 38088 3996 38148 5026
rect 38208 3934 38268 4966
rect 38328 4872 38394 4962
rect 38328 4808 38329 4872
rect 38393 4808 38394 4872
rect 38328 4792 38394 4808
rect 38328 4728 38329 4792
rect 38393 4728 38394 4792
rect 38328 4712 38394 4728
rect 38328 4648 38329 4712
rect 38393 4648 38394 4712
rect 38328 4632 38394 4648
rect 38328 4568 38329 4632
rect 38393 4568 38394 4632
rect 38328 4552 38394 4568
rect 38328 4488 38329 4552
rect 38393 4488 38394 4552
rect 38328 4472 38394 4488
rect 38328 4408 38329 4472
rect 38393 4408 38394 4472
rect 38328 4392 38394 4408
rect 38328 4328 38329 4392
rect 38393 4328 38394 4392
rect 38328 4312 38394 4328
rect 38328 4248 38329 4312
rect 38393 4248 38394 4312
rect 38328 4232 38394 4248
rect 38328 4168 38329 4232
rect 38393 4168 38394 4232
rect 38328 4152 38394 4168
rect 38328 4088 38329 4152
rect 38393 4088 38394 4152
rect 38328 3934 38394 4088
rect 38454 3996 38514 5026
rect 38574 3934 38634 4966
rect 38694 3996 38754 5026
rect 38814 3934 38874 4966
rect 38934 4872 39000 4962
rect 38934 4808 38935 4872
rect 38999 4808 39000 4872
rect 38934 4792 39000 4808
rect 38934 4728 38935 4792
rect 38999 4728 39000 4792
rect 38934 4712 39000 4728
rect 38934 4648 38935 4712
rect 38999 4648 39000 4712
rect 38934 4632 39000 4648
rect 38934 4568 38935 4632
rect 38999 4568 39000 4632
rect 38934 4552 39000 4568
rect 38934 4488 38935 4552
rect 38999 4488 39000 4552
rect 38934 4472 39000 4488
rect 38934 4408 38935 4472
rect 38999 4408 39000 4472
rect 38934 4392 39000 4408
rect 38934 4328 38935 4392
rect 38999 4328 39000 4392
rect 38934 4312 39000 4328
rect 38934 4248 38935 4312
rect 38999 4248 39000 4312
rect 38934 4232 39000 4248
rect 38934 4168 38935 4232
rect 38999 4168 39000 4232
rect 38934 4152 39000 4168
rect 38934 4088 38935 4152
rect 38999 4088 39000 4152
rect 38934 3934 39000 4088
rect 39060 3996 39120 5026
rect 39180 3934 39240 4966
rect 39300 3996 39360 5026
rect 39420 3934 39480 4966
rect 39540 4872 39606 4962
rect 39540 4808 39541 4872
rect 39605 4808 39606 4872
rect 39540 4792 39606 4808
rect 39540 4728 39541 4792
rect 39605 4728 39606 4792
rect 39540 4712 39606 4728
rect 39540 4648 39541 4712
rect 39605 4648 39606 4712
rect 39540 4632 39606 4648
rect 39540 4568 39541 4632
rect 39605 4568 39606 4632
rect 39540 4552 39606 4568
rect 39540 4488 39541 4552
rect 39605 4488 39606 4552
rect 39540 4472 39606 4488
rect 39540 4408 39541 4472
rect 39605 4408 39606 4472
rect 39540 4392 39606 4408
rect 39540 4328 39541 4392
rect 39605 4328 39606 4392
rect 39540 4312 39606 4328
rect 39540 4248 39541 4312
rect 39605 4248 39606 4312
rect 39540 4232 39606 4248
rect 39540 4168 39541 4232
rect 39605 4168 39606 4232
rect 39540 4152 39606 4168
rect 39540 4088 39541 4152
rect 39605 4088 39606 4152
rect 39540 3934 39606 4088
rect 20148 3932 39606 3934
rect 20148 3868 20252 3932
rect 20316 3868 20332 3932
rect 20396 3868 20412 3932
rect 20476 3868 20492 3932
rect 20556 3868 20572 3932
rect 20636 3868 20652 3932
rect 20716 3868 20858 3932
rect 20922 3868 20938 3932
rect 21002 3868 21018 3932
rect 21082 3868 21098 3932
rect 21162 3868 21178 3932
rect 21242 3868 21258 3932
rect 21322 3868 21464 3932
rect 21528 3868 21544 3932
rect 21608 3868 21624 3932
rect 21688 3868 21704 3932
rect 21768 3868 21784 3932
rect 21848 3868 21864 3932
rect 21928 3868 22070 3932
rect 22134 3868 22150 3932
rect 22214 3868 22230 3932
rect 22294 3868 22310 3932
rect 22374 3868 22390 3932
rect 22454 3868 22470 3932
rect 22534 3868 22676 3932
rect 22740 3868 22756 3932
rect 22820 3868 22836 3932
rect 22900 3868 22916 3932
rect 22980 3868 22996 3932
rect 23060 3868 23076 3932
rect 23140 3868 23282 3932
rect 23346 3868 23362 3932
rect 23426 3868 23442 3932
rect 23506 3868 23522 3932
rect 23586 3868 23602 3932
rect 23666 3868 23682 3932
rect 23746 3868 23888 3932
rect 23952 3868 23968 3932
rect 24032 3868 24048 3932
rect 24112 3868 24128 3932
rect 24192 3868 24208 3932
rect 24272 3868 24288 3932
rect 24352 3868 24494 3932
rect 24558 3868 24574 3932
rect 24638 3868 24654 3932
rect 24718 3868 24734 3932
rect 24798 3868 24814 3932
rect 24878 3868 24894 3932
rect 24958 3868 25100 3932
rect 25164 3868 25180 3932
rect 25244 3868 25260 3932
rect 25324 3868 25340 3932
rect 25404 3868 25420 3932
rect 25484 3868 25500 3932
rect 25564 3868 25706 3932
rect 25770 3868 25786 3932
rect 25850 3868 25866 3932
rect 25930 3868 25946 3932
rect 26010 3868 26026 3932
rect 26090 3868 26106 3932
rect 26170 3868 26312 3932
rect 26376 3868 26392 3932
rect 26456 3868 26472 3932
rect 26536 3868 26552 3932
rect 26616 3868 26632 3932
rect 26696 3868 26712 3932
rect 26776 3868 26918 3932
rect 26982 3868 26998 3932
rect 27062 3868 27078 3932
rect 27142 3868 27158 3932
rect 27222 3868 27238 3932
rect 27302 3868 27318 3932
rect 27382 3868 27524 3932
rect 27588 3868 27604 3932
rect 27668 3868 27684 3932
rect 27748 3868 27764 3932
rect 27828 3868 27844 3932
rect 27908 3868 27924 3932
rect 27988 3868 28130 3932
rect 28194 3868 28210 3932
rect 28274 3868 28290 3932
rect 28354 3868 28370 3932
rect 28434 3868 28450 3932
rect 28514 3868 28530 3932
rect 28594 3868 28736 3932
rect 28800 3868 28816 3932
rect 28880 3868 28896 3932
rect 28960 3868 28976 3932
rect 29040 3868 29056 3932
rect 29120 3868 29136 3932
rect 29200 3868 29342 3932
rect 29406 3868 29422 3932
rect 29486 3868 29502 3932
rect 29566 3868 29582 3932
rect 29646 3868 29662 3932
rect 29726 3868 29742 3932
rect 29806 3868 29948 3932
rect 30012 3868 30028 3932
rect 30092 3868 30108 3932
rect 30172 3868 30188 3932
rect 30252 3868 30268 3932
rect 30332 3868 30348 3932
rect 30412 3868 30554 3932
rect 30618 3868 30634 3932
rect 30698 3868 30714 3932
rect 30778 3868 30794 3932
rect 30858 3868 30874 3932
rect 30938 3868 30954 3932
rect 31018 3868 31160 3932
rect 31224 3868 31240 3932
rect 31304 3868 31320 3932
rect 31384 3868 31400 3932
rect 31464 3868 31480 3932
rect 31544 3868 31560 3932
rect 31624 3868 31766 3932
rect 31830 3868 31846 3932
rect 31910 3868 31926 3932
rect 31990 3868 32006 3932
rect 32070 3868 32086 3932
rect 32150 3868 32166 3932
rect 32230 3868 32372 3932
rect 32436 3868 32452 3932
rect 32516 3868 32532 3932
rect 32596 3868 32612 3932
rect 32676 3868 32692 3932
rect 32756 3868 32772 3932
rect 32836 3868 32978 3932
rect 33042 3868 33058 3932
rect 33122 3868 33138 3932
rect 33202 3868 33218 3932
rect 33282 3868 33298 3932
rect 33362 3868 33378 3932
rect 33442 3868 33584 3932
rect 33648 3868 33664 3932
rect 33728 3868 33744 3932
rect 33808 3868 33824 3932
rect 33888 3868 33904 3932
rect 33968 3868 33984 3932
rect 34048 3868 34190 3932
rect 34254 3868 34270 3932
rect 34334 3868 34350 3932
rect 34414 3868 34430 3932
rect 34494 3868 34510 3932
rect 34574 3868 34590 3932
rect 34654 3868 34796 3932
rect 34860 3868 34876 3932
rect 34940 3868 34956 3932
rect 35020 3868 35036 3932
rect 35100 3868 35116 3932
rect 35180 3868 35196 3932
rect 35260 3868 35402 3932
rect 35466 3868 35482 3932
rect 35546 3868 35562 3932
rect 35626 3868 35642 3932
rect 35706 3868 35722 3932
rect 35786 3868 35802 3932
rect 35866 3868 36008 3932
rect 36072 3868 36088 3932
rect 36152 3868 36168 3932
rect 36232 3868 36248 3932
rect 36312 3868 36328 3932
rect 36392 3868 36408 3932
rect 36472 3868 36614 3932
rect 36678 3868 36694 3932
rect 36758 3868 36774 3932
rect 36838 3868 36854 3932
rect 36918 3868 36934 3932
rect 36998 3868 37014 3932
rect 37078 3868 37220 3932
rect 37284 3868 37300 3932
rect 37364 3868 37380 3932
rect 37444 3868 37460 3932
rect 37524 3868 37540 3932
rect 37604 3868 37620 3932
rect 37684 3868 37826 3932
rect 37890 3868 37906 3932
rect 37970 3868 37986 3932
rect 38050 3868 38066 3932
rect 38130 3868 38146 3932
rect 38210 3868 38226 3932
rect 38290 3868 38432 3932
rect 38496 3868 38512 3932
rect 38576 3868 38592 3932
rect 38656 3868 38672 3932
rect 38736 3868 38752 3932
rect 38816 3868 38832 3932
rect 38896 3868 39038 3932
rect 39102 3868 39118 3932
rect 39182 3868 39198 3932
rect 39262 3868 39278 3932
rect 39342 3868 39358 3932
rect 39422 3868 39438 3932
rect 39502 3868 39606 3932
rect 20148 3866 39606 3868
rect 20148 3712 20214 3866
rect 20148 3648 20149 3712
rect 20213 3648 20214 3712
rect 20148 3632 20214 3648
rect 20148 3568 20149 3632
rect 20213 3568 20214 3632
rect 20148 3552 20214 3568
rect 20148 3488 20149 3552
rect 20213 3488 20214 3552
rect 20148 3472 20214 3488
rect 20148 3408 20149 3472
rect 20213 3408 20214 3472
rect 20148 3392 20214 3408
rect 20148 3328 20149 3392
rect 20213 3328 20214 3392
rect 20148 3312 20214 3328
rect 20148 3248 20149 3312
rect 20213 3248 20214 3312
rect 20148 3232 20214 3248
rect 20148 3168 20149 3232
rect 20213 3168 20214 3232
rect 20148 3152 20214 3168
rect 20148 3088 20149 3152
rect 20213 3088 20214 3152
rect 20148 3072 20214 3088
rect 20148 3008 20149 3072
rect 20213 3008 20214 3072
rect 20148 2992 20214 3008
rect 20148 2928 20149 2992
rect 20213 2928 20214 2992
rect 20148 2838 20214 2928
rect 20274 2834 20334 3866
rect 20394 2774 20454 3804
rect 20514 2834 20574 3866
rect 20634 2774 20694 3804
rect 20754 3712 20820 3866
rect 20754 3648 20755 3712
rect 20819 3648 20820 3712
rect 20754 3632 20820 3648
rect 20754 3568 20755 3632
rect 20819 3568 20820 3632
rect 20754 3552 20820 3568
rect 20754 3488 20755 3552
rect 20819 3488 20820 3552
rect 20754 3472 20820 3488
rect 20754 3408 20755 3472
rect 20819 3408 20820 3472
rect 20754 3392 20820 3408
rect 20754 3328 20755 3392
rect 20819 3328 20820 3392
rect 20754 3312 20820 3328
rect 20754 3248 20755 3312
rect 20819 3248 20820 3312
rect 20754 3232 20820 3248
rect 20754 3168 20755 3232
rect 20819 3168 20820 3232
rect 20754 3152 20820 3168
rect 20754 3088 20755 3152
rect 20819 3088 20820 3152
rect 20754 3072 20820 3088
rect 20754 3008 20755 3072
rect 20819 3008 20820 3072
rect 20754 2992 20820 3008
rect 20754 2928 20755 2992
rect 20819 2928 20820 2992
rect 20754 2838 20820 2928
rect 20880 2834 20940 3866
rect 21000 2774 21060 3804
rect 21120 2834 21180 3866
rect 21240 2774 21300 3804
rect 21360 3712 21426 3866
rect 21360 3648 21361 3712
rect 21425 3648 21426 3712
rect 21360 3632 21426 3648
rect 21360 3568 21361 3632
rect 21425 3568 21426 3632
rect 21360 3552 21426 3568
rect 21360 3488 21361 3552
rect 21425 3488 21426 3552
rect 21360 3472 21426 3488
rect 21360 3408 21361 3472
rect 21425 3408 21426 3472
rect 21360 3392 21426 3408
rect 21360 3328 21361 3392
rect 21425 3328 21426 3392
rect 21360 3312 21426 3328
rect 21360 3248 21361 3312
rect 21425 3248 21426 3312
rect 21360 3232 21426 3248
rect 21360 3168 21361 3232
rect 21425 3168 21426 3232
rect 21360 3152 21426 3168
rect 21360 3088 21361 3152
rect 21425 3088 21426 3152
rect 21360 3072 21426 3088
rect 21360 3008 21361 3072
rect 21425 3008 21426 3072
rect 21360 2992 21426 3008
rect 21360 2928 21361 2992
rect 21425 2928 21426 2992
rect 21360 2838 21426 2928
rect 21486 2834 21546 3866
rect 21606 2774 21666 3804
rect 21726 2834 21786 3866
rect 21846 2774 21906 3804
rect 21966 3712 22032 3866
rect 21966 3648 21967 3712
rect 22031 3648 22032 3712
rect 21966 3632 22032 3648
rect 21966 3568 21967 3632
rect 22031 3568 22032 3632
rect 21966 3552 22032 3568
rect 21966 3488 21967 3552
rect 22031 3488 22032 3552
rect 21966 3472 22032 3488
rect 21966 3408 21967 3472
rect 22031 3408 22032 3472
rect 21966 3392 22032 3408
rect 21966 3328 21967 3392
rect 22031 3328 22032 3392
rect 21966 3312 22032 3328
rect 21966 3248 21967 3312
rect 22031 3248 22032 3312
rect 21966 3232 22032 3248
rect 21966 3168 21967 3232
rect 22031 3168 22032 3232
rect 21966 3152 22032 3168
rect 21966 3088 21967 3152
rect 22031 3088 22032 3152
rect 21966 3072 22032 3088
rect 21966 3008 21967 3072
rect 22031 3008 22032 3072
rect 21966 2992 22032 3008
rect 21966 2928 21967 2992
rect 22031 2928 22032 2992
rect 21966 2838 22032 2928
rect 22092 2834 22152 3866
rect 22212 2774 22272 3804
rect 22332 2834 22392 3866
rect 22452 2774 22512 3804
rect 22572 3712 22638 3866
rect 22572 3648 22573 3712
rect 22637 3648 22638 3712
rect 22572 3632 22638 3648
rect 22572 3568 22573 3632
rect 22637 3568 22638 3632
rect 22572 3552 22638 3568
rect 22572 3488 22573 3552
rect 22637 3488 22638 3552
rect 22572 3472 22638 3488
rect 22572 3408 22573 3472
rect 22637 3408 22638 3472
rect 22572 3392 22638 3408
rect 22572 3328 22573 3392
rect 22637 3328 22638 3392
rect 22572 3312 22638 3328
rect 22572 3248 22573 3312
rect 22637 3248 22638 3312
rect 22572 3232 22638 3248
rect 22572 3168 22573 3232
rect 22637 3168 22638 3232
rect 22572 3152 22638 3168
rect 22572 3088 22573 3152
rect 22637 3088 22638 3152
rect 22572 3072 22638 3088
rect 22572 3008 22573 3072
rect 22637 3008 22638 3072
rect 22572 2992 22638 3008
rect 22572 2928 22573 2992
rect 22637 2928 22638 2992
rect 22572 2838 22638 2928
rect 22698 2834 22758 3866
rect 22818 2774 22878 3804
rect 22938 2834 22998 3866
rect 23058 2774 23118 3804
rect 23178 3712 23244 3866
rect 23178 3648 23179 3712
rect 23243 3648 23244 3712
rect 23178 3632 23244 3648
rect 23178 3568 23179 3632
rect 23243 3568 23244 3632
rect 23178 3552 23244 3568
rect 23178 3488 23179 3552
rect 23243 3488 23244 3552
rect 23178 3472 23244 3488
rect 23178 3408 23179 3472
rect 23243 3408 23244 3472
rect 23178 3392 23244 3408
rect 23178 3328 23179 3392
rect 23243 3328 23244 3392
rect 23178 3312 23244 3328
rect 23178 3248 23179 3312
rect 23243 3248 23244 3312
rect 23178 3232 23244 3248
rect 23178 3168 23179 3232
rect 23243 3168 23244 3232
rect 23178 3152 23244 3168
rect 23178 3088 23179 3152
rect 23243 3088 23244 3152
rect 23178 3072 23244 3088
rect 23178 3008 23179 3072
rect 23243 3008 23244 3072
rect 23178 2992 23244 3008
rect 23178 2928 23179 2992
rect 23243 2928 23244 2992
rect 23178 2838 23244 2928
rect 23304 2834 23364 3866
rect 23424 2774 23484 3804
rect 23544 2834 23604 3866
rect 23664 2774 23724 3804
rect 23784 3712 23850 3866
rect 23784 3648 23785 3712
rect 23849 3648 23850 3712
rect 23784 3632 23850 3648
rect 23784 3568 23785 3632
rect 23849 3568 23850 3632
rect 23784 3552 23850 3568
rect 23784 3488 23785 3552
rect 23849 3488 23850 3552
rect 23784 3472 23850 3488
rect 23784 3408 23785 3472
rect 23849 3408 23850 3472
rect 23784 3392 23850 3408
rect 23784 3328 23785 3392
rect 23849 3328 23850 3392
rect 23784 3312 23850 3328
rect 23784 3248 23785 3312
rect 23849 3248 23850 3312
rect 23784 3232 23850 3248
rect 23784 3168 23785 3232
rect 23849 3168 23850 3232
rect 23784 3152 23850 3168
rect 23784 3088 23785 3152
rect 23849 3088 23850 3152
rect 23784 3072 23850 3088
rect 23784 3008 23785 3072
rect 23849 3008 23850 3072
rect 23784 2992 23850 3008
rect 23784 2928 23785 2992
rect 23849 2928 23850 2992
rect 23784 2838 23850 2928
rect 23910 2834 23970 3866
rect 24030 2774 24090 3804
rect 24150 2834 24210 3866
rect 24270 2774 24330 3804
rect 24390 3712 24456 3866
rect 24390 3648 24391 3712
rect 24455 3648 24456 3712
rect 24390 3632 24456 3648
rect 24390 3568 24391 3632
rect 24455 3568 24456 3632
rect 24390 3552 24456 3568
rect 24390 3488 24391 3552
rect 24455 3488 24456 3552
rect 24390 3472 24456 3488
rect 24390 3408 24391 3472
rect 24455 3408 24456 3472
rect 24390 3392 24456 3408
rect 24390 3328 24391 3392
rect 24455 3328 24456 3392
rect 24390 3312 24456 3328
rect 24390 3248 24391 3312
rect 24455 3248 24456 3312
rect 24390 3232 24456 3248
rect 24390 3168 24391 3232
rect 24455 3168 24456 3232
rect 24390 3152 24456 3168
rect 24390 3088 24391 3152
rect 24455 3088 24456 3152
rect 24390 3072 24456 3088
rect 24390 3008 24391 3072
rect 24455 3008 24456 3072
rect 24390 2992 24456 3008
rect 24390 2928 24391 2992
rect 24455 2928 24456 2992
rect 24390 2838 24456 2928
rect 24516 2834 24576 3866
rect 24636 2774 24696 3804
rect 24756 2834 24816 3866
rect 24876 2774 24936 3804
rect 24996 3712 25062 3866
rect 24996 3648 24997 3712
rect 25061 3648 25062 3712
rect 24996 3632 25062 3648
rect 24996 3568 24997 3632
rect 25061 3568 25062 3632
rect 24996 3552 25062 3568
rect 24996 3488 24997 3552
rect 25061 3488 25062 3552
rect 24996 3472 25062 3488
rect 24996 3408 24997 3472
rect 25061 3408 25062 3472
rect 24996 3392 25062 3408
rect 24996 3328 24997 3392
rect 25061 3328 25062 3392
rect 24996 3312 25062 3328
rect 24996 3248 24997 3312
rect 25061 3248 25062 3312
rect 24996 3232 25062 3248
rect 24996 3168 24997 3232
rect 25061 3168 25062 3232
rect 24996 3152 25062 3168
rect 24996 3088 24997 3152
rect 25061 3088 25062 3152
rect 24996 3072 25062 3088
rect 24996 3008 24997 3072
rect 25061 3008 25062 3072
rect 24996 2992 25062 3008
rect 24996 2928 24997 2992
rect 25061 2928 25062 2992
rect 24996 2838 25062 2928
rect 25122 2834 25182 3866
rect 25242 2774 25302 3804
rect 25362 2834 25422 3866
rect 25482 2774 25542 3804
rect 25602 3712 25668 3866
rect 25602 3648 25603 3712
rect 25667 3648 25668 3712
rect 25602 3632 25668 3648
rect 25602 3568 25603 3632
rect 25667 3568 25668 3632
rect 25602 3552 25668 3568
rect 25602 3488 25603 3552
rect 25667 3488 25668 3552
rect 25602 3472 25668 3488
rect 25602 3408 25603 3472
rect 25667 3408 25668 3472
rect 25602 3392 25668 3408
rect 25602 3328 25603 3392
rect 25667 3328 25668 3392
rect 25602 3312 25668 3328
rect 25602 3248 25603 3312
rect 25667 3248 25668 3312
rect 25602 3232 25668 3248
rect 25602 3168 25603 3232
rect 25667 3168 25668 3232
rect 25602 3152 25668 3168
rect 25602 3088 25603 3152
rect 25667 3088 25668 3152
rect 25602 3072 25668 3088
rect 25602 3008 25603 3072
rect 25667 3008 25668 3072
rect 25602 2992 25668 3008
rect 25602 2928 25603 2992
rect 25667 2928 25668 2992
rect 25602 2838 25668 2928
rect 25728 2834 25788 3866
rect 25848 2774 25908 3804
rect 25968 2834 26028 3866
rect 26088 2774 26148 3804
rect 26208 3712 26274 3866
rect 26208 3648 26209 3712
rect 26273 3648 26274 3712
rect 26208 3632 26274 3648
rect 26208 3568 26209 3632
rect 26273 3568 26274 3632
rect 26208 3552 26274 3568
rect 26208 3488 26209 3552
rect 26273 3488 26274 3552
rect 26208 3472 26274 3488
rect 26208 3408 26209 3472
rect 26273 3408 26274 3472
rect 26208 3392 26274 3408
rect 26208 3328 26209 3392
rect 26273 3328 26274 3392
rect 26208 3312 26274 3328
rect 26208 3248 26209 3312
rect 26273 3248 26274 3312
rect 26208 3232 26274 3248
rect 26208 3168 26209 3232
rect 26273 3168 26274 3232
rect 26208 3152 26274 3168
rect 26208 3088 26209 3152
rect 26273 3088 26274 3152
rect 26208 3072 26274 3088
rect 26208 3008 26209 3072
rect 26273 3008 26274 3072
rect 26208 2992 26274 3008
rect 26208 2928 26209 2992
rect 26273 2928 26274 2992
rect 26208 2838 26274 2928
rect 26334 2834 26394 3866
rect 26454 2774 26514 3804
rect 26574 2834 26634 3866
rect 26694 2774 26754 3804
rect 26814 3712 26880 3866
rect 26814 3648 26815 3712
rect 26879 3648 26880 3712
rect 26814 3632 26880 3648
rect 26814 3568 26815 3632
rect 26879 3568 26880 3632
rect 26814 3552 26880 3568
rect 26814 3488 26815 3552
rect 26879 3488 26880 3552
rect 26814 3472 26880 3488
rect 26814 3408 26815 3472
rect 26879 3408 26880 3472
rect 26814 3392 26880 3408
rect 26814 3328 26815 3392
rect 26879 3328 26880 3392
rect 26814 3312 26880 3328
rect 26814 3248 26815 3312
rect 26879 3248 26880 3312
rect 26814 3232 26880 3248
rect 26814 3168 26815 3232
rect 26879 3168 26880 3232
rect 26814 3152 26880 3168
rect 26814 3088 26815 3152
rect 26879 3088 26880 3152
rect 26814 3072 26880 3088
rect 26814 3008 26815 3072
rect 26879 3008 26880 3072
rect 26814 2992 26880 3008
rect 26814 2928 26815 2992
rect 26879 2928 26880 2992
rect 26814 2838 26880 2928
rect 26940 2834 27000 3866
rect 27060 2774 27120 3804
rect 27180 2834 27240 3866
rect 27300 2774 27360 3804
rect 27420 3712 27486 3866
rect 27420 3648 27421 3712
rect 27485 3648 27486 3712
rect 27420 3632 27486 3648
rect 27420 3568 27421 3632
rect 27485 3568 27486 3632
rect 27420 3552 27486 3568
rect 27420 3488 27421 3552
rect 27485 3488 27486 3552
rect 27420 3472 27486 3488
rect 27420 3408 27421 3472
rect 27485 3408 27486 3472
rect 27420 3392 27486 3408
rect 27420 3328 27421 3392
rect 27485 3328 27486 3392
rect 27420 3312 27486 3328
rect 27420 3248 27421 3312
rect 27485 3248 27486 3312
rect 27420 3232 27486 3248
rect 27420 3168 27421 3232
rect 27485 3168 27486 3232
rect 27420 3152 27486 3168
rect 27420 3088 27421 3152
rect 27485 3088 27486 3152
rect 27420 3072 27486 3088
rect 27420 3008 27421 3072
rect 27485 3008 27486 3072
rect 27420 2992 27486 3008
rect 27420 2928 27421 2992
rect 27485 2928 27486 2992
rect 27420 2838 27486 2928
rect 27546 2834 27606 3866
rect 27666 2774 27726 3804
rect 27786 2834 27846 3866
rect 27906 2774 27966 3804
rect 28026 3712 28092 3866
rect 28026 3648 28027 3712
rect 28091 3648 28092 3712
rect 28026 3632 28092 3648
rect 28026 3568 28027 3632
rect 28091 3568 28092 3632
rect 28026 3552 28092 3568
rect 28026 3488 28027 3552
rect 28091 3488 28092 3552
rect 28026 3472 28092 3488
rect 28026 3408 28027 3472
rect 28091 3408 28092 3472
rect 28026 3392 28092 3408
rect 28026 3328 28027 3392
rect 28091 3328 28092 3392
rect 28026 3312 28092 3328
rect 28026 3248 28027 3312
rect 28091 3248 28092 3312
rect 28026 3232 28092 3248
rect 28026 3168 28027 3232
rect 28091 3168 28092 3232
rect 28026 3152 28092 3168
rect 28026 3088 28027 3152
rect 28091 3088 28092 3152
rect 28026 3072 28092 3088
rect 28026 3008 28027 3072
rect 28091 3008 28092 3072
rect 28026 2992 28092 3008
rect 28026 2928 28027 2992
rect 28091 2928 28092 2992
rect 28026 2838 28092 2928
rect 28152 2834 28212 3866
rect 28272 2774 28332 3804
rect 28392 2834 28452 3866
rect 28512 2774 28572 3804
rect 28632 3712 28698 3866
rect 28632 3648 28633 3712
rect 28697 3648 28698 3712
rect 28632 3632 28698 3648
rect 28632 3568 28633 3632
rect 28697 3568 28698 3632
rect 28632 3552 28698 3568
rect 28632 3488 28633 3552
rect 28697 3488 28698 3552
rect 28632 3472 28698 3488
rect 28632 3408 28633 3472
rect 28697 3408 28698 3472
rect 28632 3392 28698 3408
rect 28632 3328 28633 3392
rect 28697 3328 28698 3392
rect 28632 3312 28698 3328
rect 28632 3248 28633 3312
rect 28697 3248 28698 3312
rect 28632 3232 28698 3248
rect 28632 3168 28633 3232
rect 28697 3168 28698 3232
rect 28632 3152 28698 3168
rect 28632 3088 28633 3152
rect 28697 3088 28698 3152
rect 28632 3072 28698 3088
rect 28632 3008 28633 3072
rect 28697 3008 28698 3072
rect 28632 2992 28698 3008
rect 28632 2928 28633 2992
rect 28697 2928 28698 2992
rect 28632 2838 28698 2928
rect 28758 2834 28818 3866
rect 28878 2774 28938 3804
rect 28998 2834 29058 3866
rect 29118 2774 29178 3804
rect 29238 3712 29304 3866
rect 29238 3648 29239 3712
rect 29303 3648 29304 3712
rect 29238 3632 29304 3648
rect 29238 3568 29239 3632
rect 29303 3568 29304 3632
rect 29238 3552 29304 3568
rect 29238 3488 29239 3552
rect 29303 3488 29304 3552
rect 29238 3472 29304 3488
rect 29238 3408 29239 3472
rect 29303 3408 29304 3472
rect 29238 3392 29304 3408
rect 29238 3328 29239 3392
rect 29303 3328 29304 3392
rect 29238 3312 29304 3328
rect 29238 3248 29239 3312
rect 29303 3248 29304 3312
rect 29238 3232 29304 3248
rect 29238 3168 29239 3232
rect 29303 3168 29304 3232
rect 29238 3152 29304 3168
rect 29238 3088 29239 3152
rect 29303 3088 29304 3152
rect 29238 3072 29304 3088
rect 29238 3008 29239 3072
rect 29303 3008 29304 3072
rect 29238 2992 29304 3008
rect 29238 2928 29239 2992
rect 29303 2928 29304 2992
rect 29238 2838 29304 2928
rect 29364 2834 29424 3866
rect 29484 2774 29544 3804
rect 29604 2834 29664 3866
rect 29724 2774 29784 3804
rect 29844 3712 29910 3866
rect 29844 3648 29845 3712
rect 29909 3648 29910 3712
rect 29844 3632 29910 3648
rect 29844 3568 29845 3632
rect 29909 3568 29910 3632
rect 29844 3552 29910 3568
rect 29844 3488 29845 3552
rect 29909 3488 29910 3552
rect 29844 3472 29910 3488
rect 29844 3408 29845 3472
rect 29909 3408 29910 3472
rect 29844 3392 29910 3408
rect 29844 3328 29845 3392
rect 29909 3328 29910 3392
rect 29844 3312 29910 3328
rect 29844 3248 29845 3312
rect 29909 3248 29910 3312
rect 29844 3232 29910 3248
rect 29844 3168 29845 3232
rect 29909 3168 29910 3232
rect 29844 3152 29910 3168
rect 29844 3088 29845 3152
rect 29909 3088 29910 3152
rect 29844 3072 29910 3088
rect 29844 3008 29845 3072
rect 29909 3008 29910 3072
rect 29844 2992 29910 3008
rect 29844 2928 29845 2992
rect 29909 2928 29910 2992
rect 29844 2838 29910 2928
rect 29970 2834 30030 3866
rect 30090 2774 30150 3804
rect 30210 2834 30270 3866
rect 30330 2774 30390 3804
rect 30450 3712 30516 3866
rect 30450 3648 30451 3712
rect 30515 3648 30516 3712
rect 30450 3632 30516 3648
rect 30450 3568 30451 3632
rect 30515 3568 30516 3632
rect 30450 3552 30516 3568
rect 30450 3488 30451 3552
rect 30515 3488 30516 3552
rect 30450 3472 30516 3488
rect 30450 3408 30451 3472
rect 30515 3408 30516 3472
rect 30450 3392 30516 3408
rect 30450 3328 30451 3392
rect 30515 3328 30516 3392
rect 30450 3312 30516 3328
rect 30450 3248 30451 3312
rect 30515 3248 30516 3312
rect 30450 3232 30516 3248
rect 30450 3168 30451 3232
rect 30515 3168 30516 3232
rect 30450 3152 30516 3168
rect 30450 3088 30451 3152
rect 30515 3088 30516 3152
rect 30450 3072 30516 3088
rect 30450 3008 30451 3072
rect 30515 3008 30516 3072
rect 30450 2992 30516 3008
rect 30450 2928 30451 2992
rect 30515 2928 30516 2992
rect 30450 2838 30516 2928
rect 30576 2834 30636 3866
rect 30696 2774 30756 3804
rect 30816 2834 30876 3866
rect 30936 2774 30996 3804
rect 31056 3712 31122 3866
rect 31056 3648 31057 3712
rect 31121 3648 31122 3712
rect 31056 3632 31122 3648
rect 31056 3568 31057 3632
rect 31121 3568 31122 3632
rect 31056 3552 31122 3568
rect 31056 3488 31057 3552
rect 31121 3488 31122 3552
rect 31056 3472 31122 3488
rect 31056 3408 31057 3472
rect 31121 3408 31122 3472
rect 31056 3392 31122 3408
rect 31056 3328 31057 3392
rect 31121 3328 31122 3392
rect 31056 3312 31122 3328
rect 31056 3248 31057 3312
rect 31121 3248 31122 3312
rect 31056 3232 31122 3248
rect 31056 3168 31057 3232
rect 31121 3168 31122 3232
rect 31056 3152 31122 3168
rect 31056 3088 31057 3152
rect 31121 3088 31122 3152
rect 31056 3072 31122 3088
rect 31056 3008 31057 3072
rect 31121 3008 31122 3072
rect 31056 2992 31122 3008
rect 31056 2928 31057 2992
rect 31121 2928 31122 2992
rect 31056 2838 31122 2928
rect 31182 2834 31242 3866
rect 31302 2774 31362 3804
rect 31422 2834 31482 3866
rect 31542 2774 31602 3804
rect 31662 3712 31728 3866
rect 31662 3648 31663 3712
rect 31727 3648 31728 3712
rect 31662 3632 31728 3648
rect 31662 3568 31663 3632
rect 31727 3568 31728 3632
rect 31662 3552 31728 3568
rect 31662 3488 31663 3552
rect 31727 3488 31728 3552
rect 31662 3472 31728 3488
rect 31662 3408 31663 3472
rect 31727 3408 31728 3472
rect 31662 3392 31728 3408
rect 31662 3328 31663 3392
rect 31727 3328 31728 3392
rect 31662 3312 31728 3328
rect 31662 3248 31663 3312
rect 31727 3248 31728 3312
rect 31662 3232 31728 3248
rect 31662 3168 31663 3232
rect 31727 3168 31728 3232
rect 31662 3152 31728 3168
rect 31662 3088 31663 3152
rect 31727 3088 31728 3152
rect 31662 3072 31728 3088
rect 31662 3008 31663 3072
rect 31727 3008 31728 3072
rect 31662 2992 31728 3008
rect 31662 2928 31663 2992
rect 31727 2928 31728 2992
rect 31662 2838 31728 2928
rect 31788 2834 31848 3866
rect 31908 2774 31968 3804
rect 32028 2834 32088 3866
rect 32148 2774 32208 3804
rect 32268 3712 32334 3866
rect 32268 3648 32269 3712
rect 32333 3648 32334 3712
rect 32268 3632 32334 3648
rect 32268 3568 32269 3632
rect 32333 3568 32334 3632
rect 32268 3552 32334 3568
rect 32268 3488 32269 3552
rect 32333 3488 32334 3552
rect 32268 3472 32334 3488
rect 32268 3408 32269 3472
rect 32333 3408 32334 3472
rect 32268 3392 32334 3408
rect 32268 3328 32269 3392
rect 32333 3328 32334 3392
rect 32268 3312 32334 3328
rect 32268 3248 32269 3312
rect 32333 3248 32334 3312
rect 32268 3232 32334 3248
rect 32268 3168 32269 3232
rect 32333 3168 32334 3232
rect 32268 3152 32334 3168
rect 32268 3088 32269 3152
rect 32333 3088 32334 3152
rect 32268 3072 32334 3088
rect 32268 3008 32269 3072
rect 32333 3008 32334 3072
rect 32268 2992 32334 3008
rect 32268 2928 32269 2992
rect 32333 2928 32334 2992
rect 32268 2838 32334 2928
rect 32394 2834 32454 3866
rect 32514 2774 32574 3804
rect 32634 2834 32694 3866
rect 32754 2774 32814 3804
rect 32874 3712 32940 3866
rect 32874 3648 32875 3712
rect 32939 3648 32940 3712
rect 32874 3632 32940 3648
rect 32874 3568 32875 3632
rect 32939 3568 32940 3632
rect 32874 3552 32940 3568
rect 32874 3488 32875 3552
rect 32939 3488 32940 3552
rect 32874 3472 32940 3488
rect 32874 3408 32875 3472
rect 32939 3408 32940 3472
rect 32874 3392 32940 3408
rect 32874 3328 32875 3392
rect 32939 3328 32940 3392
rect 32874 3312 32940 3328
rect 32874 3248 32875 3312
rect 32939 3248 32940 3312
rect 32874 3232 32940 3248
rect 32874 3168 32875 3232
rect 32939 3168 32940 3232
rect 32874 3152 32940 3168
rect 32874 3088 32875 3152
rect 32939 3088 32940 3152
rect 32874 3072 32940 3088
rect 32874 3008 32875 3072
rect 32939 3008 32940 3072
rect 32874 2992 32940 3008
rect 32874 2928 32875 2992
rect 32939 2928 32940 2992
rect 32874 2838 32940 2928
rect 33000 2834 33060 3866
rect 33120 2774 33180 3804
rect 33240 2834 33300 3866
rect 33360 2774 33420 3804
rect 33480 3712 33546 3866
rect 33480 3648 33481 3712
rect 33545 3648 33546 3712
rect 33480 3632 33546 3648
rect 33480 3568 33481 3632
rect 33545 3568 33546 3632
rect 33480 3552 33546 3568
rect 33480 3488 33481 3552
rect 33545 3488 33546 3552
rect 33480 3472 33546 3488
rect 33480 3408 33481 3472
rect 33545 3408 33546 3472
rect 33480 3392 33546 3408
rect 33480 3328 33481 3392
rect 33545 3328 33546 3392
rect 33480 3312 33546 3328
rect 33480 3248 33481 3312
rect 33545 3248 33546 3312
rect 33480 3232 33546 3248
rect 33480 3168 33481 3232
rect 33545 3168 33546 3232
rect 33480 3152 33546 3168
rect 33480 3088 33481 3152
rect 33545 3088 33546 3152
rect 33480 3072 33546 3088
rect 33480 3008 33481 3072
rect 33545 3008 33546 3072
rect 33480 2992 33546 3008
rect 33480 2928 33481 2992
rect 33545 2928 33546 2992
rect 33480 2838 33546 2928
rect 33606 2834 33666 3866
rect 33726 2774 33786 3804
rect 33846 2834 33906 3866
rect 33966 2774 34026 3804
rect 34086 3712 34152 3866
rect 34086 3648 34087 3712
rect 34151 3648 34152 3712
rect 34086 3632 34152 3648
rect 34086 3568 34087 3632
rect 34151 3568 34152 3632
rect 34086 3552 34152 3568
rect 34086 3488 34087 3552
rect 34151 3488 34152 3552
rect 34086 3472 34152 3488
rect 34086 3408 34087 3472
rect 34151 3408 34152 3472
rect 34086 3392 34152 3408
rect 34086 3328 34087 3392
rect 34151 3328 34152 3392
rect 34086 3312 34152 3328
rect 34086 3248 34087 3312
rect 34151 3248 34152 3312
rect 34086 3232 34152 3248
rect 34086 3168 34087 3232
rect 34151 3168 34152 3232
rect 34086 3152 34152 3168
rect 34086 3088 34087 3152
rect 34151 3088 34152 3152
rect 34086 3072 34152 3088
rect 34086 3008 34087 3072
rect 34151 3008 34152 3072
rect 34086 2992 34152 3008
rect 34086 2928 34087 2992
rect 34151 2928 34152 2992
rect 34086 2838 34152 2928
rect 34212 2834 34272 3866
rect 34332 2774 34392 3804
rect 34452 2834 34512 3866
rect 34572 2774 34632 3804
rect 34692 3712 34758 3866
rect 34692 3648 34693 3712
rect 34757 3648 34758 3712
rect 34692 3632 34758 3648
rect 34692 3568 34693 3632
rect 34757 3568 34758 3632
rect 34692 3552 34758 3568
rect 34692 3488 34693 3552
rect 34757 3488 34758 3552
rect 34692 3472 34758 3488
rect 34692 3408 34693 3472
rect 34757 3408 34758 3472
rect 34692 3392 34758 3408
rect 34692 3328 34693 3392
rect 34757 3328 34758 3392
rect 34692 3312 34758 3328
rect 34692 3248 34693 3312
rect 34757 3248 34758 3312
rect 34692 3232 34758 3248
rect 34692 3168 34693 3232
rect 34757 3168 34758 3232
rect 34692 3152 34758 3168
rect 34692 3088 34693 3152
rect 34757 3088 34758 3152
rect 34692 3072 34758 3088
rect 34692 3008 34693 3072
rect 34757 3008 34758 3072
rect 34692 2992 34758 3008
rect 34692 2928 34693 2992
rect 34757 2928 34758 2992
rect 34692 2838 34758 2928
rect 34818 2834 34878 3866
rect 34938 2774 34998 3804
rect 35058 2834 35118 3866
rect 35178 2774 35238 3804
rect 35298 3712 35364 3866
rect 35298 3648 35299 3712
rect 35363 3648 35364 3712
rect 35298 3632 35364 3648
rect 35298 3568 35299 3632
rect 35363 3568 35364 3632
rect 35298 3552 35364 3568
rect 35298 3488 35299 3552
rect 35363 3488 35364 3552
rect 35298 3472 35364 3488
rect 35298 3408 35299 3472
rect 35363 3408 35364 3472
rect 35298 3392 35364 3408
rect 35298 3328 35299 3392
rect 35363 3328 35364 3392
rect 35298 3312 35364 3328
rect 35298 3248 35299 3312
rect 35363 3248 35364 3312
rect 35298 3232 35364 3248
rect 35298 3168 35299 3232
rect 35363 3168 35364 3232
rect 35298 3152 35364 3168
rect 35298 3088 35299 3152
rect 35363 3088 35364 3152
rect 35298 3072 35364 3088
rect 35298 3008 35299 3072
rect 35363 3008 35364 3072
rect 35298 2992 35364 3008
rect 35298 2928 35299 2992
rect 35363 2928 35364 2992
rect 35298 2838 35364 2928
rect 35424 2834 35484 3866
rect 35544 2774 35604 3804
rect 35664 2834 35724 3866
rect 35784 2774 35844 3804
rect 35904 3712 35970 3866
rect 35904 3648 35905 3712
rect 35969 3648 35970 3712
rect 35904 3632 35970 3648
rect 35904 3568 35905 3632
rect 35969 3568 35970 3632
rect 35904 3552 35970 3568
rect 35904 3488 35905 3552
rect 35969 3488 35970 3552
rect 35904 3472 35970 3488
rect 35904 3408 35905 3472
rect 35969 3408 35970 3472
rect 35904 3392 35970 3408
rect 35904 3328 35905 3392
rect 35969 3328 35970 3392
rect 35904 3312 35970 3328
rect 35904 3248 35905 3312
rect 35969 3248 35970 3312
rect 35904 3232 35970 3248
rect 35904 3168 35905 3232
rect 35969 3168 35970 3232
rect 35904 3152 35970 3168
rect 35904 3088 35905 3152
rect 35969 3088 35970 3152
rect 35904 3072 35970 3088
rect 35904 3008 35905 3072
rect 35969 3008 35970 3072
rect 35904 2992 35970 3008
rect 35904 2928 35905 2992
rect 35969 2928 35970 2992
rect 35904 2838 35970 2928
rect 36030 2834 36090 3866
rect 36150 2774 36210 3804
rect 36270 2834 36330 3866
rect 36390 2774 36450 3804
rect 36510 3712 36576 3866
rect 36510 3648 36511 3712
rect 36575 3648 36576 3712
rect 36510 3632 36576 3648
rect 36510 3568 36511 3632
rect 36575 3568 36576 3632
rect 36510 3552 36576 3568
rect 36510 3488 36511 3552
rect 36575 3488 36576 3552
rect 36510 3472 36576 3488
rect 36510 3408 36511 3472
rect 36575 3408 36576 3472
rect 36510 3392 36576 3408
rect 36510 3328 36511 3392
rect 36575 3328 36576 3392
rect 36510 3312 36576 3328
rect 36510 3248 36511 3312
rect 36575 3248 36576 3312
rect 36510 3232 36576 3248
rect 36510 3168 36511 3232
rect 36575 3168 36576 3232
rect 36510 3152 36576 3168
rect 36510 3088 36511 3152
rect 36575 3088 36576 3152
rect 36510 3072 36576 3088
rect 36510 3008 36511 3072
rect 36575 3008 36576 3072
rect 36510 2992 36576 3008
rect 36510 2928 36511 2992
rect 36575 2928 36576 2992
rect 36510 2838 36576 2928
rect 36636 2834 36696 3866
rect 36756 2774 36816 3804
rect 36876 2834 36936 3866
rect 36996 2774 37056 3804
rect 37116 3712 37182 3866
rect 37116 3648 37117 3712
rect 37181 3648 37182 3712
rect 37116 3632 37182 3648
rect 37116 3568 37117 3632
rect 37181 3568 37182 3632
rect 37116 3552 37182 3568
rect 37116 3488 37117 3552
rect 37181 3488 37182 3552
rect 37116 3472 37182 3488
rect 37116 3408 37117 3472
rect 37181 3408 37182 3472
rect 37116 3392 37182 3408
rect 37116 3328 37117 3392
rect 37181 3328 37182 3392
rect 37116 3312 37182 3328
rect 37116 3248 37117 3312
rect 37181 3248 37182 3312
rect 37116 3232 37182 3248
rect 37116 3168 37117 3232
rect 37181 3168 37182 3232
rect 37116 3152 37182 3168
rect 37116 3088 37117 3152
rect 37181 3088 37182 3152
rect 37116 3072 37182 3088
rect 37116 3008 37117 3072
rect 37181 3008 37182 3072
rect 37116 2992 37182 3008
rect 37116 2928 37117 2992
rect 37181 2928 37182 2992
rect 37116 2838 37182 2928
rect 37242 2834 37302 3866
rect 37362 2774 37422 3804
rect 37482 2834 37542 3866
rect 37602 2774 37662 3804
rect 37722 3712 37788 3866
rect 37722 3648 37723 3712
rect 37787 3648 37788 3712
rect 37722 3632 37788 3648
rect 37722 3568 37723 3632
rect 37787 3568 37788 3632
rect 37722 3552 37788 3568
rect 37722 3488 37723 3552
rect 37787 3488 37788 3552
rect 37722 3472 37788 3488
rect 37722 3408 37723 3472
rect 37787 3408 37788 3472
rect 37722 3392 37788 3408
rect 37722 3328 37723 3392
rect 37787 3328 37788 3392
rect 37722 3312 37788 3328
rect 37722 3248 37723 3312
rect 37787 3248 37788 3312
rect 37722 3232 37788 3248
rect 37722 3168 37723 3232
rect 37787 3168 37788 3232
rect 37722 3152 37788 3168
rect 37722 3088 37723 3152
rect 37787 3088 37788 3152
rect 37722 3072 37788 3088
rect 37722 3008 37723 3072
rect 37787 3008 37788 3072
rect 37722 2992 37788 3008
rect 37722 2928 37723 2992
rect 37787 2928 37788 2992
rect 37722 2838 37788 2928
rect 37848 2834 37908 3866
rect 37968 2774 38028 3804
rect 38088 2834 38148 3866
rect 38208 2774 38268 3804
rect 38328 3712 38394 3866
rect 38328 3648 38329 3712
rect 38393 3648 38394 3712
rect 38328 3632 38394 3648
rect 38328 3568 38329 3632
rect 38393 3568 38394 3632
rect 38328 3552 38394 3568
rect 38328 3488 38329 3552
rect 38393 3488 38394 3552
rect 38328 3472 38394 3488
rect 38328 3408 38329 3472
rect 38393 3408 38394 3472
rect 38328 3392 38394 3408
rect 38328 3328 38329 3392
rect 38393 3328 38394 3392
rect 38328 3312 38394 3328
rect 38328 3248 38329 3312
rect 38393 3248 38394 3312
rect 38328 3232 38394 3248
rect 38328 3168 38329 3232
rect 38393 3168 38394 3232
rect 38328 3152 38394 3168
rect 38328 3088 38329 3152
rect 38393 3088 38394 3152
rect 38328 3072 38394 3088
rect 38328 3008 38329 3072
rect 38393 3008 38394 3072
rect 38328 2992 38394 3008
rect 38328 2928 38329 2992
rect 38393 2928 38394 2992
rect 38328 2838 38394 2928
rect 38454 2834 38514 3866
rect 38574 2774 38634 3804
rect 38694 2834 38754 3866
rect 38814 2774 38874 3804
rect 38934 3712 39000 3866
rect 38934 3648 38935 3712
rect 38999 3648 39000 3712
rect 38934 3632 39000 3648
rect 38934 3568 38935 3632
rect 38999 3568 39000 3632
rect 38934 3552 39000 3568
rect 38934 3488 38935 3552
rect 38999 3488 39000 3552
rect 38934 3472 39000 3488
rect 38934 3408 38935 3472
rect 38999 3408 39000 3472
rect 38934 3392 39000 3408
rect 38934 3328 38935 3392
rect 38999 3328 39000 3392
rect 38934 3312 39000 3328
rect 38934 3248 38935 3312
rect 38999 3248 39000 3312
rect 38934 3232 39000 3248
rect 38934 3168 38935 3232
rect 38999 3168 39000 3232
rect 38934 3152 39000 3168
rect 38934 3088 38935 3152
rect 38999 3088 39000 3152
rect 38934 3072 39000 3088
rect 38934 3008 38935 3072
rect 38999 3008 39000 3072
rect 38934 2992 39000 3008
rect 38934 2928 38935 2992
rect 38999 2928 39000 2992
rect 38934 2838 39000 2928
rect 39060 2834 39120 3866
rect 39180 2774 39240 3804
rect 39300 2834 39360 3866
rect 39420 2774 39480 3804
rect 39540 3712 39606 3866
rect 39540 3648 39541 3712
rect 39605 3648 39606 3712
rect 39540 3632 39606 3648
rect 39540 3568 39541 3632
rect 39605 3568 39606 3632
rect 39540 3552 39606 3568
rect 39540 3488 39541 3552
rect 39605 3488 39606 3552
rect 39540 3472 39606 3488
rect 39540 3408 39541 3472
rect 39605 3408 39606 3472
rect 39540 3392 39606 3408
rect 39540 3328 39541 3392
rect 39605 3328 39606 3392
rect 39540 3312 39606 3328
rect 39540 3248 39541 3312
rect 39605 3248 39606 3312
rect 39540 3232 39606 3248
rect 39540 3168 39541 3232
rect 39605 3168 39606 3232
rect 39540 3152 39606 3168
rect 39540 3088 39541 3152
rect 39605 3088 39606 3152
rect 39540 3072 39606 3088
rect 39540 3008 39541 3072
rect 39605 3008 39606 3072
rect 39540 2992 39606 3008
rect 39540 2928 39541 2992
rect 39605 2928 39606 2992
rect 39540 2838 39606 2928
rect -459 2772 213 2774
rect -459 2708 -355 2772
rect -291 2708 -275 2772
rect -211 2708 -195 2772
rect -131 2708 -115 2772
rect -51 2708 -35 2772
rect 29 2708 45 2772
rect 109 2708 213 2772
rect -459 2706 213 2708
rect 524 2772 1027 2774
rect 524 2708 539 2772
rect 603 2708 619 2772
rect 683 2708 699 2772
rect 763 2708 779 2772
rect 843 2708 859 2772
rect 923 2708 1027 2772
rect -93 2606 -33 2615
rect -459 2604 213 2606
rect -459 2540 -355 2604
rect -291 2540 -275 2604
rect -211 2540 -195 2604
rect -131 2540 -115 2604
rect -51 2540 -35 2604
rect 29 2540 45 2604
rect 109 2540 213 2604
rect -459 2538 213 2540
rect 524 2706 1027 2708
rect 1267 2772 1717 2774
rect 1954 2772 2545 2774
rect 1267 2708 1371 2772
rect 1435 2708 1451 2772
rect 1515 2708 1531 2772
rect 1595 2708 1611 2772
rect 1675 2708 1691 2772
rect 1954 2708 1977 2772
rect 2041 2708 2057 2772
rect 2121 2708 2137 2772
rect 2201 2708 2217 2772
rect 2281 2708 2297 2772
rect 2361 2708 2377 2772
rect 2441 2708 2545 2772
rect 1267 2706 1717 2708
rect 524 2604 1027 2606
rect 524 2540 539 2604
rect 603 2540 619 2604
rect 683 2540 699 2604
rect 763 2540 779 2604
rect 843 2540 859 2604
rect 923 2540 1027 2604
rect 524 2538 1027 2540
rect 1267 2604 1717 2606
rect 1954 2706 2545 2708
rect 2801 2772 3301 2774
rect 3538 2772 5291 2774
rect 2801 2708 2905 2772
rect 2969 2708 2985 2772
rect 3049 2708 3065 2772
rect 3129 2708 3145 2772
rect 3209 2708 3225 2772
rect 3289 2708 3301 2772
rect 3575 2708 3591 2772
rect 3655 2708 3671 2772
rect 3735 2708 3751 2772
rect 3815 2708 3831 2772
rect 3895 2708 3911 2772
rect 3975 2708 4117 2772
rect 4181 2708 4197 2772
rect 4261 2708 4277 2772
rect 4341 2708 4357 2772
rect 4421 2708 4437 2772
rect 4501 2708 4517 2772
rect 4581 2708 4723 2772
rect 4787 2708 4803 2772
rect 4867 2708 4883 2772
rect 4947 2708 4963 2772
rect 5027 2708 5043 2772
rect 5107 2708 5123 2772
rect 5187 2708 5291 2772
rect 2801 2706 3301 2708
rect 1954 2604 2545 2606
rect 1267 2540 1371 2604
rect 1435 2540 1451 2604
rect 1515 2540 1531 2604
rect 1595 2540 1611 2604
rect 1675 2540 1691 2604
rect 1954 2540 1977 2604
rect 2041 2540 2057 2604
rect 2121 2540 2137 2604
rect 2201 2540 2217 2604
rect 2281 2540 2297 2604
rect 2361 2540 2377 2604
rect 2441 2540 2545 2604
rect 1267 2538 1717 2540
rect 1954 2538 2545 2540
rect 2801 2604 3301 2606
rect 3538 2706 5291 2708
rect 5352 2706 5394 2774
rect 5631 2772 10266 2774
rect 5680 2708 5696 2772
rect 5760 2708 5776 2772
rect 5840 2708 5856 2772
rect 5920 2708 6062 2772
rect 6126 2708 6142 2772
rect 6206 2708 6222 2772
rect 6286 2708 6302 2772
rect 6366 2708 6382 2772
rect 6446 2708 6462 2772
rect 6526 2708 6668 2772
rect 6732 2708 6748 2772
rect 6812 2708 6828 2772
rect 6892 2708 6908 2772
rect 6972 2708 6988 2772
rect 7052 2708 7068 2772
rect 7132 2708 7274 2772
rect 7338 2708 7354 2772
rect 7418 2708 7434 2772
rect 7498 2708 7514 2772
rect 7578 2708 7594 2772
rect 7658 2708 7674 2772
rect 7738 2708 7880 2772
rect 7944 2708 7960 2772
rect 8024 2708 8040 2772
rect 8104 2708 8120 2772
rect 8184 2708 8200 2772
rect 8264 2708 8280 2772
rect 8344 2708 8486 2772
rect 8550 2708 8566 2772
rect 8630 2708 8646 2772
rect 8710 2708 8726 2772
rect 8790 2708 8806 2772
rect 8870 2708 8886 2772
rect 8950 2708 9092 2772
rect 9156 2708 9172 2772
rect 9236 2708 9252 2772
rect 9316 2708 9332 2772
rect 9396 2708 9412 2772
rect 9476 2708 9492 2772
rect 9556 2708 9698 2772
rect 9762 2708 9778 2772
rect 9842 2708 9858 2772
rect 9922 2708 9938 2772
rect 10002 2708 10018 2772
rect 10082 2708 10098 2772
rect 10162 2708 10266 2772
rect 3538 2604 5291 2606
rect 2801 2540 2905 2604
rect 2969 2540 2985 2604
rect 3049 2540 3065 2604
rect 3129 2540 3145 2604
rect 3209 2540 3225 2604
rect 3289 2540 3301 2604
rect 3575 2540 3591 2604
rect 3655 2540 3671 2604
rect 3735 2540 3751 2604
rect 3815 2540 3831 2604
rect 3895 2540 3911 2604
rect 3975 2540 4117 2604
rect 4181 2540 4197 2604
rect 4261 2540 4277 2604
rect 4341 2540 4357 2604
rect 4421 2540 4437 2604
rect 4501 2540 4517 2604
rect 4581 2540 4723 2604
rect 4787 2540 4803 2604
rect 4867 2540 4883 2604
rect 4947 2540 4963 2604
rect 5027 2540 5043 2604
rect 5107 2540 5123 2604
rect 5187 2540 5291 2604
rect 2801 2538 3301 2540
rect 3538 2538 5291 2540
rect 5352 2538 5394 2606
rect 5631 2706 10266 2708
rect 10326 2706 10368 2774
rect 10605 2772 20088 2774
rect 10654 2708 10670 2772
rect 10734 2708 10750 2772
rect 10814 2708 10830 2772
rect 10894 2708 11036 2772
rect 11100 2708 11116 2772
rect 11180 2708 11196 2772
rect 11260 2708 11276 2772
rect 11340 2708 11356 2772
rect 11420 2708 11436 2772
rect 11500 2708 11642 2772
rect 11706 2708 11722 2772
rect 11786 2708 11802 2772
rect 11866 2708 11882 2772
rect 11946 2708 11962 2772
rect 12026 2708 12042 2772
rect 12106 2708 12248 2772
rect 12312 2708 12328 2772
rect 12392 2708 12408 2772
rect 12472 2708 12488 2772
rect 12552 2708 12568 2772
rect 12632 2708 12648 2772
rect 12712 2708 12854 2772
rect 12918 2708 12934 2772
rect 12998 2708 13014 2772
rect 13078 2708 13094 2772
rect 13158 2708 13174 2772
rect 13238 2708 13254 2772
rect 13318 2708 13460 2772
rect 13524 2708 13540 2772
rect 13604 2708 13620 2772
rect 13684 2708 13700 2772
rect 13764 2708 13780 2772
rect 13844 2708 13860 2772
rect 13924 2708 14066 2772
rect 14130 2708 14146 2772
rect 14210 2708 14226 2772
rect 14290 2708 14306 2772
rect 14370 2708 14386 2772
rect 14450 2708 14466 2772
rect 14530 2708 14672 2772
rect 14736 2708 14752 2772
rect 14816 2708 14832 2772
rect 14896 2708 14912 2772
rect 14976 2708 14992 2772
rect 15056 2708 15072 2772
rect 15136 2708 15278 2772
rect 15342 2708 15358 2772
rect 15422 2708 15438 2772
rect 15502 2708 15518 2772
rect 15582 2708 15598 2772
rect 15662 2708 15678 2772
rect 15742 2708 15884 2772
rect 15948 2708 15964 2772
rect 16028 2708 16044 2772
rect 16108 2708 16124 2772
rect 16188 2708 16204 2772
rect 16268 2708 16284 2772
rect 16348 2708 16490 2772
rect 16554 2708 16570 2772
rect 16634 2708 16650 2772
rect 16714 2708 16730 2772
rect 16794 2708 16810 2772
rect 16874 2708 16890 2772
rect 16954 2708 17096 2772
rect 17160 2708 17176 2772
rect 17240 2708 17256 2772
rect 17320 2708 17336 2772
rect 17400 2708 17416 2772
rect 17480 2708 17496 2772
rect 17560 2708 17702 2772
rect 17766 2708 17782 2772
rect 17846 2708 17862 2772
rect 17926 2708 17942 2772
rect 18006 2708 18022 2772
rect 18086 2708 18102 2772
rect 18166 2708 18308 2772
rect 18372 2708 18388 2772
rect 18452 2708 18468 2772
rect 18532 2708 18548 2772
rect 18612 2708 18628 2772
rect 18692 2708 18708 2772
rect 18772 2708 18914 2772
rect 18978 2708 18994 2772
rect 19058 2708 19074 2772
rect 19138 2708 19154 2772
rect 19218 2708 19234 2772
rect 19298 2708 19314 2772
rect 19378 2708 19520 2772
rect 19584 2708 19600 2772
rect 19664 2708 19680 2772
rect 19744 2708 19760 2772
rect 19824 2708 19840 2772
rect 19904 2708 19920 2772
rect 19984 2708 20088 2772
rect 5631 2604 10266 2606
rect 5680 2540 5696 2604
rect 5760 2540 5776 2604
rect 5840 2540 5856 2604
rect 5920 2540 6062 2604
rect 6126 2540 6142 2604
rect 6206 2540 6222 2604
rect 6286 2540 6302 2604
rect 6366 2540 6382 2604
rect 6446 2540 6462 2604
rect 6526 2540 6668 2604
rect 6732 2540 6748 2604
rect 6812 2540 6828 2604
rect 6892 2540 6908 2604
rect 6972 2540 6988 2604
rect 7052 2540 7068 2604
rect 7132 2540 7274 2604
rect 7338 2540 7354 2604
rect 7418 2540 7434 2604
rect 7498 2540 7514 2604
rect 7578 2540 7594 2604
rect 7658 2540 7674 2604
rect 7738 2540 7880 2604
rect 7944 2540 7960 2604
rect 8024 2540 8040 2604
rect 8104 2540 8120 2604
rect 8184 2540 8200 2604
rect 8264 2540 8280 2604
rect 8344 2540 8486 2604
rect 8550 2540 8566 2604
rect 8630 2540 8646 2604
rect 8710 2540 8726 2604
rect 8790 2540 8806 2604
rect 8870 2540 8886 2604
rect 8950 2540 9092 2604
rect 9156 2540 9172 2604
rect 9236 2540 9252 2604
rect 9316 2540 9332 2604
rect 9396 2540 9412 2604
rect 9476 2540 9492 2604
rect 9556 2540 9698 2604
rect 9762 2540 9778 2604
rect 9842 2540 9858 2604
rect 9922 2540 9938 2604
rect 10002 2540 10018 2604
rect 10082 2540 10098 2604
rect 10162 2540 10266 2604
rect 5631 2538 10266 2540
rect 10326 2538 10368 2606
rect 10605 2706 20088 2708
rect 20148 2772 39298 2774
rect 20148 2708 20252 2772
rect 20316 2708 20332 2772
rect 20396 2708 20412 2772
rect 20476 2708 20492 2772
rect 20556 2708 20572 2772
rect 20636 2708 20652 2772
rect 20716 2708 20858 2772
rect 20922 2708 20938 2772
rect 21002 2708 21018 2772
rect 21082 2708 21098 2772
rect 21162 2708 21178 2772
rect 21242 2708 21258 2772
rect 21322 2708 21464 2772
rect 21528 2708 21544 2772
rect 21608 2708 21624 2772
rect 21688 2708 21704 2772
rect 21768 2708 21784 2772
rect 21848 2708 21864 2772
rect 21928 2708 22070 2772
rect 22134 2708 22150 2772
rect 22214 2708 22230 2772
rect 22294 2708 22310 2772
rect 22374 2708 22390 2772
rect 22454 2708 22470 2772
rect 22534 2708 22676 2772
rect 22740 2708 22756 2772
rect 22820 2708 22836 2772
rect 22900 2708 22916 2772
rect 22980 2708 22996 2772
rect 23060 2708 23076 2772
rect 23140 2708 23282 2772
rect 23346 2708 23362 2772
rect 23426 2708 23442 2772
rect 23506 2708 23522 2772
rect 23586 2708 23602 2772
rect 23666 2708 23682 2772
rect 23746 2708 23888 2772
rect 23952 2708 23968 2772
rect 24032 2708 24048 2772
rect 24112 2708 24128 2772
rect 24192 2708 24208 2772
rect 24272 2708 24288 2772
rect 24352 2708 24494 2772
rect 24558 2708 24574 2772
rect 24638 2708 24654 2772
rect 24718 2708 24734 2772
rect 24798 2708 24814 2772
rect 24878 2708 24894 2772
rect 24958 2708 25100 2772
rect 25164 2708 25180 2772
rect 25244 2708 25260 2772
rect 25324 2708 25340 2772
rect 25404 2708 25420 2772
rect 25484 2708 25500 2772
rect 25564 2708 25706 2772
rect 25770 2708 25786 2772
rect 25850 2708 25866 2772
rect 25930 2708 25946 2772
rect 26010 2708 26026 2772
rect 26090 2708 26106 2772
rect 26170 2708 26312 2772
rect 26376 2708 26392 2772
rect 26456 2708 26472 2772
rect 26536 2708 26552 2772
rect 26616 2708 26632 2772
rect 26696 2708 26712 2772
rect 26776 2708 26918 2772
rect 26982 2708 26998 2772
rect 27062 2708 27078 2772
rect 27142 2708 27158 2772
rect 27222 2708 27238 2772
rect 27302 2708 27318 2772
rect 27382 2708 27524 2772
rect 27588 2708 27604 2772
rect 27668 2708 27684 2772
rect 27748 2708 27764 2772
rect 27828 2708 27844 2772
rect 27908 2708 27924 2772
rect 27988 2708 28130 2772
rect 28194 2708 28210 2772
rect 28274 2708 28290 2772
rect 28354 2708 28370 2772
rect 28434 2708 28450 2772
rect 28514 2708 28530 2772
rect 28594 2708 28736 2772
rect 28800 2708 28816 2772
rect 28880 2708 28896 2772
rect 28960 2708 28976 2772
rect 29040 2708 29056 2772
rect 29120 2708 29136 2772
rect 29200 2708 29342 2772
rect 29406 2708 29422 2772
rect 29486 2708 29502 2772
rect 29566 2708 29582 2772
rect 29646 2708 29662 2772
rect 29726 2708 29742 2772
rect 29806 2708 29948 2772
rect 30012 2708 30028 2772
rect 30092 2708 30108 2772
rect 30172 2708 30188 2772
rect 30252 2708 30268 2772
rect 30332 2708 30348 2772
rect 30412 2708 30554 2772
rect 30618 2708 30634 2772
rect 30698 2708 30714 2772
rect 30778 2708 30794 2772
rect 30858 2708 30874 2772
rect 30938 2708 30954 2772
rect 31018 2708 31160 2772
rect 31224 2708 31240 2772
rect 31304 2708 31320 2772
rect 31384 2708 31400 2772
rect 31464 2708 31480 2772
rect 31544 2708 31560 2772
rect 31624 2708 31766 2772
rect 31830 2708 31846 2772
rect 31910 2708 31926 2772
rect 31990 2708 32006 2772
rect 32070 2708 32086 2772
rect 32150 2708 32166 2772
rect 32230 2708 32372 2772
rect 32436 2708 32452 2772
rect 32516 2708 32532 2772
rect 32596 2708 32612 2772
rect 32676 2708 32692 2772
rect 32756 2708 32772 2772
rect 32836 2708 32978 2772
rect 33042 2708 33058 2772
rect 33122 2708 33138 2772
rect 33202 2708 33218 2772
rect 33282 2708 33298 2772
rect 33362 2708 33378 2772
rect 33442 2708 33584 2772
rect 33648 2708 33664 2772
rect 33728 2708 33744 2772
rect 33808 2708 33824 2772
rect 33888 2708 33904 2772
rect 33968 2708 33984 2772
rect 34048 2708 34190 2772
rect 34254 2708 34270 2772
rect 34334 2708 34350 2772
rect 34414 2708 34430 2772
rect 34494 2708 34510 2772
rect 34574 2708 34590 2772
rect 34654 2708 34796 2772
rect 34860 2708 34876 2772
rect 34940 2708 34956 2772
rect 35020 2708 35036 2772
rect 35100 2708 35116 2772
rect 35180 2708 35196 2772
rect 35260 2708 35402 2772
rect 35466 2708 35482 2772
rect 35546 2708 35562 2772
rect 35626 2708 35642 2772
rect 35706 2708 35722 2772
rect 35786 2708 35802 2772
rect 35866 2708 36008 2772
rect 36072 2708 36088 2772
rect 36152 2708 36168 2772
rect 36232 2708 36248 2772
rect 36312 2708 36328 2772
rect 36392 2708 36408 2772
rect 36472 2708 36614 2772
rect 36678 2708 36694 2772
rect 36758 2708 36774 2772
rect 36838 2708 36854 2772
rect 36918 2708 36934 2772
rect 36998 2708 37014 2772
rect 37078 2708 37220 2772
rect 37284 2708 37300 2772
rect 37364 2708 37380 2772
rect 37444 2708 37460 2772
rect 37524 2708 37540 2772
rect 37604 2708 37620 2772
rect 37684 2708 37826 2772
rect 37890 2708 37906 2772
rect 37970 2708 37986 2772
rect 38050 2708 38066 2772
rect 38130 2708 38146 2772
rect 38210 2708 38226 2772
rect 38290 2708 38432 2772
rect 38496 2708 38512 2772
rect 38576 2708 38592 2772
rect 38656 2708 38672 2772
rect 38736 2708 38752 2772
rect 38816 2708 38832 2772
rect 38896 2708 39038 2772
rect 39102 2708 39118 2772
rect 39182 2708 39198 2772
rect 39262 2708 39278 2772
rect 20148 2706 39298 2708
rect 10605 2604 20088 2606
rect 10654 2540 10670 2604
rect 10734 2540 10750 2604
rect 10814 2540 10830 2604
rect 10894 2540 11036 2604
rect 11100 2540 11116 2604
rect 11180 2540 11196 2604
rect 11260 2540 11276 2604
rect 11340 2540 11356 2604
rect 11420 2540 11436 2604
rect 11500 2540 11642 2604
rect 11706 2540 11722 2604
rect 11786 2540 11802 2604
rect 11866 2540 11882 2604
rect 11946 2540 11962 2604
rect 12026 2540 12042 2604
rect 12106 2540 12248 2604
rect 12312 2540 12328 2604
rect 12392 2540 12408 2604
rect 12472 2540 12488 2604
rect 12552 2540 12568 2604
rect 12632 2540 12648 2604
rect 12712 2540 12854 2604
rect 12918 2540 12934 2604
rect 12998 2540 13014 2604
rect 13078 2540 13094 2604
rect 13158 2540 13174 2604
rect 13238 2540 13254 2604
rect 13318 2540 13460 2604
rect 13524 2540 13540 2604
rect 13604 2540 13620 2604
rect 13684 2540 13700 2604
rect 13764 2540 13780 2604
rect 13844 2540 13860 2604
rect 13924 2540 14066 2604
rect 14130 2540 14146 2604
rect 14210 2540 14226 2604
rect 14290 2540 14306 2604
rect 14370 2540 14386 2604
rect 14450 2540 14466 2604
rect 14530 2540 14672 2604
rect 14736 2540 14752 2604
rect 14816 2540 14832 2604
rect 14896 2540 14912 2604
rect 14976 2540 14992 2604
rect 15056 2540 15072 2604
rect 15136 2540 15278 2604
rect 15342 2540 15358 2604
rect 15422 2540 15438 2604
rect 15502 2540 15518 2604
rect 15582 2540 15598 2604
rect 15662 2540 15678 2604
rect 15742 2540 15884 2604
rect 15948 2540 15964 2604
rect 16028 2540 16044 2604
rect 16108 2540 16124 2604
rect 16188 2540 16204 2604
rect 16268 2540 16284 2604
rect 16348 2540 16490 2604
rect 16554 2540 16570 2604
rect 16634 2540 16650 2604
rect 16714 2540 16730 2604
rect 16794 2540 16810 2604
rect 16874 2540 16890 2604
rect 16954 2540 17096 2604
rect 17160 2540 17176 2604
rect 17240 2540 17256 2604
rect 17320 2540 17336 2604
rect 17400 2540 17416 2604
rect 17480 2540 17496 2604
rect 17560 2540 17702 2604
rect 17766 2540 17782 2604
rect 17846 2540 17862 2604
rect 17926 2540 17942 2604
rect 18006 2540 18022 2604
rect 18086 2540 18102 2604
rect 18166 2540 18308 2604
rect 18372 2540 18388 2604
rect 18452 2540 18468 2604
rect 18532 2540 18548 2604
rect 18612 2540 18628 2604
rect 18692 2540 18708 2604
rect 18772 2540 18914 2604
rect 18978 2540 18994 2604
rect 19058 2540 19074 2604
rect 19138 2540 19154 2604
rect 19218 2540 19234 2604
rect 19298 2540 19314 2604
rect 19378 2540 19520 2604
rect 19584 2540 19600 2604
rect 19664 2540 19680 2604
rect 19744 2540 19760 2604
rect 19824 2540 19840 2604
rect 19904 2540 19920 2604
rect 19984 2540 20088 2604
rect 10605 2538 20088 2540
rect 20148 2604 39298 2606
rect 39534 2706 39606 2774
rect 20148 2540 20252 2604
rect 20316 2540 20332 2604
rect 20396 2540 20412 2604
rect 20476 2540 20492 2604
rect 20556 2540 20572 2604
rect 20636 2540 20652 2604
rect 20716 2540 20858 2604
rect 20922 2540 20938 2604
rect 21002 2540 21018 2604
rect 21082 2540 21098 2604
rect 21162 2540 21178 2604
rect 21242 2540 21258 2604
rect 21322 2540 21464 2604
rect 21528 2540 21544 2604
rect 21608 2540 21624 2604
rect 21688 2540 21704 2604
rect 21768 2540 21784 2604
rect 21848 2540 21864 2604
rect 21928 2540 22070 2604
rect 22134 2540 22150 2604
rect 22214 2540 22230 2604
rect 22294 2540 22310 2604
rect 22374 2540 22390 2604
rect 22454 2540 22470 2604
rect 22534 2540 22676 2604
rect 22740 2540 22756 2604
rect 22820 2540 22836 2604
rect 22900 2540 22916 2604
rect 22980 2540 22996 2604
rect 23060 2540 23076 2604
rect 23140 2540 23282 2604
rect 23346 2540 23362 2604
rect 23426 2540 23442 2604
rect 23506 2540 23522 2604
rect 23586 2540 23602 2604
rect 23666 2540 23682 2604
rect 23746 2540 23888 2604
rect 23952 2540 23968 2604
rect 24032 2540 24048 2604
rect 24112 2540 24128 2604
rect 24192 2540 24208 2604
rect 24272 2540 24288 2604
rect 24352 2540 24494 2604
rect 24558 2540 24574 2604
rect 24638 2540 24654 2604
rect 24718 2540 24734 2604
rect 24798 2540 24814 2604
rect 24878 2540 24894 2604
rect 24958 2540 25100 2604
rect 25164 2540 25180 2604
rect 25244 2540 25260 2604
rect 25324 2540 25340 2604
rect 25404 2540 25420 2604
rect 25484 2540 25500 2604
rect 25564 2540 25706 2604
rect 25770 2540 25786 2604
rect 25850 2540 25866 2604
rect 25930 2540 25946 2604
rect 26010 2540 26026 2604
rect 26090 2540 26106 2604
rect 26170 2540 26312 2604
rect 26376 2540 26392 2604
rect 26456 2540 26472 2604
rect 26536 2540 26552 2604
rect 26616 2540 26632 2604
rect 26696 2540 26712 2604
rect 26776 2540 26918 2604
rect 26982 2540 26998 2604
rect 27062 2540 27078 2604
rect 27142 2540 27158 2604
rect 27222 2540 27238 2604
rect 27302 2540 27318 2604
rect 27382 2540 27524 2604
rect 27588 2540 27604 2604
rect 27668 2540 27684 2604
rect 27748 2540 27764 2604
rect 27828 2540 27844 2604
rect 27908 2540 27924 2604
rect 27988 2540 28130 2604
rect 28194 2540 28210 2604
rect 28274 2540 28290 2604
rect 28354 2540 28370 2604
rect 28434 2540 28450 2604
rect 28514 2540 28530 2604
rect 28594 2540 28736 2604
rect 28800 2540 28816 2604
rect 28880 2540 28896 2604
rect 28960 2540 28976 2604
rect 29040 2540 29056 2604
rect 29120 2540 29136 2604
rect 29200 2540 29342 2604
rect 29406 2540 29422 2604
rect 29486 2540 29502 2604
rect 29566 2540 29582 2604
rect 29646 2540 29662 2604
rect 29726 2540 29742 2604
rect 29806 2540 29948 2604
rect 30012 2540 30028 2604
rect 30092 2540 30108 2604
rect 30172 2540 30188 2604
rect 30252 2540 30268 2604
rect 30332 2540 30348 2604
rect 30412 2540 30554 2604
rect 30618 2540 30634 2604
rect 30698 2540 30714 2604
rect 30778 2540 30794 2604
rect 30858 2540 30874 2604
rect 30938 2540 30954 2604
rect 31018 2540 31160 2604
rect 31224 2540 31240 2604
rect 31304 2540 31320 2604
rect 31384 2540 31400 2604
rect 31464 2540 31480 2604
rect 31544 2540 31560 2604
rect 31624 2540 31766 2604
rect 31830 2540 31846 2604
rect 31910 2540 31926 2604
rect 31990 2540 32006 2604
rect 32070 2540 32086 2604
rect 32150 2540 32166 2604
rect 32230 2540 32372 2604
rect 32436 2540 32452 2604
rect 32516 2540 32532 2604
rect 32596 2540 32612 2604
rect 32676 2540 32692 2604
rect 32756 2540 32772 2604
rect 32836 2540 32978 2604
rect 33042 2540 33058 2604
rect 33122 2540 33138 2604
rect 33202 2540 33218 2604
rect 33282 2540 33298 2604
rect 33362 2540 33378 2604
rect 33442 2540 33584 2604
rect 33648 2540 33664 2604
rect 33728 2540 33744 2604
rect 33808 2540 33824 2604
rect 33888 2540 33904 2604
rect 33968 2540 33984 2604
rect 34048 2540 34190 2604
rect 34254 2540 34270 2604
rect 34334 2540 34350 2604
rect 34414 2540 34430 2604
rect 34494 2540 34510 2604
rect 34574 2540 34590 2604
rect 34654 2540 34796 2604
rect 34860 2540 34876 2604
rect 34940 2540 34956 2604
rect 35020 2540 35036 2604
rect 35100 2540 35116 2604
rect 35180 2540 35196 2604
rect 35260 2540 35402 2604
rect 35466 2540 35482 2604
rect 35546 2540 35562 2604
rect 35626 2540 35642 2604
rect 35706 2540 35722 2604
rect 35786 2540 35802 2604
rect 35866 2540 36008 2604
rect 36072 2540 36088 2604
rect 36152 2540 36168 2604
rect 36232 2540 36248 2604
rect 36312 2540 36328 2604
rect 36392 2540 36408 2604
rect 36472 2540 36614 2604
rect 36678 2540 36694 2604
rect 36758 2540 36774 2604
rect 36838 2540 36854 2604
rect 36918 2540 36934 2604
rect 36998 2540 37014 2604
rect 37078 2540 37220 2604
rect 37284 2540 37300 2604
rect 37364 2540 37380 2604
rect 37444 2540 37460 2604
rect 37524 2540 37540 2604
rect 37604 2540 37620 2604
rect 37684 2540 37826 2604
rect 37890 2540 37906 2604
rect 37970 2540 37986 2604
rect 38050 2540 38066 2604
rect 38130 2540 38146 2604
rect 38210 2540 38226 2604
rect 38290 2540 38432 2604
rect 38496 2540 38512 2604
rect 38576 2540 38592 2604
rect 38656 2540 38672 2604
rect 38736 2540 38752 2604
rect 38816 2540 38832 2604
rect 38896 2540 39038 2604
rect 39102 2540 39118 2604
rect 39182 2540 39198 2604
rect 39262 2540 39278 2604
rect 20148 2538 39298 2540
rect 39534 2538 39606 2606
rect -459 2384 -393 2538
rect -459 2320 -458 2384
rect -394 2320 -393 2384
rect -459 2304 -393 2320
rect -459 2240 -458 2304
rect -394 2240 -393 2304
rect -459 2224 -393 2240
rect -459 2160 -458 2224
rect -394 2160 -393 2224
rect -459 2144 -393 2160
rect -459 2080 -458 2144
rect -394 2080 -393 2144
rect -459 2064 -393 2080
rect -459 2000 -458 2064
rect -394 2000 -393 2064
rect -459 1984 -393 2000
rect -459 1920 -458 1984
rect -394 1920 -393 1984
rect -459 1904 -393 1920
rect -459 1840 -458 1904
rect -394 1840 -393 1904
rect -459 1824 -393 1840
rect -459 1760 -458 1824
rect -394 1760 -393 1824
rect -459 1744 -393 1760
rect -459 1680 -458 1744
rect -394 1680 -393 1744
rect -459 1664 -393 1680
rect -459 1600 -458 1664
rect -394 1600 -393 1664
rect -459 1510 -393 1600
rect -333 1506 -273 2538
rect -213 1446 -153 2476
rect -93 1506 -33 2538
rect 27 1446 87 2476
rect 147 2384 213 2538
rect 147 2320 148 2384
rect 212 2320 213 2384
rect 147 2304 213 2320
rect 147 2240 148 2304
rect 212 2240 213 2304
rect 147 2224 213 2240
rect 147 2160 148 2224
rect 212 2160 213 2224
rect 147 2144 213 2160
rect 147 2080 148 2144
rect 212 2080 213 2144
rect 147 2064 213 2080
rect 147 2000 148 2064
rect 212 2000 213 2064
rect 147 1984 213 2000
rect 147 1920 148 1984
rect 212 1920 213 1984
rect 147 1904 213 1920
rect 147 1840 148 1904
rect 212 1840 213 1904
rect 147 1824 213 1840
rect 147 1760 148 1824
rect 212 1760 213 1824
rect 147 1744 213 1760
rect 147 1680 148 1744
rect 212 1680 213 1744
rect 147 1664 213 1680
rect 147 1600 148 1664
rect 212 1600 213 1664
rect 147 1510 213 1600
rect 355 2384 421 2474
rect 355 2320 356 2384
rect 420 2320 421 2384
rect 355 2304 421 2320
rect 355 2240 356 2304
rect 420 2240 421 2304
rect 355 2224 421 2240
rect 355 2160 356 2224
rect 420 2160 421 2224
rect 355 2144 421 2160
rect 355 2080 356 2144
rect 420 2080 421 2144
rect 355 2064 421 2080
rect 355 2000 356 2064
rect 420 2000 421 2064
rect 355 1984 421 2000
rect 355 1920 356 1984
rect 420 1920 421 1984
rect 355 1904 421 1920
rect 355 1840 356 1904
rect 420 1840 421 1904
rect 355 1824 421 1840
rect 355 1760 356 1824
rect 420 1760 421 1824
rect 355 1744 421 1760
rect 355 1680 356 1744
rect 420 1680 421 1744
rect 355 1664 421 1680
rect 355 1600 356 1664
rect 420 1600 421 1664
rect 355 1446 421 1600
rect 481 1508 541 2538
rect 601 1446 661 2478
rect 721 1508 781 2538
rect 841 1446 901 2478
rect 961 2465 1027 2474
rect 961 2401 962 2465
rect 1026 2401 1027 2465
rect 961 2384 1027 2401
rect 961 2320 962 2384
rect 1026 2320 1027 2384
rect 961 2304 1027 2320
rect 961 2240 962 2304
rect 1026 2240 1027 2304
rect 961 2224 1027 2240
rect 961 2160 962 2224
rect 1026 2160 1027 2224
rect 961 2144 1027 2160
rect 961 2080 962 2144
rect 1026 2080 1027 2144
rect 961 2064 1027 2080
rect 961 2000 962 2064
rect 1026 2000 1027 2064
rect 961 1984 1027 2000
rect 961 1920 962 1984
rect 1026 1920 1027 1984
rect 961 1904 1027 1920
rect 961 1840 962 1904
rect 1026 1840 1027 1904
rect 961 1824 1027 1840
rect 961 1760 962 1824
rect 1026 1760 1027 1824
rect 961 1744 1027 1760
rect 961 1680 962 1744
rect 1026 1680 1027 1744
rect 961 1664 1027 1680
rect 961 1600 962 1664
rect 1026 1600 1027 1664
rect 961 1446 1027 1600
rect -459 1444 213 1446
rect -459 1380 -355 1444
rect -291 1380 -275 1444
rect -211 1380 -195 1444
rect -131 1380 -115 1444
rect -51 1380 -35 1444
rect 29 1380 45 1444
rect 109 1380 213 1444
rect -459 1378 213 1380
rect 355 1444 1027 1446
rect 355 1380 459 1444
rect 523 1380 539 1444
rect 603 1380 619 1444
rect 683 1380 699 1444
rect 763 1380 779 1444
rect 843 1380 859 1444
rect 923 1380 1027 1444
rect 355 1378 1027 1380
rect -459 1224 -393 1314
rect -459 1160 -458 1224
rect -394 1160 -393 1224
rect -459 1144 -393 1160
rect -459 1080 -458 1144
rect -394 1080 -393 1144
rect -459 1064 -393 1080
rect -459 1000 -458 1064
rect -394 1000 -393 1064
rect -459 984 -393 1000
rect -459 920 -458 984
rect -394 920 -393 984
rect -459 904 -393 920
rect -459 840 -458 904
rect -394 840 -393 904
rect -459 824 -393 840
rect -459 760 -458 824
rect -394 760 -393 824
rect -459 744 -393 760
rect -459 680 -458 744
rect -394 680 -393 744
rect -459 664 -393 680
rect -459 600 -458 664
rect -394 600 -393 664
rect -459 584 -393 600
rect -459 520 -458 584
rect -394 520 -393 584
rect -459 504 -393 520
rect -459 440 -458 504
rect -394 440 -393 504
rect -459 286 -393 440
rect -333 348 -273 1378
rect -213 286 -153 1318
rect -93 348 -33 1378
rect 27 286 87 1318
rect 147 1224 213 1314
rect 147 1160 148 1224
rect 212 1160 213 1224
rect 147 1144 213 1160
rect 147 1080 148 1144
rect 212 1080 213 1144
rect 147 1064 213 1080
rect 147 1000 148 1064
rect 212 1000 213 1064
rect 147 984 213 1000
rect 147 920 148 984
rect 212 920 213 984
rect 147 904 213 920
rect 147 840 148 904
rect 212 840 213 904
rect 147 824 213 840
rect 147 760 148 824
rect 212 760 213 824
rect 147 744 213 760
rect 147 680 148 744
rect 212 680 213 744
rect 147 664 213 680
rect 147 600 148 664
rect 212 600 213 664
rect 147 584 213 600
rect 147 520 148 584
rect 212 520 213 584
rect 147 504 213 520
rect 147 440 148 504
rect 212 440 213 504
rect 147 286 213 440
rect 355 1224 421 1378
rect 355 1160 356 1224
rect 420 1160 421 1224
rect 355 1144 421 1160
rect 355 1080 356 1144
rect 420 1080 421 1144
rect 355 1064 421 1080
rect 355 1000 356 1064
rect 420 1000 421 1064
rect 355 984 421 1000
rect 355 920 356 984
rect 420 920 421 984
rect 355 904 421 920
rect 355 840 356 904
rect 420 840 421 904
rect 355 824 421 840
rect 355 760 356 824
rect 420 760 421 824
rect 355 744 421 760
rect 355 680 356 744
rect 420 680 421 744
rect 355 664 421 680
rect 355 600 356 664
rect 420 600 421 664
rect 355 584 421 600
rect 355 520 356 584
rect 420 520 421 584
rect 355 504 421 520
rect 355 440 356 504
rect 420 440 421 504
rect 355 350 421 440
rect 481 346 541 1378
rect 601 286 661 1316
rect 721 346 781 1378
rect 841 286 901 1316
rect 961 1224 1027 1378
rect 961 1160 962 1224
rect 1026 1160 1027 1224
rect 961 1144 1027 1160
rect 961 1080 962 1144
rect 1026 1080 1027 1144
rect 961 1064 1027 1080
rect 961 1000 962 1064
rect 1026 1000 1027 1064
rect 961 984 1027 1000
rect 961 920 962 984
rect 1026 920 1027 984
rect 961 904 1027 920
rect 961 840 962 904
rect 1026 840 1027 904
rect 961 824 1027 840
rect 961 760 962 824
rect 1026 760 1027 824
rect 961 744 1027 760
rect 961 680 962 744
rect 1026 680 1027 744
rect 961 664 1027 680
rect 961 600 962 664
rect 1026 600 1027 664
rect 961 584 1027 600
rect 961 520 962 584
rect 1026 520 1027 584
rect 961 504 1027 520
rect 961 440 962 504
rect 1026 440 1027 504
rect 961 350 1027 440
rect 1267 2384 1333 2474
rect 1267 2320 1268 2384
rect 1332 2320 1333 2384
rect 1267 2304 1333 2320
rect 1267 2240 1268 2304
rect 1332 2240 1333 2304
rect 1267 2224 1333 2240
rect 1267 2160 1268 2224
rect 1332 2160 1333 2224
rect 1267 2144 1333 2160
rect 1267 2080 1268 2144
rect 1332 2080 1333 2144
rect 1267 2064 1333 2080
rect 1267 2000 1268 2064
rect 1332 2000 1333 2064
rect 1267 1984 1333 2000
rect 1267 1920 1268 1984
rect 1332 1920 1333 1984
rect 1267 1904 1333 1920
rect 1267 1840 1268 1904
rect 1332 1840 1333 1904
rect 1267 1824 1333 1840
rect 1267 1760 1268 1824
rect 1332 1760 1333 1824
rect 1267 1744 1333 1760
rect 1267 1680 1268 1744
rect 1332 1680 1333 1744
rect 1267 1664 1333 1680
rect 1267 1600 1268 1664
rect 1332 1600 1333 1664
rect 1267 1446 1333 1600
rect 1393 1508 1453 2538
rect 1513 1446 1573 2478
rect 1633 1508 1693 2538
rect 1753 1446 1813 2478
rect 1873 2384 1939 2474
rect 1873 2320 1874 2384
rect 1938 2320 1939 2384
rect 1873 2304 1939 2320
rect 1873 2240 1874 2304
rect 1938 2240 1939 2304
rect 1873 2224 1939 2240
rect 1873 2160 1874 2224
rect 1938 2160 1939 2224
rect 1873 2144 1939 2160
rect 1873 2080 1874 2144
rect 1938 2080 1939 2144
rect 1873 2064 1939 2080
rect 1873 2000 1874 2064
rect 1938 2000 1939 2064
rect 1873 1984 1939 2000
rect 1873 1920 1874 1984
rect 1938 1920 1939 1984
rect 1873 1904 1939 1920
rect 1873 1840 1874 1904
rect 1938 1840 1939 1904
rect 1873 1824 1939 1840
rect 1873 1760 1874 1824
rect 1938 1760 1939 1824
rect 1873 1744 1939 1760
rect 1873 1680 1874 1744
rect 1938 1680 1939 1744
rect 1873 1664 1939 1680
rect 1873 1600 1874 1664
rect 1938 1600 1939 1664
rect 1873 1446 1939 1600
rect 1999 1508 2059 2538
rect 2119 1446 2179 2478
rect 2239 1508 2299 2538
rect 2359 1446 2419 2478
rect 2479 2465 2545 2474
rect 2479 2401 2480 2465
rect 2544 2401 2545 2465
rect 2479 2384 2545 2401
rect 2479 2320 2480 2384
rect 2544 2320 2545 2384
rect 2479 2304 2545 2320
rect 2479 2240 2480 2304
rect 2544 2240 2545 2304
rect 2479 2224 2545 2240
rect 2479 2160 2480 2224
rect 2544 2160 2545 2224
rect 2479 2144 2545 2160
rect 2479 2080 2480 2144
rect 2544 2080 2545 2144
rect 2479 2064 2545 2080
rect 2479 2000 2480 2064
rect 2544 2000 2545 2064
rect 2479 1984 2545 2000
rect 2479 1920 2480 1984
rect 2544 1920 2545 1984
rect 2479 1904 2545 1920
rect 2479 1840 2480 1904
rect 2544 1840 2545 1904
rect 2479 1824 2545 1840
rect 2479 1760 2480 1824
rect 2544 1760 2545 1824
rect 2479 1744 2545 1760
rect 2479 1680 2480 1744
rect 2544 1680 2545 1744
rect 2479 1664 2545 1680
rect 2479 1600 2480 1664
rect 2544 1600 2545 1664
rect 2479 1446 2545 1600
rect 1267 1444 2545 1446
rect 1267 1380 1371 1444
rect 1435 1380 1451 1444
rect 1515 1380 1531 1444
rect 1595 1380 1611 1444
rect 1675 1380 1691 1444
rect 1755 1380 1771 1444
rect 1835 1380 1977 1444
rect 2041 1380 2057 1444
rect 2121 1380 2137 1444
rect 2201 1380 2217 1444
rect 2281 1380 2297 1444
rect 2361 1380 2377 1444
rect 2441 1380 2545 1444
rect 1267 1378 2545 1380
rect 1267 1224 1333 1378
rect 1267 1160 1268 1224
rect 1332 1160 1333 1224
rect 1267 1144 1333 1160
rect 1267 1080 1268 1144
rect 1332 1080 1333 1144
rect 1267 1064 1333 1080
rect 1267 1000 1268 1064
rect 1332 1000 1333 1064
rect 1267 984 1333 1000
rect 1267 920 1268 984
rect 1332 920 1333 984
rect 1267 904 1333 920
rect 1267 840 1268 904
rect 1332 840 1333 904
rect 1267 824 1333 840
rect 1267 760 1268 824
rect 1332 760 1333 824
rect 1267 744 1333 760
rect 1267 680 1268 744
rect 1332 680 1333 744
rect 1267 664 1333 680
rect 1267 600 1268 664
rect 1332 600 1333 664
rect 1267 584 1333 600
rect 1267 520 1268 584
rect 1332 520 1333 584
rect 1267 504 1333 520
rect 1267 440 1268 504
rect 1332 440 1333 504
rect 1267 350 1333 440
rect 1393 346 1453 1378
rect 1513 286 1573 1316
rect 1633 346 1693 1378
rect 1753 286 1813 1316
rect 1873 1224 1939 1378
rect 1873 1160 1874 1224
rect 1938 1160 1939 1224
rect 1873 1144 1939 1160
rect 1873 1080 1874 1144
rect 1938 1080 1939 1144
rect 1873 1064 1939 1080
rect 1873 1000 1874 1064
rect 1938 1000 1939 1064
rect 1873 984 1939 1000
rect 1873 920 1874 984
rect 1938 920 1939 984
rect 1873 904 1939 920
rect 1873 840 1874 904
rect 1938 840 1939 904
rect 1873 824 1939 840
rect 1873 760 1874 824
rect 1938 760 1939 824
rect 1873 744 1939 760
rect 1873 680 1874 744
rect 1938 680 1939 744
rect 1873 664 1939 680
rect 1873 600 1874 664
rect 1938 600 1939 664
rect 1873 584 1939 600
rect 1873 520 1874 584
rect 1938 520 1939 584
rect 1873 504 1939 520
rect 1873 440 1874 504
rect 1938 440 1939 504
rect 1873 350 1939 440
rect 1999 346 2059 1378
rect 2119 286 2179 1316
rect 2239 346 2299 1378
rect 2359 286 2419 1316
rect 2479 1224 2545 1378
rect 2479 1160 2480 1224
rect 2544 1160 2545 1224
rect 2479 1144 2545 1160
rect 2479 1080 2480 1144
rect 2544 1080 2545 1144
rect 2479 1064 2545 1080
rect 2479 1000 2480 1064
rect 2544 1000 2545 1064
rect 2479 984 2545 1000
rect 2479 920 2480 984
rect 2544 920 2545 984
rect 2479 904 2545 920
rect 2479 840 2480 904
rect 2544 840 2545 904
rect 2479 824 2545 840
rect 2479 760 2480 824
rect 2544 760 2545 824
rect 2479 744 2545 760
rect 2479 680 2480 744
rect 2544 680 2545 744
rect 2479 664 2545 680
rect 2479 600 2480 664
rect 2544 600 2545 664
rect 2479 584 2545 600
rect 2479 520 2480 584
rect 2544 520 2545 584
rect 2479 504 2545 520
rect 2479 440 2480 504
rect 2544 440 2545 504
rect 2479 350 2545 440
rect 2801 2384 2867 2474
rect 2801 2320 2802 2384
rect 2866 2320 2867 2384
rect 2801 2304 2867 2320
rect 2801 2240 2802 2304
rect 2866 2240 2867 2304
rect 2801 2224 2867 2240
rect 2801 2160 2802 2224
rect 2866 2160 2867 2224
rect 2801 2144 2867 2160
rect 2801 2080 2802 2144
rect 2866 2080 2867 2144
rect 2801 2064 2867 2080
rect 2801 2000 2802 2064
rect 2866 2000 2867 2064
rect 2801 1984 2867 2000
rect 2801 1920 2802 1984
rect 2866 1920 2867 1984
rect 2801 1904 2867 1920
rect 2801 1840 2802 1904
rect 2866 1840 2867 1904
rect 2801 1824 2867 1840
rect 2801 1760 2802 1824
rect 2866 1760 2867 1824
rect 2801 1744 2867 1760
rect 2801 1680 2802 1744
rect 2866 1680 2867 1744
rect 2801 1664 2867 1680
rect 2801 1600 2802 1664
rect 2866 1600 2867 1664
rect 2801 1446 2867 1600
rect 2927 1508 2987 2538
rect 3047 1446 3107 2478
rect 3167 1508 3227 2538
rect 3287 1446 3347 2478
rect 3407 2384 3473 2474
rect 3407 2320 3408 2384
rect 3472 2320 3473 2384
rect 3407 2304 3473 2320
rect 3407 2240 3408 2304
rect 3472 2240 3473 2304
rect 3407 2224 3473 2240
rect 3407 2160 3408 2224
rect 3472 2160 3473 2224
rect 3407 2144 3473 2160
rect 3407 2080 3408 2144
rect 3472 2080 3473 2144
rect 3407 2064 3473 2080
rect 3407 2000 3408 2064
rect 3472 2000 3473 2064
rect 3407 1984 3473 2000
rect 3407 1920 3408 1984
rect 3472 1920 3473 1984
rect 3407 1904 3473 1920
rect 3407 1840 3408 1904
rect 3472 1840 3473 1904
rect 3407 1824 3473 1840
rect 3407 1760 3408 1824
rect 3472 1760 3473 1824
rect 3407 1744 3473 1760
rect 3407 1680 3408 1744
rect 3472 1680 3473 1744
rect 3407 1664 3473 1680
rect 3407 1600 3408 1664
rect 3472 1600 3473 1664
rect 3407 1446 3473 1600
rect 3533 1508 3593 2538
rect 3653 1446 3713 2478
rect 3773 1508 3833 2538
rect 3893 1446 3953 2478
rect 4013 2384 4079 2474
rect 4013 2320 4014 2384
rect 4078 2320 4079 2384
rect 4013 2304 4079 2320
rect 4013 2240 4014 2304
rect 4078 2240 4079 2304
rect 4013 2224 4079 2240
rect 4013 2160 4014 2224
rect 4078 2160 4079 2224
rect 4013 2144 4079 2160
rect 4013 2080 4014 2144
rect 4078 2080 4079 2144
rect 4013 2064 4079 2080
rect 4013 2000 4014 2064
rect 4078 2000 4079 2064
rect 4013 1984 4079 2000
rect 4013 1920 4014 1984
rect 4078 1920 4079 1984
rect 4013 1904 4079 1920
rect 4013 1840 4014 1904
rect 4078 1840 4079 1904
rect 4013 1824 4079 1840
rect 4013 1760 4014 1824
rect 4078 1760 4079 1824
rect 4013 1744 4079 1760
rect 4013 1680 4014 1744
rect 4078 1680 4079 1744
rect 4013 1664 4079 1680
rect 4013 1600 4014 1664
rect 4078 1600 4079 1664
rect 4013 1446 4079 1600
rect 4139 1508 4199 2538
rect 4259 1446 4319 2478
rect 4379 1508 4439 2538
rect 4499 1446 4559 2478
rect 4619 2384 4685 2474
rect 4619 2320 4620 2384
rect 4684 2320 4685 2384
rect 4619 2304 4685 2320
rect 4619 2240 4620 2304
rect 4684 2240 4685 2304
rect 4619 2224 4685 2240
rect 4619 2160 4620 2224
rect 4684 2160 4685 2224
rect 4619 2144 4685 2160
rect 4619 2080 4620 2144
rect 4684 2080 4685 2144
rect 4619 2064 4685 2080
rect 4619 2000 4620 2064
rect 4684 2000 4685 2064
rect 4619 1984 4685 2000
rect 4619 1920 4620 1984
rect 4684 1920 4685 1984
rect 4619 1904 4685 1920
rect 4619 1840 4620 1904
rect 4684 1840 4685 1904
rect 4619 1824 4685 1840
rect 4619 1760 4620 1824
rect 4684 1760 4685 1824
rect 4619 1744 4685 1760
rect 4619 1680 4620 1744
rect 4684 1680 4685 1744
rect 4619 1664 4685 1680
rect 4619 1600 4620 1664
rect 4684 1600 4685 1664
rect 4619 1446 4685 1600
rect 4745 1508 4805 2538
rect 4865 1446 4925 2478
rect 4985 1508 5045 2538
rect 5105 1446 5165 2478
rect 5225 2384 5291 2474
rect 5225 2320 5226 2384
rect 5290 2320 5291 2384
rect 5225 2304 5291 2320
rect 5225 2240 5226 2304
rect 5290 2240 5291 2304
rect 5225 2224 5291 2240
rect 5225 2160 5226 2224
rect 5290 2160 5291 2224
rect 5225 2144 5291 2160
rect 5225 2080 5226 2144
rect 5290 2080 5291 2144
rect 5225 2064 5291 2080
rect 5225 2000 5226 2064
rect 5290 2000 5291 2064
rect 5225 1984 5291 2000
rect 5225 1920 5226 1984
rect 5290 1920 5291 1984
rect 5225 1904 5291 1920
rect 5225 1840 5226 1904
rect 5290 1840 5291 1904
rect 5225 1824 5291 1840
rect 5225 1760 5226 1824
rect 5290 1760 5291 1824
rect 5225 1744 5291 1760
rect 5225 1680 5226 1744
rect 5290 1680 5291 1744
rect 5225 1664 5291 1680
rect 5225 1600 5226 1664
rect 5290 1600 5291 1664
rect 5225 1446 5291 1600
rect 2801 1444 5291 1446
rect 2801 1380 2905 1444
rect 2969 1380 2985 1444
rect 3049 1380 3065 1444
rect 3129 1380 3145 1444
rect 3209 1380 3225 1444
rect 3289 1380 3305 1444
rect 3369 1380 3511 1444
rect 3575 1380 3591 1444
rect 3655 1380 3671 1444
rect 3735 1380 3751 1444
rect 3815 1380 3831 1444
rect 3895 1380 3911 1444
rect 3975 1380 4117 1444
rect 4181 1380 4197 1444
rect 4261 1380 4277 1444
rect 4341 1380 4357 1444
rect 4421 1380 4437 1444
rect 4501 1380 4517 1444
rect 4581 1380 4723 1444
rect 4787 1380 4803 1444
rect 4867 1380 4883 1444
rect 4947 1380 4963 1444
rect 5027 1380 5043 1444
rect 5107 1380 5123 1444
rect 5187 1380 5291 1444
rect 2801 1378 5291 1380
rect 2801 1224 2867 1378
rect 2801 1160 2802 1224
rect 2866 1160 2867 1224
rect 2801 1144 2867 1160
rect 2801 1080 2802 1144
rect 2866 1080 2867 1144
rect 2801 1064 2867 1080
rect 2801 1000 2802 1064
rect 2866 1000 2867 1064
rect 2801 984 2867 1000
rect 2801 920 2802 984
rect 2866 920 2867 984
rect 2801 904 2867 920
rect 2801 840 2802 904
rect 2866 840 2867 904
rect 2801 824 2867 840
rect 2801 760 2802 824
rect 2866 760 2867 824
rect 2801 744 2867 760
rect 2801 680 2802 744
rect 2866 680 2867 744
rect 2801 664 2867 680
rect 2801 600 2802 664
rect 2866 600 2867 664
rect 2801 584 2867 600
rect 2801 520 2802 584
rect 2866 520 2867 584
rect 2801 504 2867 520
rect 2801 440 2802 504
rect 2866 440 2867 504
rect 2801 350 2867 440
rect 2927 346 2987 1378
rect 3047 286 3107 1316
rect 3167 346 3227 1378
rect 3287 286 3347 1316
rect 3407 1224 3473 1378
rect 3407 1160 3408 1224
rect 3472 1160 3473 1224
rect 3407 1144 3473 1160
rect 3407 1080 3408 1144
rect 3472 1080 3473 1144
rect 3407 1064 3473 1080
rect 3407 1000 3408 1064
rect 3472 1000 3473 1064
rect 3407 984 3473 1000
rect 3407 920 3408 984
rect 3472 920 3473 984
rect 3407 904 3473 920
rect 3407 840 3408 904
rect 3472 840 3473 904
rect 3407 824 3473 840
rect 3407 760 3408 824
rect 3472 760 3473 824
rect 3407 744 3473 760
rect 3407 680 3408 744
rect 3472 680 3473 744
rect 3407 664 3473 680
rect 3407 600 3408 664
rect 3472 600 3473 664
rect 3407 584 3473 600
rect 3407 520 3408 584
rect 3472 520 3473 584
rect 3407 504 3473 520
rect 3407 440 3408 504
rect 3472 440 3473 504
rect 3407 350 3473 440
rect 3533 346 3593 1378
rect 3653 286 3713 1316
rect 3773 346 3833 1378
rect 3893 286 3953 1316
rect 4013 1224 4079 1378
rect 4013 1160 4014 1224
rect 4078 1160 4079 1224
rect 4013 1144 4079 1160
rect 4013 1080 4014 1144
rect 4078 1080 4079 1144
rect 4013 1064 4079 1080
rect 4013 1000 4014 1064
rect 4078 1000 4079 1064
rect 4013 984 4079 1000
rect 4013 920 4014 984
rect 4078 920 4079 984
rect 4013 904 4079 920
rect 4013 840 4014 904
rect 4078 840 4079 904
rect 4013 824 4079 840
rect 4013 760 4014 824
rect 4078 760 4079 824
rect 4013 744 4079 760
rect 4013 680 4014 744
rect 4078 680 4079 744
rect 4013 664 4079 680
rect 4013 600 4014 664
rect 4078 600 4079 664
rect 4013 584 4079 600
rect 4013 520 4014 584
rect 4078 520 4079 584
rect 4013 504 4079 520
rect 4013 440 4014 504
rect 4078 440 4079 504
rect 4013 350 4079 440
rect 4139 346 4199 1378
rect 4259 286 4319 1316
rect 4379 346 4439 1378
rect 4499 286 4559 1316
rect 4619 1224 4685 1378
rect 4619 1160 4620 1224
rect 4684 1160 4685 1224
rect 4619 1144 4685 1160
rect 4619 1080 4620 1144
rect 4684 1080 4685 1144
rect 4619 1064 4685 1080
rect 4619 1000 4620 1064
rect 4684 1000 4685 1064
rect 4619 984 4685 1000
rect 4619 920 4620 984
rect 4684 920 4685 984
rect 4619 904 4685 920
rect 4619 840 4620 904
rect 4684 840 4685 904
rect 4619 824 4685 840
rect 4619 760 4620 824
rect 4684 760 4685 824
rect 4619 744 4685 760
rect 4619 680 4620 744
rect 4684 680 4685 744
rect 4619 664 4685 680
rect 4619 600 4620 664
rect 4684 600 4685 664
rect 4619 584 4685 600
rect 4619 520 4620 584
rect 4684 520 4685 584
rect 4619 504 4685 520
rect 4619 440 4620 504
rect 4684 440 4685 504
rect 4619 350 4685 440
rect 4745 346 4805 1378
rect 4865 286 4925 1316
rect 4985 346 5045 1378
rect 5105 286 5165 1316
rect 5225 1224 5291 1378
rect 5225 1160 5226 1224
rect 5290 1160 5291 1224
rect 5225 1144 5291 1160
rect 5225 1080 5226 1144
rect 5290 1080 5291 1144
rect 5225 1064 5291 1080
rect 5225 1000 5226 1064
rect 5290 1000 5291 1064
rect 5225 984 5291 1000
rect 5225 920 5226 984
rect 5290 920 5291 984
rect 5225 904 5291 920
rect 5225 840 5226 904
rect 5290 840 5291 904
rect 5225 824 5291 840
rect 5225 760 5226 824
rect 5290 760 5291 824
rect 5225 744 5291 760
rect 5225 680 5226 744
rect 5290 680 5291 744
rect 5225 664 5291 680
rect 5225 600 5226 664
rect 5290 600 5291 664
rect 5225 584 5291 600
rect 5225 520 5226 584
rect 5290 520 5291 584
rect 5225 504 5291 520
rect 5225 440 5226 504
rect 5290 440 5291 504
rect 5225 350 5291 440
rect 5352 2384 5418 2474
rect 5352 2320 5353 2384
rect 5417 2320 5418 2384
rect 5352 2304 5418 2320
rect 5352 2240 5353 2304
rect 5417 2240 5418 2304
rect 5352 2224 5418 2240
rect 5352 2160 5353 2224
rect 5417 2160 5418 2224
rect 5352 2144 5418 2160
rect 5352 2080 5353 2144
rect 5417 2080 5418 2144
rect 5352 2064 5418 2080
rect 5352 2000 5353 2064
rect 5417 2000 5418 2064
rect 5352 1984 5418 2000
rect 5352 1920 5353 1984
rect 5417 1920 5418 1984
rect 5352 1904 5418 1920
rect 5352 1840 5353 1904
rect 5417 1840 5418 1904
rect 5352 1824 5418 1840
rect 5352 1760 5353 1824
rect 5417 1760 5418 1824
rect 5352 1744 5418 1760
rect 5352 1680 5353 1744
rect 5417 1680 5418 1744
rect 5352 1664 5418 1680
rect 5352 1600 5353 1664
rect 5417 1600 5418 1664
rect 5352 1446 5418 1600
rect 5478 1508 5538 2538
rect 5598 1446 5658 2478
rect 5718 1508 5778 2538
rect 5838 1446 5898 2478
rect 5958 2384 6024 2474
rect 5958 2320 5959 2384
rect 6023 2320 6024 2384
rect 5958 2304 6024 2320
rect 5958 2240 5959 2304
rect 6023 2240 6024 2304
rect 5958 2224 6024 2240
rect 5958 2160 5959 2224
rect 6023 2160 6024 2224
rect 5958 2144 6024 2160
rect 5958 2080 5959 2144
rect 6023 2080 6024 2144
rect 5958 2064 6024 2080
rect 5958 2000 5959 2064
rect 6023 2000 6024 2064
rect 5958 1984 6024 2000
rect 5958 1920 5959 1984
rect 6023 1920 6024 1984
rect 5958 1904 6024 1920
rect 5958 1840 5959 1904
rect 6023 1840 6024 1904
rect 5958 1824 6024 1840
rect 5958 1760 5959 1824
rect 6023 1760 6024 1824
rect 5958 1744 6024 1760
rect 5958 1680 5959 1744
rect 6023 1680 6024 1744
rect 5958 1664 6024 1680
rect 5958 1600 5959 1664
rect 6023 1600 6024 1664
rect 5958 1446 6024 1600
rect 6084 1508 6144 2538
rect 6204 1446 6264 2478
rect 6324 1508 6384 2538
rect 6444 1446 6504 2478
rect 6564 2384 6630 2474
rect 6564 2320 6565 2384
rect 6629 2320 6630 2384
rect 6564 2304 6630 2320
rect 6564 2240 6565 2304
rect 6629 2240 6630 2304
rect 6564 2224 6630 2240
rect 6564 2160 6565 2224
rect 6629 2160 6630 2224
rect 6564 2144 6630 2160
rect 6564 2080 6565 2144
rect 6629 2080 6630 2144
rect 6564 2064 6630 2080
rect 6564 2000 6565 2064
rect 6629 2000 6630 2064
rect 6564 1984 6630 2000
rect 6564 1920 6565 1984
rect 6629 1920 6630 1984
rect 6564 1904 6630 1920
rect 6564 1840 6565 1904
rect 6629 1840 6630 1904
rect 6564 1824 6630 1840
rect 6564 1760 6565 1824
rect 6629 1760 6630 1824
rect 6564 1744 6630 1760
rect 6564 1680 6565 1744
rect 6629 1680 6630 1744
rect 6564 1664 6630 1680
rect 6564 1600 6565 1664
rect 6629 1600 6630 1664
rect 6564 1446 6630 1600
rect 6690 1508 6750 2538
rect 6810 1446 6870 2478
rect 6930 1508 6990 2538
rect 7050 1446 7110 2478
rect 7170 2384 7236 2474
rect 7170 2320 7171 2384
rect 7235 2320 7236 2384
rect 7170 2304 7236 2320
rect 7170 2240 7171 2304
rect 7235 2240 7236 2304
rect 7170 2224 7236 2240
rect 7170 2160 7171 2224
rect 7235 2160 7236 2224
rect 7170 2144 7236 2160
rect 7170 2080 7171 2144
rect 7235 2080 7236 2144
rect 7170 2064 7236 2080
rect 7170 2000 7171 2064
rect 7235 2000 7236 2064
rect 7170 1984 7236 2000
rect 7170 1920 7171 1984
rect 7235 1920 7236 1984
rect 7170 1904 7236 1920
rect 7170 1840 7171 1904
rect 7235 1840 7236 1904
rect 7170 1824 7236 1840
rect 7170 1760 7171 1824
rect 7235 1760 7236 1824
rect 7170 1744 7236 1760
rect 7170 1680 7171 1744
rect 7235 1680 7236 1744
rect 7170 1664 7236 1680
rect 7170 1600 7171 1664
rect 7235 1600 7236 1664
rect 7170 1446 7236 1600
rect 7296 1508 7356 2538
rect 7416 1446 7476 2478
rect 7536 1508 7596 2538
rect 7656 1446 7716 2478
rect 7776 2384 7842 2474
rect 7776 2320 7777 2384
rect 7841 2320 7842 2384
rect 7776 2304 7842 2320
rect 7776 2240 7777 2304
rect 7841 2240 7842 2304
rect 7776 2224 7842 2240
rect 7776 2160 7777 2224
rect 7841 2160 7842 2224
rect 7776 2144 7842 2160
rect 7776 2080 7777 2144
rect 7841 2080 7842 2144
rect 7776 2064 7842 2080
rect 7776 2000 7777 2064
rect 7841 2000 7842 2064
rect 7776 1984 7842 2000
rect 7776 1920 7777 1984
rect 7841 1920 7842 1984
rect 7776 1904 7842 1920
rect 7776 1840 7777 1904
rect 7841 1840 7842 1904
rect 7776 1824 7842 1840
rect 7776 1760 7777 1824
rect 7841 1760 7842 1824
rect 7776 1744 7842 1760
rect 7776 1680 7777 1744
rect 7841 1680 7842 1744
rect 7776 1664 7842 1680
rect 7776 1600 7777 1664
rect 7841 1600 7842 1664
rect 7776 1446 7842 1600
rect 7902 1508 7962 2538
rect 8022 1446 8082 2478
rect 8142 1508 8202 2538
rect 8262 1446 8322 2478
rect 8382 2384 8448 2474
rect 8382 2320 8383 2384
rect 8447 2320 8448 2384
rect 8382 2304 8448 2320
rect 8382 2240 8383 2304
rect 8447 2240 8448 2304
rect 8382 2224 8448 2240
rect 8382 2160 8383 2224
rect 8447 2160 8448 2224
rect 8382 2144 8448 2160
rect 8382 2080 8383 2144
rect 8447 2080 8448 2144
rect 8382 2064 8448 2080
rect 8382 2000 8383 2064
rect 8447 2000 8448 2064
rect 8382 1984 8448 2000
rect 8382 1920 8383 1984
rect 8447 1920 8448 1984
rect 8382 1904 8448 1920
rect 8382 1840 8383 1904
rect 8447 1840 8448 1904
rect 8382 1824 8448 1840
rect 8382 1760 8383 1824
rect 8447 1760 8448 1824
rect 8382 1744 8448 1760
rect 8382 1680 8383 1744
rect 8447 1680 8448 1744
rect 8382 1664 8448 1680
rect 8382 1600 8383 1664
rect 8447 1600 8448 1664
rect 8382 1446 8448 1600
rect 8508 1508 8568 2538
rect 8628 1446 8688 2478
rect 8748 1508 8808 2538
rect 8868 1446 8928 2478
rect 8988 2384 9054 2474
rect 8988 2320 8989 2384
rect 9053 2320 9054 2384
rect 8988 2304 9054 2320
rect 8988 2240 8989 2304
rect 9053 2240 9054 2304
rect 8988 2224 9054 2240
rect 8988 2160 8989 2224
rect 9053 2160 9054 2224
rect 8988 2144 9054 2160
rect 8988 2080 8989 2144
rect 9053 2080 9054 2144
rect 8988 2064 9054 2080
rect 8988 2000 8989 2064
rect 9053 2000 9054 2064
rect 8988 1984 9054 2000
rect 8988 1920 8989 1984
rect 9053 1920 9054 1984
rect 8988 1904 9054 1920
rect 8988 1840 8989 1904
rect 9053 1840 9054 1904
rect 8988 1824 9054 1840
rect 8988 1760 8989 1824
rect 9053 1760 9054 1824
rect 8988 1744 9054 1760
rect 8988 1680 8989 1744
rect 9053 1680 9054 1744
rect 8988 1664 9054 1680
rect 8988 1600 8989 1664
rect 9053 1600 9054 1664
rect 8988 1446 9054 1600
rect 9114 1508 9174 2538
rect 9234 1446 9294 2478
rect 9354 1508 9414 2538
rect 9474 1446 9534 2478
rect 9594 2384 9660 2474
rect 9594 2320 9595 2384
rect 9659 2320 9660 2384
rect 9594 2304 9660 2320
rect 9594 2240 9595 2304
rect 9659 2240 9660 2304
rect 9594 2224 9660 2240
rect 9594 2160 9595 2224
rect 9659 2160 9660 2224
rect 9594 2144 9660 2160
rect 9594 2080 9595 2144
rect 9659 2080 9660 2144
rect 9594 2064 9660 2080
rect 9594 2000 9595 2064
rect 9659 2000 9660 2064
rect 9594 1984 9660 2000
rect 9594 1920 9595 1984
rect 9659 1920 9660 1984
rect 9594 1904 9660 1920
rect 9594 1840 9595 1904
rect 9659 1840 9660 1904
rect 9594 1824 9660 1840
rect 9594 1760 9595 1824
rect 9659 1760 9660 1824
rect 9594 1744 9660 1760
rect 9594 1680 9595 1744
rect 9659 1680 9660 1744
rect 9594 1664 9660 1680
rect 9594 1600 9595 1664
rect 9659 1600 9660 1664
rect 9594 1446 9660 1600
rect 9720 1508 9780 2538
rect 9840 1446 9900 2478
rect 9960 1508 10020 2538
rect 10080 1446 10140 2478
rect 10200 2384 10266 2474
rect 10200 2320 10201 2384
rect 10265 2320 10266 2384
rect 10200 2304 10266 2320
rect 10200 2240 10201 2304
rect 10265 2240 10266 2304
rect 10200 2224 10266 2240
rect 10200 2160 10201 2224
rect 10265 2160 10266 2224
rect 10200 2144 10266 2160
rect 10200 2080 10201 2144
rect 10265 2080 10266 2144
rect 10200 2064 10266 2080
rect 10200 2000 10201 2064
rect 10265 2000 10266 2064
rect 10200 1984 10266 2000
rect 10200 1920 10201 1984
rect 10265 1920 10266 1984
rect 10200 1904 10266 1920
rect 10200 1840 10201 1904
rect 10265 1840 10266 1904
rect 10200 1824 10266 1840
rect 10200 1760 10201 1824
rect 10265 1760 10266 1824
rect 10200 1744 10266 1760
rect 10200 1680 10201 1744
rect 10265 1680 10266 1744
rect 10200 1664 10266 1680
rect 10200 1600 10201 1664
rect 10265 1600 10266 1664
rect 10200 1446 10266 1600
rect 5352 1444 10266 1446
rect 5352 1380 5456 1444
rect 5520 1380 5536 1444
rect 5600 1380 5616 1444
rect 5680 1380 5696 1444
rect 5760 1380 5776 1444
rect 5840 1380 5856 1444
rect 5920 1380 6062 1444
rect 6126 1380 6142 1444
rect 6206 1380 6222 1444
rect 6286 1380 6302 1444
rect 6366 1380 6382 1444
rect 6446 1380 6462 1444
rect 6526 1380 6668 1444
rect 6732 1380 6748 1444
rect 6812 1380 6828 1444
rect 6892 1380 6908 1444
rect 6972 1380 6988 1444
rect 7052 1380 7068 1444
rect 7132 1380 7274 1444
rect 7338 1380 7354 1444
rect 7418 1380 7434 1444
rect 7498 1380 7514 1444
rect 7578 1380 7594 1444
rect 7658 1380 7674 1444
rect 7738 1380 7880 1444
rect 7944 1380 7960 1444
rect 8024 1380 8040 1444
rect 8104 1380 8120 1444
rect 8184 1380 8200 1444
rect 8264 1380 8280 1444
rect 8344 1380 8486 1444
rect 8550 1380 8566 1444
rect 8630 1380 8646 1444
rect 8710 1380 8726 1444
rect 8790 1380 8806 1444
rect 8870 1380 8886 1444
rect 8950 1380 9092 1444
rect 9156 1380 9172 1444
rect 9236 1380 9252 1444
rect 9316 1380 9332 1444
rect 9396 1380 9412 1444
rect 9476 1380 9492 1444
rect 9556 1380 9698 1444
rect 9762 1380 9778 1444
rect 9842 1380 9858 1444
rect 9922 1380 9938 1444
rect 10002 1380 10018 1444
rect 10082 1380 10098 1444
rect 10162 1380 10266 1444
rect 5352 1378 10266 1380
rect 5352 1224 5418 1378
rect 5352 1160 5353 1224
rect 5417 1160 5418 1224
rect 5352 1144 5418 1160
rect 5352 1080 5353 1144
rect 5417 1080 5418 1144
rect 5352 1064 5418 1080
rect 5352 1000 5353 1064
rect 5417 1000 5418 1064
rect 5352 984 5418 1000
rect 5352 920 5353 984
rect 5417 920 5418 984
rect 5352 904 5418 920
rect 5352 840 5353 904
rect 5417 840 5418 904
rect 5352 824 5418 840
rect 5352 760 5353 824
rect 5417 760 5418 824
rect 5352 744 5418 760
rect 5352 680 5353 744
rect 5417 680 5418 744
rect 5352 664 5418 680
rect 5352 600 5353 664
rect 5417 600 5418 664
rect 5352 584 5418 600
rect 5352 520 5353 584
rect 5417 520 5418 584
rect 5352 504 5418 520
rect 5352 440 5353 504
rect 5417 440 5418 504
rect 5352 350 5418 440
rect 5478 346 5538 1378
rect 5598 286 5658 1316
rect 5718 346 5778 1378
rect 5838 286 5898 1316
rect 5958 1224 6024 1378
rect 5958 1160 5959 1224
rect 6023 1160 6024 1224
rect 5958 1144 6024 1160
rect 5958 1080 5959 1144
rect 6023 1080 6024 1144
rect 5958 1064 6024 1080
rect 5958 1000 5959 1064
rect 6023 1000 6024 1064
rect 5958 984 6024 1000
rect 5958 920 5959 984
rect 6023 920 6024 984
rect 5958 904 6024 920
rect 5958 840 5959 904
rect 6023 840 6024 904
rect 5958 824 6024 840
rect 5958 760 5959 824
rect 6023 760 6024 824
rect 5958 744 6024 760
rect 5958 680 5959 744
rect 6023 680 6024 744
rect 5958 664 6024 680
rect 5958 600 5959 664
rect 6023 600 6024 664
rect 5958 584 6024 600
rect 5958 520 5959 584
rect 6023 520 6024 584
rect 5958 504 6024 520
rect 5958 440 5959 504
rect 6023 440 6024 504
rect 5958 350 6024 440
rect 6084 346 6144 1378
rect 6204 286 6264 1316
rect 6324 346 6384 1378
rect 6444 286 6504 1316
rect 6564 1224 6630 1378
rect 6564 1160 6565 1224
rect 6629 1160 6630 1224
rect 6564 1144 6630 1160
rect 6564 1080 6565 1144
rect 6629 1080 6630 1144
rect 6564 1064 6630 1080
rect 6564 1000 6565 1064
rect 6629 1000 6630 1064
rect 6564 984 6630 1000
rect 6564 920 6565 984
rect 6629 920 6630 984
rect 6564 904 6630 920
rect 6564 840 6565 904
rect 6629 840 6630 904
rect 6564 824 6630 840
rect 6564 760 6565 824
rect 6629 760 6630 824
rect 6564 744 6630 760
rect 6564 680 6565 744
rect 6629 680 6630 744
rect 6564 664 6630 680
rect 6564 600 6565 664
rect 6629 600 6630 664
rect 6564 584 6630 600
rect 6564 520 6565 584
rect 6629 520 6630 584
rect 6564 504 6630 520
rect 6564 440 6565 504
rect 6629 440 6630 504
rect 6564 350 6630 440
rect 6690 346 6750 1378
rect 6810 286 6870 1316
rect 6930 346 6990 1378
rect 7050 286 7110 1316
rect 7170 1224 7236 1378
rect 7170 1160 7171 1224
rect 7235 1160 7236 1224
rect 7170 1144 7236 1160
rect 7170 1080 7171 1144
rect 7235 1080 7236 1144
rect 7170 1064 7236 1080
rect 7170 1000 7171 1064
rect 7235 1000 7236 1064
rect 7170 984 7236 1000
rect 7170 920 7171 984
rect 7235 920 7236 984
rect 7170 904 7236 920
rect 7170 840 7171 904
rect 7235 840 7236 904
rect 7170 824 7236 840
rect 7170 760 7171 824
rect 7235 760 7236 824
rect 7170 744 7236 760
rect 7170 680 7171 744
rect 7235 680 7236 744
rect 7170 664 7236 680
rect 7170 600 7171 664
rect 7235 600 7236 664
rect 7170 584 7236 600
rect 7170 520 7171 584
rect 7235 520 7236 584
rect 7170 504 7236 520
rect 7170 440 7171 504
rect 7235 440 7236 504
rect 7170 350 7236 440
rect 7296 346 7356 1378
rect 7416 286 7476 1316
rect 7536 346 7596 1378
rect 7656 286 7716 1316
rect 7776 1224 7842 1378
rect 7776 1160 7777 1224
rect 7841 1160 7842 1224
rect 7776 1144 7842 1160
rect 7776 1080 7777 1144
rect 7841 1080 7842 1144
rect 7776 1064 7842 1080
rect 7776 1000 7777 1064
rect 7841 1000 7842 1064
rect 7776 984 7842 1000
rect 7776 920 7777 984
rect 7841 920 7842 984
rect 7776 904 7842 920
rect 7776 840 7777 904
rect 7841 840 7842 904
rect 7776 824 7842 840
rect 7776 760 7777 824
rect 7841 760 7842 824
rect 7776 744 7842 760
rect 7776 680 7777 744
rect 7841 680 7842 744
rect 7776 664 7842 680
rect 7776 600 7777 664
rect 7841 600 7842 664
rect 7776 584 7842 600
rect 7776 520 7777 584
rect 7841 520 7842 584
rect 7776 504 7842 520
rect 7776 440 7777 504
rect 7841 440 7842 504
rect 7776 350 7842 440
rect 7902 346 7962 1378
rect 8022 286 8082 1316
rect 8142 346 8202 1378
rect 8262 286 8322 1316
rect 8382 1224 8448 1378
rect 8382 1160 8383 1224
rect 8447 1160 8448 1224
rect 8382 1144 8448 1160
rect 8382 1080 8383 1144
rect 8447 1080 8448 1144
rect 8382 1064 8448 1080
rect 8382 1000 8383 1064
rect 8447 1000 8448 1064
rect 8382 984 8448 1000
rect 8382 920 8383 984
rect 8447 920 8448 984
rect 8382 904 8448 920
rect 8382 840 8383 904
rect 8447 840 8448 904
rect 8382 824 8448 840
rect 8382 760 8383 824
rect 8447 760 8448 824
rect 8382 744 8448 760
rect 8382 680 8383 744
rect 8447 680 8448 744
rect 8382 664 8448 680
rect 8382 600 8383 664
rect 8447 600 8448 664
rect 8382 584 8448 600
rect 8382 520 8383 584
rect 8447 520 8448 584
rect 8382 504 8448 520
rect 8382 440 8383 504
rect 8447 440 8448 504
rect 8382 350 8448 440
rect 8508 346 8568 1378
rect 8628 286 8688 1316
rect 8748 346 8808 1378
rect 8868 286 8928 1316
rect 8988 1224 9054 1378
rect 8988 1160 8989 1224
rect 9053 1160 9054 1224
rect 8988 1144 9054 1160
rect 8988 1080 8989 1144
rect 9053 1080 9054 1144
rect 8988 1064 9054 1080
rect 8988 1000 8989 1064
rect 9053 1000 9054 1064
rect 8988 984 9054 1000
rect 8988 920 8989 984
rect 9053 920 9054 984
rect 8988 904 9054 920
rect 8988 840 8989 904
rect 9053 840 9054 904
rect 8988 824 9054 840
rect 8988 760 8989 824
rect 9053 760 9054 824
rect 8988 744 9054 760
rect 8988 680 8989 744
rect 9053 680 9054 744
rect 8988 664 9054 680
rect 8988 600 8989 664
rect 9053 600 9054 664
rect 8988 584 9054 600
rect 8988 520 8989 584
rect 9053 520 9054 584
rect 8988 504 9054 520
rect 8988 440 8989 504
rect 9053 440 9054 504
rect 8988 350 9054 440
rect 9114 346 9174 1378
rect 9234 286 9294 1316
rect 9354 346 9414 1378
rect 9474 286 9534 1316
rect 9594 1224 9660 1378
rect 9594 1160 9595 1224
rect 9659 1160 9660 1224
rect 9594 1144 9660 1160
rect 9594 1080 9595 1144
rect 9659 1080 9660 1144
rect 9594 1064 9660 1080
rect 9594 1000 9595 1064
rect 9659 1000 9660 1064
rect 9594 984 9660 1000
rect 9594 920 9595 984
rect 9659 920 9660 984
rect 9594 904 9660 920
rect 9594 840 9595 904
rect 9659 840 9660 904
rect 9594 824 9660 840
rect 9594 760 9595 824
rect 9659 760 9660 824
rect 9594 744 9660 760
rect 9594 680 9595 744
rect 9659 680 9660 744
rect 9594 664 9660 680
rect 9594 600 9595 664
rect 9659 600 9660 664
rect 9594 584 9660 600
rect 9594 520 9595 584
rect 9659 520 9660 584
rect 9594 504 9660 520
rect 9594 440 9595 504
rect 9659 440 9660 504
rect 9594 350 9660 440
rect 9720 346 9780 1378
rect 9840 286 9900 1316
rect 9960 346 10020 1378
rect 10080 286 10140 1316
rect 10200 1224 10266 1378
rect 10200 1160 10201 1224
rect 10265 1160 10266 1224
rect 10200 1144 10266 1160
rect 10200 1080 10201 1144
rect 10265 1080 10266 1144
rect 10200 1064 10266 1080
rect 10200 1000 10201 1064
rect 10265 1000 10266 1064
rect 10200 984 10266 1000
rect 10200 920 10201 984
rect 10265 920 10266 984
rect 10200 904 10266 920
rect 10200 840 10201 904
rect 10265 840 10266 904
rect 10200 824 10266 840
rect 10200 760 10201 824
rect 10265 760 10266 824
rect 10200 744 10266 760
rect 10200 680 10201 744
rect 10265 680 10266 744
rect 10200 664 10266 680
rect 10200 600 10201 664
rect 10265 600 10266 664
rect 10200 584 10266 600
rect 10200 520 10201 584
rect 10265 520 10266 584
rect 10200 504 10266 520
rect 10200 440 10201 504
rect 10265 440 10266 504
rect 10200 350 10266 440
rect 10326 2384 10392 2474
rect 10326 2320 10327 2384
rect 10391 2320 10392 2384
rect 10326 2304 10392 2320
rect 10326 2240 10327 2304
rect 10391 2240 10392 2304
rect 10326 2224 10392 2240
rect 10326 2160 10327 2224
rect 10391 2160 10392 2224
rect 10326 2144 10392 2160
rect 10326 2080 10327 2144
rect 10391 2080 10392 2144
rect 10326 2064 10392 2080
rect 10326 2000 10327 2064
rect 10391 2000 10392 2064
rect 10326 1984 10392 2000
rect 10326 1920 10327 1984
rect 10391 1920 10392 1984
rect 10326 1904 10392 1920
rect 10326 1840 10327 1904
rect 10391 1840 10392 1904
rect 10326 1824 10392 1840
rect 10326 1760 10327 1824
rect 10391 1760 10392 1824
rect 10326 1744 10392 1760
rect 10326 1680 10327 1744
rect 10391 1680 10392 1744
rect 10326 1664 10392 1680
rect 10326 1600 10327 1664
rect 10391 1600 10392 1664
rect 10326 1446 10392 1600
rect 10452 1508 10512 2538
rect 10572 1446 10632 2478
rect 10692 1508 10752 2538
rect 10812 1446 10872 2478
rect 10932 2384 10998 2474
rect 10932 2320 10933 2384
rect 10997 2320 10998 2384
rect 10932 2304 10998 2320
rect 10932 2240 10933 2304
rect 10997 2240 10998 2304
rect 10932 2224 10998 2240
rect 10932 2160 10933 2224
rect 10997 2160 10998 2224
rect 10932 2144 10998 2160
rect 10932 2080 10933 2144
rect 10997 2080 10998 2144
rect 10932 2064 10998 2080
rect 10932 2000 10933 2064
rect 10997 2000 10998 2064
rect 10932 1984 10998 2000
rect 10932 1920 10933 1984
rect 10997 1920 10998 1984
rect 10932 1904 10998 1920
rect 10932 1840 10933 1904
rect 10997 1840 10998 1904
rect 10932 1824 10998 1840
rect 10932 1760 10933 1824
rect 10997 1760 10998 1824
rect 10932 1744 10998 1760
rect 10932 1680 10933 1744
rect 10997 1680 10998 1744
rect 10932 1664 10998 1680
rect 10932 1600 10933 1664
rect 10997 1600 10998 1664
rect 10932 1446 10998 1600
rect 11058 1508 11118 2538
rect 11178 1446 11238 2478
rect 11298 1508 11358 2538
rect 11418 1446 11478 2478
rect 11538 2384 11604 2474
rect 11538 2320 11539 2384
rect 11603 2320 11604 2384
rect 11538 2304 11604 2320
rect 11538 2240 11539 2304
rect 11603 2240 11604 2304
rect 11538 2224 11604 2240
rect 11538 2160 11539 2224
rect 11603 2160 11604 2224
rect 11538 2144 11604 2160
rect 11538 2080 11539 2144
rect 11603 2080 11604 2144
rect 11538 2064 11604 2080
rect 11538 2000 11539 2064
rect 11603 2000 11604 2064
rect 11538 1984 11604 2000
rect 11538 1920 11539 1984
rect 11603 1920 11604 1984
rect 11538 1904 11604 1920
rect 11538 1840 11539 1904
rect 11603 1840 11604 1904
rect 11538 1824 11604 1840
rect 11538 1760 11539 1824
rect 11603 1760 11604 1824
rect 11538 1744 11604 1760
rect 11538 1680 11539 1744
rect 11603 1680 11604 1744
rect 11538 1664 11604 1680
rect 11538 1600 11539 1664
rect 11603 1600 11604 1664
rect 11538 1446 11604 1600
rect 11664 1508 11724 2538
rect 11784 1446 11844 2478
rect 11904 1508 11964 2538
rect 12024 1446 12084 2478
rect 12144 2384 12210 2474
rect 12144 2320 12145 2384
rect 12209 2320 12210 2384
rect 12144 2304 12210 2320
rect 12144 2240 12145 2304
rect 12209 2240 12210 2304
rect 12144 2224 12210 2240
rect 12144 2160 12145 2224
rect 12209 2160 12210 2224
rect 12144 2144 12210 2160
rect 12144 2080 12145 2144
rect 12209 2080 12210 2144
rect 12144 2064 12210 2080
rect 12144 2000 12145 2064
rect 12209 2000 12210 2064
rect 12144 1984 12210 2000
rect 12144 1920 12145 1984
rect 12209 1920 12210 1984
rect 12144 1904 12210 1920
rect 12144 1840 12145 1904
rect 12209 1840 12210 1904
rect 12144 1824 12210 1840
rect 12144 1760 12145 1824
rect 12209 1760 12210 1824
rect 12144 1744 12210 1760
rect 12144 1680 12145 1744
rect 12209 1680 12210 1744
rect 12144 1664 12210 1680
rect 12144 1600 12145 1664
rect 12209 1600 12210 1664
rect 12144 1446 12210 1600
rect 12270 1508 12330 2538
rect 12390 1446 12450 2478
rect 12510 1508 12570 2538
rect 12630 1446 12690 2478
rect 12750 2384 12816 2474
rect 12750 2320 12751 2384
rect 12815 2320 12816 2384
rect 12750 2304 12816 2320
rect 12750 2240 12751 2304
rect 12815 2240 12816 2304
rect 12750 2224 12816 2240
rect 12750 2160 12751 2224
rect 12815 2160 12816 2224
rect 12750 2144 12816 2160
rect 12750 2080 12751 2144
rect 12815 2080 12816 2144
rect 12750 2064 12816 2080
rect 12750 2000 12751 2064
rect 12815 2000 12816 2064
rect 12750 1984 12816 2000
rect 12750 1920 12751 1984
rect 12815 1920 12816 1984
rect 12750 1904 12816 1920
rect 12750 1840 12751 1904
rect 12815 1840 12816 1904
rect 12750 1824 12816 1840
rect 12750 1760 12751 1824
rect 12815 1760 12816 1824
rect 12750 1744 12816 1760
rect 12750 1680 12751 1744
rect 12815 1680 12816 1744
rect 12750 1664 12816 1680
rect 12750 1600 12751 1664
rect 12815 1600 12816 1664
rect 12750 1446 12816 1600
rect 12876 1508 12936 2538
rect 12996 1446 13056 2478
rect 13116 1508 13176 2538
rect 13236 1446 13296 2478
rect 13356 2384 13422 2474
rect 13356 2320 13357 2384
rect 13421 2320 13422 2384
rect 13356 2304 13422 2320
rect 13356 2240 13357 2304
rect 13421 2240 13422 2304
rect 13356 2224 13422 2240
rect 13356 2160 13357 2224
rect 13421 2160 13422 2224
rect 13356 2144 13422 2160
rect 13356 2080 13357 2144
rect 13421 2080 13422 2144
rect 13356 2064 13422 2080
rect 13356 2000 13357 2064
rect 13421 2000 13422 2064
rect 13356 1984 13422 2000
rect 13356 1920 13357 1984
rect 13421 1920 13422 1984
rect 13356 1904 13422 1920
rect 13356 1840 13357 1904
rect 13421 1840 13422 1904
rect 13356 1824 13422 1840
rect 13356 1760 13357 1824
rect 13421 1760 13422 1824
rect 13356 1744 13422 1760
rect 13356 1680 13357 1744
rect 13421 1680 13422 1744
rect 13356 1664 13422 1680
rect 13356 1600 13357 1664
rect 13421 1600 13422 1664
rect 13356 1446 13422 1600
rect 13482 1508 13542 2538
rect 13602 1446 13662 2478
rect 13722 1508 13782 2538
rect 13842 1446 13902 2478
rect 13962 2384 14028 2474
rect 13962 2320 13963 2384
rect 14027 2320 14028 2384
rect 13962 2304 14028 2320
rect 13962 2240 13963 2304
rect 14027 2240 14028 2304
rect 13962 2224 14028 2240
rect 13962 2160 13963 2224
rect 14027 2160 14028 2224
rect 13962 2144 14028 2160
rect 13962 2080 13963 2144
rect 14027 2080 14028 2144
rect 13962 2064 14028 2080
rect 13962 2000 13963 2064
rect 14027 2000 14028 2064
rect 13962 1984 14028 2000
rect 13962 1920 13963 1984
rect 14027 1920 14028 1984
rect 13962 1904 14028 1920
rect 13962 1840 13963 1904
rect 14027 1840 14028 1904
rect 13962 1824 14028 1840
rect 13962 1760 13963 1824
rect 14027 1760 14028 1824
rect 13962 1744 14028 1760
rect 13962 1680 13963 1744
rect 14027 1680 14028 1744
rect 13962 1664 14028 1680
rect 13962 1600 13963 1664
rect 14027 1600 14028 1664
rect 13962 1446 14028 1600
rect 14088 1508 14148 2538
rect 14208 1446 14268 2478
rect 14328 1508 14388 2538
rect 14448 1446 14508 2478
rect 14568 2384 14634 2474
rect 14568 2320 14569 2384
rect 14633 2320 14634 2384
rect 14568 2304 14634 2320
rect 14568 2240 14569 2304
rect 14633 2240 14634 2304
rect 14568 2224 14634 2240
rect 14568 2160 14569 2224
rect 14633 2160 14634 2224
rect 14568 2144 14634 2160
rect 14568 2080 14569 2144
rect 14633 2080 14634 2144
rect 14568 2064 14634 2080
rect 14568 2000 14569 2064
rect 14633 2000 14634 2064
rect 14568 1984 14634 2000
rect 14568 1920 14569 1984
rect 14633 1920 14634 1984
rect 14568 1904 14634 1920
rect 14568 1840 14569 1904
rect 14633 1840 14634 1904
rect 14568 1824 14634 1840
rect 14568 1760 14569 1824
rect 14633 1760 14634 1824
rect 14568 1744 14634 1760
rect 14568 1680 14569 1744
rect 14633 1680 14634 1744
rect 14568 1664 14634 1680
rect 14568 1600 14569 1664
rect 14633 1600 14634 1664
rect 14568 1446 14634 1600
rect 14694 1508 14754 2538
rect 14814 1446 14874 2478
rect 14934 1508 14994 2538
rect 15054 1446 15114 2478
rect 15174 2384 15240 2474
rect 15174 2320 15175 2384
rect 15239 2320 15240 2384
rect 15174 2304 15240 2320
rect 15174 2240 15175 2304
rect 15239 2240 15240 2304
rect 15174 2224 15240 2240
rect 15174 2160 15175 2224
rect 15239 2160 15240 2224
rect 15174 2144 15240 2160
rect 15174 2080 15175 2144
rect 15239 2080 15240 2144
rect 15174 2064 15240 2080
rect 15174 2000 15175 2064
rect 15239 2000 15240 2064
rect 15174 1984 15240 2000
rect 15174 1920 15175 1984
rect 15239 1920 15240 1984
rect 15174 1904 15240 1920
rect 15174 1840 15175 1904
rect 15239 1840 15240 1904
rect 15174 1824 15240 1840
rect 15174 1760 15175 1824
rect 15239 1760 15240 1824
rect 15174 1744 15240 1760
rect 15174 1680 15175 1744
rect 15239 1680 15240 1744
rect 15174 1664 15240 1680
rect 15174 1600 15175 1664
rect 15239 1600 15240 1664
rect 15174 1446 15240 1600
rect 15300 1508 15360 2538
rect 15420 1446 15480 2478
rect 15540 1508 15600 2538
rect 15660 1446 15720 2478
rect 15780 2384 15846 2474
rect 15780 2320 15781 2384
rect 15845 2320 15846 2384
rect 15780 2304 15846 2320
rect 15780 2240 15781 2304
rect 15845 2240 15846 2304
rect 15780 2224 15846 2240
rect 15780 2160 15781 2224
rect 15845 2160 15846 2224
rect 15780 2144 15846 2160
rect 15780 2080 15781 2144
rect 15845 2080 15846 2144
rect 15780 2064 15846 2080
rect 15780 2000 15781 2064
rect 15845 2000 15846 2064
rect 15780 1984 15846 2000
rect 15780 1920 15781 1984
rect 15845 1920 15846 1984
rect 15780 1904 15846 1920
rect 15780 1840 15781 1904
rect 15845 1840 15846 1904
rect 15780 1824 15846 1840
rect 15780 1760 15781 1824
rect 15845 1760 15846 1824
rect 15780 1744 15846 1760
rect 15780 1680 15781 1744
rect 15845 1680 15846 1744
rect 15780 1664 15846 1680
rect 15780 1600 15781 1664
rect 15845 1600 15846 1664
rect 15780 1446 15846 1600
rect 15906 1508 15966 2538
rect 16026 1446 16086 2478
rect 16146 1508 16206 2538
rect 16266 1446 16326 2478
rect 16386 2384 16452 2474
rect 16386 2320 16387 2384
rect 16451 2320 16452 2384
rect 16386 2304 16452 2320
rect 16386 2240 16387 2304
rect 16451 2240 16452 2304
rect 16386 2224 16452 2240
rect 16386 2160 16387 2224
rect 16451 2160 16452 2224
rect 16386 2144 16452 2160
rect 16386 2080 16387 2144
rect 16451 2080 16452 2144
rect 16386 2064 16452 2080
rect 16386 2000 16387 2064
rect 16451 2000 16452 2064
rect 16386 1984 16452 2000
rect 16386 1920 16387 1984
rect 16451 1920 16452 1984
rect 16386 1904 16452 1920
rect 16386 1840 16387 1904
rect 16451 1840 16452 1904
rect 16386 1824 16452 1840
rect 16386 1760 16387 1824
rect 16451 1760 16452 1824
rect 16386 1744 16452 1760
rect 16386 1680 16387 1744
rect 16451 1680 16452 1744
rect 16386 1664 16452 1680
rect 16386 1600 16387 1664
rect 16451 1600 16452 1664
rect 16386 1446 16452 1600
rect 16512 1508 16572 2538
rect 16632 1446 16692 2478
rect 16752 1508 16812 2538
rect 16872 1446 16932 2478
rect 16992 2384 17058 2474
rect 16992 2320 16993 2384
rect 17057 2320 17058 2384
rect 16992 2304 17058 2320
rect 16992 2240 16993 2304
rect 17057 2240 17058 2304
rect 16992 2224 17058 2240
rect 16992 2160 16993 2224
rect 17057 2160 17058 2224
rect 16992 2144 17058 2160
rect 16992 2080 16993 2144
rect 17057 2080 17058 2144
rect 16992 2064 17058 2080
rect 16992 2000 16993 2064
rect 17057 2000 17058 2064
rect 16992 1984 17058 2000
rect 16992 1920 16993 1984
rect 17057 1920 17058 1984
rect 16992 1904 17058 1920
rect 16992 1840 16993 1904
rect 17057 1840 17058 1904
rect 16992 1824 17058 1840
rect 16992 1760 16993 1824
rect 17057 1760 17058 1824
rect 16992 1744 17058 1760
rect 16992 1680 16993 1744
rect 17057 1680 17058 1744
rect 16992 1664 17058 1680
rect 16992 1600 16993 1664
rect 17057 1600 17058 1664
rect 16992 1446 17058 1600
rect 17118 1508 17178 2538
rect 17238 1446 17298 2478
rect 17358 1508 17418 2538
rect 17478 1446 17538 2478
rect 17598 2384 17664 2474
rect 17598 2320 17599 2384
rect 17663 2320 17664 2384
rect 17598 2304 17664 2320
rect 17598 2240 17599 2304
rect 17663 2240 17664 2304
rect 17598 2224 17664 2240
rect 17598 2160 17599 2224
rect 17663 2160 17664 2224
rect 17598 2144 17664 2160
rect 17598 2080 17599 2144
rect 17663 2080 17664 2144
rect 17598 2064 17664 2080
rect 17598 2000 17599 2064
rect 17663 2000 17664 2064
rect 17598 1984 17664 2000
rect 17598 1920 17599 1984
rect 17663 1920 17664 1984
rect 17598 1904 17664 1920
rect 17598 1840 17599 1904
rect 17663 1840 17664 1904
rect 17598 1824 17664 1840
rect 17598 1760 17599 1824
rect 17663 1760 17664 1824
rect 17598 1744 17664 1760
rect 17598 1680 17599 1744
rect 17663 1680 17664 1744
rect 17598 1664 17664 1680
rect 17598 1600 17599 1664
rect 17663 1600 17664 1664
rect 17598 1446 17664 1600
rect 17724 1508 17784 2538
rect 17844 1446 17904 2478
rect 17964 1508 18024 2538
rect 18084 1446 18144 2478
rect 18204 2384 18270 2474
rect 18204 2320 18205 2384
rect 18269 2320 18270 2384
rect 18204 2304 18270 2320
rect 18204 2240 18205 2304
rect 18269 2240 18270 2304
rect 18204 2224 18270 2240
rect 18204 2160 18205 2224
rect 18269 2160 18270 2224
rect 18204 2144 18270 2160
rect 18204 2080 18205 2144
rect 18269 2080 18270 2144
rect 18204 2064 18270 2080
rect 18204 2000 18205 2064
rect 18269 2000 18270 2064
rect 18204 1984 18270 2000
rect 18204 1920 18205 1984
rect 18269 1920 18270 1984
rect 18204 1904 18270 1920
rect 18204 1840 18205 1904
rect 18269 1840 18270 1904
rect 18204 1824 18270 1840
rect 18204 1760 18205 1824
rect 18269 1760 18270 1824
rect 18204 1744 18270 1760
rect 18204 1680 18205 1744
rect 18269 1680 18270 1744
rect 18204 1664 18270 1680
rect 18204 1600 18205 1664
rect 18269 1600 18270 1664
rect 18204 1446 18270 1600
rect 18330 1508 18390 2538
rect 18450 1446 18510 2478
rect 18570 1508 18630 2538
rect 18690 1446 18750 2478
rect 18810 2384 18876 2474
rect 18810 2320 18811 2384
rect 18875 2320 18876 2384
rect 18810 2304 18876 2320
rect 18810 2240 18811 2304
rect 18875 2240 18876 2304
rect 18810 2224 18876 2240
rect 18810 2160 18811 2224
rect 18875 2160 18876 2224
rect 18810 2144 18876 2160
rect 18810 2080 18811 2144
rect 18875 2080 18876 2144
rect 18810 2064 18876 2080
rect 18810 2000 18811 2064
rect 18875 2000 18876 2064
rect 18810 1984 18876 2000
rect 18810 1920 18811 1984
rect 18875 1920 18876 1984
rect 18810 1904 18876 1920
rect 18810 1840 18811 1904
rect 18875 1840 18876 1904
rect 18810 1824 18876 1840
rect 18810 1760 18811 1824
rect 18875 1760 18876 1824
rect 18810 1744 18876 1760
rect 18810 1680 18811 1744
rect 18875 1680 18876 1744
rect 18810 1664 18876 1680
rect 18810 1600 18811 1664
rect 18875 1600 18876 1664
rect 18810 1446 18876 1600
rect 18936 1508 18996 2538
rect 19056 1446 19116 2478
rect 19176 1508 19236 2538
rect 19296 1446 19356 2478
rect 19416 2384 19482 2474
rect 19416 2320 19417 2384
rect 19481 2320 19482 2384
rect 19416 2304 19482 2320
rect 19416 2240 19417 2304
rect 19481 2240 19482 2304
rect 19416 2224 19482 2240
rect 19416 2160 19417 2224
rect 19481 2160 19482 2224
rect 19416 2144 19482 2160
rect 19416 2080 19417 2144
rect 19481 2080 19482 2144
rect 19416 2064 19482 2080
rect 19416 2000 19417 2064
rect 19481 2000 19482 2064
rect 19416 1984 19482 2000
rect 19416 1920 19417 1984
rect 19481 1920 19482 1984
rect 19416 1904 19482 1920
rect 19416 1840 19417 1904
rect 19481 1840 19482 1904
rect 19416 1824 19482 1840
rect 19416 1760 19417 1824
rect 19481 1760 19482 1824
rect 19416 1744 19482 1760
rect 19416 1680 19417 1744
rect 19481 1680 19482 1744
rect 19416 1664 19482 1680
rect 19416 1600 19417 1664
rect 19481 1600 19482 1664
rect 19416 1446 19482 1600
rect 19542 1508 19602 2538
rect 19662 1446 19722 2478
rect 19782 1508 19842 2538
rect 19902 1446 19962 2478
rect 20022 2384 20088 2474
rect 20022 2320 20023 2384
rect 20087 2320 20088 2384
rect 20022 2304 20088 2320
rect 20022 2240 20023 2304
rect 20087 2240 20088 2304
rect 20022 2224 20088 2240
rect 20022 2160 20023 2224
rect 20087 2160 20088 2224
rect 20022 2144 20088 2160
rect 20022 2080 20023 2144
rect 20087 2080 20088 2144
rect 20022 2064 20088 2080
rect 20022 2000 20023 2064
rect 20087 2000 20088 2064
rect 20022 1984 20088 2000
rect 20022 1920 20023 1984
rect 20087 1920 20088 1984
rect 20022 1904 20088 1920
rect 20022 1840 20023 1904
rect 20087 1840 20088 1904
rect 20022 1824 20088 1840
rect 20022 1760 20023 1824
rect 20087 1760 20088 1824
rect 20022 1744 20088 1760
rect 20022 1680 20023 1744
rect 20087 1680 20088 1744
rect 20022 1664 20088 1680
rect 20022 1600 20023 1664
rect 20087 1600 20088 1664
rect 20022 1446 20088 1600
rect 10326 1444 20088 1446
rect 10326 1380 10430 1444
rect 10494 1380 10510 1444
rect 10574 1380 10590 1444
rect 10654 1380 10670 1444
rect 10734 1380 10750 1444
rect 10814 1380 10830 1444
rect 10894 1380 11036 1444
rect 11100 1380 11116 1444
rect 11180 1380 11196 1444
rect 11260 1380 11276 1444
rect 11340 1380 11356 1444
rect 11420 1380 11436 1444
rect 11500 1380 11642 1444
rect 11706 1380 11722 1444
rect 11786 1380 11802 1444
rect 11866 1380 11882 1444
rect 11946 1380 11962 1444
rect 12026 1380 12042 1444
rect 12106 1380 12248 1444
rect 12312 1380 12328 1444
rect 12392 1380 12408 1444
rect 12472 1380 12488 1444
rect 12552 1380 12568 1444
rect 12632 1380 12648 1444
rect 12712 1380 12854 1444
rect 12918 1380 12934 1444
rect 12998 1380 13014 1444
rect 13078 1380 13094 1444
rect 13158 1380 13174 1444
rect 13238 1380 13254 1444
rect 13318 1380 13460 1444
rect 13524 1380 13540 1444
rect 13604 1380 13620 1444
rect 13684 1380 13700 1444
rect 13764 1380 13780 1444
rect 13844 1380 13860 1444
rect 13924 1380 14066 1444
rect 14130 1380 14146 1444
rect 14210 1380 14226 1444
rect 14290 1380 14306 1444
rect 14370 1380 14386 1444
rect 14450 1380 14466 1444
rect 14530 1380 14672 1444
rect 14736 1380 14752 1444
rect 14816 1380 14832 1444
rect 14896 1380 14912 1444
rect 14976 1380 14992 1444
rect 15056 1380 15072 1444
rect 15136 1380 15278 1444
rect 15342 1380 15358 1444
rect 15422 1380 15438 1444
rect 15502 1380 15518 1444
rect 15582 1380 15598 1444
rect 15662 1380 15678 1444
rect 15742 1380 15884 1444
rect 15948 1380 15964 1444
rect 16028 1380 16044 1444
rect 16108 1380 16124 1444
rect 16188 1380 16204 1444
rect 16268 1380 16284 1444
rect 16348 1380 16490 1444
rect 16554 1380 16570 1444
rect 16634 1380 16650 1444
rect 16714 1380 16730 1444
rect 16794 1380 16810 1444
rect 16874 1380 16890 1444
rect 16954 1380 17096 1444
rect 17160 1380 17176 1444
rect 17240 1380 17256 1444
rect 17320 1380 17336 1444
rect 17400 1380 17416 1444
rect 17480 1380 17496 1444
rect 17560 1380 17702 1444
rect 17766 1380 17782 1444
rect 17846 1380 17862 1444
rect 17926 1380 17942 1444
rect 18006 1380 18022 1444
rect 18086 1380 18102 1444
rect 18166 1380 18308 1444
rect 18372 1380 18388 1444
rect 18452 1380 18468 1444
rect 18532 1380 18548 1444
rect 18612 1380 18628 1444
rect 18692 1380 18708 1444
rect 18772 1380 18914 1444
rect 18978 1380 18994 1444
rect 19058 1380 19074 1444
rect 19138 1380 19154 1444
rect 19218 1380 19234 1444
rect 19298 1380 19314 1444
rect 19378 1380 19520 1444
rect 19584 1380 19600 1444
rect 19664 1380 19680 1444
rect 19744 1380 19760 1444
rect 19824 1380 19840 1444
rect 19904 1380 19920 1444
rect 19984 1380 20088 1444
rect 10326 1378 20088 1380
rect 10326 1224 10392 1378
rect 10326 1160 10327 1224
rect 10391 1160 10392 1224
rect 10326 1144 10392 1160
rect 10326 1080 10327 1144
rect 10391 1080 10392 1144
rect 10326 1064 10392 1080
rect 10326 1000 10327 1064
rect 10391 1000 10392 1064
rect 10326 984 10392 1000
rect 10326 920 10327 984
rect 10391 920 10392 984
rect 10326 904 10392 920
rect 10326 840 10327 904
rect 10391 840 10392 904
rect 10326 824 10392 840
rect 10326 760 10327 824
rect 10391 760 10392 824
rect 10326 744 10392 760
rect 10326 680 10327 744
rect 10391 680 10392 744
rect 10326 664 10392 680
rect 10326 600 10327 664
rect 10391 600 10392 664
rect 10326 584 10392 600
rect 10326 520 10327 584
rect 10391 520 10392 584
rect 10326 504 10392 520
rect 10326 440 10327 504
rect 10391 440 10392 504
rect 10326 350 10392 440
rect 10452 346 10512 1378
rect 10572 286 10632 1316
rect 10692 346 10752 1378
rect 10812 286 10872 1316
rect 10932 1224 10998 1378
rect 10932 1160 10933 1224
rect 10997 1160 10998 1224
rect 10932 1144 10998 1160
rect 10932 1080 10933 1144
rect 10997 1080 10998 1144
rect 10932 1064 10998 1080
rect 10932 1000 10933 1064
rect 10997 1000 10998 1064
rect 10932 984 10998 1000
rect 10932 920 10933 984
rect 10997 920 10998 984
rect 10932 904 10998 920
rect 10932 840 10933 904
rect 10997 840 10998 904
rect 10932 824 10998 840
rect 10932 760 10933 824
rect 10997 760 10998 824
rect 10932 744 10998 760
rect 10932 680 10933 744
rect 10997 680 10998 744
rect 10932 664 10998 680
rect 10932 600 10933 664
rect 10997 600 10998 664
rect 10932 584 10998 600
rect 10932 520 10933 584
rect 10997 520 10998 584
rect 10932 504 10998 520
rect 10932 440 10933 504
rect 10997 440 10998 504
rect 10932 350 10998 440
rect 11058 346 11118 1378
rect 11178 286 11238 1316
rect 11298 346 11358 1378
rect 11418 286 11478 1316
rect 11538 1224 11604 1378
rect 11538 1160 11539 1224
rect 11603 1160 11604 1224
rect 11538 1144 11604 1160
rect 11538 1080 11539 1144
rect 11603 1080 11604 1144
rect 11538 1064 11604 1080
rect 11538 1000 11539 1064
rect 11603 1000 11604 1064
rect 11538 984 11604 1000
rect 11538 920 11539 984
rect 11603 920 11604 984
rect 11538 904 11604 920
rect 11538 840 11539 904
rect 11603 840 11604 904
rect 11538 824 11604 840
rect 11538 760 11539 824
rect 11603 760 11604 824
rect 11538 744 11604 760
rect 11538 680 11539 744
rect 11603 680 11604 744
rect 11538 664 11604 680
rect 11538 600 11539 664
rect 11603 600 11604 664
rect 11538 584 11604 600
rect 11538 520 11539 584
rect 11603 520 11604 584
rect 11538 504 11604 520
rect 11538 440 11539 504
rect 11603 440 11604 504
rect 11538 350 11604 440
rect 11664 346 11724 1378
rect 11784 286 11844 1316
rect 11904 346 11964 1378
rect 12024 286 12084 1316
rect 12144 1224 12210 1378
rect 12144 1160 12145 1224
rect 12209 1160 12210 1224
rect 12144 1144 12210 1160
rect 12144 1080 12145 1144
rect 12209 1080 12210 1144
rect 12144 1064 12210 1080
rect 12144 1000 12145 1064
rect 12209 1000 12210 1064
rect 12144 984 12210 1000
rect 12144 920 12145 984
rect 12209 920 12210 984
rect 12144 904 12210 920
rect 12144 840 12145 904
rect 12209 840 12210 904
rect 12144 824 12210 840
rect 12144 760 12145 824
rect 12209 760 12210 824
rect 12144 744 12210 760
rect 12144 680 12145 744
rect 12209 680 12210 744
rect 12144 664 12210 680
rect 12144 600 12145 664
rect 12209 600 12210 664
rect 12144 584 12210 600
rect 12144 520 12145 584
rect 12209 520 12210 584
rect 12144 504 12210 520
rect 12144 440 12145 504
rect 12209 440 12210 504
rect 12144 350 12210 440
rect 12270 346 12330 1378
rect 12390 286 12450 1316
rect 12510 346 12570 1378
rect 12630 286 12690 1316
rect 12750 1224 12816 1378
rect 12750 1160 12751 1224
rect 12815 1160 12816 1224
rect 12750 1144 12816 1160
rect 12750 1080 12751 1144
rect 12815 1080 12816 1144
rect 12750 1064 12816 1080
rect 12750 1000 12751 1064
rect 12815 1000 12816 1064
rect 12750 984 12816 1000
rect 12750 920 12751 984
rect 12815 920 12816 984
rect 12750 904 12816 920
rect 12750 840 12751 904
rect 12815 840 12816 904
rect 12750 824 12816 840
rect 12750 760 12751 824
rect 12815 760 12816 824
rect 12750 744 12816 760
rect 12750 680 12751 744
rect 12815 680 12816 744
rect 12750 664 12816 680
rect 12750 600 12751 664
rect 12815 600 12816 664
rect 12750 584 12816 600
rect 12750 520 12751 584
rect 12815 520 12816 584
rect 12750 504 12816 520
rect 12750 440 12751 504
rect 12815 440 12816 504
rect 12750 350 12816 440
rect 12876 346 12936 1378
rect 12996 286 13056 1316
rect 13116 346 13176 1378
rect 13236 286 13296 1316
rect 13356 1224 13422 1378
rect 13356 1160 13357 1224
rect 13421 1160 13422 1224
rect 13356 1144 13422 1160
rect 13356 1080 13357 1144
rect 13421 1080 13422 1144
rect 13356 1064 13422 1080
rect 13356 1000 13357 1064
rect 13421 1000 13422 1064
rect 13356 984 13422 1000
rect 13356 920 13357 984
rect 13421 920 13422 984
rect 13356 904 13422 920
rect 13356 840 13357 904
rect 13421 840 13422 904
rect 13356 824 13422 840
rect 13356 760 13357 824
rect 13421 760 13422 824
rect 13356 744 13422 760
rect 13356 680 13357 744
rect 13421 680 13422 744
rect 13356 664 13422 680
rect 13356 600 13357 664
rect 13421 600 13422 664
rect 13356 584 13422 600
rect 13356 520 13357 584
rect 13421 520 13422 584
rect 13356 504 13422 520
rect 13356 440 13357 504
rect 13421 440 13422 504
rect 13356 350 13422 440
rect 13482 346 13542 1378
rect 13602 286 13662 1316
rect 13722 346 13782 1378
rect 13842 286 13902 1316
rect 13962 1224 14028 1378
rect 13962 1160 13963 1224
rect 14027 1160 14028 1224
rect 13962 1144 14028 1160
rect 13962 1080 13963 1144
rect 14027 1080 14028 1144
rect 13962 1064 14028 1080
rect 13962 1000 13963 1064
rect 14027 1000 14028 1064
rect 13962 984 14028 1000
rect 13962 920 13963 984
rect 14027 920 14028 984
rect 13962 904 14028 920
rect 13962 840 13963 904
rect 14027 840 14028 904
rect 13962 824 14028 840
rect 13962 760 13963 824
rect 14027 760 14028 824
rect 13962 744 14028 760
rect 13962 680 13963 744
rect 14027 680 14028 744
rect 13962 664 14028 680
rect 13962 600 13963 664
rect 14027 600 14028 664
rect 13962 584 14028 600
rect 13962 520 13963 584
rect 14027 520 14028 584
rect 13962 504 14028 520
rect 13962 440 13963 504
rect 14027 440 14028 504
rect 13962 350 14028 440
rect 14088 346 14148 1378
rect 14208 286 14268 1316
rect 14328 346 14388 1378
rect 14448 286 14508 1316
rect 14568 1224 14634 1378
rect 14568 1160 14569 1224
rect 14633 1160 14634 1224
rect 14568 1144 14634 1160
rect 14568 1080 14569 1144
rect 14633 1080 14634 1144
rect 14568 1064 14634 1080
rect 14568 1000 14569 1064
rect 14633 1000 14634 1064
rect 14568 984 14634 1000
rect 14568 920 14569 984
rect 14633 920 14634 984
rect 14568 904 14634 920
rect 14568 840 14569 904
rect 14633 840 14634 904
rect 14568 824 14634 840
rect 14568 760 14569 824
rect 14633 760 14634 824
rect 14568 744 14634 760
rect 14568 680 14569 744
rect 14633 680 14634 744
rect 14568 664 14634 680
rect 14568 600 14569 664
rect 14633 600 14634 664
rect 14568 584 14634 600
rect 14568 520 14569 584
rect 14633 520 14634 584
rect 14568 504 14634 520
rect 14568 440 14569 504
rect 14633 440 14634 504
rect 14568 350 14634 440
rect 14694 346 14754 1378
rect 14814 286 14874 1316
rect 14934 346 14994 1378
rect 15054 286 15114 1316
rect 15174 1224 15240 1378
rect 15174 1160 15175 1224
rect 15239 1160 15240 1224
rect 15174 1144 15240 1160
rect 15174 1080 15175 1144
rect 15239 1080 15240 1144
rect 15174 1064 15240 1080
rect 15174 1000 15175 1064
rect 15239 1000 15240 1064
rect 15174 984 15240 1000
rect 15174 920 15175 984
rect 15239 920 15240 984
rect 15174 904 15240 920
rect 15174 840 15175 904
rect 15239 840 15240 904
rect 15174 824 15240 840
rect 15174 760 15175 824
rect 15239 760 15240 824
rect 15174 744 15240 760
rect 15174 680 15175 744
rect 15239 680 15240 744
rect 15174 664 15240 680
rect 15174 600 15175 664
rect 15239 600 15240 664
rect 15174 584 15240 600
rect 15174 520 15175 584
rect 15239 520 15240 584
rect 15174 504 15240 520
rect 15174 440 15175 504
rect 15239 440 15240 504
rect 15174 350 15240 440
rect 15300 346 15360 1378
rect 15420 286 15480 1316
rect 15540 346 15600 1378
rect 15660 286 15720 1316
rect 15780 1224 15846 1378
rect 15780 1160 15781 1224
rect 15845 1160 15846 1224
rect 15780 1144 15846 1160
rect 15780 1080 15781 1144
rect 15845 1080 15846 1144
rect 15780 1064 15846 1080
rect 15780 1000 15781 1064
rect 15845 1000 15846 1064
rect 15780 984 15846 1000
rect 15780 920 15781 984
rect 15845 920 15846 984
rect 15780 904 15846 920
rect 15780 840 15781 904
rect 15845 840 15846 904
rect 15780 824 15846 840
rect 15780 760 15781 824
rect 15845 760 15846 824
rect 15780 744 15846 760
rect 15780 680 15781 744
rect 15845 680 15846 744
rect 15780 664 15846 680
rect 15780 600 15781 664
rect 15845 600 15846 664
rect 15780 584 15846 600
rect 15780 520 15781 584
rect 15845 520 15846 584
rect 15780 504 15846 520
rect 15780 440 15781 504
rect 15845 440 15846 504
rect 15780 350 15846 440
rect 15906 346 15966 1378
rect 16026 286 16086 1316
rect 16146 346 16206 1378
rect 16266 286 16326 1316
rect 16386 1224 16452 1378
rect 16386 1160 16387 1224
rect 16451 1160 16452 1224
rect 16386 1144 16452 1160
rect 16386 1080 16387 1144
rect 16451 1080 16452 1144
rect 16386 1064 16452 1080
rect 16386 1000 16387 1064
rect 16451 1000 16452 1064
rect 16386 984 16452 1000
rect 16386 920 16387 984
rect 16451 920 16452 984
rect 16386 904 16452 920
rect 16386 840 16387 904
rect 16451 840 16452 904
rect 16386 824 16452 840
rect 16386 760 16387 824
rect 16451 760 16452 824
rect 16386 744 16452 760
rect 16386 680 16387 744
rect 16451 680 16452 744
rect 16386 664 16452 680
rect 16386 600 16387 664
rect 16451 600 16452 664
rect 16386 584 16452 600
rect 16386 520 16387 584
rect 16451 520 16452 584
rect 16386 504 16452 520
rect 16386 440 16387 504
rect 16451 440 16452 504
rect 16386 350 16452 440
rect 16512 346 16572 1378
rect 16632 286 16692 1316
rect 16752 346 16812 1378
rect 16872 286 16932 1316
rect 16992 1224 17058 1378
rect 16992 1160 16993 1224
rect 17057 1160 17058 1224
rect 16992 1144 17058 1160
rect 16992 1080 16993 1144
rect 17057 1080 17058 1144
rect 16992 1064 17058 1080
rect 16992 1000 16993 1064
rect 17057 1000 17058 1064
rect 16992 984 17058 1000
rect 16992 920 16993 984
rect 17057 920 17058 984
rect 16992 904 17058 920
rect 16992 840 16993 904
rect 17057 840 17058 904
rect 16992 824 17058 840
rect 16992 760 16993 824
rect 17057 760 17058 824
rect 16992 744 17058 760
rect 16992 680 16993 744
rect 17057 680 17058 744
rect 16992 664 17058 680
rect 16992 600 16993 664
rect 17057 600 17058 664
rect 16992 584 17058 600
rect 16992 520 16993 584
rect 17057 520 17058 584
rect 16992 504 17058 520
rect 16992 440 16993 504
rect 17057 440 17058 504
rect 16992 350 17058 440
rect 17118 346 17178 1378
rect 17238 286 17298 1316
rect 17358 346 17418 1378
rect 17478 286 17538 1316
rect 17598 1224 17664 1378
rect 17598 1160 17599 1224
rect 17663 1160 17664 1224
rect 17598 1144 17664 1160
rect 17598 1080 17599 1144
rect 17663 1080 17664 1144
rect 17598 1064 17664 1080
rect 17598 1000 17599 1064
rect 17663 1000 17664 1064
rect 17598 984 17664 1000
rect 17598 920 17599 984
rect 17663 920 17664 984
rect 17598 904 17664 920
rect 17598 840 17599 904
rect 17663 840 17664 904
rect 17598 824 17664 840
rect 17598 760 17599 824
rect 17663 760 17664 824
rect 17598 744 17664 760
rect 17598 680 17599 744
rect 17663 680 17664 744
rect 17598 664 17664 680
rect 17598 600 17599 664
rect 17663 600 17664 664
rect 17598 584 17664 600
rect 17598 520 17599 584
rect 17663 520 17664 584
rect 17598 504 17664 520
rect 17598 440 17599 504
rect 17663 440 17664 504
rect 17598 350 17664 440
rect 17724 346 17784 1378
rect 17844 286 17904 1316
rect 17964 346 18024 1378
rect 18084 286 18144 1316
rect 18204 1224 18270 1378
rect 18204 1160 18205 1224
rect 18269 1160 18270 1224
rect 18204 1144 18270 1160
rect 18204 1080 18205 1144
rect 18269 1080 18270 1144
rect 18204 1064 18270 1080
rect 18204 1000 18205 1064
rect 18269 1000 18270 1064
rect 18204 984 18270 1000
rect 18204 920 18205 984
rect 18269 920 18270 984
rect 18204 904 18270 920
rect 18204 840 18205 904
rect 18269 840 18270 904
rect 18204 824 18270 840
rect 18204 760 18205 824
rect 18269 760 18270 824
rect 18204 744 18270 760
rect 18204 680 18205 744
rect 18269 680 18270 744
rect 18204 664 18270 680
rect 18204 600 18205 664
rect 18269 600 18270 664
rect 18204 584 18270 600
rect 18204 520 18205 584
rect 18269 520 18270 584
rect 18204 504 18270 520
rect 18204 440 18205 504
rect 18269 440 18270 504
rect 18204 350 18270 440
rect 18330 346 18390 1378
rect 18450 286 18510 1316
rect 18570 346 18630 1378
rect 18690 286 18750 1316
rect 18810 1224 18876 1378
rect 18810 1160 18811 1224
rect 18875 1160 18876 1224
rect 18810 1144 18876 1160
rect 18810 1080 18811 1144
rect 18875 1080 18876 1144
rect 18810 1064 18876 1080
rect 18810 1000 18811 1064
rect 18875 1000 18876 1064
rect 18810 984 18876 1000
rect 18810 920 18811 984
rect 18875 920 18876 984
rect 18810 904 18876 920
rect 18810 840 18811 904
rect 18875 840 18876 904
rect 18810 824 18876 840
rect 18810 760 18811 824
rect 18875 760 18876 824
rect 18810 744 18876 760
rect 18810 680 18811 744
rect 18875 680 18876 744
rect 18810 664 18876 680
rect 18810 600 18811 664
rect 18875 600 18876 664
rect 18810 584 18876 600
rect 18810 520 18811 584
rect 18875 520 18876 584
rect 18810 504 18876 520
rect 18810 440 18811 504
rect 18875 440 18876 504
rect 18810 350 18876 440
rect 18936 346 18996 1378
rect 19056 286 19116 1316
rect 19176 346 19236 1378
rect 19296 286 19356 1316
rect 19416 1224 19482 1378
rect 19416 1160 19417 1224
rect 19481 1160 19482 1224
rect 19416 1144 19482 1160
rect 19416 1080 19417 1144
rect 19481 1080 19482 1144
rect 19416 1064 19482 1080
rect 19416 1000 19417 1064
rect 19481 1000 19482 1064
rect 19416 984 19482 1000
rect 19416 920 19417 984
rect 19481 920 19482 984
rect 19416 904 19482 920
rect 19416 840 19417 904
rect 19481 840 19482 904
rect 19416 824 19482 840
rect 19416 760 19417 824
rect 19481 760 19482 824
rect 19416 744 19482 760
rect 19416 680 19417 744
rect 19481 680 19482 744
rect 19416 664 19482 680
rect 19416 600 19417 664
rect 19481 600 19482 664
rect 19416 584 19482 600
rect 19416 520 19417 584
rect 19481 520 19482 584
rect 19416 504 19482 520
rect 19416 440 19417 504
rect 19481 440 19482 504
rect 19416 350 19482 440
rect 19542 346 19602 1378
rect 19662 286 19722 1316
rect 19782 346 19842 1378
rect 19902 286 19962 1316
rect 20022 1224 20088 1378
rect 20022 1160 20023 1224
rect 20087 1160 20088 1224
rect 20022 1144 20088 1160
rect 20022 1080 20023 1144
rect 20087 1080 20088 1144
rect 20022 1064 20088 1080
rect 20022 1000 20023 1064
rect 20087 1000 20088 1064
rect 20022 984 20088 1000
rect 20022 920 20023 984
rect 20087 920 20088 984
rect 20022 904 20088 920
rect 20022 840 20023 904
rect 20087 840 20088 904
rect 20022 824 20088 840
rect 20022 760 20023 824
rect 20087 760 20088 824
rect 20022 744 20088 760
rect 20022 680 20023 744
rect 20087 680 20088 744
rect 20022 664 20088 680
rect 20022 600 20023 664
rect 20087 600 20088 664
rect 20022 584 20088 600
rect 20022 520 20023 584
rect 20087 520 20088 584
rect 20022 504 20088 520
rect 20022 440 20023 504
rect 20087 440 20088 504
rect 20022 350 20088 440
rect 20148 2384 20214 2475
rect 20148 2320 20149 2384
rect 20213 2320 20214 2384
rect 20148 2304 20214 2320
rect 20148 2240 20149 2304
rect 20213 2240 20214 2304
rect 20148 2224 20214 2240
rect 20148 2160 20149 2224
rect 20213 2160 20214 2224
rect 20148 2144 20214 2160
rect 20148 2080 20149 2144
rect 20213 2080 20214 2144
rect 20148 2064 20214 2080
rect 20148 2000 20149 2064
rect 20213 2000 20214 2064
rect 20148 1984 20214 2000
rect 20148 1920 20149 1984
rect 20213 1920 20214 1984
rect 20148 1904 20214 1920
rect 20148 1840 20149 1904
rect 20213 1840 20214 1904
rect 20148 1824 20214 1840
rect 20148 1760 20149 1824
rect 20213 1760 20214 1824
rect 20148 1744 20214 1760
rect 20148 1680 20149 1744
rect 20213 1680 20214 1744
rect 20148 1664 20214 1680
rect 20148 1600 20149 1664
rect 20213 1600 20214 1664
rect 20148 1446 20214 1600
rect 20274 1508 20334 2538
rect 20394 1446 20454 2478
rect 20514 1508 20574 2538
rect 20634 1446 20694 2478
rect 20754 2384 20820 2474
rect 20754 2320 20755 2384
rect 20819 2320 20820 2384
rect 20754 2304 20820 2320
rect 20754 2240 20755 2304
rect 20819 2240 20820 2304
rect 20754 2224 20820 2240
rect 20754 2160 20755 2224
rect 20819 2160 20820 2224
rect 20754 2144 20820 2160
rect 20754 2080 20755 2144
rect 20819 2080 20820 2144
rect 20754 2064 20820 2080
rect 20754 2000 20755 2064
rect 20819 2000 20820 2064
rect 20754 1984 20820 2000
rect 20754 1920 20755 1984
rect 20819 1920 20820 1984
rect 20754 1904 20820 1920
rect 20754 1840 20755 1904
rect 20819 1840 20820 1904
rect 20754 1824 20820 1840
rect 20754 1760 20755 1824
rect 20819 1760 20820 1824
rect 20754 1744 20820 1760
rect 20754 1680 20755 1744
rect 20819 1680 20820 1744
rect 20754 1664 20820 1680
rect 20754 1600 20755 1664
rect 20819 1600 20820 1664
rect 20754 1446 20820 1600
rect 20880 1508 20940 2538
rect 21000 1446 21060 2478
rect 21120 1508 21180 2538
rect 21240 1446 21300 2478
rect 21360 2384 21426 2474
rect 21360 2320 21361 2384
rect 21425 2320 21426 2384
rect 21360 2304 21426 2320
rect 21360 2240 21361 2304
rect 21425 2240 21426 2304
rect 21360 2224 21426 2240
rect 21360 2160 21361 2224
rect 21425 2160 21426 2224
rect 21360 2144 21426 2160
rect 21360 2080 21361 2144
rect 21425 2080 21426 2144
rect 21360 2064 21426 2080
rect 21360 2000 21361 2064
rect 21425 2000 21426 2064
rect 21360 1984 21426 2000
rect 21360 1920 21361 1984
rect 21425 1920 21426 1984
rect 21360 1904 21426 1920
rect 21360 1840 21361 1904
rect 21425 1840 21426 1904
rect 21360 1824 21426 1840
rect 21360 1760 21361 1824
rect 21425 1760 21426 1824
rect 21360 1744 21426 1760
rect 21360 1680 21361 1744
rect 21425 1680 21426 1744
rect 21360 1664 21426 1680
rect 21360 1600 21361 1664
rect 21425 1600 21426 1664
rect 21360 1446 21426 1600
rect 21486 1508 21546 2538
rect 21606 1446 21666 2478
rect 21726 1508 21786 2538
rect 21846 1446 21906 2478
rect 21966 2384 22032 2474
rect 21966 2320 21967 2384
rect 22031 2320 22032 2384
rect 21966 2304 22032 2320
rect 21966 2240 21967 2304
rect 22031 2240 22032 2304
rect 21966 2224 22032 2240
rect 21966 2160 21967 2224
rect 22031 2160 22032 2224
rect 21966 2144 22032 2160
rect 21966 2080 21967 2144
rect 22031 2080 22032 2144
rect 21966 2064 22032 2080
rect 21966 2000 21967 2064
rect 22031 2000 22032 2064
rect 21966 1984 22032 2000
rect 21966 1920 21967 1984
rect 22031 1920 22032 1984
rect 21966 1904 22032 1920
rect 21966 1840 21967 1904
rect 22031 1840 22032 1904
rect 21966 1824 22032 1840
rect 21966 1760 21967 1824
rect 22031 1760 22032 1824
rect 21966 1744 22032 1760
rect 21966 1680 21967 1744
rect 22031 1680 22032 1744
rect 21966 1664 22032 1680
rect 21966 1600 21967 1664
rect 22031 1600 22032 1664
rect 21966 1446 22032 1600
rect 22092 1508 22152 2538
rect 22212 1446 22272 2478
rect 22332 1508 22392 2538
rect 22452 1446 22512 2478
rect 22572 2384 22638 2474
rect 22572 2320 22573 2384
rect 22637 2320 22638 2384
rect 22572 2304 22638 2320
rect 22572 2240 22573 2304
rect 22637 2240 22638 2304
rect 22572 2224 22638 2240
rect 22572 2160 22573 2224
rect 22637 2160 22638 2224
rect 22572 2144 22638 2160
rect 22572 2080 22573 2144
rect 22637 2080 22638 2144
rect 22572 2064 22638 2080
rect 22572 2000 22573 2064
rect 22637 2000 22638 2064
rect 22572 1984 22638 2000
rect 22572 1920 22573 1984
rect 22637 1920 22638 1984
rect 22572 1904 22638 1920
rect 22572 1840 22573 1904
rect 22637 1840 22638 1904
rect 22572 1824 22638 1840
rect 22572 1760 22573 1824
rect 22637 1760 22638 1824
rect 22572 1744 22638 1760
rect 22572 1680 22573 1744
rect 22637 1680 22638 1744
rect 22572 1664 22638 1680
rect 22572 1600 22573 1664
rect 22637 1600 22638 1664
rect 22572 1446 22638 1600
rect 22698 1508 22758 2538
rect 22818 1446 22878 2478
rect 22938 1508 22998 2538
rect 23058 1446 23118 2478
rect 23178 2384 23244 2474
rect 23178 2320 23179 2384
rect 23243 2320 23244 2384
rect 23178 2304 23244 2320
rect 23178 2240 23179 2304
rect 23243 2240 23244 2304
rect 23178 2224 23244 2240
rect 23178 2160 23179 2224
rect 23243 2160 23244 2224
rect 23178 2144 23244 2160
rect 23178 2080 23179 2144
rect 23243 2080 23244 2144
rect 23178 2064 23244 2080
rect 23178 2000 23179 2064
rect 23243 2000 23244 2064
rect 23178 1984 23244 2000
rect 23178 1920 23179 1984
rect 23243 1920 23244 1984
rect 23178 1904 23244 1920
rect 23178 1840 23179 1904
rect 23243 1840 23244 1904
rect 23178 1824 23244 1840
rect 23178 1760 23179 1824
rect 23243 1760 23244 1824
rect 23178 1744 23244 1760
rect 23178 1680 23179 1744
rect 23243 1680 23244 1744
rect 23178 1664 23244 1680
rect 23178 1600 23179 1664
rect 23243 1600 23244 1664
rect 23178 1446 23244 1600
rect 23304 1508 23364 2538
rect 23424 1446 23484 2478
rect 23544 1508 23604 2538
rect 23664 1446 23724 2478
rect 23784 2384 23850 2474
rect 23784 2320 23785 2384
rect 23849 2320 23850 2384
rect 23784 2304 23850 2320
rect 23784 2240 23785 2304
rect 23849 2240 23850 2304
rect 23784 2224 23850 2240
rect 23784 2160 23785 2224
rect 23849 2160 23850 2224
rect 23784 2144 23850 2160
rect 23784 2080 23785 2144
rect 23849 2080 23850 2144
rect 23784 2064 23850 2080
rect 23784 2000 23785 2064
rect 23849 2000 23850 2064
rect 23784 1984 23850 2000
rect 23784 1920 23785 1984
rect 23849 1920 23850 1984
rect 23784 1904 23850 1920
rect 23784 1840 23785 1904
rect 23849 1840 23850 1904
rect 23784 1824 23850 1840
rect 23784 1760 23785 1824
rect 23849 1760 23850 1824
rect 23784 1744 23850 1760
rect 23784 1680 23785 1744
rect 23849 1680 23850 1744
rect 23784 1664 23850 1680
rect 23784 1600 23785 1664
rect 23849 1600 23850 1664
rect 23784 1446 23850 1600
rect 23910 1508 23970 2538
rect 24030 1446 24090 2478
rect 24150 1508 24210 2538
rect 24270 1446 24330 2478
rect 24390 2384 24456 2474
rect 24390 2320 24391 2384
rect 24455 2320 24456 2384
rect 24390 2304 24456 2320
rect 24390 2240 24391 2304
rect 24455 2240 24456 2304
rect 24390 2224 24456 2240
rect 24390 2160 24391 2224
rect 24455 2160 24456 2224
rect 24390 2144 24456 2160
rect 24390 2080 24391 2144
rect 24455 2080 24456 2144
rect 24390 2064 24456 2080
rect 24390 2000 24391 2064
rect 24455 2000 24456 2064
rect 24390 1984 24456 2000
rect 24390 1920 24391 1984
rect 24455 1920 24456 1984
rect 24390 1904 24456 1920
rect 24390 1840 24391 1904
rect 24455 1840 24456 1904
rect 24390 1824 24456 1840
rect 24390 1760 24391 1824
rect 24455 1760 24456 1824
rect 24390 1744 24456 1760
rect 24390 1680 24391 1744
rect 24455 1680 24456 1744
rect 24390 1664 24456 1680
rect 24390 1600 24391 1664
rect 24455 1600 24456 1664
rect 24390 1446 24456 1600
rect 24516 1508 24576 2538
rect 24636 1446 24696 2478
rect 24756 1508 24816 2538
rect 24876 1446 24936 2478
rect 24996 2384 25062 2474
rect 24996 2320 24997 2384
rect 25061 2320 25062 2384
rect 24996 2304 25062 2320
rect 24996 2240 24997 2304
rect 25061 2240 25062 2304
rect 24996 2224 25062 2240
rect 24996 2160 24997 2224
rect 25061 2160 25062 2224
rect 24996 2144 25062 2160
rect 24996 2080 24997 2144
rect 25061 2080 25062 2144
rect 24996 2064 25062 2080
rect 24996 2000 24997 2064
rect 25061 2000 25062 2064
rect 24996 1984 25062 2000
rect 24996 1920 24997 1984
rect 25061 1920 25062 1984
rect 24996 1904 25062 1920
rect 24996 1840 24997 1904
rect 25061 1840 25062 1904
rect 24996 1824 25062 1840
rect 24996 1760 24997 1824
rect 25061 1760 25062 1824
rect 24996 1744 25062 1760
rect 24996 1680 24997 1744
rect 25061 1680 25062 1744
rect 24996 1664 25062 1680
rect 24996 1600 24997 1664
rect 25061 1600 25062 1664
rect 24996 1446 25062 1600
rect 25122 1508 25182 2538
rect 25242 1446 25302 2478
rect 25362 1508 25422 2538
rect 25482 1446 25542 2478
rect 25602 2384 25668 2474
rect 25602 2320 25603 2384
rect 25667 2320 25668 2384
rect 25602 2304 25668 2320
rect 25602 2240 25603 2304
rect 25667 2240 25668 2304
rect 25602 2224 25668 2240
rect 25602 2160 25603 2224
rect 25667 2160 25668 2224
rect 25602 2144 25668 2160
rect 25602 2080 25603 2144
rect 25667 2080 25668 2144
rect 25602 2064 25668 2080
rect 25602 2000 25603 2064
rect 25667 2000 25668 2064
rect 25602 1984 25668 2000
rect 25602 1920 25603 1984
rect 25667 1920 25668 1984
rect 25602 1904 25668 1920
rect 25602 1840 25603 1904
rect 25667 1840 25668 1904
rect 25602 1824 25668 1840
rect 25602 1760 25603 1824
rect 25667 1760 25668 1824
rect 25602 1744 25668 1760
rect 25602 1680 25603 1744
rect 25667 1680 25668 1744
rect 25602 1664 25668 1680
rect 25602 1600 25603 1664
rect 25667 1600 25668 1664
rect 25602 1446 25668 1600
rect 25728 1508 25788 2538
rect 25848 1446 25908 2478
rect 25968 1508 26028 2538
rect 26088 1446 26148 2478
rect 26208 2384 26274 2474
rect 26208 2320 26209 2384
rect 26273 2320 26274 2384
rect 26208 2304 26274 2320
rect 26208 2240 26209 2304
rect 26273 2240 26274 2304
rect 26208 2224 26274 2240
rect 26208 2160 26209 2224
rect 26273 2160 26274 2224
rect 26208 2144 26274 2160
rect 26208 2080 26209 2144
rect 26273 2080 26274 2144
rect 26208 2064 26274 2080
rect 26208 2000 26209 2064
rect 26273 2000 26274 2064
rect 26208 1984 26274 2000
rect 26208 1920 26209 1984
rect 26273 1920 26274 1984
rect 26208 1904 26274 1920
rect 26208 1840 26209 1904
rect 26273 1840 26274 1904
rect 26208 1824 26274 1840
rect 26208 1760 26209 1824
rect 26273 1760 26274 1824
rect 26208 1744 26274 1760
rect 26208 1680 26209 1744
rect 26273 1680 26274 1744
rect 26208 1664 26274 1680
rect 26208 1600 26209 1664
rect 26273 1600 26274 1664
rect 26208 1446 26274 1600
rect 26334 1508 26394 2538
rect 26454 1446 26514 2478
rect 26574 1508 26634 2538
rect 26694 1446 26754 2478
rect 26814 2384 26880 2474
rect 26814 2320 26815 2384
rect 26879 2320 26880 2384
rect 26814 2304 26880 2320
rect 26814 2240 26815 2304
rect 26879 2240 26880 2304
rect 26814 2224 26880 2240
rect 26814 2160 26815 2224
rect 26879 2160 26880 2224
rect 26814 2144 26880 2160
rect 26814 2080 26815 2144
rect 26879 2080 26880 2144
rect 26814 2064 26880 2080
rect 26814 2000 26815 2064
rect 26879 2000 26880 2064
rect 26814 1984 26880 2000
rect 26814 1920 26815 1984
rect 26879 1920 26880 1984
rect 26814 1904 26880 1920
rect 26814 1840 26815 1904
rect 26879 1840 26880 1904
rect 26814 1824 26880 1840
rect 26814 1760 26815 1824
rect 26879 1760 26880 1824
rect 26814 1744 26880 1760
rect 26814 1680 26815 1744
rect 26879 1680 26880 1744
rect 26814 1664 26880 1680
rect 26814 1600 26815 1664
rect 26879 1600 26880 1664
rect 26814 1446 26880 1600
rect 26940 1508 27000 2538
rect 27060 1446 27120 2478
rect 27180 1508 27240 2538
rect 27300 1446 27360 2478
rect 27420 2384 27486 2474
rect 27420 2320 27421 2384
rect 27485 2320 27486 2384
rect 27420 2304 27486 2320
rect 27420 2240 27421 2304
rect 27485 2240 27486 2304
rect 27420 2224 27486 2240
rect 27420 2160 27421 2224
rect 27485 2160 27486 2224
rect 27420 2144 27486 2160
rect 27420 2080 27421 2144
rect 27485 2080 27486 2144
rect 27420 2064 27486 2080
rect 27420 2000 27421 2064
rect 27485 2000 27486 2064
rect 27420 1984 27486 2000
rect 27420 1920 27421 1984
rect 27485 1920 27486 1984
rect 27420 1904 27486 1920
rect 27420 1840 27421 1904
rect 27485 1840 27486 1904
rect 27420 1824 27486 1840
rect 27420 1760 27421 1824
rect 27485 1760 27486 1824
rect 27420 1744 27486 1760
rect 27420 1680 27421 1744
rect 27485 1680 27486 1744
rect 27420 1664 27486 1680
rect 27420 1600 27421 1664
rect 27485 1600 27486 1664
rect 27420 1446 27486 1600
rect 27546 1508 27606 2538
rect 27666 1446 27726 2478
rect 27786 1508 27846 2538
rect 27906 1446 27966 2478
rect 28026 2384 28092 2474
rect 28026 2320 28027 2384
rect 28091 2320 28092 2384
rect 28026 2304 28092 2320
rect 28026 2240 28027 2304
rect 28091 2240 28092 2304
rect 28026 2224 28092 2240
rect 28026 2160 28027 2224
rect 28091 2160 28092 2224
rect 28026 2144 28092 2160
rect 28026 2080 28027 2144
rect 28091 2080 28092 2144
rect 28026 2064 28092 2080
rect 28026 2000 28027 2064
rect 28091 2000 28092 2064
rect 28026 1984 28092 2000
rect 28026 1920 28027 1984
rect 28091 1920 28092 1984
rect 28026 1904 28092 1920
rect 28026 1840 28027 1904
rect 28091 1840 28092 1904
rect 28026 1824 28092 1840
rect 28026 1760 28027 1824
rect 28091 1760 28092 1824
rect 28026 1744 28092 1760
rect 28026 1680 28027 1744
rect 28091 1680 28092 1744
rect 28026 1664 28092 1680
rect 28026 1600 28027 1664
rect 28091 1600 28092 1664
rect 28026 1446 28092 1600
rect 28152 1508 28212 2538
rect 28272 1446 28332 2478
rect 28392 1508 28452 2538
rect 28512 1446 28572 2478
rect 28632 2384 28698 2474
rect 28632 2320 28633 2384
rect 28697 2320 28698 2384
rect 28632 2304 28698 2320
rect 28632 2240 28633 2304
rect 28697 2240 28698 2304
rect 28632 2224 28698 2240
rect 28632 2160 28633 2224
rect 28697 2160 28698 2224
rect 28632 2144 28698 2160
rect 28632 2080 28633 2144
rect 28697 2080 28698 2144
rect 28632 2064 28698 2080
rect 28632 2000 28633 2064
rect 28697 2000 28698 2064
rect 28632 1984 28698 2000
rect 28632 1920 28633 1984
rect 28697 1920 28698 1984
rect 28632 1904 28698 1920
rect 28632 1840 28633 1904
rect 28697 1840 28698 1904
rect 28632 1824 28698 1840
rect 28632 1760 28633 1824
rect 28697 1760 28698 1824
rect 28632 1744 28698 1760
rect 28632 1680 28633 1744
rect 28697 1680 28698 1744
rect 28632 1664 28698 1680
rect 28632 1600 28633 1664
rect 28697 1600 28698 1664
rect 28632 1446 28698 1600
rect 28758 1508 28818 2538
rect 28878 1446 28938 2478
rect 28998 1508 29058 2538
rect 29118 1446 29178 2478
rect 29238 2384 29304 2474
rect 29238 2320 29239 2384
rect 29303 2320 29304 2384
rect 29238 2304 29304 2320
rect 29238 2240 29239 2304
rect 29303 2240 29304 2304
rect 29238 2224 29304 2240
rect 29238 2160 29239 2224
rect 29303 2160 29304 2224
rect 29238 2144 29304 2160
rect 29238 2080 29239 2144
rect 29303 2080 29304 2144
rect 29238 2064 29304 2080
rect 29238 2000 29239 2064
rect 29303 2000 29304 2064
rect 29238 1984 29304 2000
rect 29238 1920 29239 1984
rect 29303 1920 29304 1984
rect 29238 1904 29304 1920
rect 29238 1840 29239 1904
rect 29303 1840 29304 1904
rect 29238 1824 29304 1840
rect 29238 1760 29239 1824
rect 29303 1760 29304 1824
rect 29238 1744 29304 1760
rect 29238 1680 29239 1744
rect 29303 1680 29304 1744
rect 29238 1664 29304 1680
rect 29238 1600 29239 1664
rect 29303 1600 29304 1664
rect 29238 1446 29304 1600
rect 29364 1508 29424 2538
rect 29484 1446 29544 2478
rect 29604 1508 29664 2538
rect 29724 1446 29784 2478
rect 29844 2384 29910 2474
rect 29844 2320 29845 2384
rect 29909 2320 29910 2384
rect 29844 2304 29910 2320
rect 29844 2240 29845 2304
rect 29909 2240 29910 2304
rect 29844 2224 29910 2240
rect 29844 2160 29845 2224
rect 29909 2160 29910 2224
rect 29844 2144 29910 2160
rect 29844 2080 29845 2144
rect 29909 2080 29910 2144
rect 29844 2064 29910 2080
rect 29844 2000 29845 2064
rect 29909 2000 29910 2064
rect 29844 1984 29910 2000
rect 29844 1920 29845 1984
rect 29909 1920 29910 1984
rect 29844 1904 29910 1920
rect 29844 1840 29845 1904
rect 29909 1840 29910 1904
rect 29844 1824 29910 1840
rect 29844 1760 29845 1824
rect 29909 1760 29910 1824
rect 29844 1744 29910 1760
rect 29844 1680 29845 1744
rect 29909 1680 29910 1744
rect 29844 1664 29910 1680
rect 29844 1600 29845 1664
rect 29909 1600 29910 1664
rect 29844 1446 29910 1600
rect 29970 1508 30030 2538
rect 30090 1446 30150 2478
rect 30210 1508 30270 2538
rect 30330 1446 30390 2478
rect 30450 2384 30516 2474
rect 30450 2320 30451 2384
rect 30515 2320 30516 2384
rect 30450 2304 30516 2320
rect 30450 2240 30451 2304
rect 30515 2240 30516 2304
rect 30450 2224 30516 2240
rect 30450 2160 30451 2224
rect 30515 2160 30516 2224
rect 30450 2144 30516 2160
rect 30450 2080 30451 2144
rect 30515 2080 30516 2144
rect 30450 2064 30516 2080
rect 30450 2000 30451 2064
rect 30515 2000 30516 2064
rect 30450 1984 30516 2000
rect 30450 1920 30451 1984
rect 30515 1920 30516 1984
rect 30450 1904 30516 1920
rect 30450 1840 30451 1904
rect 30515 1840 30516 1904
rect 30450 1824 30516 1840
rect 30450 1760 30451 1824
rect 30515 1760 30516 1824
rect 30450 1744 30516 1760
rect 30450 1680 30451 1744
rect 30515 1680 30516 1744
rect 30450 1664 30516 1680
rect 30450 1600 30451 1664
rect 30515 1600 30516 1664
rect 30450 1446 30516 1600
rect 30576 1508 30636 2538
rect 30696 1446 30756 2478
rect 30816 1508 30876 2538
rect 30936 1446 30996 2478
rect 31056 2384 31122 2474
rect 31056 2320 31057 2384
rect 31121 2320 31122 2384
rect 31056 2304 31122 2320
rect 31056 2240 31057 2304
rect 31121 2240 31122 2304
rect 31056 2224 31122 2240
rect 31056 2160 31057 2224
rect 31121 2160 31122 2224
rect 31056 2144 31122 2160
rect 31056 2080 31057 2144
rect 31121 2080 31122 2144
rect 31056 2064 31122 2080
rect 31056 2000 31057 2064
rect 31121 2000 31122 2064
rect 31056 1984 31122 2000
rect 31056 1920 31057 1984
rect 31121 1920 31122 1984
rect 31056 1904 31122 1920
rect 31056 1840 31057 1904
rect 31121 1840 31122 1904
rect 31056 1824 31122 1840
rect 31056 1760 31057 1824
rect 31121 1760 31122 1824
rect 31056 1744 31122 1760
rect 31056 1680 31057 1744
rect 31121 1680 31122 1744
rect 31056 1664 31122 1680
rect 31056 1600 31057 1664
rect 31121 1600 31122 1664
rect 31056 1446 31122 1600
rect 31182 1508 31242 2538
rect 31302 1446 31362 2478
rect 31422 1508 31482 2538
rect 31542 1446 31602 2478
rect 31662 2384 31728 2474
rect 31662 2320 31663 2384
rect 31727 2320 31728 2384
rect 31662 2304 31728 2320
rect 31662 2240 31663 2304
rect 31727 2240 31728 2304
rect 31662 2224 31728 2240
rect 31662 2160 31663 2224
rect 31727 2160 31728 2224
rect 31662 2144 31728 2160
rect 31662 2080 31663 2144
rect 31727 2080 31728 2144
rect 31662 2064 31728 2080
rect 31662 2000 31663 2064
rect 31727 2000 31728 2064
rect 31662 1984 31728 2000
rect 31662 1920 31663 1984
rect 31727 1920 31728 1984
rect 31662 1904 31728 1920
rect 31662 1840 31663 1904
rect 31727 1840 31728 1904
rect 31662 1824 31728 1840
rect 31662 1760 31663 1824
rect 31727 1760 31728 1824
rect 31662 1744 31728 1760
rect 31662 1680 31663 1744
rect 31727 1680 31728 1744
rect 31662 1664 31728 1680
rect 31662 1600 31663 1664
rect 31727 1600 31728 1664
rect 31662 1446 31728 1600
rect 31788 1508 31848 2538
rect 31908 1446 31968 2478
rect 32028 1508 32088 2538
rect 32148 1446 32208 2478
rect 32268 2384 32334 2474
rect 32268 2320 32269 2384
rect 32333 2320 32334 2384
rect 32268 2304 32334 2320
rect 32268 2240 32269 2304
rect 32333 2240 32334 2304
rect 32268 2224 32334 2240
rect 32268 2160 32269 2224
rect 32333 2160 32334 2224
rect 32268 2144 32334 2160
rect 32268 2080 32269 2144
rect 32333 2080 32334 2144
rect 32268 2064 32334 2080
rect 32268 2000 32269 2064
rect 32333 2000 32334 2064
rect 32268 1984 32334 2000
rect 32268 1920 32269 1984
rect 32333 1920 32334 1984
rect 32268 1904 32334 1920
rect 32268 1840 32269 1904
rect 32333 1840 32334 1904
rect 32268 1824 32334 1840
rect 32268 1760 32269 1824
rect 32333 1760 32334 1824
rect 32268 1744 32334 1760
rect 32268 1680 32269 1744
rect 32333 1680 32334 1744
rect 32268 1664 32334 1680
rect 32268 1600 32269 1664
rect 32333 1600 32334 1664
rect 32268 1446 32334 1600
rect 32394 1508 32454 2538
rect 32514 1446 32574 2478
rect 32634 1508 32694 2538
rect 32754 1446 32814 2478
rect 32874 2384 32940 2474
rect 32874 2320 32875 2384
rect 32939 2320 32940 2384
rect 32874 2304 32940 2320
rect 32874 2240 32875 2304
rect 32939 2240 32940 2304
rect 32874 2224 32940 2240
rect 32874 2160 32875 2224
rect 32939 2160 32940 2224
rect 32874 2144 32940 2160
rect 32874 2080 32875 2144
rect 32939 2080 32940 2144
rect 32874 2064 32940 2080
rect 32874 2000 32875 2064
rect 32939 2000 32940 2064
rect 32874 1984 32940 2000
rect 32874 1920 32875 1984
rect 32939 1920 32940 1984
rect 32874 1904 32940 1920
rect 32874 1840 32875 1904
rect 32939 1840 32940 1904
rect 32874 1824 32940 1840
rect 32874 1760 32875 1824
rect 32939 1760 32940 1824
rect 32874 1744 32940 1760
rect 32874 1680 32875 1744
rect 32939 1680 32940 1744
rect 32874 1664 32940 1680
rect 32874 1600 32875 1664
rect 32939 1600 32940 1664
rect 32874 1446 32940 1600
rect 33000 1508 33060 2538
rect 33120 1446 33180 2478
rect 33240 1508 33300 2538
rect 33360 1446 33420 2478
rect 33480 2384 33546 2474
rect 33480 2320 33481 2384
rect 33545 2320 33546 2384
rect 33480 2304 33546 2320
rect 33480 2240 33481 2304
rect 33545 2240 33546 2304
rect 33480 2224 33546 2240
rect 33480 2160 33481 2224
rect 33545 2160 33546 2224
rect 33480 2144 33546 2160
rect 33480 2080 33481 2144
rect 33545 2080 33546 2144
rect 33480 2064 33546 2080
rect 33480 2000 33481 2064
rect 33545 2000 33546 2064
rect 33480 1984 33546 2000
rect 33480 1920 33481 1984
rect 33545 1920 33546 1984
rect 33480 1904 33546 1920
rect 33480 1840 33481 1904
rect 33545 1840 33546 1904
rect 33480 1824 33546 1840
rect 33480 1760 33481 1824
rect 33545 1760 33546 1824
rect 33480 1744 33546 1760
rect 33480 1680 33481 1744
rect 33545 1680 33546 1744
rect 33480 1664 33546 1680
rect 33480 1600 33481 1664
rect 33545 1600 33546 1664
rect 33480 1446 33546 1600
rect 33606 1508 33666 2538
rect 33726 1446 33786 2478
rect 33846 1508 33906 2538
rect 33966 1446 34026 2478
rect 34086 2384 34152 2474
rect 34086 2320 34087 2384
rect 34151 2320 34152 2384
rect 34086 2304 34152 2320
rect 34086 2240 34087 2304
rect 34151 2240 34152 2304
rect 34086 2224 34152 2240
rect 34086 2160 34087 2224
rect 34151 2160 34152 2224
rect 34086 2144 34152 2160
rect 34086 2080 34087 2144
rect 34151 2080 34152 2144
rect 34086 2064 34152 2080
rect 34086 2000 34087 2064
rect 34151 2000 34152 2064
rect 34086 1984 34152 2000
rect 34086 1920 34087 1984
rect 34151 1920 34152 1984
rect 34086 1904 34152 1920
rect 34086 1840 34087 1904
rect 34151 1840 34152 1904
rect 34086 1824 34152 1840
rect 34086 1760 34087 1824
rect 34151 1760 34152 1824
rect 34086 1744 34152 1760
rect 34086 1680 34087 1744
rect 34151 1680 34152 1744
rect 34086 1664 34152 1680
rect 34086 1600 34087 1664
rect 34151 1600 34152 1664
rect 34086 1446 34152 1600
rect 34212 1508 34272 2538
rect 34332 1446 34392 2478
rect 34452 1508 34512 2538
rect 34572 1446 34632 2478
rect 34692 2384 34758 2474
rect 34692 2320 34693 2384
rect 34757 2320 34758 2384
rect 34692 2304 34758 2320
rect 34692 2240 34693 2304
rect 34757 2240 34758 2304
rect 34692 2224 34758 2240
rect 34692 2160 34693 2224
rect 34757 2160 34758 2224
rect 34692 2144 34758 2160
rect 34692 2080 34693 2144
rect 34757 2080 34758 2144
rect 34692 2064 34758 2080
rect 34692 2000 34693 2064
rect 34757 2000 34758 2064
rect 34692 1984 34758 2000
rect 34692 1920 34693 1984
rect 34757 1920 34758 1984
rect 34692 1904 34758 1920
rect 34692 1840 34693 1904
rect 34757 1840 34758 1904
rect 34692 1824 34758 1840
rect 34692 1760 34693 1824
rect 34757 1760 34758 1824
rect 34692 1744 34758 1760
rect 34692 1680 34693 1744
rect 34757 1680 34758 1744
rect 34692 1664 34758 1680
rect 34692 1600 34693 1664
rect 34757 1600 34758 1664
rect 34692 1446 34758 1600
rect 34818 1508 34878 2538
rect 34938 1446 34998 2478
rect 35058 1508 35118 2538
rect 35178 1446 35238 2478
rect 35298 2384 35364 2474
rect 35298 2320 35299 2384
rect 35363 2320 35364 2384
rect 35298 2304 35364 2320
rect 35298 2240 35299 2304
rect 35363 2240 35364 2304
rect 35298 2224 35364 2240
rect 35298 2160 35299 2224
rect 35363 2160 35364 2224
rect 35298 2144 35364 2160
rect 35298 2080 35299 2144
rect 35363 2080 35364 2144
rect 35298 2064 35364 2080
rect 35298 2000 35299 2064
rect 35363 2000 35364 2064
rect 35298 1984 35364 2000
rect 35298 1920 35299 1984
rect 35363 1920 35364 1984
rect 35298 1904 35364 1920
rect 35298 1840 35299 1904
rect 35363 1840 35364 1904
rect 35298 1824 35364 1840
rect 35298 1760 35299 1824
rect 35363 1760 35364 1824
rect 35298 1744 35364 1760
rect 35298 1680 35299 1744
rect 35363 1680 35364 1744
rect 35298 1664 35364 1680
rect 35298 1600 35299 1664
rect 35363 1600 35364 1664
rect 35298 1446 35364 1600
rect 35424 1508 35484 2538
rect 35544 1446 35604 2478
rect 35664 1508 35724 2538
rect 35784 1446 35844 2478
rect 35904 2384 35970 2474
rect 35904 2320 35905 2384
rect 35969 2320 35970 2384
rect 35904 2304 35970 2320
rect 35904 2240 35905 2304
rect 35969 2240 35970 2304
rect 35904 2224 35970 2240
rect 35904 2160 35905 2224
rect 35969 2160 35970 2224
rect 35904 2144 35970 2160
rect 35904 2080 35905 2144
rect 35969 2080 35970 2144
rect 35904 2064 35970 2080
rect 35904 2000 35905 2064
rect 35969 2000 35970 2064
rect 35904 1984 35970 2000
rect 35904 1920 35905 1984
rect 35969 1920 35970 1984
rect 35904 1904 35970 1920
rect 35904 1840 35905 1904
rect 35969 1840 35970 1904
rect 35904 1824 35970 1840
rect 35904 1760 35905 1824
rect 35969 1760 35970 1824
rect 35904 1744 35970 1760
rect 35904 1680 35905 1744
rect 35969 1680 35970 1744
rect 35904 1664 35970 1680
rect 35904 1600 35905 1664
rect 35969 1600 35970 1664
rect 35904 1446 35970 1600
rect 36030 1508 36090 2538
rect 36150 1446 36210 2478
rect 36270 1508 36330 2538
rect 36390 1446 36450 2478
rect 36510 2384 36576 2474
rect 36510 2320 36511 2384
rect 36575 2320 36576 2384
rect 36510 2304 36576 2320
rect 36510 2240 36511 2304
rect 36575 2240 36576 2304
rect 36510 2224 36576 2240
rect 36510 2160 36511 2224
rect 36575 2160 36576 2224
rect 36510 2144 36576 2160
rect 36510 2080 36511 2144
rect 36575 2080 36576 2144
rect 36510 2064 36576 2080
rect 36510 2000 36511 2064
rect 36575 2000 36576 2064
rect 36510 1984 36576 2000
rect 36510 1920 36511 1984
rect 36575 1920 36576 1984
rect 36510 1904 36576 1920
rect 36510 1840 36511 1904
rect 36575 1840 36576 1904
rect 36510 1824 36576 1840
rect 36510 1760 36511 1824
rect 36575 1760 36576 1824
rect 36510 1744 36576 1760
rect 36510 1680 36511 1744
rect 36575 1680 36576 1744
rect 36510 1664 36576 1680
rect 36510 1600 36511 1664
rect 36575 1600 36576 1664
rect 36510 1446 36576 1600
rect 36636 1508 36696 2538
rect 36756 1446 36816 2478
rect 36876 1508 36936 2538
rect 36996 1446 37056 2478
rect 37116 2384 37182 2474
rect 37116 2320 37117 2384
rect 37181 2320 37182 2384
rect 37116 2304 37182 2320
rect 37116 2240 37117 2304
rect 37181 2240 37182 2304
rect 37116 2224 37182 2240
rect 37116 2160 37117 2224
rect 37181 2160 37182 2224
rect 37116 2144 37182 2160
rect 37116 2080 37117 2144
rect 37181 2080 37182 2144
rect 37116 2064 37182 2080
rect 37116 2000 37117 2064
rect 37181 2000 37182 2064
rect 37116 1984 37182 2000
rect 37116 1920 37117 1984
rect 37181 1920 37182 1984
rect 37116 1904 37182 1920
rect 37116 1840 37117 1904
rect 37181 1840 37182 1904
rect 37116 1824 37182 1840
rect 37116 1760 37117 1824
rect 37181 1760 37182 1824
rect 37116 1744 37182 1760
rect 37116 1680 37117 1744
rect 37181 1680 37182 1744
rect 37116 1664 37182 1680
rect 37116 1600 37117 1664
rect 37181 1600 37182 1664
rect 37116 1446 37182 1600
rect 37242 1508 37302 2538
rect 37362 1446 37422 2478
rect 37482 1508 37542 2538
rect 37602 1446 37662 2478
rect 37722 2384 37788 2474
rect 37722 2320 37723 2384
rect 37787 2320 37788 2384
rect 37722 2304 37788 2320
rect 37722 2240 37723 2304
rect 37787 2240 37788 2304
rect 37722 2224 37788 2240
rect 37722 2160 37723 2224
rect 37787 2160 37788 2224
rect 37722 2144 37788 2160
rect 37722 2080 37723 2144
rect 37787 2080 37788 2144
rect 37722 2064 37788 2080
rect 37722 2000 37723 2064
rect 37787 2000 37788 2064
rect 37722 1984 37788 2000
rect 37722 1920 37723 1984
rect 37787 1920 37788 1984
rect 37722 1904 37788 1920
rect 37722 1840 37723 1904
rect 37787 1840 37788 1904
rect 37722 1824 37788 1840
rect 37722 1760 37723 1824
rect 37787 1760 37788 1824
rect 37722 1744 37788 1760
rect 37722 1680 37723 1744
rect 37787 1680 37788 1744
rect 37722 1664 37788 1680
rect 37722 1600 37723 1664
rect 37787 1600 37788 1664
rect 37722 1446 37788 1600
rect 37848 1508 37908 2538
rect 37968 1446 38028 2478
rect 38088 1508 38148 2538
rect 38208 1446 38268 2478
rect 38328 2384 38394 2474
rect 38328 2320 38329 2384
rect 38393 2320 38394 2384
rect 38328 2304 38394 2320
rect 38328 2240 38329 2304
rect 38393 2240 38394 2304
rect 38328 2224 38394 2240
rect 38328 2160 38329 2224
rect 38393 2160 38394 2224
rect 38328 2144 38394 2160
rect 38328 2080 38329 2144
rect 38393 2080 38394 2144
rect 38328 2064 38394 2080
rect 38328 2000 38329 2064
rect 38393 2000 38394 2064
rect 38328 1984 38394 2000
rect 38328 1920 38329 1984
rect 38393 1920 38394 1984
rect 38328 1904 38394 1920
rect 38328 1840 38329 1904
rect 38393 1840 38394 1904
rect 38328 1824 38394 1840
rect 38328 1760 38329 1824
rect 38393 1760 38394 1824
rect 38328 1744 38394 1760
rect 38328 1680 38329 1744
rect 38393 1680 38394 1744
rect 38328 1664 38394 1680
rect 38328 1600 38329 1664
rect 38393 1600 38394 1664
rect 38328 1446 38394 1600
rect 38454 1508 38514 2538
rect 38574 1446 38634 2478
rect 38694 1508 38754 2538
rect 38814 1446 38874 2478
rect 38934 2384 39000 2474
rect 38934 2320 38935 2384
rect 38999 2320 39000 2384
rect 38934 2304 39000 2320
rect 38934 2240 38935 2304
rect 38999 2240 39000 2304
rect 38934 2224 39000 2240
rect 38934 2160 38935 2224
rect 38999 2160 39000 2224
rect 38934 2144 39000 2160
rect 38934 2080 38935 2144
rect 38999 2080 39000 2144
rect 38934 2064 39000 2080
rect 38934 2000 38935 2064
rect 38999 2000 39000 2064
rect 38934 1984 39000 2000
rect 38934 1920 38935 1984
rect 38999 1920 39000 1984
rect 38934 1904 39000 1920
rect 38934 1840 38935 1904
rect 38999 1840 39000 1904
rect 38934 1824 39000 1840
rect 38934 1760 38935 1824
rect 38999 1760 39000 1824
rect 38934 1744 39000 1760
rect 38934 1680 38935 1744
rect 38999 1680 39000 1744
rect 38934 1664 39000 1680
rect 38934 1600 38935 1664
rect 38999 1600 39000 1664
rect 38934 1446 39000 1600
rect 39060 1508 39120 2538
rect 39180 1446 39240 2478
rect 39300 1508 39360 2538
rect 39420 1446 39480 2478
rect 39540 2384 39606 2474
rect 39540 2320 39541 2384
rect 39605 2320 39606 2384
rect 39540 2304 39606 2320
rect 39540 2240 39541 2304
rect 39605 2240 39606 2304
rect 39540 2224 39606 2240
rect 39540 2160 39541 2224
rect 39605 2160 39606 2224
rect 39540 2144 39606 2160
rect 39540 2080 39541 2144
rect 39605 2080 39606 2144
rect 39540 2064 39606 2080
rect 39540 2000 39541 2064
rect 39605 2000 39606 2064
rect 39540 1984 39606 2000
rect 39540 1920 39541 1984
rect 39605 1920 39606 1984
rect 39540 1904 39606 1920
rect 39540 1840 39541 1904
rect 39605 1840 39606 1904
rect 39540 1824 39606 1840
rect 39540 1760 39541 1824
rect 39605 1760 39606 1824
rect 39540 1744 39606 1760
rect 39540 1680 39541 1744
rect 39605 1680 39606 1744
rect 39540 1664 39606 1680
rect 39540 1600 39541 1664
rect 39605 1600 39606 1664
rect 39540 1446 39606 1600
rect 20148 1444 39606 1446
rect 20148 1380 20252 1444
rect 20316 1380 20332 1444
rect 20396 1380 20412 1444
rect 20476 1380 20492 1444
rect 20556 1380 20572 1444
rect 20636 1380 20652 1444
rect 20716 1380 20858 1444
rect 20922 1380 20938 1444
rect 21002 1380 21018 1444
rect 21082 1380 21098 1444
rect 21162 1380 21178 1444
rect 21242 1380 21258 1444
rect 21322 1380 21464 1444
rect 21528 1380 21544 1444
rect 21608 1380 21624 1444
rect 21688 1380 21704 1444
rect 21768 1380 21784 1444
rect 21848 1380 21864 1444
rect 21928 1380 22070 1444
rect 22134 1380 22150 1444
rect 22214 1380 22230 1444
rect 22294 1380 22310 1444
rect 22374 1380 22390 1444
rect 22454 1380 22470 1444
rect 22534 1380 22676 1444
rect 22740 1380 22756 1444
rect 22820 1380 22836 1444
rect 22900 1380 22916 1444
rect 22980 1380 22996 1444
rect 23060 1380 23076 1444
rect 23140 1380 23282 1444
rect 23346 1380 23362 1444
rect 23426 1380 23442 1444
rect 23506 1380 23522 1444
rect 23586 1380 23602 1444
rect 23666 1380 23682 1444
rect 23746 1380 23888 1444
rect 23952 1380 23968 1444
rect 24032 1380 24048 1444
rect 24112 1380 24128 1444
rect 24192 1380 24208 1444
rect 24272 1380 24288 1444
rect 24352 1380 24494 1444
rect 24558 1380 24574 1444
rect 24638 1380 24654 1444
rect 24718 1380 24734 1444
rect 24798 1380 24814 1444
rect 24878 1380 24894 1444
rect 24958 1380 25100 1444
rect 25164 1380 25180 1444
rect 25244 1380 25260 1444
rect 25324 1380 25340 1444
rect 25404 1380 25420 1444
rect 25484 1380 25500 1444
rect 25564 1380 25706 1444
rect 25770 1380 25786 1444
rect 25850 1380 25866 1444
rect 25930 1380 25946 1444
rect 26010 1380 26026 1444
rect 26090 1380 26106 1444
rect 26170 1380 26312 1444
rect 26376 1380 26392 1444
rect 26456 1380 26472 1444
rect 26536 1380 26552 1444
rect 26616 1380 26632 1444
rect 26696 1380 26712 1444
rect 26776 1380 26918 1444
rect 26982 1380 26998 1444
rect 27062 1380 27078 1444
rect 27142 1380 27158 1444
rect 27222 1380 27238 1444
rect 27302 1380 27318 1444
rect 27382 1380 27524 1444
rect 27588 1380 27604 1444
rect 27668 1380 27684 1444
rect 27748 1380 27764 1444
rect 27828 1380 27844 1444
rect 27908 1380 27924 1444
rect 27988 1380 28130 1444
rect 28194 1380 28210 1444
rect 28274 1380 28290 1444
rect 28354 1380 28370 1444
rect 28434 1380 28450 1444
rect 28514 1380 28530 1444
rect 28594 1380 28736 1444
rect 28800 1380 28816 1444
rect 28880 1380 28896 1444
rect 28960 1380 28976 1444
rect 29040 1380 29056 1444
rect 29120 1380 29136 1444
rect 29200 1380 29342 1444
rect 29406 1380 29422 1444
rect 29486 1380 29502 1444
rect 29566 1380 29582 1444
rect 29646 1380 29662 1444
rect 29726 1380 29742 1444
rect 29806 1380 29948 1444
rect 30012 1380 30028 1444
rect 30092 1380 30108 1444
rect 30172 1380 30188 1444
rect 30252 1380 30268 1444
rect 30332 1380 30348 1444
rect 30412 1380 30554 1444
rect 30618 1380 30634 1444
rect 30698 1380 30714 1444
rect 30778 1380 30794 1444
rect 30858 1380 30874 1444
rect 30938 1380 30954 1444
rect 31018 1380 31160 1444
rect 31224 1380 31240 1444
rect 31304 1380 31320 1444
rect 31384 1380 31400 1444
rect 31464 1380 31480 1444
rect 31544 1380 31560 1444
rect 31624 1380 31766 1444
rect 31830 1380 31846 1444
rect 31910 1380 31926 1444
rect 31990 1380 32006 1444
rect 32070 1380 32086 1444
rect 32150 1380 32166 1444
rect 32230 1380 32372 1444
rect 32436 1380 32452 1444
rect 32516 1380 32532 1444
rect 32596 1380 32612 1444
rect 32676 1380 32692 1444
rect 32756 1380 32772 1444
rect 32836 1380 32978 1444
rect 33042 1380 33058 1444
rect 33122 1380 33138 1444
rect 33202 1380 33218 1444
rect 33282 1380 33298 1444
rect 33362 1380 33378 1444
rect 33442 1380 33584 1444
rect 33648 1380 33664 1444
rect 33728 1380 33744 1444
rect 33808 1380 33824 1444
rect 33888 1380 33904 1444
rect 33968 1380 33984 1444
rect 34048 1380 34190 1444
rect 34254 1380 34270 1444
rect 34334 1380 34350 1444
rect 34414 1380 34430 1444
rect 34494 1380 34510 1444
rect 34574 1380 34590 1444
rect 34654 1380 34796 1444
rect 34860 1380 34876 1444
rect 34940 1380 34956 1444
rect 35020 1380 35036 1444
rect 35100 1380 35116 1444
rect 35180 1380 35196 1444
rect 35260 1380 35402 1444
rect 35466 1380 35482 1444
rect 35546 1380 35562 1444
rect 35626 1380 35642 1444
rect 35706 1380 35722 1444
rect 35786 1380 35802 1444
rect 35866 1380 36008 1444
rect 36072 1380 36088 1444
rect 36152 1380 36168 1444
rect 36232 1380 36248 1444
rect 36312 1380 36328 1444
rect 36392 1380 36408 1444
rect 36472 1380 36614 1444
rect 36678 1380 36694 1444
rect 36758 1380 36774 1444
rect 36838 1380 36854 1444
rect 36918 1380 36934 1444
rect 36998 1380 37014 1444
rect 37078 1380 37220 1444
rect 37284 1380 37300 1444
rect 37364 1380 37380 1444
rect 37444 1380 37460 1444
rect 37524 1380 37540 1444
rect 37604 1380 37620 1444
rect 37684 1380 37826 1444
rect 37890 1380 37906 1444
rect 37970 1380 37986 1444
rect 38050 1380 38066 1444
rect 38130 1380 38146 1444
rect 38210 1380 38226 1444
rect 38290 1380 38432 1444
rect 38496 1380 38512 1444
rect 38576 1380 38592 1444
rect 38656 1380 38672 1444
rect 38736 1380 38752 1444
rect 38816 1380 38832 1444
rect 38896 1380 39038 1444
rect 39102 1380 39118 1444
rect 39182 1380 39198 1444
rect 39262 1380 39278 1444
rect 39342 1380 39358 1444
rect 39422 1380 39438 1444
rect 39502 1380 39606 1444
rect 20148 1378 39606 1380
rect 20148 1224 20214 1378
rect 20148 1160 20149 1224
rect 20213 1160 20214 1224
rect 20148 1144 20214 1160
rect 20148 1080 20149 1144
rect 20213 1080 20214 1144
rect 20148 1064 20214 1080
rect 20148 1000 20149 1064
rect 20213 1000 20214 1064
rect 20148 984 20214 1000
rect 20148 920 20149 984
rect 20213 920 20214 984
rect 20148 904 20214 920
rect 20148 840 20149 904
rect 20213 840 20214 904
rect 20148 824 20214 840
rect 20148 760 20149 824
rect 20213 760 20214 824
rect 20148 744 20214 760
rect 20148 680 20149 744
rect 20213 680 20214 744
rect 20148 664 20214 680
rect 20148 600 20149 664
rect 20213 600 20214 664
rect 20148 584 20214 600
rect 20148 520 20149 584
rect 20213 520 20214 584
rect 20148 504 20214 520
rect 20148 440 20149 504
rect 20213 440 20214 504
rect 20148 350 20214 440
rect 20274 346 20334 1378
rect 20394 286 20454 1316
rect 20514 346 20574 1378
rect 20634 286 20694 1316
rect 20754 1224 20820 1378
rect 20754 1160 20755 1224
rect 20819 1160 20820 1224
rect 20754 1144 20820 1160
rect 20754 1080 20755 1144
rect 20819 1080 20820 1144
rect 20754 1064 20820 1080
rect 20754 1000 20755 1064
rect 20819 1000 20820 1064
rect 20754 984 20820 1000
rect 20754 920 20755 984
rect 20819 920 20820 984
rect 20754 904 20820 920
rect 20754 840 20755 904
rect 20819 840 20820 904
rect 20754 824 20820 840
rect 20754 760 20755 824
rect 20819 760 20820 824
rect 20754 744 20820 760
rect 20754 680 20755 744
rect 20819 680 20820 744
rect 20754 664 20820 680
rect 20754 600 20755 664
rect 20819 600 20820 664
rect 20754 584 20820 600
rect 20754 520 20755 584
rect 20819 520 20820 584
rect 20754 504 20820 520
rect 20754 440 20755 504
rect 20819 440 20820 504
rect 20754 350 20820 440
rect 20880 346 20940 1378
rect 21000 286 21060 1316
rect 21120 346 21180 1378
rect 21240 286 21300 1316
rect 21360 1224 21426 1378
rect 21360 1160 21361 1224
rect 21425 1160 21426 1224
rect 21360 1144 21426 1160
rect 21360 1080 21361 1144
rect 21425 1080 21426 1144
rect 21360 1064 21426 1080
rect 21360 1000 21361 1064
rect 21425 1000 21426 1064
rect 21360 984 21426 1000
rect 21360 920 21361 984
rect 21425 920 21426 984
rect 21360 904 21426 920
rect 21360 840 21361 904
rect 21425 840 21426 904
rect 21360 824 21426 840
rect 21360 760 21361 824
rect 21425 760 21426 824
rect 21360 744 21426 760
rect 21360 680 21361 744
rect 21425 680 21426 744
rect 21360 664 21426 680
rect 21360 600 21361 664
rect 21425 600 21426 664
rect 21360 584 21426 600
rect 21360 520 21361 584
rect 21425 520 21426 584
rect 21360 504 21426 520
rect 21360 440 21361 504
rect 21425 440 21426 504
rect 21360 350 21426 440
rect 21486 346 21546 1378
rect 21606 286 21666 1316
rect 21726 346 21786 1378
rect 21846 286 21906 1316
rect 21966 1224 22032 1378
rect 21966 1160 21967 1224
rect 22031 1160 22032 1224
rect 21966 1144 22032 1160
rect 21966 1080 21967 1144
rect 22031 1080 22032 1144
rect 21966 1064 22032 1080
rect 21966 1000 21967 1064
rect 22031 1000 22032 1064
rect 21966 984 22032 1000
rect 21966 920 21967 984
rect 22031 920 22032 984
rect 21966 904 22032 920
rect 21966 840 21967 904
rect 22031 840 22032 904
rect 21966 824 22032 840
rect 21966 760 21967 824
rect 22031 760 22032 824
rect 21966 744 22032 760
rect 21966 680 21967 744
rect 22031 680 22032 744
rect 21966 664 22032 680
rect 21966 600 21967 664
rect 22031 600 22032 664
rect 21966 584 22032 600
rect 21966 520 21967 584
rect 22031 520 22032 584
rect 21966 504 22032 520
rect 21966 440 21967 504
rect 22031 440 22032 504
rect 21966 350 22032 440
rect 22092 346 22152 1378
rect 22212 286 22272 1316
rect 22332 346 22392 1378
rect 22452 286 22512 1316
rect 22572 1224 22638 1378
rect 22572 1160 22573 1224
rect 22637 1160 22638 1224
rect 22572 1144 22638 1160
rect 22572 1080 22573 1144
rect 22637 1080 22638 1144
rect 22572 1064 22638 1080
rect 22572 1000 22573 1064
rect 22637 1000 22638 1064
rect 22572 984 22638 1000
rect 22572 920 22573 984
rect 22637 920 22638 984
rect 22572 904 22638 920
rect 22572 840 22573 904
rect 22637 840 22638 904
rect 22572 824 22638 840
rect 22572 760 22573 824
rect 22637 760 22638 824
rect 22572 744 22638 760
rect 22572 680 22573 744
rect 22637 680 22638 744
rect 22572 664 22638 680
rect 22572 600 22573 664
rect 22637 600 22638 664
rect 22572 584 22638 600
rect 22572 520 22573 584
rect 22637 520 22638 584
rect 22572 504 22638 520
rect 22572 440 22573 504
rect 22637 440 22638 504
rect 22572 350 22638 440
rect 22698 346 22758 1378
rect 22818 286 22878 1316
rect 22938 346 22998 1378
rect 23058 286 23118 1316
rect 23178 1224 23244 1378
rect 23178 1160 23179 1224
rect 23243 1160 23244 1224
rect 23178 1144 23244 1160
rect 23178 1080 23179 1144
rect 23243 1080 23244 1144
rect 23178 1064 23244 1080
rect 23178 1000 23179 1064
rect 23243 1000 23244 1064
rect 23178 984 23244 1000
rect 23178 920 23179 984
rect 23243 920 23244 984
rect 23178 904 23244 920
rect 23178 840 23179 904
rect 23243 840 23244 904
rect 23178 824 23244 840
rect 23178 760 23179 824
rect 23243 760 23244 824
rect 23178 744 23244 760
rect 23178 680 23179 744
rect 23243 680 23244 744
rect 23178 664 23244 680
rect 23178 600 23179 664
rect 23243 600 23244 664
rect 23178 584 23244 600
rect 23178 520 23179 584
rect 23243 520 23244 584
rect 23178 504 23244 520
rect 23178 440 23179 504
rect 23243 440 23244 504
rect 23178 350 23244 440
rect 23304 346 23364 1378
rect 23424 286 23484 1316
rect 23544 346 23604 1378
rect 23664 286 23724 1316
rect 23784 1224 23850 1378
rect 23784 1160 23785 1224
rect 23849 1160 23850 1224
rect 23784 1144 23850 1160
rect 23784 1080 23785 1144
rect 23849 1080 23850 1144
rect 23784 1064 23850 1080
rect 23784 1000 23785 1064
rect 23849 1000 23850 1064
rect 23784 984 23850 1000
rect 23784 920 23785 984
rect 23849 920 23850 984
rect 23784 904 23850 920
rect 23784 840 23785 904
rect 23849 840 23850 904
rect 23784 824 23850 840
rect 23784 760 23785 824
rect 23849 760 23850 824
rect 23784 744 23850 760
rect 23784 680 23785 744
rect 23849 680 23850 744
rect 23784 664 23850 680
rect 23784 600 23785 664
rect 23849 600 23850 664
rect 23784 584 23850 600
rect 23784 520 23785 584
rect 23849 520 23850 584
rect 23784 504 23850 520
rect 23784 440 23785 504
rect 23849 440 23850 504
rect 23784 350 23850 440
rect 23910 346 23970 1378
rect 24030 286 24090 1316
rect 24150 346 24210 1378
rect 24270 286 24330 1316
rect 24390 1224 24456 1378
rect 24390 1160 24391 1224
rect 24455 1160 24456 1224
rect 24390 1144 24456 1160
rect 24390 1080 24391 1144
rect 24455 1080 24456 1144
rect 24390 1064 24456 1080
rect 24390 1000 24391 1064
rect 24455 1000 24456 1064
rect 24390 984 24456 1000
rect 24390 920 24391 984
rect 24455 920 24456 984
rect 24390 904 24456 920
rect 24390 840 24391 904
rect 24455 840 24456 904
rect 24390 824 24456 840
rect 24390 760 24391 824
rect 24455 760 24456 824
rect 24390 744 24456 760
rect 24390 680 24391 744
rect 24455 680 24456 744
rect 24390 664 24456 680
rect 24390 600 24391 664
rect 24455 600 24456 664
rect 24390 584 24456 600
rect 24390 520 24391 584
rect 24455 520 24456 584
rect 24390 504 24456 520
rect 24390 440 24391 504
rect 24455 440 24456 504
rect 24390 350 24456 440
rect 24516 346 24576 1378
rect 24636 286 24696 1316
rect 24756 346 24816 1378
rect 24876 286 24936 1316
rect 24996 1224 25062 1378
rect 24996 1160 24997 1224
rect 25061 1160 25062 1224
rect 24996 1144 25062 1160
rect 24996 1080 24997 1144
rect 25061 1080 25062 1144
rect 24996 1064 25062 1080
rect 24996 1000 24997 1064
rect 25061 1000 25062 1064
rect 24996 984 25062 1000
rect 24996 920 24997 984
rect 25061 920 25062 984
rect 24996 904 25062 920
rect 24996 840 24997 904
rect 25061 840 25062 904
rect 24996 824 25062 840
rect 24996 760 24997 824
rect 25061 760 25062 824
rect 24996 744 25062 760
rect 24996 680 24997 744
rect 25061 680 25062 744
rect 24996 664 25062 680
rect 24996 600 24997 664
rect 25061 600 25062 664
rect 24996 584 25062 600
rect 24996 520 24997 584
rect 25061 520 25062 584
rect 24996 504 25062 520
rect 24996 440 24997 504
rect 25061 440 25062 504
rect 24996 350 25062 440
rect 25122 346 25182 1378
rect 25242 286 25302 1316
rect 25362 346 25422 1378
rect 25482 286 25542 1316
rect 25602 1224 25668 1378
rect 25602 1160 25603 1224
rect 25667 1160 25668 1224
rect 25602 1144 25668 1160
rect 25602 1080 25603 1144
rect 25667 1080 25668 1144
rect 25602 1064 25668 1080
rect 25602 1000 25603 1064
rect 25667 1000 25668 1064
rect 25602 984 25668 1000
rect 25602 920 25603 984
rect 25667 920 25668 984
rect 25602 904 25668 920
rect 25602 840 25603 904
rect 25667 840 25668 904
rect 25602 824 25668 840
rect 25602 760 25603 824
rect 25667 760 25668 824
rect 25602 744 25668 760
rect 25602 680 25603 744
rect 25667 680 25668 744
rect 25602 664 25668 680
rect 25602 600 25603 664
rect 25667 600 25668 664
rect 25602 584 25668 600
rect 25602 520 25603 584
rect 25667 520 25668 584
rect 25602 504 25668 520
rect 25602 440 25603 504
rect 25667 440 25668 504
rect 25602 350 25668 440
rect 25728 346 25788 1378
rect 25848 286 25908 1316
rect 25968 346 26028 1378
rect 26088 286 26148 1316
rect 26208 1224 26274 1378
rect 26208 1160 26209 1224
rect 26273 1160 26274 1224
rect 26208 1144 26274 1160
rect 26208 1080 26209 1144
rect 26273 1080 26274 1144
rect 26208 1064 26274 1080
rect 26208 1000 26209 1064
rect 26273 1000 26274 1064
rect 26208 984 26274 1000
rect 26208 920 26209 984
rect 26273 920 26274 984
rect 26208 904 26274 920
rect 26208 840 26209 904
rect 26273 840 26274 904
rect 26208 824 26274 840
rect 26208 760 26209 824
rect 26273 760 26274 824
rect 26208 744 26274 760
rect 26208 680 26209 744
rect 26273 680 26274 744
rect 26208 664 26274 680
rect 26208 600 26209 664
rect 26273 600 26274 664
rect 26208 584 26274 600
rect 26208 520 26209 584
rect 26273 520 26274 584
rect 26208 504 26274 520
rect 26208 440 26209 504
rect 26273 440 26274 504
rect 26208 350 26274 440
rect 26334 346 26394 1378
rect 26454 286 26514 1316
rect 26574 346 26634 1378
rect 26694 286 26754 1316
rect 26814 1224 26880 1378
rect 26814 1160 26815 1224
rect 26879 1160 26880 1224
rect 26814 1144 26880 1160
rect 26814 1080 26815 1144
rect 26879 1080 26880 1144
rect 26814 1064 26880 1080
rect 26814 1000 26815 1064
rect 26879 1000 26880 1064
rect 26814 984 26880 1000
rect 26814 920 26815 984
rect 26879 920 26880 984
rect 26814 904 26880 920
rect 26814 840 26815 904
rect 26879 840 26880 904
rect 26814 824 26880 840
rect 26814 760 26815 824
rect 26879 760 26880 824
rect 26814 744 26880 760
rect 26814 680 26815 744
rect 26879 680 26880 744
rect 26814 664 26880 680
rect 26814 600 26815 664
rect 26879 600 26880 664
rect 26814 584 26880 600
rect 26814 520 26815 584
rect 26879 520 26880 584
rect 26814 504 26880 520
rect 26814 440 26815 504
rect 26879 440 26880 504
rect 26814 350 26880 440
rect 26940 346 27000 1378
rect 27060 286 27120 1316
rect 27180 346 27240 1378
rect 27300 286 27360 1316
rect 27420 1224 27486 1378
rect 27420 1160 27421 1224
rect 27485 1160 27486 1224
rect 27420 1144 27486 1160
rect 27420 1080 27421 1144
rect 27485 1080 27486 1144
rect 27420 1064 27486 1080
rect 27420 1000 27421 1064
rect 27485 1000 27486 1064
rect 27420 984 27486 1000
rect 27420 920 27421 984
rect 27485 920 27486 984
rect 27420 904 27486 920
rect 27420 840 27421 904
rect 27485 840 27486 904
rect 27420 824 27486 840
rect 27420 760 27421 824
rect 27485 760 27486 824
rect 27420 744 27486 760
rect 27420 680 27421 744
rect 27485 680 27486 744
rect 27420 664 27486 680
rect 27420 600 27421 664
rect 27485 600 27486 664
rect 27420 584 27486 600
rect 27420 520 27421 584
rect 27485 520 27486 584
rect 27420 504 27486 520
rect 27420 440 27421 504
rect 27485 440 27486 504
rect 27420 350 27486 440
rect 27546 346 27606 1378
rect 27666 286 27726 1316
rect 27786 346 27846 1378
rect 27906 286 27966 1316
rect 28026 1224 28092 1378
rect 28026 1160 28027 1224
rect 28091 1160 28092 1224
rect 28026 1144 28092 1160
rect 28026 1080 28027 1144
rect 28091 1080 28092 1144
rect 28026 1064 28092 1080
rect 28026 1000 28027 1064
rect 28091 1000 28092 1064
rect 28026 984 28092 1000
rect 28026 920 28027 984
rect 28091 920 28092 984
rect 28026 904 28092 920
rect 28026 840 28027 904
rect 28091 840 28092 904
rect 28026 824 28092 840
rect 28026 760 28027 824
rect 28091 760 28092 824
rect 28026 744 28092 760
rect 28026 680 28027 744
rect 28091 680 28092 744
rect 28026 664 28092 680
rect 28026 600 28027 664
rect 28091 600 28092 664
rect 28026 584 28092 600
rect 28026 520 28027 584
rect 28091 520 28092 584
rect 28026 504 28092 520
rect 28026 440 28027 504
rect 28091 440 28092 504
rect 28026 350 28092 440
rect 28152 346 28212 1378
rect 28272 286 28332 1316
rect 28392 346 28452 1378
rect 28512 286 28572 1316
rect 28632 1224 28698 1378
rect 28632 1160 28633 1224
rect 28697 1160 28698 1224
rect 28632 1144 28698 1160
rect 28632 1080 28633 1144
rect 28697 1080 28698 1144
rect 28632 1064 28698 1080
rect 28632 1000 28633 1064
rect 28697 1000 28698 1064
rect 28632 984 28698 1000
rect 28632 920 28633 984
rect 28697 920 28698 984
rect 28632 904 28698 920
rect 28632 840 28633 904
rect 28697 840 28698 904
rect 28632 824 28698 840
rect 28632 760 28633 824
rect 28697 760 28698 824
rect 28632 744 28698 760
rect 28632 680 28633 744
rect 28697 680 28698 744
rect 28632 664 28698 680
rect 28632 600 28633 664
rect 28697 600 28698 664
rect 28632 584 28698 600
rect 28632 520 28633 584
rect 28697 520 28698 584
rect 28632 504 28698 520
rect 28632 440 28633 504
rect 28697 440 28698 504
rect 28632 350 28698 440
rect 28758 346 28818 1378
rect 28878 286 28938 1316
rect 28998 346 29058 1378
rect 29118 286 29178 1316
rect 29238 1224 29304 1378
rect 29238 1160 29239 1224
rect 29303 1160 29304 1224
rect 29238 1144 29304 1160
rect 29238 1080 29239 1144
rect 29303 1080 29304 1144
rect 29238 1064 29304 1080
rect 29238 1000 29239 1064
rect 29303 1000 29304 1064
rect 29238 984 29304 1000
rect 29238 920 29239 984
rect 29303 920 29304 984
rect 29238 904 29304 920
rect 29238 840 29239 904
rect 29303 840 29304 904
rect 29238 824 29304 840
rect 29238 760 29239 824
rect 29303 760 29304 824
rect 29238 744 29304 760
rect 29238 680 29239 744
rect 29303 680 29304 744
rect 29238 664 29304 680
rect 29238 600 29239 664
rect 29303 600 29304 664
rect 29238 584 29304 600
rect 29238 520 29239 584
rect 29303 520 29304 584
rect 29238 504 29304 520
rect 29238 440 29239 504
rect 29303 440 29304 504
rect 29238 350 29304 440
rect 29364 346 29424 1378
rect 29484 286 29544 1316
rect 29604 346 29664 1378
rect 29724 286 29784 1316
rect 29844 1224 29910 1378
rect 29844 1160 29845 1224
rect 29909 1160 29910 1224
rect 29844 1144 29910 1160
rect 29844 1080 29845 1144
rect 29909 1080 29910 1144
rect 29844 1064 29910 1080
rect 29844 1000 29845 1064
rect 29909 1000 29910 1064
rect 29844 984 29910 1000
rect 29844 920 29845 984
rect 29909 920 29910 984
rect 29844 904 29910 920
rect 29844 840 29845 904
rect 29909 840 29910 904
rect 29844 824 29910 840
rect 29844 760 29845 824
rect 29909 760 29910 824
rect 29844 744 29910 760
rect 29844 680 29845 744
rect 29909 680 29910 744
rect 29844 664 29910 680
rect 29844 600 29845 664
rect 29909 600 29910 664
rect 29844 584 29910 600
rect 29844 520 29845 584
rect 29909 520 29910 584
rect 29844 504 29910 520
rect 29844 440 29845 504
rect 29909 440 29910 504
rect 29844 350 29910 440
rect 29970 346 30030 1378
rect 30090 286 30150 1316
rect 30210 346 30270 1378
rect 30330 286 30390 1316
rect 30450 1224 30516 1378
rect 30450 1160 30451 1224
rect 30515 1160 30516 1224
rect 30450 1144 30516 1160
rect 30450 1080 30451 1144
rect 30515 1080 30516 1144
rect 30450 1064 30516 1080
rect 30450 1000 30451 1064
rect 30515 1000 30516 1064
rect 30450 984 30516 1000
rect 30450 920 30451 984
rect 30515 920 30516 984
rect 30450 904 30516 920
rect 30450 840 30451 904
rect 30515 840 30516 904
rect 30450 824 30516 840
rect 30450 760 30451 824
rect 30515 760 30516 824
rect 30450 744 30516 760
rect 30450 680 30451 744
rect 30515 680 30516 744
rect 30450 664 30516 680
rect 30450 600 30451 664
rect 30515 600 30516 664
rect 30450 584 30516 600
rect 30450 520 30451 584
rect 30515 520 30516 584
rect 30450 504 30516 520
rect 30450 440 30451 504
rect 30515 440 30516 504
rect 30450 350 30516 440
rect 30576 346 30636 1378
rect 30696 286 30756 1316
rect 30816 346 30876 1378
rect 30936 286 30996 1316
rect 31056 1224 31122 1378
rect 31056 1160 31057 1224
rect 31121 1160 31122 1224
rect 31056 1144 31122 1160
rect 31056 1080 31057 1144
rect 31121 1080 31122 1144
rect 31056 1064 31122 1080
rect 31056 1000 31057 1064
rect 31121 1000 31122 1064
rect 31056 984 31122 1000
rect 31056 920 31057 984
rect 31121 920 31122 984
rect 31056 904 31122 920
rect 31056 840 31057 904
rect 31121 840 31122 904
rect 31056 824 31122 840
rect 31056 760 31057 824
rect 31121 760 31122 824
rect 31056 744 31122 760
rect 31056 680 31057 744
rect 31121 680 31122 744
rect 31056 664 31122 680
rect 31056 600 31057 664
rect 31121 600 31122 664
rect 31056 584 31122 600
rect 31056 520 31057 584
rect 31121 520 31122 584
rect 31056 504 31122 520
rect 31056 440 31057 504
rect 31121 440 31122 504
rect 31056 350 31122 440
rect 31182 346 31242 1378
rect 31302 286 31362 1316
rect 31422 346 31482 1378
rect 31542 286 31602 1316
rect 31662 1224 31728 1378
rect 31662 1160 31663 1224
rect 31727 1160 31728 1224
rect 31662 1144 31728 1160
rect 31662 1080 31663 1144
rect 31727 1080 31728 1144
rect 31662 1064 31728 1080
rect 31662 1000 31663 1064
rect 31727 1000 31728 1064
rect 31662 984 31728 1000
rect 31662 920 31663 984
rect 31727 920 31728 984
rect 31662 904 31728 920
rect 31662 840 31663 904
rect 31727 840 31728 904
rect 31662 824 31728 840
rect 31662 760 31663 824
rect 31727 760 31728 824
rect 31662 744 31728 760
rect 31662 680 31663 744
rect 31727 680 31728 744
rect 31662 664 31728 680
rect 31662 600 31663 664
rect 31727 600 31728 664
rect 31662 584 31728 600
rect 31662 520 31663 584
rect 31727 520 31728 584
rect 31662 504 31728 520
rect 31662 440 31663 504
rect 31727 440 31728 504
rect 31662 350 31728 440
rect 31788 346 31848 1378
rect 31908 286 31968 1316
rect 32028 346 32088 1378
rect 32148 286 32208 1316
rect 32268 1224 32334 1378
rect 32268 1160 32269 1224
rect 32333 1160 32334 1224
rect 32268 1144 32334 1160
rect 32268 1080 32269 1144
rect 32333 1080 32334 1144
rect 32268 1064 32334 1080
rect 32268 1000 32269 1064
rect 32333 1000 32334 1064
rect 32268 984 32334 1000
rect 32268 920 32269 984
rect 32333 920 32334 984
rect 32268 904 32334 920
rect 32268 840 32269 904
rect 32333 840 32334 904
rect 32268 824 32334 840
rect 32268 760 32269 824
rect 32333 760 32334 824
rect 32268 744 32334 760
rect 32268 680 32269 744
rect 32333 680 32334 744
rect 32268 664 32334 680
rect 32268 600 32269 664
rect 32333 600 32334 664
rect 32268 584 32334 600
rect 32268 520 32269 584
rect 32333 520 32334 584
rect 32268 504 32334 520
rect 32268 440 32269 504
rect 32333 440 32334 504
rect 32268 350 32334 440
rect 32394 346 32454 1378
rect 32514 286 32574 1316
rect 32634 346 32694 1378
rect 32754 286 32814 1316
rect 32874 1224 32940 1378
rect 32874 1160 32875 1224
rect 32939 1160 32940 1224
rect 32874 1144 32940 1160
rect 32874 1080 32875 1144
rect 32939 1080 32940 1144
rect 32874 1064 32940 1080
rect 32874 1000 32875 1064
rect 32939 1000 32940 1064
rect 32874 984 32940 1000
rect 32874 920 32875 984
rect 32939 920 32940 984
rect 32874 904 32940 920
rect 32874 840 32875 904
rect 32939 840 32940 904
rect 32874 824 32940 840
rect 32874 760 32875 824
rect 32939 760 32940 824
rect 32874 744 32940 760
rect 32874 680 32875 744
rect 32939 680 32940 744
rect 32874 664 32940 680
rect 32874 600 32875 664
rect 32939 600 32940 664
rect 32874 584 32940 600
rect 32874 520 32875 584
rect 32939 520 32940 584
rect 32874 504 32940 520
rect 32874 440 32875 504
rect 32939 440 32940 504
rect 32874 350 32940 440
rect 33000 346 33060 1378
rect 33120 286 33180 1316
rect 33240 346 33300 1378
rect 33360 286 33420 1316
rect 33480 1224 33546 1378
rect 33480 1160 33481 1224
rect 33545 1160 33546 1224
rect 33480 1144 33546 1160
rect 33480 1080 33481 1144
rect 33545 1080 33546 1144
rect 33480 1064 33546 1080
rect 33480 1000 33481 1064
rect 33545 1000 33546 1064
rect 33480 984 33546 1000
rect 33480 920 33481 984
rect 33545 920 33546 984
rect 33480 904 33546 920
rect 33480 840 33481 904
rect 33545 840 33546 904
rect 33480 824 33546 840
rect 33480 760 33481 824
rect 33545 760 33546 824
rect 33480 744 33546 760
rect 33480 680 33481 744
rect 33545 680 33546 744
rect 33480 664 33546 680
rect 33480 600 33481 664
rect 33545 600 33546 664
rect 33480 584 33546 600
rect 33480 520 33481 584
rect 33545 520 33546 584
rect 33480 504 33546 520
rect 33480 440 33481 504
rect 33545 440 33546 504
rect 33480 350 33546 440
rect 33606 346 33666 1378
rect 33726 286 33786 1316
rect 33846 346 33906 1378
rect 33966 286 34026 1316
rect 34086 1224 34152 1378
rect 34086 1160 34087 1224
rect 34151 1160 34152 1224
rect 34086 1144 34152 1160
rect 34086 1080 34087 1144
rect 34151 1080 34152 1144
rect 34086 1064 34152 1080
rect 34086 1000 34087 1064
rect 34151 1000 34152 1064
rect 34086 984 34152 1000
rect 34086 920 34087 984
rect 34151 920 34152 984
rect 34086 904 34152 920
rect 34086 840 34087 904
rect 34151 840 34152 904
rect 34086 824 34152 840
rect 34086 760 34087 824
rect 34151 760 34152 824
rect 34086 744 34152 760
rect 34086 680 34087 744
rect 34151 680 34152 744
rect 34086 664 34152 680
rect 34086 600 34087 664
rect 34151 600 34152 664
rect 34086 584 34152 600
rect 34086 520 34087 584
rect 34151 520 34152 584
rect 34086 504 34152 520
rect 34086 440 34087 504
rect 34151 440 34152 504
rect 34086 350 34152 440
rect 34212 346 34272 1378
rect 34332 286 34392 1316
rect 34452 346 34512 1378
rect 34572 286 34632 1316
rect 34692 1224 34758 1378
rect 34692 1160 34693 1224
rect 34757 1160 34758 1224
rect 34692 1144 34758 1160
rect 34692 1080 34693 1144
rect 34757 1080 34758 1144
rect 34692 1064 34758 1080
rect 34692 1000 34693 1064
rect 34757 1000 34758 1064
rect 34692 984 34758 1000
rect 34692 920 34693 984
rect 34757 920 34758 984
rect 34692 904 34758 920
rect 34692 840 34693 904
rect 34757 840 34758 904
rect 34692 824 34758 840
rect 34692 760 34693 824
rect 34757 760 34758 824
rect 34692 744 34758 760
rect 34692 680 34693 744
rect 34757 680 34758 744
rect 34692 664 34758 680
rect 34692 600 34693 664
rect 34757 600 34758 664
rect 34692 584 34758 600
rect 34692 520 34693 584
rect 34757 520 34758 584
rect 34692 504 34758 520
rect 34692 440 34693 504
rect 34757 440 34758 504
rect 34692 350 34758 440
rect 34818 346 34878 1378
rect 34938 286 34998 1316
rect 35058 346 35118 1378
rect 35178 286 35238 1316
rect 35298 1224 35364 1378
rect 35298 1160 35299 1224
rect 35363 1160 35364 1224
rect 35298 1144 35364 1160
rect 35298 1080 35299 1144
rect 35363 1080 35364 1144
rect 35298 1064 35364 1080
rect 35298 1000 35299 1064
rect 35363 1000 35364 1064
rect 35298 984 35364 1000
rect 35298 920 35299 984
rect 35363 920 35364 984
rect 35298 904 35364 920
rect 35298 840 35299 904
rect 35363 840 35364 904
rect 35298 824 35364 840
rect 35298 760 35299 824
rect 35363 760 35364 824
rect 35298 744 35364 760
rect 35298 680 35299 744
rect 35363 680 35364 744
rect 35298 664 35364 680
rect 35298 600 35299 664
rect 35363 600 35364 664
rect 35298 584 35364 600
rect 35298 520 35299 584
rect 35363 520 35364 584
rect 35298 504 35364 520
rect 35298 440 35299 504
rect 35363 440 35364 504
rect 35298 350 35364 440
rect 35424 346 35484 1378
rect 35544 286 35604 1316
rect 35664 346 35724 1378
rect 35784 286 35844 1316
rect 35904 1224 35970 1378
rect 35904 1160 35905 1224
rect 35969 1160 35970 1224
rect 35904 1144 35970 1160
rect 35904 1080 35905 1144
rect 35969 1080 35970 1144
rect 35904 1064 35970 1080
rect 35904 1000 35905 1064
rect 35969 1000 35970 1064
rect 35904 984 35970 1000
rect 35904 920 35905 984
rect 35969 920 35970 984
rect 35904 904 35970 920
rect 35904 840 35905 904
rect 35969 840 35970 904
rect 35904 824 35970 840
rect 35904 760 35905 824
rect 35969 760 35970 824
rect 35904 744 35970 760
rect 35904 680 35905 744
rect 35969 680 35970 744
rect 35904 664 35970 680
rect 35904 600 35905 664
rect 35969 600 35970 664
rect 35904 584 35970 600
rect 35904 520 35905 584
rect 35969 520 35970 584
rect 35904 504 35970 520
rect 35904 440 35905 504
rect 35969 440 35970 504
rect 35904 350 35970 440
rect 36030 346 36090 1378
rect 36150 286 36210 1316
rect 36270 346 36330 1378
rect 36390 286 36450 1316
rect 36510 1224 36576 1378
rect 36510 1160 36511 1224
rect 36575 1160 36576 1224
rect 36510 1144 36576 1160
rect 36510 1080 36511 1144
rect 36575 1080 36576 1144
rect 36510 1064 36576 1080
rect 36510 1000 36511 1064
rect 36575 1000 36576 1064
rect 36510 984 36576 1000
rect 36510 920 36511 984
rect 36575 920 36576 984
rect 36510 904 36576 920
rect 36510 840 36511 904
rect 36575 840 36576 904
rect 36510 824 36576 840
rect 36510 760 36511 824
rect 36575 760 36576 824
rect 36510 744 36576 760
rect 36510 680 36511 744
rect 36575 680 36576 744
rect 36510 664 36576 680
rect 36510 600 36511 664
rect 36575 600 36576 664
rect 36510 584 36576 600
rect 36510 520 36511 584
rect 36575 520 36576 584
rect 36510 504 36576 520
rect 36510 440 36511 504
rect 36575 440 36576 504
rect 36510 350 36576 440
rect 36636 346 36696 1378
rect 36756 286 36816 1316
rect 36876 346 36936 1378
rect 36996 286 37056 1316
rect 37116 1224 37182 1378
rect 37116 1160 37117 1224
rect 37181 1160 37182 1224
rect 37116 1144 37182 1160
rect 37116 1080 37117 1144
rect 37181 1080 37182 1144
rect 37116 1064 37182 1080
rect 37116 1000 37117 1064
rect 37181 1000 37182 1064
rect 37116 984 37182 1000
rect 37116 920 37117 984
rect 37181 920 37182 984
rect 37116 904 37182 920
rect 37116 840 37117 904
rect 37181 840 37182 904
rect 37116 824 37182 840
rect 37116 760 37117 824
rect 37181 760 37182 824
rect 37116 744 37182 760
rect 37116 680 37117 744
rect 37181 680 37182 744
rect 37116 664 37182 680
rect 37116 600 37117 664
rect 37181 600 37182 664
rect 37116 584 37182 600
rect 37116 520 37117 584
rect 37181 520 37182 584
rect 37116 504 37182 520
rect 37116 440 37117 504
rect 37181 440 37182 504
rect 37116 350 37182 440
rect 37242 346 37302 1378
rect 37362 286 37422 1316
rect 37482 346 37542 1378
rect 37602 286 37662 1316
rect 37722 1224 37788 1378
rect 37722 1160 37723 1224
rect 37787 1160 37788 1224
rect 37722 1144 37788 1160
rect 37722 1080 37723 1144
rect 37787 1080 37788 1144
rect 37722 1064 37788 1080
rect 37722 1000 37723 1064
rect 37787 1000 37788 1064
rect 37722 984 37788 1000
rect 37722 920 37723 984
rect 37787 920 37788 984
rect 37722 904 37788 920
rect 37722 840 37723 904
rect 37787 840 37788 904
rect 37722 824 37788 840
rect 37722 760 37723 824
rect 37787 760 37788 824
rect 37722 744 37788 760
rect 37722 680 37723 744
rect 37787 680 37788 744
rect 37722 664 37788 680
rect 37722 600 37723 664
rect 37787 600 37788 664
rect 37722 584 37788 600
rect 37722 520 37723 584
rect 37787 520 37788 584
rect 37722 504 37788 520
rect 37722 440 37723 504
rect 37787 440 37788 504
rect 37722 350 37788 440
rect 37848 346 37908 1378
rect 37968 286 38028 1316
rect 38088 346 38148 1378
rect 38208 286 38268 1316
rect 38328 1224 38394 1378
rect 38328 1160 38329 1224
rect 38393 1160 38394 1224
rect 38328 1144 38394 1160
rect 38328 1080 38329 1144
rect 38393 1080 38394 1144
rect 38328 1064 38394 1080
rect 38328 1000 38329 1064
rect 38393 1000 38394 1064
rect 38328 984 38394 1000
rect 38328 920 38329 984
rect 38393 920 38394 984
rect 38328 904 38394 920
rect 38328 840 38329 904
rect 38393 840 38394 904
rect 38328 824 38394 840
rect 38328 760 38329 824
rect 38393 760 38394 824
rect 38328 744 38394 760
rect 38328 680 38329 744
rect 38393 680 38394 744
rect 38328 664 38394 680
rect 38328 600 38329 664
rect 38393 600 38394 664
rect 38328 584 38394 600
rect 38328 520 38329 584
rect 38393 520 38394 584
rect 38328 504 38394 520
rect 38328 440 38329 504
rect 38393 440 38394 504
rect 38328 350 38394 440
rect 38454 346 38514 1378
rect 38574 286 38634 1316
rect 38694 346 38754 1378
rect 38814 286 38874 1316
rect 38934 1224 39000 1378
rect 38934 1160 38935 1224
rect 38999 1160 39000 1224
rect 38934 1144 39000 1160
rect 38934 1080 38935 1144
rect 38999 1080 39000 1144
rect 38934 1064 39000 1080
rect 38934 1000 38935 1064
rect 38999 1000 39000 1064
rect 38934 984 39000 1000
rect 38934 920 38935 984
rect 38999 920 39000 984
rect 38934 904 39000 920
rect 38934 840 38935 904
rect 38999 840 39000 904
rect 38934 824 39000 840
rect 38934 760 38935 824
rect 38999 760 39000 824
rect 38934 744 39000 760
rect 38934 680 38935 744
rect 38999 680 39000 744
rect 38934 664 39000 680
rect 38934 600 38935 664
rect 38999 600 39000 664
rect 38934 584 39000 600
rect 38934 520 38935 584
rect 38999 520 39000 584
rect 38934 504 39000 520
rect 38934 440 38935 504
rect 38999 440 39000 504
rect 38934 350 39000 440
rect 39060 346 39120 1378
rect 39180 286 39240 1316
rect 39300 346 39360 1378
rect 39420 286 39480 1316
rect 39540 1224 39606 1378
rect 39540 1160 39541 1224
rect 39605 1160 39606 1224
rect 39540 1144 39606 1160
rect 39540 1080 39541 1144
rect 39605 1080 39606 1144
rect 39540 1064 39606 1080
rect 39540 1000 39541 1064
rect 39605 1000 39606 1064
rect 39540 984 39606 1000
rect 39540 920 39541 984
rect 39605 920 39606 984
rect 39540 904 39606 920
rect 39540 840 39541 904
rect 39605 840 39606 904
rect 39540 824 39606 840
rect 39540 760 39541 824
rect 39605 760 39606 824
rect 39540 744 39606 760
rect 39540 680 39541 744
rect 39605 680 39606 744
rect 39540 664 39606 680
rect 39540 600 39541 664
rect 39605 600 39606 664
rect 39540 584 39606 600
rect 39540 520 39541 584
rect 39605 520 39606 584
rect 39540 504 39606 520
rect 39540 440 39541 504
rect 39605 440 39606 504
rect 39540 350 39606 440
rect -459 284 213 286
rect -459 220 -355 284
rect -291 220 -275 284
rect -211 220 -195 284
rect -131 220 -115 284
rect -51 220 -35 284
rect 29 220 45 284
rect 109 220 213 284
rect -459 218 213 220
rect 524 284 1027 286
rect 524 220 539 284
rect 603 220 619 284
rect 683 220 699 284
rect 763 220 779 284
rect 843 220 859 284
rect 923 220 1027 284
rect 524 218 1027 220
rect 1267 284 1717 286
rect 1954 284 2545 286
rect 1267 220 1371 284
rect 1435 220 1451 284
rect 1515 220 1531 284
rect 1595 220 1611 284
rect 1675 220 1691 284
rect 1954 220 1977 284
rect 2041 220 2057 284
rect 2121 220 2137 284
rect 2201 220 2217 284
rect 2281 220 2297 284
rect 2361 220 2377 284
rect 2441 220 2545 284
rect 1267 218 1717 220
rect 1954 218 2545 220
rect 2801 284 3301 286
rect 3538 284 5291 286
rect 2801 220 2905 284
rect 2969 220 2985 284
rect 3049 220 3065 284
rect 3129 220 3145 284
rect 3209 220 3225 284
rect 3289 220 3301 284
rect 3575 220 3591 284
rect 3655 220 3671 284
rect 3735 220 3751 284
rect 3815 220 3831 284
rect 3895 220 3911 284
rect 3975 220 4117 284
rect 4181 220 4197 284
rect 4261 220 4277 284
rect 4341 220 4357 284
rect 4421 220 4437 284
rect 4501 220 4517 284
rect 4581 220 4723 284
rect 4787 220 4803 284
rect 4867 220 4883 284
rect 4947 220 4963 284
rect 5027 220 5043 284
rect 5107 220 5123 284
rect 5187 220 5291 284
rect 2801 218 3301 220
rect 3538 218 5291 220
rect 5352 218 5394 286
rect 5631 284 10266 286
rect 5680 220 5696 284
rect 5760 220 5776 284
rect 5840 220 5856 284
rect 5920 220 6062 284
rect 6126 220 6142 284
rect 6206 220 6222 284
rect 6286 220 6302 284
rect 6366 220 6382 284
rect 6446 220 6462 284
rect 6526 220 6668 284
rect 6732 220 6748 284
rect 6812 220 6828 284
rect 6892 220 6908 284
rect 6972 220 6988 284
rect 7052 220 7068 284
rect 7132 220 7274 284
rect 7338 220 7354 284
rect 7418 220 7434 284
rect 7498 220 7514 284
rect 7578 220 7594 284
rect 7658 220 7674 284
rect 7738 220 7880 284
rect 7944 220 7960 284
rect 8024 220 8040 284
rect 8104 220 8120 284
rect 8184 220 8200 284
rect 8264 220 8280 284
rect 8344 220 8486 284
rect 8550 220 8566 284
rect 8630 220 8646 284
rect 8710 220 8726 284
rect 8790 220 8806 284
rect 8870 220 8886 284
rect 8950 220 9092 284
rect 9156 220 9172 284
rect 9236 220 9252 284
rect 9316 220 9332 284
rect 9396 220 9412 284
rect 9476 220 9492 284
rect 9556 220 9698 284
rect 9762 220 9778 284
rect 9842 220 9858 284
rect 9922 220 9938 284
rect 10002 220 10018 284
rect 10082 220 10098 284
rect 10162 220 10266 284
rect 5631 218 10266 220
rect 10326 218 10368 286
rect 10605 284 20088 286
rect 10654 220 10670 284
rect 10734 220 10750 284
rect 10814 220 10830 284
rect 10894 220 11036 284
rect 11100 220 11116 284
rect 11180 220 11196 284
rect 11260 220 11276 284
rect 11340 220 11356 284
rect 11420 220 11436 284
rect 11500 220 11642 284
rect 11706 220 11722 284
rect 11786 220 11802 284
rect 11866 220 11882 284
rect 11946 220 11962 284
rect 12026 220 12042 284
rect 12106 220 12248 284
rect 12312 220 12328 284
rect 12392 220 12408 284
rect 12472 220 12488 284
rect 12552 220 12568 284
rect 12632 220 12648 284
rect 12712 220 12854 284
rect 12918 220 12934 284
rect 12998 220 13014 284
rect 13078 220 13094 284
rect 13158 220 13174 284
rect 13238 220 13254 284
rect 13318 220 13460 284
rect 13524 220 13540 284
rect 13604 220 13620 284
rect 13684 220 13700 284
rect 13764 220 13780 284
rect 13844 220 13860 284
rect 13924 220 14066 284
rect 14130 220 14146 284
rect 14210 220 14226 284
rect 14290 220 14306 284
rect 14370 220 14386 284
rect 14450 220 14466 284
rect 14530 220 14672 284
rect 14736 220 14752 284
rect 14816 220 14832 284
rect 14896 220 14912 284
rect 14976 220 14992 284
rect 15056 220 15072 284
rect 15136 220 15278 284
rect 15342 220 15358 284
rect 15422 220 15438 284
rect 15502 220 15518 284
rect 15582 220 15598 284
rect 15662 220 15678 284
rect 15742 220 15884 284
rect 15948 220 15964 284
rect 16028 220 16044 284
rect 16108 220 16124 284
rect 16188 220 16204 284
rect 16268 220 16284 284
rect 16348 220 16490 284
rect 16554 220 16570 284
rect 16634 220 16650 284
rect 16714 220 16730 284
rect 16794 220 16810 284
rect 16874 220 16890 284
rect 16954 220 17096 284
rect 17160 220 17176 284
rect 17240 220 17256 284
rect 17320 220 17336 284
rect 17400 220 17416 284
rect 17480 220 17496 284
rect 17560 220 17702 284
rect 17766 220 17782 284
rect 17846 220 17862 284
rect 17926 220 17942 284
rect 18006 220 18022 284
rect 18086 220 18102 284
rect 18166 220 18308 284
rect 18372 220 18388 284
rect 18452 220 18468 284
rect 18532 220 18548 284
rect 18612 220 18628 284
rect 18692 220 18708 284
rect 18772 220 18914 284
rect 18978 220 18994 284
rect 19058 220 19074 284
rect 19138 220 19154 284
rect 19218 220 19234 284
rect 19298 220 19314 284
rect 19378 220 19520 284
rect 19584 220 19600 284
rect 19664 220 19680 284
rect 19744 220 19760 284
rect 19824 220 19840 284
rect 19904 220 19920 284
rect 19984 220 20088 284
rect 10605 218 20088 220
rect 20148 284 39298 286
rect 20148 220 20252 284
rect 20316 220 20332 284
rect 20396 220 20412 284
rect 20476 220 20492 284
rect 20556 220 20572 284
rect 20636 220 20652 284
rect 20716 220 20858 284
rect 20922 220 20938 284
rect 21002 220 21018 284
rect 21082 220 21098 284
rect 21162 220 21178 284
rect 21242 220 21258 284
rect 21322 220 21464 284
rect 21528 220 21544 284
rect 21608 220 21624 284
rect 21688 220 21704 284
rect 21768 220 21784 284
rect 21848 220 21864 284
rect 21928 220 22070 284
rect 22134 220 22150 284
rect 22214 220 22230 284
rect 22294 220 22310 284
rect 22374 220 22390 284
rect 22454 220 22470 284
rect 22534 220 22676 284
rect 22740 220 22756 284
rect 22820 220 22836 284
rect 22900 220 22916 284
rect 22980 220 22996 284
rect 23060 220 23076 284
rect 23140 220 23282 284
rect 23346 220 23362 284
rect 23426 220 23442 284
rect 23506 220 23522 284
rect 23586 220 23602 284
rect 23666 220 23682 284
rect 23746 220 23888 284
rect 23952 220 23968 284
rect 24032 220 24048 284
rect 24112 220 24128 284
rect 24192 220 24208 284
rect 24272 220 24288 284
rect 24352 220 24494 284
rect 24558 220 24574 284
rect 24638 220 24654 284
rect 24718 220 24734 284
rect 24798 220 24814 284
rect 24878 220 24894 284
rect 24958 220 25100 284
rect 25164 220 25180 284
rect 25244 220 25260 284
rect 25324 220 25340 284
rect 25404 220 25420 284
rect 25484 220 25500 284
rect 25564 220 25706 284
rect 25770 220 25786 284
rect 25850 220 25866 284
rect 25930 220 25946 284
rect 26010 220 26026 284
rect 26090 220 26106 284
rect 26170 220 26312 284
rect 26376 220 26392 284
rect 26456 220 26472 284
rect 26536 220 26552 284
rect 26616 220 26632 284
rect 26696 220 26712 284
rect 26776 220 26918 284
rect 26982 220 26998 284
rect 27062 220 27078 284
rect 27142 220 27158 284
rect 27222 220 27238 284
rect 27302 220 27318 284
rect 27382 220 27524 284
rect 27588 220 27604 284
rect 27668 220 27684 284
rect 27748 220 27764 284
rect 27828 220 27844 284
rect 27908 220 27924 284
rect 27988 220 28130 284
rect 28194 220 28210 284
rect 28274 220 28290 284
rect 28354 220 28370 284
rect 28434 220 28450 284
rect 28514 220 28530 284
rect 28594 220 28736 284
rect 28800 220 28816 284
rect 28880 220 28896 284
rect 28960 220 28976 284
rect 29040 220 29056 284
rect 29120 220 29136 284
rect 29200 220 29342 284
rect 29406 220 29422 284
rect 29486 220 29502 284
rect 29566 220 29582 284
rect 29646 220 29662 284
rect 29726 220 29742 284
rect 29806 220 29948 284
rect 30012 220 30028 284
rect 30092 220 30108 284
rect 30172 220 30188 284
rect 30252 220 30268 284
rect 30332 220 30348 284
rect 30412 220 30554 284
rect 30618 220 30634 284
rect 30698 220 30714 284
rect 30778 220 30794 284
rect 30858 220 30874 284
rect 30938 220 30954 284
rect 31018 220 31160 284
rect 31224 220 31240 284
rect 31304 220 31320 284
rect 31384 220 31400 284
rect 31464 220 31480 284
rect 31544 220 31560 284
rect 31624 220 31766 284
rect 31830 220 31846 284
rect 31910 220 31926 284
rect 31990 220 32006 284
rect 32070 220 32086 284
rect 32150 220 32166 284
rect 32230 220 32372 284
rect 32436 220 32452 284
rect 32516 220 32532 284
rect 32596 220 32612 284
rect 32676 220 32692 284
rect 32756 220 32772 284
rect 32836 220 32978 284
rect 33042 220 33058 284
rect 33122 220 33138 284
rect 33202 220 33218 284
rect 33282 220 33298 284
rect 33362 220 33378 284
rect 33442 220 33584 284
rect 33648 220 33664 284
rect 33728 220 33744 284
rect 33808 220 33824 284
rect 33888 220 33904 284
rect 33968 220 33984 284
rect 34048 220 34190 284
rect 34254 220 34270 284
rect 34334 220 34350 284
rect 34414 220 34430 284
rect 34494 220 34510 284
rect 34574 220 34590 284
rect 34654 220 34796 284
rect 34860 220 34876 284
rect 34940 220 34956 284
rect 35020 220 35036 284
rect 35100 220 35116 284
rect 35180 220 35196 284
rect 35260 220 35402 284
rect 35466 220 35482 284
rect 35546 220 35562 284
rect 35626 220 35642 284
rect 35706 220 35722 284
rect 35786 220 35802 284
rect 35866 220 36008 284
rect 36072 220 36088 284
rect 36152 220 36168 284
rect 36232 220 36248 284
rect 36312 220 36328 284
rect 36392 220 36408 284
rect 36472 220 36614 284
rect 36678 220 36694 284
rect 36758 220 36774 284
rect 36838 220 36854 284
rect 36918 220 36934 284
rect 36998 220 37014 284
rect 37078 220 37220 284
rect 37284 220 37300 284
rect 37364 220 37380 284
rect 37444 220 37460 284
rect 37524 220 37540 284
rect 37604 220 37620 284
rect 37684 220 37826 284
rect 37890 220 37906 284
rect 37970 220 37986 284
rect 38050 220 38066 284
rect 38130 220 38146 284
rect 38210 220 38226 284
rect 38290 220 38432 284
rect 38496 220 38512 284
rect 38576 220 38592 284
rect 38656 220 38672 284
rect 38736 220 38752 284
rect 38816 220 38832 284
rect 38896 220 39038 284
rect 39102 220 39118 284
rect 39182 220 39198 284
rect 39262 220 39278 284
rect 20148 218 39298 220
rect 39534 218 39606 286
<< via4 >>
rect 287 5092 524 5262
rect 287 5028 459 5092
rect 459 5028 523 5092
rect 523 5028 524 5092
rect 287 5026 524 5028
rect 1717 5092 1954 5262
rect 1717 5028 1755 5092
rect 1755 5028 1771 5092
rect 1771 5028 1835 5092
rect 1835 5028 1954 5092
rect 1717 5026 1954 5028
rect 3301 5092 3538 5262
rect 3301 5028 3305 5092
rect 3305 5028 3369 5092
rect 3369 5028 3511 5092
rect 3511 5028 3538 5092
rect 3301 5026 3538 5028
rect 5394 5092 5631 5262
rect 5394 5028 5456 5092
rect 5456 5028 5520 5092
rect 5520 5028 5536 5092
rect 5536 5028 5600 5092
rect 5600 5028 5616 5092
rect 5616 5028 5631 5092
rect 5394 5026 5631 5028
rect 10368 5092 10605 5262
rect 10368 5028 10430 5092
rect 10430 5028 10494 5092
rect 10494 5028 10510 5092
rect 10510 5028 10574 5092
rect 10574 5028 10590 5092
rect 10590 5028 10605 5092
rect 10368 5026 10605 5028
rect 39298 5092 39534 5262
rect 39298 5028 39342 5092
rect 39342 5028 39358 5092
rect 39358 5028 39422 5092
rect 39422 5028 39438 5092
rect 39438 5028 39502 5092
rect 39502 5028 39534 5092
rect 39298 5026 39534 5028
rect 287 2772 524 2774
rect 287 2708 459 2772
rect 459 2708 523 2772
rect 523 2708 524 2772
rect 287 2604 524 2708
rect 1717 2772 1954 2774
rect 1717 2708 1755 2772
rect 1755 2708 1771 2772
rect 1771 2708 1835 2772
rect 1835 2708 1954 2772
rect 287 2540 459 2604
rect 459 2540 523 2604
rect 523 2540 524 2604
rect 287 2538 524 2540
rect 1717 2604 1954 2708
rect 3301 2772 3538 2774
rect 3301 2708 3305 2772
rect 3305 2708 3369 2772
rect 3369 2708 3511 2772
rect 3511 2708 3538 2772
rect 1717 2540 1755 2604
rect 1755 2540 1771 2604
rect 1771 2540 1835 2604
rect 1835 2540 1954 2604
rect 1717 2538 1954 2540
rect 3301 2604 3538 2708
rect 5394 2772 5631 2774
rect 5394 2708 5456 2772
rect 5456 2708 5520 2772
rect 5520 2708 5536 2772
rect 5536 2708 5600 2772
rect 5600 2708 5616 2772
rect 5616 2708 5631 2772
rect 3301 2540 3305 2604
rect 3305 2540 3369 2604
rect 3369 2540 3511 2604
rect 3511 2540 3538 2604
rect 3301 2538 3538 2540
rect 5394 2604 5631 2708
rect 10368 2772 10605 2774
rect 10368 2708 10430 2772
rect 10430 2708 10494 2772
rect 10494 2708 10510 2772
rect 10510 2708 10574 2772
rect 10574 2708 10590 2772
rect 10590 2708 10605 2772
rect 5394 2540 5456 2604
rect 5456 2540 5520 2604
rect 5520 2540 5536 2604
rect 5536 2540 5600 2604
rect 5600 2540 5616 2604
rect 5616 2540 5631 2604
rect 5394 2538 5631 2540
rect 10368 2604 10605 2708
rect 39298 2772 39534 2774
rect 39298 2708 39342 2772
rect 39342 2708 39358 2772
rect 39358 2708 39422 2772
rect 39422 2708 39438 2772
rect 39438 2708 39502 2772
rect 39502 2708 39534 2772
rect 10368 2540 10430 2604
rect 10430 2540 10494 2604
rect 10494 2540 10510 2604
rect 10510 2540 10574 2604
rect 10574 2540 10590 2604
rect 10590 2540 10605 2604
rect 10368 2538 10605 2540
rect 39298 2604 39534 2708
rect 39298 2540 39342 2604
rect 39342 2540 39358 2604
rect 39358 2540 39422 2604
rect 39422 2540 39438 2604
rect 39438 2540 39502 2604
rect 39502 2540 39534 2604
rect 39298 2538 39534 2540
rect 287 284 524 286
rect 287 220 459 284
rect 459 220 523 284
rect 523 220 524 284
rect 287 50 524 220
rect 1717 284 1954 286
rect 1717 220 1755 284
rect 1755 220 1771 284
rect 1771 220 1835 284
rect 1835 220 1954 284
rect 1717 50 1954 220
rect 3301 284 3538 286
rect 3301 220 3305 284
rect 3305 220 3369 284
rect 3369 220 3511 284
rect 3511 220 3538 284
rect 3301 50 3538 220
rect 5394 284 5631 286
rect 5394 220 5456 284
rect 5456 220 5520 284
rect 5520 220 5536 284
rect 5536 220 5600 284
rect 5600 220 5616 284
rect 5616 220 5631 284
rect 5394 50 5631 220
rect 10368 284 10605 286
rect 10368 220 10430 284
rect 10430 220 10494 284
rect 10494 220 10510 284
rect 10510 220 10574 284
rect 10574 220 10590 284
rect 10590 220 10605 284
rect 10368 50 10605 220
rect 39298 284 39534 286
rect 39298 220 39342 284
rect 39342 220 39358 284
rect 39358 220 39422 284
rect 39422 220 39438 284
rect 39438 220 39502 284
rect 39502 220 39534 284
rect 39298 50 39534 220
<< metal5 >>
rect 245 5262 565 5300
rect 245 5026 287 5262
rect 524 5026 565 5262
rect 245 2774 565 5026
rect 245 2538 287 2774
rect 524 2538 565 2774
rect 245 286 565 2538
rect 245 50 287 286
rect 524 50 565 286
rect 245 11 565 50
rect 1675 5262 1995 5300
rect 1675 5026 1717 5262
rect 1954 5026 1995 5262
rect 1675 2774 1995 5026
rect 1675 2538 1717 2774
rect 1954 2538 1995 2774
rect 1675 286 1995 2538
rect 1675 50 1717 286
rect 1954 50 1995 286
rect 1675 11 1995 50
rect 3259 5262 3579 5300
rect 3259 5026 3301 5262
rect 3538 5026 3579 5262
rect 3259 2774 3579 5026
rect 3259 2538 3301 2774
rect 3538 2538 3579 2774
rect 3259 286 3579 2538
rect 3259 50 3301 286
rect 3538 50 3579 286
rect 3259 11 3579 50
rect 5352 5262 5672 5300
rect 5352 5026 5394 5262
rect 5631 5026 5672 5262
rect 5352 2774 5672 5026
rect 5352 2538 5394 2774
rect 5631 2538 5672 2774
rect 5352 286 5672 2538
rect 5352 50 5394 286
rect 5631 50 5672 286
rect 5352 11 5672 50
rect 10326 5262 10646 5300
rect 10326 5026 10368 5262
rect 10605 5026 10646 5262
rect 10326 2774 10646 5026
rect 10326 2538 10368 2774
rect 10605 2538 10646 2774
rect 10326 286 10646 2538
rect 10326 50 10368 286
rect 10605 50 10646 286
rect 10326 11 10646 50
rect 39256 5262 39576 5300
rect 39256 5026 39298 5262
rect 39534 5026 39576 5262
rect 39256 2808 39576 5026
rect 39256 2774 39578 2808
rect 39256 2538 39298 2774
rect 39534 2538 39578 2774
rect 39256 2488 39578 2538
rect 39256 320 39576 2488
rect 39256 286 39578 320
rect 39256 50 39298 286
rect 39534 50 39578 286
rect 39256 0 39578 50
<< labels >>
flabel metal4 -209 4434 -158 4641 0 FreeSans 480 0 0 0 t<0>
port 27 nsew
flabel metal4 -205 2058 -161 2188 0 FreeSans 320 0 0 0 tb<0>
port 76 nsew
flabel metal4 -324 3245 -280 3393 0 FreeSans 320 0 0 0 tu
port 90 nsew
flabel poly 2970 6023 3936 6093 0 FreeSans 320 0 0 0 d<3>
port 102 nsew
flabel poly 1437 6023 1891 6093 0 FreeSans 320 0 0 0 d<2>
port 104 nsew
flabel poly 656 5978 726 6110 0 FreeSans 320 0 0 0 d<1>
port 106 nsew
flabel poly -249 5978 -179 6110 0 FreeSans 320 0 0 0 d<0>
port 109 nsew
flabel poly 5521 6023 7511 6093 0 FreeSans 320 0 0 0 d<4>
port 111 nsew
flabel poly 10608 6023 14646 6093 0 FreeSans 320 0 0 0 d<5>
port 113 nsew
flabel poly 20393 6023 28527 6093 0 FreeSans 320 0 0 0 d<6>
port 115 nsew
flabel poly -271 5290 -201 5422 0 FreeSans 320 0 0 0 db<0>
port 117 nsew
flabel poly 657 5290 727 5422 0 FreeSans 320 0 0 0 db<1>
port 119 nsew
flabel poly 1921 5335 2375 5405 0 FreeSans 320 0 0 0 db<2>
port 121 nsew
flabel poly 3540 5335 4506 5405 0 FreeSans 320 0 0 0 db<3>
port 123 nsew
flabel poly 8105 5335 10095 5405 0 FreeSans 320 0 0 0 db<4>
port 125 nsew
flabel poly 15263 5335 19301 5405 0 FreeSans 320 0 0 0 db<5>
port 127 nsew
flabel metal4 -329 832 -283 967 0 FreeSans 320 0 0 0 tub
port 131 nsew
flabel poly 20317 5335 28451 5405 0 FreeSans 320 0 0 0 db<6>
port 133 nsew
flabel metal5 287 5026 524 5262 0 FreeSans 320 0 0 0 t<1>
port 135 nsew
flabel metal5 1717 5026 1954 5262 0 FreeSans 320 0 0 0 t<2>
port 137 nsew
flabel metal5 3301 5026 3538 5262 0 FreeSans 320 0 0 0 t<3>
port 139 nsew
flabel metal5 5394 5026 5631 5262 0 FreeSans 320 0 0 0 t<4>
port 141 nsew
flabel metal5 10368 5026 10605 5262 0 FreeSans 480 0 0 0 t<5>
port 143 nsew
flabel metal5 39298 5026 39534 5262 0 FreeSans 480 0 0 0 t<6>
port 145 nsew
flabel metal5 287 50 524 286 0 FreeSans 480 0 0 0 tb<1>
port 147 nsew
flabel metal5 1717 50 1954 286 0 FreeSans 480 0 0 0 tb<2>
port 149 nsew
flabel metal5 3301 50 3538 286 0 FreeSans 480 0 0 0 tb<3>
port 151 nsew
flabel metal5 5394 50 5631 286 0 FreeSans 480 0 0 0 tb<4>
port 153 nsew
flabel metal5 10368 50 10605 286 0 FreeSans 480 0 0 0 tb<5>
port 155 nsew
flabel metal5 39298 50 39534 286 0 FreeSans 480 0 0 0 tb<6>
port 157 nsew
flabel metal4 29211 5154 29572 5639 0 FreeSans 1600 0 0 0 VSS
port 159 nsew
flabel metal4 29822 5731 30233 6365 0 FreeSans 1600 0 0 0 VDD
port 161 nsew
flabel metal4 29015 5756 29404 6320 0 FreeSans 1600 0 0 0 VREF
port 163 nsew
flabel pwell 17436 1084 17468 1134 0 FreeSans 160 0 0 0 hgu_cdac_8bit_array_2.SUB
flabel metal4 7177 1391 7228 1432 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.drv<15:0>
flabel metal4 35915 1391 35966 1432 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.drv<63:0>
flabel metal4 12152 1392 12207 1431 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.drv<31:0>
flabel via4 5429 126 5596 209 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.tah<15:0>
flabel via4 10396 107 10570 207 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.tah<31:0>
flabel via4 39332 112 39506 212 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.tah<63:0>
flabel metal4 4022 1394 4073 1435 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.drv<7:0>
flabel via4 3335 113 3509 213 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.tah<7:0>
flabel via4 287 50 524 286 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.tah<1:0>
flabel metal4 966 1394 1020 1428 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.drv<1:0>
flabel metal4 -205 1618 -156 1670 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.tah<0>
flabel metal4 -85 1742 -43 1776 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.drv<0>
flabel metal4 1883 1390 1934 1432 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.drv<3:0>
flabel via4 1745 117 1919 217 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.tah<3:0>
flabel metal4 -75 2128 -49 2160 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.x1.CBOT
flabel metal4 -193 1538 -167 1570 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.x1.CTOP
flabel psubdiff -145 1794 -107 1872 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.x1.SUB
flabel psubdiff 29070 1054 29112 1144 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.SUB
flabel metal4 28886 1130 28932 1200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.CTOP
flabel metal4 29004 1804 29050 1874 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.CTOP
flabel metal4 29126 1534 29172 1604 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.CBOT
flabel metal4 20532 968 20558 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[0].CBOT
flabel metal4 20414 378 20440 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[0].CTOP
flabel psubdiff 20462 634 20500 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[0].SUB
flabel metal4 20410 1824 20436 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[1].CBOT
flabel metal4 20528 2414 20554 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[1].CTOP
flabel psubdiff 20468 2112 20506 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[1].SUB
flabel metal4 21138 968 21164 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[2].CBOT
flabel metal4 21020 378 21046 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[2].CTOP
flabel psubdiff 21068 634 21106 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[2].SUB
flabel metal4 21016 1824 21042 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[3].CBOT
flabel metal4 21134 2414 21160 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[3].CTOP
flabel psubdiff 21074 2112 21112 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[3].SUB
flabel metal4 21744 968 21770 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[4].CBOT
flabel metal4 21626 378 21652 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[4].CTOP
flabel psubdiff 21674 634 21712 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[4].SUB
flabel metal4 21622 1824 21648 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[5].CBOT
flabel metal4 21740 2414 21766 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[5].CTOP
flabel psubdiff 21680 2112 21718 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[5].SUB
flabel metal4 22350 968 22376 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[6].CBOT
flabel metal4 22232 378 22258 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[6].CTOP
flabel psubdiff 22280 634 22318 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[6].SUB
flabel metal4 22228 1824 22254 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[7].CBOT
flabel metal4 22346 2414 22372 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[7].CTOP
flabel psubdiff 22286 2112 22324 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[7].SUB
flabel metal4 22956 968 22982 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[8].CBOT
flabel metal4 22838 378 22864 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[8].CTOP
flabel psubdiff 22886 634 22924 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[8].SUB
flabel metal4 22834 1824 22860 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[9].CBOT
flabel metal4 22952 2414 22978 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[9].CTOP
flabel psubdiff 22892 2112 22930 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[9].SUB
flabel metal4 23562 968 23588 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[10].CBOT
flabel metal4 23444 378 23470 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[10].CTOP
flabel psubdiff 23492 634 23530 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[10].SUB
flabel metal4 23440 1824 23466 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[11].CBOT
flabel metal4 23558 2414 23584 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[11].CTOP
flabel psubdiff 23498 2112 23536 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[11].SUB
flabel metal4 24168 968 24194 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[12].CBOT
flabel metal4 24050 378 24076 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[12].CTOP
flabel psubdiff 24098 634 24136 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[12].SUB
flabel metal4 24046 1824 24072 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[13].CBOT
flabel metal4 24164 2414 24190 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[13].CTOP
flabel psubdiff 24104 2112 24142 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[13].SUB
flabel metal4 24774 968 24800 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[14].CBOT
flabel metal4 24656 378 24682 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[14].CTOP
flabel psubdiff 24704 634 24742 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[14].SUB
flabel metal4 24652 1824 24678 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[15].CBOT
flabel metal4 24770 2414 24796 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[15].CTOP
flabel psubdiff 24710 2112 24748 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[15].SUB
flabel metal4 25380 968 25406 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[16].CBOT
flabel metal4 25262 378 25288 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[16].CTOP
flabel psubdiff 25310 634 25348 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[16].SUB
flabel metal4 25258 1824 25284 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[17].CBOT
flabel metal4 25376 2414 25402 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[17].CTOP
flabel psubdiff 25316 2112 25354 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[17].SUB
flabel metal4 25986 968 26012 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[18].CBOT
flabel metal4 25868 378 25894 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[18].CTOP
flabel psubdiff 25916 634 25954 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[18].SUB
flabel metal4 25864 1824 25890 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[19].CBOT
flabel metal4 25982 2414 26008 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[19].CTOP
flabel psubdiff 25922 2112 25960 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[19].SUB
flabel metal4 26592 968 26618 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[20].CBOT
flabel metal4 26474 378 26500 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[20].CTOP
flabel psubdiff 26522 634 26560 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[20].SUB
flabel metal4 26470 1824 26496 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[21].CBOT
flabel metal4 26588 2414 26614 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[21].CTOP
flabel psubdiff 26528 2112 26566 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[21].SUB
flabel metal4 27198 968 27224 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[22].CBOT
flabel metal4 27080 378 27106 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[22].CTOP
flabel psubdiff 27128 634 27166 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[22].SUB
flabel metal4 27076 1824 27102 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[23].CBOT
flabel metal4 27194 2414 27220 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[23].CTOP
flabel psubdiff 27134 2112 27172 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[23].SUB
flabel metal4 27804 968 27830 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[24].CBOT
flabel metal4 27686 378 27712 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[24].CTOP
flabel psubdiff 27734 634 27772 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[24].SUB
flabel metal4 27682 1824 27708 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[25].CBOT
flabel metal4 27800 2414 27826 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[25].CTOP
flabel psubdiff 27740 2112 27778 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[25].SUB
flabel metal4 28410 968 28436 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[26].CBOT
flabel metal4 28292 378 28318 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[26].CTOP
flabel psubdiff 28340 634 28378 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[26].SUB
flabel metal4 28288 1824 28314 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[27].CBOT
flabel metal4 28406 2414 28432 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[27].CTOP
flabel psubdiff 28346 2112 28384 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[27].SUB
flabel metal4 29016 968 29042 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[28].CBOT
flabel metal4 28898 378 28924 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[28].CTOP
flabel psubdiff 28946 634 28984 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[28].SUB
flabel metal4 28894 1824 28920 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[29].CBOT
flabel metal4 29012 2414 29038 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[29].CTOP
flabel psubdiff 28952 2112 28990 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[29].SUB
flabel metal4 29622 968 29648 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[30].CBOT
flabel metal4 29504 378 29530 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[30].CTOP
flabel psubdiff 29552 634 29590 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[30].SUB
flabel metal4 29500 1824 29526 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[31].CBOT
flabel metal4 29618 2414 29644 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[31].CTOP
flabel psubdiff 29558 2112 29596 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[31].SUB
flabel metal4 30228 968 30254 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[32].CBOT
flabel metal4 30110 378 30136 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[32].CTOP
flabel psubdiff 30158 634 30196 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[32].SUB
flabel metal4 30106 1824 30132 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[33].CBOT
flabel metal4 30224 2414 30250 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[33].CTOP
flabel psubdiff 30164 2112 30202 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[33].SUB
flabel metal4 30834 968 30860 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[34].CBOT
flabel metal4 30716 378 30742 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[34].CTOP
flabel psubdiff 30764 634 30802 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[34].SUB
flabel metal4 30712 1824 30738 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[35].CBOT
flabel metal4 30830 2414 30856 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[35].CTOP
flabel psubdiff 30770 2112 30808 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[35].SUB
flabel metal4 31440 968 31466 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[36].CBOT
flabel metal4 31322 378 31348 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[36].CTOP
flabel psubdiff 31370 634 31408 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[36].SUB
flabel metal4 31318 1824 31344 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[37].CBOT
flabel metal4 31436 2414 31462 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[37].CTOP
flabel psubdiff 31376 2112 31414 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[37].SUB
flabel metal4 32046 968 32072 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[38].CBOT
flabel metal4 31928 378 31954 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[38].CTOP
flabel psubdiff 31976 634 32014 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[38].SUB
flabel metal4 31924 1824 31950 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[39].CBOT
flabel metal4 32042 2414 32068 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[39].CTOP
flabel psubdiff 31982 2112 32020 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[39].SUB
flabel metal4 32652 968 32678 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[40].CBOT
flabel metal4 32534 378 32560 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[40].CTOP
flabel psubdiff 32582 634 32620 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[40].SUB
flabel metal4 32530 1824 32556 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[41].CBOT
flabel metal4 32648 2414 32674 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[41].CTOP
flabel psubdiff 32588 2112 32626 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[41].SUB
flabel metal4 33258 968 33284 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[42].CBOT
flabel metal4 33140 378 33166 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[42].CTOP
flabel psubdiff 33188 634 33226 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[42].SUB
flabel metal4 33136 1824 33162 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[43].CBOT
flabel metal4 33254 2414 33280 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[43].CTOP
flabel psubdiff 33194 2112 33232 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[43].SUB
flabel metal4 33864 968 33890 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[44].CBOT
flabel metal4 33746 378 33772 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[44].CTOP
flabel psubdiff 33794 634 33832 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[44].SUB
flabel metal4 33742 1824 33768 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[45].CBOT
flabel metal4 33860 2414 33886 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[45].CTOP
flabel psubdiff 33800 2112 33838 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[45].SUB
flabel metal4 34470 968 34496 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[46].CBOT
flabel metal4 34352 378 34378 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[46].CTOP
flabel psubdiff 34400 634 34438 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[46].SUB
flabel metal4 34348 1824 34374 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[47].CBOT
flabel metal4 34466 2414 34492 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[47].CTOP
flabel psubdiff 34406 2112 34444 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[47].SUB
flabel metal4 35076 968 35102 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[48].CBOT
flabel metal4 34958 378 34984 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[48].CTOP
flabel psubdiff 35006 634 35044 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[48].SUB
flabel metal4 34954 1824 34980 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[49].CBOT
flabel metal4 35072 2414 35098 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[49].CTOP
flabel psubdiff 35012 2112 35050 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[49].SUB
flabel metal4 35682 968 35708 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[50].CBOT
flabel metal4 35564 378 35590 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[50].CTOP
flabel psubdiff 35612 634 35650 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[50].SUB
flabel metal4 35560 1824 35586 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[51].CBOT
flabel metal4 35678 2414 35704 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[51].CTOP
flabel psubdiff 35618 2112 35656 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[51].SUB
flabel metal4 36288 968 36314 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[52].CBOT
flabel metal4 36170 378 36196 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[52].CTOP
flabel psubdiff 36218 634 36256 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[52].SUB
flabel metal4 36166 1824 36192 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[53].CBOT
flabel metal4 36284 2414 36310 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[53].CTOP
flabel psubdiff 36224 2112 36262 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[53].SUB
flabel metal4 36894 968 36920 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[54].CBOT
flabel metal4 36776 378 36802 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[54].CTOP
flabel psubdiff 36824 634 36862 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[54].SUB
flabel metal4 36772 1824 36798 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[55].CBOT
flabel metal4 36890 2414 36916 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[55].CTOP
flabel psubdiff 36830 2112 36868 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[55].SUB
flabel metal4 37500 968 37526 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[56].CBOT
flabel metal4 37382 378 37408 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[56].CTOP
flabel psubdiff 37430 634 37468 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[56].SUB
flabel metal4 37378 1824 37404 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[57].CBOT
flabel metal4 37496 2414 37522 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[57].CTOP
flabel psubdiff 37436 2112 37474 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[57].SUB
flabel metal4 38106 968 38132 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[58].CBOT
flabel metal4 37988 378 38014 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[58].CTOP
flabel psubdiff 38036 634 38074 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[58].SUB
flabel metal4 37984 1824 38010 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[59].CBOT
flabel metal4 38102 2414 38128 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[59].CTOP
flabel psubdiff 38042 2112 38080 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[59].SUB
flabel metal4 38712 968 38738 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[60].CBOT
flabel metal4 38594 378 38620 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[60].CTOP
flabel psubdiff 38642 634 38680 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[60].SUB
flabel metal4 38590 1824 38616 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[61].CBOT
flabel metal4 38708 2414 38734 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[61].CTOP
flabel psubdiff 38648 2112 38686 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[61].SUB
flabel metal4 39318 968 39344 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[62].CBOT
flabel metal4 39200 378 39226 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[62].CTOP
flabel psubdiff 39248 634 39286 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[62].SUB
flabel metal4 39196 1824 39222 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[63].CBOT
flabel metal4 39314 2414 39340 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[63].CTOP
flabel psubdiff 39254 2112 39292 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_64_0.x1[63].SUB
flabel psubdiff 14766 1266 14810 1358 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.SUB
flabel metal4 14336 1062 14380 1154 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.CBOT
flabel metal4 14824 1066 14868 1158 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.CTOP
flabel metal4 14702 1586 14746 1678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.CTOP
flabel metal4 19800 968 19826 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[31].CBOT
flabel metal4 19682 378 19708 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[31].CTOP
flabel psubdiff 19730 634 19768 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[31].SUB
flabel metal4 19678 1824 19704 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[30].CBOT
flabel metal4 19796 2414 19822 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[30].CTOP
flabel psubdiff 19736 2112 19774 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[30].SUB
flabel metal4 19194 968 19220 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[29].CBOT
flabel metal4 19076 378 19102 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[29].CTOP
flabel psubdiff 19124 634 19162 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[29].SUB
flabel metal4 19072 1824 19098 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[28].CBOT
flabel metal4 19190 2414 19216 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[28].CTOP
flabel psubdiff 19130 2112 19168 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[28].SUB
flabel metal4 18588 968 18614 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[27].CBOT
flabel metal4 18470 378 18496 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[27].CTOP
flabel psubdiff 18518 634 18556 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[27].SUB
flabel metal4 18466 1824 18492 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[26].CBOT
flabel metal4 18584 2414 18610 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[26].CTOP
flabel psubdiff 18524 2112 18562 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[26].SUB
flabel metal4 17982 968 18008 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[25].CBOT
flabel metal4 17864 378 17890 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[25].CTOP
flabel psubdiff 17912 634 17950 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[25].SUB
flabel metal4 17860 1824 17886 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[24].CBOT
flabel metal4 17978 2414 18004 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[24].CTOP
flabel psubdiff 17918 2112 17956 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[24].SUB
flabel metal4 17376 968 17402 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[23].CBOT
flabel metal4 17258 378 17284 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[23].CTOP
flabel psubdiff 17306 634 17344 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[23].SUB
flabel metal4 17254 1824 17280 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[22].CBOT
flabel metal4 17372 2414 17398 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[22].CTOP
flabel psubdiff 17312 2112 17350 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[22].SUB
flabel metal4 16770 968 16796 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[21].CBOT
flabel metal4 16652 378 16678 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[21].CTOP
flabel psubdiff 16700 634 16738 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[21].SUB
flabel metal4 16648 1824 16674 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[20].CBOT
flabel metal4 16766 2414 16792 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[20].CTOP
flabel psubdiff 16706 2112 16744 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[20].SUB
flabel metal4 16164 968 16190 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[19].CBOT
flabel metal4 16046 378 16072 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[19].CTOP
flabel psubdiff 16094 634 16132 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[19].SUB
flabel metal4 16042 1824 16068 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[18].CBOT
flabel metal4 16160 2414 16186 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[18].CTOP
flabel psubdiff 16100 2112 16138 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[18].SUB
flabel metal4 15558 968 15584 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[17].CBOT
flabel metal4 15440 378 15466 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[17].CTOP
flabel psubdiff 15488 634 15526 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[17].SUB
flabel metal4 15436 1824 15462 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[16].CBOT
flabel metal4 15554 2414 15580 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[16].CTOP
flabel psubdiff 15494 2112 15532 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[16].SUB
flabel metal4 14952 968 14978 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[15].CBOT
flabel metal4 14834 378 14860 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[15].CTOP
flabel psubdiff 14882 634 14920 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[15].SUB
flabel metal4 14830 1824 14856 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[14].CBOT
flabel metal4 14948 2414 14974 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[14].CTOP
flabel psubdiff 14888 2112 14926 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[14].SUB
flabel metal4 14346 968 14372 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[13].CBOT
flabel metal4 14228 378 14254 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[13].CTOP
flabel psubdiff 14276 634 14314 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[13].SUB
flabel metal4 14224 1824 14250 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[12].CBOT
flabel metal4 14342 2414 14368 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[12].CTOP
flabel psubdiff 14282 2112 14320 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[12].SUB
flabel metal4 13740 968 13766 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[11].CBOT
flabel metal4 13622 378 13648 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[11].CTOP
flabel psubdiff 13670 634 13708 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[11].SUB
flabel metal4 13618 1824 13644 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[10].CBOT
flabel metal4 13736 2414 13762 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[10].CTOP
flabel psubdiff 13676 2112 13714 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[10].SUB
flabel metal4 13134 968 13160 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[9].CBOT
flabel metal4 13016 378 13042 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[9].CTOP
flabel psubdiff 13064 634 13102 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[9].SUB
flabel metal4 13012 1824 13038 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[8].CBOT
flabel metal4 13130 2414 13156 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[8].CTOP
flabel psubdiff 13070 2112 13108 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[8].SUB
flabel metal4 12528 968 12554 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[7].CBOT
flabel metal4 12410 378 12436 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[7].CTOP
flabel psubdiff 12458 634 12496 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[7].SUB
flabel metal4 12406 1824 12432 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[6].CBOT
flabel metal4 12524 2414 12550 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[6].CTOP
flabel psubdiff 12464 2112 12502 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[6].SUB
flabel metal4 11922 968 11948 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[5].CBOT
flabel metal4 11804 378 11830 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[5].CTOP
flabel psubdiff 11852 634 11890 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[5].SUB
flabel metal4 11800 1824 11826 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[4].CBOT
flabel metal4 11918 2414 11944 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[4].CTOP
flabel psubdiff 11858 2112 11896 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[4].SUB
flabel metal4 11316 968 11342 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[3].CBOT
flabel metal4 11198 378 11224 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[3].CTOP
flabel psubdiff 11246 634 11284 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[3].SUB
flabel metal4 11194 1824 11220 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[2].CBOT
flabel metal4 11312 2414 11338 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[2].CTOP
flabel psubdiff 11252 2112 11290 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[2].SUB
flabel metal4 10710 968 10736 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[1].CBOT
flabel metal4 10592 378 10618 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[1].CTOP
flabel psubdiff 10640 634 10678 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[1].SUB
flabel metal4 10588 1824 10614 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[0].CBOT
flabel metal4 10706 2414 10732 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[0].CTOP
flabel psubdiff 10646 2112 10684 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_32_0.x1[0].SUB
flabel metal4 8156 1228 8192 1308 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.CBOT
flabel metal4 7432 1198 7468 1278 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.CTOP
flabel metal4 7546 1570 7590 1652 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.CTOP
flabel psubdiff 7850 1470 7894 1552 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.SUB
flabel metal4 9978 968 10004 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[15].CBOT
flabel metal4 9860 378 9886 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[15].CTOP
flabel psubdiff 9908 634 9946 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[15].SUB
flabel metal4 9856 1824 9882 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[14].CBOT
flabel metal4 9974 2414 10000 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[14].CTOP
flabel psubdiff 9914 2112 9952 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[14].SUB
flabel metal4 9372 968 9398 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[13].CBOT
flabel metal4 9254 378 9280 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[13].CTOP
flabel psubdiff 9302 634 9340 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[13].SUB
flabel metal4 9250 1824 9276 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[12].CBOT
flabel metal4 9368 2414 9394 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[12].CTOP
flabel psubdiff 9308 2112 9346 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[12].SUB
flabel metal4 8766 968 8792 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[11].CBOT
flabel metal4 8648 378 8674 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[11].CTOP
flabel psubdiff 8696 634 8734 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[11].SUB
flabel metal4 8644 1824 8670 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[10].CBOT
flabel metal4 8762 2414 8788 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[10].CTOP
flabel psubdiff 8702 2112 8740 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[10].SUB
flabel metal4 8160 968 8186 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[9].CBOT
flabel metal4 8042 378 8068 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[9].CTOP
flabel psubdiff 8090 634 8128 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[9].SUB
flabel metal4 8038 1824 8064 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[8].CBOT
flabel metal4 8156 2414 8182 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[8].CTOP
flabel psubdiff 8096 2112 8134 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[8].SUB
flabel metal4 7554 968 7580 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[7].CBOT
flabel metal4 7436 378 7462 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[7].CTOP
flabel psubdiff 7484 634 7522 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[7].SUB
flabel metal4 7432 1824 7458 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[6].CBOT
flabel metal4 7550 2414 7576 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[6].CTOP
flabel psubdiff 7490 2112 7528 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[6].SUB
flabel metal4 6948 968 6974 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[5].CBOT
flabel metal4 6830 378 6856 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[5].CTOP
flabel psubdiff 6878 634 6916 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[5].SUB
flabel metal4 6826 1824 6852 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[4].CBOT
flabel metal4 6944 2414 6970 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[4].CTOP
flabel psubdiff 6884 2112 6922 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[4].SUB
flabel metal4 6342 968 6368 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[3].CBOT
flabel metal4 6224 378 6250 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[3].CTOP
flabel psubdiff 6272 634 6310 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[3].SUB
flabel metal4 6220 1824 6246 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[2].CBOT
flabel metal4 6338 2414 6364 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[2].CTOP
flabel psubdiff 6278 2112 6316 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[2].SUB
flabel metal4 5736 968 5762 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[1].CBOT
flabel metal4 5618 378 5644 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[1].CTOP
flabel psubdiff 5666 634 5704 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[1].SUB
flabel metal4 5614 1824 5640 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[0].CBOT
flabel metal4 5732 2414 5758 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[0].CTOP
flabel psubdiff 5672 2112 5710 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_16_0.x1[0].SUB
flabel psubdiff 4207 1266 4251 1366 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.SUB
flabel metal4 4387 1098 4433 1190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.CBOT
flabel metal4 3659 1120 3705 1212 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.CTOP
flabel metal4 3787 1958 3827 2042 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.CTOP
flabel metal4 5003 968 5029 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[7].CBOT
flabel metal4 4885 378 4911 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[7].CTOP
flabel psubdiff 4933 634 4971 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[7].SUB
flabel metal4 4881 1824 4907 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[6].CBOT
flabel metal4 4999 2414 5025 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[6].CTOP
flabel psubdiff 4939 2112 4977 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[6].SUB
flabel metal4 4397 968 4423 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[5].CBOT
flabel metal4 4279 378 4305 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[5].CTOP
flabel psubdiff 4327 634 4365 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[5].SUB
flabel metal4 4275 1824 4301 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[4].CBOT
flabel metal4 4393 2414 4419 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[4].CTOP
flabel psubdiff 4333 2112 4371 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[4].SUB
flabel metal4 3791 968 3817 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[3].CBOT
flabel metal4 3673 378 3699 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[3].CTOP
flabel psubdiff 3721 634 3759 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[3].SUB
flabel metal4 3669 1824 3695 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[2].CBOT
flabel metal4 3787 2414 3813 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[2].CTOP
flabel psubdiff 3727 2112 3765 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[2].SUB
flabel metal4 3185 968 3211 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[1].CBOT
flabel metal4 3067 378 3093 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[1].CTOP
flabel psubdiff 3115 634 3153 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[1].SUB
flabel metal4 3063 1824 3089 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[0].CBOT
flabel metal4 3181 2414 3207 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[0].CTOP
flabel psubdiff 3121 2112 3159 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_8_0.x1[0].SUB
flabel metal4 2245 1326 2297 1366 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT
flabel metal4 1519 1210 1571 1250 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CTOP
flabel psubdiff 2069 1220 2109 1330 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.SUB
flabel metal4 1643 1548 1681 1630 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CTOP
flabel metal4 2257 968 2283 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[3].CBOT
flabel metal4 2139 378 2165 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[3].CTOP
flabel psubdiff 2187 634 2225 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[3].SUB
flabel metal4 2135 1824 2161 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[2].CBOT
flabel metal4 2253 2414 2279 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[2].CTOP
flabel psubdiff 2193 2112 2231 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[2].SUB
flabel metal4 1651 968 1677 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[1].CBOT
flabel metal4 1533 378 1559 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[1].CTOP
flabel psubdiff 1581 634 1619 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[1].SUB
flabel metal4 1529 1824 1555 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[0].CBOT
flabel metal4 1647 2414 1673 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[0].CTOP
flabel psubdiff 1587 2112 1625 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.x1[0].SUB
flabel psubdiff 669 1127 717 1241 0 FreeSans 160 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_2_0.SUB
flabel metal4 733 1122 769 1212 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_2_0.CBOT
flabel metal4 613 680 649 782 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_2_0.CTOP
flabel metal4 731 2264 771 2342 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_2_0.CTOP
flabel metal4 739 968 765 1000 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_2_0.x2.CBOT
flabel metal4 621 378 647 410 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_2_0.x2.CTOP
flabel psubdiff 669 634 707 712 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_2_0.x2.SUB
flabel metal4 617 1824 643 1856 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_2_0.x1.CBOT
flabel metal4 735 2414 761 2446 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_2_0.x1.CTOP
flabel psubdiff 675 2112 713 2190 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_2.hgu_cdac_cap_2_0.x1.SUB
flabel pwell 17436 3572 17468 3622 0 FreeSans 160 0 0 0 hgu_cdac_8bit_array_3.SUB
flabel metal4 7177 3879 7228 3920 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.drv<15:0>
flabel metal4 35915 3879 35966 3920 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.drv<63:0>
flabel metal4 12152 3880 12207 3919 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.drv<31:0>
flabel via4 5429 2614 5596 2697 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.tah<15:0>
flabel via4 10396 2595 10570 2695 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.tah<31:0>
flabel via4 39332 2600 39506 2700 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.tah<63:0>
flabel metal4 4022 3882 4073 3923 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.drv<7:0>
flabel via4 3335 2601 3509 2701 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.tah<7:0>
flabel via4 287 2538 524 2774 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.tah<1:0>
flabel metal4 966 3882 1020 3916 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.drv<1:0>
flabel metal4 -205 4106 -156 4158 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.tah<0>
flabel metal4 -85 4230 -43 4264 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.drv<0>
flabel metal4 1883 3878 1934 3920 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.drv<3:0>
flabel via4 1745 2605 1919 2705 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.tah<3:0>
flabel metal4 -75 4616 -49 4648 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.x1.CBOT
flabel metal4 -193 4026 -167 4058 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.x1.CTOP
flabel psubdiff -145 4282 -107 4360 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.x1.SUB
flabel psubdiff 29070 3542 29112 3632 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.SUB
flabel metal4 28886 3618 28932 3688 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.CTOP
flabel metal4 29004 4292 29050 4362 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.CTOP
flabel metal4 29126 4022 29172 4092 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.CBOT
flabel metal4 20532 3456 20558 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[0].CBOT
flabel metal4 20414 2866 20440 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[0].CTOP
flabel psubdiff 20462 3122 20500 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[0].SUB
flabel metal4 20410 4312 20436 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[1].CBOT
flabel metal4 20528 4902 20554 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[1].CTOP
flabel psubdiff 20468 4600 20506 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[1].SUB
flabel metal4 21138 3456 21164 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[2].CBOT
flabel metal4 21020 2866 21046 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[2].CTOP
flabel psubdiff 21068 3122 21106 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[2].SUB
flabel metal4 21016 4312 21042 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[3].CBOT
flabel metal4 21134 4902 21160 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[3].CTOP
flabel psubdiff 21074 4600 21112 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[3].SUB
flabel metal4 21744 3456 21770 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[4].CBOT
flabel metal4 21626 2866 21652 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[4].CTOP
flabel psubdiff 21674 3122 21712 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[4].SUB
flabel metal4 21622 4312 21648 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[5].CBOT
flabel metal4 21740 4902 21766 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[5].CTOP
flabel psubdiff 21680 4600 21718 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[5].SUB
flabel metal4 22350 3456 22376 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[6].CBOT
flabel metal4 22232 2866 22258 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[6].CTOP
flabel psubdiff 22280 3122 22318 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[6].SUB
flabel metal4 22228 4312 22254 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[7].CBOT
flabel metal4 22346 4902 22372 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[7].CTOP
flabel psubdiff 22286 4600 22324 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[7].SUB
flabel metal4 22956 3456 22982 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[8].CBOT
flabel metal4 22838 2866 22864 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[8].CTOP
flabel psubdiff 22886 3122 22924 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[8].SUB
flabel metal4 22834 4312 22860 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[9].CBOT
flabel metal4 22952 4902 22978 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[9].CTOP
flabel psubdiff 22892 4600 22930 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[9].SUB
flabel metal4 23562 3456 23588 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[10].CBOT
flabel metal4 23444 2866 23470 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[10].CTOP
flabel psubdiff 23492 3122 23530 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[10].SUB
flabel metal4 23440 4312 23466 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[11].CBOT
flabel metal4 23558 4902 23584 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[11].CTOP
flabel psubdiff 23498 4600 23536 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[11].SUB
flabel metal4 24168 3456 24194 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[12].CBOT
flabel metal4 24050 2866 24076 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[12].CTOP
flabel psubdiff 24098 3122 24136 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[12].SUB
flabel metal4 24046 4312 24072 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[13].CBOT
flabel metal4 24164 4902 24190 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[13].CTOP
flabel psubdiff 24104 4600 24142 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[13].SUB
flabel metal4 24774 3456 24800 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[14].CBOT
flabel metal4 24656 2866 24682 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[14].CTOP
flabel psubdiff 24704 3122 24742 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[14].SUB
flabel metal4 24652 4312 24678 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[15].CBOT
flabel metal4 24770 4902 24796 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[15].CTOP
flabel psubdiff 24710 4600 24748 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[15].SUB
flabel metal4 25380 3456 25406 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[16].CBOT
flabel metal4 25262 2866 25288 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[16].CTOP
flabel psubdiff 25310 3122 25348 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[16].SUB
flabel metal4 25258 4312 25284 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[17].CBOT
flabel metal4 25376 4902 25402 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[17].CTOP
flabel psubdiff 25316 4600 25354 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[17].SUB
flabel metal4 25986 3456 26012 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[18].CBOT
flabel metal4 25868 2866 25894 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[18].CTOP
flabel psubdiff 25916 3122 25954 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[18].SUB
flabel metal4 25864 4312 25890 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[19].CBOT
flabel metal4 25982 4902 26008 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[19].CTOP
flabel psubdiff 25922 4600 25960 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[19].SUB
flabel metal4 26592 3456 26618 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[20].CBOT
flabel metal4 26474 2866 26500 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[20].CTOP
flabel psubdiff 26522 3122 26560 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[20].SUB
flabel metal4 26470 4312 26496 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[21].CBOT
flabel metal4 26588 4902 26614 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[21].CTOP
flabel psubdiff 26528 4600 26566 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[21].SUB
flabel metal4 27198 3456 27224 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[22].CBOT
flabel metal4 27080 2866 27106 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[22].CTOP
flabel psubdiff 27128 3122 27166 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[22].SUB
flabel metal4 27076 4312 27102 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[23].CBOT
flabel metal4 27194 4902 27220 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[23].CTOP
flabel psubdiff 27134 4600 27172 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[23].SUB
flabel metal4 27804 3456 27830 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[24].CBOT
flabel metal4 27686 2866 27712 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[24].CTOP
flabel psubdiff 27734 3122 27772 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[24].SUB
flabel metal4 27682 4312 27708 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[25].CBOT
flabel metal4 27800 4902 27826 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[25].CTOP
flabel psubdiff 27740 4600 27778 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[25].SUB
flabel metal4 28410 3456 28436 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[26].CBOT
flabel metal4 28292 2866 28318 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[26].CTOP
flabel psubdiff 28340 3122 28378 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[26].SUB
flabel metal4 28288 4312 28314 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[27].CBOT
flabel metal4 28406 4902 28432 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[27].CTOP
flabel psubdiff 28346 4600 28384 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[27].SUB
flabel metal4 29016 3456 29042 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[28].CBOT
flabel metal4 28898 2866 28924 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[28].CTOP
flabel psubdiff 28946 3122 28984 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[28].SUB
flabel metal4 28894 4312 28920 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[29].CBOT
flabel metal4 29012 4902 29038 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[29].CTOP
flabel psubdiff 28952 4600 28990 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[29].SUB
flabel metal4 29622 3456 29648 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[30].CBOT
flabel metal4 29504 2866 29530 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[30].CTOP
flabel psubdiff 29552 3122 29590 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[30].SUB
flabel metal4 29500 4312 29526 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[31].CBOT
flabel metal4 29618 4902 29644 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[31].CTOP
flabel psubdiff 29558 4600 29596 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[31].SUB
flabel metal4 30228 3456 30254 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[32].CBOT
flabel metal4 30110 2866 30136 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[32].CTOP
flabel psubdiff 30158 3122 30196 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[32].SUB
flabel metal4 30106 4312 30132 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[33].CBOT
flabel metal4 30224 4902 30250 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[33].CTOP
flabel psubdiff 30164 4600 30202 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[33].SUB
flabel metal4 30834 3456 30860 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[34].CBOT
flabel metal4 30716 2866 30742 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[34].CTOP
flabel psubdiff 30764 3122 30802 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[34].SUB
flabel metal4 30712 4312 30738 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[35].CBOT
flabel metal4 30830 4902 30856 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[35].CTOP
flabel psubdiff 30770 4600 30808 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[35].SUB
flabel metal4 31440 3456 31466 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[36].CBOT
flabel metal4 31322 2866 31348 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[36].CTOP
flabel psubdiff 31370 3122 31408 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[36].SUB
flabel metal4 31318 4312 31344 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[37].CBOT
flabel metal4 31436 4902 31462 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[37].CTOP
flabel psubdiff 31376 4600 31414 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[37].SUB
flabel metal4 32046 3456 32072 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[38].CBOT
flabel metal4 31928 2866 31954 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[38].CTOP
flabel psubdiff 31976 3122 32014 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[38].SUB
flabel metal4 31924 4312 31950 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[39].CBOT
flabel metal4 32042 4902 32068 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[39].CTOP
flabel psubdiff 31982 4600 32020 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[39].SUB
flabel metal4 32652 3456 32678 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[40].CBOT
flabel metal4 32534 2866 32560 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[40].CTOP
flabel psubdiff 32582 3122 32620 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[40].SUB
flabel metal4 32530 4312 32556 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[41].CBOT
flabel metal4 32648 4902 32674 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[41].CTOP
flabel psubdiff 32588 4600 32626 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[41].SUB
flabel metal4 33258 3456 33284 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[42].CBOT
flabel metal4 33140 2866 33166 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[42].CTOP
flabel psubdiff 33188 3122 33226 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[42].SUB
flabel metal4 33136 4312 33162 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[43].CBOT
flabel metal4 33254 4902 33280 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[43].CTOP
flabel psubdiff 33194 4600 33232 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[43].SUB
flabel metal4 33864 3456 33890 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[44].CBOT
flabel metal4 33746 2866 33772 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[44].CTOP
flabel psubdiff 33794 3122 33832 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[44].SUB
flabel metal4 33742 4312 33768 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[45].CBOT
flabel metal4 33860 4902 33886 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[45].CTOP
flabel psubdiff 33800 4600 33838 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[45].SUB
flabel metal4 34470 3456 34496 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[46].CBOT
flabel metal4 34352 2866 34378 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[46].CTOP
flabel psubdiff 34400 3122 34438 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[46].SUB
flabel metal4 34348 4312 34374 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[47].CBOT
flabel metal4 34466 4902 34492 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[47].CTOP
flabel psubdiff 34406 4600 34444 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[47].SUB
flabel metal4 35076 3456 35102 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[48].CBOT
flabel metal4 34958 2866 34984 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[48].CTOP
flabel psubdiff 35006 3122 35044 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[48].SUB
flabel metal4 34954 4312 34980 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[49].CBOT
flabel metal4 35072 4902 35098 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[49].CTOP
flabel psubdiff 35012 4600 35050 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[49].SUB
flabel metal4 35682 3456 35708 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[50].CBOT
flabel metal4 35564 2866 35590 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[50].CTOP
flabel psubdiff 35612 3122 35650 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[50].SUB
flabel metal4 35560 4312 35586 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[51].CBOT
flabel metal4 35678 4902 35704 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[51].CTOP
flabel psubdiff 35618 4600 35656 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[51].SUB
flabel metal4 36288 3456 36314 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[52].CBOT
flabel metal4 36170 2866 36196 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[52].CTOP
flabel psubdiff 36218 3122 36256 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[52].SUB
flabel metal4 36166 4312 36192 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[53].CBOT
flabel metal4 36284 4902 36310 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[53].CTOP
flabel psubdiff 36224 4600 36262 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[53].SUB
flabel metal4 36894 3456 36920 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[54].CBOT
flabel metal4 36776 2866 36802 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[54].CTOP
flabel psubdiff 36824 3122 36862 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[54].SUB
flabel metal4 36772 4312 36798 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[55].CBOT
flabel metal4 36890 4902 36916 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[55].CTOP
flabel psubdiff 36830 4600 36868 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[55].SUB
flabel metal4 37500 3456 37526 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[56].CBOT
flabel metal4 37382 2866 37408 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[56].CTOP
flabel psubdiff 37430 3122 37468 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[56].SUB
flabel metal4 37378 4312 37404 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[57].CBOT
flabel metal4 37496 4902 37522 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[57].CTOP
flabel psubdiff 37436 4600 37474 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[57].SUB
flabel metal4 38106 3456 38132 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[58].CBOT
flabel metal4 37988 2866 38014 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[58].CTOP
flabel psubdiff 38036 3122 38074 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[58].SUB
flabel metal4 37984 4312 38010 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[59].CBOT
flabel metal4 38102 4902 38128 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[59].CTOP
flabel psubdiff 38042 4600 38080 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[59].SUB
flabel metal4 38712 3456 38738 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[60].CBOT
flabel metal4 38594 2866 38620 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[60].CTOP
flabel psubdiff 38642 3122 38680 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[60].SUB
flabel metal4 38590 4312 38616 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[61].CBOT
flabel metal4 38708 4902 38734 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[61].CTOP
flabel psubdiff 38648 4600 38686 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[61].SUB
flabel metal4 39318 3456 39344 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[62].CBOT
flabel metal4 39200 2866 39226 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[62].CTOP
flabel psubdiff 39248 3122 39286 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[62].SUB
flabel metal4 39196 4312 39222 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[63].CBOT
flabel metal4 39314 4902 39340 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[63].CTOP
flabel psubdiff 39254 4600 39292 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_64_0.x1[63].SUB
flabel psubdiff 14766 3754 14810 3846 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.SUB
flabel metal4 14336 3550 14380 3642 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.CBOT
flabel metal4 14824 3554 14868 3646 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.CTOP
flabel metal4 14702 4074 14746 4166 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.CTOP
flabel metal4 19800 3456 19826 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[31].CBOT
flabel metal4 19682 2866 19708 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[31].CTOP
flabel psubdiff 19730 3122 19768 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[31].SUB
flabel metal4 19678 4312 19704 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[30].CBOT
flabel metal4 19796 4902 19822 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[30].CTOP
flabel psubdiff 19736 4600 19774 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[30].SUB
flabel metal4 19194 3456 19220 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[29].CBOT
flabel metal4 19076 2866 19102 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[29].CTOP
flabel psubdiff 19124 3122 19162 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[29].SUB
flabel metal4 19072 4312 19098 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[28].CBOT
flabel metal4 19190 4902 19216 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[28].CTOP
flabel psubdiff 19130 4600 19168 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[28].SUB
flabel metal4 18588 3456 18614 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[27].CBOT
flabel metal4 18470 2866 18496 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[27].CTOP
flabel psubdiff 18518 3122 18556 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[27].SUB
flabel metal4 18466 4312 18492 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[26].CBOT
flabel metal4 18584 4902 18610 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[26].CTOP
flabel psubdiff 18524 4600 18562 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[26].SUB
flabel metal4 17982 3456 18008 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[25].CBOT
flabel metal4 17864 2866 17890 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[25].CTOP
flabel psubdiff 17912 3122 17950 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[25].SUB
flabel metal4 17860 4312 17886 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[24].CBOT
flabel metal4 17978 4902 18004 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[24].CTOP
flabel psubdiff 17918 4600 17956 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[24].SUB
flabel metal4 17376 3456 17402 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[23].CBOT
flabel metal4 17258 2866 17284 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[23].CTOP
flabel psubdiff 17306 3122 17344 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[23].SUB
flabel metal4 17254 4312 17280 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[22].CBOT
flabel metal4 17372 4902 17398 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[22].CTOP
flabel psubdiff 17312 4600 17350 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[22].SUB
flabel metal4 16770 3456 16796 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[21].CBOT
flabel metal4 16652 2866 16678 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[21].CTOP
flabel psubdiff 16700 3122 16738 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[21].SUB
flabel metal4 16648 4312 16674 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[20].CBOT
flabel metal4 16766 4902 16792 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[20].CTOP
flabel psubdiff 16706 4600 16744 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[20].SUB
flabel metal4 16164 3456 16190 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[19].CBOT
flabel metal4 16046 2866 16072 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[19].CTOP
flabel psubdiff 16094 3122 16132 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[19].SUB
flabel metal4 16042 4312 16068 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[18].CBOT
flabel metal4 16160 4902 16186 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[18].CTOP
flabel psubdiff 16100 4600 16138 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[18].SUB
flabel metal4 15558 3456 15584 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[17].CBOT
flabel metal4 15440 2866 15466 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[17].CTOP
flabel psubdiff 15488 3122 15526 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[17].SUB
flabel metal4 15436 4312 15462 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[16].CBOT
flabel metal4 15554 4902 15580 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[16].CTOP
flabel psubdiff 15494 4600 15532 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[16].SUB
flabel metal4 14952 3456 14978 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[15].CBOT
flabel metal4 14834 2866 14860 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[15].CTOP
flabel psubdiff 14882 3122 14920 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[15].SUB
flabel metal4 14830 4312 14856 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[14].CBOT
flabel metal4 14948 4902 14974 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[14].CTOP
flabel psubdiff 14888 4600 14926 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[14].SUB
flabel metal4 14346 3456 14372 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[13].CBOT
flabel metal4 14228 2866 14254 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[13].CTOP
flabel psubdiff 14276 3122 14314 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[13].SUB
flabel metal4 14224 4312 14250 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[12].CBOT
flabel metal4 14342 4902 14368 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[12].CTOP
flabel psubdiff 14282 4600 14320 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[12].SUB
flabel metal4 13740 3456 13766 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[11].CBOT
flabel metal4 13622 2866 13648 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[11].CTOP
flabel psubdiff 13670 3122 13708 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[11].SUB
flabel metal4 13618 4312 13644 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[10].CBOT
flabel metal4 13736 4902 13762 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[10].CTOP
flabel psubdiff 13676 4600 13714 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[10].SUB
flabel metal4 13134 3456 13160 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[9].CBOT
flabel metal4 13016 2866 13042 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[9].CTOP
flabel psubdiff 13064 3122 13102 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[9].SUB
flabel metal4 13012 4312 13038 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[8].CBOT
flabel metal4 13130 4902 13156 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[8].CTOP
flabel psubdiff 13070 4600 13108 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[8].SUB
flabel metal4 12528 3456 12554 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[7].CBOT
flabel metal4 12410 2866 12436 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[7].CTOP
flabel psubdiff 12458 3122 12496 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[7].SUB
flabel metal4 12406 4312 12432 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[6].CBOT
flabel metal4 12524 4902 12550 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[6].CTOP
flabel psubdiff 12464 4600 12502 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[6].SUB
flabel metal4 11922 3456 11948 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[5].CBOT
flabel metal4 11804 2866 11830 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[5].CTOP
flabel psubdiff 11852 3122 11890 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[5].SUB
flabel metal4 11800 4312 11826 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[4].CBOT
flabel metal4 11918 4902 11944 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[4].CTOP
flabel psubdiff 11858 4600 11896 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[4].SUB
flabel metal4 11316 3456 11342 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[3].CBOT
flabel metal4 11198 2866 11224 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[3].CTOP
flabel psubdiff 11246 3122 11284 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[3].SUB
flabel metal4 11194 4312 11220 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[2].CBOT
flabel metal4 11312 4902 11338 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[2].CTOP
flabel psubdiff 11252 4600 11290 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[2].SUB
flabel metal4 10710 3456 10736 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[1].CBOT
flabel metal4 10592 2866 10618 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[1].CTOP
flabel psubdiff 10640 3122 10678 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[1].SUB
flabel metal4 10588 4312 10614 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[0].CBOT
flabel metal4 10706 4902 10732 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[0].CTOP
flabel psubdiff 10646 4600 10684 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_32_0.x1[0].SUB
flabel metal4 8156 3716 8192 3796 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.CBOT
flabel metal4 7432 3686 7468 3766 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.CTOP
flabel metal4 7546 4058 7590 4140 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.CTOP
flabel psubdiff 7850 3958 7894 4040 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.SUB
flabel metal4 9978 3456 10004 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[15].CBOT
flabel metal4 9860 2866 9886 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[15].CTOP
flabel psubdiff 9908 3122 9946 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[15].SUB
flabel metal4 9856 4312 9882 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[14].CBOT
flabel metal4 9974 4902 10000 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[14].CTOP
flabel psubdiff 9914 4600 9952 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[14].SUB
flabel metal4 9372 3456 9398 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[13].CBOT
flabel metal4 9254 2866 9280 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[13].CTOP
flabel psubdiff 9302 3122 9340 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[13].SUB
flabel metal4 9250 4312 9276 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[12].CBOT
flabel metal4 9368 4902 9394 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[12].CTOP
flabel psubdiff 9308 4600 9346 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[12].SUB
flabel metal4 8766 3456 8792 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[11].CBOT
flabel metal4 8648 2866 8674 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[11].CTOP
flabel psubdiff 8696 3122 8734 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[11].SUB
flabel metal4 8644 4312 8670 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[10].CBOT
flabel metal4 8762 4902 8788 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[10].CTOP
flabel psubdiff 8702 4600 8740 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[10].SUB
flabel metal4 8160 3456 8186 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[9].CBOT
flabel metal4 8042 2866 8068 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[9].CTOP
flabel psubdiff 8090 3122 8128 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[9].SUB
flabel metal4 8038 4312 8064 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[8].CBOT
flabel metal4 8156 4902 8182 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[8].CTOP
flabel psubdiff 8096 4600 8134 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[8].SUB
flabel metal4 7554 3456 7580 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[7].CBOT
flabel metal4 7436 2866 7462 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[7].CTOP
flabel psubdiff 7484 3122 7522 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[7].SUB
flabel metal4 7432 4312 7458 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[6].CBOT
flabel metal4 7550 4902 7576 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[6].CTOP
flabel psubdiff 7490 4600 7528 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[6].SUB
flabel metal4 6948 3456 6974 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[5].CBOT
flabel metal4 6830 2866 6856 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[5].CTOP
flabel psubdiff 6878 3122 6916 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[5].SUB
flabel metal4 6826 4312 6852 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[4].CBOT
flabel metal4 6944 4902 6970 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[4].CTOP
flabel psubdiff 6884 4600 6922 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[4].SUB
flabel metal4 6342 3456 6368 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[3].CBOT
flabel metal4 6224 2866 6250 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[3].CTOP
flabel psubdiff 6272 3122 6310 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[3].SUB
flabel metal4 6220 4312 6246 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[2].CBOT
flabel metal4 6338 4902 6364 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[2].CTOP
flabel psubdiff 6278 4600 6316 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[2].SUB
flabel metal4 5736 3456 5762 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[1].CBOT
flabel metal4 5618 2866 5644 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[1].CTOP
flabel psubdiff 5666 3122 5704 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[1].SUB
flabel metal4 5614 4312 5640 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[0].CBOT
flabel metal4 5732 4902 5758 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[0].CTOP
flabel psubdiff 5672 4600 5710 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_16_0.x1[0].SUB
flabel psubdiff 4207 3754 4251 3854 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.SUB
flabel metal4 4387 3586 4433 3678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.CBOT
flabel metal4 3659 3608 3705 3700 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.CTOP
flabel metal4 3787 4446 3827 4530 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.CTOP
flabel metal4 5003 3456 5029 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[7].CBOT
flabel metal4 4885 2866 4911 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[7].CTOP
flabel psubdiff 4933 3122 4971 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[7].SUB
flabel metal4 4881 4312 4907 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[6].CBOT
flabel metal4 4999 4902 5025 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[6].CTOP
flabel psubdiff 4939 4600 4977 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[6].SUB
flabel metal4 4397 3456 4423 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[5].CBOT
flabel metal4 4279 2866 4305 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[5].CTOP
flabel psubdiff 4327 3122 4365 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[5].SUB
flabel metal4 4275 4312 4301 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[4].CBOT
flabel metal4 4393 4902 4419 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[4].CTOP
flabel psubdiff 4333 4600 4371 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[4].SUB
flabel metal4 3791 3456 3817 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[3].CBOT
flabel metal4 3673 2866 3699 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[3].CTOP
flabel psubdiff 3721 3122 3759 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[3].SUB
flabel metal4 3669 4312 3695 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[2].CBOT
flabel metal4 3787 4902 3813 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[2].CTOP
flabel psubdiff 3727 4600 3765 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[2].SUB
flabel metal4 3185 3456 3211 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[1].CBOT
flabel metal4 3067 2866 3093 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[1].CTOP
flabel psubdiff 3115 3122 3153 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[1].SUB
flabel metal4 3063 4312 3089 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[0].CBOT
flabel metal4 3181 4902 3207 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[0].CTOP
flabel psubdiff 3121 4600 3159 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_8_0.x1[0].SUB
flabel metal4 2245 3814 2297 3854 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT
flabel metal4 1519 3698 1571 3738 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CTOP
flabel psubdiff 2069 3708 2109 3818 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.SUB
flabel metal4 1643 4036 1681 4118 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CTOP
flabel metal4 2257 3456 2283 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[3].CBOT
flabel metal4 2139 2866 2165 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[3].CTOP
flabel psubdiff 2187 3122 2225 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[3].SUB
flabel metal4 2135 4312 2161 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[2].CBOT
flabel metal4 2253 4902 2279 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[2].CTOP
flabel psubdiff 2193 4600 2231 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[2].SUB
flabel metal4 1651 3456 1677 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[1].CBOT
flabel metal4 1533 2866 1559 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[1].CTOP
flabel psubdiff 1581 3122 1619 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[1].SUB
flabel metal4 1529 4312 1555 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[0].CBOT
flabel metal4 1647 4902 1673 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[0].CTOP
flabel psubdiff 1587 4600 1625 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.x1[0].SUB
flabel psubdiff 669 3615 717 3729 0 FreeSans 160 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_2_0.SUB
flabel metal4 733 3610 769 3700 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_2_0.CBOT
flabel metal4 613 3168 649 3270 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_2_0.CTOP
flabel metal4 731 4752 771 4830 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_2_0.CTOP
flabel metal4 739 3456 765 3488 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_2_0.x2.CBOT
flabel metal4 621 2866 647 2898 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_2_0.x2.CTOP
flabel psubdiff 669 3122 707 3200 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_2_0.x2.SUB
flabel metal4 617 4312 643 4344 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_2_0.x1.CBOT
flabel metal4 735 4902 761 4934 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_2_0.x1.CTOP
flabel psubdiff 675 4600 713 4678 0 FreeSans 320 0 0 0 hgu_cdac_8bit_array_3.hgu_cdac_cap_2_0.x1.SUB
flabel metal4 -197 664 -171 696 0 FreeSans 320 0 0 0 hgu_cdac_unit_0.CBOT
flabel metal4 -79 1254 -53 1286 0 FreeSans 320 0 0 0 hgu_cdac_unit_0.CTOP
flabel psubdiff -139 952 -101 1030 0 FreeSans 320 0 0 0 hgu_cdac_unit_0.SUB
flabel metal4 -197 3152 -171 3184 0 FreeSans 320 0 0 0 hgu_cdac_unit_1.CBOT
flabel metal4 -79 3742 -53 3774 0 FreeSans 320 0 0 0 hgu_cdac_unit_1.CTOP
flabel psubdiff -139 3440 -101 3518 0 FreeSans 320 0 0 0 hgu_cdac_unit_1.SUB
flabel metal1 -318 5633 -291 5648 0 FreeSans 160 0 0 0 hgu_inverter_0.VREF
flabel metal1 -355 5694 -329 5722 0 FreeSans 160 0 0 0 hgu_inverter_0.VDD
flabel metal1 -357 5114 -333 5144 0 FreeSans 160 0 0 0 hgu_inverter_0.VSS
flabel metal1 875 5633 902 5648 0 FreeSans 160 0 0 0 inv_2_test_0/x2.VREF
flabel metal1 913 5694 939 5722 0 FreeSans 160 0 0 0 inv_2_test_0/x2.VDD
flabel metal1 917 5114 941 5144 0 FreeSans 160 0 0 0 inv_2_test_0/x2.VSS
flabel metal1 610 5633 637 5648 0 FreeSans 160 0 0 0 inv_2_test_0/x1.VREF
flabel metal1 573 5694 599 5722 0 FreeSans 160 0 0 0 inv_2_test_0/x1.VDD
flabel metal1 571 5114 595 5144 0 FreeSans 160 0 0 0 inv_2_test_0/x1.VSS
flabel metal1 2139 5633 2166 5648 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 2177 5694 2203 5722 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 2181 5114 2205 5144 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 1874 5633 1901 5648 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 1837 5694 1863 5722 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 1835 5114 1859 5144 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 2395 5633 2422 5648 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 2433 5694 2459 5722 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 2437 5114 2461 5144 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 2130 5633 2157 5648 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 2093 5694 2119 5722 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 2091 5114 2115 5144 0 FreeSans 160 0 0 0 inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 3758 5633 3785 5648 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 3796 5694 3822 5722 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 3800 5114 3824 5144 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 3493 5633 3520 5648 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 3456 5694 3482 5722 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 3454 5114 3478 5144 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 4014 5633 4041 5648 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 4052 5694 4078 5722 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 4056 5114 4080 5144 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 3749 5633 3776 5648 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 3712 5694 3738 5722 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 3710 5114 3734 5144 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 4270 5633 4297 5648 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 4308 5694 4334 5722 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 4312 5114 4336 5144 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 4005 5633 4032 5648 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 3968 5694 3994 5722 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 3966 5114 3990 5144 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 4526 5633 4553 5648 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 4564 5694 4590 5722 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 4568 5114 4592 5144 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 4261 5633 4288 5648 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 4224 5694 4250 5722 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 4222 5114 4246 5144 0 FreeSans 160 0 0 0 inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 8323 5633 8350 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 8361 5694 8387 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 8365 5114 8389 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 8058 5633 8085 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 8021 5694 8047 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 8019 5114 8043 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 8579 5633 8606 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 8617 5694 8643 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 8621 5114 8645 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 8314 5633 8341 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 8277 5694 8303 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 8275 5114 8299 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 8835 5633 8862 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 8873 5694 8899 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 8877 5114 8901 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 8570 5633 8597 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 8533 5694 8559 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 8531 5114 8555 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 9091 5633 9118 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 9129 5694 9155 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 9133 5114 9157 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 8826 5633 8853 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 8789 5694 8815 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 8787 5114 8811 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 9347 5633 9374 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 9385 5694 9411 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 9389 5114 9413 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 9082 5633 9109 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 9045 5694 9071 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 9043 5114 9067 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 9603 5633 9630 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 9641 5694 9667 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 9645 5114 9669 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 9338 5633 9365 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 9301 5694 9327 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 9299 5114 9323 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 9859 5633 9886 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 9897 5694 9923 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 9901 5114 9925 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 9594 5633 9621 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 9557 5694 9583 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 9555 5114 9579 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 10115 5633 10142 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 10153 5694 10179 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 10157 5114 10181 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 9850 5633 9877 5648 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 9813 5694 9839 5722 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 9811 5114 9835 5144 0 FreeSans 160 0 0 0 inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 15481 5633 15508 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 15519 5694 15545 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 15523 5114 15547 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 15216 5633 15243 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 15179 5694 15205 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 15177 5114 15201 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 15737 5633 15764 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 15775 5694 15801 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 15779 5114 15803 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 15472 5633 15499 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 15435 5694 15461 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 15433 5114 15457 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 15993 5633 16020 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 16031 5694 16057 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 16035 5114 16059 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 15728 5633 15755 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 15691 5694 15717 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 15689 5114 15713 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 16249 5633 16276 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 16287 5694 16313 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 16291 5114 16315 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 15984 5633 16011 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 15947 5694 15973 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 15945 5114 15969 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 16505 5633 16532 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 16543 5694 16569 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 16547 5114 16571 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 16240 5633 16267 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 16203 5694 16229 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 16201 5114 16225 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 16761 5633 16788 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 16799 5694 16825 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 16803 5114 16827 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 16496 5633 16523 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 16459 5694 16485 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 16457 5114 16481 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 17017 5633 17044 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 17055 5694 17081 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 17059 5114 17083 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 16752 5633 16779 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 16715 5694 16741 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 16713 5114 16737 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 17273 5633 17300 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 17311 5694 17337 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 17315 5114 17339 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 17008 5633 17035 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 16971 5694 16997 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 16969 5114 16993 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 17529 5633 17556 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 17567 5694 17593 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 17571 5114 17595 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 17264 5633 17291 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 17227 5694 17253 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 17225 5114 17249 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 17785 5633 17812 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 17823 5694 17849 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 17827 5114 17851 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 17520 5633 17547 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 17483 5694 17509 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 17481 5114 17505 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 18041 5633 18068 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 18079 5694 18105 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 18083 5114 18107 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 17776 5633 17803 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 17739 5694 17765 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 17737 5114 17761 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 18297 5633 18324 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 18335 5694 18361 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 18339 5114 18363 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 18032 5633 18059 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 17995 5694 18021 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 17993 5114 18017 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 18553 5633 18580 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 18591 5694 18617 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 18595 5114 18619 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 18288 5633 18315 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 18251 5694 18277 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 18249 5114 18273 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 18809 5633 18836 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 18847 5694 18873 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 18851 5114 18875 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 18544 5633 18571 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 18507 5694 18533 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 18505 5114 18529 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 19065 5633 19092 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 19103 5694 19129 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 19107 5114 19131 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 18800 5633 18827 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 18763 5694 18789 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 18761 5114 18785 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 19321 5633 19348 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 19359 5694 19385 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 19363 5114 19387 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 19056 5633 19083 5648 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 19019 5694 19045 5722 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 19017 5114 19041 5144 0 FreeSans 160 0 0 0 inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 24631 5633 24658 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 24669 5694 24695 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 24673 5114 24697 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 24366 5633 24393 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 24329 5694 24355 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 24327 5114 24351 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 24887 5633 24914 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 24925 5694 24951 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 24929 5114 24953 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 24622 5633 24649 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 24585 5694 24611 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 24583 5114 24607 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 25143 5633 25170 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 25181 5694 25207 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 25185 5114 25209 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 24878 5633 24905 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 24841 5694 24867 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 24839 5114 24863 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 25399 5633 25426 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 25437 5694 25463 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 25441 5114 25465 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 25134 5633 25161 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 25097 5694 25123 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 25095 5114 25119 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 25655 5633 25682 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 25693 5694 25719 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 25697 5114 25721 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 25390 5633 25417 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 25353 5694 25379 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 25351 5114 25375 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 25911 5633 25938 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 25949 5694 25975 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 25953 5114 25977 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 25646 5633 25673 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 25609 5694 25635 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 25607 5114 25631 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 26167 5633 26194 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 26205 5694 26231 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 26209 5114 26233 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 25902 5633 25929 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 25865 5694 25891 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 25863 5114 25887 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 26423 5633 26450 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 26461 5694 26487 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 26465 5114 26489 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 26158 5633 26185 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 26121 5694 26147 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 26119 5114 26143 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 26679 5633 26706 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 26717 5694 26743 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 26721 5114 26745 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 26414 5633 26441 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 26377 5694 26403 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 26375 5114 26399 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 26935 5633 26962 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 26973 5694 26999 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 26977 5114 27001 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 26670 5633 26697 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 26633 5694 26659 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 26631 5114 26655 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 27191 5633 27218 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 27229 5694 27255 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 27233 5114 27257 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 26926 5633 26953 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 26889 5694 26915 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 26887 5114 26911 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 27447 5633 27474 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 27485 5694 27511 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 27489 5114 27513 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 27182 5633 27209 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 27145 5694 27171 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 27143 5114 27167 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 27703 5633 27730 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 27741 5694 27767 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 27745 5114 27769 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 27438 5633 27465 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 27401 5694 27427 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 27399 5114 27423 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 27959 5633 27986 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 27997 5694 28023 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 28001 5114 28025 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 27694 5633 27721 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 27657 5694 27683 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 27655 5114 27679 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 28215 5633 28242 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 28253 5694 28279 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 28257 5114 28281 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 27950 5633 27977 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 27913 5694 27939 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 27911 5114 27935 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 28471 5633 28498 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 28509 5694 28535 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 28513 5114 28537 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 28206 5633 28233 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 28169 5694 28195 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 28167 5114 28191 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 20535 5633 20562 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 20573 5694 20599 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 20577 5114 20601 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 20270 5633 20297 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 20233 5694 20259 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 20231 5114 20255 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 20791 5633 20818 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 20829 5694 20855 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 20833 5114 20857 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 20526 5633 20553 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 20489 5694 20515 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 20487 5114 20511 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 21047 5633 21074 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 21085 5694 21111 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 21089 5114 21113 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 20782 5633 20809 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 20745 5694 20771 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 20743 5114 20767 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 21303 5633 21330 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 21341 5694 21367 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 21345 5114 21369 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 21038 5633 21065 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 21001 5694 21027 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 20999 5114 21023 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 21559 5633 21586 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 21597 5694 21623 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 21601 5114 21625 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 21294 5633 21321 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 21257 5694 21283 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 21255 5114 21279 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 21815 5633 21842 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 21853 5694 21879 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 21857 5114 21881 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 21550 5633 21577 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 21513 5694 21539 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 21511 5114 21535 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 22071 5633 22098 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 22109 5694 22135 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 22113 5114 22137 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 21806 5633 21833 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 21769 5694 21795 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 21767 5114 21791 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 22327 5633 22354 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 22365 5694 22391 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 22369 5114 22393 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 22062 5633 22089 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 22025 5694 22051 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 22023 5114 22047 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 22583 5633 22610 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 22621 5694 22647 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 22625 5114 22649 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 22318 5633 22345 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 22281 5694 22307 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 22279 5114 22303 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 22839 5633 22866 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 22877 5694 22903 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 22881 5114 22905 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 22574 5633 22601 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 22537 5694 22563 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 22535 5114 22559 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 23095 5633 23122 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 23133 5694 23159 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 23137 5114 23161 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 22830 5633 22857 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 22793 5694 22819 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 22791 5114 22815 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 23351 5633 23378 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 23389 5694 23415 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 23393 5114 23417 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 23086 5633 23113 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 23049 5694 23075 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 23047 5114 23071 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 23607 5633 23634 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 23645 5694 23671 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 23649 5114 23673 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 23342 5633 23369 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 23305 5694 23331 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 23303 5114 23327 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 23863 5633 23890 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 23901 5694 23927 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 23905 5114 23929 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 23598 5633 23625 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 23561 5694 23587 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 23559 5114 23583 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 24119 5633 24146 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 24157 5694 24183 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 24161 5114 24185 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 23854 5633 23881 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 23817 5694 23843 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 23815 5114 23839 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 24375 5633 24402 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 24413 5694 24439 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 24417 5114 24441 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 24110 5633 24137 5648 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 24073 5694 24099 5722 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 24071 5114 24095 5144 0 FreeSans 160 0 0 0 inv_64_test_0/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 -296 6321 -269 6336 0 FreeSans 160 0 0 0 hgu_inverter_1.VREF
flabel metal1 -333 6382 -307 6410 0 FreeSans 160 0 0 0 hgu_inverter_1.VDD
flabel metal1 -335 5802 -311 5832 0 FreeSans 160 0 0 0 hgu_inverter_1.VSS
flabel metal1 746 6321 773 6336 0 FreeSans 160 0 0 0 inv_2_test_1/x2.VREF
flabel metal1 784 6382 810 6410 0 FreeSans 160 0 0 0 inv_2_test_1/x2.VDD
flabel metal1 788 5802 812 5832 0 FreeSans 160 0 0 0 inv_2_test_1/x2.VSS
flabel metal1 481 6321 508 6336 0 FreeSans 160 0 0 0 inv_2_test_1/x1.VREF
flabel metal1 444 6382 470 6410 0 FreeSans 160 0 0 0 inv_2_test_1/x1.VDD
flabel metal1 442 5802 466 5832 0 FreeSans 160 0 0 0 inv_2_test_1/x1.VSS
flabel metal1 1655 6321 1682 6336 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_1/x2.VREF
flabel metal1 1693 6382 1719 6410 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_1/x2.VDD
flabel metal1 1697 5802 1721 5832 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_1/x2.VSS
flabel metal1 1390 6321 1417 6336 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_1/x1.VREF
flabel metal1 1353 6382 1379 6410 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_1/x1.VDD
flabel metal1 1351 5802 1375 5832 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_1/x1.VSS
flabel metal1 1911 6321 1938 6336 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_0/x2.VREF
flabel metal1 1949 6382 1975 6410 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_0/x2.VDD
flabel metal1 1953 5802 1977 5832 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_0/x2.VSS
flabel metal1 1646 6321 1673 6336 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_0/x1.VREF
flabel metal1 1609 6382 1635 6410 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_0/x1.VDD
flabel metal1 1607 5802 1631 5832 0 FreeSans 160 0 0 0 inv_4_test_2/inv_2_test_0/x1.VSS
flabel metal1 3188 6321 3215 6336 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 3226 6382 3252 6410 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 3230 5802 3254 5832 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 2923 6321 2950 6336 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 2886 6382 2912 6410 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 2884 5802 2908 5832 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 3444 6321 3471 6336 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 3482 6382 3508 6410 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 3486 5802 3510 5832 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 3179 6321 3206 6336 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 3142 6382 3168 6410 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 3140 5802 3164 5832 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 3700 6321 3727 6336 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 3738 6382 3764 6410 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 3742 5802 3766 5832 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 3435 6321 3462 6336 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 3398 6382 3424 6410 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 3396 5802 3420 5832 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 3956 6321 3983 6336 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 3994 6382 4020 6410 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 3998 5802 4022 5832 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 3691 6321 3718 6336 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 3654 6382 3680 6410 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 3652 5802 3676 5832 0 FreeSans 160 0 0 0 inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 5739 6321 5766 6336 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 5777 6382 5803 6410 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 5781 5802 5805 5832 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 5474 6321 5501 6336 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 5437 6382 5463 6410 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 5435 5802 5459 5832 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 5995 6321 6022 6336 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 6033 6382 6059 6410 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 6037 5802 6061 5832 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 5730 6321 5757 6336 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 5693 6382 5719 6410 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 5691 5802 5715 5832 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 6251 6321 6278 6336 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 6289 6382 6315 6410 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 6293 5802 6317 5832 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 5986 6321 6013 6336 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 5949 6382 5975 6410 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 5947 5802 5971 5832 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 6507 6321 6534 6336 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 6545 6382 6571 6410 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 6549 5802 6573 5832 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 6242 6321 6269 6336 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 6205 6382 6231 6410 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 6203 5802 6227 5832 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 6763 6321 6790 6336 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 6801 6382 6827 6410 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 6805 5802 6829 5832 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 6498 6321 6525 6336 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 6461 6382 6487 6410 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 6459 5802 6483 5832 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 7019 6321 7046 6336 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 7057 6382 7083 6410 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 7061 5802 7085 5832 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 6754 6321 6781 6336 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 6717 6382 6743 6410 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 6715 5802 6739 5832 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 7275 6321 7302 6336 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 7313 6382 7339 6410 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 7317 5802 7341 5832 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 7010 6321 7037 6336 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 6973 6382 6999 6410 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 6971 5802 6995 5832 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 7531 6321 7558 6336 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 7569 6382 7595 6410 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 7573 5802 7597 5832 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 7266 6321 7293 6336 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 7229 6382 7255 6410 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 7227 5802 7251 5832 0 FreeSans 160 0 0 0 inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 10826 6321 10853 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 10864 6382 10890 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 10868 5802 10892 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 10561 6321 10588 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 10524 6382 10550 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 10522 5802 10546 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 11082 6321 11109 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 11120 6382 11146 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 11124 5802 11148 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 10817 6321 10844 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 10780 6382 10806 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 10778 5802 10802 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 11338 6321 11365 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 11376 6382 11402 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 11380 5802 11404 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 11073 6321 11100 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 11036 6382 11062 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 11034 5802 11058 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 11594 6321 11621 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 11632 6382 11658 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 11636 5802 11660 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 11329 6321 11356 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 11292 6382 11318 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 11290 5802 11314 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 11850 6321 11877 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 11888 6382 11914 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 11892 5802 11916 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 11585 6321 11612 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 11548 6382 11574 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 11546 5802 11570 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 12106 6321 12133 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 12144 6382 12170 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 12148 5802 12172 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 11841 6321 11868 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 11804 6382 11830 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 11802 5802 11826 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 12362 6321 12389 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 12400 6382 12426 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 12404 5802 12428 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 12097 6321 12124 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 12060 6382 12086 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 12058 5802 12082 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 12618 6321 12645 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 12656 6382 12682 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 12660 5802 12684 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 12353 6321 12380 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 12316 6382 12342 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 12314 5802 12338 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 12874 6321 12901 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 12912 6382 12938 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 12916 5802 12940 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 12609 6321 12636 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 12572 6382 12598 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 12570 5802 12594 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 13130 6321 13157 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 13168 6382 13194 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 13172 5802 13196 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 12865 6321 12892 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 12828 6382 12854 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 12826 5802 12850 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 13386 6321 13413 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 13424 6382 13450 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 13428 5802 13452 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 13121 6321 13148 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 13084 6382 13110 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 13082 5802 13106 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 13642 6321 13669 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 13680 6382 13706 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 13684 5802 13708 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 13377 6321 13404 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 13340 6382 13366 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 13338 5802 13362 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 13898 6321 13925 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 13936 6382 13962 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 13940 5802 13964 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 13633 6321 13660 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 13596 6382 13622 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 13594 5802 13618 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 14154 6321 14181 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 14192 6382 14218 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 14196 5802 14220 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 13889 6321 13916 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 13852 6382 13878 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 13850 5802 13874 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 14410 6321 14437 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 14448 6382 14474 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 14452 5802 14476 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 14145 6321 14172 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 14108 6382 14134 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 14106 5802 14130 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 14666 6321 14693 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 14704 6382 14730 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 14708 5802 14732 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 14401 6321 14428 6336 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 14364 6382 14390 6410 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 14362 5802 14386 5832 0 FreeSans 160 0 0 0 inv_32_test_0/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 24707 6321 24734 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 24745 6382 24771 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 24749 5802 24773 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 24442 6321 24469 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 24405 6382 24431 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 24403 5802 24427 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 24963 6321 24990 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 25001 6382 25027 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 25005 5802 25029 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 24698 6321 24725 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 24661 6382 24687 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 24659 5802 24683 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 25219 6321 25246 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 25257 6382 25283 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 25261 5802 25285 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 24954 6321 24981 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 24917 6382 24943 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 24915 5802 24939 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 25475 6321 25502 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 25513 6382 25539 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 25517 5802 25541 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 25210 6321 25237 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 25173 6382 25199 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 25171 5802 25195 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 25731 6321 25758 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 25769 6382 25795 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 25773 5802 25797 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 25466 6321 25493 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 25429 6382 25455 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 25427 5802 25451 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 25987 6321 26014 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 26025 6382 26051 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 26029 5802 26053 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 25722 6321 25749 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 25685 6382 25711 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 25683 5802 25707 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 26243 6321 26270 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 26281 6382 26307 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 26285 5802 26309 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 25978 6321 26005 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 25941 6382 25967 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 25939 5802 25963 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 26499 6321 26526 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 26537 6382 26563 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 26541 5802 26565 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 26234 6321 26261 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 26197 6382 26223 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 26195 5802 26219 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 26755 6321 26782 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 26793 6382 26819 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 26797 5802 26821 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 26490 6321 26517 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 26453 6382 26479 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 26451 5802 26475 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 27011 6321 27038 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 27049 6382 27075 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 27053 5802 27077 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 26746 6321 26773 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 26709 6382 26735 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 26707 5802 26731 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 27267 6321 27294 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 27305 6382 27331 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 27309 5802 27333 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 27002 6321 27029 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 26965 6382 26991 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 26963 5802 26987 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 27523 6321 27550 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 27561 6382 27587 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 27565 5802 27589 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 27258 6321 27285 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 27221 6382 27247 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 27219 5802 27243 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 27779 6321 27806 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 27817 6382 27843 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 27821 5802 27845 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 27514 6321 27541 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 27477 6382 27503 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 27475 5802 27499 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 28035 6321 28062 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 28073 6382 28099 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 28077 5802 28101 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 27770 6321 27797 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 27733 6382 27759 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 27731 5802 27755 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 28291 6321 28318 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 28329 6382 28355 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 28333 5802 28357 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 28026 6321 28053 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 27989 6382 28015 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 27987 5802 28011 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 28547 6321 28574 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 28585 6382 28611 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 28589 5802 28613 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 28282 6321 28309 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 28245 6382 28271 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 28243 5802 28267 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_2/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 20611 6321 20638 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 20649 6382 20675 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 20653 5802 20677 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 20346 6321 20373 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 20309 6382 20335 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 20307 5802 20331 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 20867 6321 20894 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 20905 6382 20931 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 20909 5802 20933 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 20602 6321 20629 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 20565 6382 20591 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 20563 5802 20587 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 21123 6321 21150 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 21161 6382 21187 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 21165 5802 21189 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 20858 6321 20885 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 20821 6382 20847 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 20819 5802 20843 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 21379 6321 21406 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 21417 6382 21443 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 21421 5802 21445 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 21114 6321 21141 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 21077 6382 21103 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 21075 5802 21099 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 21635 6321 21662 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 21673 6382 21699 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 21677 5802 21701 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 21370 6321 21397 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 21333 6382 21359 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 21331 5802 21355 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 21891 6321 21918 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 21929 6382 21955 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 21933 5802 21957 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 21626 6321 21653 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 21589 6382 21615 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 21587 5802 21611 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 22147 6321 22174 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 22185 6382 22211 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 22189 5802 22213 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 21882 6321 21909 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 21845 6382 21871 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 21843 5802 21867 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 22403 6321 22430 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 22441 6382 22467 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 22445 5802 22469 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 22138 6321 22165 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 22101 6382 22127 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 22099 5802 22123 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_1/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 22659 6321 22686 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 22697 6382 22723 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 22701 5802 22725 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 22394 6321 22421 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 22357 6382 22383 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 22355 5802 22379 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 22915 6321 22942 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 22953 6382 22979 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 22957 5802 22981 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 22650 6321 22677 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 22613 6382 22639 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 22611 5802 22635 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 23171 6321 23198 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 23209 6382 23235 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 23213 5802 23237 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 22906 6321 22933 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 22869 6382 22895 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 22867 5802 22891 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 23427 6321 23454 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 23465 6382 23491 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 23469 5802 23493 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 23162 6321 23189 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 23125 6382 23151 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 23123 5802 23147 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_1/inv_4_test_0/inv_2_test_0/x1.VSS
flabel metal1 23683 6321 23710 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VREF
flabel metal1 23721 6382 23747 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VDD
flabel metal1 23725 5802 23749 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x2.VSS
flabel metal1 23418 6321 23445 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VREF
flabel metal1 23381 6382 23407 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VDD
flabel metal1 23379 5802 23403 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_1/x1.VSS
flabel metal1 23939 6321 23966 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VREF
flabel metal1 23977 6382 24003 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VDD
flabel metal1 23981 5802 24005 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x2.VSS
flabel metal1 23674 6321 23701 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VREF
flabel metal1 23637 6382 23663 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VDD
flabel metal1 23635 5802 23659 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_1/inv_2_test_0/x1.VSS
flabel metal1 24195 6321 24222 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VREF
flabel metal1 24233 6382 24259 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VDD
flabel metal1 24237 5802 24261 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x2.VSS
flabel metal1 23930 6321 23957 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VREF
flabel metal1 23893 6382 23919 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VDD
flabel metal1 23891 5802 23915 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_1/x1.VSS
flabel metal1 24451 6321 24478 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VREF
flabel metal1 24489 6382 24515 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VDD
flabel metal1 24493 5802 24517 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x2.VSS
flabel metal1 24186 6321 24213 6336 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VREF
flabel metal1 24149 6382 24175 6410 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VDD
flabel metal1 24147 5802 24171 5832 0 FreeSans 160 0 0 0 inv_64_test_1/inv_32_test_1/inv_16_test_0/inv_8_test_0/inv_4_test_0/inv_2_test_0/x1.VSS
<< end >>
