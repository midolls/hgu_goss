magic
tech sky130A
magscale 1 2
timestamp 1701237156
<< nwell >>
rect 991 5890 4184 6250
rect 992 5888 4176 5890
rect 984 5014 13040 5375
rect 544 4321 13040 4686
rect 589 3773 1492 3822
rect 588 3452 1492 3773
rect 3130 3457 13034 3821
rect 3130 3453 13031 3457
rect 996 2901 13031 2940
rect 995 2580 13031 2901
<< pwell >>
rect 993 5576 4167 5849
rect 1030 4706 12994 4978
rect 597 4242 12994 4282
rect 595 4086 12994 4242
rect 597 4016 12994 4086
rect 627 3212 901 3368
rect 903 3212 1425 3394
rect 657 3174 691 3212
rect 932 3174 966 3212
rect 3210 3209 12993 3404
rect 3197 3175 12993 3209
rect 3210 3144 12993 3175
rect 1034 2271 12993 2555
<< scnmos >>
rect 1114 5674 1144 5778
rect 1202 5674 1232 5778
rect 1390 5674 1420 5804
rect 1474 5674 1504 5804
rect 1558 5674 1588 5804
rect 1642 5674 1672 5804
rect 1726 5674 1756 5804
rect 2389 5674 2419 5804
rect 2473 5674 2503 5804
rect 2573 5674 2603 5804
rect 2657 5674 2687 5804
rect 2758 5674 2788 5758
rect 2853 5674 2883 5746
rect 2963 5674 2993 5746
rect 3070 5674 3100 5758
rect 3258 5674 3288 5758
rect 3343 5674 3373 5758
rect 3533 5674 3563 5758
rect 3641 5674 3671 5758
rect 3737 5674 3767 5746
rect 3847 5674 3877 5746
rect 3942 5674 3972 5758
rect 4026 5674 4056 5758
rect 1113 4801 1143 4885
rect 1197 4801 1227 4885
rect 1385 4801 1415 4885
rect 1480 4801 1510 4873
rect 1586 4801 1616 4873
rect 1682 4801 1712 4885
rect 1792 4801 1822 4885
rect 1892 4801 1922 4929
rect 1976 4801 2006 4929
rect 2164 4801 2194 4929
rect 2259 4801 2289 4873
rect 2368 4801 2398 4873
rect 2463 4801 2493 4885
rect 2549 4801 2579 4885
rect 2667 4801 2697 4929
rect 2751 4801 2781 4929
rect 2939 4801 2969 4885
rect 3034 4801 3064 4931
rect 3222 4801 3252 4885
rect 3317 4801 3347 4931
rect 3505 4801 3535 4885
rect 3589 4801 3619 4885
rect 3777 4801 3807 4885
rect 3872 4801 3902 4873
rect 3978 4801 4008 4873
rect 4074 4801 4104 4885
rect 4184 4801 4214 4885
rect 4284 4801 4314 4929
rect 4368 4801 4398 4929
rect 4556 4801 4586 4929
rect 4651 4801 4681 4873
rect 4760 4801 4790 4873
rect 4855 4801 4885 4885
rect 4941 4801 4971 4885
rect 5059 4801 5089 4929
rect 5143 4801 5173 4929
rect 5331 4801 5361 4885
rect 5426 4801 5456 4931
rect 5614 4801 5644 4885
rect 5709 4801 5739 4931
rect 5897 4801 5927 4885
rect 5981 4801 6011 4885
rect 6169 4801 6199 4885
rect 6264 4801 6294 4873
rect 6370 4801 6400 4873
rect 6466 4801 6496 4885
rect 6576 4801 6606 4885
rect 6676 4801 6706 4929
rect 6760 4801 6790 4929
rect 6948 4801 6978 4929
rect 7043 4801 7073 4873
rect 7152 4801 7182 4873
rect 7247 4801 7277 4885
rect 7333 4801 7363 4885
rect 7451 4801 7481 4929
rect 7535 4801 7565 4929
rect 7723 4801 7753 4885
rect 7818 4801 7848 4931
rect 8006 4801 8036 4885
rect 8101 4801 8131 4931
rect 8289 4801 8319 4885
rect 8373 4801 8403 4885
rect 8561 4801 8591 4885
rect 8656 4801 8686 4873
rect 8762 4801 8792 4873
rect 8858 4801 8888 4885
rect 8968 4801 8998 4885
rect 9068 4801 9098 4929
rect 9152 4801 9182 4929
rect 9340 4801 9370 4929
rect 9435 4801 9465 4873
rect 9544 4801 9574 4873
rect 9639 4801 9669 4885
rect 9725 4801 9755 4885
rect 9843 4801 9873 4929
rect 9927 4801 9957 4929
rect 10115 4801 10145 4885
rect 10210 4801 10240 4931
rect 10398 4801 10428 4885
rect 10493 4801 10523 4931
rect 10681 4801 10711 4885
rect 10765 4801 10795 4885
rect 10953 4801 10983 4885
rect 11048 4801 11078 4873
rect 11154 4801 11184 4873
rect 11250 4801 11280 4885
rect 11360 4801 11390 4885
rect 11460 4801 11490 4929
rect 11544 4801 11574 4929
rect 11732 4801 11762 4929
rect 11827 4801 11857 4873
rect 11936 4801 11966 4873
rect 12031 4801 12061 4885
rect 12117 4801 12147 4885
rect 12235 4801 12265 4929
rect 12319 4801 12349 4929
rect 12507 4801 12537 4885
rect 12602 4801 12632 4931
rect 12790 4801 12820 4885
rect 12885 4801 12915 4931
rect 673 4112 703 4216
rect 761 4112 791 4216
rect 949 4112 979 4242
rect 1033 4112 1063 4242
rect 1117 4112 1147 4242
rect 1201 4112 1231 4242
rect 1285 4112 1315 4242
rect 1481 4112 1511 4242
rect 1565 4112 1595 4242
rect 1649 4112 1679 4242
rect 1733 4112 1763 4242
rect 1817 4112 1847 4242
rect 1901 4112 1931 4242
rect 1985 4112 2015 4242
rect 2069 4112 2099 4242
rect 2153 4112 2183 4242
rect 2237 4112 2267 4242
rect 2321 4112 2351 4242
rect 2405 4112 2435 4242
rect 2489 4112 2519 4242
rect 2573 4112 2603 4242
rect 2657 4112 2687 4242
rect 2741 4112 2771 4242
rect 2825 4112 2855 4242
rect 2909 4112 2939 4242
rect 2993 4112 3023 4242
rect 3077 4112 3107 4242
rect 3161 4112 3191 4242
rect 3245 4112 3275 4242
rect 3505 4112 3535 4242
rect 3600 4112 3630 4196
rect 3788 4112 3818 4242
rect 3883 4112 3913 4196
rect 4071 4112 4101 4240
rect 4155 4112 4185 4240
rect 4273 4112 4303 4196
rect 4359 4112 4389 4196
rect 4454 4112 4484 4184
rect 4563 4112 4593 4184
rect 4658 4112 4688 4240
rect 4846 4112 4876 4240
rect 4930 4112 4960 4240
rect 5030 4112 5060 4196
rect 5140 4112 5170 4196
rect 5236 4112 5266 4184
rect 5342 4112 5372 4184
rect 5437 4112 5467 4196
rect 5625 4112 5655 4196
rect 5709 4112 5739 4196
rect 5897 4112 5927 4242
rect 5992 4112 6022 4196
rect 6180 4112 6210 4242
rect 6275 4112 6305 4196
rect 6463 4112 6493 4240
rect 6547 4112 6577 4240
rect 6665 4112 6695 4196
rect 6751 4112 6781 4196
rect 6846 4112 6876 4184
rect 6955 4112 6985 4184
rect 7050 4112 7080 4240
rect 7238 4112 7268 4240
rect 7322 4112 7352 4240
rect 7422 4112 7452 4196
rect 7532 4112 7562 4196
rect 7628 4112 7658 4184
rect 7734 4112 7764 4184
rect 7829 4112 7859 4196
rect 8017 4112 8047 4196
rect 8101 4112 8131 4196
rect 8289 4112 8319 4242
rect 8384 4112 8414 4196
rect 8572 4112 8602 4242
rect 8667 4112 8697 4196
rect 8855 4112 8885 4240
rect 8939 4112 8969 4240
rect 9057 4112 9087 4196
rect 9143 4112 9173 4196
rect 9238 4112 9268 4184
rect 9347 4112 9377 4184
rect 9442 4112 9472 4240
rect 9630 4112 9660 4240
rect 9714 4112 9744 4240
rect 9814 4112 9844 4196
rect 9924 4112 9954 4196
rect 10020 4112 10050 4184
rect 10126 4112 10156 4184
rect 10221 4112 10251 4196
rect 10409 4112 10439 4196
rect 10493 4112 10523 4196
rect 10681 4112 10711 4242
rect 10776 4112 10806 4196
rect 10964 4112 10994 4242
rect 11059 4112 11089 4196
rect 11247 4112 11277 4240
rect 11331 4112 11361 4240
rect 11449 4112 11479 4196
rect 11535 4112 11565 4196
rect 11630 4112 11660 4184
rect 11739 4112 11769 4184
rect 11834 4112 11864 4240
rect 12022 4112 12052 4240
rect 12106 4112 12136 4240
rect 12206 4112 12236 4196
rect 12316 4112 12346 4196
rect 12412 4112 12442 4184
rect 12518 4112 12548 4184
rect 12613 4112 12643 4196
rect 12801 4112 12831 4196
rect 12885 4112 12915 4196
rect 705 3238 735 3342
rect 793 3238 823 3342
rect 981 3238 1011 3368
rect 1065 3238 1095 3368
rect 1149 3238 1179 3368
rect 1233 3238 1263 3368
rect 1317 3238 1347 3368
rect 3288 3239 3318 3369
rect 3504 3239 3534 3323
rect 3588 3239 3618 3323
rect 3776 3239 3806 3323
rect 3871 3239 3901 3311
rect 3977 3239 4007 3311
rect 4073 3239 4103 3323
rect 4183 3239 4213 3323
rect 4283 3239 4313 3367
rect 4367 3239 4397 3367
rect 4555 3239 4585 3367
rect 4650 3239 4680 3311
rect 4759 3239 4789 3311
rect 4854 3239 4884 3323
rect 4940 3239 4970 3323
rect 5058 3239 5088 3367
rect 5142 3239 5172 3367
rect 5330 3239 5360 3323
rect 5425 3239 5455 3369
rect 5613 3239 5643 3323
rect 5708 3239 5738 3369
rect 5896 3239 5926 3323
rect 5980 3239 6010 3323
rect 6168 3239 6198 3323
rect 6263 3239 6293 3311
rect 6369 3239 6399 3311
rect 6465 3239 6495 3323
rect 6575 3239 6605 3323
rect 6675 3239 6705 3367
rect 6759 3239 6789 3367
rect 6947 3239 6977 3367
rect 7042 3239 7072 3311
rect 7151 3239 7181 3311
rect 7246 3239 7276 3323
rect 7332 3239 7362 3323
rect 7450 3239 7480 3367
rect 7534 3239 7564 3367
rect 7722 3239 7752 3323
rect 7817 3239 7847 3369
rect 8005 3239 8035 3323
rect 8100 3239 8130 3369
rect 8288 3239 8318 3323
rect 8372 3239 8402 3323
rect 8560 3239 8590 3323
rect 8655 3239 8685 3311
rect 8761 3239 8791 3311
rect 8857 3239 8887 3323
rect 8967 3239 8997 3323
rect 9067 3239 9097 3367
rect 9151 3239 9181 3367
rect 9339 3239 9369 3367
rect 9434 3239 9464 3311
rect 9543 3239 9573 3311
rect 9638 3239 9668 3323
rect 9724 3239 9754 3323
rect 9842 3239 9872 3367
rect 9926 3239 9956 3367
rect 10114 3239 10144 3323
rect 10209 3239 10239 3369
rect 10397 3239 10427 3323
rect 10492 3239 10522 3369
rect 10680 3239 10710 3323
rect 10764 3239 10794 3323
rect 10952 3239 10982 3323
rect 11047 3239 11077 3311
rect 11153 3239 11183 3311
rect 11249 3239 11279 3323
rect 11359 3239 11389 3323
rect 11459 3239 11489 3367
rect 11543 3239 11573 3367
rect 11731 3239 11761 3367
rect 11826 3239 11856 3311
rect 11935 3239 11965 3311
rect 12030 3239 12060 3323
rect 12116 3239 12146 3323
rect 12234 3239 12264 3367
rect 12318 3239 12348 3367
rect 12506 3239 12536 3323
rect 12601 3239 12631 3369
rect 12789 3239 12819 3323
rect 12884 3239 12914 3369
rect 1112 2366 1142 2496
rect 1207 2366 1237 2450
rect 1395 2366 1425 2496
rect 1490 2366 1520 2450
rect 1678 2366 1708 2494
rect 1762 2366 1792 2494
rect 1880 2366 1910 2450
rect 1966 2366 1996 2450
rect 2061 2366 2091 2438
rect 2170 2366 2200 2438
rect 2265 2366 2295 2494
rect 2453 2366 2483 2494
rect 2537 2366 2567 2494
rect 2637 2366 2667 2450
rect 2747 2366 2777 2450
rect 2843 2366 2873 2438
rect 2949 2366 2979 2438
rect 3044 2366 3074 2450
rect 3232 2366 3262 2450
rect 3316 2366 3346 2450
rect 3504 2366 3534 2496
rect 3599 2366 3629 2450
rect 3787 2366 3817 2496
rect 3882 2366 3912 2450
rect 4070 2366 4100 2494
rect 4154 2366 4184 2494
rect 4272 2366 4302 2450
rect 4358 2366 4388 2450
rect 4453 2366 4483 2438
rect 4562 2366 4592 2438
rect 4657 2366 4687 2494
rect 4845 2366 4875 2494
rect 4929 2366 4959 2494
rect 5029 2366 5059 2450
rect 5139 2366 5169 2450
rect 5235 2366 5265 2438
rect 5341 2366 5371 2438
rect 5436 2366 5466 2450
rect 5624 2366 5654 2450
rect 5708 2366 5738 2450
rect 5896 2366 5926 2496
rect 5991 2366 6021 2450
rect 6179 2366 6209 2496
rect 6274 2366 6304 2450
rect 6462 2366 6492 2494
rect 6546 2366 6576 2494
rect 6664 2366 6694 2450
rect 6750 2366 6780 2450
rect 6845 2366 6875 2438
rect 6954 2366 6984 2438
rect 7049 2366 7079 2494
rect 7237 2366 7267 2494
rect 7321 2366 7351 2494
rect 7421 2366 7451 2450
rect 7531 2366 7561 2450
rect 7627 2366 7657 2438
rect 7733 2366 7763 2438
rect 7828 2366 7858 2450
rect 8016 2366 8046 2450
rect 8100 2366 8130 2450
rect 8288 2366 8318 2496
rect 8383 2366 8413 2450
rect 8571 2366 8601 2496
rect 8666 2366 8696 2450
rect 8854 2366 8884 2494
rect 8938 2366 8968 2494
rect 9056 2366 9086 2450
rect 9142 2366 9172 2450
rect 9237 2366 9267 2438
rect 9346 2366 9376 2438
rect 9441 2366 9471 2494
rect 9629 2366 9659 2494
rect 9713 2366 9743 2494
rect 9813 2366 9843 2450
rect 9923 2366 9953 2450
rect 10019 2366 10049 2438
rect 10125 2366 10155 2438
rect 10220 2366 10250 2450
rect 10408 2366 10438 2450
rect 10492 2366 10522 2450
rect 10680 2366 10710 2496
rect 10775 2366 10805 2450
rect 10963 2366 10993 2496
rect 11058 2366 11088 2450
rect 11246 2366 11276 2494
rect 11330 2366 11360 2494
rect 11448 2366 11478 2450
rect 11534 2366 11564 2450
rect 11629 2366 11659 2438
rect 11738 2366 11768 2438
rect 11833 2366 11863 2494
rect 12021 2366 12051 2494
rect 12105 2366 12135 2494
rect 12205 2366 12235 2450
rect 12315 2366 12345 2450
rect 12411 2366 12441 2438
rect 12517 2366 12547 2438
rect 12612 2366 12642 2450
rect 12800 2366 12830 2450
rect 12884 2366 12914 2450
<< scpmoshvt >>
rect 1114 5966 1144 6124
rect 1202 5966 1232 6124
rect 1390 5924 1420 6124
rect 1474 5924 1504 6124
rect 1558 5924 1588 6124
rect 1642 5924 1672 6124
rect 1726 5924 1756 6124
rect 2389 5924 2419 6124
rect 2473 5924 2503 6124
rect 2573 5924 2603 6124
rect 2657 5924 2687 6124
rect 2754 5996 2784 6124
rect 2855 6040 2885 6124
rect 2939 6040 2969 6124
rect 3074 5996 3104 6124
rect 3262 5943 3292 6051
rect 3346 5943 3376 6051
rect 3534 5972 3564 6100
rect 3618 5972 3648 6100
rect 3762 6040 3792 6124
rect 3846 6040 3876 6124
rect 3942 5996 3972 6124
rect 4026 5996 4056 6124
rect 1113 5117 1143 5245
rect 1197 5117 1227 5245
rect 1385 5167 1415 5251
rect 1478 5167 1508 5251
rect 1562 5167 1592 5251
rect 1682 5167 1712 5251
rect 1788 5167 1818 5251
rect 1896 5083 1926 5251
rect 1980 5083 2010 5251
rect 2117 5083 2147 5251
rect 2261 5167 2291 5251
rect 2345 5167 2375 5251
rect 2463 5167 2493 5251
rect 2571 5167 2601 5251
rect 2667 5083 2697 5251
rect 2739 5083 2769 5251
rect 2937 5055 2967 5183
rect 3034 5051 3064 5251
rect 3222 5107 3252 5235
rect 3317 5051 3347 5251
rect 3505 5117 3535 5245
rect 3589 5117 3619 5245
rect 3777 5167 3807 5251
rect 3870 5167 3900 5251
rect 3954 5167 3984 5251
rect 4074 5167 4104 5251
rect 4180 5167 4210 5251
rect 4288 5083 4318 5251
rect 4372 5083 4402 5251
rect 4509 5083 4539 5251
rect 4653 5167 4683 5251
rect 4737 5167 4767 5251
rect 4855 5167 4885 5251
rect 4963 5167 4993 5251
rect 5059 5083 5089 5251
rect 5131 5083 5161 5251
rect 5329 5055 5359 5183
rect 5426 5051 5456 5251
rect 5614 5107 5644 5235
rect 5709 5051 5739 5251
rect 5897 5117 5927 5245
rect 5981 5117 6011 5245
rect 6169 5167 6199 5251
rect 6262 5167 6292 5251
rect 6346 5167 6376 5251
rect 6466 5167 6496 5251
rect 6572 5167 6602 5251
rect 6680 5083 6710 5251
rect 6764 5083 6794 5251
rect 6901 5083 6931 5251
rect 7045 5167 7075 5251
rect 7129 5167 7159 5251
rect 7247 5167 7277 5251
rect 7355 5167 7385 5251
rect 7451 5083 7481 5251
rect 7523 5083 7553 5251
rect 7721 5055 7751 5183
rect 7818 5051 7848 5251
rect 8006 5107 8036 5235
rect 8101 5051 8131 5251
rect 8289 5117 8319 5245
rect 8373 5117 8403 5245
rect 8561 5167 8591 5251
rect 8654 5167 8684 5251
rect 8738 5167 8768 5251
rect 8858 5167 8888 5251
rect 8964 5167 8994 5251
rect 9072 5083 9102 5251
rect 9156 5083 9186 5251
rect 9293 5083 9323 5251
rect 9437 5167 9467 5251
rect 9521 5167 9551 5251
rect 9639 5167 9669 5251
rect 9747 5167 9777 5251
rect 9843 5083 9873 5251
rect 9915 5083 9945 5251
rect 10113 5055 10143 5183
rect 10210 5051 10240 5251
rect 10398 5107 10428 5235
rect 10493 5051 10523 5251
rect 10681 5117 10711 5245
rect 10765 5117 10795 5245
rect 10953 5167 10983 5251
rect 11046 5167 11076 5251
rect 11130 5167 11160 5251
rect 11250 5167 11280 5251
rect 11356 5167 11386 5251
rect 11464 5083 11494 5251
rect 11548 5083 11578 5251
rect 11685 5083 11715 5251
rect 11829 5167 11859 5251
rect 11913 5167 11943 5251
rect 12031 5167 12061 5251
rect 12139 5167 12169 5251
rect 12235 5083 12265 5251
rect 12307 5083 12337 5251
rect 12505 5055 12535 5183
rect 12602 5051 12632 5251
rect 12790 5107 12820 5235
rect 12885 5051 12915 5251
rect 673 4404 703 4562
rect 761 4404 791 4562
rect 949 4362 979 4562
rect 1033 4362 1063 4562
rect 1117 4362 1147 4562
rect 1201 4362 1231 4562
rect 1285 4362 1315 4562
rect 1481 4362 1511 4562
rect 1565 4362 1595 4562
rect 1649 4362 1679 4562
rect 1733 4362 1763 4562
rect 1817 4362 1847 4562
rect 1901 4362 1931 4562
rect 1985 4362 2015 4562
rect 2069 4362 2099 4562
rect 2153 4362 2183 4562
rect 2237 4362 2267 4562
rect 2321 4362 2351 4562
rect 2405 4362 2435 4562
rect 2489 4362 2519 4562
rect 2573 4362 2603 4562
rect 2657 4362 2687 4562
rect 2741 4362 2771 4562
rect 2825 4362 2855 4562
rect 2909 4362 2939 4562
rect 2993 4362 3023 4562
rect 3077 4362 3107 4562
rect 3161 4362 3191 4562
rect 3245 4362 3275 4562
rect 3505 4362 3535 4562
rect 3600 4418 3630 4546
rect 3788 4362 3818 4562
rect 3885 4366 3915 4494
rect 4083 4394 4113 4562
rect 4155 4394 4185 4562
rect 4251 4478 4281 4562
rect 4359 4478 4389 4562
rect 4477 4478 4507 4562
rect 4561 4478 4591 4562
rect 4705 4394 4735 4562
rect 4842 4394 4872 4562
rect 4926 4394 4956 4562
rect 5034 4478 5064 4562
rect 5140 4478 5170 4562
rect 5260 4478 5290 4562
rect 5344 4478 5374 4562
rect 5437 4478 5467 4562
rect 5625 4428 5655 4556
rect 5709 4428 5739 4556
rect 5897 4362 5927 4562
rect 5992 4418 6022 4546
rect 6180 4362 6210 4562
rect 6277 4366 6307 4494
rect 6475 4394 6505 4562
rect 6547 4394 6577 4562
rect 6643 4478 6673 4562
rect 6751 4478 6781 4562
rect 6869 4478 6899 4562
rect 6953 4478 6983 4562
rect 7097 4394 7127 4562
rect 7234 4394 7264 4562
rect 7318 4394 7348 4562
rect 7426 4478 7456 4562
rect 7532 4478 7562 4562
rect 7652 4478 7682 4562
rect 7736 4478 7766 4562
rect 7829 4478 7859 4562
rect 8017 4428 8047 4556
rect 8101 4428 8131 4556
rect 8289 4362 8319 4562
rect 8384 4418 8414 4546
rect 8572 4362 8602 4562
rect 8669 4366 8699 4494
rect 8867 4394 8897 4562
rect 8939 4394 8969 4562
rect 9035 4478 9065 4562
rect 9143 4478 9173 4562
rect 9261 4478 9291 4562
rect 9345 4478 9375 4562
rect 9489 4394 9519 4562
rect 9626 4394 9656 4562
rect 9710 4394 9740 4562
rect 9818 4478 9848 4562
rect 9924 4478 9954 4562
rect 10044 4478 10074 4562
rect 10128 4478 10158 4562
rect 10221 4478 10251 4562
rect 10409 4428 10439 4556
rect 10493 4428 10523 4556
rect 10681 4362 10711 4562
rect 10776 4418 10806 4546
rect 10964 4362 10994 4562
rect 11061 4366 11091 4494
rect 11259 4394 11289 4562
rect 11331 4394 11361 4562
rect 11427 4478 11457 4562
rect 11535 4478 11565 4562
rect 11653 4478 11683 4562
rect 11737 4478 11767 4562
rect 11881 4394 11911 4562
rect 12018 4394 12048 4562
rect 12102 4394 12132 4562
rect 12210 4478 12240 4562
rect 12316 4478 12346 4562
rect 12436 4478 12466 4562
rect 12520 4478 12550 4562
rect 12613 4478 12643 4562
rect 12801 4428 12831 4556
rect 12885 4428 12915 4556
rect 705 3530 735 3688
rect 793 3530 823 3688
rect 981 3488 1011 3688
rect 1065 3488 1095 3688
rect 1149 3488 1179 3688
rect 1233 3488 1263 3688
rect 1317 3488 1347 3688
rect 3288 3489 3318 3689
rect 3504 3555 3534 3683
rect 3588 3555 3618 3683
rect 3776 3605 3806 3689
rect 3869 3605 3899 3689
rect 3953 3605 3983 3689
rect 4073 3605 4103 3689
rect 4179 3605 4209 3689
rect 4287 3521 4317 3689
rect 4371 3521 4401 3689
rect 4508 3521 4538 3689
rect 4652 3605 4682 3689
rect 4736 3605 4766 3689
rect 4854 3605 4884 3689
rect 4962 3605 4992 3689
rect 5058 3521 5088 3689
rect 5130 3521 5160 3689
rect 5328 3493 5358 3621
rect 5425 3489 5455 3689
rect 5613 3545 5643 3673
rect 5708 3489 5738 3689
rect 5896 3555 5926 3683
rect 5980 3555 6010 3683
rect 6168 3605 6198 3689
rect 6261 3605 6291 3689
rect 6345 3605 6375 3689
rect 6465 3605 6495 3689
rect 6571 3605 6601 3689
rect 6679 3521 6709 3689
rect 6763 3521 6793 3689
rect 6900 3521 6930 3689
rect 7044 3605 7074 3689
rect 7128 3605 7158 3689
rect 7246 3605 7276 3689
rect 7354 3605 7384 3689
rect 7450 3521 7480 3689
rect 7522 3521 7552 3689
rect 7720 3493 7750 3621
rect 7817 3489 7847 3689
rect 8005 3545 8035 3673
rect 8100 3489 8130 3689
rect 8288 3555 8318 3683
rect 8372 3555 8402 3683
rect 8560 3605 8590 3689
rect 8653 3605 8683 3689
rect 8737 3605 8767 3689
rect 8857 3605 8887 3689
rect 8963 3605 8993 3689
rect 9071 3521 9101 3689
rect 9155 3521 9185 3689
rect 9292 3521 9322 3689
rect 9436 3605 9466 3689
rect 9520 3605 9550 3689
rect 9638 3605 9668 3689
rect 9746 3605 9776 3689
rect 9842 3521 9872 3689
rect 9914 3521 9944 3689
rect 10112 3493 10142 3621
rect 10209 3489 10239 3689
rect 10397 3545 10427 3673
rect 10492 3489 10522 3689
rect 10680 3555 10710 3683
rect 10764 3555 10794 3683
rect 10952 3605 10982 3689
rect 11045 3605 11075 3689
rect 11129 3605 11159 3689
rect 11249 3605 11279 3689
rect 11355 3605 11385 3689
rect 11463 3521 11493 3689
rect 11547 3521 11577 3689
rect 11684 3521 11714 3689
rect 11828 3605 11858 3689
rect 11912 3605 11942 3689
rect 12030 3605 12060 3689
rect 12138 3605 12168 3689
rect 12234 3521 12264 3689
rect 12306 3521 12336 3689
rect 12504 3493 12534 3621
rect 12601 3489 12631 3689
rect 12789 3545 12819 3673
rect 12884 3489 12914 3689
rect 1112 2616 1142 2816
rect 1207 2672 1237 2800
rect 1395 2616 1425 2816
rect 1492 2620 1522 2748
rect 1690 2648 1720 2816
rect 1762 2648 1792 2816
rect 1858 2732 1888 2816
rect 1966 2732 1996 2816
rect 2084 2732 2114 2816
rect 2168 2732 2198 2816
rect 2312 2648 2342 2816
rect 2449 2648 2479 2816
rect 2533 2648 2563 2816
rect 2641 2732 2671 2816
rect 2747 2732 2777 2816
rect 2867 2732 2897 2816
rect 2951 2732 2981 2816
rect 3044 2732 3074 2816
rect 3232 2682 3262 2810
rect 3316 2682 3346 2810
rect 3504 2616 3534 2816
rect 3599 2672 3629 2800
rect 3787 2616 3817 2816
rect 3884 2620 3914 2748
rect 4082 2648 4112 2816
rect 4154 2648 4184 2816
rect 4250 2732 4280 2816
rect 4358 2732 4388 2816
rect 4476 2732 4506 2816
rect 4560 2732 4590 2816
rect 4704 2648 4734 2816
rect 4841 2648 4871 2816
rect 4925 2648 4955 2816
rect 5033 2732 5063 2816
rect 5139 2732 5169 2816
rect 5259 2732 5289 2816
rect 5343 2732 5373 2816
rect 5436 2732 5466 2816
rect 5624 2682 5654 2810
rect 5708 2682 5738 2810
rect 5896 2616 5926 2816
rect 5991 2672 6021 2800
rect 6179 2616 6209 2816
rect 6276 2620 6306 2748
rect 6474 2648 6504 2816
rect 6546 2648 6576 2816
rect 6642 2732 6672 2816
rect 6750 2732 6780 2816
rect 6868 2732 6898 2816
rect 6952 2732 6982 2816
rect 7096 2648 7126 2816
rect 7233 2648 7263 2816
rect 7317 2648 7347 2816
rect 7425 2732 7455 2816
rect 7531 2732 7561 2816
rect 7651 2732 7681 2816
rect 7735 2732 7765 2816
rect 7828 2732 7858 2816
rect 8016 2682 8046 2810
rect 8100 2682 8130 2810
rect 8288 2616 8318 2816
rect 8383 2672 8413 2800
rect 8571 2616 8601 2816
rect 8668 2620 8698 2748
rect 8866 2648 8896 2816
rect 8938 2648 8968 2816
rect 9034 2732 9064 2816
rect 9142 2732 9172 2816
rect 9260 2732 9290 2816
rect 9344 2732 9374 2816
rect 9488 2648 9518 2816
rect 9625 2648 9655 2816
rect 9709 2648 9739 2816
rect 9817 2732 9847 2816
rect 9923 2732 9953 2816
rect 10043 2732 10073 2816
rect 10127 2732 10157 2816
rect 10220 2732 10250 2816
rect 10408 2682 10438 2810
rect 10492 2682 10522 2810
rect 10680 2616 10710 2816
rect 10775 2672 10805 2800
rect 10963 2616 10993 2816
rect 11060 2620 11090 2748
rect 11258 2648 11288 2816
rect 11330 2648 11360 2816
rect 11426 2732 11456 2816
rect 11534 2732 11564 2816
rect 11652 2732 11682 2816
rect 11736 2732 11766 2816
rect 11880 2648 11910 2816
rect 12017 2648 12047 2816
rect 12101 2648 12131 2816
rect 12209 2732 12239 2816
rect 12315 2732 12345 2816
rect 12435 2732 12465 2816
rect 12519 2732 12549 2816
rect 12612 2732 12642 2816
rect 12800 2682 12830 2810
rect 12884 2682 12914 2810
<< ndiff >>
rect 1062 5733 1114 5778
rect 1062 5699 1070 5733
rect 1104 5699 1114 5733
rect 1062 5674 1114 5699
rect 1144 5720 1202 5778
rect 1144 5686 1156 5720
rect 1190 5686 1202 5720
rect 1144 5674 1202 5686
rect 1232 5750 1284 5778
rect 1232 5716 1242 5750
rect 1276 5716 1284 5750
rect 1232 5674 1284 5716
rect 1338 5756 1390 5804
rect 1338 5722 1346 5756
rect 1380 5722 1390 5756
rect 1338 5674 1390 5722
rect 1420 5724 1474 5804
rect 1420 5690 1430 5724
rect 1464 5690 1474 5724
rect 1420 5674 1474 5690
rect 1504 5756 1558 5804
rect 1504 5722 1514 5756
rect 1548 5722 1558 5756
rect 1504 5674 1558 5722
rect 1588 5724 1642 5804
rect 1588 5690 1598 5724
rect 1632 5690 1642 5724
rect 1588 5674 1642 5690
rect 1672 5756 1726 5804
rect 1672 5722 1682 5756
rect 1716 5722 1726 5756
rect 1672 5674 1726 5722
rect 1756 5788 1808 5804
rect 1756 5754 1766 5788
rect 1800 5754 1808 5788
rect 1756 5720 1808 5754
rect 1756 5686 1766 5720
rect 1800 5686 1808 5720
rect 1756 5674 1808 5686
rect 2322 5788 2389 5804
rect 2322 5754 2330 5788
rect 2364 5754 2389 5788
rect 2322 5720 2389 5754
rect 2322 5686 2330 5720
rect 2364 5686 2389 5720
rect 2322 5674 2389 5686
rect 2419 5756 2473 5804
rect 2419 5722 2429 5756
rect 2463 5722 2473 5756
rect 2419 5674 2473 5722
rect 2503 5788 2573 5804
rect 2503 5754 2513 5788
rect 2547 5754 2573 5788
rect 2503 5720 2573 5754
rect 2503 5686 2513 5720
rect 2547 5686 2573 5720
rect 2503 5674 2573 5686
rect 2603 5756 2657 5804
rect 2603 5722 2613 5756
rect 2647 5722 2657 5756
rect 2603 5674 2657 5722
rect 2687 5758 2743 5804
rect 2687 5746 2758 5758
rect 2687 5712 2697 5746
rect 2731 5712 2758 5746
rect 2687 5674 2758 5712
rect 2788 5746 2838 5758
rect 3008 5746 3070 5758
rect 2788 5674 2853 5746
rect 2883 5720 2963 5746
rect 2883 5686 2906 5720
rect 2940 5686 2963 5720
rect 2883 5674 2963 5686
rect 2993 5674 3070 5746
rect 3100 5720 3152 5758
rect 3100 5686 3110 5720
rect 3144 5686 3152 5720
rect 3100 5674 3152 5686
rect 3206 5728 3258 5758
rect 3206 5694 3214 5728
rect 3248 5694 3258 5728
rect 3206 5674 3258 5694
rect 3288 5746 3343 5758
rect 3288 5712 3298 5746
rect 3332 5712 3343 5746
rect 3288 5674 3343 5712
rect 3373 5746 3425 5758
rect 3373 5712 3383 5746
rect 3417 5712 3425 5746
rect 3373 5674 3425 5712
rect 3479 5720 3533 5758
rect 3479 5686 3487 5720
rect 3521 5686 3533 5720
rect 3479 5674 3533 5686
rect 3563 5720 3641 5758
rect 3563 5686 3586 5720
rect 3620 5686 3641 5720
rect 3563 5674 3641 5686
rect 3671 5746 3722 5758
rect 3892 5746 3942 5758
rect 3671 5674 3737 5746
rect 3767 5734 3847 5746
rect 3767 5700 3790 5734
rect 3824 5700 3847 5734
rect 3767 5674 3847 5700
rect 3877 5674 3942 5746
rect 3972 5720 4026 5758
rect 3972 5686 3982 5720
rect 4016 5686 4026 5720
rect 3972 5674 4026 5686
rect 4056 5746 4108 5758
rect 4056 5712 4066 5746
rect 4100 5712 4108 5746
rect 4056 5674 4108 5712
rect 1061 4873 1113 4885
rect 1061 4839 1069 4873
rect 1103 4839 1113 4873
rect 1061 4801 1113 4839
rect 1143 4847 1197 4885
rect 1143 4813 1153 4847
rect 1187 4813 1197 4847
rect 1143 4801 1197 4813
rect 1227 4873 1279 4885
rect 1227 4839 1237 4873
rect 1271 4839 1279 4873
rect 1227 4801 1279 4839
rect 1333 4847 1385 4885
rect 1333 4813 1341 4847
rect 1375 4813 1385 4847
rect 1333 4801 1385 4813
rect 1415 4873 1465 4885
rect 1842 4885 1892 4929
rect 1631 4873 1682 4885
rect 1415 4865 1480 4873
rect 1415 4831 1425 4865
rect 1459 4831 1480 4865
rect 1415 4801 1480 4831
rect 1510 4847 1586 4873
rect 1510 4813 1531 4847
rect 1565 4813 1586 4847
rect 1510 4801 1586 4813
rect 1616 4801 1682 4873
rect 1712 4843 1792 4885
rect 1712 4809 1748 4843
rect 1782 4809 1792 4843
rect 1712 4801 1792 4809
rect 1822 4863 1892 4885
rect 1822 4829 1832 4863
rect 1866 4829 1892 4863
rect 1822 4801 1892 4829
rect 1922 4907 1976 4929
rect 1922 4873 1932 4907
rect 1966 4873 1976 4907
rect 1922 4801 1976 4873
rect 2006 4881 2058 4929
rect 2006 4847 2016 4881
rect 2050 4847 2058 4881
rect 2006 4801 2058 4847
rect 2112 4847 2164 4929
rect 2112 4813 2120 4847
rect 2154 4813 2164 4847
rect 2112 4801 2164 4813
rect 2194 4873 2244 4929
rect 2617 4885 2667 4929
rect 2413 4873 2463 4885
rect 2194 4801 2259 4873
rect 2289 4847 2368 4873
rect 2289 4813 2314 4847
rect 2348 4813 2368 4847
rect 2289 4801 2368 4813
rect 2398 4801 2463 4873
rect 2493 4843 2549 4885
rect 2493 4809 2505 4843
rect 2539 4809 2549 4843
rect 2493 4801 2549 4809
rect 2579 4863 2667 4885
rect 2579 4829 2607 4863
rect 2641 4829 2667 4863
rect 2579 4801 2667 4829
rect 2697 4907 2751 4929
rect 2697 4873 2707 4907
rect 2741 4873 2751 4907
rect 2697 4801 2751 4873
rect 2781 4855 2833 4929
rect 2984 4885 3034 4931
rect 2781 4821 2791 4855
rect 2825 4821 2833 4855
rect 2781 4801 2833 4821
rect 2887 4857 2939 4885
rect 2887 4823 2895 4857
rect 2929 4823 2939 4857
rect 2887 4801 2939 4823
rect 2969 4847 3034 4885
rect 2969 4813 2990 4847
rect 3024 4813 3034 4847
rect 2969 4801 3034 4813
rect 3064 4881 3116 4931
rect 3267 4885 3317 4931
rect 3064 4847 3074 4881
rect 3108 4847 3116 4881
rect 3064 4801 3116 4847
rect 3170 4873 3222 4885
rect 3170 4839 3178 4873
rect 3212 4839 3222 4873
rect 3170 4801 3222 4839
rect 3252 4847 3317 4885
rect 3252 4813 3273 4847
rect 3307 4813 3317 4847
rect 3252 4801 3317 4813
rect 3347 4883 3399 4931
rect 3347 4849 3357 4883
rect 3391 4849 3399 4883
rect 3347 4801 3399 4849
rect 3453 4873 3505 4885
rect 3453 4839 3461 4873
rect 3495 4839 3505 4873
rect 3453 4801 3505 4839
rect 3535 4847 3589 4885
rect 3535 4813 3545 4847
rect 3579 4813 3589 4847
rect 3535 4801 3589 4813
rect 3619 4873 3671 4885
rect 3619 4839 3629 4873
rect 3663 4839 3671 4873
rect 3619 4801 3671 4839
rect 3725 4847 3777 4885
rect 3725 4813 3733 4847
rect 3767 4813 3777 4847
rect 3725 4801 3777 4813
rect 3807 4873 3857 4885
rect 4234 4885 4284 4929
rect 4023 4873 4074 4885
rect 3807 4865 3872 4873
rect 3807 4831 3817 4865
rect 3851 4831 3872 4865
rect 3807 4801 3872 4831
rect 3902 4847 3978 4873
rect 3902 4813 3923 4847
rect 3957 4813 3978 4847
rect 3902 4801 3978 4813
rect 4008 4801 4074 4873
rect 4104 4843 4184 4885
rect 4104 4809 4140 4843
rect 4174 4809 4184 4843
rect 4104 4801 4184 4809
rect 4214 4863 4284 4885
rect 4214 4829 4224 4863
rect 4258 4829 4284 4863
rect 4214 4801 4284 4829
rect 4314 4907 4368 4929
rect 4314 4873 4324 4907
rect 4358 4873 4368 4907
rect 4314 4801 4368 4873
rect 4398 4881 4450 4929
rect 4398 4847 4408 4881
rect 4442 4847 4450 4881
rect 4398 4801 4450 4847
rect 4504 4847 4556 4929
rect 4504 4813 4512 4847
rect 4546 4813 4556 4847
rect 4504 4801 4556 4813
rect 4586 4873 4636 4929
rect 5009 4885 5059 4929
rect 4805 4873 4855 4885
rect 4586 4801 4651 4873
rect 4681 4847 4760 4873
rect 4681 4813 4706 4847
rect 4740 4813 4760 4847
rect 4681 4801 4760 4813
rect 4790 4801 4855 4873
rect 4885 4843 4941 4885
rect 4885 4809 4897 4843
rect 4931 4809 4941 4843
rect 4885 4801 4941 4809
rect 4971 4863 5059 4885
rect 4971 4829 4999 4863
rect 5033 4829 5059 4863
rect 4971 4801 5059 4829
rect 5089 4907 5143 4929
rect 5089 4873 5099 4907
rect 5133 4873 5143 4907
rect 5089 4801 5143 4873
rect 5173 4855 5225 4929
rect 5376 4885 5426 4931
rect 5173 4821 5183 4855
rect 5217 4821 5225 4855
rect 5173 4801 5225 4821
rect 5279 4857 5331 4885
rect 5279 4823 5287 4857
rect 5321 4823 5331 4857
rect 5279 4801 5331 4823
rect 5361 4847 5426 4885
rect 5361 4813 5382 4847
rect 5416 4813 5426 4847
rect 5361 4801 5426 4813
rect 5456 4881 5508 4931
rect 5659 4885 5709 4931
rect 5456 4847 5466 4881
rect 5500 4847 5508 4881
rect 5456 4801 5508 4847
rect 5562 4873 5614 4885
rect 5562 4839 5570 4873
rect 5604 4839 5614 4873
rect 5562 4801 5614 4839
rect 5644 4847 5709 4885
rect 5644 4813 5665 4847
rect 5699 4813 5709 4847
rect 5644 4801 5709 4813
rect 5739 4883 5791 4931
rect 5739 4849 5749 4883
rect 5783 4849 5791 4883
rect 5739 4801 5791 4849
rect 5845 4873 5897 4885
rect 5845 4839 5853 4873
rect 5887 4839 5897 4873
rect 5845 4801 5897 4839
rect 5927 4847 5981 4885
rect 5927 4813 5937 4847
rect 5971 4813 5981 4847
rect 5927 4801 5981 4813
rect 6011 4873 6063 4885
rect 6011 4839 6021 4873
rect 6055 4839 6063 4873
rect 6011 4801 6063 4839
rect 6117 4847 6169 4885
rect 6117 4813 6125 4847
rect 6159 4813 6169 4847
rect 6117 4801 6169 4813
rect 6199 4873 6249 4885
rect 6626 4885 6676 4929
rect 6415 4873 6466 4885
rect 6199 4865 6264 4873
rect 6199 4831 6209 4865
rect 6243 4831 6264 4865
rect 6199 4801 6264 4831
rect 6294 4847 6370 4873
rect 6294 4813 6315 4847
rect 6349 4813 6370 4847
rect 6294 4801 6370 4813
rect 6400 4801 6466 4873
rect 6496 4843 6576 4885
rect 6496 4809 6532 4843
rect 6566 4809 6576 4843
rect 6496 4801 6576 4809
rect 6606 4863 6676 4885
rect 6606 4829 6616 4863
rect 6650 4829 6676 4863
rect 6606 4801 6676 4829
rect 6706 4907 6760 4929
rect 6706 4873 6716 4907
rect 6750 4873 6760 4907
rect 6706 4801 6760 4873
rect 6790 4881 6842 4929
rect 6790 4847 6800 4881
rect 6834 4847 6842 4881
rect 6790 4801 6842 4847
rect 6896 4847 6948 4929
rect 6896 4813 6904 4847
rect 6938 4813 6948 4847
rect 6896 4801 6948 4813
rect 6978 4873 7028 4929
rect 7401 4885 7451 4929
rect 7197 4873 7247 4885
rect 6978 4801 7043 4873
rect 7073 4847 7152 4873
rect 7073 4813 7098 4847
rect 7132 4813 7152 4847
rect 7073 4801 7152 4813
rect 7182 4801 7247 4873
rect 7277 4843 7333 4885
rect 7277 4809 7289 4843
rect 7323 4809 7333 4843
rect 7277 4801 7333 4809
rect 7363 4863 7451 4885
rect 7363 4829 7391 4863
rect 7425 4829 7451 4863
rect 7363 4801 7451 4829
rect 7481 4907 7535 4929
rect 7481 4873 7491 4907
rect 7525 4873 7535 4907
rect 7481 4801 7535 4873
rect 7565 4855 7617 4929
rect 7768 4885 7818 4931
rect 7565 4821 7575 4855
rect 7609 4821 7617 4855
rect 7565 4801 7617 4821
rect 7671 4857 7723 4885
rect 7671 4823 7679 4857
rect 7713 4823 7723 4857
rect 7671 4801 7723 4823
rect 7753 4847 7818 4885
rect 7753 4813 7774 4847
rect 7808 4813 7818 4847
rect 7753 4801 7818 4813
rect 7848 4881 7900 4931
rect 8051 4885 8101 4931
rect 7848 4847 7858 4881
rect 7892 4847 7900 4881
rect 7848 4801 7900 4847
rect 7954 4873 8006 4885
rect 7954 4839 7962 4873
rect 7996 4839 8006 4873
rect 7954 4801 8006 4839
rect 8036 4847 8101 4885
rect 8036 4813 8057 4847
rect 8091 4813 8101 4847
rect 8036 4801 8101 4813
rect 8131 4883 8183 4931
rect 8131 4849 8141 4883
rect 8175 4849 8183 4883
rect 8131 4801 8183 4849
rect 8237 4873 8289 4885
rect 8237 4839 8245 4873
rect 8279 4839 8289 4873
rect 8237 4801 8289 4839
rect 8319 4847 8373 4885
rect 8319 4813 8329 4847
rect 8363 4813 8373 4847
rect 8319 4801 8373 4813
rect 8403 4873 8455 4885
rect 8403 4839 8413 4873
rect 8447 4839 8455 4873
rect 8403 4801 8455 4839
rect 8509 4847 8561 4885
rect 8509 4813 8517 4847
rect 8551 4813 8561 4847
rect 8509 4801 8561 4813
rect 8591 4873 8641 4885
rect 9018 4885 9068 4929
rect 8807 4873 8858 4885
rect 8591 4865 8656 4873
rect 8591 4831 8601 4865
rect 8635 4831 8656 4865
rect 8591 4801 8656 4831
rect 8686 4847 8762 4873
rect 8686 4813 8707 4847
rect 8741 4813 8762 4847
rect 8686 4801 8762 4813
rect 8792 4801 8858 4873
rect 8888 4843 8968 4885
rect 8888 4809 8924 4843
rect 8958 4809 8968 4843
rect 8888 4801 8968 4809
rect 8998 4863 9068 4885
rect 8998 4829 9008 4863
rect 9042 4829 9068 4863
rect 8998 4801 9068 4829
rect 9098 4907 9152 4929
rect 9098 4873 9108 4907
rect 9142 4873 9152 4907
rect 9098 4801 9152 4873
rect 9182 4881 9234 4929
rect 9182 4847 9192 4881
rect 9226 4847 9234 4881
rect 9182 4801 9234 4847
rect 9288 4847 9340 4929
rect 9288 4813 9296 4847
rect 9330 4813 9340 4847
rect 9288 4801 9340 4813
rect 9370 4873 9420 4929
rect 9793 4885 9843 4929
rect 9589 4873 9639 4885
rect 9370 4801 9435 4873
rect 9465 4847 9544 4873
rect 9465 4813 9490 4847
rect 9524 4813 9544 4847
rect 9465 4801 9544 4813
rect 9574 4801 9639 4873
rect 9669 4843 9725 4885
rect 9669 4809 9681 4843
rect 9715 4809 9725 4843
rect 9669 4801 9725 4809
rect 9755 4863 9843 4885
rect 9755 4829 9783 4863
rect 9817 4829 9843 4863
rect 9755 4801 9843 4829
rect 9873 4907 9927 4929
rect 9873 4873 9883 4907
rect 9917 4873 9927 4907
rect 9873 4801 9927 4873
rect 9957 4855 10009 4929
rect 10160 4885 10210 4931
rect 9957 4821 9967 4855
rect 10001 4821 10009 4855
rect 9957 4801 10009 4821
rect 10063 4857 10115 4885
rect 10063 4823 10071 4857
rect 10105 4823 10115 4857
rect 10063 4801 10115 4823
rect 10145 4847 10210 4885
rect 10145 4813 10166 4847
rect 10200 4813 10210 4847
rect 10145 4801 10210 4813
rect 10240 4881 10292 4931
rect 10443 4885 10493 4931
rect 10240 4847 10250 4881
rect 10284 4847 10292 4881
rect 10240 4801 10292 4847
rect 10346 4873 10398 4885
rect 10346 4839 10354 4873
rect 10388 4839 10398 4873
rect 10346 4801 10398 4839
rect 10428 4847 10493 4885
rect 10428 4813 10449 4847
rect 10483 4813 10493 4847
rect 10428 4801 10493 4813
rect 10523 4883 10575 4931
rect 10523 4849 10533 4883
rect 10567 4849 10575 4883
rect 10523 4801 10575 4849
rect 10629 4873 10681 4885
rect 10629 4839 10637 4873
rect 10671 4839 10681 4873
rect 10629 4801 10681 4839
rect 10711 4847 10765 4885
rect 10711 4813 10721 4847
rect 10755 4813 10765 4847
rect 10711 4801 10765 4813
rect 10795 4873 10847 4885
rect 10795 4839 10805 4873
rect 10839 4839 10847 4873
rect 10795 4801 10847 4839
rect 10901 4847 10953 4885
rect 10901 4813 10909 4847
rect 10943 4813 10953 4847
rect 10901 4801 10953 4813
rect 10983 4873 11033 4885
rect 11410 4885 11460 4929
rect 11199 4873 11250 4885
rect 10983 4865 11048 4873
rect 10983 4831 10993 4865
rect 11027 4831 11048 4865
rect 10983 4801 11048 4831
rect 11078 4847 11154 4873
rect 11078 4813 11099 4847
rect 11133 4813 11154 4847
rect 11078 4801 11154 4813
rect 11184 4801 11250 4873
rect 11280 4843 11360 4885
rect 11280 4809 11316 4843
rect 11350 4809 11360 4843
rect 11280 4801 11360 4809
rect 11390 4863 11460 4885
rect 11390 4829 11400 4863
rect 11434 4829 11460 4863
rect 11390 4801 11460 4829
rect 11490 4907 11544 4929
rect 11490 4873 11500 4907
rect 11534 4873 11544 4907
rect 11490 4801 11544 4873
rect 11574 4881 11626 4929
rect 11574 4847 11584 4881
rect 11618 4847 11626 4881
rect 11574 4801 11626 4847
rect 11680 4847 11732 4929
rect 11680 4813 11688 4847
rect 11722 4813 11732 4847
rect 11680 4801 11732 4813
rect 11762 4873 11812 4929
rect 12185 4885 12235 4929
rect 11981 4873 12031 4885
rect 11762 4801 11827 4873
rect 11857 4847 11936 4873
rect 11857 4813 11882 4847
rect 11916 4813 11936 4847
rect 11857 4801 11936 4813
rect 11966 4801 12031 4873
rect 12061 4843 12117 4885
rect 12061 4809 12073 4843
rect 12107 4809 12117 4843
rect 12061 4801 12117 4809
rect 12147 4863 12235 4885
rect 12147 4829 12175 4863
rect 12209 4829 12235 4863
rect 12147 4801 12235 4829
rect 12265 4907 12319 4929
rect 12265 4873 12275 4907
rect 12309 4873 12319 4907
rect 12265 4801 12319 4873
rect 12349 4855 12401 4929
rect 12552 4885 12602 4931
rect 12349 4821 12359 4855
rect 12393 4821 12401 4855
rect 12349 4801 12401 4821
rect 12455 4857 12507 4885
rect 12455 4823 12463 4857
rect 12497 4823 12507 4857
rect 12455 4801 12507 4823
rect 12537 4847 12602 4885
rect 12537 4813 12558 4847
rect 12592 4813 12602 4847
rect 12537 4801 12602 4813
rect 12632 4881 12684 4931
rect 12835 4885 12885 4931
rect 12632 4847 12642 4881
rect 12676 4847 12684 4881
rect 12632 4801 12684 4847
rect 12738 4873 12790 4885
rect 12738 4839 12746 4873
rect 12780 4839 12790 4873
rect 12738 4801 12790 4839
rect 12820 4847 12885 4885
rect 12820 4813 12841 4847
rect 12875 4813 12885 4847
rect 12820 4801 12885 4813
rect 12915 4883 12967 4931
rect 12915 4849 12925 4883
rect 12959 4849 12967 4883
rect 12915 4801 12967 4849
rect 621 4171 673 4216
rect 621 4137 629 4171
rect 663 4137 673 4171
rect 621 4112 673 4137
rect 703 4158 761 4216
rect 703 4124 715 4158
rect 749 4124 761 4158
rect 703 4112 761 4124
rect 791 4188 843 4216
rect 791 4154 801 4188
rect 835 4154 843 4188
rect 791 4112 843 4154
rect 897 4194 949 4242
rect 897 4160 905 4194
rect 939 4160 949 4194
rect 897 4112 949 4160
rect 979 4162 1033 4242
rect 979 4128 989 4162
rect 1023 4128 1033 4162
rect 979 4112 1033 4128
rect 1063 4194 1117 4242
rect 1063 4160 1073 4194
rect 1107 4160 1117 4194
rect 1063 4112 1117 4160
rect 1147 4162 1201 4242
rect 1147 4128 1157 4162
rect 1191 4128 1201 4162
rect 1147 4112 1201 4128
rect 1231 4194 1285 4242
rect 1231 4160 1241 4194
rect 1275 4160 1285 4194
rect 1231 4112 1285 4160
rect 1315 4226 1367 4242
rect 1315 4192 1325 4226
rect 1359 4192 1367 4226
rect 1315 4158 1367 4192
rect 1315 4124 1325 4158
rect 1359 4124 1367 4158
rect 1315 4112 1367 4124
rect 1429 4230 1481 4242
rect 1429 4196 1437 4230
rect 1471 4196 1481 4230
rect 1429 4162 1481 4196
rect 1429 4128 1437 4162
rect 1471 4128 1481 4162
rect 1429 4112 1481 4128
rect 1511 4230 1565 4242
rect 1511 4196 1521 4230
rect 1555 4196 1565 4230
rect 1511 4162 1565 4196
rect 1511 4128 1521 4162
rect 1555 4128 1565 4162
rect 1511 4112 1565 4128
rect 1595 4162 1649 4242
rect 1595 4128 1605 4162
rect 1639 4128 1649 4162
rect 1595 4112 1649 4128
rect 1679 4230 1733 4242
rect 1679 4196 1689 4230
rect 1723 4196 1733 4230
rect 1679 4162 1733 4196
rect 1679 4128 1689 4162
rect 1723 4128 1733 4162
rect 1679 4112 1733 4128
rect 1763 4162 1817 4242
rect 1763 4128 1773 4162
rect 1807 4128 1817 4162
rect 1763 4112 1817 4128
rect 1847 4230 1901 4242
rect 1847 4196 1857 4230
rect 1891 4196 1901 4230
rect 1847 4162 1901 4196
rect 1847 4128 1857 4162
rect 1891 4128 1901 4162
rect 1847 4112 1901 4128
rect 1931 4162 1985 4242
rect 1931 4128 1941 4162
rect 1975 4128 1985 4162
rect 1931 4112 1985 4128
rect 2015 4230 2069 4242
rect 2015 4196 2025 4230
rect 2059 4196 2069 4230
rect 2015 4162 2069 4196
rect 2015 4128 2025 4162
rect 2059 4128 2069 4162
rect 2015 4112 2069 4128
rect 2099 4162 2153 4242
rect 2099 4128 2109 4162
rect 2143 4128 2153 4162
rect 2099 4112 2153 4128
rect 2183 4230 2237 4242
rect 2183 4196 2193 4230
rect 2227 4196 2237 4230
rect 2183 4162 2237 4196
rect 2183 4128 2193 4162
rect 2227 4128 2237 4162
rect 2183 4112 2237 4128
rect 2267 4162 2321 4242
rect 2267 4128 2277 4162
rect 2311 4128 2321 4162
rect 2267 4112 2321 4128
rect 2351 4230 2405 4242
rect 2351 4196 2361 4230
rect 2395 4196 2405 4230
rect 2351 4162 2405 4196
rect 2351 4128 2361 4162
rect 2395 4128 2405 4162
rect 2351 4112 2405 4128
rect 2435 4162 2489 4242
rect 2435 4128 2445 4162
rect 2479 4128 2489 4162
rect 2435 4112 2489 4128
rect 2519 4230 2573 4242
rect 2519 4196 2529 4230
rect 2563 4196 2573 4230
rect 2519 4162 2573 4196
rect 2519 4128 2529 4162
rect 2563 4128 2573 4162
rect 2519 4112 2573 4128
rect 2603 4162 2657 4242
rect 2603 4128 2613 4162
rect 2647 4128 2657 4162
rect 2603 4112 2657 4128
rect 2687 4230 2741 4242
rect 2687 4196 2697 4230
rect 2731 4196 2741 4230
rect 2687 4162 2741 4196
rect 2687 4128 2697 4162
rect 2731 4128 2741 4162
rect 2687 4112 2741 4128
rect 2771 4162 2825 4242
rect 2771 4128 2781 4162
rect 2815 4128 2825 4162
rect 2771 4112 2825 4128
rect 2855 4230 2909 4242
rect 2855 4196 2865 4230
rect 2899 4196 2909 4230
rect 2855 4162 2909 4196
rect 2855 4128 2865 4162
rect 2899 4128 2909 4162
rect 2855 4112 2909 4128
rect 2939 4162 2993 4242
rect 2939 4128 2949 4162
rect 2983 4128 2993 4162
rect 2939 4112 2993 4128
rect 3023 4230 3077 4242
rect 3023 4196 3033 4230
rect 3067 4196 3077 4230
rect 3023 4162 3077 4196
rect 3023 4128 3033 4162
rect 3067 4128 3077 4162
rect 3023 4112 3077 4128
rect 3107 4162 3161 4242
rect 3107 4128 3117 4162
rect 3151 4128 3161 4162
rect 3107 4112 3161 4128
rect 3191 4230 3245 4242
rect 3191 4196 3201 4230
rect 3235 4196 3245 4230
rect 3191 4162 3245 4196
rect 3191 4128 3201 4162
rect 3235 4128 3245 4162
rect 3191 4112 3245 4128
rect 3275 4162 3327 4242
rect 3275 4128 3285 4162
rect 3319 4128 3327 4162
rect 3275 4112 3327 4128
rect 3453 4194 3505 4242
rect 3453 4160 3461 4194
rect 3495 4160 3505 4194
rect 3453 4112 3505 4160
rect 3535 4196 3585 4242
rect 3535 4158 3600 4196
rect 3535 4124 3545 4158
rect 3579 4124 3600 4158
rect 3535 4112 3600 4124
rect 3630 4184 3682 4196
rect 3630 4150 3640 4184
rect 3674 4150 3682 4184
rect 3630 4112 3682 4150
rect 3736 4192 3788 4242
rect 3736 4158 3744 4192
rect 3778 4158 3788 4192
rect 3736 4112 3788 4158
rect 3818 4196 3868 4242
rect 3818 4158 3883 4196
rect 3818 4124 3828 4158
rect 3862 4124 3883 4158
rect 3818 4112 3883 4124
rect 3913 4168 3965 4196
rect 3913 4134 3923 4168
rect 3957 4134 3965 4168
rect 3913 4112 3965 4134
rect 4019 4166 4071 4240
rect 4019 4132 4027 4166
rect 4061 4132 4071 4166
rect 4019 4112 4071 4132
rect 4101 4218 4155 4240
rect 4101 4184 4111 4218
rect 4145 4184 4155 4218
rect 4101 4112 4155 4184
rect 4185 4196 4235 4240
rect 4185 4174 4273 4196
rect 4185 4140 4211 4174
rect 4245 4140 4273 4174
rect 4185 4112 4273 4140
rect 4303 4154 4359 4196
rect 4303 4120 4313 4154
rect 4347 4120 4359 4154
rect 4303 4112 4359 4120
rect 4389 4184 4439 4196
rect 4608 4184 4658 4240
rect 4389 4112 4454 4184
rect 4484 4158 4563 4184
rect 4484 4124 4504 4158
rect 4538 4124 4563 4158
rect 4484 4112 4563 4124
rect 4593 4112 4658 4184
rect 4688 4158 4740 4240
rect 4688 4124 4698 4158
rect 4732 4124 4740 4158
rect 4688 4112 4740 4124
rect 4794 4192 4846 4240
rect 4794 4158 4802 4192
rect 4836 4158 4846 4192
rect 4794 4112 4846 4158
rect 4876 4218 4930 4240
rect 4876 4184 4886 4218
rect 4920 4184 4930 4218
rect 4876 4112 4930 4184
rect 4960 4196 5010 4240
rect 4960 4174 5030 4196
rect 4960 4140 4986 4174
rect 5020 4140 5030 4174
rect 4960 4112 5030 4140
rect 5060 4154 5140 4196
rect 5060 4120 5070 4154
rect 5104 4120 5140 4154
rect 5060 4112 5140 4120
rect 5170 4184 5221 4196
rect 5387 4184 5437 4196
rect 5170 4112 5236 4184
rect 5266 4158 5342 4184
rect 5266 4124 5287 4158
rect 5321 4124 5342 4158
rect 5266 4112 5342 4124
rect 5372 4176 5437 4184
rect 5372 4142 5393 4176
rect 5427 4142 5437 4176
rect 5372 4112 5437 4142
rect 5467 4158 5519 4196
rect 5467 4124 5477 4158
rect 5511 4124 5519 4158
rect 5467 4112 5519 4124
rect 5573 4184 5625 4196
rect 5573 4150 5581 4184
rect 5615 4150 5625 4184
rect 5573 4112 5625 4150
rect 5655 4158 5709 4196
rect 5655 4124 5665 4158
rect 5699 4124 5709 4158
rect 5655 4112 5709 4124
rect 5739 4184 5791 4196
rect 5739 4150 5749 4184
rect 5783 4150 5791 4184
rect 5739 4112 5791 4150
rect 5845 4194 5897 4242
rect 5845 4160 5853 4194
rect 5887 4160 5897 4194
rect 5845 4112 5897 4160
rect 5927 4196 5977 4242
rect 5927 4158 5992 4196
rect 5927 4124 5937 4158
rect 5971 4124 5992 4158
rect 5927 4112 5992 4124
rect 6022 4184 6074 4196
rect 6022 4150 6032 4184
rect 6066 4150 6074 4184
rect 6022 4112 6074 4150
rect 6128 4192 6180 4242
rect 6128 4158 6136 4192
rect 6170 4158 6180 4192
rect 6128 4112 6180 4158
rect 6210 4196 6260 4242
rect 6210 4158 6275 4196
rect 6210 4124 6220 4158
rect 6254 4124 6275 4158
rect 6210 4112 6275 4124
rect 6305 4168 6357 4196
rect 6305 4134 6315 4168
rect 6349 4134 6357 4168
rect 6305 4112 6357 4134
rect 6411 4166 6463 4240
rect 6411 4132 6419 4166
rect 6453 4132 6463 4166
rect 6411 4112 6463 4132
rect 6493 4218 6547 4240
rect 6493 4184 6503 4218
rect 6537 4184 6547 4218
rect 6493 4112 6547 4184
rect 6577 4196 6627 4240
rect 6577 4174 6665 4196
rect 6577 4140 6603 4174
rect 6637 4140 6665 4174
rect 6577 4112 6665 4140
rect 6695 4154 6751 4196
rect 6695 4120 6705 4154
rect 6739 4120 6751 4154
rect 6695 4112 6751 4120
rect 6781 4184 6831 4196
rect 7000 4184 7050 4240
rect 6781 4112 6846 4184
rect 6876 4158 6955 4184
rect 6876 4124 6896 4158
rect 6930 4124 6955 4158
rect 6876 4112 6955 4124
rect 6985 4112 7050 4184
rect 7080 4158 7132 4240
rect 7080 4124 7090 4158
rect 7124 4124 7132 4158
rect 7080 4112 7132 4124
rect 7186 4192 7238 4240
rect 7186 4158 7194 4192
rect 7228 4158 7238 4192
rect 7186 4112 7238 4158
rect 7268 4218 7322 4240
rect 7268 4184 7278 4218
rect 7312 4184 7322 4218
rect 7268 4112 7322 4184
rect 7352 4196 7402 4240
rect 7352 4174 7422 4196
rect 7352 4140 7378 4174
rect 7412 4140 7422 4174
rect 7352 4112 7422 4140
rect 7452 4154 7532 4196
rect 7452 4120 7462 4154
rect 7496 4120 7532 4154
rect 7452 4112 7532 4120
rect 7562 4184 7613 4196
rect 7779 4184 7829 4196
rect 7562 4112 7628 4184
rect 7658 4158 7734 4184
rect 7658 4124 7679 4158
rect 7713 4124 7734 4158
rect 7658 4112 7734 4124
rect 7764 4176 7829 4184
rect 7764 4142 7785 4176
rect 7819 4142 7829 4176
rect 7764 4112 7829 4142
rect 7859 4158 7911 4196
rect 7859 4124 7869 4158
rect 7903 4124 7911 4158
rect 7859 4112 7911 4124
rect 7965 4184 8017 4196
rect 7965 4150 7973 4184
rect 8007 4150 8017 4184
rect 7965 4112 8017 4150
rect 8047 4158 8101 4196
rect 8047 4124 8057 4158
rect 8091 4124 8101 4158
rect 8047 4112 8101 4124
rect 8131 4184 8183 4196
rect 8131 4150 8141 4184
rect 8175 4150 8183 4184
rect 8131 4112 8183 4150
rect 8237 4194 8289 4242
rect 8237 4160 8245 4194
rect 8279 4160 8289 4194
rect 8237 4112 8289 4160
rect 8319 4196 8369 4242
rect 8319 4158 8384 4196
rect 8319 4124 8329 4158
rect 8363 4124 8384 4158
rect 8319 4112 8384 4124
rect 8414 4184 8466 4196
rect 8414 4150 8424 4184
rect 8458 4150 8466 4184
rect 8414 4112 8466 4150
rect 8520 4192 8572 4242
rect 8520 4158 8528 4192
rect 8562 4158 8572 4192
rect 8520 4112 8572 4158
rect 8602 4196 8652 4242
rect 8602 4158 8667 4196
rect 8602 4124 8612 4158
rect 8646 4124 8667 4158
rect 8602 4112 8667 4124
rect 8697 4168 8749 4196
rect 8697 4134 8707 4168
rect 8741 4134 8749 4168
rect 8697 4112 8749 4134
rect 8803 4166 8855 4240
rect 8803 4132 8811 4166
rect 8845 4132 8855 4166
rect 8803 4112 8855 4132
rect 8885 4218 8939 4240
rect 8885 4184 8895 4218
rect 8929 4184 8939 4218
rect 8885 4112 8939 4184
rect 8969 4196 9019 4240
rect 8969 4174 9057 4196
rect 8969 4140 8995 4174
rect 9029 4140 9057 4174
rect 8969 4112 9057 4140
rect 9087 4154 9143 4196
rect 9087 4120 9097 4154
rect 9131 4120 9143 4154
rect 9087 4112 9143 4120
rect 9173 4184 9223 4196
rect 9392 4184 9442 4240
rect 9173 4112 9238 4184
rect 9268 4158 9347 4184
rect 9268 4124 9288 4158
rect 9322 4124 9347 4158
rect 9268 4112 9347 4124
rect 9377 4112 9442 4184
rect 9472 4158 9524 4240
rect 9472 4124 9482 4158
rect 9516 4124 9524 4158
rect 9472 4112 9524 4124
rect 9578 4192 9630 4240
rect 9578 4158 9586 4192
rect 9620 4158 9630 4192
rect 9578 4112 9630 4158
rect 9660 4218 9714 4240
rect 9660 4184 9670 4218
rect 9704 4184 9714 4218
rect 9660 4112 9714 4184
rect 9744 4196 9794 4240
rect 9744 4174 9814 4196
rect 9744 4140 9770 4174
rect 9804 4140 9814 4174
rect 9744 4112 9814 4140
rect 9844 4154 9924 4196
rect 9844 4120 9854 4154
rect 9888 4120 9924 4154
rect 9844 4112 9924 4120
rect 9954 4184 10005 4196
rect 10171 4184 10221 4196
rect 9954 4112 10020 4184
rect 10050 4158 10126 4184
rect 10050 4124 10071 4158
rect 10105 4124 10126 4158
rect 10050 4112 10126 4124
rect 10156 4176 10221 4184
rect 10156 4142 10177 4176
rect 10211 4142 10221 4176
rect 10156 4112 10221 4142
rect 10251 4158 10303 4196
rect 10251 4124 10261 4158
rect 10295 4124 10303 4158
rect 10251 4112 10303 4124
rect 10357 4184 10409 4196
rect 10357 4150 10365 4184
rect 10399 4150 10409 4184
rect 10357 4112 10409 4150
rect 10439 4158 10493 4196
rect 10439 4124 10449 4158
rect 10483 4124 10493 4158
rect 10439 4112 10493 4124
rect 10523 4184 10575 4196
rect 10523 4150 10533 4184
rect 10567 4150 10575 4184
rect 10523 4112 10575 4150
rect 10629 4194 10681 4242
rect 10629 4160 10637 4194
rect 10671 4160 10681 4194
rect 10629 4112 10681 4160
rect 10711 4196 10761 4242
rect 10711 4158 10776 4196
rect 10711 4124 10721 4158
rect 10755 4124 10776 4158
rect 10711 4112 10776 4124
rect 10806 4184 10858 4196
rect 10806 4150 10816 4184
rect 10850 4150 10858 4184
rect 10806 4112 10858 4150
rect 10912 4192 10964 4242
rect 10912 4158 10920 4192
rect 10954 4158 10964 4192
rect 10912 4112 10964 4158
rect 10994 4196 11044 4242
rect 10994 4158 11059 4196
rect 10994 4124 11004 4158
rect 11038 4124 11059 4158
rect 10994 4112 11059 4124
rect 11089 4168 11141 4196
rect 11089 4134 11099 4168
rect 11133 4134 11141 4168
rect 11089 4112 11141 4134
rect 11195 4166 11247 4240
rect 11195 4132 11203 4166
rect 11237 4132 11247 4166
rect 11195 4112 11247 4132
rect 11277 4218 11331 4240
rect 11277 4184 11287 4218
rect 11321 4184 11331 4218
rect 11277 4112 11331 4184
rect 11361 4196 11411 4240
rect 11361 4174 11449 4196
rect 11361 4140 11387 4174
rect 11421 4140 11449 4174
rect 11361 4112 11449 4140
rect 11479 4154 11535 4196
rect 11479 4120 11489 4154
rect 11523 4120 11535 4154
rect 11479 4112 11535 4120
rect 11565 4184 11615 4196
rect 11784 4184 11834 4240
rect 11565 4112 11630 4184
rect 11660 4158 11739 4184
rect 11660 4124 11680 4158
rect 11714 4124 11739 4158
rect 11660 4112 11739 4124
rect 11769 4112 11834 4184
rect 11864 4158 11916 4240
rect 11864 4124 11874 4158
rect 11908 4124 11916 4158
rect 11864 4112 11916 4124
rect 11970 4192 12022 4240
rect 11970 4158 11978 4192
rect 12012 4158 12022 4192
rect 11970 4112 12022 4158
rect 12052 4218 12106 4240
rect 12052 4184 12062 4218
rect 12096 4184 12106 4218
rect 12052 4112 12106 4184
rect 12136 4196 12186 4240
rect 12136 4174 12206 4196
rect 12136 4140 12162 4174
rect 12196 4140 12206 4174
rect 12136 4112 12206 4140
rect 12236 4154 12316 4196
rect 12236 4120 12246 4154
rect 12280 4120 12316 4154
rect 12236 4112 12316 4120
rect 12346 4184 12397 4196
rect 12563 4184 12613 4196
rect 12346 4112 12412 4184
rect 12442 4158 12518 4184
rect 12442 4124 12463 4158
rect 12497 4124 12518 4158
rect 12442 4112 12518 4124
rect 12548 4176 12613 4184
rect 12548 4142 12569 4176
rect 12603 4142 12613 4176
rect 12548 4112 12613 4142
rect 12643 4158 12695 4196
rect 12643 4124 12653 4158
rect 12687 4124 12695 4158
rect 12643 4112 12695 4124
rect 12749 4184 12801 4196
rect 12749 4150 12757 4184
rect 12791 4150 12801 4184
rect 12749 4112 12801 4150
rect 12831 4158 12885 4196
rect 12831 4124 12841 4158
rect 12875 4124 12885 4158
rect 12831 4112 12885 4124
rect 12915 4184 12967 4196
rect 12915 4150 12925 4184
rect 12959 4150 12967 4184
rect 12915 4112 12967 4150
rect 653 3297 705 3342
rect 653 3263 661 3297
rect 695 3263 705 3297
rect 653 3238 705 3263
rect 735 3284 793 3342
rect 735 3250 747 3284
rect 781 3250 793 3284
rect 735 3238 793 3250
rect 823 3314 875 3342
rect 823 3280 833 3314
rect 867 3280 875 3314
rect 823 3238 875 3280
rect 929 3320 981 3368
rect 929 3286 937 3320
rect 971 3286 981 3320
rect 929 3238 981 3286
rect 1011 3288 1065 3368
rect 1011 3254 1021 3288
rect 1055 3254 1065 3288
rect 1011 3238 1065 3254
rect 1095 3320 1149 3368
rect 1095 3286 1105 3320
rect 1139 3286 1149 3320
rect 1095 3238 1149 3286
rect 1179 3288 1233 3368
rect 1179 3254 1189 3288
rect 1223 3254 1233 3288
rect 1179 3238 1233 3254
rect 1263 3320 1317 3368
rect 1263 3286 1273 3320
rect 1307 3286 1317 3320
rect 1263 3238 1317 3286
rect 1347 3352 1399 3368
rect 1347 3318 1357 3352
rect 1391 3318 1399 3352
rect 1347 3284 1399 3318
rect 1347 3250 1357 3284
rect 1391 3250 1399 3284
rect 1347 3238 1399 3250
rect 3236 3357 3288 3369
rect 3236 3323 3244 3357
rect 3278 3323 3288 3357
rect 3236 3289 3288 3323
rect 3236 3255 3244 3289
rect 3278 3255 3288 3289
rect 3236 3239 3288 3255
rect 3318 3357 3370 3369
rect 3318 3323 3328 3357
rect 3362 3323 3370 3357
rect 3318 3289 3370 3323
rect 3318 3255 3328 3289
rect 3362 3255 3370 3289
rect 3318 3239 3370 3255
rect 3452 3311 3504 3323
rect 3452 3277 3460 3311
rect 3494 3277 3504 3311
rect 3452 3239 3504 3277
rect 3534 3285 3588 3323
rect 3534 3251 3544 3285
rect 3578 3251 3588 3285
rect 3534 3239 3588 3251
rect 3618 3311 3670 3323
rect 3618 3277 3628 3311
rect 3662 3277 3670 3311
rect 3618 3239 3670 3277
rect 3724 3285 3776 3323
rect 3724 3251 3732 3285
rect 3766 3251 3776 3285
rect 3724 3239 3776 3251
rect 3806 3311 3856 3323
rect 4233 3323 4283 3367
rect 4022 3311 4073 3323
rect 3806 3303 3871 3311
rect 3806 3269 3816 3303
rect 3850 3269 3871 3303
rect 3806 3239 3871 3269
rect 3901 3285 3977 3311
rect 3901 3251 3922 3285
rect 3956 3251 3977 3285
rect 3901 3239 3977 3251
rect 4007 3239 4073 3311
rect 4103 3281 4183 3323
rect 4103 3247 4139 3281
rect 4173 3247 4183 3281
rect 4103 3239 4183 3247
rect 4213 3301 4283 3323
rect 4213 3267 4223 3301
rect 4257 3267 4283 3301
rect 4213 3239 4283 3267
rect 4313 3345 4367 3367
rect 4313 3311 4323 3345
rect 4357 3311 4367 3345
rect 4313 3239 4367 3311
rect 4397 3319 4449 3367
rect 4397 3285 4407 3319
rect 4441 3285 4449 3319
rect 4397 3239 4449 3285
rect 4503 3285 4555 3367
rect 4503 3251 4511 3285
rect 4545 3251 4555 3285
rect 4503 3239 4555 3251
rect 4585 3311 4635 3367
rect 5008 3323 5058 3367
rect 4804 3311 4854 3323
rect 4585 3239 4650 3311
rect 4680 3285 4759 3311
rect 4680 3251 4705 3285
rect 4739 3251 4759 3285
rect 4680 3239 4759 3251
rect 4789 3239 4854 3311
rect 4884 3281 4940 3323
rect 4884 3247 4896 3281
rect 4930 3247 4940 3281
rect 4884 3239 4940 3247
rect 4970 3301 5058 3323
rect 4970 3267 4998 3301
rect 5032 3267 5058 3301
rect 4970 3239 5058 3267
rect 5088 3345 5142 3367
rect 5088 3311 5098 3345
rect 5132 3311 5142 3345
rect 5088 3239 5142 3311
rect 5172 3293 5224 3367
rect 5375 3323 5425 3369
rect 5172 3259 5182 3293
rect 5216 3259 5224 3293
rect 5172 3239 5224 3259
rect 5278 3295 5330 3323
rect 5278 3261 5286 3295
rect 5320 3261 5330 3295
rect 5278 3239 5330 3261
rect 5360 3285 5425 3323
rect 5360 3251 5381 3285
rect 5415 3251 5425 3285
rect 5360 3239 5425 3251
rect 5455 3319 5507 3369
rect 5658 3323 5708 3369
rect 5455 3285 5465 3319
rect 5499 3285 5507 3319
rect 5455 3239 5507 3285
rect 5561 3311 5613 3323
rect 5561 3277 5569 3311
rect 5603 3277 5613 3311
rect 5561 3239 5613 3277
rect 5643 3285 5708 3323
rect 5643 3251 5664 3285
rect 5698 3251 5708 3285
rect 5643 3239 5708 3251
rect 5738 3321 5790 3369
rect 5738 3287 5748 3321
rect 5782 3287 5790 3321
rect 5738 3239 5790 3287
rect 5844 3311 5896 3323
rect 5844 3277 5852 3311
rect 5886 3277 5896 3311
rect 5844 3239 5896 3277
rect 5926 3285 5980 3323
rect 5926 3251 5936 3285
rect 5970 3251 5980 3285
rect 5926 3239 5980 3251
rect 6010 3311 6062 3323
rect 6010 3277 6020 3311
rect 6054 3277 6062 3311
rect 6010 3239 6062 3277
rect 6116 3285 6168 3323
rect 6116 3251 6124 3285
rect 6158 3251 6168 3285
rect 6116 3239 6168 3251
rect 6198 3311 6248 3323
rect 6625 3323 6675 3367
rect 6414 3311 6465 3323
rect 6198 3303 6263 3311
rect 6198 3269 6208 3303
rect 6242 3269 6263 3303
rect 6198 3239 6263 3269
rect 6293 3285 6369 3311
rect 6293 3251 6314 3285
rect 6348 3251 6369 3285
rect 6293 3239 6369 3251
rect 6399 3239 6465 3311
rect 6495 3281 6575 3323
rect 6495 3247 6531 3281
rect 6565 3247 6575 3281
rect 6495 3239 6575 3247
rect 6605 3301 6675 3323
rect 6605 3267 6615 3301
rect 6649 3267 6675 3301
rect 6605 3239 6675 3267
rect 6705 3345 6759 3367
rect 6705 3311 6715 3345
rect 6749 3311 6759 3345
rect 6705 3239 6759 3311
rect 6789 3319 6841 3367
rect 6789 3285 6799 3319
rect 6833 3285 6841 3319
rect 6789 3239 6841 3285
rect 6895 3285 6947 3367
rect 6895 3251 6903 3285
rect 6937 3251 6947 3285
rect 6895 3239 6947 3251
rect 6977 3311 7027 3367
rect 7400 3323 7450 3367
rect 7196 3311 7246 3323
rect 6977 3239 7042 3311
rect 7072 3285 7151 3311
rect 7072 3251 7097 3285
rect 7131 3251 7151 3285
rect 7072 3239 7151 3251
rect 7181 3239 7246 3311
rect 7276 3281 7332 3323
rect 7276 3247 7288 3281
rect 7322 3247 7332 3281
rect 7276 3239 7332 3247
rect 7362 3301 7450 3323
rect 7362 3267 7390 3301
rect 7424 3267 7450 3301
rect 7362 3239 7450 3267
rect 7480 3345 7534 3367
rect 7480 3311 7490 3345
rect 7524 3311 7534 3345
rect 7480 3239 7534 3311
rect 7564 3293 7616 3367
rect 7767 3323 7817 3369
rect 7564 3259 7574 3293
rect 7608 3259 7616 3293
rect 7564 3239 7616 3259
rect 7670 3295 7722 3323
rect 7670 3261 7678 3295
rect 7712 3261 7722 3295
rect 7670 3239 7722 3261
rect 7752 3285 7817 3323
rect 7752 3251 7773 3285
rect 7807 3251 7817 3285
rect 7752 3239 7817 3251
rect 7847 3319 7899 3369
rect 8050 3323 8100 3369
rect 7847 3285 7857 3319
rect 7891 3285 7899 3319
rect 7847 3239 7899 3285
rect 7953 3311 8005 3323
rect 7953 3277 7961 3311
rect 7995 3277 8005 3311
rect 7953 3239 8005 3277
rect 8035 3285 8100 3323
rect 8035 3251 8056 3285
rect 8090 3251 8100 3285
rect 8035 3239 8100 3251
rect 8130 3321 8182 3369
rect 8130 3287 8140 3321
rect 8174 3287 8182 3321
rect 8130 3239 8182 3287
rect 8236 3311 8288 3323
rect 8236 3277 8244 3311
rect 8278 3277 8288 3311
rect 8236 3239 8288 3277
rect 8318 3285 8372 3323
rect 8318 3251 8328 3285
rect 8362 3251 8372 3285
rect 8318 3239 8372 3251
rect 8402 3311 8454 3323
rect 8402 3277 8412 3311
rect 8446 3277 8454 3311
rect 8402 3239 8454 3277
rect 8508 3285 8560 3323
rect 8508 3251 8516 3285
rect 8550 3251 8560 3285
rect 8508 3239 8560 3251
rect 8590 3311 8640 3323
rect 9017 3323 9067 3367
rect 8806 3311 8857 3323
rect 8590 3303 8655 3311
rect 8590 3269 8600 3303
rect 8634 3269 8655 3303
rect 8590 3239 8655 3269
rect 8685 3285 8761 3311
rect 8685 3251 8706 3285
rect 8740 3251 8761 3285
rect 8685 3239 8761 3251
rect 8791 3239 8857 3311
rect 8887 3281 8967 3323
rect 8887 3247 8923 3281
rect 8957 3247 8967 3281
rect 8887 3239 8967 3247
rect 8997 3301 9067 3323
rect 8997 3267 9007 3301
rect 9041 3267 9067 3301
rect 8997 3239 9067 3267
rect 9097 3345 9151 3367
rect 9097 3311 9107 3345
rect 9141 3311 9151 3345
rect 9097 3239 9151 3311
rect 9181 3319 9233 3367
rect 9181 3285 9191 3319
rect 9225 3285 9233 3319
rect 9181 3239 9233 3285
rect 9287 3285 9339 3367
rect 9287 3251 9295 3285
rect 9329 3251 9339 3285
rect 9287 3239 9339 3251
rect 9369 3311 9419 3367
rect 9792 3323 9842 3367
rect 9588 3311 9638 3323
rect 9369 3239 9434 3311
rect 9464 3285 9543 3311
rect 9464 3251 9489 3285
rect 9523 3251 9543 3285
rect 9464 3239 9543 3251
rect 9573 3239 9638 3311
rect 9668 3281 9724 3323
rect 9668 3247 9680 3281
rect 9714 3247 9724 3281
rect 9668 3239 9724 3247
rect 9754 3301 9842 3323
rect 9754 3267 9782 3301
rect 9816 3267 9842 3301
rect 9754 3239 9842 3267
rect 9872 3345 9926 3367
rect 9872 3311 9882 3345
rect 9916 3311 9926 3345
rect 9872 3239 9926 3311
rect 9956 3293 10008 3367
rect 10159 3323 10209 3369
rect 9956 3259 9966 3293
rect 10000 3259 10008 3293
rect 9956 3239 10008 3259
rect 10062 3295 10114 3323
rect 10062 3261 10070 3295
rect 10104 3261 10114 3295
rect 10062 3239 10114 3261
rect 10144 3285 10209 3323
rect 10144 3251 10165 3285
rect 10199 3251 10209 3285
rect 10144 3239 10209 3251
rect 10239 3319 10291 3369
rect 10442 3323 10492 3369
rect 10239 3285 10249 3319
rect 10283 3285 10291 3319
rect 10239 3239 10291 3285
rect 10345 3311 10397 3323
rect 10345 3277 10353 3311
rect 10387 3277 10397 3311
rect 10345 3239 10397 3277
rect 10427 3285 10492 3323
rect 10427 3251 10448 3285
rect 10482 3251 10492 3285
rect 10427 3239 10492 3251
rect 10522 3321 10574 3369
rect 10522 3287 10532 3321
rect 10566 3287 10574 3321
rect 10522 3239 10574 3287
rect 10628 3311 10680 3323
rect 10628 3277 10636 3311
rect 10670 3277 10680 3311
rect 10628 3239 10680 3277
rect 10710 3285 10764 3323
rect 10710 3251 10720 3285
rect 10754 3251 10764 3285
rect 10710 3239 10764 3251
rect 10794 3311 10846 3323
rect 10794 3277 10804 3311
rect 10838 3277 10846 3311
rect 10794 3239 10846 3277
rect 10900 3285 10952 3323
rect 10900 3251 10908 3285
rect 10942 3251 10952 3285
rect 10900 3239 10952 3251
rect 10982 3311 11032 3323
rect 11409 3323 11459 3367
rect 11198 3311 11249 3323
rect 10982 3303 11047 3311
rect 10982 3269 10992 3303
rect 11026 3269 11047 3303
rect 10982 3239 11047 3269
rect 11077 3285 11153 3311
rect 11077 3251 11098 3285
rect 11132 3251 11153 3285
rect 11077 3239 11153 3251
rect 11183 3239 11249 3311
rect 11279 3281 11359 3323
rect 11279 3247 11315 3281
rect 11349 3247 11359 3281
rect 11279 3239 11359 3247
rect 11389 3301 11459 3323
rect 11389 3267 11399 3301
rect 11433 3267 11459 3301
rect 11389 3239 11459 3267
rect 11489 3345 11543 3367
rect 11489 3311 11499 3345
rect 11533 3311 11543 3345
rect 11489 3239 11543 3311
rect 11573 3319 11625 3367
rect 11573 3285 11583 3319
rect 11617 3285 11625 3319
rect 11573 3239 11625 3285
rect 11679 3285 11731 3367
rect 11679 3251 11687 3285
rect 11721 3251 11731 3285
rect 11679 3239 11731 3251
rect 11761 3311 11811 3367
rect 12184 3323 12234 3367
rect 11980 3311 12030 3323
rect 11761 3239 11826 3311
rect 11856 3285 11935 3311
rect 11856 3251 11881 3285
rect 11915 3251 11935 3285
rect 11856 3239 11935 3251
rect 11965 3239 12030 3311
rect 12060 3281 12116 3323
rect 12060 3247 12072 3281
rect 12106 3247 12116 3281
rect 12060 3239 12116 3247
rect 12146 3301 12234 3323
rect 12146 3267 12174 3301
rect 12208 3267 12234 3301
rect 12146 3239 12234 3267
rect 12264 3345 12318 3367
rect 12264 3311 12274 3345
rect 12308 3311 12318 3345
rect 12264 3239 12318 3311
rect 12348 3293 12400 3367
rect 12551 3323 12601 3369
rect 12348 3259 12358 3293
rect 12392 3259 12400 3293
rect 12348 3239 12400 3259
rect 12454 3295 12506 3323
rect 12454 3261 12462 3295
rect 12496 3261 12506 3295
rect 12454 3239 12506 3261
rect 12536 3285 12601 3323
rect 12536 3251 12557 3285
rect 12591 3251 12601 3285
rect 12536 3239 12601 3251
rect 12631 3319 12683 3369
rect 12834 3323 12884 3369
rect 12631 3285 12641 3319
rect 12675 3285 12683 3319
rect 12631 3239 12683 3285
rect 12737 3311 12789 3323
rect 12737 3277 12745 3311
rect 12779 3277 12789 3311
rect 12737 3239 12789 3277
rect 12819 3285 12884 3323
rect 12819 3251 12840 3285
rect 12874 3251 12884 3285
rect 12819 3239 12884 3251
rect 12914 3321 12966 3369
rect 12914 3287 12924 3321
rect 12958 3287 12966 3321
rect 12914 3239 12966 3287
rect 1060 2448 1112 2496
rect 1060 2414 1068 2448
rect 1102 2414 1112 2448
rect 1060 2366 1112 2414
rect 1142 2450 1192 2496
rect 1142 2412 1207 2450
rect 1142 2378 1152 2412
rect 1186 2378 1207 2412
rect 1142 2366 1207 2378
rect 1237 2438 1289 2450
rect 1237 2404 1247 2438
rect 1281 2404 1289 2438
rect 1237 2366 1289 2404
rect 1343 2446 1395 2496
rect 1343 2412 1351 2446
rect 1385 2412 1395 2446
rect 1343 2366 1395 2412
rect 1425 2450 1475 2496
rect 1425 2412 1490 2450
rect 1425 2378 1435 2412
rect 1469 2378 1490 2412
rect 1425 2366 1490 2378
rect 1520 2422 1572 2450
rect 1520 2388 1530 2422
rect 1564 2388 1572 2422
rect 1520 2366 1572 2388
rect 1626 2420 1678 2494
rect 1626 2386 1634 2420
rect 1668 2386 1678 2420
rect 1626 2366 1678 2386
rect 1708 2472 1762 2494
rect 1708 2438 1718 2472
rect 1752 2438 1762 2472
rect 1708 2366 1762 2438
rect 1792 2450 1842 2494
rect 1792 2428 1880 2450
rect 1792 2394 1818 2428
rect 1852 2394 1880 2428
rect 1792 2366 1880 2394
rect 1910 2408 1966 2450
rect 1910 2374 1920 2408
rect 1954 2374 1966 2408
rect 1910 2366 1966 2374
rect 1996 2438 2046 2450
rect 2215 2438 2265 2494
rect 1996 2366 2061 2438
rect 2091 2412 2170 2438
rect 2091 2378 2111 2412
rect 2145 2378 2170 2412
rect 2091 2366 2170 2378
rect 2200 2366 2265 2438
rect 2295 2412 2347 2494
rect 2295 2378 2305 2412
rect 2339 2378 2347 2412
rect 2295 2366 2347 2378
rect 2401 2446 2453 2494
rect 2401 2412 2409 2446
rect 2443 2412 2453 2446
rect 2401 2366 2453 2412
rect 2483 2472 2537 2494
rect 2483 2438 2493 2472
rect 2527 2438 2537 2472
rect 2483 2366 2537 2438
rect 2567 2450 2617 2494
rect 2567 2428 2637 2450
rect 2567 2394 2593 2428
rect 2627 2394 2637 2428
rect 2567 2366 2637 2394
rect 2667 2408 2747 2450
rect 2667 2374 2677 2408
rect 2711 2374 2747 2408
rect 2667 2366 2747 2374
rect 2777 2438 2828 2450
rect 2994 2438 3044 2450
rect 2777 2366 2843 2438
rect 2873 2412 2949 2438
rect 2873 2378 2894 2412
rect 2928 2378 2949 2412
rect 2873 2366 2949 2378
rect 2979 2430 3044 2438
rect 2979 2396 3000 2430
rect 3034 2396 3044 2430
rect 2979 2366 3044 2396
rect 3074 2412 3126 2450
rect 3074 2378 3084 2412
rect 3118 2378 3126 2412
rect 3074 2366 3126 2378
rect 3180 2438 3232 2450
rect 3180 2404 3188 2438
rect 3222 2404 3232 2438
rect 3180 2366 3232 2404
rect 3262 2412 3316 2450
rect 3262 2378 3272 2412
rect 3306 2378 3316 2412
rect 3262 2366 3316 2378
rect 3346 2438 3398 2450
rect 3346 2404 3356 2438
rect 3390 2404 3398 2438
rect 3346 2366 3398 2404
rect 3452 2448 3504 2496
rect 3452 2414 3460 2448
rect 3494 2414 3504 2448
rect 3452 2366 3504 2414
rect 3534 2450 3584 2496
rect 3534 2412 3599 2450
rect 3534 2378 3544 2412
rect 3578 2378 3599 2412
rect 3534 2366 3599 2378
rect 3629 2438 3681 2450
rect 3629 2404 3639 2438
rect 3673 2404 3681 2438
rect 3629 2366 3681 2404
rect 3735 2446 3787 2496
rect 3735 2412 3743 2446
rect 3777 2412 3787 2446
rect 3735 2366 3787 2412
rect 3817 2450 3867 2496
rect 3817 2412 3882 2450
rect 3817 2378 3827 2412
rect 3861 2378 3882 2412
rect 3817 2366 3882 2378
rect 3912 2422 3964 2450
rect 3912 2388 3922 2422
rect 3956 2388 3964 2422
rect 3912 2366 3964 2388
rect 4018 2420 4070 2494
rect 4018 2386 4026 2420
rect 4060 2386 4070 2420
rect 4018 2366 4070 2386
rect 4100 2472 4154 2494
rect 4100 2438 4110 2472
rect 4144 2438 4154 2472
rect 4100 2366 4154 2438
rect 4184 2450 4234 2494
rect 4184 2428 4272 2450
rect 4184 2394 4210 2428
rect 4244 2394 4272 2428
rect 4184 2366 4272 2394
rect 4302 2408 4358 2450
rect 4302 2374 4312 2408
rect 4346 2374 4358 2408
rect 4302 2366 4358 2374
rect 4388 2438 4438 2450
rect 4607 2438 4657 2494
rect 4388 2366 4453 2438
rect 4483 2412 4562 2438
rect 4483 2378 4503 2412
rect 4537 2378 4562 2412
rect 4483 2366 4562 2378
rect 4592 2366 4657 2438
rect 4687 2412 4739 2494
rect 4687 2378 4697 2412
rect 4731 2378 4739 2412
rect 4687 2366 4739 2378
rect 4793 2446 4845 2494
rect 4793 2412 4801 2446
rect 4835 2412 4845 2446
rect 4793 2366 4845 2412
rect 4875 2472 4929 2494
rect 4875 2438 4885 2472
rect 4919 2438 4929 2472
rect 4875 2366 4929 2438
rect 4959 2450 5009 2494
rect 4959 2428 5029 2450
rect 4959 2394 4985 2428
rect 5019 2394 5029 2428
rect 4959 2366 5029 2394
rect 5059 2408 5139 2450
rect 5059 2374 5069 2408
rect 5103 2374 5139 2408
rect 5059 2366 5139 2374
rect 5169 2438 5220 2450
rect 5386 2438 5436 2450
rect 5169 2366 5235 2438
rect 5265 2412 5341 2438
rect 5265 2378 5286 2412
rect 5320 2378 5341 2412
rect 5265 2366 5341 2378
rect 5371 2430 5436 2438
rect 5371 2396 5392 2430
rect 5426 2396 5436 2430
rect 5371 2366 5436 2396
rect 5466 2412 5518 2450
rect 5466 2378 5476 2412
rect 5510 2378 5518 2412
rect 5466 2366 5518 2378
rect 5572 2438 5624 2450
rect 5572 2404 5580 2438
rect 5614 2404 5624 2438
rect 5572 2366 5624 2404
rect 5654 2412 5708 2450
rect 5654 2378 5664 2412
rect 5698 2378 5708 2412
rect 5654 2366 5708 2378
rect 5738 2438 5790 2450
rect 5738 2404 5748 2438
rect 5782 2404 5790 2438
rect 5738 2366 5790 2404
rect 5844 2448 5896 2496
rect 5844 2414 5852 2448
rect 5886 2414 5896 2448
rect 5844 2366 5896 2414
rect 5926 2450 5976 2496
rect 5926 2412 5991 2450
rect 5926 2378 5936 2412
rect 5970 2378 5991 2412
rect 5926 2366 5991 2378
rect 6021 2438 6073 2450
rect 6021 2404 6031 2438
rect 6065 2404 6073 2438
rect 6021 2366 6073 2404
rect 6127 2446 6179 2496
rect 6127 2412 6135 2446
rect 6169 2412 6179 2446
rect 6127 2366 6179 2412
rect 6209 2450 6259 2496
rect 6209 2412 6274 2450
rect 6209 2378 6219 2412
rect 6253 2378 6274 2412
rect 6209 2366 6274 2378
rect 6304 2422 6356 2450
rect 6304 2388 6314 2422
rect 6348 2388 6356 2422
rect 6304 2366 6356 2388
rect 6410 2420 6462 2494
rect 6410 2386 6418 2420
rect 6452 2386 6462 2420
rect 6410 2366 6462 2386
rect 6492 2472 6546 2494
rect 6492 2438 6502 2472
rect 6536 2438 6546 2472
rect 6492 2366 6546 2438
rect 6576 2450 6626 2494
rect 6576 2428 6664 2450
rect 6576 2394 6602 2428
rect 6636 2394 6664 2428
rect 6576 2366 6664 2394
rect 6694 2408 6750 2450
rect 6694 2374 6704 2408
rect 6738 2374 6750 2408
rect 6694 2366 6750 2374
rect 6780 2438 6830 2450
rect 6999 2438 7049 2494
rect 6780 2366 6845 2438
rect 6875 2412 6954 2438
rect 6875 2378 6895 2412
rect 6929 2378 6954 2412
rect 6875 2366 6954 2378
rect 6984 2366 7049 2438
rect 7079 2412 7131 2494
rect 7079 2378 7089 2412
rect 7123 2378 7131 2412
rect 7079 2366 7131 2378
rect 7185 2446 7237 2494
rect 7185 2412 7193 2446
rect 7227 2412 7237 2446
rect 7185 2366 7237 2412
rect 7267 2472 7321 2494
rect 7267 2438 7277 2472
rect 7311 2438 7321 2472
rect 7267 2366 7321 2438
rect 7351 2450 7401 2494
rect 7351 2428 7421 2450
rect 7351 2394 7377 2428
rect 7411 2394 7421 2428
rect 7351 2366 7421 2394
rect 7451 2408 7531 2450
rect 7451 2374 7461 2408
rect 7495 2374 7531 2408
rect 7451 2366 7531 2374
rect 7561 2438 7612 2450
rect 7778 2438 7828 2450
rect 7561 2366 7627 2438
rect 7657 2412 7733 2438
rect 7657 2378 7678 2412
rect 7712 2378 7733 2412
rect 7657 2366 7733 2378
rect 7763 2430 7828 2438
rect 7763 2396 7784 2430
rect 7818 2396 7828 2430
rect 7763 2366 7828 2396
rect 7858 2412 7910 2450
rect 7858 2378 7868 2412
rect 7902 2378 7910 2412
rect 7858 2366 7910 2378
rect 7964 2438 8016 2450
rect 7964 2404 7972 2438
rect 8006 2404 8016 2438
rect 7964 2366 8016 2404
rect 8046 2412 8100 2450
rect 8046 2378 8056 2412
rect 8090 2378 8100 2412
rect 8046 2366 8100 2378
rect 8130 2438 8182 2450
rect 8130 2404 8140 2438
rect 8174 2404 8182 2438
rect 8130 2366 8182 2404
rect 8236 2448 8288 2496
rect 8236 2414 8244 2448
rect 8278 2414 8288 2448
rect 8236 2366 8288 2414
rect 8318 2450 8368 2496
rect 8318 2412 8383 2450
rect 8318 2378 8328 2412
rect 8362 2378 8383 2412
rect 8318 2366 8383 2378
rect 8413 2438 8465 2450
rect 8413 2404 8423 2438
rect 8457 2404 8465 2438
rect 8413 2366 8465 2404
rect 8519 2446 8571 2496
rect 8519 2412 8527 2446
rect 8561 2412 8571 2446
rect 8519 2366 8571 2412
rect 8601 2450 8651 2496
rect 8601 2412 8666 2450
rect 8601 2378 8611 2412
rect 8645 2378 8666 2412
rect 8601 2366 8666 2378
rect 8696 2422 8748 2450
rect 8696 2388 8706 2422
rect 8740 2388 8748 2422
rect 8696 2366 8748 2388
rect 8802 2420 8854 2494
rect 8802 2386 8810 2420
rect 8844 2386 8854 2420
rect 8802 2366 8854 2386
rect 8884 2472 8938 2494
rect 8884 2438 8894 2472
rect 8928 2438 8938 2472
rect 8884 2366 8938 2438
rect 8968 2450 9018 2494
rect 8968 2428 9056 2450
rect 8968 2394 8994 2428
rect 9028 2394 9056 2428
rect 8968 2366 9056 2394
rect 9086 2408 9142 2450
rect 9086 2374 9096 2408
rect 9130 2374 9142 2408
rect 9086 2366 9142 2374
rect 9172 2438 9222 2450
rect 9391 2438 9441 2494
rect 9172 2366 9237 2438
rect 9267 2412 9346 2438
rect 9267 2378 9287 2412
rect 9321 2378 9346 2412
rect 9267 2366 9346 2378
rect 9376 2366 9441 2438
rect 9471 2412 9523 2494
rect 9471 2378 9481 2412
rect 9515 2378 9523 2412
rect 9471 2366 9523 2378
rect 9577 2446 9629 2494
rect 9577 2412 9585 2446
rect 9619 2412 9629 2446
rect 9577 2366 9629 2412
rect 9659 2472 9713 2494
rect 9659 2438 9669 2472
rect 9703 2438 9713 2472
rect 9659 2366 9713 2438
rect 9743 2450 9793 2494
rect 9743 2428 9813 2450
rect 9743 2394 9769 2428
rect 9803 2394 9813 2428
rect 9743 2366 9813 2394
rect 9843 2408 9923 2450
rect 9843 2374 9853 2408
rect 9887 2374 9923 2408
rect 9843 2366 9923 2374
rect 9953 2438 10004 2450
rect 10170 2438 10220 2450
rect 9953 2366 10019 2438
rect 10049 2412 10125 2438
rect 10049 2378 10070 2412
rect 10104 2378 10125 2412
rect 10049 2366 10125 2378
rect 10155 2430 10220 2438
rect 10155 2396 10176 2430
rect 10210 2396 10220 2430
rect 10155 2366 10220 2396
rect 10250 2412 10302 2450
rect 10250 2378 10260 2412
rect 10294 2378 10302 2412
rect 10250 2366 10302 2378
rect 10356 2438 10408 2450
rect 10356 2404 10364 2438
rect 10398 2404 10408 2438
rect 10356 2366 10408 2404
rect 10438 2412 10492 2450
rect 10438 2378 10448 2412
rect 10482 2378 10492 2412
rect 10438 2366 10492 2378
rect 10522 2438 10574 2450
rect 10522 2404 10532 2438
rect 10566 2404 10574 2438
rect 10522 2366 10574 2404
rect 10628 2448 10680 2496
rect 10628 2414 10636 2448
rect 10670 2414 10680 2448
rect 10628 2366 10680 2414
rect 10710 2450 10760 2496
rect 10710 2412 10775 2450
rect 10710 2378 10720 2412
rect 10754 2378 10775 2412
rect 10710 2366 10775 2378
rect 10805 2438 10857 2450
rect 10805 2404 10815 2438
rect 10849 2404 10857 2438
rect 10805 2366 10857 2404
rect 10911 2446 10963 2496
rect 10911 2412 10919 2446
rect 10953 2412 10963 2446
rect 10911 2366 10963 2412
rect 10993 2450 11043 2496
rect 10993 2412 11058 2450
rect 10993 2378 11003 2412
rect 11037 2378 11058 2412
rect 10993 2366 11058 2378
rect 11088 2422 11140 2450
rect 11088 2388 11098 2422
rect 11132 2388 11140 2422
rect 11088 2366 11140 2388
rect 11194 2420 11246 2494
rect 11194 2386 11202 2420
rect 11236 2386 11246 2420
rect 11194 2366 11246 2386
rect 11276 2472 11330 2494
rect 11276 2438 11286 2472
rect 11320 2438 11330 2472
rect 11276 2366 11330 2438
rect 11360 2450 11410 2494
rect 11360 2428 11448 2450
rect 11360 2394 11386 2428
rect 11420 2394 11448 2428
rect 11360 2366 11448 2394
rect 11478 2408 11534 2450
rect 11478 2374 11488 2408
rect 11522 2374 11534 2408
rect 11478 2366 11534 2374
rect 11564 2438 11614 2450
rect 11783 2438 11833 2494
rect 11564 2366 11629 2438
rect 11659 2412 11738 2438
rect 11659 2378 11679 2412
rect 11713 2378 11738 2412
rect 11659 2366 11738 2378
rect 11768 2366 11833 2438
rect 11863 2412 11915 2494
rect 11863 2378 11873 2412
rect 11907 2378 11915 2412
rect 11863 2366 11915 2378
rect 11969 2446 12021 2494
rect 11969 2412 11977 2446
rect 12011 2412 12021 2446
rect 11969 2366 12021 2412
rect 12051 2472 12105 2494
rect 12051 2438 12061 2472
rect 12095 2438 12105 2472
rect 12051 2366 12105 2438
rect 12135 2450 12185 2494
rect 12135 2428 12205 2450
rect 12135 2394 12161 2428
rect 12195 2394 12205 2428
rect 12135 2366 12205 2394
rect 12235 2408 12315 2450
rect 12235 2374 12245 2408
rect 12279 2374 12315 2408
rect 12235 2366 12315 2374
rect 12345 2438 12396 2450
rect 12562 2438 12612 2450
rect 12345 2366 12411 2438
rect 12441 2412 12517 2438
rect 12441 2378 12462 2412
rect 12496 2378 12517 2412
rect 12441 2366 12517 2378
rect 12547 2430 12612 2438
rect 12547 2396 12568 2430
rect 12602 2396 12612 2430
rect 12547 2366 12612 2396
rect 12642 2412 12694 2450
rect 12642 2378 12652 2412
rect 12686 2378 12694 2412
rect 12642 2366 12694 2378
rect 12748 2438 12800 2450
rect 12748 2404 12756 2438
rect 12790 2404 12800 2438
rect 12748 2366 12800 2404
rect 12830 2412 12884 2450
rect 12830 2378 12840 2412
rect 12874 2378 12884 2412
rect 12830 2366 12884 2378
rect 12914 2438 12966 2450
rect 12914 2404 12924 2438
rect 12958 2404 12966 2438
rect 12914 2366 12966 2404
<< pdiff >>
rect 1062 6104 1114 6124
rect 1062 6070 1070 6104
rect 1104 6070 1114 6104
rect 1062 6036 1114 6070
rect 1062 6002 1070 6036
rect 1104 6002 1114 6036
rect 1062 5966 1114 6002
rect 1144 6104 1202 6124
rect 1144 6070 1156 6104
rect 1190 6070 1202 6104
rect 1144 6036 1202 6070
rect 1144 6002 1156 6036
rect 1190 6002 1202 6036
rect 1144 5966 1202 6002
rect 1232 6104 1284 6124
rect 1232 6070 1242 6104
rect 1276 6070 1284 6104
rect 1232 6023 1284 6070
rect 1232 5989 1242 6023
rect 1276 5989 1284 6023
rect 1232 5966 1284 5989
rect 1338 6106 1390 6124
rect 1338 6072 1346 6106
rect 1380 6072 1390 6106
rect 1338 6038 1390 6072
rect 1338 6004 1346 6038
rect 1380 6004 1390 6038
rect 1338 5970 1390 6004
rect 1338 5936 1346 5970
rect 1380 5936 1390 5970
rect 1338 5924 1390 5936
rect 1420 6112 1474 6124
rect 1420 6078 1430 6112
rect 1464 6078 1474 6112
rect 1420 6044 1474 6078
rect 1420 6010 1430 6044
rect 1464 6010 1474 6044
rect 1420 5924 1474 6010
rect 1504 6090 1558 6124
rect 1504 6056 1514 6090
rect 1548 6056 1558 6090
rect 1504 5995 1558 6056
rect 1504 5961 1514 5995
rect 1548 5961 1558 5995
rect 1504 5924 1558 5961
rect 1588 6112 1642 6124
rect 1588 6078 1598 6112
rect 1632 6078 1642 6112
rect 1588 6044 1642 6078
rect 1588 6010 1598 6044
rect 1632 6010 1642 6044
rect 1588 5924 1642 6010
rect 1672 6090 1726 6124
rect 1672 6056 1682 6090
rect 1716 6056 1726 6090
rect 1672 5995 1726 6056
rect 1672 5961 1682 5995
rect 1716 5961 1726 5995
rect 1672 5924 1726 5961
rect 1756 6112 1808 6124
rect 1756 6078 1766 6112
rect 1800 6078 1808 6112
rect 1756 6044 1808 6078
rect 1756 6010 1766 6044
rect 1800 6010 1808 6044
rect 1756 5976 1808 6010
rect 1756 5942 1766 5976
rect 1800 5942 1808 5976
rect 1756 5924 1808 5942
rect 2322 6112 2389 6124
rect 2322 6078 2330 6112
rect 2364 6078 2389 6112
rect 2322 6044 2389 6078
rect 2322 6010 2330 6044
rect 2364 6010 2389 6044
rect 2322 5976 2389 6010
rect 2322 5942 2330 5976
rect 2364 5942 2389 5976
rect 2322 5924 2389 5942
rect 2419 6102 2473 6124
rect 2419 6068 2429 6102
rect 2463 6068 2473 6102
rect 2419 5976 2473 6068
rect 2419 5942 2429 5976
rect 2463 5942 2473 5976
rect 2419 5924 2473 5942
rect 2503 6112 2573 6124
rect 2503 6078 2513 6112
rect 2547 6078 2573 6112
rect 2503 6044 2573 6078
rect 2503 6010 2513 6044
rect 2547 6010 2573 6044
rect 2503 5976 2573 6010
rect 2503 5942 2513 5976
rect 2547 5942 2573 5976
rect 2503 5924 2573 5942
rect 2603 6102 2657 6124
rect 2603 6068 2613 6102
rect 2647 6068 2657 6102
rect 2603 6028 2657 6068
rect 2603 5994 2613 6028
rect 2647 5994 2657 6028
rect 2603 5924 2657 5994
rect 2687 6112 2754 6124
rect 2687 6078 2697 6112
rect 2731 6078 2754 6112
rect 2687 6044 2754 6078
rect 2687 6010 2697 6044
rect 2731 6010 2754 6044
rect 2687 5996 2754 6010
rect 2784 6040 2855 6124
rect 2885 6092 2939 6124
rect 2885 6058 2895 6092
rect 2929 6058 2939 6092
rect 2885 6040 2939 6058
rect 2969 6040 3074 6124
rect 2784 5996 2840 6040
rect 2687 5924 2739 5996
rect 3024 5996 3074 6040
rect 3104 6078 3156 6124
rect 3104 6044 3114 6078
rect 3148 6044 3156 6078
rect 3663 6100 3762 6124
rect 3104 5996 3156 6044
rect 3210 5990 3262 6051
rect 3210 5956 3218 5990
rect 3252 5956 3262 5990
rect 3210 5943 3262 5956
rect 3292 5989 3346 6051
rect 3292 5955 3302 5989
rect 3336 5955 3346 5989
rect 3292 5943 3346 5955
rect 3376 6039 3428 6051
rect 3376 6005 3386 6039
rect 3420 6005 3428 6039
rect 3376 5943 3428 6005
rect 3482 6018 3534 6100
rect 3482 5984 3490 6018
rect 3524 5984 3534 6018
rect 3482 5972 3534 5984
rect 3564 6088 3618 6100
rect 3564 6054 3574 6088
rect 3608 6054 3618 6088
rect 3564 5972 3618 6054
rect 3648 6040 3762 6100
rect 3792 6086 3846 6124
rect 3792 6052 3802 6086
rect 3836 6052 3846 6086
rect 3792 6040 3846 6052
rect 3876 6040 3942 6124
rect 3648 5972 3706 6040
rect 3891 5996 3942 6040
rect 3972 6112 4026 6124
rect 3972 6078 3982 6112
rect 4016 6078 4026 6112
rect 3972 5996 4026 6078
rect 4056 6086 4108 6124
rect 4056 6052 4066 6086
rect 4100 6052 4108 6086
rect 4056 5996 4108 6052
rect 1061 5231 1113 5245
rect 1061 5197 1069 5231
rect 1103 5197 1113 5231
rect 1061 5163 1113 5197
rect 1061 5129 1069 5163
rect 1103 5129 1113 5163
rect 1061 5117 1113 5129
rect 1143 5215 1197 5245
rect 1143 5181 1153 5215
rect 1187 5181 1197 5215
rect 1143 5117 1197 5181
rect 1227 5231 1279 5245
rect 1227 5197 1237 5231
rect 1271 5197 1279 5231
rect 1227 5163 1279 5197
rect 1333 5215 1385 5251
rect 1333 5181 1341 5215
rect 1375 5181 1385 5215
rect 1333 5167 1385 5181
rect 1415 5231 1478 5251
rect 1415 5197 1425 5231
rect 1459 5197 1478 5231
rect 1415 5167 1478 5197
rect 1508 5238 1562 5251
rect 1508 5204 1518 5238
rect 1552 5204 1562 5238
rect 1508 5167 1562 5204
rect 1592 5167 1682 5251
rect 1712 5229 1788 5251
rect 1712 5195 1732 5229
rect 1766 5195 1788 5229
rect 1712 5167 1788 5195
rect 1818 5213 1896 5251
rect 1818 5179 1852 5213
rect 1886 5179 1896 5213
rect 1818 5167 1896 5179
rect 1227 5129 1237 5163
rect 1271 5129 1279 5163
rect 1227 5117 1279 5129
rect 1834 5145 1896 5167
rect 1834 5111 1852 5145
rect 1886 5111 1896 5145
rect 1834 5083 1896 5111
rect 1926 5083 1980 5251
rect 2010 5239 2117 5251
rect 2010 5205 2026 5239
rect 2060 5205 2117 5239
rect 2010 5171 2117 5205
rect 2010 5137 2026 5171
rect 2060 5137 2117 5171
rect 2010 5083 2117 5137
rect 2147 5167 2261 5251
rect 2291 5238 2345 5251
rect 2291 5204 2301 5238
rect 2335 5204 2345 5238
rect 2291 5167 2345 5204
rect 2375 5167 2463 5251
rect 2493 5239 2571 5251
rect 2493 5205 2515 5239
rect 2549 5205 2571 5239
rect 2493 5167 2571 5205
rect 2601 5213 2667 5251
rect 2601 5179 2623 5213
rect 2657 5179 2667 5213
rect 2601 5167 2667 5179
rect 2147 5083 2199 5167
rect 2616 5083 2667 5167
rect 2697 5083 2739 5251
rect 2769 5239 2821 5251
rect 2769 5205 2779 5239
rect 2813 5205 2821 5239
rect 2769 5083 2821 5205
rect 2982 5239 3034 5251
rect 2982 5205 2990 5239
rect 3024 5205 3034 5239
rect 2982 5183 3034 5205
rect 2885 5103 2937 5183
rect 2885 5069 2893 5103
rect 2927 5069 2937 5103
rect 2885 5055 2937 5069
rect 2967 5055 3034 5183
rect 2984 5051 3034 5055
rect 3064 5202 3116 5251
rect 3267 5235 3317 5251
rect 3064 5168 3074 5202
rect 3108 5168 3116 5202
rect 3064 5134 3116 5168
rect 3064 5100 3074 5134
rect 3108 5100 3116 5134
rect 3170 5221 3222 5235
rect 3170 5187 3178 5221
rect 3212 5187 3222 5221
rect 3170 5153 3222 5187
rect 3170 5119 3178 5153
rect 3212 5119 3222 5153
rect 3170 5107 3222 5119
rect 3252 5227 3317 5235
rect 3252 5193 3273 5227
rect 3307 5193 3317 5227
rect 3252 5159 3317 5193
rect 3252 5125 3273 5159
rect 3307 5125 3317 5159
rect 3252 5107 3317 5125
rect 3064 5051 3116 5100
rect 3267 5051 3317 5107
rect 3347 5203 3399 5251
rect 3347 5169 3357 5203
rect 3391 5169 3399 5203
rect 3347 5135 3399 5169
rect 3347 5101 3357 5135
rect 3391 5101 3399 5135
rect 3453 5231 3505 5245
rect 3453 5197 3461 5231
rect 3495 5197 3505 5231
rect 3453 5163 3505 5197
rect 3453 5129 3461 5163
rect 3495 5129 3505 5163
rect 3453 5117 3505 5129
rect 3535 5215 3589 5245
rect 3535 5181 3545 5215
rect 3579 5181 3589 5215
rect 3535 5117 3589 5181
rect 3619 5231 3671 5245
rect 3619 5197 3629 5231
rect 3663 5197 3671 5231
rect 3619 5163 3671 5197
rect 3725 5215 3777 5251
rect 3725 5181 3733 5215
rect 3767 5181 3777 5215
rect 3725 5167 3777 5181
rect 3807 5231 3870 5251
rect 3807 5197 3817 5231
rect 3851 5197 3870 5231
rect 3807 5167 3870 5197
rect 3900 5238 3954 5251
rect 3900 5204 3910 5238
rect 3944 5204 3954 5238
rect 3900 5167 3954 5204
rect 3984 5167 4074 5251
rect 4104 5229 4180 5251
rect 4104 5195 4124 5229
rect 4158 5195 4180 5229
rect 4104 5167 4180 5195
rect 4210 5213 4288 5251
rect 4210 5179 4244 5213
rect 4278 5179 4288 5213
rect 4210 5167 4288 5179
rect 3619 5129 3629 5163
rect 3663 5129 3671 5163
rect 3619 5117 3671 5129
rect 3347 5051 3399 5101
rect 4226 5145 4288 5167
rect 4226 5111 4244 5145
rect 4278 5111 4288 5145
rect 4226 5083 4288 5111
rect 4318 5083 4372 5251
rect 4402 5239 4509 5251
rect 4402 5205 4418 5239
rect 4452 5205 4509 5239
rect 4402 5171 4509 5205
rect 4402 5137 4418 5171
rect 4452 5137 4509 5171
rect 4402 5083 4509 5137
rect 4539 5167 4653 5251
rect 4683 5238 4737 5251
rect 4683 5204 4693 5238
rect 4727 5204 4737 5238
rect 4683 5167 4737 5204
rect 4767 5167 4855 5251
rect 4885 5239 4963 5251
rect 4885 5205 4907 5239
rect 4941 5205 4963 5239
rect 4885 5167 4963 5205
rect 4993 5213 5059 5251
rect 4993 5179 5015 5213
rect 5049 5179 5059 5213
rect 4993 5167 5059 5179
rect 4539 5083 4591 5167
rect 5008 5083 5059 5167
rect 5089 5083 5131 5251
rect 5161 5239 5213 5251
rect 5161 5205 5171 5239
rect 5205 5205 5213 5239
rect 5374 5239 5426 5251
rect 5161 5083 5213 5205
rect 5374 5205 5382 5239
rect 5416 5205 5426 5239
rect 5374 5183 5426 5205
rect 5277 5103 5329 5183
rect 5277 5069 5285 5103
rect 5319 5069 5329 5103
rect 5277 5055 5329 5069
rect 5359 5055 5426 5183
rect 5376 5051 5426 5055
rect 5456 5202 5508 5251
rect 5659 5235 5709 5251
rect 5456 5168 5466 5202
rect 5500 5168 5508 5202
rect 5456 5134 5508 5168
rect 5456 5100 5466 5134
rect 5500 5100 5508 5134
rect 5562 5221 5614 5235
rect 5562 5187 5570 5221
rect 5604 5187 5614 5221
rect 5562 5153 5614 5187
rect 5562 5119 5570 5153
rect 5604 5119 5614 5153
rect 5562 5107 5614 5119
rect 5644 5227 5709 5235
rect 5644 5193 5665 5227
rect 5699 5193 5709 5227
rect 5644 5159 5709 5193
rect 5644 5125 5665 5159
rect 5699 5125 5709 5159
rect 5644 5107 5709 5125
rect 5456 5051 5508 5100
rect 5659 5051 5709 5107
rect 5739 5203 5791 5251
rect 5739 5169 5749 5203
rect 5783 5169 5791 5203
rect 5739 5135 5791 5169
rect 5739 5101 5749 5135
rect 5783 5101 5791 5135
rect 5845 5231 5897 5245
rect 5845 5197 5853 5231
rect 5887 5197 5897 5231
rect 5845 5163 5897 5197
rect 5845 5129 5853 5163
rect 5887 5129 5897 5163
rect 5845 5117 5897 5129
rect 5927 5215 5981 5245
rect 5927 5181 5937 5215
rect 5971 5181 5981 5215
rect 5927 5117 5981 5181
rect 6011 5231 6063 5245
rect 6011 5197 6021 5231
rect 6055 5197 6063 5231
rect 6011 5163 6063 5197
rect 6117 5215 6169 5251
rect 6117 5181 6125 5215
rect 6159 5181 6169 5215
rect 6117 5167 6169 5181
rect 6199 5231 6262 5251
rect 6199 5197 6209 5231
rect 6243 5197 6262 5231
rect 6199 5167 6262 5197
rect 6292 5238 6346 5251
rect 6292 5204 6302 5238
rect 6336 5204 6346 5238
rect 6292 5167 6346 5204
rect 6376 5167 6466 5251
rect 6496 5229 6572 5251
rect 6496 5195 6516 5229
rect 6550 5195 6572 5229
rect 6496 5167 6572 5195
rect 6602 5213 6680 5251
rect 6602 5179 6636 5213
rect 6670 5179 6680 5213
rect 6602 5167 6680 5179
rect 6011 5129 6021 5163
rect 6055 5129 6063 5163
rect 6011 5117 6063 5129
rect 5739 5051 5791 5101
rect 6618 5145 6680 5167
rect 6618 5111 6636 5145
rect 6670 5111 6680 5145
rect 6618 5083 6680 5111
rect 6710 5083 6764 5251
rect 6794 5239 6901 5251
rect 6794 5205 6810 5239
rect 6844 5205 6901 5239
rect 6794 5171 6901 5205
rect 6794 5137 6810 5171
rect 6844 5137 6901 5171
rect 6794 5083 6901 5137
rect 6931 5167 7045 5251
rect 7075 5238 7129 5251
rect 7075 5204 7085 5238
rect 7119 5204 7129 5238
rect 7075 5167 7129 5204
rect 7159 5167 7247 5251
rect 7277 5239 7355 5251
rect 7277 5205 7299 5239
rect 7333 5205 7355 5239
rect 7277 5167 7355 5205
rect 7385 5213 7451 5251
rect 7385 5179 7407 5213
rect 7441 5179 7451 5213
rect 7385 5167 7451 5179
rect 6931 5083 6983 5167
rect 7400 5083 7451 5167
rect 7481 5083 7523 5251
rect 7553 5239 7605 5251
rect 7553 5205 7563 5239
rect 7597 5205 7605 5239
rect 7766 5239 7818 5251
rect 7553 5083 7605 5205
rect 7766 5205 7774 5239
rect 7808 5205 7818 5239
rect 7766 5183 7818 5205
rect 7669 5103 7721 5183
rect 7669 5069 7677 5103
rect 7711 5069 7721 5103
rect 7669 5055 7721 5069
rect 7751 5055 7818 5183
rect 7768 5051 7818 5055
rect 7848 5202 7900 5251
rect 8051 5235 8101 5251
rect 7848 5168 7858 5202
rect 7892 5168 7900 5202
rect 7848 5134 7900 5168
rect 7848 5100 7858 5134
rect 7892 5100 7900 5134
rect 7954 5221 8006 5235
rect 7954 5187 7962 5221
rect 7996 5187 8006 5221
rect 7954 5153 8006 5187
rect 7954 5119 7962 5153
rect 7996 5119 8006 5153
rect 7954 5107 8006 5119
rect 8036 5227 8101 5235
rect 8036 5193 8057 5227
rect 8091 5193 8101 5227
rect 8036 5159 8101 5193
rect 8036 5125 8057 5159
rect 8091 5125 8101 5159
rect 8036 5107 8101 5125
rect 7848 5051 7900 5100
rect 8051 5051 8101 5107
rect 8131 5203 8183 5251
rect 8131 5169 8141 5203
rect 8175 5169 8183 5203
rect 8131 5135 8183 5169
rect 8131 5101 8141 5135
rect 8175 5101 8183 5135
rect 8237 5231 8289 5245
rect 8237 5197 8245 5231
rect 8279 5197 8289 5231
rect 8237 5163 8289 5197
rect 8237 5129 8245 5163
rect 8279 5129 8289 5163
rect 8237 5117 8289 5129
rect 8319 5215 8373 5245
rect 8319 5181 8329 5215
rect 8363 5181 8373 5215
rect 8319 5117 8373 5181
rect 8403 5231 8455 5245
rect 8403 5197 8413 5231
rect 8447 5197 8455 5231
rect 8403 5163 8455 5197
rect 8509 5215 8561 5251
rect 8509 5181 8517 5215
rect 8551 5181 8561 5215
rect 8509 5167 8561 5181
rect 8591 5231 8654 5251
rect 8591 5197 8601 5231
rect 8635 5197 8654 5231
rect 8591 5167 8654 5197
rect 8684 5238 8738 5251
rect 8684 5204 8694 5238
rect 8728 5204 8738 5238
rect 8684 5167 8738 5204
rect 8768 5167 8858 5251
rect 8888 5229 8964 5251
rect 8888 5195 8908 5229
rect 8942 5195 8964 5229
rect 8888 5167 8964 5195
rect 8994 5213 9072 5251
rect 8994 5179 9028 5213
rect 9062 5179 9072 5213
rect 8994 5167 9072 5179
rect 8403 5129 8413 5163
rect 8447 5129 8455 5163
rect 8403 5117 8455 5129
rect 8131 5051 8183 5101
rect 9010 5145 9072 5167
rect 9010 5111 9028 5145
rect 9062 5111 9072 5145
rect 9010 5083 9072 5111
rect 9102 5083 9156 5251
rect 9186 5239 9293 5251
rect 9186 5205 9202 5239
rect 9236 5205 9293 5239
rect 9186 5171 9293 5205
rect 9186 5137 9202 5171
rect 9236 5137 9293 5171
rect 9186 5083 9293 5137
rect 9323 5167 9437 5251
rect 9467 5238 9521 5251
rect 9467 5204 9477 5238
rect 9511 5204 9521 5238
rect 9467 5167 9521 5204
rect 9551 5167 9639 5251
rect 9669 5239 9747 5251
rect 9669 5205 9691 5239
rect 9725 5205 9747 5239
rect 9669 5167 9747 5205
rect 9777 5213 9843 5251
rect 9777 5179 9799 5213
rect 9833 5179 9843 5213
rect 9777 5167 9843 5179
rect 9323 5083 9375 5167
rect 9792 5083 9843 5167
rect 9873 5083 9915 5251
rect 9945 5239 9997 5251
rect 9945 5205 9955 5239
rect 9989 5205 9997 5239
rect 10158 5239 10210 5251
rect 9945 5083 9997 5205
rect 10158 5205 10166 5239
rect 10200 5205 10210 5239
rect 10158 5183 10210 5205
rect 10061 5103 10113 5183
rect 10061 5069 10069 5103
rect 10103 5069 10113 5103
rect 10061 5055 10113 5069
rect 10143 5055 10210 5183
rect 10160 5051 10210 5055
rect 10240 5202 10292 5251
rect 10443 5235 10493 5251
rect 10240 5168 10250 5202
rect 10284 5168 10292 5202
rect 10240 5134 10292 5168
rect 10240 5100 10250 5134
rect 10284 5100 10292 5134
rect 10346 5221 10398 5235
rect 10346 5187 10354 5221
rect 10388 5187 10398 5221
rect 10346 5153 10398 5187
rect 10346 5119 10354 5153
rect 10388 5119 10398 5153
rect 10346 5107 10398 5119
rect 10428 5227 10493 5235
rect 10428 5193 10449 5227
rect 10483 5193 10493 5227
rect 10428 5159 10493 5193
rect 10428 5125 10449 5159
rect 10483 5125 10493 5159
rect 10428 5107 10493 5125
rect 10240 5051 10292 5100
rect 10443 5051 10493 5107
rect 10523 5203 10575 5251
rect 10523 5169 10533 5203
rect 10567 5169 10575 5203
rect 10523 5135 10575 5169
rect 10523 5101 10533 5135
rect 10567 5101 10575 5135
rect 10629 5231 10681 5245
rect 10629 5197 10637 5231
rect 10671 5197 10681 5231
rect 10629 5163 10681 5197
rect 10629 5129 10637 5163
rect 10671 5129 10681 5163
rect 10629 5117 10681 5129
rect 10711 5215 10765 5245
rect 10711 5181 10721 5215
rect 10755 5181 10765 5215
rect 10711 5117 10765 5181
rect 10795 5231 10847 5245
rect 10795 5197 10805 5231
rect 10839 5197 10847 5231
rect 10795 5163 10847 5197
rect 10901 5215 10953 5251
rect 10901 5181 10909 5215
rect 10943 5181 10953 5215
rect 10901 5167 10953 5181
rect 10983 5231 11046 5251
rect 10983 5197 10993 5231
rect 11027 5197 11046 5231
rect 10983 5167 11046 5197
rect 11076 5238 11130 5251
rect 11076 5204 11086 5238
rect 11120 5204 11130 5238
rect 11076 5167 11130 5204
rect 11160 5167 11250 5251
rect 11280 5229 11356 5251
rect 11280 5195 11300 5229
rect 11334 5195 11356 5229
rect 11280 5167 11356 5195
rect 11386 5213 11464 5251
rect 11386 5179 11420 5213
rect 11454 5179 11464 5213
rect 11386 5167 11464 5179
rect 10795 5129 10805 5163
rect 10839 5129 10847 5163
rect 10795 5117 10847 5129
rect 10523 5051 10575 5101
rect 11402 5145 11464 5167
rect 11402 5111 11420 5145
rect 11454 5111 11464 5145
rect 11402 5083 11464 5111
rect 11494 5083 11548 5251
rect 11578 5239 11685 5251
rect 11578 5205 11594 5239
rect 11628 5205 11685 5239
rect 11578 5171 11685 5205
rect 11578 5137 11594 5171
rect 11628 5137 11685 5171
rect 11578 5083 11685 5137
rect 11715 5167 11829 5251
rect 11859 5238 11913 5251
rect 11859 5204 11869 5238
rect 11903 5204 11913 5238
rect 11859 5167 11913 5204
rect 11943 5167 12031 5251
rect 12061 5239 12139 5251
rect 12061 5205 12083 5239
rect 12117 5205 12139 5239
rect 12061 5167 12139 5205
rect 12169 5213 12235 5251
rect 12169 5179 12191 5213
rect 12225 5179 12235 5213
rect 12169 5167 12235 5179
rect 11715 5083 11767 5167
rect 12184 5083 12235 5167
rect 12265 5083 12307 5251
rect 12337 5239 12389 5251
rect 12337 5205 12347 5239
rect 12381 5205 12389 5239
rect 12550 5239 12602 5251
rect 12337 5083 12389 5205
rect 12550 5205 12558 5239
rect 12592 5205 12602 5239
rect 12550 5183 12602 5205
rect 12453 5103 12505 5183
rect 12453 5069 12461 5103
rect 12495 5069 12505 5103
rect 12453 5055 12505 5069
rect 12535 5055 12602 5183
rect 12552 5051 12602 5055
rect 12632 5202 12684 5251
rect 12835 5235 12885 5251
rect 12632 5168 12642 5202
rect 12676 5168 12684 5202
rect 12632 5134 12684 5168
rect 12632 5100 12642 5134
rect 12676 5100 12684 5134
rect 12738 5221 12790 5235
rect 12738 5187 12746 5221
rect 12780 5187 12790 5221
rect 12738 5153 12790 5187
rect 12738 5119 12746 5153
rect 12780 5119 12790 5153
rect 12738 5107 12790 5119
rect 12820 5227 12885 5235
rect 12820 5193 12841 5227
rect 12875 5193 12885 5227
rect 12820 5159 12885 5193
rect 12820 5125 12841 5159
rect 12875 5125 12885 5159
rect 12820 5107 12885 5125
rect 12632 5051 12684 5100
rect 12835 5051 12885 5107
rect 12915 5203 12967 5251
rect 12915 5169 12925 5203
rect 12959 5169 12967 5203
rect 12915 5135 12967 5169
rect 12915 5101 12925 5135
rect 12959 5101 12967 5135
rect 12915 5051 12967 5101
rect 621 4542 673 4562
rect 621 4508 629 4542
rect 663 4508 673 4542
rect 621 4474 673 4508
rect 621 4440 629 4474
rect 663 4440 673 4474
rect 621 4404 673 4440
rect 703 4542 761 4562
rect 703 4508 715 4542
rect 749 4508 761 4542
rect 703 4474 761 4508
rect 703 4440 715 4474
rect 749 4440 761 4474
rect 703 4404 761 4440
rect 791 4542 843 4562
rect 791 4508 801 4542
rect 835 4508 843 4542
rect 791 4461 843 4508
rect 791 4427 801 4461
rect 835 4427 843 4461
rect 791 4404 843 4427
rect 897 4544 949 4562
rect 897 4510 905 4544
rect 939 4510 949 4544
rect 897 4476 949 4510
rect 897 4442 905 4476
rect 939 4442 949 4476
rect 897 4408 949 4442
rect 897 4374 905 4408
rect 939 4374 949 4408
rect 897 4362 949 4374
rect 979 4550 1033 4562
rect 979 4516 989 4550
rect 1023 4516 1033 4550
rect 979 4482 1033 4516
rect 979 4448 989 4482
rect 1023 4448 1033 4482
rect 979 4362 1033 4448
rect 1063 4528 1117 4562
rect 1063 4494 1073 4528
rect 1107 4494 1117 4528
rect 1063 4433 1117 4494
rect 1063 4399 1073 4433
rect 1107 4399 1117 4433
rect 1063 4362 1117 4399
rect 1147 4550 1201 4562
rect 1147 4516 1157 4550
rect 1191 4516 1201 4550
rect 1147 4482 1201 4516
rect 1147 4448 1157 4482
rect 1191 4448 1201 4482
rect 1147 4362 1201 4448
rect 1231 4528 1285 4562
rect 1231 4494 1241 4528
rect 1275 4494 1285 4528
rect 1231 4433 1285 4494
rect 1231 4399 1241 4433
rect 1275 4399 1285 4433
rect 1231 4362 1285 4399
rect 1315 4550 1367 4562
rect 1315 4516 1325 4550
rect 1359 4516 1367 4550
rect 1315 4482 1367 4516
rect 1315 4448 1325 4482
rect 1359 4448 1367 4482
rect 1315 4414 1367 4448
rect 1315 4380 1325 4414
rect 1359 4380 1367 4414
rect 1315 4362 1367 4380
rect 1429 4550 1481 4562
rect 1429 4516 1437 4550
rect 1471 4516 1481 4550
rect 1429 4482 1481 4516
rect 1429 4448 1437 4482
rect 1471 4448 1481 4482
rect 1429 4414 1481 4448
rect 1429 4380 1437 4414
rect 1471 4380 1481 4414
rect 1429 4362 1481 4380
rect 1511 4544 1565 4562
rect 1511 4510 1521 4544
rect 1555 4510 1565 4544
rect 1511 4476 1565 4510
rect 1511 4442 1521 4476
rect 1555 4442 1565 4476
rect 1511 4408 1565 4442
rect 1511 4374 1521 4408
rect 1555 4374 1565 4408
rect 1511 4362 1565 4374
rect 1595 4550 1649 4562
rect 1595 4516 1605 4550
rect 1639 4516 1649 4550
rect 1595 4482 1649 4516
rect 1595 4448 1605 4482
rect 1639 4448 1649 4482
rect 1595 4362 1649 4448
rect 1679 4544 1733 4562
rect 1679 4510 1689 4544
rect 1723 4510 1733 4544
rect 1679 4476 1733 4510
rect 1679 4442 1689 4476
rect 1723 4442 1733 4476
rect 1679 4408 1733 4442
rect 1679 4374 1689 4408
rect 1723 4374 1733 4408
rect 1679 4362 1733 4374
rect 1763 4550 1817 4562
rect 1763 4516 1773 4550
rect 1807 4516 1817 4550
rect 1763 4482 1817 4516
rect 1763 4448 1773 4482
rect 1807 4448 1817 4482
rect 1763 4362 1817 4448
rect 1847 4544 1901 4562
rect 1847 4510 1857 4544
rect 1891 4510 1901 4544
rect 1847 4476 1901 4510
rect 1847 4442 1857 4476
rect 1891 4442 1901 4476
rect 1847 4408 1901 4442
rect 1847 4374 1857 4408
rect 1891 4374 1901 4408
rect 1847 4362 1901 4374
rect 1931 4550 1985 4562
rect 1931 4516 1941 4550
rect 1975 4516 1985 4550
rect 1931 4482 1985 4516
rect 1931 4448 1941 4482
rect 1975 4448 1985 4482
rect 1931 4362 1985 4448
rect 2015 4544 2069 4562
rect 2015 4510 2025 4544
rect 2059 4510 2069 4544
rect 2015 4476 2069 4510
rect 2015 4442 2025 4476
rect 2059 4442 2069 4476
rect 2015 4408 2069 4442
rect 2015 4374 2025 4408
rect 2059 4374 2069 4408
rect 2015 4362 2069 4374
rect 2099 4550 2153 4562
rect 2099 4516 2109 4550
rect 2143 4516 2153 4550
rect 2099 4482 2153 4516
rect 2099 4448 2109 4482
rect 2143 4448 2153 4482
rect 2099 4362 2153 4448
rect 2183 4544 2237 4562
rect 2183 4510 2193 4544
rect 2227 4510 2237 4544
rect 2183 4476 2237 4510
rect 2183 4442 2193 4476
rect 2227 4442 2237 4476
rect 2183 4408 2237 4442
rect 2183 4374 2193 4408
rect 2227 4374 2237 4408
rect 2183 4362 2237 4374
rect 2267 4550 2321 4562
rect 2267 4516 2277 4550
rect 2311 4516 2321 4550
rect 2267 4482 2321 4516
rect 2267 4448 2277 4482
rect 2311 4448 2321 4482
rect 2267 4362 2321 4448
rect 2351 4544 2405 4562
rect 2351 4510 2361 4544
rect 2395 4510 2405 4544
rect 2351 4476 2405 4510
rect 2351 4442 2361 4476
rect 2395 4442 2405 4476
rect 2351 4408 2405 4442
rect 2351 4374 2361 4408
rect 2395 4374 2405 4408
rect 2351 4362 2405 4374
rect 2435 4550 2489 4562
rect 2435 4516 2445 4550
rect 2479 4516 2489 4550
rect 2435 4482 2489 4516
rect 2435 4448 2445 4482
rect 2479 4448 2489 4482
rect 2435 4362 2489 4448
rect 2519 4544 2573 4562
rect 2519 4510 2529 4544
rect 2563 4510 2573 4544
rect 2519 4476 2573 4510
rect 2519 4442 2529 4476
rect 2563 4442 2573 4476
rect 2519 4408 2573 4442
rect 2519 4374 2529 4408
rect 2563 4374 2573 4408
rect 2519 4362 2573 4374
rect 2603 4550 2657 4562
rect 2603 4516 2613 4550
rect 2647 4516 2657 4550
rect 2603 4482 2657 4516
rect 2603 4448 2613 4482
rect 2647 4448 2657 4482
rect 2603 4362 2657 4448
rect 2687 4544 2741 4562
rect 2687 4510 2697 4544
rect 2731 4510 2741 4544
rect 2687 4476 2741 4510
rect 2687 4442 2697 4476
rect 2731 4442 2741 4476
rect 2687 4408 2741 4442
rect 2687 4374 2697 4408
rect 2731 4374 2741 4408
rect 2687 4362 2741 4374
rect 2771 4550 2825 4562
rect 2771 4516 2781 4550
rect 2815 4516 2825 4550
rect 2771 4482 2825 4516
rect 2771 4448 2781 4482
rect 2815 4448 2825 4482
rect 2771 4362 2825 4448
rect 2855 4544 2909 4562
rect 2855 4510 2865 4544
rect 2899 4510 2909 4544
rect 2855 4476 2909 4510
rect 2855 4442 2865 4476
rect 2899 4442 2909 4476
rect 2855 4408 2909 4442
rect 2855 4374 2865 4408
rect 2899 4374 2909 4408
rect 2855 4362 2909 4374
rect 2939 4550 2993 4562
rect 2939 4516 2949 4550
rect 2983 4516 2993 4550
rect 2939 4482 2993 4516
rect 2939 4448 2949 4482
rect 2983 4448 2993 4482
rect 2939 4362 2993 4448
rect 3023 4544 3077 4562
rect 3023 4510 3033 4544
rect 3067 4510 3077 4544
rect 3023 4476 3077 4510
rect 3023 4442 3033 4476
rect 3067 4442 3077 4476
rect 3023 4408 3077 4442
rect 3023 4374 3033 4408
rect 3067 4374 3077 4408
rect 3023 4362 3077 4374
rect 3107 4550 3161 4562
rect 3107 4516 3117 4550
rect 3151 4516 3161 4550
rect 3107 4482 3161 4516
rect 3107 4448 3117 4482
rect 3151 4448 3161 4482
rect 3107 4362 3161 4448
rect 3191 4544 3245 4562
rect 3191 4510 3201 4544
rect 3235 4510 3245 4544
rect 3191 4476 3245 4510
rect 3191 4442 3201 4476
rect 3235 4442 3245 4476
rect 3191 4408 3245 4442
rect 3191 4374 3201 4408
rect 3235 4374 3245 4408
rect 3191 4362 3245 4374
rect 3275 4550 3327 4562
rect 3275 4516 3285 4550
rect 3319 4516 3327 4550
rect 3275 4482 3327 4516
rect 3275 4448 3285 4482
rect 3319 4448 3327 4482
rect 3275 4362 3327 4448
rect 3453 4514 3505 4562
rect 3453 4480 3461 4514
rect 3495 4480 3505 4514
rect 3453 4446 3505 4480
rect 3453 4412 3461 4446
rect 3495 4412 3505 4446
rect 3453 4362 3505 4412
rect 3535 4546 3585 4562
rect 3535 4538 3600 4546
rect 3535 4504 3545 4538
rect 3579 4504 3600 4538
rect 3535 4470 3600 4504
rect 3535 4436 3545 4470
rect 3579 4436 3600 4470
rect 3535 4418 3600 4436
rect 3630 4532 3682 4546
rect 3630 4498 3640 4532
rect 3674 4498 3682 4532
rect 3630 4464 3682 4498
rect 3630 4430 3640 4464
rect 3674 4430 3682 4464
rect 3630 4418 3682 4430
rect 3736 4513 3788 4562
rect 3736 4479 3744 4513
rect 3778 4479 3788 4513
rect 3736 4445 3788 4479
rect 3535 4362 3585 4418
rect 3736 4411 3744 4445
rect 3778 4411 3788 4445
rect 3736 4362 3788 4411
rect 3818 4550 3870 4562
rect 3818 4516 3828 4550
rect 3862 4516 3870 4550
rect 4031 4550 4083 4562
rect 3818 4494 3870 4516
rect 4031 4516 4039 4550
rect 4073 4516 4083 4550
rect 3818 4366 3885 4494
rect 3915 4414 3967 4494
rect 3915 4380 3925 4414
rect 3959 4380 3967 4414
rect 4031 4394 4083 4516
rect 4113 4394 4155 4562
rect 4185 4524 4251 4562
rect 4185 4490 4195 4524
rect 4229 4490 4251 4524
rect 4185 4478 4251 4490
rect 4281 4550 4359 4562
rect 4281 4516 4303 4550
rect 4337 4516 4359 4550
rect 4281 4478 4359 4516
rect 4389 4478 4477 4562
rect 4507 4549 4561 4562
rect 4507 4515 4517 4549
rect 4551 4515 4561 4549
rect 4507 4478 4561 4515
rect 4591 4478 4705 4562
rect 4185 4394 4236 4478
rect 3915 4366 3967 4380
rect 3818 4362 3868 4366
rect 4653 4394 4705 4478
rect 4735 4550 4842 4562
rect 4735 4516 4792 4550
rect 4826 4516 4842 4550
rect 4735 4482 4842 4516
rect 4735 4448 4792 4482
rect 4826 4448 4842 4482
rect 4735 4394 4842 4448
rect 4872 4394 4926 4562
rect 4956 4524 5034 4562
rect 4956 4490 4966 4524
rect 5000 4490 5034 4524
rect 4956 4478 5034 4490
rect 5064 4540 5140 4562
rect 5064 4506 5086 4540
rect 5120 4506 5140 4540
rect 5064 4478 5140 4506
rect 5170 4478 5260 4562
rect 5290 4549 5344 4562
rect 5290 4515 5300 4549
rect 5334 4515 5344 4549
rect 5290 4478 5344 4515
rect 5374 4542 5437 4562
rect 5374 4508 5393 4542
rect 5427 4508 5437 4542
rect 5374 4478 5437 4508
rect 5467 4526 5519 4562
rect 5467 4492 5477 4526
rect 5511 4492 5519 4526
rect 5467 4478 5519 4492
rect 5573 4542 5625 4556
rect 5573 4508 5581 4542
rect 5615 4508 5625 4542
rect 4956 4456 5018 4478
rect 4956 4422 4966 4456
rect 5000 4422 5018 4456
rect 4956 4394 5018 4422
rect 5573 4474 5625 4508
rect 5573 4440 5581 4474
rect 5615 4440 5625 4474
rect 5573 4428 5625 4440
rect 5655 4526 5709 4556
rect 5655 4492 5665 4526
rect 5699 4492 5709 4526
rect 5655 4428 5709 4492
rect 5739 4542 5791 4556
rect 5739 4508 5749 4542
rect 5783 4508 5791 4542
rect 5739 4474 5791 4508
rect 5739 4440 5749 4474
rect 5783 4440 5791 4474
rect 5739 4428 5791 4440
rect 5845 4514 5897 4562
rect 5845 4480 5853 4514
rect 5887 4480 5897 4514
rect 5845 4446 5897 4480
rect 5845 4412 5853 4446
rect 5887 4412 5897 4446
rect 5845 4362 5897 4412
rect 5927 4546 5977 4562
rect 5927 4538 5992 4546
rect 5927 4504 5937 4538
rect 5971 4504 5992 4538
rect 5927 4470 5992 4504
rect 5927 4436 5937 4470
rect 5971 4436 5992 4470
rect 5927 4418 5992 4436
rect 6022 4532 6074 4546
rect 6022 4498 6032 4532
rect 6066 4498 6074 4532
rect 6022 4464 6074 4498
rect 6022 4430 6032 4464
rect 6066 4430 6074 4464
rect 6022 4418 6074 4430
rect 6128 4513 6180 4562
rect 6128 4479 6136 4513
rect 6170 4479 6180 4513
rect 6128 4445 6180 4479
rect 5927 4362 5977 4418
rect 6128 4411 6136 4445
rect 6170 4411 6180 4445
rect 6128 4362 6180 4411
rect 6210 4550 6262 4562
rect 6210 4516 6220 4550
rect 6254 4516 6262 4550
rect 6423 4550 6475 4562
rect 6210 4494 6262 4516
rect 6423 4516 6431 4550
rect 6465 4516 6475 4550
rect 6210 4366 6277 4494
rect 6307 4414 6359 4494
rect 6307 4380 6317 4414
rect 6351 4380 6359 4414
rect 6423 4394 6475 4516
rect 6505 4394 6547 4562
rect 6577 4524 6643 4562
rect 6577 4490 6587 4524
rect 6621 4490 6643 4524
rect 6577 4478 6643 4490
rect 6673 4550 6751 4562
rect 6673 4516 6695 4550
rect 6729 4516 6751 4550
rect 6673 4478 6751 4516
rect 6781 4478 6869 4562
rect 6899 4549 6953 4562
rect 6899 4515 6909 4549
rect 6943 4515 6953 4549
rect 6899 4478 6953 4515
rect 6983 4478 7097 4562
rect 6577 4394 6628 4478
rect 6307 4366 6359 4380
rect 6210 4362 6260 4366
rect 7045 4394 7097 4478
rect 7127 4550 7234 4562
rect 7127 4516 7184 4550
rect 7218 4516 7234 4550
rect 7127 4482 7234 4516
rect 7127 4448 7184 4482
rect 7218 4448 7234 4482
rect 7127 4394 7234 4448
rect 7264 4394 7318 4562
rect 7348 4524 7426 4562
rect 7348 4490 7358 4524
rect 7392 4490 7426 4524
rect 7348 4478 7426 4490
rect 7456 4540 7532 4562
rect 7456 4506 7478 4540
rect 7512 4506 7532 4540
rect 7456 4478 7532 4506
rect 7562 4478 7652 4562
rect 7682 4549 7736 4562
rect 7682 4515 7692 4549
rect 7726 4515 7736 4549
rect 7682 4478 7736 4515
rect 7766 4542 7829 4562
rect 7766 4508 7785 4542
rect 7819 4508 7829 4542
rect 7766 4478 7829 4508
rect 7859 4526 7911 4562
rect 7859 4492 7869 4526
rect 7903 4492 7911 4526
rect 7859 4478 7911 4492
rect 7965 4542 8017 4556
rect 7965 4508 7973 4542
rect 8007 4508 8017 4542
rect 7348 4456 7410 4478
rect 7348 4422 7358 4456
rect 7392 4422 7410 4456
rect 7348 4394 7410 4422
rect 7965 4474 8017 4508
rect 7965 4440 7973 4474
rect 8007 4440 8017 4474
rect 7965 4428 8017 4440
rect 8047 4526 8101 4556
rect 8047 4492 8057 4526
rect 8091 4492 8101 4526
rect 8047 4428 8101 4492
rect 8131 4542 8183 4556
rect 8131 4508 8141 4542
rect 8175 4508 8183 4542
rect 8131 4474 8183 4508
rect 8131 4440 8141 4474
rect 8175 4440 8183 4474
rect 8131 4428 8183 4440
rect 8237 4514 8289 4562
rect 8237 4480 8245 4514
rect 8279 4480 8289 4514
rect 8237 4446 8289 4480
rect 8237 4412 8245 4446
rect 8279 4412 8289 4446
rect 8237 4362 8289 4412
rect 8319 4546 8369 4562
rect 8319 4538 8384 4546
rect 8319 4504 8329 4538
rect 8363 4504 8384 4538
rect 8319 4470 8384 4504
rect 8319 4436 8329 4470
rect 8363 4436 8384 4470
rect 8319 4418 8384 4436
rect 8414 4532 8466 4546
rect 8414 4498 8424 4532
rect 8458 4498 8466 4532
rect 8414 4464 8466 4498
rect 8414 4430 8424 4464
rect 8458 4430 8466 4464
rect 8414 4418 8466 4430
rect 8520 4513 8572 4562
rect 8520 4479 8528 4513
rect 8562 4479 8572 4513
rect 8520 4445 8572 4479
rect 8319 4362 8369 4418
rect 8520 4411 8528 4445
rect 8562 4411 8572 4445
rect 8520 4362 8572 4411
rect 8602 4550 8654 4562
rect 8602 4516 8612 4550
rect 8646 4516 8654 4550
rect 8815 4550 8867 4562
rect 8602 4494 8654 4516
rect 8815 4516 8823 4550
rect 8857 4516 8867 4550
rect 8602 4366 8669 4494
rect 8699 4414 8751 4494
rect 8699 4380 8709 4414
rect 8743 4380 8751 4414
rect 8815 4394 8867 4516
rect 8897 4394 8939 4562
rect 8969 4524 9035 4562
rect 8969 4490 8979 4524
rect 9013 4490 9035 4524
rect 8969 4478 9035 4490
rect 9065 4550 9143 4562
rect 9065 4516 9087 4550
rect 9121 4516 9143 4550
rect 9065 4478 9143 4516
rect 9173 4478 9261 4562
rect 9291 4549 9345 4562
rect 9291 4515 9301 4549
rect 9335 4515 9345 4549
rect 9291 4478 9345 4515
rect 9375 4478 9489 4562
rect 8969 4394 9020 4478
rect 8699 4366 8751 4380
rect 8602 4362 8652 4366
rect 9437 4394 9489 4478
rect 9519 4550 9626 4562
rect 9519 4516 9576 4550
rect 9610 4516 9626 4550
rect 9519 4482 9626 4516
rect 9519 4448 9576 4482
rect 9610 4448 9626 4482
rect 9519 4394 9626 4448
rect 9656 4394 9710 4562
rect 9740 4524 9818 4562
rect 9740 4490 9750 4524
rect 9784 4490 9818 4524
rect 9740 4478 9818 4490
rect 9848 4540 9924 4562
rect 9848 4506 9870 4540
rect 9904 4506 9924 4540
rect 9848 4478 9924 4506
rect 9954 4478 10044 4562
rect 10074 4549 10128 4562
rect 10074 4515 10084 4549
rect 10118 4515 10128 4549
rect 10074 4478 10128 4515
rect 10158 4542 10221 4562
rect 10158 4508 10177 4542
rect 10211 4508 10221 4542
rect 10158 4478 10221 4508
rect 10251 4526 10303 4562
rect 10251 4492 10261 4526
rect 10295 4492 10303 4526
rect 10251 4478 10303 4492
rect 10357 4542 10409 4556
rect 10357 4508 10365 4542
rect 10399 4508 10409 4542
rect 9740 4456 9802 4478
rect 9740 4422 9750 4456
rect 9784 4422 9802 4456
rect 9740 4394 9802 4422
rect 10357 4474 10409 4508
rect 10357 4440 10365 4474
rect 10399 4440 10409 4474
rect 10357 4428 10409 4440
rect 10439 4526 10493 4556
rect 10439 4492 10449 4526
rect 10483 4492 10493 4526
rect 10439 4428 10493 4492
rect 10523 4542 10575 4556
rect 10523 4508 10533 4542
rect 10567 4508 10575 4542
rect 10523 4474 10575 4508
rect 10523 4440 10533 4474
rect 10567 4440 10575 4474
rect 10523 4428 10575 4440
rect 10629 4514 10681 4562
rect 10629 4480 10637 4514
rect 10671 4480 10681 4514
rect 10629 4446 10681 4480
rect 10629 4412 10637 4446
rect 10671 4412 10681 4446
rect 10629 4362 10681 4412
rect 10711 4546 10761 4562
rect 10711 4538 10776 4546
rect 10711 4504 10721 4538
rect 10755 4504 10776 4538
rect 10711 4470 10776 4504
rect 10711 4436 10721 4470
rect 10755 4436 10776 4470
rect 10711 4418 10776 4436
rect 10806 4532 10858 4546
rect 10806 4498 10816 4532
rect 10850 4498 10858 4532
rect 10806 4464 10858 4498
rect 10806 4430 10816 4464
rect 10850 4430 10858 4464
rect 10806 4418 10858 4430
rect 10912 4513 10964 4562
rect 10912 4479 10920 4513
rect 10954 4479 10964 4513
rect 10912 4445 10964 4479
rect 10711 4362 10761 4418
rect 10912 4411 10920 4445
rect 10954 4411 10964 4445
rect 10912 4362 10964 4411
rect 10994 4550 11046 4562
rect 10994 4516 11004 4550
rect 11038 4516 11046 4550
rect 11207 4550 11259 4562
rect 10994 4494 11046 4516
rect 11207 4516 11215 4550
rect 11249 4516 11259 4550
rect 10994 4366 11061 4494
rect 11091 4414 11143 4494
rect 11091 4380 11101 4414
rect 11135 4380 11143 4414
rect 11207 4394 11259 4516
rect 11289 4394 11331 4562
rect 11361 4524 11427 4562
rect 11361 4490 11371 4524
rect 11405 4490 11427 4524
rect 11361 4478 11427 4490
rect 11457 4550 11535 4562
rect 11457 4516 11479 4550
rect 11513 4516 11535 4550
rect 11457 4478 11535 4516
rect 11565 4478 11653 4562
rect 11683 4549 11737 4562
rect 11683 4515 11693 4549
rect 11727 4515 11737 4549
rect 11683 4478 11737 4515
rect 11767 4478 11881 4562
rect 11361 4394 11412 4478
rect 11091 4366 11143 4380
rect 10994 4362 11044 4366
rect 11829 4394 11881 4478
rect 11911 4550 12018 4562
rect 11911 4516 11968 4550
rect 12002 4516 12018 4550
rect 11911 4482 12018 4516
rect 11911 4448 11968 4482
rect 12002 4448 12018 4482
rect 11911 4394 12018 4448
rect 12048 4394 12102 4562
rect 12132 4524 12210 4562
rect 12132 4490 12142 4524
rect 12176 4490 12210 4524
rect 12132 4478 12210 4490
rect 12240 4540 12316 4562
rect 12240 4506 12262 4540
rect 12296 4506 12316 4540
rect 12240 4478 12316 4506
rect 12346 4478 12436 4562
rect 12466 4549 12520 4562
rect 12466 4515 12476 4549
rect 12510 4515 12520 4549
rect 12466 4478 12520 4515
rect 12550 4542 12613 4562
rect 12550 4508 12569 4542
rect 12603 4508 12613 4542
rect 12550 4478 12613 4508
rect 12643 4526 12695 4562
rect 12643 4492 12653 4526
rect 12687 4492 12695 4526
rect 12643 4478 12695 4492
rect 12749 4542 12801 4556
rect 12749 4508 12757 4542
rect 12791 4508 12801 4542
rect 12132 4456 12194 4478
rect 12132 4422 12142 4456
rect 12176 4422 12194 4456
rect 12132 4394 12194 4422
rect 12749 4474 12801 4508
rect 12749 4440 12757 4474
rect 12791 4440 12801 4474
rect 12749 4428 12801 4440
rect 12831 4526 12885 4556
rect 12831 4492 12841 4526
rect 12875 4492 12885 4526
rect 12831 4428 12885 4492
rect 12915 4542 12967 4556
rect 12915 4508 12925 4542
rect 12959 4508 12967 4542
rect 12915 4474 12967 4508
rect 12915 4440 12925 4474
rect 12959 4440 12967 4474
rect 12915 4428 12967 4440
rect 653 3668 705 3688
rect 653 3634 661 3668
rect 695 3634 705 3668
rect 653 3600 705 3634
rect 653 3566 661 3600
rect 695 3566 705 3600
rect 653 3530 705 3566
rect 735 3668 793 3688
rect 735 3634 747 3668
rect 781 3634 793 3668
rect 735 3600 793 3634
rect 735 3566 747 3600
rect 781 3566 793 3600
rect 735 3530 793 3566
rect 823 3668 875 3688
rect 823 3634 833 3668
rect 867 3634 875 3668
rect 823 3587 875 3634
rect 823 3553 833 3587
rect 867 3553 875 3587
rect 823 3530 875 3553
rect 929 3670 981 3688
rect 929 3636 937 3670
rect 971 3636 981 3670
rect 929 3602 981 3636
rect 929 3568 937 3602
rect 971 3568 981 3602
rect 929 3534 981 3568
rect 929 3500 937 3534
rect 971 3500 981 3534
rect 929 3488 981 3500
rect 1011 3676 1065 3688
rect 1011 3642 1021 3676
rect 1055 3642 1065 3676
rect 1011 3608 1065 3642
rect 1011 3574 1021 3608
rect 1055 3574 1065 3608
rect 1011 3488 1065 3574
rect 1095 3654 1149 3688
rect 1095 3620 1105 3654
rect 1139 3620 1149 3654
rect 1095 3559 1149 3620
rect 1095 3525 1105 3559
rect 1139 3525 1149 3559
rect 1095 3488 1149 3525
rect 1179 3676 1233 3688
rect 1179 3642 1189 3676
rect 1223 3642 1233 3676
rect 1179 3608 1233 3642
rect 1179 3574 1189 3608
rect 1223 3574 1233 3608
rect 1179 3488 1233 3574
rect 1263 3654 1317 3688
rect 1263 3620 1273 3654
rect 1307 3620 1317 3654
rect 1263 3559 1317 3620
rect 1263 3525 1273 3559
rect 1307 3525 1317 3559
rect 1263 3488 1317 3525
rect 1347 3676 1399 3688
rect 1347 3642 1357 3676
rect 1391 3642 1399 3676
rect 1347 3608 1399 3642
rect 1347 3574 1357 3608
rect 1391 3574 1399 3608
rect 1347 3540 1399 3574
rect 1347 3506 1357 3540
rect 1391 3506 1399 3540
rect 1347 3488 1399 3506
rect 3236 3677 3288 3689
rect 3236 3643 3244 3677
rect 3278 3643 3288 3677
rect 3236 3609 3288 3643
rect 3236 3575 3244 3609
rect 3278 3575 3288 3609
rect 3236 3541 3288 3575
rect 3236 3507 3244 3541
rect 3278 3507 3288 3541
rect 3236 3489 3288 3507
rect 3318 3677 3370 3689
rect 3318 3643 3328 3677
rect 3362 3643 3370 3677
rect 3318 3609 3370 3643
rect 3318 3575 3328 3609
rect 3362 3575 3370 3609
rect 3318 3541 3370 3575
rect 3452 3669 3504 3683
rect 3452 3635 3460 3669
rect 3494 3635 3504 3669
rect 3452 3601 3504 3635
rect 3452 3567 3460 3601
rect 3494 3567 3504 3601
rect 3452 3555 3504 3567
rect 3534 3653 3588 3683
rect 3534 3619 3544 3653
rect 3578 3619 3588 3653
rect 3534 3555 3588 3619
rect 3618 3669 3670 3683
rect 3618 3635 3628 3669
rect 3662 3635 3670 3669
rect 3618 3601 3670 3635
rect 3724 3653 3776 3689
rect 3724 3619 3732 3653
rect 3766 3619 3776 3653
rect 3724 3605 3776 3619
rect 3806 3669 3869 3689
rect 3806 3635 3816 3669
rect 3850 3635 3869 3669
rect 3806 3605 3869 3635
rect 3899 3676 3953 3689
rect 3899 3642 3909 3676
rect 3943 3642 3953 3676
rect 3899 3605 3953 3642
rect 3983 3605 4073 3689
rect 4103 3667 4179 3689
rect 4103 3633 4123 3667
rect 4157 3633 4179 3667
rect 4103 3605 4179 3633
rect 4209 3651 4287 3689
rect 4209 3617 4243 3651
rect 4277 3617 4287 3651
rect 4209 3605 4287 3617
rect 3618 3567 3628 3601
rect 3662 3567 3670 3601
rect 3618 3555 3670 3567
rect 3318 3507 3328 3541
rect 3362 3507 3370 3541
rect 3318 3489 3370 3507
rect 4225 3583 4287 3605
rect 4225 3549 4243 3583
rect 4277 3549 4287 3583
rect 4225 3521 4287 3549
rect 4317 3521 4371 3689
rect 4401 3677 4508 3689
rect 4401 3643 4417 3677
rect 4451 3643 4508 3677
rect 4401 3609 4508 3643
rect 4401 3575 4417 3609
rect 4451 3575 4508 3609
rect 4401 3521 4508 3575
rect 4538 3605 4652 3689
rect 4682 3676 4736 3689
rect 4682 3642 4692 3676
rect 4726 3642 4736 3676
rect 4682 3605 4736 3642
rect 4766 3605 4854 3689
rect 4884 3677 4962 3689
rect 4884 3643 4906 3677
rect 4940 3643 4962 3677
rect 4884 3605 4962 3643
rect 4992 3651 5058 3689
rect 4992 3617 5014 3651
rect 5048 3617 5058 3651
rect 4992 3605 5058 3617
rect 4538 3521 4590 3605
rect 5007 3521 5058 3605
rect 5088 3521 5130 3689
rect 5160 3677 5212 3689
rect 5160 3643 5170 3677
rect 5204 3643 5212 3677
rect 5373 3677 5425 3689
rect 5160 3521 5212 3643
rect 5373 3643 5381 3677
rect 5415 3643 5425 3677
rect 5373 3621 5425 3643
rect 5276 3541 5328 3621
rect 5276 3507 5284 3541
rect 5318 3507 5328 3541
rect 5276 3493 5328 3507
rect 5358 3493 5425 3621
rect 5375 3489 5425 3493
rect 5455 3640 5507 3689
rect 5658 3673 5708 3689
rect 5455 3606 5465 3640
rect 5499 3606 5507 3640
rect 5455 3572 5507 3606
rect 5455 3538 5465 3572
rect 5499 3538 5507 3572
rect 5561 3659 5613 3673
rect 5561 3625 5569 3659
rect 5603 3625 5613 3659
rect 5561 3591 5613 3625
rect 5561 3557 5569 3591
rect 5603 3557 5613 3591
rect 5561 3545 5613 3557
rect 5643 3665 5708 3673
rect 5643 3631 5664 3665
rect 5698 3631 5708 3665
rect 5643 3597 5708 3631
rect 5643 3563 5664 3597
rect 5698 3563 5708 3597
rect 5643 3545 5708 3563
rect 5455 3489 5507 3538
rect 5658 3489 5708 3545
rect 5738 3641 5790 3689
rect 5738 3607 5748 3641
rect 5782 3607 5790 3641
rect 5738 3573 5790 3607
rect 5738 3539 5748 3573
rect 5782 3539 5790 3573
rect 5844 3669 5896 3683
rect 5844 3635 5852 3669
rect 5886 3635 5896 3669
rect 5844 3601 5896 3635
rect 5844 3567 5852 3601
rect 5886 3567 5896 3601
rect 5844 3555 5896 3567
rect 5926 3653 5980 3683
rect 5926 3619 5936 3653
rect 5970 3619 5980 3653
rect 5926 3555 5980 3619
rect 6010 3669 6062 3683
rect 6010 3635 6020 3669
rect 6054 3635 6062 3669
rect 6010 3601 6062 3635
rect 6116 3653 6168 3689
rect 6116 3619 6124 3653
rect 6158 3619 6168 3653
rect 6116 3605 6168 3619
rect 6198 3669 6261 3689
rect 6198 3635 6208 3669
rect 6242 3635 6261 3669
rect 6198 3605 6261 3635
rect 6291 3676 6345 3689
rect 6291 3642 6301 3676
rect 6335 3642 6345 3676
rect 6291 3605 6345 3642
rect 6375 3605 6465 3689
rect 6495 3667 6571 3689
rect 6495 3633 6515 3667
rect 6549 3633 6571 3667
rect 6495 3605 6571 3633
rect 6601 3651 6679 3689
rect 6601 3617 6635 3651
rect 6669 3617 6679 3651
rect 6601 3605 6679 3617
rect 6010 3567 6020 3601
rect 6054 3567 6062 3601
rect 6010 3555 6062 3567
rect 5738 3489 5790 3539
rect 6617 3583 6679 3605
rect 6617 3549 6635 3583
rect 6669 3549 6679 3583
rect 6617 3521 6679 3549
rect 6709 3521 6763 3689
rect 6793 3677 6900 3689
rect 6793 3643 6809 3677
rect 6843 3643 6900 3677
rect 6793 3609 6900 3643
rect 6793 3575 6809 3609
rect 6843 3575 6900 3609
rect 6793 3521 6900 3575
rect 6930 3605 7044 3689
rect 7074 3676 7128 3689
rect 7074 3642 7084 3676
rect 7118 3642 7128 3676
rect 7074 3605 7128 3642
rect 7158 3605 7246 3689
rect 7276 3677 7354 3689
rect 7276 3643 7298 3677
rect 7332 3643 7354 3677
rect 7276 3605 7354 3643
rect 7384 3651 7450 3689
rect 7384 3617 7406 3651
rect 7440 3617 7450 3651
rect 7384 3605 7450 3617
rect 6930 3521 6982 3605
rect 7399 3521 7450 3605
rect 7480 3521 7522 3689
rect 7552 3677 7604 3689
rect 7552 3643 7562 3677
rect 7596 3643 7604 3677
rect 7765 3677 7817 3689
rect 7552 3521 7604 3643
rect 7765 3643 7773 3677
rect 7807 3643 7817 3677
rect 7765 3621 7817 3643
rect 7668 3541 7720 3621
rect 7668 3507 7676 3541
rect 7710 3507 7720 3541
rect 7668 3493 7720 3507
rect 7750 3493 7817 3621
rect 7767 3489 7817 3493
rect 7847 3640 7899 3689
rect 8050 3673 8100 3689
rect 7847 3606 7857 3640
rect 7891 3606 7899 3640
rect 7847 3572 7899 3606
rect 7847 3538 7857 3572
rect 7891 3538 7899 3572
rect 7953 3659 8005 3673
rect 7953 3625 7961 3659
rect 7995 3625 8005 3659
rect 7953 3591 8005 3625
rect 7953 3557 7961 3591
rect 7995 3557 8005 3591
rect 7953 3545 8005 3557
rect 8035 3665 8100 3673
rect 8035 3631 8056 3665
rect 8090 3631 8100 3665
rect 8035 3597 8100 3631
rect 8035 3563 8056 3597
rect 8090 3563 8100 3597
rect 8035 3545 8100 3563
rect 7847 3489 7899 3538
rect 8050 3489 8100 3545
rect 8130 3641 8182 3689
rect 8130 3607 8140 3641
rect 8174 3607 8182 3641
rect 8130 3573 8182 3607
rect 8130 3539 8140 3573
rect 8174 3539 8182 3573
rect 8236 3669 8288 3683
rect 8236 3635 8244 3669
rect 8278 3635 8288 3669
rect 8236 3601 8288 3635
rect 8236 3567 8244 3601
rect 8278 3567 8288 3601
rect 8236 3555 8288 3567
rect 8318 3653 8372 3683
rect 8318 3619 8328 3653
rect 8362 3619 8372 3653
rect 8318 3555 8372 3619
rect 8402 3669 8454 3683
rect 8402 3635 8412 3669
rect 8446 3635 8454 3669
rect 8402 3601 8454 3635
rect 8508 3653 8560 3689
rect 8508 3619 8516 3653
rect 8550 3619 8560 3653
rect 8508 3605 8560 3619
rect 8590 3669 8653 3689
rect 8590 3635 8600 3669
rect 8634 3635 8653 3669
rect 8590 3605 8653 3635
rect 8683 3676 8737 3689
rect 8683 3642 8693 3676
rect 8727 3642 8737 3676
rect 8683 3605 8737 3642
rect 8767 3605 8857 3689
rect 8887 3667 8963 3689
rect 8887 3633 8907 3667
rect 8941 3633 8963 3667
rect 8887 3605 8963 3633
rect 8993 3651 9071 3689
rect 8993 3617 9027 3651
rect 9061 3617 9071 3651
rect 8993 3605 9071 3617
rect 8402 3567 8412 3601
rect 8446 3567 8454 3601
rect 8402 3555 8454 3567
rect 8130 3489 8182 3539
rect 9009 3583 9071 3605
rect 9009 3549 9027 3583
rect 9061 3549 9071 3583
rect 9009 3521 9071 3549
rect 9101 3521 9155 3689
rect 9185 3677 9292 3689
rect 9185 3643 9201 3677
rect 9235 3643 9292 3677
rect 9185 3609 9292 3643
rect 9185 3575 9201 3609
rect 9235 3575 9292 3609
rect 9185 3521 9292 3575
rect 9322 3605 9436 3689
rect 9466 3676 9520 3689
rect 9466 3642 9476 3676
rect 9510 3642 9520 3676
rect 9466 3605 9520 3642
rect 9550 3605 9638 3689
rect 9668 3677 9746 3689
rect 9668 3643 9690 3677
rect 9724 3643 9746 3677
rect 9668 3605 9746 3643
rect 9776 3651 9842 3689
rect 9776 3617 9798 3651
rect 9832 3617 9842 3651
rect 9776 3605 9842 3617
rect 9322 3521 9374 3605
rect 9791 3521 9842 3605
rect 9872 3521 9914 3689
rect 9944 3677 9996 3689
rect 9944 3643 9954 3677
rect 9988 3643 9996 3677
rect 10157 3677 10209 3689
rect 9944 3521 9996 3643
rect 10157 3643 10165 3677
rect 10199 3643 10209 3677
rect 10157 3621 10209 3643
rect 10060 3541 10112 3621
rect 10060 3507 10068 3541
rect 10102 3507 10112 3541
rect 10060 3493 10112 3507
rect 10142 3493 10209 3621
rect 10159 3489 10209 3493
rect 10239 3640 10291 3689
rect 10442 3673 10492 3689
rect 10239 3606 10249 3640
rect 10283 3606 10291 3640
rect 10239 3572 10291 3606
rect 10239 3538 10249 3572
rect 10283 3538 10291 3572
rect 10345 3659 10397 3673
rect 10345 3625 10353 3659
rect 10387 3625 10397 3659
rect 10345 3591 10397 3625
rect 10345 3557 10353 3591
rect 10387 3557 10397 3591
rect 10345 3545 10397 3557
rect 10427 3665 10492 3673
rect 10427 3631 10448 3665
rect 10482 3631 10492 3665
rect 10427 3597 10492 3631
rect 10427 3563 10448 3597
rect 10482 3563 10492 3597
rect 10427 3545 10492 3563
rect 10239 3489 10291 3538
rect 10442 3489 10492 3545
rect 10522 3641 10574 3689
rect 10522 3607 10532 3641
rect 10566 3607 10574 3641
rect 10522 3573 10574 3607
rect 10522 3539 10532 3573
rect 10566 3539 10574 3573
rect 10628 3669 10680 3683
rect 10628 3635 10636 3669
rect 10670 3635 10680 3669
rect 10628 3601 10680 3635
rect 10628 3567 10636 3601
rect 10670 3567 10680 3601
rect 10628 3555 10680 3567
rect 10710 3653 10764 3683
rect 10710 3619 10720 3653
rect 10754 3619 10764 3653
rect 10710 3555 10764 3619
rect 10794 3669 10846 3683
rect 10794 3635 10804 3669
rect 10838 3635 10846 3669
rect 10794 3601 10846 3635
rect 10900 3653 10952 3689
rect 10900 3619 10908 3653
rect 10942 3619 10952 3653
rect 10900 3605 10952 3619
rect 10982 3669 11045 3689
rect 10982 3635 10992 3669
rect 11026 3635 11045 3669
rect 10982 3605 11045 3635
rect 11075 3676 11129 3689
rect 11075 3642 11085 3676
rect 11119 3642 11129 3676
rect 11075 3605 11129 3642
rect 11159 3605 11249 3689
rect 11279 3667 11355 3689
rect 11279 3633 11299 3667
rect 11333 3633 11355 3667
rect 11279 3605 11355 3633
rect 11385 3651 11463 3689
rect 11385 3617 11419 3651
rect 11453 3617 11463 3651
rect 11385 3605 11463 3617
rect 10794 3567 10804 3601
rect 10838 3567 10846 3601
rect 10794 3555 10846 3567
rect 10522 3489 10574 3539
rect 11401 3583 11463 3605
rect 11401 3549 11419 3583
rect 11453 3549 11463 3583
rect 11401 3521 11463 3549
rect 11493 3521 11547 3689
rect 11577 3677 11684 3689
rect 11577 3643 11593 3677
rect 11627 3643 11684 3677
rect 11577 3609 11684 3643
rect 11577 3575 11593 3609
rect 11627 3575 11684 3609
rect 11577 3521 11684 3575
rect 11714 3605 11828 3689
rect 11858 3676 11912 3689
rect 11858 3642 11868 3676
rect 11902 3642 11912 3676
rect 11858 3605 11912 3642
rect 11942 3605 12030 3689
rect 12060 3677 12138 3689
rect 12060 3643 12082 3677
rect 12116 3643 12138 3677
rect 12060 3605 12138 3643
rect 12168 3651 12234 3689
rect 12168 3617 12190 3651
rect 12224 3617 12234 3651
rect 12168 3605 12234 3617
rect 11714 3521 11766 3605
rect 12183 3521 12234 3605
rect 12264 3521 12306 3689
rect 12336 3677 12388 3689
rect 12336 3643 12346 3677
rect 12380 3643 12388 3677
rect 12549 3677 12601 3689
rect 12336 3521 12388 3643
rect 12549 3643 12557 3677
rect 12591 3643 12601 3677
rect 12549 3621 12601 3643
rect 12452 3541 12504 3621
rect 12452 3507 12460 3541
rect 12494 3507 12504 3541
rect 12452 3493 12504 3507
rect 12534 3493 12601 3621
rect 12551 3489 12601 3493
rect 12631 3640 12683 3689
rect 12834 3673 12884 3689
rect 12631 3606 12641 3640
rect 12675 3606 12683 3640
rect 12631 3572 12683 3606
rect 12631 3538 12641 3572
rect 12675 3538 12683 3572
rect 12737 3659 12789 3673
rect 12737 3625 12745 3659
rect 12779 3625 12789 3659
rect 12737 3591 12789 3625
rect 12737 3557 12745 3591
rect 12779 3557 12789 3591
rect 12737 3545 12789 3557
rect 12819 3665 12884 3673
rect 12819 3631 12840 3665
rect 12874 3631 12884 3665
rect 12819 3597 12884 3631
rect 12819 3563 12840 3597
rect 12874 3563 12884 3597
rect 12819 3545 12884 3563
rect 12631 3489 12683 3538
rect 12834 3489 12884 3545
rect 12914 3641 12966 3689
rect 12914 3607 12924 3641
rect 12958 3607 12966 3641
rect 12914 3573 12966 3607
rect 12914 3539 12924 3573
rect 12958 3539 12966 3573
rect 12914 3489 12966 3539
rect 1060 2768 1112 2816
rect 1060 2734 1068 2768
rect 1102 2734 1112 2768
rect 1060 2700 1112 2734
rect 1060 2666 1068 2700
rect 1102 2666 1112 2700
rect 1060 2616 1112 2666
rect 1142 2800 1192 2816
rect 1142 2792 1207 2800
rect 1142 2758 1152 2792
rect 1186 2758 1207 2792
rect 1142 2724 1207 2758
rect 1142 2690 1152 2724
rect 1186 2690 1207 2724
rect 1142 2672 1207 2690
rect 1237 2786 1289 2800
rect 1237 2752 1247 2786
rect 1281 2752 1289 2786
rect 1237 2718 1289 2752
rect 1237 2684 1247 2718
rect 1281 2684 1289 2718
rect 1237 2672 1289 2684
rect 1343 2767 1395 2816
rect 1343 2733 1351 2767
rect 1385 2733 1395 2767
rect 1343 2699 1395 2733
rect 1142 2616 1192 2672
rect 1343 2665 1351 2699
rect 1385 2665 1395 2699
rect 1343 2616 1395 2665
rect 1425 2804 1477 2816
rect 1425 2770 1435 2804
rect 1469 2770 1477 2804
rect 1638 2804 1690 2816
rect 1425 2748 1477 2770
rect 1638 2770 1646 2804
rect 1680 2770 1690 2804
rect 1425 2620 1492 2748
rect 1522 2668 1574 2748
rect 1522 2634 1532 2668
rect 1566 2634 1574 2668
rect 1638 2648 1690 2770
rect 1720 2648 1762 2816
rect 1792 2778 1858 2816
rect 1792 2744 1802 2778
rect 1836 2744 1858 2778
rect 1792 2732 1858 2744
rect 1888 2804 1966 2816
rect 1888 2770 1910 2804
rect 1944 2770 1966 2804
rect 1888 2732 1966 2770
rect 1996 2732 2084 2816
rect 2114 2803 2168 2816
rect 2114 2769 2124 2803
rect 2158 2769 2168 2803
rect 2114 2732 2168 2769
rect 2198 2732 2312 2816
rect 1792 2648 1843 2732
rect 1522 2620 1574 2634
rect 1425 2616 1475 2620
rect 2260 2648 2312 2732
rect 2342 2804 2449 2816
rect 2342 2770 2399 2804
rect 2433 2770 2449 2804
rect 2342 2736 2449 2770
rect 2342 2702 2399 2736
rect 2433 2702 2449 2736
rect 2342 2648 2449 2702
rect 2479 2648 2533 2816
rect 2563 2778 2641 2816
rect 2563 2744 2573 2778
rect 2607 2744 2641 2778
rect 2563 2732 2641 2744
rect 2671 2794 2747 2816
rect 2671 2760 2693 2794
rect 2727 2760 2747 2794
rect 2671 2732 2747 2760
rect 2777 2732 2867 2816
rect 2897 2803 2951 2816
rect 2897 2769 2907 2803
rect 2941 2769 2951 2803
rect 2897 2732 2951 2769
rect 2981 2796 3044 2816
rect 2981 2762 3000 2796
rect 3034 2762 3044 2796
rect 2981 2732 3044 2762
rect 3074 2780 3126 2816
rect 3074 2746 3084 2780
rect 3118 2746 3126 2780
rect 3074 2732 3126 2746
rect 3180 2796 3232 2810
rect 3180 2762 3188 2796
rect 3222 2762 3232 2796
rect 2563 2710 2625 2732
rect 2563 2676 2573 2710
rect 2607 2676 2625 2710
rect 2563 2648 2625 2676
rect 3180 2728 3232 2762
rect 3180 2694 3188 2728
rect 3222 2694 3232 2728
rect 3180 2682 3232 2694
rect 3262 2780 3316 2810
rect 3262 2746 3272 2780
rect 3306 2746 3316 2780
rect 3262 2682 3316 2746
rect 3346 2796 3398 2810
rect 3346 2762 3356 2796
rect 3390 2762 3398 2796
rect 3346 2728 3398 2762
rect 3346 2694 3356 2728
rect 3390 2694 3398 2728
rect 3346 2682 3398 2694
rect 3452 2768 3504 2816
rect 3452 2734 3460 2768
rect 3494 2734 3504 2768
rect 3452 2700 3504 2734
rect 3452 2666 3460 2700
rect 3494 2666 3504 2700
rect 3452 2616 3504 2666
rect 3534 2800 3584 2816
rect 3534 2792 3599 2800
rect 3534 2758 3544 2792
rect 3578 2758 3599 2792
rect 3534 2724 3599 2758
rect 3534 2690 3544 2724
rect 3578 2690 3599 2724
rect 3534 2672 3599 2690
rect 3629 2786 3681 2800
rect 3629 2752 3639 2786
rect 3673 2752 3681 2786
rect 3629 2718 3681 2752
rect 3629 2684 3639 2718
rect 3673 2684 3681 2718
rect 3629 2672 3681 2684
rect 3735 2767 3787 2816
rect 3735 2733 3743 2767
rect 3777 2733 3787 2767
rect 3735 2699 3787 2733
rect 3534 2616 3584 2672
rect 3735 2665 3743 2699
rect 3777 2665 3787 2699
rect 3735 2616 3787 2665
rect 3817 2804 3869 2816
rect 3817 2770 3827 2804
rect 3861 2770 3869 2804
rect 4030 2804 4082 2816
rect 3817 2748 3869 2770
rect 4030 2770 4038 2804
rect 4072 2770 4082 2804
rect 3817 2620 3884 2748
rect 3914 2668 3966 2748
rect 3914 2634 3924 2668
rect 3958 2634 3966 2668
rect 4030 2648 4082 2770
rect 4112 2648 4154 2816
rect 4184 2778 4250 2816
rect 4184 2744 4194 2778
rect 4228 2744 4250 2778
rect 4184 2732 4250 2744
rect 4280 2804 4358 2816
rect 4280 2770 4302 2804
rect 4336 2770 4358 2804
rect 4280 2732 4358 2770
rect 4388 2732 4476 2816
rect 4506 2803 4560 2816
rect 4506 2769 4516 2803
rect 4550 2769 4560 2803
rect 4506 2732 4560 2769
rect 4590 2732 4704 2816
rect 4184 2648 4235 2732
rect 3914 2620 3966 2634
rect 3817 2616 3867 2620
rect 4652 2648 4704 2732
rect 4734 2804 4841 2816
rect 4734 2770 4791 2804
rect 4825 2770 4841 2804
rect 4734 2736 4841 2770
rect 4734 2702 4791 2736
rect 4825 2702 4841 2736
rect 4734 2648 4841 2702
rect 4871 2648 4925 2816
rect 4955 2778 5033 2816
rect 4955 2744 4965 2778
rect 4999 2744 5033 2778
rect 4955 2732 5033 2744
rect 5063 2794 5139 2816
rect 5063 2760 5085 2794
rect 5119 2760 5139 2794
rect 5063 2732 5139 2760
rect 5169 2732 5259 2816
rect 5289 2803 5343 2816
rect 5289 2769 5299 2803
rect 5333 2769 5343 2803
rect 5289 2732 5343 2769
rect 5373 2796 5436 2816
rect 5373 2762 5392 2796
rect 5426 2762 5436 2796
rect 5373 2732 5436 2762
rect 5466 2780 5518 2816
rect 5466 2746 5476 2780
rect 5510 2746 5518 2780
rect 5466 2732 5518 2746
rect 5572 2796 5624 2810
rect 5572 2762 5580 2796
rect 5614 2762 5624 2796
rect 4955 2710 5017 2732
rect 4955 2676 4965 2710
rect 4999 2676 5017 2710
rect 4955 2648 5017 2676
rect 5572 2728 5624 2762
rect 5572 2694 5580 2728
rect 5614 2694 5624 2728
rect 5572 2682 5624 2694
rect 5654 2780 5708 2810
rect 5654 2746 5664 2780
rect 5698 2746 5708 2780
rect 5654 2682 5708 2746
rect 5738 2796 5790 2810
rect 5738 2762 5748 2796
rect 5782 2762 5790 2796
rect 5738 2728 5790 2762
rect 5738 2694 5748 2728
rect 5782 2694 5790 2728
rect 5738 2682 5790 2694
rect 5844 2768 5896 2816
rect 5844 2734 5852 2768
rect 5886 2734 5896 2768
rect 5844 2700 5896 2734
rect 5844 2666 5852 2700
rect 5886 2666 5896 2700
rect 5844 2616 5896 2666
rect 5926 2800 5976 2816
rect 5926 2792 5991 2800
rect 5926 2758 5936 2792
rect 5970 2758 5991 2792
rect 5926 2724 5991 2758
rect 5926 2690 5936 2724
rect 5970 2690 5991 2724
rect 5926 2672 5991 2690
rect 6021 2786 6073 2800
rect 6021 2752 6031 2786
rect 6065 2752 6073 2786
rect 6021 2718 6073 2752
rect 6021 2684 6031 2718
rect 6065 2684 6073 2718
rect 6021 2672 6073 2684
rect 6127 2767 6179 2816
rect 6127 2733 6135 2767
rect 6169 2733 6179 2767
rect 6127 2699 6179 2733
rect 5926 2616 5976 2672
rect 6127 2665 6135 2699
rect 6169 2665 6179 2699
rect 6127 2616 6179 2665
rect 6209 2804 6261 2816
rect 6209 2770 6219 2804
rect 6253 2770 6261 2804
rect 6422 2804 6474 2816
rect 6209 2748 6261 2770
rect 6422 2770 6430 2804
rect 6464 2770 6474 2804
rect 6209 2620 6276 2748
rect 6306 2668 6358 2748
rect 6306 2634 6316 2668
rect 6350 2634 6358 2668
rect 6422 2648 6474 2770
rect 6504 2648 6546 2816
rect 6576 2778 6642 2816
rect 6576 2744 6586 2778
rect 6620 2744 6642 2778
rect 6576 2732 6642 2744
rect 6672 2804 6750 2816
rect 6672 2770 6694 2804
rect 6728 2770 6750 2804
rect 6672 2732 6750 2770
rect 6780 2732 6868 2816
rect 6898 2803 6952 2816
rect 6898 2769 6908 2803
rect 6942 2769 6952 2803
rect 6898 2732 6952 2769
rect 6982 2732 7096 2816
rect 6576 2648 6627 2732
rect 6306 2620 6358 2634
rect 6209 2616 6259 2620
rect 7044 2648 7096 2732
rect 7126 2804 7233 2816
rect 7126 2770 7183 2804
rect 7217 2770 7233 2804
rect 7126 2736 7233 2770
rect 7126 2702 7183 2736
rect 7217 2702 7233 2736
rect 7126 2648 7233 2702
rect 7263 2648 7317 2816
rect 7347 2778 7425 2816
rect 7347 2744 7357 2778
rect 7391 2744 7425 2778
rect 7347 2732 7425 2744
rect 7455 2794 7531 2816
rect 7455 2760 7477 2794
rect 7511 2760 7531 2794
rect 7455 2732 7531 2760
rect 7561 2732 7651 2816
rect 7681 2803 7735 2816
rect 7681 2769 7691 2803
rect 7725 2769 7735 2803
rect 7681 2732 7735 2769
rect 7765 2796 7828 2816
rect 7765 2762 7784 2796
rect 7818 2762 7828 2796
rect 7765 2732 7828 2762
rect 7858 2780 7910 2816
rect 7858 2746 7868 2780
rect 7902 2746 7910 2780
rect 7858 2732 7910 2746
rect 7964 2796 8016 2810
rect 7964 2762 7972 2796
rect 8006 2762 8016 2796
rect 7347 2710 7409 2732
rect 7347 2676 7357 2710
rect 7391 2676 7409 2710
rect 7347 2648 7409 2676
rect 7964 2728 8016 2762
rect 7964 2694 7972 2728
rect 8006 2694 8016 2728
rect 7964 2682 8016 2694
rect 8046 2780 8100 2810
rect 8046 2746 8056 2780
rect 8090 2746 8100 2780
rect 8046 2682 8100 2746
rect 8130 2796 8182 2810
rect 8130 2762 8140 2796
rect 8174 2762 8182 2796
rect 8130 2728 8182 2762
rect 8130 2694 8140 2728
rect 8174 2694 8182 2728
rect 8130 2682 8182 2694
rect 8236 2768 8288 2816
rect 8236 2734 8244 2768
rect 8278 2734 8288 2768
rect 8236 2700 8288 2734
rect 8236 2666 8244 2700
rect 8278 2666 8288 2700
rect 8236 2616 8288 2666
rect 8318 2800 8368 2816
rect 8318 2792 8383 2800
rect 8318 2758 8328 2792
rect 8362 2758 8383 2792
rect 8318 2724 8383 2758
rect 8318 2690 8328 2724
rect 8362 2690 8383 2724
rect 8318 2672 8383 2690
rect 8413 2786 8465 2800
rect 8413 2752 8423 2786
rect 8457 2752 8465 2786
rect 8413 2718 8465 2752
rect 8413 2684 8423 2718
rect 8457 2684 8465 2718
rect 8413 2672 8465 2684
rect 8519 2767 8571 2816
rect 8519 2733 8527 2767
rect 8561 2733 8571 2767
rect 8519 2699 8571 2733
rect 8318 2616 8368 2672
rect 8519 2665 8527 2699
rect 8561 2665 8571 2699
rect 8519 2616 8571 2665
rect 8601 2804 8653 2816
rect 8601 2770 8611 2804
rect 8645 2770 8653 2804
rect 8814 2804 8866 2816
rect 8601 2748 8653 2770
rect 8814 2770 8822 2804
rect 8856 2770 8866 2804
rect 8601 2620 8668 2748
rect 8698 2668 8750 2748
rect 8698 2634 8708 2668
rect 8742 2634 8750 2668
rect 8814 2648 8866 2770
rect 8896 2648 8938 2816
rect 8968 2778 9034 2816
rect 8968 2744 8978 2778
rect 9012 2744 9034 2778
rect 8968 2732 9034 2744
rect 9064 2804 9142 2816
rect 9064 2770 9086 2804
rect 9120 2770 9142 2804
rect 9064 2732 9142 2770
rect 9172 2732 9260 2816
rect 9290 2803 9344 2816
rect 9290 2769 9300 2803
rect 9334 2769 9344 2803
rect 9290 2732 9344 2769
rect 9374 2732 9488 2816
rect 8968 2648 9019 2732
rect 8698 2620 8750 2634
rect 8601 2616 8651 2620
rect 9436 2648 9488 2732
rect 9518 2804 9625 2816
rect 9518 2770 9575 2804
rect 9609 2770 9625 2804
rect 9518 2736 9625 2770
rect 9518 2702 9575 2736
rect 9609 2702 9625 2736
rect 9518 2648 9625 2702
rect 9655 2648 9709 2816
rect 9739 2778 9817 2816
rect 9739 2744 9749 2778
rect 9783 2744 9817 2778
rect 9739 2732 9817 2744
rect 9847 2794 9923 2816
rect 9847 2760 9869 2794
rect 9903 2760 9923 2794
rect 9847 2732 9923 2760
rect 9953 2732 10043 2816
rect 10073 2803 10127 2816
rect 10073 2769 10083 2803
rect 10117 2769 10127 2803
rect 10073 2732 10127 2769
rect 10157 2796 10220 2816
rect 10157 2762 10176 2796
rect 10210 2762 10220 2796
rect 10157 2732 10220 2762
rect 10250 2780 10302 2816
rect 10250 2746 10260 2780
rect 10294 2746 10302 2780
rect 10250 2732 10302 2746
rect 10356 2796 10408 2810
rect 10356 2762 10364 2796
rect 10398 2762 10408 2796
rect 9739 2710 9801 2732
rect 9739 2676 9749 2710
rect 9783 2676 9801 2710
rect 9739 2648 9801 2676
rect 10356 2728 10408 2762
rect 10356 2694 10364 2728
rect 10398 2694 10408 2728
rect 10356 2682 10408 2694
rect 10438 2780 10492 2810
rect 10438 2746 10448 2780
rect 10482 2746 10492 2780
rect 10438 2682 10492 2746
rect 10522 2796 10574 2810
rect 10522 2762 10532 2796
rect 10566 2762 10574 2796
rect 10522 2728 10574 2762
rect 10522 2694 10532 2728
rect 10566 2694 10574 2728
rect 10522 2682 10574 2694
rect 10628 2768 10680 2816
rect 10628 2734 10636 2768
rect 10670 2734 10680 2768
rect 10628 2700 10680 2734
rect 10628 2666 10636 2700
rect 10670 2666 10680 2700
rect 10628 2616 10680 2666
rect 10710 2800 10760 2816
rect 10710 2792 10775 2800
rect 10710 2758 10720 2792
rect 10754 2758 10775 2792
rect 10710 2724 10775 2758
rect 10710 2690 10720 2724
rect 10754 2690 10775 2724
rect 10710 2672 10775 2690
rect 10805 2786 10857 2800
rect 10805 2752 10815 2786
rect 10849 2752 10857 2786
rect 10805 2718 10857 2752
rect 10805 2684 10815 2718
rect 10849 2684 10857 2718
rect 10805 2672 10857 2684
rect 10911 2767 10963 2816
rect 10911 2733 10919 2767
rect 10953 2733 10963 2767
rect 10911 2699 10963 2733
rect 10710 2616 10760 2672
rect 10911 2665 10919 2699
rect 10953 2665 10963 2699
rect 10911 2616 10963 2665
rect 10993 2804 11045 2816
rect 10993 2770 11003 2804
rect 11037 2770 11045 2804
rect 11206 2804 11258 2816
rect 10993 2748 11045 2770
rect 11206 2770 11214 2804
rect 11248 2770 11258 2804
rect 10993 2620 11060 2748
rect 11090 2668 11142 2748
rect 11090 2634 11100 2668
rect 11134 2634 11142 2668
rect 11206 2648 11258 2770
rect 11288 2648 11330 2816
rect 11360 2778 11426 2816
rect 11360 2744 11370 2778
rect 11404 2744 11426 2778
rect 11360 2732 11426 2744
rect 11456 2804 11534 2816
rect 11456 2770 11478 2804
rect 11512 2770 11534 2804
rect 11456 2732 11534 2770
rect 11564 2732 11652 2816
rect 11682 2803 11736 2816
rect 11682 2769 11692 2803
rect 11726 2769 11736 2803
rect 11682 2732 11736 2769
rect 11766 2732 11880 2816
rect 11360 2648 11411 2732
rect 11090 2620 11142 2634
rect 10993 2616 11043 2620
rect 11828 2648 11880 2732
rect 11910 2804 12017 2816
rect 11910 2770 11967 2804
rect 12001 2770 12017 2804
rect 11910 2736 12017 2770
rect 11910 2702 11967 2736
rect 12001 2702 12017 2736
rect 11910 2648 12017 2702
rect 12047 2648 12101 2816
rect 12131 2778 12209 2816
rect 12131 2744 12141 2778
rect 12175 2744 12209 2778
rect 12131 2732 12209 2744
rect 12239 2794 12315 2816
rect 12239 2760 12261 2794
rect 12295 2760 12315 2794
rect 12239 2732 12315 2760
rect 12345 2732 12435 2816
rect 12465 2803 12519 2816
rect 12465 2769 12475 2803
rect 12509 2769 12519 2803
rect 12465 2732 12519 2769
rect 12549 2796 12612 2816
rect 12549 2762 12568 2796
rect 12602 2762 12612 2796
rect 12549 2732 12612 2762
rect 12642 2780 12694 2816
rect 12642 2746 12652 2780
rect 12686 2746 12694 2780
rect 12642 2732 12694 2746
rect 12748 2796 12800 2810
rect 12748 2762 12756 2796
rect 12790 2762 12800 2796
rect 12131 2710 12193 2732
rect 12131 2676 12141 2710
rect 12175 2676 12193 2710
rect 12131 2648 12193 2676
rect 12748 2728 12800 2762
rect 12748 2694 12756 2728
rect 12790 2694 12800 2728
rect 12748 2682 12800 2694
rect 12830 2780 12884 2810
rect 12830 2746 12840 2780
rect 12874 2746 12884 2780
rect 12830 2682 12884 2746
rect 12914 2796 12966 2810
rect 12914 2762 12924 2796
rect 12958 2762 12966 2796
rect 12914 2728 12966 2762
rect 12914 2694 12924 2728
rect 12958 2694 12966 2728
rect 12914 2682 12966 2694
<< ndiffc >>
rect 1070 5699 1104 5733
rect 1156 5686 1190 5720
rect 1242 5716 1276 5750
rect 1346 5722 1380 5756
rect 1430 5690 1464 5724
rect 1514 5722 1548 5756
rect 1598 5690 1632 5724
rect 1682 5722 1716 5756
rect 1766 5754 1800 5788
rect 1766 5686 1800 5720
rect 2330 5754 2364 5788
rect 2330 5686 2364 5720
rect 2429 5722 2463 5756
rect 2513 5754 2547 5788
rect 2513 5686 2547 5720
rect 2613 5722 2647 5756
rect 2697 5712 2731 5746
rect 2906 5686 2940 5720
rect 3110 5686 3144 5720
rect 3214 5694 3248 5728
rect 3298 5712 3332 5746
rect 3383 5712 3417 5746
rect 3487 5686 3521 5720
rect 3586 5686 3620 5720
rect 3790 5700 3824 5734
rect 3982 5686 4016 5720
rect 4066 5712 4100 5746
rect 1069 4839 1103 4873
rect 1153 4813 1187 4847
rect 1237 4839 1271 4873
rect 1341 4813 1375 4847
rect 1425 4831 1459 4865
rect 1531 4813 1565 4847
rect 1748 4809 1782 4843
rect 1832 4829 1866 4863
rect 1932 4873 1966 4907
rect 2016 4847 2050 4881
rect 2120 4813 2154 4847
rect 2314 4813 2348 4847
rect 2505 4809 2539 4843
rect 2607 4829 2641 4863
rect 2707 4873 2741 4907
rect 2791 4821 2825 4855
rect 2895 4823 2929 4857
rect 2990 4813 3024 4847
rect 3074 4847 3108 4881
rect 3178 4839 3212 4873
rect 3273 4813 3307 4847
rect 3357 4849 3391 4883
rect 3461 4839 3495 4873
rect 3545 4813 3579 4847
rect 3629 4839 3663 4873
rect 3733 4813 3767 4847
rect 3817 4831 3851 4865
rect 3923 4813 3957 4847
rect 4140 4809 4174 4843
rect 4224 4829 4258 4863
rect 4324 4873 4358 4907
rect 4408 4847 4442 4881
rect 4512 4813 4546 4847
rect 4706 4813 4740 4847
rect 4897 4809 4931 4843
rect 4999 4829 5033 4863
rect 5099 4873 5133 4907
rect 5183 4821 5217 4855
rect 5287 4823 5321 4857
rect 5382 4813 5416 4847
rect 5466 4847 5500 4881
rect 5570 4839 5604 4873
rect 5665 4813 5699 4847
rect 5749 4849 5783 4883
rect 5853 4839 5887 4873
rect 5937 4813 5971 4847
rect 6021 4839 6055 4873
rect 6125 4813 6159 4847
rect 6209 4831 6243 4865
rect 6315 4813 6349 4847
rect 6532 4809 6566 4843
rect 6616 4829 6650 4863
rect 6716 4873 6750 4907
rect 6800 4847 6834 4881
rect 6904 4813 6938 4847
rect 7098 4813 7132 4847
rect 7289 4809 7323 4843
rect 7391 4829 7425 4863
rect 7491 4873 7525 4907
rect 7575 4821 7609 4855
rect 7679 4823 7713 4857
rect 7774 4813 7808 4847
rect 7858 4847 7892 4881
rect 7962 4839 7996 4873
rect 8057 4813 8091 4847
rect 8141 4849 8175 4883
rect 8245 4839 8279 4873
rect 8329 4813 8363 4847
rect 8413 4839 8447 4873
rect 8517 4813 8551 4847
rect 8601 4831 8635 4865
rect 8707 4813 8741 4847
rect 8924 4809 8958 4843
rect 9008 4829 9042 4863
rect 9108 4873 9142 4907
rect 9192 4847 9226 4881
rect 9296 4813 9330 4847
rect 9490 4813 9524 4847
rect 9681 4809 9715 4843
rect 9783 4829 9817 4863
rect 9883 4873 9917 4907
rect 9967 4821 10001 4855
rect 10071 4823 10105 4857
rect 10166 4813 10200 4847
rect 10250 4847 10284 4881
rect 10354 4839 10388 4873
rect 10449 4813 10483 4847
rect 10533 4849 10567 4883
rect 10637 4839 10671 4873
rect 10721 4813 10755 4847
rect 10805 4839 10839 4873
rect 10909 4813 10943 4847
rect 10993 4831 11027 4865
rect 11099 4813 11133 4847
rect 11316 4809 11350 4843
rect 11400 4829 11434 4863
rect 11500 4873 11534 4907
rect 11584 4847 11618 4881
rect 11688 4813 11722 4847
rect 11882 4813 11916 4847
rect 12073 4809 12107 4843
rect 12175 4829 12209 4863
rect 12275 4873 12309 4907
rect 12359 4821 12393 4855
rect 12463 4823 12497 4857
rect 12558 4813 12592 4847
rect 12642 4847 12676 4881
rect 12746 4839 12780 4873
rect 12841 4813 12875 4847
rect 12925 4849 12959 4883
rect 629 4137 663 4171
rect 715 4124 749 4158
rect 801 4154 835 4188
rect 905 4160 939 4194
rect 989 4128 1023 4162
rect 1073 4160 1107 4194
rect 1157 4128 1191 4162
rect 1241 4160 1275 4194
rect 1325 4192 1359 4226
rect 1325 4124 1359 4158
rect 1437 4196 1471 4230
rect 1437 4128 1471 4162
rect 1521 4196 1555 4230
rect 1521 4128 1555 4162
rect 1605 4128 1639 4162
rect 1689 4196 1723 4230
rect 1689 4128 1723 4162
rect 1773 4128 1807 4162
rect 1857 4196 1891 4230
rect 1857 4128 1891 4162
rect 1941 4128 1975 4162
rect 2025 4196 2059 4230
rect 2025 4128 2059 4162
rect 2109 4128 2143 4162
rect 2193 4196 2227 4230
rect 2193 4128 2227 4162
rect 2277 4128 2311 4162
rect 2361 4196 2395 4230
rect 2361 4128 2395 4162
rect 2445 4128 2479 4162
rect 2529 4196 2563 4230
rect 2529 4128 2563 4162
rect 2613 4128 2647 4162
rect 2697 4196 2731 4230
rect 2697 4128 2731 4162
rect 2781 4128 2815 4162
rect 2865 4196 2899 4230
rect 2865 4128 2899 4162
rect 2949 4128 2983 4162
rect 3033 4196 3067 4230
rect 3033 4128 3067 4162
rect 3117 4128 3151 4162
rect 3201 4196 3235 4230
rect 3201 4128 3235 4162
rect 3285 4128 3319 4162
rect 3461 4160 3495 4194
rect 3545 4124 3579 4158
rect 3640 4150 3674 4184
rect 3744 4158 3778 4192
rect 3828 4124 3862 4158
rect 3923 4134 3957 4168
rect 4027 4132 4061 4166
rect 4111 4184 4145 4218
rect 4211 4140 4245 4174
rect 4313 4120 4347 4154
rect 4504 4124 4538 4158
rect 4698 4124 4732 4158
rect 4802 4158 4836 4192
rect 4886 4184 4920 4218
rect 4986 4140 5020 4174
rect 5070 4120 5104 4154
rect 5287 4124 5321 4158
rect 5393 4142 5427 4176
rect 5477 4124 5511 4158
rect 5581 4150 5615 4184
rect 5665 4124 5699 4158
rect 5749 4150 5783 4184
rect 5853 4160 5887 4194
rect 5937 4124 5971 4158
rect 6032 4150 6066 4184
rect 6136 4158 6170 4192
rect 6220 4124 6254 4158
rect 6315 4134 6349 4168
rect 6419 4132 6453 4166
rect 6503 4184 6537 4218
rect 6603 4140 6637 4174
rect 6705 4120 6739 4154
rect 6896 4124 6930 4158
rect 7090 4124 7124 4158
rect 7194 4158 7228 4192
rect 7278 4184 7312 4218
rect 7378 4140 7412 4174
rect 7462 4120 7496 4154
rect 7679 4124 7713 4158
rect 7785 4142 7819 4176
rect 7869 4124 7903 4158
rect 7973 4150 8007 4184
rect 8057 4124 8091 4158
rect 8141 4150 8175 4184
rect 8245 4160 8279 4194
rect 8329 4124 8363 4158
rect 8424 4150 8458 4184
rect 8528 4158 8562 4192
rect 8612 4124 8646 4158
rect 8707 4134 8741 4168
rect 8811 4132 8845 4166
rect 8895 4184 8929 4218
rect 8995 4140 9029 4174
rect 9097 4120 9131 4154
rect 9288 4124 9322 4158
rect 9482 4124 9516 4158
rect 9586 4158 9620 4192
rect 9670 4184 9704 4218
rect 9770 4140 9804 4174
rect 9854 4120 9888 4154
rect 10071 4124 10105 4158
rect 10177 4142 10211 4176
rect 10261 4124 10295 4158
rect 10365 4150 10399 4184
rect 10449 4124 10483 4158
rect 10533 4150 10567 4184
rect 10637 4160 10671 4194
rect 10721 4124 10755 4158
rect 10816 4150 10850 4184
rect 10920 4158 10954 4192
rect 11004 4124 11038 4158
rect 11099 4134 11133 4168
rect 11203 4132 11237 4166
rect 11287 4184 11321 4218
rect 11387 4140 11421 4174
rect 11489 4120 11523 4154
rect 11680 4124 11714 4158
rect 11874 4124 11908 4158
rect 11978 4158 12012 4192
rect 12062 4184 12096 4218
rect 12162 4140 12196 4174
rect 12246 4120 12280 4154
rect 12463 4124 12497 4158
rect 12569 4142 12603 4176
rect 12653 4124 12687 4158
rect 12757 4150 12791 4184
rect 12841 4124 12875 4158
rect 12925 4150 12959 4184
rect 661 3263 695 3297
rect 747 3250 781 3284
rect 833 3280 867 3314
rect 937 3286 971 3320
rect 1021 3254 1055 3288
rect 1105 3286 1139 3320
rect 1189 3254 1223 3288
rect 1273 3286 1307 3320
rect 1357 3318 1391 3352
rect 1357 3250 1391 3284
rect 3244 3323 3278 3357
rect 3244 3255 3278 3289
rect 3328 3323 3362 3357
rect 3328 3255 3362 3289
rect 3460 3277 3494 3311
rect 3544 3251 3578 3285
rect 3628 3277 3662 3311
rect 3732 3251 3766 3285
rect 3816 3269 3850 3303
rect 3922 3251 3956 3285
rect 4139 3247 4173 3281
rect 4223 3267 4257 3301
rect 4323 3311 4357 3345
rect 4407 3285 4441 3319
rect 4511 3251 4545 3285
rect 4705 3251 4739 3285
rect 4896 3247 4930 3281
rect 4998 3267 5032 3301
rect 5098 3311 5132 3345
rect 5182 3259 5216 3293
rect 5286 3261 5320 3295
rect 5381 3251 5415 3285
rect 5465 3285 5499 3319
rect 5569 3277 5603 3311
rect 5664 3251 5698 3285
rect 5748 3287 5782 3321
rect 5852 3277 5886 3311
rect 5936 3251 5970 3285
rect 6020 3277 6054 3311
rect 6124 3251 6158 3285
rect 6208 3269 6242 3303
rect 6314 3251 6348 3285
rect 6531 3247 6565 3281
rect 6615 3267 6649 3301
rect 6715 3311 6749 3345
rect 6799 3285 6833 3319
rect 6903 3251 6937 3285
rect 7097 3251 7131 3285
rect 7288 3247 7322 3281
rect 7390 3267 7424 3301
rect 7490 3311 7524 3345
rect 7574 3259 7608 3293
rect 7678 3261 7712 3295
rect 7773 3251 7807 3285
rect 7857 3285 7891 3319
rect 7961 3277 7995 3311
rect 8056 3251 8090 3285
rect 8140 3287 8174 3321
rect 8244 3277 8278 3311
rect 8328 3251 8362 3285
rect 8412 3277 8446 3311
rect 8516 3251 8550 3285
rect 8600 3269 8634 3303
rect 8706 3251 8740 3285
rect 8923 3247 8957 3281
rect 9007 3267 9041 3301
rect 9107 3311 9141 3345
rect 9191 3285 9225 3319
rect 9295 3251 9329 3285
rect 9489 3251 9523 3285
rect 9680 3247 9714 3281
rect 9782 3267 9816 3301
rect 9882 3311 9916 3345
rect 9966 3259 10000 3293
rect 10070 3261 10104 3295
rect 10165 3251 10199 3285
rect 10249 3285 10283 3319
rect 10353 3277 10387 3311
rect 10448 3251 10482 3285
rect 10532 3287 10566 3321
rect 10636 3277 10670 3311
rect 10720 3251 10754 3285
rect 10804 3277 10838 3311
rect 10908 3251 10942 3285
rect 10992 3269 11026 3303
rect 11098 3251 11132 3285
rect 11315 3247 11349 3281
rect 11399 3267 11433 3301
rect 11499 3311 11533 3345
rect 11583 3285 11617 3319
rect 11687 3251 11721 3285
rect 11881 3251 11915 3285
rect 12072 3247 12106 3281
rect 12174 3267 12208 3301
rect 12274 3311 12308 3345
rect 12358 3259 12392 3293
rect 12462 3261 12496 3295
rect 12557 3251 12591 3285
rect 12641 3285 12675 3319
rect 12745 3277 12779 3311
rect 12840 3251 12874 3285
rect 12924 3287 12958 3321
rect 1068 2414 1102 2448
rect 1152 2378 1186 2412
rect 1247 2404 1281 2438
rect 1351 2412 1385 2446
rect 1435 2378 1469 2412
rect 1530 2388 1564 2422
rect 1634 2386 1668 2420
rect 1718 2438 1752 2472
rect 1818 2394 1852 2428
rect 1920 2374 1954 2408
rect 2111 2378 2145 2412
rect 2305 2378 2339 2412
rect 2409 2412 2443 2446
rect 2493 2438 2527 2472
rect 2593 2394 2627 2428
rect 2677 2374 2711 2408
rect 2894 2378 2928 2412
rect 3000 2396 3034 2430
rect 3084 2378 3118 2412
rect 3188 2404 3222 2438
rect 3272 2378 3306 2412
rect 3356 2404 3390 2438
rect 3460 2414 3494 2448
rect 3544 2378 3578 2412
rect 3639 2404 3673 2438
rect 3743 2412 3777 2446
rect 3827 2378 3861 2412
rect 3922 2388 3956 2422
rect 4026 2386 4060 2420
rect 4110 2438 4144 2472
rect 4210 2394 4244 2428
rect 4312 2374 4346 2408
rect 4503 2378 4537 2412
rect 4697 2378 4731 2412
rect 4801 2412 4835 2446
rect 4885 2438 4919 2472
rect 4985 2394 5019 2428
rect 5069 2374 5103 2408
rect 5286 2378 5320 2412
rect 5392 2396 5426 2430
rect 5476 2378 5510 2412
rect 5580 2404 5614 2438
rect 5664 2378 5698 2412
rect 5748 2404 5782 2438
rect 5852 2414 5886 2448
rect 5936 2378 5970 2412
rect 6031 2404 6065 2438
rect 6135 2412 6169 2446
rect 6219 2378 6253 2412
rect 6314 2388 6348 2422
rect 6418 2386 6452 2420
rect 6502 2438 6536 2472
rect 6602 2394 6636 2428
rect 6704 2374 6738 2408
rect 6895 2378 6929 2412
rect 7089 2378 7123 2412
rect 7193 2412 7227 2446
rect 7277 2438 7311 2472
rect 7377 2394 7411 2428
rect 7461 2374 7495 2408
rect 7678 2378 7712 2412
rect 7784 2396 7818 2430
rect 7868 2378 7902 2412
rect 7972 2404 8006 2438
rect 8056 2378 8090 2412
rect 8140 2404 8174 2438
rect 8244 2414 8278 2448
rect 8328 2378 8362 2412
rect 8423 2404 8457 2438
rect 8527 2412 8561 2446
rect 8611 2378 8645 2412
rect 8706 2388 8740 2422
rect 8810 2386 8844 2420
rect 8894 2438 8928 2472
rect 8994 2394 9028 2428
rect 9096 2374 9130 2408
rect 9287 2378 9321 2412
rect 9481 2378 9515 2412
rect 9585 2412 9619 2446
rect 9669 2438 9703 2472
rect 9769 2394 9803 2428
rect 9853 2374 9887 2408
rect 10070 2378 10104 2412
rect 10176 2396 10210 2430
rect 10260 2378 10294 2412
rect 10364 2404 10398 2438
rect 10448 2378 10482 2412
rect 10532 2404 10566 2438
rect 10636 2414 10670 2448
rect 10720 2378 10754 2412
rect 10815 2404 10849 2438
rect 10919 2412 10953 2446
rect 11003 2378 11037 2412
rect 11098 2388 11132 2422
rect 11202 2386 11236 2420
rect 11286 2438 11320 2472
rect 11386 2394 11420 2428
rect 11488 2374 11522 2408
rect 11679 2378 11713 2412
rect 11873 2378 11907 2412
rect 11977 2412 12011 2446
rect 12061 2438 12095 2472
rect 12161 2394 12195 2428
rect 12245 2374 12279 2408
rect 12462 2378 12496 2412
rect 12568 2396 12602 2430
rect 12652 2378 12686 2412
rect 12756 2404 12790 2438
rect 12840 2378 12874 2412
rect 12924 2404 12958 2438
<< pdiffc >>
rect 1070 6070 1104 6104
rect 1070 6002 1104 6036
rect 1156 6070 1190 6104
rect 1156 6002 1190 6036
rect 1242 6070 1276 6104
rect 1242 5989 1276 6023
rect 1346 6072 1380 6106
rect 1346 6004 1380 6038
rect 1346 5936 1380 5970
rect 1430 6078 1464 6112
rect 1430 6010 1464 6044
rect 1514 6056 1548 6090
rect 1514 5961 1548 5995
rect 1598 6078 1632 6112
rect 1598 6010 1632 6044
rect 1682 6056 1716 6090
rect 1682 5961 1716 5995
rect 1766 6078 1800 6112
rect 1766 6010 1800 6044
rect 1766 5942 1800 5976
rect 2330 6078 2364 6112
rect 2330 6010 2364 6044
rect 2330 5942 2364 5976
rect 2429 6068 2463 6102
rect 2429 5942 2463 5976
rect 2513 6078 2547 6112
rect 2513 6010 2547 6044
rect 2513 5942 2547 5976
rect 2613 6068 2647 6102
rect 2613 5994 2647 6028
rect 2697 6078 2731 6112
rect 2697 6010 2731 6044
rect 2895 6058 2929 6092
rect 3114 6044 3148 6078
rect 3218 5956 3252 5990
rect 3302 5955 3336 5989
rect 3386 6005 3420 6039
rect 3490 5984 3524 6018
rect 3574 6054 3608 6088
rect 3802 6052 3836 6086
rect 3982 6078 4016 6112
rect 4066 6052 4100 6086
rect 1069 5197 1103 5231
rect 1069 5129 1103 5163
rect 1153 5181 1187 5215
rect 1237 5197 1271 5231
rect 1341 5181 1375 5215
rect 1425 5197 1459 5231
rect 1518 5204 1552 5238
rect 1732 5195 1766 5229
rect 1852 5179 1886 5213
rect 1237 5129 1271 5163
rect 1852 5111 1886 5145
rect 2026 5205 2060 5239
rect 2026 5137 2060 5171
rect 2301 5204 2335 5238
rect 2515 5205 2549 5239
rect 2623 5179 2657 5213
rect 2779 5205 2813 5239
rect 2990 5205 3024 5239
rect 2893 5069 2927 5103
rect 3074 5168 3108 5202
rect 3074 5100 3108 5134
rect 3178 5187 3212 5221
rect 3178 5119 3212 5153
rect 3273 5193 3307 5227
rect 3273 5125 3307 5159
rect 3357 5169 3391 5203
rect 3357 5101 3391 5135
rect 3461 5197 3495 5231
rect 3461 5129 3495 5163
rect 3545 5181 3579 5215
rect 3629 5197 3663 5231
rect 3733 5181 3767 5215
rect 3817 5197 3851 5231
rect 3910 5204 3944 5238
rect 4124 5195 4158 5229
rect 4244 5179 4278 5213
rect 3629 5129 3663 5163
rect 4244 5111 4278 5145
rect 4418 5205 4452 5239
rect 4418 5137 4452 5171
rect 4693 5204 4727 5238
rect 4907 5205 4941 5239
rect 5015 5179 5049 5213
rect 5171 5205 5205 5239
rect 5382 5205 5416 5239
rect 5285 5069 5319 5103
rect 5466 5168 5500 5202
rect 5466 5100 5500 5134
rect 5570 5187 5604 5221
rect 5570 5119 5604 5153
rect 5665 5193 5699 5227
rect 5665 5125 5699 5159
rect 5749 5169 5783 5203
rect 5749 5101 5783 5135
rect 5853 5197 5887 5231
rect 5853 5129 5887 5163
rect 5937 5181 5971 5215
rect 6021 5197 6055 5231
rect 6125 5181 6159 5215
rect 6209 5197 6243 5231
rect 6302 5204 6336 5238
rect 6516 5195 6550 5229
rect 6636 5179 6670 5213
rect 6021 5129 6055 5163
rect 6636 5111 6670 5145
rect 6810 5205 6844 5239
rect 6810 5137 6844 5171
rect 7085 5204 7119 5238
rect 7299 5205 7333 5239
rect 7407 5179 7441 5213
rect 7563 5205 7597 5239
rect 7774 5205 7808 5239
rect 7677 5069 7711 5103
rect 7858 5168 7892 5202
rect 7858 5100 7892 5134
rect 7962 5187 7996 5221
rect 7962 5119 7996 5153
rect 8057 5193 8091 5227
rect 8057 5125 8091 5159
rect 8141 5169 8175 5203
rect 8141 5101 8175 5135
rect 8245 5197 8279 5231
rect 8245 5129 8279 5163
rect 8329 5181 8363 5215
rect 8413 5197 8447 5231
rect 8517 5181 8551 5215
rect 8601 5197 8635 5231
rect 8694 5204 8728 5238
rect 8908 5195 8942 5229
rect 9028 5179 9062 5213
rect 8413 5129 8447 5163
rect 9028 5111 9062 5145
rect 9202 5205 9236 5239
rect 9202 5137 9236 5171
rect 9477 5204 9511 5238
rect 9691 5205 9725 5239
rect 9799 5179 9833 5213
rect 9955 5205 9989 5239
rect 10166 5205 10200 5239
rect 10069 5069 10103 5103
rect 10250 5168 10284 5202
rect 10250 5100 10284 5134
rect 10354 5187 10388 5221
rect 10354 5119 10388 5153
rect 10449 5193 10483 5227
rect 10449 5125 10483 5159
rect 10533 5169 10567 5203
rect 10533 5101 10567 5135
rect 10637 5197 10671 5231
rect 10637 5129 10671 5163
rect 10721 5181 10755 5215
rect 10805 5197 10839 5231
rect 10909 5181 10943 5215
rect 10993 5197 11027 5231
rect 11086 5204 11120 5238
rect 11300 5195 11334 5229
rect 11420 5179 11454 5213
rect 10805 5129 10839 5163
rect 11420 5111 11454 5145
rect 11594 5205 11628 5239
rect 11594 5137 11628 5171
rect 11869 5204 11903 5238
rect 12083 5205 12117 5239
rect 12191 5179 12225 5213
rect 12347 5205 12381 5239
rect 12558 5205 12592 5239
rect 12461 5069 12495 5103
rect 12642 5168 12676 5202
rect 12642 5100 12676 5134
rect 12746 5187 12780 5221
rect 12746 5119 12780 5153
rect 12841 5193 12875 5227
rect 12841 5125 12875 5159
rect 12925 5169 12959 5203
rect 12925 5101 12959 5135
rect 629 4508 663 4542
rect 629 4440 663 4474
rect 715 4508 749 4542
rect 715 4440 749 4474
rect 801 4508 835 4542
rect 801 4427 835 4461
rect 905 4510 939 4544
rect 905 4442 939 4476
rect 905 4374 939 4408
rect 989 4516 1023 4550
rect 989 4448 1023 4482
rect 1073 4494 1107 4528
rect 1073 4399 1107 4433
rect 1157 4516 1191 4550
rect 1157 4448 1191 4482
rect 1241 4494 1275 4528
rect 1241 4399 1275 4433
rect 1325 4516 1359 4550
rect 1325 4448 1359 4482
rect 1325 4380 1359 4414
rect 1437 4516 1471 4550
rect 1437 4448 1471 4482
rect 1437 4380 1471 4414
rect 1521 4510 1555 4544
rect 1521 4442 1555 4476
rect 1521 4374 1555 4408
rect 1605 4516 1639 4550
rect 1605 4448 1639 4482
rect 1689 4510 1723 4544
rect 1689 4442 1723 4476
rect 1689 4374 1723 4408
rect 1773 4516 1807 4550
rect 1773 4448 1807 4482
rect 1857 4510 1891 4544
rect 1857 4442 1891 4476
rect 1857 4374 1891 4408
rect 1941 4516 1975 4550
rect 1941 4448 1975 4482
rect 2025 4510 2059 4544
rect 2025 4442 2059 4476
rect 2025 4374 2059 4408
rect 2109 4516 2143 4550
rect 2109 4448 2143 4482
rect 2193 4510 2227 4544
rect 2193 4442 2227 4476
rect 2193 4374 2227 4408
rect 2277 4516 2311 4550
rect 2277 4448 2311 4482
rect 2361 4510 2395 4544
rect 2361 4442 2395 4476
rect 2361 4374 2395 4408
rect 2445 4516 2479 4550
rect 2445 4448 2479 4482
rect 2529 4510 2563 4544
rect 2529 4442 2563 4476
rect 2529 4374 2563 4408
rect 2613 4516 2647 4550
rect 2613 4448 2647 4482
rect 2697 4510 2731 4544
rect 2697 4442 2731 4476
rect 2697 4374 2731 4408
rect 2781 4516 2815 4550
rect 2781 4448 2815 4482
rect 2865 4510 2899 4544
rect 2865 4442 2899 4476
rect 2865 4374 2899 4408
rect 2949 4516 2983 4550
rect 2949 4448 2983 4482
rect 3033 4510 3067 4544
rect 3033 4442 3067 4476
rect 3033 4374 3067 4408
rect 3117 4516 3151 4550
rect 3117 4448 3151 4482
rect 3201 4510 3235 4544
rect 3201 4442 3235 4476
rect 3201 4374 3235 4408
rect 3285 4516 3319 4550
rect 3285 4448 3319 4482
rect 3461 4480 3495 4514
rect 3461 4412 3495 4446
rect 3545 4504 3579 4538
rect 3545 4436 3579 4470
rect 3640 4498 3674 4532
rect 3640 4430 3674 4464
rect 3744 4479 3778 4513
rect 3744 4411 3778 4445
rect 3828 4516 3862 4550
rect 4039 4516 4073 4550
rect 3925 4380 3959 4414
rect 4195 4490 4229 4524
rect 4303 4516 4337 4550
rect 4517 4515 4551 4549
rect 4792 4516 4826 4550
rect 4792 4448 4826 4482
rect 4966 4490 5000 4524
rect 5086 4506 5120 4540
rect 5300 4515 5334 4549
rect 5393 4508 5427 4542
rect 5477 4492 5511 4526
rect 5581 4508 5615 4542
rect 4966 4422 5000 4456
rect 5581 4440 5615 4474
rect 5665 4492 5699 4526
rect 5749 4508 5783 4542
rect 5749 4440 5783 4474
rect 5853 4480 5887 4514
rect 5853 4412 5887 4446
rect 5937 4504 5971 4538
rect 5937 4436 5971 4470
rect 6032 4498 6066 4532
rect 6032 4430 6066 4464
rect 6136 4479 6170 4513
rect 6136 4411 6170 4445
rect 6220 4516 6254 4550
rect 6431 4516 6465 4550
rect 6317 4380 6351 4414
rect 6587 4490 6621 4524
rect 6695 4516 6729 4550
rect 6909 4515 6943 4549
rect 7184 4516 7218 4550
rect 7184 4448 7218 4482
rect 7358 4490 7392 4524
rect 7478 4506 7512 4540
rect 7692 4515 7726 4549
rect 7785 4508 7819 4542
rect 7869 4492 7903 4526
rect 7973 4508 8007 4542
rect 7358 4422 7392 4456
rect 7973 4440 8007 4474
rect 8057 4492 8091 4526
rect 8141 4508 8175 4542
rect 8141 4440 8175 4474
rect 8245 4480 8279 4514
rect 8245 4412 8279 4446
rect 8329 4504 8363 4538
rect 8329 4436 8363 4470
rect 8424 4498 8458 4532
rect 8424 4430 8458 4464
rect 8528 4479 8562 4513
rect 8528 4411 8562 4445
rect 8612 4516 8646 4550
rect 8823 4516 8857 4550
rect 8709 4380 8743 4414
rect 8979 4490 9013 4524
rect 9087 4516 9121 4550
rect 9301 4515 9335 4549
rect 9576 4516 9610 4550
rect 9576 4448 9610 4482
rect 9750 4490 9784 4524
rect 9870 4506 9904 4540
rect 10084 4515 10118 4549
rect 10177 4508 10211 4542
rect 10261 4492 10295 4526
rect 10365 4508 10399 4542
rect 9750 4422 9784 4456
rect 10365 4440 10399 4474
rect 10449 4492 10483 4526
rect 10533 4508 10567 4542
rect 10533 4440 10567 4474
rect 10637 4480 10671 4514
rect 10637 4412 10671 4446
rect 10721 4504 10755 4538
rect 10721 4436 10755 4470
rect 10816 4498 10850 4532
rect 10816 4430 10850 4464
rect 10920 4479 10954 4513
rect 10920 4411 10954 4445
rect 11004 4516 11038 4550
rect 11215 4516 11249 4550
rect 11101 4380 11135 4414
rect 11371 4490 11405 4524
rect 11479 4516 11513 4550
rect 11693 4515 11727 4549
rect 11968 4516 12002 4550
rect 11968 4448 12002 4482
rect 12142 4490 12176 4524
rect 12262 4506 12296 4540
rect 12476 4515 12510 4549
rect 12569 4508 12603 4542
rect 12653 4492 12687 4526
rect 12757 4508 12791 4542
rect 12142 4422 12176 4456
rect 12757 4440 12791 4474
rect 12841 4492 12875 4526
rect 12925 4508 12959 4542
rect 12925 4440 12959 4474
rect 661 3634 695 3668
rect 661 3566 695 3600
rect 747 3634 781 3668
rect 747 3566 781 3600
rect 833 3634 867 3668
rect 833 3553 867 3587
rect 937 3636 971 3670
rect 937 3568 971 3602
rect 937 3500 971 3534
rect 1021 3642 1055 3676
rect 1021 3574 1055 3608
rect 1105 3620 1139 3654
rect 1105 3525 1139 3559
rect 1189 3642 1223 3676
rect 1189 3574 1223 3608
rect 1273 3620 1307 3654
rect 1273 3525 1307 3559
rect 1357 3642 1391 3676
rect 1357 3574 1391 3608
rect 1357 3506 1391 3540
rect 3244 3643 3278 3677
rect 3244 3575 3278 3609
rect 3244 3507 3278 3541
rect 3328 3643 3362 3677
rect 3328 3575 3362 3609
rect 3460 3635 3494 3669
rect 3460 3567 3494 3601
rect 3544 3619 3578 3653
rect 3628 3635 3662 3669
rect 3732 3619 3766 3653
rect 3816 3635 3850 3669
rect 3909 3642 3943 3676
rect 4123 3633 4157 3667
rect 4243 3617 4277 3651
rect 3628 3567 3662 3601
rect 3328 3507 3362 3541
rect 4243 3549 4277 3583
rect 4417 3643 4451 3677
rect 4417 3575 4451 3609
rect 4692 3642 4726 3676
rect 4906 3643 4940 3677
rect 5014 3617 5048 3651
rect 5170 3643 5204 3677
rect 5381 3643 5415 3677
rect 5284 3507 5318 3541
rect 5465 3606 5499 3640
rect 5465 3538 5499 3572
rect 5569 3625 5603 3659
rect 5569 3557 5603 3591
rect 5664 3631 5698 3665
rect 5664 3563 5698 3597
rect 5748 3607 5782 3641
rect 5748 3539 5782 3573
rect 5852 3635 5886 3669
rect 5852 3567 5886 3601
rect 5936 3619 5970 3653
rect 6020 3635 6054 3669
rect 6124 3619 6158 3653
rect 6208 3635 6242 3669
rect 6301 3642 6335 3676
rect 6515 3633 6549 3667
rect 6635 3617 6669 3651
rect 6020 3567 6054 3601
rect 6635 3549 6669 3583
rect 6809 3643 6843 3677
rect 6809 3575 6843 3609
rect 7084 3642 7118 3676
rect 7298 3643 7332 3677
rect 7406 3617 7440 3651
rect 7562 3643 7596 3677
rect 7773 3643 7807 3677
rect 7676 3507 7710 3541
rect 7857 3606 7891 3640
rect 7857 3538 7891 3572
rect 7961 3625 7995 3659
rect 7961 3557 7995 3591
rect 8056 3631 8090 3665
rect 8056 3563 8090 3597
rect 8140 3607 8174 3641
rect 8140 3539 8174 3573
rect 8244 3635 8278 3669
rect 8244 3567 8278 3601
rect 8328 3619 8362 3653
rect 8412 3635 8446 3669
rect 8516 3619 8550 3653
rect 8600 3635 8634 3669
rect 8693 3642 8727 3676
rect 8907 3633 8941 3667
rect 9027 3617 9061 3651
rect 8412 3567 8446 3601
rect 9027 3549 9061 3583
rect 9201 3643 9235 3677
rect 9201 3575 9235 3609
rect 9476 3642 9510 3676
rect 9690 3643 9724 3677
rect 9798 3617 9832 3651
rect 9954 3643 9988 3677
rect 10165 3643 10199 3677
rect 10068 3507 10102 3541
rect 10249 3606 10283 3640
rect 10249 3538 10283 3572
rect 10353 3625 10387 3659
rect 10353 3557 10387 3591
rect 10448 3631 10482 3665
rect 10448 3563 10482 3597
rect 10532 3607 10566 3641
rect 10532 3539 10566 3573
rect 10636 3635 10670 3669
rect 10636 3567 10670 3601
rect 10720 3619 10754 3653
rect 10804 3635 10838 3669
rect 10908 3619 10942 3653
rect 10992 3635 11026 3669
rect 11085 3642 11119 3676
rect 11299 3633 11333 3667
rect 11419 3617 11453 3651
rect 10804 3567 10838 3601
rect 11419 3549 11453 3583
rect 11593 3643 11627 3677
rect 11593 3575 11627 3609
rect 11868 3642 11902 3676
rect 12082 3643 12116 3677
rect 12190 3617 12224 3651
rect 12346 3643 12380 3677
rect 12557 3643 12591 3677
rect 12460 3507 12494 3541
rect 12641 3606 12675 3640
rect 12641 3538 12675 3572
rect 12745 3625 12779 3659
rect 12745 3557 12779 3591
rect 12840 3631 12874 3665
rect 12840 3563 12874 3597
rect 12924 3607 12958 3641
rect 12924 3539 12958 3573
rect 1068 2734 1102 2768
rect 1068 2666 1102 2700
rect 1152 2758 1186 2792
rect 1152 2690 1186 2724
rect 1247 2752 1281 2786
rect 1247 2684 1281 2718
rect 1351 2733 1385 2767
rect 1351 2665 1385 2699
rect 1435 2770 1469 2804
rect 1646 2770 1680 2804
rect 1532 2634 1566 2668
rect 1802 2744 1836 2778
rect 1910 2770 1944 2804
rect 2124 2769 2158 2803
rect 2399 2770 2433 2804
rect 2399 2702 2433 2736
rect 2573 2744 2607 2778
rect 2693 2760 2727 2794
rect 2907 2769 2941 2803
rect 3000 2762 3034 2796
rect 3084 2746 3118 2780
rect 3188 2762 3222 2796
rect 2573 2676 2607 2710
rect 3188 2694 3222 2728
rect 3272 2746 3306 2780
rect 3356 2762 3390 2796
rect 3356 2694 3390 2728
rect 3460 2734 3494 2768
rect 3460 2666 3494 2700
rect 3544 2758 3578 2792
rect 3544 2690 3578 2724
rect 3639 2752 3673 2786
rect 3639 2684 3673 2718
rect 3743 2733 3777 2767
rect 3743 2665 3777 2699
rect 3827 2770 3861 2804
rect 4038 2770 4072 2804
rect 3924 2634 3958 2668
rect 4194 2744 4228 2778
rect 4302 2770 4336 2804
rect 4516 2769 4550 2803
rect 4791 2770 4825 2804
rect 4791 2702 4825 2736
rect 4965 2744 4999 2778
rect 5085 2760 5119 2794
rect 5299 2769 5333 2803
rect 5392 2762 5426 2796
rect 5476 2746 5510 2780
rect 5580 2762 5614 2796
rect 4965 2676 4999 2710
rect 5580 2694 5614 2728
rect 5664 2746 5698 2780
rect 5748 2762 5782 2796
rect 5748 2694 5782 2728
rect 5852 2734 5886 2768
rect 5852 2666 5886 2700
rect 5936 2758 5970 2792
rect 5936 2690 5970 2724
rect 6031 2752 6065 2786
rect 6031 2684 6065 2718
rect 6135 2733 6169 2767
rect 6135 2665 6169 2699
rect 6219 2770 6253 2804
rect 6430 2770 6464 2804
rect 6316 2634 6350 2668
rect 6586 2744 6620 2778
rect 6694 2770 6728 2804
rect 6908 2769 6942 2803
rect 7183 2770 7217 2804
rect 7183 2702 7217 2736
rect 7357 2744 7391 2778
rect 7477 2760 7511 2794
rect 7691 2769 7725 2803
rect 7784 2762 7818 2796
rect 7868 2746 7902 2780
rect 7972 2762 8006 2796
rect 7357 2676 7391 2710
rect 7972 2694 8006 2728
rect 8056 2746 8090 2780
rect 8140 2762 8174 2796
rect 8140 2694 8174 2728
rect 8244 2734 8278 2768
rect 8244 2666 8278 2700
rect 8328 2758 8362 2792
rect 8328 2690 8362 2724
rect 8423 2752 8457 2786
rect 8423 2684 8457 2718
rect 8527 2733 8561 2767
rect 8527 2665 8561 2699
rect 8611 2770 8645 2804
rect 8822 2770 8856 2804
rect 8708 2634 8742 2668
rect 8978 2744 9012 2778
rect 9086 2770 9120 2804
rect 9300 2769 9334 2803
rect 9575 2770 9609 2804
rect 9575 2702 9609 2736
rect 9749 2744 9783 2778
rect 9869 2760 9903 2794
rect 10083 2769 10117 2803
rect 10176 2762 10210 2796
rect 10260 2746 10294 2780
rect 10364 2762 10398 2796
rect 9749 2676 9783 2710
rect 10364 2694 10398 2728
rect 10448 2746 10482 2780
rect 10532 2762 10566 2796
rect 10532 2694 10566 2728
rect 10636 2734 10670 2768
rect 10636 2666 10670 2700
rect 10720 2758 10754 2792
rect 10720 2690 10754 2724
rect 10815 2752 10849 2786
rect 10815 2684 10849 2718
rect 10919 2733 10953 2767
rect 10919 2665 10953 2699
rect 11003 2770 11037 2804
rect 11214 2770 11248 2804
rect 11100 2634 11134 2668
rect 11370 2744 11404 2778
rect 11478 2770 11512 2804
rect 11692 2769 11726 2803
rect 11967 2770 12001 2804
rect 11967 2702 12001 2736
rect 12141 2744 12175 2778
rect 12261 2760 12295 2794
rect 12475 2769 12509 2803
rect 12568 2762 12602 2796
rect 12652 2746 12686 2780
rect 12756 2762 12790 2796
rect 12141 2676 12175 2710
rect 12756 2694 12790 2728
rect 12840 2746 12874 2780
rect 12924 2762 12958 2796
rect 12924 2694 12958 2728
<< psubdiff >>
rect 1035 5586 1064 5620
rect 1098 5586 1156 5620
rect 1190 5586 1248 5620
rect 1282 5586 1340 5620
rect 1374 5586 1432 5620
rect 1466 5586 1524 5620
rect 1558 5586 1616 5620
rect 1650 5586 1708 5620
rect 1742 5586 1800 5620
rect 1834 5586 1892 5620
rect 1926 5586 1984 5620
rect 2018 5586 2076 5620
rect 2110 5586 2168 5620
rect 2202 5586 2260 5620
rect 2294 5586 2352 5620
rect 2386 5586 2444 5620
rect 2478 5586 2536 5620
rect 2570 5586 2628 5620
rect 2662 5586 2720 5620
rect 2754 5586 2812 5620
rect 2846 5586 2904 5620
rect 2938 5586 2996 5620
rect 3030 5586 3088 5620
rect 3122 5586 3180 5620
rect 3214 5586 3272 5620
rect 3306 5586 3364 5620
rect 3398 5586 3456 5620
rect 3490 5586 3548 5620
rect 3582 5586 3640 5620
rect 3674 5586 3732 5620
rect 3766 5586 3824 5620
rect 3858 5586 3916 5620
rect 3950 5586 4008 5620
rect 4042 5586 4135 5620
rect 1034 4713 1063 4747
rect 1097 4713 1155 4747
rect 1189 4713 1247 4747
rect 1281 4713 1339 4747
rect 1373 4713 1431 4747
rect 1465 4713 1523 4747
rect 1557 4713 1615 4747
rect 1649 4713 1707 4747
rect 1741 4713 1799 4747
rect 1833 4713 1891 4747
rect 1925 4713 1983 4747
rect 2017 4713 2075 4747
rect 2109 4713 2167 4747
rect 2201 4713 2259 4747
rect 2293 4713 2351 4747
rect 2385 4713 2443 4747
rect 2477 4713 2535 4747
rect 2569 4713 2627 4747
rect 2661 4713 2719 4747
rect 2753 4713 2811 4747
rect 2845 4713 2903 4747
rect 2937 4713 2995 4747
rect 3029 4713 3087 4747
rect 3121 4713 3179 4747
rect 3213 4713 3271 4747
rect 3305 4713 3363 4747
rect 3397 4713 3455 4747
rect 3489 4713 3547 4747
rect 3581 4713 3639 4747
rect 3673 4713 3731 4747
rect 3765 4713 3823 4747
rect 3857 4713 3915 4747
rect 3949 4713 4007 4747
rect 4041 4713 4099 4747
rect 4133 4713 4191 4747
rect 4225 4713 4283 4747
rect 4317 4713 4375 4747
rect 4409 4713 4467 4747
rect 4501 4713 4559 4747
rect 4593 4713 4651 4747
rect 4685 4713 4743 4747
rect 4777 4713 4835 4747
rect 4869 4713 4927 4747
rect 4961 4713 5019 4747
rect 5053 4713 5111 4747
rect 5145 4713 5203 4747
rect 5237 4713 5295 4747
rect 5329 4713 5387 4747
rect 5421 4713 5479 4747
rect 5513 4713 5571 4747
rect 5605 4713 5663 4747
rect 5697 4713 5755 4747
rect 5789 4713 5847 4747
rect 5881 4713 5939 4747
rect 5973 4713 6031 4747
rect 6065 4713 6123 4747
rect 6157 4713 6215 4747
rect 6249 4713 6307 4747
rect 6341 4713 6399 4747
rect 6433 4713 6491 4747
rect 6525 4713 6583 4747
rect 6617 4713 6675 4747
rect 6709 4713 6767 4747
rect 6801 4713 6859 4747
rect 6893 4713 6951 4747
rect 6985 4713 7043 4747
rect 7077 4713 7135 4747
rect 7169 4713 7227 4747
rect 7261 4713 7319 4747
rect 7353 4713 7411 4747
rect 7445 4713 7503 4747
rect 7537 4713 7595 4747
rect 7629 4713 7687 4747
rect 7721 4713 7779 4747
rect 7813 4713 7871 4747
rect 7905 4713 7963 4747
rect 7997 4713 8055 4747
rect 8089 4713 8147 4747
rect 8181 4713 8239 4747
rect 8273 4713 8331 4747
rect 8365 4713 8423 4747
rect 8457 4713 8515 4747
rect 8549 4713 8607 4747
rect 8641 4713 8699 4747
rect 8733 4713 8791 4747
rect 8825 4713 8883 4747
rect 8917 4713 8975 4747
rect 9009 4713 9067 4747
rect 9101 4713 9159 4747
rect 9193 4713 9251 4747
rect 9285 4713 9343 4747
rect 9377 4713 9435 4747
rect 9469 4713 9527 4747
rect 9561 4713 9619 4747
rect 9653 4713 9711 4747
rect 9745 4713 9803 4747
rect 9837 4713 9895 4747
rect 9929 4713 9987 4747
rect 10021 4713 10079 4747
rect 10113 4713 10171 4747
rect 10205 4713 10263 4747
rect 10297 4713 10355 4747
rect 10389 4713 10447 4747
rect 10481 4713 10539 4747
rect 10573 4713 10631 4747
rect 10665 4713 10723 4747
rect 10757 4713 10815 4747
rect 10849 4713 10907 4747
rect 10941 4713 10999 4747
rect 11033 4713 11091 4747
rect 11125 4713 11183 4747
rect 11217 4713 11275 4747
rect 11309 4713 11367 4747
rect 11401 4713 11459 4747
rect 11493 4713 11551 4747
rect 11585 4713 11643 4747
rect 11677 4713 11735 4747
rect 11769 4713 11827 4747
rect 11861 4713 11919 4747
rect 11953 4713 12011 4747
rect 12045 4713 12103 4747
rect 12137 4713 12195 4747
rect 12229 4713 12287 4747
rect 12321 4713 12379 4747
rect 12413 4713 12471 4747
rect 12505 4713 12563 4747
rect 12597 4713 12655 4747
rect 12689 4713 12747 4747
rect 12781 4713 12839 4747
rect 12873 4713 12931 4747
rect 12965 4713 12994 4747
rect 594 4024 623 4058
rect 657 4024 715 4058
rect 749 4024 807 4058
rect 841 4024 899 4058
rect 933 4024 991 4058
rect 1025 4024 1083 4058
rect 1117 4024 1175 4058
rect 1209 4024 1267 4058
rect 1301 4024 1359 4058
rect 1393 4024 1451 4058
rect 1485 4024 1543 4058
rect 1577 4024 1635 4058
rect 1669 4024 1727 4058
rect 1761 4024 1819 4058
rect 1853 4024 1911 4058
rect 1945 4024 2003 4058
rect 2037 4024 2095 4058
rect 2129 4024 2187 4058
rect 2221 4024 2279 4058
rect 2313 4024 2371 4058
rect 2405 4024 2463 4058
rect 2497 4024 2555 4058
rect 2589 4024 2647 4058
rect 2681 4024 2739 4058
rect 2773 4024 2831 4058
rect 2865 4024 2923 4058
rect 2957 4024 3015 4058
rect 3049 4024 3107 4058
rect 3141 4024 3199 4058
rect 3233 4024 3291 4058
rect 3325 4024 3383 4058
rect 3417 4024 3475 4058
rect 3509 4024 3567 4058
rect 3601 4024 3659 4058
rect 3693 4024 3751 4058
rect 3785 4024 3843 4058
rect 3877 4024 3935 4058
rect 3969 4024 4027 4058
rect 4061 4024 4119 4058
rect 4153 4024 4211 4058
rect 4245 4024 4303 4058
rect 4337 4024 4395 4058
rect 4429 4024 4487 4058
rect 4521 4024 4579 4058
rect 4613 4024 4671 4058
rect 4705 4024 4763 4058
rect 4797 4024 4855 4058
rect 4889 4024 4947 4058
rect 4981 4024 5039 4058
rect 5073 4024 5131 4058
rect 5165 4024 5223 4058
rect 5257 4024 5315 4058
rect 5349 4024 5407 4058
rect 5441 4024 5499 4058
rect 5533 4024 5591 4058
rect 5625 4024 5683 4058
rect 5717 4024 5775 4058
rect 5809 4024 5867 4058
rect 5901 4024 5959 4058
rect 5993 4024 6051 4058
rect 6085 4024 6143 4058
rect 6177 4024 6235 4058
rect 6269 4024 6327 4058
rect 6361 4024 6419 4058
rect 6453 4024 6511 4058
rect 6545 4024 6603 4058
rect 6637 4024 6695 4058
rect 6729 4024 6787 4058
rect 6821 4024 6879 4058
rect 6913 4024 6971 4058
rect 7005 4024 7063 4058
rect 7097 4024 7155 4058
rect 7189 4024 7247 4058
rect 7281 4024 7339 4058
rect 7373 4024 7431 4058
rect 7465 4024 7523 4058
rect 7557 4024 7615 4058
rect 7649 4024 7707 4058
rect 7741 4024 7799 4058
rect 7833 4024 7891 4058
rect 7925 4024 7983 4058
rect 8017 4024 8075 4058
rect 8109 4024 8167 4058
rect 8201 4024 8259 4058
rect 8293 4024 8351 4058
rect 8385 4024 8443 4058
rect 8477 4024 8535 4058
rect 8569 4024 8627 4058
rect 8661 4024 8719 4058
rect 8753 4024 8811 4058
rect 8845 4024 8903 4058
rect 8937 4024 8995 4058
rect 9029 4024 9087 4058
rect 9121 4024 9179 4058
rect 9213 4024 9271 4058
rect 9305 4024 9363 4058
rect 9397 4024 9435 4058
rect 9469 4024 9527 4058
rect 9561 4024 9619 4058
rect 9653 4024 9711 4058
rect 9745 4024 9803 4058
rect 9837 4024 9895 4058
rect 9929 4024 9987 4058
rect 10021 4024 10079 4058
rect 10113 4024 10171 4058
rect 10205 4024 10263 4058
rect 10297 4024 10355 4058
rect 10389 4024 10447 4058
rect 10481 4024 10539 4058
rect 10573 4024 10631 4058
rect 10665 4024 10723 4058
rect 10757 4024 10815 4058
rect 10849 4024 10907 4058
rect 10941 4024 10999 4058
rect 11033 4024 11091 4058
rect 11125 4024 11183 4058
rect 11217 4024 11275 4058
rect 11309 4024 11367 4058
rect 11401 4024 11459 4058
rect 11493 4024 11551 4058
rect 11585 4024 11643 4058
rect 11677 4024 11735 4058
rect 11769 4024 11827 4058
rect 11861 4024 11919 4058
rect 11953 4024 12011 4058
rect 12045 4024 12103 4058
rect 12137 4024 12195 4058
rect 12229 4024 12287 4058
rect 12321 4024 12379 4058
rect 12413 4024 12471 4058
rect 12505 4024 12563 4058
rect 12597 4024 12655 4058
rect 12689 4024 12747 4058
rect 12781 4024 12839 4058
rect 12873 4024 12931 4058
rect 12965 4024 12994 4058
rect 626 3139 654 3173
rect 688 3139 747 3173
rect 781 3139 839 3173
rect 873 3139 931 3173
rect 965 3139 1023 3173
rect 1057 3139 1115 3173
rect 1149 3139 1207 3173
rect 1241 3139 1299 3173
rect 1333 3139 1391 3173
rect 1425 3139 1454 3173
rect 3167 3151 3197 3185
rect 3231 3151 3289 3185
rect 3323 3151 3381 3185
rect 3415 3151 3473 3185
rect 3507 3151 3565 3185
rect 3599 3151 3657 3185
rect 3691 3151 3749 3185
rect 3783 3151 3841 3185
rect 3875 3151 3933 3185
rect 3967 3151 4025 3185
rect 4059 3151 4117 3185
rect 4151 3151 4209 3185
rect 4243 3151 4301 3185
rect 4335 3151 4393 3185
rect 4427 3151 4485 3185
rect 4519 3151 4577 3185
rect 4611 3151 4669 3185
rect 4703 3151 4761 3185
rect 4795 3151 4853 3185
rect 4887 3151 4945 3185
rect 4979 3151 5037 3185
rect 5071 3151 5129 3185
rect 5163 3151 5221 3185
rect 5255 3151 5313 3185
rect 5347 3151 5405 3185
rect 5439 3151 5497 3185
rect 5531 3151 5589 3185
rect 5623 3151 5681 3185
rect 5715 3151 5773 3185
rect 5807 3151 5865 3185
rect 5899 3151 5957 3185
rect 5991 3151 6049 3185
rect 6083 3151 6141 3185
rect 6175 3151 6233 3185
rect 6267 3151 6325 3185
rect 6359 3151 6417 3185
rect 6451 3151 6509 3185
rect 6543 3151 6601 3185
rect 6635 3151 6693 3185
rect 6727 3151 6785 3185
rect 6819 3151 6877 3185
rect 6911 3151 6969 3185
rect 7003 3151 7061 3185
rect 7095 3151 7153 3185
rect 7187 3151 7245 3185
rect 7279 3151 7337 3185
rect 7371 3151 7429 3185
rect 7463 3151 7521 3185
rect 7555 3151 7613 3185
rect 7647 3151 7705 3185
rect 7739 3151 7797 3185
rect 7831 3151 7889 3185
rect 7923 3151 7981 3185
rect 8015 3151 8073 3185
rect 8107 3151 8165 3185
rect 8199 3151 8257 3185
rect 8291 3151 8349 3185
rect 8383 3151 8441 3185
rect 8475 3151 8533 3185
rect 8567 3151 8625 3185
rect 8659 3151 8717 3185
rect 8751 3151 8809 3185
rect 8843 3151 8901 3185
rect 8935 3151 8993 3185
rect 9027 3151 9085 3185
rect 9119 3151 9177 3185
rect 9211 3151 9269 3185
rect 9303 3151 9361 3185
rect 9395 3151 9453 3185
rect 9487 3151 9545 3185
rect 9579 3151 9637 3185
rect 9671 3151 9729 3185
rect 9763 3151 9821 3185
rect 9855 3151 9894 3185
rect 9947 3151 9986 3185
rect 10039 3151 10078 3185
rect 10131 3151 10170 3185
rect 10223 3151 10262 3185
rect 10315 3151 10354 3185
rect 10407 3151 10446 3185
rect 10499 3151 10538 3185
rect 10591 3151 10630 3185
rect 10683 3151 10722 3185
rect 10775 3151 10814 3185
rect 10867 3151 10906 3185
rect 10959 3151 10998 3185
rect 11051 3151 11090 3185
rect 11143 3151 11182 3185
rect 11235 3151 11274 3185
rect 11327 3151 11366 3185
rect 11419 3151 11458 3185
rect 11511 3151 11550 3185
rect 11603 3151 11642 3185
rect 11695 3151 11734 3185
rect 11787 3151 11826 3185
rect 11879 3151 11918 3185
rect 11971 3151 12010 3185
rect 12044 3151 12102 3185
rect 12136 3151 12194 3185
rect 12228 3151 12286 3185
rect 12320 3151 12378 3185
rect 12412 3151 12470 3185
rect 12504 3151 12562 3185
rect 12596 3151 12654 3185
rect 12688 3151 12746 3185
rect 12780 3151 12838 3185
rect 12872 3151 12930 3185
rect 12964 3151 12992 3185
rect 1033 2278 1062 2312
rect 1096 2278 1154 2312
rect 1188 2278 1246 2312
rect 1280 2278 1338 2312
rect 1372 2278 1430 2312
rect 1464 2278 1522 2312
rect 1556 2278 1614 2312
rect 1648 2278 1706 2312
rect 1740 2278 1798 2312
rect 1832 2278 1890 2312
rect 1924 2278 1982 2312
rect 2016 2278 2074 2312
rect 2108 2278 2166 2312
rect 2200 2278 2258 2312
rect 2292 2278 2350 2312
rect 2384 2278 2442 2312
rect 2476 2278 2534 2312
rect 2568 2278 2626 2312
rect 2660 2278 2718 2312
rect 2752 2278 2810 2312
rect 2844 2278 2902 2312
rect 2936 2278 2994 2312
rect 3028 2278 3086 2312
rect 3120 2278 3178 2312
rect 3212 2278 3270 2312
rect 3304 2278 3362 2312
rect 3396 2278 3454 2312
rect 3488 2278 3546 2312
rect 3580 2278 3638 2312
rect 3672 2278 3730 2312
rect 3764 2278 3822 2312
rect 3856 2278 3914 2312
rect 3948 2278 4006 2312
rect 4040 2278 4098 2312
rect 4132 2278 4190 2312
rect 4224 2278 4282 2312
rect 4316 2278 4374 2312
rect 4408 2278 4466 2312
rect 4500 2278 4558 2312
rect 4592 2278 4650 2312
rect 4684 2278 4742 2312
rect 4776 2278 4834 2312
rect 4868 2278 4926 2312
rect 4960 2278 5018 2312
rect 5052 2278 5110 2312
rect 5144 2278 5202 2312
rect 5236 2278 5294 2312
rect 5328 2278 5386 2312
rect 5420 2278 5478 2312
rect 5512 2278 5570 2312
rect 5604 2278 5662 2312
rect 5696 2278 5754 2312
rect 5788 2278 5846 2312
rect 5880 2278 5938 2312
rect 5972 2278 6030 2312
rect 6064 2278 6122 2312
rect 6156 2278 6214 2312
rect 6248 2278 6306 2312
rect 6340 2278 6398 2312
rect 6432 2278 6490 2312
rect 6524 2278 6582 2312
rect 6616 2278 6674 2312
rect 6708 2278 6766 2312
rect 6800 2278 6858 2312
rect 6892 2278 6950 2312
rect 6984 2278 7042 2312
rect 7076 2278 7134 2312
rect 7168 2278 7226 2312
rect 7260 2278 7318 2312
rect 7352 2278 7410 2312
rect 7444 2278 7502 2312
rect 7536 2278 7594 2312
rect 7628 2278 7686 2312
rect 7720 2278 7778 2312
rect 7812 2278 7870 2312
rect 7904 2278 7962 2312
rect 7996 2278 8054 2312
rect 8088 2278 8146 2312
rect 8180 2278 8238 2312
rect 8272 2278 8330 2312
rect 8364 2278 8422 2312
rect 8456 2278 8514 2312
rect 8548 2278 8606 2312
rect 8640 2278 8698 2312
rect 8732 2278 8790 2312
rect 8824 2278 8882 2312
rect 8916 2278 8974 2312
rect 9008 2278 9066 2312
rect 9100 2278 9158 2312
rect 9192 2278 9250 2312
rect 9284 2278 9342 2312
rect 9376 2278 9434 2312
rect 9468 2278 9526 2312
rect 9560 2278 9618 2312
rect 9652 2278 9710 2312
rect 9744 2278 9802 2312
rect 9836 2278 9894 2312
rect 9928 2278 9986 2312
rect 10020 2278 10078 2312
rect 10112 2278 10170 2312
rect 10204 2278 10262 2312
rect 10296 2278 10354 2312
rect 10388 2278 10446 2312
rect 10480 2278 10538 2312
rect 10572 2278 10630 2312
rect 10664 2278 10722 2312
rect 10756 2278 10814 2312
rect 10848 2278 10906 2312
rect 10940 2278 10998 2312
rect 11032 2278 11090 2312
rect 11124 2278 11182 2312
rect 11216 2278 11274 2312
rect 11308 2278 11366 2312
rect 11400 2278 11458 2312
rect 11492 2278 11550 2312
rect 11584 2278 11642 2312
rect 11676 2278 11734 2312
rect 11768 2278 11826 2312
rect 11860 2278 11918 2312
rect 11952 2278 12010 2312
rect 12044 2278 12102 2312
rect 12136 2278 12194 2312
rect 12228 2278 12286 2312
rect 12320 2278 12378 2312
rect 12412 2278 12470 2312
rect 12504 2278 12562 2312
rect 12596 2278 12654 2312
rect 12688 2278 12746 2312
rect 12780 2278 12838 2312
rect 12872 2278 12930 2312
rect 12964 2278 12993 2312
<< nsubdiff >>
rect 1035 6178 1064 6212
rect 1098 6178 1156 6212
rect 1190 6178 1248 6212
rect 1282 6178 1340 6212
rect 1374 6178 1432 6212
rect 1466 6178 1524 6212
rect 1558 6178 1616 6212
rect 1650 6178 1679 6212
rect 2295 6178 2324 6212
rect 2358 6178 2416 6212
rect 2450 6178 2508 6212
rect 2542 6178 2600 6212
rect 2634 6178 2692 6212
rect 2726 6178 2784 6212
rect 2818 6178 2876 6212
rect 2910 6178 2968 6212
rect 3002 6178 3060 6212
rect 3094 6178 3152 6212
rect 3186 6178 3244 6212
rect 3278 6178 3336 6212
rect 3370 6178 3428 6212
rect 3462 6178 3520 6212
rect 3554 6178 3612 6212
rect 3646 6178 3704 6212
rect 3738 6178 3796 6212
rect 3830 6178 3888 6212
rect 3922 6178 3980 6212
rect 4014 6178 4072 6212
rect 4106 6178 4135 6212
rect 1034 5305 1063 5339
rect 1097 5305 1155 5339
rect 1189 5305 1247 5339
rect 1281 5305 1339 5339
rect 1373 5305 1431 5339
rect 1465 5305 1523 5339
rect 1557 5305 1615 5339
rect 1649 5305 1707 5339
rect 1741 5305 1799 5339
rect 1833 5305 1891 5339
rect 1925 5305 1983 5339
rect 2017 5305 2075 5339
rect 2109 5305 2167 5339
rect 2201 5305 2259 5339
rect 2293 5305 2351 5339
rect 2385 5305 2443 5339
rect 2477 5305 2535 5339
rect 2569 5305 2627 5339
rect 2661 5305 2719 5339
rect 2753 5305 2811 5339
rect 2845 5305 2895 5339
rect 3007 5305 3087 5339
rect 3121 5305 3179 5339
rect 3213 5305 3271 5339
rect 3305 5305 3363 5339
rect 3397 5305 3455 5339
rect 3489 5305 3547 5339
rect 3581 5305 3640 5339
rect 3674 5305 3731 5339
rect 3765 5305 3823 5339
rect 3857 5305 3915 5339
rect 3949 5305 4007 5339
rect 4041 5305 4139 5339
rect 4249 5305 4283 5339
rect 4317 5305 4375 5339
rect 4409 5305 4467 5339
rect 4501 5305 4559 5339
rect 4593 5305 4651 5339
rect 4685 5305 4743 5339
rect 4777 5305 4835 5339
rect 4869 5305 4927 5339
rect 4961 5305 5019 5339
rect 5053 5305 5111 5339
rect 5145 5305 5203 5339
rect 5237 5305 5295 5339
rect 5329 5305 5387 5339
rect 5421 5305 5479 5339
rect 5513 5305 5571 5339
rect 5605 5305 5663 5339
rect 5697 5305 5755 5339
rect 5789 5305 5847 5339
rect 5881 5305 5939 5339
rect 5973 5305 6031 5339
rect 6065 5305 6123 5339
rect 6157 5305 6215 5339
rect 6249 5305 6307 5339
rect 6341 5305 6399 5339
rect 6433 5305 6531 5339
rect 6641 5305 6675 5339
rect 6709 5305 6767 5339
rect 6801 5305 6859 5339
rect 6893 5305 6951 5339
rect 6985 5305 7043 5339
rect 7077 5305 7135 5339
rect 7169 5305 7227 5339
rect 7261 5305 7319 5339
rect 7353 5305 7411 5339
rect 7445 5305 7503 5339
rect 7537 5305 7595 5339
rect 7629 5305 7687 5339
rect 7721 5305 7779 5339
rect 7813 5305 7871 5339
rect 7905 5305 7963 5339
rect 7997 5305 8055 5339
rect 8089 5305 8147 5339
rect 8181 5305 8239 5339
rect 8273 5305 8331 5339
rect 8365 5305 8423 5339
rect 8457 5305 8515 5339
rect 8549 5305 8607 5339
rect 8641 5305 8699 5339
rect 8733 5305 8791 5339
rect 8825 5305 8923 5339
rect 9033 5305 9067 5339
rect 9101 5305 9159 5339
rect 9193 5305 9251 5339
rect 9285 5305 9343 5339
rect 9377 5305 9435 5339
rect 9469 5305 9527 5339
rect 9561 5305 9619 5339
rect 9653 5305 9711 5339
rect 9745 5305 9803 5339
rect 9837 5305 9895 5339
rect 9929 5305 9987 5339
rect 10021 5305 10079 5339
rect 10113 5305 10171 5339
rect 10205 5305 10263 5339
rect 10297 5305 10355 5339
rect 10389 5305 10447 5339
rect 10481 5305 10539 5339
rect 10573 5305 10631 5339
rect 10665 5305 10723 5339
rect 10757 5305 10815 5339
rect 10849 5305 10907 5339
rect 10941 5305 10999 5339
rect 11033 5305 11091 5339
rect 11125 5305 11183 5339
rect 11217 5305 11315 5339
rect 11425 5305 11459 5339
rect 11493 5305 11551 5339
rect 11585 5305 11643 5339
rect 11677 5305 11735 5339
rect 11769 5305 11827 5339
rect 11861 5305 11919 5339
rect 11953 5305 12011 5339
rect 12045 5305 12103 5339
rect 12137 5305 12195 5339
rect 12229 5305 12287 5339
rect 12321 5305 12379 5339
rect 12413 5305 12471 5339
rect 12505 5305 12563 5339
rect 12597 5305 12655 5339
rect 12689 5305 12747 5339
rect 12781 5305 12839 5339
rect 12873 5305 12931 5339
rect 12965 5305 12994 5339
rect 594 4616 623 4650
rect 657 4616 715 4650
rect 749 4616 807 4650
rect 841 4616 899 4650
rect 933 4616 991 4650
rect 1025 4616 1083 4650
rect 1117 4616 1175 4650
rect 1209 4616 1267 4650
rect 1301 4616 1359 4650
rect 1393 4616 1451 4650
rect 1485 4616 1543 4650
rect 1577 4616 1635 4650
rect 1669 4616 1727 4650
rect 1761 4616 1819 4650
rect 1853 4616 1911 4650
rect 1945 4616 2003 4650
rect 2037 4616 2095 4650
rect 2129 4616 2187 4650
rect 2221 4616 2279 4650
rect 2313 4616 2351 4650
rect 2405 4616 2443 4650
rect 2477 4616 2535 4650
rect 2569 4616 2627 4650
rect 2661 4616 2719 4650
rect 2753 4616 2811 4650
rect 2845 4616 2903 4650
rect 2937 4616 2995 4650
rect 3029 4616 3087 4650
rect 3121 4616 3179 4650
rect 3213 4616 3271 4650
rect 3305 4616 3363 4650
rect 3397 4616 3455 4650
rect 3489 4616 3547 4650
rect 3581 4616 3639 4650
rect 3673 4616 3731 4650
rect 3765 4616 3823 4650
rect 3857 4616 3915 4650
rect 3949 4616 4007 4650
rect 4041 4616 4099 4650
rect 4133 4616 4210 4650
rect 4320 4616 4375 4650
rect 4409 4616 4467 4650
rect 4501 4616 4559 4650
rect 4593 4616 4651 4650
rect 4685 4616 4743 4650
rect 4777 4616 4835 4650
rect 4869 4616 4927 4650
rect 4961 4616 5019 4650
rect 5053 4616 5111 4650
rect 5145 4616 5203 4650
rect 5237 4616 5295 4650
rect 5329 4616 5387 4650
rect 5421 4616 5479 4650
rect 5513 4616 5571 4650
rect 5605 4616 5663 4650
rect 5697 4616 5755 4650
rect 5789 4616 5847 4650
rect 5881 4616 5939 4650
rect 5973 4616 6031 4650
rect 6065 4616 6123 4650
rect 6157 4616 6215 4650
rect 6249 4616 6307 4650
rect 6341 4616 6399 4650
rect 6433 4616 6491 4650
rect 6525 4616 6602 4650
rect 6712 4616 6767 4650
rect 6801 4616 6859 4650
rect 6893 4616 6951 4650
rect 6985 4616 7043 4650
rect 7077 4616 7135 4650
rect 7169 4616 7227 4650
rect 7261 4616 7319 4650
rect 7353 4616 7411 4650
rect 7445 4616 7503 4650
rect 7537 4616 7595 4650
rect 7629 4616 7687 4650
rect 7721 4616 7779 4650
rect 7813 4616 7871 4650
rect 7905 4616 7963 4650
rect 7997 4616 8055 4650
rect 8089 4616 8147 4650
rect 8181 4616 8239 4650
rect 8273 4616 8331 4650
rect 8365 4616 8423 4650
rect 8457 4616 8515 4650
rect 8549 4616 8607 4650
rect 8641 4616 8699 4650
rect 8733 4616 8791 4650
rect 8825 4616 8883 4650
rect 8917 4616 8994 4650
rect 9104 4616 9159 4650
rect 9193 4616 9251 4650
rect 9285 4616 9343 4650
rect 9377 4616 9435 4650
rect 9469 4616 9527 4650
rect 9561 4616 9619 4650
rect 9653 4616 9711 4650
rect 9745 4616 9803 4650
rect 9837 4616 9895 4650
rect 9929 4616 9987 4650
rect 10021 4616 10079 4650
rect 10113 4616 10171 4650
rect 10205 4616 10263 4650
rect 10297 4616 10355 4650
rect 10389 4616 10447 4650
rect 10481 4616 10539 4650
rect 10573 4616 10631 4650
rect 10665 4616 10723 4650
rect 10757 4616 10815 4650
rect 10849 4616 10907 4650
rect 10941 4616 10999 4650
rect 11033 4616 11091 4650
rect 11125 4616 11183 4650
rect 11217 4616 11275 4650
rect 11309 4616 11386 4650
rect 11496 4616 11551 4650
rect 11585 4616 11643 4650
rect 11677 4616 11735 4650
rect 11769 4616 11827 4650
rect 11861 4616 11919 4650
rect 11953 4616 12011 4650
rect 12045 4616 12103 4650
rect 12137 4616 12195 4650
rect 12229 4616 12287 4650
rect 12321 4616 12379 4650
rect 12413 4616 12471 4650
rect 12505 4616 12563 4650
rect 12597 4616 12655 4650
rect 12689 4616 12747 4650
rect 12781 4616 12839 4650
rect 12873 4616 12931 4650
rect 12965 4616 12996 4650
rect 626 3752 655 3786
rect 689 3752 747 3786
rect 781 3752 839 3786
rect 873 3752 931 3786
rect 965 3752 1023 3786
rect 1057 3752 1114 3786
rect 1148 3752 1206 3786
rect 1240 3752 1299 3786
rect 1333 3752 1391 3786
rect 1425 3752 1455 3786
rect 626 3751 1455 3752
rect 3168 3743 3197 3777
rect 3231 3743 3289 3777
rect 3323 3743 3381 3777
rect 3415 3743 3473 3777
rect 3507 3743 3565 3777
rect 3599 3743 3657 3777
rect 3691 3743 3749 3777
rect 3783 3743 3841 3777
rect 3875 3743 3933 3777
rect 3967 3743 4025 3777
rect 4059 3743 4117 3777
rect 4151 3743 4209 3777
rect 4243 3743 4301 3777
rect 4335 3743 4393 3777
rect 4427 3743 4485 3777
rect 4519 3743 4577 3777
rect 4611 3743 4669 3777
rect 4703 3743 4761 3777
rect 4795 3743 4853 3777
rect 4887 3743 4945 3777
rect 4979 3743 5018 3777
rect 5052 3743 5110 3777
rect 5144 3743 5202 3777
rect 5236 3743 5294 3777
rect 5328 3743 5386 3777
rect 5420 3743 5478 3777
rect 5512 3743 5570 3777
rect 5604 3743 5662 3777
rect 5696 3743 5754 3777
rect 5788 3743 5846 3777
rect 5880 3743 5938 3777
rect 5972 3743 6030 3777
rect 6064 3743 6122 3777
rect 6156 3743 6214 3777
rect 6248 3743 6306 3777
rect 6340 3743 6398 3777
rect 6432 3743 6490 3777
rect 6524 3743 6582 3777
rect 6616 3743 6674 3777
rect 6708 3743 6766 3777
rect 6800 3743 6858 3777
rect 6892 3743 6950 3777
rect 6984 3743 7042 3777
rect 7076 3743 7134 3777
rect 7168 3743 7226 3777
rect 7260 3743 7318 3777
rect 7352 3743 7410 3777
rect 7444 3743 7502 3777
rect 7536 3743 7594 3777
rect 7628 3743 7686 3777
rect 7720 3743 7778 3777
rect 7812 3743 7870 3777
rect 7904 3743 7962 3777
rect 7996 3743 8054 3777
rect 8088 3743 8146 3777
rect 8180 3743 8238 3777
rect 8272 3743 8330 3777
rect 8364 3743 8422 3777
rect 8456 3743 8514 3777
rect 8548 3743 8606 3777
rect 8640 3743 8698 3777
rect 8732 3743 8790 3777
rect 8824 3743 8882 3777
rect 8916 3743 8974 3777
rect 9008 3743 9066 3777
rect 9100 3743 9158 3777
rect 9192 3743 9250 3777
rect 9284 3743 9342 3777
rect 9376 3743 9434 3777
rect 9468 3743 9526 3777
rect 9560 3743 9618 3777
rect 9652 3743 9710 3777
rect 9744 3743 9802 3777
rect 9836 3743 9894 3777
rect 9928 3743 9986 3777
rect 10020 3743 10078 3777
rect 10112 3743 10170 3777
rect 10204 3743 10262 3777
rect 10296 3743 10354 3777
rect 10388 3743 10446 3777
rect 10480 3743 10538 3777
rect 10572 3743 10630 3777
rect 10664 3743 10722 3777
rect 10756 3743 10814 3777
rect 10848 3743 10906 3777
rect 10940 3743 10998 3777
rect 11032 3743 11090 3777
rect 11124 3743 11182 3777
rect 11216 3743 11274 3777
rect 11308 3743 11366 3777
rect 11400 3743 11458 3777
rect 11492 3743 11550 3777
rect 11584 3743 11642 3777
rect 11676 3743 11734 3777
rect 11768 3743 11826 3777
rect 11860 3743 11918 3777
rect 11952 3743 12010 3777
rect 12044 3743 12102 3777
rect 12136 3743 12194 3777
rect 12228 3743 12286 3777
rect 12320 3743 12378 3777
rect 12412 3743 12470 3777
rect 12504 3743 12562 3777
rect 12596 3743 12654 3777
rect 12688 3743 12746 3777
rect 12780 3743 12838 3777
rect 12872 3743 12930 3777
rect 12964 3743 12993 3777
rect 1033 2870 1062 2904
rect 1096 2870 1154 2904
rect 1188 2870 1246 2904
rect 1280 2870 1338 2904
rect 1372 2870 1430 2904
rect 1464 2870 1522 2904
rect 1556 2870 1614 2904
rect 1648 2870 1706 2904
rect 1740 2870 1798 2904
rect 1832 2870 1890 2904
rect 1924 2870 1982 2904
rect 2016 2870 2074 2904
rect 2108 2870 2166 2904
rect 2200 2870 2258 2904
rect 2292 2870 2350 2904
rect 2384 2870 2442 2904
rect 2476 2870 2534 2904
rect 2568 2870 2626 2904
rect 2660 2870 2718 2904
rect 2752 2870 2810 2904
rect 2844 2870 2902 2904
rect 2936 2870 2994 2904
rect 3028 2870 3086 2904
rect 3120 2870 3178 2904
rect 3212 2870 3270 2904
rect 3304 2870 3362 2904
rect 3396 2870 3454 2904
rect 3488 2870 3546 2904
rect 3580 2870 3638 2904
rect 3672 2870 3730 2904
rect 3764 2870 3822 2904
rect 3856 2870 3914 2904
rect 3948 2870 4006 2904
rect 4040 2870 4098 2904
rect 4132 2870 4190 2904
rect 4224 2870 4282 2904
rect 4316 2870 4374 2904
rect 4408 2870 4466 2904
rect 4500 2870 4558 2904
rect 4592 2870 4650 2904
rect 4684 2870 4742 2904
rect 4776 2870 4834 2904
rect 4868 2870 4926 2904
rect 4960 2870 5018 2904
rect 5052 2870 5110 2904
rect 5144 2870 5202 2904
rect 5236 2870 5294 2904
rect 5328 2870 5386 2904
rect 5420 2870 5478 2904
rect 5512 2870 5570 2904
rect 5604 2870 5662 2904
rect 5696 2870 5754 2904
rect 5788 2870 5846 2904
rect 5880 2870 5938 2904
rect 5972 2870 6030 2904
rect 6064 2870 6122 2904
rect 6156 2870 6214 2904
rect 6248 2870 6306 2904
rect 6340 2870 6398 2904
rect 6432 2870 6490 2904
rect 6524 2870 6582 2904
rect 6616 2870 6674 2904
rect 6708 2870 6766 2904
rect 6800 2870 6858 2904
rect 6892 2870 6950 2904
rect 6984 2870 7042 2904
rect 7076 2870 7134 2904
rect 7168 2870 7226 2904
rect 7260 2870 7318 2904
rect 7352 2870 7410 2904
rect 7444 2870 7502 2904
rect 7536 2870 7594 2904
rect 7628 2870 7686 2904
rect 7720 2870 7778 2904
rect 7812 2870 7870 2904
rect 7904 2870 7962 2904
rect 7996 2870 8054 2904
rect 8088 2870 8146 2904
rect 8180 2870 8238 2904
rect 8272 2870 8330 2904
rect 8364 2870 8422 2904
rect 8456 2870 8514 2904
rect 8548 2870 8606 2904
rect 8640 2870 8698 2904
rect 8732 2870 8790 2904
rect 8824 2870 8882 2904
rect 8916 2870 8974 2904
rect 9008 2870 9066 2904
rect 9100 2870 9158 2904
rect 9192 2870 9250 2904
rect 9284 2870 9342 2904
rect 9376 2870 9434 2904
rect 9468 2870 9526 2904
rect 9560 2870 9618 2904
rect 9652 2870 9710 2904
rect 9744 2870 9802 2904
rect 9836 2870 9894 2904
rect 9928 2870 9986 2904
rect 10020 2870 10078 2904
rect 10112 2870 10170 2904
rect 10204 2870 10262 2904
rect 10296 2870 10354 2904
rect 10388 2870 10446 2904
rect 10480 2870 10538 2904
rect 10572 2870 10630 2904
rect 10664 2870 10722 2904
rect 10756 2870 10814 2904
rect 10848 2870 10906 2904
rect 10940 2870 10998 2904
rect 11032 2870 11090 2904
rect 11124 2870 11182 2904
rect 11216 2870 11274 2904
rect 11308 2870 11366 2904
rect 11400 2870 11458 2904
rect 11492 2870 11550 2904
rect 11584 2870 11642 2904
rect 11676 2870 11734 2904
rect 11768 2870 11826 2904
rect 11860 2870 11918 2904
rect 11952 2870 12010 2904
rect 12044 2870 12102 2904
rect 12136 2870 12194 2904
rect 12228 2870 12286 2904
rect 12320 2870 12378 2904
rect 12412 2870 12470 2904
rect 12504 2870 12562 2904
rect 12596 2870 12654 2904
rect 12688 2870 12746 2904
rect 12780 2870 12838 2904
rect 12872 2870 12930 2904
rect 12964 2870 12993 2904
<< psubdiffcont >>
rect 1064 5586 1098 5620
rect 1156 5586 1190 5620
rect 1248 5586 1282 5620
rect 1340 5586 1374 5620
rect 1432 5586 1466 5620
rect 1524 5586 1558 5620
rect 1616 5586 1650 5620
rect 1708 5586 1742 5620
rect 1800 5586 1834 5620
rect 1892 5586 1926 5620
rect 1984 5586 2018 5620
rect 2076 5586 2110 5620
rect 2168 5586 2202 5620
rect 2260 5586 2294 5620
rect 2352 5586 2386 5620
rect 2444 5586 2478 5620
rect 2536 5586 2570 5620
rect 2628 5586 2662 5620
rect 2720 5586 2754 5620
rect 2812 5586 2846 5620
rect 2904 5586 2938 5620
rect 2996 5586 3030 5620
rect 3088 5586 3122 5620
rect 3180 5586 3214 5620
rect 3272 5586 3306 5620
rect 3364 5586 3398 5620
rect 3456 5586 3490 5620
rect 3548 5586 3582 5620
rect 3640 5586 3674 5620
rect 3732 5586 3766 5620
rect 3824 5586 3858 5620
rect 3916 5586 3950 5620
rect 4008 5586 4042 5620
rect 1063 4713 1097 4747
rect 1155 4713 1189 4747
rect 1247 4713 1281 4747
rect 1339 4713 1373 4747
rect 1431 4713 1465 4747
rect 1523 4713 1557 4747
rect 1615 4713 1649 4747
rect 1707 4713 1741 4747
rect 1799 4713 1833 4747
rect 1891 4713 1925 4747
rect 1983 4713 2017 4747
rect 2075 4713 2109 4747
rect 2167 4713 2201 4747
rect 2259 4713 2293 4747
rect 2351 4713 2385 4747
rect 2443 4713 2477 4747
rect 2535 4713 2569 4747
rect 2627 4713 2661 4747
rect 2719 4713 2753 4747
rect 2811 4713 2845 4747
rect 2903 4713 2937 4747
rect 2995 4713 3029 4747
rect 3087 4713 3121 4747
rect 3179 4713 3213 4747
rect 3271 4713 3305 4747
rect 3363 4713 3397 4747
rect 3455 4713 3489 4747
rect 3547 4713 3581 4747
rect 3639 4713 3673 4747
rect 3731 4713 3765 4747
rect 3823 4713 3857 4747
rect 3915 4713 3949 4747
rect 4007 4713 4041 4747
rect 4099 4713 4133 4747
rect 4191 4713 4225 4747
rect 4283 4713 4317 4747
rect 4375 4713 4409 4747
rect 4467 4713 4501 4747
rect 4559 4713 4593 4747
rect 4651 4713 4685 4747
rect 4743 4713 4777 4747
rect 4835 4713 4869 4747
rect 4927 4713 4961 4747
rect 5019 4713 5053 4747
rect 5111 4713 5145 4747
rect 5203 4713 5237 4747
rect 5295 4713 5329 4747
rect 5387 4713 5421 4747
rect 5479 4713 5513 4747
rect 5571 4713 5605 4747
rect 5663 4713 5697 4747
rect 5755 4713 5789 4747
rect 5847 4713 5881 4747
rect 5939 4713 5973 4747
rect 6031 4713 6065 4747
rect 6123 4713 6157 4747
rect 6215 4713 6249 4747
rect 6307 4713 6341 4747
rect 6399 4713 6433 4747
rect 6491 4713 6525 4747
rect 6583 4713 6617 4747
rect 6675 4713 6709 4747
rect 6767 4713 6801 4747
rect 6859 4713 6893 4747
rect 6951 4713 6985 4747
rect 7043 4713 7077 4747
rect 7135 4713 7169 4747
rect 7227 4713 7261 4747
rect 7319 4713 7353 4747
rect 7411 4713 7445 4747
rect 7503 4713 7537 4747
rect 7595 4713 7629 4747
rect 7687 4713 7721 4747
rect 7779 4713 7813 4747
rect 7871 4713 7905 4747
rect 7963 4713 7997 4747
rect 8055 4713 8089 4747
rect 8147 4713 8181 4747
rect 8239 4713 8273 4747
rect 8331 4713 8365 4747
rect 8423 4713 8457 4747
rect 8515 4713 8549 4747
rect 8607 4713 8641 4747
rect 8699 4713 8733 4747
rect 8791 4713 8825 4747
rect 8883 4713 8917 4747
rect 8975 4713 9009 4747
rect 9067 4713 9101 4747
rect 9159 4713 9193 4747
rect 9251 4713 9285 4747
rect 9343 4713 9377 4747
rect 9435 4713 9469 4747
rect 9527 4713 9561 4747
rect 9619 4713 9653 4747
rect 9711 4713 9745 4747
rect 9803 4713 9837 4747
rect 9895 4713 9929 4747
rect 9987 4713 10021 4747
rect 10079 4713 10113 4747
rect 10171 4713 10205 4747
rect 10263 4713 10297 4747
rect 10355 4713 10389 4747
rect 10447 4713 10481 4747
rect 10539 4713 10573 4747
rect 10631 4713 10665 4747
rect 10723 4713 10757 4747
rect 10815 4713 10849 4747
rect 10907 4713 10941 4747
rect 10999 4713 11033 4747
rect 11091 4713 11125 4747
rect 11183 4713 11217 4747
rect 11275 4713 11309 4747
rect 11367 4713 11401 4747
rect 11459 4713 11493 4747
rect 11551 4713 11585 4747
rect 11643 4713 11677 4747
rect 11735 4713 11769 4747
rect 11827 4713 11861 4747
rect 11919 4713 11953 4747
rect 12011 4713 12045 4747
rect 12103 4713 12137 4747
rect 12195 4713 12229 4747
rect 12287 4713 12321 4747
rect 12379 4713 12413 4747
rect 12471 4713 12505 4747
rect 12563 4713 12597 4747
rect 12655 4713 12689 4747
rect 12747 4713 12781 4747
rect 12839 4713 12873 4747
rect 12931 4713 12965 4747
rect 623 4024 657 4058
rect 715 4024 749 4058
rect 807 4024 841 4058
rect 899 4024 933 4058
rect 991 4024 1025 4058
rect 1083 4024 1117 4058
rect 1175 4024 1209 4058
rect 1267 4024 1301 4058
rect 1359 4024 1393 4058
rect 1451 4024 1485 4058
rect 1543 4024 1577 4058
rect 1635 4024 1669 4058
rect 1727 4024 1761 4058
rect 1819 4024 1853 4058
rect 1911 4024 1945 4058
rect 2003 4024 2037 4058
rect 2095 4024 2129 4058
rect 2187 4024 2221 4058
rect 2279 4024 2313 4058
rect 2371 4024 2405 4058
rect 2463 4024 2497 4058
rect 2555 4024 2589 4058
rect 2647 4024 2681 4058
rect 2739 4024 2773 4058
rect 2831 4024 2865 4058
rect 2923 4024 2957 4058
rect 3015 4024 3049 4058
rect 3107 4024 3141 4058
rect 3199 4024 3233 4058
rect 3291 4024 3325 4058
rect 3383 4024 3417 4058
rect 3475 4024 3509 4058
rect 3567 4024 3601 4058
rect 3659 4024 3693 4058
rect 3751 4024 3785 4058
rect 3843 4024 3877 4058
rect 3935 4024 3969 4058
rect 4027 4024 4061 4058
rect 4119 4024 4153 4058
rect 4211 4024 4245 4058
rect 4303 4024 4337 4058
rect 4395 4024 4429 4058
rect 4487 4024 4521 4058
rect 4579 4024 4613 4058
rect 4671 4024 4705 4058
rect 4763 4024 4797 4058
rect 4855 4024 4889 4058
rect 4947 4024 4981 4058
rect 5039 4024 5073 4058
rect 5131 4024 5165 4058
rect 5223 4024 5257 4058
rect 5315 4024 5349 4058
rect 5407 4024 5441 4058
rect 5499 4024 5533 4058
rect 5591 4024 5625 4058
rect 5683 4024 5717 4058
rect 5775 4024 5809 4058
rect 5867 4024 5901 4058
rect 5959 4024 5993 4058
rect 6051 4024 6085 4058
rect 6143 4024 6177 4058
rect 6235 4024 6269 4058
rect 6327 4024 6361 4058
rect 6419 4024 6453 4058
rect 6511 4024 6545 4058
rect 6603 4024 6637 4058
rect 6695 4024 6729 4058
rect 6787 4024 6821 4058
rect 6879 4024 6913 4058
rect 6971 4024 7005 4058
rect 7063 4024 7097 4058
rect 7155 4024 7189 4058
rect 7247 4024 7281 4058
rect 7339 4024 7373 4058
rect 7431 4024 7465 4058
rect 7523 4024 7557 4058
rect 7615 4024 7649 4058
rect 7707 4024 7741 4058
rect 7799 4024 7833 4058
rect 7891 4024 7925 4058
rect 7983 4024 8017 4058
rect 8075 4024 8109 4058
rect 8167 4024 8201 4058
rect 8259 4024 8293 4058
rect 8351 4024 8385 4058
rect 8443 4024 8477 4058
rect 8535 4024 8569 4058
rect 8627 4024 8661 4058
rect 8719 4024 8753 4058
rect 8811 4024 8845 4058
rect 8903 4024 8937 4058
rect 8995 4024 9029 4058
rect 9087 4024 9121 4058
rect 9179 4024 9213 4058
rect 9271 4024 9305 4058
rect 9363 4024 9397 4058
rect 9435 4024 9469 4058
rect 9527 4024 9561 4058
rect 9619 4024 9653 4058
rect 9711 4024 9745 4058
rect 9803 4024 9837 4058
rect 9895 4024 9929 4058
rect 9987 4024 10021 4058
rect 10079 4024 10113 4058
rect 10171 4024 10205 4058
rect 10263 4024 10297 4058
rect 10355 4024 10389 4058
rect 10447 4024 10481 4058
rect 10539 4024 10573 4058
rect 10631 4024 10665 4058
rect 10723 4024 10757 4058
rect 10815 4024 10849 4058
rect 10907 4024 10941 4058
rect 10999 4024 11033 4058
rect 11091 4024 11125 4058
rect 11183 4024 11217 4058
rect 11275 4024 11309 4058
rect 11367 4024 11401 4058
rect 11459 4024 11493 4058
rect 11551 4024 11585 4058
rect 11643 4024 11677 4058
rect 11735 4024 11769 4058
rect 11827 4024 11861 4058
rect 11919 4024 11953 4058
rect 12011 4024 12045 4058
rect 12103 4024 12137 4058
rect 12195 4024 12229 4058
rect 12287 4024 12321 4058
rect 12379 4024 12413 4058
rect 12471 4024 12505 4058
rect 12563 4024 12597 4058
rect 12655 4024 12689 4058
rect 12747 4024 12781 4058
rect 12839 4024 12873 4058
rect 12931 4024 12965 4058
rect 654 3139 688 3173
rect 747 3139 781 3173
rect 839 3139 873 3173
rect 931 3139 965 3173
rect 1023 3139 1057 3173
rect 1115 3139 1149 3173
rect 1207 3139 1241 3173
rect 1299 3139 1333 3173
rect 1391 3139 1425 3173
rect 3197 3151 3231 3185
rect 3289 3151 3323 3185
rect 3381 3151 3415 3185
rect 3473 3151 3507 3185
rect 3565 3151 3599 3185
rect 3657 3151 3691 3185
rect 3749 3151 3783 3185
rect 3841 3151 3875 3185
rect 3933 3151 3967 3185
rect 4025 3151 4059 3185
rect 4117 3151 4151 3185
rect 4209 3151 4243 3185
rect 4301 3151 4335 3185
rect 4393 3151 4427 3185
rect 4485 3151 4519 3185
rect 4577 3151 4611 3185
rect 4669 3151 4703 3185
rect 4761 3151 4795 3185
rect 4853 3151 4887 3185
rect 4945 3151 4979 3185
rect 5037 3151 5071 3185
rect 5129 3151 5163 3185
rect 5221 3151 5255 3185
rect 5313 3151 5347 3185
rect 5405 3151 5439 3185
rect 5497 3151 5531 3185
rect 5589 3151 5623 3185
rect 5681 3151 5715 3185
rect 5773 3151 5807 3185
rect 5865 3151 5899 3185
rect 5957 3151 5991 3185
rect 6049 3151 6083 3185
rect 6141 3151 6175 3185
rect 6233 3151 6267 3185
rect 6325 3151 6359 3185
rect 6417 3151 6451 3185
rect 6509 3151 6543 3185
rect 6601 3151 6635 3185
rect 6693 3151 6727 3185
rect 6785 3151 6819 3185
rect 6877 3151 6911 3185
rect 6969 3151 7003 3185
rect 7061 3151 7095 3185
rect 7153 3151 7187 3185
rect 7245 3151 7279 3185
rect 7337 3151 7371 3185
rect 7429 3151 7463 3185
rect 7521 3151 7555 3185
rect 7613 3151 7647 3185
rect 7705 3151 7739 3185
rect 7797 3151 7831 3185
rect 7889 3151 7923 3185
rect 7981 3151 8015 3185
rect 8073 3151 8107 3185
rect 8165 3151 8199 3185
rect 8257 3151 8291 3185
rect 8349 3151 8383 3185
rect 8441 3151 8475 3185
rect 8533 3151 8567 3185
rect 8625 3151 8659 3185
rect 8717 3151 8751 3185
rect 8809 3151 8843 3185
rect 8901 3151 8935 3185
rect 8993 3151 9027 3185
rect 9085 3151 9119 3185
rect 9177 3151 9211 3185
rect 9269 3151 9303 3185
rect 9361 3151 9395 3185
rect 9453 3151 9487 3185
rect 9545 3151 9579 3185
rect 9637 3151 9671 3185
rect 9729 3151 9763 3185
rect 9821 3151 9855 3185
rect 9894 3151 9947 3185
rect 9986 3151 10039 3185
rect 10078 3151 10131 3185
rect 10170 3151 10223 3185
rect 10262 3151 10315 3185
rect 10354 3151 10407 3185
rect 10446 3151 10499 3185
rect 10538 3151 10591 3185
rect 10630 3151 10683 3185
rect 10722 3151 10775 3185
rect 10814 3151 10867 3185
rect 10906 3151 10959 3185
rect 10998 3151 11051 3185
rect 11090 3151 11143 3185
rect 11182 3151 11235 3185
rect 11274 3151 11327 3185
rect 11366 3151 11419 3185
rect 11458 3151 11511 3185
rect 11550 3151 11603 3185
rect 11642 3151 11695 3185
rect 11734 3151 11787 3185
rect 11826 3151 11879 3185
rect 11918 3151 11971 3185
rect 12010 3151 12044 3185
rect 12102 3151 12136 3185
rect 12194 3151 12228 3185
rect 12286 3151 12320 3185
rect 12378 3151 12412 3185
rect 12470 3151 12504 3185
rect 12562 3151 12596 3185
rect 12654 3151 12688 3185
rect 12746 3151 12780 3185
rect 12838 3151 12872 3185
rect 12930 3151 12964 3185
rect 1062 2278 1096 2312
rect 1154 2278 1188 2312
rect 1246 2278 1280 2312
rect 1338 2278 1372 2312
rect 1430 2278 1464 2312
rect 1522 2278 1556 2312
rect 1614 2278 1648 2312
rect 1706 2278 1740 2312
rect 1798 2278 1832 2312
rect 1890 2278 1924 2312
rect 1982 2278 2016 2312
rect 2074 2278 2108 2312
rect 2166 2278 2200 2312
rect 2258 2278 2292 2312
rect 2350 2278 2384 2312
rect 2442 2278 2476 2312
rect 2534 2278 2568 2312
rect 2626 2278 2660 2312
rect 2718 2278 2752 2312
rect 2810 2278 2844 2312
rect 2902 2278 2936 2312
rect 2994 2278 3028 2312
rect 3086 2278 3120 2312
rect 3178 2278 3212 2312
rect 3270 2278 3304 2312
rect 3362 2278 3396 2312
rect 3454 2278 3488 2312
rect 3546 2278 3580 2312
rect 3638 2278 3672 2312
rect 3730 2278 3764 2312
rect 3822 2278 3856 2312
rect 3914 2278 3948 2312
rect 4006 2278 4040 2312
rect 4098 2278 4132 2312
rect 4190 2278 4224 2312
rect 4282 2278 4316 2312
rect 4374 2278 4408 2312
rect 4466 2278 4500 2312
rect 4558 2278 4592 2312
rect 4650 2278 4684 2312
rect 4742 2278 4776 2312
rect 4834 2278 4868 2312
rect 4926 2278 4960 2312
rect 5018 2278 5052 2312
rect 5110 2278 5144 2312
rect 5202 2278 5236 2312
rect 5294 2278 5328 2312
rect 5386 2278 5420 2312
rect 5478 2278 5512 2312
rect 5570 2278 5604 2312
rect 5662 2278 5696 2312
rect 5754 2278 5788 2312
rect 5846 2278 5880 2312
rect 5938 2278 5972 2312
rect 6030 2278 6064 2312
rect 6122 2278 6156 2312
rect 6214 2278 6248 2312
rect 6306 2278 6340 2312
rect 6398 2278 6432 2312
rect 6490 2278 6524 2312
rect 6582 2278 6616 2312
rect 6674 2278 6708 2312
rect 6766 2278 6800 2312
rect 6858 2278 6892 2312
rect 6950 2278 6984 2312
rect 7042 2278 7076 2312
rect 7134 2278 7168 2312
rect 7226 2278 7260 2312
rect 7318 2278 7352 2312
rect 7410 2278 7444 2312
rect 7502 2278 7536 2312
rect 7594 2278 7628 2312
rect 7686 2278 7720 2312
rect 7778 2278 7812 2312
rect 7870 2278 7904 2312
rect 7962 2278 7996 2312
rect 8054 2278 8088 2312
rect 8146 2278 8180 2312
rect 8238 2278 8272 2312
rect 8330 2278 8364 2312
rect 8422 2278 8456 2312
rect 8514 2278 8548 2312
rect 8606 2278 8640 2312
rect 8698 2278 8732 2312
rect 8790 2278 8824 2312
rect 8882 2278 8916 2312
rect 8974 2278 9008 2312
rect 9066 2278 9100 2312
rect 9158 2278 9192 2312
rect 9250 2278 9284 2312
rect 9342 2278 9376 2312
rect 9434 2278 9468 2312
rect 9526 2278 9560 2312
rect 9618 2278 9652 2312
rect 9710 2278 9744 2312
rect 9802 2278 9836 2312
rect 9894 2278 9928 2312
rect 9986 2278 10020 2312
rect 10078 2278 10112 2312
rect 10170 2278 10204 2312
rect 10262 2278 10296 2312
rect 10354 2278 10388 2312
rect 10446 2278 10480 2312
rect 10538 2278 10572 2312
rect 10630 2278 10664 2312
rect 10722 2278 10756 2312
rect 10814 2278 10848 2312
rect 10906 2278 10940 2312
rect 10998 2278 11032 2312
rect 11090 2278 11124 2312
rect 11182 2278 11216 2312
rect 11274 2278 11308 2312
rect 11366 2278 11400 2312
rect 11458 2278 11492 2312
rect 11550 2278 11584 2312
rect 11642 2278 11676 2312
rect 11734 2278 11768 2312
rect 11826 2278 11860 2312
rect 11918 2278 11952 2312
rect 12010 2278 12044 2312
rect 12102 2278 12136 2312
rect 12194 2278 12228 2312
rect 12286 2278 12320 2312
rect 12378 2278 12412 2312
rect 12470 2278 12504 2312
rect 12562 2278 12596 2312
rect 12654 2278 12688 2312
rect 12746 2278 12780 2312
rect 12838 2278 12872 2312
rect 12930 2278 12964 2312
<< nsubdiffcont >>
rect 1064 6178 1098 6212
rect 1156 6178 1190 6212
rect 1248 6178 1282 6212
rect 1340 6178 1374 6212
rect 1432 6178 1466 6212
rect 1524 6178 1558 6212
rect 1616 6178 1650 6212
rect 2324 6178 2358 6212
rect 2416 6178 2450 6212
rect 2508 6178 2542 6212
rect 2600 6178 2634 6212
rect 2692 6178 2726 6212
rect 2784 6178 2818 6212
rect 2876 6178 2910 6212
rect 2968 6178 3002 6212
rect 3060 6178 3094 6212
rect 3152 6178 3186 6212
rect 3244 6178 3278 6212
rect 3336 6178 3370 6212
rect 3428 6178 3462 6212
rect 3520 6178 3554 6212
rect 3612 6178 3646 6212
rect 3704 6178 3738 6212
rect 3796 6178 3830 6212
rect 3888 6178 3922 6212
rect 3980 6178 4014 6212
rect 4072 6178 4106 6212
rect 1063 5305 1097 5339
rect 1155 5305 1189 5339
rect 1247 5305 1281 5339
rect 1339 5305 1373 5339
rect 1431 5305 1465 5339
rect 1523 5305 1557 5339
rect 1615 5305 1649 5339
rect 1707 5305 1741 5339
rect 1799 5305 1833 5339
rect 1891 5305 1925 5339
rect 1983 5305 2017 5339
rect 2075 5305 2109 5339
rect 2167 5305 2201 5339
rect 2259 5305 2293 5339
rect 2351 5305 2385 5339
rect 2443 5305 2477 5339
rect 2535 5305 2569 5339
rect 2627 5305 2661 5339
rect 2719 5305 2753 5339
rect 2811 5305 2845 5339
rect 3087 5305 3121 5339
rect 3179 5305 3213 5339
rect 3271 5305 3305 5339
rect 3363 5305 3397 5339
rect 3455 5305 3489 5339
rect 3547 5305 3581 5339
rect 3640 5305 3674 5339
rect 3731 5305 3765 5339
rect 3823 5305 3857 5339
rect 3915 5305 3949 5339
rect 4007 5305 4041 5339
rect 4283 5305 4317 5339
rect 4375 5305 4409 5339
rect 4467 5305 4501 5339
rect 4559 5305 4593 5339
rect 4651 5305 4685 5339
rect 4743 5305 4777 5339
rect 4835 5305 4869 5339
rect 4927 5305 4961 5339
rect 5019 5305 5053 5339
rect 5111 5305 5145 5339
rect 5203 5305 5237 5339
rect 5295 5305 5329 5339
rect 5387 5305 5421 5339
rect 5479 5305 5513 5339
rect 5571 5305 5605 5339
rect 5663 5305 5697 5339
rect 5755 5305 5789 5339
rect 5847 5305 5881 5339
rect 5939 5305 5973 5339
rect 6031 5305 6065 5339
rect 6123 5305 6157 5339
rect 6215 5305 6249 5339
rect 6307 5305 6341 5339
rect 6399 5305 6433 5339
rect 6675 5305 6709 5339
rect 6767 5305 6801 5339
rect 6859 5305 6893 5339
rect 6951 5305 6985 5339
rect 7043 5305 7077 5339
rect 7135 5305 7169 5339
rect 7227 5305 7261 5339
rect 7319 5305 7353 5339
rect 7411 5305 7445 5339
rect 7503 5305 7537 5339
rect 7595 5305 7629 5339
rect 7687 5305 7721 5339
rect 7779 5305 7813 5339
rect 7871 5305 7905 5339
rect 7963 5305 7997 5339
rect 8055 5305 8089 5339
rect 8147 5305 8181 5339
rect 8239 5305 8273 5339
rect 8331 5305 8365 5339
rect 8423 5305 8457 5339
rect 8515 5305 8549 5339
rect 8607 5305 8641 5339
rect 8699 5305 8733 5339
rect 8791 5305 8825 5339
rect 9067 5305 9101 5339
rect 9159 5305 9193 5339
rect 9251 5305 9285 5339
rect 9343 5305 9377 5339
rect 9435 5305 9469 5339
rect 9527 5305 9561 5339
rect 9619 5305 9653 5339
rect 9711 5305 9745 5339
rect 9803 5305 9837 5339
rect 9895 5305 9929 5339
rect 9987 5305 10021 5339
rect 10079 5305 10113 5339
rect 10171 5305 10205 5339
rect 10263 5305 10297 5339
rect 10355 5305 10389 5339
rect 10447 5305 10481 5339
rect 10539 5305 10573 5339
rect 10631 5305 10665 5339
rect 10723 5305 10757 5339
rect 10815 5305 10849 5339
rect 10907 5305 10941 5339
rect 10999 5305 11033 5339
rect 11091 5305 11125 5339
rect 11183 5305 11217 5339
rect 11459 5305 11493 5339
rect 11551 5305 11585 5339
rect 11643 5305 11677 5339
rect 11735 5305 11769 5339
rect 11827 5305 11861 5339
rect 11919 5305 11953 5339
rect 12011 5305 12045 5339
rect 12103 5305 12137 5339
rect 12195 5305 12229 5339
rect 12287 5305 12321 5339
rect 12379 5305 12413 5339
rect 12471 5305 12505 5339
rect 12563 5305 12597 5339
rect 12655 5305 12689 5339
rect 12747 5305 12781 5339
rect 12839 5305 12873 5339
rect 12931 5305 12965 5339
rect 623 4616 657 4650
rect 715 4616 749 4650
rect 807 4616 841 4650
rect 899 4616 933 4650
rect 991 4616 1025 4650
rect 1083 4616 1117 4650
rect 1175 4616 1209 4650
rect 1267 4616 1301 4650
rect 1359 4616 1393 4650
rect 1451 4616 1485 4650
rect 1543 4616 1577 4650
rect 1635 4616 1669 4650
rect 1727 4616 1761 4650
rect 1819 4616 1853 4650
rect 1911 4616 1945 4650
rect 2003 4616 2037 4650
rect 2095 4616 2129 4650
rect 2187 4616 2221 4650
rect 2279 4616 2313 4650
rect 2351 4616 2405 4650
rect 2443 4616 2477 4650
rect 2535 4616 2569 4650
rect 2627 4616 2661 4650
rect 2719 4616 2753 4650
rect 2811 4616 2845 4650
rect 2903 4616 2937 4650
rect 2995 4616 3029 4650
rect 3087 4616 3121 4650
rect 3179 4616 3213 4650
rect 3271 4616 3305 4650
rect 3363 4616 3397 4650
rect 3455 4616 3489 4650
rect 3547 4616 3581 4650
rect 3639 4616 3673 4650
rect 3731 4616 3765 4650
rect 3823 4616 3857 4650
rect 3915 4616 3949 4650
rect 4007 4616 4041 4650
rect 4099 4616 4133 4650
rect 4375 4616 4409 4650
rect 4467 4616 4501 4650
rect 4559 4616 4593 4650
rect 4651 4616 4685 4650
rect 4743 4616 4777 4650
rect 4835 4616 4869 4650
rect 4927 4616 4961 4650
rect 5019 4616 5053 4650
rect 5111 4616 5145 4650
rect 5203 4616 5237 4650
rect 5295 4616 5329 4650
rect 5387 4616 5421 4650
rect 5479 4616 5513 4650
rect 5571 4616 5605 4650
rect 5663 4616 5697 4650
rect 5755 4616 5789 4650
rect 5847 4616 5881 4650
rect 5939 4616 5973 4650
rect 6031 4616 6065 4650
rect 6123 4616 6157 4650
rect 6215 4616 6249 4650
rect 6307 4616 6341 4650
rect 6399 4616 6433 4650
rect 6491 4616 6525 4650
rect 6767 4616 6801 4650
rect 6859 4616 6893 4650
rect 6951 4616 6985 4650
rect 7043 4616 7077 4650
rect 7135 4616 7169 4650
rect 7227 4616 7261 4650
rect 7319 4616 7353 4650
rect 7411 4616 7445 4650
rect 7503 4616 7537 4650
rect 7595 4616 7629 4650
rect 7687 4616 7721 4650
rect 7779 4616 7813 4650
rect 7871 4616 7905 4650
rect 7963 4616 7997 4650
rect 8055 4616 8089 4650
rect 8147 4616 8181 4650
rect 8239 4616 8273 4650
rect 8331 4616 8365 4650
rect 8423 4616 8457 4650
rect 8515 4616 8549 4650
rect 8607 4616 8641 4650
rect 8699 4616 8733 4650
rect 8791 4616 8825 4650
rect 8883 4616 8917 4650
rect 9159 4616 9193 4650
rect 9251 4616 9285 4650
rect 9343 4616 9377 4650
rect 9435 4616 9469 4650
rect 9527 4616 9561 4650
rect 9619 4616 9653 4650
rect 9711 4616 9745 4650
rect 9803 4616 9837 4650
rect 9895 4616 9929 4650
rect 9987 4616 10021 4650
rect 10079 4616 10113 4650
rect 10171 4616 10205 4650
rect 10263 4616 10297 4650
rect 10355 4616 10389 4650
rect 10447 4616 10481 4650
rect 10539 4616 10573 4650
rect 10631 4616 10665 4650
rect 10723 4616 10757 4650
rect 10815 4616 10849 4650
rect 10907 4616 10941 4650
rect 10999 4616 11033 4650
rect 11091 4616 11125 4650
rect 11183 4616 11217 4650
rect 11275 4616 11309 4650
rect 11551 4616 11585 4650
rect 11643 4616 11677 4650
rect 11735 4616 11769 4650
rect 11827 4616 11861 4650
rect 11919 4616 11953 4650
rect 12011 4616 12045 4650
rect 12103 4616 12137 4650
rect 12195 4616 12229 4650
rect 12287 4616 12321 4650
rect 12379 4616 12413 4650
rect 12471 4616 12505 4650
rect 12563 4616 12597 4650
rect 12655 4616 12689 4650
rect 12747 4616 12781 4650
rect 12839 4616 12873 4650
rect 12931 4616 12965 4650
rect 655 3752 689 3786
rect 747 3752 781 3786
rect 839 3752 873 3786
rect 931 3752 965 3786
rect 1023 3752 1057 3786
rect 1114 3752 1148 3786
rect 1206 3752 1240 3786
rect 1299 3752 1333 3786
rect 1391 3752 1425 3786
rect 3197 3743 3231 3777
rect 3289 3743 3323 3777
rect 3381 3743 3415 3777
rect 3473 3743 3507 3777
rect 3565 3743 3599 3777
rect 3657 3743 3691 3777
rect 3749 3743 3783 3777
rect 3841 3743 3875 3777
rect 3933 3743 3967 3777
rect 4025 3743 4059 3777
rect 4117 3743 4151 3777
rect 4209 3743 4243 3777
rect 4301 3743 4335 3777
rect 4393 3743 4427 3777
rect 4485 3743 4519 3777
rect 4577 3743 4611 3777
rect 4669 3743 4703 3777
rect 4761 3743 4795 3777
rect 4853 3743 4887 3777
rect 4945 3743 4979 3777
rect 5018 3743 5052 3777
rect 5110 3743 5144 3777
rect 5202 3743 5236 3777
rect 5294 3743 5328 3777
rect 5386 3743 5420 3777
rect 5478 3743 5512 3777
rect 5570 3743 5604 3777
rect 5662 3743 5696 3777
rect 5754 3743 5788 3777
rect 5846 3743 5880 3777
rect 5938 3743 5972 3777
rect 6030 3743 6064 3777
rect 6122 3743 6156 3777
rect 6214 3743 6248 3777
rect 6306 3743 6340 3777
rect 6398 3743 6432 3777
rect 6490 3743 6524 3777
rect 6582 3743 6616 3777
rect 6674 3743 6708 3777
rect 6766 3743 6800 3777
rect 6858 3743 6892 3777
rect 6950 3743 6984 3777
rect 7042 3743 7076 3777
rect 7134 3743 7168 3777
rect 7226 3743 7260 3777
rect 7318 3743 7352 3777
rect 7410 3743 7444 3777
rect 7502 3743 7536 3777
rect 7594 3743 7628 3777
rect 7686 3743 7720 3777
rect 7778 3743 7812 3777
rect 7870 3743 7904 3777
rect 7962 3743 7996 3777
rect 8054 3743 8088 3777
rect 8146 3743 8180 3777
rect 8238 3743 8272 3777
rect 8330 3743 8364 3777
rect 8422 3743 8456 3777
rect 8514 3743 8548 3777
rect 8606 3743 8640 3777
rect 8698 3743 8732 3777
rect 8790 3743 8824 3777
rect 8882 3743 8916 3777
rect 8974 3743 9008 3777
rect 9066 3743 9100 3777
rect 9158 3743 9192 3777
rect 9250 3743 9284 3777
rect 9342 3743 9376 3777
rect 9434 3743 9468 3777
rect 9526 3743 9560 3777
rect 9618 3743 9652 3777
rect 9710 3743 9744 3777
rect 9802 3743 9836 3777
rect 9894 3743 9928 3777
rect 9986 3743 10020 3777
rect 10078 3743 10112 3777
rect 10170 3743 10204 3777
rect 10262 3743 10296 3777
rect 10354 3743 10388 3777
rect 10446 3743 10480 3777
rect 10538 3743 10572 3777
rect 10630 3743 10664 3777
rect 10722 3743 10756 3777
rect 10814 3743 10848 3777
rect 10906 3743 10940 3777
rect 10998 3743 11032 3777
rect 11090 3743 11124 3777
rect 11182 3743 11216 3777
rect 11274 3743 11308 3777
rect 11366 3743 11400 3777
rect 11458 3743 11492 3777
rect 11550 3743 11584 3777
rect 11642 3743 11676 3777
rect 11734 3743 11768 3777
rect 11826 3743 11860 3777
rect 11918 3743 11952 3777
rect 12010 3743 12044 3777
rect 12102 3743 12136 3777
rect 12194 3743 12228 3777
rect 12286 3743 12320 3777
rect 12378 3743 12412 3777
rect 12470 3743 12504 3777
rect 12562 3743 12596 3777
rect 12654 3743 12688 3777
rect 12746 3743 12780 3777
rect 12838 3743 12872 3777
rect 12930 3743 12964 3777
rect 1062 2870 1096 2904
rect 1154 2870 1188 2904
rect 1246 2870 1280 2904
rect 1338 2870 1372 2904
rect 1430 2870 1464 2904
rect 1522 2870 1556 2904
rect 1614 2870 1648 2904
rect 1706 2870 1740 2904
rect 1798 2870 1832 2904
rect 1890 2870 1924 2904
rect 1982 2870 2016 2904
rect 2074 2870 2108 2904
rect 2166 2870 2200 2904
rect 2258 2870 2292 2904
rect 2350 2870 2384 2904
rect 2442 2870 2476 2904
rect 2534 2870 2568 2904
rect 2626 2870 2660 2904
rect 2718 2870 2752 2904
rect 2810 2870 2844 2904
rect 2902 2870 2936 2904
rect 2994 2870 3028 2904
rect 3086 2870 3120 2904
rect 3178 2870 3212 2904
rect 3270 2870 3304 2904
rect 3362 2870 3396 2904
rect 3454 2870 3488 2904
rect 3546 2870 3580 2904
rect 3638 2870 3672 2904
rect 3730 2870 3764 2904
rect 3822 2870 3856 2904
rect 3914 2870 3948 2904
rect 4006 2870 4040 2904
rect 4098 2870 4132 2904
rect 4190 2870 4224 2904
rect 4282 2870 4316 2904
rect 4374 2870 4408 2904
rect 4466 2870 4500 2904
rect 4558 2870 4592 2904
rect 4650 2870 4684 2904
rect 4742 2870 4776 2904
rect 4834 2870 4868 2904
rect 4926 2870 4960 2904
rect 5018 2870 5052 2904
rect 5110 2870 5144 2904
rect 5202 2870 5236 2904
rect 5294 2870 5328 2904
rect 5386 2870 5420 2904
rect 5478 2870 5512 2904
rect 5570 2870 5604 2904
rect 5662 2870 5696 2904
rect 5754 2870 5788 2904
rect 5846 2870 5880 2904
rect 5938 2870 5972 2904
rect 6030 2870 6064 2904
rect 6122 2870 6156 2904
rect 6214 2870 6248 2904
rect 6306 2870 6340 2904
rect 6398 2870 6432 2904
rect 6490 2870 6524 2904
rect 6582 2870 6616 2904
rect 6674 2870 6708 2904
rect 6766 2870 6800 2904
rect 6858 2870 6892 2904
rect 6950 2870 6984 2904
rect 7042 2870 7076 2904
rect 7134 2870 7168 2904
rect 7226 2870 7260 2904
rect 7318 2870 7352 2904
rect 7410 2870 7444 2904
rect 7502 2870 7536 2904
rect 7594 2870 7628 2904
rect 7686 2870 7720 2904
rect 7778 2870 7812 2904
rect 7870 2870 7904 2904
rect 7962 2870 7996 2904
rect 8054 2870 8088 2904
rect 8146 2870 8180 2904
rect 8238 2870 8272 2904
rect 8330 2870 8364 2904
rect 8422 2870 8456 2904
rect 8514 2870 8548 2904
rect 8606 2870 8640 2904
rect 8698 2870 8732 2904
rect 8790 2870 8824 2904
rect 8882 2870 8916 2904
rect 8974 2870 9008 2904
rect 9066 2870 9100 2904
rect 9158 2870 9192 2904
rect 9250 2870 9284 2904
rect 9342 2870 9376 2904
rect 9434 2870 9468 2904
rect 9526 2870 9560 2904
rect 9618 2870 9652 2904
rect 9710 2870 9744 2904
rect 9802 2870 9836 2904
rect 9894 2870 9928 2904
rect 9986 2870 10020 2904
rect 10078 2870 10112 2904
rect 10170 2870 10204 2904
rect 10262 2870 10296 2904
rect 10354 2870 10388 2904
rect 10446 2870 10480 2904
rect 10538 2870 10572 2904
rect 10630 2870 10664 2904
rect 10722 2870 10756 2904
rect 10814 2870 10848 2904
rect 10906 2870 10940 2904
rect 10998 2870 11032 2904
rect 11090 2870 11124 2904
rect 11182 2870 11216 2904
rect 11274 2870 11308 2904
rect 11366 2870 11400 2904
rect 11458 2870 11492 2904
rect 11550 2870 11584 2904
rect 11642 2870 11676 2904
rect 11734 2870 11768 2904
rect 11826 2870 11860 2904
rect 11918 2870 11952 2904
rect 12010 2870 12044 2904
rect 12102 2870 12136 2904
rect 12194 2870 12228 2904
rect 12286 2870 12320 2904
rect 12378 2870 12412 2904
rect 12470 2870 12504 2904
rect 12562 2870 12596 2904
rect 12654 2870 12688 2904
rect 12746 2870 12780 2904
rect 12838 2870 12872 2904
rect 12930 2870 12964 2904
<< poly >>
rect 1114 6124 1144 6150
rect 1202 6124 1232 6150
rect 1390 6124 1420 6150
rect 1474 6124 1504 6150
rect 1558 6124 1588 6150
rect 1642 6124 1672 6150
rect 1726 6124 1756 6150
rect 2389 6124 2419 6150
rect 2473 6124 2503 6150
rect 2573 6124 2603 6150
rect 2657 6124 2687 6150
rect 2754 6124 2784 6150
rect 2855 6124 2885 6150
rect 2939 6124 2969 6150
rect 3074 6124 3104 6150
rect 1114 5951 1144 5966
rect 1108 5927 1144 5951
rect 1108 5892 1138 5927
rect 1202 5905 1232 5966
rect 1062 5876 1138 5892
rect 1062 5842 1072 5876
rect 1106 5842 1138 5876
rect 1062 5826 1138 5842
rect 1180 5889 1234 5905
rect 1180 5855 1190 5889
rect 1224 5855 1234 5889
rect 1390 5888 1420 5924
rect 1180 5839 1234 5855
rect 1339 5876 1420 5888
rect 1474 5886 1504 5924
rect 1558 5886 1588 5924
rect 1642 5886 1672 5924
rect 1726 5886 1756 5924
rect 1339 5842 1355 5876
rect 1389 5842 1420 5876
rect 1108 5817 1138 5826
rect 1108 5793 1144 5817
rect 1114 5778 1144 5793
rect 1202 5778 1232 5839
rect 1339 5830 1420 5842
rect 1473 5876 1756 5886
rect 1473 5842 1489 5876
rect 1523 5842 1756 5876
rect 1473 5832 1756 5842
rect 1390 5804 1420 5830
rect 1474 5804 1504 5832
rect 1558 5804 1588 5832
rect 1642 5804 1672 5832
rect 1726 5804 1756 5832
rect 2389 5892 2419 5924
rect 2473 5892 2503 5924
rect 2573 5892 2603 5924
rect 2657 5892 2687 5924
rect 2754 5892 2784 5996
rect 2855 5942 2885 6040
rect 2939 6002 2969 6040
rect 2927 5992 2993 6002
rect 3262 6120 3564 6150
rect 3262 6051 3292 6120
rect 3534 6100 3564 6120
rect 3618 6100 3648 6150
rect 3762 6124 3792 6150
rect 3846 6124 3876 6150
rect 3942 6124 3972 6150
rect 4026 6124 4056 6150
rect 3346 6051 3376 6077
rect 2927 5958 2943 5992
rect 2977 5958 2993 5992
rect 2927 5948 2993 5958
rect 2831 5926 2885 5942
rect 2831 5892 2841 5926
rect 2875 5906 2885 5926
rect 3074 5906 3104 5996
rect 3762 6002 3792 6040
rect 3738 5992 3804 6002
rect 3262 5917 3292 5943
rect 2875 5892 2993 5906
rect 2389 5876 2693 5892
rect 2389 5842 2649 5876
rect 2683 5842 2693 5876
rect 2389 5826 2693 5842
rect 2735 5876 2789 5892
rect 2831 5876 2993 5892
rect 2735 5842 2745 5876
rect 2779 5842 2789 5876
rect 2735 5826 2789 5842
rect 2389 5804 2419 5826
rect 2473 5804 2503 5826
rect 2573 5804 2603 5826
rect 2657 5804 2687 5826
rect 2758 5758 2788 5826
rect 2853 5818 2921 5834
rect 2853 5784 2877 5818
rect 2911 5784 2921 5818
rect 2853 5768 2921 5784
rect 2853 5746 2883 5768
rect 2963 5746 2993 5876
rect 3074 5890 3155 5906
rect 3074 5870 3111 5890
rect 3070 5856 3111 5870
rect 3145 5856 3155 5890
rect 3346 5899 3376 5943
rect 3346 5889 3488 5899
rect 3346 5875 3438 5889
rect 3070 5840 3155 5856
rect 3258 5855 3438 5875
rect 3472 5855 3488 5889
rect 3258 5845 3488 5855
rect 3534 5846 3564 5972
rect 3618 5957 3648 5972
rect 3738 5958 3754 5992
rect 3788 5958 3804 5992
rect 3618 5927 3671 5957
rect 3738 5948 3804 5958
rect 3846 5950 3876 6040
rect 3641 5846 3671 5927
rect 3846 5934 3900 5950
rect 3846 5906 3856 5934
rect 3737 5900 3856 5906
rect 3890 5900 3900 5934
rect 3737 5884 3900 5900
rect 3737 5876 3876 5884
rect 3070 5758 3100 5840
rect 3258 5758 3288 5845
rect 3530 5830 3584 5846
rect 3530 5803 3540 5830
rect 3343 5796 3540 5803
rect 3574 5796 3584 5830
rect 3343 5780 3584 5796
rect 3626 5830 3680 5846
rect 3626 5796 3636 5830
rect 3670 5796 3680 5830
rect 3626 5780 3680 5796
rect 3343 5773 3565 5780
rect 3343 5758 3373 5773
rect 3533 5758 3563 5773
rect 3641 5758 3671 5780
rect 3737 5746 3767 5876
rect 3942 5846 3972 5996
rect 4026 5892 4056 5996
rect 4026 5876 4114 5892
rect 3809 5818 3877 5834
rect 3809 5784 3819 5818
rect 3853 5784 3877 5818
rect 3809 5768 3877 5784
rect 3923 5830 3977 5846
rect 3923 5796 3933 5830
rect 3967 5796 3977 5830
rect 3923 5780 3977 5796
rect 4026 5842 4069 5876
rect 4103 5842 4114 5876
rect 4026 5826 4114 5842
rect 3847 5746 3877 5768
rect 3942 5758 3972 5780
rect 4026 5758 4056 5826
rect 1114 5648 1144 5674
rect 1202 5648 1232 5674
rect 1390 5648 1420 5674
rect 1474 5648 1504 5674
rect 1558 5648 1588 5674
rect 1642 5648 1672 5674
rect 1726 5648 1756 5674
rect 2389 5648 2419 5674
rect 2473 5648 2503 5674
rect 2573 5648 2603 5674
rect 2657 5648 2687 5674
rect 2758 5648 2788 5674
rect 2853 5648 2883 5674
rect 2963 5648 2993 5674
rect 3070 5648 3100 5674
rect 3258 5648 3288 5674
rect 3343 5648 3373 5674
rect 3533 5648 3563 5674
rect 3641 5648 3671 5674
rect 3737 5648 3767 5674
rect 3847 5648 3877 5674
rect 3942 5648 3972 5674
rect 4026 5648 4056 5674
rect 2918 5330 2984 5340
rect 2918 5296 2934 5330
rect 2968 5296 2984 5330
rect 4161 5333 4227 5343
rect 2918 5286 2984 5296
rect 4161 5299 4177 5333
rect 4211 5299 4227 5333
rect 6553 5335 6619 5345
rect 4161 5289 4227 5299
rect 6553 5301 6569 5335
rect 6603 5301 6619 5335
rect 8945 5335 9011 5345
rect 6553 5291 6619 5301
rect 8945 5301 8961 5335
rect 8995 5301 9011 5335
rect 11337 5336 11403 5346
rect 8945 5291 9011 5301
rect 11337 5302 11353 5336
rect 11387 5302 11403 5336
rect 11337 5292 11403 5302
rect 1113 5245 1143 5271
rect 1197 5245 1227 5271
rect 1385 5251 1415 5277
rect 1478 5251 1508 5277
rect 1562 5251 1592 5277
rect 1682 5251 1712 5277
rect 1788 5251 1818 5277
rect 1896 5251 1926 5277
rect 1980 5251 2010 5277
rect 2117 5251 2147 5277
rect 2261 5251 2291 5277
rect 2345 5251 2375 5277
rect 2463 5251 2493 5277
rect 2571 5251 2601 5277
rect 2667 5251 2697 5277
rect 2739 5251 2769 5277
rect 1113 5102 1143 5117
rect 1080 5072 1143 5102
rect 1080 5034 1110 5072
rect 1055 5018 1110 5034
rect 1197 5028 1227 5117
rect 1055 4984 1066 5018
rect 1100 4984 1110 5018
rect 1055 4968 1110 4984
rect 1152 5018 1227 5028
rect 1385 5021 1415 5167
rect 1478 5033 1508 5167
rect 1562 5129 1592 5167
rect 1682 5135 1712 5167
rect 1550 5119 1616 5129
rect 1550 5085 1566 5119
rect 1600 5085 1616 5119
rect 1550 5075 1616 5085
rect 1682 5119 1746 5135
rect 1682 5085 1702 5119
rect 1736 5085 1746 5119
rect 1682 5069 1746 5085
rect 1152 4984 1168 5018
rect 1202 4984 1227 5018
rect 1152 4974 1227 4984
rect 1080 4930 1110 4968
rect 1080 4900 1143 4930
rect 1113 4885 1143 4900
rect 1197 4885 1227 4974
rect 1374 5005 1428 5021
rect 1374 4971 1384 5005
rect 1418 4971 1428 5005
rect 1478 5003 1616 5033
rect 1374 4955 1428 4971
rect 1586 4973 1616 5003
rect 1385 4885 1415 4955
rect 1480 4945 1544 4961
rect 1480 4911 1500 4945
rect 1534 4911 1544 4945
rect 1480 4895 1544 4911
rect 1586 4957 1640 4973
rect 1586 4923 1596 4957
rect 1630 4923 1640 4957
rect 1586 4907 1640 4923
rect 1480 4873 1510 4895
rect 1586 4873 1616 4907
rect 1682 4885 1712 5069
rect 1788 4983 1818 5167
rect 2261 5135 2291 5167
rect 2237 5119 2291 5135
rect 2345 5129 2375 5167
rect 2463 5135 2493 5167
rect 2237 5085 2247 5119
rect 2281 5085 2291 5119
rect 1896 5051 1926 5083
rect 1980 5051 2010 5083
rect 1860 5035 1926 5051
rect 1860 5001 1870 5035
rect 1904 5001 1926 5035
rect 1860 4985 1926 5001
rect 1976 5035 2066 5051
rect 1976 5001 2022 5035
rect 2056 5001 2066 5035
rect 1976 4985 2066 5001
rect 2117 5017 2147 5083
rect 2237 5069 2291 5085
rect 2333 5119 2399 5129
rect 2333 5085 2349 5119
rect 2383 5085 2399 5119
rect 2333 5075 2399 5085
rect 2463 5119 2529 5135
rect 2463 5085 2485 5119
rect 2519 5085 2529 5119
rect 2261 5033 2291 5069
rect 2463 5069 2529 5085
rect 2117 5001 2194 5017
rect 2261 5003 2398 5033
rect 2117 4987 2150 5001
rect 1758 4967 1818 4983
rect 1758 4933 1768 4967
rect 1802 4947 1818 4967
rect 1802 4933 1822 4947
rect 1758 4917 1822 4933
rect 1892 4929 1922 4985
rect 1976 4929 2006 4985
rect 2140 4967 2150 4987
rect 2184 4967 2194 5001
rect 2140 4951 2194 4967
rect 2164 4929 2194 4951
rect 2259 4945 2326 4961
rect 1792 4885 1822 4917
rect 2259 4911 2282 4945
rect 2316 4911 2326 4945
rect 2259 4895 2326 4911
rect 2259 4873 2289 4895
rect 2368 4873 2398 5003
rect 2463 4885 2493 5069
rect 2571 4983 2601 5167
rect 2937 5183 2967 5286
rect 3034 5251 3064 5277
rect 2667 5035 2697 5083
rect 2535 4967 2601 4983
rect 2643 5019 2697 5035
rect 2739 5051 2769 5083
rect 2739 5035 2835 5051
rect 2739 5021 2791 5035
rect 2643 4985 2653 5019
rect 2687 4985 2697 5019
rect 2643 4969 2697 4985
rect 2535 4933 2545 4967
rect 2579 4933 2601 4967
rect 2535 4917 2601 4933
rect 2667 4929 2697 4969
rect 2751 5001 2791 5021
rect 2825 5001 2835 5035
rect 2937 5023 2967 5055
rect 3222 5235 3252 5261
rect 3317 5251 3347 5277
rect 3222 5091 3252 5107
rect 3196 5061 3252 5091
rect 2751 4985 2835 5001
rect 2906 5007 2970 5023
rect 3034 5019 3064 5051
rect 2751 4929 2781 4985
rect 2906 4973 2922 5007
rect 2956 4973 2970 5007
rect 2906 4957 2970 4973
rect 3012 5013 3064 5019
rect 3196 5013 3226 5061
rect 3505 5245 3535 5271
rect 3589 5245 3619 5271
rect 3777 5251 3807 5277
rect 3870 5251 3900 5277
rect 3954 5251 3984 5277
rect 4074 5251 4104 5277
rect 4180 5251 4210 5289
rect 4288 5251 4318 5277
rect 4372 5251 4402 5277
rect 4509 5251 4539 5277
rect 4653 5251 4683 5277
rect 4737 5251 4767 5277
rect 4855 5251 4885 5277
rect 4963 5251 4993 5277
rect 5059 5251 5089 5277
rect 5131 5251 5161 5277
rect 5426 5251 5456 5277
rect 3505 5102 3535 5117
rect 3472 5072 3535 5102
rect 3317 5019 3347 5051
rect 3472 5034 3502 5072
rect 3012 5003 3226 5013
rect 3012 4969 3022 5003
rect 3056 4969 3226 5003
rect 3012 4959 3226 4969
rect 2549 4885 2579 4917
rect 2939 4885 2969 4957
rect 3012 4953 3064 4959
rect 3034 4931 3064 4953
rect 3196 4930 3226 4959
rect 3288 5003 3347 5019
rect 3288 4969 3298 5003
rect 3332 4969 3347 5003
rect 3288 4953 3347 4969
rect 3447 5018 3502 5034
rect 3589 5028 3619 5117
rect 3447 4984 3458 5018
rect 3492 4984 3502 5018
rect 3447 4968 3502 4984
rect 3544 5018 3619 5028
rect 3777 5021 3807 5167
rect 3870 5033 3900 5167
rect 3954 5129 3984 5167
rect 4074 5135 4104 5167
rect 3942 5119 4008 5129
rect 3942 5085 3958 5119
rect 3992 5085 4008 5119
rect 3942 5075 4008 5085
rect 4074 5119 4138 5135
rect 4074 5085 4094 5119
rect 4128 5085 4138 5119
rect 4074 5069 4138 5085
rect 3544 4984 3560 5018
rect 3594 4984 3619 5018
rect 3544 4974 3619 4984
rect 3317 4931 3347 4953
rect 3196 4900 3252 4930
rect 3222 4885 3252 4900
rect 3472 4930 3502 4968
rect 3472 4900 3535 4930
rect 3505 4885 3535 4900
rect 3589 4885 3619 4974
rect 3766 5005 3820 5021
rect 3766 4971 3776 5005
rect 3810 4971 3820 5005
rect 3870 5003 4008 5033
rect 3766 4955 3820 4971
rect 3978 4973 4008 5003
rect 3777 4885 3807 4955
rect 3872 4945 3936 4961
rect 3872 4911 3892 4945
rect 3926 4911 3936 4945
rect 3872 4895 3936 4911
rect 3978 4957 4032 4973
rect 3978 4923 3988 4957
rect 4022 4923 4032 4957
rect 3978 4907 4032 4923
rect 3872 4873 3902 4895
rect 3978 4873 4008 4907
rect 4074 4885 4104 5069
rect 4180 4983 4210 5167
rect 4653 5135 4683 5167
rect 4629 5119 4683 5135
rect 4737 5129 4767 5167
rect 4855 5135 4885 5167
rect 4629 5085 4639 5119
rect 4673 5085 4683 5119
rect 4288 5051 4318 5083
rect 4372 5051 4402 5083
rect 4252 5035 4318 5051
rect 4252 5001 4262 5035
rect 4296 5001 4318 5035
rect 4252 4985 4318 5001
rect 4368 5035 4458 5051
rect 4368 5001 4414 5035
rect 4448 5001 4458 5035
rect 4368 4985 4458 5001
rect 4509 5017 4539 5083
rect 4629 5069 4683 5085
rect 4725 5119 4791 5129
rect 4725 5085 4741 5119
rect 4775 5085 4791 5119
rect 4725 5075 4791 5085
rect 4855 5119 4921 5135
rect 4855 5085 4877 5119
rect 4911 5085 4921 5119
rect 4653 5033 4683 5069
rect 4855 5069 4921 5085
rect 4509 5001 4586 5017
rect 4653 5003 4790 5033
rect 4509 4987 4542 5001
rect 4150 4967 4210 4983
rect 4150 4933 4160 4967
rect 4194 4947 4210 4967
rect 4194 4933 4214 4947
rect 4150 4917 4214 4933
rect 4284 4929 4314 4985
rect 4368 4929 4398 4985
rect 4532 4967 4542 4987
rect 4576 4967 4586 5001
rect 4532 4951 4586 4967
rect 4556 4929 4586 4951
rect 4651 4945 4718 4961
rect 4184 4885 4214 4917
rect 4651 4911 4674 4945
rect 4708 4911 4718 4945
rect 4651 4895 4718 4911
rect 4651 4873 4681 4895
rect 4760 4873 4790 5003
rect 4855 4885 4885 5069
rect 4963 4983 4993 5167
rect 5329 5183 5359 5209
rect 5059 5035 5089 5083
rect 4927 4967 4993 4983
rect 5035 5019 5089 5035
rect 5131 5051 5161 5083
rect 5131 5035 5227 5051
rect 5131 5021 5183 5035
rect 5035 4985 5045 5019
rect 5079 4985 5089 5019
rect 5035 4969 5089 4985
rect 4927 4933 4937 4967
rect 4971 4933 4993 4967
rect 4927 4917 4993 4933
rect 5059 4929 5089 4969
rect 5143 5001 5183 5021
rect 5217 5001 5227 5035
rect 5329 5023 5359 5055
rect 5614 5235 5644 5261
rect 5709 5251 5739 5277
rect 5614 5091 5644 5107
rect 5588 5061 5644 5091
rect 5143 4985 5227 5001
rect 5298 5007 5362 5023
rect 5426 5019 5456 5051
rect 5143 4929 5173 4985
rect 5298 4973 5314 5007
rect 5348 4973 5362 5007
rect 5298 4957 5362 4973
rect 5404 5013 5456 5019
rect 5588 5013 5618 5061
rect 5897 5245 5927 5271
rect 5981 5245 6011 5271
rect 6169 5251 6199 5277
rect 6262 5251 6292 5277
rect 6346 5251 6376 5277
rect 6466 5251 6496 5277
rect 6572 5251 6602 5291
rect 6680 5251 6710 5277
rect 6764 5251 6794 5277
rect 6901 5251 6931 5277
rect 7045 5251 7075 5277
rect 7129 5251 7159 5277
rect 7247 5251 7277 5277
rect 7355 5251 7385 5277
rect 7451 5251 7481 5277
rect 7523 5251 7553 5277
rect 7818 5251 7848 5277
rect 5897 5102 5927 5117
rect 5864 5072 5927 5102
rect 5709 5019 5739 5051
rect 5864 5034 5894 5072
rect 5404 5003 5618 5013
rect 5404 4969 5414 5003
rect 5448 4969 5618 5003
rect 5404 4959 5618 4969
rect 4941 4885 4971 4917
rect 5331 4885 5361 4957
rect 5404 4953 5456 4959
rect 5426 4931 5456 4953
rect 5588 4930 5618 4959
rect 5680 5003 5739 5019
rect 5680 4969 5690 5003
rect 5724 4969 5739 5003
rect 5680 4953 5739 4969
rect 5839 5018 5894 5034
rect 5981 5028 6011 5117
rect 5839 4984 5850 5018
rect 5884 4984 5894 5018
rect 5839 4968 5894 4984
rect 5936 5018 6011 5028
rect 6169 5021 6199 5167
rect 6262 5033 6292 5167
rect 6346 5129 6376 5167
rect 6466 5135 6496 5167
rect 6334 5119 6400 5129
rect 6334 5085 6350 5119
rect 6384 5085 6400 5119
rect 6334 5075 6400 5085
rect 6466 5119 6530 5135
rect 6466 5085 6486 5119
rect 6520 5085 6530 5119
rect 6466 5069 6530 5085
rect 5936 4984 5952 5018
rect 5986 4984 6011 5018
rect 5936 4974 6011 4984
rect 5709 4931 5739 4953
rect 5588 4900 5644 4930
rect 5614 4885 5644 4900
rect 5864 4930 5894 4968
rect 5864 4900 5927 4930
rect 5897 4885 5927 4900
rect 5981 4885 6011 4974
rect 6158 5005 6212 5021
rect 6158 4971 6168 5005
rect 6202 4971 6212 5005
rect 6262 5003 6400 5033
rect 6158 4955 6212 4971
rect 6370 4973 6400 5003
rect 6169 4885 6199 4955
rect 6264 4945 6328 4961
rect 6264 4911 6284 4945
rect 6318 4911 6328 4945
rect 6264 4895 6328 4911
rect 6370 4957 6424 4973
rect 6370 4923 6380 4957
rect 6414 4923 6424 4957
rect 6370 4907 6424 4923
rect 6264 4873 6294 4895
rect 6370 4873 6400 4907
rect 6466 4885 6496 5069
rect 6572 4983 6602 5167
rect 7045 5135 7075 5167
rect 7021 5119 7075 5135
rect 7129 5129 7159 5167
rect 7247 5135 7277 5167
rect 7021 5085 7031 5119
rect 7065 5085 7075 5119
rect 6680 5051 6710 5083
rect 6764 5051 6794 5083
rect 6644 5035 6710 5051
rect 6644 5001 6654 5035
rect 6688 5001 6710 5035
rect 6644 4985 6710 5001
rect 6760 5035 6850 5051
rect 6760 5001 6806 5035
rect 6840 5001 6850 5035
rect 6760 4985 6850 5001
rect 6901 5017 6931 5083
rect 7021 5069 7075 5085
rect 7117 5119 7183 5129
rect 7117 5085 7133 5119
rect 7167 5085 7183 5119
rect 7117 5075 7183 5085
rect 7247 5119 7313 5135
rect 7247 5085 7269 5119
rect 7303 5085 7313 5119
rect 7045 5033 7075 5069
rect 7247 5069 7313 5085
rect 6901 5001 6978 5017
rect 7045 5003 7182 5033
rect 6901 4987 6934 5001
rect 6542 4967 6602 4983
rect 6542 4933 6552 4967
rect 6586 4947 6602 4967
rect 6586 4933 6606 4947
rect 6542 4917 6606 4933
rect 6676 4929 6706 4985
rect 6760 4929 6790 4985
rect 6924 4967 6934 4987
rect 6968 4967 6978 5001
rect 6924 4951 6978 4967
rect 6948 4929 6978 4951
rect 7043 4945 7110 4961
rect 6576 4885 6606 4917
rect 7043 4911 7066 4945
rect 7100 4911 7110 4945
rect 7043 4895 7110 4911
rect 7043 4873 7073 4895
rect 7152 4873 7182 5003
rect 7247 4885 7277 5069
rect 7355 4983 7385 5167
rect 7721 5183 7751 5209
rect 7451 5035 7481 5083
rect 7319 4967 7385 4983
rect 7427 5019 7481 5035
rect 7523 5051 7553 5083
rect 7523 5035 7619 5051
rect 7523 5021 7575 5035
rect 7427 4985 7437 5019
rect 7471 4985 7481 5019
rect 7427 4969 7481 4985
rect 7319 4933 7329 4967
rect 7363 4933 7385 4967
rect 7319 4917 7385 4933
rect 7451 4929 7481 4969
rect 7535 5001 7575 5021
rect 7609 5001 7619 5035
rect 7721 5023 7751 5055
rect 8006 5235 8036 5261
rect 8101 5251 8131 5277
rect 8006 5091 8036 5107
rect 7980 5061 8036 5091
rect 7535 4985 7619 5001
rect 7690 5007 7754 5023
rect 7818 5019 7848 5051
rect 7535 4929 7565 4985
rect 7690 4973 7706 5007
rect 7740 4973 7754 5007
rect 7690 4957 7754 4973
rect 7796 5013 7848 5019
rect 7980 5013 8010 5061
rect 8289 5245 8319 5271
rect 8373 5245 8403 5271
rect 8561 5251 8591 5277
rect 8654 5251 8684 5277
rect 8738 5251 8768 5277
rect 8858 5251 8888 5277
rect 8964 5251 8994 5291
rect 9072 5251 9102 5277
rect 9156 5251 9186 5277
rect 9293 5251 9323 5277
rect 9437 5251 9467 5277
rect 9521 5251 9551 5277
rect 9639 5251 9669 5277
rect 9747 5251 9777 5277
rect 9843 5251 9873 5277
rect 9915 5251 9945 5277
rect 10210 5251 10240 5277
rect 8289 5102 8319 5117
rect 8256 5072 8319 5102
rect 8101 5019 8131 5051
rect 8256 5034 8286 5072
rect 7796 5003 8010 5013
rect 7796 4969 7806 5003
rect 7840 4969 8010 5003
rect 7796 4959 8010 4969
rect 7333 4885 7363 4917
rect 7723 4885 7753 4957
rect 7796 4953 7848 4959
rect 7818 4931 7848 4953
rect 7980 4930 8010 4959
rect 8072 5003 8131 5019
rect 8072 4969 8082 5003
rect 8116 4969 8131 5003
rect 8072 4953 8131 4969
rect 8231 5018 8286 5034
rect 8373 5028 8403 5117
rect 8231 4984 8242 5018
rect 8276 4984 8286 5018
rect 8231 4968 8286 4984
rect 8328 5018 8403 5028
rect 8561 5021 8591 5167
rect 8654 5033 8684 5167
rect 8738 5129 8768 5167
rect 8858 5135 8888 5167
rect 8726 5119 8792 5129
rect 8726 5085 8742 5119
rect 8776 5085 8792 5119
rect 8726 5075 8792 5085
rect 8858 5119 8922 5135
rect 8858 5085 8878 5119
rect 8912 5085 8922 5119
rect 8858 5069 8922 5085
rect 8328 4984 8344 5018
rect 8378 4984 8403 5018
rect 8328 4974 8403 4984
rect 8101 4931 8131 4953
rect 7980 4900 8036 4930
rect 8006 4885 8036 4900
rect 8256 4930 8286 4968
rect 8256 4900 8319 4930
rect 8289 4885 8319 4900
rect 8373 4885 8403 4974
rect 8550 5005 8604 5021
rect 8550 4971 8560 5005
rect 8594 4971 8604 5005
rect 8654 5003 8792 5033
rect 8550 4955 8604 4971
rect 8762 4973 8792 5003
rect 8561 4885 8591 4955
rect 8656 4945 8720 4961
rect 8656 4911 8676 4945
rect 8710 4911 8720 4945
rect 8656 4895 8720 4911
rect 8762 4957 8816 4973
rect 8762 4923 8772 4957
rect 8806 4923 8816 4957
rect 8762 4907 8816 4923
rect 8656 4873 8686 4895
rect 8762 4873 8792 4907
rect 8858 4885 8888 5069
rect 8964 4983 8994 5167
rect 9437 5135 9467 5167
rect 9413 5119 9467 5135
rect 9521 5129 9551 5167
rect 9639 5135 9669 5167
rect 9413 5085 9423 5119
rect 9457 5085 9467 5119
rect 9072 5051 9102 5083
rect 9156 5051 9186 5083
rect 9036 5035 9102 5051
rect 9036 5001 9046 5035
rect 9080 5001 9102 5035
rect 9036 4985 9102 5001
rect 9152 5035 9242 5051
rect 9152 5001 9198 5035
rect 9232 5001 9242 5035
rect 9152 4985 9242 5001
rect 9293 5017 9323 5083
rect 9413 5069 9467 5085
rect 9509 5119 9575 5129
rect 9509 5085 9525 5119
rect 9559 5085 9575 5119
rect 9509 5075 9575 5085
rect 9639 5119 9705 5135
rect 9639 5085 9661 5119
rect 9695 5085 9705 5119
rect 9437 5033 9467 5069
rect 9639 5069 9705 5085
rect 9293 5001 9370 5017
rect 9437 5003 9574 5033
rect 9293 4987 9326 5001
rect 8934 4967 8994 4983
rect 8934 4933 8944 4967
rect 8978 4947 8994 4967
rect 8978 4933 8998 4947
rect 8934 4917 8998 4933
rect 9068 4929 9098 4985
rect 9152 4929 9182 4985
rect 9316 4967 9326 4987
rect 9360 4967 9370 5001
rect 9316 4951 9370 4967
rect 9340 4929 9370 4951
rect 9435 4945 9502 4961
rect 8968 4885 8998 4917
rect 9435 4911 9458 4945
rect 9492 4911 9502 4945
rect 9435 4895 9502 4911
rect 9435 4873 9465 4895
rect 9544 4873 9574 5003
rect 9639 4885 9669 5069
rect 9747 4983 9777 5167
rect 10113 5183 10143 5209
rect 9843 5035 9873 5083
rect 9711 4967 9777 4983
rect 9819 5019 9873 5035
rect 9915 5051 9945 5083
rect 9915 5035 10011 5051
rect 9915 5021 9967 5035
rect 9819 4985 9829 5019
rect 9863 4985 9873 5019
rect 9819 4969 9873 4985
rect 9711 4933 9721 4967
rect 9755 4933 9777 4967
rect 9711 4917 9777 4933
rect 9843 4929 9873 4969
rect 9927 5001 9967 5021
rect 10001 5001 10011 5035
rect 10113 5023 10143 5055
rect 10398 5235 10428 5261
rect 10493 5251 10523 5277
rect 10398 5091 10428 5107
rect 10372 5061 10428 5091
rect 9927 4985 10011 5001
rect 10082 5007 10146 5023
rect 10210 5019 10240 5051
rect 9927 4929 9957 4985
rect 10082 4973 10098 5007
rect 10132 4973 10146 5007
rect 10082 4957 10146 4973
rect 10188 5013 10240 5019
rect 10372 5013 10402 5061
rect 10681 5245 10711 5271
rect 10765 5245 10795 5271
rect 10953 5251 10983 5277
rect 11046 5251 11076 5277
rect 11130 5251 11160 5277
rect 11250 5251 11280 5277
rect 11356 5251 11386 5292
rect 11464 5251 11494 5277
rect 11548 5251 11578 5277
rect 11685 5251 11715 5277
rect 11829 5251 11859 5277
rect 11913 5251 11943 5277
rect 12031 5251 12061 5277
rect 12139 5251 12169 5277
rect 12235 5251 12265 5277
rect 12307 5251 12337 5277
rect 12602 5251 12632 5277
rect 10681 5102 10711 5117
rect 10648 5072 10711 5102
rect 10493 5019 10523 5051
rect 10648 5034 10678 5072
rect 10188 5003 10402 5013
rect 10188 4969 10198 5003
rect 10232 4969 10402 5003
rect 10188 4959 10402 4969
rect 9725 4885 9755 4917
rect 10115 4885 10145 4957
rect 10188 4953 10240 4959
rect 10210 4931 10240 4953
rect 10372 4930 10402 4959
rect 10464 5003 10523 5019
rect 10464 4969 10474 5003
rect 10508 4969 10523 5003
rect 10464 4953 10523 4969
rect 10623 5018 10678 5034
rect 10765 5028 10795 5117
rect 10623 4984 10634 5018
rect 10668 4984 10678 5018
rect 10623 4968 10678 4984
rect 10720 5018 10795 5028
rect 10953 5021 10983 5167
rect 11046 5033 11076 5167
rect 11130 5129 11160 5167
rect 11250 5135 11280 5167
rect 11118 5119 11184 5129
rect 11118 5085 11134 5119
rect 11168 5085 11184 5119
rect 11118 5075 11184 5085
rect 11250 5119 11314 5135
rect 11250 5085 11270 5119
rect 11304 5085 11314 5119
rect 11250 5069 11314 5085
rect 10720 4984 10736 5018
rect 10770 4984 10795 5018
rect 10720 4974 10795 4984
rect 10493 4931 10523 4953
rect 10372 4900 10428 4930
rect 10398 4885 10428 4900
rect 10648 4930 10678 4968
rect 10648 4900 10711 4930
rect 10681 4885 10711 4900
rect 10765 4885 10795 4974
rect 10942 5005 10996 5021
rect 10942 4971 10952 5005
rect 10986 4971 10996 5005
rect 11046 5003 11184 5033
rect 10942 4955 10996 4971
rect 11154 4973 11184 5003
rect 10953 4885 10983 4955
rect 11048 4945 11112 4961
rect 11048 4911 11068 4945
rect 11102 4911 11112 4945
rect 11048 4895 11112 4911
rect 11154 4957 11208 4973
rect 11154 4923 11164 4957
rect 11198 4923 11208 4957
rect 11154 4907 11208 4923
rect 11048 4873 11078 4895
rect 11154 4873 11184 4907
rect 11250 4885 11280 5069
rect 11356 4983 11386 5167
rect 11829 5135 11859 5167
rect 11805 5119 11859 5135
rect 11913 5129 11943 5167
rect 12031 5135 12061 5167
rect 11805 5085 11815 5119
rect 11849 5085 11859 5119
rect 11464 5051 11494 5083
rect 11548 5051 11578 5083
rect 11428 5035 11494 5051
rect 11428 5001 11438 5035
rect 11472 5001 11494 5035
rect 11428 4985 11494 5001
rect 11544 5035 11634 5051
rect 11544 5001 11590 5035
rect 11624 5001 11634 5035
rect 11544 4985 11634 5001
rect 11685 5017 11715 5083
rect 11805 5069 11859 5085
rect 11901 5119 11967 5129
rect 11901 5085 11917 5119
rect 11951 5085 11967 5119
rect 11901 5075 11967 5085
rect 12031 5119 12097 5135
rect 12031 5085 12053 5119
rect 12087 5085 12097 5119
rect 11829 5033 11859 5069
rect 12031 5069 12097 5085
rect 11685 5001 11762 5017
rect 11829 5003 11966 5033
rect 11685 4987 11718 5001
rect 11326 4967 11386 4983
rect 11326 4933 11336 4967
rect 11370 4947 11386 4967
rect 11370 4933 11390 4947
rect 11326 4917 11390 4933
rect 11460 4929 11490 4985
rect 11544 4929 11574 4985
rect 11708 4967 11718 4987
rect 11752 4967 11762 5001
rect 11708 4951 11762 4967
rect 11732 4929 11762 4951
rect 11827 4945 11894 4961
rect 11360 4885 11390 4917
rect 11827 4911 11850 4945
rect 11884 4911 11894 4945
rect 11827 4895 11894 4911
rect 11827 4873 11857 4895
rect 11936 4873 11966 5003
rect 12031 4885 12061 5069
rect 12139 4983 12169 5167
rect 12505 5183 12535 5209
rect 12235 5035 12265 5083
rect 12103 4967 12169 4983
rect 12211 5019 12265 5035
rect 12307 5051 12337 5083
rect 12307 5035 12403 5051
rect 12307 5021 12359 5035
rect 12211 4985 12221 5019
rect 12255 4985 12265 5019
rect 12211 4969 12265 4985
rect 12103 4933 12113 4967
rect 12147 4933 12169 4967
rect 12103 4917 12169 4933
rect 12235 4929 12265 4969
rect 12319 5001 12359 5021
rect 12393 5001 12403 5035
rect 12505 5023 12535 5055
rect 12790 5235 12820 5261
rect 12885 5251 12915 5277
rect 12790 5091 12820 5107
rect 12764 5061 12820 5091
rect 12319 4985 12403 5001
rect 12474 5007 12538 5023
rect 12602 5019 12632 5051
rect 12319 4929 12349 4985
rect 12474 4973 12490 5007
rect 12524 4973 12538 5007
rect 12474 4957 12538 4973
rect 12580 5013 12632 5019
rect 12764 5013 12794 5061
rect 12885 5019 12915 5051
rect 12580 5003 12794 5013
rect 12580 4969 12590 5003
rect 12624 4969 12794 5003
rect 12580 4959 12794 4969
rect 12117 4885 12147 4917
rect 12507 4885 12537 4957
rect 12580 4953 12632 4959
rect 12602 4931 12632 4953
rect 12764 4930 12794 4959
rect 12856 5003 12915 5019
rect 12856 4969 12866 5003
rect 12900 4969 12915 5003
rect 12856 4953 12915 4969
rect 12885 4931 12915 4953
rect 12764 4900 12820 4930
rect 12790 4885 12820 4900
rect 1113 4775 1143 4801
rect 1197 4775 1227 4801
rect 1385 4775 1415 4801
rect 1480 4775 1510 4801
rect 1586 4775 1616 4801
rect 1682 4775 1712 4801
rect 1792 4775 1822 4801
rect 1892 4775 1922 4801
rect 1976 4775 2006 4801
rect 2164 4775 2194 4801
rect 2259 4775 2289 4801
rect 2368 4775 2398 4801
rect 2463 4775 2493 4801
rect 2549 4775 2579 4801
rect 2667 4775 2697 4801
rect 2751 4775 2781 4801
rect 2939 4775 2969 4801
rect 3034 4775 3064 4801
rect 3222 4775 3252 4801
rect 3317 4775 3347 4801
rect 3505 4775 3535 4801
rect 3589 4775 3619 4801
rect 3777 4775 3807 4801
rect 3872 4775 3902 4801
rect 3978 4775 4008 4801
rect 4074 4775 4104 4801
rect 4184 4775 4214 4801
rect 4284 4775 4314 4801
rect 4368 4775 4398 4801
rect 4556 4775 4586 4801
rect 4651 4775 4681 4801
rect 4760 4775 4790 4801
rect 4855 4775 4885 4801
rect 4941 4775 4971 4801
rect 5059 4775 5089 4801
rect 5143 4775 5173 4801
rect 5331 4775 5361 4801
rect 5426 4775 5456 4801
rect 5614 4775 5644 4801
rect 5709 4775 5739 4801
rect 5897 4775 5927 4801
rect 5981 4775 6011 4801
rect 6169 4775 6199 4801
rect 6264 4775 6294 4801
rect 6370 4775 6400 4801
rect 6466 4775 6496 4801
rect 6576 4775 6606 4801
rect 6676 4775 6706 4801
rect 6760 4775 6790 4801
rect 6948 4775 6978 4801
rect 7043 4775 7073 4801
rect 7152 4775 7182 4801
rect 7247 4775 7277 4801
rect 7333 4775 7363 4801
rect 7451 4775 7481 4801
rect 7535 4775 7565 4801
rect 7723 4775 7753 4801
rect 7818 4775 7848 4801
rect 8006 4775 8036 4801
rect 8101 4775 8131 4801
rect 8289 4775 8319 4801
rect 8373 4775 8403 4801
rect 8561 4775 8591 4801
rect 8656 4775 8686 4801
rect 8762 4775 8792 4801
rect 8858 4775 8888 4801
rect 8968 4775 8998 4801
rect 9068 4775 9098 4801
rect 9152 4775 9182 4801
rect 9340 4775 9370 4801
rect 9435 4775 9465 4801
rect 9544 4775 9574 4801
rect 9639 4775 9669 4801
rect 9725 4775 9755 4801
rect 9843 4775 9873 4801
rect 9927 4775 9957 4801
rect 10115 4775 10145 4801
rect 10210 4775 10240 4801
rect 10398 4775 10428 4801
rect 10493 4775 10523 4801
rect 10681 4775 10711 4801
rect 10765 4775 10795 4801
rect 10953 4775 10983 4801
rect 11048 4775 11078 4801
rect 11154 4775 11184 4801
rect 11250 4775 11280 4801
rect 11360 4775 11390 4801
rect 11460 4775 11490 4801
rect 11544 4775 11574 4801
rect 11732 4775 11762 4801
rect 11827 4775 11857 4801
rect 11936 4775 11966 4801
rect 12031 4775 12061 4801
rect 12117 4775 12147 4801
rect 12235 4775 12265 4801
rect 12319 4775 12349 4801
rect 12507 4775 12537 4801
rect 12602 4775 12632 4801
rect 12790 4775 12820 4801
rect 12885 4775 12915 4801
rect 4232 4647 4298 4657
rect 4232 4613 4248 4647
rect 4282 4613 4298 4647
rect 6624 4647 6690 4657
rect 4232 4603 4298 4613
rect 6624 4613 6640 4647
rect 6674 4613 6690 4647
rect 9016 4647 9082 4657
rect 6624 4603 6690 4613
rect 9016 4613 9032 4647
rect 9066 4613 9082 4647
rect 11408 4647 11474 4657
rect 9016 4603 9082 4613
rect 11408 4613 11424 4647
rect 11458 4613 11474 4647
rect 11408 4603 11474 4613
rect 673 4562 703 4588
rect 761 4562 791 4588
rect 949 4562 979 4588
rect 1033 4562 1063 4588
rect 1117 4562 1147 4588
rect 1201 4562 1231 4588
rect 1285 4562 1315 4588
rect 1481 4562 1511 4588
rect 1565 4562 1595 4588
rect 1649 4562 1679 4588
rect 1733 4562 1763 4588
rect 1817 4562 1847 4588
rect 1901 4562 1931 4588
rect 1985 4562 2015 4588
rect 2069 4562 2099 4588
rect 2153 4562 2183 4588
rect 2237 4562 2267 4588
rect 2321 4562 2351 4588
rect 2405 4562 2435 4588
rect 2489 4562 2519 4588
rect 2573 4562 2603 4588
rect 2657 4562 2687 4588
rect 2741 4562 2771 4588
rect 2825 4562 2855 4588
rect 2909 4562 2939 4588
rect 2993 4562 3023 4588
rect 3077 4562 3107 4588
rect 3161 4562 3191 4588
rect 3245 4562 3275 4588
rect 3505 4562 3535 4588
rect 673 4389 703 4404
rect 667 4365 703 4389
rect 667 4330 697 4365
rect 761 4343 791 4404
rect 3600 4546 3630 4572
rect 3788 4562 3818 4588
rect 4083 4562 4113 4588
rect 4155 4562 4185 4588
rect 4251 4562 4281 4603
rect 4359 4562 4389 4588
rect 4477 4562 4507 4588
rect 4561 4562 4591 4588
rect 4705 4562 4735 4588
rect 4842 4562 4872 4588
rect 4926 4562 4956 4588
rect 5034 4562 5064 4588
rect 5140 4562 5170 4588
rect 5260 4562 5290 4588
rect 5344 4562 5374 4588
rect 5437 4562 5467 4588
rect 3600 4402 3630 4418
rect 3600 4372 3656 4402
rect 621 4314 697 4330
rect 621 4280 631 4314
rect 665 4280 697 4314
rect 621 4264 697 4280
rect 739 4327 793 4343
rect 739 4293 749 4327
rect 783 4293 793 4327
rect 949 4326 979 4362
rect 739 4277 793 4293
rect 898 4314 979 4326
rect 1033 4324 1063 4362
rect 1117 4324 1147 4362
rect 1201 4324 1231 4362
rect 1285 4324 1315 4362
rect 898 4280 914 4314
rect 948 4280 979 4314
rect 667 4255 697 4264
rect 667 4231 703 4255
rect 673 4216 703 4231
rect 761 4216 791 4277
rect 898 4268 979 4280
rect 1032 4314 1315 4324
rect 1032 4280 1048 4314
rect 1082 4280 1315 4314
rect 1032 4270 1315 4280
rect 949 4242 979 4268
rect 1033 4242 1063 4270
rect 1117 4242 1147 4270
rect 1201 4242 1231 4270
rect 1285 4242 1315 4270
rect 1481 4324 1511 4362
rect 1565 4324 1595 4362
rect 1649 4324 1679 4362
rect 1733 4324 1763 4362
rect 1817 4324 1847 4362
rect 1901 4324 1931 4362
rect 1481 4314 1931 4324
rect 1481 4280 1505 4314
rect 1539 4280 1573 4314
rect 1607 4280 1641 4314
rect 1675 4280 1709 4314
rect 1743 4280 1777 4314
rect 1811 4280 1845 4314
rect 1879 4280 1931 4314
rect 1481 4270 1931 4280
rect 1481 4242 1511 4270
rect 1565 4242 1595 4270
rect 1649 4242 1679 4270
rect 1733 4242 1763 4270
rect 1817 4242 1847 4270
rect 1901 4242 1931 4270
rect 1985 4324 2015 4362
rect 2069 4324 2099 4362
rect 2153 4324 2183 4362
rect 2237 4324 2267 4362
rect 2321 4324 2351 4362
rect 2405 4324 2435 4362
rect 2489 4324 2519 4362
rect 2573 4324 2603 4362
rect 2657 4324 2687 4362
rect 2741 4324 2771 4362
rect 2825 4324 2855 4362
rect 2909 4324 2939 4362
rect 2993 4324 3023 4362
rect 3077 4324 3107 4362
rect 3161 4324 3191 4362
rect 3245 4324 3275 4362
rect 3505 4330 3535 4362
rect 1985 4314 3279 4324
rect 1985 4280 2005 4314
rect 2039 4280 2073 4314
rect 2107 4280 2141 4314
rect 2175 4280 2209 4314
rect 2243 4280 2277 4314
rect 2311 4280 2345 4314
rect 2379 4280 2413 4314
rect 2447 4280 2481 4314
rect 2515 4280 2549 4314
rect 2583 4280 2617 4314
rect 2651 4280 2685 4314
rect 2719 4280 2753 4314
rect 2787 4280 2821 4314
rect 2855 4280 2889 4314
rect 2923 4280 2957 4314
rect 2991 4280 3025 4314
rect 3059 4280 3093 4314
rect 3127 4280 3161 4314
rect 3195 4280 3229 4314
rect 3263 4280 3279 4314
rect 1985 4270 3279 4280
rect 3505 4314 3564 4330
rect 3505 4280 3520 4314
rect 3554 4280 3564 4314
rect 1985 4242 2015 4270
rect 2069 4242 2099 4270
rect 2153 4242 2183 4270
rect 2237 4242 2267 4270
rect 2321 4242 2351 4270
rect 2405 4242 2435 4270
rect 2489 4242 2519 4270
rect 2573 4242 2603 4270
rect 2657 4242 2687 4270
rect 2741 4242 2771 4270
rect 2825 4242 2855 4270
rect 2909 4242 2939 4270
rect 2993 4242 3023 4270
rect 3077 4242 3107 4270
rect 3161 4242 3191 4270
rect 3245 4242 3275 4270
rect 3505 4264 3564 4280
rect 3626 4324 3656 4372
rect 3885 4494 3915 4520
rect 3788 4330 3818 4362
rect 3885 4334 3915 4366
rect 4083 4362 4113 4394
rect 4017 4346 4113 4362
rect 3788 4324 3840 4330
rect 3626 4314 3840 4324
rect 3626 4280 3796 4314
rect 3830 4280 3840 4314
rect 3626 4270 3840 4280
rect 3505 4242 3535 4264
rect 3626 4241 3656 4270
rect 3788 4264 3840 4270
rect 3882 4318 3946 4334
rect 3882 4284 3896 4318
rect 3930 4284 3946 4318
rect 4017 4312 4027 4346
rect 4061 4332 4113 4346
rect 4155 4346 4185 4394
rect 4061 4312 4101 4332
rect 4017 4296 4101 4312
rect 3882 4268 3946 4284
rect 3788 4242 3818 4264
rect 3600 4211 3656 4241
rect 3600 4196 3630 4211
rect 3883 4196 3913 4268
rect 4071 4240 4101 4296
rect 4155 4330 4209 4346
rect 4155 4296 4165 4330
rect 4199 4296 4209 4330
rect 4155 4280 4209 4296
rect 4251 4294 4281 4478
rect 4359 4446 4389 4478
rect 4323 4430 4389 4446
rect 4477 4440 4507 4478
rect 4561 4446 4591 4478
rect 4323 4396 4333 4430
rect 4367 4396 4389 4430
rect 4323 4380 4389 4396
rect 4453 4430 4519 4440
rect 4453 4396 4469 4430
rect 4503 4396 4519 4430
rect 4453 4386 4519 4396
rect 4561 4430 4615 4446
rect 4561 4396 4571 4430
rect 4605 4396 4615 4430
rect 4155 4240 4185 4280
rect 4251 4278 4317 4294
rect 4251 4244 4273 4278
rect 4307 4244 4317 4278
rect 4251 4228 4317 4244
rect 4273 4196 4303 4228
rect 4359 4196 4389 4380
rect 4561 4380 4615 4396
rect 5625 4556 5655 4582
rect 5709 4556 5739 4582
rect 5897 4562 5927 4588
rect 4561 4344 4591 4380
rect 4454 4314 4591 4344
rect 4705 4328 4735 4394
rect 4842 4362 4872 4394
rect 4926 4362 4956 4394
rect 4454 4184 4484 4314
rect 4658 4312 4735 4328
rect 4658 4278 4668 4312
rect 4702 4298 4735 4312
rect 4786 4346 4876 4362
rect 4786 4312 4796 4346
rect 4830 4312 4876 4346
rect 4702 4278 4712 4298
rect 4786 4296 4876 4312
rect 4926 4346 4992 4362
rect 4926 4312 4948 4346
rect 4982 4312 4992 4346
rect 4926 4296 4992 4312
rect 4526 4256 4593 4272
rect 4526 4222 4536 4256
rect 4570 4222 4593 4256
rect 4658 4262 4712 4278
rect 4658 4240 4688 4262
rect 4846 4240 4876 4296
rect 4930 4240 4960 4296
rect 5034 4294 5064 4478
rect 5140 4446 5170 4478
rect 5106 4430 5170 4446
rect 5260 4440 5290 4478
rect 5106 4396 5116 4430
rect 5150 4396 5170 4430
rect 5106 4380 5170 4396
rect 5236 4430 5302 4440
rect 5236 4396 5252 4430
rect 5286 4396 5302 4430
rect 5236 4386 5302 4396
rect 5034 4278 5094 4294
rect 5034 4258 5050 4278
rect 5030 4244 5050 4258
rect 5084 4244 5094 4278
rect 4526 4206 4593 4222
rect 4563 4184 4593 4206
rect 5030 4228 5094 4244
rect 5030 4196 5060 4228
rect 5140 4196 5170 4380
rect 5344 4344 5374 4478
rect 5236 4314 5374 4344
rect 5437 4332 5467 4478
rect 5625 4339 5655 4428
rect 5709 4413 5739 4428
rect 5709 4383 5772 4413
rect 5742 4345 5772 4383
rect 5992 4546 6022 4572
rect 6180 4562 6210 4588
rect 6475 4562 6505 4588
rect 6547 4562 6577 4588
rect 6643 4562 6673 4603
rect 6751 4562 6781 4588
rect 6869 4562 6899 4588
rect 6953 4562 6983 4588
rect 7097 4562 7127 4588
rect 7234 4562 7264 4588
rect 7318 4562 7348 4588
rect 7426 4562 7456 4588
rect 7532 4562 7562 4588
rect 7652 4562 7682 4588
rect 7736 4562 7766 4588
rect 7829 4562 7859 4588
rect 5992 4402 6022 4418
rect 5992 4372 6048 4402
rect 5424 4316 5478 4332
rect 5236 4284 5266 4314
rect 5212 4268 5266 4284
rect 5424 4282 5434 4316
rect 5468 4282 5478 4316
rect 5212 4234 5222 4268
rect 5256 4234 5266 4268
rect 5212 4218 5266 4234
rect 5236 4184 5266 4218
rect 5308 4256 5372 4272
rect 5424 4266 5478 4282
rect 5625 4329 5700 4339
rect 5625 4295 5650 4329
rect 5684 4295 5700 4329
rect 5625 4285 5700 4295
rect 5742 4329 5797 4345
rect 5742 4295 5752 4329
rect 5786 4295 5797 4329
rect 5308 4222 5318 4256
rect 5352 4222 5372 4256
rect 5308 4206 5372 4222
rect 5342 4184 5372 4206
rect 5437 4196 5467 4266
rect 5625 4196 5655 4285
rect 5742 4279 5797 4295
rect 5897 4330 5927 4362
rect 5897 4314 5956 4330
rect 5897 4280 5912 4314
rect 5946 4280 5956 4314
rect 5742 4241 5772 4279
rect 5897 4264 5956 4280
rect 6018 4324 6048 4372
rect 6277 4494 6307 4520
rect 6180 4330 6210 4362
rect 6277 4334 6307 4366
rect 6475 4362 6505 4394
rect 6409 4346 6505 4362
rect 6180 4324 6232 4330
rect 6018 4314 6232 4324
rect 6018 4280 6188 4314
rect 6222 4280 6232 4314
rect 6018 4270 6232 4280
rect 5897 4242 5927 4264
rect 5709 4211 5772 4241
rect 5709 4196 5739 4211
rect 6018 4241 6048 4270
rect 6180 4264 6232 4270
rect 6274 4318 6338 4334
rect 6274 4284 6288 4318
rect 6322 4284 6338 4318
rect 6409 4312 6419 4346
rect 6453 4332 6505 4346
rect 6547 4346 6577 4394
rect 6453 4312 6493 4332
rect 6409 4296 6493 4312
rect 6274 4268 6338 4284
rect 6180 4242 6210 4264
rect 5992 4211 6048 4241
rect 5992 4196 6022 4211
rect 6275 4196 6305 4268
rect 6463 4240 6493 4296
rect 6547 4330 6601 4346
rect 6547 4296 6557 4330
rect 6591 4296 6601 4330
rect 6547 4280 6601 4296
rect 6643 4294 6673 4478
rect 6751 4446 6781 4478
rect 6715 4430 6781 4446
rect 6869 4440 6899 4478
rect 6953 4446 6983 4478
rect 6715 4396 6725 4430
rect 6759 4396 6781 4430
rect 6715 4380 6781 4396
rect 6845 4430 6911 4440
rect 6845 4396 6861 4430
rect 6895 4396 6911 4430
rect 6845 4386 6911 4396
rect 6953 4430 7007 4446
rect 6953 4396 6963 4430
rect 6997 4396 7007 4430
rect 6547 4240 6577 4280
rect 6643 4278 6709 4294
rect 6643 4244 6665 4278
rect 6699 4244 6709 4278
rect 6643 4228 6709 4244
rect 6665 4196 6695 4228
rect 6751 4196 6781 4380
rect 6953 4380 7007 4396
rect 8017 4556 8047 4582
rect 8101 4556 8131 4582
rect 8289 4562 8319 4588
rect 6953 4344 6983 4380
rect 6846 4314 6983 4344
rect 7097 4328 7127 4394
rect 7234 4362 7264 4394
rect 7318 4362 7348 4394
rect 6846 4184 6876 4314
rect 7050 4312 7127 4328
rect 7050 4278 7060 4312
rect 7094 4298 7127 4312
rect 7178 4346 7268 4362
rect 7178 4312 7188 4346
rect 7222 4312 7268 4346
rect 7094 4278 7104 4298
rect 7178 4296 7268 4312
rect 7318 4346 7384 4362
rect 7318 4312 7340 4346
rect 7374 4312 7384 4346
rect 7318 4296 7384 4312
rect 6918 4256 6985 4272
rect 6918 4222 6928 4256
rect 6962 4222 6985 4256
rect 7050 4262 7104 4278
rect 7050 4240 7080 4262
rect 7238 4240 7268 4296
rect 7322 4240 7352 4296
rect 7426 4294 7456 4478
rect 7532 4446 7562 4478
rect 7498 4430 7562 4446
rect 7652 4440 7682 4478
rect 7498 4396 7508 4430
rect 7542 4396 7562 4430
rect 7498 4380 7562 4396
rect 7628 4430 7694 4440
rect 7628 4396 7644 4430
rect 7678 4396 7694 4430
rect 7628 4386 7694 4396
rect 7426 4278 7486 4294
rect 7426 4258 7442 4278
rect 7422 4244 7442 4258
rect 7476 4244 7486 4278
rect 6918 4206 6985 4222
rect 6955 4184 6985 4206
rect 7422 4228 7486 4244
rect 7422 4196 7452 4228
rect 7532 4196 7562 4380
rect 7736 4344 7766 4478
rect 7628 4314 7766 4344
rect 7829 4332 7859 4478
rect 8017 4339 8047 4428
rect 8101 4413 8131 4428
rect 8101 4383 8164 4413
rect 8134 4345 8164 4383
rect 8384 4546 8414 4572
rect 8572 4562 8602 4588
rect 8867 4562 8897 4588
rect 8939 4562 8969 4588
rect 9035 4562 9065 4603
rect 9143 4562 9173 4588
rect 9261 4562 9291 4588
rect 9345 4562 9375 4588
rect 9489 4562 9519 4588
rect 9626 4562 9656 4588
rect 9710 4562 9740 4588
rect 9818 4562 9848 4588
rect 9924 4562 9954 4588
rect 10044 4562 10074 4588
rect 10128 4562 10158 4588
rect 10221 4562 10251 4588
rect 8384 4402 8414 4418
rect 8384 4372 8440 4402
rect 7816 4316 7870 4332
rect 7628 4284 7658 4314
rect 7604 4268 7658 4284
rect 7816 4282 7826 4316
rect 7860 4282 7870 4316
rect 7604 4234 7614 4268
rect 7648 4234 7658 4268
rect 7604 4218 7658 4234
rect 7628 4184 7658 4218
rect 7700 4256 7764 4272
rect 7816 4266 7870 4282
rect 8017 4329 8092 4339
rect 8017 4295 8042 4329
rect 8076 4295 8092 4329
rect 8017 4285 8092 4295
rect 8134 4329 8189 4345
rect 8134 4295 8144 4329
rect 8178 4295 8189 4329
rect 7700 4222 7710 4256
rect 7744 4222 7764 4256
rect 7700 4206 7764 4222
rect 7734 4184 7764 4206
rect 7829 4196 7859 4266
rect 8017 4196 8047 4285
rect 8134 4279 8189 4295
rect 8289 4330 8319 4362
rect 8289 4314 8348 4330
rect 8289 4280 8304 4314
rect 8338 4280 8348 4314
rect 8134 4241 8164 4279
rect 8289 4264 8348 4280
rect 8410 4324 8440 4372
rect 8669 4494 8699 4520
rect 8572 4330 8602 4362
rect 8669 4334 8699 4366
rect 8867 4362 8897 4394
rect 8801 4346 8897 4362
rect 8572 4324 8624 4330
rect 8410 4314 8624 4324
rect 8410 4280 8580 4314
rect 8614 4280 8624 4314
rect 8410 4270 8624 4280
rect 8289 4242 8319 4264
rect 8101 4211 8164 4241
rect 8101 4196 8131 4211
rect 8410 4241 8440 4270
rect 8572 4264 8624 4270
rect 8666 4318 8730 4334
rect 8666 4284 8680 4318
rect 8714 4284 8730 4318
rect 8801 4312 8811 4346
rect 8845 4332 8897 4346
rect 8939 4346 8969 4394
rect 8845 4312 8885 4332
rect 8801 4296 8885 4312
rect 8666 4268 8730 4284
rect 8572 4242 8602 4264
rect 8384 4211 8440 4241
rect 8384 4196 8414 4211
rect 8667 4196 8697 4268
rect 8855 4240 8885 4296
rect 8939 4330 8993 4346
rect 8939 4296 8949 4330
rect 8983 4296 8993 4330
rect 8939 4280 8993 4296
rect 9035 4294 9065 4478
rect 9143 4446 9173 4478
rect 9107 4430 9173 4446
rect 9261 4440 9291 4478
rect 9345 4446 9375 4478
rect 9107 4396 9117 4430
rect 9151 4396 9173 4430
rect 9107 4380 9173 4396
rect 9237 4430 9303 4440
rect 9237 4396 9253 4430
rect 9287 4396 9303 4430
rect 9237 4386 9303 4396
rect 9345 4430 9399 4446
rect 9345 4396 9355 4430
rect 9389 4396 9399 4430
rect 8939 4240 8969 4280
rect 9035 4278 9101 4294
rect 9035 4244 9057 4278
rect 9091 4244 9101 4278
rect 9035 4228 9101 4244
rect 9057 4196 9087 4228
rect 9143 4196 9173 4380
rect 9345 4380 9399 4396
rect 10409 4556 10439 4582
rect 10493 4556 10523 4582
rect 10681 4562 10711 4588
rect 9345 4344 9375 4380
rect 9238 4314 9375 4344
rect 9489 4328 9519 4394
rect 9626 4362 9656 4394
rect 9710 4362 9740 4394
rect 9238 4184 9268 4314
rect 9442 4312 9519 4328
rect 9442 4278 9452 4312
rect 9486 4298 9519 4312
rect 9570 4346 9660 4362
rect 9570 4312 9580 4346
rect 9614 4312 9660 4346
rect 9486 4278 9496 4298
rect 9570 4296 9660 4312
rect 9710 4346 9776 4362
rect 9710 4312 9732 4346
rect 9766 4312 9776 4346
rect 9710 4296 9776 4312
rect 9310 4256 9377 4272
rect 9310 4222 9320 4256
rect 9354 4222 9377 4256
rect 9442 4262 9496 4278
rect 9442 4240 9472 4262
rect 9630 4240 9660 4296
rect 9714 4240 9744 4296
rect 9818 4294 9848 4478
rect 9924 4446 9954 4478
rect 9890 4430 9954 4446
rect 10044 4440 10074 4478
rect 9890 4396 9900 4430
rect 9934 4396 9954 4430
rect 9890 4380 9954 4396
rect 10020 4430 10086 4440
rect 10020 4396 10036 4430
rect 10070 4396 10086 4430
rect 10020 4386 10086 4396
rect 9818 4278 9878 4294
rect 9818 4258 9834 4278
rect 9814 4244 9834 4258
rect 9868 4244 9878 4278
rect 9310 4206 9377 4222
rect 9347 4184 9377 4206
rect 9814 4228 9878 4244
rect 9814 4196 9844 4228
rect 9924 4196 9954 4380
rect 10128 4344 10158 4478
rect 10020 4314 10158 4344
rect 10221 4332 10251 4478
rect 10409 4339 10439 4428
rect 10493 4413 10523 4428
rect 10493 4383 10556 4413
rect 10526 4345 10556 4383
rect 10776 4546 10806 4572
rect 10964 4562 10994 4588
rect 11259 4562 11289 4588
rect 11331 4562 11361 4588
rect 11427 4562 11457 4603
rect 11535 4562 11565 4588
rect 11653 4562 11683 4588
rect 11737 4562 11767 4588
rect 11881 4562 11911 4588
rect 12018 4562 12048 4588
rect 12102 4562 12132 4588
rect 12210 4562 12240 4588
rect 12316 4562 12346 4588
rect 12436 4562 12466 4588
rect 12520 4562 12550 4588
rect 12613 4562 12643 4588
rect 10776 4402 10806 4418
rect 10776 4372 10832 4402
rect 10208 4316 10262 4332
rect 10020 4284 10050 4314
rect 9996 4268 10050 4284
rect 10208 4282 10218 4316
rect 10252 4282 10262 4316
rect 9996 4234 10006 4268
rect 10040 4234 10050 4268
rect 9996 4218 10050 4234
rect 10020 4184 10050 4218
rect 10092 4256 10156 4272
rect 10208 4266 10262 4282
rect 10409 4329 10484 4339
rect 10409 4295 10434 4329
rect 10468 4295 10484 4329
rect 10409 4285 10484 4295
rect 10526 4329 10581 4345
rect 10526 4295 10536 4329
rect 10570 4295 10581 4329
rect 10092 4222 10102 4256
rect 10136 4222 10156 4256
rect 10092 4206 10156 4222
rect 10126 4184 10156 4206
rect 10221 4196 10251 4266
rect 10409 4196 10439 4285
rect 10526 4279 10581 4295
rect 10681 4330 10711 4362
rect 10681 4314 10740 4330
rect 10681 4280 10696 4314
rect 10730 4280 10740 4314
rect 10526 4241 10556 4279
rect 10681 4264 10740 4280
rect 10802 4324 10832 4372
rect 11061 4494 11091 4520
rect 10964 4330 10994 4362
rect 11061 4334 11091 4366
rect 11259 4362 11289 4394
rect 11193 4346 11289 4362
rect 10964 4324 11016 4330
rect 10802 4314 11016 4324
rect 10802 4280 10972 4314
rect 11006 4280 11016 4314
rect 10802 4270 11016 4280
rect 10681 4242 10711 4264
rect 10493 4211 10556 4241
rect 10493 4196 10523 4211
rect 10802 4241 10832 4270
rect 10964 4264 11016 4270
rect 11058 4318 11122 4334
rect 11058 4284 11072 4318
rect 11106 4284 11122 4318
rect 11193 4312 11203 4346
rect 11237 4332 11289 4346
rect 11331 4346 11361 4394
rect 11237 4312 11277 4332
rect 11193 4296 11277 4312
rect 11058 4268 11122 4284
rect 10964 4242 10994 4264
rect 10776 4211 10832 4241
rect 10776 4196 10806 4211
rect 11059 4196 11089 4268
rect 11247 4240 11277 4296
rect 11331 4330 11385 4346
rect 11331 4296 11341 4330
rect 11375 4296 11385 4330
rect 11331 4280 11385 4296
rect 11427 4294 11457 4478
rect 11535 4446 11565 4478
rect 11499 4430 11565 4446
rect 11653 4440 11683 4478
rect 11737 4446 11767 4478
rect 11499 4396 11509 4430
rect 11543 4396 11565 4430
rect 11499 4380 11565 4396
rect 11629 4430 11695 4440
rect 11629 4396 11645 4430
rect 11679 4396 11695 4430
rect 11629 4386 11695 4396
rect 11737 4430 11791 4446
rect 11737 4396 11747 4430
rect 11781 4396 11791 4430
rect 11331 4240 11361 4280
rect 11427 4278 11493 4294
rect 11427 4244 11449 4278
rect 11483 4244 11493 4278
rect 11427 4228 11493 4244
rect 11449 4196 11479 4228
rect 11535 4196 11565 4380
rect 11737 4380 11791 4396
rect 12801 4556 12831 4582
rect 12885 4556 12915 4582
rect 11737 4344 11767 4380
rect 11630 4314 11767 4344
rect 11881 4328 11911 4394
rect 12018 4362 12048 4394
rect 12102 4362 12132 4394
rect 11630 4184 11660 4314
rect 11834 4312 11911 4328
rect 11834 4278 11844 4312
rect 11878 4298 11911 4312
rect 11962 4346 12052 4362
rect 11962 4312 11972 4346
rect 12006 4312 12052 4346
rect 11878 4278 11888 4298
rect 11962 4296 12052 4312
rect 12102 4346 12168 4362
rect 12102 4312 12124 4346
rect 12158 4312 12168 4346
rect 12102 4296 12168 4312
rect 11702 4256 11769 4272
rect 11702 4222 11712 4256
rect 11746 4222 11769 4256
rect 11834 4262 11888 4278
rect 11834 4240 11864 4262
rect 12022 4240 12052 4296
rect 12106 4240 12136 4296
rect 12210 4294 12240 4478
rect 12316 4446 12346 4478
rect 12282 4430 12346 4446
rect 12436 4440 12466 4478
rect 12282 4396 12292 4430
rect 12326 4396 12346 4430
rect 12282 4380 12346 4396
rect 12412 4430 12478 4440
rect 12412 4396 12428 4430
rect 12462 4396 12478 4430
rect 12412 4386 12478 4396
rect 12210 4278 12270 4294
rect 12210 4258 12226 4278
rect 12206 4244 12226 4258
rect 12260 4244 12270 4278
rect 11702 4206 11769 4222
rect 11739 4184 11769 4206
rect 12206 4228 12270 4244
rect 12206 4196 12236 4228
rect 12316 4196 12346 4380
rect 12520 4344 12550 4478
rect 12412 4314 12550 4344
rect 12613 4332 12643 4478
rect 12801 4339 12831 4428
rect 12885 4413 12915 4428
rect 12885 4383 12948 4413
rect 12918 4345 12948 4383
rect 12600 4316 12654 4332
rect 12412 4284 12442 4314
rect 12388 4268 12442 4284
rect 12600 4282 12610 4316
rect 12644 4282 12654 4316
rect 12388 4234 12398 4268
rect 12432 4234 12442 4268
rect 12388 4218 12442 4234
rect 12412 4184 12442 4218
rect 12484 4256 12548 4272
rect 12600 4266 12654 4282
rect 12801 4329 12876 4339
rect 12801 4295 12826 4329
rect 12860 4295 12876 4329
rect 12801 4285 12876 4295
rect 12918 4329 12973 4345
rect 12918 4295 12928 4329
rect 12962 4295 12973 4329
rect 12484 4222 12494 4256
rect 12528 4222 12548 4256
rect 12484 4206 12548 4222
rect 12518 4184 12548 4206
rect 12613 4196 12643 4266
rect 12801 4196 12831 4285
rect 12918 4279 12973 4295
rect 12918 4241 12948 4279
rect 12885 4211 12948 4241
rect 12885 4196 12915 4211
rect 673 4086 703 4112
rect 761 4086 791 4112
rect 949 4086 979 4112
rect 1033 4086 1063 4112
rect 1117 4086 1147 4112
rect 1201 4086 1231 4112
rect 1285 4086 1315 4112
rect 1481 4086 1511 4112
rect 1565 4086 1595 4112
rect 1649 4086 1679 4112
rect 1733 4086 1763 4112
rect 1817 4086 1847 4112
rect 1901 4086 1931 4112
rect 1985 4086 2015 4112
rect 2069 4086 2099 4112
rect 2153 4086 2183 4112
rect 2237 4086 2267 4112
rect 2321 4086 2351 4112
rect 2405 4086 2435 4112
rect 2489 4086 2519 4112
rect 2573 4086 2603 4112
rect 2657 4086 2687 4112
rect 2741 4086 2771 4112
rect 2825 4086 2855 4112
rect 2909 4086 2939 4112
rect 2993 4086 3023 4112
rect 3077 4086 3107 4112
rect 3161 4086 3191 4112
rect 3245 4086 3275 4112
rect 3505 4086 3535 4112
rect 3600 4086 3630 4112
rect 3788 4086 3818 4112
rect 3883 4086 3913 4112
rect 4071 4086 4101 4112
rect 4155 4086 4185 4112
rect 4273 4086 4303 4112
rect 4359 4086 4389 4112
rect 4454 4086 4484 4112
rect 4563 4086 4593 4112
rect 4658 4086 4688 4112
rect 4846 4086 4876 4112
rect 4930 4086 4960 4112
rect 5030 4086 5060 4112
rect 5140 4086 5170 4112
rect 5236 4086 5266 4112
rect 5342 4086 5372 4112
rect 5437 4086 5467 4112
rect 5625 4086 5655 4112
rect 5709 4086 5739 4112
rect 5897 4086 5927 4112
rect 5992 4086 6022 4112
rect 6180 4086 6210 4112
rect 6275 4086 6305 4112
rect 6463 4086 6493 4112
rect 6547 4086 6577 4112
rect 6665 4086 6695 4112
rect 6751 4086 6781 4112
rect 6846 4086 6876 4112
rect 6955 4086 6985 4112
rect 7050 4086 7080 4112
rect 7238 4086 7268 4112
rect 7322 4086 7352 4112
rect 7422 4086 7452 4112
rect 7532 4086 7562 4112
rect 7628 4086 7658 4112
rect 7734 4086 7764 4112
rect 7829 4086 7859 4112
rect 8017 4086 8047 4112
rect 8101 4086 8131 4112
rect 8289 4086 8319 4112
rect 8384 4086 8414 4112
rect 8572 4086 8602 4112
rect 8667 4086 8697 4112
rect 8855 4086 8885 4112
rect 8939 4086 8969 4112
rect 9057 4086 9087 4112
rect 9143 4086 9173 4112
rect 9238 4086 9268 4112
rect 9347 4086 9377 4112
rect 9442 4086 9472 4112
rect 9630 4086 9660 4112
rect 9714 4086 9744 4112
rect 9814 4086 9844 4112
rect 9924 4086 9954 4112
rect 10020 4086 10050 4112
rect 10126 4086 10156 4112
rect 10221 4086 10251 4112
rect 10409 4086 10439 4112
rect 10493 4086 10523 4112
rect 10681 4086 10711 4112
rect 10776 4086 10806 4112
rect 10964 4086 10994 4112
rect 11059 4086 11089 4112
rect 11247 4086 11277 4112
rect 11331 4086 11361 4112
rect 11449 4086 11479 4112
rect 11535 4086 11565 4112
rect 11630 4086 11660 4112
rect 11739 4086 11769 4112
rect 11834 4086 11864 4112
rect 12022 4086 12052 4112
rect 12106 4086 12136 4112
rect 12206 4086 12236 4112
rect 12316 4086 12346 4112
rect 12412 4086 12442 4112
rect 12518 4086 12548 4112
rect 12613 4086 12643 4112
rect 12801 4086 12831 4112
rect 12885 4086 12915 4112
rect 705 3688 735 3714
rect 793 3688 823 3714
rect 981 3688 1011 3714
rect 1065 3688 1095 3714
rect 1149 3688 1179 3714
rect 1233 3688 1263 3714
rect 1317 3688 1347 3714
rect 3288 3689 3318 3715
rect 705 3515 735 3530
rect 699 3491 735 3515
rect 699 3456 729 3491
rect 793 3469 823 3530
rect 3504 3683 3534 3709
rect 3588 3683 3618 3709
rect 3776 3689 3806 3715
rect 3869 3689 3899 3715
rect 3953 3689 3983 3715
rect 4073 3689 4103 3715
rect 4179 3689 4209 3715
rect 4287 3689 4317 3715
rect 4371 3689 4401 3715
rect 4508 3689 4538 3715
rect 4652 3689 4682 3715
rect 4736 3689 4766 3715
rect 4854 3689 4884 3715
rect 4962 3689 4992 3715
rect 5058 3689 5088 3715
rect 5130 3689 5160 3715
rect 5425 3689 5455 3715
rect 3504 3540 3534 3555
rect 3471 3510 3534 3540
rect 653 3440 729 3456
rect 653 3406 663 3440
rect 697 3406 729 3440
rect 653 3390 729 3406
rect 771 3453 825 3469
rect 771 3419 781 3453
rect 815 3419 825 3453
rect 981 3452 1011 3488
rect 771 3403 825 3419
rect 930 3440 1011 3452
rect 1065 3450 1095 3488
rect 1149 3450 1179 3488
rect 1233 3450 1263 3488
rect 1317 3450 1347 3488
rect 3288 3457 3318 3489
rect 3471 3472 3501 3510
rect 930 3406 946 3440
rect 980 3406 1011 3440
rect 699 3381 729 3390
rect 699 3357 735 3381
rect 705 3342 735 3357
rect 793 3342 823 3403
rect 930 3394 1011 3406
rect 1064 3440 1347 3450
rect 1064 3406 1080 3440
rect 1114 3406 1347 3440
rect 1064 3396 1347 3406
rect 981 3368 1011 3394
rect 1065 3368 1095 3396
rect 1149 3368 1179 3396
rect 1233 3368 1263 3396
rect 1317 3368 1347 3396
rect 3232 3441 3318 3457
rect 3232 3407 3248 3441
rect 3282 3407 3318 3441
rect 3232 3391 3318 3407
rect 3446 3456 3501 3472
rect 3588 3466 3618 3555
rect 3446 3422 3457 3456
rect 3491 3422 3501 3456
rect 3446 3406 3501 3422
rect 3543 3456 3618 3466
rect 3776 3459 3806 3605
rect 3869 3471 3899 3605
rect 3953 3567 3983 3605
rect 4073 3573 4103 3605
rect 3941 3557 4007 3567
rect 3941 3523 3957 3557
rect 3991 3523 4007 3557
rect 3941 3513 4007 3523
rect 4073 3557 4137 3573
rect 4073 3523 4093 3557
rect 4127 3523 4137 3557
rect 4073 3507 4137 3523
rect 3543 3422 3559 3456
rect 3593 3422 3618 3456
rect 3543 3412 3618 3422
rect 3288 3369 3318 3391
rect 3471 3368 3501 3406
rect 3471 3338 3534 3368
rect 3504 3323 3534 3338
rect 3588 3323 3618 3412
rect 3765 3443 3819 3459
rect 3765 3409 3775 3443
rect 3809 3409 3819 3443
rect 3869 3441 4007 3471
rect 3765 3393 3819 3409
rect 3977 3411 4007 3441
rect 3776 3323 3806 3393
rect 3871 3383 3935 3399
rect 3871 3349 3891 3383
rect 3925 3349 3935 3383
rect 3871 3333 3935 3349
rect 3977 3395 4031 3411
rect 3977 3361 3987 3395
rect 4021 3361 4031 3395
rect 3977 3345 4031 3361
rect 3871 3311 3901 3333
rect 3977 3311 4007 3345
rect 4073 3323 4103 3507
rect 4179 3421 4209 3605
rect 4652 3573 4682 3605
rect 4628 3557 4682 3573
rect 4736 3567 4766 3605
rect 4854 3573 4884 3605
rect 4628 3523 4638 3557
rect 4672 3523 4682 3557
rect 4287 3489 4317 3521
rect 4371 3489 4401 3521
rect 4251 3473 4317 3489
rect 4251 3439 4261 3473
rect 4295 3439 4317 3473
rect 4251 3423 4317 3439
rect 4367 3473 4457 3489
rect 4367 3439 4413 3473
rect 4447 3439 4457 3473
rect 4367 3423 4457 3439
rect 4508 3455 4538 3521
rect 4628 3507 4682 3523
rect 4724 3557 4790 3567
rect 4724 3523 4740 3557
rect 4774 3523 4790 3557
rect 4724 3513 4790 3523
rect 4854 3557 4920 3573
rect 4854 3523 4876 3557
rect 4910 3523 4920 3557
rect 4652 3471 4682 3507
rect 4854 3507 4920 3523
rect 4508 3439 4585 3455
rect 4652 3441 4789 3471
rect 4508 3425 4541 3439
rect 4149 3405 4209 3421
rect 4149 3371 4159 3405
rect 4193 3385 4209 3405
rect 4193 3371 4213 3385
rect 4149 3355 4213 3371
rect 4283 3367 4313 3423
rect 4367 3367 4397 3423
rect 4531 3405 4541 3425
rect 4575 3405 4585 3439
rect 4531 3389 4585 3405
rect 4555 3367 4585 3389
rect 4650 3383 4717 3399
rect 4183 3323 4213 3355
rect 4650 3349 4673 3383
rect 4707 3349 4717 3383
rect 4650 3333 4717 3349
rect 4650 3311 4680 3333
rect 4759 3311 4789 3441
rect 4854 3323 4884 3507
rect 4962 3421 4992 3605
rect 5328 3621 5358 3647
rect 5058 3473 5088 3521
rect 4926 3405 4992 3421
rect 5034 3457 5088 3473
rect 5130 3489 5160 3521
rect 5130 3473 5226 3489
rect 5130 3459 5182 3473
rect 5034 3423 5044 3457
rect 5078 3423 5088 3457
rect 5034 3407 5088 3423
rect 4926 3371 4936 3405
rect 4970 3371 4992 3405
rect 4926 3355 4992 3371
rect 5058 3367 5088 3407
rect 5142 3439 5182 3459
rect 5216 3439 5226 3473
rect 5328 3461 5358 3493
rect 5613 3673 5643 3699
rect 5708 3689 5738 3715
rect 5613 3529 5643 3545
rect 5587 3499 5643 3529
rect 5142 3423 5226 3439
rect 5297 3445 5361 3461
rect 5425 3457 5455 3489
rect 5142 3367 5172 3423
rect 5297 3411 5313 3445
rect 5347 3411 5361 3445
rect 5297 3395 5361 3411
rect 5403 3451 5455 3457
rect 5587 3451 5617 3499
rect 5896 3683 5926 3709
rect 5980 3683 6010 3709
rect 6168 3689 6198 3715
rect 6261 3689 6291 3715
rect 6345 3689 6375 3715
rect 6465 3689 6495 3715
rect 6571 3689 6601 3715
rect 6679 3689 6709 3715
rect 6763 3689 6793 3715
rect 6900 3689 6930 3715
rect 7044 3689 7074 3715
rect 7128 3689 7158 3715
rect 7246 3689 7276 3715
rect 7354 3689 7384 3715
rect 7450 3689 7480 3715
rect 7522 3689 7552 3715
rect 7817 3689 7847 3715
rect 5896 3540 5926 3555
rect 5863 3510 5926 3540
rect 5708 3457 5738 3489
rect 5863 3472 5893 3510
rect 5403 3441 5617 3451
rect 5403 3407 5413 3441
rect 5447 3407 5617 3441
rect 5403 3397 5617 3407
rect 4940 3323 4970 3355
rect 5330 3323 5360 3395
rect 5403 3391 5455 3397
rect 5425 3369 5455 3391
rect 5587 3368 5617 3397
rect 5679 3441 5738 3457
rect 5679 3407 5689 3441
rect 5723 3407 5738 3441
rect 5679 3391 5738 3407
rect 5838 3456 5893 3472
rect 5980 3466 6010 3555
rect 5838 3422 5849 3456
rect 5883 3422 5893 3456
rect 5838 3406 5893 3422
rect 5935 3456 6010 3466
rect 6168 3459 6198 3605
rect 6261 3471 6291 3605
rect 6345 3567 6375 3605
rect 6465 3573 6495 3605
rect 6333 3557 6399 3567
rect 6333 3523 6349 3557
rect 6383 3523 6399 3557
rect 6333 3513 6399 3523
rect 6465 3557 6529 3573
rect 6465 3523 6485 3557
rect 6519 3523 6529 3557
rect 6465 3507 6529 3523
rect 5935 3422 5951 3456
rect 5985 3422 6010 3456
rect 5935 3412 6010 3422
rect 5708 3369 5738 3391
rect 5587 3338 5643 3368
rect 5613 3323 5643 3338
rect 5863 3368 5893 3406
rect 5863 3338 5926 3368
rect 5896 3323 5926 3338
rect 5980 3323 6010 3412
rect 6157 3443 6211 3459
rect 6157 3409 6167 3443
rect 6201 3409 6211 3443
rect 6261 3441 6399 3471
rect 6157 3393 6211 3409
rect 6369 3411 6399 3441
rect 6168 3323 6198 3393
rect 6263 3383 6327 3399
rect 6263 3349 6283 3383
rect 6317 3349 6327 3383
rect 6263 3333 6327 3349
rect 6369 3395 6423 3411
rect 6369 3361 6379 3395
rect 6413 3361 6423 3395
rect 6369 3345 6423 3361
rect 6263 3311 6293 3333
rect 6369 3311 6399 3345
rect 6465 3323 6495 3507
rect 6571 3421 6601 3605
rect 7044 3573 7074 3605
rect 7020 3557 7074 3573
rect 7128 3567 7158 3605
rect 7246 3573 7276 3605
rect 7020 3523 7030 3557
rect 7064 3523 7074 3557
rect 6679 3489 6709 3521
rect 6763 3489 6793 3521
rect 6643 3473 6709 3489
rect 6643 3439 6653 3473
rect 6687 3439 6709 3473
rect 6643 3423 6709 3439
rect 6759 3473 6849 3489
rect 6759 3439 6805 3473
rect 6839 3439 6849 3473
rect 6759 3423 6849 3439
rect 6900 3455 6930 3521
rect 7020 3507 7074 3523
rect 7116 3557 7182 3567
rect 7116 3523 7132 3557
rect 7166 3523 7182 3557
rect 7116 3513 7182 3523
rect 7246 3557 7312 3573
rect 7246 3523 7268 3557
rect 7302 3523 7312 3557
rect 7044 3471 7074 3507
rect 7246 3507 7312 3523
rect 6900 3439 6977 3455
rect 7044 3441 7181 3471
rect 6900 3425 6933 3439
rect 6541 3405 6601 3421
rect 6541 3371 6551 3405
rect 6585 3385 6601 3405
rect 6585 3371 6605 3385
rect 6541 3355 6605 3371
rect 6675 3367 6705 3423
rect 6759 3367 6789 3423
rect 6923 3405 6933 3425
rect 6967 3405 6977 3439
rect 6923 3389 6977 3405
rect 6947 3367 6977 3389
rect 7042 3383 7109 3399
rect 6575 3323 6605 3355
rect 7042 3349 7065 3383
rect 7099 3349 7109 3383
rect 7042 3333 7109 3349
rect 7042 3311 7072 3333
rect 7151 3311 7181 3441
rect 7246 3323 7276 3507
rect 7354 3421 7384 3605
rect 7720 3621 7750 3647
rect 7450 3473 7480 3521
rect 7318 3405 7384 3421
rect 7426 3457 7480 3473
rect 7522 3489 7552 3521
rect 7522 3473 7618 3489
rect 7522 3459 7574 3473
rect 7426 3423 7436 3457
rect 7470 3423 7480 3457
rect 7426 3407 7480 3423
rect 7318 3371 7328 3405
rect 7362 3371 7384 3405
rect 7318 3355 7384 3371
rect 7450 3367 7480 3407
rect 7534 3439 7574 3459
rect 7608 3439 7618 3473
rect 7720 3461 7750 3493
rect 8005 3673 8035 3699
rect 8100 3689 8130 3715
rect 8005 3529 8035 3545
rect 7979 3499 8035 3529
rect 7534 3423 7618 3439
rect 7689 3445 7753 3461
rect 7817 3457 7847 3489
rect 7534 3367 7564 3423
rect 7689 3411 7705 3445
rect 7739 3411 7753 3445
rect 7689 3395 7753 3411
rect 7795 3451 7847 3457
rect 7979 3451 8009 3499
rect 8288 3683 8318 3709
rect 8372 3683 8402 3709
rect 8560 3689 8590 3715
rect 8653 3689 8683 3715
rect 8737 3689 8767 3715
rect 8857 3689 8887 3715
rect 8963 3689 8993 3715
rect 9071 3689 9101 3715
rect 9155 3689 9185 3715
rect 9292 3689 9322 3715
rect 9436 3689 9466 3715
rect 9520 3689 9550 3715
rect 9638 3689 9668 3715
rect 9746 3689 9776 3715
rect 9842 3689 9872 3715
rect 9914 3689 9944 3715
rect 10209 3689 10239 3715
rect 8288 3540 8318 3555
rect 8255 3510 8318 3540
rect 8100 3457 8130 3489
rect 8255 3472 8285 3510
rect 7795 3441 8009 3451
rect 7795 3407 7805 3441
rect 7839 3407 8009 3441
rect 7795 3397 8009 3407
rect 7332 3323 7362 3355
rect 7722 3323 7752 3395
rect 7795 3391 7847 3397
rect 7817 3369 7847 3391
rect 7979 3368 8009 3397
rect 8071 3441 8130 3457
rect 8071 3407 8081 3441
rect 8115 3407 8130 3441
rect 8071 3391 8130 3407
rect 8230 3456 8285 3472
rect 8372 3466 8402 3555
rect 8230 3422 8241 3456
rect 8275 3422 8285 3456
rect 8230 3406 8285 3422
rect 8327 3456 8402 3466
rect 8560 3459 8590 3605
rect 8653 3471 8683 3605
rect 8737 3567 8767 3605
rect 8857 3573 8887 3605
rect 8725 3557 8791 3567
rect 8725 3523 8741 3557
rect 8775 3523 8791 3557
rect 8725 3513 8791 3523
rect 8857 3557 8921 3573
rect 8857 3523 8877 3557
rect 8911 3523 8921 3557
rect 8857 3507 8921 3523
rect 8327 3422 8343 3456
rect 8377 3422 8402 3456
rect 8327 3412 8402 3422
rect 8100 3369 8130 3391
rect 7979 3338 8035 3368
rect 8005 3323 8035 3338
rect 8255 3368 8285 3406
rect 8255 3338 8318 3368
rect 8288 3323 8318 3338
rect 8372 3323 8402 3412
rect 8549 3443 8603 3459
rect 8549 3409 8559 3443
rect 8593 3409 8603 3443
rect 8653 3441 8791 3471
rect 8549 3393 8603 3409
rect 8761 3411 8791 3441
rect 8560 3323 8590 3393
rect 8655 3383 8719 3399
rect 8655 3349 8675 3383
rect 8709 3349 8719 3383
rect 8655 3333 8719 3349
rect 8761 3395 8815 3411
rect 8761 3361 8771 3395
rect 8805 3361 8815 3395
rect 8761 3345 8815 3361
rect 8655 3311 8685 3333
rect 8761 3311 8791 3345
rect 8857 3323 8887 3507
rect 8963 3421 8993 3605
rect 9436 3573 9466 3605
rect 9412 3557 9466 3573
rect 9520 3567 9550 3605
rect 9638 3573 9668 3605
rect 9412 3523 9422 3557
rect 9456 3523 9466 3557
rect 9071 3489 9101 3521
rect 9155 3489 9185 3521
rect 9035 3473 9101 3489
rect 9035 3439 9045 3473
rect 9079 3439 9101 3473
rect 9035 3423 9101 3439
rect 9151 3473 9241 3489
rect 9151 3439 9197 3473
rect 9231 3439 9241 3473
rect 9151 3423 9241 3439
rect 9292 3455 9322 3521
rect 9412 3507 9466 3523
rect 9508 3557 9574 3567
rect 9508 3523 9524 3557
rect 9558 3523 9574 3557
rect 9508 3513 9574 3523
rect 9638 3557 9704 3573
rect 9638 3523 9660 3557
rect 9694 3523 9704 3557
rect 9436 3471 9466 3507
rect 9638 3507 9704 3523
rect 9292 3439 9369 3455
rect 9436 3441 9573 3471
rect 9292 3425 9325 3439
rect 8933 3405 8993 3421
rect 8933 3371 8943 3405
rect 8977 3385 8993 3405
rect 8977 3371 8997 3385
rect 8933 3355 8997 3371
rect 9067 3367 9097 3423
rect 9151 3367 9181 3423
rect 9315 3405 9325 3425
rect 9359 3405 9369 3439
rect 9315 3389 9369 3405
rect 9339 3367 9369 3389
rect 9434 3383 9501 3399
rect 8967 3323 8997 3355
rect 9434 3349 9457 3383
rect 9491 3349 9501 3383
rect 9434 3333 9501 3349
rect 9434 3311 9464 3333
rect 9543 3311 9573 3441
rect 9638 3323 9668 3507
rect 9746 3421 9776 3605
rect 10112 3621 10142 3647
rect 9842 3473 9872 3521
rect 9710 3405 9776 3421
rect 9818 3457 9872 3473
rect 9914 3489 9944 3521
rect 9914 3473 10010 3489
rect 9914 3459 9966 3473
rect 9818 3423 9828 3457
rect 9862 3423 9872 3457
rect 9818 3407 9872 3423
rect 9710 3371 9720 3405
rect 9754 3371 9776 3405
rect 9710 3355 9776 3371
rect 9842 3367 9872 3407
rect 9926 3439 9966 3459
rect 10000 3439 10010 3473
rect 10112 3461 10142 3493
rect 10397 3673 10427 3699
rect 10492 3689 10522 3715
rect 10397 3529 10427 3545
rect 10371 3499 10427 3529
rect 9926 3423 10010 3439
rect 10081 3445 10145 3461
rect 10209 3457 10239 3489
rect 9926 3367 9956 3423
rect 10081 3411 10097 3445
rect 10131 3411 10145 3445
rect 10081 3395 10145 3411
rect 10187 3451 10239 3457
rect 10371 3451 10401 3499
rect 10680 3683 10710 3709
rect 10764 3683 10794 3709
rect 10952 3689 10982 3715
rect 11045 3689 11075 3715
rect 11129 3689 11159 3715
rect 11249 3689 11279 3715
rect 11355 3689 11385 3715
rect 11463 3689 11493 3715
rect 11547 3689 11577 3715
rect 11684 3689 11714 3715
rect 11828 3689 11858 3715
rect 11912 3689 11942 3715
rect 12030 3689 12060 3715
rect 12138 3689 12168 3715
rect 12234 3689 12264 3715
rect 12306 3689 12336 3715
rect 12601 3689 12631 3715
rect 10680 3540 10710 3555
rect 10647 3510 10710 3540
rect 10492 3457 10522 3489
rect 10647 3472 10677 3510
rect 10187 3441 10401 3451
rect 10187 3407 10197 3441
rect 10231 3407 10401 3441
rect 10187 3397 10401 3407
rect 9724 3323 9754 3355
rect 10114 3323 10144 3395
rect 10187 3391 10239 3397
rect 10209 3369 10239 3391
rect 10371 3368 10401 3397
rect 10463 3441 10522 3457
rect 10463 3407 10473 3441
rect 10507 3407 10522 3441
rect 10463 3391 10522 3407
rect 10622 3456 10677 3472
rect 10764 3466 10794 3555
rect 10622 3422 10633 3456
rect 10667 3422 10677 3456
rect 10622 3406 10677 3422
rect 10719 3456 10794 3466
rect 10952 3459 10982 3605
rect 11045 3471 11075 3605
rect 11129 3567 11159 3605
rect 11249 3573 11279 3605
rect 11117 3557 11183 3567
rect 11117 3523 11133 3557
rect 11167 3523 11183 3557
rect 11117 3513 11183 3523
rect 11249 3557 11313 3573
rect 11249 3523 11269 3557
rect 11303 3523 11313 3557
rect 11249 3507 11313 3523
rect 10719 3422 10735 3456
rect 10769 3422 10794 3456
rect 10719 3412 10794 3422
rect 10492 3369 10522 3391
rect 10371 3338 10427 3368
rect 10397 3323 10427 3338
rect 10647 3368 10677 3406
rect 10647 3338 10710 3368
rect 10680 3323 10710 3338
rect 10764 3323 10794 3412
rect 10941 3443 10995 3459
rect 10941 3409 10951 3443
rect 10985 3409 10995 3443
rect 11045 3441 11183 3471
rect 10941 3393 10995 3409
rect 11153 3411 11183 3441
rect 10952 3323 10982 3393
rect 11047 3383 11111 3399
rect 11047 3349 11067 3383
rect 11101 3349 11111 3383
rect 11047 3333 11111 3349
rect 11153 3395 11207 3411
rect 11153 3361 11163 3395
rect 11197 3361 11207 3395
rect 11153 3345 11207 3361
rect 11047 3311 11077 3333
rect 11153 3311 11183 3345
rect 11249 3323 11279 3507
rect 11355 3421 11385 3605
rect 11828 3573 11858 3605
rect 11804 3557 11858 3573
rect 11912 3567 11942 3605
rect 12030 3573 12060 3605
rect 11804 3523 11814 3557
rect 11848 3523 11858 3557
rect 11463 3489 11493 3521
rect 11547 3489 11577 3521
rect 11427 3473 11493 3489
rect 11427 3439 11437 3473
rect 11471 3439 11493 3473
rect 11427 3423 11493 3439
rect 11543 3473 11633 3489
rect 11543 3439 11589 3473
rect 11623 3439 11633 3473
rect 11543 3423 11633 3439
rect 11684 3455 11714 3521
rect 11804 3507 11858 3523
rect 11900 3557 11966 3567
rect 11900 3523 11916 3557
rect 11950 3523 11966 3557
rect 11900 3513 11966 3523
rect 12030 3557 12096 3573
rect 12030 3523 12052 3557
rect 12086 3523 12096 3557
rect 11828 3471 11858 3507
rect 12030 3507 12096 3523
rect 11684 3439 11761 3455
rect 11828 3441 11965 3471
rect 11684 3425 11717 3439
rect 11325 3405 11385 3421
rect 11325 3371 11335 3405
rect 11369 3385 11385 3405
rect 11369 3371 11389 3385
rect 11325 3355 11389 3371
rect 11459 3367 11489 3423
rect 11543 3367 11573 3423
rect 11707 3405 11717 3425
rect 11751 3405 11761 3439
rect 11707 3389 11761 3405
rect 11731 3367 11761 3389
rect 11826 3383 11893 3399
rect 11359 3323 11389 3355
rect 11826 3349 11849 3383
rect 11883 3349 11893 3383
rect 11826 3333 11893 3349
rect 11826 3311 11856 3333
rect 11935 3311 11965 3441
rect 12030 3323 12060 3507
rect 12138 3421 12168 3605
rect 12504 3621 12534 3647
rect 12234 3473 12264 3521
rect 12102 3405 12168 3421
rect 12210 3457 12264 3473
rect 12306 3489 12336 3521
rect 12306 3473 12402 3489
rect 12306 3459 12358 3473
rect 12210 3423 12220 3457
rect 12254 3423 12264 3457
rect 12210 3407 12264 3423
rect 12102 3371 12112 3405
rect 12146 3371 12168 3405
rect 12102 3355 12168 3371
rect 12234 3367 12264 3407
rect 12318 3439 12358 3459
rect 12392 3439 12402 3473
rect 12504 3461 12534 3493
rect 12789 3673 12819 3699
rect 12884 3689 12914 3715
rect 12789 3529 12819 3545
rect 12763 3499 12819 3529
rect 12318 3423 12402 3439
rect 12473 3445 12537 3461
rect 12601 3457 12631 3489
rect 12318 3367 12348 3423
rect 12473 3411 12489 3445
rect 12523 3411 12537 3445
rect 12473 3395 12537 3411
rect 12579 3451 12631 3457
rect 12763 3451 12793 3499
rect 12884 3457 12914 3489
rect 12579 3441 12793 3451
rect 12579 3407 12589 3441
rect 12623 3407 12793 3441
rect 12579 3397 12793 3407
rect 12116 3323 12146 3355
rect 12506 3323 12536 3395
rect 12579 3391 12631 3397
rect 12601 3369 12631 3391
rect 12763 3368 12793 3397
rect 12855 3441 12914 3457
rect 12855 3407 12865 3441
rect 12899 3407 12914 3441
rect 12855 3391 12914 3407
rect 12884 3369 12914 3391
rect 12763 3338 12819 3368
rect 12789 3323 12819 3338
rect 705 3212 735 3238
rect 793 3212 823 3238
rect 981 3212 1011 3238
rect 1065 3212 1095 3238
rect 1149 3212 1179 3238
rect 1233 3212 1263 3238
rect 1317 3212 1347 3238
rect 3288 3213 3318 3239
rect 3504 3213 3534 3239
rect 3588 3213 3618 3239
rect 3776 3213 3806 3239
rect 3871 3213 3901 3239
rect 3977 3213 4007 3239
rect 4073 3213 4103 3239
rect 4183 3213 4213 3239
rect 4283 3213 4313 3239
rect 4367 3213 4397 3239
rect 4555 3213 4585 3239
rect 4650 3213 4680 3239
rect 4759 3213 4789 3239
rect 4854 3213 4884 3239
rect 4940 3213 4970 3239
rect 5058 3213 5088 3239
rect 5142 3213 5172 3239
rect 5330 3213 5360 3239
rect 5425 3213 5455 3239
rect 5613 3213 5643 3239
rect 5708 3213 5738 3239
rect 5896 3213 5926 3239
rect 5980 3213 6010 3239
rect 6168 3213 6198 3239
rect 6263 3213 6293 3239
rect 6369 3213 6399 3239
rect 6465 3213 6495 3239
rect 6575 3213 6605 3239
rect 6675 3213 6705 3239
rect 6759 3213 6789 3239
rect 6947 3213 6977 3239
rect 7042 3213 7072 3239
rect 7151 3213 7181 3239
rect 7246 3213 7276 3239
rect 7332 3213 7362 3239
rect 7450 3213 7480 3239
rect 7534 3213 7564 3239
rect 7722 3213 7752 3239
rect 7817 3213 7847 3239
rect 8005 3213 8035 3239
rect 8100 3213 8130 3239
rect 8288 3213 8318 3239
rect 8372 3213 8402 3239
rect 8560 3213 8590 3239
rect 8655 3213 8685 3239
rect 8761 3213 8791 3239
rect 8857 3213 8887 3239
rect 8967 3213 8997 3239
rect 9067 3213 9097 3239
rect 9151 3213 9181 3239
rect 9339 3213 9369 3239
rect 9434 3213 9464 3239
rect 9543 3213 9573 3239
rect 9638 3213 9668 3239
rect 9724 3213 9754 3239
rect 9842 3213 9872 3239
rect 9926 3213 9956 3239
rect 10114 3213 10144 3239
rect 10209 3213 10239 3239
rect 10397 3213 10427 3239
rect 10492 3213 10522 3239
rect 10680 3213 10710 3239
rect 10764 3213 10794 3239
rect 10952 3213 10982 3239
rect 11047 3213 11077 3239
rect 11153 3213 11183 3239
rect 11249 3213 11279 3239
rect 11359 3213 11389 3239
rect 11459 3213 11489 3239
rect 11543 3213 11573 3239
rect 11731 3213 11761 3239
rect 11826 3213 11856 3239
rect 11935 3213 11965 3239
rect 12030 3213 12060 3239
rect 12116 3213 12146 3239
rect 12234 3213 12264 3239
rect 12318 3213 12348 3239
rect 12506 3213 12536 3239
rect 12601 3213 12631 3239
rect 12789 3213 12819 3239
rect 12884 3213 12914 3239
rect 1112 2816 1142 2842
rect 1207 2800 1237 2826
rect 1395 2816 1425 2842
rect 1690 2816 1720 2842
rect 1762 2816 1792 2842
rect 1858 2816 1888 2842
rect 1966 2816 1996 2842
rect 2084 2816 2114 2842
rect 2168 2816 2198 2842
rect 2312 2816 2342 2842
rect 2449 2816 2479 2842
rect 2533 2816 2563 2842
rect 2641 2816 2671 2842
rect 2747 2816 2777 2842
rect 2867 2816 2897 2842
rect 2951 2816 2981 2842
rect 3044 2816 3074 2842
rect 1207 2656 1237 2672
rect 1207 2626 1263 2656
rect 1112 2584 1142 2616
rect 1112 2568 1171 2584
rect 1112 2534 1127 2568
rect 1161 2534 1171 2568
rect 1112 2518 1171 2534
rect 1233 2578 1263 2626
rect 1492 2748 1522 2774
rect 1395 2584 1425 2616
rect 1492 2588 1522 2620
rect 1690 2616 1720 2648
rect 1624 2600 1720 2616
rect 1395 2578 1447 2584
rect 1233 2568 1447 2578
rect 1233 2534 1403 2568
rect 1437 2534 1447 2568
rect 1233 2524 1447 2534
rect 1112 2496 1142 2518
rect 1233 2495 1263 2524
rect 1395 2518 1447 2524
rect 1489 2572 1553 2588
rect 1489 2538 1503 2572
rect 1537 2538 1553 2572
rect 1624 2566 1634 2600
rect 1668 2586 1720 2600
rect 1762 2600 1792 2648
rect 1668 2566 1708 2586
rect 1624 2550 1708 2566
rect 1489 2522 1553 2538
rect 1395 2496 1425 2518
rect 1207 2465 1263 2495
rect 1207 2450 1237 2465
rect 1490 2450 1520 2522
rect 1678 2494 1708 2550
rect 1762 2584 1816 2600
rect 1762 2550 1772 2584
rect 1806 2550 1816 2584
rect 1762 2534 1816 2550
rect 1858 2548 1888 2732
rect 1966 2700 1996 2732
rect 1930 2684 1996 2700
rect 2084 2694 2114 2732
rect 2168 2700 2198 2732
rect 1930 2650 1940 2684
rect 1974 2650 1996 2684
rect 1930 2634 1996 2650
rect 2060 2684 2126 2694
rect 2060 2650 2076 2684
rect 2110 2650 2126 2684
rect 2060 2640 2126 2650
rect 2168 2684 2222 2700
rect 2168 2650 2178 2684
rect 2212 2650 2222 2684
rect 1762 2494 1792 2534
rect 1858 2532 1924 2548
rect 1858 2498 1880 2532
rect 1914 2498 1924 2532
rect 1858 2482 1924 2498
rect 1880 2450 1910 2482
rect 1966 2450 1996 2634
rect 2168 2634 2222 2650
rect 3232 2810 3262 2836
rect 3316 2810 3346 2836
rect 3504 2816 3534 2842
rect 2168 2598 2198 2634
rect 2061 2568 2198 2598
rect 2312 2582 2342 2648
rect 2449 2616 2479 2648
rect 2533 2616 2563 2648
rect 2061 2438 2091 2568
rect 2265 2566 2342 2582
rect 2265 2532 2275 2566
rect 2309 2552 2342 2566
rect 2393 2600 2483 2616
rect 2393 2566 2403 2600
rect 2437 2566 2483 2600
rect 2309 2532 2319 2552
rect 2393 2550 2483 2566
rect 2533 2600 2599 2616
rect 2533 2566 2555 2600
rect 2589 2566 2599 2600
rect 2533 2550 2599 2566
rect 2133 2510 2200 2526
rect 2133 2476 2143 2510
rect 2177 2476 2200 2510
rect 2265 2516 2319 2532
rect 2265 2494 2295 2516
rect 2453 2494 2483 2550
rect 2537 2494 2567 2550
rect 2641 2548 2671 2732
rect 2747 2700 2777 2732
rect 2713 2684 2777 2700
rect 2867 2694 2897 2732
rect 2713 2650 2723 2684
rect 2757 2650 2777 2684
rect 2713 2634 2777 2650
rect 2843 2684 2909 2694
rect 2843 2650 2859 2684
rect 2893 2650 2909 2684
rect 2843 2640 2909 2650
rect 2641 2532 2701 2548
rect 2641 2512 2657 2532
rect 2637 2498 2657 2512
rect 2691 2498 2701 2532
rect 2133 2460 2200 2476
rect 2170 2438 2200 2460
rect 2637 2482 2701 2498
rect 2637 2450 2667 2482
rect 2747 2450 2777 2634
rect 2951 2598 2981 2732
rect 2843 2568 2981 2598
rect 3044 2586 3074 2732
rect 3232 2593 3262 2682
rect 3316 2667 3346 2682
rect 3316 2637 3379 2667
rect 3349 2599 3379 2637
rect 3599 2800 3629 2826
rect 3787 2816 3817 2842
rect 4082 2816 4112 2842
rect 4154 2816 4184 2842
rect 4250 2816 4280 2842
rect 4358 2816 4388 2842
rect 4476 2816 4506 2842
rect 4560 2816 4590 2842
rect 4704 2816 4734 2842
rect 4841 2816 4871 2842
rect 4925 2816 4955 2842
rect 5033 2816 5063 2842
rect 5139 2816 5169 2842
rect 5259 2816 5289 2842
rect 5343 2816 5373 2842
rect 5436 2816 5466 2842
rect 3599 2656 3629 2672
rect 3599 2626 3655 2656
rect 3031 2570 3085 2586
rect 2843 2538 2873 2568
rect 2819 2522 2873 2538
rect 3031 2536 3041 2570
rect 3075 2536 3085 2570
rect 2819 2488 2829 2522
rect 2863 2488 2873 2522
rect 2819 2472 2873 2488
rect 2843 2438 2873 2472
rect 2915 2510 2979 2526
rect 3031 2520 3085 2536
rect 3232 2583 3307 2593
rect 3232 2549 3257 2583
rect 3291 2549 3307 2583
rect 3232 2539 3307 2549
rect 3349 2583 3404 2599
rect 3349 2549 3359 2583
rect 3393 2549 3404 2583
rect 2915 2476 2925 2510
rect 2959 2476 2979 2510
rect 2915 2460 2979 2476
rect 2949 2438 2979 2460
rect 3044 2450 3074 2520
rect 3232 2450 3262 2539
rect 3349 2533 3404 2549
rect 3504 2584 3534 2616
rect 3504 2568 3563 2584
rect 3504 2534 3519 2568
rect 3553 2534 3563 2568
rect 3349 2495 3379 2533
rect 3504 2518 3563 2534
rect 3625 2578 3655 2626
rect 3884 2748 3914 2774
rect 3787 2584 3817 2616
rect 3884 2588 3914 2620
rect 4082 2616 4112 2648
rect 4016 2600 4112 2616
rect 3787 2578 3839 2584
rect 3625 2568 3839 2578
rect 3625 2534 3795 2568
rect 3829 2534 3839 2568
rect 3625 2524 3839 2534
rect 3504 2496 3534 2518
rect 3316 2465 3379 2495
rect 3316 2450 3346 2465
rect 3625 2495 3655 2524
rect 3787 2518 3839 2524
rect 3881 2572 3945 2588
rect 3881 2538 3895 2572
rect 3929 2538 3945 2572
rect 4016 2566 4026 2600
rect 4060 2586 4112 2600
rect 4154 2600 4184 2648
rect 4060 2566 4100 2586
rect 4016 2550 4100 2566
rect 3881 2522 3945 2538
rect 3787 2496 3817 2518
rect 3599 2465 3655 2495
rect 3599 2450 3629 2465
rect 3882 2450 3912 2522
rect 4070 2494 4100 2550
rect 4154 2584 4208 2600
rect 4154 2550 4164 2584
rect 4198 2550 4208 2584
rect 4154 2534 4208 2550
rect 4250 2548 4280 2732
rect 4358 2700 4388 2732
rect 4322 2684 4388 2700
rect 4476 2694 4506 2732
rect 4560 2700 4590 2732
rect 4322 2650 4332 2684
rect 4366 2650 4388 2684
rect 4322 2634 4388 2650
rect 4452 2684 4518 2694
rect 4452 2650 4468 2684
rect 4502 2650 4518 2684
rect 4452 2640 4518 2650
rect 4560 2684 4614 2700
rect 4560 2650 4570 2684
rect 4604 2650 4614 2684
rect 4154 2494 4184 2534
rect 4250 2532 4316 2548
rect 4250 2498 4272 2532
rect 4306 2498 4316 2532
rect 4250 2482 4316 2498
rect 4272 2450 4302 2482
rect 4358 2450 4388 2634
rect 4560 2634 4614 2650
rect 5624 2810 5654 2836
rect 5708 2810 5738 2836
rect 5896 2816 5926 2842
rect 4560 2598 4590 2634
rect 4453 2568 4590 2598
rect 4704 2582 4734 2648
rect 4841 2616 4871 2648
rect 4925 2616 4955 2648
rect 4453 2438 4483 2568
rect 4657 2566 4734 2582
rect 4657 2532 4667 2566
rect 4701 2552 4734 2566
rect 4785 2600 4875 2616
rect 4785 2566 4795 2600
rect 4829 2566 4875 2600
rect 4701 2532 4711 2552
rect 4785 2550 4875 2566
rect 4925 2600 4991 2616
rect 4925 2566 4947 2600
rect 4981 2566 4991 2600
rect 4925 2550 4991 2566
rect 4525 2510 4592 2526
rect 4525 2476 4535 2510
rect 4569 2476 4592 2510
rect 4657 2516 4711 2532
rect 4657 2494 4687 2516
rect 4845 2494 4875 2550
rect 4929 2494 4959 2550
rect 5033 2548 5063 2732
rect 5139 2700 5169 2732
rect 5105 2684 5169 2700
rect 5259 2694 5289 2732
rect 5105 2650 5115 2684
rect 5149 2650 5169 2684
rect 5105 2634 5169 2650
rect 5235 2684 5301 2694
rect 5235 2650 5251 2684
rect 5285 2650 5301 2684
rect 5235 2640 5301 2650
rect 5033 2532 5093 2548
rect 5033 2512 5049 2532
rect 5029 2498 5049 2512
rect 5083 2498 5093 2532
rect 4525 2460 4592 2476
rect 4562 2438 4592 2460
rect 5029 2482 5093 2498
rect 5029 2450 5059 2482
rect 5139 2450 5169 2634
rect 5343 2598 5373 2732
rect 5235 2568 5373 2598
rect 5436 2586 5466 2732
rect 5624 2593 5654 2682
rect 5708 2667 5738 2682
rect 5708 2637 5771 2667
rect 5741 2599 5771 2637
rect 5991 2800 6021 2826
rect 6179 2816 6209 2842
rect 6474 2816 6504 2842
rect 6546 2816 6576 2842
rect 6642 2816 6672 2842
rect 6750 2816 6780 2842
rect 6868 2816 6898 2842
rect 6952 2816 6982 2842
rect 7096 2816 7126 2842
rect 7233 2816 7263 2842
rect 7317 2816 7347 2842
rect 7425 2816 7455 2842
rect 7531 2816 7561 2842
rect 7651 2816 7681 2842
rect 7735 2816 7765 2842
rect 7828 2816 7858 2842
rect 5991 2656 6021 2672
rect 5991 2626 6047 2656
rect 5423 2570 5477 2586
rect 5235 2538 5265 2568
rect 5211 2522 5265 2538
rect 5423 2536 5433 2570
rect 5467 2536 5477 2570
rect 5211 2488 5221 2522
rect 5255 2488 5265 2522
rect 5211 2472 5265 2488
rect 5235 2438 5265 2472
rect 5307 2510 5371 2526
rect 5423 2520 5477 2536
rect 5624 2583 5699 2593
rect 5624 2549 5649 2583
rect 5683 2549 5699 2583
rect 5624 2539 5699 2549
rect 5741 2583 5796 2599
rect 5741 2549 5751 2583
rect 5785 2549 5796 2583
rect 5307 2476 5317 2510
rect 5351 2476 5371 2510
rect 5307 2460 5371 2476
rect 5341 2438 5371 2460
rect 5436 2450 5466 2520
rect 5624 2450 5654 2539
rect 5741 2533 5796 2549
rect 5896 2584 5926 2616
rect 5896 2568 5955 2584
rect 5896 2534 5911 2568
rect 5945 2534 5955 2568
rect 5741 2495 5771 2533
rect 5896 2518 5955 2534
rect 6017 2578 6047 2626
rect 6276 2748 6306 2774
rect 6179 2584 6209 2616
rect 6276 2588 6306 2620
rect 6474 2616 6504 2648
rect 6408 2600 6504 2616
rect 6179 2578 6231 2584
rect 6017 2568 6231 2578
rect 6017 2534 6187 2568
rect 6221 2534 6231 2568
rect 6017 2524 6231 2534
rect 5896 2496 5926 2518
rect 5708 2465 5771 2495
rect 5708 2450 5738 2465
rect 6017 2495 6047 2524
rect 6179 2518 6231 2524
rect 6273 2572 6337 2588
rect 6273 2538 6287 2572
rect 6321 2538 6337 2572
rect 6408 2566 6418 2600
rect 6452 2586 6504 2600
rect 6546 2600 6576 2648
rect 6452 2566 6492 2586
rect 6408 2550 6492 2566
rect 6273 2522 6337 2538
rect 6179 2496 6209 2518
rect 5991 2465 6047 2495
rect 5991 2450 6021 2465
rect 6274 2450 6304 2522
rect 6462 2494 6492 2550
rect 6546 2584 6600 2600
rect 6546 2550 6556 2584
rect 6590 2550 6600 2584
rect 6546 2534 6600 2550
rect 6642 2548 6672 2732
rect 6750 2700 6780 2732
rect 6714 2684 6780 2700
rect 6868 2694 6898 2732
rect 6952 2700 6982 2732
rect 6714 2650 6724 2684
rect 6758 2650 6780 2684
rect 6714 2634 6780 2650
rect 6844 2684 6910 2694
rect 6844 2650 6860 2684
rect 6894 2650 6910 2684
rect 6844 2640 6910 2650
rect 6952 2684 7006 2700
rect 6952 2650 6962 2684
rect 6996 2650 7006 2684
rect 6546 2494 6576 2534
rect 6642 2532 6708 2548
rect 6642 2498 6664 2532
rect 6698 2498 6708 2532
rect 6642 2482 6708 2498
rect 6664 2450 6694 2482
rect 6750 2450 6780 2634
rect 6952 2634 7006 2650
rect 8016 2810 8046 2836
rect 8100 2810 8130 2836
rect 8288 2816 8318 2842
rect 6952 2598 6982 2634
rect 6845 2568 6982 2598
rect 7096 2582 7126 2648
rect 7233 2616 7263 2648
rect 7317 2616 7347 2648
rect 6845 2438 6875 2568
rect 7049 2566 7126 2582
rect 7049 2532 7059 2566
rect 7093 2552 7126 2566
rect 7177 2600 7267 2616
rect 7177 2566 7187 2600
rect 7221 2566 7267 2600
rect 7093 2532 7103 2552
rect 7177 2550 7267 2566
rect 7317 2600 7383 2616
rect 7317 2566 7339 2600
rect 7373 2566 7383 2600
rect 7317 2550 7383 2566
rect 6917 2510 6984 2526
rect 6917 2476 6927 2510
rect 6961 2476 6984 2510
rect 7049 2516 7103 2532
rect 7049 2494 7079 2516
rect 7237 2494 7267 2550
rect 7321 2494 7351 2550
rect 7425 2548 7455 2732
rect 7531 2700 7561 2732
rect 7497 2684 7561 2700
rect 7651 2694 7681 2732
rect 7497 2650 7507 2684
rect 7541 2650 7561 2684
rect 7497 2634 7561 2650
rect 7627 2684 7693 2694
rect 7627 2650 7643 2684
rect 7677 2650 7693 2684
rect 7627 2640 7693 2650
rect 7425 2532 7485 2548
rect 7425 2512 7441 2532
rect 7421 2498 7441 2512
rect 7475 2498 7485 2532
rect 6917 2460 6984 2476
rect 6954 2438 6984 2460
rect 7421 2482 7485 2498
rect 7421 2450 7451 2482
rect 7531 2450 7561 2634
rect 7735 2598 7765 2732
rect 7627 2568 7765 2598
rect 7828 2586 7858 2732
rect 8016 2593 8046 2682
rect 8100 2667 8130 2682
rect 8100 2637 8163 2667
rect 8133 2599 8163 2637
rect 8383 2800 8413 2826
rect 8571 2816 8601 2842
rect 8866 2816 8896 2842
rect 8938 2816 8968 2842
rect 9034 2816 9064 2842
rect 9142 2816 9172 2842
rect 9260 2816 9290 2842
rect 9344 2816 9374 2842
rect 9488 2816 9518 2842
rect 9625 2816 9655 2842
rect 9709 2816 9739 2842
rect 9817 2816 9847 2842
rect 9923 2816 9953 2842
rect 10043 2816 10073 2842
rect 10127 2816 10157 2842
rect 10220 2816 10250 2842
rect 8383 2656 8413 2672
rect 8383 2626 8439 2656
rect 7815 2570 7869 2586
rect 7627 2538 7657 2568
rect 7603 2522 7657 2538
rect 7815 2536 7825 2570
rect 7859 2536 7869 2570
rect 7603 2488 7613 2522
rect 7647 2488 7657 2522
rect 7603 2472 7657 2488
rect 7627 2438 7657 2472
rect 7699 2510 7763 2526
rect 7815 2520 7869 2536
rect 8016 2583 8091 2593
rect 8016 2549 8041 2583
rect 8075 2549 8091 2583
rect 8016 2539 8091 2549
rect 8133 2583 8188 2599
rect 8133 2549 8143 2583
rect 8177 2549 8188 2583
rect 7699 2476 7709 2510
rect 7743 2476 7763 2510
rect 7699 2460 7763 2476
rect 7733 2438 7763 2460
rect 7828 2450 7858 2520
rect 8016 2450 8046 2539
rect 8133 2533 8188 2549
rect 8288 2584 8318 2616
rect 8288 2568 8347 2584
rect 8288 2534 8303 2568
rect 8337 2534 8347 2568
rect 8133 2495 8163 2533
rect 8288 2518 8347 2534
rect 8409 2578 8439 2626
rect 8668 2748 8698 2774
rect 8571 2584 8601 2616
rect 8668 2588 8698 2620
rect 8866 2616 8896 2648
rect 8800 2600 8896 2616
rect 8571 2578 8623 2584
rect 8409 2568 8623 2578
rect 8409 2534 8579 2568
rect 8613 2534 8623 2568
rect 8409 2524 8623 2534
rect 8288 2496 8318 2518
rect 8100 2465 8163 2495
rect 8100 2450 8130 2465
rect 8409 2495 8439 2524
rect 8571 2518 8623 2524
rect 8665 2572 8729 2588
rect 8665 2538 8679 2572
rect 8713 2538 8729 2572
rect 8800 2566 8810 2600
rect 8844 2586 8896 2600
rect 8938 2600 8968 2648
rect 8844 2566 8884 2586
rect 8800 2550 8884 2566
rect 8665 2522 8729 2538
rect 8571 2496 8601 2518
rect 8383 2465 8439 2495
rect 8383 2450 8413 2465
rect 8666 2450 8696 2522
rect 8854 2494 8884 2550
rect 8938 2584 8992 2600
rect 8938 2550 8948 2584
rect 8982 2550 8992 2584
rect 8938 2534 8992 2550
rect 9034 2548 9064 2732
rect 9142 2700 9172 2732
rect 9106 2684 9172 2700
rect 9260 2694 9290 2732
rect 9344 2700 9374 2732
rect 9106 2650 9116 2684
rect 9150 2650 9172 2684
rect 9106 2634 9172 2650
rect 9236 2684 9302 2694
rect 9236 2650 9252 2684
rect 9286 2650 9302 2684
rect 9236 2640 9302 2650
rect 9344 2684 9398 2700
rect 9344 2650 9354 2684
rect 9388 2650 9398 2684
rect 8938 2494 8968 2534
rect 9034 2532 9100 2548
rect 9034 2498 9056 2532
rect 9090 2498 9100 2532
rect 9034 2482 9100 2498
rect 9056 2450 9086 2482
rect 9142 2450 9172 2634
rect 9344 2634 9398 2650
rect 10408 2810 10438 2836
rect 10492 2810 10522 2836
rect 10680 2816 10710 2842
rect 9344 2598 9374 2634
rect 9237 2568 9374 2598
rect 9488 2582 9518 2648
rect 9625 2616 9655 2648
rect 9709 2616 9739 2648
rect 9237 2438 9267 2568
rect 9441 2566 9518 2582
rect 9441 2532 9451 2566
rect 9485 2552 9518 2566
rect 9569 2600 9659 2616
rect 9569 2566 9579 2600
rect 9613 2566 9659 2600
rect 9485 2532 9495 2552
rect 9569 2550 9659 2566
rect 9709 2600 9775 2616
rect 9709 2566 9731 2600
rect 9765 2566 9775 2600
rect 9709 2550 9775 2566
rect 9309 2510 9376 2526
rect 9309 2476 9319 2510
rect 9353 2476 9376 2510
rect 9441 2516 9495 2532
rect 9441 2494 9471 2516
rect 9629 2494 9659 2550
rect 9713 2494 9743 2550
rect 9817 2548 9847 2732
rect 9923 2700 9953 2732
rect 9889 2684 9953 2700
rect 10043 2694 10073 2732
rect 9889 2650 9899 2684
rect 9933 2650 9953 2684
rect 9889 2634 9953 2650
rect 10019 2684 10085 2694
rect 10019 2650 10035 2684
rect 10069 2650 10085 2684
rect 10019 2640 10085 2650
rect 9817 2532 9877 2548
rect 9817 2512 9833 2532
rect 9813 2498 9833 2512
rect 9867 2498 9877 2532
rect 9309 2460 9376 2476
rect 9346 2438 9376 2460
rect 9813 2482 9877 2498
rect 9813 2450 9843 2482
rect 9923 2450 9953 2634
rect 10127 2598 10157 2732
rect 10019 2568 10157 2598
rect 10220 2586 10250 2732
rect 10408 2593 10438 2682
rect 10492 2667 10522 2682
rect 10492 2637 10555 2667
rect 10525 2599 10555 2637
rect 10775 2800 10805 2826
rect 10963 2816 10993 2842
rect 11258 2816 11288 2842
rect 11330 2816 11360 2842
rect 11426 2816 11456 2842
rect 11534 2816 11564 2842
rect 11652 2816 11682 2842
rect 11736 2816 11766 2842
rect 11880 2816 11910 2842
rect 12017 2816 12047 2842
rect 12101 2816 12131 2842
rect 12209 2816 12239 2842
rect 12315 2816 12345 2842
rect 12435 2816 12465 2842
rect 12519 2816 12549 2842
rect 12612 2816 12642 2842
rect 10775 2656 10805 2672
rect 10775 2626 10831 2656
rect 10207 2570 10261 2586
rect 10019 2538 10049 2568
rect 9995 2522 10049 2538
rect 10207 2536 10217 2570
rect 10251 2536 10261 2570
rect 9995 2488 10005 2522
rect 10039 2488 10049 2522
rect 9995 2472 10049 2488
rect 10019 2438 10049 2472
rect 10091 2510 10155 2526
rect 10207 2520 10261 2536
rect 10408 2583 10483 2593
rect 10408 2549 10433 2583
rect 10467 2549 10483 2583
rect 10408 2539 10483 2549
rect 10525 2583 10580 2599
rect 10525 2549 10535 2583
rect 10569 2549 10580 2583
rect 10091 2476 10101 2510
rect 10135 2476 10155 2510
rect 10091 2460 10155 2476
rect 10125 2438 10155 2460
rect 10220 2450 10250 2520
rect 10408 2450 10438 2539
rect 10525 2533 10580 2549
rect 10680 2584 10710 2616
rect 10680 2568 10739 2584
rect 10680 2534 10695 2568
rect 10729 2534 10739 2568
rect 10525 2495 10555 2533
rect 10680 2518 10739 2534
rect 10801 2578 10831 2626
rect 11060 2748 11090 2774
rect 10963 2584 10993 2616
rect 11060 2588 11090 2620
rect 11258 2616 11288 2648
rect 11192 2600 11288 2616
rect 10963 2578 11015 2584
rect 10801 2568 11015 2578
rect 10801 2534 10971 2568
rect 11005 2534 11015 2568
rect 10801 2524 11015 2534
rect 10680 2496 10710 2518
rect 10492 2465 10555 2495
rect 10492 2450 10522 2465
rect 10801 2495 10831 2524
rect 10963 2518 11015 2524
rect 11057 2572 11121 2588
rect 11057 2538 11071 2572
rect 11105 2538 11121 2572
rect 11192 2566 11202 2600
rect 11236 2586 11288 2600
rect 11330 2600 11360 2648
rect 11236 2566 11276 2586
rect 11192 2550 11276 2566
rect 11057 2522 11121 2538
rect 10963 2496 10993 2518
rect 10775 2465 10831 2495
rect 10775 2450 10805 2465
rect 11058 2450 11088 2522
rect 11246 2494 11276 2550
rect 11330 2584 11384 2600
rect 11330 2550 11340 2584
rect 11374 2550 11384 2584
rect 11330 2534 11384 2550
rect 11426 2548 11456 2732
rect 11534 2700 11564 2732
rect 11498 2684 11564 2700
rect 11652 2694 11682 2732
rect 11736 2700 11766 2732
rect 11498 2650 11508 2684
rect 11542 2650 11564 2684
rect 11498 2634 11564 2650
rect 11628 2684 11694 2694
rect 11628 2650 11644 2684
rect 11678 2650 11694 2684
rect 11628 2640 11694 2650
rect 11736 2684 11790 2700
rect 11736 2650 11746 2684
rect 11780 2650 11790 2684
rect 11330 2494 11360 2534
rect 11426 2532 11492 2548
rect 11426 2498 11448 2532
rect 11482 2498 11492 2532
rect 11426 2482 11492 2498
rect 11448 2450 11478 2482
rect 11534 2450 11564 2634
rect 11736 2634 11790 2650
rect 12800 2810 12830 2836
rect 12884 2810 12914 2836
rect 11736 2598 11766 2634
rect 11629 2568 11766 2598
rect 11880 2582 11910 2648
rect 12017 2616 12047 2648
rect 12101 2616 12131 2648
rect 11629 2438 11659 2568
rect 11833 2566 11910 2582
rect 11833 2532 11843 2566
rect 11877 2552 11910 2566
rect 11961 2600 12051 2616
rect 11961 2566 11971 2600
rect 12005 2566 12051 2600
rect 11877 2532 11887 2552
rect 11961 2550 12051 2566
rect 12101 2600 12167 2616
rect 12101 2566 12123 2600
rect 12157 2566 12167 2600
rect 12101 2550 12167 2566
rect 11701 2510 11768 2526
rect 11701 2476 11711 2510
rect 11745 2476 11768 2510
rect 11833 2516 11887 2532
rect 11833 2494 11863 2516
rect 12021 2494 12051 2550
rect 12105 2494 12135 2550
rect 12209 2548 12239 2732
rect 12315 2700 12345 2732
rect 12281 2684 12345 2700
rect 12435 2694 12465 2732
rect 12281 2650 12291 2684
rect 12325 2650 12345 2684
rect 12281 2634 12345 2650
rect 12411 2684 12477 2694
rect 12411 2650 12427 2684
rect 12461 2650 12477 2684
rect 12411 2640 12477 2650
rect 12209 2532 12269 2548
rect 12209 2512 12225 2532
rect 12205 2498 12225 2512
rect 12259 2498 12269 2532
rect 11701 2460 11768 2476
rect 11738 2438 11768 2460
rect 12205 2482 12269 2498
rect 12205 2450 12235 2482
rect 12315 2450 12345 2634
rect 12519 2598 12549 2732
rect 12411 2568 12549 2598
rect 12612 2586 12642 2732
rect 12800 2593 12830 2682
rect 12884 2667 12914 2682
rect 12884 2637 12947 2667
rect 12917 2599 12947 2637
rect 12599 2570 12653 2586
rect 12411 2538 12441 2568
rect 12387 2522 12441 2538
rect 12599 2536 12609 2570
rect 12643 2536 12653 2570
rect 12387 2488 12397 2522
rect 12431 2488 12441 2522
rect 12387 2472 12441 2488
rect 12411 2438 12441 2472
rect 12483 2510 12547 2526
rect 12599 2520 12653 2536
rect 12800 2583 12875 2593
rect 12800 2549 12825 2583
rect 12859 2549 12875 2583
rect 12800 2539 12875 2549
rect 12917 2583 12972 2599
rect 12917 2549 12927 2583
rect 12961 2549 12972 2583
rect 12483 2476 12493 2510
rect 12527 2476 12547 2510
rect 12483 2460 12547 2476
rect 12517 2438 12547 2460
rect 12612 2450 12642 2520
rect 12800 2450 12830 2539
rect 12917 2533 12972 2549
rect 12917 2495 12947 2533
rect 12884 2465 12947 2495
rect 12884 2450 12914 2465
rect 1112 2340 1142 2366
rect 1207 2340 1237 2366
rect 1395 2340 1425 2366
rect 1490 2340 1520 2366
rect 1678 2340 1708 2366
rect 1762 2340 1792 2366
rect 1880 2340 1910 2366
rect 1966 2340 1996 2366
rect 2061 2340 2091 2366
rect 2170 2340 2200 2366
rect 2265 2340 2295 2366
rect 2453 2340 2483 2366
rect 2537 2340 2567 2366
rect 2637 2340 2667 2366
rect 2747 2340 2777 2366
rect 2843 2340 2873 2366
rect 2949 2340 2979 2366
rect 3044 2340 3074 2366
rect 3232 2340 3262 2366
rect 3316 2340 3346 2366
rect 3504 2340 3534 2366
rect 3599 2340 3629 2366
rect 3787 2340 3817 2366
rect 3882 2340 3912 2366
rect 4070 2340 4100 2366
rect 4154 2340 4184 2366
rect 4272 2340 4302 2366
rect 4358 2340 4388 2366
rect 4453 2340 4483 2366
rect 4562 2340 4592 2366
rect 4657 2340 4687 2366
rect 4845 2340 4875 2366
rect 4929 2340 4959 2366
rect 5029 2340 5059 2366
rect 5139 2340 5169 2366
rect 5235 2340 5265 2366
rect 5341 2340 5371 2366
rect 5436 2340 5466 2366
rect 5624 2340 5654 2366
rect 5708 2340 5738 2366
rect 5896 2340 5926 2366
rect 5991 2340 6021 2366
rect 6179 2340 6209 2366
rect 6274 2340 6304 2366
rect 6462 2340 6492 2366
rect 6546 2340 6576 2366
rect 6664 2340 6694 2366
rect 6750 2340 6780 2366
rect 6845 2340 6875 2366
rect 6954 2340 6984 2366
rect 7049 2340 7079 2366
rect 7237 2340 7267 2366
rect 7321 2340 7351 2366
rect 7421 2340 7451 2366
rect 7531 2340 7561 2366
rect 7627 2340 7657 2366
rect 7733 2340 7763 2366
rect 7828 2340 7858 2366
rect 8016 2340 8046 2366
rect 8100 2340 8130 2366
rect 8288 2340 8318 2366
rect 8383 2340 8413 2366
rect 8571 2340 8601 2366
rect 8666 2340 8696 2366
rect 8854 2340 8884 2366
rect 8938 2340 8968 2366
rect 9056 2340 9086 2366
rect 9142 2340 9172 2366
rect 9237 2340 9267 2366
rect 9346 2340 9376 2366
rect 9441 2340 9471 2366
rect 9629 2340 9659 2366
rect 9713 2340 9743 2366
rect 9813 2340 9843 2366
rect 9923 2340 9953 2366
rect 10019 2340 10049 2366
rect 10125 2340 10155 2366
rect 10220 2340 10250 2366
rect 10408 2340 10438 2366
rect 10492 2340 10522 2366
rect 10680 2340 10710 2366
rect 10775 2340 10805 2366
rect 10963 2340 10993 2366
rect 11058 2340 11088 2366
rect 11246 2340 11276 2366
rect 11330 2340 11360 2366
rect 11448 2340 11478 2366
rect 11534 2340 11564 2366
rect 11629 2340 11659 2366
rect 11738 2340 11768 2366
rect 11833 2340 11863 2366
rect 12021 2340 12051 2366
rect 12105 2340 12135 2366
rect 12205 2340 12235 2366
rect 12315 2340 12345 2366
rect 12411 2340 12441 2366
rect 12517 2340 12547 2366
rect 12612 2340 12642 2366
rect 12800 2340 12830 2366
rect 12884 2340 12914 2366
<< polycont >>
rect 1072 5842 1106 5876
rect 1190 5855 1224 5889
rect 1355 5842 1389 5876
rect 1489 5842 1523 5876
rect 2943 5958 2977 5992
rect 2841 5892 2875 5926
rect 2649 5842 2683 5876
rect 2745 5842 2779 5876
rect 2877 5784 2911 5818
rect 3111 5856 3145 5890
rect 3438 5855 3472 5889
rect 3754 5958 3788 5992
rect 3856 5900 3890 5934
rect 3540 5796 3574 5830
rect 3636 5796 3670 5830
rect 3819 5784 3853 5818
rect 3933 5796 3967 5830
rect 4069 5842 4103 5876
rect 2934 5296 2968 5330
rect 4177 5299 4211 5333
rect 6569 5301 6603 5335
rect 8961 5301 8995 5335
rect 11353 5302 11387 5336
rect 1066 4984 1100 5018
rect 1566 5085 1600 5119
rect 1702 5085 1736 5119
rect 1168 4984 1202 5018
rect 1384 4971 1418 5005
rect 1500 4911 1534 4945
rect 1596 4923 1630 4957
rect 2247 5085 2281 5119
rect 1870 5001 1904 5035
rect 2022 5001 2056 5035
rect 2349 5085 2383 5119
rect 2485 5085 2519 5119
rect 1768 4933 1802 4967
rect 2150 4967 2184 5001
rect 2282 4911 2316 4945
rect 2653 4985 2687 5019
rect 2545 4933 2579 4967
rect 2791 5001 2825 5035
rect 2922 4973 2956 5007
rect 3022 4969 3056 5003
rect 3298 4969 3332 5003
rect 3458 4984 3492 5018
rect 3958 5085 3992 5119
rect 4094 5085 4128 5119
rect 3560 4984 3594 5018
rect 3776 4971 3810 5005
rect 3892 4911 3926 4945
rect 3988 4923 4022 4957
rect 4639 5085 4673 5119
rect 4262 5001 4296 5035
rect 4414 5001 4448 5035
rect 4741 5085 4775 5119
rect 4877 5085 4911 5119
rect 4160 4933 4194 4967
rect 4542 4967 4576 5001
rect 4674 4911 4708 4945
rect 5045 4985 5079 5019
rect 4937 4933 4971 4967
rect 5183 5001 5217 5035
rect 5314 4973 5348 5007
rect 5414 4969 5448 5003
rect 5690 4969 5724 5003
rect 5850 4984 5884 5018
rect 6350 5085 6384 5119
rect 6486 5085 6520 5119
rect 5952 4984 5986 5018
rect 6168 4971 6202 5005
rect 6284 4911 6318 4945
rect 6380 4923 6414 4957
rect 7031 5085 7065 5119
rect 6654 5001 6688 5035
rect 6806 5001 6840 5035
rect 7133 5085 7167 5119
rect 7269 5085 7303 5119
rect 6552 4933 6586 4967
rect 6934 4967 6968 5001
rect 7066 4911 7100 4945
rect 7437 4985 7471 5019
rect 7329 4933 7363 4967
rect 7575 5001 7609 5035
rect 7706 4973 7740 5007
rect 7806 4969 7840 5003
rect 8082 4969 8116 5003
rect 8242 4984 8276 5018
rect 8742 5085 8776 5119
rect 8878 5085 8912 5119
rect 8344 4984 8378 5018
rect 8560 4971 8594 5005
rect 8676 4911 8710 4945
rect 8772 4923 8806 4957
rect 9423 5085 9457 5119
rect 9046 5001 9080 5035
rect 9198 5001 9232 5035
rect 9525 5085 9559 5119
rect 9661 5085 9695 5119
rect 8944 4933 8978 4967
rect 9326 4967 9360 5001
rect 9458 4911 9492 4945
rect 9829 4985 9863 5019
rect 9721 4933 9755 4967
rect 9967 5001 10001 5035
rect 10098 4973 10132 5007
rect 10198 4969 10232 5003
rect 10474 4969 10508 5003
rect 10634 4984 10668 5018
rect 11134 5085 11168 5119
rect 11270 5085 11304 5119
rect 10736 4984 10770 5018
rect 10952 4971 10986 5005
rect 11068 4911 11102 4945
rect 11164 4923 11198 4957
rect 11815 5085 11849 5119
rect 11438 5001 11472 5035
rect 11590 5001 11624 5035
rect 11917 5085 11951 5119
rect 12053 5085 12087 5119
rect 11336 4933 11370 4967
rect 11718 4967 11752 5001
rect 11850 4911 11884 4945
rect 12221 4985 12255 5019
rect 12113 4933 12147 4967
rect 12359 5001 12393 5035
rect 12490 4973 12524 5007
rect 12590 4969 12624 5003
rect 12866 4969 12900 5003
rect 4248 4613 4282 4647
rect 6640 4613 6674 4647
rect 9032 4613 9066 4647
rect 11424 4613 11458 4647
rect 631 4280 665 4314
rect 749 4293 783 4327
rect 914 4280 948 4314
rect 1048 4280 1082 4314
rect 1505 4280 1539 4314
rect 1573 4280 1607 4314
rect 1641 4280 1675 4314
rect 1709 4280 1743 4314
rect 1777 4280 1811 4314
rect 1845 4280 1879 4314
rect 2005 4280 2039 4314
rect 2073 4280 2107 4314
rect 2141 4280 2175 4314
rect 2209 4280 2243 4314
rect 2277 4280 2311 4314
rect 2345 4280 2379 4314
rect 2413 4280 2447 4314
rect 2481 4280 2515 4314
rect 2549 4280 2583 4314
rect 2617 4280 2651 4314
rect 2685 4280 2719 4314
rect 2753 4280 2787 4314
rect 2821 4280 2855 4314
rect 2889 4280 2923 4314
rect 2957 4280 2991 4314
rect 3025 4280 3059 4314
rect 3093 4280 3127 4314
rect 3161 4280 3195 4314
rect 3229 4280 3263 4314
rect 3520 4280 3554 4314
rect 3796 4280 3830 4314
rect 3896 4284 3930 4318
rect 4027 4312 4061 4346
rect 4165 4296 4199 4330
rect 4333 4396 4367 4430
rect 4469 4396 4503 4430
rect 4571 4396 4605 4430
rect 4273 4244 4307 4278
rect 4668 4278 4702 4312
rect 4796 4312 4830 4346
rect 4948 4312 4982 4346
rect 4536 4222 4570 4256
rect 5116 4396 5150 4430
rect 5252 4396 5286 4430
rect 5050 4244 5084 4278
rect 5434 4282 5468 4316
rect 5222 4234 5256 4268
rect 5650 4295 5684 4329
rect 5752 4295 5786 4329
rect 5318 4222 5352 4256
rect 5912 4280 5946 4314
rect 6188 4280 6222 4314
rect 6288 4284 6322 4318
rect 6419 4312 6453 4346
rect 6557 4296 6591 4330
rect 6725 4396 6759 4430
rect 6861 4396 6895 4430
rect 6963 4396 6997 4430
rect 6665 4244 6699 4278
rect 7060 4278 7094 4312
rect 7188 4312 7222 4346
rect 7340 4312 7374 4346
rect 6928 4222 6962 4256
rect 7508 4396 7542 4430
rect 7644 4396 7678 4430
rect 7442 4244 7476 4278
rect 7826 4282 7860 4316
rect 7614 4234 7648 4268
rect 8042 4295 8076 4329
rect 8144 4295 8178 4329
rect 7710 4222 7744 4256
rect 8304 4280 8338 4314
rect 8580 4280 8614 4314
rect 8680 4284 8714 4318
rect 8811 4312 8845 4346
rect 8949 4296 8983 4330
rect 9117 4396 9151 4430
rect 9253 4396 9287 4430
rect 9355 4396 9389 4430
rect 9057 4244 9091 4278
rect 9452 4278 9486 4312
rect 9580 4312 9614 4346
rect 9732 4312 9766 4346
rect 9320 4222 9354 4256
rect 9900 4396 9934 4430
rect 10036 4396 10070 4430
rect 9834 4244 9868 4278
rect 10218 4282 10252 4316
rect 10006 4234 10040 4268
rect 10434 4295 10468 4329
rect 10536 4295 10570 4329
rect 10102 4222 10136 4256
rect 10696 4280 10730 4314
rect 10972 4280 11006 4314
rect 11072 4284 11106 4318
rect 11203 4312 11237 4346
rect 11341 4296 11375 4330
rect 11509 4396 11543 4430
rect 11645 4396 11679 4430
rect 11747 4396 11781 4430
rect 11449 4244 11483 4278
rect 11844 4278 11878 4312
rect 11972 4312 12006 4346
rect 12124 4312 12158 4346
rect 11712 4222 11746 4256
rect 12292 4396 12326 4430
rect 12428 4396 12462 4430
rect 12226 4244 12260 4278
rect 12610 4282 12644 4316
rect 12398 4234 12432 4268
rect 12826 4295 12860 4329
rect 12928 4295 12962 4329
rect 12494 4222 12528 4256
rect 663 3406 697 3440
rect 781 3419 815 3453
rect 946 3406 980 3440
rect 1080 3406 1114 3440
rect 3248 3407 3282 3441
rect 3457 3422 3491 3456
rect 3957 3523 3991 3557
rect 4093 3523 4127 3557
rect 3559 3422 3593 3456
rect 3775 3409 3809 3443
rect 3891 3349 3925 3383
rect 3987 3361 4021 3395
rect 4638 3523 4672 3557
rect 4261 3439 4295 3473
rect 4413 3439 4447 3473
rect 4740 3523 4774 3557
rect 4876 3523 4910 3557
rect 4159 3371 4193 3405
rect 4541 3405 4575 3439
rect 4673 3349 4707 3383
rect 5044 3423 5078 3457
rect 4936 3371 4970 3405
rect 5182 3439 5216 3473
rect 5313 3411 5347 3445
rect 5413 3407 5447 3441
rect 5689 3407 5723 3441
rect 5849 3422 5883 3456
rect 6349 3523 6383 3557
rect 6485 3523 6519 3557
rect 5951 3422 5985 3456
rect 6167 3409 6201 3443
rect 6283 3349 6317 3383
rect 6379 3361 6413 3395
rect 7030 3523 7064 3557
rect 6653 3439 6687 3473
rect 6805 3439 6839 3473
rect 7132 3523 7166 3557
rect 7268 3523 7302 3557
rect 6551 3371 6585 3405
rect 6933 3405 6967 3439
rect 7065 3349 7099 3383
rect 7436 3423 7470 3457
rect 7328 3371 7362 3405
rect 7574 3439 7608 3473
rect 7705 3411 7739 3445
rect 7805 3407 7839 3441
rect 8081 3407 8115 3441
rect 8241 3422 8275 3456
rect 8741 3523 8775 3557
rect 8877 3523 8911 3557
rect 8343 3422 8377 3456
rect 8559 3409 8593 3443
rect 8675 3349 8709 3383
rect 8771 3361 8805 3395
rect 9422 3523 9456 3557
rect 9045 3439 9079 3473
rect 9197 3439 9231 3473
rect 9524 3523 9558 3557
rect 9660 3523 9694 3557
rect 8943 3371 8977 3405
rect 9325 3405 9359 3439
rect 9457 3349 9491 3383
rect 9828 3423 9862 3457
rect 9720 3371 9754 3405
rect 9966 3439 10000 3473
rect 10097 3411 10131 3445
rect 10197 3407 10231 3441
rect 10473 3407 10507 3441
rect 10633 3422 10667 3456
rect 11133 3523 11167 3557
rect 11269 3523 11303 3557
rect 10735 3422 10769 3456
rect 10951 3409 10985 3443
rect 11067 3349 11101 3383
rect 11163 3361 11197 3395
rect 11814 3523 11848 3557
rect 11437 3439 11471 3473
rect 11589 3439 11623 3473
rect 11916 3523 11950 3557
rect 12052 3523 12086 3557
rect 11335 3371 11369 3405
rect 11717 3405 11751 3439
rect 11849 3349 11883 3383
rect 12220 3423 12254 3457
rect 12112 3371 12146 3405
rect 12358 3439 12392 3473
rect 12489 3411 12523 3445
rect 12589 3407 12623 3441
rect 12865 3407 12899 3441
rect 1127 2534 1161 2568
rect 1403 2534 1437 2568
rect 1503 2538 1537 2572
rect 1634 2566 1668 2600
rect 1772 2550 1806 2584
rect 1940 2650 1974 2684
rect 2076 2650 2110 2684
rect 2178 2650 2212 2684
rect 1880 2498 1914 2532
rect 2275 2532 2309 2566
rect 2403 2566 2437 2600
rect 2555 2566 2589 2600
rect 2143 2476 2177 2510
rect 2723 2650 2757 2684
rect 2859 2650 2893 2684
rect 2657 2498 2691 2532
rect 3041 2536 3075 2570
rect 2829 2488 2863 2522
rect 3257 2549 3291 2583
rect 3359 2549 3393 2583
rect 2925 2476 2959 2510
rect 3519 2534 3553 2568
rect 3795 2534 3829 2568
rect 3895 2538 3929 2572
rect 4026 2566 4060 2600
rect 4164 2550 4198 2584
rect 4332 2650 4366 2684
rect 4468 2650 4502 2684
rect 4570 2650 4604 2684
rect 4272 2498 4306 2532
rect 4667 2532 4701 2566
rect 4795 2566 4829 2600
rect 4947 2566 4981 2600
rect 4535 2476 4569 2510
rect 5115 2650 5149 2684
rect 5251 2650 5285 2684
rect 5049 2498 5083 2532
rect 5433 2536 5467 2570
rect 5221 2488 5255 2522
rect 5649 2549 5683 2583
rect 5751 2549 5785 2583
rect 5317 2476 5351 2510
rect 5911 2534 5945 2568
rect 6187 2534 6221 2568
rect 6287 2538 6321 2572
rect 6418 2566 6452 2600
rect 6556 2550 6590 2584
rect 6724 2650 6758 2684
rect 6860 2650 6894 2684
rect 6962 2650 6996 2684
rect 6664 2498 6698 2532
rect 7059 2532 7093 2566
rect 7187 2566 7221 2600
rect 7339 2566 7373 2600
rect 6927 2476 6961 2510
rect 7507 2650 7541 2684
rect 7643 2650 7677 2684
rect 7441 2498 7475 2532
rect 7825 2536 7859 2570
rect 7613 2488 7647 2522
rect 8041 2549 8075 2583
rect 8143 2549 8177 2583
rect 7709 2476 7743 2510
rect 8303 2534 8337 2568
rect 8579 2534 8613 2568
rect 8679 2538 8713 2572
rect 8810 2566 8844 2600
rect 8948 2550 8982 2584
rect 9116 2650 9150 2684
rect 9252 2650 9286 2684
rect 9354 2650 9388 2684
rect 9056 2498 9090 2532
rect 9451 2532 9485 2566
rect 9579 2566 9613 2600
rect 9731 2566 9765 2600
rect 9319 2476 9353 2510
rect 9899 2650 9933 2684
rect 10035 2650 10069 2684
rect 9833 2498 9867 2532
rect 10217 2536 10251 2570
rect 10005 2488 10039 2522
rect 10433 2549 10467 2583
rect 10535 2549 10569 2583
rect 10101 2476 10135 2510
rect 10695 2534 10729 2568
rect 10971 2534 11005 2568
rect 11071 2538 11105 2572
rect 11202 2566 11236 2600
rect 11340 2550 11374 2584
rect 11508 2650 11542 2684
rect 11644 2650 11678 2684
rect 11746 2650 11780 2684
rect 11448 2498 11482 2532
rect 11843 2532 11877 2566
rect 11971 2566 12005 2600
rect 12123 2566 12157 2600
rect 11711 2476 11745 2510
rect 12291 2650 12325 2684
rect 12427 2650 12461 2684
rect 12225 2498 12259 2532
rect 12609 2536 12643 2570
rect 12397 2488 12431 2522
rect 12825 2549 12859 2583
rect 12927 2549 12961 2583
rect 12493 2476 12527 2510
<< locali >>
rect 1035 6154 1064 6212
rect 1098 6154 1156 6212
rect 1190 6154 1248 6212
rect 1282 6154 1340 6212
rect 1374 6154 1432 6212
rect 1466 6154 1524 6212
rect 1558 6154 1616 6212
rect 1650 6188 1679 6212
rect 1650 6154 1708 6188
rect 1742 6154 1800 6188
rect 1834 6154 1863 6188
rect 2295 6154 2324 6212
rect 2358 6154 2416 6212
rect 2450 6154 2508 6212
rect 2542 6154 2600 6212
rect 2634 6154 2692 6212
rect 2726 6154 2784 6212
rect 2818 6154 2876 6212
rect 2910 6154 2968 6212
rect 3002 6154 3060 6212
rect 3094 6154 3152 6212
rect 3186 6154 3244 6212
rect 3278 6154 3336 6212
rect 3370 6154 3428 6212
rect 3462 6154 3520 6212
rect 3554 6154 3612 6212
rect 3646 6154 3704 6212
rect 3738 6154 3796 6212
rect 3830 6154 3888 6212
rect 3922 6154 3980 6212
rect 4014 6154 4072 6212
rect 4106 6154 4135 6212
rect 1068 6104 1104 6120
rect 1068 6070 1070 6104
rect 1068 6036 1104 6070
rect 1068 6002 1070 6036
rect 1140 6104 1206 6154
rect 1140 6070 1156 6104
rect 1190 6070 1206 6104
rect 1140 6036 1206 6070
rect 1140 6002 1156 6036
rect 1190 6002 1206 6036
rect 1240 6104 1294 6120
rect 1240 6070 1242 6104
rect 1276 6070 1294 6104
rect 1240 6023 1294 6070
rect 1068 5968 1104 6002
rect 1240 5989 1242 6023
rect 1276 5989 1294 6023
rect 1068 5934 1203 5968
rect 1240 5939 1294 5989
rect 1169 5905 1203 5934
rect 1056 5883 1124 5898
rect 1056 5849 1068 5883
rect 1102 5876 1124 5883
rect 1056 5842 1072 5849
rect 1106 5842 1124 5876
rect 1056 5824 1124 5842
rect 1169 5889 1224 5905
rect 1169 5855 1190 5889
rect 1169 5839 1224 5855
rect 1258 5884 1294 5939
rect 1330 6106 1396 6120
rect 1330 6072 1346 6106
rect 1380 6072 1396 6106
rect 1330 6038 1396 6072
rect 1330 6004 1346 6038
rect 1380 6004 1396 6038
rect 1330 5970 1396 6004
rect 1430 6112 1478 6154
rect 1464 6078 1478 6112
rect 1430 6044 1478 6078
rect 1464 6010 1478 6044
rect 1430 5994 1478 6010
rect 1514 6090 1548 6120
rect 1514 5995 1548 6056
rect 1330 5936 1346 5970
rect 1380 5958 1396 5970
rect 1582 6112 1648 6154
rect 1582 6078 1598 6112
rect 1632 6078 1648 6112
rect 1582 6044 1648 6078
rect 1582 6010 1598 6044
rect 1632 6010 1648 6044
rect 1582 5994 1648 6010
rect 1682 6090 1716 6120
rect 1682 5995 1716 6056
rect 1380 5936 1473 5958
rect 1330 5924 1473 5936
rect 1329 5884 1405 5890
rect 1258 5876 1405 5884
rect 1258 5846 1355 5876
rect 1169 5788 1203 5839
rect 1070 5754 1203 5788
rect 1258 5779 1294 5846
rect 1329 5842 1355 5846
rect 1389 5842 1405 5876
rect 1439 5876 1473 5924
rect 1514 5950 1548 5961
rect 1682 5950 1716 5961
rect 1514 5916 1716 5950
rect 1750 6112 1816 6154
rect 1750 6078 1766 6112
rect 1800 6078 1816 6112
rect 1750 6044 1816 6078
rect 1750 6010 1766 6044
rect 1800 6010 1816 6044
rect 1750 5976 1816 6010
rect 1750 5942 1766 5976
rect 1800 5942 1816 5976
rect 1750 5924 1816 5942
rect 2314 6112 2364 6154
rect 2314 6078 2330 6112
rect 2314 6044 2364 6078
rect 2314 6010 2330 6044
rect 2314 5976 2364 6010
rect 2314 5942 2330 5976
rect 2314 5926 2364 5942
rect 2398 6102 2463 6118
rect 2398 6068 2429 6102
rect 2398 5976 2463 6068
rect 2398 5942 2429 5976
rect 1617 5883 1716 5916
rect 2398 5888 2463 5942
rect 2497 6112 2547 6154
rect 2497 6078 2513 6112
rect 2497 6044 2547 6078
rect 2497 6010 2513 6044
rect 2497 5976 2547 6010
rect 2497 5942 2513 5976
rect 2497 5926 2547 5942
rect 2581 6102 2663 6118
rect 2581 6068 2613 6102
rect 2647 6068 2663 6102
rect 2581 6028 2663 6068
rect 2581 5994 2613 6028
rect 2647 5994 2663 6028
rect 2697 6112 2731 6154
rect 2697 6044 2731 6078
rect 2697 5994 2731 6010
rect 2765 6052 2783 6086
rect 2817 6052 2829 6086
rect 2879 6058 2895 6092
rect 2929 6058 3069 6092
rect 2581 5926 2643 5994
rect 2765 5960 2799 6052
rect 2677 5926 2799 5960
rect 2943 6018 3001 6024
rect 2943 5992 2967 6018
rect 2977 5958 3001 5984
rect 2841 5950 2909 5956
rect 2841 5926 2875 5950
rect 2581 5888 2615 5926
rect 2677 5892 2711 5926
rect 2875 5892 2909 5916
rect 1439 5842 1489 5876
rect 1523 5842 1539 5876
rect 1617 5849 1712 5883
rect 1746 5849 1756 5883
rect 2398 5880 2615 5888
rect 1439 5808 1473 5842
rect 1617 5808 1716 5849
rect 1070 5733 1104 5754
rect 1242 5750 1294 5779
rect 1070 5678 1104 5699
rect 1140 5686 1156 5720
rect 1190 5686 1206 5720
rect 1140 5644 1206 5686
rect 1276 5716 1294 5750
rect 1242 5678 1294 5716
rect 1346 5774 1473 5808
rect 1514 5774 1716 5808
rect 2398 5846 2410 5880
rect 2444 5846 2615 5880
rect 2398 5840 2615 5846
rect 1346 5756 1380 5774
rect 1514 5756 1548 5774
rect 1346 5678 1380 5722
rect 1416 5724 1464 5740
rect 1416 5690 1430 5724
rect 1416 5644 1464 5690
rect 1682 5756 1716 5774
rect 1514 5678 1548 5722
rect 1582 5724 1648 5740
rect 1582 5690 1598 5724
rect 1632 5690 1648 5724
rect 1582 5644 1648 5690
rect 1682 5678 1716 5722
rect 1750 5788 1816 5804
rect 1750 5754 1766 5788
rect 1800 5754 1816 5788
rect 1750 5720 1816 5754
rect 1750 5686 1766 5720
rect 1800 5686 1816 5720
rect 1750 5644 1816 5686
rect 2314 5788 2364 5804
rect 2314 5754 2330 5788
rect 2314 5720 2364 5754
rect 2314 5686 2330 5720
rect 2314 5644 2364 5686
rect 2398 5756 2463 5840
rect 2398 5722 2429 5756
rect 2398 5680 2463 5722
rect 2497 5788 2547 5804
rect 2497 5754 2513 5788
rect 2497 5720 2547 5754
rect 2497 5686 2513 5720
rect 2497 5644 2547 5686
rect 2581 5772 2615 5840
rect 2649 5876 2711 5892
rect 2683 5842 2711 5876
rect 2649 5826 2711 5842
rect 2745 5876 2807 5892
rect 2841 5876 2909 5892
rect 2779 5842 2807 5876
rect 2745 5826 2827 5842
rect 2943 5834 3001 5958
rect 2581 5756 2647 5772
rect 2581 5722 2613 5756
rect 2581 5680 2647 5722
rect 2681 5746 2731 5790
rect 2681 5712 2697 5746
rect 2681 5644 2731 5712
rect 2765 5743 2827 5826
rect 2877 5818 3001 5834
rect 2911 5784 3001 5818
rect 2877 5768 3001 5784
rect 3035 5974 3069 6058
rect 3114 6078 3183 6154
rect 3569 6088 3615 6154
rect 3148 6044 3183 6078
rect 3231 6052 3243 6086
rect 3277 6052 3336 6086
rect 3114 6028 3183 6044
rect 3217 5990 3255 6006
rect 3217 5974 3218 5990
rect 3035 5956 3218 5974
rect 3252 5956 3255 5990
rect 3035 5940 3255 5956
rect 2765 5709 2778 5743
rect 2812 5709 2827 5743
rect 3035 5720 3069 5940
rect 3111 5890 3185 5906
rect 3145 5884 3185 5890
rect 3111 5850 3138 5856
rect 3172 5850 3185 5884
rect 3111 5770 3185 5850
rect 3221 5744 3255 5940
rect 2765 5702 2827 5709
rect 2890 5686 2906 5720
rect 2940 5686 3069 5720
rect 3109 5720 3175 5736
rect 3109 5686 3110 5720
rect 3144 5686 3175 5720
rect 3109 5644 3175 5686
rect 3214 5728 3255 5744
rect 3248 5694 3255 5728
rect 3298 5989 3336 6052
rect 3298 5955 3302 5989
rect 3298 5746 3336 5955
rect 3332 5712 3336 5746
rect 3298 5696 3336 5712
rect 3370 6052 3427 6086
rect 3461 6052 3473 6086
rect 3569 6054 3574 6088
rect 3608 6054 3615 6088
rect 3966 6112 4032 6154
rect 3370 6039 3420 6052
rect 3370 6005 3386 6039
rect 3569 6038 3615 6054
rect 3686 6052 3703 6086
rect 3737 6052 3802 6086
rect 3836 6052 3852 6086
rect 3966 6078 3982 6112
rect 4016 6078 4032 6112
rect 4066 6086 4108 6102
rect 4100 6052 4108 6086
rect 3370 5989 3420 6005
rect 3370 5762 3404 5989
rect 3471 5984 3490 6018
rect 3524 5984 3540 6018
rect 3471 5959 3505 5984
rect 3451 5925 3505 5959
rect 3451 5905 3485 5925
rect 3438 5889 3485 5905
rect 3686 5908 3720 6052
rect 4066 6044 4108 6052
rect 4001 6018 4108 6044
rect 3754 5992 3795 6018
rect 3788 5984 3795 5992
rect 3829 6010 4108 6018
rect 3829 5984 4035 6010
rect 3788 5958 3822 5984
rect 3754 5942 3822 5958
rect 3472 5855 3485 5889
rect 3438 5839 3485 5855
rect 3370 5746 3417 5762
rect 3370 5712 3383 5746
rect 3370 5696 3417 5712
rect 3451 5720 3485 5839
rect 3519 5830 3577 5891
rect 3519 5813 3540 5830
rect 3574 5796 3577 5830
rect 3553 5779 3577 5796
rect 3519 5770 3577 5779
rect 3611 5830 3652 5891
rect 3686 5874 3754 5908
rect 3611 5813 3636 5830
rect 3611 5779 3613 5813
rect 3670 5796 3686 5830
rect 3647 5779 3686 5796
rect 3611 5770 3686 5779
rect 3578 5720 3644 5736
rect 3214 5678 3255 5694
rect 3451 5686 3487 5720
rect 3521 5686 3537 5720
rect 3578 5686 3586 5720
rect 3620 5686 3644 5720
rect 3720 5734 3754 5874
rect 3788 5834 3822 5942
rect 3856 5934 3887 5950
rect 3921 5916 3933 5950
rect 3856 5884 3890 5900
rect 3788 5818 3853 5834
rect 3788 5784 3819 5818
rect 3788 5768 3853 5784
rect 3887 5830 3967 5846
rect 3887 5796 3933 5830
rect 3887 5780 3967 5796
rect 4001 5788 4035 5984
rect 4069 5950 4105 5976
rect 4069 5916 4071 5950
rect 4069 5876 4105 5916
rect 4103 5842 4105 5876
rect 4069 5822 4105 5842
rect 3887 5752 3930 5780
rect 4001 5754 4108 5788
rect 3720 5700 3790 5734
rect 3824 5700 3840 5734
rect 3887 5718 3891 5752
rect 3925 5718 3930 5752
rect 4066 5746 4108 5754
rect 3887 5706 3930 5718
rect 3578 5644 3644 5686
rect 3966 5686 3982 5720
rect 4016 5686 4032 5720
rect 4100 5712 4108 5746
rect 4066 5696 4108 5712
rect 3966 5644 4032 5686
rect 1035 5586 1064 5644
rect 1098 5586 1156 5644
rect 1190 5586 1248 5644
rect 1282 5586 1340 5644
rect 1374 5586 1432 5644
rect 1466 5586 1524 5644
rect 1558 5586 1616 5644
rect 1650 5586 1708 5644
rect 1742 5586 1800 5644
rect 1834 5625 1863 5644
rect 2295 5625 2324 5644
rect 1834 5620 2324 5625
rect 2358 5620 2416 5644
rect 2450 5620 2508 5644
rect 2542 5620 2600 5644
rect 2634 5620 2692 5644
rect 2726 5620 2784 5644
rect 2818 5620 2876 5644
rect 2910 5620 2968 5644
rect 3002 5620 3060 5644
rect 3094 5620 3152 5644
rect 3186 5620 3244 5644
rect 3278 5620 3336 5644
rect 3370 5620 3428 5644
rect 3462 5620 3520 5644
rect 3554 5620 3612 5644
rect 3646 5620 3704 5644
rect 3738 5620 3796 5644
rect 3830 5620 3888 5644
rect 3922 5620 3980 5644
rect 4014 5620 4072 5644
rect 1834 5586 1892 5620
rect 1926 5586 1984 5620
rect 2018 5586 2076 5620
rect 2110 5586 2168 5620
rect 2202 5586 2260 5620
rect 2294 5610 2324 5620
rect 2386 5610 2416 5620
rect 2478 5610 2508 5620
rect 2570 5610 2600 5620
rect 2662 5610 2692 5620
rect 2754 5610 2784 5620
rect 2846 5610 2876 5620
rect 2938 5610 2968 5620
rect 3030 5610 3060 5620
rect 3122 5610 3152 5620
rect 3214 5610 3244 5620
rect 3306 5610 3336 5620
rect 3398 5610 3428 5620
rect 3490 5610 3520 5620
rect 3582 5610 3612 5620
rect 3674 5610 3704 5620
rect 3766 5610 3796 5620
rect 3858 5610 3888 5620
rect 3950 5610 3980 5620
rect 4042 5610 4072 5620
rect 4106 5610 4136 5644
rect 2294 5586 2352 5610
rect 2386 5586 2444 5610
rect 2478 5586 2536 5610
rect 2570 5586 2628 5610
rect 2662 5586 2720 5610
rect 2754 5586 2812 5610
rect 2846 5586 2904 5610
rect 2938 5586 2996 5610
rect 3030 5586 3088 5610
rect 3122 5586 3180 5610
rect 3214 5586 3272 5610
rect 3306 5586 3364 5610
rect 3398 5586 3456 5610
rect 3490 5586 3548 5610
rect 3582 5586 3640 5610
rect 3674 5586 3732 5610
rect 3766 5586 3824 5610
rect 3858 5586 3916 5610
rect 3950 5586 4008 5610
rect 4042 5586 4136 5610
rect 1034 5281 1063 5339
rect 1097 5281 1155 5339
rect 1189 5281 1247 5339
rect 1281 5281 1339 5339
rect 1373 5281 1431 5339
rect 1465 5281 1523 5339
rect 1557 5281 1615 5339
rect 1649 5281 1707 5339
rect 1741 5281 1799 5339
rect 1833 5281 1891 5339
rect 1925 5281 1983 5339
rect 2017 5281 2075 5339
rect 2109 5281 2167 5339
rect 2201 5281 2259 5339
rect 2293 5281 2351 5339
rect 2385 5281 2443 5339
rect 2477 5281 2535 5339
rect 2569 5281 2627 5339
rect 2661 5281 2719 5339
rect 2753 5281 2811 5339
rect 2845 5330 3087 5339
rect 2845 5315 2934 5330
rect 2968 5315 3087 5330
rect 2845 5281 2903 5315
rect 2968 5296 2995 5315
rect 2937 5281 2995 5296
rect 3029 5281 3087 5315
rect 3121 5281 3179 5339
rect 3213 5281 3271 5339
rect 3305 5281 3363 5339
rect 3397 5281 3455 5339
rect 3489 5281 3547 5339
rect 3581 5315 3640 5339
rect 3581 5281 3639 5315
rect 3674 5305 3731 5339
rect 3673 5281 3731 5305
rect 3765 5281 3823 5339
rect 3857 5281 3915 5339
rect 3949 5281 4007 5339
rect 4041 5333 4283 5339
rect 4041 5315 4177 5333
rect 4211 5315 4283 5333
rect 4041 5281 4099 5315
rect 4133 5299 4177 5315
rect 4133 5281 4191 5299
rect 4225 5281 4283 5315
rect 4317 5281 4375 5339
rect 4409 5281 4467 5339
rect 4501 5281 4559 5339
rect 4593 5281 4651 5339
rect 4685 5281 4743 5339
rect 4777 5281 4835 5339
rect 4869 5281 4927 5339
rect 4961 5281 5019 5339
rect 5053 5281 5111 5339
rect 5145 5281 5203 5339
rect 5237 5281 5295 5339
rect 5329 5281 5387 5339
rect 5421 5281 5479 5339
rect 5513 5281 5571 5339
rect 5605 5281 5663 5339
rect 5697 5281 5755 5339
rect 5789 5281 5847 5339
rect 5881 5281 5939 5339
rect 5973 5281 6031 5339
rect 6065 5281 6123 5339
rect 6157 5281 6215 5339
rect 6249 5281 6307 5339
rect 6341 5281 6399 5339
rect 6433 5335 6675 5339
rect 6433 5315 6569 5335
rect 6603 5315 6675 5335
rect 6433 5281 6491 5315
rect 6525 5301 6569 5315
rect 6525 5281 6583 5301
rect 6617 5281 6675 5315
rect 6709 5281 6767 5339
rect 6801 5281 6859 5339
rect 6893 5281 6951 5339
rect 6985 5281 7043 5339
rect 7077 5281 7135 5339
rect 7169 5281 7227 5339
rect 7261 5281 7319 5339
rect 7353 5281 7411 5339
rect 7445 5281 7503 5339
rect 7537 5281 7595 5339
rect 7629 5281 7687 5339
rect 7721 5281 7779 5339
rect 7813 5281 7871 5339
rect 7905 5281 7963 5339
rect 7997 5281 8055 5339
rect 8089 5281 8147 5339
rect 8181 5281 8239 5339
rect 8273 5281 8331 5339
rect 8365 5281 8423 5339
rect 8457 5281 8515 5339
rect 8549 5281 8607 5339
rect 8641 5281 8699 5339
rect 8733 5281 8791 5339
rect 8825 5335 9067 5339
rect 8825 5315 8961 5335
rect 8995 5315 9067 5335
rect 8825 5281 8883 5315
rect 8917 5301 8961 5315
rect 8917 5281 8975 5301
rect 9009 5281 9067 5315
rect 9101 5281 9159 5339
rect 9193 5281 9251 5339
rect 9285 5281 9343 5339
rect 9377 5281 9435 5339
rect 9469 5281 9527 5339
rect 9561 5281 9619 5339
rect 9653 5281 9711 5339
rect 9745 5281 9803 5339
rect 9837 5281 9895 5339
rect 9929 5281 9987 5339
rect 10021 5281 10079 5339
rect 10113 5281 10171 5339
rect 10205 5281 10263 5339
rect 10297 5281 10355 5339
rect 10389 5281 10447 5339
rect 10481 5281 10539 5339
rect 10573 5281 10631 5339
rect 10665 5281 10723 5339
rect 10757 5281 10815 5339
rect 10849 5281 10907 5339
rect 10941 5281 10999 5339
rect 11033 5281 11091 5339
rect 11125 5281 11183 5339
rect 11217 5336 11459 5339
rect 11217 5315 11353 5336
rect 11387 5315 11459 5336
rect 11217 5281 11275 5315
rect 11309 5302 11353 5315
rect 11309 5281 11367 5302
rect 11401 5281 11459 5315
rect 11493 5281 11551 5339
rect 11585 5281 11643 5339
rect 11677 5281 11735 5339
rect 11769 5281 11827 5339
rect 11861 5281 11919 5339
rect 11953 5281 12011 5339
rect 12045 5281 12103 5339
rect 12137 5281 12195 5339
rect 12229 5281 12287 5339
rect 12321 5281 12379 5339
rect 12413 5281 12471 5339
rect 12505 5281 12563 5339
rect 12597 5281 12655 5339
rect 12689 5281 12747 5339
rect 12781 5281 12839 5339
rect 12873 5281 12931 5339
rect 12965 5281 12994 5339
rect 1051 5231 1103 5247
rect 1051 5197 1069 5231
rect 1051 5163 1103 5197
rect 1137 5215 1203 5281
rect 1137 5181 1153 5215
rect 1187 5181 1203 5215
rect 1237 5231 1282 5247
rect 1271 5197 1282 5231
rect 1051 5129 1069 5163
rect 1237 5163 1282 5197
rect 1321 5215 1391 5281
rect 1321 5181 1341 5215
rect 1375 5181 1391 5215
rect 1425 5231 1459 5247
rect 1502 5204 1518 5238
rect 1552 5204 1668 5238
rect 1103 5145 1202 5147
rect 1103 5129 1156 5145
rect 1051 5113 1156 5129
rect 1190 5111 1202 5145
rect 1051 5018 1122 5079
rect 1051 4984 1066 5018
rect 1100 4994 1122 5018
rect 1051 4960 1067 4984
rect 1101 4960 1122 4994
rect 1051 4949 1122 4960
rect 1156 5018 1202 5111
rect 1156 4984 1168 5018
rect 1156 4915 1202 4984
rect 1051 4881 1202 4915
rect 1271 5129 1282 5163
rect 1425 5147 1459 5197
rect 1237 4941 1282 5129
rect 1237 4907 1248 4941
rect 1051 4873 1103 4881
rect 1051 4839 1069 4873
rect 1237 4873 1282 4907
rect 1316 5113 1459 5147
rect 1316 4919 1350 5113
rect 1500 5111 1524 5145
rect 1558 5119 1600 5145
rect 1558 5111 1566 5119
rect 1500 5085 1566 5111
rect 1384 5074 1466 5079
rect 1384 5040 1428 5074
rect 1462 5040 1466 5074
rect 1384 5005 1466 5040
rect 1418 4971 1466 5005
rect 1384 4955 1466 4971
rect 1500 5069 1600 5085
rect 1500 4945 1544 5069
rect 1634 5035 1668 5204
rect 1716 5229 1792 5281
rect 2010 5239 2076 5281
rect 1716 5195 1732 5229
rect 1766 5195 1792 5229
rect 1852 5213 1886 5229
rect 1852 5161 1886 5179
rect 2010 5205 2026 5239
rect 2060 5205 2076 5239
rect 2499 5239 2575 5281
rect 2010 5171 2076 5205
rect 2285 5204 2301 5238
rect 2335 5204 2451 5238
rect 2499 5205 2515 5239
rect 2549 5205 2575 5239
rect 2763 5239 3040 5281
rect 2623 5213 2657 5229
rect 1702 5145 1972 5161
rect 1702 5119 1852 5145
rect 1736 5111 1852 5119
rect 1886 5111 1972 5145
rect 2010 5137 2026 5171
rect 2060 5137 2076 5171
rect 2247 5145 2294 5151
rect 1736 5085 1752 5111
rect 1702 5069 1752 5085
rect 1854 5035 1904 5051
rect 1634 5001 1870 5035
rect 1634 4993 1714 5001
rect 1316 4881 1459 4919
rect 1534 4911 1544 4945
rect 1500 4895 1544 4911
rect 1580 4923 1596 4957
rect 1630 4941 1646 4957
rect 1580 4907 1612 4923
rect 1580 4883 1646 4907
rect 1051 4823 1103 4839
rect 1137 4813 1153 4847
rect 1187 4813 1203 4847
rect 1271 4839 1282 4873
rect 1425 4865 1459 4881
rect 1237 4823 1282 4839
rect 1137 4771 1203 4813
rect 1321 4813 1341 4847
rect 1375 4813 1391 4847
rect 1680 4847 1714 4993
rect 1860 4985 1904 5001
rect 1938 4967 1972 5111
rect 2247 5119 2260 5145
rect 2281 5085 2294 5111
rect 2006 5077 2207 5085
rect 2006 5043 2168 5077
rect 2202 5043 2207 5077
rect 2247 5069 2294 5085
rect 2342 5119 2383 5135
rect 2342 5085 2349 5119
rect 2006 5037 2207 5043
rect 2006 5035 2072 5037
rect 2006 5001 2022 5035
rect 2056 5001 2072 5035
rect 2342 5015 2383 5085
rect 2259 5009 2383 5015
rect 2134 4967 2150 5001
rect 2184 4967 2200 5001
rect 1752 4933 1768 4967
rect 1802 4947 1818 4967
rect 1802 4941 1834 4947
rect 1752 4907 1800 4933
rect 1938 4933 2200 4967
rect 2259 4975 2260 5009
rect 2294 4979 2383 5009
rect 2417 5035 2451 5204
rect 2763 5205 2779 5239
rect 2813 5205 2990 5239
rect 3024 5205 3040 5239
rect 2623 5171 2657 5179
rect 3074 5202 3131 5247
rect 2485 5137 3040 5171
rect 2485 5119 2535 5137
rect 2519 5085 2535 5119
rect 2485 5069 2535 5085
rect 2417 5019 2687 5035
rect 2417 5001 2653 5019
rect 2294 4975 2316 4979
rect 2259 4945 2316 4975
rect 1938 4907 1982 4933
rect 1752 4901 1834 4907
rect 1916 4873 1932 4907
rect 1966 4873 1982 4907
rect 2259 4911 2282 4945
rect 2016 4881 2050 4897
rect 2259 4895 2316 4911
rect 1425 4815 1459 4831
rect 1321 4771 1391 4813
rect 1515 4813 1531 4847
rect 1565 4813 1714 4847
rect 1515 4807 1714 4813
rect 1748 4843 1782 4859
rect 1748 4771 1782 4809
rect 1816 4829 1832 4863
rect 1866 4839 1882 4863
rect 2417 4847 2451 5001
rect 2643 4985 2653 5001
rect 2643 4969 2687 4985
rect 2526 4941 2545 4967
rect 2526 4907 2536 4941
rect 2579 4933 2601 4967
rect 2570 4907 2601 4933
rect 2721 4910 2757 5137
rect 2526 4901 2601 4907
rect 2691 4907 2757 4910
rect 2691 4873 2707 4907
rect 2741 4873 2757 4907
rect 2791 5077 2893 5103
rect 2791 5043 2812 5077
rect 2846 5069 2893 5077
rect 2927 5069 2943 5103
rect 2791 5035 2846 5043
rect 2825 5001 2846 5035
rect 3006 5019 3040 5137
rect 3108 5168 3131 5202
rect 3074 5134 3131 5168
rect 3108 5100 3131 5134
rect 3074 5080 3131 5100
rect 2791 4939 2846 5001
rect 2897 5007 2972 5019
rect 2897 4973 2922 5007
rect 2956 4973 2972 5007
rect 3006 5003 3056 5019
rect 3006 4969 3022 5003
rect 3006 4953 3056 4969
rect 2791 4905 2929 4939
rect 2016 4839 2050 4847
rect 1866 4829 2050 4839
rect 1816 4805 2050 4829
rect 2104 4813 2120 4847
rect 2154 4813 2170 4847
rect 2104 4771 2170 4813
rect 2298 4813 2314 4847
rect 2348 4813 2451 4847
rect 2298 4807 2451 4813
rect 2487 4843 2539 4859
rect 2487 4809 2505 4843
rect 2487 4771 2539 4809
rect 2591 4829 2607 4863
rect 2641 4839 2657 4863
rect 2791 4855 2825 4871
rect 2641 4829 2791 4839
rect 2591 4821 2791 4829
rect 2591 4805 2825 4821
rect 2882 4857 2929 4905
rect 2882 4823 2895 4857
rect 2882 4807 2929 4823
rect 2974 4847 3040 4915
rect 3090 4897 3131 5080
rect 2974 4813 2990 4847
rect 3024 4813 3040 4847
rect 2974 4771 3040 4813
rect 3074 4883 3131 4897
rect 3074 4881 3087 4883
rect 3121 4849 3131 4883
rect 3108 4847 3131 4849
rect 3074 4805 3131 4847
rect 3165 5221 3228 5237
rect 3165 5187 3178 5221
rect 3212 5187 3228 5221
rect 3165 5153 3228 5187
rect 3165 5119 3178 5153
rect 3212 5119 3228 5153
rect 3165 5019 3228 5119
rect 3264 5227 3323 5281
rect 3264 5193 3273 5227
rect 3307 5193 3323 5227
rect 3264 5159 3323 5193
rect 3264 5125 3273 5159
rect 3307 5125 3323 5159
rect 3264 5107 3323 5125
rect 3357 5203 3409 5247
rect 3391 5169 3409 5203
rect 3357 5135 3409 5169
rect 3391 5101 3409 5135
rect 3443 5231 3495 5247
rect 3443 5197 3461 5231
rect 3443 5163 3495 5197
rect 3529 5215 3595 5281
rect 3529 5181 3545 5215
rect 3579 5181 3595 5215
rect 3629 5231 3674 5247
rect 3663 5197 3674 5231
rect 3443 5129 3461 5163
rect 3629 5163 3674 5197
rect 3713 5215 3783 5281
rect 3713 5181 3733 5215
rect 3767 5181 3783 5215
rect 3817 5231 3851 5247
rect 3894 5204 3910 5238
rect 3944 5204 4060 5238
rect 3495 5145 3594 5147
rect 3495 5129 3548 5145
rect 3443 5113 3548 5129
rect 3357 5081 3409 5101
rect 3357 5047 3368 5081
rect 3402 5047 3409 5081
rect 3582 5111 3594 5145
rect 3357 5043 3409 5047
rect 3165 5003 3332 5019
rect 3165 4969 3298 5003
rect 3165 4953 3332 4969
rect 3165 4873 3228 4953
rect 3366 4919 3409 5043
rect 3443 5018 3514 5079
rect 3443 4994 3458 5018
rect 3443 4960 3457 4994
rect 3492 4984 3514 5018
rect 3491 4960 3514 4984
rect 3443 4949 3514 4960
rect 3548 5018 3594 5111
rect 3548 4984 3560 5018
rect 3165 4839 3178 4873
rect 3212 4839 3228 4873
rect 3357 4883 3409 4919
rect 3548 4915 3594 4984
rect 3165 4805 3228 4839
rect 3264 4847 3323 4863
rect 3264 4813 3273 4847
rect 3307 4813 3323 4847
rect 3264 4771 3323 4813
rect 3391 4849 3409 4883
rect 3357 4805 3409 4849
rect 3443 4881 3594 4915
rect 3663 5129 3674 5163
rect 3817 5147 3851 5197
rect 3629 4941 3674 5129
rect 3629 4907 3640 4941
rect 3443 4873 3495 4881
rect 3443 4839 3461 4873
rect 3629 4873 3674 4907
rect 3708 5113 3851 5147
rect 3708 4919 3742 5113
rect 3892 5111 3916 5145
rect 3950 5119 3992 5145
rect 3950 5111 3958 5119
rect 3892 5085 3958 5111
rect 3776 5077 3858 5079
rect 3776 5043 3779 5077
rect 3813 5043 3858 5077
rect 3776 5005 3858 5043
rect 3810 4971 3858 5005
rect 3776 4955 3858 4971
rect 3892 5069 3992 5085
rect 3892 4945 3936 5069
rect 4026 5035 4060 5204
rect 4108 5229 4184 5281
rect 4402 5239 4468 5281
rect 4108 5195 4124 5229
rect 4158 5195 4184 5229
rect 4244 5213 4278 5229
rect 4244 5161 4278 5179
rect 4402 5205 4418 5239
rect 4452 5205 4468 5239
rect 4891 5239 4967 5281
rect 4402 5171 4468 5205
rect 4677 5204 4693 5238
rect 4727 5204 4843 5238
rect 4891 5205 4907 5239
rect 4941 5205 4967 5239
rect 5155 5239 5432 5281
rect 5015 5213 5049 5229
rect 4094 5145 4364 5161
rect 4094 5119 4244 5145
rect 4128 5111 4244 5119
rect 4278 5111 4364 5145
rect 4402 5137 4418 5171
rect 4452 5137 4468 5171
rect 4639 5145 4686 5151
rect 4128 5085 4144 5111
rect 4094 5069 4144 5085
rect 4246 5035 4296 5051
rect 4026 5001 4262 5035
rect 4026 4993 4106 5001
rect 3708 4881 3851 4919
rect 3926 4911 3936 4945
rect 3892 4895 3936 4911
rect 3972 4923 3988 4957
rect 4022 4941 4038 4957
rect 3972 4907 4004 4923
rect 3972 4883 4038 4907
rect 3443 4823 3495 4839
rect 3529 4813 3545 4847
rect 3579 4813 3595 4847
rect 3663 4839 3674 4873
rect 3817 4865 3851 4881
rect 3629 4823 3674 4839
rect 3529 4771 3595 4813
rect 3713 4813 3733 4847
rect 3767 4813 3783 4847
rect 4072 4847 4106 4993
rect 4252 4985 4296 5001
rect 4330 4967 4364 5111
rect 4639 5119 4652 5145
rect 4673 5085 4686 5111
rect 4398 5077 4599 5085
rect 4398 5043 4560 5077
rect 4594 5043 4599 5077
rect 4639 5069 4686 5085
rect 4734 5119 4775 5135
rect 4734 5085 4741 5119
rect 4398 5037 4599 5043
rect 4398 5035 4464 5037
rect 4398 5001 4414 5035
rect 4448 5001 4464 5035
rect 4734 5015 4775 5085
rect 4651 5009 4775 5015
rect 4526 4967 4542 5001
rect 4576 4967 4592 5001
rect 4144 4933 4160 4967
rect 4194 4947 4210 4967
rect 4194 4941 4226 4947
rect 4144 4907 4192 4933
rect 4330 4933 4592 4967
rect 4651 4975 4652 5009
rect 4686 4979 4775 5009
rect 4809 5035 4843 5204
rect 5155 5205 5171 5239
rect 5205 5205 5382 5239
rect 5416 5205 5432 5239
rect 5015 5171 5049 5179
rect 5466 5202 5523 5247
rect 4877 5137 5432 5171
rect 4877 5119 4927 5137
rect 4911 5085 4927 5119
rect 4877 5069 4927 5085
rect 4809 5019 5079 5035
rect 4809 5001 5045 5019
rect 4686 4975 4708 4979
rect 4651 4945 4708 4975
rect 4330 4907 4374 4933
rect 4144 4901 4226 4907
rect 4308 4873 4324 4907
rect 4358 4873 4374 4907
rect 4651 4911 4674 4945
rect 4408 4881 4442 4897
rect 4651 4895 4708 4911
rect 3817 4815 3851 4831
rect 3713 4771 3783 4813
rect 3907 4813 3923 4847
rect 3957 4813 4106 4847
rect 3907 4807 4106 4813
rect 4140 4843 4174 4859
rect 4140 4771 4174 4809
rect 4208 4829 4224 4863
rect 4258 4839 4274 4863
rect 4809 4847 4843 5001
rect 5035 4985 5045 5001
rect 5035 4969 5079 4985
rect 4918 4941 4937 4967
rect 4918 4907 4928 4941
rect 4971 4933 4993 4967
rect 4962 4907 4993 4933
rect 5113 4910 5149 5137
rect 4918 4901 4993 4907
rect 5083 4907 5149 4910
rect 5083 4873 5099 4907
rect 5133 4873 5149 4907
rect 5183 5077 5285 5103
rect 5183 5043 5204 5077
rect 5238 5069 5285 5077
rect 5319 5069 5335 5103
rect 5183 5035 5238 5043
rect 5217 5001 5238 5035
rect 5398 5019 5432 5137
rect 5500 5168 5523 5202
rect 5466 5134 5523 5168
rect 5500 5100 5523 5134
rect 5466 5080 5523 5100
rect 5183 4939 5238 5001
rect 5289 5011 5364 5019
rect 5289 4977 5305 5011
rect 5339 5007 5364 5011
rect 5289 4973 5314 4977
rect 5348 4973 5364 5007
rect 5398 5003 5448 5019
rect 5398 4969 5414 5003
rect 5398 4953 5448 4969
rect 5183 4905 5321 4939
rect 4408 4839 4442 4847
rect 4258 4829 4442 4839
rect 4208 4805 4442 4829
rect 4496 4813 4512 4847
rect 4546 4813 4562 4847
rect 4496 4771 4562 4813
rect 4690 4813 4706 4847
rect 4740 4813 4843 4847
rect 4690 4807 4843 4813
rect 4879 4843 4931 4859
rect 4879 4809 4897 4843
rect 4879 4771 4931 4809
rect 4983 4829 4999 4863
rect 5033 4839 5049 4863
rect 5183 4855 5217 4871
rect 5033 4829 5183 4839
rect 4983 4821 5183 4829
rect 4983 4805 5217 4821
rect 5274 4857 5321 4905
rect 5274 4823 5287 4857
rect 5274 4807 5321 4823
rect 5366 4847 5432 4915
rect 5482 4897 5523 5080
rect 5366 4813 5382 4847
rect 5416 4813 5432 4847
rect 5366 4771 5432 4813
rect 5466 4894 5523 4897
rect 5466 4881 5476 4894
rect 5510 4860 5523 4894
rect 5500 4847 5523 4860
rect 5466 4805 5523 4847
rect 5557 5221 5620 5237
rect 5557 5187 5570 5221
rect 5604 5187 5620 5221
rect 5557 5153 5620 5187
rect 5557 5119 5570 5153
rect 5604 5119 5620 5153
rect 5557 5019 5620 5119
rect 5656 5227 5715 5281
rect 5656 5193 5665 5227
rect 5699 5193 5715 5227
rect 5656 5159 5715 5193
rect 5656 5125 5665 5159
rect 5699 5125 5715 5159
rect 5656 5107 5715 5125
rect 5749 5203 5801 5247
rect 5783 5169 5801 5203
rect 5749 5135 5801 5169
rect 5783 5101 5801 5135
rect 5835 5231 5887 5247
rect 5835 5197 5853 5231
rect 5835 5163 5887 5197
rect 5921 5215 5987 5281
rect 5921 5181 5937 5215
rect 5971 5181 5987 5215
rect 6021 5231 6066 5247
rect 6055 5197 6066 5231
rect 5835 5129 5853 5163
rect 6021 5163 6066 5197
rect 6105 5215 6175 5281
rect 6105 5181 6125 5215
rect 6159 5181 6175 5215
rect 6209 5231 6243 5247
rect 6286 5204 6302 5238
rect 6336 5204 6452 5238
rect 5887 5145 5986 5147
rect 5887 5129 5940 5145
rect 5835 5113 5940 5129
rect 5749 5080 5801 5101
rect 5749 5046 5757 5080
rect 5791 5046 5801 5080
rect 5974 5111 5986 5145
rect 5749 5043 5801 5046
rect 5557 5003 5724 5019
rect 5557 4969 5690 5003
rect 5557 4953 5724 4969
rect 5557 4873 5620 4953
rect 5758 4919 5801 5043
rect 5835 5018 5906 5079
rect 5835 4961 5850 5018
rect 5884 4961 5906 5018
rect 5835 4949 5906 4961
rect 5940 5018 5986 5111
rect 5940 4984 5952 5018
rect 5749 4906 5801 4919
rect 5940 4915 5986 4984
rect 5557 4839 5570 4873
rect 5604 4839 5620 4873
rect 5782 4883 5801 4906
rect 5557 4805 5620 4839
rect 5656 4847 5715 4863
rect 5656 4813 5665 4847
rect 5699 4813 5715 4847
rect 5656 4771 5715 4813
rect 5783 4849 5801 4883
rect 5749 4805 5801 4849
rect 5835 4881 5986 4915
rect 6055 5129 6066 5163
rect 6209 5147 6243 5197
rect 6021 4941 6066 5129
rect 6021 4907 6032 4941
rect 5835 4873 5887 4881
rect 5835 4839 5853 4873
rect 6021 4873 6066 4907
rect 6100 5113 6243 5147
rect 6100 4919 6134 5113
rect 6284 5111 6308 5145
rect 6342 5119 6384 5145
rect 6342 5111 6350 5119
rect 6284 5085 6350 5111
rect 6168 5076 6250 5079
rect 6202 5042 6250 5076
rect 6168 5005 6250 5042
rect 6202 4971 6250 5005
rect 6168 4955 6250 4971
rect 6284 5069 6384 5085
rect 6284 4945 6328 5069
rect 6418 5035 6452 5204
rect 6500 5229 6576 5281
rect 6794 5239 6860 5281
rect 6500 5195 6516 5229
rect 6550 5195 6576 5229
rect 6636 5213 6670 5229
rect 6636 5161 6670 5179
rect 6794 5205 6810 5239
rect 6844 5205 6860 5239
rect 7283 5239 7359 5281
rect 6794 5171 6860 5205
rect 7069 5204 7085 5238
rect 7119 5204 7235 5238
rect 7283 5205 7299 5239
rect 7333 5205 7359 5239
rect 7547 5239 7824 5281
rect 7407 5213 7441 5229
rect 6486 5145 6756 5161
rect 6486 5119 6636 5145
rect 6520 5111 6636 5119
rect 6670 5111 6756 5145
rect 6794 5137 6810 5171
rect 6844 5137 6860 5171
rect 7031 5145 7078 5151
rect 6520 5085 6536 5111
rect 6486 5069 6536 5085
rect 6638 5035 6688 5051
rect 6418 5001 6654 5035
rect 6418 4993 6498 5001
rect 6100 4881 6243 4919
rect 6318 4911 6328 4945
rect 6284 4895 6328 4911
rect 6364 4923 6380 4957
rect 6414 4941 6430 4957
rect 6364 4907 6396 4923
rect 6364 4883 6430 4907
rect 5835 4823 5887 4839
rect 5921 4813 5937 4847
rect 5971 4813 5987 4847
rect 6055 4839 6066 4873
rect 6209 4865 6243 4881
rect 6021 4823 6066 4839
rect 5921 4771 5987 4813
rect 6105 4813 6125 4847
rect 6159 4813 6175 4847
rect 6464 4847 6498 4993
rect 6644 4985 6688 5001
rect 6722 4967 6756 5111
rect 7031 5119 7044 5145
rect 7065 5085 7078 5111
rect 6790 5077 6991 5085
rect 6790 5043 6952 5077
rect 6986 5043 6991 5077
rect 7031 5069 7078 5085
rect 7126 5119 7167 5135
rect 7126 5085 7133 5119
rect 6790 5037 6991 5043
rect 6790 5035 6856 5037
rect 6790 5001 6806 5035
rect 6840 5001 6856 5035
rect 7126 5015 7167 5085
rect 7043 5009 7167 5015
rect 6918 4967 6934 5001
rect 6968 4967 6984 5001
rect 6536 4933 6552 4967
rect 6586 4947 6602 4967
rect 6586 4941 6618 4947
rect 6536 4907 6584 4933
rect 6722 4933 6984 4967
rect 7043 4975 7044 5009
rect 7078 4979 7167 5009
rect 7201 5035 7235 5204
rect 7547 5205 7563 5239
rect 7597 5205 7774 5239
rect 7808 5205 7824 5239
rect 7407 5171 7441 5179
rect 7858 5202 7915 5247
rect 7269 5137 7824 5171
rect 7269 5119 7319 5137
rect 7303 5085 7319 5119
rect 7269 5069 7319 5085
rect 7201 5019 7471 5035
rect 7201 5001 7437 5019
rect 7078 4975 7100 4979
rect 7043 4945 7100 4975
rect 6722 4907 6766 4933
rect 6536 4901 6618 4907
rect 6700 4873 6716 4907
rect 6750 4873 6766 4907
rect 7043 4911 7066 4945
rect 6800 4881 6834 4897
rect 7043 4895 7100 4911
rect 6209 4815 6243 4831
rect 6105 4771 6175 4813
rect 6299 4813 6315 4847
rect 6349 4813 6498 4847
rect 6299 4807 6498 4813
rect 6532 4843 6566 4859
rect 6532 4771 6566 4809
rect 6600 4829 6616 4863
rect 6650 4839 6666 4863
rect 7201 4847 7235 5001
rect 7427 4985 7437 5001
rect 7427 4969 7471 4985
rect 7310 4941 7329 4967
rect 7310 4907 7320 4941
rect 7363 4933 7385 4967
rect 7354 4907 7385 4933
rect 7505 4910 7541 5137
rect 7310 4901 7385 4907
rect 7475 4907 7541 4910
rect 7475 4873 7491 4907
rect 7525 4873 7541 4907
rect 7575 5077 7677 5103
rect 7575 5043 7596 5077
rect 7630 5069 7677 5077
rect 7711 5069 7727 5103
rect 7575 5035 7630 5043
rect 7609 5001 7630 5035
rect 7790 5019 7824 5137
rect 7892 5168 7915 5202
rect 7858 5134 7915 5168
rect 7892 5100 7915 5134
rect 7858 5080 7915 5100
rect 7575 4939 7630 5001
rect 7681 5012 7756 5019
rect 7681 4978 7695 5012
rect 7729 5007 7756 5012
rect 7681 4973 7706 4978
rect 7740 4973 7756 5007
rect 7790 5003 7840 5019
rect 7790 4969 7806 5003
rect 7790 4953 7840 4969
rect 7575 4905 7713 4939
rect 6800 4839 6834 4847
rect 6650 4829 6834 4839
rect 6600 4805 6834 4829
rect 6888 4813 6904 4847
rect 6938 4813 6954 4847
rect 6888 4771 6954 4813
rect 7082 4813 7098 4847
rect 7132 4813 7235 4847
rect 7082 4807 7235 4813
rect 7271 4843 7323 4859
rect 7271 4809 7289 4843
rect 7271 4771 7323 4809
rect 7375 4829 7391 4863
rect 7425 4839 7441 4863
rect 7575 4855 7609 4871
rect 7425 4829 7575 4839
rect 7375 4821 7575 4829
rect 7375 4805 7609 4821
rect 7666 4857 7713 4905
rect 7666 4823 7679 4857
rect 7666 4807 7713 4823
rect 7758 4847 7824 4915
rect 7874 4897 7915 5080
rect 7758 4813 7774 4847
rect 7808 4813 7824 4847
rect 7758 4771 7824 4813
rect 7858 4881 7864 4897
rect 7898 4863 7915 4897
rect 7892 4847 7915 4863
rect 7858 4805 7915 4847
rect 7949 5221 8012 5237
rect 7949 5187 7962 5221
rect 7996 5187 8012 5221
rect 7949 5153 8012 5187
rect 7949 5119 7962 5153
rect 7996 5119 8012 5153
rect 7949 5019 8012 5119
rect 8048 5227 8107 5281
rect 8048 5193 8057 5227
rect 8091 5193 8107 5227
rect 8048 5159 8107 5193
rect 8048 5125 8057 5159
rect 8091 5125 8107 5159
rect 8048 5107 8107 5125
rect 8141 5203 8193 5247
rect 8175 5169 8193 5203
rect 8141 5135 8193 5169
rect 8175 5101 8193 5135
rect 8227 5231 8279 5247
rect 8227 5197 8245 5231
rect 8227 5163 8279 5197
rect 8313 5215 8379 5281
rect 8313 5181 8329 5215
rect 8363 5181 8379 5215
rect 8413 5231 8458 5247
rect 8447 5197 8458 5231
rect 8227 5129 8245 5163
rect 8413 5163 8458 5197
rect 8497 5215 8567 5281
rect 8497 5181 8517 5215
rect 8551 5181 8567 5215
rect 8601 5231 8635 5247
rect 8678 5204 8694 5238
rect 8728 5204 8844 5238
rect 8279 5145 8378 5147
rect 8279 5129 8332 5145
rect 8227 5113 8332 5129
rect 8141 5078 8193 5101
rect 8366 5111 8378 5145
rect 8141 5044 8152 5078
rect 8186 5044 8193 5078
rect 8141 5043 8193 5044
rect 7949 5003 8116 5019
rect 7949 4969 8082 5003
rect 7949 4953 8116 4969
rect 7949 4873 8012 4953
rect 8150 4919 8193 5043
rect 8227 5018 8298 5079
rect 8227 4960 8242 5018
rect 8276 4960 8298 5018
rect 8227 4949 8298 4960
rect 8332 5018 8378 5111
rect 8332 4984 8344 5018
rect 7949 4839 7962 4873
rect 7996 4839 8012 4873
rect 8141 4895 8193 4919
rect 8332 4915 8378 4984
rect 8141 4883 8144 4895
rect 7949 4805 8012 4839
rect 8048 4847 8107 4863
rect 8048 4813 8057 4847
rect 8091 4813 8107 4847
rect 8048 4771 8107 4813
rect 8178 4861 8193 4895
rect 8175 4849 8193 4861
rect 8141 4805 8193 4849
rect 8227 4881 8378 4915
rect 8447 5129 8458 5163
rect 8601 5147 8635 5197
rect 8413 4941 8458 5129
rect 8413 4907 8424 4941
rect 8227 4873 8279 4881
rect 8227 4839 8245 4873
rect 8413 4873 8458 4907
rect 8492 5113 8635 5147
rect 8492 4919 8526 5113
rect 8676 5111 8700 5145
rect 8734 5119 8776 5145
rect 8734 5111 8742 5119
rect 8676 5085 8742 5111
rect 8560 5074 8642 5079
rect 8560 5040 8563 5074
rect 8597 5040 8642 5074
rect 8560 5005 8642 5040
rect 8594 4971 8642 5005
rect 8560 4955 8642 4971
rect 8676 5069 8776 5085
rect 8676 4945 8720 5069
rect 8810 5035 8844 5204
rect 8892 5229 8968 5281
rect 9186 5239 9252 5281
rect 8892 5195 8908 5229
rect 8942 5195 8968 5229
rect 9028 5213 9062 5229
rect 9028 5161 9062 5179
rect 9186 5205 9202 5239
rect 9236 5205 9252 5239
rect 9675 5239 9751 5281
rect 9186 5171 9252 5205
rect 9461 5204 9477 5238
rect 9511 5204 9627 5238
rect 9675 5205 9691 5239
rect 9725 5205 9751 5239
rect 9939 5239 10216 5281
rect 9799 5213 9833 5229
rect 8878 5145 9148 5161
rect 8878 5119 9028 5145
rect 8912 5111 9028 5119
rect 9062 5111 9148 5145
rect 9186 5137 9202 5171
rect 9236 5137 9252 5171
rect 9423 5145 9470 5151
rect 8912 5085 8928 5111
rect 8878 5069 8928 5085
rect 9030 5035 9080 5051
rect 8810 5001 9046 5035
rect 8810 4993 8890 5001
rect 8492 4881 8635 4919
rect 8710 4911 8720 4945
rect 8676 4895 8720 4911
rect 8756 4923 8772 4957
rect 8806 4941 8822 4957
rect 8756 4907 8788 4923
rect 8756 4883 8822 4907
rect 8227 4823 8279 4839
rect 8313 4813 8329 4847
rect 8363 4813 8379 4847
rect 8447 4839 8458 4873
rect 8601 4865 8635 4881
rect 8413 4823 8458 4839
rect 8313 4771 8379 4813
rect 8497 4813 8517 4847
rect 8551 4813 8567 4847
rect 8856 4847 8890 4993
rect 9036 4985 9080 5001
rect 9114 4967 9148 5111
rect 9423 5119 9436 5145
rect 9457 5085 9470 5111
rect 9182 5077 9383 5085
rect 9182 5043 9344 5077
rect 9378 5043 9383 5077
rect 9423 5069 9470 5085
rect 9518 5119 9559 5135
rect 9518 5085 9525 5119
rect 9182 5037 9383 5043
rect 9182 5035 9248 5037
rect 9182 5001 9198 5035
rect 9232 5001 9248 5035
rect 9518 5015 9559 5085
rect 9435 5009 9559 5015
rect 9310 4967 9326 5001
rect 9360 4967 9376 5001
rect 8928 4933 8944 4967
rect 8978 4947 8994 4967
rect 8978 4941 9010 4947
rect 8928 4907 8976 4933
rect 9114 4933 9376 4967
rect 9435 4975 9436 5009
rect 9470 4979 9559 5009
rect 9593 5035 9627 5204
rect 9939 5205 9955 5239
rect 9989 5205 10166 5239
rect 10200 5205 10216 5239
rect 9799 5171 9833 5179
rect 10250 5202 10307 5247
rect 9661 5137 10216 5171
rect 9661 5119 9711 5137
rect 9695 5085 9711 5119
rect 9661 5069 9711 5085
rect 9593 5019 9863 5035
rect 9593 5001 9829 5019
rect 9470 4975 9492 4979
rect 9435 4945 9492 4975
rect 9114 4907 9158 4933
rect 8928 4901 9010 4907
rect 9092 4873 9108 4907
rect 9142 4873 9158 4907
rect 9435 4911 9458 4945
rect 9192 4881 9226 4897
rect 9435 4895 9492 4911
rect 8601 4815 8635 4831
rect 8497 4771 8567 4813
rect 8691 4813 8707 4847
rect 8741 4813 8890 4847
rect 8691 4807 8890 4813
rect 8924 4843 8958 4859
rect 8924 4771 8958 4809
rect 8992 4829 9008 4863
rect 9042 4839 9058 4863
rect 9593 4847 9627 5001
rect 9819 4985 9829 5001
rect 9819 4969 9863 4985
rect 9702 4941 9721 4967
rect 9702 4907 9712 4941
rect 9755 4933 9777 4967
rect 9746 4907 9777 4933
rect 9897 4910 9933 5137
rect 9702 4901 9777 4907
rect 9867 4907 9933 4910
rect 9867 4873 9883 4907
rect 9917 4873 9933 4907
rect 9967 5077 10069 5103
rect 9967 5043 9988 5077
rect 10022 5069 10069 5077
rect 10103 5069 10119 5103
rect 9967 5035 10022 5043
rect 10001 5001 10022 5035
rect 10182 5019 10216 5137
rect 10284 5168 10307 5202
rect 10250 5134 10307 5168
rect 10284 5100 10307 5134
rect 10250 5080 10307 5100
rect 9967 4939 10022 5001
rect 10073 5014 10148 5019
rect 10073 4980 10086 5014
rect 10120 5007 10148 5014
rect 10073 4973 10098 4980
rect 10132 4973 10148 5007
rect 10182 5003 10232 5019
rect 10182 4969 10198 5003
rect 10182 4953 10232 4969
rect 9967 4905 10105 4939
rect 9192 4839 9226 4847
rect 9042 4829 9226 4839
rect 8992 4805 9226 4829
rect 9280 4813 9296 4847
rect 9330 4813 9346 4847
rect 9280 4771 9346 4813
rect 9474 4813 9490 4847
rect 9524 4813 9627 4847
rect 9474 4807 9627 4813
rect 9663 4843 9715 4859
rect 9663 4809 9681 4843
rect 9663 4771 9715 4809
rect 9767 4829 9783 4863
rect 9817 4839 9833 4863
rect 9967 4855 10001 4871
rect 9817 4829 9967 4839
rect 9767 4821 9967 4829
rect 9767 4805 10001 4821
rect 10058 4857 10105 4905
rect 10058 4823 10071 4857
rect 10058 4807 10105 4823
rect 10150 4847 10216 4915
rect 10266 4897 10307 5080
rect 10150 4813 10166 4847
rect 10200 4813 10216 4847
rect 10150 4771 10216 4813
rect 10250 4881 10307 4897
rect 10284 4880 10307 4881
rect 10250 4846 10261 4847
rect 10295 4846 10307 4880
rect 10250 4805 10307 4846
rect 10341 5221 10404 5237
rect 10341 5187 10354 5221
rect 10388 5187 10404 5221
rect 10341 5153 10404 5187
rect 10341 5119 10354 5153
rect 10388 5119 10404 5153
rect 10341 5019 10404 5119
rect 10440 5227 10499 5281
rect 10440 5193 10449 5227
rect 10483 5193 10499 5227
rect 10440 5159 10499 5193
rect 10440 5125 10449 5159
rect 10483 5125 10499 5159
rect 10440 5107 10499 5125
rect 10533 5203 10585 5247
rect 10567 5169 10585 5203
rect 10533 5135 10585 5169
rect 10567 5101 10585 5135
rect 10619 5231 10671 5247
rect 10619 5197 10637 5231
rect 10619 5163 10671 5197
rect 10705 5215 10771 5281
rect 10705 5181 10721 5215
rect 10755 5181 10771 5215
rect 10805 5231 10850 5247
rect 10839 5197 10850 5231
rect 10619 5129 10637 5163
rect 10805 5163 10850 5197
rect 10889 5215 10959 5281
rect 10889 5181 10909 5215
rect 10943 5181 10959 5215
rect 10993 5231 11027 5247
rect 11070 5204 11086 5238
rect 11120 5204 11236 5238
rect 10671 5145 10770 5147
rect 10671 5129 10724 5145
rect 10619 5113 10724 5129
rect 10533 5077 10585 5101
rect 10758 5111 10770 5145
rect 10533 5043 10543 5077
rect 10577 5043 10585 5077
rect 10341 5003 10508 5019
rect 10341 4969 10474 5003
rect 10341 4953 10508 4969
rect 10341 4873 10404 4953
rect 10542 4919 10585 5043
rect 10619 5018 10690 5079
rect 10619 4984 10634 5018
rect 10668 4996 10690 5018
rect 10619 4962 10637 4984
rect 10671 4962 10690 4996
rect 10619 4949 10690 4962
rect 10724 5018 10770 5111
rect 10724 4984 10736 5018
rect 10341 4839 10354 4873
rect 10388 4839 10404 4873
rect 10533 4911 10585 4919
rect 10724 4915 10770 4984
rect 10533 4883 10544 4911
rect 10578 4877 10585 4911
rect 10341 4805 10404 4839
rect 10440 4847 10499 4863
rect 10440 4813 10449 4847
rect 10483 4813 10499 4847
rect 10440 4771 10499 4813
rect 10567 4849 10585 4877
rect 10533 4805 10585 4849
rect 10619 4881 10770 4915
rect 10839 5129 10850 5163
rect 10993 5147 11027 5197
rect 10805 4941 10850 5129
rect 10805 4907 10816 4941
rect 10619 4873 10671 4881
rect 10619 4839 10637 4873
rect 10805 4873 10850 4907
rect 10884 5113 11027 5147
rect 10884 4919 10918 5113
rect 11068 5111 11092 5145
rect 11126 5119 11168 5145
rect 11126 5111 11134 5119
rect 11068 5085 11134 5111
rect 10952 5073 11034 5079
rect 10952 5039 10954 5073
rect 10988 5039 11034 5073
rect 10952 5005 11034 5039
rect 10986 4971 11034 5005
rect 10952 4955 11034 4971
rect 11068 5069 11168 5085
rect 11068 4945 11112 5069
rect 11202 5035 11236 5204
rect 11284 5229 11360 5281
rect 11578 5239 11644 5281
rect 11284 5195 11300 5229
rect 11334 5195 11360 5229
rect 11420 5213 11454 5229
rect 11420 5161 11454 5179
rect 11578 5205 11594 5239
rect 11628 5205 11644 5239
rect 12067 5239 12143 5281
rect 11578 5171 11644 5205
rect 11853 5204 11869 5238
rect 11903 5204 12019 5238
rect 12067 5205 12083 5239
rect 12117 5205 12143 5239
rect 12331 5239 12608 5281
rect 12191 5213 12225 5229
rect 11270 5145 11540 5161
rect 11270 5119 11420 5145
rect 11304 5111 11420 5119
rect 11454 5111 11540 5145
rect 11578 5137 11594 5171
rect 11628 5137 11644 5171
rect 11815 5145 11862 5151
rect 11304 5085 11320 5111
rect 11270 5069 11320 5085
rect 11422 5035 11472 5051
rect 11202 5001 11438 5035
rect 11202 4993 11282 5001
rect 10884 4881 11027 4919
rect 11102 4911 11112 4945
rect 11068 4895 11112 4911
rect 11148 4923 11164 4957
rect 11198 4941 11214 4957
rect 11148 4907 11180 4923
rect 11148 4883 11214 4907
rect 10619 4823 10671 4839
rect 10705 4813 10721 4847
rect 10755 4813 10771 4847
rect 10839 4839 10850 4873
rect 10993 4865 11027 4881
rect 10805 4823 10850 4839
rect 10705 4771 10771 4813
rect 10889 4813 10909 4847
rect 10943 4813 10959 4847
rect 11248 4847 11282 4993
rect 11428 4985 11472 5001
rect 11506 4967 11540 5111
rect 11815 5119 11828 5145
rect 11849 5085 11862 5111
rect 11574 5077 11775 5085
rect 11574 5043 11736 5077
rect 11770 5043 11775 5077
rect 11815 5069 11862 5085
rect 11910 5119 11951 5135
rect 11910 5085 11917 5119
rect 11574 5037 11775 5043
rect 11574 5035 11640 5037
rect 11574 5001 11590 5035
rect 11624 5001 11640 5035
rect 11910 5015 11951 5085
rect 11827 5009 11951 5015
rect 11702 4967 11718 5001
rect 11752 4967 11768 5001
rect 11320 4933 11336 4967
rect 11370 4947 11386 4967
rect 11370 4941 11402 4947
rect 11320 4907 11368 4933
rect 11506 4933 11768 4967
rect 11827 4975 11828 5009
rect 11862 4979 11951 5009
rect 11985 5035 12019 5204
rect 12331 5205 12347 5239
rect 12381 5205 12558 5239
rect 12592 5205 12608 5239
rect 12191 5171 12225 5179
rect 12642 5202 12699 5247
rect 12053 5137 12608 5171
rect 12053 5119 12103 5137
rect 12087 5085 12103 5119
rect 12053 5069 12103 5085
rect 11985 5019 12255 5035
rect 11985 5001 12221 5019
rect 11862 4975 11884 4979
rect 11827 4945 11884 4975
rect 11506 4907 11550 4933
rect 11320 4901 11402 4907
rect 11484 4873 11500 4907
rect 11534 4873 11550 4907
rect 11827 4911 11850 4945
rect 11584 4881 11618 4897
rect 11827 4895 11884 4911
rect 10993 4815 11027 4831
rect 10889 4771 10959 4813
rect 11083 4813 11099 4847
rect 11133 4813 11282 4847
rect 11083 4807 11282 4813
rect 11316 4843 11350 4859
rect 11316 4771 11350 4809
rect 11384 4829 11400 4863
rect 11434 4839 11450 4863
rect 11985 4847 12019 5001
rect 12211 4985 12221 5001
rect 12211 4969 12255 4985
rect 12094 4941 12113 4967
rect 12094 4907 12104 4941
rect 12147 4933 12169 4967
rect 12138 4907 12169 4933
rect 12289 4910 12325 5137
rect 12094 4901 12169 4907
rect 12259 4907 12325 4910
rect 12259 4873 12275 4907
rect 12309 4873 12325 4907
rect 12359 5077 12461 5103
rect 12359 5043 12380 5077
rect 12414 5069 12461 5077
rect 12495 5069 12511 5103
rect 12359 5035 12414 5043
rect 12393 5001 12414 5035
rect 12574 5019 12608 5137
rect 12676 5168 12699 5202
rect 12642 5134 12699 5168
rect 12676 5100 12699 5134
rect 12642 5080 12699 5100
rect 12359 4939 12414 5001
rect 12465 5012 12540 5019
rect 12465 4978 12477 5012
rect 12511 5007 12540 5012
rect 12465 4973 12490 4978
rect 12524 4973 12540 5007
rect 12574 5003 12624 5019
rect 12574 4969 12590 5003
rect 12574 4953 12624 4969
rect 12359 4905 12497 4939
rect 11584 4839 11618 4847
rect 11434 4829 11618 4839
rect 11384 4805 11618 4829
rect 11672 4813 11688 4847
rect 11722 4813 11738 4847
rect 11672 4771 11738 4813
rect 11866 4813 11882 4847
rect 11916 4813 12019 4847
rect 11866 4807 12019 4813
rect 12055 4843 12107 4859
rect 12055 4809 12073 4843
rect 12055 4771 12107 4809
rect 12159 4829 12175 4863
rect 12209 4839 12225 4863
rect 12359 4855 12393 4871
rect 12209 4829 12359 4839
rect 12159 4821 12359 4829
rect 12159 4805 12393 4821
rect 12450 4857 12497 4905
rect 12450 4823 12463 4857
rect 12450 4807 12497 4823
rect 12542 4847 12608 4915
rect 12658 4897 12699 5080
rect 12542 4813 12558 4847
rect 12592 4813 12608 4847
rect 12542 4771 12608 4813
rect 12642 4881 12699 4897
rect 12686 4847 12699 4881
rect 12642 4805 12699 4847
rect 12733 5221 12796 5237
rect 12733 5187 12746 5221
rect 12780 5187 12796 5221
rect 12733 5153 12796 5187
rect 12733 5119 12746 5153
rect 12780 5119 12796 5153
rect 12733 5019 12796 5119
rect 12832 5227 12891 5281
rect 12832 5193 12841 5227
rect 12875 5193 12891 5227
rect 12832 5159 12891 5193
rect 12832 5125 12841 5159
rect 12875 5125 12891 5159
rect 12832 5107 12891 5125
rect 12925 5203 12977 5247
rect 12959 5201 12977 5203
rect 12925 5167 12931 5169
rect 12965 5167 12977 5201
rect 12925 5135 12977 5167
rect 12959 5101 12977 5135
rect 12925 5043 12977 5101
rect 12733 5003 12900 5019
rect 12733 4969 12866 5003
rect 12733 4953 12900 4969
rect 12733 4873 12796 4953
rect 12934 4919 12977 5043
rect 12733 4839 12746 4873
rect 12780 4839 12796 4873
rect 12925 4911 12977 4919
rect 12925 4883 12939 4911
rect 12973 4877 12977 4911
rect 12733 4805 12796 4839
rect 12832 4847 12891 4863
rect 12832 4813 12841 4847
rect 12875 4813 12891 4847
rect 12832 4771 12891 4813
rect 12959 4849 12977 4877
rect 12925 4805 12977 4849
rect 1034 4713 1063 4771
rect 1097 4713 1155 4771
rect 1189 4713 1247 4771
rect 1281 4713 1339 4771
rect 1373 4713 1431 4771
rect 1465 4713 1523 4771
rect 1557 4713 1615 4771
rect 1649 4713 1707 4771
rect 1741 4713 1799 4771
rect 1833 4713 1891 4771
rect 1925 4713 1983 4771
rect 2017 4713 2075 4771
rect 2109 4713 2167 4771
rect 2201 4713 2259 4771
rect 2293 4713 2351 4771
rect 2385 4713 2443 4771
rect 2477 4713 2535 4771
rect 2569 4713 2627 4771
rect 2661 4713 2719 4771
rect 2753 4713 2811 4771
rect 2845 4713 2903 4771
rect 2937 4713 2995 4771
rect 3029 4713 3087 4771
rect 3121 4713 3179 4771
rect 3213 4713 3271 4771
rect 3305 4713 3363 4771
rect 3397 4713 3455 4771
rect 3489 4713 3547 4771
rect 3581 4713 3639 4771
rect 3673 4713 3731 4771
rect 3765 4713 3823 4771
rect 3857 4713 3915 4771
rect 3949 4713 4007 4771
rect 4041 4713 4099 4771
rect 4133 4713 4191 4771
rect 4225 4713 4283 4771
rect 4317 4713 4375 4771
rect 4409 4713 4467 4771
rect 4501 4713 4559 4771
rect 4593 4713 4651 4771
rect 4685 4713 4743 4771
rect 4777 4713 4835 4771
rect 4869 4713 4927 4771
rect 4961 4713 5019 4771
rect 5053 4713 5111 4771
rect 5145 4713 5203 4771
rect 5237 4713 5295 4771
rect 5329 4713 5387 4771
rect 5421 4713 5479 4771
rect 5513 4713 5571 4771
rect 5605 4713 5663 4771
rect 5697 4713 5755 4771
rect 5789 4713 5847 4771
rect 5881 4713 5939 4771
rect 5973 4713 6031 4771
rect 6065 4713 6123 4771
rect 6157 4713 6215 4771
rect 6249 4713 6307 4771
rect 6341 4713 6399 4771
rect 6433 4713 6491 4771
rect 6525 4713 6583 4771
rect 6617 4713 6675 4771
rect 6709 4713 6767 4771
rect 6801 4713 6859 4771
rect 6893 4713 6951 4771
rect 6985 4713 7043 4771
rect 7077 4713 7135 4771
rect 7169 4713 7227 4771
rect 7261 4713 7319 4771
rect 7353 4713 7411 4771
rect 7445 4713 7503 4771
rect 7537 4713 7595 4771
rect 7629 4713 7687 4771
rect 7721 4713 7779 4771
rect 7813 4713 7871 4771
rect 7905 4713 7963 4771
rect 7997 4713 8055 4771
rect 8089 4713 8147 4771
rect 8181 4713 8239 4771
rect 8273 4713 8331 4771
rect 8365 4713 8423 4771
rect 8457 4713 8515 4771
rect 8549 4713 8607 4771
rect 8641 4713 8699 4771
rect 8733 4713 8791 4771
rect 8825 4713 8883 4771
rect 8917 4713 8975 4771
rect 9009 4713 9067 4771
rect 9101 4713 9159 4771
rect 9193 4713 9251 4771
rect 9285 4713 9343 4771
rect 9377 4713 9435 4771
rect 9469 4713 9527 4771
rect 9561 4713 9619 4771
rect 9653 4713 9711 4771
rect 9745 4713 9803 4771
rect 9837 4713 9895 4771
rect 9929 4713 9987 4771
rect 10021 4713 10079 4771
rect 10113 4713 10171 4771
rect 10205 4713 10263 4771
rect 10297 4713 10355 4771
rect 10389 4713 10447 4771
rect 10481 4713 10539 4771
rect 10573 4713 10631 4771
rect 10665 4713 10723 4771
rect 10757 4713 10815 4771
rect 10849 4713 10907 4771
rect 10941 4713 10999 4771
rect 11033 4713 11091 4771
rect 11125 4713 11183 4771
rect 11217 4713 11275 4771
rect 11309 4713 11367 4771
rect 11401 4713 11459 4771
rect 11493 4713 11551 4771
rect 11585 4713 11643 4771
rect 11677 4713 11735 4771
rect 11769 4713 11827 4771
rect 11861 4713 11919 4771
rect 11953 4713 12011 4771
rect 12045 4713 12103 4771
rect 12137 4713 12195 4771
rect 12229 4713 12287 4771
rect 12321 4713 12379 4771
rect 12413 4713 12471 4771
rect 12505 4713 12563 4771
rect 12597 4713 12655 4771
rect 12689 4713 12747 4771
rect 12781 4713 12839 4771
rect 12873 4713 12931 4771
rect 12965 4713 12994 4771
rect 594 4592 623 4650
rect 657 4592 715 4650
rect 749 4592 807 4650
rect 841 4592 899 4650
rect 933 4592 991 4650
rect 1025 4592 1083 4650
rect 1117 4592 1175 4650
rect 1209 4592 1267 4650
rect 1301 4592 1359 4650
rect 1393 4626 1451 4650
rect 1485 4626 1543 4650
rect 1577 4626 1635 4650
rect 1669 4626 1727 4650
rect 1761 4626 1819 4650
rect 1853 4626 1911 4650
rect 1945 4626 2003 4650
rect 2037 4626 2095 4650
rect 2129 4626 2187 4650
rect 2221 4626 2279 4650
rect 1393 4592 1431 4626
rect 1485 4616 1523 4626
rect 1577 4616 1615 4626
rect 1669 4616 1707 4626
rect 1761 4616 1799 4626
rect 1853 4616 1891 4626
rect 1945 4616 1983 4626
rect 2037 4616 2075 4626
rect 2129 4616 2167 4626
rect 2221 4616 2259 4626
rect 2313 4616 2351 4650
rect 2405 4616 2443 4650
rect 1465 4592 1523 4616
rect 1557 4592 1615 4616
rect 1649 4592 1707 4616
rect 1741 4592 1799 4616
rect 1833 4592 1891 4616
rect 1925 4592 1983 4616
rect 2017 4592 2075 4616
rect 2109 4592 2167 4616
rect 2201 4592 2259 4616
rect 2293 4592 2351 4616
rect 2385 4592 2443 4616
rect 2477 4592 2535 4650
rect 2569 4592 2627 4650
rect 2661 4592 2719 4650
rect 2753 4592 2811 4650
rect 2845 4592 2903 4650
rect 2937 4592 2995 4650
rect 3029 4592 3087 4650
rect 3121 4592 3179 4650
rect 3213 4592 3271 4650
rect 3305 4592 3363 4650
rect 3397 4592 3455 4650
rect 3489 4592 3547 4650
rect 3581 4592 3639 4650
rect 3673 4592 3731 4650
rect 3765 4592 3823 4650
rect 3857 4592 3915 4650
rect 3949 4592 4007 4650
rect 4041 4592 4099 4650
rect 4133 4647 4375 4650
rect 4133 4626 4248 4647
rect 4133 4592 4191 4626
rect 4225 4613 4248 4626
rect 4282 4626 4375 4647
rect 4282 4613 4283 4626
rect 4225 4592 4283 4613
rect 4317 4592 4375 4626
rect 4409 4592 4467 4650
rect 4501 4592 4559 4650
rect 4593 4592 4651 4650
rect 4685 4592 4743 4650
rect 4777 4592 4835 4650
rect 4869 4592 4927 4650
rect 4961 4592 5019 4650
rect 5053 4592 5111 4650
rect 5145 4592 5203 4650
rect 5237 4592 5295 4650
rect 5329 4592 5387 4650
rect 5421 4592 5479 4650
rect 5513 4592 5571 4650
rect 5605 4592 5663 4650
rect 5697 4592 5755 4650
rect 5789 4592 5847 4650
rect 5881 4592 5939 4650
rect 5973 4592 6031 4650
rect 6065 4592 6123 4650
rect 6157 4592 6215 4650
rect 6249 4592 6307 4650
rect 6341 4592 6399 4650
rect 6433 4592 6491 4650
rect 6525 4647 6767 4650
rect 6525 4626 6640 4647
rect 6525 4592 6583 4626
rect 6617 4613 6640 4626
rect 6674 4626 6767 4647
rect 6674 4613 6675 4626
rect 6617 4592 6675 4613
rect 6709 4592 6767 4626
rect 6801 4592 6859 4650
rect 6893 4592 6951 4650
rect 6985 4592 7043 4650
rect 7077 4592 7135 4650
rect 7169 4592 7227 4650
rect 7261 4592 7319 4650
rect 7353 4592 7411 4650
rect 7445 4592 7503 4650
rect 7537 4592 7595 4650
rect 7629 4592 7687 4650
rect 7721 4592 7779 4650
rect 7813 4592 7871 4650
rect 7905 4592 7963 4650
rect 7997 4592 8055 4650
rect 8089 4592 8147 4650
rect 8181 4592 8239 4650
rect 8273 4592 8331 4650
rect 8365 4592 8423 4650
rect 8457 4592 8515 4650
rect 8549 4592 8607 4650
rect 8641 4592 8699 4650
rect 8733 4592 8791 4650
rect 8825 4592 8883 4650
rect 8917 4647 9159 4650
rect 8917 4626 9032 4647
rect 8917 4592 8975 4626
rect 9009 4613 9032 4626
rect 9066 4626 9159 4647
rect 9066 4613 9067 4626
rect 9009 4592 9067 4613
rect 9101 4592 9159 4626
rect 9193 4592 9251 4650
rect 9285 4592 9343 4650
rect 9377 4592 9435 4650
rect 9469 4592 9527 4650
rect 9561 4592 9619 4650
rect 9653 4592 9711 4650
rect 9745 4592 9803 4650
rect 9837 4592 9895 4650
rect 9929 4592 9987 4650
rect 10021 4592 10079 4650
rect 10113 4592 10171 4650
rect 10205 4592 10263 4650
rect 10297 4592 10355 4650
rect 10389 4592 10447 4650
rect 10481 4592 10539 4650
rect 10573 4592 10631 4650
rect 10665 4592 10723 4650
rect 10757 4592 10815 4650
rect 10849 4592 10907 4650
rect 10941 4592 10999 4650
rect 11033 4592 11091 4650
rect 11125 4592 11183 4650
rect 11217 4592 11275 4650
rect 11309 4647 11551 4650
rect 11309 4626 11424 4647
rect 11309 4592 11367 4626
rect 11401 4613 11424 4626
rect 11458 4626 11551 4647
rect 11458 4613 11459 4626
rect 11401 4592 11459 4613
rect 11493 4592 11551 4626
rect 11585 4592 11643 4650
rect 11677 4592 11735 4650
rect 11769 4592 11827 4650
rect 11861 4592 11919 4650
rect 11953 4592 12011 4650
rect 12045 4592 12103 4650
rect 12137 4592 12195 4650
rect 12229 4592 12287 4650
rect 12321 4592 12379 4650
rect 12413 4592 12471 4650
rect 12505 4592 12563 4650
rect 12597 4592 12655 4650
rect 12689 4592 12747 4650
rect 12781 4592 12839 4650
rect 12873 4592 12931 4650
rect 12965 4592 12994 4650
rect 627 4542 663 4558
rect 627 4508 629 4542
rect 627 4474 663 4508
rect 627 4440 629 4474
rect 699 4542 765 4592
rect 699 4508 715 4542
rect 749 4508 765 4542
rect 699 4474 765 4508
rect 699 4440 715 4474
rect 749 4440 765 4474
rect 799 4542 853 4558
rect 799 4508 801 4542
rect 835 4508 853 4542
rect 799 4461 853 4508
rect 627 4406 663 4440
rect 799 4427 801 4461
rect 835 4427 853 4461
rect 627 4372 762 4406
rect 799 4377 853 4427
rect 728 4343 762 4372
rect 615 4318 683 4336
rect 615 4284 625 4318
rect 659 4314 683 4318
rect 615 4280 631 4284
rect 665 4280 683 4314
rect 615 4262 683 4280
rect 728 4327 783 4343
rect 728 4293 749 4327
rect 728 4277 783 4293
rect 817 4327 853 4377
rect 889 4544 955 4558
rect 889 4510 905 4544
rect 939 4510 955 4544
rect 889 4476 955 4510
rect 889 4442 905 4476
rect 939 4442 955 4476
rect 889 4408 955 4442
rect 989 4550 1037 4592
rect 1023 4516 1037 4550
rect 989 4482 1037 4516
rect 1023 4448 1037 4482
rect 989 4432 1037 4448
rect 1073 4528 1107 4558
rect 1073 4433 1107 4494
rect 889 4374 905 4408
rect 939 4396 955 4408
rect 1141 4550 1207 4592
rect 1141 4516 1157 4550
rect 1191 4516 1207 4550
rect 1141 4482 1207 4516
rect 1141 4448 1157 4482
rect 1191 4448 1207 4482
rect 1141 4432 1207 4448
rect 1241 4528 1275 4558
rect 1241 4433 1275 4494
rect 939 4374 1032 4396
rect 889 4362 1032 4374
rect 888 4327 964 4328
rect 817 4314 964 4327
rect 817 4282 914 4314
rect 728 4226 762 4277
rect 629 4192 762 4226
rect 817 4217 853 4282
rect 888 4280 914 4282
rect 948 4280 964 4314
rect 998 4314 1032 4362
rect 1073 4388 1107 4399
rect 1241 4388 1275 4399
rect 1073 4354 1275 4388
rect 1309 4550 1375 4592
rect 1309 4516 1325 4550
rect 1359 4516 1375 4550
rect 1309 4482 1375 4516
rect 1309 4448 1325 4482
rect 1359 4448 1375 4482
rect 1309 4414 1375 4448
rect 1309 4380 1325 4414
rect 1359 4380 1375 4414
rect 1309 4362 1375 4380
rect 1437 4550 1471 4592
rect 1437 4482 1471 4516
rect 1437 4414 1471 4448
rect 1437 4354 1471 4380
rect 1505 4544 1571 4558
rect 1505 4510 1521 4544
rect 1555 4510 1571 4544
rect 1505 4476 1571 4510
rect 1505 4442 1521 4476
rect 1555 4442 1571 4476
rect 1505 4408 1571 4442
rect 1605 4550 1639 4592
rect 1605 4482 1639 4516
rect 1605 4432 1639 4448
rect 1673 4544 1739 4558
rect 1673 4510 1689 4544
rect 1723 4510 1739 4544
rect 1673 4476 1739 4510
rect 1673 4442 1689 4476
rect 1723 4442 1739 4476
rect 1505 4374 1521 4408
rect 1555 4388 1571 4408
rect 1673 4408 1739 4442
rect 1773 4550 1807 4592
rect 1773 4482 1807 4516
rect 1773 4432 1807 4448
rect 1841 4544 1907 4558
rect 1841 4510 1857 4544
rect 1891 4510 1907 4544
rect 1841 4476 1907 4510
rect 1841 4442 1857 4476
rect 1891 4442 1907 4476
rect 1673 4388 1689 4408
rect 1555 4374 1689 4388
rect 1723 4388 1739 4408
rect 1841 4408 1907 4442
rect 1941 4550 1975 4592
rect 1941 4482 1975 4516
rect 1941 4432 1975 4448
rect 2009 4544 2075 4558
rect 2009 4510 2025 4544
rect 2059 4510 2075 4544
rect 2009 4476 2075 4510
rect 2009 4442 2025 4476
rect 2059 4442 2075 4476
rect 1841 4388 1857 4408
rect 1723 4374 1857 4388
rect 1891 4388 1907 4408
rect 2009 4408 2075 4442
rect 2109 4550 2143 4592
rect 2109 4482 2143 4516
rect 2109 4432 2143 4448
rect 2177 4544 2243 4558
rect 2177 4510 2193 4544
rect 2227 4510 2243 4544
rect 2177 4476 2243 4510
rect 2177 4442 2193 4476
rect 2227 4442 2243 4476
rect 1891 4374 1975 4388
rect 1505 4354 1975 4374
rect 2009 4374 2025 4408
rect 2059 4388 2075 4408
rect 2177 4408 2243 4442
rect 2277 4550 2311 4592
rect 2277 4482 2311 4516
rect 2277 4432 2311 4448
rect 2345 4544 2411 4558
rect 2345 4510 2361 4544
rect 2395 4510 2411 4544
rect 2345 4476 2411 4510
rect 2345 4442 2361 4476
rect 2395 4442 2411 4476
rect 2177 4388 2193 4408
rect 2059 4374 2193 4388
rect 2227 4388 2243 4408
rect 2345 4408 2411 4442
rect 2445 4550 2479 4592
rect 2445 4482 2479 4516
rect 2445 4432 2479 4448
rect 2513 4544 2579 4558
rect 2513 4510 2529 4544
rect 2563 4510 2579 4544
rect 2513 4488 2579 4510
rect 2513 4476 2538 4488
rect 2513 4442 2529 4476
rect 2572 4454 2579 4488
rect 2563 4442 2579 4454
rect 2345 4388 2361 4408
rect 2227 4374 2361 4388
rect 2395 4388 2411 4408
rect 2513 4408 2579 4442
rect 2613 4550 2647 4592
rect 2613 4482 2647 4516
rect 2613 4432 2647 4448
rect 2681 4544 2747 4558
rect 2681 4510 2697 4544
rect 2731 4510 2747 4544
rect 2681 4476 2747 4510
rect 2681 4442 2697 4476
rect 2731 4442 2747 4476
rect 2513 4388 2529 4408
rect 2395 4374 2529 4388
rect 2563 4388 2579 4408
rect 2681 4408 2747 4442
rect 2781 4550 2815 4592
rect 2781 4482 2815 4516
rect 2781 4432 2815 4448
rect 2849 4544 2915 4558
rect 2849 4510 2865 4544
rect 2899 4510 2915 4544
rect 2849 4476 2915 4510
rect 2849 4442 2865 4476
rect 2899 4442 2915 4476
rect 2681 4388 2697 4408
rect 2563 4374 2697 4388
rect 2731 4388 2747 4408
rect 2849 4408 2915 4442
rect 2949 4550 2983 4592
rect 2949 4482 2983 4516
rect 2949 4432 2983 4448
rect 3017 4544 3083 4558
rect 3017 4510 3033 4544
rect 3067 4510 3083 4544
rect 3017 4476 3083 4510
rect 3017 4442 3033 4476
rect 3067 4442 3083 4476
rect 2849 4388 2865 4408
rect 2731 4374 2865 4388
rect 2899 4388 2915 4408
rect 3017 4408 3083 4442
rect 3117 4550 3151 4592
rect 3117 4482 3151 4516
rect 3117 4432 3151 4448
rect 3185 4544 3251 4558
rect 3185 4510 3201 4544
rect 3235 4510 3251 4544
rect 3185 4476 3251 4510
rect 3185 4442 3201 4476
rect 3235 4442 3251 4476
rect 3017 4388 3033 4408
rect 2899 4374 3033 4388
rect 3067 4388 3083 4408
rect 3185 4408 3251 4442
rect 3285 4550 3319 4592
rect 3285 4482 3319 4516
rect 3285 4432 3319 4448
rect 3185 4388 3201 4408
rect 3067 4374 3201 4388
rect 3235 4388 3251 4408
rect 3354 4388 3409 4537
rect 3235 4374 3409 4388
rect 2009 4354 3409 4374
rect 1176 4320 1275 4354
rect 1940 4320 1975 4354
rect 1176 4314 1899 4320
rect 998 4280 1048 4314
rect 1082 4280 1098 4314
rect 1176 4280 1505 4314
rect 1539 4280 1573 4314
rect 1607 4280 1641 4314
rect 1675 4280 1709 4314
rect 1743 4280 1777 4314
rect 1811 4280 1845 4314
rect 1879 4280 1899 4314
rect 1940 4314 3284 4320
rect 1940 4280 2005 4314
rect 2039 4280 2073 4314
rect 2107 4280 2141 4314
rect 2175 4280 2209 4314
rect 2243 4280 2277 4314
rect 2311 4280 2345 4314
rect 2379 4280 2413 4314
rect 2447 4280 2481 4314
rect 2515 4280 2549 4314
rect 2583 4280 2617 4314
rect 2651 4280 2685 4314
rect 2719 4280 2753 4314
rect 2787 4280 2821 4314
rect 2855 4280 2889 4314
rect 2923 4280 2957 4314
rect 2991 4280 3025 4314
rect 3059 4280 3093 4314
rect 3127 4280 3161 4314
rect 3195 4280 3229 4314
rect 3263 4280 3284 4314
rect 998 4246 1032 4280
rect 1176 4246 1275 4280
rect 1940 4246 1975 4280
rect 3333 4246 3409 4354
rect 629 4171 663 4192
rect 801 4188 853 4217
rect 629 4116 663 4137
rect 699 4124 715 4158
rect 749 4124 765 4158
rect 699 4082 765 4124
rect 835 4154 853 4188
rect 801 4116 853 4154
rect 905 4212 1032 4246
rect 1073 4212 1275 4246
rect 905 4194 939 4212
rect 1073 4194 1107 4212
rect 905 4116 939 4160
rect 975 4162 1023 4178
rect 975 4128 989 4162
rect 975 4082 1023 4128
rect 1241 4194 1275 4212
rect 1073 4116 1107 4160
rect 1141 4162 1207 4178
rect 1141 4128 1157 4162
rect 1191 4128 1207 4162
rect 1141 4082 1207 4128
rect 1241 4116 1275 4160
rect 1309 4226 1375 4242
rect 1309 4192 1325 4226
rect 1359 4192 1375 4226
rect 1309 4158 1375 4192
rect 1309 4124 1325 4158
rect 1359 4124 1375 4158
rect 1309 4082 1375 4124
rect 1437 4230 1471 4246
rect 1437 4162 1471 4196
rect 1437 4082 1471 4128
rect 1505 4230 1975 4246
rect 1505 4196 1521 4230
rect 1555 4212 1689 4230
rect 1555 4196 1571 4212
rect 1505 4162 1571 4196
rect 1673 4196 1689 4212
rect 1723 4212 1857 4230
rect 1723 4196 1739 4212
rect 1505 4128 1521 4162
rect 1555 4128 1571 4162
rect 1505 4117 1571 4128
rect 1605 4162 1639 4178
rect 1605 4082 1639 4128
rect 1673 4162 1739 4196
rect 1841 4196 1857 4212
rect 1891 4212 1975 4230
rect 2009 4230 3409 4246
rect 1891 4196 1907 4212
rect 1673 4128 1689 4162
rect 1723 4128 1739 4162
rect 1673 4117 1739 4128
rect 1773 4162 1807 4178
rect 1773 4082 1807 4128
rect 1841 4162 1907 4196
rect 2009 4196 2025 4230
rect 2059 4212 2193 4230
rect 2059 4196 2075 4212
rect 1841 4128 1857 4162
rect 1891 4128 1907 4162
rect 1841 4117 1907 4128
rect 1941 4162 1975 4178
rect 1941 4082 1975 4128
rect 2009 4162 2075 4196
rect 2177 4196 2193 4212
rect 2227 4212 2361 4230
rect 2227 4196 2243 4212
rect 2009 4128 2025 4162
rect 2059 4128 2075 4162
rect 2009 4117 2075 4128
rect 2109 4162 2143 4178
rect 2009 4116 2059 4117
rect 2109 4082 2143 4128
rect 2177 4162 2243 4196
rect 2345 4196 2361 4212
rect 2395 4212 2529 4230
rect 2395 4196 2411 4212
rect 2177 4128 2193 4162
rect 2227 4128 2243 4162
rect 2177 4117 2243 4128
rect 2277 4162 2311 4178
rect 2193 4116 2227 4117
rect 2277 4082 2311 4128
rect 2345 4162 2411 4196
rect 2513 4196 2529 4212
rect 2563 4212 2697 4230
rect 2563 4196 2579 4212
rect 2345 4128 2361 4162
rect 2395 4128 2411 4162
rect 2345 4117 2411 4128
rect 2445 4162 2479 4178
rect 2361 4116 2395 4117
rect 2445 4082 2479 4128
rect 2513 4162 2579 4196
rect 2681 4196 2697 4212
rect 2731 4212 2865 4230
rect 2731 4196 2747 4212
rect 2513 4128 2529 4162
rect 2563 4128 2579 4162
rect 2513 4117 2579 4128
rect 2613 4162 2647 4178
rect 2613 4082 2647 4128
rect 2681 4162 2747 4196
rect 2849 4196 2865 4212
rect 2899 4212 3033 4230
rect 2899 4196 2915 4212
rect 2681 4128 2697 4162
rect 2731 4128 2747 4162
rect 2681 4117 2747 4128
rect 2781 4162 2815 4178
rect 2781 4082 2815 4128
rect 2849 4162 2915 4196
rect 3017 4196 3033 4212
rect 3067 4212 3201 4230
rect 3067 4196 3083 4212
rect 2849 4128 2865 4162
rect 2899 4128 2915 4162
rect 2849 4117 2915 4128
rect 2949 4162 2983 4178
rect 2949 4082 2983 4128
rect 3017 4162 3083 4196
rect 3185 4196 3201 4212
rect 3235 4212 3409 4230
rect 3235 4196 3251 4212
rect 3017 4128 3033 4162
rect 3067 4128 3083 4162
rect 3017 4117 3083 4128
rect 3117 4162 3151 4178
rect 3117 4082 3151 4128
rect 3185 4162 3251 4196
rect 3354 4187 3409 4212
rect 3185 4128 3201 4162
rect 3235 4128 3251 4162
rect 3185 4117 3251 4128
rect 3285 4162 3319 4178
rect 3354 4153 3366 4187
rect 3400 4153 3409 4187
rect 3354 4138 3409 4153
rect 3443 4524 3495 4558
rect 3443 4490 3452 4524
rect 3486 4514 3495 4524
rect 3443 4480 3461 4490
rect 3443 4446 3495 4480
rect 3443 4412 3461 4446
rect 3529 4538 3588 4592
rect 3529 4504 3545 4538
rect 3579 4504 3588 4538
rect 3529 4470 3588 4504
rect 3529 4436 3545 4470
rect 3579 4436 3588 4470
rect 3529 4418 3588 4436
rect 3624 4532 3687 4548
rect 3624 4498 3640 4532
rect 3674 4498 3687 4532
rect 3624 4464 3687 4498
rect 3624 4430 3640 4464
rect 3674 4430 3687 4464
rect 3443 4354 3495 4412
rect 3443 4230 3486 4354
rect 3624 4330 3687 4430
rect 3520 4314 3687 4330
rect 3554 4280 3687 4314
rect 3520 4264 3687 4280
rect 3443 4194 3495 4230
rect 3443 4160 3461 4194
rect 3624 4184 3687 4264
rect 3285 4082 3319 4128
rect 3443 4116 3495 4160
rect 3529 4158 3588 4174
rect 3529 4124 3545 4158
rect 3579 4124 3588 4158
rect 3529 4082 3588 4124
rect 3624 4150 3640 4184
rect 3674 4150 3687 4184
rect 3624 4116 3687 4150
rect 3721 4513 3778 4558
rect 3812 4550 4089 4592
rect 3812 4516 3828 4550
rect 3862 4516 4039 4550
rect 4073 4516 4089 4550
rect 4277 4550 4353 4592
rect 4195 4524 4229 4540
rect 3721 4479 3744 4513
rect 4277 4516 4303 4550
rect 4337 4516 4353 4550
rect 4776 4550 4842 4592
rect 4195 4482 4229 4490
rect 4401 4515 4517 4549
rect 4551 4515 4567 4549
rect 4776 4516 4792 4550
rect 4826 4516 4842 4550
rect 5060 4540 5136 4592
rect 3721 4445 3778 4479
rect 3721 4411 3744 4445
rect 3721 4391 3778 4411
rect 3812 4448 4367 4482
rect 3721 4208 3762 4391
rect 3812 4330 3846 4448
rect 3909 4380 3925 4414
rect 3959 4388 4061 4414
rect 3959 4380 4006 4388
rect 4040 4354 4061 4388
rect 4006 4346 4061 4354
rect 3796 4314 3846 4330
rect 3830 4280 3846 4314
rect 3880 4322 3955 4330
rect 3880 4318 3898 4322
rect 3880 4284 3896 4318
rect 3932 4288 3955 4322
rect 3930 4284 3955 4288
rect 4006 4312 4027 4346
rect 3796 4264 3846 4280
rect 4006 4250 4061 4312
rect 3721 4192 3778 4208
rect 3721 4158 3744 4192
rect 3721 4116 3778 4158
rect 3812 4158 3878 4226
rect 3812 4124 3828 4158
rect 3862 4124 3878 4158
rect 3812 4082 3878 4124
rect 3923 4216 4061 4250
rect 4095 4221 4131 4448
rect 4317 4430 4367 4448
rect 4317 4396 4333 4430
rect 4317 4380 4367 4396
rect 4401 4346 4435 4515
rect 4776 4482 4842 4516
rect 4558 4456 4605 4462
rect 4165 4330 4435 4346
rect 4199 4312 4435 4330
rect 4199 4296 4209 4312
rect 4165 4280 4209 4296
rect 4251 4244 4273 4278
rect 4307 4252 4326 4278
rect 4095 4218 4161 4221
rect 3923 4168 3970 4216
rect 4095 4184 4111 4218
rect 4145 4184 4161 4218
rect 4251 4218 4282 4244
rect 4316 4218 4326 4252
rect 4251 4212 4326 4218
rect 3957 4134 3970 4168
rect 3923 4118 3970 4134
rect 4027 4166 4061 4182
rect 4195 4150 4211 4174
rect 4061 4140 4211 4150
rect 4245 4140 4261 4174
rect 4061 4132 4261 4140
rect 4027 4116 4261 4132
rect 4313 4154 4365 4170
rect 4347 4120 4365 4154
rect 4313 4082 4365 4120
rect 4401 4158 4435 4312
rect 4469 4430 4510 4446
rect 4503 4396 4510 4430
rect 4469 4326 4510 4396
rect 4592 4430 4605 4456
rect 4776 4448 4792 4482
rect 4826 4448 4842 4482
rect 4966 4524 5000 4540
rect 5060 4506 5086 4540
rect 5120 4506 5136 4540
rect 5184 4515 5300 4549
rect 5334 4515 5350 4549
rect 5393 4542 5427 4558
rect 4966 4472 5000 4490
rect 4880 4456 5150 4472
rect 4558 4396 4571 4422
rect 4880 4422 4966 4456
rect 5000 4430 5150 4456
rect 5000 4422 5116 4430
rect 4558 4380 4605 4396
rect 4645 4388 4846 4396
rect 4645 4354 4650 4388
rect 4684 4354 4846 4388
rect 4645 4348 4846 4354
rect 4780 4346 4846 4348
rect 4469 4320 4593 4326
rect 4469 4290 4558 4320
rect 4536 4286 4558 4290
rect 4592 4286 4593 4320
rect 4780 4312 4796 4346
rect 4830 4312 4846 4346
rect 4536 4256 4593 4286
rect 4570 4222 4593 4256
rect 4652 4278 4668 4312
rect 4702 4278 4718 4312
rect 4880 4278 4914 4422
rect 5100 4396 5116 4422
rect 5100 4380 5150 4396
rect 4948 4346 4998 4362
rect 5184 4346 5218 4515
rect 5393 4458 5427 4508
rect 5461 4526 5531 4592
rect 5461 4492 5477 4526
rect 5511 4492 5531 4526
rect 5570 4542 5615 4558
rect 5570 4508 5581 4542
rect 5570 4474 5615 4508
rect 5649 4526 5715 4592
rect 5649 4492 5665 4526
rect 5699 4492 5715 4526
rect 5749 4542 5801 4558
rect 5783 4508 5801 4542
rect 5252 4430 5294 4456
rect 5286 4422 5294 4430
rect 5328 4422 5352 4456
rect 5393 4424 5536 4458
rect 5286 4396 5352 4422
rect 5252 4380 5352 4396
rect 4982 4312 5218 4346
rect 4948 4296 4992 4312
rect 5138 4304 5218 4312
rect 4652 4244 4914 4278
rect 5034 4258 5050 4278
rect 4536 4206 4593 4222
rect 4870 4218 4914 4244
rect 5018 4252 5050 4258
rect 5084 4244 5100 4278
rect 5052 4218 5100 4244
rect 4802 4192 4836 4208
rect 4870 4184 4886 4218
rect 4920 4184 4936 4218
rect 5018 4212 5100 4218
rect 4401 4124 4504 4158
rect 4538 4124 4554 4158
rect 4401 4118 4554 4124
rect 4682 4124 4698 4158
rect 4732 4124 4748 4158
rect 4682 4082 4748 4124
rect 4802 4150 4836 4158
rect 4970 4150 4986 4174
rect 4802 4140 4986 4150
rect 5020 4140 5036 4174
rect 4802 4116 5036 4140
rect 5070 4154 5104 4170
rect 5070 4082 5104 4120
rect 5138 4158 5172 4304
rect 5206 4252 5222 4268
rect 5256 4234 5272 4268
rect 5240 4218 5272 4234
rect 5206 4194 5272 4218
rect 5308 4256 5352 4380
rect 5386 4386 5468 4390
rect 5386 4352 5430 4386
rect 5464 4352 5468 4386
rect 5386 4316 5468 4352
rect 5386 4282 5434 4316
rect 5386 4266 5468 4282
rect 5308 4222 5318 4256
rect 5502 4230 5536 4424
rect 5308 4206 5352 4222
rect 5393 4192 5536 4230
rect 5570 4440 5581 4474
rect 5749 4474 5801 4508
rect 5570 4252 5615 4440
rect 5604 4218 5615 4252
rect 5393 4176 5427 4192
rect 5138 4124 5287 4158
rect 5321 4124 5337 4158
rect 5570 4184 5615 4218
rect 5650 4456 5749 4458
rect 5650 4422 5662 4456
rect 5696 4440 5749 4456
rect 5783 4440 5801 4474
rect 5696 4424 5801 4440
rect 5835 4514 5887 4558
rect 5835 4480 5853 4514
rect 5835 4446 5887 4480
rect 5650 4329 5696 4422
rect 5835 4412 5853 4446
rect 5921 4538 5980 4592
rect 5921 4504 5937 4538
rect 5971 4504 5980 4538
rect 5921 4470 5980 4504
rect 5921 4436 5937 4470
rect 5971 4436 5980 4470
rect 5921 4418 5980 4436
rect 6016 4532 6079 4548
rect 6016 4498 6032 4532
rect 6066 4498 6079 4532
rect 6016 4464 6079 4498
rect 6016 4430 6032 4464
rect 6066 4430 6079 4464
rect 5835 4390 5887 4412
rect 5684 4295 5696 4329
rect 5650 4226 5696 4295
rect 5730 4329 5801 4390
rect 5730 4301 5752 4329
rect 5730 4267 5750 4301
rect 5786 4295 5801 4329
rect 5784 4267 5801 4295
rect 5730 4260 5801 4267
rect 5835 4356 5841 4390
rect 5875 4356 5887 4390
rect 5835 4354 5887 4356
rect 5835 4230 5878 4354
rect 6016 4330 6079 4430
rect 5912 4314 6079 4330
rect 5946 4280 6079 4314
rect 5912 4264 6079 4280
rect 5650 4192 5801 4226
rect 5393 4126 5427 4142
rect 5138 4118 5337 4124
rect 5461 4124 5477 4158
rect 5511 4124 5531 4158
rect 5570 4150 5581 4184
rect 5749 4184 5801 4192
rect 5570 4134 5615 4150
rect 5461 4082 5531 4124
rect 5649 4124 5665 4158
rect 5699 4124 5715 4158
rect 5783 4150 5801 4184
rect 5749 4134 5801 4150
rect 5835 4222 5887 4230
rect 5835 4188 5845 4222
rect 5879 4194 5887 4222
rect 5835 4160 5853 4188
rect 6016 4184 6079 4264
rect 5649 4082 5715 4124
rect 5835 4116 5887 4160
rect 5921 4158 5980 4174
rect 5921 4124 5937 4158
rect 5971 4124 5980 4158
rect 5921 4082 5980 4124
rect 6016 4150 6032 4184
rect 6066 4150 6079 4184
rect 6016 4116 6079 4150
rect 6113 4513 6170 4558
rect 6204 4550 6481 4592
rect 6204 4516 6220 4550
rect 6254 4516 6431 4550
rect 6465 4516 6481 4550
rect 6669 4550 6745 4592
rect 6587 4524 6621 4540
rect 6113 4479 6136 4513
rect 6669 4516 6695 4550
rect 6729 4516 6745 4550
rect 7168 4550 7234 4592
rect 6587 4482 6621 4490
rect 6793 4515 6909 4549
rect 6943 4515 6959 4549
rect 7168 4516 7184 4550
rect 7218 4516 7234 4550
rect 7452 4540 7528 4592
rect 6113 4445 6170 4479
rect 6113 4411 6136 4445
rect 6113 4391 6170 4411
rect 6204 4448 6759 4482
rect 6113 4208 6154 4391
rect 6204 4330 6238 4448
rect 6301 4380 6317 4414
rect 6351 4388 6453 4414
rect 6351 4380 6398 4388
rect 6432 4354 6453 4388
rect 6398 4346 6453 4354
rect 6188 4314 6238 4330
rect 6222 4280 6238 4314
rect 6272 4324 6347 4330
rect 6272 4318 6292 4324
rect 6272 4284 6288 4318
rect 6326 4290 6347 4324
rect 6322 4284 6347 4290
rect 6398 4312 6419 4346
rect 6188 4264 6238 4280
rect 6398 4250 6453 4312
rect 6113 4192 6170 4208
rect 6113 4183 6136 4192
rect 6113 4149 6131 4183
rect 6165 4149 6170 4158
rect 6113 4116 6170 4149
rect 6204 4158 6270 4226
rect 6204 4124 6220 4158
rect 6254 4124 6270 4158
rect 6204 4082 6270 4124
rect 6315 4216 6453 4250
rect 6487 4221 6523 4448
rect 6709 4430 6759 4448
rect 6709 4396 6725 4430
rect 6709 4380 6759 4396
rect 6793 4346 6827 4515
rect 7168 4482 7234 4516
rect 6950 4456 6997 4462
rect 6557 4330 6827 4346
rect 6591 4312 6827 4330
rect 6591 4296 6601 4312
rect 6557 4280 6601 4296
rect 6643 4244 6665 4278
rect 6699 4252 6718 4278
rect 6487 4218 6553 4221
rect 6315 4168 6362 4216
rect 6487 4184 6503 4218
rect 6537 4184 6553 4218
rect 6643 4218 6674 4244
rect 6708 4218 6718 4252
rect 6643 4212 6718 4218
rect 6349 4134 6362 4168
rect 6315 4118 6362 4134
rect 6419 4166 6453 4182
rect 6587 4150 6603 4174
rect 6453 4140 6603 4150
rect 6637 4140 6653 4174
rect 6453 4132 6653 4140
rect 6419 4116 6653 4132
rect 6705 4154 6757 4170
rect 6739 4120 6757 4154
rect 6705 4082 6757 4120
rect 6793 4158 6827 4312
rect 6861 4430 6902 4446
rect 6895 4396 6902 4430
rect 6861 4326 6902 4396
rect 6984 4430 6997 4456
rect 7168 4448 7184 4482
rect 7218 4448 7234 4482
rect 7358 4524 7392 4540
rect 7452 4506 7478 4540
rect 7512 4506 7528 4540
rect 7576 4515 7692 4549
rect 7726 4515 7742 4549
rect 7785 4542 7819 4558
rect 7358 4472 7392 4490
rect 7272 4456 7542 4472
rect 6950 4396 6963 4422
rect 7272 4422 7358 4456
rect 7392 4430 7542 4456
rect 7392 4422 7508 4430
rect 6950 4380 6997 4396
rect 7037 4388 7238 4396
rect 7037 4354 7042 4388
rect 7076 4354 7238 4388
rect 7037 4348 7238 4354
rect 7172 4346 7238 4348
rect 6861 4320 6985 4326
rect 6861 4290 6950 4320
rect 6928 4286 6950 4290
rect 6984 4286 6985 4320
rect 7172 4312 7188 4346
rect 7222 4312 7238 4346
rect 6928 4256 6985 4286
rect 6962 4222 6985 4256
rect 7044 4278 7060 4312
rect 7094 4278 7110 4312
rect 7272 4278 7306 4422
rect 7492 4396 7508 4422
rect 7492 4380 7542 4396
rect 7340 4346 7390 4362
rect 7576 4346 7610 4515
rect 7785 4458 7819 4508
rect 7853 4526 7923 4592
rect 7853 4492 7869 4526
rect 7903 4492 7923 4526
rect 7962 4542 8007 4558
rect 7962 4508 7973 4542
rect 7962 4474 8007 4508
rect 8041 4526 8107 4592
rect 8041 4492 8057 4526
rect 8091 4492 8107 4526
rect 8141 4542 8193 4558
rect 8175 4508 8193 4542
rect 7644 4430 7686 4456
rect 7678 4422 7686 4430
rect 7720 4422 7744 4456
rect 7785 4424 7928 4458
rect 7678 4396 7744 4422
rect 7644 4380 7744 4396
rect 7374 4312 7610 4346
rect 7340 4296 7384 4312
rect 7530 4304 7610 4312
rect 7044 4244 7306 4278
rect 7426 4258 7442 4278
rect 6928 4206 6985 4222
rect 7262 4218 7306 4244
rect 7410 4252 7442 4258
rect 7476 4244 7492 4278
rect 7444 4218 7492 4244
rect 7194 4192 7228 4208
rect 7262 4184 7278 4218
rect 7312 4184 7328 4218
rect 7410 4212 7492 4218
rect 6793 4124 6896 4158
rect 6930 4124 6946 4158
rect 6793 4118 6946 4124
rect 7074 4124 7090 4158
rect 7124 4124 7140 4158
rect 7074 4082 7140 4124
rect 7194 4150 7228 4158
rect 7362 4150 7378 4174
rect 7194 4140 7378 4150
rect 7412 4140 7428 4174
rect 7194 4116 7428 4140
rect 7462 4154 7496 4170
rect 7462 4082 7496 4120
rect 7530 4158 7564 4304
rect 7598 4252 7614 4268
rect 7648 4234 7664 4268
rect 7632 4218 7664 4234
rect 7598 4194 7664 4218
rect 7700 4256 7744 4380
rect 7778 4386 7860 4390
rect 7778 4352 7822 4386
rect 7856 4352 7860 4386
rect 7778 4316 7860 4352
rect 7778 4282 7826 4316
rect 7778 4266 7860 4282
rect 7700 4222 7710 4256
rect 7894 4230 7928 4424
rect 7700 4206 7744 4222
rect 7785 4192 7928 4230
rect 7962 4440 7973 4474
rect 8141 4474 8193 4508
rect 7962 4252 8007 4440
rect 7996 4218 8007 4252
rect 7785 4176 7819 4192
rect 7530 4124 7679 4158
rect 7713 4124 7729 4158
rect 7962 4184 8007 4218
rect 8042 4456 8141 4458
rect 8042 4422 8054 4456
rect 8088 4440 8141 4456
rect 8175 4440 8193 4474
rect 8088 4424 8193 4440
rect 8227 4514 8279 4558
rect 8227 4480 8245 4514
rect 8227 4446 8279 4480
rect 8042 4329 8088 4422
rect 8227 4412 8245 4446
rect 8313 4538 8372 4592
rect 8313 4504 8329 4538
rect 8363 4504 8372 4538
rect 8313 4470 8372 4504
rect 8313 4436 8329 4470
rect 8363 4436 8372 4470
rect 8313 4418 8372 4436
rect 8408 4532 8471 4548
rect 8408 4498 8424 4532
rect 8458 4498 8471 4532
rect 8408 4464 8471 4498
rect 8408 4430 8424 4464
rect 8458 4430 8471 4464
rect 8227 4390 8279 4412
rect 8076 4295 8088 4329
rect 8042 4226 8088 4295
rect 8122 4329 8193 4390
rect 8122 4295 8144 4329
rect 8178 4302 8193 4329
rect 8122 4268 8147 4295
rect 8181 4268 8193 4302
rect 8122 4260 8193 4268
rect 8227 4356 8233 4390
rect 8267 4356 8279 4390
rect 8227 4354 8279 4356
rect 8227 4230 8270 4354
rect 8408 4330 8471 4430
rect 8304 4314 8471 4330
rect 8338 4280 8471 4314
rect 8304 4264 8471 4280
rect 8042 4192 8193 4226
rect 7785 4126 7819 4142
rect 7530 4118 7729 4124
rect 7853 4124 7869 4158
rect 7903 4124 7923 4158
rect 7962 4150 7973 4184
rect 8141 4184 8193 4192
rect 7962 4134 8007 4150
rect 7853 4082 7923 4124
rect 8041 4124 8057 4158
rect 8091 4124 8107 4158
rect 8175 4150 8193 4184
rect 8141 4134 8193 4150
rect 8227 4209 8279 4230
rect 8227 4160 8245 4209
rect 8408 4184 8471 4264
rect 8041 4082 8107 4124
rect 8227 4116 8279 4160
rect 8313 4158 8372 4174
rect 8313 4124 8329 4158
rect 8363 4124 8372 4158
rect 8313 4082 8372 4124
rect 8408 4150 8424 4184
rect 8458 4150 8471 4184
rect 8408 4116 8471 4150
rect 8505 4513 8562 4558
rect 8596 4550 8873 4592
rect 8596 4516 8612 4550
rect 8646 4516 8823 4550
rect 8857 4516 8873 4550
rect 9061 4550 9137 4592
rect 8979 4524 9013 4540
rect 8505 4479 8528 4513
rect 9061 4516 9087 4550
rect 9121 4516 9137 4550
rect 9560 4550 9626 4592
rect 8979 4482 9013 4490
rect 9185 4515 9301 4549
rect 9335 4515 9351 4549
rect 9560 4516 9576 4550
rect 9610 4516 9626 4550
rect 9844 4540 9920 4592
rect 8505 4445 8562 4479
rect 8505 4411 8528 4445
rect 8505 4391 8562 4411
rect 8596 4448 9151 4482
rect 8505 4208 8546 4391
rect 8596 4330 8630 4448
rect 8693 4380 8709 4414
rect 8743 4388 8845 4414
rect 8743 4380 8790 4388
rect 8824 4354 8845 4388
rect 8790 4346 8845 4354
rect 8580 4314 8630 4330
rect 8614 4280 8630 4314
rect 8664 4325 8739 4330
rect 8664 4318 8682 4325
rect 8664 4284 8680 4318
rect 8716 4291 8739 4325
rect 8714 4284 8739 4291
rect 8790 4312 8811 4346
rect 8580 4264 8630 4280
rect 8790 4250 8845 4312
rect 8505 4192 8562 4208
rect 8505 4182 8528 4192
rect 8505 4148 8519 4182
rect 8553 4148 8562 4158
rect 8505 4116 8562 4148
rect 8596 4158 8662 4226
rect 8596 4124 8612 4158
rect 8646 4124 8662 4158
rect 8596 4082 8662 4124
rect 8707 4216 8845 4250
rect 8879 4221 8915 4448
rect 9101 4430 9151 4448
rect 9101 4396 9117 4430
rect 9101 4380 9151 4396
rect 9185 4346 9219 4515
rect 9560 4482 9626 4516
rect 9342 4456 9389 4462
rect 8949 4330 9219 4346
rect 8983 4312 9219 4330
rect 8983 4296 8993 4312
rect 8949 4280 8993 4296
rect 9035 4244 9057 4278
rect 9091 4252 9110 4278
rect 8879 4218 8945 4221
rect 8707 4168 8754 4216
rect 8879 4184 8895 4218
rect 8929 4184 8945 4218
rect 9035 4218 9066 4244
rect 9100 4218 9110 4252
rect 9035 4212 9110 4218
rect 8741 4134 8754 4168
rect 8707 4118 8754 4134
rect 8811 4166 8845 4182
rect 8979 4150 8995 4174
rect 8845 4140 8995 4150
rect 9029 4140 9045 4174
rect 8845 4132 9045 4140
rect 8811 4116 9045 4132
rect 9097 4154 9149 4170
rect 9131 4120 9149 4154
rect 9097 4082 9149 4120
rect 9185 4158 9219 4312
rect 9253 4430 9294 4446
rect 9287 4396 9294 4430
rect 9253 4326 9294 4396
rect 9376 4430 9389 4456
rect 9560 4448 9576 4482
rect 9610 4448 9626 4482
rect 9750 4524 9784 4540
rect 9844 4506 9870 4540
rect 9904 4506 9920 4540
rect 9968 4515 10084 4549
rect 10118 4515 10134 4549
rect 10177 4542 10211 4558
rect 9750 4472 9784 4490
rect 9664 4456 9934 4472
rect 9342 4396 9355 4422
rect 9664 4422 9750 4456
rect 9784 4430 9934 4456
rect 9784 4422 9900 4430
rect 9342 4380 9389 4396
rect 9429 4388 9630 4396
rect 9429 4354 9434 4388
rect 9468 4354 9630 4388
rect 9429 4348 9630 4354
rect 9564 4346 9630 4348
rect 9253 4320 9377 4326
rect 9253 4290 9342 4320
rect 9320 4286 9342 4290
rect 9376 4286 9377 4320
rect 9564 4312 9580 4346
rect 9614 4312 9630 4346
rect 9320 4256 9377 4286
rect 9354 4222 9377 4256
rect 9436 4278 9452 4312
rect 9486 4278 9502 4312
rect 9664 4278 9698 4422
rect 9884 4396 9900 4422
rect 9884 4380 9934 4396
rect 9732 4346 9782 4362
rect 9968 4346 10002 4515
rect 10177 4458 10211 4508
rect 10245 4526 10315 4592
rect 10245 4492 10261 4526
rect 10295 4492 10315 4526
rect 10354 4542 10399 4558
rect 10354 4508 10365 4542
rect 10354 4474 10399 4508
rect 10433 4526 10499 4592
rect 10433 4492 10449 4526
rect 10483 4492 10499 4526
rect 10533 4542 10585 4558
rect 10567 4508 10585 4542
rect 10036 4430 10078 4456
rect 10070 4422 10078 4430
rect 10112 4422 10136 4456
rect 10177 4424 10320 4458
rect 10070 4396 10136 4422
rect 10036 4380 10136 4396
rect 9766 4312 10002 4346
rect 9732 4296 9776 4312
rect 9922 4304 10002 4312
rect 9436 4244 9698 4278
rect 9818 4258 9834 4278
rect 9320 4206 9377 4222
rect 9654 4218 9698 4244
rect 9802 4252 9834 4258
rect 9868 4244 9884 4278
rect 9836 4218 9884 4244
rect 9586 4192 9620 4208
rect 9654 4184 9670 4218
rect 9704 4184 9720 4218
rect 9802 4212 9884 4218
rect 9185 4124 9288 4158
rect 9322 4124 9338 4158
rect 9185 4118 9338 4124
rect 9466 4124 9482 4158
rect 9516 4124 9532 4158
rect 9466 4082 9532 4124
rect 9586 4150 9620 4158
rect 9754 4150 9770 4174
rect 9586 4140 9770 4150
rect 9804 4140 9820 4174
rect 9586 4116 9820 4140
rect 9854 4154 9888 4170
rect 9854 4082 9888 4120
rect 9922 4158 9956 4304
rect 9990 4252 10006 4268
rect 10040 4234 10056 4268
rect 10024 4218 10056 4234
rect 9990 4194 10056 4218
rect 10092 4256 10136 4380
rect 10170 4387 10252 4390
rect 10170 4353 10214 4387
rect 10248 4353 10252 4387
rect 10170 4316 10252 4353
rect 10170 4282 10218 4316
rect 10170 4266 10252 4282
rect 10092 4222 10102 4256
rect 10286 4230 10320 4424
rect 10092 4206 10136 4222
rect 10177 4192 10320 4230
rect 10354 4440 10365 4474
rect 10533 4474 10585 4508
rect 10354 4252 10399 4440
rect 10388 4218 10399 4252
rect 10177 4176 10211 4192
rect 9922 4124 10071 4158
rect 10105 4124 10121 4158
rect 10354 4184 10399 4218
rect 10434 4456 10533 4458
rect 10434 4422 10446 4456
rect 10480 4440 10533 4456
rect 10567 4440 10585 4474
rect 10480 4424 10585 4440
rect 10619 4514 10671 4558
rect 10619 4480 10637 4514
rect 10619 4446 10671 4480
rect 10434 4329 10480 4422
rect 10619 4412 10637 4446
rect 10705 4538 10764 4592
rect 10705 4504 10721 4538
rect 10755 4504 10764 4538
rect 10705 4470 10764 4504
rect 10705 4436 10721 4470
rect 10755 4436 10764 4470
rect 10705 4418 10764 4436
rect 10800 4532 10863 4548
rect 10800 4498 10816 4532
rect 10850 4498 10863 4532
rect 10800 4464 10863 4498
rect 10800 4430 10816 4464
rect 10850 4430 10863 4464
rect 10619 4391 10671 4412
rect 10468 4295 10480 4329
rect 10434 4226 10480 4295
rect 10514 4329 10585 4390
rect 10514 4295 10536 4329
rect 10570 4302 10585 4329
rect 10514 4268 10538 4295
rect 10572 4268 10585 4302
rect 10514 4260 10585 4268
rect 10619 4357 10625 4391
rect 10659 4357 10671 4391
rect 10619 4354 10671 4357
rect 10619 4230 10662 4354
rect 10800 4330 10863 4430
rect 10696 4314 10863 4330
rect 10730 4280 10863 4314
rect 10696 4264 10863 4280
rect 10434 4192 10585 4226
rect 10177 4126 10211 4142
rect 9922 4118 10121 4124
rect 10245 4124 10261 4158
rect 10295 4124 10315 4158
rect 10354 4150 10365 4184
rect 10533 4184 10585 4192
rect 10354 4134 10399 4150
rect 10245 4082 10315 4124
rect 10433 4124 10449 4158
rect 10483 4124 10499 4158
rect 10567 4150 10585 4184
rect 10533 4134 10585 4150
rect 10619 4217 10671 4230
rect 10619 4183 10633 4217
rect 10667 4194 10671 4217
rect 10619 4160 10637 4183
rect 10800 4184 10863 4264
rect 10433 4082 10499 4124
rect 10619 4116 10671 4160
rect 10705 4158 10764 4174
rect 10705 4124 10721 4158
rect 10755 4124 10764 4158
rect 10705 4082 10764 4124
rect 10800 4150 10816 4184
rect 10850 4150 10863 4184
rect 10800 4116 10863 4150
rect 10897 4513 10954 4558
rect 10988 4550 11265 4592
rect 10988 4516 11004 4550
rect 11038 4516 11215 4550
rect 11249 4516 11265 4550
rect 11453 4550 11529 4592
rect 11371 4524 11405 4540
rect 10897 4479 10920 4513
rect 11453 4516 11479 4550
rect 11513 4516 11529 4550
rect 11952 4550 12018 4592
rect 11371 4482 11405 4490
rect 11577 4515 11693 4549
rect 11727 4515 11743 4549
rect 11952 4516 11968 4550
rect 12002 4516 12018 4550
rect 12236 4540 12312 4592
rect 10897 4445 10954 4479
rect 10897 4411 10920 4445
rect 10897 4391 10954 4411
rect 10988 4448 11543 4482
rect 10897 4208 10938 4391
rect 10988 4330 11022 4448
rect 11085 4380 11101 4414
rect 11135 4388 11237 4414
rect 11135 4380 11182 4388
rect 11216 4354 11237 4388
rect 11182 4346 11237 4354
rect 10972 4314 11022 4330
rect 11006 4280 11022 4314
rect 11056 4322 11131 4330
rect 11056 4318 11076 4322
rect 11056 4284 11072 4318
rect 11110 4288 11131 4322
rect 11106 4284 11131 4288
rect 11182 4312 11203 4346
rect 10972 4264 11022 4280
rect 11182 4250 11237 4312
rect 10897 4192 10954 4208
rect 10897 4188 10920 4192
rect 10897 4154 10913 4188
rect 10947 4154 10954 4158
rect 10897 4116 10954 4154
rect 10988 4158 11054 4226
rect 10988 4124 11004 4158
rect 11038 4124 11054 4158
rect 10988 4082 11054 4124
rect 11099 4216 11237 4250
rect 11271 4221 11307 4448
rect 11493 4430 11543 4448
rect 11493 4396 11509 4430
rect 11493 4380 11543 4396
rect 11577 4346 11611 4515
rect 11952 4482 12018 4516
rect 11734 4456 11781 4462
rect 11341 4330 11611 4346
rect 11375 4312 11611 4330
rect 11375 4296 11385 4312
rect 11341 4280 11385 4296
rect 11427 4244 11449 4278
rect 11483 4252 11502 4278
rect 11271 4218 11337 4221
rect 11099 4168 11146 4216
rect 11271 4184 11287 4218
rect 11321 4184 11337 4218
rect 11427 4218 11458 4244
rect 11492 4218 11502 4252
rect 11427 4212 11502 4218
rect 11133 4134 11146 4168
rect 11099 4118 11146 4134
rect 11203 4166 11237 4182
rect 11371 4150 11387 4174
rect 11237 4140 11387 4150
rect 11421 4140 11437 4174
rect 11237 4132 11437 4140
rect 11203 4116 11437 4132
rect 11489 4154 11541 4170
rect 11523 4120 11541 4154
rect 11489 4082 11541 4120
rect 11577 4158 11611 4312
rect 11645 4430 11686 4446
rect 11679 4396 11686 4430
rect 11645 4326 11686 4396
rect 11768 4430 11781 4456
rect 11952 4448 11968 4482
rect 12002 4448 12018 4482
rect 12142 4524 12176 4540
rect 12236 4506 12262 4540
rect 12296 4506 12312 4540
rect 12360 4515 12476 4549
rect 12510 4515 12526 4549
rect 12569 4542 12603 4558
rect 12142 4472 12176 4490
rect 12056 4456 12326 4472
rect 11734 4396 11747 4422
rect 12056 4422 12142 4456
rect 12176 4430 12326 4456
rect 12176 4422 12292 4430
rect 11734 4380 11781 4396
rect 11821 4388 12022 4396
rect 11821 4354 11826 4388
rect 11860 4354 12022 4388
rect 11821 4348 12022 4354
rect 11956 4346 12022 4348
rect 11645 4320 11769 4326
rect 11645 4290 11734 4320
rect 11712 4286 11734 4290
rect 11768 4286 11769 4320
rect 11956 4312 11972 4346
rect 12006 4312 12022 4346
rect 11712 4256 11769 4286
rect 11746 4222 11769 4256
rect 11828 4278 11844 4312
rect 11878 4278 11894 4312
rect 12056 4278 12090 4422
rect 12276 4396 12292 4422
rect 12276 4380 12326 4396
rect 12124 4346 12174 4362
rect 12360 4346 12394 4515
rect 12569 4458 12603 4508
rect 12637 4526 12707 4592
rect 12637 4492 12653 4526
rect 12687 4492 12707 4526
rect 12746 4542 12791 4558
rect 12746 4508 12757 4542
rect 12746 4474 12791 4508
rect 12825 4526 12891 4592
rect 12825 4492 12841 4526
rect 12875 4492 12891 4526
rect 12925 4542 12977 4558
rect 12959 4508 12977 4542
rect 12428 4430 12470 4456
rect 12462 4422 12470 4430
rect 12504 4422 12528 4456
rect 12569 4424 12712 4458
rect 12462 4396 12528 4422
rect 12428 4380 12528 4396
rect 12158 4312 12394 4346
rect 12124 4296 12168 4312
rect 12314 4304 12394 4312
rect 11828 4244 12090 4278
rect 12210 4258 12226 4278
rect 11712 4206 11769 4222
rect 12046 4218 12090 4244
rect 12194 4252 12226 4258
rect 12260 4244 12276 4278
rect 12228 4218 12276 4244
rect 11978 4192 12012 4208
rect 12046 4184 12062 4218
rect 12096 4184 12112 4218
rect 12194 4212 12276 4218
rect 11577 4124 11680 4158
rect 11714 4124 11730 4158
rect 11577 4118 11730 4124
rect 11858 4124 11874 4158
rect 11908 4124 11924 4158
rect 11858 4082 11924 4124
rect 11978 4150 12012 4158
rect 12146 4150 12162 4174
rect 11978 4140 12162 4150
rect 12196 4140 12212 4174
rect 11978 4116 12212 4140
rect 12246 4154 12280 4170
rect 12246 4082 12280 4120
rect 12314 4158 12348 4304
rect 12382 4252 12398 4268
rect 12432 4234 12448 4268
rect 12416 4218 12448 4234
rect 12382 4194 12448 4218
rect 12484 4256 12528 4380
rect 12562 4383 12644 4390
rect 12562 4349 12575 4383
rect 12609 4349 12644 4383
rect 12562 4316 12644 4349
rect 12562 4282 12610 4316
rect 12562 4266 12644 4282
rect 12484 4222 12494 4256
rect 12678 4230 12712 4424
rect 12484 4206 12528 4222
rect 12569 4192 12712 4230
rect 12746 4440 12757 4474
rect 12925 4474 12977 4508
rect 12746 4252 12791 4440
rect 12780 4218 12791 4252
rect 12569 4176 12603 4192
rect 12314 4124 12463 4158
rect 12497 4124 12513 4158
rect 12746 4184 12791 4218
rect 12826 4456 12925 4458
rect 12826 4422 12838 4456
rect 12872 4440 12925 4456
rect 12959 4440 12977 4474
rect 12872 4424 12977 4440
rect 12826 4329 12872 4422
rect 12860 4295 12872 4329
rect 12826 4226 12872 4295
rect 12906 4375 12977 4390
rect 12906 4341 12930 4375
rect 12964 4341 12977 4375
rect 12906 4329 12977 4341
rect 12906 4295 12928 4329
rect 12962 4295 12977 4329
rect 12906 4260 12977 4295
rect 12826 4192 12977 4226
rect 12569 4126 12603 4142
rect 12314 4118 12513 4124
rect 12637 4124 12653 4158
rect 12687 4124 12707 4158
rect 12746 4150 12757 4184
rect 12925 4184 12977 4192
rect 12746 4134 12791 4150
rect 12637 4082 12707 4124
rect 12825 4124 12841 4158
rect 12875 4124 12891 4158
rect 12959 4150 12977 4184
rect 12925 4134 12977 4150
rect 12825 4082 12891 4124
rect 594 4024 623 4082
rect 657 4024 715 4082
rect 749 4024 807 4082
rect 841 4024 899 4082
rect 933 4024 991 4082
rect 1025 4024 1083 4082
rect 1117 4024 1175 4082
rect 1209 4024 1267 4082
rect 1301 4024 1359 4082
rect 1393 4048 1431 4082
rect 1465 4058 1523 4082
rect 1557 4058 1615 4082
rect 1649 4058 1707 4082
rect 1741 4058 1799 4082
rect 1833 4058 1891 4082
rect 1925 4058 1983 4082
rect 2017 4058 2075 4082
rect 2109 4058 2167 4082
rect 2201 4058 2259 4082
rect 2293 4058 2351 4082
rect 2385 4058 2443 4082
rect 2477 4058 2535 4082
rect 2569 4058 2627 4082
rect 2661 4058 2719 4082
rect 2753 4058 2811 4082
rect 2845 4058 2903 4082
rect 2937 4058 2995 4082
rect 3029 4058 3087 4082
rect 3121 4058 3179 4082
rect 3213 4058 3271 4082
rect 3305 4058 3363 4082
rect 3397 4058 3455 4082
rect 3489 4058 3547 4082
rect 3581 4058 3639 4082
rect 3673 4058 3731 4082
rect 3765 4058 3823 4082
rect 3857 4058 3915 4082
rect 3949 4058 4007 4082
rect 4041 4058 4099 4082
rect 4133 4058 4191 4082
rect 4225 4058 4283 4082
rect 4317 4058 4375 4082
rect 4409 4058 4467 4082
rect 4501 4058 4559 4082
rect 4593 4058 4651 4082
rect 4685 4058 4743 4082
rect 4777 4058 4835 4082
rect 4869 4058 4927 4082
rect 4961 4058 5019 4082
rect 5053 4058 5111 4082
rect 5145 4058 5203 4082
rect 5237 4058 5295 4082
rect 5329 4058 5387 4082
rect 5421 4058 5479 4082
rect 5513 4058 5571 4082
rect 5605 4058 5663 4082
rect 5697 4058 5755 4082
rect 5789 4058 5847 4082
rect 5881 4058 5939 4082
rect 5973 4058 6031 4082
rect 6065 4058 6123 4082
rect 6157 4058 6215 4082
rect 6249 4058 6307 4082
rect 6341 4058 6399 4082
rect 6433 4058 6491 4082
rect 6525 4058 6583 4082
rect 6617 4058 6675 4082
rect 6709 4058 6767 4082
rect 6801 4058 6859 4082
rect 6893 4058 6951 4082
rect 6985 4058 7043 4082
rect 7077 4058 7135 4082
rect 7169 4058 7227 4082
rect 7261 4058 7319 4082
rect 7353 4058 7411 4082
rect 7445 4058 7503 4082
rect 7537 4058 7595 4082
rect 7629 4058 7687 4082
rect 7721 4058 7779 4082
rect 7813 4058 7871 4082
rect 7905 4058 7963 4082
rect 7997 4058 8055 4082
rect 8089 4058 8147 4082
rect 8181 4058 8239 4082
rect 8273 4058 8331 4082
rect 8365 4058 8423 4082
rect 8457 4058 8515 4082
rect 8549 4058 8607 4082
rect 8641 4058 8699 4082
rect 8733 4058 8791 4082
rect 8825 4058 8883 4082
rect 8917 4058 8975 4082
rect 9009 4058 9067 4082
rect 9101 4058 9159 4082
rect 9193 4058 9251 4082
rect 9285 4058 9343 4082
rect 9377 4058 9435 4082
rect 1485 4048 1523 4058
rect 1577 4048 1615 4058
rect 1669 4048 1707 4058
rect 1761 4048 1799 4058
rect 1853 4048 1891 4058
rect 1945 4048 1983 4058
rect 2037 4048 2075 4058
rect 2129 4048 2167 4058
rect 2221 4048 2259 4058
rect 2313 4048 2351 4058
rect 2405 4048 2443 4058
rect 2497 4048 2535 4058
rect 2589 4048 2627 4058
rect 2681 4048 2719 4058
rect 2773 4048 2811 4058
rect 2865 4048 2903 4058
rect 2957 4048 2995 4058
rect 3049 4048 3087 4058
rect 3141 4048 3179 4058
rect 3233 4048 3271 4058
rect 3325 4048 3363 4058
rect 3417 4048 3455 4058
rect 3509 4048 3547 4058
rect 3601 4048 3639 4058
rect 3693 4048 3731 4058
rect 3785 4048 3823 4058
rect 3877 4048 3915 4058
rect 3969 4048 4007 4058
rect 4061 4048 4099 4058
rect 4153 4048 4191 4058
rect 4245 4048 4283 4058
rect 4337 4048 4375 4058
rect 4429 4048 4467 4058
rect 4521 4048 4559 4058
rect 4613 4048 4651 4058
rect 4705 4048 4743 4058
rect 4797 4048 4835 4058
rect 4889 4048 4927 4058
rect 4981 4048 5019 4058
rect 5073 4048 5111 4058
rect 5165 4048 5203 4058
rect 5257 4048 5295 4058
rect 5349 4048 5387 4058
rect 5441 4048 5479 4058
rect 5533 4048 5571 4058
rect 5625 4048 5663 4058
rect 5717 4048 5755 4058
rect 5809 4048 5847 4058
rect 5901 4048 5939 4058
rect 5993 4048 6031 4058
rect 6085 4048 6123 4058
rect 6177 4048 6215 4058
rect 6269 4048 6307 4058
rect 6361 4048 6399 4058
rect 6453 4048 6491 4058
rect 6545 4048 6583 4058
rect 6637 4048 6675 4058
rect 6729 4048 6767 4058
rect 6821 4048 6859 4058
rect 6913 4048 6951 4058
rect 7005 4048 7043 4058
rect 7097 4048 7135 4058
rect 7189 4048 7227 4058
rect 7281 4048 7319 4058
rect 7373 4048 7411 4058
rect 7465 4048 7503 4058
rect 7557 4048 7595 4058
rect 7649 4048 7687 4058
rect 7741 4048 7779 4058
rect 7833 4048 7871 4058
rect 7925 4048 7963 4058
rect 8017 4048 8055 4058
rect 8109 4048 8147 4058
rect 8201 4048 8239 4058
rect 8293 4048 8331 4058
rect 8385 4048 8423 4058
rect 8477 4048 8515 4058
rect 8569 4048 8607 4058
rect 8661 4048 8699 4058
rect 8753 4048 8791 4058
rect 8845 4048 8883 4058
rect 8937 4048 8975 4058
rect 9029 4048 9067 4058
rect 9121 4048 9159 4058
rect 9213 4048 9251 4058
rect 9305 4048 9343 4058
rect 1393 4024 1451 4048
rect 1485 4024 1543 4048
rect 1577 4024 1635 4048
rect 1669 4024 1727 4048
rect 1761 4024 1819 4048
rect 1853 4024 1911 4048
rect 1945 4024 2003 4048
rect 2037 4024 2095 4048
rect 2129 4024 2187 4048
rect 2221 4024 2279 4048
rect 2313 4024 2371 4048
rect 2405 4024 2463 4048
rect 2497 4024 2555 4048
rect 2589 4024 2647 4048
rect 2681 4024 2739 4048
rect 2773 4024 2831 4048
rect 2865 4024 2923 4048
rect 2957 4024 3015 4048
rect 3049 4024 3107 4048
rect 3141 4024 3199 4048
rect 3233 4024 3291 4048
rect 3325 4024 3383 4048
rect 3417 4024 3475 4048
rect 3509 4024 3567 4048
rect 3601 4024 3659 4048
rect 3693 4024 3751 4048
rect 3785 4024 3843 4048
rect 3877 4024 3935 4048
rect 3969 4024 4027 4048
rect 4061 4024 4119 4048
rect 4153 4024 4211 4048
rect 4245 4024 4303 4048
rect 4337 4024 4395 4048
rect 4429 4024 4487 4048
rect 4521 4024 4579 4048
rect 4613 4024 4671 4048
rect 4705 4024 4763 4048
rect 4797 4024 4855 4048
rect 4889 4024 4947 4048
rect 4981 4024 5039 4048
rect 5073 4024 5131 4048
rect 5165 4024 5223 4048
rect 5257 4024 5315 4048
rect 5349 4024 5407 4048
rect 5441 4024 5499 4048
rect 5533 4024 5591 4048
rect 5625 4024 5683 4048
rect 5717 4024 5775 4048
rect 5809 4024 5867 4048
rect 5901 4024 5959 4048
rect 5993 4024 6051 4048
rect 6085 4024 6143 4048
rect 6177 4024 6235 4048
rect 6269 4024 6327 4048
rect 6361 4024 6419 4048
rect 6453 4024 6511 4048
rect 6545 4024 6603 4048
rect 6637 4024 6695 4048
rect 6729 4024 6787 4048
rect 6821 4024 6879 4048
rect 6913 4024 6971 4048
rect 7005 4024 7063 4048
rect 7097 4024 7155 4048
rect 7189 4024 7247 4048
rect 7281 4024 7339 4048
rect 7373 4024 7431 4048
rect 7465 4024 7523 4048
rect 7557 4024 7615 4048
rect 7649 4024 7707 4048
rect 7741 4024 7799 4048
rect 7833 4024 7891 4048
rect 7925 4024 7983 4048
rect 8017 4024 8075 4048
rect 8109 4024 8167 4048
rect 8201 4024 8259 4048
rect 8293 4024 8351 4048
rect 8385 4024 8443 4048
rect 8477 4024 8535 4048
rect 8569 4024 8627 4048
rect 8661 4024 8719 4048
rect 8753 4024 8811 4048
rect 8845 4024 8903 4048
rect 8937 4024 8995 4048
rect 9029 4024 9087 4048
rect 9121 4024 9179 4048
rect 9213 4024 9271 4048
rect 9305 4024 9363 4048
rect 9397 4024 9435 4058
rect 9469 4024 9527 4082
rect 9561 4024 9619 4082
rect 9653 4024 9711 4082
rect 9745 4024 9803 4082
rect 9837 4024 9895 4082
rect 9929 4024 9987 4082
rect 10021 4024 10079 4082
rect 10113 4024 10171 4082
rect 10205 4024 10263 4082
rect 10297 4024 10355 4082
rect 10389 4024 10447 4082
rect 10481 4024 10539 4082
rect 10573 4024 10631 4082
rect 10665 4024 10723 4082
rect 10757 4024 10815 4082
rect 10849 4024 10907 4082
rect 10941 4024 10999 4082
rect 11033 4024 11091 4082
rect 11125 4024 11183 4082
rect 11217 4024 11275 4082
rect 11309 4024 11367 4082
rect 11401 4024 11459 4082
rect 11493 4024 11551 4082
rect 11585 4024 11643 4082
rect 11677 4024 11735 4082
rect 11769 4024 11827 4082
rect 11861 4024 11919 4082
rect 11953 4024 12011 4082
rect 12045 4024 12103 4082
rect 12137 4024 12195 4082
rect 12229 4024 12287 4082
rect 12321 4024 12379 4082
rect 12413 4024 12471 4082
rect 12505 4024 12563 4082
rect 12597 4024 12655 4082
rect 12689 4024 12747 4082
rect 12781 4024 12839 4082
rect 12873 4024 12931 4082
rect 12965 4024 12994 4082
rect 626 3718 655 3786
rect 689 3718 747 3786
rect 781 3718 839 3786
rect 873 3718 931 3786
rect 965 3718 1023 3786
rect 1057 3752 1114 3786
rect 1148 3752 1206 3786
rect 1240 3752 1299 3786
rect 1057 3718 1115 3752
rect 1149 3718 1207 3752
rect 1241 3718 1299 3752
rect 1333 3718 1391 3786
rect 1425 3751 1455 3786
rect 1425 3718 1454 3751
rect 3168 3719 3197 3777
rect 3231 3719 3289 3777
rect 3323 3719 3381 3777
rect 3415 3753 3473 3777
rect 3507 3753 3565 3777
rect 3599 3753 3657 3777
rect 3691 3753 3749 3777
rect 3783 3753 3841 3777
rect 3875 3753 3933 3777
rect 3967 3753 4025 3777
rect 4059 3753 4117 3777
rect 4151 3753 4209 3777
rect 4243 3753 4301 3777
rect 4335 3753 4393 3777
rect 4427 3753 4485 3777
rect 4519 3753 4577 3777
rect 4611 3753 4669 3777
rect 4703 3753 4761 3777
rect 4795 3753 4853 3777
rect 4887 3753 4945 3777
rect 3415 3719 3454 3753
rect 3507 3743 3546 3753
rect 3599 3743 3638 3753
rect 3691 3743 3730 3753
rect 3783 3743 3822 3753
rect 3875 3743 3914 3753
rect 3967 3743 4006 3753
rect 4059 3743 4098 3753
rect 4151 3743 4190 3753
rect 4243 3743 4282 3753
rect 4335 3743 4374 3753
rect 4427 3743 4466 3753
rect 4519 3743 4558 3753
rect 4611 3743 4650 3753
rect 4703 3743 4742 3753
rect 4795 3743 4834 3753
rect 4887 3743 4926 3753
rect 4979 3743 5018 3777
rect 3488 3719 3546 3743
rect 3580 3719 3638 3743
rect 3672 3719 3730 3743
rect 3764 3719 3822 3743
rect 3856 3719 3914 3743
rect 3948 3719 4006 3743
rect 4040 3719 4098 3743
rect 4132 3719 4190 3743
rect 4224 3719 4282 3743
rect 4316 3719 4374 3743
rect 4408 3719 4466 3743
rect 4500 3719 4558 3743
rect 4592 3719 4650 3743
rect 4684 3719 4742 3743
rect 4776 3719 4834 3743
rect 4868 3719 4926 3743
rect 4960 3719 5018 3743
rect 5052 3719 5110 3777
rect 5144 3719 5202 3777
rect 5236 3719 5294 3777
rect 5328 3719 5386 3777
rect 5420 3719 5478 3777
rect 5512 3719 5570 3777
rect 5604 3719 5662 3777
rect 5696 3719 5754 3777
rect 5788 3719 5846 3777
rect 5880 3719 5938 3777
rect 5972 3719 6030 3777
rect 6064 3719 6122 3777
rect 6156 3719 6214 3777
rect 6248 3719 6306 3777
rect 6340 3719 6398 3777
rect 6432 3719 6490 3777
rect 6524 3719 6582 3777
rect 6616 3719 6674 3777
rect 6708 3719 6766 3777
rect 6800 3719 6858 3777
rect 6892 3719 6950 3777
rect 6984 3719 7042 3777
rect 7076 3719 7134 3777
rect 7168 3719 7226 3777
rect 7260 3719 7318 3777
rect 7352 3719 7410 3777
rect 7444 3719 7502 3777
rect 7536 3719 7594 3777
rect 7628 3719 7686 3777
rect 7720 3719 7778 3777
rect 7812 3719 7870 3777
rect 7904 3719 7962 3777
rect 7996 3719 8054 3777
rect 8088 3719 8146 3777
rect 8180 3719 8238 3777
rect 8272 3719 8330 3777
rect 8364 3719 8422 3777
rect 8456 3719 8514 3777
rect 8548 3719 8606 3777
rect 8640 3719 8698 3777
rect 8732 3719 8790 3777
rect 8824 3719 8882 3777
rect 8916 3719 8974 3777
rect 9008 3719 9066 3777
rect 9100 3719 9158 3777
rect 9192 3719 9250 3777
rect 9284 3719 9342 3777
rect 9376 3719 9434 3777
rect 9468 3719 9526 3777
rect 9560 3719 9618 3777
rect 9652 3719 9710 3777
rect 9744 3719 9802 3777
rect 9836 3719 9894 3777
rect 9928 3719 9986 3777
rect 10020 3719 10078 3777
rect 10112 3719 10170 3777
rect 10204 3719 10262 3777
rect 10296 3719 10354 3777
rect 10388 3719 10446 3777
rect 10480 3719 10538 3777
rect 10572 3719 10630 3777
rect 10664 3719 10722 3777
rect 10756 3719 10814 3777
rect 10848 3719 10906 3777
rect 10940 3719 10998 3777
rect 11032 3719 11090 3777
rect 11124 3719 11182 3777
rect 11216 3719 11274 3777
rect 11308 3719 11366 3777
rect 11400 3719 11458 3777
rect 11492 3719 11550 3777
rect 11584 3719 11642 3777
rect 11676 3719 11734 3777
rect 11768 3719 11826 3777
rect 11860 3719 11918 3777
rect 11952 3719 12010 3777
rect 12044 3719 12102 3777
rect 12136 3719 12194 3777
rect 12228 3719 12286 3777
rect 12320 3719 12378 3777
rect 12412 3719 12470 3777
rect 12504 3719 12562 3777
rect 12596 3719 12654 3777
rect 12688 3719 12746 3777
rect 12780 3719 12838 3777
rect 12872 3719 12930 3777
rect 12964 3719 12993 3777
rect 659 3668 695 3684
rect 659 3634 661 3668
rect 659 3600 695 3634
rect 659 3566 661 3600
rect 731 3668 797 3718
rect 731 3634 747 3668
rect 781 3634 797 3668
rect 731 3600 797 3634
rect 731 3566 747 3600
rect 781 3566 797 3600
rect 831 3668 885 3684
rect 831 3634 833 3668
rect 867 3634 885 3668
rect 831 3587 885 3634
rect 659 3532 695 3566
rect 831 3553 833 3587
rect 867 3553 885 3587
rect 659 3498 794 3532
rect 831 3503 885 3553
rect 760 3469 794 3498
rect 647 3440 715 3462
rect 647 3406 663 3440
rect 697 3439 715 3440
rect 647 3405 665 3406
rect 699 3405 715 3439
rect 647 3388 715 3405
rect 760 3453 815 3469
rect 760 3419 781 3453
rect 760 3403 815 3419
rect 849 3454 885 3503
rect 921 3670 987 3684
rect 921 3636 937 3670
rect 971 3636 987 3670
rect 921 3602 987 3636
rect 921 3568 937 3602
rect 971 3568 987 3602
rect 921 3534 987 3568
rect 1021 3676 1069 3718
rect 1055 3642 1069 3676
rect 1021 3608 1069 3642
rect 1055 3574 1069 3608
rect 1021 3558 1069 3574
rect 1105 3654 1139 3684
rect 1105 3559 1139 3620
rect 921 3500 937 3534
rect 971 3522 987 3534
rect 1173 3676 1239 3718
rect 1173 3642 1189 3676
rect 1223 3642 1239 3676
rect 1173 3608 1239 3642
rect 1173 3574 1189 3608
rect 1223 3574 1239 3608
rect 1173 3558 1239 3574
rect 1273 3654 1307 3684
rect 1273 3559 1307 3620
rect 971 3500 1064 3522
rect 921 3488 1064 3500
rect 849 3440 996 3454
rect 849 3406 946 3440
rect 980 3406 996 3440
rect 1030 3440 1064 3488
rect 1105 3514 1139 3525
rect 1273 3514 1307 3525
rect 1105 3480 1307 3514
rect 1341 3676 1407 3718
rect 1341 3642 1357 3676
rect 1391 3642 1407 3676
rect 1341 3608 1407 3642
rect 1341 3574 1357 3608
rect 1391 3574 1407 3608
rect 1341 3540 1407 3574
rect 1341 3506 1357 3540
rect 1391 3506 1407 3540
rect 1341 3488 1407 3506
rect 3236 3677 3278 3719
rect 3236 3643 3244 3677
rect 3236 3609 3278 3643
rect 3236 3575 3244 3609
rect 3236 3541 3278 3575
rect 3236 3507 3244 3541
rect 3236 3491 3278 3507
rect 3312 3677 3378 3685
rect 3312 3643 3328 3677
rect 3362 3643 3378 3677
rect 3312 3609 3378 3643
rect 3312 3575 3328 3609
rect 3362 3575 3378 3609
rect 3312 3541 3378 3575
rect 3442 3669 3494 3685
rect 3442 3635 3460 3669
rect 3442 3601 3494 3635
rect 3528 3653 3594 3719
rect 3528 3619 3544 3653
rect 3578 3619 3594 3653
rect 3628 3669 3673 3685
rect 3662 3635 3673 3669
rect 3442 3567 3460 3601
rect 3628 3601 3673 3635
rect 3712 3653 3782 3719
rect 3712 3619 3732 3653
rect 3766 3619 3782 3653
rect 3816 3669 3850 3685
rect 3893 3642 3909 3676
rect 3943 3642 4059 3676
rect 3494 3583 3593 3585
rect 3494 3567 3547 3583
rect 3442 3551 3547 3567
rect 3312 3507 3328 3541
rect 3362 3520 3378 3541
rect 3581 3549 3593 3583
rect 3312 3489 3347 3507
rect 1208 3440 1307 3480
rect 3332 3486 3347 3489
rect 1030 3406 1080 3440
rect 1114 3406 1130 3440
rect 1208 3406 1270 3440
rect 1304 3406 1307 3440
rect 3160 3446 3298 3455
rect 3160 3412 3162 3446
rect 3196 3441 3298 3446
rect 3196 3412 3248 3441
rect 3160 3407 3248 3412
rect 3282 3407 3298 3441
rect 760 3352 794 3403
rect 661 3318 794 3352
rect 849 3343 885 3406
rect 1030 3372 1064 3406
rect 1208 3372 1307 3406
rect 661 3297 695 3318
rect 833 3314 885 3343
rect 661 3242 695 3263
rect 731 3250 747 3284
rect 781 3250 797 3284
rect 731 3208 797 3250
rect 867 3280 885 3314
rect 833 3242 885 3280
rect 937 3338 1064 3372
rect 1105 3338 1307 3372
rect 937 3320 971 3338
rect 1105 3320 1139 3338
rect 937 3242 971 3286
rect 1007 3288 1055 3304
rect 1007 3254 1021 3288
rect 1007 3208 1055 3254
rect 1273 3320 1307 3338
rect 1105 3242 1139 3286
rect 1173 3288 1239 3304
rect 1173 3254 1189 3288
rect 1223 3254 1239 3288
rect 1173 3208 1239 3254
rect 1273 3242 1307 3286
rect 1341 3352 1407 3368
rect 1341 3318 1357 3352
rect 1391 3318 1407 3352
rect 1341 3284 1407 3318
rect 1341 3250 1357 3284
rect 1391 3250 1407 3284
rect 1341 3208 1407 3250
rect 3232 3357 3278 3373
rect 3332 3369 3378 3486
rect 3442 3456 3513 3517
rect 3442 3445 3457 3456
rect 3442 3411 3455 3445
rect 3491 3422 3513 3456
rect 3489 3411 3513 3422
rect 3442 3387 3513 3411
rect 3547 3456 3593 3549
rect 3547 3422 3559 3456
rect 3232 3323 3244 3357
rect 3232 3289 3278 3323
rect 3232 3255 3244 3289
rect 3232 3209 3278 3255
rect 3312 3357 3378 3369
rect 3312 3323 3328 3357
rect 3362 3323 3378 3357
rect 3547 3353 3593 3422
rect 3312 3289 3378 3323
rect 3312 3255 3328 3289
rect 3362 3255 3378 3289
rect 3442 3319 3593 3353
rect 3662 3567 3673 3601
rect 3816 3585 3850 3635
rect 3628 3379 3673 3567
rect 3628 3345 3639 3379
rect 3442 3311 3494 3319
rect 3442 3277 3460 3311
rect 3628 3311 3673 3345
rect 3707 3551 3850 3585
rect 3707 3357 3741 3551
rect 3891 3549 3915 3583
rect 3949 3557 3991 3583
rect 3949 3549 3957 3557
rect 3891 3523 3957 3549
rect 3775 3453 3857 3517
rect 3775 3443 3784 3453
rect 3818 3419 3857 3453
rect 3809 3409 3857 3419
rect 3775 3393 3857 3409
rect 3891 3507 3991 3523
rect 3891 3383 3935 3507
rect 4025 3473 4059 3642
rect 4107 3667 4183 3719
rect 4401 3677 4467 3719
rect 4107 3633 4123 3667
rect 4157 3633 4183 3667
rect 4243 3651 4277 3667
rect 4243 3599 4277 3617
rect 4401 3643 4417 3677
rect 4451 3643 4467 3677
rect 4890 3677 4966 3719
rect 4401 3609 4467 3643
rect 4676 3642 4692 3676
rect 4726 3642 4842 3676
rect 4890 3643 4906 3677
rect 4940 3643 4966 3677
rect 5154 3677 5431 3719
rect 5014 3651 5048 3667
rect 4093 3583 4363 3599
rect 4093 3557 4243 3583
rect 4127 3549 4243 3557
rect 4277 3549 4363 3583
rect 4401 3575 4417 3609
rect 4451 3575 4467 3609
rect 4638 3583 4685 3589
rect 4127 3523 4143 3549
rect 4093 3507 4143 3523
rect 4245 3473 4295 3489
rect 4025 3439 4261 3473
rect 4025 3431 4105 3439
rect 3707 3319 3850 3357
rect 3925 3349 3935 3383
rect 3891 3333 3935 3349
rect 3971 3361 3987 3395
rect 4021 3379 4037 3395
rect 3971 3345 4003 3361
rect 3971 3321 4037 3345
rect 3442 3261 3494 3277
rect 3312 3243 3378 3255
rect 3528 3251 3544 3285
rect 3578 3251 3594 3285
rect 3662 3277 3673 3311
rect 3816 3303 3850 3319
rect 3628 3261 3673 3277
rect 3528 3209 3594 3251
rect 3712 3251 3732 3285
rect 3766 3251 3782 3285
rect 4071 3285 4105 3431
rect 4251 3423 4295 3439
rect 4329 3405 4363 3549
rect 4638 3557 4651 3583
rect 4672 3523 4685 3549
rect 4397 3515 4598 3523
rect 4397 3481 4559 3515
rect 4593 3481 4598 3515
rect 4638 3507 4685 3523
rect 4733 3557 4774 3573
rect 4733 3523 4740 3557
rect 4397 3475 4598 3481
rect 4397 3473 4463 3475
rect 4397 3439 4413 3473
rect 4447 3439 4463 3473
rect 4733 3453 4774 3523
rect 4650 3447 4774 3453
rect 4525 3405 4541 3439
rect 4575 3405 4591 3439
rect 4143 3371 4159 3405
rect 4193 3385 4209 3405
rect 4193 3379 4225 3385
rect 4143 3345 4191 3371
rect 4329 3371 4591 3405
rect 4650 3413 4651 3447
rect 4685 3417 4774 3447
rect 4808 3473 4842 3642
rect 5154 3643 5170 3677
rect 5204 3643 5381 3677
rect 5415 3643 5431 3677
rect 5014 3609 5048 3617
rect 5465 3640 5522 3685
rect 4876 3575 5431 3609
rect 4876 3557 4926 3575
rect 4910 3523 4926 3557
rect 4876 3507 4926 3523
rect 4808 3457 5078 3473
rect 4808 3439 5044 3457
rect 4685 3413 4707 3417
rect 4650 3383 4707 3413
rect 4329 3345 4373 3371
rect 4143 3339 4225 3345
rect 4307 3311 4323 3345
rect 4357 3311 4373 3345
rect 4650 3349 4673 3383
rect 4407 3319 4441 3335
rect 4650 3333 4707 3349
rect 3816 3253 3850 3269
rect 3712 3209 3782 3251
rect 3906 3251 3922 3285
rect 3956 3251 4105 3285
rect 3906 3245 4105 3251
rect 4139 3281 4173 3297
rect 4139 3209 4173 3247
rect 4207 3267 4223 3301
rect 4257 3277 4273 3301
rect 4808 3285 4842 3439
rect 5034 3423 5044 3439
rect 5034 3407 5078 3423
rect 4917 3379 4936 3405
rect 4917 3345 4927 3379
rect 4970 3371 4992 3405
rect 4961 3345 4992 3371
rect 5112 3348 5148 3575
rect 4917 3339 4992 3345
rect 5082 3345 5148 3348
rect 5082 3311 5098 3345
rect 5132 3311 5148 3345
rect 5182 3515 5284 3541
rect 5182 3481 5203 3515
rect 5237 3507 5284 3515
rect 5318 3507 5334 3541
rect 5182 3473 5237 3481
rect 5216 3439 5237 3473
rect 5397 3457 5431 3575
rect 5499 3606 5522 3640
rect 5465 3572 5522 3606
rect 5499 3538 5522 3572
rect 5465 3518 5522 3538
rect 5182 3377 5237 3439
rect 5288 3446 5363 3457
rect 5288 3412 5303 3446
rect 5337 3445 5363 3446
rect 5288 3411 5313 3412
rect 5347 3411 5363 3445
rect 5397 3441 5447 3457
rect 5397 3407 5413 3441
rect 5397 3391 5447 3407
rect 5182 3343 5320 3377
rect 4407 3277 4441 3285
rect 4257 3267 4441 3277
rect 4207 3243 4441 3267
rect 4495 3251 4511 3285
rect 4545 3251 4561 3285
rect 4495 3209 4561 3251
rect 4689 3251 4705 3285
rect 4739 3251 4842 3285
rect 4689 3245 4842 3251
rect 4878 3281 4930 3297
rect 4878 3247 4896 3281
rect 4878 3209 4930 3247
rect 4982 3267 4998 3301
rect 5032 3277 5048 3301
rect 5182 3293 5216 3309
rect 5032 3267 5182 3277
rect 4982 3259 5182 3267
rect 4982 3243 5216 3259
rect 5273 3295 5320 3343
rect 5273 3261 5286 3295
rect 5273 3245 5320 3261
rect 5365 3285 5431 3353
rect 5481 3335 5522 3518
rect 5365 3251 5381 3285
rect 5415 3251 5431 3285
rect 5365 3209 5431 3251
rect 5465 3319 5522 3335
rect 5499 3285 5522 3319
rect 5465 3243 5522 3285
rect 5556 3659 5619 3675
rect 5556 3625 5569 3659
rect 5603 3625 5619 3659
rect 5556 3591 5619 3625
rect 5556 3557 5569 3591
rect 5603 3557 5619 3591
rect 5556 3457 5619 3557
rect 5655 3665 5714 3719
rect 5655 3631 5664 3665
rect 5698 3631 5714 3665
rect 5655 3597 5714 3631
rect 5655 3563 5664 3597
rect 5698 3563 5714 3597
rect 5655 3545 5714 3563
rect 5748 3641 5800 3685
rect 5782 3607 5800 3641
rect 5748 3573 5800 3607
rect 5782 3539 5800 3573
rect 5834 3669 5886 3685
rect 5834 3635 5852 3669
rect 5834 3601 5886 3635
rect 5920 3653 5986 3719
rect 5920 3619 5936 3653
rect 5970 3619 5986 3653
rect 6020 3669 6065 3685
rect 6054 3635 6065 3669
rect 5834 3567 5852 3601
rect 6020 3601 6065 3635
rect 6104 3653 6174 3719
rect 6104 3619 6124 3653
rect 6158 3619 6174 3653
rect 6208 3669 6242 3685
rect 6285 3642 6301 3676
rect 6335 3642 6451 3676
rect 5886 3583 5985 3585
rect 5886 3567 5939 3583
rect 5834 3551 5939 3567
rect 5748 3481 5800 3539
rect 5973 3549 5985 3583
rect 5757 3471 5800 3481
rect 5834 3471 5905 3517
rect 5556 3441 5723 3457
rect 5556 3407 5689 3441
rect 5556 3391 5723 3407
rect 5757 3456 5905 3471
rect 5757 3423 5849 3456
rect 5556 3311 5619 3391
rect 5757 3357 5800 3423
rect 5834 3422 5849 3423
rect 5883 3422 5905 3456
rect 5834 3387 5905 3422
rect 5939 3456 5985 3549
rect 5939 3422 5951 3456
rect 5556 3277 5569 3311
rect 5603 3277 5619 3311
rect 5748 3321 5800 3357
rect 5939 3353 5985 3422
rect 5556 3243 5619 3277
rect 5655 3285 5714 3301
rect 5655 3251 5664 3285
rect 5698 3251 5714 3285
rect 5655 3209 5714 3251
rect 5782 3287 5800 3321
rect 5748 3243 5800 3287
rect 5834 3319 5985 3353
rect 6054 3567 6065 3601
rect 6208 3585 6242 3635
rect 6020 3379 6065 3567
rect 6020 3345 6031 3379
rect 5834 3311 5886 3319
rect 5834 3277 5852 3311
rect 6020 3311 6065 3345
rect 6099 3551 6242 3585
rect 6099 3357 6133 3551
rect 6283 3549 6307 3583
rect 6341 3557 6383 3583
rect 6341 3549 6349 3557
rect 6283 3523 6349 3549
rect 6167 3449 6249 3517
rect 6167 3443 6200 3449
rect 6234 3415 6249 3449
rect 6201 3409 6249 3415
rect 6167 3393 6249 3409
rect 6283 3507 6383 3523
rect 6283 3383 6327 3507
rect 6417 3473 6451 3642
rect 6499 3667 6575 3719
rect 6793 3677 6859 3719
rect 6499 3633 6515 3667
rect 6549 3633 6575 3667
rect 6635 3651 6669 3667
rect 6635 3599 6669 3617
rect 6793 3643 6809 3677
rect 6843 3643 6859 3677
rect 7282 3677 7358 3719
rect 6793 3609 6859 3643
rect 7068 3642 7084 3676
rect 7118 3642 7234 3676
rect 7282 3643 7298 3677
rect 7332 3643 7358 3677
rect 7546 3677 7823 3719
rect 7406 3651 7440 3667
rect 6485 3583 6755 3599
rect 6485 3557 6635 3583
rect 6519 3549 6635 3557
rect 6669 3549 6755 3583
rect 6793 3575 6809 3609
rect 6843 3575 6859 3609
rect 7030 3583 7077 3589
rect 6519 3523 6535 3549
rect 6485 3507 6535 3523
rect 6637 3473 6687 3489
rect 6417 3439 6653 3473
rect 6417 3431 6497 3439
rect 6099 3319 6242 3357
rect 6317 3349 6327 3383
rect 6283 3333 6327 3349
rect 6363 3361 6379 3395
rect 6413 3379 6429 3395
rect 6363 3345 6395 3361
rect 6363 3321 6429 3345
rect 5834 3261 5886 3277
rect 5920 3251 5936 3285
rect 5970 3251 5986 3285
rect 6054 3277 6065 3311
rect 6208 3303 6242 3319
rect 6020 3261 6065 3277
rect 5920 3209 5986 3251
rect 6104 3251 6124 3285
rect 6158 3251 6174 3285
rect 6463 3285 6497 3431
rect 6643 3423 6687 3439
rect 6721 3405 6755 3549
rect 7030 3557 7043 3583
rect 7064 3523 7077 3549
rect 6789 3515 6990 3523
rect 6789 3481 6951 3515
rect 6985 3481 6990 3515
rect 7030 3507 7077 3523
rect 7125 3557 7166 3573
rect 7125 3523 7132 3557
rect 6789 3475 6990 3481
rect 6789 3473 6855 3475
rect 6789 3439 6805 3473
rect 6839 3439 6855 3473
rect 7125 3453 7166 3523
rect 7042 3447 7166 3453
rect 6917 3405 6933 3439
rect 6967 3405 6983 3439
rect 6535 3371 6551 3405
rect 6585 3385 6601 3405
rect 6585 3379 6617 3385
rect 6535 3345 6583 3371
rect 6721 3371 6983 3405
rect 7042 3413 7043 3447
rect 7077 3417 7166 3447
rect 7200 3473 7234 3642
rect 7546 3643 7562 3677
rect 7596 3643 7773 3677
rect 7807 3643 7823 3677
rect 7406 3609 7440 3617
rect 7857 3640 7914 3685
rect 7268 3575 7823 3609
rect 7268 3557 7318 3575
rect 7302 3523 7318 3557
rect 7268 3507 7318 3523
rect 7200 3457 7470 3473
rect 7200 3439 7436 3457
rect 7077 3413 7099 3417
rect 7042 3383 7099 3413
rect 6721 3345 6765 3371
rect 6535 3339 6617 3345
rect 6699 3311 6715 3345
rect 6749 3311 6765 3345
rect 7042 3349 7065 3383
rect 6799 3319 6833 3335
rect 7042 3333 7099 3349
rect 6208 3253 6242 3269
rect 6104 3209 6174 3251
rect 6298 3251 6314 3285
rect 6348 3251 6497 3285
rect 6298 3245 6497 3251
rect 6531 3281 6565 3297
rect 6531 3209 6565 3247
rect 6599 3267 6615 3301
rect 6649 3277 6665 3301
rect 7200 3285 7234 3439
rect 7426 3423 7436 3439
rect 7426 3407 7470 3423
rect 7309 3379 7328 3405
rect 7309 3345 7319 3379
rect 7362 3371 7384 3405
rect 7353 3345 7384 3371
rect 7504 3348 7540 3575
rect 7309 3339 7384 3345
rect 7474 3345 7540 3348
rect 7474 3311 7490 3345
rect 7524 3311 7540 3345
rect 7574 3515 7676 3541
rect 7574 3481 7595 3515
rect 7629 3507 7676 3515
rect 7710 3507 7726 3541
rect 7574 3473 7629 3481
rect 7608 3439 7629 3473
rect 7789 3457 7823 3575
rect 7891 3606 7914 3640
rect 7857 3572 7914 3606
rect 7891 3538 7914 3572
rect 7857 3518 7914 3538
rect 7574 3377 7629 3439
rect 7680 3454 7755 3457
rect 7680 3420 7693 3454
rect 7727 3445 7755 3454
rect 7680 3411 7705 3420
rect 7739 3411 7755 3445
rect 7789 3441 7839 3457
rect 7789 3407 7805 3441
rect 7789 3391 7839 3407
rect 7574 3343 7712 3377
rect 6799 3277 6833 3285
rect 6649 3267 6833 3277
rect 6599 3243 6833 3267
rect 6887 3251 6903 3285
rect 6937 3251 6953 3285
rect 6887 3209 6953 3251
rect 7081 3251 7097 3285
rect 7131 3251 7234 3285
rect 7081 3245 7234 3251
rect 7270 3281 7322 3297
rect 7270 3247 7288 3281
rect 7270 3209 7322 3247
rect 7374 3267 7390 3301
rect 7424 3277 7440 3301
rect 7574 3293 7608 3309
rect 7424 3267 7574 3277
rect 7374 3259 7574 3267
rect 7374 3243 7608 3259
rect 7665 3295 7712 3343
rect 7665 3261 7678 3295
rect 7665 3245 7712 3261
rect 7757 3285 7823 3353
rect 7873 3335 7914 3518
rect 7757 3251 7773 3285
rect 7807 3251 7823 3285
rect 7757 3209 7823 3251
rect 7857 3319 7914 3335
rect 7891 3285 7914 3319
rect 7857 3243 7914 3285
rect 7948 3659 8011 3675
rect 7948 3625 7961 3659
rect 7995 3625 8011 3659
rect 7948 3591 8011 3625
rect 7948 3557 7961 3591
rect 7995 3557 8011 3591
rect 7948 3457 8011 3557
rect 8047 3665 8106 3719
rect 8047 3631 8056 3665
rect 8090 3631 8106 3665
rect 8047 3597 8106 3631
rect 8047 3563 8056 3597
rect 8090 3563 8106 3597
rect 8047 3545 8106 3563
rect 8140 3641 8192 3685
rect 8174 3607 8192 3641
rect 8140 3573 8192 3607
rect 8174 3539 8192 3573
rect 8226 3669 8278 3685
rect 8226 3635 8244 3669
rect 8226 3601 8278 3635
rect 8312 3653 8378 3719
rect 8312 3619 8328 3653
rect 8362 3619 8378 3653
rect 8412 3669 8457 3685
rect 8446 3635 8457 3669
rect 8226 3567 8244 3601
rect 8412 3601 8457 3635
rect 8496 3653 8566 3719
rect 8496 3619 8516 3653
rect 8550 3619 8566 3653
rect 8600 3669 8634 3685
rect 8677 3642 8693 3676
rect 8727 3642 8843 3676
rect 8278 3583 8377 3585
rect 8278 3567 8331 3583
rect 8226 3551 8331 3567
rect 8140 3481 8192 3539
rect 8365 3549 8377 3583
rect 8149 3472 8192 3481
rect 8226 3472 8297 3517
rect 7948 3441 8115 3457
rect 7948 3407 8081 3441
rect 7948 3391 8115 3407
rect 8149 3456 8297 3472
rect 8149 3424 8241 3456
rect 7948 3311 8011 3391
rect 8149 3357 8192 3424
rect 8226 3422 8241 3424
rect 8275 3422 8297 3456
rect 8226 3387 8297 3422
rect 8331 3456 8377 3549
rect 8331 3422 8343 3456
rect 7948 3277 7961 3311
rect 7995 3277 8011 3311
rect 8140 3347 8192 3357
rect 8331 3353 8377 3422
rect 8140 3321 8149 3347
rect 8183 3313 8192 3347
rect 7948 3243 8011 3277
rect 8047 3285 8106 3301
rect 8047 3251 8056 3285
rect 8090 3251 8106 3285
rect 8047 3209 8106 3251
rect 8174 3287 8192 3313
rect 8140 3243 8192 3287
rect 8226 3319 8377 3353
rect 8446 3567 8457 3601
rect 8600 3585 8634 3635
rect 8412 3379 8457 3567
rect 8412 3345 8423 3379
rect 8226 3311 8278 3319
rect 8226 3277 8244 3311
rect 8412 3311 8457 3345
rect 8491 3551 8634 3585
rect 8491 3357 8525 3551
rect 8675 3549 8699 3583
rect 8733 3557 8775 3583
rect 8733 3549 8741 3557
rect 8675 3523 8741 3549
rect 8559 3449 8641 3517
rect 8559 3443 8587 3449
rect 8621 3415 8641 3449
rect 8593 3409 8641 3415
rect 8559 3393 8641 3409
rect 8675 3507 8775 3523
rect 8675 3383 8719 3507
rect 8809 3473 8843 3642
rect 8891 3667 8967 3719
rect 9185 3677 9251 3719
rect 8891 3633 8907 3667
rect 8941 3633 8967 3667
rect 9027 3651 9061 3667
rect 9027 3599 9061 3617
rect 9185 3643 9201 3677
rect 9235 3643 9251 3677
rect 9674 3677 9750 3719
rect 9185 3609 9251 3643
rect 9460 3642 9476 3676
rect 9510 3642 9626 3676
rect 9674 3643 9690 3677
rect 9724 3643 9750 3677
rect 9938 3677 10215 3719
rect 9798 3651 9832 3667
rect 8877 3583 9147 3599
rect 8877 3557 9027 3583
rect 8911 3549 9027 3557
rect 9061 3549 9147 3583
rect 9185 3575 9201 3609
rect 9235 3575 9251 3609
rect 9422 3583 9469 3589
rect 8911 3523 8927 3549
rect 8877 3507 8927 3523
rect 9029 3473 9079 3489
rect 8809 3439 9045 3473
rect 8809 3431 8889 3439
rect 8491 3319 8634 3357
rect 8709 3349 8719 3383
rect 8675 3333 8719 3349
rect 8755 3361 8771 3395
rect 8805 3379 8821 3395
rect 8755 3345 8787 3361
rect 8755 3321 8821 3345
rect 8226 3261 8278 3277
rect 8312 3251 8328 3285
rect 8362 3251 8378 3285
rect 8446 3277 8457 3311
rect 8600 3303 8634 3319
rect 8412 3261 8457 3277
rect 8312 3209 8378 3251
rect 8496 3251 8516 3285
rect 8550 3251 8566 3285
rect 8855 3285 8889 3431
rect 9035 3423 9079 3439
rect 9113 3405 9147 3549
rect 9422 3557 9435 3583
rect 9456 3523 9469 3549
rect 9181 3515 9382 3523
rect 9181 3481 9343 3515
rect 9377 3481 9382 3515
rect 9422 3507 9469 3523
rect 9517 3557 9558 3573
rect 9517 3523 9524 3557
rect 9181 3475 9382 3481
rect 9181 3473 9247 3475
rect 9181 3439 9197 3473
rect 9231 3439 9247 3473
rect 9517 3453 9558 3523
rect 9434 3447 9558 3453
rect 9309 3405 9325 3439
rect 9359 3405 9375 3439
rect 8927 3371 8943 3405
rect 8977 3385 8993 3405
rect 8977 3379 9009 3385
rect 8927 3345 8975 3371
rect 9113 3371 9375 3405
rect 9434 3413 9435 3447
rect 9469 3417 9558 3447
rect 9592 3473 9626 3642
rect 9938 3643 9954 3677
rect 9988 3643 10165 3677
rect 10199 3643 10215 3677
rect 9798 3609 9832 3617
rect 10249 3640 10306 3685
rect 9660 3575 10215 3609
rect 9660 3557 9710 3575
rect 9694 3523 9710 3557
rect 9660 3507 9710 3523
rect 9592 3457 9862 3473
rect 9592 3439 9828 3457
rect 9469 3413 9491 3417
rect 9434 3383 9491 3413
rect 9113 3345 9157 3371
rect 8927 3339 9009 3345
rect 9091 3311 9107 3345
rect 9141 3311 9157 3345
rect 9434 3349 9457 3383
rect 9191 3319 9225 3335
rect 9434 3333 9491 3349
rect 8600 3253 8634 3269
rect 8496 3209 8566 3251
rect 8690 3251 8706 3285
rect 8740 3251 8889 3285
rect 8690 3245 8889 3251
rect 8923 3281 8957 3297
rect 8923 3209 8957 3247
rect 8991 3267 9007 3301
rect 9041 3277 9057 3301
rect 9592 3285 9626 3439
rect 9818 3423 9828 3439
rect 9818 3407 9862 3423
rect 9701 3379 9720 3405
rect 9701 3345 9711 3379
rect 9754 3371 9776 3405
rect 9745 3345 9776 3371
rect 9896 3348 9932 3575
rect 9701 3339 9776 3345
rect 9866 3345 9932 3348
rect 9866 3311 9882 3345
rect 9916 3311 9932 3345
rect 9966 3515 10068 3541
rect 9966 3481 9987 3515
rect 10021 3507 10068 3515
rect 10102 3507 10118 3541
rect 9966 3473 10021 3481
rect 10000 3439 10021 3473
rect 10181 3457 10215 3575
rect 10283 3606 10306 3640
rect 10249 3572 10306 3606
rect 10283 3538 10306 3572
rect 10249 3518 10306 3538
rect 9966 3377 10021 3439
rect 10072 3450 10147 3457
rect 10072 3416 10084 3450
rect 10118 3445 10147 3450
rect 10072 3411 10097 3416
rect 10131 3411 10147 3445
rect 10181 3441 10231 3457
rect 10181 3407 10197 3441
rect 10181 3391 10231 3407
rect 9966 3343 10104 3377
rect 9191 3277 9225 3285
rect 9041 3267 9225 3277
rect 8991 3243 9225 3267
rect 9279 3251 9295 3285
rect 9329 3251 9345 3285
rect 9279 3209 9345 3251
rect 9473 3251 9489 3285
rect 9523 3251 9626 3285
rect 9473 3245 9626 3251
rect 9662 3281 9714 3297
rect 9662 3247 9680 3281
rect 9662 3209 9714 3247
rect 9766 3267 9782 3301
rect 9816 3277 9832 3301
rect 9966 3293 10000 3309
rect 9816 3267 9966 3277
rect 9766 3259 9966 3267
rect 9766 3243 10000 3259
rect 10057 3295 10104 3343
rect 10057 3261 10070 3295
rect 10057 3245 10104 3261
rect 10149 3285 10215 3353
rect 10265 3335 10306 3518
rect 10149 3251 10165 3285
rect 10199 3251 10215 3285
rect 10149 3209 10215 3251
rect 10249 3319 10306 3335
rect 10283 3285 10306 3319
rect 10249 3243 10306 3285
rect 10340 3659 10403 3675
rect 10340 3625 10353 3659
rect 10387 3625 10403 3659
rect 10340 3591 10403 3625
rect 10340 3557 10353 3591
rect 10387 3557 10403 3591
rect 10340 3457 10403 3557
rect 10439 3665 10498 3719
rect 10439 3631 10448 3665
rect 10482 3631 10498 3665
rect 10439 3597 10498 3631
rect 10439 3563 10448 3597
rect 10482 3563 10498 3597
rect 10439 3545 10498 3563
rect 10532 3641 10584 3685
rect 10566 3607 10584 3641
rect 10532 3573 10584 3607
rect 10566 3539 10584 3573
rect 10618 3669 10670 3685
rect 10618 3635 10636 3669
rect 10618 3601 10670 3635
rect 10704 3653 10770 3719
rect 10704 3619 10720 3653
rect 10754 3619 10770 3653
rect 10804 3669 10849 3685
rect 10838 3635 10849 3669
rect 10618 3567 10636 3601
rect 10804 3601 10849 3635
rect 10888 3653 10958 3719
rect 10888 3619 10908 3653
rect 10942 3619 10958 3653
rect 10992 3669 11026 3685
rect 11069 3642 11085 3676
rect 11119 3642 11235 3676
rect 10670 3583 10769 3585
rect 10670 3567 10723 3583
rect 10618 3551 10723 3567
rect 10532 3481 10584 3539
rect 10757 3549 10769 3583
rect 10541 3463 10584 3481
rect 10618 3463 10689 3517
rect 10340 3441 10507 3457
rect 10340 3407 10473 3441
rect 10340 3391 10507 3407
rect 10541 3456 10689 3463
rect 10541 3422 10633 3456
rect 10667 3422 10689 3456
rect 10541 3415 10689 3422
rect 10340 3311 10403 3391
rect 10541 3357 10584 3415
rect 10618 3387 10689 3415
rect 10723 3456 10769 3549
rect 10723 3422 10735 3456
rect 10340 3277 10353 3311
rect 10387 3277 10403 3311
rect 10532 3348 10584 3357
rect 10723 3353 10769 3422
rect 10532 3321 10541 3348
rect 10575 3314 10584 3348
rect 10340 3243 10403 3277
rect 10439 3285 10498 3301
rect 10439 3251 10448 3285
rect 10482 3251 10498 3285
rect 10439 3209 10498 3251
rect 10566 3287 10584 3314
rect 10532 3243 10584 3287
rect 10618 3319 10769 3353
rect 10838 3567 10849 3601
rect 10992 3585 11026 3635
rect 10804 3379 10849 3567
rect 10804 3345 10815 3379
rect 10618 3311 10670 3319
rect 10618 3277 10636 3311
rect 10804 3311 10849 3345
rect 10883 3551 11026 3585
rect 10883 3357 10917 3551
rect 11067 3549 11091 3583
rect 11125 3557 11167 3583
rect 11125 3549 11133 3557
rect 11067 3523 11133 3549
rect 10951 3448 11033 3517
rect 10951 3443 10990 3448
rect 10985 3414 10990 3443
rect 11024 3414 11033 3448
rect 10985 3409 11033 3414
rect 10951 3393 11033 3409
rect 11067 3507 11167 3523
rect 11067 3383 11111 3507
rect 11201 3473 11235 3642
rect 11283 3667 11359 3719
rect 11577 3677 11643 3719
rect 11283 3633 11299 3667
rect 11333 3633 11359 3667
rect 11419 3651 11453 3667
rect 11419 3599 11453 3617
rect 11577 3643 11593 3677
rect 11627 3643 11643 3677
rect 12066 3677 12142 3719
rect 11577 3609 11643 3643
rect 11852 3642 11868 3676
rect 11902 3642 12018 3676
rect 12066 3643 12082 3677
rect 12116 3643 12142 3677
rect 12330 3677 12607 3719
rect 12190 3651 12224 3667
rect 11269 3583 11539 3599
rect 11269 3557 11419 3583
rect 11303 3549 11419 3557
rect 11453 3549 11539 3583
rect 11577 3575 11593 3609
rect 11627 3575 11643 3609
rect 11814 3583 11861 3589
rect 11303 3523 11319 3549
rect 11269 3507 11319 3523
rect 11421 3473 11471 3489
rect 11201 3439 11437 3473
rect 11201 3431 11281 3439
rect 10883 3319 11026 3357
rect 11101 3349 11111 3383
rect 11067 3333 11111 3349
rect 11147 3361 11163 3395
rect 11197 3379 11213 3395
rect 11147 3345 11179 3361
rect 11147 3321 11213 3345
rect 10618 3261 10670 3277
rect 10704 3251 10720 3285
rect 10754 3251 10770 3285
rect 10838 3277 10849 3311
rect 10992 3303 11026 3319
rect 10804 3261 10849 3277
rect 10704 3209 10770 3251
rect 10888 3251 10908 3285
rect 10942 3251 10958 3285
rect 11247 3285 11281 3431
rect 11427 3423 11471 3439
rect 11505 3405 11539 3549
rect 11814 3557 11827 3583
rect 11848 3523 11861 3549
rect 11573 3515 11774 3523
rect 11573 3481 11735 3515
rect 11769 3481 11774 3515
rect 11814 3507 11861 3523
rect 11909 3557 11950 3573
rect 11909 3523 11916 3557
rect 11573 3475 11774 3481
rect 11573 3473 11639 3475
rect 11573 3439 11589 3473
rect 11623 3439 11639 3473
rect 11909 3453 11950 3523
rect 11826 3447 11950 3453
rect 11701 3405 11717 3439
rect 11751 3405 11767 3439
rect 11319 3371 11335 3405
rect 11369 3385 11385 3405
rect 11369 3379 11401 3385
rect 11319 3345 11367 3371
rect 11505 3371 11767 3405
rect 11826 3413 11827 3447
rect 11861 3417 11950 3447
rect 11984 3473 12018 3642
rect 12330 3643 12346 3677
rect 12380 3643 12557 3677
rect 12591 3643 12607 3677
rect 12190 3609 12224 3617
rect 12641 3640 12698 3685
rect 12052 3575 12607 3609
rect 12052 3557 12102 3575
rect 12086 3523 12102 3557
rect 12052 3507 12102 3523
rect 11984 3457 12254 3473
rect 11984 3439 12220 3457
rect 11861 3413 11883 3417
rect 11826 3383 11883 3413
rect 11505 3345 11549 3371
rect 11319 3339 11401 3345
rect 11483 3311 11499 3345
rect 11533 3311 11549 3345
rect 11826 3349 11849 3383
rect 11583 3319 11617 3335
rect 11826 3333 11883 3349
rect 10992 3253 11026 3269
rect 10888 3209 10958 3251
rect 11082 3251 11098 3285
rect 11132 3251 11281 3285
rect 11082 3245 11281 3251
rect 11315 3281 11349 3297
rect 11315 3209 11349 3247
rect 11383 3267 11399 3301
rect 11433 3277 11449 3301
rect 11984 3285 12018 3439
rect 12210 3423 12220 3439
rect 12210 3407 12254 3423
rect 12093 3379 12112 3405
rect 12093 3345 12103 3379
rect 12146 3371 12168 3405
rect 12137 3345 12168 3371
rect 12288 3348 12324 3575
rect 12093 3339 12168 3345
rect 12258 3345 12324 3348
rect 12258 3311 12274 3345
rect 12308 3311 12324 3345
rect 12358 3515 12460 3541
rect 12358 3481 12379 3515
rect 12413 3507 12460 3515
rect 12494 3507 12510 3541
rect 12358 3473 12413 3481
rect 12392 3439 12413 3473
rect 12573 3457 12607 3575
rect 12675 3606 12698 3640
rect 12641 3572 12698 3606
rect 12675 3538 12698 3572
rect 12641 3518 12698 3538
rect 12358 3377 12413 3439
rect 12464 3449 12539 3457
rect 12464 3415 12476 3449
rect 12510 3445 12539 3449
rect 12464 3411 12489 3415
rect 12523 3411 12539 3445
rect 12573 3441 12623 3457
rect 12573 3407 12589 3441
rect 12573 3391 12623 3407
rect 12358 3343 12496 3377
rect 11583 3277 11617 3285
rect 11433 3267 11617 3277
rect 11383 3243 11617 3267
rect 11671 3251 11687 3285
rect 11721 3251 11737 3285
rect 11671 3209 11737 3251
rect 11865 3251 11881 3285
rect 11915 3251 12018 3285
rect 11865 3245 12018 3251
rect 12054 3281 12106 3297
rect 12054 3247 12072 3281
rect 12054 3209 12106 3247
rect 12158 3267 12174 3301
rect 12208 3277 12224 3301
rect 12358 3293 12392 3309
rect 12208 3267 12358 3277
rect 12158 3259 12358 3267
rect 12158 3243 12392 3259
rect 12449 3295 12496 3343
rect 12449 3261 12462 3295
rect 12449 3245 12496 3261
rect 12541 3285 12607 3353
rect 12657 3335 12698 3518
rect 12541 3251 12557 3285
rect 12591 3251 12607 3285
rect 12541 3209 12607 3251
rect 12641 3319 12698 3335
rect 12675 3285 12698 3319
rect 12641 3243 12698 3285
rect 12732 3659 12795 3675
rect 12732 3625 12745 3659
rect 12779 3625 12795 3659
rect 12732 3591 12795 3625
rect 12732 3557 12745 3591
rect 12779 3557 12795 3591
rect 12732 3457 12795 3557
rect 12831 3665 12890 3719
rect 12831 3631 12840 3665
rect 12874 3631 12890 3665
rect 12831 3597 12890 3631
rect 12831 3563 12840 3597
rect 12874 3563 12890 3597
rect 12831 3545 12890 3563
rect 12924 3641 12976 3685
rect 12958 3607 12976 3641
rect 12924 3573 12976 3607
rect 12958 3539 12976 3573
rect 12924 3481 12976 3539
rect 12732 3441 12899 3457
rect 12732 3407 12865 3441
rect 12732 3391 12899 3407
rect 12732 3311 12795 3391
rect 12933 3357 12976 3481
rect 12732 3277 12745 3311
rect 12779 3277 12795 3311
rect 12924 3351 12976 3357
rect 12924 3321 12931 3351
rect 12965 3317 12976 3351
rect 12732 3243 12795 3277
rect 12831 3285 12890 3301
rect 12831 3251 12840 3285
rect 12874 3251 12890 3285
rect 12831 3209 12890 3251
rect 12958 3287 12976 3317
rect 12924 3243 12976 3287
rect 626 3174 655 3208
rect 689 3174 747 3208
rect 781 3174 839 3208
rect 873 3174 931 3208
rect 965 3174 1023 3208
rect 1057 3174 1115 3208
rect 1149 3174 1207 3208
rect 1241 3174 1299 3208
rect 1333 3174 1391 3208
rect 1425 3174 1454 3208
rect 3168 3185 3197 3209
rect 626 3173 1454 3174
rect 626 3139 654 3173
rect 688 3139 747 3173
rect 781 3139 839 3173
rect 873 3139 931 3173
rect 965 3139 1023 3173
rect 1057 3139 1115 3173
rect 1149 3139 1207 3173
rect 1241 3139 1299 3173
rect 1333 3139 1391 3173
rect 1425 3139 1454 3173
rect 3167 3151 3197 3185
rect 3231 3151 3289 3209
rect 3323 3151 3381 3209
rect 3415 3175 3454 3209
rect 3488 3185 3546 3209
rect 3580 3185 3638 3209
rect 3672 3185 3730 3209
rect 3764 3185 3822 3209
rect 3856 3185 3914 3209
rect 3948 3185 4006 3209
rect 4040 3185 4098 3209
rect 4132 3185 4190 3209
rect 4224 3185 4282 3209
rect 4316 3185 4374 3209
rect 4408 3185 4466 3209
rect 4500 3185 4558 3209
rect 4592 3185 4650 3209
rect 4684 3185 4742 3209
rect 4776 3185 4834 3209
rect 4868 3185 4926 3209
rect 4960 3185 5018 3209
rect 5052 3185 5110 3209
rect 5144 3185 5202 3209
rect 5236 3185 5294 3209
rect 5328 3185 5386 3209
rect 5420 3185 5478 3209
rect 5512 3185 5570 3209
rect 5604 3185 5662 3209
rect 5696 3185 5754 3209
rect 5788 3185 5846 3209
rect 5880 3185 5938 3209
rect 5972 3185 6030 3209
rect 6064 3185 6122 3209
rect 6156 3185 6214 3209
rect 6248 3185 6306 3209
rect 6340 3185 6398 3209
rect 6432 3185 6490 3209
rect 6524 3185 6582 3209
rect 6616 3185 6674 3209
rect 6708 3185 6766 3209
rect 6800 3185 6858 3209
rect 6892 3185 6950 3209
rect 6984 3185 7042 3209
rect 7076 3185 7134 3209
rect 7168 3185 7226 3209
rect 7260 3185 7318 3209
rect 7352 3185 7410 3209
rect 7444 3185 7502 3209
rect 7536 3185 7594 3209
rect 7628 3185 7686 3209
rect 7720 3185 7778 3209
rect 7812 3185 7870 3209
rect 7904 3185 7962 3209
rect 7996 3185 8054 3209
rect 8088 3185 8146 3209
rect 8180 3185 8238 3209
rect 8272 3185 8330 3209
rect 8364 3185 8422 3209
rect 8456 3185 8514 3209
rect 8548 3185 8606 3209
rect 8640 3185 8698 3209
rect 8732 3185 8790 3209
rect 8824 3185 8882 3209
rect 8916 3185 8974 3209
rect 9008 3185 9066 3209
rect 9100 3185 9158 3209
rect 9192 3185 9250 3209
rect 9284 3185 9342 3209
rect 9376 3185 9434 3209
rect 9468 3185 9526 3209
rect 9560 3185 9618 3209
rect 9652 3185 9710 3209
rect 9744 3185 9802 3209
rect 9836 3185 9894 3209
rect 9928 3185 9986 3209
rect 10020 3185 10078 3209
rect 10112 3185 10170 3209
rect 10204 3185 10262 3209
rect 10296 3185 10354 3209
rect 10388 3185 10446 3209
rect 10480 3185 10538 3209
rect 10572 3185 10630 3209
rect 10664 3185 10722 3209
rect 10756 3185 10814 3209
rect 10848 3185 10906 3209
rect 10940 3185 10998 3209
rect 11032 3185 11090 3209
rect 11124 3185 11182 3209
rect 11216 3185 11274 3209
rect 11308 3185 11366 3209
rect 11400 3185 11458 3209
rect 11492 3185 11550 3209
rect 11584 3185 11642 3209
rect 11676 3185 11734 3209
rect 11768 3185 11826 3209
rect 11860 3185 11918 3209
rect 11952 3185 12010 3209
rect 3507 3175 3546 3185
rect 3599 3175 3638 3185
rect 3691 3175 3730 3185
rect 3783 3175 3822 3185
rect 3875 3175 3914 3185
rect 3967 3175 4006 3185
rect 4059 3175 4098 3185
rect 4151 3175 4190 3185
rect 4243 3175 4282 3185
rect 4335 3175 4374 3185
rect 4427 3175 4466 3185
rect 4519 3175 4558 3185
rect 4611 3175 4650 3185
rect 4703 3175 4742 3185
rect 4795 3175 4834 3185
rect 4887 3175 4926 3185
rect 4979 3175 5018 3185
rect 5071 3175 5110 3185
rect 5163 3175 5202 3185
rect 5255 3175 5294 3185
rect 5347 3175 5386 3185
rect 5439 3175 5478 3185
rect 5531 3175 5570 3185
rect 5623 3175 5662 3185
rect 5715 3175 5754 3185
rect 5807 3175 5846 3185
rect 5899 3175 5938 3185
rect 5991 3175 6030 3185
rect 6083 3175 6122 3185
rect 6175 3175 6214 3185
rect 6267 3175 6306 3185
rect 6359 3175 6398 3185
rect 6451 3175 6490 3185
rect 6543 3175 6582 3185
rect 6635 3175 6674 3185
rect 6727 3175 6766 3185
rect 6819 3175 6858 3185
rect 6911 3175 6950 3185
rect 7003 3175 7042 3185
rect 7095 3175 7134 3185
rect 7187 3175 7226 3185
rect 7279 3175 7318 3185
rect 7371 3175 7410 3185
rect 7463 3175 7502 3185
rect 7555 3175 7594 3185
rect 7647 3175 7686 3185
rect 7739 3175 7778 3185
rect 7831 3175 7870 3185
rect 7923 3175 7962 3185
rect 8015 3175 8054 3185
rect 8107 3175 8146 3185
rect 8199 3175 8238 3185
rect 8291 3175 8330 3185
rect 8383 3175 8422 3185
rect 8475 3175 8514 3185
rect 8567 3175 8606 3185
rect 8659 3175 8698 3185
rect 8751 3175 8790 3185
rect 8843 3175 8882 3185
rect 8935 3175 8974 3185
rect 9027 3175 9066 3185
rect 9119 3175 9158 3185
rect 9211 3175 9250 3185
rect 9303 3175 9342 3185
rect 9395 3175 9434 3185
rect 9487 3175 9526 3185
rect 9579 3175 9618 3185
rect 9671 3175 9710 3185
rect 9763 3175 9802 3185
rect 3415 3151 3473 3175
rect 3507 3151 3565 3175
rect 3599 3151 3657 3175
rect 3691 3151 3749 3175
rect 3783 3151 3841 3175
rect 3875 3151 3933 3175
rect 3967 3151 4025 3175
rect 4059 3151 4117 3175
rect 4151 3151 4209 3175
rect 4243 3151 4301 3175
rect 4335 3151 4393 3175
rect 4427 3151 4485 3175
rect 4519 3151 4577 3175
rect 4611 3151 4669 3175
rect 4703 3151 4761 3175
rect 4795 3151 4853 3175
rect 4887 3151 4945 3175
rect 4979 3151 5037 3175
rect 5071 3151 5129 3175
rect 5163 3151 5221 3175
rect 5255 3151 5313 3175
rect 5347 3151 5405 3175
rect 5439 3151 5497 3175
rect 5531 3151 5589 3175
rect 5623 3151 5681 3175
rect 5715 3151 5773 3175
rect 5807 3151 5865 3175
rect 5899 3151 5957 3175
rect 5991 3151 6049 3175
rect 6083 3151 6141 3175
rect 6175 3151 6233 3175
rect 6267 3151 6325 3175
rect 6359 3151 6417 3175
rect 6451 3151 6509 3175
rect 6543 3151 6601 3175
rect 6635 3151 6693 3175
rect 6727 3151 6785 3175
rect 6819 3151 6877 3175
rect 6911 3151 6969 3175
rect 7003 3151 7061 3175
rect 7095 3151 7153 3175
rect 7187 3151 7245 3175
rect 7279 3151 7337 3175
rect 7371 3151 7429 3175
rect 7463 3151 7521 3175
rect 7555 3151 7613 3175
rect 7647 3151 7705 3175
rect 7739 3151 7797 3175
rect 7831 3151 7889 3175
rect 7923 3151 7981 3175
rect 8015 3151 8073 3175
rect 8107 3151 8165 3175
rect 8199 3151 8257 3175
rect 8291 3151 8349 3175
rect 8383 3151 8441 3175
rect 8475 3151 8533 3175
rect 8567 3151 8625 3175
rect 8659 3151 8717 3175
rect 8751 3151 8809 3175
rect 8843 3151 8901 3175
rect 8935 3151 8993 3175
rect 9027 3151 9085 3175
rect 9119 3151 9177 3175
rect 9211 3151 9269 3175
rect 9303 3151 9361 3175
rect 9395 3151 9453 3175
rect 9487 3151 9545 3175
rect 9579 3151 9637 3175
rect 9671 3151 9729 3175
rect 9763 3151 9821 3175
rect 9855 3151 9894 3185
rect 9947 3151 9986 3185
rect 10039 3151 10078 3185
rect 10131 3151 10170 3185
rect 10223 3151 10262 3185
rect 10315 3151 10354 3185
rect 10407 3151 10446 3185
rect 10499 3151 10538 3185
rect 10591 3151 10630 3185
rect 10683 3151 10722 3185
rect 10775 3151 10814 3185
rect 10867 3151 10906 3185
rect 10959 3151 10998 3185
rect 11051 3151 11090 3185
rect 11143 3151 11182 3185
rect 11235 3151 11274 3185
rect 11327 3151 11366 3185
rect 11419 3151 11458 3185
rect 11511 3151 11550 3185
rect 11603 3151 11642 3185
rect 11695 3151 11734 3185
rect 11787 3151 11826 3185
rect 11879 3151 11918 3185
rect 11971 3151 12010 3185
rect 12044 3151 12102 3209
rect 12136 3151 12194 3209
rect 12228 3151 12286 3209
rect 12320 3151 12378 3209
rect 12412 3151 12470 3209
rect 12504 3151 12562 3209
rect 12596 3151 12654 3209
rect 12688 3151 12746 3209
rect 12780 3151 12838 3209
rect 12872 3151 12930 3209
rect 12964 3175 12993 3209
rect 12964 3151 12992 3175
rect 1033 2846 1062 2904
rect 1096 2846 1154 2904
rect 1188 2846 1246 2904
rect 1280 2846 1338 2904
rect 1372 2846 1430 2904
rect 1464 2846 1522 2904
rect 1556 2846 1614 2904
rect 1648 2846 1706 2904
rect 1740 2846 1798 2904
rect 1832 2846 1890 2904
rect 1924 2846 1982 2904
rect 2016 2846 2074 2904
rect 2108 2846 2166 2904
rect 2200 2846 2258 2904
rect 2292 2846 2350 2904
rect 2384 2846 2442 2904
rect 2476 2846 2534 2904
rect 2568 2846 2626 2904
rect 2660 2846 2718 2904
rect 2752 2846 2810 2904
rect 2844 2846 2902 2904
rect 2936 2846 2994 2904
rect 3028 2846 3086 2904
rect 3120 2846 3178 2904
rect 3212 2846 3270 2904
rect 3304 2846 3362 2904
rect 3396 2846 3454 2904
rect 3488 2846 3546 2904
rect 3580 2846 3638 2904
rect 3672 2846 3730 2904
rect 3764 2846 3822 2904
rect 3856 2846 3914 2904
rect 3948 2846 4006 2904
rect 4040 2846 4098 2904
rect 4132 2846 4190 2904
rect 4224 2846 4282 2904
rect 4316 2846 4374 2904
rect 4408 2846 4466 2904
rect 4500 2846 4558 2904
rect 4592 2846 4650 2904
rect 4684 2846 4742 2904
rect 4776 2846 4834 2904
rect 4868 2846 4926 2904
rect 4960 2846 5018 2904
rect 5052 2846 5110 2904
rect 5144 2846 5202 2904
rect 5236 2846 5294 2904
rect 5328 2846 5386 2904
rect 5420 2846 5478 2904
rect 5512 2846 5570 2904
rect 5604 2846 5662 2904
rect 5696 2846 5754 2904
rect 5788 2846 5846 2904
rect 5880 2846 5938 2904
rect 5972 2846 6030 2904
rect 6064 2846 6122 2904
rect 6156 2846 6214 2904
rect 6248 2846 6306 2904
rect 6340 2846 6398 2904
rect 6432 2846 6490 2904
rect 6524 2846 6582 2904
rect 6616 2846 6674 2904
rect 6708 2846 6766 2904
rect 6800 2846 6858 2904
rect 6892 2846 6950 2904
rect 6984 2846 7042 2904
rect 7076 2846 7134 2904
rect 7168 2846 7226 2904
rect 7260 2846 7318 2904
rect 7352 2846 7410 2904
rect 7444 2846 7502 2904
rect 7536 2846 7594 2904
rect 7628 2846 7686 2904
rect 7720 2846 7778 2904
rect 7812 2846 7870 2904
rect 7904 2846 7962 2904
rect 7996 2846 8054 2904
rect 8088 2846 8146 2904
rect 8180 2846 8238 2904
rect 8272 2846 8330 2904
rect 8364 2846 8422 2904
rect 8456 2846 8514 2904
rect 8548 2846 8606 2904
rect 8640 2846 8698 2904
rect 8732 2846 8790 2904
rect 8824 2846 8882 2904
rect 8916 2846 8974 2904
rect 9008 2846 9066 2904
rect 9100 2846 9158 2904
rect 9192 2846 9250 2904
rect 9284 2846 9342 2904
rect 9376 2846 9434 2904
rect 9468 2846 9526 2904
rect 9560 2846 9618 2904
rect 9652 2846 9710 2904
rect 9744 2846 9802 2904
rect 9836 2846 9894 2904
rect 9928 2846 9986 2904
rect 10020 2846 10078 2904
rect 10112 2846 10170 2904
rect 10204 2846 10262 2904
rect 10296 2846 10354 2904
rect 10388 2846 10446 2904
rect 10480 2846 10538 2904
rect 10572 2846 10630 2904
rect 10664 2846 10722 2904
rect 10756 2846 10814 2904
rect 10848 2846 10906 2904
rect 10940 2846 10998 2904
rect 11032 2846 11090 2904
rect 11124 2846 11182 2904
rect 11216 2846 11274 2904
rect 11308 2846 11366 2904
rect 11400 2846 11458 2904
rect 11492 2846 11550 2904
rect 11584 2846 11642 2904
rect 11676 2846 11734 2904
rect 11768 2846 11826 2904
rect 11860 2846 11918 2904
rect 11952 2846 12010 2904
rect 12044 2846 12102 2904
rect 12136 2846 12194 2904
rect 12228 2846 12286 2904
rect 12320 2846 12378 2904
rect 12412 2846 12470 2904
rect 12504 2846 12562 2904
rect 12596 2846 12654 2904
rect 12688 2846 12746 2904
rect 12780 2846 12838 2904
rect 12872 2846 12930 2904
rect 12964 2846 12993 2904
rect 1050 2768 1102 2812
rect 1050 2734 1068 2768
rect 1050 2700 1102 2734
rect 1050 2666 1068 2700
rect 1136 2792 1195 2846
rect 1136 2758 1152 2792
rect 1186 2758 1195 2792
rect 1136 2724 1195 2758
rect 1136 2690 1152 2724
rect 1186 2690 1195 2724
rect 1136 2672 1195 2690
rect 1231 2786 1294 2802
rect 1231 2752 1247 2786
rect 1281 2752 1294 2786
rect 1231 2718 1294 2752
rect 1231 2684 1247 2718
rect 1281 2684 1294 2718
rect 1050 2608 1102 2666
rect 1050 2484 1093 2608
rect 1231 2584 1294 2684
rect 1127 2568 1294 2584
rect 1161 2534 1294 2568
rect 1127 2518 1294 2534
rect 1050 2448 1102 2484
rect 1050 2447 1068 2448
rect 1050 2413 1059 2447
rect 1231 2438 1294 2518
rect 1093 2413 1102 2414
rect 1050 2370 1102 2413
rect 1136 2412 1195 2428
rect 1136 2378 1152 2412
rect 1186 2378 1195 2412
rect 1136 2336 1195 2378
rect 1231 2404 1247 2438
rect 1281 2404 1294 2438
rect 1231 2370 1294 2404
rect 1328 2767 1385 2812
rect 1419 2804 1696 2846
rect 1419 2770 1435 2804
rect 1469 2770 1646 2804
rect 1680 2770 1696 2804
rect 1884 2804 1960 2846
rect 1802 2778 1836 2794
rect 1328 2733 1351 2767
rect 1884 2770 1910 2804
rect 1944 2770 1960 2804
rect 2383 2804 2449 2846
rect 1802 2736 1836 2744
rect 2008 2769 2124 2803
rect 2158 2769 2174 2803
rect 2383 2770 2399 2804
rect 2433 2770 2449 2804
rect 2667 2794 2743 2846
rect 1328 2699 1385 2733
rect 1328 2665 1351 2699
rect 1328 2645 1385 2665
rect 1419 2702 1974 2736
rect 1328 2462 1369 2645
rect 1419 2584 1453 2702
rect 1516 2634 1532 2668
rect 1566 2642 1668 2668
rect 1566 2634 1613 2642
rect 1647 2608 1668 2642
rect 1613 2600 1668 2608
rect 1403 2568 1453 2584
rect 1437 2534 1453 2568
rect 1487 2572 1562 2584
rect 1487 2538 1503 2572
rect 1537 2538 1562 2572
rect 1613 2566 1634 2600
rect 1403 2518 1453 2534
rect 1613 2504 1668 2566
rect 1328 2446 1385 2462
rect 1328 2412 1351 2446
rect 1328 2370 1385 2412
rect 1419 2412 1485 2480
rect 1419 2378 1435 2412
rect 1469 2378 1485 2412
rect 1419 2336 1485 2378
rect 1530 2470 1668 2504
rect 1702 2475 1738 2702
rect 1924 2684 1974 2702
rect 1924 2650 1940 2684
rect 1924 2634 1974 2650
rect 2008 2600 2042 2769
rect 2383 2736 2449 2770
rect 2165 2710 2212 2716
rect 1772 2584 2042 2600
rect 1806 2566 2042 2584
rect 1806 2550 1816 2566
rect 1772 2534 1816 2550
rect 1858 2498 1880 2532
rect 1914 2506 1933 2532
rect 1702 2472 1768 2475
rect 1530 2422 1577 2470
rect 1702 2438 1718 2472
rect 1752 2438 1768 2472
rect 1858 2472 1889 2498
rect 1923 2472 1933 2506
rect 1858 2466 1933 2472
rect 1564 2388 1577 2422
rect 1530 2372 1577 2388
rect 1634 2420 1668 2436
rect 1802 2404 1818 2428
rect 1668 2394 1818 2404
rect 1852 2394 1868 2428
rect 1668 2386 1868 2394
rect 1634 2370 1868 2386
rect 1920 2408 1972 2424
rect 1954 2374 1972 2408
rect 1920 2336 1972 2374
rect 2008 2412 2042 2566
rect 2076 2684 2117 2700
rect 2110 2650 2117 2684
rect 2076 2580 2117 2650
rect 2199 2684 2212 2710
rect 2383 2702 2399 2736
rect 2433 2702 2449 2736
rect 2573 2778 2607 2794
rect 2667 2760 2693 2794
rect 2727 2760 2743 2794
rect 2791 2769 2907 2803
rect 2941 2769 2957 2803
rect 3000 2796 3034 2812
rect 2573 2726 2607 2744
rect 2487 2710 2757 2726
rect 2165 2650 2178 2676
rect 2487 2676 2573 2710
rect 2607 2684 2757 2710
rect 2607 2676 2723 2684
rect 2165 2634 2212 2650
rect 2252 2642 2453 2650
rect 2252 2608 2257 2642
rect 2291 2608 2453 2642
rect 2252 2602 2453 2608
rect 2387 2600 2453 2602
rect 2076 2574 2200 2580
rect 2076 2544 2165 2574
rect 2143 2540 2165 2544
rect 2199 2540 2200 2574
rect 2387 2566 2403 2600
rect 2437 2566 2453 2600
rect 2143 2510 2200 2540
rect 2177 2476 2200 2510
rect 2259 2532 2275 2566
rect 2309 2532 2325 2566
rect 2487 2532 2521 2676
rect 2707 2650 2723 2676
rect 2707 2634 2757 2650
rect 2555 2600 2605 2616
rect 2791 2600 2825 2769
rect 3000 2712 3034 2762
rect 3068 2780 3138 2846
rect 3068 2746 3084 2780
rect 3118 2746 3138 2780
rect 3177 2796 3222 2812
rect 3177 2762 3188 2796
rect 3177 2728 3222 2762
rect 3256 2780 3322 2846
rect 3256 2746 3272 2780
rect 3306 2746 3322 2780
rect 3356 2796 3408 2812
rect 3390 2762 3408 2796
rect 2859 2684 2901 2710
rect 2893 2676 2901 2684
rect 2935 2676 2959 2710
rect 3000 2678 3143 2712
rect 2893 2650 2959 2676
rect 2859 2634 2959 2650
rect 2589 2566 2825 2600
rect 2555 2550 2599 2566
rect 2745 2558 2825 2566
rect 2259 2498 2521 2532
rect 2641 2512 2657 2532
rect 2143 2460 2200 2476
rect 2477 2472 2521 2498
rect 2625 2506 2657 2512
rect 2691 2498 2707 2532
rect 2659 2472 2707 2498
rect 2409 2446 2443 2462
rect 2477 2438 2493 2472
rect 2527 2438 2543 2472
rect 2625 2466 2707 2472
rect 2008 2378 2111 2412
rect 2145 2378 2161 2412
rect 2008 2372 2161 2378
rect 2289 2378 2305 2412
rect 2339 2378 2355 2412
rect 2289 2336 2355 2378
rect 2409 2404 2443 2412
rect 2577 2404 2593 2428
rect 2409 2394 2593 2404
rect 2627 2394 2643 2428
rect 2409 2370 2643 2394
rect 2677 2408 2711 2424
rect 2677 2336 2711 2374
rect 2745 2412 2779 2558
rect 2813 2506 2829 2522
rect 2863 2488 2879 2522
rect 2847 2472 2879 2488
rect 2813 2448 2879 2472
rect 2915 2510 2959 2634
rect 2993 2632 3075 2644
rect 2993 2598 3015 2632
rect 3049 2598 3075 2632
rect 2993 2570 3075 2598
rect 2993 2536 3041 2570
rect 2993 2520 3075 2536
rect 2915 2476 2925 2510
rect 3109 2484 3143 2678
rect 2915 2460 2959 2476
rect 3000 2446 3143 2484
rect 3177 2694 3188 2728
rect 3356 2728 3408 2762
rect 3177 2506 3222 2694
rect 3211 2472 3222 2506
rect 3000 2430 3034 2446
rect 2745 2378 2894 2412
rect 2928 2378 2944 2412
rect 3177 2438 3222 2472
rect 3257 2710 3356 2712
rect 3257 2676 3269 2710
rect 3303 2694 3356 2710
rect 3390 2694 3408 2728
rect 3303 2678 3408 2694
rect 3442 2768 3494 2812
rect 3442 2734 3460 2768
rect 3442 2700 3494 2734
rect 3257 2583 3303 2676
rect 3442 2666 3460 2700
rect 3528 2792 3587 2846
rect 3528 2758 3544 2792
rect 3578 2758 3587 2792
rect 3528 2724 3587 2758
rect 3528 2690 3544 2724
rect 3578 2690 3587 2724
rect 3528 2672 3587 2690
rect 3623 2786 3686 2802
rect 3623 2752 3639 2786
rect 3673 2752 3686 2786
rect 3623 2718 3686 2752
rect 3623 2684 3639 2718
rect 3673 2684 3686 2718
rect 3291 2549 3303 2583
rect 3257 2480 3303 2549
rect 3337 2583 3408 2644
rect 3337 2549 3359 2583
rect 3393 2582 3408 2583
rect 3442 2608 3494 2666
rect 3442 2582 3485 2608
rect 3623 2584 3686 2684
rect 3393 2549 3485 2582
rect 3337 2534 3485 2549
rect 3337 2514 3408 2534
rect 3442 2484 3485 2534
rect 3519 2568 3686 2584
rect 3553 2534 3686 2568
rect 3519 2518 3686 2534
rect 3257 2446 3408 2480
rect 3000 2380 3034 2396
rect 2745 2372 2944 2378
rect 3068 2378 3084 2412
rect 3118 2378 3138 2412
rect 3177 2404 3188 2438
rect 3356 2438 3408 2446
rect 3177 2388 3222 2404
rect 3068 2336 3138 2378
rect 3256 2378 3272 2412
rect 3306 2378 3322 2412
rect 3390 2404 3408 2438
rect 3356 2388 3408 2404
rect 3442 2470 3494 2484
rect 3442 2436 3450 2470
rect 3484 2448 3494 2470
rect 3442 2414 3460 2436
rect 3623 2438 3686 2518
rect 3256 2336 3322 2378
rect 3442 2370 3494 2414
rect 3528 2412 3587 2428
rect 3528 2378 3544 2412
rect 3578 2378 3587 2412
rect 3528 2336 3587 2378
rect 3623 2404 3639 2438
rect 3673 2404 3686 2438
rect 3623 2370 3686 2404
rect 3720 2767 3777 2812
rect 3811 2804 4088 2846
rect 3811 2770 3827 2804
rect 3861 2770 4038 2804
rect 4072 2770 4088 2804
rect 4276 2804 4352 2846
rect 4194 2778 4228 2794
rect 3720 2733 3743 2767
rect 4276 2770 4302 2804
rect 4336 2770 4352 2804
rect 4775 2804 4841 2846
rect 4194 2736 4228 2744
rect 4400 2769 4516 2803
rect 4550 2769 4566 2803
rect 4775 2770 4791 2804
rect 4825 2770 4841 2804
rect 5059 2794 5135 2846
rect 3720 2699 3777 2733
rect 3720 2665 3743 2699
rect 3720 2645 3777 2665
rect 3811 2702 4366 2736
rect 3720 2462 3761 2645
rect 3811 2584 3845 2702
rect 3908 2634 3924 2668
rect 3958 2642 4060 2668
rect 3958 2634 4005 2642
rect 4039 2608 4060 2642
rect 4005 2600 4060 2608
rect 3795 2568 3845 2584
rect 3829 2534 3845 2568
rect 3879 2577 3954 2584
rect 3879 2572 3896 2577
rect 3879 2538 3895 2572
rect 3930 2543 3954 2577
rect 3929 2538 3954 2543
rect 4005 2566 4026 2600
rect 3795 2518 3845 2534
rect 4005 2504 4060 2566
rect 3720 2446 3777 2462
rect 3720 2412 3743 2446
rect 3720 2370 3777 2412
rect 3811 2412 3877 2480
rect 3811 2378 3827 2412
rect 3861 2378 3877 2412
rect 3811 2336 3877 2378
rect 3922 2470 4060 2504
rect 4094 2475 4130 2702
rect 4316 2684 4366 2702
rect 4316 2650 4332 2684
rect 4316 2634 4366 2650
rect 4400 2600 4434 2769
rect 4775 2736 4841 2770
rect 4557 2710 4604 2716
rect 4164 2584 4434 2600
rect 4198 2566 4434 2584
rect 4198 2550 4208 2566
rect 4164 2534 4208 2550
rect 4250 2498 4272 2532
rect 4306 2506 4325 2532
rect 4094 2472 4160 2475
rect 3922 2422 3969 2470
rect 4094 2438 4110 2472
rect 4144 2438 4160 2472
rect 4250 2472 4281 2498
rect 4315 2472 4325 2506
rect 4250 2466 4325 2472
rect 3956 2388 3969 2422
rect 3922 2372 3969 2388
rect 4026 2420 4060 2436
rect 4194 2404 4210 2428
rect 4060 2394 4210 2404
rect 4244 2394 4260 2428
rect 4060 2386 4260 2394
rect 4026 2370 4260 2386
rect 4312 2408 4364 2424
rect 4346 2374 4364 2408
rect 4312 2336 4364 2374
rect 4400 2412 4434 2566
rect 4468 2684 4509 2700
rect 4502 2650 4509 2684
rect 4468 2580 4509 2650
rect 4591 2684 4604 2710
rect 4775 2702 4791 2736
rect 4825 2702 4841 2736
rect 4965 2778 4999 2794
rect 5059 2760 5085 2794
rect 5119 2760 5135 2794
rect 5183 2769 5299 2803
rect 5333 2769 5349 2803
rect 5392 2796 5426 2812
rect 4965 2726 4999 2744
rect 4879 2710 5149 2726
rect 4557 2650 4570 2676
rect 4879 2676 4965 2710
rect 4999 2684 5149 2710
rect 4999 2676 5115 2684
rect 4557 2634 4604 2650
rect 4644 2642 4845 2650
rect 4644 2608 4649 2642
rect 4683 2608 4845 2642
rect 4644 2602 4845 2608
rect 4779 2600 4845 2602
rect 4468 2574 4592 2580
rect 4468 2544 4557 2574
rect 4535 2540 4557 2544
rect 4591 2540 4592 2574
rect 4779 2566 4795 2600
rect 4829 2566 4845 2600
rect 4535 2510 4592 2540
rect 4569 2476 4592 2510
rect 4651 2532 4667 2566
rect 4701 2532 4717 2566
rect 4879 2532 4913 2676
rect 5099 2650 5115 2676
rect 5099 2634 5149 2650
rect 4947 2600 4997 2616
rect 5183 2600 5217 2769
rect 5392 2712 5426 2762
rect 5460 2780 5530 2846
rect 5460 2746 5476 2780
rect 5510 2746 5530 2780
rect 5569 2796 5614 2812
rect 5569 2762 5580 2796
rect 5569 2728 5614 2762
rect 5648 2780 5714 2846
rect 5648 2746 5664 2780
rect 5698 2746 5714 2780
rect 5748 2796 5800 2812
rect 5782 2762 5800 2796
rect 5251 2684 5293 2710
rect 5285 2676 5293 2684
rect 5327 2676 5351 2710
rect 5392 2678 5535 2712
rect 5285 2650 5351 2676
rect 5251 2634 5351 2650
rect 4981 2566 5217 2600
rect 4947 2550 4991 2566
rect 5137 2558 5217 2566
rect 4651 2498 4913 2532
rect 5033 2512 5049 2532
rect 4535 2460 4592 2476
rect 4869 2472 4913 2498
rect 5017 2506 5049 2512
rect 5083 2498 5099 2532
rect 5051 2472 5099 2498
rect 4801 2446 4835 2462
rect 4869 2438 4885 2472
rect 4919 2438 4935 2472
rect 5017 2466 5099 2472
rect 4400 2378 4503 2412
rect 4537 2378 4553 2412
rect 4400 2372 4553 2378
rect 4681 2378 4697 2412
rect 4731 2378 4747 2412
rect 4681 2336 4747 2378
rect 4801 2404 4835 2412
rect 4969 2404 4985 2428
rect 4801 2394 4985 2404
rect 5019 2394 5035 2428
rect 4801 2370 5035 2394
rect 5069 2408 5103 2424
rect 5069 2336 5103 2374
rect 5137 2412 5171 2558
rect 5205 2506 5221 2522
rect 5255 2488 5271 2522
rect 5239 2472 5271 2488
rect 5205 2448 5271 2472
rect 5307 2510 5351 2634
rect 5385 2629 5467 2644
rect 5385 2595 5396 2629
rect 5430 2595 5467 2629
rect 5385 2570 5467 2595
rect 5385 2536 5433 2570
rect 5385 2520 5467 2536
rect 5307 2476 5317 2510
rect 5501 2484 5535 2678
rect 5307 2460 5351 2476
rect 5392 2446 5535 2484
rect 5569 2694 5580 2728
rect 5748 2728 5800 2762
rect 5569 2506 5614 2694
rect 5603 2472 5614 2506
rect 5392 2430 5426 2446
rect 5137 2378 5286 2412
rect 5320 2378 5336 2412
rect 5569 2438 5614 2472
rect 5649 2710 5748 2712
rect 5649 2676 5661 2710
rect 5695 2694 5748 2710
rect 5782 2694 5800 2728
rect 5695 2678 5800 2694
rect 5834 2768 5886 2812
rect 5834 2734 5852 2768
rect 5834 2700 5886 2734
rect 5649 2583 5695 2676
rect 5834 2666 5852 2700
rect 5920 2792 5979 2846
rect 5920 2758 5936 2792
rect 5970 2758 5979 2792
rect 5920 2724 5979 2758
rect 5920 2690 5936 2724
rect 5970 2690 5979 2724
rect 5920 2672 5979 2690
rect 6015 2786 6078 2802
rect 6015 2752 6031 2786
rect 6065 2752 6078 2786
rect 6015 2718 6078 2752
rect 6015 2684 6031 2718
rect 6065 2684 6078 2718
rect 5683 2549 5695 2583
rect 5649 2480 5695 2549
rect 5729 2585 5800 2644
rect 5834 2608 5886 2666
rect 5834 2585 5877 2608
rect 5729 2583 5877 2585
rect 6015 2584 6078 2684
rect 5729 2549 5751 2583
rect 5785 2549 5877 2583
rect 5729 2537 5877 2549
rect 5729 2514 5800 2537
rect 5834 2484 5877 2537
rect 5911 2568 6078 2584
rect 5945 2534 6078 2568
rect 5911 2518 6078 2534
rect 5649 2446 5800 2480
rect 5392 2380 5426 2396
rect 5137 2372 5336 2378
rect 5460 2378 5476 2412
rect 5510 2378 5530 2412
rect 5569 2404 5580 2438
rect 5748 2438 5800 2446
rect 5569 2388 5614 2404
rect 5460 2336 5530 2378
rect 5648 2378 5664 2412
rect 5698 2378 5714 2412
rect 5782 2404 5800 2438
rect 5748 2388 5800 2404
rect 5834 2469 5886 2484
rect 5834 2435 5841 2469
rect 5875 2448 5886 2469
rect 5834 2414 5852 2435
rect 6015 2438 6078 2518
rect 5648 2336 5714 2378
rect 5834 2370 5886 2414
rect 5920 2412 5979 2428
rect 5920 2378 5936 2412
rect 5970 2378 5979 2412
rect 5920 2336 5979 2378
rect 6015 2404 6031 2438
rect 6065 2404 6078 2438
rect 6015 2370 6078 2404
rect 6112 2767 6169 2812
rect 6203 2804 6480 2846
rect 6203 2770 6219 2804
rect 6253 2770 6430 2804
rect 6464 2770 6480 2804
rect 6668 2804 6744 2846
rect 6586 2778 6620 2794
rect 6112 2733 6135 2767
rect 6668 2770 6694 2804
rect 6728 2770 6744 2804
rect 7167 2804 7233 2846
rect 6586 2736 6620 2744
rect 6792 2769 6908 2803
rect 6942 2769 6958 2803
rect 7167 2770 7183 2804
rect 7217 2770 7233 2804
rect 7451 2794 7527 2846
rect 6112 2699 6169 2733
rect 6112 2665 6135 2699
rect 6112 2645 6169 2665
rect 6203 2702 6758 2736
rect 6112 2462 6153 2645
rect 6203 2584 6237 2702
rect 6300 2634 6316 2668
rect 6350 2642 6452 2668
rect 6350 2634 6397 2642
rect 6431 2608 6452 2642
rect 6397 2600 6452 2608
rect 6187 2568 6237 2584
rect 6221 2534 6237 2568
rect 6271 2577 6346 2584
rect 6271 2572 6290 2577
rect 6271 2538 6287 2572
rect 6324 2543 6346 2577
rect 6321 2538 6346 2543
rect 6397 2566 6418 2600
rect 6187 2518 6237 2534
rect 6397 2504 6452 2566
rect 6112 2446 6169 2462
rect 6112 2412 6135 2446
rect 6112 2370 6169 2412
rect 6203 2412 6269 2480
rect 6203 2378 6219 2412
rect 6253 2378 6269 2412
rect 6203 2336 6269 2378
rect 6314 2470 6452 2504
rect 6486 2475 6522 2702
rect 6708 2684 6758 2702
rect 6708 2650 6724 2684
rect 6708 2634 6758 2650
rect 6792 2600 6826 2769
rect 7167 2736 7233 2770
rect 6949 2710 6996 2716
rect 6556 2584 6826 2600
rect 6590 2566 6826 2584
rect 6590 2550 6600 2566
rect 6556 2534 6600 2550
rect 6642 2498 6664 2532
rect 6698 2506 6717 2532
rect 6486 2472 6552 2475
rect 6314 2422 6361 2470
rect 6486 2438 6502 2472
rect 6536 2438 6552 2472
rect 6642 2472 6673 2498
rect 6707 2472 6717 2506
rect 6642 2466 6717 2472
rect 6348 2388 6361 2422
rect 6314 2372 6361 2388
rect 6418 2420 6452 2436
rect 6586 2404 6602 2428
rect 6452 2394 6602 2404
rect 6636 2394 6652 2428
rect 6452 2386 6652 2394
rect 6418 2370 6652 2386
rect 6704 2408 6756 2424
rect 6738 2374 6756 2408
rect 6704 2336 6756 2374
rect 6792 2412 6826 2566
rect 6860 2684 6901 2700
rect 6894 2650 6901 2684
rect 6860 2580 6901 2650
rect 6983 2684 6996 2710
rect 7167 2702 7183 2736
rect 7217 2702 7233 2736
rect 7357 2778 7391 2794
rect 7451 2760 7477 2794
rect 7511 2760 7527 2794
rect 7575 2769 7691 2803
rect 7725 2769 7741 2803
rect 7784 2796 7818 2812
rect 7357 2726 7391 2744
rect 7271 2710 7541 2726
rect 6949 2650 6962 2676
rect 7271 2676 7357 2710
rect 7391 2684 7541 2710
rect 7391 2676 7507 2684
rect 6949 2634 6996 2650
rect 7036 2642 7237 2650
rect 7036 2608 7041 2642
rect 7075 2608 7237 2642
rect 7036 2602 7237 2608
rect 7171 2600 7237 2602
rect 6860 2574 6984 2580
rect 6860 2544 6949 2574
rect 6927 2540 6949 2544
rect 6983 2540 6984 2574
rect 7171 2566 7187 2600
rect 7221 2566 7237 2600
rect 6927 2510 6984 2540
rect 6961 2476 6984 2510
rect 7043 2532 7059 2566
rect 7093 2532 7109 2566
rect 7271 2532 7305 2676
rect 7491 2650 7507 2676
rect 7491 2634 7541 2650
rect 7339 2600 7389 2616
rect 7575 2600 7609 2769
rect 7784 2712 7818 2762
rect 7852 2780 7922 2846
rect 7852 2746 7868 2780
rect 7902 2746 7922 2780
rect 7961 2796 8006 2812
rect 7961 2762 7972 2796
rect 7961 2728 8006 2762
rect 8040 2780 8106 2846
rect 8040 2746 8056 2780
rect 8090 2746 8106 2780
rect 8140 2796 8192 2812
rect 8174 2762 8192 2796
rect 7643 2684 7685 2710
rect 7677 2676 7685 2684
rect 7719 2676 7743 2710
rect 7784 2678 7927 2712
rect 7677 2650 7743 2676
rect 7643 2634 7743 2650
rect 7373 2566 7609 2600
rect 7339 2550 7383 2566
rect 7529 2558 7609 2566
rect 7043 2498 7305 2532
rect 7425 2512 7441 2532
rect 6927 2460 6984 2476
rect 7261 2472 7305 2498
rect 7409 2506 7441 2512
rect 7475 2498 7491 2532
rect 7443 2472 7491 2498
rect 7193 2446 7227 2462
rect 7261 2438 7277 2472
rect 7311 2438 7327 2472
rect 7409 2466 7491 2472
rect 6792 2378 6895 2412
rect 6929 2378 6945 2412
rect 6792 2372 6945 2378
rect 7073 2378 7089 2412
rect 7123 2378 7139 2412
rect 7073 2336 7139 2378
rect 7193 2404 7227 2412
rect 7361 2404 7377 2428
rect 7193 2394 7377 2404
rect 7411 2394 7427 2428
rect 7193 2370 7427 2394
rect 7461 2408 7495 2424
rect 7461 2336 7495 2374
rect 7529 2412 7563 2558
rect 7597 2506 7613 2522
rect 7647 2488 7663 2522
rect 7631 2472 7663 2488
rect 7597 2448 7663 2472
rect 7699 2510 7743 2634
rect 7777 2633 7859 2644
rect 7777 2599 7787 2633
rect 7821 2599 7859 2633
rect 7777 2570 7859 2599
rect 7777 2536 7825 2570
rect 7777 2520 7859 2536
rect 7699 2476 7709 2510
rect 7893 2484 7927 2678
rect 7699 2460 7743 2476
rect 7784 2446 7927 2484
rect 7961 2694 7972 2728
rect 8140 2728 8192 2762
rect 7961 2506 8006 2694
rect 7995 2472 8006 2506
rect 7784 2430 7818 2446
rect 7529 2378 7678 2412
rect 7712 2378 7728 2412
rect 7961 2438 8006 2472
rect 8041 2710 8140 2712
rect 8041 2676 8053 2710
rect 8087 2694 8140 2710
rect 8174 2694 8192 2728
rect 8087 2678 8192 2694
rect 8226 2768 8278 2812
rect 8226 2734 8244 2768
rect 8226 2700 8278 2734
rect 8041 2583 8087 2676
rect 8226 2666 8244 2700
rect 8312 2792 8371 2846
rect 8312 2758 8328 2792
rect 8362 2758 8371 2792
rect 8312 2724 8371 2758
rect 8312 2690 8328 2724
rect 8362 2690 8371 2724
rect 8312 2672 8371 2690
rect 8407 2786 8470 2802
rect 8407 2752 8423 2786
rect 8457 2752 8470 2786
rect 8407 2718 8470 2752
rect 8407 2684 8423 2718
rect 8457 2684 8470 2718
rect 8075 2549 8087 2583
rect 8041 2480 8087 2549
rect 8121 2586 8192 2644
rect 8226 2608 8278 2666
rect 8226 2586 8269 2608
rect 8121 2583 8269 2586
rect 8407 2584 8470 2684
rect 8121 2549 8143 2583
rect 8177 2549 8269 2583
rect 8121 2538 8269 2549
rect 8121 2514 8192 2538
rect 8226 2484 8269 2538
rect 8303 2568 8470 2584
rect 8337 2534 8470 2568
rect 8303 2518 8470 2534
rect 8041 2446 8192 2480
rect 7784 2380 7818 2396
rect 7529 2372 7728 2378
rect 7852 2378 7868 2412
rect 7902 2378 7922 2412
rect 7961 2404 7972 2438
rect 8140 2438 8192 2446
rect 7961 2388 8006 2404
rect 7852 2336 7922 2378
rect 8040 2378 8056 2412
rect 8090 2378 8106 2412
rect 8174 2404 8192 2438
rect 8140 2388 8192 2404
rect 8226 2472 8278 2484
rect 8226 2438 8236 2472
rect 8270 2448 8278 2472
rect 8226 2414 8244 2438
rect 8407 2438 8470 2518
rect 8040 2336 8106 2378
rect 8226 2370 8278 2414
rect 8312 2412 8371 2428
rect 8312 2378 8328 2412
rect 8362 2378 8371 2412
rect 8312 2336 8371 2378
rect 8407 2404 8423 2438
rect 8457 2404 8470 2438
rect 8407 2370 8470 2404
rect 8504 2767 8561 2812
rect 8595 2804 8872 2846
rect 8595 2770 8611 2804
rect 8645 2770 8822 2804
rect 8856 2770 8872 2804
rect 9060 2804 9136 2846
rect 8978 2778 9012 2794
rect 8504 2733 8527 2767
rect 9060 2770 9086 2804
rect 9120 2770 9136 2804
rect 9559 2804 9625 2846
rect 8978 2736 9012 2744
rect 9184 2769 9300 2803
rect 9334 2769 9350 2803
rect 9559 2770 9575 2804
rect 9609 2770 9625 2804
rect 9843 2794 9919 2846
rect 8504 2699 8561 2733
rect 8504 2665 8527 2699
rect 8504 2645 8561 2665
rect 8595 2702 9150 2736
rect 8504 2462 8545 2645
rect 8595 2584 8629 2702
rect 8692 2634 8708 2668
rect 8742 2642 8844 2668
rect 8742 2634 8789 2642
rect 8823 2608 8844 2642
rect 8789 2600 8844 2608
rect 8579 2568 8629 2584
rect 8613 2534 8629 2568
rect 8663 2578 8738 2584
rect 8663 2572 8682 2578
rect 8663 2538 8679 2572
rect 8716 2544 8738 2578
rect 8713 2538 8738 2544
rect 8789 2566 8810 2600
rect 8579 2518 8629 2534
rect 8789 2504 8844 2566
rect 8504 2446 8561 2462
rect 8504 2412 8527 2446
rect 8504 2370 8561 2412
rect 8595 2412 8661 2480
rect 8595 2378 8611 2412
rect 8645 2378 8661 2412
rect 8595 2336 8661 2378
rect 8706 2470 8844 2504
rect 8878 2475 8914 2702
rect 9100 2684 9150 2702
rect 9100 2650 9116 2684
rect 9100 2634 9150 2650
rect 9184 2600 9218 2769
rect 9559 2736 9625 2770
rect 9341 2710 9388 2716
rect 8948 2584 9218 2600
rect 8982 2566 9218 2584
rect 8982 2550 8992 2566
rect 8948 2534 8992 2550
rect 9034 2498 9056 2532
rect 9090 2506 9109 2532
rect 8878 2472 8944 2475
rect 8706 2422 8753 2470
rect 8878 2438 8894 2472
rect 8928 2438 8944 2472
rect 9034 2472 9065 2498
rect 9099 2472 9109 2506
rect 9034 2466 9109 2472
rect 8740 2388 8753 2422
rect 8706 2372 8753 2388
rect 8810 2420 8844 2436
rect 8978 2404 8994 2428
rect 8844 2394 8994 2404
rect 9028 2394 9044 2428
rect 8844 2386 9044 2394
rect 8810 2370 9044 2386
rect 9096 2408 9148 2424
rect 9130 2374 9148 2408
rect 9096 2336 9148 2374
rect 9184 2412 9218 2566
rect 9252 2684 9293 2700
rect 9286 2650 9293 2684
rect 9252 2580 9293 2650
rect 9375 2684 9388 2710
rect 9559 2702 9575 2736
rect 9609 2702 9625 2736
rect 9749 2778 9783 2794
rect 9843 2760 9869 2794
rect 9903 2760 9919 2794
rect 9967 2769 10083 2803
rect 10117 2769 10133 2803
rect 10176 2796 10210 2812
rect 9749 2726 9783 2744
rect 9663 2710 9933 2726
rect 9341 2650 9354 2676
rect 9663 2676 9749 2710
rect 9783 2684 9933 2710
rect 9783 2676 9899 2684
rect 9341 2634 9388 2650
rect 9428 2642 9629 2650
rect 9428 2608 9433 2642
rect 9467 2608 9629 2642
rect 9428 2602 9629 2608
rect 9563 2600 9629 2602
rect 9252 2574 9376 2580
rect 9252 2544 9341 2574
rect 9319 2540 9341 2544
rect 9375 2540 9376 2574
rect 9563 2566 9579 2600
rect 9613 2566 9629 2600
rect 9319 2510 9376 2540
rect 9353 2476 9376 2510
rect 9435 2532 9451 2566
rect 9485 2532 9501 2566
rect 9663 2532 9697 2676
rect 9883 2650 9899 2676
rect 9883 2634 9933 2650
rect 9731 2600 9781 2616
rect 9967 2600 10001 2769
rect 10176 2712 10210 2762
rect 10244 2780 10314 2846
rect 10244 2746 10260 2780
rect 10294 2746 10314 2780
rect 10353 2796 10398 2812
rect 10353 2762 10364 2796
rect 10353 2728 10398 2762
rect 10432 2780 10498 2846
rect 10432 2746 10448 2780
rect 10482 2746 10498 2780
rect 10532 2796 10584 2812
rect 10566 2762 10584 2796
rect 10035 2684 10077 2710
rect 10069 2676 10077 2684
rect 10111 2676 10135 2710
rect 10176 2678 10319 2712
rect 10069 2650 10135 2676
rect 10035 2634 10135 2650
rect 9765 2566 10001 2600
rect 9731 2550 9775 2566
rect 9921 2558 10001 2566
rect 9435 2498 9697 2532
rect 9817 2512 9833 2532
rect 9319 2460 9376 2476
rect 9653 2472 9697 2498
rect 9801 2506 9833 2512
rect 9867 2498 9883 2532
rect 9835 2472 9883 2498
rect 9585 2446 9619 2462
rect 9653 2438 9669 2472
rect 9703 2438 9719 2472
rect 9801 2466 9883 2472
rect 9184 2378 9287 2412
rect 9321 2378 9337 2412
rect 9184 2372 9337 2378
rect 9465 2378 9481 2412
rect 9515 2378 9531 2412
rect 9465 2336 9531 2378
rect 9585 2404 9619 2412
rect 9753 2404 9769 2428
rect 9585 2394 9769 2404
rect 9803 2394 9819 2428
rect 9585 2370 9819 2394
rect 9853 2408 9887 2424
rect 9853 2336 9887 2374
rect 9921 2412 9955 2558
rect 9989 2506 10005 2522
rect 10039 2488 10055 2522
rect 10023 2472 10055 2488
rect 9989 2448 10055 2472
rect 10091 2510 10135 2634
rect 10169 2634 10251 2644
rect 10169 2600 10176 2634
rect 10210 2600 10251 2634
rect 10169 2570 10251 2600
rect 10169 2536 10217 2570
rect 10169 2520 10251 2536
rect 10091 2476 10101 2510
rect 10285 2484 10319 2678
rect 10091 2460 10135 2476
rect 10176 2446 10319 2484
rect 10353 2694 10364 2728
rect 10532 2728 10584 2762
rect 10353 2506 10398 2694
rect 10387 2472 10398 2506
rect 10176 2430 10210 2446
rect 9921 2378 10070 2412
rect 10104 2378 10120 2412
rect 10353 2438 10398 2472
rect 10433 2710 10532 2712
rect 10433 2676 10445 2710
rect 10479 2694 10532 2710
rect 10566 2694 10584 2728
rect 10479 2678 10584 2694
rect 10618 2768 10670 2812
rect 10618 2734 10636 2768
rect 10618 2700 10670 2734
rect 10433 2583 10479 2676
rect 10618 2666 10636 2700
rect 10704 2792 10763 2846
rect 10704 2758 10720 2792
rect 10754 2758 10763 2792
rect 10704 2724 10763 2758
rect 10704 2690 10720 2724
rect 10754 2690 10763 2724
rect 10704 2672 10763 2690
rect 10799 2786 10862 2802
rect 10799 2752 10815 2786
rect 10849 2752 10862 2786
rect 10799 2718 10862 2752
rect 10799 2684 10815 2718
rect 10849 2684 10862 2718
rect 10467 2549 10479 2583
rect 10433 2480 10479 2549
rect 10513 2583 10584 2644
rect 10513 2549 10535 2583
rect 10569 2575 10584 2583
rect 10618 2608 10670 2666
rect 10618 2575 10661 2608
rect 10799 2584 10862 2684
rect 10569 2549 10661 2575
rect 10513 2527 10661 2549
rect 10513 2514 10584 2527
rect 10618 2484 10661 2527
rect 10695 2568 10862 2584
rect 10729 2534 10862 2568
rect 10695 2518 10862 2534
rect 10433 2446 10584 2480
rect 10176 2380 10210 2396
rect 9921 2372 10120 2378
rect 10244 2378 10260 2412
rect 10294 2378 10314 2412
rect 10353 2404 10364 2438
rect 10532 2438 10584 2446
rect 10353 2388 10398 2404
rect 10244 2336 10314 2378
rect 10432 2378 10448 2412
rect 10482 2378 10498 2412
rect 10566 2404 10584 2438
rect 10532 2388 10584 2404
rect 10618 2470 10670 2484
rect 10618 2436 10625 2470
rect 10659 2448 10670 2470
rect 10618 2414 10636 2436
rect 10799 2438 10862 2518
rect 10432 2336 10498 2378
rect 10618 2370 10670 2414
rect 10704 2412 10763 2428
rect 10704 2378 10720 2412
rect 10754 2378 10763 2412
rect 10704 2336 10763 2378
rect 10799 2404 10815 2438
rect 10849 2404 10862 2438
rect 10799 2370 10862 2404
rect 10896 2767 10953 2812
rect 10987 2804 11264 2846
rect 10987 2770 11003 2804
rect 11037 2770 11214 2804
rect 11248 2770 11264 2804
rect 11452 2804 11528 2846
rect 11370 2778 11404 2794
rect 10896 2733 10919 2767
rect 11452 2770 11478 2804
rect 11512 2770 11528 2804
rect 11951 2804 12017 2846
rect 11370 2736 11404 2744
rect 11576 2769 11692 2803
rect 11726 2769 11742 2803
rect 11951 2770 11967 2804
rect 12001 2770 12017 2804
rect 12235 2794 12311 2846
rect 10896 2699 10953 2733
rect 10896 2665 10919 2699
rect 10896 2645 10953 2665
rect 10987 2702 11542 2736
rect 10896 2462 10937 2645
rect 10987 2584 11021 2702
rect 11084 2634 11100 2668
rect 11134 2642 11236 2668
rect 11134 2634 11181 2642
rect 11215 2608 11236 2642
rect 11181 2600 11236 2608
rect 10971 2568 11021 2584
rect 11005 2534 11021 2568
rect 11055 2579 11130 2584
rect 11055 2572 11075 2579
rect 11055 2538 11071 2572
rect 11109 2545 11130 2579
rect 11105 2538 11130 2545
rect 11181 2566 11202 2600
rect 10971 2518 11021 2534
rect 11181 2504 11236 2566
rect 10896 2446 10953 2462
rect 10896 2412 10919 2446
rect 10896 2370 10953 2412
rect 10987 2412 11053 2480
rect 10987 2378 11003 2412
rect 11037 2378 11053 2412
rect 10987 2336 11053 2378
rect 11098 2470 11236 2504
rect 11270 2475 11306 2702
rect 11492 2684 11542 2702
rect 11492 2650 11508 2684
rect 11492 2634 11542 2650
rect 11576 2600 11610 2769
rect 11951 2736 12017 2770
rect 11733 2710 11780 2716
rect 11340 2584 11610 2600
rect 11374 2566 11610 2584
rect 11374 2550 11384 2566
rect 11340 2534 11384 2550
rect 11426 2498 11448 2532
rect 11482 2506 11501 2532
rect 11270 2472 11336 2475
rect 11098 2422 11145 2470
rect 11270 2438 11286 2472
rect 11320 2438 11336 2472
rect 11426 2472 11457 2498
rect 11491 2472 11501 2506
rect 11426 2466 11501 2472
rect 11132 2388 11145 2422
rect 11098 2372 11145 2388
rect 11202 2420 11236 2436
rect 11370 2404 11386 2428
rect 11236 2394 11386 2404
rect 11420 2394 11436 2428
rect 11236 2386 11436 2394
rect 11202 2370 11436 2386
rect 11488 2408 11540 2424
rect 11522 2374 11540 2408
rect 11488 2336 11540 2374
rect 11576 2412 11610 2566
rect 11644 2684 11685 2700
rect 11678 2650 11685 2684
rect 11644 2580 11685 2650
rect 11767 2684 11780 2710
rect 11951 2702 11967 2736
rect 12001 2702 12017 2736
rect 12141 2778 12175 2794
rect 12235 2760 12261 2794
rect 12295 2760 12311 2794
rect 12359 2769 12475 2803
rect 12509 2769 12525 2803
rect 12568 2796 12602 2812
rect 12141 2726 12175 2744
rect 12055 2710 12325 2726
rect 11733 2650 11746 2676
rect 12055 2676 12141 2710
rect 12175 2684 12325 2710
rect 12175 2676 12291 2684
rect 11733 2634 11780 2650
rect 11820 2642 12021 2650
rect 11820 2608 11825 2642
rect 11859 2608 12021 2642
rect 11820 2602 12021 2608
rect 11955 2600 12021 2602
rect 11644 2574 11768 2580
rect 11644 2544 11733 2574
rect 11711 2540 11733 2544
rect 11767 2540 11768 2574
rect 11955 2566 11971 2600
rect 12005 2566 12021 2600
rect 11711 2510 11768 2540
rect 11745 2476 11768 2510
rect 11827 2532 11843 2566
rect 11877 2532 11893 2566
rect 12055 2532 12089 2676
rect 12275 2650 12291 2676
rect 12275 2634 12325 2650
rect 12123 2600 12173 2616
rect 12359 2600 12393 2769
rect 12568 2712 12602 2762
rect 12636 2780 12706 2846
rect 12636 2746 12652 2780
rect 12686 2746 12706 2780
rect 12745 2796 12790 2812
rect 12745 2762 12756 2796
rect 12745 2728 12790 2762
rect 12824 2780 12890 2846
rect 12824 2746 12840 2780
rect 12874 2746 12890 2780
rect 12924 2796 12976 2812
rect 12958 2762 12976 2796
rect 12427 2684 12469 2710
rect 12461 2676 12469 2684
rect 12503 2676 12527 2710
rect 12568 2678 12711 2712
rect 12461 2650 12527 2676
rect 12427 2634 12527 2650
rect 12157 2566 12393 2600
rect 12123 2550 12167 2566
rect 12313 2558 12393 2566
rect 11827 2498 12089 2532
rect 12209 2512 12225 2532
rect 11711 2460 11768 2476
rect 12045 2472 12089 2498
rect 12193 2506 12225 2512
rect 12259 2498 12275 2532
rect 12227 2472 12275 2498
rect 11977 2446 12011 2462
rect 12045 2438 12061 2472
rect 12095 2438 12111 2472
rect 12193 2466 12275 2472
rect 11576 2378 11679 2412
rect 11713 2378 11729 2412
rect 11576 2372 11729 2378
rect 11857 2378 11873 2412
rect 11907 2378 11923 2412
rect 11857 2336 11923 2378
rect 11977 2404 12011 2412
rect 12145 2404 12161 2428
rect 11977 2394 12161 2404
rect 12195 2394 12211 2428
rect 11977 2370 12211 2394
rect 12245 2408 12279 2424
rect 12245 2336 12279 2374
rect 12313 2412 12347 2558
rect 12381 2506 12397 2522
rect 12431 2488 12447 2522
rect 12415 2472 12447 2488
rect 12381 2448 12447 2472
rect 12483 2510 12527 2634
rect 12561 2634 12643 2644
rect 12561 2600 12570 2634
rect 12604 2600 12643 2634
rect 12561 2570 12643 2600
rect 12561 2536 12609 2570
rect 12561 2520 12643 2536
rect 12483 2476 12493 2510
rect 12677 2484 12711 2678
rect 12483 2460 12527 2476
rect 12568 2446 12711 2484
rect 12745 2694 12756 2728
rect 12924 2728 12976 2762
rect 12745 2506 12790 2694
rect 12779 2472 12790 2506
rect 12568 2430 12602 2446
rect 12313 2378 12462 2412
rect 12496 2378 12512 2412
rect 12745 2438 12790 2472
rect 12825 2710 12924 2712
rect 12825 2676 12837 2710
rect 12871 2694 12924 2710
rect 12958 2694 12976 2728
rect 12871 2678 12976 2694
rect 12825 2583 12871 2676
rect 12859 2549 12871 2583
rect 12825 2480 12871 2549
rect 12905 2583 12976 2644
rect 12905 2549 12927 2583
rect 12961 2549 12976 2583
rect 12905 2514 12976 2549
rect 12825 2446 12976 2480
rect 12568 2380 12602 2396
rect 12313 2372 12512 2378
rect 12636 2378 12652 2412
rect 12686 2378 12706 2412
rect 12745 2404 12756 2438
rect 12924 2438 12976 2446
rect 12745 2388 12790 2404
rect 12636 2336 12706 2378
rect 12824 2378 12840 2412
rect 12874 2378 12890 2412
rect 12958 2404 12976 2438
rect 12924 2388 12976 2404
rect 12824 2336 12890 2378
rect 1033 2278 1062 2336
rect 1096 2278 1154 2336
rect 1188 2278 1246 2336
rect 1280 2278 1338 2336
rect 1372 2278 1430 2336
rect 1464 2278 1522 2336
rect 1556 2278 1614 2336
rect 1648 2278 1706 2336
rect 1740 2278 1798 2336
rect 1832 2278 1890 2336
rect 1924 2278 1982 2336
rect 2016 2278 2074 2336
rect 2108 2278 2166 2336
rect 2200 2278 2258 2336
rect 2292 2278 2350 2336
rect 2384 2278 2442 2336
rect 2476 2278 2534 2336
rect 2568 2278 2626 2336
rect 2660 2278 2718 2336
rect 2752 2278 2810 2336
rect 2844 2278 2902 2336
rect 2936 2278 2994 2336
rect 3028 2278 3086 2336
rect 3120 2278 3178 2336
rect 3212 2278 3270 2336
rect 3304 2278 3362 2336
rect 3396 2278 3454 2336
rect 3488 2278 3546 2336
rect 3580 2278 3638 2336
rect 3672 2278 3730 2336
rect 3764 2278 3822 2336
rect 3856 2278 3914 2336
rect 3948 2278 4006 2336
rect 4040 2278 4098 2336
rect 4132 2278 4190 2336
rect 4224 2278 4282 2336
rect 4316 2278 4374 2336
rect 4408 2278 4466 2336
rect 4500 2278 4558 2336
rect 4592 2278 4650 2336
rect 4684 2278 4742 2336
rect 4776 2278 4834 2336
rect 4868 2278 4926 2336
rect 4960 2278 5018 2336
rect 5052 2278 5110 2336
rect 5144 2278 5202 2336
rect 5236 2278 5294 2336
rect 5328 2278 5386 2336
rect 5420 2278 5478 2336
rect 5512 2278 5570 2336
rect 5604 2278 5662 2336
rect 5696 2278 5754 2336
rect 5788 2278 5846 2336
rect 5880 2278 5938 2336
rect 5972 2278 6030 2336
rect 6064 2278 6122 2336
rect 6156 2278 6214 2336
rect 6248 2278 6306 2336
rect 6340 2278 6398 2336
rect 6432 2278 6490 2336
rect 6524 2278 6582 2336
rect 6616 2278 6674 2336
rect 6708 2278 6766 2336
rect 6800 2278 6858 2336
rect 6892 2278 6950 2336
rect 6984 2278 7042 2336
rect 7076 2278 7134 2336
rect 7168 2278 7226 2336
rect 7260 2278 7318 2336
rect 7352 2278 7410 2336
rect 7444 2278 7502 2336
rect 7536 2278 7594 2336
rect 7628 2278 7686 2336
rect 7720 2278 7778 2336
rect 7812 2278 7870 2336
rect 7904 2278 7962 2336
rect 7996 2278 8054 2336
rect 8088 2278 8146 2336
rect 8180 2278 8238 2336
rect 8272 2278 8330 2336
rect 8364 2278 8422 2336
rect 8456 2278 8514 2336
rect 8548 2278 8606 2336
rect 8640 2278 8698 2336
rect 8732 2278 8790 2336
rect 8824 2278 8882 2336
rect 8916 2278 8974 2336
rect 9008 2278 9066 2336
rect 9100 2278 9158 2336
rect 9192 2278 9250 2336
rect 9284 2278 9342 2336
rect 9376 2278 9434 2336
rect 9468 2278 9526 2336
rect 9560 2278 9618 2336
rect 9652 2278 9710 2336
rect 9744 2278 9802 2336
rect 9836 2278 9894 2336
rect 9928 2278 9986 2336
rect 10020 2278 10078 2336
rect 10112 2278 10170 2336
rect 10204 2278 10262 2336
rect 10296 2278 10354 2336
rect 10388 2278 10446 2336
rect 10480 2278 10538 2336
rect 10572 2278 10630 2336
rect 10664 2278 10722 2336
rect 10756 2278 10814 2336
rect 10848 2278 10906 2336
rect 10940 2278 10998 2336
rect 11032 2278 11090 2336
rect 11124 2278 11182 2336
rect 11216 2278 11274 2336
rect 11308 2278 11366 2336
rect 11400 2278 11458 2336
rect 11492 2278 11550 2336
rect 11584 2278 11642 2336
rect 11676 2278 11734 2336
rect 11768 2278 11826 2336
rect 11860 2278 11918 2336
rect 11952 2278 12010 2336
rect 12044 2278 12102 2336
rect 12136 2278 12194 2336
rect 12228 2278 12286 2336
rect 12320 2278 12378 2336
rect 12412 2278 12470 2336
rect 12504 2278 12562 2336
rect 12596 2278 12654 2336
rect 12688 2278 12746 2336
rect 12780 2278 12838 2336
rect 12872 2278 12930 2336
rect 12964 2278 12993 2336
<< viali >>
rect 1064 6178 1098 6188
rect 1064 6154 1098 6178
rect 1156 6178 1190 6188
rect 1156 6154 1190 6178
rect 1248 6178 1282 6188
rect 1248 6154 1282 6178
rect 1340 6178 1374 6188
rect 1340 6154 1374 6178
rect 1432 6178 1466 6188
rect 1432 6154 1466 6178
rect 1524 6178 1558 6188
rect 1524 6154 1558 6178
rect 1616 6178 1650 6188
rect 1616 6154 1650 6178
rect 1708 6154 1742 6188
rect 1800 6154 1834 6188
rect 2324 6178 2358 6188
rect 2324 6154 2358 6178
rect 2416 6178 2450 6188
rect 2416 6154 2450 6178
rect 2508 6178 2542 6188
rect 2508 6154 2542 6178
rect 2600 6178 2634 6188
rect 2600 6154 2634 6178
rect 2692 6178 2726 6188
rect 2692 6154 2726 6178
rect 2784 6178 2818 6188
rect 2784 6154 2818 6178
rect 2876 6178 2910 6188
rect 2876 6154 2910 6178
rect 2968 6178 3002 6188
rect 2968 6154 3002 6178
rect 3060 6178 3094 6188
rect 3060 6154 3094 6178
rect 3152 6178 3186 6188
rect 3152 6154 3186 6178
rect 3244 6178 3278 6188
rect 3244 6154 3278 6178
rect 3336 6178 3370 6188
rect 3336 6154 3370 6178
rect 3428 6178 3462 6188
rect 3428 6154 3462 6178
rect 3520 6178 3554 6188
rect 3520 6154 3554 6178
rect 3612 6178 3646 6188
rect 3612 6154 3646 6178
rect 3704 6178 3738 6188
rect 3704 6154 3738 6178
rect 3796 6178 3830 6188
rect 3796 6154 3830 6178
rect 3888 6178 3922 6188
rect 3888 6154 3922 6178
rect 3980 6178 4014 6188
rect 3980 6154 4014 6178
rect 4072 6178 4106 6188
rect 4072 6154 4106 6178
rect 1068 5876 1102 5883
rect 1068 5849 1072 5876
rect 1072 5849 1102 5876
rect 2783 6052 2817 6086
rect 2967 5992 3001 6018
rect 2967 5984 2977 5992
rect 2977 5984 3001 5992
rect 2875 5916 2909 5950
rect 1712 5849 1746 5883
rect 2410 5846 2444 5880
rect 3243 6052 3277 6086
rect 2778 5709 2812 5743
rect 3138 5856 3145 5884
rect 3145 5856 3172 5884
rect 3138 5850 3172 5856
rect 3427 6052 3461 6086
rect 3703 6052 3737 6086
rect 3795 5984 3829 6018
rect 3519 5796 3540 5813
rect 3540 5796 3553 5813
rect 3519 5779 3553 5796
rect 3613 5796 3636 5813
rect 3636 5796 3647 5813
rect 3613 5779 3647 5796
rect 3887 5934 3921 5950
rect 3887 5916 3890 5934
rect 3890 5916 3921 5934
rect 4071 5916 4105 5950
rect 3891 5718 3925 5752
rect 1064 5620 1098 5644
rect 1064 5610 1098 5620
rect 1156 5620 1190 5644
rect 1156 5610 1190 5620
rect 1248 5620 1282 5644
rect 1248 5610 1282 5620
rect 1340 5620 1374 5644
rect 1340 5610 1374 5620
rect 1432 5620 1466 5644
rect 1432 5610 1466 5620
rect 1524 5620 1558 5644
rect 1524 5610 1558 5620
rect 1616 5620 1650 5644
rect 1616 5610 1650 5620
rect 1708 5620 1742 5644
rect 1708 5610 1742 5620
rect 1800 5620 1834 5644
rect 2324 5620 2358 5644
rect 2416 5620 2450 5644
rect 2508 5620 2542 5644
rect 2600 5620 2634 5644
rect 2692 5620 2726 5644
rect 2784 5620 2818 5644
rect 2876 5620 2910 5644
rect 2968 5620 3002 5644
rect 3060 5620 3094 5644
rect 3152 5620 3186 5644
rect 3244 5620 3278 5644
rect 3336 5620 3370 5644
rect 3428 5620 3462 5644
rect 3520 5620 3554 5644
rect 3612 5620 3646 5644
rect 3704 5620 3738 5644
rect 3796 5620 3830 5644
rect 3888 5620 3922 5644
rect 3980 5620 4014 5644
rect 1800 5610 1834 5620
rect 2324 5610 2352 5620
rect 2352 5610 2358 5620
rect 2416 5610 2444 5620
rect 2444 5610 2450 5620
rect 2508 5610 2536 5620
rect 2536 5610 2542 5620
rect 2600 5610 2628 5620
rect 2628 5610 2634 5620
rect 2692 5610 2720 5620
rect 2720 5610 2726 5620
rect 2784 5610 2812 5620
rect 2812 5610 2818 5620
rect 2876 5610 2904 5620
rect 2904 5610 2910 5620
rect 2968 5610 2996 5620
rect 2996 5610 3002 5620
rect 3060 5610 3088 5620
rect 3088 5610 3094 5620
rect 3152 5610 3180 5620
rect 3180 5610 3186 5620
rect 3244 5610 3272 5620
rect 3272 5610 3278 5620
rect 3336 5610 3364 5620
rect 3364 5610 3370 5620
rect 3428 5610 3456 5620
rect 3456 5610 3462 5620
rect 3520 5610 3548 5620
rect 3548 5610 3554 5620
rect 3612 5610 3640 5620
rect 3640 5610 3646 5620
rect 3704 5610 3732 5620
rect 3732 5610 3738 5620
rect 3796 5610 3824 5620
rect 3824 5610 3830 5620
rect 3888 5610 3916 5620
rect 3916 5610 3922 5620
rect 3980 5610 4008 5620
rect 4008 5610 4014 5620
rect 4072 5610 4106 5644
rect 1063 5305 1097 5315
rect 1063 5281 1097 5305
rect 1155 5305 1189 5315
rect 1155 5281 1189 5305
rect 1247 5305 1281 5315
rect 1247 5281 1281 5305
rect 1339 5305 1373 5315
rect 1339 5281 1373 5305
rect 1431 5305 1465 5315
rect 1431 5281 1465 5305
rect 1523 5305 1557 5315
rect 1523 5281 1557 5305
rect 1615 5305 1649 5315
rect 1615 5281 1649 5305
rect 1707 5305 1741 5315
rect 1707 5281 1741 5305
rect 1799 5305 1833 5315
rect 1799 5281 1833 5305
rect 1891 5305 1925 5315
rect 1891 5281 1925 5305
rect 1983 5305 2017 5315
rect 1983 5281 2017 5305
rect 2075 5305 2109 5315
rect 2075 5281 2109 5305
rect 2167 5305 2201 5315
rect 2167 5281 2201 5305
rect 2259 5305 2293 5315
rect 2259 5281 2293 5305
rect 2351 5305 2385 5315
rect 2351 5281 2385 5305
rect 2443 5305 2477 5315
rect 2443 5281 2477 5305
rect 2535 5305 2569 5315
rect 2535 5281 2569 5305
rect 2627 5305 2661 5315
rect 2627 5281 2661 5305
rect 2719 5305 2753 5315
rect 2719 5281 2753 5305
rect 2811 5305 2845 5315
rect 2811 5281 2845 5305
rect 2903 5296 2934 5315
rect 2934 5296 2937 5315
rect 2903 5281 2937 5296
rect 2995 5281 3029 5315
rect 3087 5305 3121 5315
rect 3087 5281 3121 5305
rect 3179 5305 3213 5315
rect 3179 5281 3213 5305
rect 3271 5305 3305 5315
rect 3271 5281 3305 5305
rect 3363 5305 3397 5315
rect 3363 5281 3397 5305
rect 3455 5305 3489 5315
rect 3455 5281 3489 5305
rect 3547 5305 3581 5315
rect 3547 5281 3581 5305
rect 3639 5305 3640 5315
rect 3640 5305 3673 5315
rect 3731 5305 3765 5315
rect 3639 5281 3673 5305
rect 3731 5281 3765 5305
rect 3823 5305 3857 5315
rect 3823 5281 3857 5305
rect 3915 5305 3949 5315
rect 3915 5281 3949 5305
rect 4007 5305 4041 5315
rect 4007 5281 4041 5305
rect 4099 5281 4133 5315
rect 4191 5299 4211 5315
rect 4211 5299 4225 5315
rect 4191 5281 4225 5299
rect 4283 5305 4317 5315
rect 4283 5281 4317 5305
rect 4375 5305 4409 5315
rect 4375 5281 4409 5305
rect 4467 5305 4501 5315
rect 4467 5281 4501 5305
rect 4559 5305 4593 5315
rect 4559 5281 4593 5305
rect 4651 5305 4685 5315
rect 4651 5281 4685 5305
rect 4743 5305 4777 5315
rect 4743 5281 4777 5305
rect 4835 5305 4869 5315
rect 4835 5281 4869 5305
rect 4927 5305 4961 5315
rect 4927 5281 4961 5305
rect 5019 5305 5053 5315
rect 5019 5281 5053 5305
rect 5111 5305 5145 5315
rect 5111 5281 5145 5305
rect 5203 5305 5237 5315
rect 5203 5281 5237 5305
rect 5295 5305 5329 5315
rect 5295 5281 5329 5305
rect 5387 5305 5421 5315
rect 5387 5281 5421 5305
rect 5479 5305 5513 5315
rect 5479 5281 5513 5305
rect 5571 5305 5605 5315
rect 5571 5281 5605 5305
rect 5663 5305 5697 5315
rect 5663 5281 5697 5305
rect 5755 5305 5789 5315
rect 5755 5281 5789 5305
rect 5847 5305 5881 5315
rect 5847 5281 5881 5305
rect 5939 5305 5973 5315
rect 5939 5281 5973 5305
rect 6031 5305 6065 5315
rect 6031 5281 6065 5305
rect 6123 5305 6157 5315
rect 6123 5281 6157 5305
rect 6215 5305 6249 5315
rect 6215 5281 6249 5305
rect 6307 5305 6341 5315
rect 6307 5281 6341 5305
rect 6399 5305 6433 5315
rect 6399 5281 6433 5305
rect 6491 5281 6525 5315
rect 6583 5301 6603 5315
rect 6603 5301 6617 5315
rect 6583 5281 6617 5301
rect 6675 5305 6709 5315
rect 6675 5281 6709 5305
rect 6767 5305 6801 5315
rect 6767 5281 6801 5305
rect 6859 5305 6893 5315
rect 6859 5281 6893 5305
rect 6951 5305 6985 5315
rect 6951 5281 6985 5305
rect 7043 5305 7077 5315
rect 7043 5281 7077 5305
rect 7135 5305 7169 5315
rect 7135 5281 7169 5305
rect 7227 5305 7261 5315
rect 7227 5281 7261 5305
rect 7319 5305 7353 5315
rect 7319 5281 7353 5305
rect 7411 5305 7445 5315
rect 7411 5281 7445 5305
rect 7503 5305 7537 5315
rect 7503 5281 7537 5305
rect 7595 5305 7629 5315
rect 7595 5281 7629 5305
rect 7687 5305 7721 5315
rect 7687 5281 7721 5305
rect 7779 5305 7813 5315
rect 7779 5281 7813 5305
rect 7871 5305 7905 5315
rect 7871 5281 7905 5305
rect 7963 5305 7997 5315
rect 7963 5281 7997 5305
rect 8055 5305 8089 5315
rect 8055 5281 8089 5305
rect 8147 5305 8181 5315
rect 8147 5281 8181 5305
rect 8239 5305 8273 5315
rect 8239 5281 8273 5305
rect 8331 5305 8365 5315
rect 8331 5281 8365 5305
rect 8423 5305 8457 5315
rect 8423 5281 8457 5305
rect 8515 5305 8549 5315
rect 8515 5281 8549 5305
rect 8607 5305 8641 5315
rect 8607 5281 8641 5305
rect 8699 5305 8733 5315
rect 8699 5281 8733 5305
rect 8791 5305 8825 5315
rect 8791 5281 8825 5305
rect 8883 5281 8917 5315
rect 8975 5301 8995 5315
rect 8995 5301 9009 5315
rect 8975 5281 9009 5301
rect 9067 5305 9101 5315
rect 9067 5281 9101 5305
rect 9159 5305 9193 5315
rect 9159 5281 9193 5305
rect 9251 5305 9285 5315
rect 9251 5281 9285 5305
rect 9343 5305 9377 5315
rect 9343 5281 9377 5305
rect 9435 5305 9469 5315
rect 9435 5281 9469 5305
rect 9527 5305 9561 5315
rect 9527 5281 9561 5305
rect 9619 5305 9653 5315
rect 9619 5281 9653 5305
rect 9711 5305 9745 5315
rect 9711 5281 9745 5305
rect 9803 5305 9837 5315
rect 9803 5281 9837 5305
rect 9895 5305 9929 5315
rect 9895 5281 9929 5305
rect 9987 5305 10021 5315
rect 9987 5281 10021 5305
rect 10079 5305 10113 5315
rect 10079 5281 10113 5305
rect 10171 5305 10205 5315
rect 10171 5281 10205 5305
rect 10263 5305 10297 5315
rect 10263 5281 10297 5305
rect 10355 5305 10389 5315
rect 10355 5281 10389 5305
rect 10447 5305 10481 5315
rect 10447 5281 10481 5305
rect 10539 5305 10573 5315
rect 10539 5281 10573 5305
rect 10631 5305 10665 5315
rect 10631 5281 10665 5305
rect 10723 5305 10757 5315
rect 10723 5281 10757 5305
rect 10815 5305 10849 5315
rect 10815 5281 10849 5305
rect 10907 5305 10941 5315
rect 10907 5281 10941 5305
rect 10999 5305 11033 5315
rect 10999 5281 11033 5305
rect 11091 5305 11125 5315
rect 11091 5281 11125 5305
rect 11183 5305 11217 5315
rect 11183 5281 11217 5305
rect 11275 5281 11309 5315
rect 11367 5302 11387 5315
rect 11387 5302 11401 5315
rect 11367 5281 11401 5302
rect 11459 5305 11493 5315
rect 11459 5281 11493 5305
rect 11551 5305 11585 5315
rect 11551 5281 11585 5305
rect 11643 5305 11677 5315
rect 11643 5281 11677 5305
rect 11735 5305 11769 5315
rect 11735 5281 11769 5305
rect 11827 5305 11861 5315
rect 11827 5281 11861 5305
rect 11919 5305 11953 5315
rect 11919 5281 11953 5305
rect 12011 5305 12045 5315
rect 12011 5281 12045 5305
rect 12103 5305 12137 5315
rect 12103 5281 12137 5305
rect 12195 5305 12229 5315
rect 12195 5281 12229 5305
rect 12287 5305 12321 5315
rect 12287 5281 12321 5305
rect 12379 5305 12413 5315
rect 12379 5281 12413 5305
rect 12471 5305 12505 5315
rect 12471 5281 12505 5305
rect 12563 5305 12597 5315
rect 12563 5281 12597 5305
rect 12655 5305 12689 5315
rect 12655 5281 12689 5305
rect 12747 5305 12781 5315
rect 12747 5281 12781 5305
rect 12839 5305 12873 5315
rect 12839 5281 12873 5305
rect 12931 5305 12965 5315
rect 12931 5281 12965 5305
rect 1156 5111 1190 5145
rect 1067 4984 1100 4994
rect 1100 4984 1101 4994
rect 1067 4960 1101 4984
rect 1248 4907 1282 4941
rect 1524 5111 1558 5145
rect 1428 5040 1462 5074
rect 1612 4923 1630 4941
rect 1630 4923 1646 4941
rect 1612 4907 1646 4923
rect 2260 5119 2294 5145
rect 2260 5111 2281 5119
rect 2281 5111 2294 5119
rect 2168 5043 2202 5077
rect 1800 4933 1802 4941
rect 1802 4933 1834 4941
rect 1800 4907 1834 4933
rect 2260 4975 2294 5009
rect 2536 4933 2545 4941
rect 2545 4933 2570 4941
rect 2536 4907 2570 4933
rect 2812 5043 2846 5077
rect 3087 4881 3121 4883
rect 3087 4849 3108 4881
rect 3108 4849 3121 4881
rect 3368 5047 3402 5081
rect 3548 5111 3582 5145
rect 3457 4984 3458 4994
rect 3458 4984 3491 4994
rect 3457 4960 3491 4984
rect 3640 4907 3674 4941
rect 3916 5111 3950 5145
rect 3779 5043 3813 5077
rect 4004 4923 4022 4941
rect 4022 4923 4038 4941
rect 4004 4907 4038 4923
rect 4652 5119 4686 5145
rect 4652 5111 4673 5119
rect 4673 5111 4686 5119
rect 4560 5043 4594 5077
rect 4192 4933 4194 4941
rect 4194 4933 4226 4941
rect 4192 4907 4226 4933
rect 4652 4975 4686 5009
rect 4928 4933 4937 4941
rect 4937 4933 4962 4941
rect 4928 4907 4962 4933
rect 5204 5043 5238 5077
rect 5305 5007 5339 5011
rect 5305 4977 5314 5007
rect 5314 4977 5339 5007
rect 5476 4881 5510 4894
rect 5476 4860 5500 4881
rect 5500 4860 5510 4881
rect 5757 5046 5791 5080
rect 5940 5111 5974 5145
rect 5850 4984 5884 4995
rect 5850 4961 5884 4984
rect 5748 4883 5782 4906
rect 5748 4872 5749 4883
rect 5749 4872 5782 4883
rect 6032 4907 6066 4941
rect 6308 5111 6342 5145
rect 6168 5042 6202 5076
rect 6396 4923 6414 4941
rect 6414 4923 6430 4941
rect 6396 4907 6430 4923
rect 7044 5119 7078 5145
rect 7044 5111 7065 5119
rect 7065 5111 7078 5119
rect 6952 5043 6986 5077
rect 6584 4933 6586 4941
rect 6586 4933 6618 4941
rect 6584 4907 6618 4933
rect 7044 4975 7078 5009
rect 7320 4933 7329 4941
rect 7329 4933 7354 4941
rect 7320 4907 7354 4933
rect 7596 5043 7630 5077
rect 7695 5007 7729 5012
rect 7695 4978 7706 5007
rect 7706 4978 7729 5007
rect 7864 4881 7898 4897
rect 7864 4863 7892 4881
rect 7892 4863 7898 4881
rect 8332 5111 8366 5145
rect 8152 5044 8186 5078
rect 8242 4984 8276 4994
rect 8242 4960 8276 4984
rect 8144 4883 8178 4895
rect 8144 4861 8175 4883
rect 8175 4861 8178 4883
rect 8424 4907 8458 4941
rect 8700 5111 8734 5145
rect 8563 5040 8597 5074
rect 8788 4923 8806 4941
rect 8806 4923 8822 4941
rect 8788 4907 8822 4923
rect 9436 5119 9470 5145
rect 9436 5111 9457 5119
rect 9457 5111 9470 5119
rect 9344 5043 9378 5077
rect 8976 4933 8978 4941
rect 8978 4933 9010 4941
rect 8976 4907 9010 4933
rect 9436 4975 9470 5009
rect 9712 4933 9721 4941
rect 9721 4933 9746 4941
rect 9712 4907 9746 4933
rect 9988 5043 10022 5077
rect 10086 5007 10120 5014
rect 10086 4980 10098 5007
rect 10098 4980 10120 5007
rect 10261 4847 10284 4880
rect 10284 4847 10295 4880
rect 10261 4846 10295 4847
rect 10724 5111 10758 5145
rect 10543 5043 10577 5077
rect 10637 4984 10668 4996
rect 10668 4984 10671 4996
rect 10637 4962 10671 4984
rect 10544 4883 10578 4911
rect 10544 4877 10567 4883
rect 10567 4877 10578 4883
rect 10816 4907 10850 4941
rect 11092 5111 11126 5145
rect 10954 5039 10988 5073
rect 11180 4923 11198 4941
rect 11198 4923 11214 4941
rect 11180 4907 11214 4923
rect 11828 5119 11862 5145
rect 11828 5111 11849 5119
rect 11849 5111 11862 5119
rect 11736 5043 11770 5077
rect 11368 4933 11370 4941
rect 11370 4933 11402 4941
rect 11368 4907 11402 4933
rect 11828 4975 11862 5009
rect 12104 4933 12113 4941
rect 12113 4933 12138 4941
rect 12104 4907 12138 4933
rect 12380 5043 12414 5077
rect 12477 5007 12511 5012
rect 12477 4978 12490 5007
rect 12490 4978 12511 5007
rect 12652 4847 12676 4881
rect 12676 4847 12686 4881
rect 12931 5169 12959 5201
rect 12959 5169 12965 5201
rect 12931 5167 12965 5169
rect 12939 4883 12973 4911
rect 12939 4877 12959 4883
rect 12959 4877 12973 4883
rect 1063 4747 1097 4771
rect 1063 4737 1097 4747
rect 1155 4747 1189 4771
rect 1155 4737 1189 4747
rect 1247 4747 1281 4771
rect 1247 4737 1281 4747
rect 1339 4747 1373 4771
rect 1339 4737 1373 4747
rect 1431 4747 1465 4771
rect 1431 4737 1465 4747
rect 1523 4747 1557 4771
rect 1523 4737 1557 4747
rect 1615 4747 1649 4771
rect 1615 4737 1649 4747
rect 1707 4747 1741 4771
rect 1707 4737 1741 4747
rect 1799 4747 1833 4771
rect 1799 4737 1833 4747
rect 1891 4747 1925 4771
rect 1891 4737 1925 4747
rect 1983 4747 2017 4771
rect 1983 4737 2017 4747
rect 2075 4747 2109 4771
rect 2075 4737 2109 4747
rect 2167 4747 2201 4771
rect 2167 4737 2201 4747
rect 2259 4747 2293 4771
rect 2259 4737 2293 4747
rect 2351 4747 2385 4771
rect 2351 4737 2385 4747
rect 2443 4747 2477 4771
rect 2443 4737 2477 4747
rect 2535 4747 2569 4771
rect 2535 4737 2569 4747
rect 2627 4747 2661 4771
rect 2627 4737 2661 4747
rect 2719 4747 2753 4771
rect 2719 4737 2753 4747
rect 2811 4747 2845 4771
rect 2811 4737 2845 4747
rect 2903 4747 2937 4771
rect 2903 4737 2937 4747
rect 2995 4747 3029 4771
rect 2995 4737 3029 4747
rect 3087 4747 3121 4771
rect 3087 4737 3121 4747
rect 3179 4747 3213 4771
rect 3179 4737 3213 4747
rect 3271 4747 3305 4771
rect 3271 4737 3305 4747
rect 3363 4747 3397 4771
rect 3363 4737 3397 4747
rect 3455 4747 3489 4771
rect 3455 4737 3489 4747
rect 3547 4747 3581 4771
rect 3547 4737 3581 4747
rect 3639 4747 3673 4771
rect 3639 4737 3673 4747
rect 3731 4747 3765 4771
rect 3731 4737 3765 4747
rect 3823 4747 3857 4771
rect 3823 4737 3857 4747
rect 3915 4747 3949 4771
rect 3915 4737 3949 4747
rect 4007 4747 4041 4771
rect 4007 4737 4041 4747
rect 4099 4747 4133 4771
rect 4099 4737 4133 4747
rect 4191 4747 4225 4771
rect 4191 4737 4225 4747
rect 4283 4747 4317 4771
rect 4283 4737 4317 4747
rect 4375 4747 4409 4771
rect 4375 4737 4409 4747
rect 4467 4747 4501 4771
rect 4467 4737 4501 4747
rect 4559 4747 4593 4771
rect 4559 4737 4593 4747
rect 4651 4747 4685 4771
rect 4651 4737 4685 4747
rect 4743 4747 4777 4771
rect 4743 4737 4777 4747
rect 4835 4747 4869 4771
rect 4835 4737 4869 4747
rect 4927 4747 4961 4771
rect 4927 4737 4961 4747
rect 5019 4747 5053 4771
rect 5019 4737 5053 4747
rect 5111 4747 5145 4771
rect 5111 4737 5145 4747
rect 5203 4747 5237 4771
rect 5203 4737 5237 4747
rect 5295 4747 5329 4771
rect 5295 4737 5329 4747
rect 5387 4747 5421 4771
rect 5387 4737 5421 4747
rect 5479 4747 5513 4771
rect 5479 4737 5513 4747
rect 5571 4747 5605 4771
rect 5571 4737 5605 4747
rect 5663 4747 5697 4771
rect 5663 4737 5697 4747
rect 5755 4747 5789 4771
rect 5755 4737 5789 4747
rect 5847 4747 5881 4771
rect 5847 4737 5881 4747
rect 5939 4747 5973 4771
rect 5939 4737 5973 4747
rect 6031 4747 6065 4771
rect 6031 4737 6065 4747
rect 6123 4747 6157 4771
rect 6123 4737 6157 4747
rect 6215 4747 6249 4771
rect 6215 4737 6249 4747
rect 6307 4747 6341 4771
rect 6307 4737 6341 4747
rect 6399 4747 6433 4771
rect 6399 4737 6433 4747
rect 6491 4747 6525 4771
rect 6491 4737 6525 4747
rect 6583 4747 6617 4771
rect 6583 4737 6617 4747
rect 6675 4747 6709 4771
rect 6675 4737 6709 4747
rect 6767 4747 6801 4771
rect 6767 4737 6801 4747
rect 6859 4747 6893 4771
rect 6859 4737 6893 4747
rect 6951 4747 6985 4771
rect 6951 4737 6985 4747
rect 7043 4747 7077 4771
rect 7043 4737 7077 4747
rect 7135 4747 7169 4771
rect 7135 4737 7169 4747
rect 7227 4747 7261 4771
rect 7227 4737 7261 4747
rect 7319 4747 7353 4771
rect 7319 4737 7353 4747
rect 7411 4747 7445 4771
rect 7411 4737 7445 4747
rect 7503 4747 7537 4771
rect 7503 4737 7537 4747
rect 7595 4747 7629 4771
rect 7595 4737 7629 4747
rect 7687 4747 7721 4771
rect 7687 4737 7721 4747
rect 7779 4747 7813 4771
rect 7779 4737 7813 4747
rect 7871 4747 7905 4771
rect 7871 4737 7905 4747
rect 7963 4747 7997 4771
rect 7963 4737 7997 4747
rect 8055 4747 8089 4771
rect 8055 4737 8089 4747
rect 8147 4747 8181 4771
rect 8147 4737 8181 4747
rect 8239 4747 8273 4771
rect 8239 4737 8273 4747
rect 8331 4747 8365 4771
rect 8331 4737 8365 4747
rect 8423 4747 8457 4771
rect 8423 4737 8457 4747
rect 8515 4747 8549 4771
rect 8515 4737 8549 4747
rect 8607 4747 8641 4771
rect 8607 4737 8641 4747
rect 8699 4747 8733 4771
rect 8699 4737 8733 4747
rect 8791 4747 8825 4771
rect 8791 4737 8825 4747
rect 8883 4747 8917 4771
rect 8883 4737 8917 4747
rect 8975 4747 9009 4771
rect 8975 4737 9009 4747
rect 9067 4747 9101 4771
rect 9067 4737 9101 4747
rect 9159 4747 9193 4771
rect 9159 4737 9193 4747
rect 9251 4747 9285 4771
rect 9251 4737 9285 4747
rect 9343 4747 9377 4771
rect 9343 4737 9377 4747
rect 9435 4747 9469 4771
rect 9435 4737 9469 4747
rect 9527 4747 9561 4771
rect 9527 4737 9561 4747
rect 9619 4747 9653 4771
rect 9619 4737 9653 4747
rect 9711 4747 9745 4771
rect 9711 4737 9745 4747
rect 9803 4747 9837 4771
rect 9803 4737 9837 4747
rect 9895 4747 9929 4771
rect 9895 4737 9929 4747
rect 9987 4747 10021 4771
rect 9987 4737 10021 4747
rect 10079 4747 10113 4771
rect 10079 4737 10113 4747
rect 10171 4747 10205 4771
rect 10171 4737 10205 4747
rect 10263 4747 10297 4771
rect 10263 4737 10297 4747
rect 10355 4747 10389 4771
rect 10355 4737 10389 4747
rect 10447 4747 10481 4771
rect 10447 4737 10481 4747
rect 10539 4747 10573 4771
rect 10539 4737 10573 4747
rect 10631 4747 10665 4771
rect 10631 4737 10665 4747
rect 10723 4747 10757 4771
rect 10723 4737 10757 4747
rect 10815 4747 10849 4771
rect 10815 4737 10849 4747
rect 10907 4747 10941 4771
rect 10907 4737 10941 4747
rect 10999 4747 11033 4771
rect 10999 4737 11033 4747
rect 11091 4747 11125 4771
rect 11091 4737 11125 4747
rect 11183 4747 11217 4771
rect 11183 4737 11217 4747
rect 11275 4747 11309 4771
rect 11275 4737 11309 4747
rect 11367 4747 11401 4771
rect 11367 4737 11401 4747
rect 11459 4747 11493 4771
rect 11459 4737 11493 4747
rect 11551 4747 11585 4771
rect 11551 4737 11585 4747
rect 11643 4747 11677 4771
rect 11643 4737 11677 4747
rect 11735 4747 11769 4771
rect 11735 4737 11769 4747
rect 11827 4747 11861 4771
rect 11827 4737 11861 4747
rect 11919 4747 11953 4771
rect 11919 4737 11953 4747
rect 12011 4747 12045 4771
rect 12011 4737 12045 4747
rect 12103 4747 12137 4771
rect 12103 4737 12137 4747
rect 12195 4747 12229 4771
rect 12195 4737 12229 4747
rect 12287 4747 12321 4771
rect 12287 4737 12321 4747
rect 12379 4747 12413 4771
rect 12379 4737 12413 4747
rect 12471 4747 12505 4771
rect 12471 4737 12505 4747
rect 12563 4747 12597 4771
rect 12563 4737 12597 4747
rect 12655 4747 12689 4771
rect 12655 4737 12689 4747
rect 12747 4747 12781 4771
rect 12747 4737 12781 4747
rect 12839 4747 12873 4771
rect 12839 4737 12873 4747
rect 12931 4747 12965 4771
rect 12931 4737 12965 4747
rect 623 4616 657 4626
rect 623 4592 657 4616
rect 715 4616 749 4626
rect 715 4592 749 4616
rect 807 4616 841 4626
rect 807 4592 841 4616
rect 899 4616 933 4626
rect 899 4592 933 4616
rect 991 4616 1025 4626
rect 991 4592 1025 4616
rect 1083 4616 1117 4626
rect 1083 4592 1117 4616
rect 1175 4616 1209 4626
rect 1175 4592 1209 4616
rect 1267 4616 1301 4626
rect 1267 4592 1301 4616
rect 1359 4616 1393 4626
rect 1359 4592 1393 4616
rect 1431 4616 1451 4626
rect 1451 4616 1465 4626
rect 1523 4616 1543 4626
rect 1543 4616 1557 4626
rect 1615 4616 1635 4626
rect 1635 4616 1649 4626
rect 1707 4616 1727 4626
rect 1727 4616 1741 4626
rect 1799 4616 1819 4626
rect 1819 4616 1833 4626
rect 1891 4616 1911 4626
rect 1911 4616 1925 4626
rect 1983 4616 2003 4626
rect 2003 4616 2017 4626
rect 2075 4616 2095 4626
rect 2095 4616 2109 4626
rect 2167 4616 2187 4626
rect 2187 4616 2201 4626
rect 2259 4616 2279 4626
rect 2279 4616 2293 4626
rect 2351 4616 2385 4626
rect 2443 4616 2477 4626
rect 1431 4592 1465 4616
rect 1523 4592 1557 4616
rect 1615 4592 1649 4616
rect 1707 4592 1741 4616
rect 1799 4592 1833 4616
rect 1891 4592 1925 4616
rect 1983 4592 2017 4616
rect 2075 4592 2109 4616
rect 2167 4592 2201 4616
rect 2259 4592 2293 4616
rect 2351 4592 2385 4616
rect 2443 4592 2477 4616
rect 2535 4616 2569 4626
rect 2535 4592 2569 4616
rect 2627 4616 2661 4626
rect 2627 4592 2661 4616
rect 2719 4616 2753 4626
rect 2719 4592 2753 4616
rect 2811 4616 2845 4626
rect 2811 4592 2845 4616
rect 2903 4616 2937 4626
rect 2903 4592 2937 4616
rect 2995 4616 3029 4626
rect 2995 4592 3029 4616
rect 3087 4616 3121 4626
rect 3087 4592 3121 4616
rect 3179 4616 3213 4626
rect 3179 4592 3213 4616
rect 3271 4616 3305 4626
rect 3271 4592 3305 4616
rect 3363 4616 3397 4626
rect 3363 4592 3397 4616
rect 3455 4616 3489 4626
rect 3455 4592 3489 4616
rect 3547 4616 3581 4626
rect 3547 4592 3581 4616
rect 3639 4616 3673 4626
rect 3639 4592 3673 4616
rect 3731 4616 3765 4626
rect 3731 4592 3765 4616
rect 3823 4616 3857 4626
rect 3823 4592 3857 4616
rect 3915 4616 3949 4626
rect 3915 4592 3949 4616
rect 4007 4616 4041 4626
rect 4007 4592 4041 4616
rect 4099 4616 4133 4626
rect 4099 4592 4133 4616
rect 4191 4592 4225 4626
rect 4283 4592 4317 4626
rect 4375 4616 4409 4626
rect 4375 4592 4409 4616
rect 4467 4616 4501 4626
rect 4467 4592 4501 4616
rect 4559 4616 4593 4626
rect 4559 4592 4593 4616
rect 4651 4616 4685 4626
rect 4651 4592 4685 4616
rect 4743 4616 4777 4626
rect 4743 4592 4777 4616
rect 4835 4616 4869 4626
rect 4835 4592 4869 4616
rect 4927 4616 4961 4626
rect 4927 4592 4961 4616
rect 5019 4616 5053 4626
rect 5019 4592 5053 4616
rect 5111 4616 5145 4626
rect 5111 4592 5145 4616
rect 5203 4616 5237 4626
rect 5203 4592 5237 4616
rect 5295 4616 5329 4626
rect 5295 4592 5329 4616
rect 5387 4616 5421 4626
rect 5387 4592 5421 4616
rect 5479 4616 5513 4626
rect 5479 4592 5513 4616
rect 5571 4616 5605 4626
rect 5571 4592 5605 4616
rect 5663 4616 5697 4626
rect 5663 4592 5697 4616
rect 5755 4616 5789 4626
rect 5755 4592 5789 4616
rect 5847 4616 5881 4626
rect 5847 4592 5881 4616
rect 5939 4616 5973 4626
rect 5939 4592 5973 4616
rect 6031 4616 6065 4626
rect 6031 4592 6065 4616
rect 6123 4616 6157 4626
rect 6123 4592 6157 4616
rect 6215 4616 6249 4626
rect 6215 4592 6249 4616
rect 6307 4616 6341 4626
rect 6307 4592 6341 4616
rect 6399 4616 6433 4626
rect 6399 4592 6433 4616
rect 6491 4616 6525 4626
rect 6491 4592 6525 4616
rect 6583 4592 6617 4626
rect 6675 4592 6709 4626
rect 6767 4616 6801 4626
rect 6767 4592 6801 4616
rect 6859 4616 6893 4626
rect 6859 4592 6893 4616
rect 6951 4616 6985 4626
rect 6951 4592 6985 4616
rect 7043 4616 7077 4626
rect 7043 4592 7077 4616
rect 7135 4616 7169 4626
rect 7135 4592 7169 4616
rect 7227 4616 7261 4626
rect 7227 4592 7261 4616
rect 7319 4616 7353 4626
rect 7319 4592 7353 4616
rect 7411 4616 7445 4626
rect 7411 4592 7445 4616
rect 7503 4616 7537 4626
rect 7503 4592 7537 4616
rect 7595 4616 7629 4626
rect 7595 4592 7629 4616
rect 7687 4616 7721 4626
rect 7687 4592 7721 4616
rect 7779 4616 7813 4626
rect 7779 4592 7813 4616
rect 7871 4616 7905 4626
rect 7871 4592 7905 4616
rect 7963 4616 7997 4626
rect 7963 4592 7997 4616
rect 8055 4616 8089 4626
rect 8055 4592 8089 4616
rect 8147 4616 8181 4626
rect 8147 4592 8181 4616
rect 8239 4616 8273 4626
rect 8239 4592 8273 4616
rect 8331 4616 8365 4626
rect 8331 4592 8365 4616
rect 8423 4616 8457 4626
rect 8423 4592 8457 4616
rect 8515 4616 8549 4626
rect 8515 4592 8549 4616
rect 8607 4616 8641 4626
rect 8607 4592 8641 4616
rect 8699 4616 8733 4626
rect 8699 4592 8733 4616
rect 8791 4616 8825 4626
rect 8791 4592 8825 4616
rect 8883 4616 8917 4626
rect 8883 4592 8917 4616
rect 8975 4592 9009 4626
rect 9067 4592 9101 4626
rect 9159 4616 9193 4626
rect 9159 4592 9193 4616
rect 9251 4616 9285 4626
rect 9251 4592 9285 4616
rect 9343 4616 9377 4626
rect 9343 4592 9377 4616
rect 9435 4616 9469 4626
rect 9435 4592 9469 4616
rect 9527 4616 9561 4626
rect 9527 4592 9561 4616
rect 9619 4616 9653 4626
rect 9619 4592 9653 4616
rect 9711 4616 9745 4626
rect 9711 4592 9745 4616
rect 9803 4616 9837 4626
rect 9803 4592 9837 4616
rect 9895 4616 9929 4626
rect 9895 4592 9929 4616
rect 9987 4616 10021 4626
rect 9987 4592 10021 4616
rect 10079 4616 10113 4626
rect 10079 4592 10113 4616
rect 10171 4616 10205 4626
rect 10171 4592 10205 4616
rect 10263 4616 10297 4626
rect 10263 4592 10297 4616
rect 10355 4616 10389 4626
rect 10355 4592 10389 4616
rect 10447 4616 10481 4626
rect 10447 4592 10481 4616
rect 10539 4616 10573 4626
rect 10539 4592 10573 4616
rect 10631 4616 10665 4626
rect 10631 4592 10665 4616
rect 10723 4616 10757 4626
rect 10723 4592 10757 4616
rect 10815 4616 10849 4626
rect 10815 4592 10849 4616
rect 10907 4616 10941 4626
rect 10907 4592 10941 4616
rect 10999 4616 11033 4626
rect 10999 4592 11033 4616
rect 11091 4616 11125 4626
rect 11091 4592 11125 4616
rect 11183 4616 11217 4626
rect 11183 4592 11217 4616
rect 11275 4616 11309 4626
rect 11275 4592 11309 4616
rect 11367 4592 11401 4626
rect 11459 4592 11493 4626
rect 11551 4616 11585 4626
rect 11551 4592 11585 4616
rect 11643 4616 11677 4626
rect 11643 4592 11677 4616
rect 11735 4616 11769 4626
rect 11735 4592 11769 4616
rect 11827 4616 11861 4626
rect 11827 4592 11861 4616
rect 11919 4616 11953 4626
rect 11919 4592 11953 4616
rect 12011 4616 12045 4626
rect 12011 4592 12045 4616
rect 12103 4616 12137 4626
rect 12103 4592 12137 4616
rect 12195 4616 12229 4626
rect 12195 4592 12229 4616
rect 12287 4616 12321 4626
rect 12287 4592 12321 4616
rect 12379 4616 12413 4626
rect 12379 4592 12413 4616
rect 12471 4616 12505 4626
rect 12471 4592 12505 4616
rect 12563 4616 12597 4626
rect 12563 4592 12597 4616
rect 12655 4616 12689 4626
rect 12655 4592 12689 4616
rect 12747 4616 12781 4626
rect 12747 4592 12781 4616
rect 12839 4616 12873 4626
rect 12839 4592 12873 4616
rect 12931 4616 12965 4626
rect 12931 4592 12965 4616
rect 625 4314 659 4318
rect 625 4284 631 4314
rect 631 4284 659 4314
rect 2538 4476 2572 4488
rect 2538 4454 2563 4476
rect 2563 4454 2572 4476
rect 3366 4153 3400 4187
rect 3452 4514 3486 4524
rect 3452 4490 3461 4514
rect 3461 4490 3486 4514
rect 4006 4354 4040 4388
rect 3898 4318 3932 4322
rect 3898 4288 3930 4318
rect 3930 4288 3932 4318
rect 4282 4244 4307 4252
rect 4307 4244 4316 4252
rect 4282 4218 4316 4244
rect 4558 4430 4592 4456
rect 4558 4422 4571 4430
rect 4571 4422 4592 4430
rect 4650 4354 4684 4388
rect 4558 4286 4592 4320
rect 5294 4422 5328 4456
rect 5018 4244 5050 4252
rect 5050 4244 5052 4252
rect 5018 4218 5052 4244
rect 5206 4234 5222 4252
rect 5222 4234 5240 4252
rect 5206 4218 5240 4234
rect 5430 4352 5464 4386
rect 5570 4218 5604 4252
rect 5662 4422 5696 4456
rect 5750 4295 5752 4301
rect 5752 4295 5784 4301
rect 5750 4267 5784 4295
rect 5841 4356 5875 4390
rect 5845 4194 5879 4222
rect 5845 4188 5853 4194
rect 5853 4188 5879 4194
rect 6398 4354 6432 4388
rect 6292 4318 6326 4324
rect 6292 4290 6322 4318
rect 6322 4290 6326 4318
rect 6131 4158 6136 4183
rect 6136 4158 6165 4183
rect 6131 4149 6165 4158
rect 6674 4244 6699 4252
rect 6699 4244 6708 4252
rect 6674 4218 6708 4244
rect 6950 4430 6984 4456
rect 6950 4422 6963 4430
rect 6963 4422 6984 4430
rect 7042 4354 7076 4388
rect 6950 4286 6984 4320
rect 7686 4422 7720 4456
rect 7410 4244 7442 4252
rect 7442 4244 7444 4252
rect 7410 4218 7444 4244
rect 7598 4234 7614 4252
rect 7614 4234 7632 4252
rect 7598 4218 7632 4234
rect 7822 4352 7856 4386
rect 7962 4218 7996 4252
rect 8054 4422 8088 4456
rect 8147 4295 8178 4302
rect 8178 4295 8181 4302
rect 8147 4268 8181 4295
rect 8233 4356 8267 4390
rect 8245 4194 8279 4209
rect 8245 4175 8279 4194
rect 8790 4354 8824 4388
rect 8682 4318 8716 4325
rect 8682 4291 8714 4318
rect 8714 4291 8716 4318
rect 8519 4158 8528 4182
rect 8528 4158 8553 4182
rect 8519 4148 8553 4158
rect 9066 4244 9091 4252
rect 9091 4244 9100 4252
rect 9066 4218 9100 4244
rect 9342 4430 9376 4456
rect 9342 4422 9355 4430
rect 9355 4422 9376 4430
rect 9434 4354 9468 4388
rect 9342 4286 9376 4320
rect 10078 4422 10112 4456
rect 9802 4244 9834 4252
rect 9834 4244 9836 4252
rect 9802 4218 9836 4244
rect 9990 4234 10006 4252
rect 10006 4234 10024 4252
rect 9990 4218 10024 4234
rect 10214 4353 10248 4387
rect 10354 4218 10388 4252
rect 10446 4422 10480 4456
rect 10538 4295 10570 4302
rect 10570 4295 10572 4302
rect 10538 4268 10572 4295
rect 10625 4357 10659 4391
rect 10633 4194 10667 4217
rect 10633 4183 10637 4194
rect 10637 4183 10667 4194
rect 11182 4354 11216 4388
rect 11076 4318 11110 4322
rect 11076 4288 11106 4318
rect 11106 4288 11110 4318
rect 10913 4158 10920 4188
rect 10920 4158 10947 4188
rect 10913 4154 10947 4158
rect 11458 4244 11483 4252
rect 11483 4244 11492 4252
rect 11458 4218 11492 4244
rect 11734 4430 11768 4456
rect 11734 4422 11747 4430
rect 11747 4422 11768 4430
rect 11826 4354 11860 4388
rect 11734 4286 11768 4320
rect 12470 4422 12504 4456
rect 12194 4244 12226 4252
rect 12226 4244 12228 4252
rect 12194 4218 12228 4244
rect 12382 4234 12398 4252
rect 12398 4234 12416 4252
rect 12382 4218 12416 4234
rect 12575 4349 12609 4383
rect 12746 4218 12780 4252
rect 12838 4422 12872 4456
rect 12930 4341 12964 4375
rect 623 4058 657 4082
rect 623 4048 657 4058
rect 715 4058 749 4082
rect 715 4048 749 4058
rect 807 4058 841 4082
rect 807 4048 841 4058
rect 899 4058 933 4082
rect 899 4048 933 4058
rect 991 4058 1025 4082
rect 991 4048 1025 4058
rect 1083 4058 1117 4082
rect 1083 4048 1117 4058
rect 1175 4058 1209 4082
rect 1175 4048 1209 4058
rect 1267 4058 1301 4082
rect 1267 4048 1301 4058
rect 1359 4058 1393 4082
rect 1359 4048 1393 4058
rect 1431 4058 1465 4082
rect 1523 4058 1557 4082
rect 1615 4058 1649 4082
rect 1707 4058 1741 4082
rect 1799 4058 1833 4082
rect 1891 4058 1925 4082
rect 1983 4058 2017 4082
rect 2075 4058 2109 4082
rect 2167 4058 2201 4082
rect 2259 4058 2293 4082
rect 2351 4058 2385 4082
rect 2443 4058 2477 4082
rect 2535 4058 2569 4082
rect 2627 4058 2661 4082
rect 2719 4058 2753 4082
rect 2811 4058 2845 4082
rect 2903 4058 2937 4082
rect 2995 4058 3029 4082
rect 3087 4058 3121 4082
rect 3179 4058 3213 4082
rect 3271 4058 3305 4082
rect 3363 4058 3397 4082
rect 3455 4058 3489 4082
rect 3547 4058 3581 4082
rect 3639 4058 3673 4082
rect 3731 4058 3765 4082
rect 3823 4058 3857 4082
rect 3915 4058 3949 4082
rect 4007 4058 4041 4082
rect 4099 4058 4133 4082
rect 4191 4058 4225 4082
rect 4283 4058 4317 4082
rect 4375 4058 4409 4082
rect 4467 4058 4501 4082
rect 4559 4058 4593 4082
rect 4651 4058 4685 4082
rect 4743 4058 4777 4082
rect 4835 4058 4869 4082
rect 4927 4058 4961 4082
rect 5019 4058 5053 4082
rect 5111 4058 5145 4082
rect 5203 4058 5237 4082
rect 5295 4058 5329 4082
rect 5387 4058 5421 4082
rect 5479 4058 5513 4082
rect 5571 4058 5605 4082
rect 5663 4058 5697 4082
rect 5755 4058 5789 4082
rect 5847 4058 5881 4082
rect 5939 4058 5973 4082
rect 6031 4058 6065 4082
rect 6123 4058 6157 4082
rect 6215 4058 6249 4082
rect 6307 4058 6341 4082
rect 6399 4058 6433 4082
rect 6491 4058 6525 4082
rect 6583 4058 6617 4082
rect 6675 4058 6709 4082
rect 6767 4058 6801 4082
rect 6859 4058 6893 4082
rect 6951 4058 6985 4082
rect 7043 4058 7077 4082
rect 7135 4058 7169 4082
rect 7227 4058 7261 4082
rect 7319 4058 7353 4082
rect 7411 4058 7445 4082
rect 7503 4058 7537 4082
rect 7595 4058 7629 4082
rect 7687 4058 7721 4082
rect 7779 4058 7813 4082
rect 7871 4058 7905 4082
rect 7963 4058 7997 4082
rect 8055 4058 8089 4082
rect 8147 4058 8181 4082
rect 8239 4058 8273 4082
rect 8331 4058 8365 4082
rect 8423 4058 8457 4082
rect 8515 4058 8549 4082
rect 8607 4058 8641 4082
rect 8699 4058 8733 4082
rect 8791 4058 8825 4082
rect 8883 4058 8917 4082
rect 8975 4058 9009 4082
rect 9067 4058 9101 4082
rect 9159 4058 9193 4082
rect 9251 4058 9285 4082
rect 9343 4058 9377 4082
rect 9435 4058 9469 4082
rect 1431 4048 1451 4058
rect 1451 4048 1465 4058
rect 1523 4048 1543 4058
rect 1543 4048 1557 4058
rect 1615 4048 1635 4058
rect 1635 4048 1649 4058
rect 1707 4048 1727 4058
rect 1727 4048 1741 4058
rect 1799 4048 1819 4058
rect 1819 4048 1833 4058
rect 1891 4048 1911 4058
rect 1911 4048 1925 4058
rect 1983 4048 2003 4058
rect 2003 4048 2017 4058
rect 2075 4048 2095 4058
rect 2095 4048 2109 4058
rect 2167 4048 2187 4058
rect 2187 4048 2201 4058
rect 2259 4048 2279 4058
rect 2279 4048 2293 4058
rect 2351 4048 2371 4058
rect 2371 4048 2385 4058
rect 2443 4048 2463 4058
rect 2463 4048 2477 4058
rect 2535 4048 2555 4058
rect 2555 4048 2569 4058
rect 2627 4048 2647 4058
rect 2647 4048 2661 4058
rect 2719 4048 2739 4058
rect 2739 4048 2753 4058
rect 2811 4048 2831 4058
rect 2831 4048 2845 4058
rect 2903 4048 2923 4058
rect 2923 4048 2937 4058
rect 2995 4048 3015 4058
rect 3015 4048 3029 4058
rect 3087 4048 3107 4058
rect 3107 4048 3121 4058
rect 3179 4048 3199 4058
rect 3199 4048 3213 4058
rect 3271 4048 3291 4058
rect 3291 4048 3305 4058
rect 3363 4048 3383 4058
rect 3383 4048 3397 4058
rect 3455 4048 3475 4058
rect 3475 4048 3489 4058
rect 3547 4048 3567 4058
rect 3567 4048 3581 4058
rect 3639 4048 3659 4058
rect 3659 4048 3673 4058
rect 3731 4048 3751 4058
rect 3751 4048 3765 4058
rect 3823 4048 3843 4058
rect 3843 4048 3857 4058
rect 3915 4048 3935 4058
rect 3935 4048 3949 4058
rect 4007 4048 4027 4058
rect 4027 4048 4041 4058
rect 4099 4048 4119 4058
rect 4119 4048 4133 4058
rect 4191 4048 4211 4058
rect 4211 4048 4225 4058
rect 4283 4048 4303 4058
rect 4303 4048 4317 4058
rect 4375 4048 4395 4058
rect 4395 4048 4409 4058
rect 4467 4048 4487 4058
rect 4487 4048 4501 4058
rect 4559 4048 4579 4058
rect 4579 4048 4593 4058
rect 4651 4048 4671 4058
rect 4671 4048 4685 4058
rect 4743 4048 4763 4058
rect 4763 4048 4777 4058
rect 4835 4048 4855 4058
rect 4855 4048 4869 4058
rect 4927 4048 4947 4058
rect 4947 4048 4961 4058
rect 5019 4048 5039 4058
rect 5039 4048 5053 4058
rect 5111 4048 5131 4058
rect 5131 4048 5145 4058
rect 5203 4048 5223 4058
rect 5223 4048 5237 4058
rect 5295 4048 5315 4058
rect 5315 4048 5329 4058
rect 5387 4048 5407 4058
rect 5407 4048 5421 4058
rect 5479 4048 5499 4058
rect 5499 4048 5513 4058
rect 5571 4048 5591 4058
rect 5591 4048 5605 4058
rect 5663 4048 5683 4058
rect 5683 4048 5697 4058
rect 5755 4048 5775 4058
rect 5775 4048 5789 4058
rect 5847 4048 5867 4058
rect 5867 4048 5881 4058
rect 5939 4048 5959 4058
rect 5959 4048 5973 4058
rect 6031 4048 6051 4058
rect 6051 4048 6065 4058
rect 6123 4048 6143 4058
rect 6143 4048 6157 4058
rect 6215 4048 6235 4058
rect 6235 4048 6249 4058
rect 6307 4048 6327 4058
rect 6327 4048 6341 4058
rect 6399 4048 6419 4058
rect 6419 4048 6433 4058
rect 6491 4048 6511 4058
rect 6511 4048 6525 4058
rect 6583 4048 6603 4058
rect 6603 4048 6617 4058
rect 6675 4048 6695 4058
rect 6695 4048 6709 4058
rect 6767 4048 6787 4058
rect 6787 4048 6801 4058
rect 6859 4048 6879 4058
rect 6879 4048 6893 4058
rect 6951 4048 6971 4058
rect 6971 4048 6985 4058
rect 7043 4048 7063 4058
rect 7063 4048 7077 4058
rect 7135 4048 7155 4058
rect 7155 4048 7169 4058
rect 7227 4048 7247 4058
rect 7247 4048 7261 4058
rect 7319 4048 7339 4058
rect 7339 4048 7353 4058
rect 7411 4048 7431 4058
rect 7431 4048 7445 4058
rect 7503 4048 7523 4058
rect 7523 4048 7537 4058
rect 7595 4048 7615 4058
rect 7615 4048 7629 4058
rect 7687 4048 7707 4058
rect 7707 4048 7721 4058
rect 7779 4048 7799 4058
rect 7799 4048 7813 4058
rect 7871 4048 7891 4058
rect 7891 4048 7905 4058
rect 7963 4048 7983 4058
rect 7983 4048 7997 4058
rect 8055 4048 8075 4058
rect 8075 4048 8089 4058
rect 8147 4048 8167 4058
rect 8167 4048 8181 4058
rect 8239 4048 8259 4058
rect 8259 4048 8273 4058
rect 8331 4048 8351 4058
rect 8351 4048 8365 4058
rect 8423 4048 8443 4058
rect 8443 4048 8457 4058
rect 8515 4048 8535 4058
rect 8535 4048 8549 4058
rect 8607 4048 8627 4058
rect 8627 4048 8641 4058
rect 8699 4048 8719 4058
rect 8719 4048 8733 4058
rect 8791 4048 8811 4058
rect 8811 4048 8825 4058
rect 8883 4048 8903 4058
rect 8903 4048 8917 4058
rect 8975 4048 8995 4058
rect 8995 4048 9009 4058
rect 9067 4048 9087 4058
rect 9087 4048 9101 4058
rect 9159 4048 9179 4058
rect 9179 4048 9193 4058
rect 9251 4048 9271 4058
rect 9271 4048 9285 4058
rect 9343 4048 9363 4058
rect 9363 4048 9377 4058
rect 9435 4048 9469 4058
rect 9527 4058 9561 4082
rect 9527 4048 9561 4058
rect 9619 4058 9653 4082
rect 9619 4048 9653 4058
rect 9711 4058 9745 4082
rect 9711 4048 9745 4058
rect 9803 4058 9837 4082
rect 9803 4048 9837 4058
rect 9895 4058 9929 4082
rect 9895 4048 9929 4058
rect 9987 4058 10021 4082
rect 9987 4048 10021 4058
rect 10079 4058 10113 4082
rect 10079 4048 10113 4058
rect 10171 4058 10205 4082
rect 10171 4048 10205 4058
rect 10263 4058 10297 4082
rect 10263 4048 10297 4058
rect 10355 4058 10389 4082
rect 10355 4048 10389 4058
rect 10447 4058 10481 4082
rect 10447 4048 10481 4058
rect 10539 4058 10573 4082
rect 10539 4048 10573 4058
rect 10631 4058 10665 4082
rect 10631 4048 10665 4058
rect 10723 4058 10757 4082
rect 10723 4048 10757 4058
rect 10815 4058 10849 4082
rect 10815 4048 10849 4058
rect 10907 4058 10941 4082
rect 10907 4048 10941 4058
rect 10999 4058 11033 4082
rect 10999 4048 11033 4058
rect 11091 4058 11125 4082
rect 11091 4048 11125 4058
rect 11183 4058 11217 4082
rect 11183 4048 11217 4058
rect 11275 4058 11309 4082
rect 11275 4048 11309 4058
rect 11367 4058 11401 4082
rect 11367 4048 11401 4058
rect 11459 4058 11493 4082
rect 11459 4048 11493 4058
rect 11551 4058 11585 4082
rect 11551 4048 11585 4058
rect 11643 4058 11677 4082
rect 11643 4048 11677 4058
rect 11735 4058 11769 4082
rect 11735 4048 11769 4058
rect 11827 4058 11861 4082
rect 11827 4048 11861 4058
rect 11919 4058 11953 4082
rect 11919 4048 11953 4058
rect 12011 4058 12045 4082
rect 12011 4048 12045 4058
rect 12103 4058 12137 4082
rect 12103 4048 12137 4058
rect 12195 4058 12229 4082
rect 12195 4048 12229 4058
rect 12287 4058 12321 4082
rect 12287 4048 12321 4058
rect 12379 4058 12413 4082
rect 12379 4048 12413 4058
rect 12471 4058 12505 4082
rect 12471 4048 12505 4058
rect 12563 4058 12597 4082
rect 12563 4048 12597 4058
rect 12655 4058 12689 4082
rect 12655 4048 12689 4058
rect 12747 4058 12781 4082
rect 12747 4048 12781 4058
rect 12839 4058 12873 4082
rect 12839 4048 12873 4058
rect 12931 4058 12965 4082
rect 12931 4048 12965 4058
rect 655 3718 689 3752
rect 747 3718 781 3752
rect 839 3718 873 3752
rect 931 3718 965 3752
rect 1023 3718 1057 3752
rect 1115 3718 1149 3752
rect 1207 3718 1241 3752
rect 1299 3718 1333 3752
rect 1391 3718 1425 3752
rect 3197 3743 3231 3753
rect 3197 3719 3231 3743
rect 3289 3743 3323 3753
rect 3289 3719 3323 3743
rect 3381 3743 3415 3753
rect 3381 3719 3415 3743
rect 3454 3743 3473 3753
rect 3473 3743 3488 3753
rect 3546 3743 3565 3753
rect 3565 3743 3580 3753
rect 3638 3743 3657 3753
rect 3657 3743 3672 3753
rect 3730 3743 3749 3753
rect 3749 3743 3764 3753
rect 3822 3743 3841 3753
rect 3841 3743 3856 3753
rect 3914 3743 3933 3753
rect 3933 3743 3948 3753
rect 4006 3743 4025 3753
rect 4025 3743 4040 3753
rect 4098 3743 4117 3753
rect 4117 3743 4132 3753
rect 4190 3743 4209 3753
rect 4209 3743 4224 3753
rect 4282 3743 4301 3753
rect 4301 3743 4316 3753
rect 4374 3743 4393 3753
rect 4393 3743 4408 3753
rect 4466 3743 4485 3753
rect 4485 3743 4500 3753
rect 4558 3743 4577 3753
rect 4577 3743 4592 3753
rect 4650 3743 4669 3753
rect 4669 3743 4684 3753
rect 4742 3743 4761 3753
rect 4761 3743 4776 3753
rect 4834 3743 4853 3753
rect 4853 3743 4868 3753
rect 4926 3743 4945 3753
rect 4945 3743 4960 3753
rect 5018 3743 5052 3753
rect 3454 3719 3488 3743
rect 3546 3719 3580 3743
rect 3638 3719 3672 3743
rect 3730 3719 3764 3743
rect 3822 3719 3856 3743
rect 3914 3719 3948 3743
rect 4006 3719 4040 3743
rect 4098 3719 4132 3743
rect 4190 3719 4224 3743
rect 4282 3719 4316 3743
rect 4374 3719 4408 3743
rect 4466 3719 4500 3743
rect 4558 3719 4592 3743
rect 4650 3719 4684 3743
rect 4742 3719 4776 3743
rect 4834 3719 4868 3743
rect 4926 3719 4960 3743
rect 5018 3719 5052 3743
rect 5110 3743 5144 3753
rect 5110 3719 5144 3743
rect 5202 3743 5236 3753
rect 5202 3719 5236 3743
rect 5294 3743 5328 3753
rect 5294 3719 5328 3743
rect 5386 3743 5420 3753
rect 5386 3719 5420 3743
rect 5478 3743 5512 3753
rect 5478 3719 5512 3743
rect 5570 3743 5604 3753
rect 5570 3719 5604 3743
rect 5662 3743 5696 3753
rect 5662 3719 5696 3743
rect 5754 3743 5788 3753
rect 5754 3719 5788 3743
rect 5846 3743 5880 3753
rect 5846 3719 5880 3743
rect 5938 3743 5972 3753
rect 5938 3719 5972 3743
rect 6030 3743 6064 3753
rect 6030 3719 6064 3743
rect 6122 3743 6156 3753
rect 6122 3719 6156 3743
rect 6214 3743 6248 3753
rect 6214 3719 6248 3743
rect 6306 3743 6340 3753
rect 6306 3719 6340 3743
rect 6398 3743 6432 3753
rect 6398 3719 6432 3743
rect 6490 3743 6524 3753
rect 6490 3719 6524 3743
rect 6582 3743 6616 3753
rect 6582 3719 6616 3743
rect 6674 3743 6708 3753
rect 6674 3719 6708 3743
rect 6766 3743 6800 3753
rect 6766 3719 6800 3743
rect 6858 3743 6892 3753
rect 6858 3719 6892 3743
rect 6950 3743 6984 3753
rect 6950 3719 6984 3743
rect 7042 3743 7076 3753
rect 7042 3719 7076 3743
rect 7134 3743 7168 3753
rect 7134 3719 7168 3743
rect 7226 3743 7260 3753
rect 7226 3719 7260 3743
rect 7318 3743 7352 3753
rect 7318 3719 7352 3743
rect 7410 3743 7444 3753
rect 7410 3719 7444 3743
rect 7502 3743 7536 3753
rect 7502 3719 7536 3743
rect 7594 3743 7628 3753
rect 7594 3719 7628 3743
rect 7686 3743 7720 3753
rect 7686 3719 7720 3743
rect 7778 3743 7812 3753
rect 7778 3719 7812 3743
rect 7870 3743 7904 3753
rect 7870 3719 7904 3743
rect 7962 3743 7996 3753
rect 7962 3719 7996 3743
rect 8054 3743 8088 3753
rect 8054 3719 8088 3743
rect 8146 3743 8180 3753
rect 8146 3719 8180 3743
rect 8238 3743 8272 3753
rect 8238 3719 8272 3743
rect 8330 3743 8364 3753
rect 8330 3719 8364 3743
rect 8422 3743 8456 3753
rect 8422 3719 8456 3743
rect 8514 3743 8548 3753
rect 8514 3719 8548 3743
rect 8606 3743 8640 3753
rect 8606 3719 8640 3743
rect 8698 3743 8732 3753
rect 8698 3719 8732 3743
rect 8790 3743 8824 3753
rect 8790 3719 8824 3743
rect 8882 3743 8916 3753
rect 8882 3719 8916 3743
rect 8974 3743 9008 3753
rect 8974 3719 9008 3743
rect 9066 3743 9100 3753
rect 9066 3719 9100 3743
rect 9158 3743 9192 3753
rect 9158 3719 9192 3743
rect 9250 3743 9284 3753
rect 9250 3719 9284 3743
rect 9342 3743 9376 3753
rect 9342 3719 9376 3743
rect 9434 3743 9468 3753
rect 9434 3719 9468 3743
rect 9526 3743 9560 3753
rect 9526 3719 9560 3743
rect 9618 3743 9652 3753
rect 9618 3719 9652 3743
rect 9710 3743 9744 3753
rect 9710 3719 9744 3743
rect 9802 3743 9836 3753
rect 9802 3719 9836 3743
rect 9894 3743 9928 3753
rect 9894 3719 9928 3743
rect 9986 3743 10020 3753
rect 9986 3719 10020 3743
rect 10078 3743 10112 3753
rect 10078 3719 10112 3743
rect 10170 3743 10204 3753
rect 10170 3719 10204 3743
rect 10262 3743 10296 3753
rect 10262 3719 10296 3743
rect 10354 3743 10388 3753
rect 10354 3719 10388 3743
rect 10446 3743 10480 3753
rect 10446 3719 10480 3743
rect 10538 3743 10572 3753
rect 10538 3719 10572 3743
rect 10630 3743 10664 3753
rect 10630 3719 10664 3743
rect 10722 3743 10756 3753
rect 10722 3719 10756 3743
rect 10814 3743 10848 3753
rect 10814 3719 10848 3743
rect 10906 3743 10940 3753
rect 10906 3719 10940 3743
rect 10998 3743 11032 3753
rect 10998 3719 11032 3743
rect 11090 3743 11124 3753
rect 11090 3719 11124 3743
rect 11182 3743 11216 3753
rect 11182 3719 11216 3743
rect 11274 3743 11308 3753
rect 11274 3719 11308 3743
rect 11366 3743 11400 3753
rect 11366 3719 11400 3743
rect 11458 3743 11492 3753
rect 11458 3719 11492 3743
rect 11550 3743 11584 3753
rect 11550 3719 11584 3743
rect 11642 3743 11676 3753
rect 11642 3719 11676 3743
rect 11734 3743 11768 3753
rect 11734 3719 11768 3743
rect 11826 3743 11860 3753
rect 11826 3719 11860 3743
rect 11918 3743 11952 3753
rect 11918 3719 11952 3743
rect 12010 3743 12044 3753
rect 12010 3719 12044 3743
rect 12102 3743 12136 3753
rect 12102 3719 12136 3743
rect 12194 3743 12228 3753
rect 12194 3719 12228 3743
rect 12286 3743 12320 3753
rect 12286 3719 12320 3743
rect 12378 3743 12412 3753
rect 12378 3719 12412 3743
rect 12470 3743 12504 3753
rect 12470 3719 12504 3743
rect 12562 3743 12596 3753
rect 12562 3719 12596 3743
rect 12654 3743 12688 3753
rect 12654 3719 12688 3743
rect 12746 3743 12780 3753
rect 12746 3719 12780 3743
rect 12838 3743 12872 3753
rect 12838 3719 12872 3743
rect 12930 3743 12964 3753
rect 12930 3719 12964 3743
rect 665 3406 697 3439
rect 697 3406 699 3439
rect 665 3405 699 3406
rect 3547 3549 3581 3583
rect 3347 3507 3362 3520
rect 3362 3507 3381 3520
rect 3347 3486 3381 3507
rect 1270 3406 1304 3440
rect 3162 3412 3196 3446
rect 3455 3422 3457 3445
rect 3457 3422 3489 3445
rect 3455 3411 3489 3422
rect 3639 3345 3673 3379
rect 3915 3549 3949 3583
rect 3784 3443 3818 3453
rect 3784 3419 3809 3443
rect 3809 3419 3818 3443
rect 4003 3361 4021 3379
rect 4021 3361 4037 3379
rect 4003 3345 4037 3361
rect 4651 3557 4685 3583
rect 4651 3549 4672 3557
rect 4672 3549 4685 3557
rect 4559 3481 4593 3515
rect 4191 3371 4193 3379
rect 4193 3371 4225 3379
rect 4191 3345 4225 3371
rect 4651 3413 4685 3447
rect 4927 3371 4936 3379
rect 4936 3371 4961 3379
rect 4927 3345 4961 3371
rect 5203 3481 5237 3515
rect 5303 3445 5337 3446
rect 5303 3412 5313 3445
rect 5313 3412 5337 3445
rect 5939 3549 5973 3583
rect 6031 3345 6065 3379
rect 6307 3549 6341 3583
rect 6200 3443 6234 3449
rect 6200 3415 6201 3443
rect 6201 3415 6234 3443
rect 6395 3361 6413 3379
rect 6413 3361 6429 3379
rect 6395 3345 6429 3361
rect 7043 3557 7077 3583
rect 7043 3549 7064 3557
rect 7064 3549 7077 3557
rect 6951 3481 6985 3515
rect 6583 3371 6585 3379
rect 6585 3371 6617 3379
rect 6583 3345 6617 3371
rect 7043 3413 7077 3447
rect 7319 3371 7328 3379
rect 7328 3371 7353 3379
rect 7319 3345 7353 3371
rect 7595 3481 7629 3515
rect 7693 3445 7727 3454
rect 7693 3420 7705 3445
rect 7705 3420 7727 3445
rect 8331 3549 8365 3583
rect 8149 3321 8183 3347
rect 8149 3313 8174 3321
rect 8174 3313 8183 3321
rect 8423 3345 8457 3379
rect 8699 3549 8733 3583
rect 8587 3443 8621 3449
rect 8587 3415 8593 3443
rect 8593 3415 8621 3443
rect 8787 3361 8805 3379
rect 8805 3361 8821 3379
rect 8787 3345 8821 3361
rect 9435 3557 9469 3583
rect 9435 3549 9456 3557
rect 9456 3549 9469 3557
rect 9343 3481 9377 3515
rect 8975 3371 8977 3379
rect 8977 3371 9009 3379
rect 8975 3345 9009 3371
rect 9435 3413 9469 3447
rect 9711 3371 9720 3379
rect 9720 3371 9745 3379
rect 9711 3345 9745 3371
rect 9987 3481 10021 3515
rect 10084 3445 10118 3450
rect 10084 3416 10097 3445
rect 10097 3416 10118 3445
rect 10723 3549 10757 3583
rect 10541 3321 10575 3348
rect 10541 3314 10566 3321
rect 10566 3314 10575 3321
rect 10815 3345 10849 3379
rect 11091 3549 11125 3583
rect 10990 3414 11024 3448
rect 11179 3361 11197 3379
rect 11197 3361 11213 3379
rect 11179 3345 11213 3361
rect 11827 3557 11861 3583
rect 11827 3549 11848 3557
rect 11848 3549 11861 3557
rect 11735 3481 11769 3515
rect 11367 3371 11369 3379
rect 11369 3371 11401 3379
rect 11367 3345 11401 3371
rect 11827 3413 11861 3447
rect 12103 3371 12112 3379
rect 12112 3371 12137 3379
rect 12103 3345 12137 3371
rect 12379 3481 12413 3515
rect 12476 3445 12510 3449
rect 12476 3415 12489 3445
rect 12489 3415 12510 3445
rect 12931 3321 12965 3351
rect 12931 3317 12958 3321
rect 12958 3317 12965 3321
rect 655 3174 689 3208
rect 747 3174 781 3208
rect 839 3174 873 3208
rect 931 3174 965 3208
rect 1023 3174 1057 3208
rect 1115 3174 1149 3208
rect 1207 3174 1241 3208
rect 1299 3174 1333 3208
rect 1391 3174 1425 3208
rect 3197 3185 3231 3209
rect 3197 3175 3231 3185
rect 3289 3185 3323 3209
rect 3289 3175 3323 3185
rect 3381 3185 3415 3209
rect 3381 3175 3415 3185
rect 3454 3185 3488 3209
rect 3546 3185 3580 3209
rect 3638 3185 3672 3209
rect 3730 3185 3764 3209
rect 3822 3185 3856 3209
rect 3914 3185 3948 3209
rect 4006 3185 4040 3209
rect 4098 3185 4132 3209
rect 4190 3185 4224 3209
rect 4282 3185 4316 3209
rect 4374 3185 4408 3209
rect 4466 3185 4500 3209
rect 4558 3185 4592 3209
rect 4650 3185 4684 3209
rect 4742 3185 4776 3209
rect 4834 3185 4868 3209
rect 4926 3185 4960 3209
rect 5018 3185 5052 3209
rect 5110 3185 5144 3209
rect 5202 3185 5236 3209
rect 5294 3185 5328 3209
rect 5386 3185 5420 3209
rect 5478 3185 5512 3209
rect 5570 3185 5604 3209
rect 5662 3185 5696 3209
rect 5754 3185 5788 3209
rect 5846 3185 5880 3209
rect 5938 3185 5972 3209
rect 6030 3185 6064 3209
rect 6122 3185 6156 3209
rect 6214 3185 6248 3209
rect 6306 3185 6340 3209
rect 6398 3185 6432 3209
rect 6490 3185 6524 3209
rect 6582 3185 6616 3209
rect 6674 3185 6708 3209
rect 6766 3185 6800 3209
rect 6858 3185 6892 3209
rect 6950 3185 6984 3209
rect 7042 3185 7076 3209
rect 7134 3185 7168 3209
rect 7226 3185 7260 3209
rect 7318 3185 7352 3209
rect 7410 3185 7444 3209
rect 7502 3185 7536 3209
rect 7594 3185 7628 3209
rect 7686 3185 7720 3209
rect 7778 3185 7812 3209
rect 7870 3185 7904 3209
rect 7962 3185 7996 3209
rect 8054 3185 8088 3209
rect 8146 3185 8180 3209
rect 8238 3185 8272 3209
rect 8330 3185 8364 3209
rect 8422 3185 8456 3209
rect 8514 3185 8548 3209
rect 8606 3185 8640 3209
rect 8698 3185 8732 3209
rect 8790 3185 8824 3209
rect 8882 3185 8916 3209
rect 8974 3185 9008 3209
rect 9066 3185 9100 3209
rect 9158 3185 9192 3209
rect 9250 3185 9284 3209
rect 9342 3185 9376 3209
rect 9434 3185 9468 3209
rect 9526 3185 9560 3209
rect 9618 3185 9652 3209
rect 9710 3185 9744 3209
rect 9802 3185 9836 3209
rect 9894 3185 9928 3209
rect 9986 3185 10020 3209
rect 10078 3185 10112 3209
rect 10170 3185 10204 3209
rect 10262 3185 10296 3209
rect 10354 3185 10388 3209
rect 10446 3185 10480 3209
rect 10538 3185 10572 3209
rect 10630 3185 10664 3209
rect 10722 3185 10756 3209
rect 10814 3185 10848 3209
rect 10906 3185 10940 3209
rect 10998 3185 11032 3209
rect 11090 3185 11124 3209
rect 11182 3185 11216 3209
rect 11274 3185 11308 3209
rect 11366 3185 11400 3209
rect 11458 3185 11492 3209
rect 11550 3185 11584 3209
rect 11642 3185 11676 3209
rect 11734 3185 11768 3209
rect 11826 3185 11860 3209
rect 11918 3185 11952 3209
rect 12010 3185 12044 3209
rect 3454 3175 3473 3185
rect 3473 3175 3488 3185
rect 3546 3175 3565 3185
rect 3565 3175 3580 3185
rect 3638 3175 3657 3185
rect 3657 3175 3672 3185
rect 3730 3175 3749 3185
rect 3749 3175 3764 3185
rect 3822 3175 3841 3185
rect 3841 3175 3856 3185
rect 3914 3175 3933 3185
rect 3933 3175 3948 3185
rect 4006 3175 4025 3185
rect 4025 3175 4040 3185
rect 4098 3175 4117 3185
rect 4117 3175 4132 3185
rect 4190 3175 4209 3185
rect 4209 3175 4224 3185
rect 4282 3175 4301 3185
rect 4301 3175 4316 3185
rect 4374 3175 4393 3185
rect 4393 3175 4408 3185
rect 4466 3175 4485 3185
rect 4485 3175 4500 3185
rect 4558 3175 4577 3185
rect 4577 3175 4592 3185
rect 4650 3175 4669 3185
rect 4669 3175 4684 3185
rect 4742 3175 4761 3185
rect 4761 3175 4776 3185
rect 4834 3175 4853 3185
rect 4853 3175 4868 3185
rect 4926 3175 4945 3185
rect 4945 3175 4960 3185
rect 5018 3175 5037 3185
rect 5037 3175 5052 3185
rect 5110 3175 5129 3185
rect 5129 3175 5144 3185
rect 5202 3175 5221 3185
rect 5221 3175 5236 3185
rect 5294 3175 5313 3185
rect 5313 3175 5328 3185
rect 5386 3175 5405 3185
rect 5405 3175 5420 3185
rect 5478 3175 5497 3185
rect 5497 3175 5512 3185
rect 5570 3175 5589 3185
rect 5589 3175 5604 3185
rect 5662 3175 5681 3185
rect 5681 3175 5696 3185
rect 5754 3175 5773 3185
rect 5773 3175 5788 3185
rect 5846 3175 5865 3185
rect 5865 3175 5880 3185
rect 5938 3175 5957 3185
rect 5957 3175 5972 3185
rect 6030 3175 6049 3185
rect 6049 3175 6064 3185
rect 6122 3175 6141 3185
rect 6141 3175 6156 3185
rect 6214 3175 6233 3185
rect 6233 3175 6248 3185
rect 6306 3175 6325 3185
rect 6325 3175 6340 3185
rect 6398 3175 6417 3185
rect 6417 3175 6432 3185
rect 6490 3175 6509 3185
rect 6509 3175 6524 3185
rect 6582 3175 6601 3185
rect 6601 3175 6616 3185
rect 6674 3175 6693 3185
rect 6693 3175 6708 3185
rect 6766 3175 6785 3185
rect 6785 3175 6800 3185
rect 6858 3175 6877 3185
rect 6877 3175 6892 3185
rect 6950 3175 6969 3185
rect 6969 3175 6984 3185
rect 7042 3175 7061 3185
rect 7061 3175 7076 3185
rect 7134 3175 7153 3185
rect 7153 3175 7168 3185
rect 7226 3175 7245 3185
rect 7245 3175 7260 3185
rect 7318 3175 7337 3185
rect 7337 3175 7352 3185
rect 7410 3175 7429 3185
rect 7429 3175 7444 3185
rect 7502 3175 7521 3185
rect 7521 3175 7536 3185
rect 7594 3175 7613 3185
rect 7613 3175 7628 3185
rect 7686 3175 7705 3185
rect 7705 3175 7720 3185
rect 7778 3175 7797 3185
rect 7797 3175 7812 3185
rect 7870 3175 7889 3185
rect 7889 3175 7904 3185
rect 7962 3175 7981 3185
rect 7981 3175 7996 3185
rect 8054 3175 8073 3185
rect 8073 3175 8088 3185
rect 8146 3175 8165 3185
rect 8165 3175 8180 3185
rect 8238 3175 8257 3185
rect 8257 3175 8272 3185
rect 8330 3175 8349 3185
rect 8349 3175 8364 3185
rect 8422 3175 8441 3185
rect 8441 3175 8456 3185
rect 8514 3175 8533 3185
rect 8533 3175 8548 3185
rect 8606 3175 8625 3185
rect 8625 3175 8640 3185
rect 8698 3175 8717 3185
rect 8717 3175 8732 3185
rect 8790 3175 8809 3185
rect 8809 3175 8824 3185
rect 8882 3175 8901 3185
rect 8901 3175 8916 3185
rect 8974 3175 8993 3185
rect 8993 3175 9008 3185
rect 9066 3175 9085 3185
rect 9085 3175 9100 3185
rect 9158 3175 9177 3185
rect 9177 3175 9192 3185
rect 9250 3175 9269 3185
rect 9269 3175 9284 3185
rect 9342 3175 9361 3185
rect 9361 3175 9376 3185
rect 9434 3175 9453 3185
rect 9453 3175 9468 3185
rect 9526 3175 9545 3185
rect 9545 3175 9560 3185
rect 9618 3175 9637 3185
rect 9637 3175 9652 3185
rect 9710 3175 9729 3185
rect 9729 3175 9744 3185
rect 9802 3175 9821 3185
rect 9821 3175 9836 3185
rect 9894 3175 9928 3185
rect 9986 3175 10020 3185
rect 10078 3175 10112 3185
rect 10170 3175 10204 3185
rect 10262 3175 10296 3185
rect 10354 3175 10388 3185
rect 10446 3175 10480 3185
rect 10538 3175 10572 3185
rect 10630 3175 10664 3185
rect 10722 3175 10756 3185
rect 10814 3175 10848 3185
rect 10906 3175 10940 3185
rect 10998 3175 11032 3185
rect 11090 3175 11124 3185
rect 11182 3175 11216 3185
rect 11274 3175 11308 3185
rect 11366 3175 11400 3185
rect 11458 3175 11492 3185
rect 11550 3175 11584 3185
rect 11642 3175 11676 3185
rect 11734 3175 11768 3185
rect 11826 3175 11860 3185
rect 11918 3175 11952 3185
rect 12010 3175 12044 3185
rect 12102 3185 12136 3209
rect 12102 3175 12136 3185
rect 12194 3185 12228 3209
rect 12194 3175 12228 3185
rect 12286 3185 12320 3209
rect 12286 3175 12320 3185
rect 12378 3185 12412 3209
rect 12378 3175 12412 3185
rect 12470 3185 12504 3209
rect 12470 3175 12504 3185
rect 12562 3185 12596 3209
rect 12562 3175 12596 3185
rect 12654 3185 12688 3209
rect 12654 3175 12688 3185
rect 12746 3185 12780 3209
rect 12746 3175 12780 3185
rect 12838 3185 12872 3209
rect 12838 3175 12872 3185
rect 12930 3185 12964 3209
rect 12930 3175 12964 3185
rect 1062 2870 1096 2880
rect 1062 2846 1096 2870
rect 1154 2870 1188 2880
rect 1154 2846 1188 2870
rect 1246 2870 1280 2880
rect 1246 2846 1280 2870
rect 1338 2870 1372 2880
rect 1338 2846 1372 2870
rect 1430 2870 1464 2880
rect 1430 2846 1464 2870
rect 1522 2870 1556 2880
rect 1522 2846 1556 2870
rect 1614 2870 1648 2880
rect 1614 2846 1648 2870
rect 1706 2870 1740 2880
rect 1706 2846 1740 2870
rect 1798 2870 1832 2880
rect 1798 2846 1832 2870
rect 1890 2870 1924 2880
rect 1890 2846 1924 2870
rect 1982 2870 2016 2880
rect 1982 2846 2016 2870
rect 2074 2870 2108 2880
rect 2074 2846 2108 2870
rect 2166 2870 2200 2880
rect 2166 2846 2200 2870
rect 2258 2870 2292 2880
rect 2258 2846 2292 2870
rect 2350 2870 2384 2880
rect 2350 2846 2384 2870
rect 2442 2870 2476 2880
rect 2442 2846 2476 2870
rect 2534 2870 2568 2880
rect 2534 2846 2568 2870
rect 2626 2870 2660 2880
rect 2626 2846 2660 2870
rect 2718 2870 2752 2880
rect 2718 2846 2752 2870
rect 2810 2870 2844 2880
rect 2810 2846 2844 2870
rect 2902 2870 2936 2880
rect 2902 2846 2936 2870
rect 2994 2870 3028 2880
rect 2994 2846 3028 2870
rect 3086 2870 3120 2880
rect 3086 2846 3120 2870
rect 3178 2870 3212 2880
rect 3178 2846 3212 2870
rect 3270 2870 3304 2880
rect 3270 2846 3304 2870
rect 3362 2870 3396 2880
rect 3362 2846 3396 2870
rect 3454 2870 3488 2880
rect 3454 2846 3488 2870
rect 3546 2870 3580 2880
rect 3546 2846 3580 2870
rect 3638 2870 3672 2880
rect 3638 2846 3672 2870
rect 3730 2870 3764 2880
rect 3730 2846 3764 2870
rect 3822 2870 3856 2880
rect 3822 2846 3856 2870
rect 3914 2870 3948 2880
rect 3914 2846 3948 2870
rect 4006 2870 4040 2880
rect 4006 2846 4040 2870
rect 4098 2870 4132 2880
rect 4098 2846 4132 2870
rect 4190 2870 4224 2880
rect 4190 2846 4224 2870
rect 4282 2870 4316 2880
rect 4282 2846 4316 2870
rect 4374 2870 4408 2880
rect 4374 2846 4408 2870
rect 4466 2870 4500 2880
rect 4466 2846 4500 2870
rect 4558 2870 4592 2880
rect 4558 2846 4592 2870
rect 4650 2870 4684 2880
rect 4650 2846 4684 2870
rect 4742 2870 4776 2880
rect 4742 2846 4776 2870
rect 4834 2870 4868 2880
rect 4834 2846 4868 2870
rect 4926 2870 4960 2880
rect 4926 2846 4960 2870
rect 5018 2870 5052 2880
rect 5018 2846 5052 2870
rect 5110 2870 5144 2880
rect 5110 2846 5144 2870
rect 5202 2870 5236 2880
rect 5202 2846 5236 2870
rect 5294 2870 5328 2880
rect 5294 2846 5328 2870
rect 5386 2870 5420 2880
rect 5386 2846 5420 2870
rect 5478 2870 5512 2880
rect 5478 2846 5512 2870
rect 5570 2870 5604 2880
rect 5570 2846 5604 2870
rect 5662 2870 5696 2880
rect 5662 2846 5696 2870
rect 5754 2870 5788 2880
rect 5754 2846 5788 2870
rect 5846 2870 5880 2880
rect 5846 2846 5880 2870
rect 5938 2870 5972 2880
rect 5938 2846 5972 2870
rect 6030 2870 6064 2880
rect 6030 2846 6064 2870
rect 6122 2870 6156 2880
rect 6122 2846 6156 2870
rect 6214 2870 6248 2880
rect 6214 2846 6248 2870
rect 6306 2870 6340 2880
rect 6306 2846 6340 2870
rect 6398 2870 6432 2880
rect 6398 2846 6432 2870
rect 6490 2870 6524 2880
rect 6490 2846 6524 2870
rect 6582 2870 6616 2880
rect 6582 2846 6616 2870
rect 6674 2870 6708 2880
rect 6674 2846 6708 2870
rect 6766 2870 6800 2880
rect 6766 2846 6800 2870
rect 6858 2870 6892 2880
rect 6858 2846 6892 2870
rect 6950 2870 6984 2880
rect 6950 2846 6984 2870
rect 7042 2870 7076 2880
rect 7042 2846 7076 2870
rect 7134 2870 7168 2880
rect 7134 2846 7168 2870
rect 7226 2870 7260 2880
rect 7226 2846 7260 2870
rect 7318 2870 7352 2880
rect 7318 2846 7352 2870
rect 7410 2870 7444 2880
rect 7410 2846 7444 2870
rect 7502 2870 7536 2880
rect 7502 2846 7536 2870
rect 7594 2870 7628 2880
rect 7594 2846 7628 2870
rect 7686 2870 7720 2880
rect 7686 2846 7720 2870
rect 7778 2870 7812 2880
rect 7778 2846 7812 2870
rect 7870 2870 7904 2880
rect 7870 2846 7904 2870
rect 7962 2870 7996 2880
rect 7962 2846 7996 2870
rect 8054 2870 8088 2880
rect 8054 2846 8088 2870
rect 8146 2870 8180 2880
rect 8146 2846 8180 2870
rect 8238 2870 8272 2880
rect 8238 2846 8272 2870
rect 8330 2870 8364 2880
rect 8330 2846 8364 2870
rect 8422 2870 8456 2880
rect 8422 2846 8456 2870
rect 8514 2870 8548 2880
rect 8514 2846 8548 2870
rect 8606 2870 8640 2880
rect 8606 2846 8640 2870
rect 8698 2870 8732 2880
rect 8698 2846 8732 2870
rect 8790 2870 8824 2880
rect 8790 2846 8824 2870
rect 8882 2870 8916 2880
rect 8882 2846 8916 2870
rect 8974 2870 9008 2880
rect 8974 2846 9008 2870
rect 9066 2870 9100 2880
rect 9066 2846 9100 2870
rect 9158 2870 9192 2880
rect 9158 2846 9192 2870
rect 9250 2870 9284 2880
rect 9250 2846 9284 2870
rect 9342 2870 9376 2880
rect 9342 2846 9376 2870
rect 9434 2870 9468 2880
rect 9434 2846 9468 2870
rect 9526 2870 9560 2880
rect 9526 2846 9560 2870
rect 9618 2870 9652 2880
rect 9618 2846 9652 2870
rect 9710 2870 9744 2880
rect 9710 2846 9744 2870
rect 9802 2870 9836 2880
rect 9802 2846 9836 2870
rect 9894 2870 9928 2880
rect 9894 2846 9928 2870
rect 9986 2870 10020 2880
rect 9986 2846 10020 2870
rect 10078 2870 10112 2880
rect 10078 2846 10112 2870
rect 10170 2870 10204 2880
rect 10170 2846 10204 2870
rect 10262 2870 10296 2880
rect 10262 2846 10296 2870
rect 10354 2870 10388 2880
rect 10354 2846 10388 2870
rect 10446 2870 10480 2880
rect 10446 2846 10480 2870
rect 10538 2870 10572 2880
rect 10538 2846 10572 2870
rect 10630 2870 10664 2880
rect 10630 2846 10664 2870
rect 10722 2870 10756 2880
rect 10722 2846 10756 2870
rect 10814 2870 10848 2880
rect 10814 2846 10848 2870
rect 10906 2870 10940 2880
rect 10906 2846 10940 2870
rect 10998 2870 11032 2880
rect 10998 2846 11032 2870
rect 11090 2870 11124 2880
rect 11090 2846 11124 2870
rect 11182 2870 11216 2880
rect 11182 2846 11216 2870
rect 11274 2870 11308 2880
rect 11274 2846 11308 2870
rect 11366 2870 11400 2880
rect 11366 2846 11400 2870
rect 11458 2870 11492 2880
rect 11458 2846 11492 2870
rect 11550 2870 11584 2880
rect 11550 2846 11584 2870
rect 11642 2870 11676 2880
rect 11642 2846 11676 2870
rect 11734 2870 11768 2880
rect 11734 2846 11768 2870
rect 11826 2870 11860 2880
rect 11826 2846 11860 2870
rect 11918 2870 11952 2880
rect 11918 2846 11952 2870
rect 12010 2870 12044 2880
rect 12010 2846 12044 2870
rect 12102 2870 12136 2880
rect 12102 2846 12136 2870
rect 12194 2870 12228 2880
rect 12194 2846 12228 2870
rect 12286 2870 12320 2880
rect 12286 2846 12320 2870
rect 12378 2870 12412 2880
rect 12378 2846 12412 2870
rect 12470 2870 12504 2880
rect 12470 2846 12504 2870
rect 12562 2870 12596 2880
rect 12562 2846 12596 2870
rect 12654 2870 12688 2880
rect 12654 2846 12688 2870
rect 12746 2870 12780 2880
rect 12746 2846 12780 2870
rect 12838 2870 12872 2880
rect 12838 2846 12872 2870
rect 12930 2870 12964 2880
rect 12930 2846 12964 2870
rect 1059 2414 1068 2447
rect 1068 2414 1093 2447
rect 1059 2413 1093 2414
rect 1613 2608 1647 2642
rect 1503 2538 1537 2572
rect 1889 2498 1914 2506
rect 1914 2498 1923 2506
rect 1889 2472 1923 2498
rect 2165 2684 2199 2710
rect 2165 2676 2178 2684
rect 2178 2676 2199 2684
rect 2257 2608 2291 2642
rect 2165 2540 2199 2574
rect 2901 2676 2935 2710
rect 2625 2498 2657 2506
rect 2657 2498 2659 2506
rect 2625 2472 2659 2498
rect 2813 2488 2829 2506
rect 2829 2488 2847 2506
rect 2813 2472 2847 2488
rect 3015 2598 3049 2632
rect 3177 2472 3211 2506
rect 3269 2676 3303 2710
rect 3450 2448 3484 2470
rect 3450 2436 3460 2448
rect 3460 2436 3484 2448
rect 4005 2608 4039 2642
rect 3896 2572 3930 2577
rect 3896 2543 3929 2572
rect 3929 2543 3930 2572
rect 4281 2498 4306 2506
rect 4306 2498 4315 2506
rect 4281 2472 4315 2498
rect 4557 2684 4591 2710
rect 4557 2676 4570 2684
rect 4570 2676 4591 2684
rect 4649 2608 4683 2642
rect 4557 2540 4591 2574
rect 5293 2676 5327 2710
rect 5017 2498 5049 2506
rect 5049 2498 5051 2506
rect 5017 2472 5051 2498
rect 5205 2488 5221 2506
rect 5221 2488 5239 2506
rect 5205 2472 5239 2488
rect 5396 2595 5430 2629
rect 5569 2472 5603 2506
rect 5661 2676 5695 2710
rect 5841 2448 5875 2469
rect 5841 2435 5852 2448
rect 5852 2435 5875 2448
rect 6397 2608 6431 2642
rect 6290 2572 6324 2577
rect 6290 2543 6321 2572
rect 6321 2543 6324 2572
rect 6673 2498 6698 2506
rect 6698 2498 6707 2506
rect 6673 2472 6707 2498
rect 6949 2684 6983 2710
rect 6949 2676 6962 2684
rect 6962 2676 6983 2684
rect 7041 2608 7075 2642
rect 6949 2540 6983 2574
rect 7685 2676 7719 2710
rect 7409 2498 7441 2506
rect 7441 2498 7443 2506
rect 7409 2472 7443 2498
rect 7597 2488 7613 2506
rect 7613 2488 7631 2506
rect 7597 2472 7631 2488
rect 7787 2599 7821 2633
rect 7961 2472 7995 2506
rect 8053 2676 8087 2710
rect 8236 2448 8270 2472
rect 8236 2438 8244 2448
rect 8244 2438 8270 2448
rect 8789 2608 8823 2642
rect 8682 2572 8716 2578
rect 8682 2544 8713 2572
rect 8713 2544 8716 2572
rect 9065 2498 9090 2506
rect 9090 2498 9099 2506
rect 9065 2472 9099 2498
rect 9341 2684 9375 2710
rect 9341 2676 9354 2684
rect 9354 2676 9375 2684
rect 9433 2608 9467 2642
rect 9341 2540 9375 2574
rect 10077 2676 10111 2710
rect 9801 2498 9833 2506
rect 9833 2498 9835 2506
rect 9801 2472 9835 2498
rect 9989 2488 10005 2506
rect 10005 2488 10023 2506
rect 9989 2472 10023 2488
rect 10176 2600 10210 2634
rect 10353 2472 10387 2506
rect 10445 2676 10479 2710
rect 10625 2448 10659 2470
rect 10625 2436 10636 2448
rect 10636 2436 10659 2448
rect 11181 2608 11215 2642
rect 11075 2572 11109 2579
rect 11075 2545 11105 2572
rect 11105 2545 11109 2572
rect 11457 2498 11482 2506
rect 11482 2498 11491 2506
rect 11457 2472 11491 2498
rect 11733 2684 11767 2710
rect 11733 2676 11746 2684
rect 11746 2676 11767 2684
rect 11825 2608 11859 2642
rect 11733 2540 11767 2574
rect 12469 2676 12503 2710
rect 12193 2498 12225 2506
rect 12225 2498 12227 2506
rect 12193 2472 12227 2498
rect 12381 2488 12397 2506
rect 12397 2488 12415 2506
rect 12381 2472 12415 2488
rect 12570 2600 12604 2634
rect 12745 2472 12779 2506
rect 12837 2676 12871 2710
rect 12927 2549 12961 2583
rect 1062 2312 1096 2336
rect 1062 2302 1096 2312
rect 1154 2312 1188 2336
rect 1154 2302 1188 2312
rect 1246 2312 1280 2336
rect 1246 2302 1280 2312
rect 1338 2312 1372 2336
rect 1338 2302 1372 2312
rect 1430 2312 1464 2336
rect 1430 2302 1464 2312
rect 1522 2312 1556 2336
rect 1522 2302 1556 2312
rect 1614 2312 1648 2336
rect 1614 2302 1648 2312
rect 1706 2312 1740 2336
rect 1706 2302 1740 2312
rect 1798 2312 1832 2336
rect 1798 2302 1832 2312
rect 1890 2312 1924 2336
rect 1890 2302 1924 2312
rect 1982 2312 2016 2336
rect 1982 2302 2016 2312
rect 2074 2312 2108 2336
rect 2074 2302 2108 2312
rect 2166 2312 2200 2336
rect 2166 2302 2200 2312
rect 2258 2312 2292 2336
rect 2258 2302 2292 2312
rect 2350 2312 2384 2336
rect 2350 2302 2384 2312
rect 2442 2312 2476 2336
rect 2442 2302 2476 2312
rect 2534 2312 2568 2336
rect 2534 2302 2568 2312
rect 2626 2312 2660 2336
rect 2626 2302 2660 2312
rect 2718 2312 2752 2336
rect 2718 2302 2752 2312
rect 2810 2312 2844 2336
rect 2810 2302 2844 2312
rect 2902 2312 2936 2336
rect 2902 2302 2936 2312
rect 2994 2312 3028 2336
rect 2994 2302 3028 2312
rect 3086 2312 3120 2336
rect 3086 2302 3120 2312
rect 3178 2312 3212 2336
rect 3178 2302 3212 2312
rect 3270 2312 3304 2336
rect 3270 2302 3304 2312
rect 3362 2312 3396 2336
rect 3362 2302 3396 2312
rect 3454 2312 3488 2336
rect 3454 2302 3488 2312
rect 3546 2312 3580 2336
rect 3546 2302 3580 2312
rect 3638 2312 3672 2336
rect 3638 2302 3672 2312
rect 3730 2312 3764 2336
rect 3730 2302 3764 2312
rect 3822 2312 3856 2336
rect 3822 2302 3856 2312
rect 3914 2312 3948 2336
rect 3914 2302 3948 2312
rect 4006 2312 4040 2336
rect 4006 2302 4040 2312
rect 4098 2312 4132 2336
rect 4098 2302 4132 2312
rect 4190 2312 4224 2336
rect 4190 2302 4224 2312
rect 4282 2312 4316 2336
rect 4282 2302 4316 2312
rect 4374 2312 4408 2336
rect 4374 2302 4408 2312
rect 4466 2312 4500 2336
rect 4466 2302 4500 2312
rect 4558 2312 4592 2336
rect 4558 2302 4592 2312
rect 4650 2312 4684 2336
rect 4650 2302 4684 2312
rect 4742 2312 4776 2336
rect 4742 2302 4776 2312
rect 4834 2312 4868 2336
rect 4834 2302 4868 2312
rect 4926 2312 4960 2336
rect 4926 2302 4960 2312
rect 5018 2312 5052 2336
rect 5018 2302 5052 2312
rect 5110 2312 5144 2336
rect 5110 2302 5144 2312
rect 5202 2312 5236 2336
rect 5202 2302 5236 2312
rect 5294 2312 5328 2336
rect 5294 2302 5328 2312
rect 5386 2312 5420 2336
rect 5386 2302 5420 2312
rect 5478 2312 5512 2336
rect 5478 2302 5512 2312
rect 5570 2312 5604 2336
rect 5570 2302 5604 2312
rect 5662 2312 5696 2336
rect 5662 2302 5696 2312
rect 5754 2312 5788 2336
rect 5754 2302 5788 2312
rect 5846 2312 5880 2336
rect 5846 2302 5880 2312
rect 5938 2312 5972 2336
rect 5938 2302 5972 2312
rect 6030 2312 6064 2336
rect 6030 2302 6064 2312
rect 6122 2312 6156 2336
rect 6122 2302 6156 2312
rect 6214 2312 6248 2336
rect 6214 2302 6248 2312
rect 6306 2312 6340 2336
rect 6306 2302 6340 2312
rect 6398 2312 6432 2336
rect 6398 2302 6432 2312
rect 6490 2312 6524 2336
rect 6490 2302 6524 2312
rect 6582 2312 6616 2336
rect 6582 2302 6616 2312
rect 6674 2312 6708 2336
rect 6674 2302 6708 2312
rect 6766 2312 6800 2336
rect 6766 2302 6800 2312
rect 6858 2312 6892 2336
rect 6858 2302 6892 2312
rect 6950 2312 6984 2336
rect 6950 2302 6984 2312
rect 7042 2312 7076 2336
rect 7042 2302 7076 2312
rect 7134 2312 7168 2336
rect 7134 2302 7168 2312
rect 7226 2312 7260 2336
rect 7226 2302 7260 2312
rect 7318 2312 7352 2336
rect 7318 2302 7352 2312
rect 7410 2312 7444 2336
rect 7410 2302 7444 2312
rect 7502 2312 7536 2336
rect 7502 2302 7536 2312
rect 7594 2312 7628 2336
rect 7594 2302 7628 2312
rect 7686 2312 7720 2336
rect 7686 2302 7720 2312
rect 7778 2312 7812 2336
rect 7778 2302 7812 2312
rect 7870 2312 7904 2336
rect 7870 2302 7904 2312
rect 7962 2312 7996 2336
rect 7962 2302 7996 2312
rect 8054 2312 8088 2336
rect 8054 2302 8088 2312
rect 8146 2312 8180 2336
rect 8146 2302 8180 2312
rect 8238 2312 8272 2336
rect 8238 2302 8272 2312
rect 8330 2312 8364 2336
rect 8330 2302 8364 2312
rect 8422 2312 8456 2336
rect 8422 2302 8456 2312
rect 8514 2312 8548 2336
rect 8514 2302 8548 2312
rect 8606 2312 8640 2336
rect 8606 2302 8640 2312
rect 8698 2312 8732 2336
rect 8698 2302 8732 2312
rect 8790 2312 8824 2336
rect 8790 2302 8824 2312
rect 8882 2312 8916 2336
rect 8882 2302 8916 2312
rect 8974 2312 9008 2336
rect 8974 2302 9008 2312
rect 9066 2312 9100 2336
rect 9066 2302 9100 2312
rect 9158 2312 9192 2336
rect 9158 2302 9192 2312
rect 9250 2312 9284 2336
rect 9250 2302 9284 2312
rect 9342 2312 9376 2336
rect 9342 2302 9376 2312
rect 9434 2312 9468 2336
rect 9434 2302 9468 2312
rect 9526 2312 9560 2336
rect 9526 2302 9560 2312
rect 9618 2312 9652 2336
rect 9618 2302 9652 2312
rect 9710 2312 9744 2336
rect 9710 2302 9744 2312
rect 9802 2312 9836 2336
rect 9802 2302 9836 2312
rect 9894 2312 9928 2336
rect 9894 2302 9928 2312
rect 9986 2312 10020 2336
rect 9986 2302 10020 2312
rect 10078 2312 10112 2336
rect 10078 2302 10112 2312
rect 10170 2312 10204 2336
rect 10170 2302 10204 2312
rect 10262 2312 10296 2336
rect 10262 2302 10296 2312
rect 10354 2312 10388 2336
rect 10354 2302 10388 2312
rect 10446 2312 10480 2336
rect 10446 2302 10480 2312
rect 10538 2312 10572 2336
rect 10538 2302 10572 2312
rect 10630 2312 10664 2336
rect 10630 2302 10664 2312
rect 10722 2312 10756 2336
rect 10722 2302 10756 2312
rect 10814 2312 10848 2336
rect 10814 2302 10848 2312
rect 10906 2312 10940 2336
rect 10906 2302 10940 2312
rect 10998 2312 11032 2336
rect 10998 2302 11032 2312
rect 11090 2312 11124 2336
rect 11090 2302 11124 2312
rect 11182 2312 11216 2336
rect 11182 2302 11216 2312
rect 11274 2312 11308 2336
rect 11274 2302 11308 2312
rect 11366 2312 11400 2336
rect 11366 2302 11400 2312
rect 11458 2312 11492 2336
rect 11458 2302 11492 2312
rect 11550 2312 11584 2336
rect 11550 2302 11584 2312
rect 11642 2312 11676 2336
rect 11642 2302 11676 2312
rect 11734 2312 11768 2336
rect 11734 2302 11768 2312
rect 11826 2312 11860 2336
rect 11826 2302 11860 2312
rect 11918 2312 11952 2336
rect 11918 2302 11952 2312
rect 12010 2312 12044 2336
rect 12010 2302 12044 2312
rect 12102 2312 12136 2336
rect 12102 2302 12136 2312
rect 12194 2312 12228 2336
rect 12194 2302 12228 2312
rect 12286 2312 12320 2336
rect 12286 2302 12320 2312
rect 12378 2312 12412 2336
rect 12378 2302 12412 2312
rect 12470 2312 12504 2336
rect 12470 2302 12504 2312
rect 12562 2312 12596 2336
rect 12562 2302 12596 2312
rect 12654 2312 12688 2336
rect 12654 2302 12688 2312
rect 12746 2312 12780 2336
rect 12746 2302 12780 2312
rect 12838 2312 12872 2336
rect 12838 2302 12872 2312
rect 12930 2312 12964 2336
rect 12930 2302 12964 2312
<< metal1 >>
rect 612 6218 4314 6219
rect 290 6188 4314 6218
rect 290 6174 1064 6188
rect 290 6028 428 6174
rect 578 6158 1064 6174
rect 578 6028 740 6158
rect 290 6012 740 6028
rect 890 6154 1064 6158
rect 1098 6154 1156 6188
rect 1190 6154 1248 6188
rect 1282 6154 1340 6188
rect 1374 6154 1432 6188
rect 1466 6154 1524 6188
rect 1558 6154 1616 6188
rect 1650 6154 1708 6188
rect 1742 6154 1800 6188
rect 1834 6154 2324 6188
rect 2358 6154 2416 6188
rect 2450 6154 2508 6188
rect 2542 6154 2600 6188
rect 2634 6154 2692 6188
rect 2726 6154 2784 6188
rect 2818 6154 2876 6188
rect 2910 6154 2968 6188
rect 3002 6154 3060 6188
rect 3094 6154 3152 6188
rect 3186 6154 3244 6188
rect 3278 6154 3336 6188
rect 3370 6154 3428 6188
rect 3462 6154 3520 6188
rect 3554 6154 3612 6188
rect 3646 6154 3704 6188
rect 3738 6154 3796 6188
rect 3830 6154 3888 6188
rect 3922 6154 3980 6188
rect 4014 6154 4072 6188
rect 4106 6154 4314 6188
rect 890 6123 4314 6154
rect 890 6012 954 6123
rect 2771 6086 2829 6092
rect 2771 6052 2783 6086
rect 2817 6083 2829 6086
rect 3231 6086 3289 6092
rect 3231 6083 3243 6086
rect 2817 6055 3243 6083
rect 2817 6052 2829 6055
rect 2771 6046 2829 6052
rect 3231 6052 3243 6055
rect 3277 6052 3289 6086
rect 3231 6046 3289 6052
rect 3415 6086 3473 6092
rect 3415 6052 3427 6086
rect 3461 6083 3473 6086
rect 3691 6086 3749 6092
rect 3691 6083 3703 6086
rect 3461 6055 3703 6083
rect 3461 6052 3473 6055
rect 3415 6046 3473 6052
rect 3691 6052 3703 6055
rect 3737 6052 3749 6086
rect 3691 6046 3749 6052
rect 290 5988 954 6012
rect 2955 6018 3013 6024
rect 2955 5984 2967 6018
rect 3001 6015 3013 6018
rect 3783 6018 3841 6024
rect 3783 6015 3795 6018
rect 3001 5987 3795 6015
rect 3001 5984 3013 5987
rect 2955 5978 3013 5984
rect 3783 5984 3795 5987
rect 3829 5984 3841 6018
rect 3783 5978 3841 5984
rect 459 5947 493 5952
rect 2863 5950 2921 5956
rect 2863 5947 2875 5950
rect 459 5919 2875 5947
rect 459 5918 493 5919
rect 2863 5916 2875 5919
rect 2909 5947 2921 5950
rect 3875 5950 3933 5956
rect 3875 5947 3887 5950
rect 2909 5919 3887 5947
rect 2909 5916 2921 5919
rect 2863 5910 2921 5916
rect 3875 5916 3887 5919
rect 3921 5947 3933 5950
rect 4059 5950 4118 5956
rect 4059 5947 4071 5950
rect 3921 5919 4071 5947
rect 3921 5916 3933 5919
rect 3875 5910 3933 5916
rect 4059 5916 4071 5919
rect 4105 5916 4118 5950
rect 4059 5910 4118 5916
rect 8120 5903 8173 5910
rect 1056 5883 1122 5890
rect 462 5881 496 5882
rect 1056 5881 1068 5883
rect 462 5853 1068 5881
rect 462 5848 496 5853
rect 1056 5849 1068 5853
rect 1102 5849 1122 5883
rect 1056 5838 1122 5849
rect 1690 5839 1697 5891
rect 1749 5839 1758 5891
rect 2013 5890 2079 5891
rect 2013 5838 2020 5890
rect 2072 5876 2079 5890
rect 2397 5881 2455 5886
rect 3124 5884 3184 5890
rect 2397 5880 2457 5881
rect 2397 5876 2410 5880
rect 2072 5848 2410 5876
rect 2072 5838 2079 5848
rect 2397 5846 2410 5848
rect 2444 5846 2457 5880
rect 2397 5845 2457 5846
rect 3124 5850 3138 5884
rect 3172 5881 3184 5884
rect 3172 5853 8120 5881
rect 3172 5850 3184 5853
rect 2397 5840 2455 5845
rect 3124 5840 3184 5850
rect 8172 5851 8173 5903
rect 8120 5844 8173 5851
rect 10528 5827 10581 5834
rect 464 5810 498 5816
rect 3503 5813 3566 5820
rect 3503 5810 3519 5813
rect 463 5782 3519 5810
rect 3503 5779 3519 5782
rect 3553 5779 3566 5813
rect 3503 5772 3566 5779
rect 3596 5769 3602 5821
rect 3654 5769 3660 5821
rect 3727 5787 10528 5815
rect 2766 5743 2825 5750
rect 2766 5709 2778 5743
rect 2812 5731 2825 5743
rect 3727 5741 3756 5787
rect 10580 5775 10581 5827
rect 10528 5768 10581 5775
rect 3727 5731 3755 5741
rect 2812 5709 3755 5731
rect 2766 5703 3755 5709
rect 3875 5707 3882 5759
rect 3934 5734 3941 5759
rect 5724 5734 5731 5759
rect 3934 5707 5731 5734
rect 5783 5707 5790 5759
rect 3875 5706 5790 5707
rect 502 5675 582 5676
rect 420 5665 12039 5675
rect 12278 5665 13332 5672
rect 420 5644 13332 5665
rect 420 5640 1064 5644
rect 416 5610 1064 5640
rect 1098 5610 1156 5644
rect 1190 5610 1248 5644
rect 1282 5610 1340 5644
rect 1374 5610 1432 5644
rect 1466 5610 1524 5644
rect 1558 5610 1616 5644
rect 1650 5610 1708 5644
rect 1742 5610 1800 5644
rect 1834 5610 2324 5644
rect 2358 5610 2416 5644
rect 2450 5610 2508 5644
rect 2542 5610 2600 5644
rect 2634 5610 2692 5644
rect 2726 5610 2784 5644
rect 2818 5610 2876 5644
rect 2910 5610 2968 5644
rect 3002 5610 3060 5644
rect 3094 5610 3152 5644
rect 3186 5610 3244 5644
rect 3278 5610 3336 5644
rect 3370 5610 3428 5644
rect 3462 5610 3520 5644
rect 3554 5610 3612 5644
rect 3646 5610 3704 5644
rect 3738 5610 3796 5644
rect 3830 5610 3888 5644
rect 3922 5610 3980 5644
rect 4014 5610 4072 5644
rect 4106 5610 13332 5644
rect 416 5602 13332 5610
rect 420 5589 13332 5602
rect 420 5579 12039 5589
rect 13082 5560 13332 5589
rect 1053 5516 1119 5517
rect 1053 5505 1060 5516
rect 1039 5477 1060 5505
rect 1053 5464 1060 5477
rect 1112 5505 1119 5516
rect 1714 5516 1780 5517
rect 1714 5505 1721 5516
rect 1112 5477 1721 5505
rect 1112 5464 1119 5477
rect 1714 5464 1721 5477
rect 1773 5505 1780 5516
rect 3444 5516 3510 5517
rect 3444 5505 3451 5516
rect 1773 5477 3451 5505
rect 1773 5464 1780 5477
rect 3444 5464 3451 5477
rect 3503 5505 3510 5516
rect 5827 5516 5893 5517
rect 5827 5505 5834 5516
rect 3503 5477 5834 5505
rect 3503 5464 3510 5477
rect 5827 5464 5834 5477
rect 5886 5505 5893 5516
rect 8222 5516 8288 5517
rect 8222 5505 8229 5516
rect 5886 5477 8229 5505
rect 5886 5464 5893 5477
rect 8222 5464 8229 5477
rect 8281 5505 8288 5516
rect 10617 5516 10683 5517
rect 10617 5505 10624 5516
rect 8281 5477 10624 5505
rect 8281 5464 8288 5477
rect 10617 5464 10624 5477
rect 10676 5505 10683 5516
rect 12913 5516 12979 5517
rect 12913 5505 12920 5516
rect 10676 5477 12920 5505
rect 10676 5464 10683 5477
rect 12913 5464 12920 5477
rect 12972 5464 12979 5516
rect 13082 5414 13146 5560
rect 13296 5414 13332 5560
rect 13082 5402 13332 5414
rect 412 5374 13332 5402
rect 412 5345 13030 5346
rect 290 5315 13030 5345
rect 290 5281 1063 5315
rect 1097 5281 1155 5315
rect 1189 5281 1247 5315
rect 1281 5281 1339 5315
rect 1373 5281 1431 5315
rect 1465 5281 1523 5315
rect 1557 5281 1615 5315
rect 1649 5281 1707 5315
rect 1741 5281 1799 5315
rect 1833 5281 1891 5315
rect 1925 5281 1983 5315
rect 2017 5281 2075 5315
rect 2109 5281 2167 5315
rect 2201 5281 2259 5315
rect 2293 5281 2351 5315
rect 2385 5281 2443 5315
rect 2477 5281 2535 5315
rect 2569 5281 2627 5315
rect 2661 5281 2719 5315
rect 2753 5281 2811 5315
rect 2845 5281 2903 5315
rect 2937 5281 2995 5315
rect 3029 5281 3087 5315
rect 3121 5281 3179 5315
rect 3213 5281 3271 5315
rect 3305 5281 3363 5315
rect 3397 5281 3455 5315
rect 3489 5281 3547 5315
rect 3581 5281 3639 5315
rect 3673 5281 3731 5315
rect 3765 5281 3823 5315
rect 3857 5281 3915 5315
rect 3949 5281 4007 5315
rect 4041 5281 4099 5315
rect 4133 5281 4191 5315
rect 4225 5281 4283 5315
rect 4317 5281 4375 5315
rect 4409 5281 4467 5315
rect 4501 5281 4559 5315
rect 4593 5281 4651 5315
rect 4685 5281 4743 5315
rect 4777 5281 4835 5315
rect 4869 5281 4927 5315
rect 4961 5281 5019 5315
rect 5053 5281 5111 5315
rect 5145 5281 5203 5315
rect 5237 5281 5295 5315
rect 5329 5281 5387 5315
rect 5421 5281 5479 5315
rect 5513 5281 5571 5315
rect 5605 5281 5663 5315
rect 5697 5281 5755 5315
rect 5789 5281 5847 5315
rect 5881 5281 5939 5315
rect 5973 5281 6031 5315
rect 6065 5281 6123 5315
rect 6157 5281 6215 5315
rect 6249 5281 6307 5315
rect 6341 5281 6399 5315
rect 6433 5281 6491 5315
rect 6525 5281 6583 5315
rect 6617 5281 6675 5315
rect 6709 5281 6767 5315
rect 6801 5281 6859 5315
rect 6893 5281 6951 5315
rect 6985 5281 7043 5315
rect 7077 5281 7135 5315
rect 7169 5281 7227 5315
rect 7261 5281 7319 5315
rect 7353 5281 7411 5315
rect 7445 5281 7503 5315
rect 7537 5281 7595 5315
rect 7629 5281 7687 5315
rect 7721 5281 7779 5315
rect 7813 5281 7871 5315
rect 7905 5281 7963 5315
rect 7997 5281 8055 5315
rect 8089 5281 8147 5315
rect 8181 5281 8239 5315
rect 8273 5281 8331 5315
rect 8365 5281 8423 5315
rect 8457 5281 8515 5315
rect 8549 5281 8607 5315
rect 8641 5281 8699 5315
rect 8733 5281 8791 5315
rect 8825 5281 8883 5315
rect 8917 5281 8975 5315
rect 9009 5281 9067 5315
rect 9101 5281 9159 5315
rect 9193 5281 9251 5315
rect 9285 5281 9343 5315
rect 9377 5281 9435 5315
rect 9469 5281 9527 5315
rect 9561 5281 9619 5315
rect 9653 5281 9711 5315
rect 9745 5281 9803 5315
rect 9837 5281 9895 5315
rect 9929 5281 9987 5315
rect 10021 5281 10079 5315
rect 10113 5281 10171 5315
rect 10205 5281 10263 5315
rect 10297 5281 10355 5315
rect 10389 5281 10447 5315
rect 10481 5281 10539 5315
rect 10573 5281 10631 5315
rect 10665 5281 10723 5315
rect 10757 5281 10815 5315
rect 10849 5281 10907 5315
rect 10941 5281 10999 5315
rect 11033 5281 11091 5315
rect 11125 5281 11183 5315
rect 11217 5281 11275 5315
rect 11309 5281 11367 5315
rect 11401 5281 11459 5315
rect 11493 5281 11551 5315
rect 11585 5281 11643 5315
rect 11677 5281 11735 5315
rect 11769 5281 11827 5315
rect 11861 5281 11919 5315
rect 11953 5281 12011 5315
rect 12045 5281 12103 5315
rect 12137 5281 12195 5315
rect 12229 5281 12287 5315
rect 12321 5281 12379 5315
rect 12413 5281 12471 5315
rect 12505 5281 12563 5315
rect 12597 5281 12655 5315
rect 12689 5281 12747 5315
rect 12781 5281 12839 5315
rect 12873 5281 12931 5315
rect 12965 5293 13030 5315
rect 12965 5281 13031 5293
rect 290 5250 13031 5281
rect 290 5226 966 5250
rect 290 5214 798 5226
rect 290 5068 492 5214
rect 642 5080 798 5214
rect 948 5080 966 5226
rect 12557 5215 12589 5216
rect 12557 5211 12638 5215
rect 12557 5159 12563 5211
rect 12615 5201 12638 5211
rect 12918 5201 12977 5207
rect 12615 5167 12931 5201
rect 12965 5167 12977 5201
rect 12615 5166 12977 5167
rect 12615 5159 12638 5166
rect 12918 5160 12977 5166
rect 1144 5145 1202 5151
rect 1144 5111 1156 5145
rect 1190 5142 1202 5145
rect 1512 5145 1570 5151
rect 1512 5142 1524 5145
rect 1190 5114 1524 5142
rect 1190 5111 1202 5114
rect 1144 5105 1202 5111
rect 1512 5111 1524 5114
rect 1558 5142 1570 5145
rect 2248 5145 2306 5151
rect 2248 5142 2260 5145
rect 1558 5114 2260 5142
rect 1558 5111 1570 5114
rect 1512 5105 1570 5111
rect 2248 5111 2260 5114
rect 2294 5111 2306 5145
rect 2248 5105 2306 5111
rect 3536 5145 3594 5151
rect 3536 5111 3548 5145
rect 3582 5142 3594 5145
rect 3904 5145 3962 5151
rect 3904 5142 3916 5145
rect 3582 5114 3916 5142
rect 3582 5111 3594 5114
rect 3536 5105 3594 5111
rect 3904 5111 3916 5114
rect 3950 5142 3962 5145
rect 4640 5145 4698 5151
rect 4640 5142 4652 5145
rect 3950 5114 4652 5142
rect 3950 5111 3962 5114
rect 3904 5105 3962 5111
rect 4640 5111 4652 5114
rect 4686 5111 4698 5145
rect 4640 5105 4698 5111
rect 5928 5145 5986 5151
rect 5928 5111 5940 5145
rect 5974 5142 5986 5145
rect 6296 5145 6354 5151
rect 6296 5142 6308 5145
rect 5974 5114 6308 5142
rect 5974 5111 5986 5114
rect 5928 5105 5986 5111
rect 6296 5111 6308 5114
rect 6342 5142 6354 5145
rect 7032 5145 7090 5151
rect 7032 5142 7044 5145
rect 6342 5114 7044 5142
rect 6342 5111 6354 5114
rect 6296 5105 6354 5111
rect 7032 5111 7044 5114
rect 7078 5111 7090 5145
rect 7032 5105 7090 5111
rect 8320 5145 8378 5151
rect 8320 5111 8332 5145
rect 8366 5142 8378 5145
rect 8688 5145 8746 5151
rect 8688 5142 8700 5145
rect 8366 5114 8700 5142
rect 8366 5111 8378 5114
rect 8320 5105 8378 5111
rect 8688 5111 8700 5114
rect 8734 5142 8746 5145
rect 9424 5145 9482 5151
rect 9424 5142 9436 5145
rect 8734 5114 9436 5142
rect 8734 5111 8746 5114
rect 8688 5105 8746 5111
rect 9424 5111 9436 5114
rect 9470 5111 9482 5145
rect 9424 5105 9482 5111
rect 10712 5145 10770 5151
rect 10712 5111 10724 5145
rect 10758 5142 10770 5145
rect 11080 5145 11138 5151
rect 11080 5142 11092 5145
rect 10758 5114 11092 5142
rect 10758 5111 10770 5114
rect 10712 5105 10770 5111
rect 11080 5111 11092 5114
rect 11126 5142 11138 5145
rect 11816 5145 11874 5151
rect 12557 5150 12638 5159
rect 12557 5149 12589 5150
rect 11816 5142 11828 5145
rect 11126 5114 11828 5142
rect 11126 5111 11138 5114
rect 11080 5105 11138 5111
rect 11816 5111 11828 5114
rect 11862 5111 11874 5145
rect 11816 5105 11874 5111
rect 13068 5134 13332 5226
rect 642 5068 966 5080
rect 290 4958 966 5068
rect 1411 5074 1474 5081
rect 2015 5074 2022 5086
rect 1411 5040 1428 5074
rect 1462 5046 2022 5074
rect 1462 5040 1474 5046
rect 1411 5034 1474 5040
rect 2015 5034 2022 5046
rect 2074 5034 2081 5086
rect 2156 5077 2214 5083
rect 2156 5043 2168 5077
rect 2202 5074 2214 5077
rect 2800 5077 2858 5083
rect 2800 5074 2812 5077
rect 2202 5046 2812 5074
rect 2202 5043 2214 5046
rect 2156 5037 2214 5043
rect 2800 5043 2812 5046
rect 2846 5043 2858 5077
rect 2800 5037 2858 5043
rect 3356 5081 3415 5087
rect 3356 5047 3368 5081
rect 3402 5077 3415 5081
rect 3767 5077 3826 5083
rect 3402 5049 3779 5077
rect 3402 5047 3415 5049
rect 3356 5040 3415 5047
rect 3767 5043 3779 5049
rect 3813 5043 3826 5077
rect 3767 5036 3826 5043
rect 4548 5077 4606 5083
rect 4548 5043 4560 5077
rect 4594 5074 4606 5077
rect 5192 5077 5250 5083
rect 5192 5074 5204 5077
rect 4594 5046 5204 5074
rect 4594 5043 4606 5046
rect 4548 5037 4606 5043
rect 5192 5043 5204 5046
rect 5238 5043 5250 5077
rect 5192 5037 5250 5043
rect 5745 5080 5804 5086
rect 5745 5046 5757 5080
rect 5791 5076 5804 5080
rect 6156 5076 6215 5082
rect 5791 5048 6168 5076
rect 5791 5046 5804 5048
rect 5745 5039 5804 5046
rect 6156 5042 6168 5048
rect 6202 5042 6215 5076
rect 6156 5035 6215 5042
rect 6940 5077 6998 5083
rect 6940 5043 6952 5077
rect 6986 5074 6998 5077
rect 7584 5077 7642 5083
rect 7584 5074 7596 5077
rect 6986 5046 7596 5074
rect 6986 5043 6998 5046
rect 6940 5037 6998 5043
rect 7584 5043 7596 5046
rect 7630 5043 7642 5077
rect 7584 5037 7642 5043
rect 8140 5078 8199 5084
rect 8140 5044 8152 5078
rect 8186 5074 8199 5078
rect 8551 5074 8610 5080
rect 8186 5046 8563 5074
rect 8186 5044 8199 5046
rect 8140 5037 8199 5044
rect 8551 5040 8563 5046
rect 8597 5040 8610 5074
rect 8551 5033 8610 5040
rect 9332 5077 9390 5083
rect 9332 5043 9344 5077
rect 9378 5074 9390 5077
rect 9976 5077 10034 5083
rect 9976 5074 9988 5077
rect 9378 5046 9988 5074
rect 9378 5043 9390 5046
rect 9332 5037 9390 5043
rect 9976 5043 9988 5046
rect 10022 5043 10034 5077
rect 9976 5037 10034 5043
rect 10531 5077 10590 5083
rect 10531 5043 10543 5077
rect 10577 5073 10590 5077
rect 10942 5073 11001 5079
rect 10577 5045 10954 5073
rect 10577 5043 10590 5045
rect 10531 5036 10590 5043
rect 10942 5039 10954 5045
rect 10988 5039 11001 5073
rect 10942 5032 11001 5039
rect 11724 5077 11782 5083
rect 11724 5043 11736 5077
rect 11770 5074 11782 5077
rect 12368 5077 12426 5083
rect 12368 5074 12380 5077
rect 11770 5046 12380 5074
rect 11770 5043 11782 5046
rect 11724 5037 11782 5043
rect 12368 5043 12380 5046
rect 12414 5043 12426 5077
rect 12368 5037 12426 5043
rect 2248 5009 2306 5015
rect 2248 5006 2260 5009
rect 1052 5003 1118 5004
rect 1052 4951 1059 5003
rect 1111 4951 1118 5003
rect 1619 4978 2260 5006
rect 1619 4947 1658 4978
rect 2248 4975 2260 4978
rect 2294 4975 2306 5009
rect 4640 5009 4698 5015
rect 4640 5006 4652 5009
rect 2248 4969 2306 4975
rect 3442 5003 3508 5004
rect 3442 4951 3449 5003
rect 3501 4951 3508 5003
rect 4011 4978 4652 5006
rect 2520 4948 2586 4949
rect 1236 4941 1294 4947
rect 1236 4907 1248 4941
rect 1282 4938 1294 4941
rect 1600 4941 1658 4947
rect 1600 4938 1612 4941
rect 1282 4910 1612 4938
rect 1282 4907 1294 4910
rect 1236 4901 1294 4907
rect 1600 4907 1612 4910
rect 1646 4907 1658 4941
rect 1600 4901 1658 4907
rect 1788 4941 1846 4947
rect 1788 4907 1800 4941
rect 1834 4938 1846 4941
rect 2520 4938 2527 4948
rect 1834 4910 2527 4938
rect 1834 4907 1846 4910
rect 1788 4901 1846 4907
rect 2520 4896 2527 4910
rect 2579 4896 2586 4948
rect 4011 4947 4050 4978
rect 4640 4975 4652 4978
rect 4686 4975 4698 5009
rect 4640 4969 4698 4975
rect 5286 4970 5293 5022
rect 5345 4970 5351 5022
rect 7686 5021 7739 5028
rect 7032 5009 7090 5015
rect 7032 5006 7044 5009
rect 5835 5004 5901 5005
rect 5835 4952 5842 5004
rect 5894 4952 5901 5004
rect 6403 4978 7044 5006
rect 6403 4947 6442 4978
rect 7032 4975 7044 4978
rect 7078 4975 7090 5009
rect 7032 4969 7090 4975
rect 7738 4969 7739 5021
rect 10077 5023 10130 5030
rect 9424 5009 9482 5015
rect 9424 5006 9436 5009
rect 7686 4962 7739 4969
rect 8227 5003 8293 5004
rect 8227 4951 8234 5003
rect 8286 4951 8293 5003
rect 8795 4978 9436 5006
rect 8795 4947 8834 4978
rect 9424 4975 9436 4978
rect 9470 4975 9482 5009
rect 9424 4969 9482 4975
rect 10129 4971 10130 5023
rect 12468 5021 12521 5028
rect 11816 5009 11874 5015
rect 11816 5006 11828 5009
rect 10077 4964 10130 4971
rect 10622 5005 10688 5006
rect 10622 4953 10629 5005
rect 10681 4953 10688 5005
rect 11187 4978 11828 5006
rect 11187 4947 11226 4978
rect 11816 4975 11828 4978
rect 11862 4975 11874 5009
rect 11816 4969 11874 4975
rect 12520 4969 12521 5021
rect 12468 4962 12521 4969
rect 13068 4988 13146 5134
rect 13296 4988 13332 5134
rect 3628 4941 3686 4947
rect 3628 4907 3640 4941
rect 3674 4938 3686 4941
rect 3992 4941 4050 4947
rect 3992 4938 4004 4941
rect 3674 4910 4004 4938
rect 3674 4907 3686 4910
rect 3628 4901 3686 4907
rect 3992 4907 4004 4910
rect 4038 4907 4050 4941
rect 3992 4901 4050 4907
rect 4180 4941 4238 4947
rect 4180 4907 4192 4941
rect 4226 4938 4238 4941
rect 4916 4941 4974 4947
rect 4916 4938 4928 4941
rect 4226 4910 4928 4938
rect 4226 4907 4238 4910
rect 4180 4901 4238 4907
rect 4916 4907 4928 4910
rect 4962 4907 4974 4941
rect 6020 4941 6078 4947
rect 5576 4915 5629 4922
rect 4916 4901 4974 4907
rect 5460 4904 5524 4910
rect 3070 4890 3136 4891
rect 3070 4838 3077 4890
rect 3129 4838 3136 4890
rect 5460 4852 5467 4904
rect 5519 4852 5524 4904
rect 5576 4863 5577 4915
rect 5737 4911 5798 4915
rect 5736 4906 5798 4911
rect 5629 4872 5748 4906
rect 5782 4872 5798 4906
rect 6020 4907 6032 4941
rect 6066 4938 6078 4941
rect 6384 4941 6442 4947
rect 6384 4938 6396 4941
rect 6066 4910 6396 4938
rect 6066 4907 6078 4910
rect 6020 4901 6078 4907
rect 6384 4907 6396 4910
rect 6430 4907 6442 4941
rect 6384 4901 6442 4907
rect 6572 4941 6630 4947
rect 6572 4907 6584 4941
rect 6618 4938 6630 4941
rect 7308 4941 7366 4947
rect 7308 4938 7320 4941
rect 6618 4910 7320 4938
rect 6618 4907 6630 4910
rect 6572 4901 6630 4907
rect 7308 4907 7320 4910
rect 7354 4907 7366 4941
rect 8412 4941 8470 4947
rect 7308 4901 7366 4907
rect 5736 4867 5798 4872
rect 5737 4864 5798 4867
rect 5576 4856 5629 4863
rect 7850 4860 7856 4912
rect 7908 4860 7914 4912
rect 7850 4852 7914 4860
rect 7972 4904 8025 4911
rect 8412 4907 8424 4941
rect 8458 4938 8470 4941
rect 8776 4941 8834 4947
rect 8776 4938 8788 4941
rect 8458 4910 8788 4938
rect 8458 4907 8470 4910
rect 7972 4852 7973 4904
rect 8135 4900 8196 4905
rect 8412 4901 8470 4907
rect 8776 4907 8788 4910
rect 8822 4907 8834 4941
rect 8776 4901 8834 4907
rect 8964 4941 9022 4947
rect 8964 4907 8976 4941
rect 9010 4938 9022 4941
rect 9700 4941 9758 4947
rect 9700 4938 9712 4941
rect 9010 4910 9712 4938
rect 9010 4907 9022 4910
rect 8964 4901 9022 4907
rect 9700 4907 9712 4910
rect 9746 4907 9758 4941
rect 10804 4941 10862 4947
rect 9700 4901 9758 4907
rect 10372 4920 10425 4927
rect 8132 4895 8196 4900
rect 8025 4861 8144 4895
rect 8178 4861 8196 4895
rect 8132 4856 8196 4861
rect 8135 4854 8196 4856
rect 10252 4889 10305 4896
rect 5460 4851 5524 4852
rect 5460 4846 5523 4851
rect 7972 4845 8025 4852
rect 10304 4837 10305 4889
rect 10372 4868 10373 4920
rect 10532 4911 10593 4920
rect 10425 4877 10544 4911
rect 10578 4877 10593 4911
rect 10804 4907 10816 4941
rect 10850 4938 10862 4941
rect 11168 4941 11226 4947
rect 11168 4938 11180 4941
rect 10850 4910 11180 4938
rect 10850 4907 10862 4910
rect 10804 4901 10862 4907
rect 11168 4907 11180 4910
rect 11214 4907 11226 4941
rect 11168 4901 11226 4907
rect 11356 4941 11414 4947
rect 11356 4907 11368 4941
rect 11402 4938 11414 4941
rect 12092 4941 12150 4947
rect 12092 4938 12104 4941
rect 11402 4910 12104 4938
rect 11402 4907 11414 4910
rect 11356 4901 11414 4907
rect 12092 4907 12104 4910
rect 12138 4907 12150 4941
rect 12092 4901 12150 4907
rect 12767 4920 12820 4927
rect 10532 4869 10593 4877
rect 12643 4890 12696 4897
rect 10372 4861 10425 4868
rect 10252 4830 10305 4837
rect 12695 4838 12696 4890
rect 12767 4868 12768 4920
rect 12926 4911 12987 4920
rect 12820 4877 12939 4911
rect 12973 4877 12987 4911
rect 12926 4869 12987 4877
rect 13068 4908 13332 4988
rect 12767 4861 12820 4868
rect 12643 4831 12696 4838
rect 408 4795 13027 4802
rect 13068 4795 13146 4908
rect 408 4771 13146 4795
rect 408 4737 1063 4771
rect 1097 4737 1155 4771
rect 1189 4737 1247 4771
rect 1281 4737 1339 4771
rect 1373 4737 1431 4771
rect 1465 4737 1523 4771
rect 1557 4737 1615 4771
rect 1649 4737 1707 4771
rect 1741 4737 1799 4771
rect 1833 4737 1891 4771
rect 1925 4737 1983 4771
rect 2017 4737 2075 4771
rect 2109 4737 2167 4771
rect 2201 4737 2259 4771
rect 2293 4737 2351 4771
rect 2385 4737 2443 4771
rect 2477 4737 2535 4771
rect 2569 4737 2627 4771
rect 2661 4737 2719 4771
rect 2753 4737 2811 4771
rect 2845 4737 2903 4771
rect 2937 4737 2995 4771
rect 3029 4737 3087 4771
rect 3121 4737 3179 4771
rect 3213 4737 3271 4771
rect 3305 4737 3363 4771
rect 3397 4737 3455 4771
rect 3489 4737 3547 4771
rect 3581 4737 3639 4771
rect 3673 4737 3731 4771
rect 3765 4737 3823 4771
rect 3857 4737 3915 4771
rect 3949 4737 4007 4771
rect 4041 4737 4099 4771
rect 4133 4737 4191 4771
rect 4225 4737 4283 4771
rect 4317 4737 4375 4771
rect 4409 4737 4467 4771
rect 4501 4737 4559 4771
rect 4593 4737 4651 4771
rect 4685 4737 4743 4771
rect 4777 4737 4835 4771
rect 4869 4737 4927 4771
rect 4961 4737 5019 4771
rect 5053 4737 5111 4771
rect 5145 4737 5203 4771
rect 5237 4737 5295 4771
rect 5329 4737 5387 4771
rect 5421 4737 5479 4771
rect 5513 4737 5571 4771
rect 5605 4737 5663 4771
rect 5697 4737 5755 4771
rect 5789 4737 5847 4771
rect 5881 4737 5939 4771
rect 5973 4737 6031 4771
rect 6065 4737 6123 4771
rect 6157 4737 6215 4771
rect 6249 4737 6307 4771
rect 6341 4737 6399 4771
rect 6433 4737 6491 4771
rect 6525 4737 6583 4771
rect 6617 4737 6675 4771
rect 6709 4737 6767 4771
rect 6801 4737 6859 4771
rect 6893 4737 6951 4771
rect 6985 4737 7043 4771
rect 7077 4737 7135 4771
rect 7169 4737 7227 4771
rect 7261 4737 7319 4771
rect 7353 4737 7411 4771
rect 7445 4737 7503 4771
rect 7537 4737 7595 4771
rect 7629 4737 7687 4771
rect 7721 4737 7779 4771
rect 7813 4737 7871 4771
rect 7905 4737 7963 4771
rect 7997 4737 8055 4771
rect 8089 4737 8147 4771
rect 8181 4737 8239 4771
rect 8273 4737 8331 4771
rect 8365 4737 8423 4771
rect 8457 4737 8515 4771
rect 8549 4737 8607 4771
rect 8641 4737 8699 4771
rect 8733 4737 8791 4771
rect 8825 4737 8883 4771
rect 8917 4737 8975 4771
rect 9009 4737 9067 4771
rect 9101 4737 9159 4771
rect 9193 4737 9251 4771
rect 9285 4737 9343 4771
rect 9377 4737 9435 4771
rect 9469 4737 9527 4771
rect 9561 4737 9619 4771
rect 9653 4737 9711 4771
rect 9745 4737 9803 4771
rect 9837 4737 9895 4771
rect 9929 4737 9987 4771
rect 10021 4737 10079 4771
rect 10113 4737 10171 4771
rect 10205 4737 10263 4771
rect 10297 4737 10355 4771
rect 10389 4737 10447 4771
rect 10481 4737 10539 4771
rect 10573 4737 10631 4771
rect 10665 4737 10723 4771
rect 10757 4737 10815 4771
rect 10849 4737 10907 4771
rect 10941 4737 10999 4771
rect 11033 4737 11091 4771
rect 11125 4737 11183 4771
rect 11217 4737 11275 4771
rect 11309 4737 11367 4771
rect 11401 4737 11459 4771
rect 11493 4737 11551 4771
rect 11585 4737 11643 4771
rect 11677 4737 11735 4771
rect 11769 4737 11827 4771
rect 11861 4737 11919 4771
rect 11953 4737 12011 4771
rect 12045 4737 12103 4771
rect 12137 4737 12195 4771
rect 12229 4737 12287 4771
rect 12321 4737 12379 4771
rect 12413 4737 12471 4771
rect 12505 4737 12563 4771
rect 12597 4737 12655 4771
rect 12689 4737 12747 4771
rect 12781 4737 12839 4771
rect 12873 4737 12931 4771
rect 12965 4762 13146 4771
rect 13296 4762 13332 4908
rect 12965 4737 13332 4762
rect 408 4719 13332 4737
rect 408 4706 13027 4719
rect 408 4650 13027 4657
rect 290 4626 13027 4650
rect 290 4592 623 4626
rect 657 4592 715 4626
rect 749 4592 807 4626
rect 841 4592 899 4626
rect 933 4592 991 4626
rect 1025 4592 1083 4626
rect 1117 4592 1175 4626
rect 1209 4592 1267 4626
rect 1301 4592 1359 4626
rect 1393 4592 1431 4626
rect 1465 4592 1523 4626
rect 1557 4592 1615 4626
rect 1649 4592 1707 4626
rect 1741 4592 1799 4626
rect 1833 4592 1891 4626
rect 1925 4592 1983 4626
rect 2017 4592 2075 4626
rect 2109 4592 2167 4626
rect 2201 4592 2259 4626
rect 2293 4592 2351 4626
rect 2385 4592 2443 4626
rect 2477 4592 2535 4626
rect 2569 4592 2627 4626
rect 2661 4592 2719 4626
rect 2753 4592 2811 4626
rect 2845 4592 2903 4626
rect 2937 4592 2995 4626
rect 3029 4592 3087 4626
rect 3121 4592 3179 4626
rect 3213 4592 3271 4626
rect 3305 4592 3363 4626
rect 3397 4592 3455 4626
rect 3489 4592 3547 4626
rect 3581 4592 3639 4626
rect 3673 4592 3731 4626
rect 3765 4592 3823 4626
rect 3857 4592 3915 4626
rect 3949 4592 4007 4626
rect 4041 4592 4099 4626
rect 4133 4592 4191 4626
rect 4225 4592 4283 4626
rect 4317 4592 4375 4626
rect 4409 4592 4467 4626
rect 4501 4592 4559 4626
rect 4593 4592 4651 4626
rect 4685 4592 4743 4626
rect 4777 4592 4835 4626
rect 4869 4592 4927 4626
rect 4961 4592 5019 4626
rect 5053 4592 5111 4626
rect 5145 4592 5203 4626
rect 5237 4592 5295 4626
rect 5329 4592 5387 4626
rect 5421 4592 5479 4626
rect 5513 4592 5571 4626
rect 5605 4592 5663 4626
rect 5697 4592 5755 4626
rect 5789 4592 5847 4626
rect 5881 4592 5939 4626
rect 5973 4592 6031 4626
rect 6065 4592 6123 4626
rect 6157 4592 6215 4626
rect 6249 4592 6307 4626
rect 6341 4592 6399 4626
rect 6433 4592 6491 4626
rect 6525 4592 6583 4626
rect 6617 4592 6675 4626
rect 6709 4592 6767 4626
rect 6801 4592 6859 4626
rect 6893 4592 6951 4626
rect 6985 4592 7043 4626
rect 7077 4592 7135 4626
rect 7169 4592 7227 4626
rect 7261 4592 7319 4626
rect 7353 4592 7411 4626
rect 7445 4592 7503 4626
rect 7537 4592 7595 4626
rect 7629 4592 7687 4626
rect 7721 4592 7779 4626
rect 7813 4592 7871 4626
rect 7905 4592 7963 4626
rect 7997 4592 8055 4626
rect 8089 4592 8147 4626
rect 8181 4592 8239 4626
rect 8273 4592 8331 4626
rect 8365 4592 8423 4626
rect 8457 4592 8515 4626
rect 8549 4592 8607 4626
rect 8641 4592 8699 4626
rect 8733 4592 8791 4626
rect 8825 4592 8883 4626
rect 8917 4592 8975 4626
rect 9009 4592 9067 4626
rect 9101 4592 9159 4626
rect 9193 4592 9251 4626
rect 9285 4592 9343 4626
rect 9377 4592 9435 4626
rect 9469 4592 9527 4626
rect 9561 4592 9619 4626
rect 9653 4592 9711 4626
rect 9745 4592 9803 4626
rect 9837 4592 9895 4626
rect 9929 4592 9987 4626
rect 10021 4592 10079 4626
rect 10113 4592 10171 4626
rect 10205 4592 10263 4626
rect 10297 4592 10355 4626
rect 10389 4592 10447 4626
rect 10481 4592 10539 4626
rect 10573 4592 10631 4626
rect 10665 4592 10723 4626
rect 10757 4592 10815 4626
rect 10849 4592 10907 4626
rect 10941 4592 10999 4626
rect 11033 4592 11091 4626
rect 11125 4592 11183 4626
rect 11217 4592 11275 4626
rect 11309 4592 11367 4626
rect 11401 4592 11459 4626
rect 11493 4592 11551 4626
rect 11585 4592 11643 4626
rect 11677 4592 11735 4626
rect 11769 4592 11827 4626
rect 11861 4592 11919 4626
rect 11953 4592 12011 4626
rect 12045 4592 12103 4626
rect 12137 4592 12195 4626
rect 12229 4592 12287 4626
rect 12321 4592 12379 4626
rect 12413 4592 12471 4626
rect 12505 4592 12563 4626
rect 12597 4592 12655 4626
rect 12689 4592 12747 4626
rect 12781 4592 12839 4626
rect 12873 4592 12931 4626
rect 12965 4592 13027 4626
rect 290 4586 13027 4592
rect 290 4440 324 4586
rect 474 4561 13027 4586
rect 474 4440 520 4561
rect 290 4378 520 4440
rect 2527 4498 2580 4505
rect 2527 4446 2528 4498
rect 3436 4480 3442 4532
rect 3494 4480 3500 4532
rect 5833 4514 5899 4515
rect 5833 4462 5840 4514
rect 5892 4499 5899 4514
rect 8224 4514 8290 4515
rect 5892 4462 5952 4499
rect 8224 4462 8231 4514
rect 8283 4499 8290 4514
rect 10618 4505 10671 4511
rect 8283 4462 8344 4499
rect 2527 4439 2580 4446
rect 4546 4456 4604 4462
rect 4546 4422 4558 4456
rect 4592 4453 4604 4456
rect 5282 4456 5340 4462
rect 5282 4453 5294 4456
rect 4592 4425 5294 4453
rect 4592 4422 4604 4425
rect 4546 4416 4604 4422
rect 5282 4422 5294 4425
rect 5328 4453 5340 4456
rect 5650 4456 5708 4462
rect 5650 4453 5662 4456
rect 5328 4425 5662 4453
rect 5328 4422 5340 4425
rect 5282 4416 5340 4422
rect 5650 4422 5662 4425
rect 5696 4422 5708 4456
rect 5650 4416 5708 4422
rect 5833 4397 5886 4404
rect 5833 4396 5834 4397
rect 3994 4388 4052 4394
rect 3994 4354 4006 4388
rect 4040 4385 4052 4388
rect 4638 4388 4696 4394
rect 4638 4385 4650 4388
rect 4040 4357 4650 4385
rect 4040 4354 4052 4357
rect 3994 4348 4052 4354
rect 4638 4354 4650 4357
rect 4684 4354 4696 4388
rect 4638 4348 4696 4354
rect 5417 4386 5476 4392
rect 5828 4386 5834 4396
rect 5417 4352 5430 4386
rect 5464 4358 5834 4386
rect 5464 4352 5476 4358
rect 5417 4345 5476 4352
rect 5828 4349 5834 4358
rect 5833 4345 5834 4349
rect 5886 4349 5887 4396
rect 3888 4332 3941 4339
rect 5833 4338 5886 4345
rect 617 4328 682 4329
rect 470 4319 504 4322
rect 611 4319 682 4328
rect 468 4318 682 4319
rect 468 4291 625 4318
rect 470 4288 504 4291
rect 611 4284 625 4291
rect 659 4284 682 4318
rect 611 4278 682 4284
rect 617 4277 682 4278
rect 3940 4280 3941 4332
rect 4546 4320 4604 4326
rect 4546 4286 4558 4320
rect 4592 4317 4604 4320
rect 4592 4289 5233 4317
rect 4592 4286 4604 4289
rect 4546 4280 4604 4286
rect 3888 4273 3941 4280
rect 5194 4258 5233 4289
rect 5736 4307 5786 4308
rect 5736 4305 5796 4307
rect 5915 4305 5952 4462
rect 6938 4456 6996 4462
rect 6938 4422 6950 4456
rect 6984 4453 6996 4456
rect 7674 4456 7732 4462
rect 7674 4453 7686 4456
rect 6984 4425 7686 4453
rect 6984 4422 6996 4425
rect 6938 4416 6996 4422
rect 7674 4422 7686 4425
rect 7720 4453 7732 4456
rect 8042 4456 8100 4462
rect 8042 4453 8054 4456
rect 7720 4425 8054 4453
rect 7720 4422 7732 4425
rect 7674 4416 7732 4422
rect 8042 4422 8054 4425
rect 8088 4422 8100 4456
rect 8042 4416 8100 4422
rect 8221 4396 8274 4402
rect 8220 4395 8279 4396
rect 6386 4388 6444 4394
rect 6386 4354 6398 4388
rect 6432 4385 6444 4388
rect 7030 4388 7088 4394
rect 7030 4385 7042 4388
rect 6432 4357 7042 4385
rect 6432 4354 6444 4357
rect 6386 4348 6444 4354
rect 7030 4354 7042 4357
rect 7076 4354 7088 4388
rect 7030 4348 7088 4354
rect 7809 4386 7868 4392
rect 8220 4386 8222 4395
rect 7809 4352 7822 4386
rect 7856 4358 8222 4386
rect 7856 4352 7868 4358
rect 7809 4345 7868 4352
rect 8220 4349 8222 4358
rect 8221 4343 8222 4349
rect 8274 4349 8279 4395
rect 5736 4301 5952 4305
rect 5736 4267 5750 4301
rect 5784 4268 5952 4301
rect 6283 4333 6336 4340
rect 8221 4336 8274 4343
rect 6335 4281 6336 4333
rect 6283 4274 6336 4281
rect 6938 4320 6996 4326
rect 6938 4286 6950 4320
rect 6984 4317 6996 4320
rect 6984 4289 7625 4317
rect 6984 4286 6996 4289
rect 6938 4280 6996 4286
rect 5784 4267 5796 4268
rect 5736 4260 5796 4267
rect 7586 4258 7625 4289
rect 8133 4305 8190 4308
rect 8307 4305 8344 4462
rect 9330 4456 9388 4462
rect 9330 4422 9342 4456
rect 9376 4453 9388 4456
rect 10066 4456 10124 4462
rect 10066 4453 10078 4456
rect 9376 4425 10078 4453
rect 9376 4422 9388 4425
rect 9330 4416 9388 4422
rect 10066 4422 10078 4425
rect 10112 4453 10124 4456
rect 10434 4456 10492 4462
rect 10434 4453 10446 4456
rect 10112 4425 10446 4453
rect 10112 4422 10124 4425
rect 10066 4416 10124 4422
rect 10434 4422 10446 4425
rect 10480 4422 10492 4456
rect 10618 4453 10619 4505
rect 10671 4462 10736 4499
rect 10618 4445 10671 4453
rect 10434 4416 10492 4422
rect 10613 4397 10666 4403
rect 10612 4396 10671 4397
rect 8778 4388 8836 4394
rect 8778 4354 8790 4388
rect 8824 4385 8836 4388
rect 9422 4388 9480 4394
rect 9422 4385 9434 4388
rect 8824 4357 9434 4385
rect 8824 4354 8836 4357
rect 8778 4348 8836 4354
rect 9422 4354 9434 4357
rect 9468 4354 9480 4388
rect 9422 4348 9480 4354
rect 10201 4387 10260 4393
rect 10612 4387 10614 4396
rect 10201 4353 10214 4387
rect 10248 4359 10614 4387
rect 10248 4353 10260 4359
rect 10201 4346 10260 4353
rect 10612 4350 10614 4359
rect 10613 4344 10614 4350
rect 10666 4350 10671 4396
rect 8133 4302 8344 4305
rect 8133 4268 8147 4302
rect 8181 4268 8344 4302
rect 8673 4334 8726 4341
rect 10613 4337 10666 4344
rect 8725 4282 8726 4334
rect 8673 4275 8726 4282
rect 9330 4320 9388 4326
rect 9330 4286 9342 4320
rect 9376 4317 9388 4320
rect 9376 4289 10017 4317
rect 9376 4286 9388 4289
rect 9330 4280 9388 4286
rect 4270 4252 4328 4258
rect 4270 4218 4282 4252
rect 4316 4249 4328 4252
rect 5006 4252 5064 4258
rect 5006 4249 5018 4252
rect 4316 4221 5018 4249
rect 4316 4218 4328 4221
rect 4270 4212 4328 4218
rect 5006 4218 5018 4221
rect 5052 4218 5064 4252
rect 5006 4212 5064 4218
rect 5194 4252 5252 4258
rect 5194 4218 5206 4252
rect 5240 4249 5252 4252
rect 5558 4252 5616 4258
rect 5558 4249 5570 4252
rect 5240 4221 5570 4249
rect 5240 4218 5252 4221
rect 5194 4212 5252 4218
rect 5558 4218 5570 4221
rect 5604 4218 5616 4252
rect 6662 4252 6720 4258
rect 5976 4229 6029 4236
rect 5558 4212 5616 4218
rect 5831 4222 5893 4228
rect 3349 4194 3415 4195
rect 3349 4142 3356 4194
rect 3408 4142 3415 4194
rect 5831 4188 5845 4222
rect 5879 4221 5893 4222
rect 5879 4188 5976 4221
rect 5831 4187 5976 4188
rect 5831 4182 5893 4187
rect 6028 4177 6029 4229
rect 6662 4218 6674 4252
rect 6708 4249 6720 4252
rect 7398 4252 7456 4258
rect 7398 4249 7410 4252
rect 6708 4221 7410 4249
rect 6708 4218 6720 4221
rect 6662 4212 6720 4218
rect 7398 4218 7410 4221
rect 7444 4218 7456 4252
rect 7398 4212 7456 4218
rect 7586 4252 7644 4258
rect 7586 4218 7598 4252
rect 7632 4249 7644 4252
rect 7950 4252 8008 4258
rect 8133 4255 8190 4268
rect 9978 4258 10017 4289
rect 10525 4305 10579 4309
rect 10699 4305 10736 4462
rect 11722 4456 11780 4462
rect 11722 4422 11734 4456
rect 11768 4453 11780 4456
rect 12458 4456 12516 4462
rect 12458 4453 12470 4456
rect 11768 4425 12470 4453
rect 11768 4422 11780 4425
rect 11722 4416 11780 4422
rect 12458 4422 12470 4425
rect 12504 4453 12516 4456
rect 12826 4456 12884 4462
rect 12826 4453 12838 4456
rect 12504 4425 12838 4453
rect 12504 4422 12516 4425
rect 12458 4416 12516 4422
rect 12826 4422 12838 4425
rect 12872 4422 12884 4456
rect 12826 4416 12884 4422
rect 11170 4388 11228 4394
rect 11170 4354 11182 4388
rect 11216 4385 11228 4388
rect 11814 4388 11872 4394
rect 11814 4385 11826 4388
rect 11216 4357 11826 4385
rect 11216 4354 11228 4357
rect 11170 4348 11228 4354
rect 11814 4354 11826 4357
rect 11860 4354 11872 4388
rect 11814 4348 11872 4354
rect 12558 4388 12629 4396
rect 10525 4302 10736 4305
rect 10525 4268 10538 4302
rect 10572 4268 10736 4302
rect 11067 4331 11120 4338
rect 12558 4336 12566 4388
rect 12618 4336 12629 4388
rect 11119 4279 11120 4331
rect 12914 4331 12920 4383
rect 12972 4331 12978 4383
rect 12914 4330 12978 4331
rect 11722 4320 11780 4326
rect 11722 4286 11734 4320
rect 11768 4317 11780 4320
rect 11768 4289 12409 4317
rect 11768 4286 11780 4289
rect 11722 4280 11780 4286
rect 11067 4272 11120 4279
rect 7950 4249 7962 4252
rect 7632 4221 7962 4249
rect 7632 4218 7644 4221
rect 7586 4212 7644 4218
rect 7950 4218 7962 4221
rect 7996 4218 8008 4252
rect 9054 4252 9112 4258
rect 7950 4212 8008 4218
rect 8227 4209 8294 4219
rect 8398 4218 8451 4225
rect 5976 4170 6029 4177
rect 6118 4183 6171 4195
rect 6118 4149 6131 4183
rect 6165 4174 6171 4183
rect 6567 4193 6633 4194
rect 6567 4174 6574 4193
rect 6165 4149 6574 4174
rect 6118 4146 6574 4149
rect 6118 4143 6171 4146
rect 6567 4141 6574 4146
rect 6626 4174 6633 4193
rect 8227 4175 8245 4209
rect 8279 4175 8398 4209
rect 6626 4146 6832 4174
rect 8227 4165 8294 4175
rect 8450 4166 8451 4218
rect 9054 4218 9066 4252
rect 9100 4249 9112 4252
rect 9790 4252 9848 4258
rect 9790 4249 9802 4252
rect 9100 4221 9802 4249
rect 9100 4218 9112 4221
rect 9054 4212 9112 4218
rect 9790 4218 9802 4221
rect 9836 4218 9848 4252
rect 9790 4212 9848 4218
rect 9978 4252 10036 4258
rect 9978 4218 9990 4252
rect 10024 4249 10036 4252
rect 10342 4252 10400 4258
rect 10525 4257 10579 4268
rect 12370 4258 12409 4289
rect 10342 4249 10354 4252
rect 10024 4221 10354 4249
rect 10024 4218 10036 4221
rect 9978 4212 10036 4218
rect 10342 4218 10354 4221
rect 10388 4218 10400 4252
rect 11446 4252 11504 4258
rect 10342 4212 10400 4218
rect 10615 4217 10682 4227
rect 10786 4226 10839 4233
rect 8959 4194 9025 4195
rect 8398 4159 8451 4166
rect 8507 4182 8565 4189
rect 8507 4148 8519 4182
rect 8553 4173 8565 4182
rect 8959 4173 8966 4194
rect 8553 4148 8966 4173
rect 6626 4141 6633 4146
rect 8507 4145 8966 4148
rect 8507 4142 8565 4145
rect 8959 4142 8966 4145
rect 9018 4173 9025 4194
rect 10615 4183 10633 4217
rect 10667 4183 10786 4217
rect 10615 4173 10682 4183
rect 10838 4174 10839 4226
rect 11446 4218 11458 4252
rect 11492 4249 11504 4252
rect 12182 4252 12240 4258
rect 12182 4249 12194 4252
rect 11492 4221 12194 4249
rect 11492 4218 11504 4221
rect 11446 4212 11504 4218
rect 12182 4218 12194 4221
rect 12228 4218 12240 4252
rect 12182 4212 12240 4218
rect 12370 4252 12428 4258
rect 12370 4218 12382 4252
rect 12416 4249 12428 4252
rect 12734 4252 12792 4258
rect 12734 4249 12746 4252
rect 12416 4221 12746 4249
rect 12416 4218 12428 4221
rect 12370 4212 12428 4218
rect 12734 4218 12746 4221
rect 12780 4218 12792 4252
rect 12734 4212 12792 4218
rect 11348 4195 11414 4196
rect 9018 4145 9225 4173
rect 10786 4167 10839 4174
rect 10898 4188 10959 4194
rect 10898 4154 10913 4188
rect 10947 4174 10959 4188
rect 11348 4174 11355 4195
rect 10947 4154 11355 4174
rect 10898 4146 11355 4154
rect 9018 4142 9025 4145
rect 10898 4142 10959 4146
rect 11348 4143 11355 4146
rect 11407 4174 11414 4195
rect 13080 4174 13332 4256
rect 11407 4146 11617 4174
rect 11407 4143 11414 4146
rect 13080 4113 13162 4174
rect 469 4082 13162 4113
rect 469 4048 623 4082
rect 657 4048 715 4082
rect 749 4048 807 4082
rect 841 4048 899 4082
rect 933 4048 991 4082
rect 1025 4048 1083 4082
rect 1117 4048 1175 4082
rect 1209 4048 1267 4082
rect 1301 4048 1359 4082
rect 1393 4048 1431 4082
rect 1465 4048 1523 4082
rect 1557 4048 1615 4082
rect 1649 4048 1707 4082
rect 1741 4048 1799 4082
rect 1833 4048 1891 4082
rect 1925 4048 1983 4082
rect 2017 4048 2075 4082
rect 2109 4048 2167 4082
rect 2201 4048 2259 4082
rect 2293 4048 2351 4082
rect 2385 4048 2443 4082
rect 2477 4048 2535 4082
rect 2569 4048 2627 4082
rect 2661 4048 2719 4082
rect 2753 4048 2811 4082
rect 2845 4048 2903 4082
rect 2937 4048 2995 4082
rect 3029 4048 3087 4082
rect 3121 4048 3179 4082
rect 3213 4048 3271 4082
rect 3305 4048 3363 4082
rect 3397 4048 3455 4082
rect 3489 4048 3547 4082
rect 3581 4048 3639 4082
rect 3673 4048 3731 4082
rect 3765 4048 3823 4082
rect 3857 4048 3915 4082
rect 3949 4048 4007 4082
rect 4041 4048 4099 4082
rect 4133 4048 4191 4082
rect 4225 4048 4283 4082
rect 4317 4048 4375 4082
rect 4409 4048 4467 4082
rect 4501 4048 4559 4082
rect 4593 4048 4651 4082
rect 4685 4048 4743 4082
rect 4777 4048 4835 4082
rect 4869 4048 4927 4082
rect 4961 4048 5019 4082
rect 5053 4048 5111 4082
rect 5145 4048 5203 4082
rect 5237 4048 5295 4082
rect 5329 4048 5387 4082
rect 5421 4048 5479 4082
rect 5513 4048 5571 4082
rect 5605 4048 5663 4082
rect 5697 4048 5755 4082
rect 5789 4048 5847 4082
rect 5881 4048 5939 4082
rect 5973 4048 6031 4082
rect 6065 4048 6123 4082
rect 6157 4048 6215 4082
rect 6249 4048 6307 4082
rect 6341 4048 6399 4082
rect 6433 4048 6491 4082
rect 6525 4048 6583 4082
rect 6617 4048 6675 4082
rect 6709 4048 6767 4082
rect 6801 4048 6859 4082
rect 6893 4048 6951 4082
rect 6985 4048 7043 4082
rect 7077 4048 7135 4082
rect 7169 4048 7227 4082
rect 7261 4048 7319 4082
rect 7353 4048 7411 4082
rect 7445 4048 7503 4082
rect 7537 4048 7595 4082
rect 7629 4048 7687 4082
rect 7721 4048 7779 4082
rect 7813 4048 7871 4082
rect 7905 4048 7963 4082
rect 7997 4048 8055 4082
rect 8089 4048 8147 4082
rect 8181 4048 8239 4082
rect 8273 4048 8331 4082
rect 8365 4048 8423 4082
rect 8457 4048 8515 4082
rect 8549 4048 8607 4082
rect 8641 4048 8699 4082
rect 8733 4048 8791 4082
rect 8825 4048 8883 4082
rect 8917 4048 8975 4082
rect 9009 4048 9067 4082
rect 9101 4048 9159 4082
rect 9193 4048 9251 4082
rect 9285 4048 9343 4082
rect 9377 4048 9435 4082
rect 9469 4048 9527 4082
rect 9561 4048 9619 4082
rect 9653 4048 9711 4082
rect 9745 4048 9803 4082
rect 9837 4048 9895 4082
rect 9929 4048 9987 4082
rect 10021 4048 10079 4082
rect 10113 4048 10171 4082
rect 10205 4048 10263 4082
rect 10297 4048 10355 4082
rect 10389 4048 10447 4082
rect 10481 4048 10539 4082
rect 10573 4048 10631 4082
rect 10665 4048 10723 4082
rect 10757 4048 10815 4082
rect 10849 4048 10907 4082
rect 10941 4048 10999 4082
rect 11033 4048 11091 4082
rect 11125 4048 11183 4082
rect 11217 4048 11275 4082
rect 11309 4048 11367 4082
rect 11401 4048 11459 4082
rect 11493 4048 11551 4082
rect 11585 4048 11643 4082
rect 11677 4048 11735 4082
rect 11769 4048 11827 4082
rect 11861 4048 11919 4082
rect 11953 4048 12011 4082
rect 12045 4048 12103 4082
rect 12137 4048 12195 4082
rect 12229 4048 12287 4082
rect 12321 4048 12379 4082
rect 12413 4048 12471 4082
rect 12505 4048 12563 4082
rect 12597 4048 12655 4082
rect 12689 4048 12747 4082
rect 12781 4048 12839 4082
rect 12873 4048 12931 4082
rect 12965 4048 13162 4082
rect 469 4028 13162 4048
rect 13312 4028 13332 4174
rect 469 4017 13332 4028
rect 3349 3952 3415 3953
rect 1489 3941 1496 3952
rect 1484 3912 1496 3941
rect 1489 3900 1496 3912
rect 1548 3941 1555 3952
rect 3349 3941 3356 3952
rect 1548 3912 3356 3941
rect 1548 3900 1555 3912
rect 3349 3900 3356 3912
rect 3408 3941 3415 3952
rect 3881 3952 3947 3953
rect 3881 3941 3888 3952
rect 3408 3912 3888 3941
rect 3408 3900 3415 3912
rect 3881 3900 3888 3912
rect 3940 3941 3947 3952
rect 5285 3952 5351 3953
rect 5285 3941 5292 3952
rect 3940 3913 5292 3941
rect 3940 3900 3947 3913
rect 5285 3900 5292 3913
rect 5344 3941 5351 3952
rect 6270 3952 6336 3953
rect 6270 3941 6277 3952
rect 5344 3913 6277 3941
rect 5344 3900 5351 3913
rect 6270 3900 6277 3913
rect 6329 3941 6336 3952
rect 7677 3952 7743 3953
rect 7677 3941 7684 3952
rect 6329 3913 7684 3941
rect 6329 3900 6336 3913
rect 7677 3900 7684 3913
rect 7736 3941 7743 3952
rect 8660 3952 8726 3953
rect 8660 3941 8667 3952
rect 7736 3913 8667 3941
rect 7736 3900 7743 3913
rect 8660 3900 8667 3913
rect 8719 3941 8726 3952
rect 10074 3952 10140 3953
rect 10074 3941 10081 3952
rect 8719 3913 10081 3941
rect 8719 3900 8726 3913
rect 10074 3900 10081 3913
rect 10133 3941 10140 3952
rect 11050 3952 11116 3953
rect 11050 3941 11057 3952
rect 10133 3913 11057 3941
rect 10133 3900 10140 3913
rect 11050 3900 11057 3913
rect 11109 3941 11116 3952
rect 12462 3952 12528 3953
rect 12462 3941 12469 3952
rect 11109 3913 12469 3941
rect 11109 3900 11116 3913
rect 12462 3900 12469 3913
rect 12521 3941 12528 3952
rect 12521 3913 12941 3941
rect 12521 3900 12528 3913
rect 13074 3840 13332 4017
rect 489 3812 13332 3840
rect 486 3779 13105 3784
rect 290 3753 13105 3779
rect 290 3752 3197 3753
rect 290 3740 655 3752
rect 290 3594 360 3740
rect 510 3718 655 3740
rect 689 3744 747 3752
rect 781 3744 839 3752
rect 689 3718 712 3744
rect 873 3718 931 3752
rect 965 3718 1023 3752
rect 1057 3718 1115 3752
rect 1149 3744 1207 3752
rect 1241 3744 1299 3752
rect 1149 3718 1158 3744
rect 1333 3718 1391 3752
rect 1425 3748 3197 3752
rect 1425 3718 1724 3748
rect 510 3598 712 3718
rect 862 3598 1158 3718
rect 1308 3602 1724 3718
rect 1874 3602 2390 3748
rect 2540 3732 3197 3748
rect 2540 3602 2772 3732
rect 1308 3598 2772 3602
rect 510 3594 2772 3598
rect 290 3586 2772 3594
rect 2922 3719 3197 3732
rect 3231 3719 3289 3753
rect 3323 3719 3381 3753
rect 3415 3719 3454 3753
rect 3488 3719 3546 3753
rect 3580 3719 3638 3753
rect 3672 3719 3730 3753
rect 3764 3719 3822 3753
rect 3856 3719 3914 3753
rect 3948 3719 4006 3753
rect 4040 3719 4098 3753
rect 4132 3719 4190 3753
rect 4224 3719 4282 3753
rect 4316 3719 4374 3753
rect 4408 3719 4466 3753
rect 4500 3719 4558 3753
rect 4592 3719 4650 3753
rect 4684 3719 4742 3753
rect 4776 3719 4834 3753
rect 4868 3719 4926 3753
rect 4960 3719 5018 3753
rect 5052 3719 5110 3753
rect 5144 3719 5202 3753
rect 5236 3719 5294 3753
rect 5328 3719 5386 3753
rect 5420 3719 5478 3753
rect 5512 3719 5570 3753
rect 5604 3719 5662 3753
rect 5696 3719 5754 3753
rect 5788 3719 5846 3753
rect 5880 3719 5938 3753
rect 5972 3719 6030 3753
rect 6064 3719 6122 3753
rect 6156 3719 6214 3753
rect 6248 3719 6306 3753
rect 6340 3719 6398 3753
rect 6432 3719 6490 3753
rect 6524 3719 6582 3753
rect 6616 3719 6674 3753
rect 6708 3719 6766 3753
rect 6800 3719 6858 3753
rect 6892 3719 6950 3753
rect 6984 3719 7042 3753
rect 7076 3719 7134 3753
rect 7168 3719 7226 3753
rect 7260 3719 7318 3753
rect 7352 3719 7410 3753
rect 7444 3719 7502 3753
rect 7536 3719 7594 3753
rect 7628 3719 7686 3753
rect 7720 3719 7778 3753
rect 7812 3719 7870 3753
rect 7904 3719 7962 3753
rect 7996 3719 8054 3753
rect 8088 3719 8146 3753
rect 8180 3719 8238 3753
rect 8272 3719 8330 3753
rect 8364 3719 8422 3753
rect 8456 3719 8514 3753
rect 8548 3719 8606 3753
rect 8640 3719 8698 3753
rect 8732 3719 8790 3753
rect 8824 3719 8882 3753
rect 8916 3719 8974 3753
rect 9008 3719 9066 3753
rect 9100 3719 9158 3753
rect 9192 3719 9250 3753
rect 9284 3719 9342 3753
rect 9376 3719 9434 3753
rect 9468 3719 9526 3753
rect 9560 3719 9618 3753
rect 9652 3719 9710 3753
rect 9744 3719 9802 3753
rect 9836 3719 9894 3753
rect 9928 3719 9986 3753
rect 10020 3719 10078 3753
rect 10112 3719 10170 3753
rect 10204 3719 10262 3753
rect 10296 3719 10354 3753
rect 10388 3719 10446 3753
rect 10480 3719 10538 3753
rect 10572 3719 10630 3753
rect 10664 3719 10722 3753
rect 10756 3719 10814 3753
rect 10848 3719 10906 3753
rect 10940 3719 10998 3753
rect 11032 3719 11090 3753
rect 11124 3719 11182 3753
rect 11216 3719 11274 3753
rect 11308 3719 11366 3753
rect 11400 3719 11458 3753
rect 11492 3719 11550 3753
rect 11584 3719 11642 3753
rect 11676 3719 11734 3753
rect 11768 3719 11826 3753
rect 11860 3719 11918 3753
rect 11952 3719 12010 3753
rect 12044 3719 12102 3753
rect 12136 3719 12194 3753
rect 12228 3719 12286 3753
rect 12320 3719 12378 3753
rect 12412 3719 12470 3753
rect 12504 3719 12562 3753
rect 12596 3719 12654 3753
rect 12688 3719 12746 3753
rect 12780 3719 12838 3753
rect 12872 3719 12930 3753
rect 12964 3719 13105 3753
rect 2922 3688 13105 3719
rect 2922 3586 3026 3688
rect 290 3554 3026 3586
rect 3535 3583 3593 3589
rect 3535 3549 3547 3583
rect 3581 3580 3593 3583
rect 3903 3583 3961 3589
rect 3903 3580 3915 3583
rect 3581 3552 3915 3580
rect 3581 3549 3593 3552
rect 3535 3543 3593 3549
rect 3903 3549 3915 3552
rect 3949 3580 3961 3583
rect 4639 3583 4697 3589
rect 4639 3580 4651 3583
rect 3949 3552 4651 3580
rect 3949 3549 3961 3552
rect 3903 3543 3961 3549
rect 4639 3549 4651 3552
rect 4685 3549 4697 3583
rect 4639 3543 4697 3549
rect 5927 3583 5985 3589
rect 5927 3549 5939 3583
rect 5973 3580 5985 3583
rect 6295 3583 6353 3589
rect 6295 3580 6307 3583
rect 5973 3552 6307 3580
rect 5973 3549 5985 3552
rect 5927 3543 5985 3549
rect 6295 3549 6307 3552
rect 6341 3580 6353 3583
rect 7031 3583 7089 3589
rect 7031 3580 7043 3583
rect 6341 3552 7043 3580
rect 6341 3549 6353 3552
rect 6295 3543 6353 3549
rect 7031 3549 7043 3552
rect 7077 3549 7089 3583
rect 7031 3543 7089 3549
rect 8319 3583 8377 3589
rect 8319 3549 8331 3583
rect 8365 3580 8377 3583
rect 8687 3583 8745 3589
rect 8687 3580 8699 3583
rect 8365 3552 8699 3580
rect 8365 3549 8377 3552
rect 8319 3543 8377 3549
rect 8687 3549 8699 3552
rect 8733 3580 8745 3583
rect 9423 3583 9481 3589
rect 9423 3580 9435 3583
rect 8733 3552 9435 3580
rect 8733 3549 8745 3552
rect 8687 3543 8745 3549
rect 9423 3549 9435 3552
rect 9469 3549 9481 3583
rect 9423 3543 9481 3549
rect 10711 3583 10769 3589
rect 10711 3549 10723 3583
rect 10757 3580 10769 3583
rect 11079 3583 11137 3589
rect 11079 3580 11091 3583
rect 10757 3552 11091 3580
rect 10757 3549 10769 3552
rect 10711 3543 10769 3549
rect 11079 3549 11091 3552
rect 11125 3580 11137 3583
rect 11815 3583 11873 3589
rect 11815 3580 11827 3583
rect 11125 3552 11827 3580
rect 11125 3549 11137 3552
rect 11079 3543 11137 3549
rect 11815 3549 11827 3552
rect 11861 3549 11873 3583
rect 11815 3543 11873 3549
rect 2614 3524 2681 3525
rect 468 3483 1632 3511
rect 468 3414 502 3483
rect 650 3397 656 3449
rect 708 3397 714 3449
rect 1257 3397 1263 3449
rect 1315 3397 1321 3449
rect 1598 3443 1632 3483
rect 2614 3472 2622 3524
rect 2674 3499 2681 3524
rect 3060 3523 3126 3524
rect 3060 3499 3067 3523
rect 2674 3472 3067 3499
rect 2622 3471 3067 3472
rect 3119 3471 3126 3523
rect 3333 3520 3394 3527
rect 3333 3486 3347 3520
rect 3381 3515 3394 3520
rect 4181 3515 4189 3524
rect 3381 3487 4189 3515
rect 3381 3486 3394 3487
rect 3333 3480 3394 3486
rect 4181 3472 4189 3487
rect 4241 3472 4248 3524
rect 4547 3515 4605 3521
rect 4547 3481 4559 3515
rect 4593 3512 4605 3515
rect 5191 3515 5249 3521
rect 5191 3512 5203 3515
rect 4593 3484 5203 3512
rect 4593 3481 4605 3484
rect 4547 3475 4605 3481
rect 5191 3481 5203 3484
rect 5237 3481 5249 3515
rect 5191 3475 5249 3481
rect 6939 3515 6997 3521
rect 6939 3481 6951 3515
rect 6985 3512 6997 3515
rect 7583 3515 7641 3521
rect 7583 3512 7595 3515
rect 6985 3484 7595 3512
rect 6985 3481 6997 3484
rect 6939 3475 6997 3481
rect 7583 3481 7595 3484
rect 7629 3481 7641 3515
rect 7583 3475 7641 3481
rect 9331 3515 9389 3521
rect 9331 3481 9343 3515
rect 9377 3512 9389 3515
rect 9975 3515 10033 3521
rect 9975 3512 9987 3515
rect 9377 3484 9987 3512
rect 9377 3481 9389 3484
rect 9331 3475 9389 3481
rect 9975 3481 9987 3484
rect 10021 3481 10033 3515
rect 9975 3475 10033 3481
rect 11723 3515 11781 3521
rect 11723 3481 11735 3515
rect 11769 3512 11781 3515
rect 12367 3515 12425 3521
rect 12367 3512 12379 3515
rect 11769 3484 12379 3512
rect 11769 3481 11781 3484
rect 11723 3475 11781 3481
rect 12367 3481 12379 3484
rect 12413 3481 12425 3515
rect 12367 3475 12425 3481
rect 7684 3463 7737 3470
rect 2012 3451 2078 3452
rect 2012 3443 2019 3451
rect 1598 3415 2019 3443
rect 2012 3399 2019 3415
rect 2071 3443 2078 3451
rect 3156 3446 3202 3458
rect 3156 3443 3162 3446
rect 2071 3415 3162 3443
rect 2071 3399 2078 3415
rect 3156 3412 3162 3415
rect 3196 3412 3202 3446
rect 3156 3400 3202 3412
rect 3446 3445 3495 3458
rect 3446 3411 3455 3445
rect 3489 3411 3495 3445
rect 3446 3404 3495 3411
rect 3541 3453 3837 3459
rect 5293 3453 5346 3460
rect 3541 3420 3784 3453
rect 3453 3240 3492 3404
rect 3541 3240 3580 3420
rect 3776 3419 3784 3420
rect 3818 3419 3837 3453
rect 4639 3447 4697 3453
rect 4639 3444 4651 3447
rect 3776 3407 3837 3419
rect 4010 3416 4651 3444
rect 4010 3385 4049 3416
rect 4639 3413 4651 3416
rect 4685 3413 4697 3447
rect 4639 3407 4697 3413
rect 5345 3401 5346 3453
rect 6184 3405 6191 3457
rect 6243 3405 6250 3457
rect 7031 3447 7089 3453
rect 7031 3444 7043 3447
rect 6402 3416 7043 3444
rect 5293 3394 5346 3401
rect 3627 3379 3685 3385
rect 3627 3345 3639 3379
rect 3673 3376 3685 3379
rect 3991 3379 4049 3385
rect 3991 3376 4003 3379
rect 3673 3348 4003 3376
rect 3673 3345 3685 3348
rect 3627 3339 3685 3345
rect 3991 3345 4003 3348
rect 4037 3345 4049 3379
rect 3991 3339 4049 3345
rect 4175 3387 4239 3388
rect 4175 3335 4181 3387
rect 4233 3376 4239 3387
rect 6402 3385 6441 3416
rect 7031 3413 7043 3416
rect 7077 3413 7089 3447
rect 7031 3407 7089 3413
rect 7736 3411 7737 3463
rect 10075 3459 10128 3466
rect 7684 3404 7737 3411
rect 8571 3405 8578 3457
rect 8630 3405 8637 3457
rect 9423 3447 9481 3453
rect 9423 3444 9435 3447
rect 8794 3416 9435 3444
rect 4915 3379 4973 3385
rect 4915 3376 4927 3379
rect 4233 3348 4927 3376
rect 4233 3335 4239 3348
rect 4915 3345 4927 3348
rect 4961 3345 4973 3379
rect 4915 3339 4973 3345
rect 6019 3379 6077 3385
rect 6019 3345 6031 3379
rect 6065 3376 6077 3379
rect 6383 3379 6441 3385
rect 6383 3376 6395 3379
rect 6065 3348 6395 3376
rect 6065 3345 6077 3348
rect 6019 3339 6077 3345
rect 6383 3345 6395 3348
rect 6429 3345 6441 3379
rect 6383 3339 6441 3345
rect 6568 3386 6634 3387
rect 6568 3334 6575 3386
rect 6627 3376 6634 3386
rect 8794 3385 8833 3416
rect 9423 3413 9435 3416
rect 9469 3413 9481 3447
rect 9423 3407 9481 3413
rect 10127 3407 10128 3459
rect 12467 3458 12520 3465
rect 10075 3400 10128 3407
rect 10974 3404 10981 3456
rect 11033 3404 11040 3456
rect 11815 3447 11873 3453
rect 11815 3444 11827 3447
rect 11186 3416 11827 3444
rect 7307 3379 7365 3385
rect 7307 3376 7319 3379
rect 6627 3348 7319 3376
rect 6627 3334 6634 3348
rect 7307 3345 7319 3348
rect 7353 3345 7365 3379
rect 8411 3379 8469 3385
rect 7307 3339 7365 3345
rect 8141 3355 8194 3362
rect 8193 3303 8194 3355
rect 8411 3345 8423 3379
rect 8457 3376 8469 3379
rect 8775 3379 8833 3385
rect 8775 3376 8787 3379
rect 8457 3348 8787 3376
rect 8457 3345 8469 3348
rect 8411 3339 8469 3345
rect 8775 3345 8787 3348
rect 8821 3345 8833 3379
rect 8775 3339 8833 3345
rect 8962 3385 9028 3386
rect 11186 3385 11225 3416
rect 11815 3413 11827 3416
rect 11861 3413 11873 3447
rect 11815 3407 11873 3413
rect 12519 3406 12520 3458
rect 12467 3399 12520 3406
rect 8962 3333 8969 3385
rect 9021 3376 9028 3385
rect 9699 3379 9757 3385
rect 9699 3376 9711 3379
rect 9021 3348 9711 3376
rect 9021 3333 9028 3348
rect 9699 3345 9711 3348
rect 9745 3345 9757 3379
rect 10803 3379 10861 3385
rect 9699 3339 9757 3345
rect 10533 3356 10586 3363
rect 8141 3296 8194 3303
rect 10585 3304 10586 3356
rect 10803 3345 10815 3379
rect 10849 3376 10861 3379
rect 11167 3379 11225 3385
rect 11167 3376 11179 3379
rect 10849 3348 11179 3376
rect 10849 3345 10861 3348
rect 10803 3339 10861 3345
rect 11167 3345 11179 3348
rect 11213 3345 11225 3379
rect 11167 3339 11225 3345
rect 11348 3386 11414 3387
rect 11348 3334 11355 3386
rect 11407 3376 11414 3386
rect 12091 3379 12149 3385
rect 12091 3376 12103 3379
rect 11407 3348 12103 3376
rect 11407 3334 11414 3348
rect 12091 3345 12103 3348
rect 12137 3345 12149 3379
rect 12091 3339 12149 3345
rect 12923 3359 12976 3366
rect 10533 3297 10586 3304
rect 12975 3307 12976 3359
rect 12923 3300 12976 3307
rect 13066 3240 13332 3310
rect 465 3209 13332 3240
rect 465 3208 3197 3209
rect 465 3174 655 3208
rect 689 3174 747 3208
rect 781 3174 839 3208
rect 873 3174 931 3208
rect 965 3174 1023 3208
rect 1057 3174 1115 3208
rect 1149 3174 1207 3208
rect 1241 3174 1299 3208
rect 1333 3174 1391 3208
rect 1425 3175 3197 3208
rect 3231 3175 3289 3209
rect 3323 3175 3381 3209
rect 3415 3175 3454 3209
rect 3488 3175 3546 3209
rect 3580 3175 3638 3209
rect 3672 3175 3730 3209
rect 3764 3175 3822 3209
rect 3856 3175 3914 3209
rect 3948 3175 4006 3209
rect 4040 3175 4098 3209
rect 4132 3175 4190 3209
rect 4224 3175 4282 3209
rect 4316 3175 4374 3209
rect 4408 3175 4466 3209
rect 4500 3175 4558 3209
rect 4592 3175 4650 3209
rect 4684 3175 4742 3209
rect 4776 3175 4834 3209
rect 4868 3175 4926 3209
rect 4960 3175 5018 3209
rect 5052 3175 5110 3209
rect 5144 3175 5202 3209
rect 5236 3175 5294 3209
rect 5328 3175 5386 3209
rect 5420 3175 5478 3209
rect 5512 3175 5570 3209
rect 5604 3175 5662 3209
rect 5696 3175 5754 3209
rect 5788 3175 5846 3209
rect 5880 3175 5938 3209
rect 5972 3175 6030 3209
rect 6064 3175 6122 3209
rect 6156 3175 6214 3209
rect 6248 3175 6306 3209
rect 6340 3175 6398 3209
rect 6432 3175 6490 3209
rect 6524 3175 6582 3209
rect 6616 3175 6674 3209
rect 6708 3175 6766 3209
rect 6800 3175 6858 3209
rect 6892 3175 6950 3209
rect 6984 3175 7042 3209
rect 7076 3175 7134 3209
rect 7168 3175 7226 3209
rect 7260 3175 7318 3209
rect 7352 3175 7410 3209
rect 7444 3175 7502 3209
rect 7536 3175 7594 3209
rect 7628 3175 7686 3209
rect 7720 3175 7778 3209
rect 7812 3175 7870 3209
rect 7904 3175 7962 3209
rect 7996 3175 8054 3209
rect 8088 3175 8146 3209
rect 8180 3175 8238 3209
rect 8272 3175 8330 3209
rect 8364 3175 8422 3209
rect 8456 3175 8514 3209
rect 8548 3175 8606 3209
rect 8640 3175 8698 3209
rect 8732 3175 8790 3209
rect 8824 3175 8882 3209
rect 8916 3175 8974 3209
rect 9008 3175 9066 3209
rect 9100 3175 9158 3209
rect 9192 3175 9250 3209
rect 9284 3175 9342 3209
rect 9376 3175 9434 3209
rect 9468 3175 9526 3209
rect 9560 3175 9618 3209
rect 9652 3175 9710 3209
rect 9744 3175 9802 3209
rect 9836 3175 9894 3209
rect 9928 3175 9986 3209
rect 10020 3175 10078 3209
rect 10112 3175 10170 3209
rect 10204 3175 10262 3209
rect 10296 3175 10354 3209
rect 10388 3175 10446 3209
rect 10480 3175 10538 3209
rect 10572 3175 10630 3209
rect 10664 3175 10722 3209
rect 10756 3175 10814 3209
rect 10848 3175 10906 3209
rect 10940 3175 10998 3209
rect 11032 3175 11090 3209
rect 11124 3175 11182 3209
rect 11216 3175 11274 3209
rect 11308 3175 11366 3209
rect 11400 3175 11458 3209
rect 11492 3175 11550 3209
rect 11584 3175 11642 3209
rect 11676 3175 11734 3209
rect 11768 3175 11826 3209
rect 11860 3175 11918 3209
rect 11952 3175 12010 3209
rect 12044 3175 12102 3209
rect 12136 3175 12194 3209
rect 12228 3175 12286 3209
rect 12320 3175 12378 3209
rect 12412 3175 12470 3209
rect 12504 3175 12562 3209
rect 12596 3175 12654 3209
rect 12688 3175 12746 3209
rect 12780 3175 12838 3209
rect 12872 3175 12930 3209
rect 12964 3182 13332 3209
rect 12964 3175 13142 3182
rect 1425 3174 13142 3175
rect 465 3144 13142 3174
rect 626 3143 1454 3144
rect 470 3066 504 3071
rect 640 3066 646 3082
rect 468 3038 646 3066
rect 470 3037 504 3038
rect 640 3030 646 3038
rect 698 3030 704 3082
rect 1260 3027 1266 3079
rect 1318 3066 1324 3079
rect 3000 3066 3007 3077
rect 1318 3038 3007 3066
rect 1318 3027 1324 3038
rect 3000 3025 3007 3038
rect 3059 3066 3066 3077
rect 5380 3066 5387 3078
rect 3059 3038 5387 3066
rect 3059 3025 3066 3038
rect 5380 3026 5387 3038
rect 5439 3066 5446 3078
rect 6179 3066 6186 3077
rect 5439 3038 6186 3066
rect 5439 3026 5446 3038
rect 6179 3025 6186 3038
rect 6238 3066 6245 3077
rect 7773 3066 7780 3077
rect 6238 3038 7780 3066
rect 6238 3025 6245 3038
rect 7773 3025 7780 3038
rect 7832 3066 7839 3077
rect 8568 3066 8575 3078
rect 7832 3038 8575 3066
rect 7832 3025 7839 3038
rect 8568 3026 8575 3038
rect 8627 3066 8634 3078
rect 10160 3066 10167 3077
rect 8627 3038 10167 3066
rect 8627 3026 8634 3038
rect 10160 3025 10167 3038
rect 10219 3066 10226 3077
rect 10977 3066 10984 3078
rect 10219 3038 10984 3066
rect 10219 3025 10226 3038
rect 10977 3026 10984 3038
rect 11036 3066 11043 3078
rect 12555 3066 12562 3078
rect 11036 3038 12562 3066
rect 11036 3026 11043 3038
rect 12555 3026 12562 3038
rect 12614 3066 12621 3078
rect 12614 3038 12998 3066
rect 12614 3026 12621 3038
rect 13062 3036 13142 3144
rect 13292 3036 13332 3182
rect 13062 2968 13332 3036
rect 555 2940 13332 2968
rect 555 2939 13058 2940
rect 363 2907 13212 2911
rect 290 2894 13212 2907
rect 290 2886 792 2894
rect 290 2740 442 2886
rect 592 2748 792 2886
rect 942 2880 13212 2894
rect 942 2846 1062 2880
rect 1096 2846 1154 2880
rect 1188 2846 1246 2880
rect 1280 2846 1338 2880
rect 1372 2846 1430 2880
rect 1464 2846 1522 2880
rect 1556 2846 1614 2880
rect 1648 2846 1706 2880
rect 1740 2846 1798 2880
rect 1832 2846 1890 2880
rect 1924 2846 1982 2880
rect 2016 2846 2074 2880
rect 2108 2846 2166 2880
rect 2200 2846 2258 2880
rect 2292 2846 2350 2880
rect 2384 2846 2442 2880
rect 2476 2846 2534 2880
rect 2568 2846 2626 2880
rect 2660 2846 2718 2880
rect 2752 2846 2810 2880
rect 2844 2846 2902 2880
rect 2936 2846 2994 2880
rect 3028 2846 3086 2880
rect 3120 2846 3178 2880
rect 3212 2846 3270 2880
rect 3304 2846 3362 2880
rect 3396 2846 3454 2880
rect 3488 2846 3546 2880
rect 3580 2846 3638 2880
rect 3672 2846 3730 2880
rect 3764 2846 3822 2880
rect 3856 2846 3914 2880
rect 3948 2846 4006 2880
rect 4040 2846 4098 2880
rect 4132 2846 4190 2880
rect 4224 2846 4282 2880
rect 4316 2846 4374 2880
rect 4408 2846 4466 2880
rect 4500 2846 4558 2880
rect 4592 2846 4650 2880
rect 4684 2846 4742 2880
rect 4776 2846 4834 2880
rect 4868 2846 4926 2880
rect 4960 2846 5018 2880
rect 5052 2846 5110 2880
rect 5144 2846 5202 2880
rect 5236 2846 5294 2880
rect 5328 2846 5386 2880
rect 5420 2846 5478 2880
rect 5512 2846 5570 2880
rect 5604 2846 5662 2880
rect 5696 2846 5754 2880
rect 5788 2846 5846 2880
rect 5880 2846 5938 2880
rect 5972 2846 6030 2880
rect 6064 2846 6122 2880
rect 6156 2846 6214 2880
rect 6248 2846 6306 2880
rect 6340 2846 6398 2880
rect 6432 2846 6490 2880
rect 6524 2846 6582 2880
rect 6616 2846 6674 2880
rect 6708 2846 6766 2880
rect 6800 2846 6858 2880
rect 6892 2846 6950 2880
rect 6984 2846 7042 2880
rect 7076 2846 7134 2880
rect 7168 2846 7226 2880
rect 7260 2846 7318 2880
rect 7352 2846 7410 2880
rect 7444 2846 7502 2880
rect 7536 2846 7594 2880
rect 7628 2846 7686 2880
rect 7720 2846 7778 2880
rect 7812 2846 7870 2880
rect 7904 2846 7962 2880
rect 7996 2846 8054 2880
rect 8088 2846 8146 2880
rect 8180 2846 8238 2880
rect 8272 2846 8330 2880
rect 8364 2846 8422 2880
rect 8456 2846 8514 2880
rect 8548 2846 8606 2880
rect 8640 2846 8698 2880
rect 8732 2846 8790 2880
rect 8824 2846 8882 2880
rect 8916 2846 8974 2880
rect 9008 2846 9066 2880
rect 9100 2846 9158 2880
rect 9192 2846 9250 2880
rect 9284 2846 9342 2880
rect 9376 2846 9434 2880
rect 9468 2846 9526 2880
rect 9560 2846 9618 2880
rect 9652 2846 9710 2880
rect 9744 2846 9802 2880
rect 9836 2846 9894 2880
rect 9928 2846 9986 2880
rect 10020 2846 10078 2880
rect 10112 2846 10170 2880
rect 10204 2846 10262 2880
rect 10296 2846 10354 2880
rect 10388 2846 10446 2880
rect 10480 2846 10538 2880
rect 10572 2846 10630 2880
rect 10664 2846 10722 2880
rect 10756 2846 10814 2880
rect 10848 2846 10906 2880
rect 10940 2846 10998 2880
rect 11032 2846 11090 2880
rect 11124 2846 11182 2880
rect 11216 2846 11274 2880
rect 11308 2846 11366 2880
rect 11400 2846 11458 2880
rect 11492 2846 11550 2880
rect 11584 2846 11642 2880
rect 11676 2846 11734 2880
rect 11768 2846 11826 2880
rect 11860 2846 11918 2880
rect 11952 2846 12010 2880
rect 12044 2846 12102 2880
rect 12136 2846 12194 2880
rect 12228 2846 12286 2880
rect 12320 2846 12378 2880
rect 12412 2846 12470 2880
rect 12504 2846 12562 2880
rect 12596 2846 12654 2880
rect 12688 2846 12746 2880
rect 12780 2846 12838 2880
rect 12872 2846 12930 2880
rect 12964 2846 13212 2880
rect 942 2815 13212 2846
rect 942 2748 974 2815
rect 592 2740 974 2748
rect 290 2466 974 2740
rect 2153 2710 2211 2716
rect 2153 2676 2165 2710
rect 2199 2707 2211 2710
rect 2889 2710 2947 2716
rect 2889 2707 2901 2710
rect 2199 2679 2901 2707
rect 2199 2676 2211 2679
rect 2153 2670 2211 2676
rect 2889 2676 2901 2679
rect 2935 2707 2947 2710
rect 3257 2710 3315 2716
rect 3257 2707 3269 2710
rect 2935 2679 3269 2707
rect 2935 2676 2947 2679
rect 2889 2670 2947 2676
rect 3257 2676 3269 2679
rect 3303 2676 3315 2710
rect 3257 2670 3315 2676
rect 4545 2710 4603 2716
rect 4545 2676 4557 2710
rect 4591 2707 4603 2710
rect 5281 2710 5339 2716
rect 5281 2707 5293 2710
rect 4591 2679 5293 2707
rect 4591 2676 4603 2679
rect 4545 2670 4603 2676
rect 5281 2676 5293 2679
rect 5327 2707 5339 2710
rect 5649 2710 5707 2716
rect 5649 2707 5661 2710
rect 5327 2679 5661 2707
rect 5327 2676 5339 2679
rect 5281 2670 5339 2676
rect 5649 2676 5661 2679
rect 5695 2676 5707 2710
rect 5649 2670 5707 2676
rect 6937 2710 6995 2716
rect 6937 2676 6949 2710
rect 6983 2707 6995 2710
rect 7673 2710 7731 2716
rect 7673 2707 7685 2710
rect 6983 2679 7685 2707
rect 6983 2676 6995 2679
rect 6937 2670 6995 2676
rect 7673 2676 7685 2679
rect 7719 2707 7731 2710
rect 8041 2710 8099 2716
rect 8041 2707 8053 2710
rect 7719 2679 8053 2707
rect 7719 2676 7731 2679
rect 7673 2670 7731 2676
rect 8041 2676 8053 2679
rect 8087 2676 8099 2710
rect 8041 2670 8099 2676
rect 9329 2710 9387 2716
rect 9329 2676 9341 2710
rect 9375 2707 9387 2710
rect 10065 2710 10123 2716
rect 10065 2707 10077 2710
rect 9375 2679 10077 2707
rect 9375 2676 9387 2679
rect 9329 2670 9387 2676
rect 10065 2676 10077 2679
rect 10111 2707 10123 2710
rect 10433 2710 10491 2716
rect 10433 2707 10445 2710
rect 10111 2679 10445 2707
rect 10111 2676 10123 2679
rect 10065 2670 10123 2676
rect 10433 2676 10445 2679
rect 10479 2676 10491 2710
rect 10433 2670 10491 2676
rect 11721 2710 11779 2716
rect 11721 2676 11733 2710
rect 11767 2707 11779 2710
rect 12457 2710 12515 2716
rect 12457 2707 12469 2710
rect 11767 2679 12469 2707
rect 11767 2676 11779 2679
rect 11721 2670 11779 2676
rect 12457 2676 12469 2679
rect 12503 2707 12515 2710
rect 12825 2710 12883 2716
rect 12825 2707 12837 2710
rect 12503 2679 12837 2707
rect 12503 2676 12515 2679
rect 12457 2670 12515 2676
rect 12825 2676 12837 2679
rect 12871 2676 12883 2710
rect 12825 2670 12883 2676
rect 1601 2642 1659 2648
rect 1601 2608 1613 2642
rect 1647 2639 1659 2642
rect 2245 2642 2303 2648
rect 2245 2639 2257 2642
rect 1647 2611 2257 2639
rect 1647 2608 1659 2611
rect 1601 2602 1659 2608
rect 2245 2608 2257 2611
rect 2291 2608 2303 2642
rect 3993 2642 4051 2648
rect 2245 2602 2303 2608
rect 2999 2588 3006 2640
rect 3058 2588 3065 2640
rect 3993 2608 4005 2642
rect 4039 2639 4051 2642
rect 4637 2642 4695 2648
rect 4637 2639 4649 2642
rect 4039 2611 4649 2639
rect 4039 2608 4051 2611
rect 3993 2602 4051 2608
rect 4637 2608 4649 2611
rect 4683 2608 4695 2642
rect 6385 2642 6443 2648
rect 4637 2602 4695 2608
rect 3887 2588 3940 2595
rect 1488 2530 1498 2582
rect 1550 2530 1562 2582
rect 2153 2574 2211 2580
rect 2153 2540 2165 2574
rect 2199 2571 2211 2574
rect 2199 2543 2840 2571
rect 2199 2540 2211 2543
rect 2153 2534 2211 2540
rect 1488 2528 1562 2530
rect 2612 2514 2678 2515
rect 1877 2506 1935 2512
rect 1877 2472 1889 2506
rect 1923 2503 1935 2506
rect 2612 2503 2619 2514
rect 1923 2475 2619 2503
rect 1923 2472 1935 2475
rect 1877 2466 1935 2472
rect 2612 2462 2619 2475
rect 2671 2462 2678 2514
rect 2801 2512 2840 2543
rect 3887 2536 3888 2588
rect 5380 2585 5387 2637
rect 5439 2585 5446 2637
rect 6385 2608 6397 2642
rect 6431 2639 6443 2642
rect 7029 2642 7087 2648
rect 7029 2639 7041 2642
rect 6431 2611 7041 2639
rect 6431 2608 6443 2611
rect 6385 2602 6443 2608
rect 7029 2608 7041 2611
rect 7075 2608 7087 2642
rect 8777 2642 8835 2648
rect 7029 2602 7087 2608
rect 6281 2586 6334 2593
rect 7771 2589 7778 2641
rect 7830 2589 7837 2641
rect 8777 2608 8789 2642
rect 8823 2639 8835 2642
rect 9421 2642 9479 2648
rect 11169 2642 11227 2648
rect 9421 2639 9433 2642
rect 8823 2611 9433 2639
rect 8823 2608 8835 2611
rect 8777 2602 8835 2608
rect 9421 2608 9433 2611
rect 9467 2608 9479 2642
rect 9421 2602 9479 2608
rect 3887 2529 3940 2536
rect 4545 2574 4603 2580
rect 4545 2540 4557 2574
rect 4591 2571 4603 2574
rect 4591 2543 5232 2571
rect 4591 2540 4603 2543
rect 4545 2534 4603 2540
rect 5193 2512 5232 2543
rect 6333 2534 6334 2586
rect 8673 2587 8726 2594
rect 10160 2590 10167 2642
rect 10219 2590 10226 2642
rect 11169 2608 11181 2642
rect 11215 2639 11227 2642
rect 11813 2642 11871 2648
rect 11813 2639 11825 2642
rect 11215 2611 11825 2639
rect 11215 2608 11227 2611
rect 11169 2602 11227 2608
rect 11813 2608 11825 2611
rect 11859 2608 11871 2642
rect 11813 2602 11871 2608
rect 6937 2574 6995 2580
rect 6937 2540 6949 2574
rect 6983 2571 6995 2574
rect 6983 2543 7624 2571
rect 6983 2540 6995 2543
rect 6937 2534 6995 2540
rect 6281 2527 6334 2534
rect 7585 2512 7624 2543
rect 8725 2535 8726 2587
rect 11066 2588 11119 2595
rect 12554 2590 12561 2642
rect 12613 2590 12620 2642
rect 12919 2595 12971 2597
rect 12916 2591 12973 2595
rect 8673 2528 8726 2535
rect 9329 2574 9387 2580
rect 9329 2540 9341 2574
rect 9375 2571 9387 2574
rect 9375 2543 10016 2571
rect 9375 2540 9387 2543
rect 9329 2534 9387 2540
rect 9977 2512 10016 2543
rect 11118 2536 11119 2588
rect 11066 2529 11119 2536
rect 11721 2574 11779 2580
rect 11721 2540 11733 2574
rect 11767 2571 11779 2574
rect 11767 2543 12408 2571
rect 11767 2540 11779 2543
rect 11721 2534 11779 2540
rect 12369 2512 12408 2543
rect 12916 2539 12919 2591
rect 12971 2539 12973 2591
rect 12916 2536 12973 2539
rect 12919 2533 12971 2536
rect 2801 2506 2859 2512
rect 2801 2472 2813 2506
rect 2847 2503 2859 2506
rect 3165 2506 3223 2512
rect 3165 2503 3177 2506
rect 2847 2475 3177 2503
rect 2847 2472 2859 2475
rect 2801 2466 2859 2472
rect 3165 2472 3177 2475
rect 3211 2472 3223 2506
rect 4269 2506 4327 2512
rect 3165 2466 3223 2472
rect 3442 2478 3495 2485
rect 1051 2455 1104 2462
rect 1103 2403 1104 2455
rect 3494 2426 3495 2478
rect 4269 2472 4281 2506
rect 4315 2503 4327 2506
rect 5005 2506 5063 2512
rect 5005 2503 5017 2506
rect 4315 2475 5017 2503
rect 4315 2472 4327 2475
rect 4269 2466 4327 2472
rect 5005 2472 5017 2475
rect 5051 2472 5063 2506
rect 5005 2466 5063 2472
rect 5193 2506 5251 2512
rect 5193 2472 5205 2506
rect 5239 2503 5251 2506
rect 5557 2506 5615 2512
rect 5557 2503 5569 2506
rect 5239 2475 5569 2503
rect 5239 2472 5251 2475
rect 5193 2466 5251 2472
rect 5557 2472 5569 2475
rect 5603 2472 5615 2506
rect 6661 2506 6719 2512
rect 5557 2466 5615 2472
rect 5833 2477 5886 2484
rect 3442 2419 3495 2426
rect 5017 2438 5051 2466
rect 5460 2438 5466 2447
rect 5017 2410 5466 2438
rect 1051 2396 1104 2403
rect 5460 2395 5466 2410
rect 5518 2395 5524 2447
rect 5885 2425 5886 2477
rect 6661 2472 6673 2506
rect 6707 2503 6719 2506
rect 7397 2506 7455 2512
rect 7397 2503 7409 2506
rect 6707 2475 7409 2503
rect 6707 2472 6719 2475
rect 6661 2466 6719 2472
rect 7397 2472 7409 2475
rect 7443 2472 7455 2506
rect 7397 2466 7455 2472
rect 7585 2506 7643 2512
rect 7585 2472 7597 2506
rect 7631 2503 7643 2506
rect 7949 2506 8007 2512
rect 7949 2503 7961 2506
rect 7631 2475 7961 2503
rect 7631 2472 7643 2475
rect 7585 2466 7643 2472
rect 7949 2472 7961 2475
rect 7995 2472 8007 2506
rect 9053 2506 9111 2512
rect 7949 2466 8007 2472
rect 8228 2480 8281 2487
rect 5833 2418 5886 2425
rect 7409 2438 7443 2466
rect 7852 2438 7858 2447
rect 7409 2410 7858 2438
rect 7852 2395 7858 2410
rect 7910 2395 7916 2447
rect 8280 2428 8281 2480
rect 9053 2472 9065 2506
rect 9099 2503 9111 2506
rect 9789 2506 9847 2512
rect 9789 2503 9801 2506
rect 9099 2475 9801 2503
rect 9099 2472 9111 2475
rect 9053 2466 9111 2472
rect 9789 2472 9801 2475
rect 9835 2472 9847 2506
rect 9789 2466 9847 2472
rect 9977 2506 10035 2512
rect 9977 2472 9989 2506
rect 10023 2503 10035 2506
rect 10341 2506 10399 2512
rect 10341 2503 10353 2506
rect 10023 2475 10353 2503
rect 10023 2472 10035 2475
rect 9977 2466 10035 2472
rect 10341 2472 10353 2475
rect 10387 2472 10399 2506
rect 11445 2506 11503 2512
rect 10341 2466 10399 2472
rect 10617 2478 10670 2485
rect 8228 2421 8281 2428
rect 9801 2438 9835 2466
rect 10244 2438 10250 2447
rect 9801 2410 10250 2438
rect 10244 2395 10250 2410
rect 10302 2395 10308 2447
rect 10669 2426 10670 2478
rect 11445 2472 11457 2506
rect 11491 2503 11503 2506
rect 12181 2506 12239 2512
rect 12181 2503 12193 2506
rect 11491 2475 12193 2503
rect 11491 2472 11503 2475
rect 11445 2466 11503 2472
rect 12181 2472 12193 2475
rect 12227 2472 12239 2506
rect 12181 2466 12239 2472
rect 12369 2506 12427 2512
rect 12369 2472 12381 2506
rect 12415 2503 12427 2506
rect 12733 2506 12791 2512
rect 12733 2503 12745 2506
rect 12415 2475 12745 2503
rect 12415 2472 12427 2475
rect 12369 2466 12427 2472
rect 12733 2472 12745 2475
rect 12779 2472 12791 2506
rect 12733 2466 12791 2472
rect 13072 2504 13332 2666
rect 10617 2419 10670 2426
rect 12193 2438 12227 2466
rect 12635 2438 12641 2447
rect 12193 2410 12641 2438
rect 12635 2395 12641 2410
rect 12693 2395 12699 2447
rect 13072 2367 13148 2504
rect 390 2358 13148 2367
rect 13298 2358 13332 2504
rect 390 2336 13332 2358
rect 390 2302 1062 2336
rect 1096 2302 1154 2336
rect 1188 2302 1246 2336
rect 1280 2302 1338 2336
rect 1372 2302 1430 2336
rect 1464 2302 1522 2336
rect 1556 2302 1614 2336
rect 1648 2302 1706 2336
rect 1740 2302 1798 2336
rect 1832 2302 1890 2336
rect 1924 2302 1982 2336
rect 2016 2302 2074 2336
rect 2108 2302 2166 2336
rect 2200 2302 2258 2336
rect 2292 2302 2350 2336
rect 2384 2302 2442 2336
rect 2476 2302 2534 2336
rect 2568 2302 2626 2336
rect 2660 2302 2718 2336
rect 2752 2302 2810 2336
rect 2844 2302 2902 2336
rect 2936 2302 2994 2336
rect 3028 2302 3086 2336
rect 3120 2302 3178 2336
rect 3212 2302 3270 2336
rect 3304 2302 3362 2336
rect 3396 2302 3454 2336
rect 3488 2302 3546 2336
rect 3580 2302 3638 2336
rect 3672 2302 3730 2336
rect 3764 2302 3822 2336
rect 3856 2302 3914 2336
rect 3948 2302 4006 2336
rect 4040 2302 4098 2336
rect 4132 2302 4190 2336
rect 4224 2302 4282 2336
rect 4316 2302 4374 2336
rect 4408 2302 4466 2336
rect 4500 2302 4558 2336
rect 4592 2302 4650 2336
rect 4684 2302 4742 2336
rect 4776 2302 4834 2336
rect 4868 2302 4926 2336
rect 4960 2302 5018 2336
rect 5052 2302 5110 2336
rect 5144 2302 5202 2336
rect 5236 2302 5294 2336
rect 5328 2302 5386 2336
rect 5420 2302 5478 2336
rect 5512 2302 5570 2336
rect 5604 2302 5662 2336
rect 5696 2302 5754 2336
rect 5788 2302 5846 2336
rect 5880 2302 5938 2336
rect 5972 2302 6030 2336
rect 6064 2302 6122 2336
rect 6156 2302 6214 2336
rect 6248 2302 6306 2336
rect 6340 2302 6398 2336
rect 6432 2302 6490 2336
rect 6524 2302 6582 2336
rect 6616 2302 6674 2336
rect 6708 2302 6766 2336
rect 6800 2302 6858 2336
rect 6892 2302 6950 2336
rect 6984 2302 7042 2336
rect 7076 2302 7134 2336
rect 7168 2302 7226 2336
rect 7260 2302 7318 2336
rect 7352 2302 7410 2336
rect 7444 2302 7502 2336
rect 7536 2302 7594 2336
rect 7628 2302 7686 2336
rect 7720 2302 7778 2336
rect 7812 2302 7870 2336
rect 7904 2302 7962 2336
rect 7996 2302 8054 2336
rect 8088 2302 8146 2336
rect 8180 2302 8238 2336
rect 8272 2302 8330 2336
rect 8364 2302 8422 2336
rect 8456 2302 8514 2336
rect 8548 2302 8606 2336
rect 8640 2302 8698 2336
rect 8732 2302 8790 2336
rect 8824 2302 8882 2336
rect 8916 2302 8974 2336
rect 9008 2302 9066 2336
rect 9100 2302 9158 2336
rect 9192 2302 9250 2336
rect 9284 2302 9342 2336
rect 9376 2302 9434 2336
rect 9468 2302 9526 2336
rect 9560 2302 9618 2336
rect 9652 2302 9710 2336
rect 9744 2302 9802 2336
rect 9836 2302 9894 2336
rect 9928 2302 9986 2336
rect 10020 2302 10078 2336
rect 10112 2302 10170 2336
rect 10204 2302 10262 2336
rect 10296 2302 10354 2336
rect 10388 2302 10446 2336
rect 10480 2302 10538 2336
rect 10572 2302 10630 2336
rect 10664 2302 10722 2336
rect 10756 2302 10814 2336
rect 10848 2302 10906 2336
rect 10940 2302 10998 2336
rect 11032 2302 11090 2336
rect 11124 2302 11182 2336
rect 11216 2302 11274 2336
rect 11308 2302 11366 2336
rect 11400 2302 11458 2336
rect 11492 2302 11550 2336
rect 11584 2302 11642 2336
rect 11676 2302 11734 2336
rect 11768 2302 11826 2336
rect 11860 2302 11918 2336
rect 11952 2302 12010 2336
rect 12044 2302 12102 2336
rect 12136 2302 12194 2336
rect 12228 2302 12286 2336
rect 12320 2302 12378 2336
rect 12412 2302 12470 2336
rect 12504 2302 12562 2336
rect 12596 2302 12654 2336
rect 12688 2302 12746 2336
rect 12780 2302 12838 2336
rect 12872 2302 12930 2336
rect 12964 2302 13332 2336
rect 390 2271 13332 2302
rect 13072 2270 13332 2271
<< via1 >>
rect 428 6028 578 6174
rect 740 6012 890 6158
rect 1697 5883 1749 5891
rect 1697 5849 1712 5883
rect 1712 5849 1746 5883
rect 1746 5849 1749 5883
rect 1697 5839 1749 5849
rect 2020 5838 2072 5890
rect 8120 5851 8172 5903
rect 3602 5813 3654 5821
rect 3602 5779 3613 5813
rect 3613 5779 3647 5813
rect 3647 5779 3654 5813
rect 3602 5769 3654 5779
rect 10528 5775 10580 5827
rect 3882 5752 3934 5759
rect 3882 5718 3891 5752
rect 3891 5718 3925 5752
rect 3925 5718 3934 5752
rect 3882 5707 3934 5718
rect 5731 5707 5783 5759
rect 1060 5464 1112 5516
rect 1721 5464 1773 5516
rect 3451 5464 3503 5516
rect 5834 5464 5886 5516
rect 8229 5464 8281 5516
rect 10624 5464 10676 5516
rect 12920 5464 12972 5516
rect 13146 5414 13296 5560
rect 492 5068 642 5214
rect 798 5080 948 5226
rect 12563 5159 12615 5211
rect 2022 5034 2074 5086
rect 1059 4994 1111 5003
rect 1059 4960 1067 4994
rect 1067 4960 1101 4994
rect 1101 4960 1111 4994
rect 1059 4951 1111 4960
rect 3449 4994 3501 5003
rect 3449 4960 3457 4994
rect 3457 4960 3491 4994
rect 3491 4960 3501 4994
rect 3449 4951 3501 4960
rect 2527 4941 2579 4948
rect 2527 4907 2536 4941
rect 2536 4907 2570 4941
rect 2570 4907 2579 4941
rect 2527 4896 2579 4907
rect 5293 5011 5345 5022
rect 5293 4977 5305 5011
rect 5305 4977 5339 5011
rect 5339 4977 5345 5011
rect 5293 4970 5345 4977
rect 5842 4995 5894 5004
rect 5842 4961 5850 4995
rect 5850 4961 5884 4995
rect 5884 4961 5894 4995
rect 5842 4952 5894 4961
rect 7686 5012 7738 5021
rect 7686 4978 7695 5012
rect 7695 4978 7729 5012
rect 7729 4978 7738 5012
rect 7686 4969 7738 4978
rect 8234 4994 8286 5003
rect 8234 4960 8242 4994
rect 8242 4960 8276 4994
rect 8276 4960 8286 4994
rect 8234 4951 8286 4960
rect 10077 5014 10129 5023
rect 10077 4980 10086 5014
rect 10086 4980 10120 5014
rect 10120 4980 10129 5014
rect 10077 4971 10129 4980
rect 10629 4996 10681 5005
rect 10629 4962 10637 4996
rect 10637 4962 10671 4996
rect 10671 4962 10681 4996
rect 10629 4953 10681 4962
rect 12468 5012 12520 5021
rect 12468 4978 12477 5012
rect 12477 4978 12511 5012
rect 12511 4978 12520 5012
rect 12468 4969 12520 4978
rect 13146 4988 13296 5134
rect 3077 4883 3129 4890
rect 3077 4849 3087 4883
rect 3087 4849 3121 4883
rect 3121 4849 3129 4883
rect 3077 4838 3129 4849
rect 5467 4894 5519 4904
rect 5467 4860 5476 4894
rect 5476 4860 5510 4894
rect 5510 4860 5519 4894
rect 5467 4852 5519 4860
rect 5577 4863 5629 4915
rect 7856 4897 7908 4912
rect 7856 4863 7864 4897
rect 7864 4863 7898 4897
rect 7898 4863 7908 4897
rect 7856 4860 7908 4863
rect 7973 4852 8025 4904
rect 10252 4880 10304 4889
rect 10252 4846 10261 4880
rect 10261 4846 10295 4880
rect 10295 4846 10304 4880
rect 10252 4837 10304 4846
rect 10373 4868 10425 4920
rect 12643 4881 12695 4890
rect 12643 4847 12652 4881
rect 12652 4847 12686 4881
rect 12686 4847 12695 4881
rect 12643 4838 12695 4847
rect 12768 4868 12820 4920
rect 13146 4762 13296 4908
rect 324 4440 474 4586
rect 2528 4488 2580 4498
rect 2528 4454 2538 4488
rect 2538 4454 2572 4488
rect 2572 4454 2580 4488
rect 3442 4524 3494 4532
rect 3442 4490 3452 4524
rect 3452 4490 3486 4524
rect 3486 4490 3494 4524
rect 3442 4480 3494 4490
rect 5840 4462 5892 4514
rect 8231 4462 8283 4514
rect 2528 4446 2580 4454
rect 5834 4390 5886 4397
rect 5834 4356 5841 4390
rect 5841 4356 5875 4390
rect 5875 4356 5886 4390
rect 5834 4345 5886 4356
rect 3888 4322 3940 4332
rect 3888 4288 3898 4322
rect 3898 4288 3932 4322
rect 3932 4288 3940 4322
rect 3888 4280 3940 4288
rect 8222 4390 8274 4395
rect 8222 4356 8233 4390
rect 8233 4356 8267 4390
rect 8267 4356 8274 4390
rect 8222 4343 8274 4356
rect 6283 4324 6335 4333
rect 6283 4290 6292 4324
rect 6292 4290 6326 4324
rect 6326 4290 6335 4324
rect 6283 4281 6335 4290
rect 10619 4453 10671 4505
rect 10614 4391 10666 4396
rect 10614 4357 10625 4391
rect 10625 4357 10659 4391
rect 10659 4357 10666 4391
rect 10614 4344 10666 4357
rect 8673 4325 8725 4334
rect 8673 4291 8682 4325
rect 8682 4291 8716 4325
rect 8716 4291 8725 4325
rect 8673 4282 8725 4291
rect 3356 4187 3408 4194
rect 3356 4153 3366 4187
rect 3366 4153 3400 4187
rect 3400 4153 3408 4187
rect 3356 4142 3408 4153
rect 5976 4177 6028 4229
rect 12566 4383 12618 4388
rect 12566 4349 12575 4383
rect 12575 4349 12609 4383
rect 12609 4349 12618 4383
rect 12566 4336 12618 4349
rect 11067 4322 11119 4331
rect 11067 4288 11076 4322
rect 11076 4288 11110 4322
rect 11110 4288 11119 4322
rect 11067 4279 11119 4288
rect 12920 4375 12972 4383
rect 12920 4341 12930 4375
rect 12930 4341 12964 4375
rect 12964 4341 12972 4375
rect 12920 4331 12972 4341
rect 6574 4141 6626 4193
rect 8398 4166 8450 4218
rect 8966 4142 9018 4194
rect 10786 4174 10838 4226
rect 11355 4143 11407 4195
rect 13162 4028 13312 4174
rect 1496 3900 1548 3952
rect 3356 3900 3408 3952
rect 3888 3900 3940 3952
rect 5292 3900 5344 3952
rect 6277 3900 6329 3952
rect 7684 3900 7736 3952
rect 8667 3900 8719 3952
rect 10081 3900 10133 3952
rect 11057 3900 11109 3952
rect 12469 3900 12521 3952
rect 360 3594 510 3740
rect 712 3718 747 3744
rect 747 3718 781 3744
rect 781 3718 839 3744
rect 839 3718 862 3744
rect 1158 3718 1207 3744
rect 1207 3718 1241 3744
rect 1241 3718 1299 3744
rect 1299 3718 1308 3744
rect 712 3598 862 3718
rect 1158 3598 1308 3718
rect 1724 3602 1874 3748
rect 2390 3602 2540 3748
rect 2772 3586 2922 3732
rect 656 3439 708 3449
rect 656 3405 665 3439
rect 665 3405 699 3439
rect 699 3405 708 3439
rect 656 3397 708 3405
rect 1263 3440 1315 3449
rect 1263 3406 1270 3440
rect 1270 3406 1304 3440
rect 1304 3406 1315 3440
rect 1263 3397 1315 3406
rect 2622 3472 2674 3524
rect 3067 3471 3119 3523
rect 4189 3472 4241 3524
rect 2019 3399 2071 3451
rect 5293 3446 5345 3453
rect 5293 3412 5303 3446
rect 5303 3412 5337 3446
rect 5337 3412 5345 3446
rect 5293 3401 5345 3412
rect 6191 3449 6243 3457
rect 6191 3415 6200 3449
rect 6200 3415 6234 3449
rect 6234 3415 6243 3449
rect 6191 3405 6243 3415
rect 7684 3454 7736 3463
rect 4181 3379 4233 3387
rect 4181 3345 4191 3379
rect 4191 3345 4225 3379
rect 4225 3345 4233 3379
rect 7684 3420 7693 3454
rect 7693 3420 7727 3454
rect 7727 3420 7736 3454
rect 7684 3411 7736 3420
rect 8578 3449 8630 3457
rect 8578 3415 8587 3449
rect 8587 3415 8621 3449
rect 8621 3415 8630 3449
rect 8578 3405 8630 3415
rect 4181 3335 4233 3345
rect 6575 3379 6627 3386
rect 6575 3345 6583 3379
rect 6583 3345 6617 3379
rect 6617 3345 6627 3379
rect 10075 3450 10127 3459
rect 10075 3416 10084 3450
rect 10084 3416 10118 3450
rect 10118 3416 10127 3450
rect 10075 3407 10127 3416
rect 10981 3448 11033 3456
rect 10981 3414 10990 3448
rect 10990 3414 11024 3448
rect 11024 3414 11033 3448
rect 10981 3404 11033 3414
rect 6575 3334 6627 3345
rect 8141 3347 8193 3355
rect 8141 3313 8149 3347
rect 8149 3313 8183 3347
rect 8183 3313 8193 3347
rect 8141 3303 8193 3313
rect 12467 3449 12519 3458
rect 12467 3415 12476 3449
rect 12476 3415 12510 3449
rect 12510 3415 12519 3449
rect 12467 3406 12519 3415
rect 8969 3379 9021 3385
rect 8969 3345 8975 3379
rect 8975 3345 9009 3379
rect 9009 3345 9021 3379
rect 8969 3333 9021 3345
rect 10533 3348 10585 3356
rect 10533 3314 10541 3348
rect 10541 3314 10575 3348
rect 10575 3314 10585 3348
rect 10533 3304 10585 3314
rect 11355 3379 11407 3386
rect 11355 3345 11367 3379
rect 11367 3345 11401 3379
rect 11401 3345 11407 3379
rect 11355 3334 11407 3345
rect 12923 3351 12975 3359
rect 12923 3317 12931 3351
rect 12931 3317 12965 3351
rect 12965 3317 12975 3351
rect 12923 3307 12975 3317
rect 646 3030 698 3082
rect 1266 3027 1318 3079
rect 3007 3025 3059 3077
rect 5387 3026 5439 3078
rect 6186 3025 6238 3077
rect 7780 3025 7832 3077
rect 8575 3026 8627 3078
rect 10167 3025 10219 3077
rect 10984 3026 11036 3078
rect 12562 3026 12614 3078
rect 13142 3036 13292 3182
rect 442 2740 592 2886
rect 792 2748 942 2894
rect 3006 2632 3058 2640
rect 3006 2598 3015 2632
rect 3015 2598 3049 2632
rect 3049 2598 3058 2632
rect 3006 2588 3058 2598
rect 1498 2572 1550 2582
rect 1498 2538 1503 2572
rect 1503 2538 1537 2572
rect 1537 2538 1550 2572
rect 1498 2530 1550 2538
rect 2619 2506 2671 2514
rect 2619 2472 2625 2506
rect 2625 2472 2659 2506
rect 2659 2472 2671 2506
rect 2619 2462 2671 2472
rect 3888 2577 3940 2588
rect 5387 2629 5439 2637
rect 5387 2595 5396 2629
rect 5396 2595 5430 2629
rect 5430 2595 5439 2629
rect 5387 2585 5439 2595
rect 7778 2633 7830 2641
rect 7778 2599 7787 2633
rect 7787 2599 7821 2633
rect 7821 2599 7830 2633
rect 7778 2589 7830 2599
rect 3888 2543 3896 2577
rect 3896 2543 3930 2577
rect 3930 2543 3940 2577
rect 3888 2536 3940 2543
rect 6281 2577 6333 2586
rect 6281 2543 6290 2577
rect 6290 2543 6324 2577
rect 6324 2543 6333 2577
rect 6281 2534 6333 2543
rect 10167 2634 10219 2642
rect 10167 2600 10176 2634
rect 10176 2600 10210 2634
rect 10210 2600 10219 2634
rect 10167 2590 10219 2600
rect 8673 2578 8725 2587
rect 8673 2544 8682 2578
rect 8682 2544 8716 2578
rect 8716 2544 8725 2578
rect 8673 2535 8725 2544
rect 12561 2634 12613 2642
rect 12561 2600 12570 2634
rect 12570 2600 12604 2634
rect 12604 2600 12613 2634
rect 12561 2590 12613 2600
rect 11066 2579 11118 2588
rect 11066 2545 11075 2579
rect 11075 2545 11109 2579
rect 11109 2545 11118 2579
rect 11066 2536 11118 2545
rect 12919 2583 12971 2591
rect 12919 2549 12927 2583
rect 12927 2549 12961 2583
rect 12961 2549 12971 2583
rect 12919 2539 12971 2549
rect 3442 2470 3494 2478
rect 1051 2447 1103 2455
rect 1051 2413 1059 2447
rect 1059 2413 1093 2447
rect 1093 2413 1103 2447
rect 1051 2403 1103 2413
rect 3442 2436 3450 2470
rect 3450 2436 3484 2470
rect 3484 2436 3494 2470
rect 3442 2426 3494 2436
rect 5833 2469 5885 2477
rect 5466 2395 5518 2447
rect 5833 2435 5841 2469
rect 5841 2435 5875 2469
rect 5875 2435 5885 2469
rect 5833 2425 5885 2435
rect 8228 2472 8280 2480
rect 7858 2395 7910 2447
rect 8228 2438 8236 2472
rect 8236 2438 8270 2472
rect 8270 2438 8280 2472
rect 8228 2428 8280 2438
rect 10617 2470 10669 2478
rect 10250 2395 10302 2447
rect 10617 2436 10625 2470
rect 10625 2436 10659 2470
rect 10659 2436 10669 2470
rect 10617 2426 10669 2436
rect 12641 2395 12693 2447
rect 13148 2358 13298 2504
<< metal2 >>
rect 418 6174 590 6184
rect 418 6028 428 6174
rect 578 6028 590 6174
rect 418 6018 590 6028
rect 730 6158 902 6168
rect 730 6012 740 6158
rect 890 6012 902 6158
rect 730 6002 902 6012
rect 8120 5903 8173 5910
rect 1690 5839 1697 5891
rect 1749 5839 1758 5891
rect 1730 5517 1758 5839
rect 2013 5890 2079 5891
rect 2013 5838 2020 5890
rect 2072 5838 2079 5890
rect 8172 5851 8173 5903
rect 8120 5844 8173 5851
rect 1053 5516 1119 5517
rect 1053 5464 1060 5516
rect 1112 5464 1119 5516
rect 1714 5516 1780 5517
rect 1714 5464 1721 5516
rect 1773 5464 1780 5516
rect 788 5226 960 5236
rect 482 5214 654 5224
rect 482 5068 492 5214
rect 642 5068 654 5214
rect 788 5080 798 5226
rect 948 5080 960 5226
rect 788 5070 960 5080
rect 482 5058 654 5068
rect 1071 5029 1099 5464
rect 2032 5086 2060 5838
rect 3596 5769 3602 5821
rect 3654 5769 3660 5821
rect 3444 5516 3510 5517
rect 3444 5464 3451 5516
rect 3503 5464 3510 5516
rect 2015 5034 2022 5086
rect 2074 5034 2081 5086
rect 1070 5004 1099 5029
rect 1052 5003 1118 5004
rect 1052 4951 1059 5003
rect 1111 4951 1118 5003
rect 314 4586 486 4596
rect 314 4440 324 4586
rect 474 4440 486 4586
rect 314 4430 486 4440
rect 1489 3900 1496 3952
rect 1548 3900 1555 3952
rect 350 3740 522 3750
rect 350 3594 360 3740
rect 510 3594 522 3740
rect 350 3584 522 3594
rect 702 3744 874 3754
rect 702 3598 712 3744
rect 862 3598 874 3744
rect 702 3588 874 3598
rect 1148 3744 1320 3754
rect 1148 3598 1158 3744
rect 1308 3598 1320 3744
rect 1148 3588 1320 3598
rect 650 3397 656 3449
rect 708 3397 714 3449
rect 1257 3397 1263 3449
rect 1315 3397 1321 3449
rect 654 3082 690 3397
rect 640 3030 646 3082
rect 698 3030 704 3082
rect 1271 3079 1307 3397
rect 1260 3027 1266 3079
rect 1318 3027 1324 3079
rect 432 2886 604 2896
rect 432 2740 442 2886
rect 592 2740 604 2886
rect 432 2730 604 2740
rect 782 2894 954 2904
rect 782 2748 792 2894
rect 942 2748 954 2894
rect 782 2738 954 2748
rect 1508 2582 1536 3900
rect 1714 3748 1886 3758
rect 1714 3602 1724 3748
rect 1874 3602 1886 3748
rect 1714 3592 1886 3602
rect 2032 3452 2060 5034
rect 3464 5004 3492 5464
rect 3442 5003 3508 5004
rect 3442 4951 3449 5003
rect 3501 4951 3508 5003
rect 2520 4948 2586 4949
rect 2520 4896 2527 4948
rect 2579 4896 2586 4948
rect 2535 4505 2568 4896
rect 3070 4890 3136 4891
rect 3070 4838 3077 4890
rect 3129 4838 3136 4890
rect 2527 4498 2580 4505
rect 2527 4446 2528 4498
rect 2527 4439 2580 4446
rect 2380 3748 2552 3758
rect 2380 3602 2390 3748
rect 2540 3602 2552 3748
rect 2380 3592 2552 3602
rect 2762 3732 2934 3742
rect 2762 3586 2772 3732
rect 2922 3586 2934 3732
rect 2762 3576 2934 3586
rect 2616 3525 2681 3526
rect 2615 3524 2681 3525
rect 3094 3524 3122 4838
rect 3436 4480 3442 4532
rect 3494 4525 3500 4532
rect 3608 4525 3641 5769
rect 3875 5707 3882 5759
rect 3934 5707 3941 5759
rect 5724 5707 5731 5759
rect 5783 5707 5790 5759
rect 3875 5706 3941 5707
rect 5286 4970 5293 5022
rect 5345 4970 5351 5022
rect 3494 4490 3641 4525
rect 3494 4480 3500 4490
rect 3888 4332 3941 4339
rect 3940 4280 3941 4332
rect 3888 4273 3941 4280
rect 3349 4194 3415 4195
rect 3349 4142 3356 4194
rect 3408 4142 3415 4194
rect 3369 3953 3397 4142
rect 3900 3953 3928 4273
rect 5305 3953 5333 4970
rect 5576 4915 5629 4922
rect 5460 4904 5524 4910
rect 5460 4852 5467 4904
rect 5519 4852 5524 4904
rect 5576 4863 5577 4915
rect 5576 4856 5629 4863
rect 5460 4851 5524 4852
rect 5460 4846 5523 4851
rect 3349 3952 3415 3953
rect 3349 3900 3356 3952
rect 3408 3900 3415 3952
rect 3881 3952 3947 3953
rect 3881 3900 3888 3952
rect 3940 3900 3947 3952
rect 5285 3952 5351 3953
rect 5285 3900 5292 3952
rect 5344 3900 5351 3952
rect 2615 3472 2622 3524
rect 2674 3472 2681 3524
rect 3060 3523 3126 3524
rect 2012 3451 2078 3452
rect 2012 3399 2019 3451
rect 2071 3399 2078 3451
rect 1488 2530 1498 2582
rect 1550 2530 1562 2582
rect 1488 2528 1562 2530
rect 2629 2515 2657 3472
rect 3060 3471 3067 3523
rect 3119 3471 3126 3523
rect 3000 3025 3007 3077
rect 3059 3025 3066 3077
rect 3020 2640 3048 3025
rect 2999 2588 3006 2640
rect 3058 2588 3065 2640
rect 3900 2595 3928 3900
rect 4181 3472 4189 3524
rect 4241 3472 4248 3524
rect 4194 3388 4222 3472
rect 5305 3460 5333 3900
rect 5293 3453 5346 3460
rect 5345 3401 5346 3453
rect 5293 3394 5346 3401
rect 4175 3387 4239 3388
rect 4175 3335 4181 3387
rect 4233 3335 4239 3387
rect 5380 3026 5387 3078
rect 5439 3026 5446 3078
rect 5400 2637 5428 3026
rect 3887 2588 3940 2595
rect 3887 2536 3888 2588
rect 5380 2585 5387 2637
rect 5439 2585 5446 2637
rect 3887 2529 3940 2536
rect 2612 2514 2678 2515
rect 2612 2462 2619 2514
rect 2671 2462 2678 2514
rect 3442 2478 3495 2485
rect 1051 2455 1104 2462
rect 1103 2403 1104 2455
rect 3494 2426 3495 2478
rect 5476 2447 5509 4846
rect 3442 2419 3495 2426
rect 1051 2396 1104 2403
rect 1063 1784 1091 2396
rect 3454 1784 3482 2419
rect 5460 2395 5466 2447
rect 5518 2395 5524 2447
rect 5476 2392 5509 2395
rect 1058 1750 1092 1784
rect 3450 1750 3484 1784
rect 5589 1782 5617 4856
rect 5739 4390 5772 5707
rect 5827 5516 5893 5517
rect 5827 5464 5834 5516
rect 5886 5464 5893 5516
rect 5847 5005 5875 5464
rect 7686 5021 7739 5028
rect 5835 5004 5901 5005
rect 5835 4952 5842 5004
rect 5894 4952 5901 5004
rect 7738 4969 7739 5021
rect 7686 4962 7739 4969
rect 5847 4515 5875 4952
rect 5833 4514 5899 4515
rect 5833 4462 5840 4514
rect 5892 4462 5899 4514
rect 5833 4397 5886 4404
rect 5833 4390 5834 4397
rect 5739 4356 5834 4390
rect 5833 4345 5834 4356
rect 5833 4338 5886 4345
rect 6283 4333 6336 4340
rect 6335 4281 6336 4333
rect 6283 4274 6336 4281
rect 5976 4229 6029 4236
rect 6028 4177 6029 4229
rect 5976 4170 6029 4177
rect 5833 2477 5886 2484
rect 5885 2425 5886 2477
rect 5833 2418 5886 2425
rect 5845 1782 5873 2418
rect 1063 1748 1091 1750
rect 3454 1748 3482 1750
rect 5586 1748 5620 1782
rect 5844 1748 5878 1782
rect 5988 1779 6016 4170
rect 6292 3953 6320 4274
rect 6567 4193 6633 4194
rect 6567 4141 6574 4193
rect 6626 4141 6633 4193
rect 6270 3952 6336 3953
rect 6270 3900 6277 3952
rect 6329 3900 6336 3952
rect 6184 3405 6191 3457
rect 6243 3405 6250 3457
rect 6197 3077 6225 3405
rect 6179 3025 6186 3077
rect 6238 3025 6245 3077
rect 6292 2593 6320 3900
rect 6584 3387 6612 4141
rect 7697 3953 7725 4962
rect 7850 4860 7856 4912
rect 7908 4860 7914 4912
rect 7850 4852 7914 4860
rect 7972 4904 8025 4911
rect 7972 4852 7973 4904
rect 7677 3952 7743 3953
rect 7677 3900 7684 3952
rect 7736 3900 7743 3952
rect 7697 3470 7725 3900
rect 7684 3463 7737 3470
rect 7736 3411 7737 3463
rect 7684 3404 7737 3411
rect 6568 3386 6634 3387
rect 6568 3334 6575 3386
rect 6627 3334 6634 3386
rect 7773 3025 7780 3077
rect 7832 3025 7839 3077
rect 7793 2641 7821 3025
rect 6281 2586 6334 2593
rect 7771 2589 7778 2641
rect 7830 2589 7837 2641
rect 6333 2534 6334 2586
rect 6281 2527 6334 2534
rect 7867 2447 7900 4852
rect 7972 4845 8025 4852
rect 7852 2395 7858 2447
rect 7910 2395 7916 2447
rect 7985 1784 8013 4845
rect 8129 4390 8162 5844
rect 10528 5827 10581 5834
rect 10580 5775 10581 5827
rect 10528 5768 10581 5775
rect 8222 5516 8288 5517
rect 8222 5464 8229 5516
rect 8281 5464 8288 5516
rect 8242 5004 8270 5464
rect 10077 5023 10130 5030
rect 8227 5003 8293 5004
rect 8227 4951 8234 5003
rect 8286 4951 8293 5003
rect 10129 4971 10130 5023
rect 10077 4964 10130 4971
rect 8242 4515 8270 4951
rect 8224 4514 8290 4515
rect 8224 4462 8231 4514
rect 8283 4462 8290 4514
rect 8221 4395 8274 4402
rect 8221 4390 8222 4395
rect 8129 4356 8222 4390
rect 8130 4355 8222 4356
rect 8221 4343 8222 4355
rect 8221 4336 8274 4343
rect 8673 4334 8726 4341
rect 8725 4282 8726 4334
rect 8673 4275 8726 4282
rect 8398 4218 8451 4225
rect 8450 4166 8451 4218
rect 8398 4159 8451 4166
rect 8141 3355 8194 3362
rect 8193 3303 8194 3355
rect 8141 3296 8194 3303
rect 8153 1898 8181 3296
rect 8228 2480 8281 2487
rect 8280 2428 8281 2480
rect 8228 2421 8281 2428
rect 8151 1864 8185 1898
rect 5986 1745 6020 1779
rect 7982 1750 8016 1784
rect 7985 1748 8013 1750
rect 8153 1748 8181 1864
rect 8240 1844 8268 2421
rect 8238 1810 8272 1844
rect 8240 1748 8268 1810
rect 8410 1779 8438 4159
rect 8684 3953 8712 4275
rect 8959 4194 9025 4195
rect 8959 4142 8966 4194
rect 9018 4142 9025 4194
rect 8660 3952 8726 3953
rect 8660 3900 8667 3952
rect 8719 3900 8726 3952
rect 8571 3405 8578 3457
rect 8630 3405 8637 3457
rect 8586 3078 8614 3405
rect 8568 3026 8575 3078
rect 8627 3026 8634 3078
rect 8684 2594 8712 3900
rect 8977 3386 9005 4142
rect 10089 3953 10117 4964
rect 10372 4920 10425 4927
rect 10252 4889 10305 4896
rect 10304 4837 10305 4889
rect 10372 4868 10373 4920
rect 10372 4861 10425 4868
rect 10252 4830 10305 4837
rect 10074 3952 10140 3953
rect 10074 3900 10081 3952
rect 10133 3900 10140 3952
rect 10089 3466 10117 3900
rect 10075 3459 10128 3466
rect 10127 3407 10128 3459
rect 10075 3400 10128 3407
rect 8962 3385 9028 3386
rect 8962 3333 8969 3385
rect 9021 3333 9028 3385
rect 10160 3025 10167 3077
rect 10219 3025 10226 3077
rect 10180 2642 10208 3025
rect 8673 2587 8726 2594
rect 10160 2590 10167 2642
rect 10219 2590 10226 2642
rect 8725 2535 8726 2587
rect 8673 2528 8726 2535
rect 10259 2447 10292 4830
rect 10244 2395 10250 2447
rect 10302 2395 10308 2447
rect 10385 1779 10413 4861
rect 10537 4391 10570 5768
rect 13136 5560 13308 5570
rect 10617 5516 10683 5517
rect 10617 5464 10624 5516
rect 10676 5464 10683 5516
rect 12913 5516 12979 5517
rect 12913 5464 12920 5516
rect 12972 5464 12979 5516
rect 10637 5006 10665 5464
rect 12557 5211 12622 5216
rect 12557 5159 12563 5211
rect 12615 5159 12622 5211
rect 12557 5149 12622 5159
rect 12468 5021 12521 5028
rect 10622 5005 10688 5006
rect 10622 4953 10629 5005
rect 10681 4953 10688 5005
rect 12520 4969 12521 5021
rect 12468 4962 12521 4969
rect 10637 4511 10665 4953
rect 10618 4505 10671 4511
rect 10618 4453 10619 4505
rect 10618 4445 10671 4453
rect 10613 4396 10666 4403
rect 10613 4391 10614 4396
rect 10537 4357 10614 4391
rect 10613 4344 10614 4357
rect 10613 4337 10666 4344
rect 11067 4331 11120 4338
rect 11119 4279 11120 4331
rect 11067 4272 11120 4279
rect 10786 4226 10839 4233
rect 10838 4174 10839 4226
rect 10786 4167 10839 4174
rect 10533 3356 10586 3363
rect 10585 3304 10586 3356
rect 10533 3297 10586 3304
rect 10545 1870 10573 3297
rect 10617 2478 10670 2485
rect 10669 2426 10670 2478
rect 10617 2419 10670 2426
rect 10629 1870 10657 2419
rect 10544 1836 10578 1870
rect 10627 1836 10661 1870
rect 8406 1745 8440 1779
rect 10382 1745 10416 1779
rect 10545 1748 10573 1836
rect 10629 1748 10657 1836
rect 10798 1782 10826 4167
rect 11076 3953 11104 4272
rect 11348 4195 11414 4196
rect 11348 4143 11355 4195
rect 11407 4143 11414 4195
rect 11050 3952 11116 3953
rect 11050 3900 11057 3952
rect 11109 3900 11116 3952
rect 10974 3404 10981 3456
rect 11033 3404 11040 3456
rect 10995 3078 11023 3404
rect 10977 3026 10984 3078
rect 11036 3026 11043 3078
rect 11076 2595 11104 3900
rect 11369 3387 11397 4143
rect 12481 3953 12509 4962
rect 12575 4388 12608 5149
rect 12933 5148 12961 5464
rect 13136 5414 13146 5560
rect 13296 5414 13308 5560
rect 13136 5404 13308 5414
rect 12767 4920 12820 4927
rect 12643 4890 12696 4897
rect 12695 4838 12696 4890
rect 12767 4868 12768 4920
rect 12767 4861 12820 4868
rect 12643 4831 12696 4838
rect 12560 4336 12566 4388
rect 12618 4336 12624 4388
rect 12462 3952 12528 3953
rect 12462 3900 12469 3952
rect 12521 3900 12528 3952
rect 12481 3465 12509 3900
rect 12467 3458 12520 3465
rect 12519 3406 12520 3458
rect 12467 3399 12520 3406
rect 11348 3386 11414 3387
rect 11348 3334 11355 3386
rect 11407 3334 11414 3386
rect 12555 3026 12562 3078
rect 12614 3026 12621 3078
rect 12575 2642 12603 3026
rect 11066 2588 11119 2595
rect 12554 2590 12561 2642
rect 12613 2590 12620 2642
rect 11118 2536 11119 2588
rect 11066 2529 11119 2536
rect 12652 2447 12685 4831
rect 12635 2395 12641 2447
rect 12693 2395 12699 2447
rect 10795 1748 10829 1782
rect 12780 1779 12808 4861
rect 12932 4383 12965 5148
rect 13136 5134 13308 5144
rect 13136 4988 13146 5134
rect 13296 4988 13308 5134
rect 13136 4978 13308 4988
rect 13136 4908 13308 4918
rect 13136 4762 13146 4908
rect 13296 4762 13308 4908
rect 13136 4752 13308 4762
rect 12914 4331 12920 4383
rect 12972 4331 12978 4383
rect 12914 4330 12978 4331
rect 13152 4174 13324 4184
rect 13152 4028 13162 4174
rect 13312 4028 13324 4174
rect 13152 4018 13324 4028
rect 12923 3359 12976 3366
rect 12975 3307 12976 3359
rect 12923 3300 12976 3307
rect 12935 2597 12963 3300
rect 13132 3182 13304 3192
rect 13132 3036 13142 3182
rect 13292 3036 13304 3182
rect 13132 3026 13304 3036
rect 12919 2591 12971 2597
rect 12919 2533 12971 2539
rect 12935 1854 12963 2533
rect 13138 2504 13310 2514
rect 13138 2358 13148 2504
rect 13298 2358 13310 2504
rect 13138 2348 13310 2358
rect 12932 1820 12966 1854
rect 12776 1745 12810 1779
rect 12935 1748 12963 1820
<< via2 >>
rect 428 6028 578 6174
rect 740 6012 890 6158
rect 492 5068 642 5214
rect 798 5080 948 5226
rect 324 4440 474 4586
rect 360 3594 510 3740
rect 712 3598 862 3744
rect 1158 3598 1308 3744
rect 442 2740 592 2886
rect 792 2748 942 2894
rect 1724 3602 1874 3748
rect 2390 3602 2540 3748
rect 2772 3586 2922 3732
rect 13146 5414 13296 5560
rect 13146 4988 13296 5134
rect 13146 4762 13296 4908
rect 13162 4028 13312 4174
rect 13142 3036 13292 3182
rect 13148 2358 13298 2504
<< metal3 >>
rect 418 6174 590 6184
rect 418 6028 428 6174
rect 578 6028 590 6174
rect 418 6018 590 6028
rect 730 6158 902 6168
rect 730 6012 740 6158
rect 890 6012 902 6158
rect 730 6002 902 6012
rect 13136 5560 13308 5570
rect 13136 5414 13146 5560
rect 13296 5414 13308 5560
rect 13136 5404 13308 5414
rect 788 5226 960 5236
rect 482 5214 654 5224
rect 482 5068 492 5214
rect 642 5068 654 5214
rect 788 5080 798 5226
rect 948 5080 960 5226
rect 788 5070 960 5080
rect 13136 5134 13308 5144
rect 482 5058 654 5068
rect 13136 4988 13146 5134
rect 13296 4988 13308 5134
rect 13136 4978 13308 4988
rect 13136 4908 13308 4918
rect 13136 4762 13146 4908
rect 13296 4762 13308 4908
rect 13136 4752 13308 4762
rect 314 4586 486 4596
rect 314 4440 324 4586
rect 474 4440 486 4586
rect 314 4430 486 4440
rect 13152 4174 13324 4184
rect 13152 4028 13162 4174
rect 13312 4028 13324 4174
rect 13152 4018 13324 4028
rect 350 3740 522 3750
rect 350 3594 360 3740
rect 510 3594 522 3740
rect 350 3584 522 3594
rect 702 3744 874 3754
rect 702 3598 712 3744
rect 862 3598 874 3744
rect 702 3588 874 3598
rect 1148 3744 1320 3754
rect 1148 3598 1158 3744
rect 1308 3598 1320 3744
rect 1148 3588 1320 3598
rect 1714 3748 1886 3758
rect 1714 3602 1724 3748
rect 1874 3602 1886 3748
rect 1714 3592 1886 3602
rect 2380 3748 2552 3758
rect 2380 3602 2390 3748
rect 2540 3602 2552 3748
rect 2380 3592 2552 3602
rect 2762 3732 2934 3742
rect 2762 3586 2772 3732
rect 2922 3586 2934 3732
rect 2762 3576 2934 3586
rect 13132 3182 13304 3192
rect 13132 3036 13142 3182
rect 13292 3036 13304 3182
rect 13132 3026 13304 3036
rect 432 2886 604 2896
rect 432 2740 442 2886
rect 592 2740 604 2886
rect 432 2730 604 2740
rect 782 2894 954 2904
rect 782 2748 792 2894
rect 942 2748 954 2894
rect 782 2738 954 2748
rect 13138 2504 13310 2514
rect 13138 2358 13148 2504
rect 13298 2358 13310 2504
rect 13138 2348 13310 2358
<< via3 >>
rect 428 6028 578 6174
rect 740 6012 890 6158
rect 13146 5414 13296 5560
rect 492 5068 642 5214
rect 798 5080 948 5226
rect 13146 4988 13296 5134
rect 13146 4762 13296 4908
rect 324 4440 474 4586
rect 13162 4028 13312 4174
rect 360 3594 510 3740
rect 712 3598 862 3744
rect 1158 3598 1308 3744
rect 1724 3602 1874 3748
rect 2390 3602 2540 3748
rect 2772 3586 2922 3732
rect 13142 3036 13292 3182
rect 442 2740 592 2886
rect 792 2748 942 2894
rect 13148 2358 13298 2504
<< metal4 >>
rect 290 6174 3896 6228
rect 290 6028 428 6174
rect 578 6158 3896 6174
rect 578 6028 740 6158
rect 290 6012 740 6028
rect 890 6012 3896 6158
rect 290 5226 3896 6012
rect 290 5214 798 5226
rect 290 5068 492 5214
rect 642 5080 798 5214
rect 948 5080 3896 5226
rect 642 5068 3896 5080
rect 290 4586 3896 5068
rect 290 4440 324 4586
rect 474 4440 3896 4586
rect 290 3748 3896 4440
rect 290 3744 1724 3748
rect 290 3740 712 3744
rect 290 3594 360 3740
rect 510 3598 712 3740
rect 862 3598 1158 3744
rect 1308 3602 1724 3744
rect 1874 3602 2390 3748
rect 2540 3732 3896 3748
rect 2540 3602 2772 3732
rect 1308 3598 2772 3602
rect 510 3594 2772 3598
rect 290 3586 2772 3594
rect 2922 3586 3896 3732
rect 290 2894 3896 3586
rect 290 2886 792 2894
rect 290 2740 442 2886
rect 592 2748 792 2886
rect 942 2748 3896 2894
rect 592 2740 3896 2748
rect 290 2258 3896 2740
rect 12894 6202 13396 6204
rect 12894 5560 13444 6202
rect 12894 5414 13146 5560
rect 13296 5414 13444 5560
rect 12894 5134 13444 5414
rect 12894 4988 13146 5134
rect 13296 4988 13444 5134
rect 12894 4908 13444 4988
rect 12894 4762 13146 4908
rect 13296 4762 13444 4908
rect 12894 4174 13444 4762
rect 12894 4028 13162 4174
rect 13312 4028 13444 4174
rect 12894 3182 13444 4028
rect 12894 3036 13142 3182
rect 13292 3036 13444 3182
rect 12894 2504 13444 3036
rect 12894 2358 13148 2504
rect 13298 2358 13444 2504
rect 12894 2246 13444 2358
rect 12972 2244 13444 2246
<< labels >>
flabel metal2 1058 1750 1092 1784 0 FreeSans 480 0 0 0 D[7]
port 9 nsew
flabel metal2 3450 1750 3484 1784 0 FreeSans 480 0 0 0 D[6]
port 10 nsew
flabel metal2 5844 1748 5878 1782 0 FreeSans 480 0 0 0 D[5]
port 12 nsew
flabel metal2 7982 1750 8016 1784 0 FreeSans 480 0 0 0 check[5]
port 14 nsew
flabel metal2 8406 1745 8440 1779 0 FreeSans 480 0 0 0 check[1]
port 15 nsew
flabel metal2 10382 1745 10416 1779 0 FreeSans 480 0 0 0 check[4]
port 16 nsew
flabel metal2 10795 1748 10829 1782 0 FreeSans 480 0 0 0 check[2]
port 17 nsew
flabel metal2 12776 1745 12810 1779 0 FreeSans 480 0 0 0 check[3]
port 18 nsew
flabel metal2 10627 1836 10661 1870 0 FreeSans 480 0 0 0 D[3]
port 20 nsew
flabel metal2 10544 1836 10578 1870 0 FreeSans 480 0 0 0 D[1]
port 21 nsew
flabel metal2 5586 1748 5620 1782 0 FreeSans 480 0 0 0 check[6]
port 11 nsew
flabel metal2 8238 1810 8272 1844 0 FreeSans 480 0 0 0 D[4]
port 22 nsew
flabel metal2 8151 1864 8185 1898 0 FreeSans 480 0 0 0 D[0]
port 24 nsew
flabel metal2 12932 1820 12966 1854 0 FreeSans 480 0 0 0 D[2]
port 19 nsew
flabel metal2 5986 1745 6020 1779 0 FreeSans 480 0 0 0 check[0]
port 13 nsew
flabel metal1 470 4288 504 4322 0 FreeSans 480 0 0 0 reset
port 6 nsew
flabel metal1 468 3414 502 3448 0 FreeSans 480 0 0 0 eob
port 7 nsew
flabel metal1 470 3037 504 3071 0 FreeSans 480 0 0 0 comparator_out
port 8 nsew
flabel metal1 462 5848 496 5882 0 FreeSans 480 0 0 0 clk_sar
port 45 nsew
flabel metal1 464 5782 498 5816 0 FreeSans 480 0 0 0 sel_bit[1]
port 5 nsew
flabel metal1 459 5918 493 5952 0 FreeSans 480 0 0 0 sel_bit[0]
port 4 nsew
flabel metal4 12894 5560 13444 6202 0 FreeSans 320 0 0 0 VSS
port 51 nsew
flabel metal4 290 5226 3896 6012 0 FreeSans 320 0 0 0 VDD
port 53 nsew
flabel locali 3332 3481 3366 3515 0 FreeSans 340 0 0 0 x77.Y
flabel locali 3332 3413 3366 3447 0 FreeSans 340 0 0 0 x77.Y
flabel locali 3240 3413 3274 3447 0 FreeSans 340 0 0 0 x77.A
flabel metal1 3197 3175 3231 3209 0 FreeSans 200 0 0 0 x77.VGND
flabel metal1 3197 3719 3231 3753 0 FreeSans 200 0 0 0 x77.VPWR
rlabel comment 3168 3192 3168 3192 4 x77.inv_1
rlabel metal1 3168 3144 3444 3240 1 x77.VGND
rlabel metal1 3168 3688 3444 3784 1 x77.VPWR
flabel pwell 3197 3175 3231 3209 0 FreeSans 200 0 0 0 x77.VNB
flabel nwell 3197 3719 3231 3753 0 FreeSans 200 0 0 0 x77.VPB
flabel locali 5288 3411 5363 3457 0 FreeSans 400 0 0 0 x75.RESET_B
flabel locali 3455 3175 3489 3209 3 FreeSans 400 0 0 0 x75.VGND
flabel locali 3455 3413 3489 3447 0 FreeSans 400 0 0 0 x75.CLK
flabel locali 3455 3481 3489 3515 0 FreeSans 400 0 0 0 x75.CLK
flabel locali 4191 3345 4225 3379 0 FreeSans 400 0 0 0 x75.SET_B
flabel locali 5753 3277 5787 3311 0 FreeSans 400 0 0 0 x75.Q
flabel locali 5753 3549 5787 3583 0 FreeSans 400 0 0 0 x75.Q
flabel locali 5753 3617 5787 3651 0 FreeSans 400 0 0 0 x75.Q
flabel locali 3455 3719 3489 3753 3 FreeSans 400 0 0 0 x75.VPWR
flabel locali 3823 3413 3857 3447 0 FreeSans 200 0 0 0 x75.D
flabel locali 3823 3481 3857 3515 0 FreeSans 200 0 0 0 x75.D
flabel locali 5473 3617 5507 3651 0 FreeSans 400 0 0 0 x75.Q_N
flabel locali 5473 3549 5507 3583 0 FreeSans 400 0 0 0 x75.Q_N
flabel locali 5473 3277 5507 3311 0 FreeSans 400 0 0 0 x75.Q_N
flabel metal1 3455 3175 3489 3209 0 FreeSans 200 0 0 0 x75.VGND
flabel metal1 3455 3719 3489 3753 0 FreeSans 200 0 0 0 x75.VPWR
flabel nwell 3455 3719 3489 3753 3 FreeSans 400 0 0 0 x75.VPB
flabel nwell 3472 3736 3472 3736 0 FreeSans 200 0 0 0 x75.VPB
flabel pwell 3455 3175 3489 3209 3 FreeSans 400 0 0 0 x75.VNB
flabel pwell 3472 3192 3472 3192 0 FreeSans 200 0 0 0 x75.VNB
rlabel comment 3425 3192 3425 3192 4 x75.dfbbp_1
rlabel locali 4917 3339 4992 3405 1 x75.SET_B
rlabel metal1 4915 3376 4973 3385 1 x75.SET_B
rlabel metal1 4915 3339 4973 3348 1 x75.SET_B
rlabel metal1 4179 3376 4237 3385 1 x75.SET_B
rlabel metal1 4179 3348 4973 3376 1 x75.SET_B
rlabel metal1 4179 3339 4237 3348 1 x75.SET_B
rlabel metal1 3425 3144 5817 3240 1 x75.VGND
rlabel metal1 3425 3688 5817 3784 1 x75.VPWR
flabel locali 7680 3411 7755 3457 0 FreeSans 400 0 0 0 x72.RESET_B
flabel locali 5847 3175 5881 3209 3 FreeSans 400 0 0 0 x72.VGND
flabel locali 5847 3413 5881 3447 0 FreeSans 400 0 0 0 x72.CLK
flabel locali 5847 3481 5881 3515 0 FreeSans 400 0 0 0 x72.CLK
flabel locali 6583 3345 6617 3379 0 FreeSans 400 0 0 0 x72.SET_B
flabel locali 8145 3277 8179 3311 0 FreeSans 400 0 0 0 x72.Q
flabel locali 8145 3549 8179 3583 0 FreeSans 400 0 0 0 x72.Q
flabel locali 8145 3617 8179 3651 0 FreeSans 400 0 0 0 x72.Q
flabel locali 5847 3719 5881 3753 3 FreeSans 400 0 0 0 x72.VPWR
flabel locali 6215 3413 6249 3447 0 FreeSans 200 0 0 0 x72.D
flabel locali 6215 3481 6249 3515 0 FreeSans 200 0 0 0 x72.D
flabel locali 7865 3617 7899 3651 0 FreeSans 400 0 0 0 x72.Q_N
flabel locali 7865 3549 7899 3583 0 FreeSans 400 0 0 0 x72.Q_N
flabel locali 7865 3277 7899 3311 0 FreeSans 400 0 0 0 x72.Q_N
flabel metal1 5847 3175 5881 3209 0 FreeSans 200 0 0 0 x72.VGND
flabel metal1 5847 3719 5881 3753 0 FreeSans 200 0 0 0 x72.VPWR
flabel nwell 5847 3719 5881 3753 3 FreeSans 400 0 0 0 x72.VPB
flabel nwell 5864 3736 5864 3736 0 FreeSans 200 0 0 0 x72.VPB
flabel pwell 5847 3175 5881 3209 3 FreeSans 400 0 0 0 x72.VNB
flabel pwell 5864 3192 5864 3192 0 FreeSans 200 0 0 0 x72.VNB
rlabel comment 5817 3192 5817 3192 4 x72.dfbbp_1
rlabel locali 7309 3339 7384 3405 1 x72.SET_B
rlabel metal1 7307 3376 7365 3385 1 x72.SET_B
rlabel metal1 7307 3339 7365 3348 1 x72.SET_B
rlabel metal1 6571 3376 6629 3385 1 x72.SET_B
rlabel metal1 6571 3348 7365 3376 1 x72.SET_B
rlabel metal1 6571 3339 6629 3348 1 x72.SET_B
rlabel metal1 5817 3144 8209 3240 1 x72.VGND
rlabel metal1 5817 3688 8209 3784 1 x72.VPWR
flabel locali 10072 3411 10147 3457 0 FreeSans 400 0 0 0 x69.RESET_B
flabel locali 8239 3175 8273 3209 3 FreeSans 400 0 0 0 x69.VGND
flabel locali 8239 3413 8273 3447 0 FreeSans 400 0 0 0 x69.CLK
flabel locali 8239 3481 8273 3515 0 FreeSans 400 0 0 0 x69.CLK
flabel locali 8975 3345 9009 3379 0 FreeSans 400 0 0 0 x69.SET_B
flabel locali 10537 3277 10571 3311 0 FreeSans 400 0 0 0 x69.Q
flabel locali 10537 3549 10571 3583 0 FreeSans 400 0 0 0 x69.Q
flabel locali 10537 3617 10571 3651 0 FreeSans 400 0 0 0 x69.Q
flabel locali 8239 3719 8273 3753 3 FreeSans 400 0 0 0 x69.VPWR
flabel locali 8607 3413 8641 3447 0 FreeSans 200 0 0 0 x69.D
flabel locali 8607 3481 8641 3515 0 FreeSans 200 0 0 0 x69.D
flabel locali 10257 3617 10291 3651 0 FreeSans 400 0 0 0 x69.Q_N
flabel locali 10257 3549 10291 3583 0 FreeSans 400 0 0 0 x69.Q_N
flabel locali 10257 3277 10291 3311 0 FreeSans 400 0 0 0 x69.Q_N
flabel metal1 8239 3175 8273 3209 0 FreeSans 200 0 0 0 x69.VGND
flabel metal1 8239 3719 8273 3753 0 FreeSans 200 0 0 0 x69.VPWR
flabel nwell 8239 3719 8273 3753 3 FreeSans 400 0 0 0 x69.VPB
flabel nwell 8256 3736 8256 3736 0 FreeSans 200 0 0 0 x69.VPB
flabel pwell 8239 3175 8273 3209 3 FreeSans 400 0 0 0 x69.VNB
flabel pwell 8256 3192 8256 3192 0 FreeSans 200 0 0 0 x69.VNB
rlabel comment 8209 3192 8209 3192 4 x69.dfbbp_1
rlabel locali 9701 3339 9776 3405 1 x69.SET_B
rlabel metal1 9699 3376 9757 3385 1 x69.SET_B
rlabel metal1 9699 3339 9757 3348 1 x69.SET_B
rlabel metal1 8963 3376 9021 3385 1 x69.SET_B
rlabel metal1 8963 3348 9757 3376 1 x69.SET_B
rlabel metal1 8963 3339 9021 3348 1 x69.SET_B
rlabel metal1 8209 3144 10601 3240 1 x69.VGND
rlabel metal1 8209 3688 10601 3784 1 x69.VPWR
flabel locali 12464 3411 12539 3457 0 FreeSans 400 0 0 0 x66.RESET_B
flabel locali 10631 3175 10665 3209 3 FreeSans 400 0 0 0 x66.VGND
flabel locali 10631 3413 10665 3447 0 FreeSans 400 0 0 0 x66.CLK
flabel locali 10631 3481 10665 3515 0 FreeSans 400 0 0 0 x66.CLK
flabel locali 11367 3345 11401 3379 0 FreeSans 400 0 0 0 x66.SET_B
flabel locali 12929 3277 12963 3311 0 FreeSans 400 0 0 0 x66.Q
flabel locali 12929 3549 12963 3583 0 FreeSans 400 0 0 0 x66.Q
flabel locali 12929 3617 12963 3651 0 FreeSans 400 0 0 0 x66.Q
flabel locali 10631 3719 10665 3753 3 FreeSans 400 0 0 0 x66.VPWR
flabel locali 10999 3413 11033 3447 0 FreeSans 200 0 0 0 x66.D
flabel locali 10999 3481 11033 3515 0 FreeSans 200 0 0 0 x66.D
flabel locali 12649 3617 12683 3651 0 FreeSans 400 0 0 0 x66.Q_N
flabel locali 12649 3549 12683 3583 0 FreeSans 400 0 0 0 x66.Q_N
flabel locali 12649 3277 12683 3311 0 FreeSans 400 0 0 0 x66.Q_N
flabel metal1 10631 3175 10665 3209 0 FreeSans 200 0 0 0 x66.VGND
flabel metal1 10631 3719 10665 3753 0 FreeSans 200 0 0 0 x66.VPWR
flabel nwell 10631 3719 10665 3753 3 FreeSans 400 0 0 0 x66.VPB
flabel nwell 10648 3736 10648 3736 0 FreeSans 200 0 0 0 x66.VPB
flabel pwell 10631 3175 10665 3209 3 FreeSans 400 0 0 0 x66.VNB
flabel pwell 10648 3192 10648 3192 0 FreeSans 200 0 0 0 x66.VNB
rlabel comment 10601 3192 10601 3192 4 x66.dfbbp_1
rlabel locali 12093 3339 12168 3405 1 x66.SET_B
rlabel metal1 12091 3376 12149 3385 1 x66.SET_B
rlabel metal1 12091 3339 12149 3348 1 x66.SET_B
rlabel metal1 11355 3376 11413 3385 1 x66.SET_B
rlabel metal1 11355 3348 12149 3376 1 x66.SET_B
rlabel metal1 11355 3339 11413 3348 1 x66.SET_B
rlabel metal1 10601 3144 12993 3240 1 x66.VGND
rlabel metal1 10601 3688 12993 3784 1 x66.VPWR
flabel locali 11055 2538 11130 2584 0 FreeSans 400 0 0 0 x63.RESET_B
flabel locali 12929 2302 12963 2336 7 FreeSans 400 0 0 0 x63.VGND
flabel locali 12929 2540 12963 2574 0 FreeSans 400 0 0 0 x63.CLK
flabel locali 12929 2608 12963 2642 0 FreeSans 400 0 0 0 x63.CLK
flabel locali 12193 2472 12227 2506 0 FreeSans 400 0 0 0 x63.SET_B
flabel locali 10631 2404 10665 2438 0 FreeSans 400 0 0 0 x63.Q
flabel locali 10631 2676 10665 2710 0 FreeSans 400 0 0 0 x63.Q
flabel locali 10631 2744 10665 2778 0 FreeSans 400 0 0 0 x63.Q
flabel locali 12929 2846 12963 2880 7 FreeSans 400 0 0 0 x63.VPWR
flabel locali 12561 2540 12595 2574 0 FreeSans 200 0 0 0 x63.D
flabel locali 12561 2608 12595 2642 0 FreeSans 200 0 0 0 x63.D
flabel locali 10911 2744 10945 2778 0 FreeSans 400 0 0 0 x63.Q_N
flabel locali 10911 2676 10945 2710 0 FreeSans 400 0 0 0 x63.Q_N
flabel locali 10911 2404 10945 2438 0 FreeSans 400 0 0 0 x63.Q_N
flabel metal1 12929 2302 12963 2336 0 FreeSans 200 0 0 0 x63.VGND
flabel metal1 12929 2846 12963 2880 0 FreeSans 200 0 0 0 x63.VPWR
flabel nwell 12929 2846 12963 2880 7 FreeSans 400 0 0 0 x63.VPB
flabel nwell 12946 2863 12946 2863 0 FreeSans 200 0 0 0 x63.VPB
flabel pwell 12929 2302 12963 2336 7 FreeSans 400 0 0 0 x63.VNB
flabel pwell 12946 2319 12946 2319 0 FreeSans 200 0 0 0 x63.VNB
rlabel comment 12993 2319 12993 2319 6 x63.dfbbp_1
rlabel locali 11426 2466 11501 2532 1 x63.SET_B
rlabel metal1 11445 2503 11503 2512 1 x63.SET_B
rlabel metal1 11445 2466 11503 2475 1 x63.SET_B
rlabel metal1 12181 2503 12239 2512 1 x63.SET_B
rlabel metal1 11445 2475 12239 2503 1 x63.SET_B
rlabel metal1 12181 2466 12239 2475 1 x63.SET_B
rlabel metal1 10601 2271 12993 2367 1 x63.VGND
rlabel metal1 10601 2815 12993 2911 1 x63.VPWR
flabel locali 8663 2538 8738 2584 0 FreeSans 400 0 0 0 x60.RESET_B
flabel locali 10537 2302 10571 2336 7 FreeSans 400 0 0 0 x60.VGND
flabel locali 10537 2540 10571 2574 0 FreeSans 400 0 0 0 x60.CLK
flabel locali 10537 2608 10571 2642 0 FreeSans 400 0 0 0 x60.CLK
flabel locali 9801 2472 9835 2506 0 FreeSans 400 0 0 0 x60.SET_B
flabel locali 8239 2404 8273 2438 0 FreeSans 400 0 0 0 x60.Q
flabel locali 8239 2676 8273 2710 0 FreeSans 400 0 0 0 x60.Q
flabel locali 8239 2744 8273 2778 0 FreeSans 400 0 0 0 x60.Q
flabel locali 10537 2846 10571 2880 7 FreeSans 400 0 0 0 x60.VPWR
flabel locali 10169 2540 10203 2574 0 FreeSans 200 0 0 0 x60.D
flabel locali 10169 2608 10203 2642 0 FreeSans 200 0 0 0 x60.D
flabel locali 8519 2744 8553 2778 0 FreeSans 400 0 0 0 x60.Q_N
flabel locali 8519 2676 8553 2710 0 FreeSans 400 0 0 0 x60.Q_N
flabel locali 8519 2404 8553 2438 0 FreeSans 400 0 0 0 x60.Q_N
flabel metal1 10537 2302 10571 2336 0 FreeSans 200 0 0 0 x60.VGND
flabel metal1 10537 2846 10571 2880 0 FreeSans 200 0 0 0 x60.VPWR
flabel nwell 10537 2846 10571 2880 7 FreeSans 400 0 0 0 x60.VPB
flabel nwell 10554 2863 10554 2863 0 FreeSans 200 0 0 0 x60.VPB
flabel pwell 10537 2302 10571 2336 7 FreeSans 400 0 0 0 x60.VNB
flabel pwell 10554 2319 10554 2319 0 FreeSans 200 0 0 0 x60.VNB
rlabel comment 10601 2319 10601 2319 6 x60.dfbbp_1
rlabel locali 9034 2466 9109 2532 1 x60.SET_B
rlabel metal1 9053 2503 9111 2512 1 x60.SET_B
rlabel metal1 9053 2466 9111 2475 1 x60.SET_B
rlabel metal1 9789 2503 9847 2512 1 x60.SET_B
rlabel metal1 9053 2475 9847 2503 1 x60.SET_B
rlabel metal1 9789 2466 9847 2475 1 x60.SET_B
rlabel metal1 8209 2271 10601 2367 1 x60.VGND
rlabel metal1 8209 2815 10601 2911 1 x60.VPWR
flabel locali 6271 2538 6346 2584 0 FreeSans 400 0 0 0 x57.RESET_B
flabel locali 8145 2302 8179 2336 7 FreeSans 400 0 0 0 x57.VGND
flabel locali 8145 2540 8179 2574 0 FreeSans 400 0 0 0 x57.CLK
flabel locali 8145 2608 8179 2642 0 FreeSans 400 0 0 0 x57.CLK
flabel locali 7409 2472 7443 2506 0 FreeSans 400 0 0 0 x57.SET_B
flabel locali 5847 2404 5881 2438 0 FreeSans 400 0 0 0 x57.Q
flabel locali 5847 2676 5881 2710 0 FreeSans 400 0 0 0 x57.Q
flabel locali 5847 2744 5881 2778 0 FreeSans 400 0 0 0 x57.Q
flabel locali 8145 2846 8179 2880 7 FreeSans 400 0 0 0 x57.VPWR
flabel locali 7777 2540 7811 2574 0 FreeSans 200 0 0 0 x57.D
flabel locali 7777 2608 7811 2642 0 FreeSans 200 0 0 0 x57.D
flabel locali 6127 2744 6161 2778 0 FreeSans 400 0 0 0 x57.Q_N
flabel locali 6127 2676 6161 2710 0 FreeSans 400 0 0 0 x57.Q_N
flabel locali 6127 2404 6161 2438 0 FreeSans 400 0 0 0 x57.Q_N
flabel metal1 8145 2302 8179 2336 0 FreeSans 200 0 0 0 x57.VGND
flabel metal1 8145 2846 8179 2880 0 FreeSans 200 0 0 0 x57.VPWR
flabel nwell 8145 2846 8179 2880 7 FreeSans 400 0 0 0 x57.VPB
flabel nwell 8162 2863 8162 2863 0 FreeSans 200 0 0 0 x57.VPB
flabel pwell 8145 2302 8179 2336 7 FreeSans 400 0 0 0 x57.VNB
flabel pwell 8162 2319 8162 2319 0 FreeSans 200 0 0 0 x57.VNB
rlabel comment 8209 2319 8209 2319 6 x57.dfbbp_1
rlabel locali 6642 2466 6717 2532 1 x57.SET_B
rlabel metal1 6661 2503 6719 2512 1 x57.SET_B
rlabel metal1 6661 2466 6719 2475 1 x57.SET_B
rlabel metal1 7397 2503 7455 2512 1 x57.SET_B
rlabel metal1 6661 2475 7455 2503 1 x57.SET_B
rlabel metal1 7397 2466 7455 2475 1 x57.SET_B
rlabel metal1 5817 2271 8209 2367 1 x57.VGND
rlabel metal1 5817 2815 8209 2911 1 x57.VPWR
flabel locali 3879 2538 3954 2584 0 FreeSans 400 0 0 0 x54.RESET_B
flabel locali 5753 2302 5787 2336 7 FreeSans 400 0 0 0 x54.VGND
flabel locali 5753 2540 5787 2574 0 FreeSans 400 0 0 0 x54.CLK
flabel locali 5753 2608 5787 2642 0 FreeSans 400 0 0 0 x54.CLK
flabel locali 5017 2472 5051 2506 0 FreeSans 400 0 0 0 x54.SET_B
flabel locali 3455 2404 3489 2438 0 FreeSans 400 0 0 0 x54.Q
flabel locali 3455 2676 3489 2710 0 FreeSans 400 0 0 0 x54.Q
flabel locali 3455 2744 3489 2778 0 FreeSans 400 0 0 0 x54.Q
flabel locali 5753 2846 5787 2880 7 FreeSans 400 0 0 0 x54.VPWR
flabel locali 5385 2540 5419 2574 0 FreeSans 200 0 0 0 x54.D
flabel locali 5385 2608 5419 2642 0 FreeSans 200 0 0 0 x54.D
flabel locali 3735 2744 3769 2778 0 FreeSans 400 0 0 0 x54.Q_N
flabel locali 3735 2676 3769 2710 0 FreeSans 400 0 0 0 x54.Q_N
flabel locali 3735 2404 3769 2438 0 FreeSans 400 0 0 0 x54.Q_N
flabel metal1 5753 2302 5787 2336 0 FreeSans 200 0 0 0 x54.VGND
flabel metal1 5753 2846 5787 2880 0 FreeSans 200 0 0 0 x54.VPWR
flabel nwell 5753 2846 5787 2880 7 FreeSans 400 0 0 0 x54.VPB
flabel nwell 5770 2863 5770 2863 0 FreeSans 200 0 0 0 x54.VPB
flabel pwell 5753 2302 5787 2336 7 FreeSans 400 0 0 0 x54.VNB
flabel pwell 5770 2319 5770 2319 0 FreeSans 200 0 0 0 x54.VNB
rlabel comment 5817 2319 5817 2319 6 x54.dfbbp_1
rlabel locali 4250 2466 4325 2532 1 x54.SET_B
rlabel metal1 4269 2503 4327 2512 1 x54.SET_B
rlabel metal1 4269 2466 4327 2475 1 x54.SET_B
rlabel metal1 5005 2503 5063 2512 1 x54.SET_B
rlabel metal1 4269 2475 5063 2503 1 x54.SET_B
rlabel metal1 5005 2466 5063 2475 1 x54.SET_B
rlabel metal1 3425 2271 5817 2367 1 x54.VGND
rlabel metal1 3425 2815 5817 2911 1 x54.VPWR
flabel locali 1487 2538 1562 2584 0 FreeSans 400 0 0 0 x51.RESET_B
flabel locali 3361 2302 3395 2336 7 FreeSans 400 0 0 0 x51.VGND
flabel locali 3361 2540 3395 2574 0 FreeSans 400 0 0 0 x51.CLK
flabel locali 3361 2608 3395 2642 0 FreeSans 400 0 0 0 x51.CLK
flabel locali 2625 2472 2659 2506 0 FreeSans 400 0 0 0 x51.SET_B
flabel locali 1063 2404 1097 2438 0 FreeSans 400 0 0 0 x51.Q
flabel locali 1063 2676 1097 2710 0 FreeSans 400 0 0 0 x51.Q
flabel locali 1063 2744 1097 2778 0 FreeSans 400 0 0 0 x51.Q
flabel locali 3361 2846 3395 2880 7 FreeSans 400 0 0 0 x51.VPWR
flabel locali 2993 2540 3027 2574 0 FreeSans 200 0 0 0 x51.D
flabel locali 2993 2608 3027 2642 0 FreeSans 200 0 0 0 x51.D
flabel locali 1343 2744 1377 2778 0 FreeSans 400 0 0 0 x51.Q_N
flabel locali 1343 2676 1377 2710 0 FreeSans 400 0 0 0 x51.Q_N
flabel locali 1343 2404 1377 2438 0 FreeSans 400 0 0 0 x51.Q_N
flabel metal1 3361 2302 3395 2336 0 FreeSans 200 0 0 0 x51.VGND
flabel metal1 3361 2846 3395 2880 0 FreeSans 200 0 0 0 x51.VPWR
flabel nwell 3361 2846 3395 2880 7 FreeSans 400 0 0 0 x51.VPB
flabel nwell 3378 2863 3378 2863 0 FreeSans 200 0 0 0 x51.VPB
flabel pwell 3361 2302 3395 2336 7 FreeSans 400 0 0 0 x51.VNB
flabel pwell 3378 2319 3378 2319 0 FreeSans 200 0 0 0 x51.VNB
rlabel comment 3425 2319 3425 2319 6 x51.dfbbp_1
rlabel locali 1858 2466 1933 2532 1 x51.SET_B
rlabel metal1 1877 2503 1935 2512 1 x51.SET_B
rlabel metal1 1877 2466 1935 2475 1 x51.SET_B
rlabel metal1 2613 2503 2671 2512 1 x51.SET_B
rlabel metal1 1877 2475 2671 2503 1 x51.SET_B
rlabel metal1 2613 2466 2671 2475 1 x51.SET_B
rlabel metal1 1033 2271 3425 2367 1 x51.VGND
rlabel metal1 1033 2815 3425 2911 1 x51.VPWR
flabel locali 3880 4284 3955 4330 0 FreeSans 400 0 0 0 x48.RESET_B
flabel locali 5754 4048 5788 4082 7 FreeSans 400 0 0 0 x48.VGND
flabel locali 5754 4286 5788 4320 0 FreeSans 400 0 0 0 x48.CLK
flabel locali 5754 4354 5788 4388 0 FreeSans 400 0 0 0 x48.CLK
flabel locali 5018 4218 5052 4252 0 FreeSans 400 0 0 0 x48.SET_B
flabel locali 3456 4150 3490 4184 0 FreeSans 400 0 0 0 x48.Q
flabel locali 3456 4422 3490 4456 0 FreeSans 400 0 0 0 x48.Q
flabel locali 3456 4490 3490 4524 0 FreeSans 400 0 0 0 x48.Q
flabel locali 5754 4592 5788 4626 7 FreeSans 400 0 0 0 x48.VPWR
flabel locali 5386 4286 5420 4320 0 FreeSans 200 0 0 0 x48.D
flabel locali 5386 4354 5420 4388 0 FreeSans 200 0 0 0 x48.D
flabel locali 3736 4490 3770 4524 0 FreeSans 400 0 0 0 x48.Q_N
flabel locali 3736 4422 3770 4456 0 FreeSans 400 0 0 0 x48.Q_N
flabel locali 3736 4150 3770 4184 0 FreeSans 400 0 0 0 x48.Q_N
flabel metal1 5754 4048 5788 4082 0 FreeSans 200 0 0 0 x48.VGND
flabel metal1 5754 4592 5788 4626 0 FreeSans 200 0 0 0 x48.VPWR
flabel nwell 5754 4592 5788 4626 7 FreeSans 400 0 0 0 x48.VPB
flabel nwell 5771 4609 5771 4609 0 FreeSans 200 0 0 0 x48.VPB
flabel pwell 5754 4048 5788 4082 7 FreeSans 400 0 0 0 x48.VNB
flabel pwell 5771 4065 5771 4065 0 FreeSans 200 0 0 0 x48.VNB
rlabel comment 5818 4065 5818 4065 6 x48.dfbbp_1
rlabel locali 4251 4212 4326 4278 1 x48.SET_B
rlabel metal1 4270 4249 4328 4258 1 x48.SET_B
rlabel metal1 4270 4212 4328 4221 1 x48.SET_B
rlabel metal1 5006 4249 5064 4258 1 x48.SET_B
rlabel metal1 4270 4221 5064 4249 1 x48.SET_B
rlabel metal1 5006 4212 5064 4221 1 x48.SET_B
rlabel metal1 3426 4017 5818 4113 1 x48.VGND
rlabel metal1 3426 4561 5818 4657 1 x48.VPWR
flabel locali 6272 4284 6347 4330 0 FreeSans 400 0 0 0 x45.RESET_B
flabel locali 8146 4048 8180 4082 7 FreeSans 400 0 0 0 x45.VGND
flabel locali 8146 4286 8180 4320 0 FreeSans 400 0 0 0 x45.CLK
flabel locali 8146 4354 8180 4388 0 FreeSans 400 0 0 0 x45.CLK
flabel locali 7410 4218 7444 4252 0 FreeSans 400 0 0 0 x45.SET_B
flabel locali 5848 4150 5882 4184 0 FreeSans 400 0 0 0 x45.Q
flabel locali 5848 4422 5882 4456 0 FreeSans 400 0 0 0 x45.Q
flabel locali 5848 4490 5882 4524 0 FreeSans 400 0 0 0 x45.Q
flabel locali 8146 4592 8180 4626 7 FreeSans 400 0 0 0 x45.VPWR
flabel locali 7778 4286 7812 4320 0 FreeSans 200 0 0 0 x45.D
flabel locali 7778 4354 7812 4388 0 FreeSans 200 0 0 0 x45.D
flabel locali 6128 4490 6162 4524 0 FreeSans 400 0 0 0 x45.Q_N
flabel locali 6128 4422 6162 4456 0 FreeSans 400 0 0 0 x45.Q_N
flabel locali 6128 4150 6162 4184 0 FreeSans 400 0 0 0 x45.Q_N
flabel metal1 8146 4048 8180 4082 0 FreeSans 200 0 0 0 x45.VGND
flabel metal1 8146 4592 8180 4626 0 FreeSans 200 0 0 0 x45.VPWR
flabel nwell 8146 4592 8180 4626 7 FreeSans 400 0 0 0 x45.VPB
flabel nwell 8163 4609 8163 4609 0 FreeSans 200 0 0 0 x45.VPB
flabel pwell 8146 4048 8180 4082 7 FreeSans 400 0 0 0 x45.VNB
flabel pwell 8163 4065 8163 4065 0 FreeSans 200 0 0 0 x45.VNB
rlabel comment 8210 4065 8210 4065 6 x45.dfbbp_1
rlabel locali 6643 4212 6718 4278 1 x45.SET_B
rlabel metal1 6662 4249 6720 4258 1 x45.SET_B
rlabel metal1 6662 4212 6720 4221 1 x45.SET_B
rlabel metal1 7398 4249 7456 4258 1 x45.SET_B
rlabel metal1 6662 4221 7456 4249 1 x45.SET_B
rlabel metal1 7398 4212 7456 4221 1 x45.SET_B
rlabel metal1 5818 4017 8210 4113 1 x45.VGND
rlabel metal1 5818 4561 8210 4657 1 x45.VPWR
flabel locali 8664 4284 8739 4330 0 FreeSans 400 0 0 0 x42.RESET_B
flabel locali 10538 4048 10572 4082 7 FreeSans 400 0 0 0 x42.VGND
flabel locali 10538 4286 10572 4320 0 FreeSans 400 0 0 0 x42.CLK
flabel locali 10538 4354 10572 4388 0 FreeSans 400 0 0 0 x42.CLK
flabel locali 9802 4218 9836 4252 0 FreeSans 400 0 0 0 x42.SET_B
flabel locali 8240 4150 8274 4184 0 FreeSans 400 0 0 0 x42.Q
flabel locali 8240 4422 8274 4456 0 FreeSans 400 0 0 0 x42.Q
flabel locali 8240 4490 8274 4524 0 FreeSans 400 0 0 0 x42.Q
flabel locali 10538 4592 10572 4626 7 FreeSans 400 0 0 0 x42.VPWR
flabel locali 10170 4286 10204 4320 0 FreeSans 200 0 0 0 x42.D
flabel locali 10170 4354 10204 4388 0 FreeSans 200 0 0 0 x42.D
flabel locali 8520 4490 8554 4524 0 FreeSans 400 0 0 0 x42.Q_N
flabel locali 8520 4422 8554 4456 0 FreeSans 400 0 0 0 x42.Q_N
flabel locali 8520 4150 8554 4184 0 FreeSans 400 0 0 0 x42.Q_N
flabel metal1 10538 4048 10572 4082 0 FreeSans 200 0 0 0 x42.VGND
flabel metal1 10538 4592 10572 4626 0 FreeSans 200 0 0 0 x42.VPWR
flabel nwell 10538 4592 10572 4626 7 FreeSans 400 0 0 0 x42.VPB
flabel nwell 10555 4609 10555 4609 0 FreeSans 200 0 0 0 x42.VPB
flabel pwell 10538 4048 10572 4082 7 FreeSans 400 0 0 0 x42.VNB
flabel pwell 10555 4065 10555 4065 0 FreeSans 200 0 0 0 x42.VNB
rlabel comment 10602 4065 10602 4065 6 x42.dfbbp_1
rlabel locali 9035 4212 9110 4278 1 x42.SET_B
rlabel metal1 9054 4249 9112 4258 1 x42.SET_B
rlabel metal1 9054 4212 9112 4221 1 x42.SET_B
rlabel metal1 9790 4249 9848 4258 1 x42.SET_B
rlabel metal1 9054 4221 9848 4249 1 x42.SET_B
rlabel metal1 9790 4212 9848 4221 1 x42.SET_B
rlabel metal1 8210 4017 10602 4113 1 x42.VGND
rlabel metal1 8210 4561 10602 4657 1 x42.VPWR
flabel locali 11056 4284 11131 4330 0 FreeSans 400 0 0 0 x39.RESET_B
flabel locali 12930 4048 12964 4082 7 FreeSans 400 0 0 0 x39.VGND
flabel locali 12930 4286 12964 4320 0 FreeSans 400 0 0 0 x39.CLK
flabel locali 12930 4354 12964 4388 0 FreeSans 400 0 0 0 x39.CLK
flabel locali 12194 4218 12228 4252 0 FreeSans 400 0 0 0 x39.SET_B
flabel locali 10632 4150 10666 4184 0 FreeSans 400 0 0 0 x39.Q
flabel locali 10632 4422 10666 4456 0 FreeSans 400 0 0 0 x39.Q
flabel locali 10632 4490 10666 4524 0 FreeSans 400 0 0 0 x39.Q
flabel locali 12930 4592 12964 4626 7 FreeSans 400 0 0 0 x39.VPWR
flabel locali 12562 4286 12596 4320 0 FreeSans 200 0 0 0 x39.D
flabel locali 12562 4354 12596 4388 0 FreeSans 200 0 0 0 x39.D
flabel locali 10912 4490 10946 4524 0 FreeSans 400 0 0 0 x39.Q_N
flabel locali 10912 4422 10946 4456 0 FreeSans 400 0 0 0 x39.Q_N
flabel locali 10912 4150 10946 4184 0 FreeSans 400 0 0 0 x39.Q_N
flabel metal1 12930 4048 12964 4082 0 FreeSans 200 0 0 0 x39.VGND
flabel metal1 12930 4592 12964 4626 0 FreeSans 200 0 0 0 x39.VPWR
flabel nwell 12930 4592 12964 4626 7 FreeSans 400 0 0 0 x39.VPB
flabel nwell 12947 4609 12947 4609 0 FreeSans 200 0 0 0 x39.VPB
flabel pwell 12930 4048 12964 4082 7 FreeSans 400 0 0 0 x39.VNB
flabel pwell 12947 4065 12947 4065 0 FreeSans 200 0 0 0 x39.VNB
rlabel comment 12994 4065 12994 4065 6 x39.dfbbp_1
rlabel locali 11427 4212 11502 4278 1 x39.SET_B
rlabel metal1 11446 4249 11504 4258 1 x39.SET_B
rlabel metal1 11446 4212 11504 4221 1 x39.SET_B
rlabel metal1 12182 4249 12240 4258 1 x39.SET_B
rlabel metal1 11446 4221 12240 4249 1 x39.SET_B
rlabel metal1 12182 4212 12240 4221 1 x39.SET_B
rlabel metal1 10602 4017 12994 4113 1 x39.VGND
rlabel metal1 10602 4561 12994 4657 1 x39.VPWR
flabel locali 12465 4973 12540 5019 0 FreeSans 400 0 0 0 x36.RESET_B
flabel locali 10632 4737 10666 4771 3 FreeSans 400 0 0 0 x36.VGND
flabel locali 10632 4975 10666 5009 0 FreeSans 400 0 0 0 x36.CLK
flabel locali 10632 5043 10666 5077 0 FreeSans 400 0 0 0 x36.CLK
flabel locali 11368 4907 11402 4941 0 FreeSans 400 0 0 0 x36.SET_B
flabel locali 12930 4839 12964 4873 0 FreeSans 400 0 0 0 x36.Q
flabel locali 12930 5111 12964 5145 0 FreeSans 400 0 0 0 x36.Q
flabel locali 12930 5179 12964 5213 0 FreeSans 400 0 0 0 x36.Q
flabel locali 10632 5281 10666 5315 3 FreeSans 400 0 0 0 x36.VPWR
flabel locali 11000 4975 11034 5009 0 FreeSans 200 0 0 0 x36.D
flabel locali 11000 5043 11034 5077 0 FreeSans 200 0 0 0 x36.D
flabel locali 12650 5179 12684 5213 0 FreeSans 400 0 0 0 x36.Q_N
flabel locali 12650 5111 12684 5145 0 FreeSans 400 0 0 0 x36.Q_N
flabel locali 12650 4839 12684 4873 0 FreeSans 400 0 0 0 x36.Q_N
flabel metal1 10632 4737 10666 4771 0 FreeSans 200 0 0 0 x36.VGND
flabel metal1 10632 5281 10666 5315 0 FreeSans 200 0 0 0 x36.VPWR
flabel nwell 10632 5281 10666 5315 3 FreeSans 400 0 0 0 x36.VPB
flabel nwell 10649 5298 10649 5298 0 FreeSans 200 0 0 0 x36.VPB
flabel pwell 10632 4737 10666 4771 3 FreeSans 400 0 0 0 x36.VNB
flabel pwell 10649 4754 10649 4754 0 FreeSans 200 0 0 0 x36.VNB
rlabel comment 10602 4754 10602 4754 4 x36.dfbbp_1
rlabel locali 12094 4901 12169 4967 1 x36.SET_B
rlabel metal1 12092 4938 12150 4947 1 x36.SET_B
rlabel metal1 12092 4901 12150 4910 1 x36.SET_B
rlabel metal1 11356 4938 11414 4947 1 x36.SET_B
rlabel metal1 11356 4910 12150 4938 1 x36.SET_B
rlabel metal1 11356 4901 11414 4910 1 x36.SET_B
rlabel metal1 10602 4706 12994 4802 1 x36.VGND
rlabel metal1 10602 5250 12994 5346 1 x36.VPWR
flabel locali 10073 4973 10148 5019 0 FreeSans 400 0 0 0 x33.RESET_B
flabel locali 8240 4737 8274 4771 3 FreeSans 400 0 0 0 x33.VGND
flabel locali 8240 4975 8274 5009 0 FreeSans 400 0 0 0 x33.CLK
flabel locali 8240 5043 8274 5077 0 FreeSans 400 0 0 0 x33.CLK
flabel locali 8976 4907 9010 4941 0 FreeSans 400 0 0 0 x33.SET_B
flabel locali 10538 4839 10572 4873 0 FreeSans 400 0 0 0 x33.Q
flabel locali 10538 5111 10572 5145 0 FreeSans 400 0 0 0 x33.Q
flabel locali 10538 5179 10572 5213 0 FreeSans 400 0 0 0 x33.Q
flabel locali 8240 5281 8274 5315 3 FreeSans 400 0 0 0 x33.VPWR
flabel locali 8608 4975 8642 5009 0 FreeSans 200 0 0 0 x33.D
flabel locali 8608 5043 8642 5077 0 FreeSans 200 0 0 0 x33.D
flabel locali 10258 5179 10292 5213 0 FreeSans 400 0 0 0 x33.Q_N
flabel locali 10258 5111 10292 5145 0 FreeSans 400 0 0 0 x33.Q_N
flabel locali 10258 4839 10292 4873 0 FreeSans 400 0 0 0 x33.Q_N
flabel metal1 8240 4737 8274 4771 0 FreeSans 200 0 0 0 x33.VGND
flabel metal1 8240 5281 8274 5315 0 FreeSans 200 0 0 0 x33.VPWR
flabel nwell 8240 5281 8274 5315 3 FreeSans 400 0 0 0 x33.VPB
flabel nwell 8257 5298 8257 5298 0 FreeSans 200 0 0 0 x33.VPB
flabel pwell 8240 4737 8274 4771 3 FreeSans 400 0 0 0 x33.VNB
flabel pwell 8257 4754 8257 4754 0 FreeSans 200 0 0 0 x33.VNB
rlabel comment 8210 4754 8210 4754 4 x33.dfbbp_1
rlabel locali 9702 4901 9777 4967 1 x33.SET_B
rlabel metal1 9700 4938 9758 4947 1 x33.SET_B
rlabel metal1 9700 4901 9758 4910 1 x33.SET_B
rlabel metal1 8964 4938 9022 4947 1 x33.SET_B
rlabel metal1 8964 4910 9758 4938 1 x33.SET_B
rlabel metal1 8964 4901 9022 4910 1 x33.SET_B
rlabel metal1 8210 4706 10602 4802 1 x33.VGND
rlabel metal1 8210 5250 10602 5346 1 x33.VPWR
flabel locali 7681 4973 7756 5019 0 FreeSans 400 0 0 0 x30.RESET_B
flabel locali 5848 4737 5882 4771 3 FreeSans 400 0 0 0 x30.VGND
flabel locali 5848 4975 5882 5009 0 FreeSans 400 0 0 0 x30.CLK
flabel locali 5848 5043 5882 5077 0 FreeSans 400 0 0 0 x30.CLK
flabel locali 6584 4907 6618 4941 0 FreeSans 400 0 0 0 x30.SET_B
flabel locali 8146 4839 8180 4873 0 FreeSans 400 0 0 0 x30.Q
flabel locali 8146 5111 8180 5145 0 FreeSans 400 0 0 0 x30.Q
flabel locali 8146 5179 8180 5213 0 FreeSans 400 0 0 0 x30.Q
flabel locali 5848 5281 5882 5315 3 FreeSans 400 0 0 0 x30.VPWR
flabel locali 6216 4975 6250 5009 0 FreeSans 200 0 0 0 x30.D
flabel locali 6216 5043 6250 5077 0 FreeSans 200 0 0 0 x30.D
flabel locali 7866 5179 7900 5213 0 FreeSans 400 0 0 0 x30.Q_N
flabel locali 7866 5111 7900 5145 0 FreeSans 400 0 0 0 x30.Q_N
flabel locali 7866 4839 7900 4873 0 FreeSans 400 0 0 0 x30.Q_N
flabel metal1 5848 4737 5882 4771 0 FreeSans 200 0 0 0 x30.VGND
flabel metal1 5848 5281 5882 5315 0 FreeSans 200 0 0 0 x30.VPWR
flabel nwell 5848 5281 5882 5315 3 FreeSans 400 0 0 0 x30.VPB
flabel nwell 5865 5298 5865 5298 0 FreeSans 200 0 0 0 x30.VPB
flabel pwell 5848 4737 5882 4771 3 FreeSans 400 0 0 0 x30.VNB
flabel pwell 5865 4754 5865 4754 0 FreeSans 200 0 0 0 x30.VNB
rlabel comment 5818 4754 5818 4754 4 x30.dfbbp_1
rlabel locali 7310 4901 7385 4967 1 x30.SET_B
rlabel metal1 7308 4938 7366 4947 1 x30.SET_B
rlabel metal1 7308 4901 7366 4910 1 x30.SET_B
rlabel metal1 6572 4938 6630 4947 1 x30.SET_B
rlabel metal1 6572 4910 7366 4938 1 x30.SET_B
rlabel metal1 6572 4901 6630 4910 1 x30.SET_B
rlabel metal1 5818 4706 8210 4802 1 x30.VGND
rlabel metal1 5818 5250 8210 5346 1 x30.VPWR
flabel locali 5289 4973 5364 5019 0 FreeSans 400 0 0 0 x27.RESET_B
flabel locali 3456 4737 3490 4771 3 FreeSans 400 0 0 0 x27.VGND
flabel locali 3456 4975 3490 5009 0 FreeSans 400 0 0 0 x27.CLK
flabel locali 3456 5043 3490 5077 0 FreeSans 400 0 0 0 x27.CLK
flabel locali 4192 4907 4226 4941 0 FreeSans 400 0 0 0 x27.SET_B
flabel locali 5754 4839 5788 4873 0 FreeSans 400 0 0 0 x27.Q
flabel locali 5754 5111 5788 5145 0 FreeSans 400 0 0 0 x27.Q
flabel locali 5754 5179 5788 5213 0 FreeSans 400 0 0 0 x27.Q
flabel locali 3456 5281 3490 5315 3 FreeSans 400 0 0 0 x27.VPWR
flabel locali 3824 4975 3858 5009 0 FreeSans 200 0 0 0 x27.D
flabel locali 3824 5043 3858 5077 0 FreeSans 200 0 0 0 x27.D
flabel locali 5474 5179 5508 5213 0 FreeSans 400 0 0 0 x27.Q_N
flabel locali 5474 5111 5508 5145 0 FreeSans 400 0 0 0 x27.Q_N
flabel locali 5474 4839 5508 4873 0 FreeSans 400 0 0 0 x27.Q_N
flabel metal1 3456 4737 3490 4771 0 FreeSans 200 0 0 0 x27.VGND
flabel metal1 3456 5281 3490 5315 0 FreeSans 200 0 0 0 x27.VPWR
flabel nwell 3456 5281 3490 5315 3 FreeSans 400 0 0 0 x27.VPB
flabel nwell 3473 5298 3473 5298 0 FreeSans 200 0 0 0 x27.VPB
flabel pwell 3456 4737 3490 4771 3 FreeSans 400 0 0 0 x27.VNB
flabel pwell 3473 4754 3473 4754 0 FreeSans 200 0 0 0 x27.VNB
rlabel comment 3426 4754 3426 4754 4 x27.dfbbp_1
rlabel locali 4918 4901 4993 4967 1 x27.SET_B
rlabel metal1 4916 4938 4974 4947 1 x27.SET_B
rlabel metal1 4916 4901 4974 4910 1 x27.SET_B
rlabel metal1 4180 4938 4238 4947 1 x27.SET_B
rlabel metal1 4180 4910 4974 4938 1 x27.SET_B
rlabel metal1 4180 4901 4238 4910 1 x27.SET_B
rlabel metal1 3426 4706 5818 4802 1 x27.VGND
rlabel metal1 3426 5250 5818 5346 1 x27.VPWR
flabel locali 2897 4973 2972 5019 0 FreeSans 400 0 0 0 x20.RESET_B
flabel locali 1064 4737 1098 4771 3 FreeSans 400 0 0 0 x20.VGND
flabel locali 1064 4975 1098 5009 0 FreeSans 400 0 0 0 x20.CLK
flabel locali 1064 5043 1098 5077 0 FreeSans 400 0 0 0 x20.CLK
flabel locali 1800 4907 1834 4941 0 FreeSans 400 0 0 0 x20.SET_B
flabel locali 3362 4839 3396 4873 0 FreeSans 400 0 0 0 x20.Q
flabel locali 3362 5111 3396 5145 0 FreeSans 400 0 0 0 x20.Q
flabel locali 3362 5179 3396 5213 0 FreeSans 400 0 0 0 x20.Q
flabel locali 1064 5281 1098 5315 3 FreeSans 400 0 0 0 x20.VPWR
flabel locali 1432 4975 1466 5009 0 FreeSans 200 0 0 0 x20.D
flabel locali 1432 5043 1466 5077 0 FreeSans 200 0 0 0 x20.D
flabel locali 3082 5179 3116 5213 0 FreeSans 400 0 0 0 x20.Q_N
flabel locali 3082 5111 3116 5145 0 FreeSans 400 0 0 0 x20.Q_N
flabel locali 3082 4839 3116 4873 0 FreeSans 400 0 0 0 x20.Q_N
flabel metal1 1064 4737 1098 4771 0 FreeSans 200 0 0 0 x20.VGND
flabel metal1 1064 5281 1098 5315 0 FreeSans 200 0 0 0 x20.VPWR
flabel nwell 1064 5281 1098 5315 3 FreeSans 400 0 0 0 x20.VPB
flabel nwell 1081 5298 1081 5298 0 FreeSans 200 0 0 0 x20.VPB
flabel pwell 1064 4737 1098 4771 3 FreeSans 400 0 0 0 x20.VNB
flabel pwell 1081 4754 1081 4754 0 FreeSans 200 0 0 0 x20.VNB
rlabel comment 1034 4754 1034 4754 4 x20.dfbbp_1
rlabel locali 2526 4901 2601 4967 1 x20.SET_B
rlabel metal1 2524 4938 2582 4947 1 x20.SET_B
rlabel metal1 2524 4901 2582 4910 1 x20.SET_B
rlabel metal1 1788 4938 1846 4947 1 x20.SET_B
rlabel metal1 1788 4910 2582 4938 1 x20.SET_B
rlabel metal1 1788 4901 1846 4910 1 x20.SET_B
rlabel metal1 1034 4706 3426 4802 1 x20.VGND
rlabel metal1 1034 5250 3426 5346 1 x20.VPWR
flabel metal1 932 3718 966 3752 0 FreeSans 200 0 0 0 x7.VPWR
flabel metal1 932 3174 966 3208 0 FreeSans 200 0 0 0 x7.VGND
flabel locali 1208 3412 1242 3446 0 FreeSans 200 0 0 0 x7.X
flabel locali 1208 3480 1242 3514 0 FreeSans 200 0 0 0 x7.X
flabel locali 1208 3344 1242 3378 0 FreeSans 200 0 0 0 x7.X
flabel locali 932 3718 966 3752 0 FreeSans 200 0 0 0 x7.VPWR
flabel locali 932 3174 966 3208 0 FreeSans 200 0 0 0 x7.VGND
flabel locali 932 3412 966 3446 0 FreeSans 200 0 0 0 x7.A
flabel nwell 932 3718 966 3752 0 FreeSans 200 0 0 0 x7.VPB
flabel pwell 932 3174 966 3208 0 FreeSans 200 0 0 0 x7.VNB
rlabel comment 902 3191 902 3191 4 x7.buf_4
rlabel metal1 902 3143 1454 3239 1 x7.VGND
rlabel metal1 902 3687 1454 3783 1 x7.VPWR
flabel metal1 657 3174 691 3208 0 FreeSans 200 0 0 0 x6.VGND
flabel metal1 655 3718 689 3752 0 FreeSans 200 0 0 0 x6.VPWR
flabel locali 655 3718 689 3752 0 FreeSans 200 0 0 0 x6.VPWR
flabel locali 657 3174 691 3208 0 FreeSans 200 0 0 0 x6.VGND
flabel locali 837 3276 871 3310 0 FreeSans 200 0 0 0 x6.X
flabel locali 837 3548 871 3582 0 FreeSans 200 0 0 0 x6.X
flabel locali 837 3616 871 3650 0 FreeSans 200 0 0 0 x6.X
flabel locali 655 3412 689 3446 0 FreeSans 200 0 0 0 x6.A
flabel nwell 655 3718 689 3752 0 FreeSans 200 0 0 0 x6.VPB
flabel pwell 657 3174 691 3208 0 FreeSans 200 0 0 0 x6.VNB
rlabel comment 626 3191 626 3191 4 x6.buf_1
rlabel metal1 626 3143 902 3239 1 x6.VGND
rlabel metal1 626 3687 902 3783 1 x6.VPWR
flabel metal1 1341 6154 1375 6188 0 FreeSans 200 0 0 0 x5.VPWR
flabel metal1 1341 5610 1375 5644 0 FreeSans 200 0 0 0 x5.VGND
flabel locali 1617 5848 1651 5882 0 FreeSans 200 0 0 0 x5.X
flabel locali 1617 5916 1651 5950 0 FreeSans 200 0 0 0 x5.X
flabel locali 1617 5780 1651 5814 0 FreeSans 200 0 0 0 x5.X
flabel locali 1341 6154 1375 6188 0 FreeSans 200 0 0 0 x5.VPWR
flabel locali 1341 5610 1375 5644 0 FreeSans 200 0 0 0 x5.VGND
flabel locali 1341 5848 1375 5882 0 FreeSans 200 0 0 0 x5.A
flabel nwell 1341 6154 1375 6188 0 FreeSans 200 0 0 0 x5.VPB
flabel pwell 1341 5610 1375 5644 0 FreeSans 200 0 0 0 x5.VNB
rlabel comment 1311 5627 1311 5627 4 x5.buf_4
rlabel metal1 1311 5579 1863 5675 1 x5.VGND
rlabel metal1 1311 6123 1863 6219 1 x5.VPWR
flabel locali 1800 4286 1834 4320 0 FreeSans 200 0 0 0 x4.A
flabel locali 1708 4286 1742 4320 0 FreeSans 200 0 0 0 x4.A
flabel locali 3363 4286 3397 4320 0 FreeSans 200 0 0 0 x4.X
flabel locali 3363 4354 3397 4388 0 FreeSans 200 0 0 0 x4.X
flabel pwell 1432 4048 1466 4082 0 FreeSans 200 0 0 0 x4.VNB
flabel nwell 1432 4592 1466 4626 0 FreeSans 200 0 0 0 x4.VPB
flabel metal1 1432 4048 1466 4082 0 FreeSans 200 0 0 0 x4.VGND
flabel metal1 1432 4592 1466 4626 0 FreeSans 200 0 0 0 x4.VPWR
rlabel comment 1402 4065 1402 4065 4 x4.buf_16
rlabel metal1 1402 4017 3426 4113 1 x4.VGND
rlabel metal1 1402 4561 3426 4657 1 x4.VPWR
flabel metal1 900 4592 934 4626 0 FreeSans 200 0 0 0 x3.VPWR
flabel metal1 900 4048 934 4082 0 FreeSans 200 0 0 0 x3.VGND
flabel locali 1176 4286 1210 4320 0 FreeSans 200 0 0 0 x3.X
flabel locali 1176 4354 1210 4388 0 FreeSans 200 0 0 0 x3.X
flabel locali 1176 4218 1210 4252 0 FreeSans 200 0 0 0 x3.X
flabel locali 900 4592 934 4626 0 FreeSans 200 0 0 0 x3.VPWR
flabel locali 900 4048 934 4082 0 FreeSans 200 0 0 0 x3.VGND
flabel locali 900 4286 934 4320 0 FreeSans 200 0 0 0 x3.A
flabel nwell 900 4592 934 4626 0 FreeSans 200 0 0 0 x3.VPB
flabel pwell 900 4048 934 4082 0 FreeSans 200 0 0 0 x3.VNB
rlabel comment 870 4065 870 4065 4 x3.buf_4
rlabel metal1 870 4017 1422 4113 1 x3.VGND
rlabel metal1 870 4561 1422 4657 1 x3.VPWR
flabel metal1 1066 5610 1100 5644 0 FreeSans 200 0 0 0 x2.VGND
flabel metal1 1064 6154 1098 6188 0 FreeSans 200 0 0 0 x2.VPWR
flabel locali 1064 6154 1098 6188 0 FreeSans 200 0 0 0 x2.VPWR
flabel locali 1066 5610 1100 5644 0 FreeSans 200 0 0 0 x2.VGND
flabel locali 1246 5712 1280 5746 0 FreeSans 200 0 0 0 x2.X
flabel locali 1246 5984 1280 6018 0 FreeSans 200 0 0 0 x2.X
flabel locali 1246 6052 1280 6086 0 FreeSans 200 0 0 0 x2.X
flabel locali 1064 5848 1098 5882 0 FreeSans 200 0 0 0 x2.A
flabel nwell 1064 6154 1098 6188 0 FreeSans 200 0 0 0 x2.VPB
flabel pwell 1066 5610 1100 5644 0 FreeSans 200 0 0 0 x2.VNB
rlabel comment 1035 5627 1035 5627 4 x2.buf_1
rlabel metal1 1035 5579 1311 5675 1 x2.VGND
rlabel metal1 1035 6123 1311 6219 1 x2.VPWR
flabel metal1 625 4048 659 4082 0 FreeSans 200 0 0 0 x1.VGND
flabel metal1 623 4592 657 4626 0 FreeSans 200 0 0 0 x1.VPWR
flabel locali 623 4592 657 4626 0 FreeSans 200 0 0 0 x1.VPWR
flabel locali 625 4048 659 4082 0 FreeSans 200 0 0 0 x1.VGND
flabel locali 805 4150 839 4184 0 FreeSans 200 0 0 0 x1.X
flabel locali 805 4422 839 4456 0 FreeSans 200 0 0 0 x1.X
flabel locali 805 4490 839 4524 0 FreeSans 200 0 0 0 x1.X
flabel locali 623 4286 657 4320 0 FreeSans 200 0 0 0 x1.A
flabel nwell 623 4592 657 4626 0 FreeSans 200 0 0 0 x1.VPB
flabel pwell 625 4048 659 4082 0 FreeSans 200 0 0 0 x1.VNB
rlabel comment 594 4065 594 4065 4 x1.buf_1
rlabel metal1 594 4017 870 4113 1 x1.VGND
rlabel metal1 594 4561 870 4657 1 x1.VPWR
flabel pwell 4071 5610 4105 5644 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__mux4_4_0.VNB
flabel nwell 4071 6154 4105 6188 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__mux4_4_0.VPB
flabel metal1 4071 5610 4105 5644 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__mux4_4_0.VGND
flabel metal1 4071 6154 4105 6188 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__mux4_4_0.VPWR
flabel locali 2415 5712 2449 5746 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__mux4_4_0.X
flabel locali 2415 5780 2449 5814 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__mux4_4_0.X
flabel locali 2415 5848 2449 5882 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__mux4_4_0.X
flabel locali 2415 5916 2449 5950 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__mux4_4_0.X
flabel locali 2415 5984 2449 6018 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__mux4_4_0.X
flabel locali 2415 6052 2449 6086 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__mux4_4_0.X
flabel locali 4071 5848 4105 5882 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__mux4_4_0.S0
flabel locali 4071 5916 4105 5950 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__mux4_4_0.S0
flabel locali 3887 5780 3921 5814 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__mux4_4_0.A2
flabel locali 3887 5712 3921 5746 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__mux4_4_0.A2
flabel locali 3611 5780 3645 5814 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__mux4_4_0.A3
flabel locali 3611 5848 3645 5882 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__mux4_4_0.A3
flabel locali 3519 5848 3553 5882 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__mux4_4_0.S1
flabel locali 3519 5780 3553 5814 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__mux4_4_0.S1
flabel locali 3151 5848 3185 5882 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__mux4_4_0.A1
flabel locali 3151 5780 3185 5814 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__mux4_4_0.A1
flabel locali 2783 5780 2817 5814 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__mux4_4_0.A0
flabel locali 2783 5712 2817 5746 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__mux4_4_0.A0
rlabel comment 4135 5627 4135 5627 6 sky130_fd_sc_hd__mux4_4_0.mux4_4
rlabel locali 3856 5884 3890 5916 1 sky130_fd_sc_hd__mux4_4_0.S0
rlabel locali 3856 5916 3933 5950 1 sky130_fd_sc_hd__mux4_4_0.S0
rlabel locali 2841 5876 2909 5956 1 sky130_fd_sc_hd__mux4_4_0.S0
rlabel metal1 2863 5947 2921 5956 1 sky130_fd_sc_hd__mux4_4_0.S0
rlabel metal1 2863 5910 2921 5919 1 sky130_fd_sc_hd__mux4_4_0.S0
rlabel metal1 3875 5947 3933 5956 1 sky130_fd_sc_hd__mux4_4_0.S0
rlabel metal1 3875 5910 3933 5919 1 sky130_fd_sc_hd__mux4_4_0.S0
rlabel metal1 4059 5947 4118 5956 1 sky130_fd_sc_hd__mux4_4_0.S0
rlabel metal1 2863 5919 4118 5947 1 sky130_fd_sc_hd__mux4_4_0.S0
rlabel metal1 4059 5910 4118 5919 1 sky130_fd_sc_hd__mux4_4_0.S0
rlabel metal1 2295 5579 4135 5675 1 sky130_fd_sc_hd__mux4_4_0.VGND
rlabel metal1 2295 6123 4135 6219 1 sky130_fd_sc_hd__mux4_4_0.VPWR
<< end >>
