magic
tech sky130A
magscale 1 2
timestamp 1698381494
<< pwell >>
rect 1006 4372 1032 4404
rect 1612 4372 1638 4404
rect 1006 3214 1032 3246
rect 1612 3214 1638 3246
<< metal3 >>
rect 686 5180 1964 5182
rect 686 5116 790 5180
rect 854 5116 870 5180
rect 934 5116 950 5180
rect 1014 5116 1030 5180
rect 1094 5116 1110 5180
rect 1174 5116 1190 5180
rect 1254 5116 1396 5180
rect 1460 5116 1476 5180
rect 1540 5116 1556 5180
rect 1620 5116 1636 5180
rect 1700 5116 1716 5180
rect 1780 5116 1796 5180
rect 1860 5116 1964 5180
rect 686 5114 1964 5116
rect 686 4932 752 5114
rect 686 4868 687 4932
rect 751 4868 752 4932
rect 686 4852 752 4868
rect 686 4788 687 4852
rect 751 4788 752 4852
rect 686 4772 752 4788
rect 686 4708 687 4772
rect 751 4708 752 4772
rect 686 4692 752 4708
rect 686 4628 687 4692
rect 751 4628 752 4692
rect 686 4612 752 4628
rect 686 4548 687 4612
rect 751 4548 752 4612
rect 686 4532 752 4548
rect 686 4468 687 4532
rect 751 4468 752 4532
rect 686 4452 752 4468
rect 686 4388 687 4452
rect 751 4388 752 4452
rect 686 4372 752 4388
rect 686 4308 687 4372
rect 751 4308 752 4372
rect 686 4292 752 4308
rect 686 4228 687 4292
rect 751 4228 752 4292
rect 686 4212 752 4228
rect 686 4148 687 4212
rect 751 4148 752 4212
rect 686 4084 752 4148
rect 812 4084 872 5114
rect 932 4024 992 5054
rect 1052 4084 1112 5114
rect 1172 4024 1232 5054
rect 1292 4932 1358 5114
rect 1292 4868 1293 4932
rect 1357 4868 1358 4932
rect 1292 4852 1358 4868
rect 1292 4788 1293 4852
rect 1357 4788 1358 4852
rect 1292 4772 1358 4788
rect 1292 4708 1293 4772
rect 1357 4708 1358 4772
rect 1292 4692 1358 4708
rect 1292 4628 1293 4692
rect 1357 4628 1358 4692
rect 1292 4612 1358 4628
rect 1292 4548 1293 4612
rect 1357 4548 1358 4612
rect 1292 4532 1358 4548
rect 1292 4468 1293 4532
rect 1357 4468 1358 4532
rect 1292 4452 1358 4468
rect 1292 4388 1293 4452
rect 1357 4388 1358 4452
rect 1292 4372 1358 4388
rect 1292 4308 1293 4372
rect 1357 4308 1358 4372
rect 1292 4292 1358 4308
rect 1292 4228 1293 4292
rect 1357 4228 1358 4292
rect 1292 4212 1358 4228
rect 1292 4148 1293 4212
rect 1357 4148 1358 4212
rect 1292 4024 1358 4148
rect 1418 4084 1478 5114
rect 1538 4024 1598 5054
rect 1658 4084 1718 5114
rect 1778 4024 1838 5054
rect 1898 4932 1964 5050
rect 1898 4868 1899 4932
rect 1963 4868 1964 4932
rect 1898 4852 1964 4868
rect 1898 4788 1899 4852
rect 1963 4788 1964 4852
rect 1898 4772 1964 4788
rect 1898 4708 1899 4772
rect 1963 4708 1964 4772
rect 1898 4692 1964 4708
rect 1898 4628 1899 4692
rect 1963 4628 1964 4692
rect 1898 4612 1964 4628
rect 1898 4548 1899 4612
rect 1963 4548 1964 4612
rect 1898 4532 1964 4548
rect 1898 4468 1899 4532
rect 1963 4468 1964 4532
rect 1898 4452 1964 4468
rect 1898 4388 1899 4452
rect 1963 4388 1964 4452
rect 1898 4372 1964 4388
rect 1898 4308 1899 4372
rect 1963 4308 1964 4372
rect 1898 4292 1964 4308
rect 1898 4228 1899 4292
rect 1963 4228 1964 4292
rect 1898 4212 1964 4228
rect 1898 4148 1899 4212
rect 1963 4148 1964 4212
rect 1898 4024 1964 4148
rect 686 4022 1964 4024
rect 686 3958 790 4022
rect 854 3958 870 4022
rect 934 3958 950 4022
rect 1014 3958 1030 4022
rect 1094 3958 1110 4022
rect 1174 3958 1190 4022
rect 1254 3958 1396 4022
rect 1460 3958 1476 4022
rect 1540 3958 1556 4022
rect 1620 3958 1636 4022
rect 1700 3958 1716 4022
rect 1780 3958 1796 4022
rect 1860 3958 1964 4022
rect 686 3956 1964 3958
rect 686 3774 752 3956
rect 686 3710 687 3774
rect 751 3710 752 3774
rect 686 3694 752 3710
rect 686 3630 687 3694
rect 751 3630 752 3694
rect 686 3614 752 3630
rect 686 3550 687 3614
rect 751 3550 752 3614
rect 686 3534 752 3550
rect 686 3470 687 3534
rect 751 3470 752 3534
rect 686 3454 752 3470
rect 686 3390 687 3454
rect 751 3390 752 3454
rect 686 3374 752 3390
rect 686 3310 687 3374
rect 751 3310 752 3374
rect 686 3294 752 3310
rect 686 3230 687 3294
rect 751 3230 752 3294
rect 686 3214 752 3230
rect 686 3150 687 3214
rect 751 3150 752 3214
rect 686 3134 752 3150
rect 686 3070 687 3134
rect 751 3070 752 3134
rect 686 3054 752 3070
rect 686 2990 687 3054
rect 751 2990 752 3054
rect 686 2926 752 2990
rect 812 2926 872 3956
rect 932 2866 992 3896
rect 1052 2926 1112 3956
rect 1172 2866 1232 3896
rect 1292 3774 1358 3956
rect 1292 3710 1293 3774
rect 1357 3710 1358 3774
rect 1292 3694 1358 3710
rect 1292 3630 1293 3694
rect 1357 3630 1358 3694
rect 1292 3614 1358 3630
rect 1292 3550 1293 3614
rect 1357 3550 1358 3614
rect 1292 3534 1358 3550
rect 1292 3470 1293 3534
rect 1357 3470 1358 3534
rect 1292 3454 1358 3470
rect 1292 3390 1293 3454
rect 1357 3390 1358 3454
rect 1292 3374 1358 3390
rect 1292 3310 1293 3374
rect 1357 3310 1358 3374
rect 1292 3294 1358 3310
rect 1292 3230 1293 3294
rect 1357 3230 1358 3294
rect 1292 3214 1358 3230
rect 1292 3150 1293 3214
rect 1357 3150 1358 3214
rect 1292 3134 1358 3150
rect 1292 3070 1293 3134
rect 1357 3070 1358 3134
rect 1292 3054 1358 3070
rect 1292 2990 1293 3054
rect 1357 2990 1358 3054
rect 1292 2866 1358 2990
rect 1418 2926 1478 3956
rect 1538 2866 1598 3896
rect 1658 2926 1718 3956
rect 1778 2866 1838 3896
rect 1898 3774 1964 3892
rect 1898 3710 1899 3774
rect 1963 3710 1964 3774
rect 1898 3694 1964 3710
rect 1898 3630 1899 3694
rect 1963 3630 1964 3694
rect 1898 3614 1964 3630
rect 1898 3550 1899 3614
rect 1963 3550 1964 3614
rect 1898 3534 1964 3550
rect 1898 3470 1899 3534
rect 1963 3470 1964 3534
rect 1898 3454 1964 3470
rect 1898 3390 1899 3454
rect 1963 3390 1964 3454
rect 1898 3374 1964 3390
rect 1898 3310 1899 3374
rect 1963 3310 1964 3374
rect 1898 3294 1964 3310
rect 1898 3230 1899 3294
rect 1963 3230 1964 3294
rect 1898 3214 1964 3230
rect 1898 3150 1899 3214
rect 1963 3150 1964 3214
rect 1898 3134 1964 3150
rect 1898 3070 1899 3134
rect 1963 3070 1964 3134
rect 1898 3054 1964 3070
rect 1898 2990 1899 3054
rect 1963 2990 1964 3054
rect 1898 2866 1964 2990
rect 686 2864 1964 2866
rect 686 2800 790 2864
rect 854 2800 870 2864
rect 934 2800 950 2864
rect 1014 2800 1030 2864
rect 1094 2800 1110 2864
rect 1174 2800 1190 2864
rect 1254 2800 1396 2864
rect 1460 2800 1476 2864
rect 1540 2800 1556 2864
rect 1620 2800 1636 2864
rect 1700 2800 1716 2864
rect 1780 2800 1796 2864
rect 1860 2800 1964 2864
rect 686 2798 1964 2800
<< via3 >>
rect 790 5116 854 5180
rect 870 5116 934 5180
rect 950 5116 1014 5180
rect 1030 5116 1094 5180
rect 1110 5116 1174 5180
rect 1190 5116 1254 5180
rect 1396 5116 1460 5180
rect 1476 5116 1540 5180
rect 1556 5116 1620 5180
rect 1636 5116 1700 5180
rect 1716 5116 1780 5180
rect 1796 5116 1860 5180
rect 687 4868 751 4932
rect 687 4788 751 4852
rect 687 4708 751 4772
rect 687 4628 751 4692
rect 687 4548 751 4612
rect 687 4468 751 4532
rect 687 4388 751 4452
rect 687 4308 751 4372
rect 687 4228 751 4292
rect 687 4148 751 4212
rect 1293 4868 1357 4932
rect 1293 4788 1357 4852
rect 1293 4708 1357 4772
rect 1293 4628 1357 4692
rect 1293 4548 1357 4612
rect 1293 4468 1357 4532
rect 1293 4388 1357 4452
rect 1293 4308 1357 4372
rect 1293 4228 1357 4292
rect 1293 4148 1357 4212
rect 1899 4868 1963 4932
rect 1899 4788 1963 4852
rect 1899 4708 1963 4772
rect 1899 4628 1963 4692
rect 1899 4548 1963 4612
rect 1899 4468 1963 4532
rect 1899 4388 1963 4452
rect 1899 4308 1963 4372
rect 1899 4228 1963 4292
rect 1899 4148 1963 4212
rect 790 3958 854 4022
rect 870 3958 934 4022
rect 950 3958 1014 4022
rect 1030 3958 1094 4022
rect 1110 3958 1174 4022
rect 1190 3958 1254 4022
rect 1396 3958 1460 4022
rect 1476 3958 1540 4022
rect 1556 3958 1620 4022
rect 1636 3958 1700 4022
rect 1716 3958 1780 4022
rect 1796 3958 1860 4022
rect 687 3710 751 3774
rect 687 3630 751 3694
rect 687 3550 751 3614
rect 687 3470 751 3534
rect 687 3390 751 3454
rect 687 3310 751 3374
rect 687 3230 751 3294
rect 687 3150 751 3214
rect 687 3070 751 3134
rect 687 2990 751 3054
rect 1293 3710 1357 3774
rect 1293 3630 1357 3694
rect 1293 3550 1357 3614
rect 1293 3470 1357 3534
rect 1293 3390 1357 3454
rect 1293 3310 1357 3374
rect 1293 3230 1357 3294
rect 1293 3150 1357 3214
rect 1293 3070 1357 3134
rect 1293 2990 1357 3054
rect 1899 3710 1963 3774
rect 1899 3630 1963 3694
rect 1899 3550 1963 3614
rect 1899 3470 1963 3534
rect 1899 3390 1963 3454
rect 1899 3310 1963 3374
rect 1899 3230 1963 3294
rect 1899 3150 1963 3214
rect 1899 3070 1963 3134
rect 1899 2990 1963 3054
rect 790 2800 854 2864
rect 870 2800 934 2864
rect 950 2800 1014 2864
rect 1030 2800 1094 2864
rect 1110 2800 1174 2864
rect 1190 2800 1254 2864
rect 1396 2800 1460 2864
rect 1476 2800 1540 2864
rect 1556 2800 1620 2864
rect 1636 2800 1700 2864
rect 1716 2800 1780 2864
rect 1796 2800 1860 2864
<< metal4 >>
rect 686 5180 1964 5182
rect 686 5116 790 5180
rect 854 5116 870 5180
rect 934 5116 950 5180
rect 1014 5116 1030 5180
rect 1094 5116 1110 5180
rect 1174 5116 1190 5180
rect 1254 5116 1396 5180
rect 1460 5116 1476 5180
rect 1540 5116 1556 5180
rect 1620 5116 1636 5180
rect 1700 5116 1716 5180
rect 1780 5116 1796 5180
rect 1860 5116 1964 5180
rect 686 5114 1964 5116
rect 686 4932 752 5114
rect 686 4868 687 4932
rect 751 4868 752 4932
rect 686 4852 752 4868
rect 686 4788 687 4852
rect 751 4788 752 4852
rect 686 4772 752 4788
rect 686 4708 687 4772
rect 751 4708 752 4772
rect 686 4692 752 4708
rect 686 4628 687 4692
rect 751 4628 752 4692
rect 686 4612 752 4628
rect 686 4548 687 4612
rect 751 4548 752 4612
rect 686 4532 752 4548
rect 686 4468 687 4532
rect 751 4468 752 4532
rect 686 4452 752 4468
rect 686 4388 687 4452
rect 751 4388 752 4452
rect 686 4372 752 4388
rect 686 4308 687 4372
rect 751 4308 752 4372
rect 686 4292 752 4308
rect 686 4228 687 4292
rect 751 4228 752 4292
rect 686 4212 752 4228
rect 686 4148 687 4212
rect 751 4148 752 4212
rect 686 4084 752 4148
rect 812 4024 872 5054
rect 932 4084 992 5114
rect 1052 4024 1112 5054
rect 1172 4084 1232 5114
rect 1292 4932 1358 5114
rect 1292 4868 1293 4932
rect 1357 4868 1358 4932
rect 1292 4852 1358 4868
rect 1292 4788 1293 4852
rect 1357 4788 1358 4852
rect 1292 4772 1358 4788
rect 1292 4708 1293 4772
rect 1357 4708 1358 4772
rect 1292 4692 1358 4708
rect 1292 4628 1293 4692
rect 1357 4628 1358 4692
rect 1292 4612 1358 4628
rect 1292 4548 1293 4612
rect 1357 4548 1358 4612
rect 1292 4532 1358 4548
rect 1292 4468 1293 4532
rect 1357 4468 1358 4532
rect 1292 4452 1358 4468
rect 1292 4388 1293 4452
rect 1357 4388 1358 4452
rect 1292 4372 1358 4388
rect 1292 4308 1293 4372
rect 1357 4308 1358 4372
rect 1292 4292 1358 4308
rect 1292 4228 1293 4292
rect 1357 4228 1358 4292
rect 1292 4212 1358 4228
rect 1292 4148 1293 4212
rect 1357 4148 1358 4212
rect 1292 4024 1358 4148
rect 1418 4024 1478 5054
rect 1538 4084 1598 5114
rect 1658 4024 1718 5054
rect 1778 4084 1838 5114
rect 1898 4932 1964 5050
rect 1898 4868 1899 4932
rect 1963 4868 1964 4932
rect 1898 4852 1964 4868
rect 1898 4788 1899 4852
rect 1963 4788 1964 4852
rect 1898 4772 1964 4788
rect 1898 4708 1899 4772
rect 1963 4708 1964 4772
rect 1898 4692 1964 4708
rect 1898 4628 1899 4692
rect 1963 4628 1964 4692
rect 1898 4612 1964 4628
rect 1898 4548 1899 4612
rect 1963 4548 1964 4612
rect 1898 4532 1964 4548
rect 1898 4468 1899 4532
rect 1963 4468 1964 4532
rect 1898 4452 1964 4468
rect 1898 4388 1899 4452
rect 1963 4388 1964 4452
rect 1898 4372 1964 4388
rect 1898 4308 1899 4372
rect 1963 4308 1964 4372
rect 1898 4292 1964 4308
rect 1898 4228 1899 4292
rect 1963 4228 1964 4292
rect 1898 4212 1964 4228
rect 1898 4148 1899 4212
rect 1963 4148 1964 4212
rect 1898 4024 1964 4148
rect 686 4022 1964 4024
rect 686 3958 790 4022
rect 854 3958 870 4022
rect 934 3958 950 4022
rect 1014 3958 1030 4022
rect 1094 3958 1110 4022
rect 1174 3958 1190 4022
rect 1254 3958 1396 4022
rect 1460 3958 1476 4022
rect 1540 3958 1556 4022
rect 1620 3958 1636 4022
rect 1700 3958 1716 4022
rect 1780 3958 1796 4022
rect 1860 3958 1964 4022
rect 686 3956 1964 3958
rect 686 3774 752 3956
rect 686 3710 687 3774
rect 751 3710 752 3774
rect 686 3694 752 3710
rect 686 3630 687 3694
rect 751 3630 752 3694
rect 686 3614 752 3630
rect 686 3550 687 3614
rect 751 3550 752 3614
rect 686 3534 752 3550
rect 686 3470 687 3534
rect 751 3470 752 3534
rect 686 3454 752 3470
rect 686 3390 687 3454
rect 751 3390 752 3454
rect 686 3374 752 3390
rect 686 3310 687 3374
rect 751 3310 752 3374
rect 686 3294 752 3310
rect 686 3230 687 3294
rect 751 3230 752 3294
rect 686 3214 752 3230
rect 686 3150 687 3214
rect 751 3150 752 3214
rect 686 3134 752 3150
rect 686 3070 687 3134
rect 751 3070 752 3134
rect 686 3054 752 3070
rect 686 2990 687 3054
rect 751 2990 752 3054
rect 686 2926 752 2990
rect 812 2866 872 3896
rect 932 2926 992 3956
rect 1052 2866 1112 3896
rect 1172 2926 1232 3956
rect 1292 3774 1358 3956
rect 1292 3710 1293 3774
rect 1357 3710 1358 3774
rect 1292 3694 1358 3710
rect 1292 3630 1293 3694
rect 1357 3630 1358 3694
rect 1292 3614 1358 3630
rect 1292 3550 1293 3614
rect 1357 3550 1358 3614
rect 1292 3534 1358 3550
rect 1292 3470 1293 3534
rect 1357 3470 1358 3534
rect 1292 3454 1358 3470
rect 1292 3390 1293 3454
rect 1357 3390 1358 3454
rect 1292 3374 1358 3390
rect 1292 3310 1293 3374
rect 1357 3310 1358 3374
rect 1292 3294 1358 3310
rect 1292 3230 1293 3294
rect 1357 3230 1358 3294
rect 1292 3214 1358 3230
rect 1292 3150 1293 3214
rect 1357 3150 1358 3214
rect 1292 3134 1358 3150
rect 1292 3070 1293 3134
rect 1357 3070 1358 3134
rect 1292 3054 1358 3070
rect 1292 2990 1293 3054
rect 1357 2990 1358 3054
rect 1292 2866 1358 2990
rect 1418 2866 1478 3896
rect 1538 2926 1598 3956
rect 1658 2866 1718 3896
rect 1778 2926 1838 3956
rect 1898 3774 1964 3892
rect 1898 3710 1899 3774
rect 1963 3710 1964 3774
rect 1898 3694 1964 3710
rect 1898 3630 1899 3694
rect 1963 3630 1964 3694
rect 1898 3614 1964 3630
rect 1898 3550 1899 3614
rect 1963 3550 1964 3614
rect 1898 3534 1964 3550
rect 1898 3470 1899 3534
rect 1963 3470 1964 3534
rect 1898 3454 1964 3470
rect 1898 3390 1899 3454
rect 1963 3390 1964 3454
rect 1898 3374 1964 3390
rect 1898 3310 1899 3374
rect 1963 3310 1964 3374
rect 1898 3294 1964 3310
rect 1898 3230 1899 3294
rect 1963 3230 1964 3294
rect 1898 3214 1964 3230
rect 1898 3150 1899 3214
rect 1963 3150 1964 3214
rect 1898 3134 1964 3150
rect 1898 3070 1899 3134
rect 1963 3070 1964 3134
rect 1898 3054 1964 3070
rect 1898 2990 1899 3054
rect 1963 2990 1964 3054
rect 1898 2866 1964 2990
rect 686 2864 1964 2866
rect 686 2800 790 2864
rect 854 2800 870 2864
rect 934 2800 950 2864
rect 1014 2800 1030 2864
rect 1094 2800 1110 2864
rect 1174 2800 1190 2864
rect 1254 2800 1396 2864
rect 1460 2800 1476 2864
rect 1540 2800 1556 2864
rect 1620 2800 1636 2864
rect 1700 2800 1716 2864
rect 1780 2800 1796 2864
rect 1860 2800 1964 2864
rect 686 2798 1964 2800
<< labels >>
flabel pwell 1612 4372 1638 4404 0 FreeSans 160 0 0 0 x1[3].SUB
flabel metal4 1554 4706 1580 4738 0 FreeSans 320 0 0 0 x1[3].CBOT
flabel metal4 1672 4116 1698 4148 0 FreeSans 320 0 0 0 x1[3].CTOP
flabel pwell 1006 4372 1032 4404 0 FreeSans 160 0 0 0 x1[1].SUB
flabel metal4 948 4706 974 4738 0 FreeSans 320 0 0 0 x1[1].CBOT
flabel metal4 1066 4116 1092 4148 0 FreeSans 320 0 0 0 x1[1].CTOP
flabel pwell 1612 3214 1638 3246 0 FreeSans 160 0 0 0 x1[2].SUB
flabel metal4 1554 3548 1580 3580 0 FreeSans 320 0 0 0 x1[2].CBOT
flabel metal4 1672 2958 1698 2990 0 FreeSans 320 0 0 0 x1[2].CTOP
flabel pwell 1006 3214 1032 3246 0 FreeSans 160 0 0 0 x1[0].SUB
flabel metal4 948 3548 974 3580 0 FreeSans 320 0 0 0 x1[0].CBOT
flabel metal4 1066 2958 1092 2990 0 FreeSans 320 0 0 0 x1[0].CTOP
<< end >>
