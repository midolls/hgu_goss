* NGSPICE file created from hgu_cdac_cap_2.ext - technology: sky130A

.subckt hgu_cdac_cap_2 SUB
C0 x2.CTOP x1.CBOT 5.11f
C1 x2.CBOT x2.CTOP 5.11f
.ends

