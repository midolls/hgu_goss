* NGSPICE file created from hgu_cdac_cap_8.ext - technology: sky130A

.subckt hgu_cdac_cap_8 SUB
C0 x1[6].CTOP x1[7].CTOP 20.2f
C1 x1[7].CTOP x1[7].CBOT 20.2f
.ends

