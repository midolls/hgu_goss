magic
tech sky130A
magscale 1 2
timestamp 1699578588
<< error_p >>
rect -15 64 15 68
rect 310 -41 368 -35
rect -29 -80 29 -74
rect 310 -75 322 -41
rect -29 -114 -17 -80
rect 310 -81 368 -75
rect -29 -120 29 -114
<< nmos >>
rect -15 -42 15 42
<< ndiff >>
rect -73 30 -15 42
rect -73 -30 -61 30
rect -27 -30 -15 30
rect -73 -42 -15 -30
rect 15 30 73 42
rect 15 -30 27 30
rect 61 -30 73 30
rect 15 -42 73 -30
<< ndiffc >>
rect -61 -30 -27 30
rect 27 -30 61 30
<< poly >>
rect -15 42 15 64
rect 306 -41 372 -25
rect -15 -64 15 -42
rect -33 -80 33 -64
rect -33 -114 -17 -80
rect 17 -114 33 -80
rect 306 -75 322 -41
rect 356 -75 372 -41
rect 306 -91 372 -75
rect -33 -130 33 -114
<< polycont >>
rect -17 -114 17 -80
rect 322 -75 356 -41
<< locali >>
rect -61 30 -27 46
rect -61 -46 -27 -30
rect 27 30 61 46
rect 27 -46 61 -30
rect 306 -75 322 -41
rect 356 -75 372 -41
rect -33 -114 -17 -80
rect 17 -114 33 -80
<< viali >>
rect -61 -30 -27 30
rect 27 -30 61 30
rect 322 -75 356 -41
rect -17 -114 17 -80
<< metal1 >>
rect -67 30 -21 42
rect -67 -30 -61 30
rect -27 -30 -21 30
rect -67 -42 -21 -30
rect 21 30 67 42
rect 21 -30 27 30
rect 61 -30 67 30
rect 21 -42 67 -30
rect 310 -41 368 -35
rect -29 -80 29 -74
rect -29 -114 -17 -80
rect 17 -114 29 -80
rect 310 -75 322 -41
rect 356 -75 368 -41
rect 310 -81 368 -75
rect -29 -120 29 -114
<< properties >>
string FIXED_BBOX -158 -199 158 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
