magic
tech sky130A
magscale 1 2
timestamp 1698047669
<< nwell >>
rect -36 1170 314 1230
rect 0 1152 276 1170
<< psubdiff >>
rect 0 590 276 592
rect 0 556 122 590
rect 156 556 276 590
<< nsubdiff >>
rect 0 1186 276 1192
rect 0 1152 120 1186
rect 154 1152 276 1186
<< psubdiffcont >>
rect 122 556 156 590
<< nsubdiffcont >>
rect 120 1152 154 1186
<< locali >>
rect 0 1186 276 1192
rect 0 1152 120 1186
rect 154 1152 276 1186
rect 0 1142 276 1152
rect 64 815 80 863
rect 164 765 210 915
rect 0 590 276 592
rect 0 556 122 590
rect 156 556 276 590
<< metal1 >>
rect 0 1142 276 1182
rect 0 617 276 648
rect 0 556 276 592
use sky130_fd_sc_hd__inv_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697965495
transform 1 0 0 0 1 600
box -38 -48 314 592
<< labels >>
flabel nsubdiffcont 120 1152 154 1186 0 FreeSans 160 0 0 0 VPB
port 1 nsew
flabel locali 0 1142 276 1192 0 FreeSans 160 0 0 0 VPWR
port 2 nsew
flabel locali 164 765 210 915 0 FreeSans 160 0 0 0 output
port 4 nsew
flabel metal1 122 556 156 590 0 FreeSans 160 0 0 0 VNB
port 5 nsew
flabel locali 64 815 80 863 0 FreeSans 160 0 0 0 input
port 3 nsew
flabel metal1 0 617 276 648 0 FreeSans 160 0 0 0 VGND
port 9 nsew
<< end >>
