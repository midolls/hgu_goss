* NGSPICE file created from hgu_cdac_half_flat.ext - technology: sky130A

.subckt hgu_cdac_half d<3> d<2> d<1> d<0> d<5> db<0> db<1> db<2> db<3> tb<1>
+ tb<2> tb<3> tb<4> VREF t<1> t<2> t<3> t<4> d<6> db<6> db<5> d<4> db<4> tb<0> tb<5>
+ t<0> t<5> t<6> tb<6> VDD VSS
X0 VREF.t235 d<3>.t0 hgu_cdac_8bit_array_3.drv<7:0>.t5 VDD.t147 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X1 VREF.t35 db<3>.t0 hgu_cdac_8bit_array_2.drv<7:0>.t15 VDD.t35 sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X2 hgu_cdac_8bit_array_2.drv<31:0>.t43 db<5>.t0 VREF.t56 VDD.t56 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X3 hgu_cdac_8bit_array_3.drv<63:0>.t89 d<6>.t0 VREF.t217 VDD.t216 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X4 VREF.t63 d<5>.t0 hgu_cdac_8bit_array_3.drv<31:0>.t46 VDD.t63 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X5 hgu_cdac_8bit_array_3.drv<63:0>.t20 d<6>.t1 VSS.t345 VSS.t344 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X6 hgu_cdac_8bit_array_3.drv<31:0>.t9 d<5>.t1 VSS.t161 VSS.t160 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X7 VSS.t397 db<6>.t0 hgu_cdac_8bit_array_2.drv<63:0>.t127 VSS.t396 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X8 VREF.t190 db<6>.t1 hgu_cdac_8bit_array_2.drv<63:0>.t63 VDD.t189 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X9 hgu_cdac_8bit_array_3.drv<63:0>.t127 d<6>.t2 VSS.t343 VSS.t342 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X10 VREF.t144 d<4>.t0 hgu_cdac_8bit_array_3.drv<15:0>.t15 VDD.t144 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X11 VSS.t63 db<5>.t1 hgu_cdac_8bit_array_2.drv<31:0>.t0 VSS.t62 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X12 hgu_cdac_8bit_array_3.drv<63:0>.t88 d<6>.t3 VREF.t121 VDD.t121 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X13 VREF.t122 d<6>.t4 hgu_cdac_8bit_array_3.drv<63:0>.t87 VDD.t122 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X14 VSS.t399 db<6>.t2 hgu_cdac_8bit_array_2.drv<63:0>.t126 VSS.t398 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X15 hgu_cdac_8bit_array_3.drv<31:0>.t45 d<5>.t2 VREF.t42 VDD.t42 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X16 VREF.t234 d<3>.t1 hgu_cdac_8bit_array_3.drv<7:0>.t4 VDD.t230 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X17 hgu_cdac_8bit_array_3.drv<1:0>.t3 d<1> VSS.t391 VSS.t390 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X18 hgu_cdac_8bit_array_3.drv<15:0>.t31 d<4>.t1 VSS.t369 VSS.t368 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X19 VSS.t193 db<6>.t3 hgu_cdac_8bit_array_2.drv<63:0>.t125 VSS.t192 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X20 hgu_cdac_8bit_array_3.drv<31:0>.t8 d<5>.t3 VSS.t159 VSS.t158 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X21 VREF.t86 db<6>.t4 hgu_cdac_8bit_array_2.drv<63:0>.t62 VDD.t86 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X22 hgu_cdac_8bit_array_2.drv<15:0>.t15 db<4>.t0 VREF.t112 VDD.t112 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X23 hgu_cdac_8bit_array_3.drv<63:0>.t126 d<6>.t5 VSS.t341 VSS.t340 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X24 VSS.t207 db<4>.t1 hgu_cdac_8bit_array_2.drv<15:0>.t31 VSS.t206 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X25 VSS.t61 db<5>.t2 hgu_cdac_8bit_array_2.drv<31:0>.t10 VSS.t60 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X26 VREF.t44 d<6>.t6 hgu_cdac_8bit_array_3.drv<63:0>.t86 VDD.t44 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X27 hgu_cdac_8bit_array_3.drv<15:0>.t14 d<4>.t2 VREF.t218 VDD.t217 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X28 hgu_cdac_8bit_array_3.drv<15:0>.t30 d<4>.t3 VSS.t439 VSS.t438 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X29 hgu_cdac_8bit_array_2.drv<63:0>.t124 db<6>.t5 VSS.t169 VSS.t168 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X30 hgu_cdac_8bit_array_2.drv<63:0>.t61 db<6>.t6 VREF.t203 VDD.t202 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X31 hgu_cdac_8bit_array_2.drv<1:0>.t3 db<1>.t0 VSS.t465 VSS.t464 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X32 VSS.t339 d<6>.t7 hgu_cdac_8bit_array_3.drv<63:0>.t125 VSS.t338 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X33 VREF.t156 db<6>.t7 hgu_cdac_8bit_array_2.drv<63:0>.t60 VDD.t156 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X34 hgu_cdac_8bit_array_3.drv<63:0>.t85 d<6>.t8 VREF.t9 VDD.t9 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X35 hgu_cdac_8bit_array_2.drv<7:0>.t3 db<3>.t1 VSS.t493 VSS.t492 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X36 hgu_cdac_8bit_array_2.drv<31:0>.t42 db<5>.t3 VREF.t174 VDD.t174 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X37 VSS.t199 db<6>.t8 hgu_cdac_8bit_array_2.drv<63:0>.t123 VSS.t198 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X38 VREF.t175 db<6>.t9 hgu_cdac_8bit_array_2.drv<63:0>.t59 VDD.t175 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X39 VREF.t48 d<6>.t9 hgu_cdac_8bit_array_3.drv<63:0>.t84 VDD.t48 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X40 hgu_cdac_8bit_array_2.drv<63:0>.t122 db<6>.t10 VSS.t201 VSS.t200 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X41 hgu_cdac_8bit_array_3.drv<63:0>.t124 d<6>.t10 VSS.t337 VSS.t336 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X42 VREF.t17 d<5>.t4 hgu_cdac_8bit_array_3.drv<31:0>.t44 VDD.t17 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X43 hgu_cdac_8bit_array_2.drv<7:0>.t14 db<3>.t2 VREF.t88 VDD.t88 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X44 VREF.t250 db<2>.t0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t3 VDD.t245 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X45 VSS.t335 d<6>.t11 hgu_cdac_8bit_array_3.drv<63:0>.t123 VSS.t334 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X46 VSS.t157 d<5>.t5 hgu_cdac_8bit_array_3.drv<31:0>.t7 VSS.t156 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X47 hgu_cdac_8bit_array_3.drv<7:0>.t10 d<3>.t2 VSS.t463 VSS.t462 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X48 hgu_cdac_8bit_array_3.drv<63:0>.t83 d<6>.t12 VREF.t143 VDD.t143 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X49 VSS.t167 db<6>.t11 hgu_cdac_8bit_array_2.drv<63:0>.t121 VSS.t166 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X50 hgu_cdac_8bit_array_3.drv<31:0>.t6 d<5>.t6 VSS.t155 VSS.t154 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X51 VREF.t221 d<6>.t13 hgu_cdac_8bit_array_3.drv<63:0>.t82 VDD.t220 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X52 hgu_cdac_8bit_array_3.drv<63:0>.t122 d<6>.t14 VSS.t333 VSS.t332 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X53 hgu_cdac_8bit_array_3.drv<63:0>.t116 d<6>.t15 VSS.t331 VSS.t330 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X54 VSS.t59 db<5>.t4 hgu_cdac_8bit_array_2.drv<31:0>.t9 VSS.t58 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X55 VREF.t85 db<6>.t12 hgu_cdac_8bit_array_2.drv<63:0>.t58 VDD.t85 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X56 VREF.t189 d<6>.t16 hgu_cdac_8bit_array_3.drv<63:0>.t81 VDD.t188 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X57 hgu_cdac_8bit_array_3.drv<31:0>.t43 d<5>.t7 VREF.t149 VDD.t149 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X58 hgu_cdac_8bit_array_2.drv<63:0>.t120 db<6>.t13 VSS.t443 VSS.t442 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X59 hgu_cdac_8bit_array_2.drv<31:0>.t41 db<5>.t5 VREF.t104 VDD.t104 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X60 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t7 db<2>.t1 VSS.t73 VSS.t72 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X61 VREF.t106 db<6>.t14 hgu_cdac_8bit_array_2.drv<63:0>.t57 VDD.t106 sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X62 hgu_cdac_8bit_array_2.drv<0>.t1 db<0>.t0 VSS.t347 VSS.t346 sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.35
X63 hgu_cdac_8bit_array_3.drv<63:0>.t115 d<6>.t17 VSS.t329 VSS.t328 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X64 VSS.t57 db<5>.t6 hgu_cdac_8bit_array_2.drv<31:0>.t8 VSS.t56 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X65 VREF.t195 db<6>.t15 hgu_cdac_8bit_array_2.drv<63:0>.t56 VDD.t194 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X66 VREF.t177 d<6>.t18 hgu_cdac_8bit_array_3.drv<63:0>.t80 VDD.t177 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X67 hgu_cdac_8bit_array_3.drv<15:0>.t13 d<4>.t4 VREF.t2 VDD.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X68 VREF.t205 d<6>.t19 hgu_cdac_8bit_array_3.drv<63:0>.t79 VDD.t204 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X69 VREF.t206 d<5>.t8 hgu_cdac_8bit_array_3.drv<31:0>.t42 VDD.t205 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X70 VSS.t379 d<4>.t5 hgu_cdac_8bit_array_3.drv<15:0>.t29 VSS.t378 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X71 hgu_cdac_8bit_array_2.drv<63:0>.t119 db<6>.t16 VSS.t409 VSS.t408 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X72 VREF.t253 db<4>.t2 hgu_cdac_8bit_array_2.drv<15:0>.t14 VDD.t248 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X73 VREF.t47 d<6>.t20 hgu_cdac_8bit_array_3.drv<63:0>.t78 VDD.t47 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X74 VREF.t161 db<5>.t7 hgu_cdac_8bit_array_2.drv<31:0>.t40 VDD.t161 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X75 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t7 d<2>.t0 VSS.t423 VSS.t422 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X76 hgu_cdac_8bit_array_2.drv<63:0>.t118 db<6>.t17 VSS.t431 VSS.t430 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X77 hgu_cdac_8bit_array_2.drv<63:0>.t55 db<6>.t18 VREF.t211 VDD.t210 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X78 VREF.t202 d<4>.t6 hgu_cdac_8bit_array_3.drv<15:0>.t12 VDD.t201 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X79 VREF.t38 db<6>.t19 hgu_cdac_8bit_array_2.drv<63:0>.t54 VDD.t38 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X80 VSS.t327 d<6>.t21 hgu_cdac_8bit_array_3.drv<63:0>.t114 VSS.t326 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X81 hgu_cdac_8bit_array_2.drv<15:0>.t30 db<4>.t3 VSS.t507 VSS.t506 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X82 VREF.t135 d<6>.t22 hgu_cdac_8bit_array_3.drv<63:0>.t77 VDD.t135 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X83 VSS.t501 d<4>.t7 hgu_cdac_8bit_array_3.drv<15:0>.t28 VSS.t500 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X84 hgu_cdac_8bit_array_3.drv<63:0>.t113 d<6>.t23 VSS.t325 VSS.t324 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X85 hgu_cdac_8bit_array_2.drv<31:0>.t39 db<5>.t8 VREF.t162 VDD.t162 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X86 VREF.t53 d<5>.t9 hgu_cdac_8bit_array_3.drv<31:0>.t41 VDD.t53 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X87 hgu_cdac_8bit_array_3.drv<31:0>.t5 d<5>.t10 VSS.t153 VSS.t152 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X88 VREF.t1 db<4>.t4 hgu_cdac_8bit_array_2.drv<15:0>.t13 VDD.t1 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X89 VREF.t91 db<5>.t9 hgu_cdac_8bit_array_2.drv<31:0>.t38 VDD.t91 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X90 VREF.t43 d<6>.t24 hgu_cdac_8bit_array_3.drv<63:0>.t76 VDD.t43 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X91 VSS.t323 d<6>.t25 hgu_cdac_8bit_array_3.drv<63:0>.t112 VSS.t322 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X92 hgu_cdac_8bit_array_2.drv<63:0>.t117 db<6>.t20 VSS.t89 VSS.t88 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X93 VSS.t151 d<5>.t11 hgu_cdac_8bit_array_3.drv<31:0>.t4 VSS.t150 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X94 hgu_cdac_8bit_array_3.drv<63:0>.t94 d<6>.t26 VSS.t321 VSS.t320 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X95 hgu_cdac_8bit_array_2.drv<63:0>.t53 db<6>.t21 VREF.t148 VDD.t148 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X96 hgu_cdac_8bit_array_3.drv<63:0>.t75 d<6>.t27 VREF.t140 VDD.t140 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X97 VSS.t371 db<6>.t22 hgu_cdac_8bit_array_2.drv<63:0>.t116 VSS.t370 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X98 hgu_cdac_8bit_array_2.drv<15:0>.t29 db<4>.t5 VSS.t429 VSS.t428 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X99 VREF.t184 d<1> hgu_cdac_8bit_array_3.drv<1:0>.t1 VDD.t155 sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X100 hgu_cdac_8bit_array_2.drv<15:0>.t28 db<4>.t6 VSS.t191 VSS.t190 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X101 hgu_cdac_8bit_array_2.drv<31:0>.t7 db<5>.t10 VSS.t55 VSS.t54 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X102 VREF.t147 db<3>.t3 hgu_cdac_8bit_array_2.drv<7:0>.t13 VDD.t147 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X103 hgu_cdac_8bit_array_3.drv<63:0>.t74 d<6>.t28 VREF.t45 VDD.t45 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X104 VREF.t55 d<5>.t12 hgu_cdac_8bit_array_3.drv<31:0>.t40 VDD.t55 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X105 hgu_cdac_8bit_array_2.drv<63:0>.t115 db<6>.t23 VSS.t355 VSS.t354 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X106 hgu_cdac_8bit_array_3.drv<63:0>.t93 d<6>.t29 VSS.t319 VSS.t318 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X107 VSS.t357 db<6>.t24 hgu_cdac_8bit_array_2.drv<63:0>.t114 VSS.t356 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X108 VSS.t461 d<3>.t3 hgu_cdac_8bit_array_3.drv<7:0>.t9 VSS.t460 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X109 hgu_cdac_8bit_array_3.drv<31:0>.t3 d<5>.t13 VSS.t149 VSS.t148 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X110 VREF.t82 db<6>.t25 hgu_cdac_8bit_array_2.drv<63:0>.t52 VDD.t82 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X111 VREF.t103 d<6>.t30 hgu_cdac_8bit_array_3.drv<63:0>.t73 VDD.t103 sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X112 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t3 d<2>.t1 VREF.t30 VDD.t30 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X113 VSS.t147 d<5>.t14 hgu_cdac_8bit_array_3.drv<31:0>.t2 VSS.t146 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X114 hgu_cdac_8bit_array_3.drv<63:0>.t92 d<6>.t31 VSS.t317 VSS.t316 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X115 VREF.t146 d<5>.t15 hgu_cdac_8bit_array_3.drv<31:0>.t39 VDD.t146 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X116 VSS.t53 db<5>.t11 hgu_cdac_8bit_array_2.drv<31:0>.t6 VSS.t52 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X117 hgu_cdac_8bit_array_2.drv<63:0>.t51 db<6>.t26 VREF.t83 VDD.t83 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X118 hgu_cdac_8bit_array_2.drv<15:0>.t27 db<4>.t7 VSS.t353 VSS.t352 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X119 VREF.t168 db<5>.t12 hgu_cdac_8bit_array_2.drv<31:0>.t37 VDD.t168 sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X120 VSS.t171 d<4>.t8 hgu_cdac_8bit_array_3.drv<15:0>.t27 VSS.t170 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X121 hgu_cdac_8bit_array_3.drv<63:0>.t91 d<6>.t32 VSS.t315 VSS.t314 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X122 VSS.t313 d<6>.t33 hgu_cdac_8bit_array_3.drv<63:0>.t90 VSS.t312 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X123 VSS.t459 d<3>.t4 hgu_cdac_8bit_array_3.drv<7:0>.t8 VSS.t458 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X124 hgu_cdac_8bit_array_3.drv<31:0>.t1 d<5>.t16 VSS.t145 VSS.t144 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X125 VREF.t239 db<6>.t27 hgu_cdac_8bit_array_2.drv<63:0>.t50 VDD.t234 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X126 hgu_cdac_8bit_array_2.drv<15:0>.t12 db<4>.t8 VREF.t248 VDD.t243 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X127 hgu_cdac_8bit_array_2.drv<7:0>.t2 db<3>.t4 VSS.t491 VSS.t490 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X128 VREF.t188 d<6>.t34 hgu_cdac_8bit_array_3.drv<63:0>.t72 VDD.t187 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X129 VREF.t98 db<5>.t13 hgu_cdac_8bit_array_2.drv<31:0>.t36 VDD.t98 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X130 hgu_cdac_8bit_array_2.drv<63:0>.t113 db<6>.t28 VSS.t475 VSS.t474 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X131 VSS.t403 db<2>.t2 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t6 VSS.t402 sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X132 hgu_cdac_8bit_array_3.drv<15:0>.t26 d<4>.t9 VSS.t393 VSS.t392 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X133 VSS.t311 d<6>.t35 hgu_cdac_8bit_array_3.drv<63:0>.t109 VSS.t310 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X134 hgu_cdac_8bit_array_2.drv<15:0>.t11 db<4>.t9 VREF.t160 VDD.t160 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X135 VREF.t176 d<5>.t17 hgu_cdac_8bit_array_3.drv<31:0>.t38 VDD.t176 sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X136 hgu_cdac_8bit_array_3.drv<0>.t0 d<0>.t0 VREF.t249 VDD.t244 sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.35
X137 VSS.t85 db<6>.t29 hgu_cdac_8bit_array_2.drv<63:0>.t112 VSS.t84 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X138 VREF.t152 d<6>.t36 hgu_cdac_8bit_array_3.drv<63:0>.t71 VDD.t152 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X139 hgu_cdac_8bit_array_2.drv<63:0>.t49 db<6>.t30 VREF.t31 VDD.t31 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X140 hgu_cdac_8bit_array_2.drv<63:0>.t111 db<6>.t31 VSS.t175 VSS.t174 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X141 hgu_cdac_8bit_array_3.drv<63:0>.t108 d<6>.t37 VSS.t309 VSS.t308 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X142 VSS.t51 db<5>.t14 hgu_cdac_8bit_array_2.drv<31:0>.t58 VSS.t50 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X143 VSS.t307 d<6>.t38 hgu_cdac_8bit_array_3.drv<63:0>.t107 VSS.t306 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X144 hgu_cdac_8bit_array_2.drv<31:0>.t57 db<5>.t15 VSS.t49 VSS.t48 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X145 VSS.t143 d<5>.t18 hgu_cdac_8bit_array_3.drv<31:0>.t0 VSS.t142 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X146 hgu_cdac_8bit_array_2.drv<63:0>.t48 db<6>.t32 VREF.t62 VDD.t62 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X147 hgu_cdac_8bit_array_2.drv<31:0>.t35 db<5>.t16 VREF.t142 VDD.t142 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X148 hgu_cdac_8bit_array_3.drv<63:0>.t70 d<6>.t39 VREF.t225 VDD.t224 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X149 hgu_cdac_8bit_array_3.drv<63:0>.t69 d<6>.t40 VREF.t0 VDD.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X150 VREF.t252 d<5>.t19 hgu_cdac_8bit_array_3.drv<31:0>.t37 VDD.t247 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X151 hgu_cdac_8bit_array_3.drv<31:0>.t36 d<5>.t20 VREF.t127 VDD.t127 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X152 VSS.t87 db<6>.t33 hgu_cdac_8bit_array_2.drv<63:0>.t110 VSS.t86 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X153 VREF.t34 db<6>.t34 hgu_cdac_8bit_array_2.drv<63:0>.t47 VDD.t34 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X154 hgu_cdac_8bit_array_3.drv<63:0>.t106 d<6>.t41 VSS.t305 VSS.t304 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X155 hgu_cdac_8bit_array_2.drv<7:0>.t1 db<3>.t5 VSS.t489 VSS.t488 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X156 hgu_cdac_8bit_array_2.drv<31:0>.t34 db<5>.t17 VREF.t163 VDD.t163 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X157 VSS.t47 db<5>.t18 hgu_cdac_8bit_array_2.drv<31:0>.t56 VSS.t46 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X158 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t5 db<2>.t3 VSS.t471 VSS.t470 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X159 VREF.t33 d<6>.t42 hgu_cdac_8bit_array_3.drv<63:0>.t68 VDD.t33 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X160 VSS.t303 d<6>.t43 hgu_cdac_8bit_array_3.drv<63:0>.t105 VSS.t302 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X161 hgu_cdac_8bit_array_3.drv<63:0>.t67 d<6>.t44 VREF.t32 VDD.t32 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X162 VSS.t417 db<6>.t35 hgu_cdac_8bit_array_2.drv<63:0>.t109 VSS.t416 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X163 hgu_cdac_8bit_array_3.drv<31:0>.t35 d<5>.t21 VREF.t61 VDD.t61 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X164 VREF.t223 d<2>.t2 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t2 VDD.t222 sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X165 VSS.t301 d<6>.t45 hgu_cdac_8bit_array_3.drv<63:0>.t9 VSS.t300 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X166 VSS.t419 db<6>.t36 hgu_cdac_8bit_array_2.drv<63:0>.t108 VSS.t418 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X167 VSS.t177 db<6>.t37 hgu_cdac_8bit_array_2.drv<63:0>.t107 VSS.t176 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X168 hgu_cdac_8bit_array_3.drv<31:0>.t14 d<5>.t22 VSS.t141 VSS.t140 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X169 VSS.t45 db<5>.t19 hgu_cdac_8bit_array_2.drv<31:0>.t55 VSS.t44 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X170 VREF.t66 db<6>.t38 hgu_cdac_8bit_array_2.drv<63:0>.t46 VDD.t66 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X171 VREF.t64 d<6>.t46 hgu_cdac_8bit_array_3.drv<63:0>.t66 VDD.t64 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X172 hgu_cdac_8bit_array_3.drv<15:0>.t11 d<4>.t10 VREF.t57 VDD.t57 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X173 VREF.t19 d<5>.t23 hgu_cdac_8bit_array_3.drv<31:0>.t34 VDD.t19 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X174 hgu_cdac_8bit_array_2.drv<63:0>.t106 db<6>.t39 VSS.t217 VSS.t216 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X175 VSS.t203 db<4>.t10 hgu_cdac_8bit_array_2.drv<15:0>.t26 VSS.t202 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X176 hgu_cdac_8bit_array_3.drv<63:0>.t65 d<6>.t47 VREF.t93 VDD.t93 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X177 hgu_cdac_8bit_array_3.drv<15:0>.t25 d<4>.t11 VSS.t497 VSS.t496 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X178 VSS.t299 d<6>.t48 hgu_cdac_8bit_array_3.drv<63:0>.t8 VSS.t298 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X179 VREF.t97 db<5>.t20 hgu_cdac_8bit_array_2.drv<31:0>.t33 VDD.t97 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X180 hgu_cdac_8bit_array_3.drv<31:0>.t33 d<5>.t24 VREF.t116 VDD.t116 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X181 VSS.t139 d<5>.t25 hgu_cdac_8bit_array_3.drv<31:0>.t13 VSS.t138 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X182 VSS.t297 d<6>.t49 hgu_cdac_8bit_array_3.drv<63:0>.t7 VSS.t296 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X183 VREF.t119 db<6>.t40 hgu_cdac_8bit_array_2.drv<63:0>.t45 VDD.t119 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X184 VSS.t487 db<3>.t6 hgu_cdac_8bit_array_2.drv<7:0>.t0 VSS.t486 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X185 VSS.t295 d<6>.t50 hgu_cdac_8bit_array_3.drv<63:0>.t6 VSS.t294 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X186 hgu_cdac_8bit_array_3.drv<15:0>.t10 d<4>.t12 VREF.t180 VDD.t180 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X187 VREF.t22 db<6>.t41 hgu_cdac_8bit_array_2.drv<63:0>.t44 VDD.t22 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X188 VSS.t469 d<4>.t13 hgu_cdac_8bit_array_3.drv<15:0>.t24 VSS.t468 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X189 hgu_cdac_8bit_array_2.drv<63:0>.t105 db<6>.t42 VSS.t69 VSS.t68 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X190 VSS.t67 db<4>.t11 hgu_cdac_8bit_array_2.drv<15:0>.t25 VSS.t66 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X191 hgu_cdac_8bit_array_3.drv<7:0>.t3 d<3>.t5 VREF.t233 VDD.t80 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X192 VREF.t178 db<4>.t12 hgu_cdac_8bit_array_2.drv<15:0>.t10 VDD.t178 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X193 VREF.t138 db<5>.t21 hgu_cdac_8bit_array_2.drv<31:0>.t32 VDD.t138 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X194 VREF.t52 d<6>.t51 hgu_cdac_8bit_array_3.drv<63:0>.t64 VDD.t52 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X195 VSS.t293 d<6>.t52 hgu_cdac_8bit_array_3.drv<63:0>.t5 VSS.t292 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X196 VSS.t137 d<5>.t26 hgu_cdac_8bit_array_3.drv<31:0>.t12 VSS.t136 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X197 hgu_cdac_8bit_array_2.drv<63:0>.t104 db<6>.t43 VSS.t363 VSS.t362 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X198 hgu_cdac_8bit_array_2.drv<63:0>.t43 db<6>.t44 VREF.t126 VDD.t126 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X199 VSS.t291 d<6>.t53 hgu_cdac_8bit_array_3.drv<63:0>.t104 VSS.t290 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X200 hgu_cdac_8bit_array_2.drv<1:0>.t1 db<1>.t1 VREF.t155 VDD.t155 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X201 hgu_cdac_8bit_array_2.drv<31:0>.t54 db<5>.t22 VSS.t43 VSS.t42 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X202 hgu_cdac_8bit_array_3.drv<63:0>.t103 d<6>.t54 VSS.t289 VSS.t288 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X203 hgu_cdac_8bit_array_3.drv<7:0>.t15 d<3>.t6 VREF.t232 VDD.t229 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X204 hgu_cdac_8bit_array_2.drv<7:0>.t12 db<3>.t7 VREF.t153 VDD.t153 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X205 VSS.t389 d<1> hgu_cdac_8bit_array_3.drv<1:0>.t2 VSS.t388 sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X206 VREF.t208 db<6>.t45 hgu_cdac_8bit_array_2.drv<63:0>.t42 VDD.t207 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X207 hgu_cdac_8bit_array_3.drv<63:0>.t102 d<6>.t55 VSS.t287 VSS.t286 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X208 hgu_cdac_8bit_array_2.drv<63:0>.t103 db<6>.t46 VSS.t425 VSS.t424 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X209 VSS.t135 d<5>.t27 hgu_cdac_8bit_array_3.drv<31:0>.t11 VSS.t134 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X210 hgu_cdac_8bit_array_2.drv<63:0>.t41 db<6>.t47 VREF.t179 VDD.t179 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X211 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t6 d<2>.t3 VSS.t187 VSS.t186 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X212 VSS.t285 d<6>.t56 hgu_cdac_8bit_array_3.drv<63:0>.t101 VSS.t284 sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X213 hgu_cdac_8bit_array_2.drv<63:0>.t102 db<6>.t48 VSS.t385 VSS.t384 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X214 VSS.t133 d<5>.t28 hgu_cdac_8bit_array_3.drv<31:0>.t10 VSS.t132 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X215 hgu_cdac_8bit_array_2.drv<31:0>.t5 db<5>.t23 VSS.t41 VSS.t40 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X216 hgu_cdac_8bit_array_3.drv<63:0>.t63 d<6>.t57 VREF.t23 VDD.t23 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X217 VSS.t39 db<5>.t24 hgu_cdac_8bit_array_2.drv<31:0>.t4 VSS.t38 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X218 VSS.t473 db<6>.t49 hgu_cdac_8bit_array_2.drv<63:0>.t101 VSS.t472 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X219 VREF.t238 db<6>.t50 hgu_cdac_8bit_array_2.drv<63:0>.t40 VDD.t233 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X220 VREF.t77 d<6>.t58 hgu_cdac_8bit_array_3.drv<63:0>.t62 VDD.t77 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X221 hgu_cdac_8bit_array_2.drv<31:0>.t3 db<5>.t25 VSS.t37 VSS.t36 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X222 VREF.t164 d<5>.t29 hgu_cdac_8bit_array_3.drv<31:0>.t32 VDD.t164 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X223 hgu_cdac_8bit_array_2.drv<63:0>.t100 db<6>.t51 VSS.t349 VSS.t348 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X224 VSS.t91 db<1>.t2 hgu_cdac_8bit_array_2.drv<1:0>.t2 VSS.t90 sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X225 hgu_cdac_8bit_array_2.drv<63:0>.t99 db<6>.t52 VSS.t351 VSS.t350 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X226 hgu_cdac_8bit_array_2.drv<63:0>.t98 db<6>.t53 VSS.t213 VSS.t212 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X227 VSS.t485 db<3>.t8 hgu_cdac_8bit_array_2.drv<7:0>.t7 VSS.t484 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X228 VREF.t92 db<5>.t26 hgu_cdac_8bit_array_2.drv<31:0>.t31 VDD.t92 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X229 VREF.t129 d<6>.t59 hgu_cdac_8bit_array_3.drv<63:0>.t61 VDD.t129 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X230 hgu_cdac_8bit_array_2.drv<63:0>.t97 db<6>.t54 VSS.t215 VSS.t214 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X231 hgu_cdac_8bit_array_2.drv<63:0>.t39 db<6>.t55 VREF.t157 VDD.t157 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X232 VSS.t283 d<6>.t60 hgu_cdac_8bit_array_3.drv<63:0>.t100 VSS.t282 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X233 hgu_cdac_8bit_array_2.drv<31:0>.t2 db<5>.t27 VSS.t35 VSS.t34 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X234 VREF.t136 d<5>.t30 hgu_cdac_8bit_array_3.drv<31:0>.t31 VDD.t136 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X235 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t2 db<2>.t4 VREF.t181 VDD.t181 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X236 hgu_cdac_8bit_array_2.drv<63:0>.t96 db<6>.t56 VSS.t377 VSS.t376 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X237 hgu_cdac_8bit_array_2.drv<0>.t0 db<0>.t1 VREF.t108 VDD.t108 sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.35
X238 VSS.t503 db<4>.t13 hgu_cdac_8bit_array_2.drv<15:0>.t24 VSS.t502 sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X239 VREF.t14 db<5>.t28 hgu_cdac_8bit_array_2.drv<31:0>.t30 VDD.t14 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X240 VREF.t96 d<6>.t61 hgu_cdac_8bit_array_3.drv<63:0>.t60 VDD.t96 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X241 hgu_cdac_8bit_array_2.drv<63:0>.t95 db<6>.t57 VSS.t71 VSS.t70 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X242 hgu_cdac_8bit_array_3.drv<0>.t1 d<0>.t1 VSS.t395 VSS.t394 sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.35
X243 VSS.t131 d<5>.t31 hgu_cdac_8bit_array_3.drv<31:0>.t56 VSS.t130 sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X244 hgu_cdac_8bit_array_2.drv<63:0>.t38 db<6>.t58 VREF.t25 VDD.t25 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X245 VSS.t281 d<6>.t62 hgu_cdac_8bit_array_3.drv<63:0>.t25 VSS.t280 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X246 hgu_cdac_8bit_array_2.drv<15:0>.t23 db<4>.t14 VSS.t93 VSS.t92 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X247 hgu_cdac_8bit_array_2.drv<31:0>.t1 db<5>.t29 VSS.t33 VSS.t32 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X248 hgu_cdac_8bit_array_2.drv<63:0>.t37 db<6>.t59 VREF.t198 VDD.t197 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X249 hgu_cdac_8bit_array_3.drv<63:0>.t59 d<6>.t63 VREF.t13 VDD.t13 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X250 VREF.t78 d<5>.t32 hgu_cdac_8bit_array_3.drv<31:0>.t30 VDD.t78 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X251 VSS.t411 db<6>.t60 hgu_cdac_8bit_array_2.drv<63:0>.t94 VSS.t410 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X252 VREF.t231 d<3>.t7 hgu_cdac_8bit_array_3.drv<7:0>.t14 VDD.t172 sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X253 hgu_cdac_8bit_array_2.drv<15:0>.t9 db<4>.t15 VREF.t67 VDD.t67 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X254 hgu_cdac_8bit_array_3.drv<63:0>.t58 d<6>.t64 VREF.t5 VDD.t5 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X255 hgu_cdac_8bit_array_3.drv<63:0>.t24 d<6>.t65 VSS.t279 VSS.t278 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X256 hgu_cdac_8bit_array_3.drv<63:0>.t23 d<6>.t66 VSS.t277 VSS.t276 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X257 VSS.t129 d<5>.t33 hgu_cdac_8bit_array_3.drv<31:0>.t55 VSS.t128 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X258 VSS.t373 db<6>.t61 hgu_cdac_8bit_array_2.drv<63:0>.t93 VSS.t372 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X259 hgu_cdac_8bit_array_3.drv<31:0>.t54 d<5>.t34 VSS.t127 VSS.t126 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X260 hgu_cdac_8bit_array_2.drv<63:0>.t92 db<6>.t62 VSS.t375 VSS.t374 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X261 hgu_cdac_8bit_array_2.drv<31:0>.t48 db<5>.t30 VSS.t31 VSS.t30 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X262 hgu_cdac_8bit_array_2.drv<63:0>.t36 db<6>.t63 VREF.t40 VDD.t40 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X263 hgu_cdac_8bit_array_3.drv<63:0>.t57 d<6>.t67 VREF.t128 VDD.t128 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X264 VREF.t70 d<4>.t14 hgu_cdac_8bit_array_3.drv<15:0>.t9 VDD.t70 sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X265 hgu_cdac_8bit_array_3.drv<31:0>.t29 d<5>.t35 VREF.t28 VDD.t28 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X266 VSS.t275 d<6>.t68 hgu_cdac_8bit_array_3.drv<63:0>.t22 VSS.t274 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X267 VSS.t95 db<6>.t64 hgu_cdac_8bit_array_2.drv<63:0>.t91 VSS.t94 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X268 VREF.t230 d<3>.t8 hgu_cdac_8bit_array_3.drv<7:0>.t13 VDD.t228 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X269 VREF.t240 db<6>.t65 hgu_cdac_8bit_array_2.drv<63:0>.t35 VDD.t235 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X270 hgu_cdac_8bit_array_2.drv<15:0>.t8 db<4>.t16 VREF.t219 VDD.t218 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X271 hgu_cdac_8bit_array_2.drv<31:0>.t47 db<5>.t31 VSS.t29 VSS.t28 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X272 hgu_cdac_8bit_array_3.drv<63:0>.t21 d<6>.t69 VSS.t273 VSS.t272 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X273 hgu_cdac_8bit_array_2.drv<15:0>.t7 db<4>.t17 VREF.t41 VDD.t41 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X274 hgu_cdac_8bit_array_3.drv<63:0>.t56 d<6>.t70 VREF.t169 VDD.t169 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X275 hgu_cdac_8bit_array_2.drv<31:0>.t29 db<5>.t32 VREF.t65 VDD.t65 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X276 VSS.t445 d<2>.t4 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t5 VSS.t444 sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X277 hgu_cdac_8bit_array_3.drv<31:0>.t53 d<5>.t36 VSS.t125 VSS.t124 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X278 hgu_cdac_8bit_array_2.drv<63:0>.t34 db<6>.t66 VREF.t241 VDD.t236 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X279 VREF.t76 db<6>.t67 hgu_cdac_8bit_array_2.drv<63:0>.t33 VDD.t76 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X280 VREF.t192 d<6>.t71 hgu_cdac_8bit_array_3.drv<63:0>.t55 VDD.t191 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X281 hgu_cdac_8bit_array_3.drv<15:0>.t8 d<4>.t15 VREF.t183 VDD.t183 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X282 hgu_cdac_8bit_array_2.drv<63:0>.t90 db<6>.t68 VSS.t185 VSS.t184 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X283 VSS.t97 db<4>.t18 hgu_cdac_8bit_array_2.drv<15:0>.t22 VSS.t96 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X284 hgu_cdac_8bit_array_3.drv<31:0>.t28 d<5>.t37 VREF.t6 VDD.t6 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X285 hgu_cdac_8bit_array_3.drv<15:0>.t23 d<4>.t16 VSS.t447 VSS.t446 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X286 VSS.t271 d<6>.t72 hgu_cdac_8bit_array_3.drv<63:0>.t99 VSS.t270 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X287 VREF.t46 db<5>.t33 hgu_cdac_8bit_array_2.drv<31:0>.t28 VDD.t46 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X288 VSS.t123 d<5>.t38 hgu_cdac_8bit_array_3.drv<31:0>.t52 VSS.t122 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X289 hgu_cdac_8bit_array_2.drv<15:0>.t6 db<4>.t19 VREF.t159 VDD.t159 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X290 hgu_cdac_8bit_array_3.drv<63:0>.t98 d<6>.t73 VSS.t269 VSS.t268 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X291 hgu_cdac_8bit_array_3.drv<31:0>.t51 d<5>.t39 VSS.t121 VSS.t120 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X292 VREF.t191 d<6>.t74 hgu_cdac_8bit_array_3.drv<63:0>.t54 VDD.t190 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X293 hgu_cdac_8bit_array_2.drv<63:0>.t89 db<6>.t69 VSS.t173 VSS.t172 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X294 VSS.t75 db<4>.t20 hgu_cdac_8bit_array_2.drv<15:0>.t21 VSS.t74 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X295 hgu_cdac_8bit_array_3.drv<15:0>.t22 d<4>.t17 VSS.t401 VSS.t400 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X296 hgu_cdac_8bit_array_2.drv<7:0>.t11 db<3>.t9 VREF.t80 VDD.t80 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X297 hgu_cdac_8bit_array_3.drv<7:0>.t7 d<3>.t9 VSS.t457 VSS.t456 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X298 hgu_cdac_8bit_array_2.drv<63:0>.t32 db<6>.t70 VREF.t60 VDD.t60 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X299 VREF.t145 d<2>.t5 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t1 VDD.t145 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X300 VREF.t193 db<2>.t5 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t1 VDD.t192 sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X301 VSS.t267 d<6>.t75 hgu_cdac_8bit_array_3.drv<63:0>.t97 VSS.t266 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X302 hgu_cdac_8bit_array_3.drv<31:0>.t27 d<5>.t40 VREF.t21 VDD.t21 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X303 VSS.t183 db<6>.t71 hgu_cdac_8bit_array_2.drv<63:0>.t88 VSS.t182 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X304 VREF.t73 db<6>.t72 hgu_cdac_8bit_array_2.drv<63:0>.t31 VDD.t73 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X305 hgu_cdac_8bit_array_3.drv<7:0>.t6 d<3>.t10 VSS.t455 VSS.t454 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X306 hgu_cdac_8bit_array_2.drv<63:0>.t30 db<6>.t73 VREF.t123 VDD.t123 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X307 hgu_cdac_8bit_array_3.drv<63:0>.t53 d<6>.t76 VREF.t71 VDD.t71 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X308 VSS.t27 db<5>.t34 hgu_cdac_8bit_array_2.drv<31:0>.t46 VSS.t26 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X309 VREF.t94 db<5>.t35 hgu_cdac_8bit_array_2.drv<31:0>.t27 VDD.t94 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X310 VREF.t50 d<6>.t77 hgu_cdac_8bit_array_3.drv<63:0>.t52 VDD.t50 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X311 hgu_cdac_8bit_array_3.drv<31:0>.t26 d<5>.t41 VREF.t101 VDD.t101 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X312 hgu_cdac_8bit_array_2.drv<63:0>.t87 db<6>.t74 VSS.t361 VSS.t360 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X313 hgu_cdac_8bit_array_3.drv<63:0>.t51 d<6>.t78 VREF.t100 VDD.t100 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X314 VSS.t433 db<6>.t75 hgu_cdac_8bit_array_2.drv<63:0>.t86 VSS.t432 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X315 hgu_cdac_8bit_array_2.drv<31:0>.t26 db<5>.t36 VREF.t95 VDD.t95 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X316 VSS.t435 db<6>.t76 hgu_cdac_8bit_array_2.drv<63:0>.t85 VSS.t434 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X317 VREF.t251 db<6>.t77 hgu_cdac_8bit_array_2.drv<63:0>.t29 VDD.t246 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X318 hgu_cdac_8bit_array_3.drv<63:0>.t96 d<6>.t79 VSS.t265 VSS.t264 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X319 VSS.t25 db<5>.t37 hgu_cdac_8bit_array_2.drv<31:0>.t45 VSS.t24 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X320 hgu_cdac_8bit_array_2.drv<7:0>.t10 db<3>.t10 VREF.t158 VDD.t158 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X321 VSS.t263 d<6>.t80 hgu_cdac_8bit_array_3.drv<63:0>.t95 VSS.t262 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X322 VREF.t199 db<5>.t38 hgu_cdac_8bit_array_2.drv<31:0>.t25 VDD.t198 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X323 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t0 db<2>.t6 VREF.t87 VDD.t87 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X324 VSS.t119 d<5>.t42 hgu_cdac_8bit_array_3.drv<31:0>.t50 VSS.t118 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X325 hgu_cdac_8bit_array_2.drv<63:0>.t84 db<6>.t78 VSS.t505 VSS.t504 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X326 hgu_cdac_8bit_array_3.drv<63:0>.t50 d<6>.t81 VREF.t20 VDD.t20 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X327 VREF.t204 db<6>.t79 hgu_cdac_8bit_array_2.drv<63:0>.t28 VDD.t203 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X328 VSS.t421 db<6>.t80 hgu_cdac_8bit_array_2.drv<63:0>.t83 VSS.t420 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X329 VSS.t261 d<6>.t82 hgu_cdac_8bit_array_3.drv<63:0>.t14 VSS.t260 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X330 VREF.t196 db<6>.t81 hgu_cdac_8bit_array_2.drv<63:0>.t27 VDD.t195 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X331 hgu_cdac_8bit_array_3.drv<15:0>.t7 d<4>.t18 VREF.t29 VDD.t29 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X332 hgu_cdac_8bit_array_2.drv<31:0>.t44 db<5>.t39 VSS.t23 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X333 VREF.t197 db<6>.t82 hgu_cdac_8bit_array_2.drv<63:0>.t26 VDD.t196 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X334 VREF.t120 d<4>.t19 hgu_cdac_8bit_array_3.drv<15:0>.t6 VDD.t120 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X335 hgu_cdac_8bit_array_2.drv<63:0>.t82 db<6>.t83 VSS.t195 VSS.t194 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X336 VREF.t37 d<5>.t43 hgu_cdac_8bit_array_3.drv<31:0>.t25 VDD.t37 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X337 hgu_cdac_8bit_array_3.drv<7:0>.t12 d<3>.t11 VREF.t229 VDD.t227 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X338 VSS.t197 db<6>.t84 hgu_cdac_8bit_array_2.drv<63:0>.t81 VSS.t196 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X339 VSS.t21 db<5>.t40 hgu_cdac_8bit_array_2.drv<31:0>.t63 VSS.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X340 VREF.t171 db<5>.t41 hgu_cdac_8bit_array_2.drv<31:0>.t24 VDD.t171 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X341 VREF.t75 d<6>.t83 hgu_cdac_8bit_array_3.drv<63:0>.t49 VDD.t75 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X342 VREF.t137 d<6>.t84 hgu_cdac_8bit_array_3.drv<63:0>.t48 VDD.t137 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X343 hgu_cdac_8bit_array_3.drv<31:0>.t24 d<5>.t44 VREF.t170 VDD.t170 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X344 VSS.t117 d<5>.t45 hgu_cdac_8bit_array_3.drv<31:0>.t49 VSS.t116 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X345 hgu_cdac_8bit_array_2.drv<63:0>.t25 db<6>.t85 VREF.t27 VDD.t27 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X346 VREF.t117 db<4>.t21 hgu_cdac_8bit_array_2.drv<15:0>.t5 VDD.t117 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X347 VSS.t259 d<6>.t85 hgu_cdac_8bit_array_3.drv<63:0>.t13 VSS.t258 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X348 VSS.t483 db<3>.t11 hgu_cdac_8bit_array_2.drv<7:0>.t6 VSS.t482 sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X349 hgu_cdac_8bit_array_2.drv<31:0>.t62 db<5>.t42 VSS.t19 VSS.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X350 VSS.t79 db<6>.t86 hgu_cdac_8bit_array_2.drv<63:0>.t80 VSS.t78 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X351 VREF.t172 db<3>.t12 hgu_cdac_8bit_array_2.drv<7:0>.t9 VDD.t172 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X352 VREF.t187 d<6>.t86 hgu_cdac_8bit_array_3.drv<63:0>.t47 VDD.t186 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X353 hgu_cdac_8bit_array_3.drv<63:0>.t12 d<6>.t87 VSS.t257 VSS.t256 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X354 VSS.t115 d<5>.t46 hgu_cdac_8bit_array_3.drv<31:0>.t48 VSS.t114 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X355 hgu_cdac_8bit_array_2.drv<63:0>.t24 db<6>.t87 VREF.t124 VDD.t124 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X356 VREF.t131 db<4>.t22 hgu_cdac_8bit_array_2.drv<15:0>.t4 VDD.t131 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X357 VSS.t453 d<3>.t12 hgu_cdac_8bit_array_3.drv<7:0>.t2 VSS.t452 sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X358 hgu_cdac_8bit_array_3.drv<63:0>.t11 d<6>.t88 VSS.t255 VSS.t254 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X359 hgu_cdac_8bit_array_2.drv<63:0>.t23 db<6>.t88 VREF.t125 VDD.t125 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X360 hgu_cdac_8bit_array_3.drv<63:0>.t46 d<6>.t89 VREF.t226 VDD.t225 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X361 VREF.t115 d<4>.t20 hgu_cdac_8bit_array_3.drv<15:0>.t5 VDD.t115 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X362 hgu_cdac_8bit_array_3.drv<31:0>.t23 d<5>.t47 VREF.t54 VDD.t54 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X363 VSS.t405 db<6>.t89 hgu_cdac_8bit_array_2.drv<63:0>.t79 VSS.t404 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X364 hgu_cdac_8bit_array_2.drv<15:0>.t20 db<4>.t23 VSS.t359 VSS.t358 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X365 VSS.t441 d<4>.t21 hgu_cdac_8bit_array_3.drv<15:0>.t21 VSS.t440 sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X366 hgu_cdac_8bit_array_3.drv<63:0>.t10 d<6>.t90 VSS.t253 VSS.t252 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X367 hgu_cdac_8bit_array_2.drv<31:0>.t23 db<5>.t43 VREF.t246 VDD.t241 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X368 hgu_cdac_8bit_array_3.drv<31:0>.t47 d<5>.t48 VSS.t113 VSS.t112 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X369 VSS.t451 d<3>.t13 hgu_cdac_8bit_array_3.drv<7:0>.t1 VSS.t450 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X370 VREF.t12 d<6>.t91 hgu_cdac_8bit_array_3.drv<63:0>.t45 VDD.t12 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X371 hgu_cdac_8bit_array_2.drv<63:0>.t78 db<6>.t90 VSS.t407 VSS.t406 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X372 hgu_cdac_8bit_array_3.drv<63:0>.t121 d<6>.t92 VSS.t251 VSS.t250 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X373 hgu_cdac_8bit_array_3.drv<63:0>.t44 d<6>.t93 VREF.t99 VDD.t99 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X374 VREF.t10 d<4>.t22 hgu_cdac_8bit_array_3.drv<15:0>.t4 VDD.t10 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X375 hgu_cdac_8bit_array_2.drv<63:0>.t22 db<6>.t91 VREF.t209 VDD.t208 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X376 VREF.t132 d<6>.t94 hgu_cdac_8bit_array_3.drv<63:0>.t43 VDD.t132 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X377 hgu_cdac_8bit_array_3.drv<15:0>.t20 d<4>.t23 VSS.t467 VSS.t466 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X378 VSS.t427 db<6>.t92 hgu_cdac_8bit_array_2.drv<63:0>.t77 VSS.t426 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X379 VSS.t249 d<6>.t95 hgu_cdac_8bit_array_3.drv<63:0>.t120 VSS.t248 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X380 hgu_cdac_8bit_array_2.drv<31:0>.t61 db<5>.t44 VSS.t17 VSS.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X381 hgu_cdac_8bit_array_2.drv<63:0>.t21 db<6>.t93 VREF.t84 VDD.t84 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X382 hgu_cdac_8bit_array_2.drv<31:0>.t22 db<5>.t45 VREF.t173 VDD.t173 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X383 VSS.t189 db<6>.t94 hgu_cdac_8bit_array_2.drv<63:0>.t76 VSS.t188 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X384 hgu_cdac_8bit_array_3.drv<31:0>.t61 d<5>.t49 VSS.t111 VSS.t110 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X385 VREF.t109 db<6>.t95 hgu_cdac_8bit_array_2.drv<63:0>.t20 VDD.t109 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X386 VREF.t4 db<5>.t46 hgu_cdac_8bit_array_2.drv<31:0>.t21 VDD.t4 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X387 VREF.t111 d<6>.t96 hgu_cdac_8bit_array_3.drv<63:0>.t42 VDD.t111 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X388 hgu_cdac_8bit_array_2.drv<7:0>.t5 db<3>.t13 VSS.t481 VSS.t480 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X389 hgu_cdac_8bit_array_2.drv<31:0>.t20 db<5>.t47 VREF.t133 VDD.t133 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X390 VSS.t413 db<2>.t7 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t4 VSS.t412 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X391 hgu_cdac_8bit_array_2.drv<63:0>.t19 db<6>.t96 VREF.t110 VDD.t110 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X392 VREF.t245 db<1>.t3 hgu_cdac_8bit_array_2.drv<1:0>.t0 VDD.t240 sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X393 VSS.t247 d<6>.t97 hgu_cdac_8bit_array_3.drv<63:0>.t119 VSS.t246 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X394 hgu_cdac_8bit_array_2.drv<63:0>.t18 db<6>.t97 VREF.t212 VDD.t211 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X395 hgu_cdac_8bit_array_2.drv<63:0>.t17 db<6>.t98 VREF.t213 VDD.t212 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X396 VREF.t222 db<3>.t14 hgu_cdac_8bit_array_2.drv<7:0>.t8 VDD.t221 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X397 hgu_cdac_8bit_array_2.drv<63:0>.t16 db<6>.t99 VREF.t18 VDD.t18 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X398 hgu_cdac_8bit_array_3.drv<63:0>.t41 d<6>.t98 VREF.t227 VDD.t226 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X399 hgu_cdac_8bit_array_3.drv<63:0>.t40 d<6>.t99 VREF.t154 VDD.t154 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X400 hgu_cdac_8bit_array_2.drv<31:0>.t19 db<5>.t48 VREF.t51 VDD.t51 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X401 VREF.t90 d<5>.t50 hgu_cdac_8bit_array_3.drv<31:0>.t22 VDD.t90 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X402 VSS.t477 d<2>.t6 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t4 VSS.t476 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X403 VSS.t65 db<6>.t100 hgu_cdac_8bit_array_2.drv<63:0>.t75 VSS.t64 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X404 hgu_cdac_8bit_array_3.drv<31:0>.t60 d<5>.t51 VSS.t109 VSS.t108 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X405 hgu_cdac_8bit_array_2.drv<63:0>.t15 db<6>.t101 VREF.t7 VDD.t7 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X406 VREF.t210 db<4>.t24 hgu_cdac_8bit_array_2.drv<15:0>.t3 VDD.t209 sky130_fd_pr__pfet_01v8_lvt ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.35
X407 hgu_cdac_8bit_array_2.drv<31:0>.t60 db<5>.t49 VSS.t15 VSS.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X408 hgu_cdac_8bit_array_2.drv<63:0>.t14 db<6>.t102 VREF.t8 VDD.t8 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X409 hgu_cdac_8bit_array_3.drv<63:0>.t39 d<6>.t100 VREF.t167 VDD.t167 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X410 hgu_cdac_8bit_array_3.drv<31:0>.t21 d<5>.t52 VREF.t74 VDD.t74 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X411 VSS.t381 db<6>.t103 hgu_cdac_8bit_array_2.drv<63:0>.t74 VSS.t380 sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X412 hgu_cdac_8bit_array_2.drv<15:0>.t2 db<4>.t25 VREF.t237 VDD.t232 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X413 hgu_cdac_8bit_array_3.drv<63:0>.t38 d<6>.t101 VREF.t11 VDD.t11 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X414 hgu_cdac_8bit_array_3.drv<63:0>.t118 d<6>.t102 VSS.t245 VSS.t244 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X415 VSS.t383 db<6>.t104 hgu_cdac_8bit_array_2.drv<63:0>.t73 VSS.t382 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X416 hgu_cdac_8bit_array_2.drv<31:0>.t18 db<5>.t50 VREF.t224 VDD.t223 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X417 hgu_cdac_8bit_array_3.drv<31:0>.t59 d<5>.t53 VSS.t107 VSS.t106 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X418 VSS.t243 d<6>.t103 hgu_cdac_8bit_array_3.drv<63:0>.t117 VSS.t242 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X419 VREF.t58 db<6>.t105 hgu_cdac_8bit_array_2.drv<63:0>.t13 VDD.t58 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X420 hgu_cdac_8bit_array_3.drv<1:0>.t0 d<1> VREF.t185 VDD.t184 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X421 hgu_cdac_8bit_array_3.drv<63:0>.t4 d<6>.t104 VSS.t241 VSS.t240 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X422 VSS.t209 db<4>.t26 hgu_cdac_8bit_array_2.drv<15:0>.t19 VSS.t208 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X423 VSS.t13 db<5>.t51 hgu_cdac_8bit_array_2.drv<31:0>.t59 VSS.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X424 hgu_cdac_8bit_array_3.drv<15:0>.t3 d<4>.t24 VREF.t105 VDD.t105 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X425 VREF.t59 db<6>.t106 hgu_cdac_8bit_array_2.drv<63:0>.t12 VDD.t59 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X426 hgu_cdac_8bit_array_3.drv<31:0>.t20 d<5>.t54 VREF.t220 VDD.t219 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X427 hgu_cdac_8bit_array_2.drv<63:0>.t72 db<6>.t107 VSS.t163 VSS.t162 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X428 VSS.t165 db<6>.t108 hgu_cdac_8bit_array_2.drv<63:0>.t71 VSS.t164 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X429 hgu_cdac_8bit_array_2.drv<63:0>.t11 db<6>.t109 VREF.t214 VDD.t213 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X430 hgu_cdac_8bit_array_2.drv<31:0>.t17 db<5>.t52 VREF.t200 VDD.t199 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X431 hgu_cdac_8bit_array_3.drv<63:0>.t37 d<6>.t105 VREF.t69 VDD.t69 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X432 hgu_cdac_8bit_array_3.drv<15:0>.t2 d<4>.t25 VREF.t49 VDD.t49 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X433 hgu_cdac_8bit_array_2.drv<31:0>.t53 db<5>.t53 VSS.t11 VSS.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X434 VREF.t215 db<6>.t110 hgu_cdac_8bit_array_2.drv<63:0>.t10 VDD.t214 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X435 hgu_cdac_8bit_array_3.drv<63:0>.t3 d<6>.t106 VSS.t239 VSS.t238 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X436 VSS.t205 db<4>.t27 hgu_cdac_8bit_array_2.drv<15:0>.t18 VSS.t204 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X437 hgu_cdac_8bit_array_2.drv<31:0>.t16 db<5>.t54 VREF.t194 VDD.t193 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X438 VSS.t9 db<5>.t55 hgu_cdac_8bit_array_2.drv<31:0>.t52 VSS.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X439 hgu_cdac_8bit_array_3.drv<15:0>.t19 d<4>.t26 VSS.t495 VSS.t494 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X440 VREF.t79 d<6>.t107 hgu_cdac_8bit_array_3.drv<63:0>.t36 VDD.t79 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X441 VSS.t365 d<4>.t27 hgu_cdac_8bit_array_3.drv<15:0>.t18 VSS.t364 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X442 hgu_cdac_8bit_array_2.drv<63:0>.t70 db<6>.t111 VSS.t367 VSS.t366 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X443 hgu_cdac_8bit_array_3.drv<7:0>.t0 d<3>.t14 VSS.t449 VSS.t448 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.35
X444 VSS.t105 d<5>.t55 hgu_cdac_8bit_array_3.drv<31:0>.t58 VSS.t104 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X445 hgu_cdac_8bit_array_2.drv<63:0>.t9 db<6>.t112 VREF.t130 VDD.t130 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X446 VREF.t113 db<4>.t28 hgu_cdac_8bit_array_2.drv<15:0>.t1 VDD.t113 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X447 VSS.t237 d<6>.t108 hgu_cdac_8bit_array_3.drv<63:0>.t2 VSS.t236 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X448 VSS.t235 d<6>.t109 hgu_cdac_8bit_array_3.drv<63:0>.t1 VSS.t234 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X449 VSS.t479 db<3>.t15 hgu_cdac_8bit_array_2.drv<7:0>.t4 VSS.t478 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X450 hgu_cdac_8bit_array_3.drv<31:0>.t57 d<5>.t56 VSS.t103 VSS.t102 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X451 hgu_cdac_8bit_array_3.drv<63:0>.t35 d<6>.t110 VREF.t102 VDD.t102 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X452 VSS.t81 db<6>.t113 hgu_cdac_8bit_array_2.drv<63:0>.t69 VSS.t80 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X453 VREF.t139 d<6>.t111 hgu_cdac_8bit_array_3.drv<63:0>.t34 VDD.t139 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X454 VREF.t182 d<5>.t57 hgu_cdac_8bit_array_3.drv<31:0>.t19 VDD.t182 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X455 hgu_cdac_8bit_array_2.drv<63:0>.t68 db<6>.t114 VSS.t83 VSS.t82 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X456 hgu_cdac_8bit_array_3.drv<7:0>.t11 d<3>.t15 VREF.t228 VDD.t88 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X457 hgu_cdac_8bit_array_2.drv<63:0>.t8 db<6>.t115 VREF.t247 VDD.t242 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X458 VREF.t81 db<4>.t29 hgu_cdac_8bit_array_2.drv<15:0>.t0 VDD.t81 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X459 VSS.t7 db<5>.t56 hgu_cdac_8bit_array_2.drv<31:0>.t51 VSS.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.35
X460 VSS.t233 d<6>.t112 hgu_cdac_8bit_array_3.drv<63:0>.t0 VSS.t232 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X461 hgu_cdac_8bit_array_3.drv<31:0>.t18 d<5>.t58 VREF.t166 VDD.t166 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X462 hgu_cdac_8bit_array_3.drv<63:0>.t33 d<6>.t113 VREF.t236 VDD.t231 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X463 hgu_cdac_8bit_array_3.drv<63:0>.t32 d<6>.t114 VREF.t134 VDD.t134 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X464 VSS.t499 db<6>.t116 hgu_cdac_8bit_array_2.drv<63:0>.t67 VSS.t498 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X465 hgu_cdac_8bit_array_2.drv<15:0>.t17 db<4>.t30 VSS.t415 VSS.t414 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X466 VSS.t387 d<4>.t28 hgu_cdac_8bit_array_3.drv<15:0>.t17 VSS.t386 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X467 hgu_cdac_8bit_array_3.drv<63:0>.t19 d<6>.t115 VSS.t231 VSS.t230 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X468 VSS.t5 db<5>.t57 hgu_cdac_8bit_array_2.drv<31:0>.t50 VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X469 hgu_cdac_8bit_array_3.drv<31:0>.t63 d<5>.t59 VSS.t101 VSS.t100 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X470 VREF.t15 db<6>.t117 hgu_cdac_8bit_array_2.drv<63:0>.t7 VDD.t15 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X471 hgu_cdac_8bit_array_3.drv<63:0>.t31 d<6>.t116 VREF.t89 VDD.t89 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X472 VSS.t229 d<6>.t117 hgu_cdac_8bit_array_3.drv<63:0>.t18 VSS.t228 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X473 hgu_cdac_8bit_array_2.drv<15:0>.t16 db<4>.t31 VSS.t77 VSS.t76 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X474 VREF.t201 db<5>.t58 hgu_cdac_8bit_array_2.drv<31:0>.t15 VDD.t200 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X475 VSS.t179 d<4>.t29 hgu_cdac_8bit_array_3.drv<15:0>.t16 VSS.t178 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X476 hgu_cdac_8bit_array_2.drv<63:0>.t6 db<6>.t118 VREF.t16 VDD.t16 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X477 VREF.t26 d<4>.t30 hgu_cdac_8bit_array_3.drv<15:0>.t1 VDD.t26 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X478 hgu_cdac_8bit_array_3.drv<63:0>.t17 d<6>.t118 VSS.t227 VSS.t226 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X479 VSS.t225 d<6>.t119 hgu_cdac_8bit_array_3.drv<63:0>.t16 VSS.t224 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X480 VREF.t114 db<6>.t119 hgu_cdac_8bit_array_2.drv<63:0>.t5 VDD.t114 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X481 hgu_cdac_8bit_array_2.drv<63:0>.t66 db<6>.t120 VSS.t211 VSS.t210 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X482 VREF.t216 db<6>.t121 hgu_cdac_8bit_array_2.drv<63:0>.t4 VDD.t215 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X483 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t0 d<2>.t7 VREF.t186 VDD.t185 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X484 VREF.t39 d<6>.t120 hgu_cdac_8bit_array_3.drv<63:0>.t30 VDD.t39 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X485 VREF.t151 db<5>.t59 hgu_cdac_8bit_array_2.drv<31:0>.t14 VDD.t151 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X486 VSS.t223 d<6>.t121 hgu_cdac_8bit_array_3.drv<63:0>.t15 VSS.t222 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X487 hgu_cdac_8bit_array_2.drv<63:0>.t65 db<6>.t122 VSS.t437 VSS.t436 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X488 hgu_cdac_8bit_array_2.drv<31:0>.t49 db<5>.t60 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X489 hgu_cdac_8bit_array_2.drv<63:0>.t3 db<6>.t123 VREF.t72 VDD.t72 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X490 hgu_cdac_8bit_array_3.drv<63:0>.t29 d<6>.t122 VREF.t3 VDD.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X491 VREF.t207 d<4>.t31 hgu_cdac_8bit_array_3.drv<15:0>.t0 VDD.t206 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X492 hgu_cdac_8bit_array_3.drv<31:0>.t17 d<5>.t60 VREF.t36 VDD.t36 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.35
X493 VSS.t181 db<6>.t124 hgu_cdac_8bit_array_2.drv<63:0>.t64 VSS.t180 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X494 VREF.t242 db<6>.t125 hgu_cdac_8bit_array_2.drv<63:0>.t2 VDD.t237 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X495 VREF.t150 d<6>.t123 hgu_cdac_8bit_array_3.drv<63:0>.t28 VDD.t150 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X496 hgu_cdac_8bit_array_2.drv<31:0>.t11 db<5>.t61 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X497 hgu_cdac_8bit_array_2.drv<31:0>.t13 db<5>.t62 VREF.t107 VDD.t107 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X498 hgu_cdac_8bit_array_3.drv<63:0>.t27 d<6>.t124 VREF.t24 VDD.t24 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X499 VREF.t68 d<5>.t61 hgu_cdac_8bit_array_3.drv<31:0>.t16 VDD.t68 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X500 hgu_cdac_8bit_array_3.drv<63:0>.t111 d<6>.t125 VSS.t221 VSS.t220 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X501 hgu_cdac_8bit_array_2.drv<63:0>.t1 db<6>.t126 VREF.t243 VDD.t238 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X502 VREF.t141 db<6>.t127 hgu_cdac_8bit_array_2.drv<63:0>.t0 VDD.t141 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X503 VREF.t118 db<5>.t63 hgu_cdac_8bit_array_2.drv<31:0>.t12 VDD.t118 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X504 VSS.t99 d<5>.t62 hgu_cdac_8bit_array_3.drv<31:0>.t62 VSS.t98 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X505 hgu_cdac_8bit_array_3.drv<63:0>.t110 d<6>.t126 VSS.t219 VSS.t218 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=0.35
X506 hgu_cdac_8bit_array_3.drv<63:0>.t26 d<6>.t127 VREF.t165 VDD.t165 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
X507 hgu_cdac_8bit_array_3.drv<31:0>.t15 d<5>.t63 VREF.t244 VDD.t239 sky130_fd_pr__pfet_01v8_lvt ad=0.122 pd=1.13 as=0.122 ps=1.13 w=0.84 l=0.35
R0 d<3>.n1 d<3>.n0 88.1376
R1 d<3>.n2 d<3>.n1 88.1376
R2 d<3>.n3 d<3>.n2 88.1376
R3 d<3>.n4 d<3>.n3 88.1376
R4 d<3>.n5 d<3>.n4 88.1376
R5 d<3>.n6 d<3>.n5 88.1376
R6 d<3>.n7 d<3>.n6 88.1376
R7 d<3>.n0 d<3>.t7 69.5462
R8 d<3>.n1 d<3>.t5 69.5462
R9 d<3>.n2 d<3>.t0 69.5462
R10 d<3>.n3 d<3>.t15 69.5462
R11 d<3>.n4 d<3>.t8 69.5462
R12 d<3>.n5 d<3>.t6 69.5462
R13 d<3>.n6 d<3>.t1 69.5462
R14 d<3>.n7 d<3>.t11 69.5462
R15 d<3>.n0 d<3>.t12 59.9062
R16 d<3>.n1 d<3>.t9 59.9062
R17 d<3>.n2 d<3>.t3 59.9062
R18 d<3>.n3 d<3>.t2 59.9062
R19 d<3>.n4 d<3>.t13 59.9062
R20 d<3>.n5 d<3>.t10 59.9062
R21 d<3>.n6 d<3>.t4 59.9062
R22 d<3>.n7 d<3>.t14 59.9062
R23 d<3> d<3>.n7 24.1005
R24 hgu_cdac_8bit_array_3.drv<7:0>.n2 hgu_cdac_8bit_array_3.drv<7:0>.t9 41.4291
R25 hgu_cdac_8bit_array_3.drv<7:0>.n2 hgu_cdac_8bit_array_3.drv<7:0>.t10 41.4291
R26 hgu_cdac_8bit_array_3.drv<7:0>.n3 hgu_cdac_8bit_array_3.drv<7:0>.t1 41.4291
R27 hgu_cdac_8bit_array_3.drv<7:0>.n3 hgu_cdac_8bit_array_3.drv<7:0>.t6 41.4291
R28 hgu_cdac_8bit_array_3.drv<7:0>.n4 hgu_cdac_8bit_array_3.drv<7:0>.t8 41.4291
R29 hgu_cdac_8bit_array_3.drv<7:0>.n4 hgu_cdac_8bit_array_3.drv<7:0>.t0 41.4291
R30 hgu_cdac_8bit_array_3.drv<7:0>.n0 hgu_cdac_8bit_array_3.drv<7:0>.t2 41.4291
R31 hgu_cdac_8bit_array_3.drv<7:0>.n0 hgu_cdac_8bit_array_3.drv<7:0>.t7 41.4291
R32 hgu_cdac_8bit_array_3.drv<7:0>.n5 hgu_cdac_8bit_array_3.drv<7:0>.t5 34.0065
R33 hgu_cdac_8bit_array_3.drv<7:0>.n5 hgu_cdac_8bit_array_3.drv<7:0>.t11 34.0065
R34 hgu_cdac_8bit_array_3.drv<7:0>.n6 hgu_cdac_8bit_array_3.drv<7:0>.t13 34.0065
R35 hgu_cdac_8bit_array_3.drv<7:0>.n6 hgu_cdac_8bit_array_3.drv<7:0>.t15 34.0065
R36 hgu_cdac_8bit_array_3.drv<7:0>.n9 hgu_cdac_8bit_array_3.drv<7:0>.t4 34.0065
R37 hgu_cdac_8bit_array_3.drv<7:0>.n9 hgu_cdac_8bit_array_3.drv<7:0>.t12 34.0065
R38 hgu_cdac_8bit_array_3.drv<7:0>.n7 hgu_cdac_8bit_array_3.drv<7:0>.t14 34.0065
R39 hgu_cdac_8bit_array_3.drv<7:0>.n7 hgu_cdac_8bit_array_3.drv<7:0>.t3 34.0065
R40 hgu_cdac_8bit_array_3.drv<7:0>.n1 hgu_cdac_8bit_array_3.drv<7:0>.n4 11.883
R41 hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_8bit_array_3.drv<7:0>.n8 8.35989
R42 hgu_cdac_8bit_array_3.drv<7:0>.n8 hgu_cdac_8bit_array_3.drv<7:0>.n0 2.68086
R43 hgu_cdac_8bit_array_3.drv<7:0>.n0 hgu_cdac_8bit_array_3.drv<7:0>.n2 0.957397
R44 hgu_cdac_8bit_array_3.drv<7:0>.n2 hgu_cdac_8bit_array_3.drv<7:0>.n3 0.957397
R45 hgu_cdac_8bit_array_3.drv<7:0>.n0 hgu_cdac_8bit_array_3.drv<7:0>.n7 0.892799
R46 hgu_cdac_8bit_array_3.drv<7:0>.n4 hgu_cdac_8bit_array_3.drv<7:0>.n9 0.85856
R47 hgu_cdac_8bit_array_3.drv<7:0>.n3 hgu_cdac_8bit_array_3.drv<7:0>.n6 0.85856
R48 hgu_cdac_8bit_array_3.drv<7:0>.n2 hgu_cdac_8bit_array_3.drv<7:0>.n5 0.85856
R49 hgu_cdac_8bit_array_3.drv<7:0> hgu_cdac_8bit_array_3.drv<7:0>.n1 0.728175
R50 hgu_cdac_8bit_array_3.drv<7:0>.n1 hgu_cdac_8bit_array_3.drv<7:0> 0.686479
R51 VREF.n254 VREF.n253 37.9198
R52 VREF VREF.n188 36.77
R53 VREF.n0 VREF.t249 34.4208
R54 VREF.n1 VREF.t185 34.4208
R55 VREF.n2 VREF.t184 34.4208
R56 VREF.n3 VREF.t30 34.4208
R57 VREF.n6 VREF.t223 34.4208
R58 VREF.n7 VREF.t229 34.4208
R59 VREF.n14 VREF.t231 34.4208
R60 VREF.n15 VREF.t218 34.4208
R61 VREF.n30 VREF.t70 34.4208
R62 VREF.n31 VREF.t36 34.4208
R63 VREF.n62 VREF.t176 34.4208
R64 VREF.n63 VREF.t217 34.4208
R65 VREF.n254 VREF.t103 34.4208
R66 VREF VREF.t108 34.3987
R67 VREF VREF.t155 34.3987
R68 VREF VREF.t245 34.3987
R69 VREF VREF.t87 34.3987
R70 VREF VREF.t193 34.3987
R71 VREF VREF.t88 34.3987
R72 VREF VREF.t35 34.3987
R73 VREF VREF.t219 34.3987
R74 VREF VREF.t210 34.3987
R75 VREF VREF.t162 34.3987
R76 VREF VREF.t168 34.3987
R77 VREF VREF.t7 34.3987
R78 VREF VREF.t106 34.3987
R79 VREF.n130 VREF.t181 34.0065
R80 VREF.n130 VREF.t250 34.0065
R81 VREF.n134 VREF.t80 34.0065
R82 VREF.n134 VREF.t147 34.0065
R83 VREF.n136 VREF.t153 34.0065
R84 VREF.n136 VREF.t172 34.0065
R85 VREF.n138 VREF.t158 34.0065
R86 VREF.n138 VREF.t222 34.0065
R87 VREF.n142 VREF.t160 34.0065
R88 VREF.n142 VREF.t81 34.0065
R89 VREF.n144 VREF.t67 34.0065
R90 VREF.n144 VREF.t178 34.0065
R91 VREF.n146 VREF.t248 34.0065
R92 VREF.n146 VREF.t113 34.0065
R93 VREF.n148 VREF.t237 34.0065
R94 VREF.n148 VREF.t131 34.0065
R95 VREF.n150 VREF.t159 34.0065
R96 VREF.n150 VREF.t1 34.0065
R97 VREF.n152 VREF.t112 34.0065
R98 VREF.n152 VREF.t117 34.0065
R99 VREF.n154 VREF.t41 34.0065
R100 VREF.n154 VREF.t253 34.0065
R101 VREF.n158 VREF.t56 34.0065
R102 VREF.n158 VREF.t46 34.0065
R103 VREF.n160 VREF.t173 34.0065
R104 VREF.n160 VREF.t138 34.0065
R105 VREF.n162 VREF.t107 34.0065
R106 VREF.n162 VREF.t94 34.0065
R107 VREF.n164 VREF.t246 34.0065
R108 VREF.n164 VREF.t97 34.0065
R109 VREF.n166 VREF.t142 34.0065
R110 VREF.n166 VREF.t91 34.0065
R111 VREF.n168 VREF.t51 34.0065
R112 VREF.n168 VREF.t171 34.0065
R113 VREF.n170 VREF.t65 34.0065
R114 VREF.n170 VREF.t161 34.0065
R115 VREF.n172 VREF.t133 34.0065
R116 VREF.n172 VREF.t199 34.0065
R117 VREF.n174 VREF.t200 34.0065
R118 VREF.n174 VREF.t14 34.0065
R119 VREF.n176 VREF.t174 34.0065
R120 VREF.n176 VREF.t151 34.0065
R121 VREF.n178 VREF.t224 34.0065
R122 VREF.n178 VREF.t92 34.0065
R123 VREF.n180 VREF.t163 34.0065
R124 VREF.n180 VREF.t201 34.0065
R125 VREF.n182 VREF.t104 34.0065
R126 VREF.n182 VREF.t4 34.0065
R127 VREF.n184 VREF.t95 34.0065
R128 VREF.n184 VREF.t98 34.0065
R129 VREF.n186 VREF.t194 34.0065
R130 VREF.n186 VREF.t118 34.0065
R131 VREF.n190 VREF.t31 34.0065
R132 VREF.n190 VREF.t38 34.0065
R133 VREF.n192 VREF.t212 34.0065
R134 VREF.n192 VREF.t204 34.0065
R135 VREF.n194 VREF.t209 34.0065
R136 VREF.n194 VREF.t22 34.0065
R137 VREF.n196 VREF.t72 34.0065
R138 VREF.n196 VREF.t73 34.0065
R139 VREF.n198 VREF.t125 34.0065
R140 VREF.n198 VREF.t66 34.0065
R141 VREF.n200 VREF.t16 34.0065
R142 VREF.n200 VREF.t59 34.0065
R143 VREF.n202 VREF.t213 34.0065
R144 VREF.n202 VREF.t197 34.0065
R145 VREF.n204 VREF.t40 34.0065
R146 VREF.n204 VREF.t195 34.0065
R147 VREF.n206 VREF.t84 34.0065
R148 VREF.n206 VREF.t251 34.0065
R149 VREF.n208 VREF.t198 34.0065
R150 VREF.n208 VREF.t85 34.0065
R151 VREF.n210 VREF.t203 34.0065
R152 VREF.n210 VREF.t114 34.0065
R153 VREF.n212 VREF.t8 34.0065
R154 VREF.n212 VREF.t238 34.0065
R155 VREF.n214 VREF.t62 34.0065
R156 VREF.n214 VREF.t15 34.0065
R157 VREF.n216 VREF.t18 34.0065
R158 VREF.n216 VREF.t208 34.0065
R159 VREF.n218 VREF.t123 34.0065
R160 VREF.n218 VREF.t239 34.0065
R161 VREF.n220 VREF.t214 34.0065
R162 VREF.n220 VREF.t242 34.0065
R163 VREF.n222 VREF.t60 34.0065
R164 VREF.n222 VREF.t82 34.0065
R165 VREF.n224 VREF.t179 34.0065
R166 VREF.n224 VREF.t216 34.0065
R167 VREF.n226 VREF.t247 34.0065
R168 VREF.n226 VREF.t240 34.0065
R169 VREF.n228 VREF.t126 34.0065
R170 VREF.n228 VREF.t190 34.0065
R171 VREF.n230 VREF.t130 34.0065
R172 VREF.n230 VREF.t109 34.0065
R173 VREF.n232 VREF.t124 34.0065
R174 VREF.n232 VREF.t141 34.0065
R175 VREF.n234 VREF.t148 34.0065
R176 VREF.n234 VREF.t156 34.0065
R177 VREF.n236 VREF.t27 34.0065
R178 VREF.n236 VREF.t34 34.0065
R179 VREF.n238 VREF.t211 34.0065
R180 VREF.n238 VREF.t86 34.0065
R181 VREF.n240 VREF.t243 34.0065
R182 VREF.n240 VREF.t76 34.0065
R183 VREF.n242 VREF.t25 34.0065
R184 VREF.n242 VREF.t119 34.0065
R185 VREF.n244 VREF.t83 34.0065
R186 VREF.n244 VREF.t215 34.0065
R187 VREF.n246 VREF.t157 34.0065
R188 VREF.n246 VREF.t175 34.0065
R189 VREF.n248 VREF.t241 34.0065
R190 VREF.n248 VREF.t58 34.0065
R191 VREF.n250 VREF.t110 34.0065
R192 VREF.n250 VREF.t196 34.0065
R193 VREF.n4 VREF.t186 34.0065
R194 VREF.n4 VREF.t145 34.0065
R195 VREF.n8 VREF.t232 34.0065
R196 VREF.n8 VREF.t234 34.0065
R197 VREF.n10 VREF.t228 34.0065
R198 VREF.n10 VREF.t230 34.0065
R199 VREF.n12 VREF.t233 34.0065
R200 VREF.n12 VREF.t235 34.0065
R201 VREF.n16 VREF.t183 34.0065
R202 VREF.n16 VREF.t202 34.0065
R203 VREF.n18 VREF.t180 34.0065
R204 VREF.n18 VREF.t120 34.0065
R205 VREF.n20 VREF.t49 34.0065
R206 VREF.n20 VREF.t10 34.0065
R207 VREF.n22 VREF.t57 34.0065
R208 VREF.n22 VREF.t207 34.0065
R209 VREF.n24 VREF.t105 34.0065
R210 VREF.n24 VREF.t115 34.0065
R211 VREF.n26 VREF.t29 34.0065
R212 VREF.n26 VREF.t26 34.0065
R213 VREF.n28 VREF.t2 34.0065
R214 VREF.n28 VREF.t144 34.0065
R215 VREF.n32 VREF.t54 34.0065
R216 VREF.n32 VREF.t19 34.0065
R217 VREF.n34 VREF.t6 34.0065
R218 VREF.n34 VREF.t17 34.0065
R219 VREF.n36 VREF.t42 34.0065
R220 VREF.n36 VREF.t37 34.0065
R221 VREF.n38 VREF.t28 34.0065
R222 VREF.n38 VREF.t206 34.0065
R223 VREF.n40 VREF.t244 34.0065
R224 VREF.n40 VREF.t182 34.0065
R225 VREF.n42 VREF.t220 34.0065
R226 VREF.n42 VREF.t136 34.0065
R227 VREF.n44 VREF.t61 34.0065
R228 VREF.n44 VREF.t55 34.0065
R229 VREF.n46 VREF.t74 34.0065
R230 VREF.n46 VREF.t164 34.0065
R231 VREF.n48 VREF.t127 34.0065
R232 VREF.n48 VREF.t53 34.0065
R233 VREF.n50 VREF.t149 34.0065
R234 VREF.n50 VREF.t63 34.0065
R235 VREF.n52 VREF.t101 34.0065
R236 VREF.n52 VREF.t78 34.0065
R237 VREF.n54 VREF.t116 34.0065
R238 VREF.n54 VREF.t68 34.0065
R239 VREF.n56 VREF.t21 34.0065
R240 VREF.n56 VREF.t146 34.0065
R241 VREF.n58 VREF.t170 34.0065
R242 VREF.n58 VREF.t252 34.0065
R243 VREF.n60 VREF.t166 34.0065
R244 VREF.n60 VREF.t90 34.0065
R245 VREF.n64 VREF.t5 34.0065
R246 VREF.n64 VREF.t52 34.0065
R247 VREF.n66 VREF.t24 34.0065
R248 VREF.n66 VREF.t50 34.0065
R249 VREF.n68 VREF.t11 34.0065
R250 VREF.n68 VREF.t187 34.0065
R251 VREF.n70 VREF.t0 34.0065
R252 VREF.n70 VREF.t43 34.0065
R253 VREF.n72 VREF.t154 34.0065
R254 VREF.n72 VREF.t137 34.0065
R255 VREF.n74 VREF.t169 34.0065
R256 VREF.n74 VREF.t47 34.0065
R257 VREF.n76 VREF.t143 34.0065
R258 VREF.n76 VREF.t12 34.0065
R259 VREF.n78 VREF.t69 34.0065
R260 VREF.n78 VREF.t96 34.0065
R261 VREF.n80 VREF.t9 34.0065
R262 VREF.n80 VREF.t39 34.0065
R263 VREF.n82 VREF.t236 34.0065
R264 VREF.n82 VREF.t129 34.0065
R265 VREF.n84 VREF.t20 34.0065
R266 VREF.n84 VREF.t152 34.0065
R267 VREF.n86 VREF.t102 34.0065
R268 VREF.n86 VREF.t111 34.0065
R269 VREF.n88 VREF.t100 34.0065
R270 VREF.n88 VREF.t188 34.0065
R271 VREF.n90 VREF.t140 34.0065
R272 VREF.n90 VREF.t132 34.0065
R273 VREF.n92 VREF.t89 34.0065
R274 VREF.n92 VREF.t191 34.0065
R275 VREF.n94 VREF.t23 34.0065
R276 VREF.n94 VREF.t44 34.0065
R277 VREF.n96 VREF.t134 34.0065
R278 VREF.n96 VREF.t192 34.0065
R279 VREF.n98 VREF.t99 34.0065
R280 VREF.n98 VREF.t122 34.0065
R281 VREF.n100 VREF.t3 34.0065
R282 VREF.n100 VREF.t221 34.0065
R283 VREF.n102 VREF.t226 34.0065
R284 VREF.n102 VREF.t64 34.0065
R285 VREF.n104 VREF.t45 34.0065
R286 VREF.n104 VREF.t48 34.0065
R287 VREF.n106 VREF.t121 34.0065
R288 VREF.n106 VREF.t33 34.0065
R289 VREF.n108 VREF.t128 34.0065
R290 VREF.n108 VREF.t177 34.0065
R291 VREF.n110 VREF.t165 34.0065
R292 VREF.n110 VREF.t139 34.0065
R293 VREF.n112 VREF.t13 34.0065
R294 VREF.n112 VREF.t189 34.0065
R295 VREF.n114 VREF.t32 34.0065
R296 VREF.n114 VREF.t79 34.0065
R297 VREF.n116 VREF.t167 34.0065
R298 VREF.n116 VREF.t77 34.0065
R299 VREF.n118 VREF.t225 34.0065
R300 VREF.n118 VREF.t135 34.0065
R301 VREF.n120 VREF.t227 34.0065
R302 VREF.n120 VREF.t75 34.0065
R303 VREF.n122 VREF.t71 34.0065
R304 VREF.n122 VREF.t205 34.0065
R305 VREF.n124 VREF.t93 34.0065
R306 VREF.n124 VREF.t150 34.0065
R307 VREF VREF.n62 22.2896
R308 VREF VREF.n156 22.1919
R309 VREF VREF.n140 13.6958
R310 VREF VREF.n30 11.7349
R311 VREF VREF.n14 5.60206
R312 VREF VREF.n132 4.188
R313 VREF VREF.n6 4.188
R314 VREF VREF.n128 3.80128
R315 VREF VREF.n126 3.48878
R316 VREF VREF.n0 2.98878
R317 VREF.n253 VREF.n252 2.8886
R318 VREF.n253 VREF 2.60824
R319 VREF VREF.n2 2.30128
R320 VREF.n128 VREF.n127 0.867688
R321 VREF.n132 VREF.n131 0.867688
R322 VREF.n140 VREF.n139 0.867688
R323 VREF.n156 VREF.n155 0.867688
R324 VREF.n188 VREF.n187 0.867688
R325 VREF.n252 VREF.n251 0.867688
R326 VREF.n2 VREF.n1 0.867688
R327 VREF.n6 VREF.n5 0.867688
R328 VREF.n14 VREF.n13 0.867688
R329 VREF.n30 VREF.n29 0.867688
R330 VREF.n62 VREF.n61 0.867688
R331 VREF.n254 VREF.n125 0.867688
R332 VREF VREF.n129 0.863781
R333 VREF VREF.n133 0.863781
R334 VREF VREF.n135 0.863781
R335 VREF VREF.n137 0.863781
R336 VREF VREF.n141 0.863781
R337 VREF VREF.n143 0.863781
R338 VREF VREF.n145 0.863781
R339 VREF VREF.n147 0.863781
R340 VREF VREF.n149 0.863781
R341 VREF VREF.n151 0.863781
R342 VREF VREF.n153 0.863781
R343 VREF VREF.n157 0.863781
R344 VREF VREF.n159 0.863781
R345 VREF VREF.n161 0.863781
R346 VREF VREF.n163 0.863781
R347 VREF VREF.n165 0.863781
R348 VREF VREF.n167 0.863781
R349 VREF VREF.n169 0.863781
R350 VREF VREF.n171 0.863781
R351 VREF VREF.n173 0.863781
R352 VREF VREF.n175 0.863781
R353 VREF VREF.n177 0.863781
R354 VREF VREF.n179 0.863781
R355 VREF VREF.n181 0.863781
R356 VREF VREF.n183 0.863781
R357 VREF VREF.n185 0.863781
R358 VREF VREF.n189 0.863781
R359 VREF VREF.n191 0.863781
R360 VREF VREF.n193 0.863781
R361 VREF VREF.n195 0.863781
R362 VREF VREF.n197 0.863781
R363 VREF VREF.n199 0.863781
R364 VREF VREF.n201 0.863781
R365 VREF VREF.n203 0.863781
R366 VREF VREF.n205 0.863781
R367 VREF VREF.n207 0.863781
R368 VREF VREF.n209 0.863781
R369 VREF VREF.n211 0.863781
R370 VREF VREF.n213 0.863781
R371 VREF VREF.n215 0.863781
R372 VREF VREF.n217 0.863781
R373 VREF VREF.n219 0.863781
R374 VREF VREF.n221 0.863781
R375 VREF VREF.n223 0.863781
R376 VREF VREF.n225 0.863781
R377 VREF VREF.n227 0.863781
R378 VREF VREF.n229 0.863781
R379 VREF VREF.n231 0.863781
R380 VREF VREF.n233 0.863781
R381 VREF VREF.n235 0.863781
R382 VREF VREF.n237 0.863781
R383 VREF VREF.n239 0.863781
R384 VREF VREF.n241 0.863781
R385 VREF VREF.n243 0.863781
R386 VREF VREF.n245 0.863781
R387 VREF VREF.n247 0.863781
R388 VREF VREF.n249 0.863781
R389 VREF VREF.n3 0.863781
R390 VREF VREF.n7 0.863781
R391 VREF VREF.n9 0.863781
R392 VREF VREF.n11 0.863781
R393 VREF VREF.n15 0.863781
R394 VREF VREF.n17 0.863781
R395 VREF VREF.n19 0.863781
R396 VREF VREF.n21 0.863781
R397 VREF VREF.n23 0.863781
R398 VREF VREF.n25 0.863781
R399 VREF VREF.n27 0.863781
R400 VREF VREF.n31 0.863781
R401 VREF VREF.n33 0.863781
R402 VREF VREF.n35 0.863781
R403 VREF VREF.n37 0.863781
R404 VREF VREF.n39 0.863781
R405 VREF VREF.n41 0.863781
R406 VREF VREF.n43 0.863781
R407 VREF VREF.n45 0.863781
R408 VREF VREF.n47 0.863781
R409 VREF VREF.n49 0.863781
R410 VREF VREF.n51 0.863781
R411 VREF VREF.n53 0.863781
R412 VREF VREF.n55 0.863781
R413 VREF VREF.n57 0.863781
R414 VREF VREF.n59 0.863781
R415 VREF VREF.n63 0.863781
R416 VREF VREF.n65 0.863781
R417 VREF VREF.n67 0.863781
R418 VREF VREF.n69 0.863781
R419 VREF VREF.n71 0.863781
R420 VREF VREF.n73 0.863781
R421 VREF VREF.n75 0.863781
R422 VREF VREF.n77 0.863781
R423 VREF VREF.n79 0.863781
R424 VREF VREF.n81 0.863781
R425 VREF VREF.n83 0.863781
R426 VREF VREF.n85 0.863781
R427 VREF VREF.n87 0.863781
R428 VREF VREF.n89 0.863781
R429 VREF VREF.n91 0.863781
R430 VREF VREF.n93 0.863781
R431 VREF VREF.n95 0.863781
R432 VREF VREF.n97 0.863781
R433 VREF VREF.n99 0.863781
R434 VREF VREF.n101 0.863781
R435 VREF VREF.n103 0.863781
R436 VREF VREF.n105 0.863781
R437 VREF VREF.n107 0.863781
R438 VREF VREF.n109 0.863781
R439 VREF VREF.n111 0.863781
R440 VREF VREF.n113 0.863781
R441 VREF VREF.n115 0.863781
R442 VREF VREF.n117 0.863781
R443 VREF VREF.n119 0.863781
R444 VREF VREF.n121 0.863781
R445 VREF VREF.n123 0.863781
R446 VREF.n5 VREF.n4 0.414822
R447 VREF.n9 VREF.n8 0.414822
R448 VREF.n11 VREF.n10 0.414822
R449 VREF.n13 VREF.n12 0.414822
R450 VREF.n17 VREF.n16 0.414822
R451 VREF.n19 VREF.n18 0.414822
R452 VREF.n21 VREF.n20 0.414822
R453 VREF.n23 VREF.n22 0.414822
R454 VREF.n25 VREF.n24 0.414822
R455 VREF.n27 VREF.n26 0.414822
R456 VREF.n29 VREF.n28 0.414822
R457 VREF.n33 VREF.n32 0.414822
R458 VREF.n35 VREF.n34 0.414822
R459 VREF.n37 VREF.n36 0.414822
R460 VREF.n39 VREF.n38 0.414822
R461 VREF.n41 VREF.n40 0.414822
R462 VREF.n43 VREF.n42 0.414822
R463 VREF.n45 VREF.n44 0.414822
R464 VREF.n47 VREF.n46 0.414822
R465 VREF.n49 VREF.n48 0.414822
R466 VREF.n51 VREF.n50 0.414822
R467 VREF.n53 VREF.n52 0.414822
R468 VREF.n55 VREF.n54 0.414822
R469 VREF.n57 VREF.n56 0.414822
R470 VREF.n59 VREF.n58 0.414822
R471 VREF.n61 VREF.n60 0.414822
R472 VREF.n65 VREF.n64 0.414822
R473 VREF.n67 VREF.n66 0.414822
R474 VREF.n69 VREF.n68 0.414822
R475 VREF.n71 VREF.n70 0.414822
R476 VREF.n73 VREF.n72 0.414822
R477 VREF.n75 VREF.n74 0.414822
R478 VREF.n77 VREF.n76 0.414822
R479 VREF.n79 VREF.n78 0.414822
R480 VREF.n81 VREF.n80 0.414822
R481 VREF.n83 VREF.n82 0.414822
R482 VREF.n85 VREF.n84 0.414822
R483 VREF.n87 VREF.n86 0.414822
R484 VREF.n89 VREF.n88 0.414822
R485 VREF.n91 VREF.n90 0.414822
R486 VREF.n93 VREF.n92 0.414822
R487 VREF.n95 VREF.n94 0.414822
R488 VREF.n97 VREF.n96 0.414822
R489 VREF.n99 VREF.n98 0.414822
R490 VREF.n101 VREF.n100 0.414822
R491 VREF.n103 VREF.n102 0.414822
R492 VREF.n105 VREF.n104 0.414822
R493 VREF.n107 VREF.n106 0.414822
R494 VREF.n109 VREF.n108 0.414822
R495 VREF.n111 VREF.n110 0.414822
R496 VREF.n113 VREF.n112 0.414822
R497 VREF.n115 VREF.n114 0.414822
R498 VREF.n117 VREF.n116 0.414822
R499 VREF.n119 VREF.n118 0.414822
R500 VREF.n121 VREF.n120 0.414822
R501 VREF.n123 VREF.n122 0.414822
R502 VREF.n125 VREF.n124 0.414822
R503 VREF VREF.n130 0.392763
R504 VREF VREF.n134 0.392763
R505 VREF VREF.n136 0.392763
R506 VREF VREF.n138 0.392763
R507 VREF VREF.n142 0.392763
R508 VREF VREF.n144 0.392763
R509 VREF VREF.n146 0.392763
R510 VREF VREF.n148 0.392763
R511 VREF VREF.n150 0.392763
R512 VREF VREF.n152 0.392763
R513 VREF VREF.n154 0.392763
R514 VREF VREF.n158 0.392763
R515 VREF VREF.n160 0.392763
R516 VREF VREF.n162 0.392763
R517 VREF VREF.n164 0.392763
R518 VREF VREF.n166 0.392763
R519 VREF VREF.n168 0.392763
R520 VREF VREF.n170 0.392763
R521 VREF VREF.n172 0.392763
R522 VREF VREF.n174 0.392763
R523 VREF VREF.n176 0.392763
R524 VREF VREF.n178 0.392763
R525 VREF VREF.n180 0.392763
R526 VREF VREF.n182 0.392763
R527 VREF VREF.n184 0.392763
R528 VREF VREF.n186 0.392763
R529 VREF VREF.n190 0.392763
R530 VREF VREF.n192 0.392763
R531 VREF VREF.n194 0.392763
R532 VREF VREF.n196 0.392763
R533 VREF VREF.n198 0.392763
R534 VREF VREF.n200 0.392763
R535 VREF VREF.n202 0.392763
R536 VREF VREF.n204 0.392763
R537 VREF VREF.n206 0.392763
R538 VREF VREF.n208 0.392763
R539 VREF VREF.n210 0.392763
R540 VREF VREF.n212 0.392763
R541 VREF VREF.n214 0.392763
R542 VREF VREF.n216 0.392763
R543 VREF VREF.n218 0.392763
R544 VREF VREF.n220 0.392763
R545 VREF VREF.n222 0.392763
R546 VREF VREF.n224 0.392763
R547 VREF VREF.n226 0.392763
R548 VREF VREF.n228 0.392763
R549 VREF VREF.n230 0.392763
R550 VREF VREF.n232 0.392763
R551 VREF VREF.n234 0.392763
R552 VREF VREF.n236 0.392763
R553 VREF VREF.n238 0.392763
R554 VREF VREF.n240 0.392763
R555 VREF VREF.n242 0.392763
R556 VREF VREF.n244 0.392763
R557 VREF VREF.n246 0.392763
R558 VREF VREF.n248 0.392763
R559 VREF VREF.n250 0.392763
R560 VREF.n128 VREF 0.102062
R561 VREF.n131 VREF 0.102062
R562 VREF.n132 VREF 0.102062
R563 VREF.n135 VREF 0.102062
R564 VREF.n137 VREF 0.102062
R565 VREF.n139 VREF 0.102062
R566 VREF.n140 VREF 0.102062
R567 VREF.n143 VREF 0.102062
R568 VREF.n145 VREF 0.102062
R569 VREF.n147 VREF 0.102062
R570 VREF.n149 VREF 0.102062
R571 VREF.n151 VREF 0.102062
R572 VREF.n153 VREF 0.102062
R573 VREF.n155 VREF 0.102062
R574 VREF.n156 VREF 0.102062
R575 VREF.n159 VREF 0.102062
R576 VREF.n161 VREF 0.102062
R577 VREF.n163 VREF 0.102062
R578 VREF.n165 VREF 0.102062
R579 VREF.n167 VREF 0.102062
R580 VREF.n169 VREF 0.102062
R581 VREF.n171 VREF 0.102062
R582 VREF.n173 VREF 0.102062
R583 VREF.n175 VREF 0.102062
R584 VREF.n177 VREF 0.102062
R585 VREF.n179 VREF 0.102062
R586 VREF.n181 VREF 0.102062
R587 VREF.n183 VREF 0.102062
R588 VREF.n185 VREF 0.102062
R589 VREF.n187 VREF 0.102062
R590 VREF.n188 VREF 0.102062
R591 VREF.n191 VREF 0.102062
R592 VREF.n193 VREF 0.102062
R593 VREF.n195 VREF 0.102062
R594 VREF.n197 VREF 0.102062
R595 VREF.n199 VREF 0.102062
R596 VREF.n201 VREF 0.102062
R597 VREF.n203 VREF 0.102062
R598 VREF.n205 VREF 0.102062
R599 VREF.n207 VREF 0.102062
R600 VREF.n209 VREF 0.102062
R601 VREF.n211 VREF 0.102062
R602 VREF.n213 VREF 0.102062
R603 VREF.n215 VREF 0.102062
R604 VREF.n217 VREF 0.102062
R605 VREF.n219 VREF 0.102062
R606 VREF.n221 VREF 0.102062
R607 VREF.n223 VREF 0.102062
R608 VREF.n225 VREF 0.102062
R609 VREF.n227 VREF 0.102062
R610 VREF.n229 VREF 0.102062
R611 VREF.n231 VREF 0.102062
R612 VREF.n233 VREF 0.102062
R613 VREF.n235 VREF 0.102062
R614 VREF.n237 VREF 0.102062
R615 VREF.n239 VREF 0.102062
R616 VREF.n241 VREF 0.102062
R617 VREF.n243 VREF 0.102062
R618 VREF.n245 VREF 0.102062
R619 VREF.n247 VREF 0.102062
R620 VREF.n249 VREF 0.102062
R621 VREF.n251 VREF 0.102062
R622 VREF.n252 VREF 0.102062
R623 VREF.n2 VREF 0.102062
R624 VREF.n5 VREF 0.102062
R625 VREF.n6 VREF 0.102062
R626 VREF.n9 VREF 0.102062
R627 VREF.n11 VREF 0.102062
R628 VREF.n13 VREF 0.102062
R629 VREF.n14 VREF 0.102062
R630 VREF.n17 VREF 0.102062
R631 VREF.n19 VREF 0.102062
R632 VREF.n21 VREF 0.102062
R633 VREF.n23 VREF 0.102062
R634 VREF.n25 VREF 0.102062
R635 VREF.n27 VREF 0.102062
R636 VREF.n29 VREF 0.102062
R637 VREF.n30 VREF 0.102062
R638 VREF.n33 VREF 0.102062
R639 VREF.n35 VREF 0.102062
R640 VREF.n37 VREF 0.102062
R641 VREF.n39 VREF 0.102062
R642 VREF.n41 VREF 0.102062
R643 VREF.n43 VREF 0.102062
R644 VREF.n45 VREF 0.102062
R645 VREF.n47 VREF 0.102062
R646 VREF.n49 VREF 0.102062
R647 VREF.n51 VREF 0.102062
R648 VREF.n53 VREF 0.102062
R649 VREF.n55 VREF 0.102062
R650 VREF.n57 VREF 0.102062
R651 VREF.n59 VREF 0.102062
R652 VREF.n61 VREF 0.102062
R653 VREF.n62 VREF 0.102062
R654 VREF.n65 VREF 0.102062
R655 VREF.n67 VREF 0.102062
R656 VREF.n69 VREF 0.102062
R657 VREF.n71 VREF 0.102062
R658 VREF.n73 VREF 0.102062
R659 VREF.n75 VREF 0.102062
R660 VREF.n77 VREF 0.102062
R661 VREF.n79 VREF 0.102062
R662 VREF.n81 VREF 0.102062
R663 VREF.n83 VREF 0.102062
R664 VREF.n85 VREF 0.102062
R665 VREF.n87 VREF 0.102062
R666 VREF.n89 VREF 0.102062
R667 VREF.n91 VREF 0.102062
R668 VREF.n93 VREF 0.102062
R669 VREF.n95 VREF 0.102062
R670 VREF.n97 VREF 0.102062
R671 VREF.n99 VREF 0.102062
R672 VREF.n101 VREF 0.102062
R673 VREF.n103 VREF 0.102062
R674 VREF.n105 VREF 0.102062
R675 VREF.n107 VREF 0.102062
R676 VREF.n109 VREF 0.102062
R677 VREF.n111 VREF 0.102062
R678 VREF.n113 VREF 0.102062
R679 VREF.n115 VREF 0.102062
R680 VREF.n117 VREF 0.102062
R681 VREF.n119 VREF 0.102062
R682 VREF.n121 VREF 0.102062
R683 VREF.n123 VREF 0.102062
R684 VREF.n125 VREF 0.102062
R685 VREF VREF.n254 0.102062
R686 VREF.n0 VREF 0.0335882
R687 VREF.n1 VREF 0.0335882
R688 VREF.n2 VREF 0.0335882
R689 VREF.n3 VREF 0.0335882
R690 VREF.n5 VREF 0.0335882
R691 VREF.n6 VREF 0.0335882
R692 VREF.n7 VREF 0.0335882
R693 VREF.n9 VREF 0.0335882
R694 VREF.n11 VREF 0.0335882
R695 VREF.n13 VREF 0.0335882
R696 VREF.n14 VREF 0.0335882
R697 VREF.n15 VREF 0.0335882
R698 VREF.n17 VREF 0.0335882
R699 VREF.n19 VREF 0.0335882
R700 VREF.n21 VREF 0.0335882
R701 VREF.n23 VREF 0.0335882
R702 VREF.n25 VREF 0.0335882
R703 VREF.n27 VREF 0.0335882
R704 VREF.n29 VREF 0.0335882
R705 VREF.n30 VREF 0.0335882
R706 VREF.n31 VREF 0.0335882
R707 VREF.n33 VREF 0.0335882
R708 VREF.n35 VREF 0.0335882
R709 VREF.n37 VREF 0.0335882
R710 VREF.n39 VREF 0.0335882
R711 VREF.n41 VREF 0.0335882
R712 VREF.n43 VREF 0.0335882
R713 VREF.n45 VREF 0.0335882
R714 VREF.n47 VREF 0.0335882
R715 VREF.n49 VREF 0.0335882
R716 VREF.n51 VREF 0.0335882
R717 VREF.n53 VREF 0.0335882
R718 VREF.n55 VREF 0.0335882
R719 VREF.n57 VREF 0.0335882
R720 VREF.n59 VREF 0.0335882
R721 VREF.n61 VREF 0.0335882
R722 VREF.n62 VREF 0.0335882
R723 VREF.n63 VREF 0.0335882
R724 VREF.n65 VREF 0.0335882
R725 VREF.n67 VREF 0.0335882
R726 VREF.n69 VREF 0.0335882
R727 VREF.n71 VREF 0.0335882
R728 VREF.n73 VREF 0.0335882
R729 VREF.n75 VREF 0.0335882
R730 VREF.n77 VREF 0.0335882
R731 VREF.n79 VREF 0.0335882
R732 VREF.n81 VREF 0.0335882
R733 VREF.n83 VREF 0.0335882
R734 VREF.n85 VREF 0.0335882
R735 VREF.n87 VREF 0.0335882
R736 VREF.n89 VREF 0.0335882
R737 VREF.n91 VREF 0.0335882
R738 VREF.n93 VREF 0.0335882
R739 VREF.n95 VREF 0.0335882
R740 VREF.n97 VREF 0.0335882
R741 VREF.n99 VREF 0.0335882
R742 VREF.n101 VREF 0.0335882
R743 VREF.n103 VREF 0.0335882
R744 VREF.n105 VREF 0.0335882
R745 VREF.n107 VREF 0.0335882
R746 VREF.n109 VREF 0.0335882
R747 VREF.n111 VREF 0.0335882
R748 VREF.n113 VREF 0.0335882
R749 VREF.n115 VREF 0.0335882
R750 VREF.n117 VREF 0.0335882
R751 VREF.n119 VREF 0.0335882
R752 VREF.n121 VREF 0.0335882
R753 VREF.n123 VREF 0.0335882
R754 VREF.n125 VREF 0.0335882
R755 VREF.n254 VREF 0.0335882
R756 VREF.n0 VREF 0.0249565
R757 VREF.n126 VREF 0.0225588
R758 VREF.n127 VREF 0.0225588
R759 VREF.n128 VREF 0.0225588
R760 VREF.n129 VREF 0.0225588
R761 VREF.n131 VREF 0.0225588
R762 VREF.n132 VREF 0.0225588
R763 VREF.n133 VREF 0.0225588
R764 VREF.n135 VREF 0.0225588
R765 VREF.n137 VREF 0.0225588
R766 VREF.n139 VREF 0.0225588
R767 VREF.n140 VREF 0.0225588
R768 VREF.n141 VREF 0.0225588
R769 VREF.n143 VREF 0.0225588
R770 VREF.n145 VREF 0.0225588
R771 VREF.n147 VREF 0.0225588
R772 VREF.n149 VREF 0.0225588
R773 VREF.n151 VREF 0.0225588
R774 VREF.n153 VREF 0.0225588
R775 VREF.n155 VREF 0.0225588
R776 VREF.n156 VREF 0.0225588
R777 VREF.n157 VREF 0.0225588
R778 VREF.n159 VREF 0.0225588
R779 VREF.n161 VREF 0.0225588
R780 VREF.n163 VREF 0.0225588
R781 VREF.n165 VREF 0.0225588
R782 VREF.n167 VREF 0.0225588
R783 VREF.n169 VREF 0.0225588
R784 VREF.n171 VREF 0.0225588
R785 VREF.n173 VREF 0.0225588
R786 VREF.n175 VREF 0.0225588
R787 VREF.n177 VREF 0.0225588
R788 VREF.n179 VREF 0.0225588
R789 VREF.n181 VREF 0.0225588
R790 VREF.n183 VREF 0.0225588
R791 VREF.n185 VREF 0.0225588
R792 VREF.n187 VREF 0.0225588
R793 VREF.n188 VREF 0.0225588
R794 VREF.n189 VREF 0.0225588
R795 VREF.n191 VREF 0.0225588
R796 VREF.n193 VREF 0.0225588
R797 VREF.n195 VREF 0.0225588
R798 VREF.n197 VREF 0.0225588
R799 VREF.n199 VREF 0.0225588
R800 VREF.n201 VREF 0.0225588
R801 VREF.n203 VREF 0.0225588
R802 VREF.n205 VREF 0.0225588
R803 VREF.n207 VREF 0.0225588
R804 VREF.n209 VREF 0.0225588
R805 VREF.n211 VREF 0.0225588
R806 VREF.n213 VREF 0.0225588
R807 VREF.n215 VREF 0.0225588
R808 VREF.n217 VREF 0.0225588
R809 VREF.n219 VREF 0.0225588
R810 VREF.n221 VREF 0.0225588
R811 VREF.n223 VREF 0.0225588
R812 VREF.n225 VREF 0.0225588
R813 VREF.n227 VREF 0.0225588
R814 VREF.n229 VREF 0.0225588
R815 VREF.n231 VREF 0.0225588
R816 VREF.n233 VREF 0.0225588
R817 VREF.n235 VREF 0.0225588
R818 VREF.n237 VREF 0.0225588
R819 VREF.n239 VREF 0.0225588
R820 VREF.n241 VREF 0.0225588
R821 VREF.n243 VREF 0.0225588
R822 VREF.n245 VREF 0.0225588
R823 VREF.n247 VREF 0.0225588
R824 VREF.n249 VREF 0.0225588
R825 VREF.n251 VREF 0.0225588
R826 VREF.n252 VREF 0.0225588
R827 VREF.n126 VREF 0.0168043
R828 VREF.n127 VREF 0.00440625
R829 VREF.n129 VREF 0.00440625
R830 VREF.n131 VREF 0.00440625
R831 VREF.n133 VREF 0.00440625
R832 VREF.n135 VREF 0.00440625
R833 VREF.n137 VREF 0.00440625
R834 VREF.n139 VREF 0.00440625
R835 VREF.n141 VREF 0.00440625
R836 VREF.n143 VREF 0.00440625
R837 VREF.n145 VREF 0.00440625
R838 VREF.n147 VREF 0.00440625
R839 VREF.n149 VREF 0.00440625
R840 VREF.n151 VREF 0.00440625
R841 VREF.n153 VREF 0.00440625
R842 VREF.n155 VREF 0.00440625
R843 VREF.n157 VREF 0.00440625
R844 VREF.n159 VREF 0.00440625
R845 VREF.n161 VREF 0.00440625
R846 VREF.n163 VREF 0.00440625
R847 VREF.n165 VREF 0.00440625
R848 VREF.n167 VREF 0.00440625
R849 VREF.n169 VREF 0.00440625
R850 VREF.n171 VREF 0.00440625
R851 VREF.n173 VREF 0.00440625
R852 VREF.n175 VREF 0.00440625
R853 VREF.n177 VREF 0.00440625
R854 VREF.n179 VREF 0.00440625
R855 VREF.n181 VREF 0.00440625
R856 VREF.n183 VREF 0.00440625
R857 VREF.n185 VREF 0.00440625
R858 VREF.n187 VREF 0.00440625
R859 VREF.n189 VREF 0.00440625
R860 VREF.n191 VREF 0.00440625
R861 VREF.n193 VREF 0.00440625
R862 VREF.n195 VREF 0.00440625
R863 VREF.n197 VREF 0.00440625
R864 VREF.n199 VREF 0.00440625
R865 VREF.n201 VREF 0.00440625
R866 VREF.n203 VREF 0.00440625
R867 VREF.n205 VREF 0.00440625
R868 VREF.n207 VREF 0.00440625
R869 VREF.n209 VREF 0.00440625
R870 VREF.n211 VREF 0.00440625
R871 VREF.n213 VREF 0.00440625
R872 VREF.n215 VREF 0.00440625
R873 VREF.n217 VREF 0.00440625
R874 VREF.n219 VREF 0.00440625
R875 VREF.n221 VREF 0.00440625
R876 VREF.n223 VREF 0.00440625
R877 VREF.n225 VREF 0.00440625
R878 VREF.n227 VREF 0.00440625
R879 VREF.n229 VREF 0.00440625
R880 VREF.n231 VREF 0.00440625
R881 VREF.n233 VREF 0.00440625
R882 VREF.n235 VREF 0.00440625
R883 VREF.n237 VREF 0.00440625
R884 VREF.n239 VREF 0.00440625
R885 VREF.n241 VREF 0.00440625
R886 VREF.n243 VREF 0.00440625
R887 VREF.n245 VREF 0.00440625
R888 VREF.n247 VREF 0.00440625
R889 VREF.n249 VREF 0.00440625
R890 VREF.n251 VREF 0.00440625
R891 VREF.n1 VREF 0.00440625
R892 VREF.n3 VREF 0.00440625
R893 VREF.n5 VREF 0.00440625
R894 VREF.n7 VREF 0.00440625
R895 VREF.n9 VREF 0.00440625
R896 VREF.n11 VREF 0.00440625
R897 VREF.n13 VREF 0.00440625
R898 VREF.n15 VREF 0.00440625
R899 VREF.n17 VREF 0.00440625
R900 VREF.n19 VREF 0.00440625
R901 VREF.n21 VREF 0.00440625
R902 VREF.n23 VREF 0.00440625
R903 VREF.n25 VREF 0.00440625
R904 VREF.n27 VREF 0.00440625
R905 VREF.n29 VREF 0.00440625
R906 VREF.n31 VREF 0.00440625
R907 VREF.n33 VREF 0.00440625
R908 VREF.n35 VREF 0.00440625
R909 VREF.n37 VREF 0.00440625
R910 VREF.n39 VREF 0.00440625
R911 VREF.n41 VREF 0.00440625
R912 VREF.n43 VREF 0.00440625
R913 VREF.n45 VREF 0.00440625
R914 VREF.n47 VREF 0.00440625
R915 VREF.n49 VREF 0.00440625
R916 VREF.n51 VREF 0.00440625
R917 VREF.n53 VREF 0.00440625
R918 VREF.n55 VREF 0.00440625
R919 VREF.n57 VREF 0.00440625
R920 VREF.n59 VREF 0.00440625
R921 VREF.n61 VREF 0.00440625
R922 VREF.n63 VREF 0.00440625
R923 VREF.n65 VREF 0.00440625
R924 VREF.n67 VREF 0.00440625
R925 VREF.n69 VREF 0.00440625
R926 VREF.n71 VREF 0.00440625
R927 VREF.n73 VREF 0.00440625
R928 VREF.n75 VREF 0.00440625
R929 VREF.n77 VREF 0.00440625
R930 VREF.n79 VREF 0.00440625
R931 VREF.n81 VREF 0.00440625
R932 VREF.n83 VREF 0.00440625
R933 VREF.n85 VREF 0.00440625
R934 VREF.n87 VREF 0.00440625
R935 VREF.n89 VREF 0.00440625
R936 VREF.n91 VREF 0.00440625
R937 VREF.n93 VREF 0.00440625
R938 VREF.n95 VREF 0.00440625
R939 VREF.n97 VREF 0.00440625
R940 VREF.n99 VREF 0.00440625
R941 VREF.n101 VREF 0.00440625
R942 VREF.n103 VREF 0.00440625
R943 VREF.n105 VREF 0.00440625
R944 VREF.n107 VREF 0.00440625
R945 VREF.n109 VREF 0.00440625
R946 VREF.n111 VREF 0.00440625
R947 VREF.n113 VREF 0.00440625
R948 VREF.n115 VREF 0.00440625
R949 VREF.n117 VREF 0.00440625
R950 VREF.n119 VREF 0.00440625
R951 VREF.n121 VREF 0.00440625
R952 VREF.n123 VREF 0.00440625
R953 VREF.n125 VREF 0.00440625
R954 VDD.n407 VDD.t244 587.957
R955 VDD.n407 VDD.t108 587.957
R956 VDD.n394 VDD.t222 332.5
R957 VDD.n390 VDD.t87 332.5
R958 VDD.n634 VDD.n633 324.175
R959 VDD.n475 VDD.n473 266.296
R960 VDD.n865 VDD.n864 215.93
R961 VDD.n413 VDD.n409 186.992
R962 VDD.n443 VDD.n442 165.565
R963 VDD.n369 VDD.t35 158.335
R964 VDD.n317 VDD.t209 158.335
R965 VDD.n215 VDD.t168 158.335
R966 VDD.n863 VDD.t103 158.335
R967 VDD.n632 VDD.t176 158.335
R968 VDD.n513 VDD.t70 158.335
R969 VDD.n441 VDD.t192 158.335
R970 VDD.n382 VDD.t229 158.333
R971 VDD.n385 VDD.t230 158.333
R972 VDD.n446 VDD.t227 158.333
R973 VDD.n468 VDD.t158 158.333
R974 VDD.n370 VDD.t221 158.333
R975 VDD.n548 VDD.t41 158.333
R976 VDD.n318 VDD.t248 158.333
R977 VDD.n320 VDD.t112 158.333
R978 VDD.n323 VDD.t117 158.333
R979 VDD.n540 VDD.t159 158.333
R980 VDD.n325 VDD.t1 158.333
R981 VDD.n534 VDD.t232 158.333
R982 VDD.n328 VDD.t131 158.333
R983 VDD.n330 VDD.t243 158.333
R984 VDD.n333 VDD.t113 158.333
R985 VDD.n526 VDD.t67 158.333
R986 VDD.n335 VDD.t178 158.333
R987 VDD.n520 VDD.t160 158.333
R988 VDD.n338 VDD.t81 158.333
R989 VDD.n340 VDD.t218 158.333
R990 VDD.n706 VDD.t193 158.333
R991 VDD.n216 VDD.t118 158.333
R992 VDD.n218 VDD.t95 158.333
R993 VDD.n221 VDD.t98 158.333
R994 VDD.n698 VDD.t104 158.333
R995 VDD.n223 VDD.t4 158.333
R996 VDD.n692 VDD.t163 158.333
R997 VDD.n226 VDD.t200 158.333
R998 VDD.n228 VDD.t223 158.333
R999 VDD.n231 VDD.t92 158.333
R1000 VDD.n684 VDD.t174 158.333
R1001 VDD.n233 VDD.t151 158.333
R1002 VDD.n678 VDD.t199 158.333
R1003 VDD.n236 VDD.t14 158.333
R1004 VDD.n238 VDD.t133 158.333
R1005 VDD.n241 VDD.t198 158.333
R1006 VDD.n670 VDD.t65 158.333
R1007 VDD.n243 VDD.t161 158.333
R1008 VDD.n664 VDD.t51 158.333
R1009 VDD.n246 VDD.t171 158.333
R1010 VDD.n248 VDD.t142 158.333
R1011 VDD.n251 VDD.t91 158.333
R1012 VDD.n656 VDD.t241 158.333
R1013 VDD.n253 VDD.t97 158.333
R1014 VDD.n650 VDD.t107 158.333
R1015 VDD.n256 VDD.t94 158.333
R1016 VDD.n258 VDD.t173 158.333
R1017 VDD.n261 VDD.t138 158.333
R1018 VDD.n642 VDD.t56 158.333
R1019 VDD.n263 VDD.t46 158.333
R1020 VDD.n636 VDD.t162 158.333
R1021 VDD.n3 VDD.t106 158.333
R1022 VDD.n7 VDD.t110 158.333
R1023 VDD.n7 VDD.t195 158.333
R1024 VDD.n1008 VDD.t236 158.333
R1025 VDD.n9 VDD.t58 158.333
R1026 VDD.n1002 VDD.t157 158.333
R1027 VDD.n12 VDD.t175 158.333
R1028 VDD.n14 VDD.t83 158.333
R1029 VDD.n17 VDD.t214 158.333
R1030 VDD.n994 VDD.t25 158.333
R1031 VDD.n19 VDD.t119 158.333
R1032 VDD.n988 VDD.t238 158.333
R1033 VDD.n22 VDD.t76 158.333
R1034 VDD.n24 VDD.t210 158.333
R1035 VDD.n27 VDD.t86 158.333
R1036 VDD.n980 VDD.t27 158.333
R1037 VDD.n29 VDD.t34 158.333
R1038 VDD.n974 VDD.t148 158.333
R1039 VDD.n32 VDD.t156 158.333
R1040 VDD.n34 VDD.t124 158.333
R1041 VDD.n37 VDD.t141 158.333
R1042 VDD.n966 VDD.t130 158.333
R1043 VDD.n39 VDD.t109 158.333
R1044 VDD.n960 VDD.t126 158.333
R1045 VDD.n42 VDD.t189 158.333
R1046 VDD.n44 VDD.t242 158.333
R1047 VDD.n47 VDD.t235 158.333
R1048 VDD.n952 VDD.t179 158.333
R1049 VDD.n49 VDD.t215 158.333
R1050 VDD.n946 VDD.t60 158.333
R1051 VDD.n52 VDD.t82 158.333
R1052 VDD.n54 VDD.t213 158.333
R1053 VDD.n57 VDD.t237 158.333
R1054 VDD.n938 VDD.t123 158.333
R1055 VDD.n59 VDD.t234 158.333
R1056 VDD.n932 VDD.t18 158.333
R1057 VDD.n62 VDD.t207 158.333
R1058 VDD.n64 VDD.t62 158.333
R1059 VDD.n67 VDD.t15 158.333
R1060 VDD.n924 VDD.t8 158.333
R1061 VDD.n69 VDD.t233 158.333
R1062 VDD.n918 VDD.t202 158.333
R1063 VDD.n72 VDD.t114 158.333
R1064 VDD.n74 VDD.t197 158.333
R1065 VDD.n77 VDD.t85 158.333
R1066 VDD.n910 VDD.t84 158.333
R1067 VDD.n79 VDD.t246 158.333
R1068 VDD.n904 VDD.t40 158.333
R1069 VDD.n82 VDD.t194 158.333
R1070 VDD.n84 VDD.t212 158.333
R1071 VDD.n87 VDD.t196 158.333
R1072 VDD.n896 VDD.t16 158.333
R1073 VDD.n89 VDD.t59 158.333
R1074 VDD.n890 VDD.t125 158.333
R1075 VDD.n92 VDD.t66 158.333
R1076 VDD.n94 VDD.t72 158.333
R1077 VDD.n97 VDD.t73 158.333
R1078 VDD.n882 VDD.t208 158.333
R1079 VDD.n99 VDD.t22 158.333
R1080 VDD.n876 VDD.t211 158.333
R1081 VDD.n102 VDD.t203 158.333
R1082 VDD.n104 VDD.t31 158.333
R1083 VDD.n107 VDD.t38 158.333
R1084 VDD.n868 VDD.t7 158.333
R1085 VDD.n110 VDD.t93 158.333
R1086 VDD.n857 VDD.t150 158.333
R1087 VDD.n112 VDD.t71 158.333
R1088 VDD.n851 VDD.t204 158.333
R1089 VDD.n115 VDD.t226 158.333
R1090 VDD.n117 VDD.t75 158.333
R1091 VDD.n120 VDD.t224 158.333
R1092 VDD.n843 VDD.t135 158.333
R1093 VDD.n122 VDD.t167 158.333
R1094 VDD.n837 VDD.t77 158.333
R1095 VDD.n125 VDD.t32 158.333
R1096 VDD.n127 VDD.t79 158.333
R1097 VDD.n130 VDD.t13 158.333
R1098 VDD.n829 VDD.t188 158.333
R1099 VDD.n132 VDD.t165 158.333
R1100 VDD.n823 VDD.t139 158.333
R1101 VDD.n135 VDD.t128 158.333
R1102 VDD.n137 VDD.t177 158.333
R1103 VDD.n140 VDD.t121 158.333
R1104 VDD.n815 VDD.t33 158.333
R1105 VDD.n142 VDD.t45 158.333
R1106 VDD.n809 VDD.t48 158.333
R1107 VDD.n145 VDD.t225 158.333
R1108 VDD.n147 VDD.t64 158.333
R1109 VDD.n150 VDD.t3 158.333
R1110 VDD.n801 VDD.t220 158.333
R1111 VDD.n152 VDD.t99 158.333
R1112 VDD.n795 VDD.t122 158.333
R1113 VDD.n155 VDD.t134 158.333
R1114 VDD.n157 VDD.t191 158.333
R1115 VDD.n160 VDD.t23 158.333
R1116 VDD.n787 VDD.t44 158.333
R1117 VDD.n162 VDD.t89 158.333
R1118 VDD.n781 VDD.t190 158.333
R1119 VDD.n165 VDD.t140 158.333
R1120 VDD.n167 VDD.t132 158.333
R1121 VDD.n170 VDD.t100 158.333
R1122 VDD.n773 VDD.t187 158.333
R1123 VDD.n172 VDD.t102 158.333
R1124 VDD.n767 VDD.t111 158.333
R1125 VDD.n175 VDD.t20 158.333
R1126 VDD.n177 VDD.t152 158.333
R1127 VDD.n180 VDD.t231 158.333
R1128 VDD.n759 VDD.t129 158.333
R1129 VDD.n182 VDD.t9 158.333
R1130 VDD.n753 VDD.t39 158.333
R1131 VDD.n185 VDD.t69 158.333
R1132 VDD.n187 VDD.t96 158.333
R1133 VDD.n190 VDD.t143 158.333
R1134 VDD.n745 VDD.t12 158.333
R1135 VDD.n192 VDD.t169 158.333
R1136 VDD.n739 VDD.t47 158.333
R1137 VDD.n195 VDD.t154 158.333
R1138 VDD.n197 VDD.t137 158.333
R1139 VDD.n200 VDD.t0 158.333
R1140 VDD.n731 VDD.t43 158.333
R1141 VDD.n202 VDD.t11 158.333
R1142 VDD.n725 VDD.t186 158.333
R1143 VDD.n205 VDD.t24 158.333
R1144 VDD.n207 VDD.t50 158.333
R1145 VDD.n210 VDD.t5 158.333
R1146 VDD.n717 VDD.t52 158.333
R1147 VDD.n212 VDD.t216 158.333
R1148 VDD.n267 VDD.t166 158.333
R1149 VDD.n626 VDD.t90 158.333
R1150 VDD.n269 VDD.t170 158.333
R1151 VDD.n620 VDD.t247 158.333
R1152 VDD.n272 VDD.t21 158.333
R1153 VDD.n274 VDD.t146 158.333
R1154 VDD.n277 VDD.t116 158.333
R1155 VDD.n612 VDD.t68 158.333
R1156 VDD.n279 VDD.t101 158.333
R1157 VDD.n606 VDD.t78 158.333
R1158 VDD.n282 VDD.t149 158.333
R1159 VDD.n284 VDD.t63 158.333
R1160 VDD.n287 VDD.t127 158.333
R1161 VDD.n598 VDD.t53 158.333
R1162 VDD.n289 VDD.t74 158.333
R1163 VDD.n592 VDD.t164 158.333
R1164 VDD.n292 VDD.t61 158.333
R1165 VDD.n294 VDD.t55 158.333
R1166 VDD.n297 VDD.t219 158.333
R1167 VDD.n584 VDD.t136 158.333
R1168 VDD.n299 VDD.t239 158.333
R1169 VDD.n578 VDD.t182 158.333
R1170 VDD.n302 VDD.t28 158.333
R1171 VDD.n304 VDD.t205 158.333
R1172 VDD.n307 VDD.t42 158.333
R1173 VDD.n570 VDD.t37 158.333
R1174 VDD.n309 VDD.t6 158.333
R1175 VDD.n564 VDD.t17 158.333
R1176 VDD.n312 VDD.t54 158.333
R1177 VDD.n314 VDD.t19 158.333
R1178 VDD.n557 VDD.t36 158.333
R1179 VDD.n344 VDD.t2 158.333
R1180 VDD.n507 VDD.t144 158.333
R1181 VDD.n346 VDD.t29 158.333
R1182 VDD.n501 VDD.t26 158.333
R1183 VDD.n349 VDD.t105 158.333
R1184 VDD.n351 VDD.t115 158.333
R1185 VDD.n354 VDD.t57 158.333
R1186 VDD.n493 VDD.t206 158.333
R1187 VDD.n356 VDD.t49 158.333
R1188 VDD.n487 VDD.t10 158.333
R1189 VDD.n359 VDD.t180 158.333
R1190 VDD.n361 VDD.t120 158.333
R1191 VDD.n364 VDD.t183 158.333
R1192 VDD.n479 VDD.t201 158.333
R1193 VDD.n366 VDD.t217 158.333
R1194 VDD.n388 VDD.t181 158.333
R1195 VDD.n435 VDD.t245 158.333
R1196 VDD.n395 VDD.t185 158.333
R1197 VDD.n397 VDD.t145 158.333
R1198 VDD.n422 VDD.t30 158.333
R1199 VDD.n515 VDD.n514 149.149
R1200 VDD.n420 VDD.n418 138.018
R1201 VDD.n713 VDD.n711 133.565
R1202 VDD.n555 VDD.n553 126.609
R1203 VDD.n372 VDD.t153 121.886
R1204 VDD.n375 VDD.t172 93.539
R1205 VDD.n460 VDD.t80 93.539
R1206 VDD.n377 VDD.t147 93.539
R1207 VDD.n454 VDD.t88 93.539
R1208 VDD.n380 VDD.t228 93.539
R1209 VDD.n401 VDD.t240 93.539
R1210 VDD.n401 VDD.t155 93.539
R1211 VDD.n404 VDD.t184 93.539
R1212 VDD.n391 VDD.n390 69.2713
R1213 VDD.n395 VDD.n394 69.2713
R1214 VDD.n1011 VDD.n1010 35.6179
R1215 VDD.n1010 VDD.n11 35.6179
R1216 VDD.n1004 VDD.n11 35.6179
R1217 VDD.n1004 VDD.n1001 35.6179
R1218 VDD.n1001 VDD.n16 35.6179
R1219 VDD.n997 VDD.n16 35.6179
R1220 VDD.n997 VDD.n996 35.6179
R1221 VDD.n996 VDD.n21 35.6179
R1222 VDD.n990 VDD.n21 35.6179
R1223 VDD.n990 VDD.n987 35.6179
R1224 VDD.n987 VDD.n26 35.6179
R1225 VDD.n983 VDD.n26 35.6179
R1226 VDD.n983 VDD.n982 35.6179
R1227 VDD.n982 VDD.n31 35.6179
R1228 VDD.n976 VDD.n31 35.6179
R1229 VDD.n976 VDD.n973 35.6179
R1230 VDD.n973 VDD.n36 35.6179
R1231 VDD.n969 VDD.n36 35.6179
R1232 VDD.n969 VDD.n968 35.6179
R1233 VDD.n968 VDD.n41 35.6179
R1234 VDD.n962 VDD.n41 35.6179
R1235 VDD.n962 VDD.n959 35.6179
R1236 VDD.n959 VDD.n46 35.6179
R1237 VDD.n955 VDD.n46 35.6179
R1238 VDD.n955 VDD.n954 35.6179
R1239 VDD.n954 VDD.n51 35.6179
R1240 VDD.n948 VDD.n51 35.6179
R1241 VDD.n948 VDD.n945 35.6179
R1242 VDD.n945 VDD.n56 35.6179
R1243 VDD.n941 VDD.n56 35.6179
R1244 VDD.n941 VDD.n940 35.6179
R1245 VDD.n940 VDD.n61 35.6179
R1246 VDD.n934 VDD.n61 35.6179
R1247 VDD.n934 VDD.n931 35.6179
R1248 VDD.n931 VDD.n66 35.6179
R1249 VDD.n927 VDD.n66 35.6179
R1250 VDD.n927 VDD.n926 35.6179
R1251 VDD.n926 VDD.n71 35.6179
R1252 VDD.n920 VDD.n71 35.6179
R1253 VDD.n920 VDD.n917 35.6179
R1254 VDD.n917 VDD.n76 35.6179
R1255 VDD.n913 VDD.n76 35.6179
R1256 VDD.n913 VDD.n912 35.6179
R1257 VDD.n912 VDD.n81 35.6179
R1258 VDD.n906 VDD.n81 35.6179
R1259 VDD.n906 VDD.n903 35.6179
R1260 VDD.n903 VDD.n86 35.6179
R1261 VDD.n899 VDD.n86 35.6179
R1262 VDD.n899 VDD.n898 35.6179
R1263 VDD.n898 VDD.n91 35.6179
R1264 VDD.n892 VDD.n91 35.6179
R1265 VDD.n892 VDD.n889 35.6179
R1266 VDD.n889 VDD.n96 35.6179
R1267 VDD.n885 VDD.n96 35.6179
R1268 VDD.n885 VDD.n884 35.6179
R1269 VDD.n884 VDD.n101 35.6179
R1270 VDD.n878 VDD.n101 35.6179
R1271 VDD.n878 VDD.n875 35.6179
R1272 VDD.n875 VDD.n106 35.6179
R1273 VDD.n871 VDD.n106 35.6179
R1274 VDD.n871 VDD.n870 35.6179
R1275 VDD.n860 VDD.n859 35.6179
R1276 VDD.n859 VDD.n114 35.6179
R1277 VDD.n853 VDD.n114 35.6179
R1278 VDD.n853 VDD.n850 35.6179
R1279 VDD.n850 VDD.n119 35.6179
R1280 VDD.n846 VDD.n119 35.6179
R1281 VDD.n846 VDD.n845 35.6179
R1282 VDD.n845 VDD.n124 35.6179
R1283 VDD.n839 VDD.n124 35.6179
R1284 VDD.n839 VDD.n836 35.6179
R1285 VDD.n836 VDD.n129 35.6179
R1286 VDD.n832 VDD.n129 35.6179
R1287 VDD.n832 VDD.n831 35.6179
R1288 VDD.n831 VDD.n134 35.6179
R1289 VDD.n825 VDD.n134 35.6179
R1290 VDD.n825 VDD.n822 35.6179
R1291 VDD.n822 VDD.n139 35.6179
R1292 VDD.n818 VDD.n139 35.6179
R1293 VDD.n818 VDD.n817 35.6179
R1294 VDD.n817 VDD.n144 35.6179
R1295 VDD.n811 VDD.n144 35.6179
R1296 VDD.n811 VDD.n808 35.6179
R1297 VDD.n808 VDD.n149 35.6179
R1298 VDD.n804 VDD.n149 35.6179
R1299 VDD.n804 VDD.n803 35.6179
R1300 VDD.n803 VDD.n154 35.6179
R1301 VDD.n797 VDD.n154 35.6179
R1302 VDD.n797 VDD.n794 35.6179
R1303 VDD.n794 VDD.n159 35.6179
R1304 VDD.n790 VDD.n159 35.6179
R1305 VDD.n790 VDD.n789 35.6179
R1306 VDD.n789 VDD.n164 35.6179
R1307 VDD.n783 VDD.n164 35.6179
R1308 VDD.n783 VDD.n780 35.6179
R1309 VDD.n780 VDD.n169 35.6179
R1310 VDD.n776 VDD.n169 35.6179
R1311 VDD.n776 VDD.n775 35.6179
R1312 VDD.n775 VDD.n174 35.6179
R1313 VDD.n769 VDD.n174 35.6179
R1314 VDD.n769 VDD.n766 35.6179
R1315 VDD.n766 VDD.n179 35.6179
R1316 VDD.n762 VDD.n179 35.6179
R1317 VDD.n762 VDD.n761 35.6179
R1318 VDD.n761 VDD.n184 35.6179
R1319 VDD.n755 VDD.n184 35.6179
R1320 VDD.n755 VDD.n752 35.6179
R1321 VDD.n752 VDD.n189 35.6179
R1322 VDD.n748 VDD.n189 35.6179
R1323 VDD.n748 VDD.n747 35.6179
R1324 VDD.n747 VDD.n194 35.6179
R1325 VDD.n741 VDD.n194 35.6179
R1326 VDD.n741 VDD.n738 35.6179
R1327 VDD.n738 VDD.n199 35.6179
R1328 VDD.n734 VDD.n199 35.6179
R1329 VDD.n734 VDD.n733 35.6179
R1330 VDD.n733 VDD.n204 35.6179
R1331 VDD.n727 VDD.n204 35.6179
R1332 VDD.n727 VDD.n724 35.6179
R1333 VDD.n724 VDD.n209 35.6179
R1334 VDD.n720 VDD.n209 35.6179
R1335 VDD.n720 VDD.n719 35.6179
R1336 VDD.n719 VDD.n214 35.6179
R1337 VDD.n708 VDD.n705 35.6179
R1338 VDD.n705 VDD.n220 35.6179
R1339 VDD.n701 VDD.n220 35.6179
R1340 VDD.n701 VDD.n700 35.6179
R1341 VDD.n700 VDD.n225 35.6179
R1342 VDD.n694 VDD.n225 35.6179
R1343 VDD.n694 VDD.n691 35.6179
R1344 VDD.n691 VDD.n230 35.6179
R1345 VDD.n687 VDD.n230 35.6179
R1346 VDD.n687 VDD.n686 35.6179
R1347 VDD.n686 VDD.n235 35.6179
R1348 VDD.n680 VDD.n235 35.6179
R1349 VDD.n680 VDD.n677 35.6179
R1350 VDD.n677 VDD.n240 35.6179
R1351 VDD.n673 VDD.n240 35.6179
R1352 VDD.n673 VDD.n672 35.6179
R1353 VDD.n672 VDD.n245 35.6179
R1354 VDD.n666 VDD.n245 35.6179
R1355 VDD.n666 VDD.n663 35.6179
R1356 VDD.n663 VDD.n250 35.6179
R1357 VDD.n659 VDD.n250 35.6179
R1358 VDD.n659 VDD.n658 35.6179
R1359 VDD.n658 VDD.n255 35.6179
R1360 VDD.n652 VDD.n255 35.6179
R1361 VDD.n652 VDD.n649 35.6179
R1362 VDD.n649 VDD.n260 35.6179
R1363 VDD.n645 VDD.n260 35.6179
R1364 VDD.n645 VDD.n644 35.6179
R1365 VDD.n644 VDD.n265 35.6179
R1366 VDD.n638 VDD.n265 35.6179
R1367 VDD.n629 VDD.n628 35.6179
R1368 VDD.n628 VDD.n271 35.6179
R1369 VDD.n622 VDD.n271 35.6179
R1370 VDD.n622 VDD.n619 35.6179
R1371 VDD.n619 VDD.n276 35.6179
R1372 VDD.n615 VDD.n276 35.6179
R1373 VDD.n615 VDD.n614 35.6179
R1374 VDD.n614 VDD.n281 35.6179
R1375 VDD.n608 VDD.n281 35.6179
R1376 VDD.n608 VDD.n605 35.6179
R1377 VDD.n605 VDD.n286 35.6179
R1378 VDD.n601 VDD.n286 35.6179
R1379 VDD.n601 VDD.n600 35.6179
R1380 VDD.n600 VDD.n291 35.6179
R1381 VDD.n594 VDD.n291 35.6179
R1382 VDD.n594 VDD.n591 35.6179
R1383 VDD.n591 VDD.n296 35.6179
R1384 VDD.n587 VDD.n296 35.6179
R1385 VDD.n587 VDD.n586 35.6179
R1386 VDD.n586 VDD.n301 35.6179
R1387 VDD.n580 VDD.n301 35.6179
R1388 VDD.n580 VDD.n577 35.6179
R1389 VDD.n577 VDD.n306 35.6179
R1390 VDD.n573 VDD.n306 35.6179
R1391 VDD.n573 VDD.n572 35.6179
R1392 VDD.n572 VDD.n311 35.6179
R1393 VDD.n566 VDD.n311 35.6179
R1394 VDD.n566 VDD.n563 35.6179
R1395 VDD.n563 VDD.n316 35.6179
R1396 VDD.n559 VDD.n316 35.6179
R1397 VDD.n550 VDD.n547 35.6179
R1398 VDD.n547 VDD.n322 35.6179
R1399 VDD.n543 VDD.n322 35.6179
R1400 VDD.n543 VDD.n542 35.6179
R1401 VDD.n542 VDD.n327 35.6179
R1402 VDD.n536 VDD.n327 35.6179
R1403 VDD.n536 VDD.n533 35.6179
R1404 VDD.n533 VDD.n332 35.6179
R1405 VDD.n529 VDD.n332 35.6179
R1406 VDD.n529 VDD.n528 35.6179
R1407 VDD.n528 VDD.n337 35.6179
R1408 VDD.n522 VDD.n337 35.6179
R1409 VDD.n522 VDD.n519 35.6179
R1410 VDD.n519 VDD.n342 35.6179
R1411 VDD.n510 VDD.n509 35.6179
R1412 VDD.n509 VDD.n348 35.6179
R1413 VDD.n503 VDD.n348 35.6179
R1414 VDD.n503 VDD.n500 35.6179
R1415 VDD.n500 VDD.n353 35.6179
R1416 VDD.n496 VDD.n353 35.6179
R1417 VDD.n496 VDD.n495 35.6179
R1418 VDD.n495 VDD.n358 35.6179
R1419 VDD.n489 VDD.n358 35.6179
R1420 VDD.n489 VDD.n486 35.6179
R1421 VDD.n486 VDD.n363 35.6179
R1422 VDD.n482 VDD.n363 35.6179
R1423 VDD.n482 VDD.n481 35.6179
R1424 VDD.n481 VDD.n368 35.6179
R1425 VDD.n470 VDD.n467 35.6179
R1426 VDD.n467 VDD.n374 35.6179
R1427 VDD.n463 VDD.n374 35.6179
R1428 VDD.n463 VDD.n462 35.6179
R1429 VDD.n462 VDD.n379 35.6179
R1430 VDD.n456 VDD.n379 35.6179
R1431 VDD.n456 VDD.n453 35.6179
R1432 VDD.n453 VDD.n384 35.6179
R1433 VDD.n449 VDD.n384 35.6179
R1434 VDD.n449 VDD.n448 35.6179
R1435 VDD.n438 VDD.n437 35.6179
R1436 VDD.n437 VDD.n393 35.6179
R1437 VDD.n431 VDD.n393 35.6179
R1438 VDD.n431 VDD.n428 35.6179
R1439 VDD.n428 VDD.n399 35.6179
R1440 VDD.n424 VDD.n399 35.6179
R1441 VDD.n418 VDD.n403 35.6179
R1442 VDD.n414 VDD.n413 35.6179
R1443 VDD VDD.n411 1.543
R1444 VDD.n710 VDD.n709 0.3205
R1445 VDD.n639 VDD.n635 0.3205
R1446 VDD.n631 VDD.n630 0.3205
R1447 VDD.n560 VDD.n556 0.3205
R1448 VDD.n552 VDD.n551 0.3205
R1449 VDD.n517 VDD.n516 0.3205
R1450 VDD.n512 VDD.n511 0.3205
R1451 VDD.n477 VDD.n476 0.3205
R1452 VDD.n472 VDD.n471 0.3205
R1453 VDD.n445 VDD.n444 0.3205
R1454 VDD.n440 VDD.n439 0.3205
R1455 VDD.n425 VDD.n421 0.3205
R1456 VDD.n416 VDD.n415 0.3205
R1457 VDD.n6 VDD.n2 0.3205
R1458 VDD.n867 VDD.n866 0.3205
R1459 VDD.n862 VDD.n861 0.3205
R1460 VDD.n715 VDD.n714 0.3205
R1461 VDD.n709 VDD 0.248
R1462 VDD.n703 VDD 0.248
R1463 VDD.n697 VDD 0.248
R1464 VDD.n695 VDD 0.248
R1465 VDD.n689 VDD 0.248
R1466 VDD.n683 VDD 0.248
R1467 VDD.n681 VDD 0.248
R1468 VDD.n675 VDD 0.248
R1469 VDD.n669 VDD 0.248
R1470 VDD.n667 VDD 0.248
R1471 VDD.n661 VDD 0.248
R1472 VDD.n655 VDD 0.248
R1473 VDD.n653 VDD 0.248
R1474 VDD.n647 VDD 0.248
R1475 VDD.n641 VDD 0.248
R1476 VDD.n630 VDD 0.248
R1477 VDD.n624 VDD 0.248
R1478 VDD.n618 VDD 0.248
R1479 VDD.n616 VDD 0.248
R1480 VDD.n610 VDD 0.248
R1481 VDD.n604 VDD 0.248
R1482 VDD.n602 VDD 0.248
R1483 VDD.n596 VDD 0.248
R1484 VDD.n590 VDD 0.248
R1485 VDD.n588 VDD 0.248
R1486 VDD.n582 VDD 0.248
R1487 VDD.n576 VDD 0.248
R1488 VDD.n574 VDD 0.248
R1489 VDD.n568 VDD 0.248
R1490 VDD.n562 VDD 0.248
R1491 VDD.n551 VDD 0.248
R1492 VDD.n545 VDD 0.248
R1493 VDD.n539 VDD 0.248
R1494 VDD.n537 VDD 0.248
R1495 VDD.n531 VDD 0.248
R1496 VDD.n525 VDD 0.248
R1497 VDD.n523 VDD 0.248
R1498 VDD.n511 VDD 0.248
R1499 VDD.n505 VDD 0.248
R1500 VDD.n499 VDD 0.248
R1501 VDD.n497 VDD 0.248
R1502 VDD.n491 VDD 0.248
R1503 VDD.n485 VDD 0.248
R1504 VDD.n483 VDD 0.248
R1505 VDD.n471 VDD 0.248
R1506 VDD.n465 VDD 0.248
R1507 VDD.n459 VDD 0.248
R1508 VDD.n457 VDD 0.248
R1509 VDD.n451 VDD 0.248
R1510 VDD.n439 VDD 0.248
R1511 VDD.n433 VDD 0.248
R1512 VDD.n427 VDD 0.248
R1513 VDD.n417 VDD 0.248
R1514 VDD VDD.n6 0.248
R1515 VDD.n1007 VDD 0.248
R1516 VDD.n1005 VDD 0.248
R1517 VDD.n999 VDD 0.248
R1518 VDD.n993 VDD 0.248
R1519 VDD.n991 VDD 0.248
R1520 VDD.n985 VDD 0.248
R1521 VDD.n979 VDD 0.248
R1522 VDD.n977 VDD 0.248
R1523 VDD.n971 VDD 0.248
R1524 VDD.n965 VDD 0.248
R1525 VDD.n963 VDD 0.248
R1526 VDD.n957 VDD 0.248
R1527 VDD.n951 VDD 0.248
R1528 VDD.n949 VDD 0.248
R1529 VDD.n943 VDD 0.248
R1530 VDD.n937 VDD 0.248
R1531 VDD.n935 VDD 0.248
R1532 VDD.n929 VDD 0.248
R1533 VDD.n923 VDD 0.248
R1534 VDD.n921 VDD 0.248
R1535 VDD.n915 VDD 0.248
R1536 VDD.n909 VDD 0.248
R1537 VDD.n907 VDD 0.248
R1538 VDD.n901 VDD 0.248
R1539 VDD.n895 VDD 0.248
R1540 VDD.n893 VDD 0.248
R1541 VDD.n887 VDD 0.248
R1542 VDD.n881 VDD 0.248
R1543 VDD.n879 VDD 0.248
R1544 VDD.n873 VDD 0.248
R1545 VDD.n861 VDD 0.248
R1546 VDD.n855 VDD 0.248
R1547 VDD.n849 VDD 0.248
R1548 VDD.n847 VDD 0.248
R1549 VDD.n841 VDD 0.248
R1550 VDD.n835 VDD 0.248
R1551 VDD.n833 VDD 0.248
R1552 VDD.n827 VDD 0.248
R1553 VDD.n821 VDD 0.248
R1554 VDD.n819 VDD 0.248
R1555 VDD.n813 VDD 0.248
R1556 VDD.n807 VDD 0.248
R1557 VDD.n805 VDD 0.248
R1558 VDD.n799 VDD 0.248
R1559 VDD.n793 VDD 0.248
R1560 VDD.n791 VDD 0.248
R1561 VDD.n785 VDD 0.248
R1562 VDD.n779 VDD 0.248
R1563 VDD.n777 VDD 0.248
R1564 VDD.n771 VDD 0.248
R1565 VDD.n765 VDD 0.248
R1566 VDD.n763 VDD 0.248
R1567 VDD.n757 VDD 0.248
R1568 VDD.n751 VDD 0.248
R1569 VDD.n749 VDD 0.248
R1570 VDD.n743 VDD 0.248
R1571 VDD.n737 VDD 0.248
R1572 VDD.n735 VDD 0.248
R1573 VDD.n729 VDD 0.248
R1574 VDD.n723 VDD 0.248
R1575 VDD.n721 VDD 0.248
R1576 VDD VDD.n703 0.183
R1577 VDD.n697 VDD 0.183
R1578 VDD VDD.n695 0.183
R1579 VDD VDD.n689 0.183
R1580 VDD.n683 VDD 0.183
R1581 VDD VDD.n681 0.183
R1582 VDD VDD.n675 0.183
R1583 VDD.n669 VDD 0.183
R1584 VDD VDD.n667 0.183
R1585 VDD VDD.n661 0.183
R1586 VDD.n655 VDD 0.183
R1587 VDD VDD.n653 0.183
R1588 VDD VDD.n647 0.183
R1589 VDD.n641 VDD 0.183
R1590 VDD VDD.n639 0.183
R1591 VDD VDD.n624 0.183
R1592 VDD.n618 VDD 0.183
R1593 VDD VDD.n616 0.183
R1594 VDD VDD.n610 0.183
R1595 VDD.n604 VDD 0.183
R1596 VDD VDD.n602 0.183
R1597 VDD VDD.n596 0.183
R1598 VDD.n590 VDD 0.183
R1599 VDD VDD.n588 0.183
R1600 VDD VDD.n582 0.183
R1601 VDD.n576 VDD 0.183
R1602 VDD VDD.n574 0.183
R1603 VDD VDD.n568 0.183
R1604 VDD.n562 VDD 0.183
R1605 VDD VDD.n560 0.183
R1606 VDD VDD.n545 0.183
R1607 VDD.n539 VDD 0.183
R1608 VDD VDD.n537 0.183
R1609 VDD VDD.n531 0.183
R1610 VDD.n525 VDD 0.183
R1611 VDD VDD.n523 0.183
R1612 VDD VDD.n517 0.183
R1613 VDD VDD.n505 0.183
R1614 VDD.n499 VDD 0.183
R1615 VDD VDD.n497 0.183
R1616 VDD VDD.n491 0.183
R1617 VDD.n485 VDD 0.183
R1618 VDD VDD.n483 0.183
R1619 VDD VDD.n477 0.183
R1620 VDD VDD.n465 0.183
R1621 VDD.n459 VDD 0.183
R1622 VDD VDD.n457 0.183
R1623 VDD VDD.n451 0.183
R1624 VDD.n445 VDD 0.183
R1625 VDD VDD.n433 0.183
R1626 VDD.n427 VDD 0.183
R1627 VDD VDD.n425 0.183
R1628 VDD.n412 VDD 0.183
R1629 VDD.n1007 VDD 0.183
R1630 VDD VDD.n1005 0.183
R1631 VDD VDD.n999 0.183
R1632 VDD.n993 VDD 0.183
R1633 VDD VDD.n991 0.183
R1634 VDD VDD.n985 0.183
R1635 VDD.n979 VDD 0.183
R1636 VDD VDD.n977 0.183
R1637 VDD VDD.n971 0.183
R1638 VDD.n965 VDD 0.183
R1639 VDD VDD.n963 0.183
R1640 VDD VDD.n957 0.183
R1641 VDD.n951 VDD 0.183
R1642 VDD VDD.n949 0.183
R1643 VDD VDD.n943 0.183
R1644 VDD.n937 VDD 0.183
R1645 VDD VDD.n935 0.183
R1646 VDD VDD.n929 0.183
R1647 VDD.n923 VDD 0.183
R1648 VDD VDD.n921 0.183
R1649 VDD VDD.n915 0.183
R1650 VDD.n909 VDD 0.183
R1651 VDD VDD.n907 0.183
R1652 VDD VDD.n901 0.183
R1653 VDD.n895 VDD 0.183
R1654 VDD VDD.n893 0.183
R1655 VDD VDD.n887 0.183
R1656 VDD.n881 VDD 0.183
R1657 VDD VDD.n879 0.183
R1658 VDD VDD.n873 0.183
R1659 VDD.n867 VDD 0.183
R1660 VDD VDD.n855 0.183
R1661 VDD.n849 VDD 0.183
R1662 VDD VDD.n847 0.183
R1663 VDD VDD.n841 0.183
R1664 VDD.n835 VDD 0.183
R1665 VDD VDD.n833 0.183
R1666 VDD VDD.n827 0.183
R1667 VDD.n821 VDD 0.183
R1668 VDD VDD.n819 0.183
R1669 VDD VDD.n813 0.183
R1670 VDD.n807 VDD 0.183
R1671 VDD VDD.n805 0.183
R1672 VDD VDD.n799 0.183
R1673 VDD.n793 VDD 0.183
R1674 VDD VDD.n791 0.183
R1675 VDD VDD.n785 0.183
R1676 VDD.n779 VDD 0.183
R1677 VDD VDD.n777 0.183
R1678 VDD VDD.n771 0.183
R1679 VDD.n765 VDD 0.183
R1680 VDD VDD.n763 0.183
R1681 VDD VDD.n757 0.183
R1682 VDD.n751 VDD 0.183
R1683 VDD VDD.n749 0.183
R1684 VDD VDD.n743 0.183
R1685 VDD.n737 VDD 0.183
R1686 VDD VDD.n735 0.183
R1687 VDD VDD.n729 0.183
R1688 VDD.n723 VDD 0.183
R1689 VDD VDD.n721 0.183
R1690 VDD VDD.n715 0.183
R1691 VDD.n704 VDD 0.138
R1692 VDD.n702 VDD 0.138
R1693 VDD.n696 VDD 0.138
R1694 VDD.n690 VDD 0.138
R1695 VDD.n688 VDD 0.138
R1696 VDD.n682 VDD 0.138
R1697 VDD.n676 VDD 0.138
R1698 VDD.n674 VDD 0.138
R1699 VDD.n668 VDD 0.138
R1700 VDD.n662 VDD 0.138
R1701 VDD.n660 VDD 0.138
R1702 VDD.n654 VDD 0.138
R1703 VDD.n648 VDD 0.138
R1704 VDD.n646 VDD 0.138
R1705 VDD.n640 VDD 0.138
R1706 VDD.n635 VDD 0.138
R1707 VDD.n625 VDD 0.138
R1708 VDD.n623 VDD 0.138
R1709 VDD.n617 VDD 0.138
R1710 VDD.n611 VDD 0.138
R1711 VDD.n609 VDD 0.138
R1712 VDD.n603 VDD 0.138
R1713 VDD.n597 VDD 0.138
R1714 VDD.n595 VDD 0.138
R1715 VDD.n589 VDD 0.138
R1716 VDD.n583 VDD 0.138
R1717 VDD.n581 VDD 0.138
R1718 VDD.n575 VDD 0.138
R1719 VDD.n569 VDD 0.138
R1720 VDD.n567 VDD 0.138
R1721 VDD.n561 VDD 0.138
R1722 VDD.n556 VDD 0.138
R1723 VDD.n546 VDD 0.138
R1724 VDD.n544 VDD 0.138
R1725 VDD.n538 VDD 0.138
R1726 VDD.n532 VDD 0.138
R1727 VDD.n530 VDD 0.138
R1728 VDD.n524 VDD 0.138
R1729 VDD.n518 VDD 0.138
R1730 VDD.n516 VDD 0.138
R1731 VDD.n506 VDD 0.138
R1732 VDD.n504 VDD 0.138
R1733 VDD.n498 VDD 0.138
R1734 VDD.n492 VDD 0.138
R1735 VDD.n490 VDD 0.138
R1736 VDD.n484 VDD 0.138
R1737 VDD.n478 VDD 0.138
R1738 VDD.n476 VDD 0.138
R1739 VDD.n466 VDD 0.138
R1740 VDD.n464 VDD 0.138
R1741 VDD.n458 VDD 0.138
R1742 VDD.n452 VDD 0.138
R1743 VDD.n450 VDD 0.138
R1744 VDD.n444 VDD 0.138
R1745 VDD.n434 VDD 0.138
R1746 VDD.n432 VDD 0.138
R1747 VDD.n426 VDD 0.138
R1748 VDD.n421 VDD 0.138
R1749 VDD.n415 VDD 0.138
R1750 VDD.n412 VDD 0.138
R1751 VDD.n406 VDD 0.138
R1752 VDD.n1012 VDD 0.138
R1753 VDD.n1006 VDD 0.138
R1754 VDD.n1000 VDD 0.138
R1755 VDD.n998 VDD 0.138
R1756 VDD.n992 VDD 0.138
R1757 VDD.n986 VDD 0.138
R1758 VDD.n984 VDD 0.138
R1759 VDD.n978 VDD 0.138
R1760 VDD.n972 VDD 0.138
R1761 VDD.n970 VDD 0.138
R1762 VDD.n964 VDD 0.138
R1763 VDD.n958 VDD 0.138
R1764 VDD.n956 VDD 0.138
R1765 VDD.n950 VDD 0.138
R1766 VDD.n944 VDD 0.138
R1767 VDD.n942 VDD 0.138
R1768 VDD.n936 VDD 0.138
R1769 VDD.n930 VDD 0.138
R1770 VDD.n928 VDD 0.138
R1771 VDD.n922 VDD 0.138
R1772 VDD.n916 VDD 0.138
R1773 VDD.n914 VDD 0.138
R1774 VDD.n908 VDD 0.138
R1775 VDD.n902 VDD 0.138
R1776 VDD.n900 VDD 0.138
R1777 VDD.n894 VDD 0.138
R1778 VDD.n888 VDD 0.138
R1779 VDD.n886 VDD 0.138
R1780 VDD.n880 VDD 0.138
R1781 VDD.n874 VDD 0.138
R1782 VDD.n872 VDD 0.138
R1783 VDD.n866 VDD 0.138
R1784 VDD.n856 VDD 0.138
R1785 VDD.n854 VDD 0.138
R1786 VDD.n848 VDD 0.138
R1787 VDD.n842 VDD 0.138
R1788 VDD.n840 VDD 0.138
R1789 VDD.n834 VDD 0.138
R1790 VDD.n828 VDD 0.138
R1791 VDD.n826 VDD 0.138
R1792 VDD.n820 VDD 0.138
R1793 VDD.n814 VDD 0.138
R1794 VDD.n812 VDD 0.138
R1795 VDD.n806 VDD 0.138
R1796 VDD.n800 VDD 0.138
R1797 VDD.n798 VDD 0.138
R1798 VDD.n792 VDD 0.138
R1799 VDD.n786 VDD 0.138
R1800 VDD.n784 VDD 0.138
R1801 VDD.n778 VDD 0.138
R1802 VDD.n772 VDD 0.138
R1803 VDD.n770 VDD 0.138
R1804 VDD.n764 VDD 0.138
R1805 VDD.n758 VDD 0.138
R1806 VDD.n756 VDD 0.138
R1807 VDD.n750 VDD 0.138
R1808 VDD.n744 VDD 0.138
R1809 VDD.n742 VDD 0.138
R1810 VDD.n736 VDD 0.138
R1811 VDD.n730 VDD 0.138
R1812 VDD.n728 VDD 0.138
R1813 VDD.n722 VDD 0.138
R1814 VDD.n716 VDD 0.138
R1815 VDD.n714 VDD 0.138
R1816 VDD.n710 VDD 0.073
R1817 VDD.n704 VDD 0.073
R1818 VDD VDD.n702 0.073
R1819 VDD VDD.n696 0.073
R1820 VDD.n690 VDD 0.073
R1821 VDD VDD.n688 0.073
R1822 VDD VDD.n682 0.073
R1823 VDD.n676 VDD 0.073
R1824 VDD VDD.n674 0.073
R1825 VDD VDD.n668 0.073
R1826 VDD.n662 VDD 0.073
R1827 VDD VDD.n660 0.073
R1828 VDD VDD.n654 0.073
R1829 VDD.n648 VDD 0.073
R1830 VDD VDD.n646 0.073
R1831 VDD VDD.n640 0.073
R1832 VDD.n631 VDD 0.073
R1833 VDD.n625 VDD 0.073
R1834 VDD VDD.n623 0.073
R1835 VDD VDD.n617 0.073
R1836 VDD.n611 VDD 0.073
R1837 VDD VDD.n609 0.073
R1838 VDD VDD.n603 0.073
R1839 VDD.n597 VDD 0.073
R1840 VDD VDD.n595 0.073
R1841 VDD VDD.n589 0.073
R1842 VDD.n583 VDD 0.073
R1843 VDD VDD.n581 0.073
R1844 VDD VDD.n575 0.073
R1845 VDD.n569 VDD 0.073
R1846 VDD VDD.n567 0.073
R1847 VDD VDD.n561 0.073
R1848 VDD.n552 VDD 0.073
R1849 VDD.n546 VDD 0.073
R1850 VDD VDD.n544 0.073
R1851 VDD VDD.n538 0.073
R1852 VDD.n532 VDD 0.073
R1853 VDD VDD.n530 0.073
R1854 VDD VDD.n524 0.073
R1855 VDD.n518 VDD 0.073
R1856 VDD.n512 VDD 0.073
R1857 VDD.n506 VDD 0.073
R1858 VDD VDD.n504 0.073
R1859 VDD VDD.n498 0.073
R1860 VDD.n492 VDD 0.073
R1861 VDD VDD.n490 0.073
R1862 VDD VDD.n484 0.073
R1863 VDD.n478 VDD 0.073
R1864 VDD.n472 VDD 0.073
R1865 VDD.n466 VDD 0.073
R1866 VDD VDD.n464 0.073
R1867 VDD VDD.n458 0.073
R1868 VDD.n452 VDD 0.073
R1869 VDD VDD.n450 0.073
R1870 VDD.n440 VDD 0.073
R1871 VDD.n434 VDD 0.073
R1872 VDD VDD.n432 0.073
R1873 VDD VDD.n426 0.073
R1874 VDD.n417 VDD 0.073
R1875 VDD VDD.n416 0.073
R1876 VDD.n2 VDD 0.073
R1877 VDD VDD.n1012 0.073
R1878 VDD VDD.n1006 0.073
R1879 VDD.n1000 VDD 0.073
R1880 VDD VDD.n998 0.073
R1881 VDD VDD.n992 0.073
R1882 VDD.n986 VDD 0.073
R1883 VDD VDD.n984 0.073
R1884 VDD VDD.n978 0.073
R1885 VDD.n972 VDD 0.073
R1886 VDD VDD.n970 0.073
R1887 VDD VDD.n964 0.073
R1888 VDD.n958 VDD 0.073
R1889 VDD VDD.n956 0.073
R1890 VDD VDD.n950 0.073
R1891 VDD.n944 VDD 0.073
R1892 VDD VDD.n942 0.073
R1893 VDD VDD.n936 0.073
R1894 VDD.n930 VDD 0.073
R1895 VDD VDD.n928 0.073
R1896 VDD VDD.n922 0.073
R1897 VDD.n916 VDD 0.073
R1898 VDD VDD.n914 0.073
R1899 VDD VDD.n908 0.073
R1900 VDD.n902 VDD 0.073
R1901 VDD VDD.n900 0.073
R1902 VDD VDD.n894 0.073
R1903 VDD.n888 VDD 0.073
R1904 VDD VDD.n886 0.073
R1905 VDD VDD.n880 0.073
R1906 VDD.n874 VDD 0.073
R1907 VDD VDD.n872 0.073
R1908 VDD.n862 VDD 0.073
R1909 VDD.n856 VDD 0.073
R1910 VDD VDD.n854 0.073
R1911 VDD VDD.n848 0.073
R1912 VDD.n842 VDD 0.073
R1913 VDD VDD.n840 0.073
R1914 VDD VDD.n834 0.073
R1915 VDD.n828 VDD 0.073
R1916 VDD VDD.n826 0.073
R1917 VDD VDD.n820 0.073
R1918 VDD.n814 VDD 0.073
R1919 VDD VDD.n812 0.073
R1920 VDD VDD.n806 0.073
R1921 VDD.n800 VDD 0.073
R1922 VDD VDD.n798 0.073
R1923 VDD VDD.n792 0.073
R1924 VDD.n786 VDD 0.073
R1925 VDD VDD.n784 0.073
R1926 VDD VDD.n778 0.073
R1927 VDD.n772 VDD 0.073
R1928 VDD VDD.n770 0.073
R1929 VDD VDD.n764 0.073
R1930 VDD.n758 VDD 0.073
R1931 VDD VDD.n756 0.073
R1932 VDD VDD.n750 0.073
R1933 VDD.n744 VDD 0.073
R1934 VDD VDD.n742 0.073
R1935 VDD VDD.n736 0.073
R1936 VDD.n730 VDD 0.073
R1937 VDD VDD.n728 0.073
R1938 VDD VDD.n722 0.073
R1939 VDD.n716 VDD 0.073
R1940 VDD.n408 VDD.n406 0.00452048
R1941 VDD.n409 VDD.n408 0.00383931
R1942 VDD.n413 VDD.n410 0.00166989
R1943 VDD.n420 VDD.n419 0.00166989
R1944 VDD.n475 VDD.n474 0.00166989
R1945 VDD.n555 VDD.n554 0.00166989
R1946 VDD.n713 VDD.n712 0.00166989
R1947 VDD.n1 VDD.n0 0.00166989
R1948 VDD.n711 VDD.n215 0.00166989
R1949 VDD.n553 VDD.n317 0.00166989
R1950 VDD.n473 VDD.n369 0.00166989
R1951 VDD.n708 VDD.n707 0.00166989
R1952 VDD.n707 VDD.n706 0.00166989
R1953 VDD.n705 VDD.n217 0.00166989
R1954 VDD.n217 VDD.n216 0.00166989
R1955 VDD.n220 VDD.n219 0.00166989
R1956 VDD.n219 VDD.n218 0.00166989
R1957 VDD.n701 VDD.n222 0.00166989
R1958 VDD.n222 VDD.n221 0.00166989
R1959 VDD.n700 VDD.n699 0.00166989
R1960 VDD.n699 VDD.n698 0.00166989
R1961 VDD.n225 VDD.n224 0.00166989
R1962 VDD.n224 VDD.n223 0.00166989
R1963 VDD.n694 VDD.n693 0.00166989
R1964 VDD.n693 VDD.n692 0.00166989
R1965 VDD.n691 VDD.n227 0.00166989
R1966 VDD.n227 VDD.n226 0.00166989
R1967 VDD.n230 VDD.n229 0.00166989
R1968 VDD.n229 VDD.n228 0.00166989
R1969 VDD.n687 VDD.n232 0.00166989
R1970 VDD.n232 VDD.n231 0.00166989
R1971 VDD.n686 VDD.n685 0.00166989
R1972 VDD.n685 VDD.n684 0.00166989
R1973 VDD.n235 VDD.n234 0.00166989
R1974 VDD.n234 VDD.n233 0.00166989
R1975 VDD.n680 VDD.n679 0.00166989
R1976 VDD.n679 VDD.n678 0.00166989
R1977 VDD.n677 VDD.n237 0.00166989
R1978 VDD.n237 VDD.n236 0.00166989
R1979 VDD.n240 VDD.n239 0.00166989
R1980 VDD.n239 VDD.n238 0.00166989
R1981 VDD.n673 VDD.n242 0.00166989
R1982 VDD.n242 VDD.n241 0.00166989
R1983 VDD.n672 VDD.n671 0.00166989
R1984 VDD.n671 VDD.n670 0.00166989
R1985 VDD.n245 VDD.n244 0.00166989
R1986 VDD.n244 VDD.n243 0.00166989
R1987 VDD.n666 VDD.n665 0.00166989
R1988 VDD.n665 VDD.n664 0.00166989
R1989 VDD.n663 VDD.n247 0.00166989
R1990 VDD.n247 VDD.n246 0.00166989
R1991 VDD.n250 VDD.n249 0.00166989
R1992 VDD.n249 VDD.n248 0.00166989
R1993 VDD.n659 VDD.n252 0.00166989
R1994 VDD.n252 VDD.n251 0.00166989
R1995 VDD.n658 VDD.n657 0.00166989
R1996 VDD.n657 VDD.n656 0.00166989
R1997 VDD.n255 VDD.n254 0.00166989
R1998 VDD.n254 VDD.n253 0.00166989
R1999 VDD.n652 VDD.n651 0.00166989
R2000 VDD.n651 VDD.n650 0.00166989
R2001 VDD.n649 VDD.n257 0.00166989
R2002 VDD.n257 VDD.n256 0.00166989
R2003 VDD.n260 VDD.n259 0.00166989
R2004 VDD.n259 VDD.n258 0.00166989
R2005 VDD.n645 VDD.n262 0.00166989
R2006 VDD.n262 VDD.n261 0.00166989
R2007 VDD.n644 VDD.n643 0.00166989
R2008 VDD.n643 VDD.n642 0.00166989
R2009 VDD.n265 VDD.n264 0.00166989
R2010 VDD.n264 VDD.n263 0.00166989
R2011 VDD.n638 VDD.n637 0.00166989
R2012 VDD.n637 VDD.n636 0.00166989
R2013 VDD.n634 VDD.n266 0.00166989
R2014 VDD.n633 VDD.n632 0.00166989
R2015 VDD.n629 VDD.n268 0.00166989
R2016 VDD.n268 VDD.n267 0.00166989
R2017 VDD.n628 VDD.n627 0.00166989
R2018 VDD.n627 VDD.n626 0.00166989
R2019 VDD.n271 VDD.n270 0.00166989
R2020 VDD.n270 VDD.n269 0.00166989
R2021 VDD.n622 VDD.n621 0.00166989
R2022 VDD.n621 VDD.n620 0.00166989
R2023 VDD.n619 VDD.n273 0.00166989
R2024 VDD.n273 VDD.n272 0.00166989
R2025 VDD.n276 VDD.n275 0.00166989
R2026 VDD.n275 VDD.n274 0.00166989
R2027 VDD.n615 VDD.n278 0.00166989
R2028 VDD.n278 VDD.n277 0.00166989
R2029 VDD.n614 VDD.n613 0.00166989
R2030 VDD.n613 VDD.n612 0.00166989
R2031 VDD.n281 VDD.n280 0.00166989
R2032 VDD.n280 VDD.n279 0.00166989
R2033 VDD.n608 VDD.n607 0.00166989
R2034 VDD.n607 VDD.n606 0.00166989
R2035 VDD.n605 VDD.n283 0.00166989
R2036 VDD.n283 VDD.n282 0.00166989
R2037 VDD.n286 VDD.n285 0.00166989
R2038 VDD.n285 VDD.n284 0.00166989
R2039 VDD.n601 VDD.n288 0.00166989
R2040 VDD.n288 VDD.n287 0.00166989
R2041 VDD.n600 VDD.n599 0.00166989
R2042 VDD.n599 VDD.n598 0.00166989
R2043 VDD.n291 VDD.n290 0.00166989
R2044 VDD.n290 VDD.n289 0.00166989
R2045 VDD.n594 VDD.n593 0.00166989
R2046 VDD.n593 VDD.n592 0.00166989
R2047 VDD.n591 VDD.n293 0.00166989
R2048 VDD.n293 VDD.n292 0.00166989
R2049 VDD.n296 VDD.n295 0.00166989
R2050 VDD.n295 VDD.n294 0.00166989
R2051 VDD.n587 VDD.n298 0.00166989
R2052 VDD.n298 VDD.n297 0.00166989
R2053 VDD.n586 VDD.n585 0.00166989
R2054 VDD.n585 VDD.n584 0.00166989
R2055 VDD.n301 VDD.n300 0.00166989
R2056 VDD.n300 VDD.n299 0.00166989
R2057 VDD.n580 VDD.n579 0.00166989
R2058 VDD.n579 VDD.n578 0.00166989
R2059 VDD.n577 VDD.n303 0.00166989
R2060 VDD.n303 VDD.n302 0.00166989
R2061 VDD.n306 VDD.n305 0.00166989
R2062 VDD.n305 VDD.n304 0.00166989
R2063 VDD.n573 VDD.n308 0.00166989
R2064 VDD.n308 VDD.n307 0.00166989
R2065 VDD.n572 VDD.n571 0.00166989
R2066 VDD.n571 VDD.n570 0.00166989
R2067 VDD.n311 VDD.n310 0.00166989
R2068 VDD.n310 VDD.n309 0.00166989
R2069 VDD.n566 VDD.n565 0.00166989
R2070 VDD.n565 VDD.n564 0.00166989
R2071 VDD.n563 VDD.n313 0.00166989
R2072 VDD.n313 VDD.n312 0.00166989
R2073 VDD.n316 VDD.n315 0.00166989
R2074 VDD.n315 VDD.n314 0.00166989
R2075 VDD.n559 VDD.n558 0.00166989
R2076 VDD.n558 VDD.n557 0.00166989
R2077 VDD.n550 VDD.n549 0.00166989
R2078 VDD.n549 VDD.n548 0.00166989
R2079 VDD.n547 VDD.n319 0.00166989
R2080 VDD.n319 VDD.n318 0.00166989
R2081 VDD.n322 VDD.n321 0.00166989
R2082 VDD.n321 VDD.n320 0.00166989
R2083 VDD.n543 VDD.n324 0.00166989
R2084 VDD.n324 VDD.n323 0.00166989
R2085 VDD.n542 VDD.n541 0.00166989
R2086 VDD.n541 VDD.n540 0.00166989
R2087 VDD.n327 VDD.n326 0.00166989
R2088 VDD.n326 VDD.n325 0.00166989
R2089 VDD.n536 VDD.n535 0.00166989
R2090 VDD.n535 VDD.n534 0.00166989
R2091 VDD.n533 VDD.n329 0.00166989
R2092 VDD.n329 VDD.n328 0.00166989
R2093 VDD.n332 VDD.n331 0.00166989
R2094 VDD.n331 VDD.n330 0.00166989
R2095 VDD.n529 VDD.n334 0.00166989
R2096 VDD.n334 VDD.n333 0.00166989
R2097 VDD.n528 VDD.n527 0.00166989
R2098 VDD.n527 VDD.n526 0.00166989
R2099 VDD.n337 VDD.n336 0.00166989
R2100 VDD.n336 VDD.n335 0.00166989
R2101 VDD.n522 VDD.n521 0.00166989
R2102 VDD.n521 VDD.n520 0.00166989
R2103 VDD.n519 VDD.n339 0.00166989
R2104 VDD.n339 VDD.n338 0.00166989
R2105 VDD.n342 VDD.n341 0.00166989
R2106 VDD.n341 VDD.n340 0.00166989
R2107 VDD.n515 VDD.n343 0.00166989
R2108 VDD.n514 VDD.n513 0.00166989
R2109 VDD.n510 VDD.n345 0.00166989
R2110 VDD.n345 VDD.n344 0.00166989
R2111 VDD.n509 VDD.n508 0.00166989
R2112 VDD.n508 VDD.n507 0.00166989
R2113 VDD.n348 VDD.n347 0.00166989
R2114 VDD.n347 VDD.n346 0.00166989
R2115 VDD.n503 VDD.n502 0.00166989
R2116 VDD.n502 VDD.n501 0.00166989
R2117 VDD.n500 VDD.n350 0.00166989
R2118 VDD.n350 VDD.n349 0.00166989
R2119 VDD.n353 VDD.n352 0.00166989
R2120 VDD.n352 VDD.n351 0.00166989
R2121 VDD.n496 VDD.n355 0.00166989
R2122 VDD.n355 VDD.n354 0.00166989
R2123 VDD.n495 VDD.n494 0.00166989
R2124 VDD.n494 VDD.n493 0.00166989
R2125 VDD.n358 VDD.n357 0.00166989
R2126 VDD.n357 VDD.n356 0.00166989
R2127 VDD.n489 VDD.n488 0.00166989
R2128 VDD.n488 VDD.n487 0.00166989
R2129 VDD.n486 VDD.n360 0.00166989
R2130 VDD.n360 VDD.n359 0.00166989
R2131 VDD.n363 VDD.n362 0.00166989
R2132 VDD.n362 VDD.n361 0.00166989
R2133 VDD.n482 VDD.n365 0.00166989
R2134 VDD.n365 VDD.n364 0.00166989
R2135 VDD.n481 VDD.n480 0.00166989
R2136 VDD.n480 VDD.n479 0.00166989
R2137 VDD.n368 VDD.n367 0.00166989
R2138 VDD.n367 VDD.n366 0.00166989
R2139 VDD.n470 VDD.n469 0.00166989
R2140 VDD.n469 VDD.n468 0.00166989
R2141 VDD.n467 VDD.n371 0.00166989
R2142 VDD.n371 VDD.n370 0.00166989
R2143 VDD.n374 VDD.n373 0.00166989
R2144 VDD.n373 VDD.n372 0.00166989
R2145 VDD.n463 VDD.n376 0.00166989
R2146 VDD.n376 VDD.n375 0.00166989
R2147 VDD.n462 VDD.n461 0.00166989
R2148 VDD.n461 VDD.n460 0.00166989
R2149 VDD.n379 VDD.n378 0.00166989
R2150 VDD.n378 VDD.n377 0.00166989
R2151 VDD.n456 VDD.n455 0.00166989
R2152 VDD.n455 VDD.n454 0.00166989
R2153 VDD.n453 VDD.n381 0.00166989
R2154 VDD.n381 VDD.n380 0.00166989
R2155 VDD.n384 VDD.n383 0.00166989
R2156 VDD.n383 VDD.n382 0.00166989
R2157 VDD.n449 VDD.n386 0.00166989
R2158 VDD.n386 VDD.n385 0.00166989
R2159 VDD.n448 VDD.n447 0.00166989
R2160 VDD.n447 VDD.n446 0.00166989
R2161 VDD.n443 VDD.n387 0.00166989
R2162 VDD.n442 VDD.n441 0.00166989
R2163 VDD.n438 VDD.n389 0.00166989
R2164 VDD.n389 VDD.n388 0.00166989
R2165 VDD.n437 VDD.n436 0.00166989
R2166 VDD.n436 VDD.n435 0.00166989
R2167 VDD.n393 VDD.n392 0.00166989
R2168 VDD.n392 VDD.n391 0.00166989
R2169 VDD.n431 VDD.n430 0.00166989
R2170 VDD.n430 VDD.n429 0.00166989
R2171 VDD.n428 VDD.n396 0.00166989
R2172 VDD.n396 VDD.n395 0.00166989
R2173 VDD.n399 VDD.n398 0.00166989
R2174 VDD.n398 VDD.n397 0.00166989
R2175 VDD.n424 VDD.n423 0.00166989
R2176 VDD.n423 VDD.n422 0.00166989
R2177 VDD.n418 VDD.n400 0.00166989
R2178 VDD.n403 VDD.n402 0.00166989
R2179 VDD.n402 VDD.n401 0.00166989
R2180 VDD.n414 VDD.n405 0.00166989
R2181 VDD.n405 VDD.n404 0.00166989
R2182 VDD.n5 VDD.n4 0.00166989
R2183 VDD.n4 VDD.n3 0.00166989
R2184 VDD.n1011 VDD.n8 0.00166989
R2185 VDD.n8 VDD.n7 0.00166989
R2186 VDD.n1010 VDD.n1009 0.00166989
R2187 VDD.n1009 VDD.n1008 0.00166989
R2188 VDD.n11 VDD.n10 0.00166989
R2189 VDD.n10 VDD.n9 0.00166989
R2190 VDD.n1004 VDD.n1003 0.00166989
R2191 VDD.n1003 VDD.n1002 0.00166989
R2192 VDD.n1001 VDD.n13 0.00166989
R2193 VDD.n13 VDD.n12 0.00166989
R2194 VDD.n16 VDD.n15 0.00166989
R2195 VDD.n15 VDD.n14 0.00166989
R2196 VDD.n997 VDD.n18 0.00166989
R2197 VDD.n18 VDD.n17 0.00166989
R2198 VDD.n996 VDD.n995 0.00166989
R2199 VDD.n995 VDD.n994 0.00166989
R2200 VDD.n21 VDD.n20 0.00166989
R2201 VDD.n20 VDD.n19 0.00166989
R2202 VDD.n990 VDD.n989 0.00166989
R2203 VDD.n989 VDD.n988 0.00166989
R2204 VDD.n987 VDD.n23 0.00166989
R2205 VDD.n23 VDD.n22 0.00166989
R2206 VDD.n26 VDD.n25 0.00166989
R2207 VDD.n25 VDD.n24 0.00166989
R2208 VDD.n983 VDD.n28 0.00166989
R2209 VDD.n28 VDD.n27 0.00166989
R2210 VDD.n982 VDD.n981 0.00166989
R2211 VDD.n981 VDD.n980 0.00166989
R2212 VDD.n31 VDD.n30 0.00166989
R2213 VDD.n30 VDD.n29 0.00166989
R2214 VDD.n976 VDD.n975 0.00166989
R2215 VDD.n975 VDD.n974 0.00166989
R2216 VDD.n973 VDD.n33 0.00166989
R2217 VDD.n33 VDD.n32 0.00166989
R2218 VDD.n36 VDD.n35 0.00166989
R2219 VDD.n35 VDD.n34 0.00166989
R2220 VDD.n969 VDD.n38 0.00166989
R2221 VDD.n38 VDD.n37 0.00166989
R2222 VDD.n968 VDD.n967 0.00166989
R2223 VDD.n967 VDD.n966 0.00166989
R2224 VDD.n41 VDD.n40 0.00166989
R2225 VDD.n40 VDD.n39 0.00166989
R2226 VDD.n962 VDD.n961 0.00166989
R2227 VDD.n961 VDD.n960 0.00166989
R2228 VDD.n959 VDD.n43 0.00166989
R2229 VDD.n43 VDD.n42 0.00166989
R2230 VDD.n46 VDD.n45 0.00166989
R2231 VDD.n45 VDD.n44 0.00166989
R2232 VDD.n955 VDD.n48 0.00166989
R2233 VDD.n48 VDD.n47 0.00166989
R2234 VDD.n954 VDD.n953 0.00166989
R2235 VDD.n953 VDD.n952 0.00166989
R2236 VDD.n51 VDD.n50 0.00166989
R2237 VDD.n50 VDD.n49 0.00166989
R2238 VDD.n948 VDD.n947 0.00166989
R2239 VDD.n947 VDD.n946 0.00166989
R2240 VDD.n945 VDD.n53 0.00166989
R2241 VDD.n53 VDD.n52 0.00166989
R2242 VDD.n56 VDD.n55 0.00166989
R2243 VDD.n55 VDD.n54 0.00166989
R2244 VDD.n941 VDD.n58 0.00166989
R2245 VDD.n58 VDD.n57 0.00166989
R2246 VDD.n940 VDD.n939 0.00166989
R2247 VDD.n939 VDD.n938 0.00166989
R2248 VDD.n61 VDD.n60 0.00166989
R2249 VDD.n60 VDD.n59 0.00166989
R2250 VDD.n934 VDD.n933 0.00166989
R2251 VDD.n933 VDD.n932 0.00166989
R2252 VDD.n931 VDD.n63 0.00166989
R2253 VDD.n63 VDD.n62 0.00166989
R2254 VDD.n66 VDD.n65 0.00166989
R2255 VDD.n65 VDD.n64 0.00166989
R2256 VDD.n927 VDD.n68 0.00166989
R2257 VDD.n68 VDD.n67 0.00166989
R2258 VDD.n926 VDD.n925 0.00166989
R2259 VDD.n925 VDD.n924 0.00166989
R2260 VDD.n71 VDD.n70 0.00166989
R2261 VDD.n70 VDD.n69 0.00166989
R2262 VDD.n920 VDD.n919 0.00166989
R2263 VDD.n919 VDD.n918 0.00166989
R2264 VDD.n917 VDD.n73 0.00166989
R2265 VDD.n73 VDD.n72 0.00166989
R2266 VDD.n76 VDD.n75 0.00166989
R2267 VDD.n75 VDD.n74 0.00166989
R2268 VDD.n913 VDD.n78 0.00166989
R2269 VDD.n78 VDD.n77 0.00166989
R2270 VDD.n912 VDD.n911 0.00166989
R2271 VDD.n911 VDD.n910 0.00166989
R2272 VDD.n81 VDD.n80 0.00166989
R2273 VDD.n80 VDD.n79 0.00166989
R2274 VDD.n906 VDD.n905 0.00166989
R2275 VDD.n905 VDD.n904 0.00166989
R2276 VDD.n903 VDD.n83 0.00166989
R2277 VDD.n83 VDD.n82 0.00166989
R2278 VDD.n86 VDD.n85 0.00166989
R2279 VDD.n85 VDD.n84 0.00166989
R2280 VDD.n899 VDD.n88 0.00166989
R2281 VDD.n88 VDD.n87 0.00166989
R2282 VDD.n898 VDD.n897 0.00166989
R2283 VDD.n897 VDD.n896 0.00166989
R2284 VDD.n91 VDD.n90 0.00166989
R2285 VDD.n90 VDD.n89 0.00166989
R2286 VDD.n892 VDD.n891 0.00166989
R2287 VDD.n891 VDD.n890 0.00166989
R2288 VDD.n889 VDD.n93 0.00166989
R2289 VDD.n93 VDD.n92 0.00166989
R2290 VDD.n96 VDD.n95 0.00166989
R2291 VDD.n95 VDD.n94 0.00166989
R2292 VDD.n885 VDD.n98 0.00166989
R2293 VDD.n98 VDD.n97 0.00166989
R2294 VDD.n884 VDD.n883 0.00166989
R2295 VDD.n883 VDD.n882 0.00166989
R2296 VDD.n101 VDD.n100 0.00166989
R2297 VDD.n100 VDD.n99 0.00166989
R2298 VDD.n878 VDD.n877 0.00166989
R2299 VDD.n877 VDD.n876 0.00166989
R2300 VDD.n875 VDD.n103 0.00166989
R2301 VDD.n103 VDD.n102 0.00166989
R2302 VDD.n106 VDD.n105 0.00166989
R2303 VDD.n105 VDD.n104 0.00166989
R2304 VDD.n871 VDD.n108 0.00166989
R2305 VDD.n108 VDD.n107 0.00166989
R2306 VDD.n870 VDD.n869 0.00166989
R2307 VDD.n869 VDD.n868 0.00166989
R2308 VDD.n865 VDD.n109 0.00166989
R2309 VDD.n864 VDD.n863 0.00166989
R2310 VDD.n860 VDD.n111 0.00166989
R2311 VDD.n111 VDD.n110 0.00166989
R2312 VDD.n859 VDD.n858 0.00166989
R2313 VDD.n858 VDD.n857 0.00166989
R2314 VDD.n114 VDD.n113 0.00166989
R2315 VDD.n113 VDD.n112 0.00166989
R2316 VDD.n853 VDD.n852 0.00166989
R2317 VDD.n852 VDD.n851 0.00166989
R2318 VDD.n850 VDD.n116 0.00166989
R2319 VDD.n116 VDD.n115 0.00166989
R2320 VDD.n119 VDD.n118 0.00166989
R2321 VDD.n118 VDD.n117 0.00166989
R2322 VDD.n846 VDD.n121 0.00166989
R2323 VDD.n121 VDD.n120 0.00166989
R2324 VDD.n845 VDD.n844 0.00166989
R2325 VDD.n844 VDD.n843 0.00166989
R2326 VDD.n124 VDD.n123 0.00166989
R2327 VDD.n123 VDD.n122 0.00166989
R2328 VDD.n839 VDD.n838 0.00166989
R2329 VDD.n838 VDD.n837 0.00166989
R2330 VDD.n836 VDD.n126 0.00166989
R2331 VDD.n126 VDD.n125 0.00166989
R2332 VDD.n129 VDD.n128 0.00166989
R2333 VDD.n128 VDD.n127 0.00166989
R2334 VDD.n832 VDD.n131 0.00166989
R2335 VDD.n131 VDD.n130 0.00166989
R2336 VDD.n831 VDD.n830 0.00166989
R2337 VDD.n830 VDD.n829 0.00166989
R2338 VDD.n134 VDD.n133 0.00166989
R2339 VDD.n133 VDD.n132 0.00166989
R2340 VDD.n825 VDD.n824 0.00166989
R2341 VDD.n824 VDD.n823 0.00166989
R2342 VDD.n822 VDD.n136 0.00166989
R2343 VDD.n136 VDD.n135 0.00166989
R2344 VDD.n139 VDD.n138 0.00166989
R2345 VDD.n138 VDD.n137 0.00166989
R2346 VDD.n818 VDD.n141 0.00166989
R2347 VDD.n141 VDD.n140 0.00166989
R2348 VDD.n817 VDD.n816 0.00166989
R2349 VDD.n816 VDD.n815 0.00166989
R2350 VDD.n144 VDD.n143 0.00166989
R2351 VDD.n143 VDD.n142 0.00166989
R2352 VDD.n811 VDD.n810 0.00166989
R2353 VDD.n810 VDD.n809 0.00166989
R2354 VDD.n808 VDD.n146 0.00166989
R2355 VDD.n146 VDD.n145 0.00166989
R2356 VDD.n149 VDD.n148 0.00166989
R2357 VDD.n148 VDD.n147 0.00166989
R2358 VDD.n804 VDD.n151 0.00166989
R2359 VDD.n151 VDD.n150 0.00166989
R2360 VDD.n803 VDD.n802 0.00166989
R2361 VDD.n802 VDD.n801 0.00166989
R2362 VDD.n154 VDD.n153 0.00166989
R2363 VDD.n153 VDD.n152 0.00166989
R2364 VDD.n797 VDD.n796 0.00166989
R2365 VDD.n796 VDD.n795 0.00166989
R2366 VDD.n794 VDD.n156 0.00166989
R2367 VDD.n156 VDD.n155 0.00166989
R2368 VDD.n159 VDD.n158 0.00166989
R2369 VDD.n158 VDD.n157 0.00166989
R2370 VDD.n790 VDD.n161 0.00166989
R2371 VDD.n161 VDD.n160 0.00166989
R2372 VDD.n789 VDD.n788 0.00166989
R2373 VDD.n788 VDD.n787 0.00166989
R2374 VDD.n164 VDD.n163 0.00166989
R2375 VDD.n163 VDD.n162 0.00166989
R2376 VDD.n783 VDD.n782 0.00166989
R2377 VDD.n782 VDD.n781 0.00166989
R2378 VDD.n780 VDD.n166 0.00166989
R2379 VDD.n166 VDD.n165 0.00166989
R2380 VDD.n169 VDD.n168 0.00166989
R2381 VDD.n168 VDD.n167 0.00166989
R2382 VDD.n776 VDD.n171 0.00166989
R2383 VDD.n171 VDD.n170 0.00166989
R2384 VDD.n775 VDD.n774 0.00166989
R2385 VDD.n774 VDD.n773 0.00166989
R2386 VDD.n174 VDD.n173 0.00166989
R2387 VDD.n173 VDD.n172 0.00166989
R2388 VDD.n769 VDD.n768 0.00166989
R2389 VDD.n768 VDD.n767 0.00166989
R2390 VDD.n766 VDD.n176 0.00166989
R2391 VDD.n176 VDD.n175 0.00166989
R2392 VDD.n179 VDD.n178 0.00166989
R2393 VDD.n178 VDD.n177 0.00166989
R2394 VDD.n762 VDD.n181 0.00166989
R2395 VDD.n181 VDD.n180 0.00166989
R2396 VDD.n761 VDD.n760 0.00166989
R2397 VDD.n760 VDD.n759 0.00166989
R2398 VDD.n184 VDD.n183 0.00166989
R2399 VDD.n183 VDD.n182 0.00166989
R2400 VDD.n755 VDD.n754 0.00166989
R2401 VDD.n754 VDD.n753 0.00166989
R2402 VDD.n752 VDD.n186 0.00166989
R2403 VDD.n186 VDD.n185 0.00166989
R2404 VDD.n189 VDD.n188 0.00166989
R2405 VDD.n188 VDD.n187 0.00166989
R2406 VDD.n748 VDD.n191 0.00166989
R2407 VDD.n191 VDD.n190 0.00166989
R2408 VDD.n747 VDD.n746 0.00166989
R2409 VDD.n746 VDD.n745 0.00166989
R2410 VDD.n194 VDD.n193 0.00166989
R2411 VDD.n193 VDD.n192 0.00166989
R2412 VDD.n741 VDD.n740 0.00166989
R2413 VDD.n740 VDD.n739 0.00166989
R2414 VDD.n738 VDD.n196 0.00166989
R2415 VDD.n196 VDD.n195 0.00166989
R2416 VDD.n199 VDD.n198 0.00166989
R2417 VDD.n198 VDD.n197 0.00166989
R2418 VDD.n734 VDD.n201 0.00166989
R2419 VDD.n201 VDD.n200 0.00166989
R2420 VDD.n733 VDD.n732 0.00166989
R2421 VDD.n732 VDD.n731 0.00166989
R2422 VDD.n204 VDD.n203 0.00166989
R2423 VDD.n203 VDD.n202 0.00166989
R2424 VDD.n727 VDD.n726 0.00166989
R2425 VDD.n726 VDD.n725 0.00166989
R2426 VDD.n724 VDD.n206 0.00166989
R2427 VDD.n206 VDD.n205 0.00166989
R2428 VDD.n209 VDD.n208 0.00166989
R2429 VDD.n208 VDD.n207 0.00166989
R2430 VDD.n720 VDD.n211 0.00166989
R2431 VDD.n211 VDD.n210 0.00166989
R2432 VDD.n719 VDD.n718 0.00166989
R2433 VDD.n718 VDD.n717 0.00166989
R2434 VDD.n214 VDD.n213 0.00166989
R2435 VDD.n213 VDD.n212 0.00166989
R2436 VDD.n408 VDD.n407 0.00150023
R2437 VDD.n711 VDD.n710 0.00118117
R2438 VDD.n709 VDD.n708 0.00118117
R2439 VDD.n705 VDD.n704 0.00118117
R2440 VDD.n703 VDD.n220 0.00118117
R2441 VDD.n702 VDD.n701 0.00118117
R2442 VDD.n700 VDD.n697 0.00118117
R2443 VDD.n696 VDD.n225 0.00118117
R2444 VDD.n695 VDD.n694 0.00118117
R2445 VDD.n691 VDD.n690 0.00118117
R2446 VDD.n689 VDD.n230 0.00118117
R2447 VDD.n688 VDD.n687 0.00118117
R2448 VDD.n686 VDD.n683 0.00118117
R2449 VDD.n682 VDD.n235 0.00118117
R2450 VDD.n681 VDD.n680 0.00118117
R2451 VDD.n677 VDD.n676 0.00118117
R2452 VDD.n675 VDD.n240 0.00118117
R2453 VDD.n674 VDD.n673 0.00118117
R2454 VDD.n672 VDD.n669 0.00118117
R2455 VDD.n668 VDD.n245 0.00118117
R2456 VDD.n667 VDD.n666 0.00118117
R2457 VDD.n663 VDD.n662 0.00118117
R2458 VDD.n661 VDD.n250 0.00118117
R2459 VDD.n660 VDD.n659 0.00118117
R2460 VDD.n658 VDD.n655 0.00118117
R2461 VDD.n654 VDD.n255 0.00118117
R2462 VDD.n653 VDD.n652 0.00118117
R2463 VDD.n649 VDD.n648 0.00118117
R2464 VDD.n647 VDD.n260 0.00118117
R2465 VDD.n646 VDD.n645 0.00118117
R2466 VDD.n644 VDD.n641 0.00118117
R2467 VDD.n640 VDD.n265 0.00118117
R2468 VDD.n639 VDD.n638 0.00118117
R2469 VDD.n635 VDD.n634 0.00118117
R2470 VDD.n633 VDD.n631 0.00118117
R2471 VDD.n630 VDD.n629 0.00118117
R2472 VDD.n628 VDD.n625 0.00118117
R2473 VDD.n624 VDD.n271 0.00118117
R2474 VDD.n623 VDD.n622 0.00118117
R2475 VDD.n619 VDD.n618 0.00118117
R2476 VDD.n617 VDD.n276 0.00118117
R2477 VDD.n616 VDD.n615 0.00118117
R2478 VDD.n614 VDD.n611 0.00118117
R2479 VDD.n610 VDD.n281 0.00118117
R2480 VDD.n609 VDD.n608 0.00118117
R2481 VDD.n605 VDD.n604 0.00118117
R2482 VDD.n603 VDD.n286 0.00118117
R2483 VDD.n602 VDD.n601 0.00118117
R2484 VDD.n600 VDD.n597 0.00118117
R2485 VDD.n596 VDD.n291 0.00118117
R2486 VDD.n595 VDD.n594 0.00118117
R2487 VDD.n591 VDD.n590 0.00118117
R2488 VDD.n589 VDD.n296 0.00118117
R2489 VDD.n588 VDD.n587 0.00118117
R2490 VDD.n586 VDD.n583 0.00118117
R2491 VDD.n582 VDD.n301 0.00118117
R2492 VDD.n581 VDD.n580 0.00118117
R2493 VDD.n577 VDD.n576 0.00118117
R2494 VDD.n575 VDD.n306 0.00118117
R2495 VDD.n574 VDD.n573 0.00118117
R2496 VDD.n572 VDD.n569 0.00118117
R2497 VDD.n568 VDD.n311 0.00118117
R2498 VDD.n567 VDD.n566 0.00118117
R2499 VDD.n563 VDD.n562 0.00118117
R2500 VDD.n561 VDD.n316 0.00118117
R2501 VDD.n560 VDD.n559 0.00118117
R2502 VDD.n556 VDD.n555 0.00118117
R2503 VDD.n553 VDD.n552 0.00118117
R2504 VDD.n551 VDD.n550 0.00118117
R2505 VDD.n547 VDD.n546 0.00118117
R2506 VDD.n545 VDD.n322 0.00118117
R2507 VDD.n544 VDD.n543 0.00118117
R2508 VDD.n542 VDD.n539 0.00118117
R2509 VDD.n538 VDD.n327 0.00118117
R2510 VDD.n537 VDD.n536 0.00118117
R2511 VDD.n533 VDD.n532 0.00118117
R2512 VDD.n531 VDD.n332 0.00118117
R2513 VDD.n530 VDD.n529 0.00118117
R2514 VDD.n528 VDD.n525 0.00118117
R2515 VDD.n524 VDD.n337 0.00118117
R2516 VDD.n523 VDD.n522 0.00118117
R2517 VDD.n519 VDD.n518 0.00118117
R2518 VDD.n517 VDD.n342 0.00118117
R2519 VDD.n516 VDD.n515 0.00118117
R2520 VDD.n514 VDD.n512 0.00118117
R2521 VDD.n511 VDD.n510 0.00118117
R2522 VDD.n509 VDD.n506 0.00118117
R2523 VDD.n505 VDD.n348 0.00118117
R2524 VDD.n504 VDD.n503 0.00118117
R2525 VDD.n500 VDD.n499 0.00118117
R2526 VDD.n498 VDD.n353 0.00118117
R2527 VDD.n497 VDD.n496 0.00118117
R2528 VDD.n495 VDD.n492 0.00118117
R2529 VDD.n491 VDD.n358 0.00118117
R2530 VDD.n490 VDD.n489 0.00118117
R2531 VDD.n486 VDD.n485 0.00118117
R2532 VDD.n484 VDD.n363 0.00118117
R2533 VDD.n483 VDD.n482 0.00118117
R2534 VDD.n481 VDD.n478 0.00118117
R2535 VDD.n477 VDD.n368 0.00118117
R2536 VDD.n476 VDD.n475 0.00118117
R2537 VDD.n473 VDD.n472 0.00118117
R2538 VDD.n471 VDD.n470 0.00118117
R2539 VDD.n467 VDD.n466 0.00118117
R2540 VDD.n465 VDD.n374 0.00118117
R2541 VDD.n464 VDD.n463 0.00118117
R2542 VDD.n462 VDD.n459 0.00118117
R2543 VDD.n458 VDD.n379 0.00118117
R2544 VDD.n457 VDD.n456 0.00118117
R2545 VDD.n453 VDD.n452 0.00118117
R2546 VDD.n451 VDD.n384 0.00118117
R2547 VDD.n450 VDD.n449 0.00118117
R2548 VDD.n448 VDD.n445 0.00118117
R2549 VDD.n444 VDD.n443 0.00118117
R2550 VDD.n442 VDD.n440 0.00118117
R2551 VDD.n439 VDD.n438 0.00118117
R2552 VDD.n437 VDD.n434 0.00118117
R2553 VDD.n433 VDD.n393 0.00118117
R2554 VDD.n432 VDD.n431 0.00118117
R2555 VDD.n428 VDD.n427 0.00118117
R2556 VDD.n426 VDD.n399 0.00118117
R2557 VDD.n425 VDD.n424 0.00118117
R2558 VDD.n421 VDD.n420 0.00118117
R2559 VDD.n418 VDD.n417 0.00118117
R2560 VDD.n416 VDD.n403 0.00118117
R2561 VDD.n415 VDD.n414 0.00118117
R2562 VDD.n413 VDD.n412 0.00118117
R2563 VDD.n411 VDD.n409 0.00118117
R2564 VDD.n2 VDD.n1 0.00118117
R2565 VDD.n6 VDD.n5 0.00118117
R2566 VDD.n1012 VDD.n1011 0.00118117
R2567 VDD.n1010 VDD.n1007 0.00118117
R2568 VDD.n1006 VDD.n11 0.00118117
R2569 VDD.n1005 VDD.n1004 0.00118117
R2570 VDD.n1001 VDD.n1000 0.00118117
R2571 VDD.n999 VDD.n16 0.00118117
R2572 VDD.n998 VDD.n997 0.00118117
R2573 VDD.n996 VDD.n993 0.00118117
R2574 VDD.n992 VDD.n21 0.00118117
R2575 VDD.n991 VDD.n990 0.00118117
R2576 VDD.n987 VDD.n986 0.00118117
R2577 VDD.n985 VDD.n26 0.00118117
R2578 VDD.n984 VDD.n983 0.00118117
R2579 VDD.n982 VDD.n979 0.00118117
R2580 VDD.n978 VDD.n31 0.00118117
R2581 VDD.n977 VDD.n976 0.00118117
R2582 VDD.n973 VDD.n972 0.00118117
R2583 VDD.n971 VDD.n36 0.00118117
R2584 VDD.n970 VDD.n969 0.00118117
R2585 VDD.n968 VDD.n965 0.00118117
R2586 VDD.n964 VDD.n41 0.00118117
R2587 VDD.n963 VDD.n962 0.00118117
R2588 VDD.n959 VDD.n958 0.00118117
R2589 VDD.n957 VDD.n46 0.00118117
R2590 VDD.n956 VDD.n955 0.00118117
R2591 VDD.n954 VDD.n951 0.00118117
R2592 VDD.n950 VDD.n51 0.00118117
R2593 VDD.n949 VDD.n948 0.00118117
R2594 VDD.n945 VDD.n944 0.00118117
R2595 VDD.n943 VDD.n56 0.00118117
R2596 VDD.n942 VDD.n941 0.00118117
R2597 VDD.n940 VDD.n937 0.00118117
R2598 VDD.n936 VDD.n61 0.00118117
R2599 VDD.n935 VDD.n934 0.00118117
R2600 VDD.n931 VDD.n930 0.00118117
R2601 VDD.n929 VDD.n66 0.00118117
R2602 VDD.n928 VDD.n927 0.00118117
R2603 VDD.n926 VDD.n923 0.00118117
R2604 VDD.n922 VDD.n71 0.00118117
R2605 VDD.n921 VDD.n920 0.00118117
R2606 VDD.n917 VDD.n916 0.00118117
R2607 VDD.n915 VDD.n76 0.00118117
R2608 VDD.n914 VDD.n913 0.00118117
R2609 VDD.n912 VDD.n909 0.00118117
R2610 VDD.n908 VDD.n81 0.00118117
R2611 VDD.n907 VDD.n906 0.00118117
R2612 VDD.n903 VDD.n902 0.00118117
R2613 VDD.n901 VDD.n86 0.00118117
R2614 VDD.n900 VDD.n899 0.00118117
R2615 VDD.n898 VDD.n895 0.00118117
R2616 VDD.n894 VDD.n91 0.00118117
R2617 VDD.n893 VDD.n892 0.00118117
R2618 VDD.n889 VDD.n888 0.00118117
R2619 VDD.n887 VDD.n96 0.00118117
R2620 VDD.n886 VDD.n885 0.00118117
R2621 VDD.n884 VDD.n881 0.00118117
R2622 VDD.n880 VDD.n101 0.00118117
R2623 VDD.n879 VDD.n878 0.00118117
R2624 VDD.n875 VDD.n874 0.00118117
R2625 VDD.n873 VDD.n106 0.00118117
R2626 VDD.n872 VDD.n871 0.00118117
R2627 VDD.n870 VDD.n867 0.00118117
R2628 VDD.n866 VDD.n865 0.00118117
R2629 VDD.n864 VDD.n862 0.00118117
R2630 VDD.n861 VDD.n860 0.00118117
R2631 VDD.n859 VDD.n856 0.00118117
R2632 VDD.n855 VDD.n114 0.00118117
R2633 VDD.n854 VDD.n853 0.00118117
R2634 VDD.n850 VDD.n849 0.00118117
R2635 VDD.n848 VDD.n119 0.00118117
R2636 VDD.n847 VDD.n846 0.00118117
R2637 VDD.n845 VDD.n842 0.00118117
R2638 VDD.n841 VDD.n124 0.00118117
R2639 VDD.n840 VDD.n839 0.00118117
R2640 VDD.n836 VDD.n835 0.00118117
R2641 VDD.n834 VDD.n129 0.00118117
R2642 VDD.n833 VDD.n832 0.00118117
R2643 VDD.n831 VDD.n828 0.00118117
R2644 VDD.n827 VDD.n134 0.00118117
R2645 VDD.n826 VDD.n825 0.00118117
R2646 VDD.n822 VDD.n821 0.00118117
R2647 VDD.n820 VDD.n139 0.00118117
R2648 VDD.n819 VDD.n818 0.00118117
R2649 VDD.n817 VDD.n814 0.00118117
R2650 VDD.n813 VDD.n144 0.00118117
R2651 VDD.n812 VDD.n811 0.00118117
R2652 VDD.n808 VDD.n807 0.00118117
R2653 VDD.n806 VDD.n149 0.00118117
R2654 VDD.n805 VDD.n804 0.00118117
R2655 VDD.n803 VDD.n800 0.00118117
R2656 VDD.n799 VDD.n154 0.00118117
R2657 VDD.n798 VDD.n797 0.00118117
R2658 VDD.n794 VDD.n793 0.00118117
R2659 VDD.n792 VDD.n159 0.00118117
R2660 VDD.n791 VDD.n790 0.00118117
R2661 VDD.n789 VDD.n786 0.00118117
R2662 VDD.n785 VDD.n164 0.00118117
R2663 VDD.n784 VDD.n783 0.00118117
R2664 VDD.n780 VDD.n779 0.00118117
R2665 VDD.n778 VDD.n169 0.00118117
R2666 VDD.n777 VDD.n776 0.00118117
R2667 VDD.n775 VDD.n772 0.00118117
R2668 VDD.n771 VDD.n174 0.00118117
R2669 VDD.n770 VDD.n769 0.00118117
R2670 VDD.n766 VDD.n765 0.00118117
R2671 VDD.n764 VDD.n179 0.00118117
R2672 VDD.n763 VDD.n762 0.00118117
R2673 VDD.n761 VDD.n758 0.00118117
R2674 VDD.n757 VDD.n184 0.00118117
R2675 VDD.n756 VDD.n755 0.00118117
R2676 VDD.n752 VDD.n751 0.00118117
R2677 VDD.n750 VDD.n189 0.00118117
R2678 VDD.n749 VDD.n748 0.00118117
R2679 VDD.n747 VDD.n744 0.00118117
R2680 VDD.n743 VDD.n194 0.00118117
R2681 VDD.n742 VDD.n741 0.00118117
R2682 VDD.n738 VDD.n737 0.00118117
R2683 VDD.n736 VDD.n199 0.00118117
R2684 VDD.n735 VDD.n734 0.00118117
R2685 VDD.n733 VDD.n730 0.00118117
R2686 VDD.n729 VDD.n204 0.00118117
R2687 VDD.n728 VDD.n727 0.00118117
R2688 VDD.n724 VDD.n723 0.00118117
R2689 VDD.n722 VDD.n209 0.00118117
R2690 VDD.n721 VDD.n720 0.00118117
R2691 VDD.n719 VDD.n716 0.00118117
R2692 VDD.n715 VDD.n214 0.00118117
R2693 VDD.n714 VDD.n713 0.00118117
R2694 db<3>.n1 db<3>.n0 88.1376
R2695 db<3>.n2 db<3>.n1 88.1376
R2696 db<3>.n3 db<3>.n2 88.1376
R2697 db<3>.n4 db<3>.n3 88.1376
R2698 db<3>.n5 db<3>.n4 88.1376
R2699 db<3>.n6 db<3>.n5 88.1376
R2700 db<3>.n7 db<3>.n6 88.1376
R2701 db<3>.n0 db<3>.t0 69.5462
R2702 db<3>.n1 db<3>.t10 69.5462
R2703 db<3>.n2 db<3>.t14 69.5462
R2704 db<3>.n3 db<3>.t7 69.5462
R2705 db<3>.n4 db<3>.t12 69.5462
R2706 db<3>.n5 db<3>.t9 69.5462
R2707 db<3>.n6 db<3>.t3 69.5462
R2708 db<3>.n7 db<3>.t2 69.5462
R2709 db<3>.n0 db<3>.t11 59.9062
R2710 db<3>.n1 db<3>.t5 59.9062
R2711 db<3>.n2 db<3>.t8 59.9062
R2712 db<3>.n3 db<3>.t1 59.9062
R2713 db<3>.n4 db<3>.t6 59.9062
R2714 db<3>.n5 db<3>.t4 59.9062
R2715 db<3>.n6 db<3>.t15 59.9062
R2716 db<3>.n7 db<3>.t13 59.9062
R2717 db<3> db<3>.n7 24.1005
R2718 hgu_cdac_8bit_array_2.drv<7:0>.n30 hgu_cdac_8bit_array_2.drv<7:0>.t0 41.4291
R2719 hgu_cdac_8bit_array_2.drv<7:0>.n30 hgu_cdac_8bit_array_2.drv<7:0>.t2 41.4291
R2720 hgu_cdac_8bit_array_2.drv<7:0>.n10 hgu_cdac_8bit_array_2.drv<7:0>.t7 41.4291
R2721 hgu_cdac_8bit_array_2.drv<7:0>.n10 hgu_cdac_8bit_array_2.drv<7:0>.t3 41.4291
R2722 hgu_cdac_8bit_array_2.drv<7:0>.n13 hgu_cdac_8bit_array_2.drv<7:0>.t6 41.4291
R2723 hgu_cdac_8bit_array_2.drv<7:0>.n13 hgu_cdac_8bit_array_2.drv<7:0>.t1 41.4291
R2724 hgu_cdac_8bit_array_2.drv<7:0>.n33 hgu_cdac_8bit_array_2.drv<7:0>.t4 41.4291
R2725 hgu_cdac_8bit_array_2.drv<7:0>.n33 hgu_cdac_8bit_array_2.drv<7:0>.t5 41.4291
R2726 hgu_cdac_8bit_array_2.drv<7:0>.n29 hgu_cdac_8bit_array_2.drv<7:0>.t9 34.0065
R2727 hgu_cdac_8bit_array_2.drv<7:0>.n29 hgu_cdac_8bit_array_2.drv<7:0>.t11 34.0065
R2728 hgu_cdac_8bit_array_2.drv<7:0>.n9 hgu_cdac_8bit_array_2.drv<7:0>.t8 34.0065
R2729 hgu_cdac_8bit_array_2.drv<7:0>.n9 hgu_cdac_8bit_array_2.drv<7:0>.t12 34.0065
R2730 hgu_cdac_8bit_array_2.drv<7:0>.n12 hgu_cdac_8bit_array_2.drv<7:0>.t15 34.0065
R2731 hgu_cdac_8bit_array_2.drv<7:0>.n12 hgu_cdac_8bit_array_2.drv<7:0>.t10 34.0065
R2732 hgu_cdac_8bit_array_2.drv<7:0>.n32 hgu_cdac_8bit_array_2.drv<7:0>.t13 34.0065
R2733 hgu_cdac_8bit_array_2.drv<7:0>.n32 hgu_cdac_8bit_array_2.drv<7:0>.t14 34.0065
R2734 hgu_cdac_8bit_array_2.drv<7:0>.n38 hgu_cdac_8bit_array_2.drv<7:0>.n34 12.4472
R2735 hgu_cdac_8bit_array_2.drv<7:0>.n15 hgu_cdac_8bit_array_2.drv<7:0>.n14 11.1146
R2736 hgu_cdac_8bit_array_2.drv<7:0>.n21 hgu_cdac_8bit_array_2.drv<7:0>.n15 1.37688
R2737 hgu_cdac_8bit_array_2.drv<7:0>.n14 hgu_cdac_8bit_array_2.drv<7:0>.n11 0.957397
R2738 hgu_cdac_8bit_array_2.drv<7:0>.n34 hgu_cdac_8bit_array_2.drv<7:0>.n31 0.957397
R2739 hgu_cdac_8bit_array_2.drv<7:0>.n31 hgu_cdac_8bit_array_2.drv<7:0>.n29 0.561881
R2740 hgu_cdac_8bit_array_2.drv<7:0>.n11 hgu_cdac_8bit_array_2.drv<7:0>.n9 0.561881
R2741 hgu_cdac_8bit_array_2.drv<7:0>.n14 hgu_cdac_8bit_array_2.drv<7:0>.n12 0.561881
R2742 hgu_cdac_8bit_array_2.drv<7:0>.n34 hgu_cdac_8bit_array_2.drv<7:0>.n32 0.561881
R2743 hgu_cdac_8bit_array_2.drv<7:0>.n0 hgu_cdac_8bit_array_2.drv<7:0> 0.321667
R2744 hgu_cdac_8bit_array_2.drv<7:0>.n6 hgu_cdac_8bit_array_2.drv<7:0> 0.321667
R2745 hgu_cdac_8bit_array_2.drv<7:0>.n1 hgu_cdac_8bit_array_2.drv<7:0> 0.321667
R2746 hgu_cdac_8bit_array_2.drv<7:0>.n39 hgu_cdac_8bit_array_2.drv<7:0> 0.313448
R2747 hgu_cdac_8bit_array_2.drv<7:0>.n31 hgu_cdac_8bit_array_2.drv<7:0>.n30 0.297179
R2748 hgu_cdac_8bit_array_2.drv<7:0>.n11 hgu_cdac_8bit_array_2.drv<7:0>.n10 0.297179
R2749 hgu_cdac_8bit_array_2.drv<7:0>.n14 hgu_cdac_8bit_array_2.drv<7:0>.n13 0.297179
R2750 hgu_cdac_8bit_array_2.drv<7:0>.n34 hgu_cdac_8bit_array_2.drv<7:0>.n33 0.297179
R2751 hgu_cdac_8bit_array_2.drv<7:0>.n2 hgu_cdac_8bit_array_2.drv<7:0> 0.2966
R2752 hgu_cdac_8bit_array_2.drv<7:0>.n5 hgu_cdac_8bit_array_2.drv<7:0> 0.2966
R2753 hgu_cdac_8bit_array_2.drv<7:0>.n8 hgu_cdac_8bit_array_2.drv<7:0> 0.2966
R2754 hgu_cdac_8bit_array_2.drv<7:0>.n1 hgu_cdac_8bit_array_2.drv<7:0>.n22 0.241293
R2755 hgu_cdac_8bit_array_2.drv<7:0>.n4 hgu_cdac_8bit_array_2.drv<7:0> 0.219833
R2756 hgu_cdac_8bit_array_2.drv<7:0>.n25 hgu_cdac_8bit_array_2.drv<7:0>.n21 0.182836
R2757 hgu_cdac_8bit_array_2.drv<7:0>.n41 hgu_cdac_8bit_array_2.drv<7:0>.n38 0.182836
R2758 hgu_cdac_8bit_array_2.drv<7:0>.n21 hgu_cdac_8bit_array_2.drv<7:0>.n20 0.149114
R2759 hgu_cdac_8bit_array_2.drv<7:0>.n38 hgu_cdac_8bit_array_2.drv<7:0>.n37 0.149114
R2760 hgu_cdac_8bit_array_2.drv<7:0>.n40 hgu_cdac_8bit_array_2.drv<7:0>.n0 0.0972647
R2761 hgu_cdac_8bit_array_2.drv<7:0>.n25 hgu_cdac_8bit_array_2.drv<7:0>.n24 0.0716912
R2762 hgu_cdac_8bit_array_2.drv<7:0>.n26 hgu_cdac_8bit_array_2.drv<7:0>.n25 0.0716912
R2763 hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_8bit_array_2.drv<7:0>.n28 0.0716912
R2764 hgu_cdac_8bit_array_2.drv<7:0>.n42 hgu_cdac_8bit_array_2.drv<7:0>.n41 0.0716912
R2765 hgu_cdac_8bit_array_2.drv<7:0>.n41 hgu_cdac_8bit_array_2.drv<7:0>.n40 0.0716912
R2766 hgu_cdac_8bit_array_2.drv<7:0>.n20 hgu_cdac_8bit_array_2.drv<7:0>.n19 0.0716912
R2767 hgu_cdac_8bit_array_2.drv<7:0>.n37 hgu_cdac_8bit_array_2.drv<7:0>.n36 0.0716912
R2768 hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_8bit_array_2.drv<7:0>.n44 0.0716912
R2769 hgu_cdac_8bit_array_2.drv<7:0>.n2 hgu_cdac_8bit_array_2.drv<7:0>.n1 0.0696176
R2770 hgu_cdac_8bit_array_2.drv<7:0>.n0 hgu_cdac_8bit_array_2.drv<7:0>.n39 0.0664894
R2771 hgu_cdac_8bit_array_2.drv<7:0>.n24 hgu_cdac_8bit_array_2.drv<7:0>.n23 0.0557941
R2772 hgu_cdac_8bit_array_2.drv<7:0>.n3 hgu_cdac_8bit_array_2.drv<7:0>.n26 0.0557941
R2773 hgu_cdac_8bit_array_2.drv<7:0>.n5 hgu_cdac_8bit_array_2.drv<7:0>.n4 0.0557941
R2774 hgu_cdac_8bit_array_2.drv<7:0>.n28 hgu_cdac_8bit_array_2.drv<7:0>.n27 0.0557941
R2775 hgu_cdac_8bit_array_2.drv<7:0>.n44 hgu_cdac_8bit_array_2.drv<7:0>.n43 0.0557941
R2776 hgu_cdac_8bit_array_2.drv<7:0>.n6 hgu_cdac_8bit_array_2.drv<7:0>.n8 0.0557941
R2777 hgu_cdac_8bit_array_2.drv<7:0>.n7 hgu_cdac_8bit_array_2.drv<7:0>.n42 0.0557941
R2778 hgu_cdac_8bit_array_2.drv<7:0>.n17 hgu_cdac_8bit_array_2.drv<7:0>.n16 0.0557941
R2779 hgu_cdac_8bit_array_2.drv<7:0>.n18 hgu_cdac_8bit_array_2.drv<7:0>.n17 0.0557941
R2780 hgu_cdac_8bit_array_2.drv<7:0>.n19 hgu_cdac_8bit_array_2.drv<7:0>.n18 0.0557941
R2781 hgu_cdac_8bit_array_2.drv<7:0>.n36 hgu_cdac_8bit_array_2.drv<7:0>.n35 0.0557941
R2782 hgu_cdac_8bit_array_2.drv<7:0>.n8 hgu_cdac_8bit_array_2.drv<7:0>.n7 0.0557941
R2783 hgu_cdac_8bit_array_2.drv<7:0>.n43 hgu_cdac_8bit_array_2.drv<7:0>.n6 0.0557941
R2784 hgu_cdac_8bit_array_2.drv<7:0>.n27 hgu_cdac_8bit_array_2.drv<7:0>.n5 0.0557941
R2785 hgu_cdac_8bit_array_2.drv<7:0>.n4 hgu_cdac_8bit_array_2.drv<7:0>.n3 0.0557941
R2786 hgu_cdac_8bit_array_2.drv<7:0>.n23 hgu_cdac_8bit_array_2.drv<7:0>.n2 0.0557941
R2787 db<5>.n1 db<5>.n0 88.1376
R2788 db<5>.n2 db<5>.n1 88.1376
R2789 db<5>.n3 db<5>.n2 88.1376
R2790 db<5>.n4 db<5>.n3 88.1376
R2791 db<5>.n5 db<5>.n4 88.1376
R2792 db<5>.n6 db<5>.n5 88.1376
R2793 db<5>.n7 db<5>.n6 88.1376
R2794 db<5>.n8 db<5>.n7 88.1376
R2795 db<5>.n9 db<5>.n8 88.1376
R2796 db<5>.n10 db<5>.n9 88.1376
R2797 db<5>.n11 db<5>.n10 88.1376
R2798 db<5>.n12 db<5>.n11 88.1376
R2799 db<5>.n13 db<5>.n12 88.1376
R2800 db<5>.n14 db<5>.n13 88.1376
R2801 db<5>.n15 db<5>.n14 88.1376
R2802 db<5>.n16 db<5>.n15 88.1376
R2803 db<5>.n17 db<5>.n16 88.1376
R2804 db<5>.n18 db<5>.n17 88.1376
R2805 db<5>.n19 db<5>.n18 88.1376
R2806 db<5>.n20 db<5>.n19 88.1376
R2807 db<5>.n21 db<5>.n20 88.1376
R2808 db<5>.n22 db<5>.n21 88.1376
R2809 db<5>.n23 db<5>.n22 88.1376
R2810 db<5>.n24 db<5>.n23 88.1376
R2811 db<5>.n25 db<5>.n24 88.1376
R2812 db<5>.n26 db<5>.n25 88.1376
R2813 db<5>.n27 db<5>.n26 88.1376
R2814 db<5>.n28 db<5>.n27 88.1376
R2815 db<5>.n29 db<5>.n28 88.1376
R2816 db<5>.n30 db<5>.n29 88.1376
R2817 db<5>.n31 db<5>.n30 88.1376
R2818 db<5>.n0 db<5>.t12 69.5462
R2819 db<5>.n1 db<5>.t54 69.5462
R2820 db<5>.n2 db<5>.t63 69.5462
R2821 db<5>.n3 db<5>.t36 69.5462
R2822 db<5>.n4 db<5>.t13 69.5462
R2823 db<5>.n5 db<5>.t5 69.5462
R2824 db<5>.n6 db<5>.t46 69.5462
R2825 db<5>.n7 db<5>.t17 69.5462
R2826 db<5>.n8 db<5>.t58 69.5462
R2827 db<5>.n9 db<5>.t50 69.5462
R2828 db<5>.n10 db<5>.t26 69.5462
R2829 db<5>.n11 db<5>.t3 69.5462
R2830 db<5>.n12 db<5>.t59 69.5462
R2831 db<5>.n13 db<5>.t52 69.5462
R2832 db<5>.n14 db<5>.t28 69.5462
R2833 db<5>.n15 db<5>.t47 69.5462
R2834 db<5>.n16 db<5>.t38 69.5462
R2835 db<5>.n17 db<5>.t32 69.5462
R2836 db<5>.n18 db<5>.t7 69.5462
R2837 db<5>.n19 db<5>.t48 69.5462
R2838 db<5>.n20 db<5>.t41 69.5462
R2839 db<5>.n21 db<5>.t16 69.5462
R2840 db<5>.n22 db<5>.t9 69.5462
R2841 db<5>.n23 db<5>.t43 69.5462
R2842 db<5>.n24 db<5>.t20 69.5462
R2843 db<5>.n25 db<5>.t62 69.5462
R2844 db<5>.n26 db<5>.t35 69.5462
R2845 db<5>.n27 db<5>.t45 69.5462
R2846 db<5>.n28 db<5>.t21 69.5462
R2847 db<5>.n29 db<5>.t0 69.5462
R2848 db<5>.n30 db<5>.t33 69.5462
R2849 db<5>.n31 db<5>.t8 69.5462
R2850 db<5>.n0 db<5>.t56 59.9062
R2851 db<5>.n1 db<5>.t31 59.9062
R2852 db<5>.n2 db<5>.t40 59.9062
R2853 db<5>.n3 db<5>.t15 59.9062
R2854 db<5>.n4 db<5>.t57 59.9062
R2855 db<5>.n5 db<5>.t49 59.9062
R2856 db<5>.n6 db<5>.t24 59.9062
R2857 db<5>.n7 db<5>.t61 59.9062
R2858 db<5>.n8 db<5>.t34 59.9062
R2859 db<5>.n9 db<5>.t29 59.9062
R2860 db<5>.n10 db<5>.t4 59.9062
R2861 db<5>.n11 db<5>.t44 59.9062
R2862 db<5>.n12 db<5>.t37 59.9062
R2863 db<5>.n13 db<5>.t30 59.9062
R2864 db<5>.n14 db<5>.t6 59.9062
R2865 db<5>.n15 db<5>.t25 59.9062
R2866 db<5>.n16 db<5>.t18 59.9062
R2867 db<5>.n17 db<5>.t10 59.9062
R2868 db<5>.n18 db<5>.t51 59.9062
R2869 db<5>.n19 db<5>.t27 59.9062
R2870 db<5>.n20 db<5>.t19 59.9062
R2871 db<5>.n21 db<5>.t60 59.9062
R2872 db<5>.n22 db<5>.t55 59.9062
R2873 db<5>.n23 db<5>.t22 59.9062
R2874 db<5>.n24 db<5>.t1 59.9062
R2875 db<5>.n25 db<5>.t39 59.9062
R2876 db<5>.n26 db<5>.t14 59.9062
R2877 db<5>.n27 db<5>.t23 59.9062
R2878 db<5>.n28 db<5>.t2 59.9062
R2879 db<5>.n29 db<5>.t42 59.9062
R2880 db<5>.n30 db<5>.t11 59.9062
R2881 db<5>.n31 db<5>.t53 59.9062
R2882 db<5> db<5>.n31 24.1005
R2883 hgu_cdac_8bit_array_2.drv<31:0>.n129 hgu_cdac_8bit_array_2.drv<31:0>.t51 41.4291
R2884 hgu_cdac_8bit_array_2.drv<31:0>.n129 hgu_cdac_8bit_array_2.drv<31:0>.t47 41.4291
R2885 hgu_cdac_8bit_array_2.drv<31:0>.n85 hgu_cdac_8bit_array_2.drv<31:0>.t63 41.4291
R2886 hgu_cdac_8bit_array_2.drv<31:0>.n85 hgu_cdac_8bit_array_2.drv<31:0>.t57 41.4291
R2887 hgu_cdac_8bit_array_2.drv<31:0>.n87 hgu_cdac_8bit_array_2.drv<31:0>.t50 41.4291
R2888 hgu_cdac_8bit_array_2.drv<31:0>.n87 hgu_cdac_8bit_array_2.drv<31:0>.t60 41.4291
R2889 hgu_cdac_8bit_array_2.drv<31:0>.n89 hgu_cdac_8bit_array_2.drv<31:0>.t4 41.4291
R2890 hgu_cdac_8bit_array_2.drv<31:0>.n89 hgu_cdac_8bit_array_2.drv<31:0>.t11 41.4291
R2891 hgu_cdac_8bit_array_2.drv<31:0>.n91 hgu_cdac_8bit_array_2.drv<31:0>.t46 41.4291
R2892 hgu_cdac_8bit_array_2.drv<31:0>.n91 hgu_cdac_8bit_array_2.drv<31:0>.t1 41.4291
R2893 hgu_cdac_8bit_array_2.drv<31:0>.n93 hgu_cdac_8bit_array_2.drv<31:0>.t9 41.4291
R2894 hgu_cdac_8bit_array_2.drv<31:0>.n93 hgu_cdac_8bit_array_2.drv<31:0>.t61 41.4291
R2895 hgu_cdac_8bit_array_2.drv<31:0>.n95 hgu_cdac_8bit_array_2.drv<31:0>.t45 41.4291
R2896 hgu_cdac_8bit_array_2.drv<31:0>.n95 hgu_cdac_8bit_array_2.drv<31:0>.t48 41.4291
R2897 hgu_cdac_8bit_array_2.drv<31:0>.n97 hgu_cdac_8bit_array_2.drv<31:0>.t8 41.4291
R2898 hgu_cdac_8bit_array_2.drv<31:0>.n97 hgu_cdac_8bit_array_2.drv<31:0>.t3 41.4291
R2899 hgu_cdac_8bit_array_2.drv<31:0>.n99 hgu_cdac_8bit_array_2.drv<31:0>.t56 41.4291
R2900 hgu_cdac_8bit_array_2.drv<31:0>.n99 hgu_cdac_8bit_array_2.drv<31:0>.t7 41.4291
R2901 hgu_cdac_8bit_array_2.drv<31:0>.n101 hgu_cdac_8bit_array_2.drv<31:0>.t59 41.4291
R2902 hgu_cdac_8bit_array_2.drv<31:0>.n101 hgu_cdac_8bit_array_2.drv<31:0>.t2 41.4291
R2903 hgu_cdac_8bit_array_2.drv<31:0>.n103 hgu_cdac_8bit_array_2.drv<31:0>.t55 41.4291
R2904 hgu_cdac_8bit_array_2.drv<31:0>.n103 hgu_cdac_8bit_array_2.drv<31:0>.t49 41.4291
R2905 hgu_cdac_8bit_array_2.drv<31:0>.n105 hgu_cdac_8bit_array_2.drv<31:0>.t52 41.4291
R2906 hgu_cdac_8bit_array_2.drv<31:0>.n105 hgu_cdac_8bit_array_2.drv<31:0>.t54 41.4291
R2907 hgu_cdac_8bit_array_2.drv<31:0>.n107 hgu_cdac_8bit_array_2.drv<31:0>.t0 41.4291
R2908 hgu_cdac_8bit_array_2.drv<31:0>.n107 hgu_cdac_8bit_array_2.drv<31:0>.t44 41.4291
R2909 hgu_cdac_8bit_array_2.drv<31:0>.n109 hgu_cdac_8bit_array_2.drv<31:0>.t58 41.4291
R2910 hgu_cdac_8bit_array_2.drv<31:0>.n109 hgu_cdac_8bit_array_2.drv<31:0>.t5 41.4291
R2911 hgu_cdac_8bit_array_2.drv<31:0>.n111 hgu_cdac_8bit_array_2.drv<31:0>.t6 41.4291
R2912 hgu_cdac_8bit_array_2.drv<31:0>.n111 hgu_cdac_8bit_array_2.drv<31:0>.t53 41.4291
R2913 hgu_cdac_8bit_array_2.drv<31:0>.n114 hgu_cdac_8bit_array_2.drv<31:0>.t10 41.4291
R2914 hgu_cdac_8bit_array_2.drv<31:0>.n114 hgu_cdac_8bit_array_2.drv<31:0>.t62 41.4291
R2915 hgu_cdac_8bit_array_2.drv<31:0>.n83 hgu_cdac_8bit_array_2.drv<31:0>.t37 34.0065
R2916 hgu_cdac_8bit_array_2.drv<31:0>.n83 hgu_cdac_8bit_array_2.drv<31:0>.t16 34.0065
R2917 hgu_cdac_8bit_array_2.drv<31:0>.n84 hgu_cdac_8bit_array_2.drv<31:0>.t12 34.0065
R2918 hgu_cdac_8bit_array_2.drv<31:0>.n84 hgu_cdac_8bit_array_2.drv<31:0>.t26 34.0065
R2919 hgu_cdac_8bit_array_2.drv<31:0>.n86 hgu_cdac_8bit_array_2.drv<31:0>.t36 34.0065
R2920 hgu_cdac_8bit_array_2.drv<31:0>.n86 hgu_cdac_8bit_array_2.drv<31:0>.t41 34.0065
R2921 hgu_cdac_8bit_array_2.drv<31:0>.n88 hgu_cdac_8bit_array_2.drv<31:0>.t21 34.0065
R2922 hgu_cdac_8bit_array_2.drv<31:0>.n88 hgu_cdac_8bit_array_2.drv<31:0>.t34 34.0065
R2923 hgu_cdac_8bit_array_2.drv<31:0>.n90 hgu_cdac_8bit_array_2.drv<31:0>.t15 34.0065
R2924 hgu_cdac_8bit_array_2.drv<31:0>.n90 hgu_cdac_8bit_array_2.drv<31:0>.t18 34.0065
R2925 hgu_cdac_8bit_array_2.drv<31:0>.n92 hgu_cdac_8bit_array_2.drv<31:0>.t31 34.0065
R2926 hgu_cdac_8bit_array_2.drv<31:0>.n92 hgu_cdac_8bit_array_2.drv<31:0>.t42 34.0065
R2927 hgu_cdac_8bit_array_2.drv<31:0>.n94 hgu_cdac_8bit_array_2.drv<31:0>.t14 34.0065
R2928 hgu_cdac_8bit_array_2.drv<31:0>.n94 hgu_cdac_8bit_array_2.drv<31:0>.t17 34.0065
R2929 hgu_cdac_8bit_array_2.drv<31:0>.n96 hgu_cdac_8bit_array_2.drv<31:0>.t30 34.0065
R2930 hgu_cdac_8bit_array_2.drv<31:0>.n96 hgu_cdac_8bit_array_2.drv<31:0>.t20 34.0065
R2931 hgu_cdac_8bit_array_2.drv<31:0>.n98 hgu_cdac_8bit_array_2.drv<31:0>.t25 34.0065
R2932 hgu_cdac_8bit_array_2.drv<31:0>.n98 hgu_cdac_8bit_array_2.drv<31:0>.t29 34.0065
R2933 hgu_cdac_8bit_array_2.drv<31:0>.n100 hgu_cdac_8bit_array_2.drv<31:0>.t40 34.0065
R2934 hgu_cdac_8bit_array_2.drv<31:0>.n100 hgu_cdac_8bit_array_2.drv<31:0>.t19 34.0065
R2935 hgu_cdac_8bit_array_2.drv<31:0>.n102 hgu_cdac_8bit_array_2.drv<31:0>.t24 34.0065
R2936 hgu_cdac_8bit_array_2.drv<31:0>.n102 hgu_cdac_8bit_array_2.drv<31:0>.t35 34.0065
R2937 hgu_cdac_8bit_array_2.drv<31:0>.n104 hgu_cdac_8bit_array_2.drv<31:0>.t38 34.0065
R2938 hgu_cdac_8bit_array_2.drv<31:0>.n104 hgu_cdac_8bit_array_2.drv<31:0>.t23 34.0065
R2939 hgu_cdac_8bit_array_2.drv<31:0>.n106 hgu_cdac_8bit_array_2.drv<31:0>.t33 34.0065
R2940 hgu_cdac_8bit_array_2.drv<31:0>.n106 hgu_cdac_8bit_array_2.drv<31:0>.t13 34.0065
R2941 hgu_cdac_8bit_array_2.drv<31:0>.n108 hgu_cdac_8bit_array_2.drv<31:0>.t27 34.0065
R2942 hgu_cdac_8bit_array_2.drv<31:0>.n108 hgu_cdac_8bit_array_2.drv<31:0>.t22 34.0065
R2943 hgu_cdac_8bit_array_2.drv<31:0>.n110 hgu_cdac_8bit_array_2.drv<31:0>.t28 34.0065
R2944 hgu_cdac_8bit_array_2.drv<31:0>.n110 hgu_cdac_8bit_array_2.drv<31:0>.t39 34.0065
R2945 hgu_cdac_8bit_array_2.drv<31:0>.n113 hgu_cdac_8bit_array_2.drv<31:0>.t32 34.0065
R2946 hgu_cdac_8bit_array_2.drv<31:0>.n113 hgu_cdac_8bit_array_2.drv<31:0>.t43 34.0065
R2947 hgu_cdac_8bit_array_2.drv<31:0>.n130 hgu_cdac_8bit_array_2.drv<31:0>.n0 12.6591
R2948 hgu_cdac_8bit_array_2.drv<31:0>.n0 hgu_cdac_8bit_array_2.drv<31:0>.n128 0.957397
R2949 hgu_cdac_8bit_array_2.drv<31:0>.n128 hgu_cdac_8bit_array_2.drv<31:0>.n127 0.957397
R2950 hgu_cdac_8bit_array_2.drv<31:0>.n127 hgu_cdac_8bit_array_2.drv<31:0>.n126 0.957397
R2951 hgu_cdac_8bit_array_2.drv<31:0>.n126 hgu_cdac_8bit_array_2.drv<31:0>.n125 0.957397
R2952 hgu_cdac_8bit_array_2.drv<31:0>.n125 hgu_cdac_8bit_array_2.drv<31:0>.n124 0.957397
R2953 hgu_cdac_8bit_array_2.drv<31:0>.n124 hgu_cdac_8bit_array_2.drv<31:0>.n123 0.957397
R2954 hgu_cdac_8bit_array_2.drv<31:0>.n123 hgu_cdac_8bit_array_2.drv<31:0>.n122 0.957397
R2955 hgu_cdac_8bit_array_2.drv<31:0>.n122 hgu_cdac_8bit_array_2.drv<31:0>.n121 0.957397
R2956 hgu_cdac_8bit_array_2.drv<31:0>.n121 hgu_cdac_8bit_array_2.drv<31:0>.n120 0.957397
R2957 hgu_cdac_8bit_array_2.drv<31:0>.n120 hgu_cdac_8bit_array_2.drv<31:0>.n119 0.957397
R2958 hgu_cdac_8bit_array_2.drv<31:0>.n119 hgu_cdac_8bit_array_2.drv<31:0>.n118 0.957397
R2959 hgu_cdac_8bit_array_2.drv<31:0>.n118 hgu_cdac_8bit_array_2.drv<31:0>.n117 0.957397
R2960 hgu_cdac_8bit_array_2.drv<31:0>.n117 hgu_cdac_8bit_array_2.drv<31:0>.n116 0.957397
R2961 hgu_cdac_8bit_array_2.drv<31:0>.n115 hgu_cdac_8bit_array_2.drv<31:0>.n112 0.957397
R2962 hgu_cdac_8bit_array_2.drv<31:0>.n116 hgu_cdac_8bit_array_2.drv<31:0>.n115 0.957397
R2963 hgu_cdac_8bit_array_2.drv<31:0>.n0 hgu_cdac_8bit_array_2.drv<31:0>.n83 0.561881
R2964 hgu_cdac_8bit_array_2.drv<31:0>.n128 hgu_cdac_8bit_array_2.drv<31:0>.n84 0.561881
R2965 hgu_cdac_8bit_array_2.drv<31:0>.n127 hgu_cdac_8bit_array_2.drv<31:0>.n86 0.561881
R2966 hgu_cdac_8bit_array_2.drv<31:0>.n126 hgu_cdac_8bit_array_2.drv<31:0>.n88 0.561881
R2967 hgu_cdac_8bit_array_2.drv<31:0>.n125 hgu_cdac_8bit_array_2.drv<31:0>.n90 0.561881
R2968 hgu_cdac_8bit_array_2.drv<31:0>.n124 hgu_cdac_8bit_array_2.drv<31:0>.n92 0.561881
R2969 hgu_cdac_8bit_array_2.drv<31:0>.n123 hgu_cdac_8bit_array_2.drv<31:0>.n94 0.561881
R2970 hgu_cdac_8bit_array_2.drv<31:0>.n122 hgu_cdac_8bit_array_2.drv<31:0>.n96 0.561881
R2971 hgu_cdac_8bit_array_2.drv<31:0>.n121 hgu_cdac_8bit_array_2.drv<31:0>.n98 0.561881
R2972 hgu_cdac_8bit_array_2.drv<31:0>.n120 hgu_cdac_8bit_array_2.drv<31:0>.n100 0.561881
R2973 hgu_cdac_8bit_array_2.drv<31:0>.n119 hgu_cdac_8bit_array_2.drv<31:0>.n102 0.561881
R2974 hgu_cdac_8bit_array_2.drv<31:0>.n118 hgu_cdac_8bit_array_2.drv<31:0>.n104 0.561881
R2975 hgu_cdac_8bit_array_2.drv<31:0>.n117 hgu_cdac_8bit_array_2.drv<31:0>.n106 0.561881
R2976 hgu_cdac_8bit_array_2.drv<31:0>.n116 hgu_cdac_8bit_array_2.drv<31:0>.n108 0.561881
R2977 hgu_cdac_8bit_array_2.drv<31:0>.n112 hgu_cdac_8bit_array_2.drv<31:0>.n110 0.561881
R2978 hgu_cdac_8bit_array_2.drv<31:0>.n115 hgu_cdac_8bit_array_2.drv<31:0>.n113 0.561881
R2979 hgu_cdac_8bit_array_2.drv<31:0>.n137 hgu_cdac_8bit_array_2.drv<31:0>.n82 0.330451
R2980 hgu_cdac_8bit_array_2.drv<31:0>.n146 hgu_cdac_8bit_array_2.drv<31:0>.n77 0.330451
R2981 hgu_cdac_8bit_array_2.drv<31:0>.n155 hgu_cdac_8bit_array_2.drv<31:0>.n70 0.330451
R2982 hgu_cdac_8bit_array_2.drv<31:0>.n164 hgu_cdac_8bit_array_2.drv<31:0>.n63 0.330451
R2983 hgu_cdac_8bit_array_2.drv<31:0>.n173 hgu_cdac_8bit_array_2.drv<31:0>.n56 0.330451
R2984 hgu_cdac_8bit_array_2.drv<31:0>.n182 hgu_cdac_8bit_array_2.drv<31:0>.n49 0.330451
R2985 hgu_cdac_8bit_array_2.drv<31:0>.n191 hgu_cdac_8bit_array_2.drv<31:0>.n42 0.330451
R2986 hgu_cdac_8bit_array_2.drv<31:0>.n200 hgu_cdac_8bit_array_2.drv<31:0>.n35 0.330451
R2987 hgu_cdac_8bit_array_2.drv<31:0>.n209 hgu_cdac_8bit_array_2.drv<31:0>.n28 0.330451
R2988 hgu_cdac_8bit_array_2.drv<31:0>.n218 hgu_cdac_8bit_array_2.drv<31:0>.n21 0.330451
R2989 hgu_cdac_8bit_array_2.drv<31:0>.n227 hgu_cdac_8bit_array_2.drv<31:0>.n14 0.330451
R2990 hgu_cdac_8bit_array_2.drv<31:0>.n236 hgu_cdac_8bit_array_2.drv<31:0>.n7 0.330451
R2991 hgu_cdac_8bit_array_2.drv<31:0>.n269 hgu_cdac_8bit_array_2.drv<31:0>.n252 0.330451
R2992 hgu_cdac_8bit_array_2.drv<31:0>.n260 hgu_cdac_8bit_array_2.drv<31:0>.n255 0.330451
R2993 hgu_cdac_8bit_array_2.drv<31:0>.n257 hgu_cdac_8bit_array_2.drv<31:0> 0.321667
R2994 hgu_cdac_8bit_array_2.drv<31:0>.n266 hgu_cdac_8bit_array_2.drv<31:0> 0.321667
R2995 hgu_cdac_8bit_array_2.drv<31:0>.n275 hgu_cdac_8bit_array_2.drv<31:0> 0.321667
R2996 hgu_cdac_8bit_array_2.drv<31:0>.n239 hgu_cdac_8bit_array_2.drv<31:0> 0.321667
R2997 hgu_cdac_8bit_array_2.drv<31:0>.n230 hgu_cdac_8bit_array_2.drv<31:0> 0.321667
R2998 hgu_cdac_8bit_array_2.drv<31:0>.n221 hgu_cdac_8bit_array_2.drv<31:0> 0.321667
R2999 hgu_cdac_8bit_array_2.drv<31:0>.n203 hgu_cdac_8bit_array_2.drv<31:0> 0.321667
R3000 hgu_cdac_8bit_array_2.drv<31:0>.n194 hgu_cdac_8bit_array_2.drv<31:0> 0.321667
R3001 hgu_cdac_8bit_array_2.drv<31:0>.n185 hgu_cdac_8bit_array_2.drv<31:0> 0.321667
R3002 hgu_cdac_8bit_array_2.drv<31:0>.n176 hgu_cdac_8bit_array_2.drv<31:0> 0.321667
R3003 hgu_cdac_8bit_array_2.drv<31:0>.n167 hgu_cdac_8bit_array_2.drv<31:0> 0.321667
R3004 hgu_cdac_8bit_array_2.drv<31:0>.n158 hgu_cdac_8bit_array_2.drv<31:0> 0.321667
R3005 hgu_cdac_8bit_array_2.drv<31:0>.n149 hgu_cdac_8bit_array_2.drv<31:0> 0.321667
R3006 hgu_cdac_8bit_array_2.drv<31:0>.n140 hgu_cdac_8bit_array_2.drv<31:0> 0.321667
R3007 hgu_cdac_8bit_array_2.drv<31:0>.n131 hgu_cdac_8bit_array_2.drv<31:0> 0.321667
R3008 hgu_cdac_8bit_array_2.drv<31:0>.n112 hgu_cdac_8bit_array_2.drv<31:0>.n111 0.314299
R3009 hgu_cdac_8bit_array_2.drv<31:0>.n0 hgu_cdac_8bit_array_2.drv<31:0>.n129 0.314299
R3010 hgu_cdac_8bit_array_2.drv<31:0>.n256 hgu_cdac_8bit_array_2.drv<31:0> 0.313448
R3011 hgu_cdac_8bit_array_2.drv<31:0>.n128 hgu_cdac_8bit_array_2.drv<31:0>.n85 0.297179
R3012 hgu_cdac_8bit_array_2.drv<31:0>.n127 hgu_cdac_8bit_array_2.drv<31:0>.n87 0.297179
R3013 hgu_cdac_8bit_array_2.drv<31:0>.n126 hgu_cdac_8bit_array_2.drv<31:0>.n89 0.297179
R3014 hgu_cdac_8bit_array_2.drv<31:0>.n125 hgu_cdac_8bit_array_2.drv<31:0>.n91 0.297179
R3015 hgu_cdac_8bit_array_2.drv<31:0>.n124 hgu_cdac_8bit_array_2.drv<31:0>.n93 0.297179
R3016 hgu_cdac_8bit_array_2.drv<31:0>.n123 hgu_cdac_8bit_array_2.drv<31:0>.n95 0.297179
R3017 hgu_cdac_8bit_array_2.drv<31:0>.n122 hgu_cdac_8bit_array_2.drv<31:0>.n97 0.297179
R3018 hgu_cdac_8bit_array_2.drv<31:0>.n121 hgu_cdac_8bit_array_2.drv<31:0>.n99 0.297179
R3019 hgu_cdac_8bit_array_2.drv<31:0>.n120 hgu_cdac_8bit_array_2.drv<31:0>.n101 0.297179
R3020 hgu_cdac_8bit_array_2.drv<31:0>.n119 hgu_cdac_8bit_array_2.drv<31:0>.n103 0.297179
R3021 hgu_cdac_8bit_array_2.drv<31:0>.n118 hgu_cdac_8bit_array_2.drv<31:0>.n105 0.297179
R3022 hgu_cdac_8bit_array_2.drv<31:0>.n117 hgu_cdac_8bit_array_2.drv<31:0>.n107 0.297179
R3023 hgu_cdac_8bit_array_2.drv<31:0>.n116 hgu_cdac_8bit_array_2.drv<31:0>.n109 0.297179
R3024 hgu_cdac_8bit_array_2.drv<31:0>.n115 hgu_cdac_8bit_array_2.drv<31:0>.n114 0.297179
R3025 hgu_cdac_8bit_array_2.drv<31:0>.n134 hgu_cdac_8bit_array_2.drv<31:0> 0.2966
R3026 hgu_cdac_8bit_array_2.drv<31:0>.n143 hgu_cdac_8bit_array_2.drv<31:0> 0.2966
R3027 hgu_cdac_8bit_array_2.drv<31:0>.n152 hgu_cdac_8bit_array_2.drv<31:0> 0.2966
R3028 hgu_cdac_8bit_array_2.drv<31:0>.n161 hgu_cdac_8bit_array_2.drv<31:0> 0.2966
R3029 hgu_cdac_8bit_array_2.drv<31:0>.n170 hgu_cdac_8bit_array_2.drv<31:0> 0.2966
R3030 hgu_cdac_8bit_array_2.drv<31:0>.n179 hgu_cdac_8bit_array_2.drv<31:0> 0.2966
R3031 hgu_cdac_8bit_array_2.drv<31:0>.n188 hgu_cdac_8bit_array_2.drv<31:0> 0.2966
R3032 hgu_cdac_8bit_array_2.drv<31:0>.n197 hgu_cdac_8bit_array_2.drv<31:0> 0.2966
R3033 hgu_cdac_8bit_array_2.drv<31:0>.n206 hgu_cdac_8bit_array_2.drv<31:0> 0.2966
R3034 hgu_cdac_8bit_array_2.drv<31:0>.n215 hgu_cdac_8bit_array_2.drv<31:0> 0.2966
R3035 hgu_cdac_8bit_array_2.drv<31:0>.n224 hgu_cdac_8bit_array_2.drv<31:0> 0.2966
R3036 hgu_cdac_8bit_array_2.drv<31:0>.n233 hgu_cdac_8bit_array_2.drv<31:0> 0.2966
R3037 hgu_cdac_8bit_array_2.drv<31:0>.n242 hgu_cdac_8bit_array_2.drv<31:0> 0.2966
R3038 hgu_cdac_8bit_array_2.drv<31:0>.n272 hgu_cdac_8bit_array_2.drv<31:0> 0.2966
R3039 hgu_cdac_8bit_array_2.drv<31:0>.n263 hgu_cdac_8bit_array_2.drv<31:0> 0.2966
R3040 hgu_cdac_8bit_array_2.drv<31:0>.n212 hgu_cdac_8bit_array_2.drv<31:0> 0.248033
R3041 hgu_cdac_8bit_array_2.drv<31:0>.n131 hgu_cdac_8bit_array_2.drv<31:0>.n130 0.240666
R3042 hgu_cdac_8bit_array_2.drv<31:0>.n137 hgu_cdac_8bit_array_2.drv<31:0>.n136 0.0716912
R3043 hgu_cdac_8bit_array_2.drv<31:0>.n138 hgu_cdac_8bit_array_2.drv<31:0>.n137 0.0716912
R3044 hgu_cdac_8bit_array_2.drv<31:0>.n146 hgu_cdac_8bit_array_2.drv<31:0>.n145 0.0716912
R3045 hgu_cdac_8bit_array_2.drv<31:0>.n147 hgu_cdac_8bit_array_2.drv<31:0>.n146 0.0716912
R3046 hgu_cdac_8bit_array_2.drv<31:0>.n155 hgu_cdac_8bit_array_2.drv<31:0>.n154 0.0716912
R3047 hgu_cdac_8bit_array_2.drv<31:0>.n156 hgu_cdac_8bit_array_2.drv<31:0>.n155 0.0716912
R3048 hgu_cdac_8bit_array_2.drv<31:0>.n164 hgu_cdac_8bit_array_2.drv<31:0>.n163 0.0716912
R3049 hgu_cdac_8bit_array_2.drv<31:0>.n165 hgu_cdac_8bit_array_2.drv<31:0>.n164 0.0716912
R3050 hgu_cdac_8bit_array_2.drv<31:0>.n173 hgu_cdac_8bit_array_2.drv<31:0>.n172 0.0716912
R3051 hgu_cdac_8bit_array_2.drv<31:0>.n174 hgu_cdac_8bit_array_2.drv<31:0>.n173 0.0716912
R3052 hgu_cdac_8bit_array_2.drv<31:0>.n182 hgu_cdac_8bit_array_2.drv<31:0>.n181 0.0716912
R3053 hgu_cdac_8bit_array_2.drv<31:0>.n183 hgu_cdac_8bit_array_2.drv<31:0>.n182 0.0716912
R3054 hgu_cdac_8bit_array_2.drv<31:0>.n191 hgu_cdac_8bit_array_2.drv<31:0>.n190 0.0716912
R3055 hgu_cdac_8bit_array_2.drv<31:0>.n192 hgu_cdac_8bit_array_2.drv<31:0>.n191 0.0716912
R3056 hgu_cdac_8bit_array_2.drv<31:0>.n200 hgu_cdac_8bit_array_2.drv<31:0>.n199 0.0716912
R3057 hgu_cdac_8bit_array_2.drv<31:0>.n201 hgu_cdac_8bit_array_2.drv<31:0>.n200 0.0716912
R3058 hgu_cdac_8bit_array_2.drv<31:0>.n209 hgu_cdac_8bit_array_2.drv<31:0>.n208 0.0716912
R3059 hgu_cdac_8bit_array_2.drv<31:0>.n210 hgu_cdac_8bit_array_2.drv<31:0>.n209 0.0716912
R3060 hgu_cdac_8bit_array_2.drv<31:0>.n218 hgu_cdac_8bit_array_2.drv<31:0>.n217 0.0716912
R3061 hgu_cdac_8bit_array_2.drv<31:0>.n219 hgu_cdac_8bit_array_2.drv<31:0>.n218 0.0716912
R3062 hgu_cdac_8bit_array_2.drv<31:0>.n227 hgu_cdac_8bit_array_2.drv<31:0>.n226 0.0716912
R3063 hgu_cdac_8bit_array_2.drv<31:0>.n228 hgu_cdac_8bit_array_2.drv<31:0>.n227 0.0716912
R3064 hgu_cdac_8bit_array_2.drv<31:0>.n236 hgu_cdac_8bit_array_2.drv<31:0>.n235 0.0716912
R3065 hgu_cdac_8bit_array_2.drv<31:0>.n237 hgu_cdac_8bit_array_2.drv<31:0>.n236 0.0716912
R3066 hgu_cdac_8bit_array_2.drv<31:0>.n245 hgu_cdac_8bit_array_2.drv<31:0>.n244 0.0716912
R3067 hgu_cdac_8bit_array_2.drv<31:0>.n270 hgu_cdac_8bit_array_2.drv<31:0>.n269 0.0716912
R3068 hgu_cdac_8bit_array_2.drv<31:0>.n269 hgu_cdac_8bit_array_2.drv<31:0>.n268 0.0716912
R3069 hgu_cdac_8bit_array_2.drv<31:0>.n261 hgu_cdac_8bit_array_2.drv<31:0>.n260 0.0716912
R3070 hgu_cdac_8bit_array_2.drv<31:0>.n260 hgu_cdac_8bit_array_2.drv<31:0>.n259 0.0716912
R3071 hgu_cdac_8bit_array_2.drv<31:0>.n82 hgu_cdac_8bit_array_2.drv<31:0>.n81 0.0716912
R3072 hgu_cdac_8bit_array_2.drv<31:0>.n77 hgu_cdac_8bit_array_2.drv<31:0>.n76 0.0716912
R3073 hgu_cdac_8bit_array_2.drv<31:0>.n70 hgu_cdac_8bit_array_2.drv<31:0>.n69 0.0716912
R3074 hgu_cdac_8bit_array_2.drv<31:0>.n63 hgu_cdac_8bit_array_2.drv<31:0>.n62 0.0716912
R3075 hgu_cdac_8bit_array_2.drv<31:0>.n56 hgu_cdac_8bit_array_2.drv<31:0>.n55 0.0716912
R3076 hgu_cdac_8bit_array_2.drv<31:0>.n49 hgu_cdac_8bit_array_2.drv<31:0>.n48 0.0716912
R3077 hgu_cdac_8bit_array_2.drv<31:0>.n42 hgu_cdac_8bit_array_2.drv<31:0>.n41 0.0716912
R3078 hgu_cdac_8bit_array_2.drv<31:0>.n35 hgu_cdac_8bit_array_2.drv<31:0>.n34 0.0716912
R3079 hgu_cdac_8bit_array_2.drv<31:0>.n28 hgu_cdac_8bit_array_2.drv<31:0>.n27 0.0716912
R3080 hgu_cdac_8bit_array_2.drv<31:0>.n21 hgu_cdac_8bit_array_2.drv<31:0>.n20 0.0716912
R3081 hgu_cdac_8bit_array_2.drv<31:0>.n14 hgu_cdac_8bit_array_2.drv<31:0>.n13 0.0716912
R3082 hgu_cdac_8bit_array_2.drv<31:0>.n7 hgu_cdac_8bit_array_2.drv<31:0>.n6 0.0716912
R3083 hgu_cdac_8bit_array_2.drv<31:0>.n252 hgu_cdac_8bit_array_2.drv<31:0>.n251 0.0716912
R3084 hgu_cdac_8bit_array_2.drv<31:0>.n255 hgu_cdac_8bit_array_2.drv<31:0>.n254 0.0716912
R3085 hgu_cdac_8bit_array_2.drv<31:0>.n257 hgu_cdac_8bit_array_2.drv<31:0>.n256 0.0664894
R3086 hgu_cdac_8bit_array_2.drv<31:0>.n133 hgu_cdac_8bit_array_2.drv<31:0>.n132 0.0557941
R3087 hgu_cdac_8bit_array_2.drv<31:0>.n136 hgu_cdac_8bit_array_2.drv<31:0>.n135 0.0557941
R3088 hgu_cdac_8bit_array_2.drv<31:0>.n139 hgu_cdac_8bit_array_2.drv<31:0>.n138 0.0557941
R3089 hgu_cdac_8bit_array_2.drv<31:0>.n142 hgu_cdac_8bit_array_2.drv<31:0>.n141 0.0557941
R3090 hgu_cdac_8bit_array_2.drv<31:0>.n145 hgu_cdac_8bit_array_2.drv<31:0>.n144 0.0557941
R3091 hgu_cdac_8bit_array_2.drv<31:0>.n148 hgu_cdac_8bit_array_2.drv<31:0>.n147 0.0557941
R3092 hgu_cdac_8bit_array_2.drv<31:0>.n151 hgu_cdac_8bit_array_2.drv<31:0>.n150 0.0557941
R3093 hgu_cdac_8bit_array_2.drv<31:0>.n154 hgu_cdac_8bit_array_2.drv<31:0>.n153 0.0557941
R3094 hgu_cdac_8bit_array_2.drv<31:0>.n157 hgu_cdac_8bit_array_2.drv<31:0>.n156 0.0557941
R3095 hgu_cdac_8bit_array_2.drv<31:0>.n160 hgu_cdac_8bit_array_2.drv<31:0>.n159 0.0557941
R3096 hgu_cdac_8bit_array_2.drv<31:0>.n163 hgu_cdac_8bit_array_2.drv<31:0>.n162 0.0557941
R3097 hgu_cdac_8bit_array_2.drv<31:0>.n166 hgu_cdac_8bit_array_2.drv<31:0>.n165 0.0557941
R3098 hgu_cdac_8bit_array_2.drv<31:0>.n169 hgu_cdac_8bit_array_2.drv<31:0>.n168 0.0557941
R3099 hgu_cdac_8bit_array_2.drv<31:0>.n172 hgu_cdac_8bit_array_2.drv<31:0>.n171 0.0557941
R3100 hgu_cdac_8bit_array_2.drv<31:0>.n175 hgu_cdac_8bit_array_2.drv<31:0>.n174 0.0557941
R3101 hgu_cdac_8bit_array_2.drv<31:0>.n178 hgu_cdac_8bit_array_2.drv<31:0>.n177 0.0557941
R3102 hgu_cdac_8bit_array_2.drv<31:0>.n181 hgu_cdac_8bit_array_2.drv<31:0>.n180 0.0557941
R3103 hgu_cdac_8bit_array_2.drv<31:0>.n184 hgu_cdac_8bit_array_2.drv<31:0>.n183 0.0557941
R3104 hgu_cdac_8bit_array_2.drv<31:0>.n187 hgu_cdac_8bit_array_2.drv<31:0>.n186 0.0557941
R3105 hgu_cdac_8bit_array_2.drv<31:0>.n190 hgu_cdac_8bit_array_2.drv<31:0>.n189 0.0557941
R3106 hgu_cdac_8bit_array_2.drv<31:0>.n193 hgu_cdac_8bit_array_2.drv<31:0>.n192 0.0557941
R3107 hgu_cdac_8bit_array_2.drv<31:0>.n196 hgu_cdac_8bit_array_2.drv<31:0>.n195 0.0557941
R3108 hgu_cdac_8bit_array_2.drv<31:0>.n199 hgu_cdac_8bit_array_2.drv<31:0>.n198 0.0557941
R3109 hgu_cdac_8bit_array_2.drv<31:0>.n202 hgu_cdac_8bit_array_2.drv<31:0>.n201 0.0557941
R3110 hgu_cdac_8bit_array_2.drv<31:0>.n205 hgu_cdac_8bit_array_2.drv<31:0>.n204 0.0557941
R3111 hgu_cdac_8bit_array_2.drv<31:0>.n208 hgu_cdac_8bit_array_2.drv<31:0>.n207 0.0557941
R3112 hgu_cdac_8bit_array_2.drv<31:0>.n211 hgu_cdac_8bit_array_2.drv<31:0>.n210 0.0557941
R3113 hgu_cdac_8bit_array_2.drv<31:0>.n214 hgu_cdac_8bit_array_2.drv<31:0>.n213 0.0557941
R3114 hgu_cdac_8bit_array_2.drv<31:0>.n217 hgu_cdac_8bit_array_2.drv<31:0>.n216 0.0557941
R3115 hgu_cdac_8bit_array_2.drv<31:0>.n220 hgu_cdac_8bit_array_2.drv<31:0>.n219 0.0557941
R3116 hgu_cdac_8bit_array_2.drv<31:0>.n223 hgu_cdac_8bit_array_2.drv<31:0>.n222 0.0557941
R3117 hgu_cdac_8bit_array_2.drv<31:0>.n226 hgu_cdac_8bit_array_2.drv<31:0>.n225 0.0557941
R3118 hgu_cdac_8bit_array_2.drv<31:0>.n229 hgu_cdac_8bit_array_2.drv<31:0>.n228 0.0557941
R3119 hgu_cdac_8bit_array_2.drv<31:0>.n232 hgu_cdac_8bit_array_2.drv<31:0>.n231 0.0557941
R3120 hgu_cdac_8bit_array_2.drv<31:0>.n235 hgu_cdac_8bit_array_2.drv<31:0>.n234 0.0557941
R3121 hgu_cdac_8bit_array_2.drv<31:0>.n238 hgu_cdac_8bit_array_2.drv<31:0>.n237 0.0557941
R3122 hgu_cdac_8bit_array_2.drv<31:0>.n241 hgu_cdac_8bit_array_2.drv<31:0>.n240 0.0557941
R3123 hgu_cdac_8bit_array_2.drv<31:0>.n244 hgu_cdac_8bit_array_2.drv<31:0>.n243 0.0557941
R3124 hgu_cdac_8bit_array_2.drv<31:0>.n277 hgu_cdac_8bit_array_2.drv<31:0>.n276 0.0557941
R3125 hgu_cdac_8bit_array_2.drv<31:0>.n274 hgu_cdac_8bit_array_2.drv<31:0>.n273 0.0557941
R3126 hgu_cdac_8bit_array_2.drv<31:0>.n271 hgu_cdac_8bit_array_2.drv<31:0>.n270 0.0557941
R3127 hgu_cdac_8bit_array_2.drv<31:0>.n268 hgu_cdac_8bit_array_2.drv<31:0>.n267 0.0557941
R3128 hgu_cdac_8bit_array_2.drv<31:0>.n265 hgu_cdac_8bit_array_2.drv<31:0>.n264 0.0557941
R3129 hgu_cdac_8bit_array_2.drv<31:0>.n262 hgu_cdac_8bit_array_2.drv<31:0>.n261 0.0557941
R3130 hgu_cdac_8bit_array_2.drv<31:0>.n259 hgu_cdac_8bit_array_2.drv<31:0>.n258 0.0557941
R3131 hgu_cdac_8bit_array_2.drv<31:0>.n79 hgu_cdac_8bit_array_2.drv<31:0>.n78 0.0557941
R3132 hgu_cdac_8bit_array_2.drv<31:0>.n80 hgu_cdac_8bit_array_2.drv<31:0>.n79 0.0557941
R3133 hgu_cdac_8bit_array_2.drv<31:0>.n81 hgu_cdac_8bit_array_2.drv<31:0>.n80 0.0557941
R3134 hgu_cdac_8bit_array_2.drv<31:0>.n72 hgu_cdac_8bit_array_2.drv<31:0>.n71 0.0557941
R3135 hgu_cdac_8bit_array_2.drv<31:0>.n73 hgu_cdac_8bit_array_2.drv<31:0>.n72 0.0557941
R3136 hgu_cdac_8bit_array_2.drv<31:0>.n74 hgu_cdac_8bit_array_2.drv<31:0>.n73 0.0557941
R3137 hgu_cdac_8bit_array_2.drv<31:0>.n75 hgu_cdac_8bit_array_2.drv<31:0>.n74 0.0557941
R3138 hgu_cdac_8bit_array_2.drv<31:0>.n76 hgu_cdac_8bit_array_2.drv<31:0>.n75 0.0557941
R3139 hgu_cdac_8bit_array_2.drv<31:0>.n65 hgu_cdac_8bit_array_2.drv<31:0>.n64 0.0557941
R3140 hgu_cdac_8bit_array_2.drv<31:0>.n66 hgu_cdac_8bit_array_2.drv<31:0>.n65 0.0557941
R3141 hgu_cdac_8bit_array_2.drv<31:0>.n67 hgu_cdac_8bit_array_2.drv<31:0>.n66 0.0557941
R3142 hgu_cdac_8bit_array_2.drv<31:0>.n68 hgu_cdac_8bit_array_2.drv<31:0>.n67 0.0557941
R3143 hgu_cdac_8bit_array_2.drv<31:0>.n69 hgu_cdac_8bit_array_2.drv<31:0>.n68 0.0557941
R3144 hgu_cdac_8bit_array_2.drv<31:0>.n58 hgu_cdac_8bit_array_2.drv<31:0>.n57 0.0557941
R3145 hgu_cdac_8bit_array_2.drv<31:0>.n59 hgu_cdac_8bit_array_2.drv<31:0>.n58 0.0557941
R3146 hgu_cdac_8bit_array_2.drv<31:0>.n60 hgu_cdac_8bit_array_2.drv<31:0>.n59 0.0557941
R3147 hgu_cdac_8bit_array_2.drv<31:0>.n61 hgu_cdac_8bit_array_2.drv<31:0>.n60 0.0557941
R3148 hgu_cdac_8bit_array_2.drv<31:0>.n62 hgu_cdac_8bit_array_2.drv<31:0>.n61 0.0557941
R3149 hgu_cdac_8bit_array_2.drv<31:0>.n51 hgu_cdac_8bit_array_2.drv<31:0>.n50 0.0557941
R3150 hgu_cdac_8bit_array_2.drv<31:0>.n52 hgu_cdac_8bit_array_2.drv<31:0>.n51 0.0557941
R3151 hgu_cdac_8bit_array_2.drv<31:0>.n53 hgu_cdac_8bit_array_2.drv<31:0>.n52 0.0557941
R3152 hgu_cdac_8bit_array_2.drv<31:0>.n54 hgu_cdac_8bit_array_2.drv<31:0>.n53 0.0557941
R3153 hgu_cdac_8bit_array_2.drv<31:0>.n55 hgu_cdac_8bit_array_2.drv<31:0>.n54 0.0557941
R3154 hgu_cdac_8bit_array_2.drv<31:0>.n44 hgu_cdac_8bit_array_2.drv<31:0>.n43 0.0557941
R3155 hgu_cdac_8bit_array_2.drv<31:0>.n45 hgu_cdac_8bit_array_2.drv<31:0>.n44 0.0557941
R3156 hgu_cdac_8bit_array_2.drv<31:0>.n46 hgu_cdac_8bit_array_2.drv<31:0>.n45 0.0557941
R3157 hgu_cdac_8bit_array_2.drv<31:0>.n47 hgu_cdac_8bit_array_2.drv<31:0>.n46 0.0557941
R3158 hgu_cdac_8bit_array_2.drv<31:0>.n48 hgu_cdac_8bit_array_2.drv<31:0>.n47 0.0557941
R3159 hgu_cdac_8bit_array_2.drv<31:0>.n37 hgu_cdac_8bit_array_2.drv<31:0>.n36 0.0557941
R3160 hgu_cdac_8bit_array_2.drv<31:0>.n38 hgu_cdac_8bit_array_2.drv<31:0>.n37 0.0557941
R3161 hgu_cdac_8bit_array_2.drv<31:0>.n39 hgu_cdac_8bit_array_2.drv<31:0>.n38 0.0557941
R3162 hgu_cdac_8bit_array_2.drv<31:0>.n40 hgu_cdac_8bit_array_2.drv<31:0>.n39 0.0557941
R3163 hgu_cdac_8bit_array_2.drv<31:0>.n41 hgu_cdac_8bit_array_2.drv<31:0>.n40 0.0557941
R3164 hgu_cdac_8bit_array_2.drv<31:0>.n30 hgu_cdac_8bit_array_2.drv<31:0>.n29 0.0557941
R3165 hgu_cdac_8bit_array_2.drv<31:0>.n31 hgu_cdac_8bit_array_2.drv<31:0>.n30 0.0557941
R3166 hgu_cdac_8bit_array_2.drv<31:0>.n32 hgu_cdac_8bit_array_2.drv<31:0>.n31 0.0557941
R3167 hgu_cdac_8bit_array_2.drv<31:0>.n33 hgu_cdac_8bit_array_2.drv<31:0>.n32 0.0557941
R3168 hgu_cdac_8bit_array_2.drv<31:0>.n34 hgu_cdac_8bit_array_2.drv<31:0>.n33 0.0557941
R3169 hgu_cdac_8bit_array_2.drv<31:0>.n23 hgu_cdac_8bit_array_2.drv<31:0>.n22 0.0557941
R3170 hgu_cdac_8bit_array_2.drv<31:0>.n24 hgu_cdac_8bit_array_2.drv<31:0>.n23 0.0557941
R3171 hgu_cdac_8bit_array_2.drv<31:0>.n25 hgu_cdac_8bit_array_2.drv<31:0>.n24 0.0557941
R3172 hgu_cdac_8bit_array_2.drv<31:0>.n26 hgu_cdac_8bit_array_2.drv<31:0>.n25 0.0557941
R3173 hgu_cdac_8bit_array_2.drv<31:0>.n27 hgu_cdac_8bit_array_2.drv<31:0>.n26 0.0557941
R3174 hgu_cdac_8bit_array_2.drv<31:0>.n16 hgu_cdac_8bit_array_2.drv<31:0>.n15 0.0557941
R3175 hgu_cdac_8bit_array_2.drv<31:0>.n17 hgu_cdac_8bit_array_2.drv<31:0>.n16 0.0557941
R3176 hgu_cdac_8bit_array_2.drv<31:0>.n18 hgu_cdac_8bit_array_2.drv<31:0>.n17 0.0557941
R3177 hgu_cdac_8bit_array_2.drv<31:0>.n19 hgu_cdac_8bit_array_2.drv<31:0>.n18 0.0557941
R3178 hgu_cdac_8bit_array_2.drv<31:0>.n20 hgu_cdac_8bit_array_2.drv<31:0>.n19 0.0557941
R3179 hgu_cdac_8bit_array_2.drv<31:0>.n9 hgu_cdac_8bit_array_2.drv<31:0>.n8 0.0557941
R3180 hgu_cdac_8bit_array_2.drv<31:0>.n10 hgu_cdac_8bit_array_2.drv<31:0>.n9 0.0557941
R3181 hgu_cdac_8bit_array_2.drv<31:0>.n11 hgu_cdac_8bit_array_2.drv<31:0>.n10 0.0557941
R3182 hgu_cdac_8bit_array_2.drv<31:0>.n12 hgu_cdac_8bit_array_2.drv<31:0>.n11 0.0557941
R3183 hgu_cdac_8bit_array_2.drv<31:0>.n13 hgu_cdac_8bit_array_2.drv<31:0>.n12 0.0557941
R3184 hgu_cdac_8bit_array_2.drv<31:0>.n2 hgu_cdac_8bit_array_2.drv<31:0>.n1 0.0557941
R3185 hgu_cdac_8bit_array_2.drv<31:0>.n3 hgu_cdac_8bit_array_2.drv<31:0>.n2 0.0557941
R3186 hgu_cdac_8bit_array_2.drv<31:0>.n4 hgu_cdac_8bit_array_2.drv<31:0>.n3 0.0557941
R3187 hgu_cdac_8bit_array_2.drv<31:0>.n5 hgu_cdac_8bit_array_2.drv<31:0>.n4 0.0557941
R3188 hgu_cdac_8bit_array_2.drv<31:0>.n6 hgu_cdac_8bit_array_2.drv<31:0>.n5 0.0557941
R3189 hgu_cdac_8bit_array_2.drv<31:0>.n251 hgu_cdac_8bit_array_2.drv<31:0>.n250 0.0557941
R3190 hgu_cdac_8bit_array_2.drv<31:0>.n250 hgu_cdac_8bit_array_2.drv<31:0>.n249 0.0557941
R3191 hgu_cdac_8bit_array_2.drv<31:0>.n249 hgu_cdac_8bit_array_2.drv<31:0>.n248 0.0557941
R3192 hgu_cdac_8bit_array_2.drv<31:0>.n248 hgu_cdac_8bit_array_2.drv<31:0>.n247 0.0557941
R3193 hgu_cdac_8bit_array_2.drv<31:0>.n247 hgu_cdac_8bit_array_2.drv<31:0>.n246 0.0557941
R3194 hgu_cdac_8bit_array_2.drv<31:0>.n254 hgu_cdac_8bit_array_2.drv<31:0>.n253 0.0557941
R3195 hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_8bit_array_2.drv<31:0>.n277 0.0544118
R3196 hgu_cdac_8bit_array_2.drv<31:0>.n135 hgu_cdac_8bit_array_2.drv<31:0>.n134 0.0419706
R3197 hgu_cdac_8bit_array_2.drv<31:0>.n140 hgu_cdac_8bit_array_2.drv<31:0>.n139 0.0419706
R3198 hgu_cdac_8bit_array_2.drv<31:0>.n144 hgu_cdac_8bit_array_2.drv<31:0>.n143 0.0419706
R3199 hgu_cdac_8bit_array_2.drv<31:0>.n149 hgu_cdac_8bit_array_2.drv<31:0>.n148 0.0419706
R3200 hgu_cdac_8bit_array_2.drv<31:0>.n153 hgu_cdac_8bit_array_2.drv<31:0>.n152 0.0419706
R3201 hgu_cdac_8bit_array_2.drv<31:0>.n158 hgu_cdac_8bit_array_2.drv<31:0>.n157 0.0419706
R3202 hgu_cdac_8bit_array_2.drv<31:0>.n162 hgu_cdac_8bit_array_2.drv<31:0>.n161 0.0419706
R3203 hgu_cdac_8bit_array_2.drv<31:0>.n167 hgu_cdac_8bit_array_2.drv<31:0>.n166 0.0419706
R3204 hgu_cdac_8bit_array_2.drv<31:0>.n171 hgu_cdac_8bit_array_2.drv<31:0>.n170 0.0419706
R3205 hgu_cdac_8bit_array_2.drv<31:0>.n176 hgu_cdac_8bit_array_2.drv<31:0>.n175 0.0419706
R3206 hgu_cdac_8bit_array_2.drv<31:0>.n180 hgu_cdac_8bit_array_2.drv<31:0>.n179 0.0419706
R3207 hgu_cdac_8bit_array_2.drv<31:0>.n185 hgu_cdac_8bit_array_2.drv<31:0>.n184 0.0419706
R3208 hgu_cdac_8bit_array_2.drv<31:0>.n189 hgu_cdac_8bit_array_2.drv<31:0>.n188 0.0419706
R3209 hgu_cdac_8bit_array_2.drv<31:0>.n194 hgu_cdac_8bit_array_2.drv<31:0>.n193 0.0419706
R3210 hgu_cdac_8bit_array_2.drv<31:0>.n198 hgu_cdac_8bit_array_2.drv<31:0>.n197 0.0419706
R3211 hgu_cdac_8bit_array_2.drv<31:0>.n203 hgu_cdac_8bit_array_2.drv<31:0>.n202 0.0419706
R3212 hgu_cdac_8bit_array_2.drv<31:0>.n207 hgu_cdac_8bit_array_2.drv<31:0>.n206 0.0419706
R3213 hgu_cdac_8bit_array_2.drv<31:0>.n212 hgu_cdac_8bit_array_2.drv<31:0>.n211 0.0419706
R3214 hgu_cdac_8bit_array_2.drv<31:0>.n216 hgu_cdac_8bit_array_2.drv<31:0>.n215 0.0419706
R3215 hgu_cdac_8bit_array_2.drv<31:0>.n221 hgu_cdac_8bit_array_2.drv<31:0>.n220 0.0419706
R3216 hgu_cdac_8bit_array_2.drv<31:0>.n225 hgu_cdac_8bit_array_2.drv<31:0>.n224 0.0419706
R3217 hgu_cdac_8bit_array_2.drv<31:0>.n230 hgu_cdac_8bit_array_2.drv<31:0>.n229 0.0419706
R3218 hgu_cdac_8bit_array_2.drv<31:0>.n234 hgu_cdac_8bit_array_2.drv<31:0>.n233 0.0419706
R3219 hgu_cdac_8bit_array_2.drv<31:0>.n239 hgu_cdac_8bit_array_2.drv<31:0>.n238 0.0419706
R3220 hgu_cdac_8bit_array_2.drv<31:0>.n243 hgu_cdac_8bit_array_2.drv<31:0>.n242 0.0419706
R3221 hgu_cdac_8bit_array_2.drv<31:0>.n276 hgu_cdac_8bit_array_2.drv<31:0>.n275 0.0419706
R3222 hgu_cdac_8bit_array_2.drv<31:0>.n272 hgu_cdac_8bit_array_2.drv<31:0>.n271 0.0419706
R3223 hgu_cdac_8bit_array_2.drv<31:0>.n267 hgu_cdac_8bit_array_2.drv<31:0>.n266 0.0419706
R3224 hgu_cdac_8bit_array_2.drv<31:0>.n263 hgu_cdac_8bit_array_2.drv<31:0>.n262 0.0419706
R3225 hgu_cdac_8bit_array_2.drv<31:0>.n258 hgu_cdac_8bit_array_2.drv<31:0>.n257 0.0419706
R3226 hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_8bit_array_2.drv<31:0>.n245 0.0177794
R3227 hgu_cdac_8bit_array_2.drv<31:0>.n132 hgu_cdac_8bit_array_2.drv<31:0>.n131 0.0143235
R3228 hgu_cdac_8bit_array_2.drv<31:0>.n134 hgu_cdac_8bit_array_2.drv<31:0>.n133 0.0143235
R3229 hgu_cdac_8bit_array_2.drv<31:0>.n141 hgu_cdac_8bit_array_2.drv<31:0>.n140 0.0143235
R3230 hgu_cdac_8bit_array_2.drv<31:0>.n143 hgu_cdac_8bit_array_2.drv<31:0>.n142 0.0143235
R3231 hgu_cdac_8bit_array_2.drv<31:0>.n150 hgu_cdac_8bit_array_2.drv<31:0>.n149 0.0143235
R3232 hgu_cdac_8bit_array_2.drv<31:0>.n152 hgu_cdac_8bit_array_2.drv<31:0>.n151 0.0143235
R3233 hgu_cdac_8bit_array_2.drv<31:0>.n159 hgu_cdac_8bit_array_2.drv<31:0>.n158 0.0143235
R3234 hgu_cdac_8bit_array_2.drv<31:0>.n161 hgu_cdac_8bit_array_2.drv<31:0>.n160 0.0143235
R3235 hgu_cdac_8bit_array_2.drv<31:0>.n168 hgu_cdac_8bit_array_2.drv<31:0>.n167 0.0143235
R3236 hgu_cdac_8bit_array_2.drv<31:0>.n170 hgu_cdac_8bit_array_2.drv<31:0>.n169 0.0143235
R3237 hgu_cdac_8bit_array_2.drv<31:0>.n177 hgu_cdac_8bit_array_2.drv<31:0>.n176 0.0143235
R3238 hgu_cdac_8bit_array_2.drv<31:0>.n179 hgu_cdac_8bit_array_2.drv<31:0>.n178 0.0143235
R3239 hgu_cdac_8bit_array_2.drv<31:0>.n186 hgu_cdac_8bit_array_2.drv<31:0>.n185 0.0143235
R3240 hgu_cdac_8bit_array_2.drv<31:0>.n188 hgu_cdac_8bit_array_2.drv<31:0>.n187 0.0143235
R3241 hgu_cdac_8bit_array_2.drv<31:0>.n195 hgu_cdac_8bit_array_2.drv<31:0>.n194 0.0143235
R3242 hgu_cdac_8bit_array_2.drv<31:0>.n197 hgu_cdac_8bit_array_2.drv<31:0>.n196 0.0143235
R3243 hgu_cdac_8bit_array_2.drv<31:0>.n204 hgu_cdac_8bit_array_2.drv<31:0>.n203 0.0143235
R3244 hgu_cdac_8bit_array_2.drv<31:0>.n206 hgu_cdac_8bit_array_2.drv<31:0>.n205 0.0143235
R3245 hgu_cdac_8bit_array_2.drv<31:0>.n213 hgu_cdac_8bit_array_2.drv<31:0>.n212 0.0143235
R3246 hgu_cdac_8bit_array_2.drv<31:0>.n215 hgu_cdac_8bit_array_2.drv<31:0>.n214 0.0143235
R3247 hgu_cdac_8bit_array_2.drv<31:0>.n222 hgu_cdac_8bit_array_2.drv<31:0>.n221 0.0143235
R3248 hgu_cdac_8bit_array_2.drv<31:0>.n224 hgu_cdac_8bit_array_2.drv<31:0>.n223 0.0143235
R3249 hgu_cdac_8bit_array_2.drv<31:0>.n231 hgu_cdac_8bit_array_2.drv<31:0>.n230 0.0143235
R3250 hgu_cdac_8bit_array_2.drv<31:0>.n233 hgu_cdac_8bit_array_2.drv<31:0>.n232 0.0143235
R3251 hgu_cdac_8bit_array_2.drv<31:0>.n240 hgu_cdac_8bit_array_2.drv<31:0>.n239 0.0143235
R3252 hgu_cdac_8bit_array_2.drv<31:0>.n242 hgu_cdac_8bit_array_2.drv<31:0>.n241 0.0143235
R3253 hgu_cdac_8bit_array_2.drv<31:0>.n275 hgu_cdac_8bit_array_2.drv<31:0>.n274 0.0143235
R3254 hgu_cdac_8bit_array_2.drv<31:0>.n273 hgu_cdac_8bit_array_2.drv<31:0>.n272 0.0143235
R3255 hgu_cdac_8bit_array_2.drv<31:0>.n266 hgu_cdac_8bit_array_2.drv<31:0>.n265 0.0143235
R3256 hgu_cdac_8bit_array_2.drv<31:0>.n264 hgu_cdac_8bit_array_2.drv<31:0>.n263 0.0143235
R3257 d<6>.n1 d<6>.n0 88.1376
R3258 d<6>.n2 d<6>.n1 88.1376
R3259 d<6>.n3 d<6>.n2 88.1376
R3260 d<6>.n4 d<6>.n3 88.1376
R3261 d<6>.n5 d<6>.n4 88.1376
R3262 d<6>.n6 d<6>.n5 88.1376
R3263 d<6>.n7 d<6>.n6 88.1376
R3264 d<6>.n8 d<6>.n7 88.1376
R3265 d<6>.n9 d<6>.n8 88.1376
R3266 d<6>.n10 d<6>.n9 88.1376
R3267 d<6>.n11 d<6>.n10 88.1376
R3268 d<6>.n12 d<6>.n11 88.1376
R3269 d<6>.n13 d<6>.n12 88.1376
R3270 d<6>.n14 d<6>.n13 88.1376
R3271 d<6>.n15 d<6>.n14 88.1376
R3272 d<6>.n16 d<6>.n15 88.1376
R3273 d<6>.n17 d<6>.n16 88.1376
R3274 d<6>.n18 d<6>.n17 88.1376
R3275 d<6>.n19 d<6>.n18 88.1376
R3276 d<6>.n20 d<6>.n19 88.1376
R3277 d<6>.n21 d<6>.n20 88.1376
R3278 d<6>.n22 d<6>.n21 88.1376
R3279 d<6>.n23 d<6>.n22 88.1376
R3280 d<6>.n24 d<6>.n23 88.1376
R3281 d<6>.n25 d<6>.n24 88.1376
R3282 d<6>.n26 d<6>.n25 88.1376
R3283 d<6>.n27 d<6>.n26 88.1376
R3284 d<6>.n28 d<6>.n27 88.1376
R3285 d<6>.n29 d<6>.n28 88.1376
R3286 d<6>.n30 d<6>.n29 88.1376
R3287 d<6>.n31 d<6>.n30 88.1376
R3288 d<6>.n32 d<6>.n31 88.1376
R3289 d<6>.n33 d<6>.n32 88.1376
R3290 d<6>.n34 d<6>.n33 88.1376
R3291 d<6>.n35 d<6>.n34 88.1376
R3292 d<6>.n36 d<6>.n35 88.1376
R3293 d<6>.n37 d<6>.n36 88.1376
R3294 d<6>.n38 d<6>.n37 88.1376
R3295 d<6>.n39 d<6>.n38 88.1376
R3296 d<6>.n40 d<6>.n39 88.1376
R3297 d<6>.n41 d<6>.n40 88.1376
R3298 d<6>.n42 d<6>.n41 88.1376
R3299 d<6>.n43 d<6>.n42 88.1376
R3300 d<6>.n44 d<6>.n43 88.1376
R3301 d<6>.n45 d<6>.n44 88.1376
R3302 d<6>.n46 d<6>.n45 88.1376
R3303 d<6>.n47 d<6>.n46 88.1376
R3304 d<6>.n48 d<6>.n47 88.1376
R3305 d<6>.n49 d<6>.n48 88.1376
R3306 d<6>.n50 d<6>.n49 88.1376
R3307 d<6>.n51 d<6>.n50 88.1376
R3308 d<6>.n52 d<6>.n51 88.1376
R3309 d<6>.n53 d<6>.n52 88.1376
R3310 d<6>.n54 d<6>.n53 88.1376
R3311 d<6>.n55 d<6>.n54 88.1376
R3312 d<6>.n56 d<6>.n55 88.1376
R3313 d<6>.n57 d<6>.n56 88.1376
R3314 d<6>.n58 d<6>.n57 88.1376
R3315 d<6>.n59 d<6>.n58 88.1376
R3316 d<6>.n60 d<6>.n59 88.1376
R3317 d<6>.n61 d<6>.n60 88.1376
R3318 d<6>.n62 d<6>.n61 88.1376
R3319 d<6>.n63 d<6>.n62 88.1376
R3320 d<6>.n0 d<6>.t30 69.5462
R3321 d<6>.n1 d<6>.t47 69.5462
R3322 d<6>.n2 d<6>.t123 69.5462
R3323 d<6>.n3 d<6>.t76 69.5462
R3324 d<6>.n4 d<6>.t19 69.5462
R3325 d<6>.n5 d<6>.t98 69.5462
R3326 d<6>.n6 d<6>.t83 69.5462
R3327 d<6>.n7 d<6>.t39 69.5462
R3328 d<6>.n8 d<6>.t22 69.5462
R3329 d<6>.n9 d<6>.t100 69.5462
R3330 d<6>.n10 d<6>.t58 69.5462
R3331 d<6>.n11 d<6>.t44 69.5462
R3332 d<6>.n12 d<6>.t107 69.5462
R3333 d<6>.n13 d<6>.t63 69.5462
R3334 d<6>.n14 d<6>.t16 69.5462
R3335 d<6>.n15 d<6>.t127 69.5462
R3336 d<6>.n16 d<6>.t111 69.5462
R3337 d<6>.n17 d<6>.t67 69.5462
R3338 d<6>.n18 d<6>.t18 69.5462
R3339 d<6>.n19 d<6>.t3 69.5462
R3340 d<6>.n20 d<6>.t42 69.5462
R3341 d<6>.n21 d<6>.t28 69.5462
R3342 d<6>.n22 d<6>.t9 69.5462
R3343 d<6>.n23 d<6>.t89 69.5462
R3344 d<6>.n24 d<6>.t46 69.5462
R3345 d<6>.n25 d<6>.t122 69.5462
R3346 d<6>.n26 d<6>.t13 69.5462
R3347 d<6>.n27 d<6>.t93 69.5462
R3348 d<6>.n28 d<6>.t4 69.5462
R3349 d<6>.n29 d<6>.t114 69.5462
R3350 d<6>.n30 d<6>.t71 69.5462
R3351 d<6>.n31 d<6>.t57 69.5462
R3352 d<6>.n32 d<6>.t6 69.5462
R3353 d<6>.n33 d<6>.t116 69.5462
R3354 d<6>.n34 d<6>.t74 69.5462
R3355 d<6>.n35 d<6>.t27 69.5462
R3356 d<6>.n36 d<6>.t94 69.5462
R3357 d<6>.n37 d<6>.t78 69.5462
R3358 d<6>.n38 d<6>.t34 69.5462
R3359 d<6>.n39 d<6>.t110 69.5462
R3360 d<6>.n40 d<6>.t96 69.5462
R3361 d<6>.n41 d<6>.t81 69.5462
R3362 d<6>.n42 d<6>.t36 69.5462
R3363 d<6>.n43 d<6>.t113 69.5462
R3364 d<6>.n44 d<6>.t59 69.5462
R3365 d<6>.n45 d<6>.t8 69.5462
R3366 d<6>.n46 d<6>.t120 69.5462
R3367 d<6>.n47 d<6>.t105 69.5462
R3368 d<6>.n48 d<6>.t61 69.5462
R3369 d<6>.n49 d<6>.t12 69.5462
R3370 d<6>.n50 d<6>.t91 69.5462
R3371 d<6>.n51 d<6>.t70 69.5462
R3372 d<6>.n52 d<6>.t20 69.5462
R3373 d<6>.n53 d<6>.t99 69.5462
R3374 d<6>.n54 d<6>.t84 69.5462
R3375 d<6>.n55 d<6>.t40 69.5462
R3376 d<6>.n56 d<6>.t24 69.5462
R3377 d<6>.n57 d<6>.t101 69.5462
R3378 d<6>.n58 d<6>.t86 69.5462
R3379 d<6>.n59 d<6>.t124 69.5462
R3380 d<6>.n60 d<6>.t77 69.5462
R3381 d<6>.n61 d<6>.t64 69.5462
R3382 d<6>.n62 d<6>.t51 69.5462
R3383 d<6>.n63 d<6>.t0 69.5462
R3384 d<6>.n0 d<6>.t56 59.9062
R3385 d<6>.n1 d<6>.t73 59.9062
R3386 d<6>.n2 d<6>.t25 59.9062
R3387 d<6>.n3 d<6>.t102 59.9062
R3388 d<6>.n4 d<6>.t49 59.9062
R3389 d<6>.n5 d<6>.t125 59.9062
R3390 d<6>.n6 d<6>.t109 59.9062
R3391 d<6>.n7 d<6>.t66 59.9062
R3392 d<6>.n8 d<6>.t52 59.9062
R3393 d<6>.n9 d<6>.t1 59.9062
R3394 d<6>.n10 d<6>.t80 59.9062
R3395 d<6>.n11 d<6>.t69 59.9062
R3396 d<6>.n12 d<6>.t7 59.9062
R3397 d<6>.n13 d<6>.t87 59.9062
R3398 d<6>.n14 d<6>.t45 59.9062
R3399 d<6>.n15 d<6>.t29 59.9062
R3400 d<6>.n16 d<6>.t11 59.9062
R3401 d<6>.n17 d<6>.t90 59.9062
R3402 d<6>.n18 d<6>.t48 59.9062
R3403 d<6>.n19 d<6>.t32 59.9062
R3404 d<6>.n20 d<6>.t68 59.9062
R3405 d<6>.n21 d<6>.t55 59.9062
R3406 d<6>.n22 d<6>.t38 59.9062
R3407 d<6>.n23 d<6>.t115 59.9062
R3408 d<6>.n24 d<6>.t72 59.9062
R3409 d<6>.n25 d<6>.t23 59.9062
R3410 d<6>.n26 d<6>.t43 59.9062
R3411 d<6>.n27 d<6>.t118 59.9062
R3412 d<6>.n28 d<6>.t33 59.9062
R3413 d<6>.n29 d<6>.t15 59.9062
R3414 d<6>.n30 d<6>.t95 59.9062
R3415 d<6>.n31 d<6>.t79 59.9062
R3416 d<6>.n32 d<6>.t35 59.9062
R3417 d<6>.n33 d<6>.t17 59.9062
R3418 d<6>.n34 d<6>.t97 59.9062
R3419 d<6>.n35 d<6>.t54 59.9062
R3420 d<6>.n36 d<6>.t119 59.9062
R3421 d<6>.n37 d<6>.t104 59.9062
R3422 d<6>.n38 d<6>.t60 59.9062
R3423 d<6>.n39 d<6>.t10 59.9062
R3424 d<6>.n40 d<6>.t121 59.9062
R3425 d<6>.n41 d<6>.t106 59.9062
R3426 d<6>.n42 d<6>.t62 59.9062
R3427 d<6>.n43 d<6>.t14 59.9062
R3428 d<6>.n44 d<6>.t82 59.9062
R3429 d<6>.n45 d<6>.t37 59.9062
R3430 d<6>.n46 d<6>.t21 59.9062
R3431 d<6>.n47 d<6>.t5 59.9062
R3432 d<6>.n48 d<6>.t85 59.9062
R3433 d<6>.n49 d<6>.t41 59.9062
R3434 d<6>.n50 d<6>.t117 59.9062
R3435 d<6>.n51 d<6>.t92 59.9062
R3436 d<6>.n52 d<6>.t50 59.9062
R3437 d<6>.n53 d<6>.t126 59.9062
R3438 d<6>.n54 d<6>.t108 59.9062
R3439 d<6>.n55 d<6>.t65 59.9062
R3440 d<6>.n56 d<6>.t53 59.9062
R3441 d<6>.n57 d<6>.t2 59.9062
R3442 d<6>.n58 d<6>.t112 59.9062
R3443 d<6>.n59 d<6>.t26 59.9062
R3444 d<6>.n60 d<6>.t103 59.9062
R3445 d<6>.n61 d<6>.t88 59.9062
R3446 d<6>.n62 d<6>.t75 59.9062
R3447 d<6>.n63 d<6>.t31 59.9062
R3448 d<6> d<6>.n63 24.1005
R3449 hgu_cdac_8bit_array_3.drv<63:0>.n159 hgu_cdac_8bit_array_3.drv<63:0>.t101 41.4291
R3450 hgu_cdac_8bit_array_3.drv<63:0>.n159 hgu_cdac_8bit_array_3.drv<63:0>.t98 41.4291
R3451 hgu_cdac_8bit_array_3.drv<63:0>.n177 hgu_cdac_8bit_array_3.drv<63:0>.t112 41.4291
R3452 hgu_cdac_8bit_array_3.drv<63:0>.n177 hgu_cdac_8bit_array_3.drv<63:0>.t118 41.4291
R3453 hgu_cdac_8bit_array_3.drv<63:0>.n180 hgu_cdac_8bit_array_3.drv<63:0>.t7 41.4291
R3454 hgu_cdac_8bit_array_3.drv<63:0>.n180 hgu_cdac_8bit_array_3.drv<63:0>.t111 41.4291
R3455 hgu_cdac_8bit_array_3.drv<63:0>.n182 hgu_cdac_8bit_array_3.drv<63:0>.t1 41.4291
R3456 hgu_cdac_8bit_array_3.drv<63:0>.n182 hgu_cdac_8bit_array_3.drv<63:0>.t23 41.4291
R3457 hgu_cdac_8bit_array_3.drv<63:0>.n195 hgu_cdac_8bit_array_3.drv<63:0>.t5 41.4291
R3458 hgu_cdac_8bit_array_3.drv<63:0>.n195 hgu_cdac_8bit_array_3.drv<63:0>.t20 41.4291
R3459 hgu_cdac_8bit_array_3.drv<63:0>.n197 hgu_cdac_8bit_array_3.drv<63:0>.t95 41.4291
R3460 hgu_cdac_8bit_array_3.drv<63:0>.n197 hgu_cdac_8bit_array_3.drv<63:0>.t21 41.4291
R3461 hgu_cdac_8bit_array_3.drv<63:0>.n201 hgu_cdac_8bit_array_3.drv<63:0>.t125 41.4291
R3462 hgu_cdac_8bit_array_3.drv<63:0>.n201 hgu_cdac_8bit_array_3.drv<63:0>.t12 41.4291
R3463 hgu_cdac_8bit_array_3.drv<63:0>.n204 hgu_cdac_8bit_array_3.drv<63:0>.t9 41.4291
R3464 hgu_cdac_8bit_array_3.drv<63:0>.n204 hgu_cdac_8bit_array_3.drv<63:0>.t93 41.4291
R3465 hgu_cdac_8bit_array_3.drv<63:0>.n216 hgu_cdac_8bit_array_3.drv<63:0>.t123 41.4291
R3466 hgu_cdac_8bit_array_3.drv<63:0>.n216 hgu_cdac_8bit_array_3.drv<63:0>.t10 41.4291
R3467 hgu_cdac_8bit_array_3.drv<63:0>.n219 hgu_cdac_8bit_array_3.drv<63:0>.t8 41.4291
R3468 hgu_cdac_8bit_array_3.drv<63:0>.n219 hgu_cdac_8bit_array_3.drv<63:0>.t91 41.4291
R3469 hgu_cdac_8bit_array_3.drv<63:0>.n221 hgu_cdac_8bit_array_3.drv<63:0>.t22 41.4291
R3470 hgu_cdac_8bit_array_3.drv<63:0>.n221 hgu_cdac_8bit_array_3.drv<63:0>.t102 41.4291
R3471 hgu_cdac_8bit_array_3.drv<63:0>.n234 hgu_cdac_8bit_array_3.drv<63:0>.t107 41.4291
R3472 hgu_cdac_8bit_array_3.drv<63:0>.n234 hgu_cdac_8bit_array_3.drv<63:0>.t19 41.4291
R3473 hgu_cdac_8bit_array_3.drv<63:0>.n237 hgu_cdac_8bit_array_3.drv<63:0>.t99 41.4291
R3474 hgu_cdac_8bit_array_3.drv<63:0>.n237 hgu_cdac_8bit_array_3.drv<63:0>.t113 41.4291
R3475 hgu_cdac_8bit_array_3.drv<63:0>.n249 hgu_cdac_8bit_array_3.drv<63:0>.t105 41.4291
R3476 hgu_cdac_8bit_array_3.drv<63:0>.n249 hgu_cdac_8bit_array_3.drv<63:0>.t17 41.4291
R3477 hgu_cdac_8bit_array_3.drv<63:0>.n252 hgu_cdac_8bit_array_3.drv<63:0>.t90 41.4291
R3478 hgu_cdac_8bit_array_3.drv<63:0>.n252 hgu_cdac_8bit_array_3.drv<63:0>.t116 41.4291
R3479 hgu_cdac_8bit_array_3.drv<63:0>.n254 hgu_cdac_8bit_array_3.drv<63:0>.t120 41.4291
R3480 hgu_cdac_8bit_array_3.drv<63:0>.n254 hgu_cdac_8bit_array_3.drv<63:0>.t96 41.4291
R3481 hgu_cdac_8bit_array_3.drv<63:0>.n256 hgu_cdac_8bit_array_3.drv<63:0>.t109 41.4291
R3482 hgu_cdac_8bit_array_3.drv<63:0>.n256 hgu_cdac_8bit_array_3.drv<63:0>.t115 41.4291
R3483 hgu_cdac_8bit_array_3.drv<63:0>.n279 hgu_cdac_8bit_array_3.drv<63:0>.t119 41.4291
R3484 hgu_cdac_8bit_array_3.drv<63:0>.n279 hgu_cdac_8bit_array_3.drv<63:0>.t103 41.4291
R3485 hgu_cdac_8bit_array_3.drv<63:0>.n277 hgu_cdac_8bit_array_3.drv<63:0>.t16 41.4291
R3486 hgu_cdac_8bit_array_3.drv<63:0>.n277 hgu_cdac_8bit_array_3.drv<63:0>.t4 41.4291
R3487 hgu_cdac_8bit_array_3.drv<63:0>.n299 hgu_cdac_8bit_array_3.drv<63:0>.t100 41.4291
R3488 hgu_cdac_8bit_array_3.drv<63:0>.n299 hgu_cdac_8bit_array_3.drv<63:0>.t124 41.4291
R3489 hgu_cdac_8bit_array_3.drv<63:0>.n302 hgu_cdac_8bit_array_3.drv<63:0>.t15 41.4291
R3490 hgu_cdac_8bit_array_3.drv<63:0>.n302 hgu_cdac_8bit_array_3.drv<63:0>.t3 41.4291
R3491 hgu_cdac_8bit_array_3.drv<63:0>.n305 hgu_cdac_8bit_array_3.drv<63:0>.t25 41.4291
R3492 hgu_cdac_8bit_array_3.drv<63:0>.n305 hgu_cdac_8bit_array_3.drv<63:0>.t122 41.4291
R3493 hgu_cdac_8bit_array_3.drv<63:0>.n310 hgu_cdac_8bit_array_3.drv<63:0>.t14 41.4291
R3494 hgu_cdac_8bit_array_3.drv<63:0>.n310 hgu_cdac_8bit_array_3.drv<63:0>.t108 41.4291
R3495 hgu_cdac_8bit_array_3.drv<63:0>.n313 hgu_cdac_8bit_array_3.drv<63:0>.t114 41.4291
R3496 hgu_cdac_8bit_array_3.drv<63:0>.n313 hgu_cdac_8bit_array_3.drv<63:0>.t126 41.4291
R3497 hgu_cdac_8bit_array_3.drv<63:0>.n325 hgu_cdac_8bit_array_3.drv<63:0>.t13 41.4291
R3498 hgu_cdac_8bit_array_3.drv<63:0>.n325 hgu_cdac_8bit_array_3.drv<63:0>.t106 41.4291
R3499 hgu_cdac_8bit_array_3.drv<63:0>.n328 hgu_cdac_8bit_array_3.drv<63:0>.t18 41.4291
R3500 hgu_cdac_8bit_array_3.drv<63:0>.n328 hgu_cdac_8bit_array_3.drv<63:0>.t121 41.4291
R3501 hgu_cdac_8bit_array_3.drv<63:0>.n331 hgu_cdac_8bit_array_3.drv<63:0>.t6 41.4291
R3502 hgu_cdac_8bit_array_3.drv<63:0>.n331 hgu_cdac_8bit_array_3.drv<63:0>.t110 41.4291
R3503 hgu_cdac_8bit_array_3.drv<63:0>.n343 hgu_cdac_8bit_array_3.drv<63:0>.t2 41.4291
R3504 hgu_cdac_8bit_array_3.drv<63:0>.n343 hgu_cdac_8bit_array_3.drv<63:0>.t24 41.4291
R3505 hgu_cdac_8bit_array_3.drv<63:0>.n346 hgu_cdac_8bit_array_3.drv<63:0>.t104 41.4291
R3506 hgu_cdac_8bit_array_3.drv<63:0>.n346 hgu_cdac_8bit_array_3.drv<63:0>.t127 41.4291
R3507 hgu_cdac_8bit_array_3.drv<63:0>.n358 hgu_cdac_8bit_array_3.drv<63:0>.t0 41.4291
R3508 hgu_cdac_8bit_array_3.drv<63:0>.n358 hgu_cdac_8bit_array_3.drv<63:0>.t94 41.4291
R3509 hgu_cdac_8bit_array_3.drv<63:0>.n361 hgu_cdac_8bit_array_3.drv<63:0>.t117 41.4291
R3510 hgu_cdac_8bit_array_3.drv<63:0>.n361 hgu_cdac_8bit_array_3.drv<63:0>.t11 41.4291
R3511 hgu_cdac_8bit_array_3.drv<63:0>.n363 hgu_cdac_8bit_array_3.drv<63:0>.t97 41.4291
R3512 hgu_cdac_8bit_array_3.drv<63:0>.n363 hgu_cdac_8bit_array_3.drv<63:0>.t92 41.4291
R3513 hgu_cdac_8bit_array_3.drv<63:0>.n160 hgu_cdac_8bit_array_3.drv<63:0>.t73 34.0065
R3514 hgu_cdac_8bit_array_3.drv<63:0>.n160 hgu_cdac_8bit_array_3.drv<63:0>.t65 34.0065
R3515 hgu_cdac_8bit_array_3.drv<63:0>.n178 hgu_cdac_8bit_array_3.drv<63:0>.t28 34.0065
R3516 hgu_cdac_8bit_array_3.drv<63:0>.n178 hgu_cdac_8bit_array_3.drv<63:0>.t53 34.0065
R3517 hgu_cdac_8bit_array_3.drv<63:0>.n181 hgu_cdac_8bit_array_3.drv<63:0>.t79 34.0065
R3518 hgu_cdac_8bit_array_3.drv<63:0>.n181 hgu_cdac_8bit_array_3.drv<63:0>.t41 34.0065
R3519 hgu_cdac_8bit_array_3.drv<63:0>.n183 hgu_cdac_8bit_array_3.drv<63:0>.t49 34.0065
R3520 hgu_cdac_8bit_array_3.drv<63:0>.n183 hgu_cdac_8bit_array_3.drv<63:0>.t70 34.0065
R3521 hgu_cdac_8bit_array_3.drv<63:0>.n196 hgu_cdac_8bit_array_3.drv<63:0>.t77 34.0065
R3522 hgu_cdac_8bit_array_3.drv<63:0>.n196 hgu_cdac_8bit_array_3.drv<63:0>.t39 34.0065
R3523 hgu_cdac_8bit_array_3.drv<63:0>.n198 hgu_cdac_8bit_array_3.drv<63:0>.t62 34.0065
R3524 hgu_cdac_8bit_array_3.drv<63:0>.n198 hgu_cdac_8bit_array_3.drv<63:0>.t67 34.0065
R3525 hgu_cdac_8bit_array_3.drv<63:0>.n202 hgu_cdac_8bit_array_3.drv<63:0>.t36 34.0065
R3526 hgu_cdac_8bit_array_3.drv<63:0>.n202 hgu_cdac_8bit_array_3.drv<63:0>.t59 34.0065
R3527 hgu_cdac_8bit_array_3.drv<63:0>.n205 hgu_cdac_8bit_array_3.drv<63:0>.t81 34.0065
R3528 hgu_cdac_8bit_array_3.drv<63:0>.n205 hgu_cdac_8bit_array_3.drv<63:0>.t26 34.0065
R3529 hgu_cdac_8bit_array_3.drv<63:0>.n217 hgu_cdac_8bit_array_3.drv<63:0>.t34 34.0065
R3530 hgu_cdac_8bit_array_3.drv<63:0>.n217 hgu_cdac_8bit_array_3.drv<63:0>.t57 34.0065
R3531 hgu_cdac_8bit_array_3.drv<63:0>.n220 hgu_cdac_8bit_array_3.drv<63:0>.t80 34.0065
R3532 hgu_cdac_8bit_array_3.drv<63:0>.n220 hgu_cdac_8bit_array_3.drv<63:0>.t88 34.0065
R3533 hgu_cdac_8bit_array_3.drv<63:0>.n222 hgu_cdac_8bit_array_3.drv<63:0>.t68 34.0065
R3534 hgu_cdac_8bit_array_3.drv<63:0>.n222 hgu_cdac_8bit_array_3.drv<63:0>.t74 34.0065
R3535 hgu_cdac_8bit_array_3.drv<63:0>.n235 hgu_cdac_8bit_array_3.drv<63:0>.t84 34.0065
R3536 hgu_cdac_8bit_array_3.drv<63:0>.n235 hgu_cdac_8bit_array_3.drv<63:0>.t46 34.0065
R3537 hgu_cdac_8bit_array_3.drv<63:0>.n238 hgu_cdac_8bit_array_3.drv<63:0>.t66 34.0065
R3538 hgu_cdac_8bit_array_3.drv<63:0>.n238 hgu_cdac_8bit_array_3.drv<63:0>.t29 34.0065
R3539 hgu_cdac_8bit_array_3.drv<63:0>.n250 hgu_cdac_8bit_array_3.drv<63:0>.t82 34.0065
R3540 hgu_cdac_8bit_array_3.drv<63:0>.n250 hgu_cdac_8bit_array_3.drv<63:0>.t44 34.0065
R3541 hgu_cdac_8bit_array_3.drv<63:0>.n253 hgu_cdac_8bit_array_3.drv<63:0>.t87 34.0065
R3542 hgu_cdac_8bit_array_3.drv<63:0>.n253 hgu_cdac_8bit_array_3.drv<63:0>.t32 34.0065
R3543 hgu_cdac_8bit_array_3.drv<63:0>.n255 hgu_cdac_8bit_array_3.drv<63:0>.t55 34.0065
R3544 hgu_cdac_8bit_array_3.drv<63:0>.n255 hgu_cdac_8bit_array_3.drv<63:0>.t63 34.0065
R3545 hgu_cdac_8bit_array_3.drv<63:0>.n257 hgu_cdac_8bit_array_3.drv<63:0>.t86 34.0065
R3546 hgu_cdac_8bit_array_3.drv<63:0>.n257 hgu_cdac_8bit_array_3.drv<63:0>.t31 34.0065
R3547 hgu_cdac_8bit_array_3.drv<63:0>.n280 hgu_cdac_8bit_array_3.drv<63:0>.t54 34.0065
R3548 hgu_cdac_8bit_array_3.drv<63:0>.n280 hgu_cdac_8bit_array_3.drv<63:0>.t75 34.0065
R3549 hgu_cdac_8bit_array_3.drv<63:0>.n278 hgu_cdac_8bit_array_3.drv<63:0>.t43 34.0065
R3550 hgu_cdac_8bit_array_3.drv<63:0>.n278 hgu_cdac_8bit_array_3.drv<63:0>.t51 34.0065
R3551 hgu_cdac_8bit_array_3.drv<63:0>.n300 hgu_cdac_8bit_array_3.drv<63:0>.t72 34.0065
R3552 hgu_cdac_8bit_array_3.drv<63:0>.n300 hgu_cdac_8bit_array_3.drv<63:0>.t35 34.0065
R3553 hgu_cdac_8bit_array_3.drv<63:0>.n303 hgu_cdac_8bit_array_3.drv<63:0>.t42 34.0065
R3554 hgu_cdac_8bit_array_3.drv<63:0>.n303 hgu_cdac_8bit_array_3.drv<63:0>.t50 34.0065
R3555 hgu_cdac_8bit_array_3.drv<63:0>.n306 hgu_cdac_8bit_array_3.drv<63:0>.t71 34.0065
R3556 hgu_cdac_8bit_array_3.drv<63:0>.n306 hgu_cdac_8bit_array_3.drv<63:0>.t33 34.0065
R3557 hgu_cdac_8bit_array_3.drv<63:0>.n311 hgu_cdac_8bit_array_3.drv<63:0>.t61 34.0065
R3558 hgu_cdac_8bit_array_3.drv<63:0>.n311 hgu_cdac_8bit_array_3.drv<63:0>.t85 34.0065
R3559 hgu_cdac_8bit_array_3.drv<63:0>.n314 hgu_cdac_8bit_array_3.drv<63:0>.t30 34.0065
R3560 hgu_cdac_8bit_array_3.drv<63:0>.n314 hgu_cdac_8bit_array_3.drv<63:0>.t37 34.0065
R3561 hgu_cdac_8bit_array_3.drv<63:0>.n326 hgu_cdac_8bit_array_3.drv<63:0>.t60 34.0065
R3562 hgu_cdac_8bit_array_3.drv<63:0>.n326 hgu_cdac_8bit_array_3.drv<63:0>.t83 34.0065
R3563 hgu_cdac_8bit_array_3.drv<63:0>.n329 hgu_cdac_8bit_array_3.drv<63:0>.t45 34.0065
R3564 hgu_cdac_8bit_array_3.drv<63:0>.n329 hgu_cdac_8bit_array_3.drv<63:0>.t56 34.0065
R3565 hgu_cdac_8bit_array_3.drv<63:0>.n332 hgu_cdac_8bit_array_3.drv<63:0>.t78 34.0065
R3566 hgu_cdac_8bit_array_3.drv<63:0>.n332 hgu_cdac_8bit_array_3.drv<63:0>.t40 34.0065
R3567 hgu_cdac_8bit_array_3.drv<63:0>.n344 hgu_cdac_8bit_array_3.drv<63:0>.t48 34.0065
R3568 hgu_cdac_8bit_array_3.drv<63:0>.n344 hgu_cdac_8bit_array_3.drv<63:0>.t69 34.0065
R3569 hgu_cdac_8bit_array_3.drv<63:0>.n347 hgu_cdac_8bit_array_3.drv<63:0>.t76 34.0065
R3570 hgu_cdac_8bit_array_3.drv<63:0>.n347 hgu_cdac_8bit_array_3.drv<63:0>.t38 34.0065
R3571 hgu_cdac_8bit_array_3.drv<63:0>.n359 hgu_cdac_8bit_array_3.drv<63:0>.t47 34.0065
R3572 hgu_cdac_8bit_array_3.drv<63:0>.n359 hgu_cdac_8bit_array_3.drv<63:0>.t27 34.0065
R3573 hgu_cdac_8bit_array_3.drv<63:0>.n367 hgu_cdac_8bit_array_3.drv<63:0>.t52 34.0065
R3574 hgu_cdac_8bit_array_3.drv<63:0>.n367 hgu_cdac_8bit_array_3.drv<63:0>.t58 34.0065
R3575 hgu_cdac_8bit_array_3.drv<63:0>.n364 hgu_cdac_8bit_array_3.drv<63:0>.t64 34.0065
R3576 hgu_cdac_8bit_array_3.drv<63:0>.n364 hgu_cdac_8bit_array_3.drv<63:0>.t89 34.0065
R3577 hgu_cdac_8bit_array_3.drv<63:0>.n169 hgu_cdac_8bit_array_3.drv<63:0>.n161 11.3459
R3578 hgu_cdac_8bit_array_3.drv<63:0>.n291 hgu_cdac_8bit_array_3.drv<63:0>.n283 11.0733
R3579 hgu_cdac_8bit_array_3.drv<63:0>.n187 hgu_cdac_8bit_array_3.drv<63:0>.n186 10.7039
R3580 hgu_cdac_8bit_array_3.drv<63:0>.n309 hgu_cdac_8bit_array_3.drv<63:0>.n308 10.7039
R3581 hgu_cdac_8bit_array_3.drv<63:0>.n200 hgu_cdac_8bit_array_3.drv<63:0>.n0 10.7015
R3582 hgu_cdac_8bit_array_3.drv<63:0>.n215 hgu_cdac_8bit_array_3.drv<63:0>.n207 10.7015
R3583 hgu_cdac_8bit_array_3.drv<63:0>.n248 hgu_cdac_8bit_array_3.drv<63:0>.n240 10.7015
R3584 hgu_cdac_8bit_array_3.drv<63:0>.n269 hgu_cdac_8bit_array_3.drv<63:0>.n261 10.7015
R3585 hgu_cdac_8bit_array_3.drv<63:0>.n324 hgu_cdac_8bit_array_3.drv<63:0>.n316 10.7015
R3586 hgu_cdac_8bit_array_3.drv<63:0>.n342 hgu_cdac_8bit_array_3.drv<63:0>.n334 10.7015
R3587 hgu_cdac_8bit_array_3.drv<63:0>.n372 hgu_cdac_8bit_array_3.drv<63:0>.n368 10.6992
R3588 hgu_cdac_8bit_array_3.drv<63:0>.n357 hgu_cdac_8bit_array_3.drv<63:0>.n349 10.6961
R3589 hgu_cdac_8bit_array_3.drv<63:0>.n233 hgu_cdac_8bit_array_3.drv<63:0>.n225 10.6886
R3590 hgu_cdac_8bit_array_3.drv<63:0>.n366 hgu_cdac_8bit_array_3.drv<63:0>.n365 1.96171
R3591 hgu_cdac_8bit_array_3.drv<63:0>.n334 hgu_cdac_8bit_array_3.drv<63:0>.n333 1.6061
R3592 hgu_cdac_8bit_array_3.drv<63:0>.n349 hgu_cdac_8bit_array_3.drv<63:0>.n348 1.32066
R3593 hgu_cdac_8bit_array_3.drv<63:0>.n308 hgu_cdac_8bit_array_3.drv<63:0>.n307 1.313
R3594 hgu_cdac_8bit_array_3.drv<63:0>.n282 hgu_cdac_8bit_array_3.drv<63:0>.n281 0.9906
R3595 hgu_cdac_8bit_array_3.drv<63:0>.n224 hgu_cdac_8bit_array_3.drv<63:0>.n223 0.990089
R3596 hgu_cdac_8bit_array_3.drv<63:0>.n185 hgu_cdac_8bit_array_3.drv<63:0>.n184 0.957397
R3597 hgu_cdac_8bit_array_3.drv<63:0>.n260 hgu_cdac_8bit_array_3.drv<63:0>.n259 0.957397
R3598 hgu_cdac_8bit_array_3.drv<63:0>.n259 hgu_cdac_8bit_array_3.drv<63:0>.n258 0.957397
R3599 hgu_cdac_8bit_array_3.drv<63:0>.n304 hgu_cdac_8bit_array_3.drv<63:0>.n301 0.957397
R3600 hgu_cdac_8bit_array_3.drv<63:0>.n330 hgu_cdac_8bit_array_3.drv<63:0>.n327 0.957397
R3601 hgu_cdac_8bit_array_3.drv<63:0>.n0 hgu_cdac_8bit_array_3.drv<63:0>.n199 0.950931
R3602 hgu_cdac_8bit_array_3.drv<63:0>.n362 hgu_cdac_8bit_array_3.drv<63:0>.n360 0.944465
R3603 hgu_cdac_8bit_array_3.drv<63:0>.n316 hgu_cdac_8bit_array_3.drv<63:0>.n312 0.894897
R3604 hgu_cdac_8bit_array_3.drv<63:0>.n240 hgu_cdac_8bit_array_3.drv<63:0>.n239 0.830241
R3605 hgu_cdac_8bit_array_3.drv<63:0>.n225 hgu_cdac_8bit_array_3.drv<63:0>.n218 0.751694
R3606 hgu_cdac_8bit_array_3.drv<63:0>.n349 hgu_cdac_8bit_array_3.drv<63:0>.n345 0.605142
R3607 hgu_cdac_8bit_array_3.drv<63:0>.n365 hgu_cdac_8bit_array_3.drv<63:0>.n364 0.592444
R3608 hgu_cdac_8bit_array_3.drv<63:0>.n186 hgu_cdac_8bit_array_3.drv<63:0>.n179 0.55869
R3609 hgu_cdac_8bit_array_3.drv<63:0>.n161 hgu_cdac_8bit_array_3.drv<63:0>.n160 0.558205
R3610 hgu_cdac_8bit_array_3.drv<63:0>.n179 hgu_cdac_8bit_array_3.drv<63:0>.n178 0.558205
R3611 hgu_cdac_8bit_array_3.drv<63:0>.n185 hgu_cdac_8bit_array_3.drv<63:0>.n181 0.558205
R3612 hgu_cdac_8bit_array_3.drv<63:0>.n184 hgu_cdac_8bit_array_3.drv<63:0>.n183 0.558205
R3613 hgu_cdac_8bit_array_3.drv<63:0>.n199 hgu_cdac_8bit_array_3.drv<63:0>.n198 0.558205
R3614 hgu_cdac_8bit_array_3.drv<63:0>.n203 hgu_cdac_8bit_array_3.drv<63:0>.n202 0.558205
R3615 hgu_cdac_8bit_array_3.drv<63:0>.n206 hgu_cdac_8bit_array_3.drv<63:0>.n205 0.558205
R3616 hgu_cdac_8bit_array_3.drv<63:0>.n218 hgu_cdac_8bit_array_3.drv<63:0>.n217 0.558205
R3617 hgu_cdac_8bit_array_3.drv<63:0>.n223 hgu_cdac_8bit_array_3.drv<63:0>.n222 0.558205
R3618 hgu_cdac_8bit_array_3.drv<63:0>.n239 hgu_cdac_8bit_array_3.drv<63:0>.n238 0.558205
R3619 hgu_cdac_8bit_array_3.drv<63:0>.n251 hgu_cdac_8bit_array_3.drv<63:0>.n250 0.558205
R3620 hgu_cdac_8bit_array_3.drv<63:0>.n260 hgu_cdac_8bit_array_3.drv<63:0>.n253 0.558205
R3621 hgu_cdac_8bit_array_3.drv<63:0>.n259 hgu_cdac_8bit_array_3.drv<63:0>.n255 0.558205
R3622 hgu_cdac_8bit_array_3.drv<63:0>.n258 hgu_cdac_8bit_array_3.drv<63:0>.n257 0.558205
R3623 hgu_cdac_8bit_array_3.drv<63:0>.n281 hgu_cdac_8bit_array_3.drv<63:0>.n280 0.558205
R3624 hgu_cdac_8bit_array_3.drv<63:0>.n301 hgu_cdac_8bit_array_3.drv<63:0>.n300 0.558205
R3625 hgu_cdac_8bit_array_3.drv<63:0>.n304 hgu_cdac_8bit_array_3.drv<63:0>.n303 0.558205
R3626 hgu_cdac_8bit_array_3.drv<63:0>.n307 hgu_cdac_8bit_array_3.drv<63:0>.n306 0.558205
R3627 hgu_cdac_8bit_array_3.drv<63:0>.n312 hgu_cdac_8bit_array_3.drv<63:0>.n311 0.558205
R3628 hgu_cdac_8bit_array_3.drv<63:0>.n327 hgu_cdac_8bit_array_3.drv<63:0>.n326 0.558205
R3629 hgu_cdac_8bit_array_3.drv<63:0>.n330 hgu_cdac_8bit_array_3.drv<63:0>.n329 0.558205
R3630 hgu_cdac_8bit_array_3.drv<63:0>.n333 hgu_cdac_8bit_array_3.drv<63:0>.n332 0.558205
R3631 hgu_cdac_8bit_array_3.drv<63:0>.n345 hgu_cdac_8bit_array_3.drv<63:0>.n344 0.558205
R3632 hgu_cdac_8bit_array_3.drv<63:0>.n348 hgu_cdac_8bit_array_3.drv<63:0>.n347 0.558205
R3633 hgu_cdac_8bit_array_3.drv<63:0>.n360 hgu_cdac_8bit_array_3.drv<63:0>.n359 0.558205
R3634 hgu_cdac_8bit_array_3.drv<63:0>.n207 hgu_cdac_8bit_array_3.drv<63:0>.n206 0.541448
R3635 hgu_cdac_8bit_array_3.drv<63:0>.n308 hgu_cdac_8bit_array_3.drv<63:0>.n304 0.489724
R3636 hgu_cdac_8bit_array_3.drv<63:0>.n368 hgu_cdac_8bit_array_3.drv<63:0>.n367 0.436881
R3637 hgu_cdac_8bit_array_3.drv<63:0>.n261 hgu_cdac_8bit_array_3.drv<63:0>.n260 0.425069
R3638 hgu_cdac_8bit_array_3.drv<63:0>.n261 hgu_cdac_8bit_array_3.drv<63:0>.n251 0.381966
R3639 hgu_cdac_8bit_array_3.drv<63:0>.n0 hgu_cdac_8bit_array_3.drv<63:0>.n196 0.378057
R3640 hgu_cdac_8bit_array_3.drv<63:0>.n236 hgu_cdac_8bit_array_3.drv<63:0>.n235 0.378057
R3641 hgu_cdac_8bit_array_3.drv<63:0>.n282 hgu_cdac_8bit_array_3.drv<63:0>.n278 0.378057
R3642 hgu_cdac_8bit_array_3.drv<63:0>.n315 hgu_cdac_8bit_array_3.drv<63:0>.n314 0.378057
R3643 hgu_cdac_8bit_array_3.drv<63:0>.n224 hgu_cdac_8bit_array_3.drv<63:0>.n220 0.374381
R3644 hgu_cdac_8bit_array_3.drv<63:0>.n32 hgu_cdac_8bit_array_3.drv<63:0> 0.338468
R3645 hgu_cdac_8bit_array_3.drv<63:0>.n36 hgu_cdac_8bit_array_3.drv<63:0>.n31 0.330451
R3646 hgu_cdac_8bit_array_3.drv<63:0>.n45 hgu_cdac_8bit_array_3.drv<63:0>.n28 0.330451
R3647 hgu_cdac_8bit_array_3.drv<63:0>.n54 hgu_cdac_8bit_array_3.drv<63:0>.n21 0.330451
R3648 hgu_cdac_8bit_array_3.drv<63:0>.n63 hgu_cdac_8bit_array_3.drv<63:0>.n14 0.330451
R3649 hgu_cdac_8bit_array_3.drv<63:0>.n72 hgu_cdac_8bit_array_3.drv<63:0>.n7 0.330451
R3650 hgu_cdac_8bit_array_3.drv<63:0>.n594 hgu_cdac_8bit_array_3.drv<63:0>.n88 0.330451
R3651 hgu_cdac_8bit_array_3.drv<63:0>.n585 hgu_cdac_8bit_array_3.drv<63:0>.n95 0.330451
R3652 hgu_cdac_8bit_array_3.drv<63:0>.n576 hgu_cdac_8bit_array_3.drv<63:0>.n102 0.330451
R3653 hgu_cdac_8bit_array_3.drv<63:0>.n567 hgu_cdac_8bit_array_3.drv<63:0>.n109 0.330451
R3654 hgu_cdac_8bit_array_3.drv<63:0>.n558 hgu_cdac_8bit_array_3.drv<63:0>.n116 0.330451
R3655 hgu_cdac_8bit_array_3.drv<63:0>.n549 hgu_cdac_8bit_array_3.drv<63:0>.n123 0.330451
R3656 hgu_cdac_8bit_array_3.drv<63:0>.n540 hgu_cdac_8bit_array_3.drv<63:0>.n130 0.330451
R3657 hgu_cdac_8bit_array_3.drv<63:0>.n531 hgu_cdac_8bit_array_3.drv<63:0>.n137 0.330451
R3658 hgu_cdac_8bit_array_3.drv<63:0>.n522 hgu_cdac_8bit_array_3.drv<63:0>.n144 0.330451
R3659 hgu_cdac_8bit_array_3.drv<63:0>.n513 hgu_cdac_8bit_array_3.drv<63:0>.n151 0.330451
R3660 hgu_cdac_8bit_array_3.drv<63:0>.n504 hgu_cdac_8bit_array_3.drv<63:0>.n158 0.330451
R3661 hgu_cdac_8bit_array_3.drv<63:0>.n431 hgu_cdac_8bit_array_3.drv<63:0>.n276 0.330451
R3662 hgu_cdac_8bit_array_3.drv<63:0>.n374 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3663 hgu_cdac_8bit_array_3.drv<63:0>.n383 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3664 hgu_cdac_8bit_array_3.drv<63:0>.n392 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3665 hgu_cdac_8bit_array_3.drv<63:0>.n401 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3666 hgu_cdac_8bit_array_3.drv<63:0>.n410 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3667 hgu_cdac_8bit_array_3.drv<63:0>.n419 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3668 hgu_cdac_8bit_array_3.drv<63:0>.n428 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3669 hgu_cdac_8bit_array_3.drv<63:0>.n437 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3670 hgu_cdac_8bit_array_3.drv<63:0>.n446 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3671 hgu_cdac_8bit_array_3.drv<63:0>.n455 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3672 hgu_cdac_8bit_array_3.drv<63:0>.n464 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3673 hgu_cdac_8bit_array_3.drv<63:0>.n473 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3674 hgu_cdac_8bit_array_3.drv<63:0>.n482 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3675 hgu_cdac_8bit_array_3.drv<63:0>.n491 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3676 hgu_cdac_8bit_array_3.drv<63:0>.n500 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3677 hgu_cdac_8bit_array_3.drv<63:0>.n510 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3678 hgu_cdac_8bit_array_3.drv<63:0>.n519 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3679 hgu_cdac_8bit_array_3.drv<63:0>.n528 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3680 hgu_cdac_8bit_array_3.drv<63:0>.n537 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3681 hgu_cdac_8bit_array_3.drv<63:0>.n546 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3682 hgu_cdac_8bit_array_3.drv<63:0>.n555 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3683 hgu_cdac_8bit_array_3.drv<63:0>.n564 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3684 hgu_cdac_8bit_array_3.drv<63:0>.n573 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3685 hgu_cdac_8bit_array_3.drv<63:0>.n582 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3686 hgu_cdac_8bit_array_3.drv<63:0>.n591 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3687 hgu_cdac_8bit_array_3.drv<63:0>.n600 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3688 hgu_cdac_8bit_array_3.drv<63:0>.n75 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3689 hgu_cdac_8bit_array_3.drv<63:0>.n66 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3690 hgu_cdac_8bit_array_3.drv<63:0>.n57 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3691 hgu_cdac_8bit_array_3.drv<63:0>.n48 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3692 hgu_cdac_8bit_array_3.drv<63:0>.n39 hgu_cdac_8bit_array_3.drv<63:0> 0.321667
R3693 hgu_cdac_8bit_array_3.drv<63:0>.n373 hgu_cdac_8bit_array_3.drv<63:0> 0.313448
R3694 hgu_cdac_8bit_array_3.drv<63:0>.n161 hgu_cdac_8bit_array_3.drv<63:0>.n159 0.300856
R3695 hgu_cdac_8bit_array_3.drv<63:0>.n179 hgu_cdac_8bit_array_3.drv<63:0>.n177 0.300856
R3696 hgu_cdac_8bit_array_3.drv<63:0>.n185 hgu_cdac_8bit_array_3.drv<63:0>.n180 0.300856
R3697 hgu_cdac_8bit_array_3.drv<63:0>.n184 hgu_cdac_8bit_array_3.drv<63:0>.n182 0.300856
R3698 hgu_cdac_8bit_array_3.drv<63:0>.n199 hgu_cdac_8bit_array_3.drv<63:0>.n197 0.300856
R3699 hgu_cdac_8bit_array_3.drv<63:0>.n203 hgu_cdac_8bit_array_3.drv<63:0>.n201 0.300856
R3700 hgu_cdac_8bit_array_3.drv<63:0>.n206 hgu_cdac_8bit_array_3.drv<63:0>.n204 0.300856
R3701 hgu_cdac_8bit_array_3.drv<63:0>.n218 hgu_cdac_8bit_array_3.drv<63:0>.n216 0.300856
R3702 hgu_cdac_8bit_array_3.drv<63:0>.n223 hgu_cdac_8bit_array_3.drv<63:0>.n221 0.300856
R3703 hgu_cdac_8bit_array_3.drv<63:0>.n239 hgu_cdac_8bit_array_3.drv<63:0>.n237 0.300856
R3704 hgu_cdac_8bit_array_3.drv<63:0>.n251 hgu_cdac_8bit_array_3.drv<63:0>.n249 0.300856
R3705 hgu_cdac_8bit_array_3.drv<63:0>.n260 hgu_cdac_8bit_array_3.drv<63:0>.n252 0.300856
R3706 hgu_cdac_8bit_array_3.drv<63:0>.n259 hgu_cdac_8bit_array_3.drv<63:0>.n254 0.300856
R3707 hgu_cdac_8bit_array_3.drv<63:0>.n258 hgu_cdac_8bit_array_3.drv<63:0>.n256 0.300856
R3708 hgu_cdac_8bit_array_3.drv<63:0>.n281 hgu_cdac_8bit_array_3.drv<63:0>.n279 0.300856
R3709 hgu_cdac_8bit_array_3.drv<63:0>.n301 hgu_cdac_8bit_array_3.drv<63:0>.n299 0.300856
R3710 hgu_cdac_8bit_array_3.drv<63:0>.n304 hgu_cdac_8bit_array_3.drv<63:0>.n302 0.300856
R3711 hgu_cdac_8bit_array_3.drv<63:0>.n307 hgu_cdac_8bit_array_3.drv<63:0>.n305 0.300856
R3712 hgu_cdac_8bit_array_3.drv<63:0>.n312 hgu_cdac_8bit_array_3.drv<63:0>.n310 0.300856
R3713 hgu_cdac_8bit_array_3.drv<63:0>.n327 hgu_cdac_8bit_array_3.drv<63:0>.n325 0.300856
R3714 hgu_cdac_8bit_array_3.drv<63:0>.n330 hgu_cdac_8bit_array_3.drv<63:0>.n328 0.300856
R3715 hgu_cdac_8bit_array_3.drv<63:0>.n333 hgu_cdac_8bit_array_3.drv<63:0>.n331 0.300856
R3716 hgu_cdac_8bit_array_3.drv<63:0>.n345 hgu_cdac_8bit_array_3.drv<63:0>.n343 0.300856
R3717 hgu_cdac_8bit_array_3.drv<63:0>.n348 hgu_cdac_8bit_array_3.drv<63:0>.n346 0.300856
R3718 hgu_cdac_8bit_array_3.drv<63:0>.n360 hgu_cdac_8bit_array_3.drv<63:0>.n358 0.300856
R3719 hgu_cdac_8bit_array_3.drv<63:0>.n365 hgu_cdac_8bit_array_3.drv<63:0>.n363 0.300856
R3720 hgu_cdac_8bit_array_3.drv<63:0>.n33 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3721 hgu_cdac_8bit_array_3.drv<63:0>.n42 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3722 hgu_cdac_8bit_array_3.drv<63:0>.n51 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3723 hgu_cdac_8bit_array_3.drv<63:0>.n60 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3724 hgu_cdac_8bit_array_3.drv<63:0>.n69 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3725 hgu_cdac_8bit_array_3.drv<63:0>.n78 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3726 hgu_cdac_8bit_array_3.drv<63:0>.n597 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3727 hgu_cdac_8bit_array_3.drv<63:0>.n588 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3728 hgu_cdac_8bit_array_3.drv<63:0>.n579 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3729 hgu_cdac_8bit_array_3.drv<63:0>.n570 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3730 hgu_cdac_8bit_array_3.drv<63:0>.n561 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3731 hgu_cdac_8bit_array_3.drv<63:0>.n552 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3732 hgu_cdac_8bit_array_3.drv<63:0>.n543 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3733 hgu_cdac_8bit_array_3.drv<63:0>.n534 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3734 hgu_cdac_8bit_array_3.drv<63:0>.n525 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3735 hgu_cdac_8bit_array_3.drv<63:0>.n516 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3736 hgu_cdac_8bit_array_3.drv<63:0>.n507 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3737 hgu_cdac_8bit_array_3.drv<63:0>.n497 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3738 hgu_cdac_8bit_array_3.drv<63:0>.n488 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3739 hgu_cdac_8bit_array_3.drv<63:0>.n479 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3740 hgu_cdac_8bit_array_3.drv<63:0>.n470 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3741 hgu_cdac_8bit_array_3.drv<63:0>.n461 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3742 hgu_cdac_8bit_array_3.drv<63:0>.n452 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3743 hgu_cdac_8bit_array_3.drv<63:0>.n443 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3744 hgu_cdac_8bit_array_3.drv<63:0>.n434 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3745 hgu_cdac_8bit_array_3.drv<63:0>.n425 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3746 hgu_cdac_8bit_array_3.drv<63:0>.n416 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3747 hgu_cdac_8bit_array_3.drv<63:0>.n407 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3748 hgu_cdac_8bit_array_3.drv<63:0>.n398 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3749 hgu_cdac_8bit_array_3.drv<63:0>.n389 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3750 hgu_cdac_8bit_array_3.drv<63:0>.n380 hgu_cdac_8bit_array_3.drv<63:0> 0.2966
R3751 hgu_cdac_8bit_array_3.drv<63:0>.n362 hgu_cdac_8bit_array_3.drv<63:0>.n361 0.275005
R3752 hgu_cdac_8bit_array_3.drv<63:0>.n207 hgu_cdac_8bit_array_3.drv<63:0>.n203 0.265586
R3753 hgu_cdac_8bit_array_3.drv<63:0>.n186 hgu_cdac_8bit_array_3.drv<63:0>.n185 0.248345
R3754 hgu_cdac_8bit_array_3.drv<63:0>.n0 hgu_cdac_8bit_array_3.drv<63:0>.n195 0.247662
R3755 hgu_cdac_8bit_array_3.drv<63:0>.n224 hgu_cdac_8bit_array_3.drv<63:0>.n219 0.245708
R3756 hgu_cdac_8bit_array_3.drv<63:0>.n236 hgu_cdac_8bit_array_3.drv<63:0>.n234 0.245708
R3757 hgu_cdac_8bit_array_3.drv<63:0>.n282 hgu_cdac_8bit_array_3.drv<63:0>.n277 0.245708
R3758 hgu_cdac_8bit_array_3.drv<63:0>.n315 hgu_cdac_8bit_array_3.drv<63:0>.n313 0.245708
R3759 hgu_cdac_8bit_array_3.drv<63:0>.n334 hgu_cdac_8bit_array_3.drv<63:0>.n330 0.196621
R3760 hgu_cdac_8bit_array_3.drv<63:0>.n494 hgu_cdac_8bit_array_3.drv<63:0>.n169 0.182836
R3761 hgu_cdac_8bit_array_3.drv<63:0>.n485 hgu_cdac_8bit_array_3.drv<63:0>.n187 0.182836
R3762 hgu_cdac_8bit_array_3.drv<63:0>.n476 hgu_cdac_8bit_array_3.drv<63:0>.n200 0.182836
R3763 hgu_cdac_8bit_array_3.drv<63:0>.n467 hgu_cdac_8bit_array_3.drv<63:0>.n215 0.182836
R3764 hgu_cdac_8bit_array_3.drv<63:0>.n458 hgu_cdac_8bit_array_3.drv<63:0>.n233 0.182836
R3765 hgu_cdac_8bit_array_3.drv<63:0>.n449 hgu_cdac_8bit_array_3.drv<63:0>.n248 0.182836
R3766 hgu_cdac_8bit_array_3.drv<63:0>.n440 hgu_cdac_8bit_array_3.drv<63:0>.n269 0.182836
R3767 hgu_cdac_8bit_array_3.drv<63:0>.n422 hgu_cdac_8bit_array_3.drv<63:0>.n291 0.182836
R3768 hgu_cdac_8bit_array_3.drv<63:0>.n413 hgu_cdac_8bit_array_3.drv<63:0>.n309 0.182836
R3769 hgu_cdac_8bit_array_3.drv<63:0>.n404 hgu_cdac_8bit_array_3.drv<63:0>.n324 0.182836
R3770 hgu_cdac_8bit_array_3.drv<63:0>.n395 hgu_cdac_8bit_array_3.drv<63:0>.n342 0.182836
R3771 hgu_cdac_8bit_array_3.drv<63:0>.n386 hgu_cdac_8bit_array_3.drv<63:0>.n357 0.182836
R3772 hgu_cdac_8bit_array_3.drv<63:0>.n377 hgu_cdac_8bit_array_3.drv<63:0>.n372 0.182836
R3773 hgu_cdac_8bit_array_3.drv<63:0>.n169 hgu_cdac_8bit_array_3.drv<63:0>.n168 0.149114
R3774 hgu_cdac_8bit_array_3.drv<63:0>.n187 hgu_cdac_8bit_array_3.drv<63:0>.n176 0.149114
R3775 hgu_cdac_8bit_array_3.drv<63:0>.n200 hgu_cdac_8bit_array_3.drv<63:0>.n194 0.149114
R3776 hgu_cdac_8bit_array_3.drv<63:0>.n215 hgu_cdac_8bit_array_3.drv<63:0>.n214 0.149114
R3777 hgu_cdac_8bit_array_3.drv<63:0>.n233 hgu_cdac_8bit_array_3.drv<63:0>.n232 0.149114
R3778 hgu_cdac_8bit_array_3.drv<63:0>.n248 hgu_cdac_8bit_array_3.drv<63:0>.n247 0.149114
R3779 hgu_cdac_8bit_array_3.drv<63:0>.n269 hgu_cdac_8bit_array_3.drv<63:0>.n268 0.149114
R3780 hgu_cdac_8bit_array_3.drv<63:0>.n291 hgu_cdac_8bit_array_3.drv<63:0>.n290 0.149114
R3781 hgu_cdac_8bit_array_3.drv<63:0>.n309 hgu_cdac_8bit_array_3.drv<63:0>.n298 0.149114
R3782 hgu_cdac_8bit_array_3.drv<63:0>.n324 hgu_cdac_8bit_array_3.drv<63:0>.n323 0.149114
R3783 hgu_cdac_8bit_array_3.drv<63:0>.n342 hgu_cdac_8bit_array_3.drv<63:0>.n341 0.149114
R3784 hgu_cdac_8bit_array_3.drv<63:0>.n357 hgu_cdac_8bit_array_3.drv<63:0>.n356 0.149114
R3785 hgu_cdac_8bit_array_3.drv<63:0>.n372 hgu_cdac_8bit_array_3.drv<63:0>.n371 0.149114
R3786 hgu_cdac_8bit_array_3.drv<63:0>.n283 hgu_cdac_8bit_array_3.drv<63:0>.n282 0.09425
R3787 hgu_cdac_8bit_array_3.drv<63:0>.n225 hgu_cdac_8bit_array_3.drv<63:0>.n224 0.0908846
R3788 hgu_cdac_8bit_array_3.drv<63:0>.n36 hgu_cdac_8bit_array_3.drv<63:0>.n35 0.0716912
R3789 hgu_cdac_8bit_array_3.drv<63:0>.n37 hgu_cdac_8bit_array_3.drv<63:0>.n36 0.0716912
R3790 hgu_cdac_8bit_array_3.drv<63:0>.n45 hgu_cdac_8bit_array_3.drv<63:0>.n44 0.0716912
R3791 hgu_cdac_8bit_array_3.drv<63:0>.n46 hgu_cdac_8bit_array_3.drv<63:0>.n45 0.0716912
R3792 hgu_cdac_8bit_array_3.drv<63:0>.n54 hgu_cdac_8bit_array_3.drv<63:0>.n53 0.0716912
R3793 hgu_cdac_8bit_array_3.drv<63:0>.n55 hgu_cdac_8bit_array_3.drv<63:0>.n54 0.0716912
R3794 hgu_cdac_8bit_array_3.drv<63:0>.n63 hgu_cdac_8bit_array_3.drv<63:0>.n62 0.0716912
R3795 hgu_cdac_8bit_array_3.drv<63:0>.n64 hgu_cdac_8bit_array_3.drv<63:0>.n63 0.0716912
R3796 hgu_cdac_8bit_array_3.drv<63:0>.n72 hgu_cdac_8bit_array_3.drv<63:0>.n71 0.0716912
R3797 hgu_cdac_8bit_array_3.drv<63:0>.n73 hgu_cdac_8bit_array_3.drv<63:0>.n72 0.0716912
R3798 hgu_cdac_8bit_array_3.drv<63:0>.n81 hgu_cdac_8bit_array_3.drv<63:0>.n80 0.0716912
R3799 hgu_cdac_8bit_array_3.drv<63:0>.n595 hgu_cdac_8bit_array_3.drv<63:0>.n594 0.0716912
R3800 hgu_cdac_8bit_array_3.drv<63:0>.n594 hgu_cdac_8bit_array_3.drv<63:0>.n593 0.0716912
R3801 hgu_cdac_8bit_array_3.drv<63:0>.n586 hgu_cdac_8bit_array_3.drv<63:0>.n585 0.0716912
R3802 hgu_cdac_8bit_array_3.drv<63:0>.n585 hgu_cdac_8bit_array_3.drv<63:0>.n584 0.0716912
R3803 hgu_cdac_8bit_array_3.drv<63:0>.n577 hgu_cdac_8bit_array_3.drv<63:0>.n576 0.0716912
R3804 hgu_cdac_8bit_array_3.drv<63:0>.n576 hgu_cdac_8bit_array_3.drv<63:0>.n575 0.0716912
R3805 hgu_cdac_8bit_array_3.drv<63:0>.n568 hgu_cdac_8bit_array_3.drv<63:0>.n567 0.0716912
R3806 hgu_cdac_8bit_array_3.drv<63:0>.n567 hgu_cdac_8bit_array_3.drv<63:0>.n566 0.0716912
R3807 hgu_cdac_8bit_array_3.drv<63:0>.n559 hgu_cdac_8bit_array_3.drv<63:0>.n558 0.0716912
R3808 hgu_cdac_8bit_array_3.drv<63:0>.n558 hgu_cdac_8bit_array_3.drv<63:0>.n557 0.0716912
R3809 hgu_cdac_8bit_array_3.drv<63:0>.n550 hgu_cdac_8bit_array_3.drv<63:0>.n549 0.0716912
R3810 hgu_cdac_8bit_array_3.drv<63:0>.n549 hgu_cdac_8bit_array_3.drv<63:0>.n548 0.0716912
R3811 hgu_cdac_8bit_array_3.drv<63:0>.n541 hgu_cdac_8bit_array_3.drv<63:0>.n540 0.0716912
R3812 hgu_cdac_8bit_array_3.drv<63:0>.n540 hgu_cdac_8bit_array_3.drv<63:0>.n539 0.0716912
R3813 hgu_cdac_8bit_array_3.drv<63:0>.n532 hgu_cdac_8bit_array_3.drv<63:0>.n531 0.0716912
R3814 hgu_cdac_8bit_array_3.drv<63:0>.n531 hgu_cdac_8bit_array_3.drv<63:0>.n530 0.0716912
R3815 hgu_cdac_8bit_array_3.drv<63:0>.n523 hgu_cdac_8bit_array_3.drv<63:0>.n522 0.0716912
R3816 hgu_cdac_8bit_array_3.drv<63:0>.n522 hgu_cdac_8bit_array_3.drv<63:0>.n521 0.0716912
R3817 hgu_cdac_8bit_array_3.drv<63:0>.n514 hgu_cdac_8bit_array_3.drv<63:0>.n513 0.0716912
R3818 hgu_cdac_8bit_array_3.drv<63:0>.n513 hgu_cdac_8bit_array_3.drv<63:0>.n512 0.0716912
R3819 hgu_cdac_8bit_array_3.drv<63:0>.n505 hgu_cdac_8bit_array_3.drv<63:0>.n504 0.0716912
R3820 hgu_cdac_8bit_array_3.drv<63:0>.n504 hgu_cdac_8bit_array_3.drv<63:0>.n503 0.0716912
R3821 hgu_cdac_8bit_array_3.drv<63:0>.n495 hgu_cdac_8bit_array_3.drv<63:0>.n494 0.0716912
R3822 hgu_cdac_8bit_array_3.drv<63:0>.n494 hgu_cdac_8bit_array_3.drv<63:0>.n493 0.0716912
R3823 hgu_cdac_8bit_array_3.drv<63:0>.n486 hgu_cdac_8bit_array_3.drv<63:0>.n485 0.0716912
R3824 hgu_cdac_8bit_array_3.drv<63:0>.n485 hgu_cdac_8bit_array_3.drv<63:0>.n484 0.0716912
R3825 hgu_cdac_8bit_array_3.drv<63:0>.n477 hgu_cdac_8bit_array_3.drv<63:0>.n476 0.0716912
R3826 hgu_cdac_8bit_array_3.drv<63:0>.n476 hgu_cdac_8bit_array_3.drv<63:0>.n475 0.0716912
R3827 hgu_cdac_8bit_array_3.drv<63:0>.n468 hgu_cdac_8bit_array_3.drv<63:0>.n467 0.0716912
R3828 hgu_cdac_8bit_array_3.drv<63:0>.n467 hgu_cdac_8bit_array_3.drv<63:0>.n466 0.0716912
R3829 hgu_cdac_8bit_array_3.drv<63:0>.n459 hgu_cdac_8bit_array_3.drv<63:0>.n458 0.0716912
R3830 hgu_cdac_8bit_array_3.drv<63:0>.n458 hgu_cdac_8bit_array_3.drv<63:0>.n457 0.0716912
R3831 hgu_cdac_8bit_array_3.drv<63:0>.n450 hgu_cdac_8bit_array_3.drv<63:0>.n449 0.0716912
R3832 hgu_cdac_8bit_array_3.drv<63:0>.n449 hgu_cdac_8bit_array_3.drv<63:0>.n448 0.0716912
R3833 hgu_cdac_8bit_array_3.drv<63:0>.n441 hgu_cdac_8bit_array_3.drv<63:0>.n440 0.0716912
R3834 hgu_cdac_8bit_array_3.drv<63:0>.n440 hgu_cdac_8bit_array_3.drv<63:0>.n439 0.0716912
R3835 hgu_cdac_8bit_array_3.drv<63:0>.n432 hgu_cdac_8bit_array_3.drv<63:0>.n431 0.0716912
R3836 hgu_cdac_8bit_array_3.drv<63:0>.n431 hgu_cdac_8bit_array_3.drv<63:0>.n430 0.0716912
R3837 hgu_cdac_8bit_array_3.drv<63:0>.n423 hgu_cdac_8bit_array_3.drv<63:0>.n422 0.0716912
R3838 hgu_cdac_8bit_array_3.drv<63:0>.n422 hgu_cdac_8bit_array_3.drv<63:0>.n421 0.0716912
R3839 hgu_cdac_8bit_array_3.drv<63:0>.n414 hgu_cdac_8bit_array_3.drv<63:0>.n413 0.0716912
R3840 hgu_cdac_8bit_array_3.drv<63:0>.n413 hgu_cdac_8bit_array_3.drv<63:0>.n412 0.0716912
R3841 hgu_cdac_8bit_array_3.drv<63:0>.n405 hgu_cdac_8bit_array_3.drv<63:0>.n404 0.0716912
R3842 hgu_cdac_8bit_array_3.drv<63:0>.n404 hgu_cdac_8bit_array_3.drv<63:0>.n403 0.0716912
R3843 hgu_cdac_8bit_array_3.drv<63:0>.n396 hgu_cdac_8bit_array_3.drv<63:0>.n395 0.0716912
R3844 hgu_cdac_8bit_array_3.drv<63:0>.n395 hgu_cdac_8bit_array_3.drv<63:0>.n394 0.0716912
R3845 hgu_cdac_8bit_array_3.drv<63:0>.n387 hgu_cdac_8bit_array_3.drv<63:0>.n386 0.0716912
R3846 hgu_cdac_8bit_array_3.drv<63:0>.n386 hgu_cdac_8bit_array_3.drv<63:0>.n385 0.0716912
R3847 hgu_cdac_8bit_array_3.drv<63:0>.n378 hgu_cdac_8bit_array_3.drv<63:0>.n377 0.0716912
R3848 hgu_cdac_8bit_array_3.drv<63:0>.n377 hgu_cdac_8bit_array_3.drv<63:0>.n376 0.0716912
R3849 hgu_cdac_8bit_array_3.drv<63:0>.n31 hgu_cdac_8bit_array_3.drv<63:0>.n30 0.0716912
R3850 hgu_cdac_8bit_array_3.drv<63:0>.n28 hgu_cdac_8bit_array_3.drv<63:0>.n27 0.0716912
R3851 hgu_cdac_8bit_array_3.drv<63:0>.n21 hgu_cdac_8bit_array_3.drv<63:0>.n20 0.0716912
R3852 hgu_cdac_8bit_array_3.drv<63:0>.n14 hgu_cdac_8bit_array_3.drv<63:0>.n13 0.0716912
R3853 hgu_cdac_8bit_array_3.drv<63:0>.n7 hgu_cdac_8bit_array_3.drv<63:0>.n6 0.0716912
R3854 hgu_cdac_8bit_array_3.drv<63:0>.n88 hgu_cdac_8bit_array_3.drv<63:0>.n87 0.0716912
R3855 hgu_cdac_8bit_array_3.drv<63:0>.n95 hgu_cdac_8bit_array_3.drv<63:0>.n94 0.0716912
R3856 hgu_cdac_8bit_array_3.drv<63:0>.n102 hgu_cdac_8bit_array_3.drv<63:0>.n101 0.0716912
R3857 hgu_cdac_8bit_array_3.drv<63:0>.n109 hgu_cdac_8bit_array_3.drv<63:0>.n108 0.0716912
R3858 hgu_cdac_8bit_array_3.drv<63:0>.n116 hgu_cdac_8bit_array_3.drv<63:0>.n115 0.0716912
R3859 hgu_cdac_8bit_array_3.drv<63:0>.n123 hgu_cdac_8bit_array_3.drv<63:0>.n122 0.0716912
R3860 hgu_cdac_8bit_array_3.drv<63:0>.n130 hgu_cdac_8bit_array_3.drv<63:0>.n129 0.0716912
R3861 hgu_cdac_8bit_array_3.drv<63:0>.n137 hgu_cdac_8bit_array_3.drv<63:0>.n136 0.0716912
R3862 hgu_cdac_8bit_array_3.drv<63:0>.n144 hgu_cdac_8bit_array_3.drv<63:0>.n143 0.0716912
R3863 hgu_cdac_8bit_array_3.drv<63:0>.n151 hgu_cdac_8bit_array_3.drv<63:0>.n150 0.0716912
R3864 hgu_cdac_8bit_array_3.drv<63:0>.n158 hgu_cdac_8bit_array_3.drv<63:0>.n157 0.0716912
R3865 hgu_cdac_8bit_array_3.drv<63:0>.n168 hgu_cdac_8bit_array_3.drv<63:0>.n167 0.0716912
R3866 hgu_cdac_8bit_array_3.drv<63:0>.n176 hgu_cdac_8bit_array_3.drv<63:0>.n175 0.0716912
R3867 hgu_cdac_8bit_array_3.drv<63:0>.n194 hgu_cdac_8bit_array_3.drv<63:0>.n193 0.0716912
R3868 hgu_cdac_8bit_array_3.drv<63:0>.n214 hgu_cdac_8bit_array_3.drv<63:0>.n213 0.0716912
R3869 hgu_cdac_8bit_array_3.drv<63:0>.n232 hgu_cdac_8bit_array_3.drv<63:0>.n231 0.0716912
R3870 hgu_cdac_8bit_array_3.drv<63:0>.n247 hgu_cdac_8bit_array_3.drv<63:0>.n246 0.0716912
R3871 hgu_cdac_8bit_array_3.drv<63:0>.n268 hgu_cdac_8bit_array_3.drv<63:0>.n267 0.0716912
R3872 hgu_cdac_8bit_array_3.drv<63:0>.n276 hgu_cdac_8bit_array_3.drv<63:0>.n275 0.0716912
R3873 hgu_cdac_8bit_array_3.drv<63:0>.n290 hgu_cdac_8bit_array_3.drv<63:0>.n289 0.0716912
R3874 hgu_cdac_8bit_array_3.drv<63:0>.n298 hgu_cdac_8bit_array_3.drv<63:0>.n297 0.0716912
R3875 hgu_cdac_8bit_array_3.drv<63:0>.n323 hgu_cdac_8bit_array_3.drv<63:0>.n322 0.0716912
R3876 hgu_cdac_8bit_array_3.drv<63:0>.n341 hgu_cdac_8bit_array_3.drv<63:0>.n340 0.0716912
R3877 hgu_cdac_8bit_array_3.drv<63:0>.n356 hgu_cdac_8bit_array_3.drv<63:0>.n355 0.0716912
R3878 hgu_cdac_8bit_array_3.drv<63:0>.n371 hgu_cdac_8bit_array_3.drv<63:0>.n370 0.0716912
R3879 hgu_cdac_8bit_array_3.drv<63:0>.n502 hgu_cdac_8bit_array_3.drv<63:0> 0.0694333
R3880 hgu_cdac_8bit_array_3.drv<63:0>.n33 hgu_cdac_8bit_array_3.drv<63:0>.n32 0.0665339
R3881 hgu_cdac_8bit_array_3.drv<63:0>.n374 hgu_cdac_8bit_array_3.drv<63:0>.n373 0.0664894
R3882 hgu_cdac_8bit_array_3.drv<63:0>.n240 hgu_cdac_8bit_array_3.drv<63:0>.n236 0.0571406
R3883 hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_8bit_array_3.drv<63:0>.n602 0.0564853
R3884 hgu_cdac_8bit_array_3.drv<63:0>.n35 hgu_cdac_8bit_array_3.drv<63:0>.n34 0.0557941
R3885 hgu_cdac_8bit_array_3.drv<63:0>.n38 hgu_cdac_8bit_array_3.drv<63:0>.n37 0.0557941
R3886 hgu_cdac_8bit_array_3.drv<63:0>.n41 hgu_cdac_8bit_array_3.drv<63:0>.n40 0.0557941
R3887 hgu_cdac_8bit_array_3.drv<63:0>.n44 hgu_cdac_8bit_array_3.drv<63:0>.n43 0.0557941
R3888 hgu_cdac_8bit_array_3.drv<63:0>.n47 hgu_cdac_8bit_array_3.drv<63:0>.n46 0.0557941
R3889 hgu_cdac_8bit_array_3.drv<63:0>.n50 hgu_cdac_8bit_array_3.drv<63:0>.n49 0.0557941
R3890 hgu_cdac_8bit_array_3.drv<63:0>.n53 hgu_cdac_8bit_array_3.drv<63:0>.n52 0.0557941
R3891 hgu_cdac_8bit_array_3.drv<63:0>.n56 hgu_cdac_8bit_array_3.drv<63:0>.n55 0.0557941
R3892 hgu_cdac_8bit_array_3.drv<63:0>.n59 hgu_cdac_8bit_array_3.drv<63:0>.n58 0.0557941
R3893 hgu_cdac_8bit_array_3.drv<63:0>.n62 hgu_cdac_8bit_array_3.drv<63:0>.n61 0.0557941
R3894 hgu_cdac_8bit_array_3.drv<63:0>.n65 hgu_cdac_8bit_array_3.drv<63:0>.n64 0.0557941
R3895 hgu_cdac_8bit_array_3.drv<63:0>.n68 hgu_cdac_8bit_array_3.drv<63:0>.n67 0.0557941
R3896 hgu_cdac_8bit_array_3.drv<63:0>.n71 hgu_cdac_8bit_array_3.drv<63:0>.n70 0.0557941
R3897 hgu_cdac_8bit_array_3.drv<63:0>.n74 hgu_cdac_8bit_array_3.drv<63:0>.n73 0.0557941
R3898 hgu_cdac_8bit_array_3.drv<63:0>.n77 hgu_cdac_8bit_array_3.drv<63:0>.n76 0.0557941
R3899 hgu_cdac_8bit_array_3.drv<63:0>.n80 hgu_cdac_8bit_array_3.drv<63:0>.n79 0.0557941
R3900 hgu_cdac_8bit_array_3.drv<63:0>.n602 hgu_cdac_8bit_array_3.drv<63:0>.n601 0.0557941
R3901 hgu_cdac_8bit_array_3.drv<63:0>.n599 hgu_cdac_8bit_array_3.drv<63:0>.n598 0.0557941
R3902 hgu_cdac_8bit_array_3.drv<63:0>.n596 hgu_cdac_8bit_array_3.drv<63:0>.n595 0.0557941
R3903 hgu_cdac_8bit_array_3.drv<63:0>.n593 hgu_cdac_8bit_array_3.drv<63:0>.n592 0.0557941
R3904 hgu_cdac_8bit_array_3.drv<63:0>.n590 hgu_cdac_8bit_array_3.drv<63:0>.n589 0.0557941
R3905 hgu_cdac_8bit_array_3.drv<63:0>.n587 hgu_cdac_8bit_array_3.drv<63:0>.n586 0.0557941
R3906 hgu_cdac_8bit_array_3.drv<63:0>.n584 hgu_cdac_8bit_array_3.drv<63:0>.n583 0.0557941
R3907 hgu_cdac_8bit_array_3.drv<63:0>.n581 hgu_cdac_8bit_array_3.drv<63:0>.n580 0.0557941
R3908 hgu_cdac_8bit_array_3.drv<63:0>.n578 hgu_cdac_8bit_array_3.drv<63:0>.n577 0.0557941
R3909 hgu_cdac_8bit_array_3.drv<63:0>.n575 hgu_cdac_8bit_array_3.drv<63:0>.n574 0.0557941
R3910 hgu_cdac_8bit_array_3.drv<63:0>.n572 hgu_cdac_8bit_array_3.drv<63:0>.n571 0.0557941
R3911 hgu_cdac_8bit_array_3.drv<63:0>.n569 hgu_cdac_8bit_array_3.drv<63:0>.n568 0.0557941
R3912 hgu_cdac_8bit_array_3.drv<63:0>.n566 hgu_cdac_8bit_array_3.drv<63:0>.n565 0.0557941
R3913 hgu_cdac_8bit_array_3.drv<63:0>.n563 hgu_cdac_8bit_array_3.drv<63:0>.n562 0.0557941
R3914 hgu_cdac_8bit_array_3.drv<63:0>.n560 hgu_cdac_8bit_array_3.drv<63:0>.n559 0.0557941
R3915 hgu_cdac_8bit_array_3.drv<63:0>.n557 hgu_cdac_8bit_array_3.drv<63:0>.n556 0.0557941
R3916 hgu_cdac_8bit_array_3.drv<63:0>.n554 hgu_cdac_8bit_array_3.drv<63:0>.n553 0.0557941
R3917 hgu_cdac_8bit_array_3.drv<63:0>.n551 hgu_cdac_8bit_array_3.drv<63:0>.n550 0.0557941
R3918 hgu_cdac_8bit_array_3.drv<63:0>.n548 hgu_cdac_8bit_array_3.drv<63:0>.n547 0.0557941
R3919 hgu_cdac_8bit_array_3.drv<63:0>.n545 hgu_cdac_8bit_array_3.drv<63:0>.n544 0.0557941
R3920 hgu_cdac_8bit_array_3.drv<63:0>.n542 hgu_cdac_8bit_array_3.drv<63:0>.n541 0.0557941
R3921 hgu_cdac_8bit_array_3.drv<63:0>.n539 hgu_cdac_8bit_array_3.drv<63:0>.n538 0.0557941
R3922 hgu_cdac_8bit_array_3.drv<63:0>.n536 hgu_cdac_8bit_array_3.drv<63:0>.n535 0.0557941
R3923 hgu_cdac_8bit_array_3.drv<63:0>.n533 hgu_cdac_8bit_array_3.drv<63:0>.n532 0.0557941
R3924 hgu_cdac_8bit_array_3.drv<63:0>.n530 hgu_cdac_8bit_array_3.drv<63:0>.n529 0.0557941
R3925 hgu_cdac_8bit_array_3.drv<63:0>.n527 hgu_cdac_8bit_array_3.drv<63:0>.n526 0.0557941
R3926 hgu_cdac_8bit_array_3.drv<63:0>.n524 hgu_cdac_8bit_array_3.drv<63:0>.n523 0.0557941
R3927 hgu_cdac_8bit_array_3.drv<63:0>.n521 hgu_cdac_8bit_array_3.drv<63:0>.n520 0.0557941
R3928 hgu_cdac_8bit_array_3.drv<63:0>.n518 hgu_cdac_8bit_array_3.drv<63:0>.n517 0.0557941
R3929 hgu_cdac_8bit_array_3.drv<63:0>.n515 hgu_cdac_8bit_array_3.drv<63:0>.n514 0.0557941
R3930 hgu_cdac_8bit_array_3.drv<63:0>.n512 hgu_cdac_8bit_array_3.drv<63:0>.n511 0.0557941
R3931 hgu_cdac_8bit_array_3.drv<63:0>.n509 hgu_cdac_8bit_array_3.drv<63:0>.n508 0.0557941
R3932 hgu_cdac_8bit_array_3.drv<63:0>.n506 hgu_cdac_8bit_array_3.drv<63:0>.n505 0.0557941
R3933 hgu_cdac_8bit_array_3.drv<63:0>.n499 hgu_cdac_8bit_array_3.drv<63:0>.n498 0.0557941
R3934 hgu_cdac_8bit_array_3.drv<63:0>.n496 hgu_cdac_8bit_array_3.drv<63:0>.n495 0.0557941
R3935 hgu_cdac_8bit_array_3.drv<63:0>.n493 hgu_cdac_8bit_array_3.drv<63:0>.n492 0.0557941
R3936 hgu_cdac_8bit_array_3.drv<63:0>.n490 hgu_cdac_8bit_array_3.drv<63:0>.n489 0.0557941
R3937 hgu_cdac_8bit_array_3.drv<63:0>.n487 hgu_cdac_8bit_array_3.drv<63:0>.n486 0.0557941
R3938 hgu_cdac_8bit_array_3.drv<63:0>.n484 hgu_cdac_8bit_array_3.drv<63:0>.n483 0.0557941
R3939 hgu_cdac_8bit_array_3.drv<63:0>.n481 hgu_cdac_8bit_array_3.drv<63:0>.n480 0.0557941
R3940 hgu_cdac_8bit_array_3.drv<63:0>.n478 hgu_cdac_8bit_array_3.drv<63:0>.n477 0.0557941
R3941 hgu_cdac_8bit_array_3.drv<63:0>.n475 hgu_cdac_8bit_array_3.drv<63:0>.n474 0.0557941
R3942 hgu_cdac_8bit_array_3.drv<63:0>.n472 hgu_cdac_8bit_array_3.drv<63:0>.n471 0.0557941
R3943 hgu_cdac_8bit_array_3.drv<63:0>.n469 hgu_cdac_8bit_array_3.drv<63:0>.n468 0.0557941
R3944 hgu_cdac_8bit_array_3.drv<63:0>.n466 hgu_cdac_8bit_array_3.drv<63:0>.n465 0.0557941
R3945 hgu_cdac_8bit_array_3.drv<63:0>.n463 hgu_cdac_8bit_array_3.drv<63:0>.n462 0.0557941
R3946 hgu_cdac_8bit_array_3.drv<63:0>.n460 hgu_cdac_8bit_array_3.drv<63:0>.n459 0.0557941
R3947 hgu_cdac_8bit_array_3.drv<63:0>.n457 hgu_cdac_8bit_array_3.drv<63:0>.n456 0.0557941
R3948 hgu_cdac_8bit_array_3.drv<63:0>.n454 hgu_cdac_8bit_array_3.drv<63:0>.n453 0.0557941
R3949 hgu_cdac_8bit_array_3.drv<63:0>.n451 hgu_cdac_8bit_array_3.drv<63:0>.n450 0.0557941
R3950 hgu_cdac_8bit_array_3.drv<63:0>.n448 hgu_cdac_8bit_array_3.drv<63:0>.n447 0.0557941
R3951 hgu_cdac_8bit_array_3.drv<63:0>.n445 hgu_cdac_8bit_array_3.drv<63:0>.n444 0.0557941
R3952 hgu_cdac_8bit_array_3.drv<63:0>.n442 hgu_cdac_8bit_array_3.drv<63:0>.n441 0.0557941
R3953 hgu_cdac_8bit_array_3.drv<63:0>.n439 hgu_cdac_8bit_array_3.drv<63:0>.n438 0.0557941
R3954 hgu_cdac_8bit_array_3.drv<63:0>.n436 hgu_cdac_8bit_array_3.drv<63:0>.n435 0.0557941
R3955 hgu_cdac_8bit_array_3.drv<63:0>.n433 hgu_cdac_8bit_array_3.drv<63:0>.n432 0.0557941
R3956 hgu_cdac_8bit_array_3.drv<63:0>.n430 hgu_cdac_8bit_array_3.drv<63:0>.n429 0.0557941
R3957 hgu_cdac_8bit_array_3.drv<63:0>.n427 hgu_cdac_8bit_array_3.drv<63:0>.n426 0.0557941
R3958 hgu_cdac_8bit_array_3.drv<63:0>.n424 hgu_cdac_8bit_array_3.drv<63:0>.n423 0.0557941
R3959 hgu_cdac_8bit_array_3.drv<63:0>.n421 hgu_cdac_8bit_array_3.drv<63:0>.n420 0.0557941
R3960 hgu_cdac_8bit_array_3.drv<63:0>.n418 hgu_cdac_8bit_array_3.drv<63:0>.n417 0.0557941
R3961 hgu_cdac_8bit_array_3.drv<63:0>.n415 hgu_cdac_8bit_array_3.drv<63:0>.n414 0.0557941
R3962 hgu_cdac_8bit_array_3.drv<63:0>.n412 hgu_cdac_8bit_array_3.drv<63:0>.n411 0.0557941
R3963 hgu_cdac_8bit_array_3.drv<63:0>.n409 hgu_cdac_8bit_array_3.drv<63:0>.n408 0.0557941
R3964 hgu_cdac_8bit_array_3.drv<63:0>.n406 hgu_cdac_8bit_array_3.drv<63:0>.n405 0.0557941
R3965 hgu_cdac_8bit_array_3.drv<63:0>.n403 hgu_cdac_8bit_array_3.drv<63:0>.n402 0.0557941
R3966 hgu_cdac_8bit_array_3.drv<63:0>.n400 hgu_cdac_8bit_array_3.drv<63:0>.n399 0.0557941
R3967 hgu_cdac_8bit_array_3.drv<63:0>.n397 hgu_cdac_8bit_array_3.drv<63:0>.n396 0.0557941
R3968 hgu_cdac_8bit_array_3.drv<63:0>.n394 hgu_cdac_8bit_array_3.drv<63:0>.n393 0.0557941
R3969 hgu_cdac_8bit_array_3.drv<63:0>.n391 hgu_cdac_8bit_array_3.drv<63:0>.n390 0.0557941
R3970 hgu_cdac_8bit_array_3.drv<63:0>.n388 hgu_cdac_8bit_array_3.drv<63:0>.n387 0.0557941
R3971 hgu_cdac_8bit_array_3.drv<63:0>.n385 hgu_cdac_8bit_array_3.drv<63:0>.n384 0.0557941
R3972 hgu_cdac_8bit_array_3.drv<63:0>.n382 hgu_cdac_8bit_array_3.drv<63:0>.n381 0.0557941
R3973 hgu_cdac_8bit_array_3.drv<63:0>.n379 hgu_cdac_8bit_array_3.drv<63:0>.n378 0.0557941
R3974 hgu_cdac_8bit_array_3.drv<63:0>.n376 hgu_cdac_8bit_array_3.drv<63:0>.n375 0.0557941
R3975 hgu_cdac_8bit_array_3.drv<63:0>.n30 hgu_cdac_8bit_array_3.drv<63:0>.n29 0.0557941
R3976 hgu_cdac_8bit_array_3.drv<63:0>.n23 hgu_cdac_8bit_array_3.drv<63:0>.n22 0.0557941
R3977 hgu_cdac_8bit_array_3.drv<63:0>.n24 hgu_cdac_8bit_array_3.drv<63:0>.n23 0.0557941
R3978 hgu_cdac_8bit_array_3.drv<63:0>.n25 hgu_cdac_8bit_array_3.drv<63:0>.n24 0.0557941
R3979 hgu_cdac_8bit_array_3.drv<63:0>.n26 hgu_cdac_8bit_array_3.drv<63:0>.n25 0.0557941
R3980 hgu_cdac_8bit_array_3.drv<63:0>.n27 hgu_cdac_8bit_array_3.drv<63:0>.n26 0.0557941
R3981 hgu_cdac_8bit_array_3.drv<63:0>.n16 hgu_cdac_8bit_array_3.drv<63:0>.n15 0.0557941
R3982 hgu_cdac_8bit_array_3.drv<63:0>.n17 hgu_cdac_8bit_array_3.drv<63:0>.n16 0.0557941
R3983 hgu_cdac_8bit_array_3.drv<63:0>.n18 hgu_cdac_8bit_array_3.drv<63:0>.n17 0.0557941
R3984 hgu_cdac_8bit_array_3.drv<63:0>.n19 hgu_cdac_8bit_array_3.drv<63:0>.n18 0.0557941
R3985 hgu_cdac_8bit_array_3.drv<63:0>.n20 hgu_cdac_8bit_array_3.drv<63:0>.n19 0.0557941
R3986 hgu_cdac_8bit_array_3.drv<63:0>.n9 hgu_cdac_8bit_array_3.drv<63:0>.n8 0.0557941
R3987 hgu_cdac_8bit_array_3.drv<63:0>.n10 hgu_cdac_8bit_array_3.drv<63:0>.n9 0.0557941
R3988 hgu_cdac_8bit_array_3.drv<63:0>.n11 hgu_cdac_8bit_array_3.drv<63:0>.n10 0.0557941
R3989 hgu_cdac_8bit_array_3.drv<63:0>.n12 hgu_cdac_8bit_array_3.drv<63:0>.n11 0.0557941
R3990 hgu_cdac_8bit_array_3.drv<63:0>.n13 hgu_cdac_8bit_array_3.drv<63:0>.n12 0.0557941
R3991 hgu_cdac_8bit_array_3.drv<63:0>.n2 hgu_cdac_8bit_array_3.drv<63:0>.n1 0.0557941
R3992 hgu_cdac_8bit_array_3.drv<63:0>.n3 hgu_cdac_8bit_array_3.drv<63:0>.n2 0.0557941
R3993 hgu_cdac_8bit_array_3.drv<63:0>.n4 hgu_cdac_8bit_array_3.drv<63:0>.n3 0.0557941
R3994 hgu_cdac_8bit_array_3.drv<63:0>.n5 hgu_cdac_8bit_array_3.drv<63:0>.n4 0.0557941
R3995 hgu_cdac_8bit_array_3.drv<63:0>.n6 hgu_cdac_8bit_array_3.drv<63:0>.n5 0.0557941
R3996 hgu_cdac_8bit_array_3.drv<63:0>.n87 hgu_cdac_8bit_array_3.drv<63:0>.n86 0.0557941
R3997 hgu_cdac_8bit_array_3.drv<63:0>.n86 hgu_cdac_8bit_array_3.drv<63:0>.n85 0.0557941
R3998 hgu_cdac_8bit_array_3.drv<63:0>.n85 hgu_cdac_8bit_array_3.drv<63:0>.n84 0.0557941
R3999 hgu_cdac_8bit_array_3.drv<63:0>.n84 hgu_cdac_8bit_array_3.drv<63:0>.n83 0.0557941
R4000 hgu_cdac_8bit_array_3.drv<63:0>.n83 hgu_cdac_8bit_array_3.drv<63:0>.n82 0.0557941
R4001 hgu_cdac_8bit_array_3.drv<63:0>.n94 hgu_cdac_8bit_array_3.drv<63:0>.n93 0.0557941
R4002 hgu_cdac_8bit_array_3.drv<63:0>.n93 hgu_cdac_8bit_array_3.drv<63:0>.n92 0.0557941
R4003 hgu_cdac_8bit_array_3.drv<63:0>.n92 hgu_cdac_8bit_array_3.drv<63:0>.n91 0.0557941
R4004 hgu_cdac_8bit_array_3.drv<63:0>.n91 hgu_cdac_8bit_array_3.drv<63:0>.n90 0.0557941
R4005 hgu_cdac_8bit_array_3.drv<63:0>.n90 hgu_cdac_8bit_array_3.drv<63:0>.n89 0.0557941
R4006 hgu_cdac_8bit_array_3.drv<63:0>.n101 hgu_cdac_8bit_array_3.drv<63:0>.n100 0.0557941
R4007 hgu_cdac_8bit_array_3.drv<63:0>.n100 hgu_cdac_8bit_array_3.drv<63:0>.n99 0.0557941
R4008 hgu_cdac_8bit_array_3.drv<63:0>.n99 hgu_cdac_8bit_array_3.drv<63:0>.n98 0.0557941
R4009 hgu_cdac_8bit_array_3.drv<63:0>.n98 hgu_cdac_8bit_array_3.drv<63:0>.n97 0.0557941
R4010 hgu_cdac_8bit_array_3.drv<63:0>.n97 hgu_cdac_8bit_array_3.drv<63:0>.n96 0.0557941
R4011 hgu_cdac_8bit_array_3.drv<63:0>.n108 hgu_cdac_8bit_array_3.drv<63:0>.n107 0.0557941
R4012 hgu_cdac_8bit_array_3.drv<63:0>.n107 hgu_cdac_8bit_array_3.drv<63:0>.n106 0.0557941
R4013 hgu_cdac_8bit_array_3.drv<63:0>.n106 hgu_cdac_8bit_array_3.drv<63:0>.n105 0.0557941
R4014 hgu_cdac_8bit_array_3.drv<63:0>.n105 hgu_cdac_8bit_array_3.drv<63:0>.n104 0.0557941
R4015 hgu_cdac_8bit_array_3.drv<63:0>.n104 hgu_cdac_8bit_array_3.drv<63:0>.n103 0.0557941
R4016 hgu_cdac_8bit_array_3.drv<63:0>.n115 hgu_cdac_8bit_array_3.drv<63:0>.n114 0.0557941
R4017 hgu_cdac_8bit_array_3.drv<63:0>.n114 hgu_cdac_8bit_array_3.drv<63:0>.n113 0.0557941
R4018 hgu_cdac_8bit_array_3.drv<63:0>.n113 hgu_cdac_8bit_array_3.drv<63:0>.n112 0.0557941
R4019 hgu_cdac_8bit_array_3.drv<63:0>.n112 hgu_cdac_8bit_array_3.drv<63:0>.n111 0.0557941
R4020 hgu_cdac_8bit_array_3.drv<63:0>.n111 hgu_cdac_8bit_array_3.drv<63:0>.n110 0.0557941
R4021 hgu_cdac_8bit_array_3.drv<63:0>.n122 hgu_cdac_8bit_array_3.drv<63:0>.n121 0.0557941
R4022 hgu_cdac_8bit_array_3.drv<63:0>.n121 hgu_cdac_8bit_array_3.drv<63:0>.n120 0.0557941
R4023 hgu_cdac_8bit_array_3.drv<63:0>.n120 hgu_cdac_8bit_array_3.drv<63:0>.n119 0.0557941
R4024 hgu_cdac_8bit_array_3.drv<63:0>.n119 hgu_cdac_8bit_array_3.drv<63:0>.n118 0.0557941
R4025 hgu_cdac_8bit_array_3.drv<63:0>.n118 hgu_cdac_8bit_array_3.drv<63:0>.n117 0.0557941
R4026 hgu_cdac_8bit_array_3.drv<63:0>.n129 hgu_cdac_8bit_array_3.drv<63:0>.n128 0.0557941
R4027 hgu_cdac_8bit_array_3.drv<63:0>.n128 hgu_cdac_8bit_array_3.drv<63:0>.n127 0.0557941
R4028 hgu_cdac_8bit_array_3.drv<63:0>.n127 hgu_cdac_8bit_array_3.drv<63:0>.n126 0.0557941
R4029 hgu_cdac_8bit_array_3.drv<63:0>.n126 hgu_cdac_8bit_array_3.drv<63:0>.n125 0.0557941
R4030 hgu_cdac_8bit_array_3.drv<63:0>.n125 hgu_cdac_8bit_array_3.drv<63:0>.n124 0.0557941
R4031 hgu_cdac_8bit_array_3.drv<63:0>.n136 hgu_cdac_8bit_array_3.drv<63:0>.n135 0.0557941
R4032 hgu_cdac_8bit_array_3.drv<63:0>.n135 hgu_cdac_8bit_array_3.drv<63:0>.n134 0.0557941
R4033 hgu_cdac_8bit_array_3.drv<63:0>.n134 hgu_cdac_8bit_array_3.drv<63:0>.n133 0.0557941
R4034 hgu_cdac_8bit_array_3.drv<63:0>.n133 hgu_cdac_8bit_array_3.drv<63:0>.n132 0.0557941
R4035 hgu_cdac_8bit_array_3.drv<63:0>.n132 hgu_cdac_8bit_array_3.drv<63:0>.n131 0.0557941
R4036 hgu_cdac_8bit_array_3.drv<63:0>.n143 hgu_cdac_8bit_array_3.drv<63:0>.n142 0.0557941
R4037 hgu_cdac_8bit_array_3.drv<63:0>.n142 hgu_cdac_8bit_array_3.drv<63:0>.n141 0.0557941
R4038 hgu_cdac_8bit_array_3.drv<63:0>.n141 hgu_cdac_8bit_array_3.drv<63:0>.n140 0.0557941
R4039 hgu_cdac_8bit_array_3.drv<63:0>.n140 hgu_cdac_8bit_array_3.drv<63:0>.n139 0.0557941
R4040 hgu_cdac_8bit_array_3.drv<63:0>.n139 hgu_cdac_8bit_array_3.drv<63:0>.n138 0.0557941
R4041 hgu_cdac_8bit_array_3.drv<63:0>.n150 hgu_cdac_8bit_array_3.drv<63:0>.n149 0.0557941
R4042 hgu_cdac_8bit_array_3.drv<63:0>.n149 hgu_cdac_8bit_array_3.drv<63:0>.n148 0.0557941
R4043 hgu_cdac_8bit_array_3.drv<63:0>.n148 hgu_cdac_8bit_array_3.drv<63:0>.n147 0.0557941
R4044 hgu_cdac_8bit_array_3.drv<63:0>.n147 hgu_cdac_8bit_array_3.drv<63:0>.n146 0.0557941
R4045 hgu_cdac_8bit_array_3.drv<63:0>.n146 hgu_cdac_8bit_array_3.drv<63:0>.n145 0.0557941
R4046 hgu_cdac_8bit_array_3.drv<63:0>.n157 hgu_cdac_8bit_array_3.drv<63:0>.n156 0.0557941
R4047 hgu_cdac_8bit_array_3.drv<63:0>.n156 hgu_cdac_8bit_array_3.drv<63:0>.n155 0.0557941
R4048 hgu_cdac_8bit_array_3.drv<63:0>.n155 hgu_cdac_8bit_array_3.drv<63:0>.n154 0.0557941
R4049 hgu_cdac_8bit_array_3.drv<63:0>.n154 hgu_cdac_8bit_array_3.drv<63:0>.n153 0.0557941
R4050 hgu_cdac_8bit_array_3.drv<63:0>.n153 hgu_cdac_8bit_array_3.drv<63:0>.n152 0.0557941
R4051 hgu_cdac_8bit_array_3.drv<63:0>.n167 hgu_cdac_8bit_array_3.drv<63:0>.n166 0.0557941
R4052 hgu_cdac_8bit_array_3.drv<63:0>.n166 hgu_cdac_8bit_array_3.drv<63:0>.n165 0.0557941
R4053 hgu_cdac_8bit_array_3.drv<63:0>.n165 hgu_cdac_8bit_array_3.drv<63:0>.n164 0.0557941
R4054 hgu_cdac_8bit_array_3.drv<63:0>.n164 hgu_cdac_8bit_array_3.drv<63:0>.n163 0.0557941
R4055 hgu_cdac_8bit_array_3.drv<63:0>.n163 hgu_cdac_8bit_array_3.drv<63:0>.n162 0.0557941
R4056 hgu_cdac_8bit_array_3.drv<63:0>.n175 hgu_cdac_8bit_array_3.drv<63:0>.n174 0.0557941
R4057 hgu_cdac_8bit_array_3.drv<63:0>.n174 hgu_cdac_8bit_array_3.drv<63:0>.n173 0.0557941
R4058 hgu_cdac_8bit_array_3.drv<63:0>.n173 hgu_cdac_8bit_array_3.drv<63:0>.n172 0.0557941
R4059 hgu_cdac_8bit_array_3.drv<63:0>.n172 hgu_cdac_8bit_array_3.drv<63:0>.n171 0.0557941
R4060 hgu_cdac_8bit_array_3.drv<63:0>.n171 hgu_cdac_8bit_array_3.drv<63:0>.n170 0.0557941
R4061 hgu_cdac_8bit_array_3.drv<63:0>.n193 hgu_cdac_8bit_array_3.drv<63:0>.n192 0.0557941
R4062 hgu_cdac_8bit_array_3.drv<63:0>.n192 hgu_cdac_8bit_array_3.drv<63:0>.n191 0.0557941
R4063 hgu_cdac_8bit_array_3.drv<63:0>.n191 hgu_cdac_8bit_array_3.drv<63:0>.n190 0.0557941
R4064 hgu_cdac_8bit_array_3.drv<63:0>.n190 hgu_cdac_8bit_array_3.drv<63:0>.n189 0.0557941
R4065 hgu_cdac_8bit_array_3.drv<63:0>.n189 hgu_cdac_8bit_array_3.drv<63:0>.n188 0.0557941
R4066 hgu_cdac_8bit_array_3.drv<63:0>.n213 hgu_cdac_8bit_array_3.drv<63:0>.n212 0.0557941
R4067 hgu_cdac_8bit_array_3.drv<63:0>.n212 hgu_cdac_8bit_array_3.drv<63:0>.n211 0.0557941
R4068 hgu_cdac_8bit_array_3.drv<63:0>.n211 hgu_cdac_8bit_array_3.drv<63:0>.n210 0.0557941
R4069 hgu_cdac_8bit_array_3.drv<63:0>.n210 hgu_cdac_8bit_array_3.drv<63:0>.n209 0.0557941
R4070 hgu_cdac_8bit_array_3.drv<63:0>.n209 hgu_cdac_8bit_array_3.drv<63:0>.n208 0.0557941
R4071 hgu_cdac_8bit_array_3.drv<63:0>.n231 hgu_cdac_8bit_array_3.drv<63:0>.n230 0.0557941
R4072 hgu_cdac_8bit_array_3.drv<63:0>.n230 hgu_cdac_8bit_array_3.drv<63:0>.n229 0.0557941
R4073 hgu_cdac_8bit_array_3.drv<63:0>.n229 hgu_cdac_8bit_array_3.drv<63:0>.n228 0.0557941
R4074 hgu_cdac_8bit_array_3.drv<63:0>.n228 hgu_cdac_8bit_array_3.drv<63:0>.n227 0.0557941
R4075 hgu_cdac_8bit_array_3.drv<63:0>.n227 hgu_cdac_8bit_array_3.drv<63:0>.n226 0.0557941
R4076 hgu_cdac_8bit_array_3.drv<63:0>.n246 hgu_cdac_8bit_array_3.drv<63:0>.n245 0.0557941
R4077 hgu_cdac_8bit_array_3.drv<63:0>.n245 hgu_cdac_8bit_array_3.drv<63:0>.n244 0.0557941
R4078 hgu_cdac_8bit_array_3.drv<63:0>.n244 hgu_cdac_8bit_array_3.drv<63:0>.n243 0.0557941
R4079 hgu_cdac_8bit_array_3.drv<63:0>.n243 hgu_cdac_8bit_array_3.drv<63:0>.n242 0.0557941
R4080 hgu_cdac_8bit_array_3.drv<63:0>.n242 hgu_cdac_8bit_array_3.drv<63:0>.n241 0.0557941
R4081 hgu_cdac_8bit_array_3.drv<63:0>.n267 hgu_cdac_8bit_array_3.drv<63:0>.n266 0.0557941
R4082 hgu_cdac_8bit_array_3.drv<63:0>.n266 hgu_cdac_8bit_array_3.drv<63:0>.n265 0.0557941
R4083 hgu_cdac_8bit_array_3.drv<63:0>.n265 hgu_cdac_8bit_array_3.drv<63:0>.n264 0.0557941
R4084 hgu_cdac_8bit_array_3.drv<63:0>.n264 hgu_cdac_8bit_array_3.drv<63:0>.n263 0.0557941
R4085 hgu_cdac_8bit_array_3.drv<63:0>.n263 hgu_cdac_8bit_array_3.drv<63:0>.n262 0.0557941
R4086 hgu_cdac_8bit_array_3.drv<63:0>.n275 hgu_cdac_8bit_array_3.drv<63:0>.n274 0.0557941
R4087 hgu_cdac_8bit_array_3.drv<63:0>.n274 hgu_cdac_8bit_array_3.drv<63:0>.n273 0.0557941
R4088 hgu_cdac_8bit_array_3.drv<63:0>.n273 hgu_cdac_8bit_array_3.drv<63:0>.n272 0.0557941
R4089 hgu_cdac_8bit_array_3.drv<63:0>.n272 hgu_cdac_8bit_array_3.drv<63:0>.n271 0.0557941
R4090 hgu_cdac_8bit_array_3.drv<63:0>.n271 hgu_cdac_8bit_array_3.drv<63:0>.n270 0.0557941
R4091 hgu_cdac_8bit_array_3.drv<63:0>.n289 hgu_cdac_8bit_array_3.drv<63:0>.n288 0.0557941
R4092 hgu_cdac_8bit_array_3.drv<63:0>.n288 hgu_cdac_8bit_array_3.drv<63:0>.n287 0.0557941
R4093 hgu_cdac_8bit_array_3.drv<63:0>.n287 hgu_cdac_8bit_array_3.drv<63:0>.n286 0.0557941
R4094 hgu_cdac_8bit_array_3.drv<63:0>.n286 hgu_cdac_8bit_array_3.drv<63:0>.n285 0.0557941
R4095 hgu_cdac_8bit_array_3.drv<63:0>.n285 hgu_cdac_8bit_array_3.drv<63:0>.n284 0.0557941
R4096 hgu_cdac_8bit_array_3.drv<63:0>.n297 hgu_cdac_8bit_array_3.drv<63:0>.n296 0.0557941
R4097 hgu_cdac_8bit_array_3.drv<63:0>.n296 hgu_cdac_8bit_array_3.drv<63:0>.n295 0.0557941
R4098 hgu_cdac_8bit_array_3.drv<63:0>.n295 hgu_cdac_8bit_array_3.drv<63:0>.n294 0.0557941
R4099 hgu_cdac_8bit_array_3.drv<63:0>.n294 hgu_cdac_8bit_array_3.drv<63:0>.n293 0.0557941
R4100 hgu_cdac_8bit_array_3.drv<63:0>.n293 hgu_cdac_8bit_array_3.drv<63:0>.n292 0.0557941
R4101 hgu_cdac_8bit_array_3.drv<63:0>.n322 hgu_cdac_8bit_array_3.drv<63:0>.n321 0.0557941
R4102 hgu_cdac_8bit_array_3.drv<63:0>.n321 hgu_cdac_8bit_array_3.drv<63:0>.n320 0.0557941
R4103 hgu_cdac_8bit_array_3.drv<63:0>.n320 hgu_cdac_8bit_array_3.drv<63:0>.n319 0.0557941
R4104 hgu_cdac_8bit_array_3.drv<63:0>.n319 hgu_cdac_8bit_array_3.drv<63:0>.n318 0.0557941
R4105 hgu_cdac_8bit_array_3.drv<63:0>.n318 hgu_cdac_8bit_array_3.drv<63:0>.n317 0.0557941
R4106 hgu_cdac_8bit_array_3.drv<63:0>.n340 hgu_cdac_8bit_array_3.drv<63:0>.n339 0.0557941
R4107 hgu_cdac_8bit_array_3.drv<63:0>.n339 hgu_cdac_8bit_array_3.drv<63:0>.n338 0.0557941
R4108 hgu_cdac_8bit_array_3.drv<63:0>.n338 hgu_cdac_8bit_array_3.drv<63:0>.n337 0.0557941
R4109 hgu_cdac_8bit_array_3.drv<63:0>.n337 hgu_cdac_8bit_array_3.drv<63:0>.n336 0.0557941
R4110 hgu_cdac_8bit_array_3.drv<63:0>.n336 hgu_cdac_8bit_array_3.drv<63:0>.n335 0.0557941
R4111 hgu_cdac_8bit_array_3.drv<63:0>.n355 hgu_cdac_8bit_array_3.drv<63:0>.n354 0.0557941
R4112 hgu_cdac_8bit_array_3.drv<63:0>.n354 hgu_cdac_8bit_array_3.drv<63:0>.n353 0.0557941
R4113 hgu_cdac_8bit_array_3.drv<63:0>.n353 hgu_cdac_8bit_array_3.drv<63:0>.n352 0.0557941
R4114 hgu_cdac_8bit_array_3.drv<63:0>.n352 hgu_cdac_8bit_array_3.drv<63:0>.n351 0.0557941
R4115 hgu_cdac_8bit_array_3.drv<63:0>.n351 hgu_cdac_8bit_array_3.drv<63:0>.n350 0.0557941
R4116 hgu_cdac_8bit_array_3.drv<63:0>.n370 hgu_cdac_8bit_array_3.drv<63:0>.n369 0.0557941
R4117 hgu_cdac_8bit_array_3.drv<63:0>.n34 hgu_cdac_8bit_array_3.drv<63:0>.n33 0.0419706
R4118 hgu_cdac_8bit_array_3.drv<63:0>.n39 hgu_cdac_8bit_array_3.drv<63:0>.n38 0.0419706
R4119 hgu_cdac_8bit_array_3.drv<63:0>.n43 hgu_cdac_8bit_array_3.drv<63:0>.n42 0.0419706
R4120 hgu_cdac_8bit_array_3.drv<63:0>.n48 hgu_cdac_8bit_array_3.drv<63:0>.n47 0.0419706
R4121 hgu_cdac_8bit_array_3.drv<63:0>.n52 hgu_cdac_8bit_array_3.drv<63:0>.n51 0.0419706
R4122 hgu_cdac_8bit_array_3.drv<63:0>.n57 hgu_cdac_8bit_array_3.drv<63:0>.n56 0.0419706
R4123 hgu_cdac_8bit_array_3.drv<63:0>.n61 hgu_cdac_8bit_array_3.drv<63:0>.n60 0.0419706
R4124 hgu_cdac_8bit_array_3.drv<63:0>.n66 hgu_cdac_8bit_array_3.drv<63:0>.n65 0.0419706
R4125 hgu_cdac_8bit_array_3.drv<63:0>.n70 hgu_cdac_8bit_array_3.drv<63:0>.n69 0.0419706
R4126 hgu_cdac_8bit_array_3.drv<63:0>.n75 hgu_cdac_8bit_array_3.drv<63:0>.n74 0.0419706
R4127 hgu_cdac_8bit_array_3.drv<63:0>.n79 hgu_cdac_8bit_array_3.drv<63:0>.n78 0.0419706
R4128 hgu_cdac_8bit_array_3.drv<63:0>.n601 hgu_cdac_8bit_array_3.drv<63:0>.n600 0.0419706
R4129 hgu_cdac_8bit_array_3.drv<63:0>.n597 hgu_cdac_8bit_array_3.drv<63:0>.n596 0.0419706
R4130 hgu_cdac_8bit_array_3.drv<63:0>.n592 hgu_cdac_8bit_array_3.drv<63:0>.n591 0.0419706
R4131 hgu_cdac_8bit_array_3.drv<63:0>.n588 hgu_cdac_8bit_array_3.drv<63:0>.n587 0.0419706
R4132 hgu_cdac_8bit_array_3.drv<63:0>.n583 hgu_cdac_8bit_array_3.drv<63:0>.n582 0.0419706
R4133 hgu_cdac_8bit_array_3.drv<63:0>.n579 hgu_cdac_8bit_array_3.drv<63:0>.n578 0.0419706
R4134 hgu_cdac_8bit_array_3.drv<63:0>.n574 hgu_cdac_8bit_array_3.drv<63:0>.n573 0.0419706
R4135 hgu_cdac_8bit_array_3.drv<63:0>.n570 hgu_cdac_8bit_array_3.drv<63:0>.n569 0.0419706
R4136 hgu_cdac_8bit_array_3.drv<63:0>.n565 hgu_cdac_8bit_array_3.drv<63:0>.n564 0.0419706
R4137 hgu_cdac_8bit_array_3.drv<63:0>.n561 hgu_cdac_8bit_array_3.drv<63:0>.n560 0.0419706
R4138 hgu_cdac_8bit_array_3.drv<63:0>.n556 hgu_cdac_8bit_array_3.drv<63:0>.n555 0.0419706
R4139 hgu_cdac_8bit_array_3.drv<63:0>.n552 hgu_cdac_8bit_array_3.drv<63:0>.n551 0.0419706
R4140 hgu_cdac_8bit_array_3.drv<63:0>.n547 hgu_cdac_8bit_array_3.drv<63:0>.n546 0.0419706
R4141 hgu_cdac_8bit_array_3.drv<63:0>.n543 hgu_cdac_8bit_array_3.drv<63:0>.n542 0.0419706
R4142 hgu_cdac_8bit_array_3.drv<63:0>.n538 hgu_cdac_8bit_array_3.drv<63:0>.n537 0.0419706
R4143 hgu_cdac_8bit_array_3.drv<63:0>.n534 hgu_cdac_8bit_array_3.drv<63:0>.n533 0.0419706
R4144 hgu_cdac_8bit_array_3.drv<63:0>.n529 hgu_cdac_8bit_array_3.drv<63:0>.n528 0.0419706
R4145 hgu_cdac_8bit_array_3.drv<63:0>.n525 hgu_cdac_8bit_array_3.drv<63:0>.n524 0.0419706
R4146 hgu_cdac_8bit_array_3.drv<63:0>.n520 hgu_cdac_8bit_array_3.drv<63:0>.n519 0.0419706
R4147 hgu_cdac_8bit_array_3.drv<63:0>.n516 hgu_cdac_8bit_array_3.drv<63:0>.n515 0.0419706
R4148 hgu_cdac_8bit_array_3.drv<63:0>.n511 hgu_cdac_8bit_array_3.drv<63:0>.n510 0.0419706
R4149 hgu_cdac_8bit_array_3.drv<63:0>.n507 hgu_cdac_8bit_array_3.drv<63:0>.n506 0.0419706
R4150 hgu_cdac_8bit_array_3.drv<63:0>.n502 hgu_cdac_8bit_array_3.drv<63:0>.n501 0.0419706
R4151 hgu_cdac_8bit_array_3.drv<63:0>.n501 hgu_cdac_8bit_array_3.drv<63:0>.n500 0.0419706
R4152 hgu_cdac_8bit_array_3.drv<63:0>.n497 hgu_cdac_8bit_array_3.drv<63:0>.n496 0.0419706
R4153 hgu_cdac_8bit_array_3.drv<63:0>.n492 hgu_cdac_8bit_array_3.drv<63:0>.n491 0.0419706
R4154 hgu_cdac_8bit_array_3.drv<63:0>.n488 hgu_cdac_8bit_array_3.drv<63:0>.n487 0.0419706
R4155 hgu_cdac_8bit_array_3.drv<63:0>.n483 hgu_cdac_8bit_array_3.drv<63:0>.n482 0.0419706
R4156 hgu_cdac_8bit_array_3.drv<63:0>.n479 hgu_cdac_8bit_array_3.drv<63:0>.n478 0.0419706
R4157 hgu_cdac_8bit_array_3.drv<63:0>.n474 hgu_cdac_8bit_array_3.drv<63:0>.n473 0.0419706
R4158 hgu_cdac_8bit_array_3.drv<63:0>.n470 hgu_cdac_8bit_array_3.drv<63:0>.n469 0.0419706
R4159 hgu_cdac_8bit_array_3.drv<63:0>.n465 hgu_cdac_8bit_array_3.drv<63:0>.n464 0.0419706
R4160 hgu_cdac_8bit_array_3.drv<63:0>.n461 hgu_cdac_8bit_array_3.drv<63:0>.n460 0.0419706
R4161 hgu_cdac_8bit_array_3.drv<63:0>.n456 hgu_cdac_8bit_array_3.drv<63:0>.n455 0.0419706
R4162 hgu_cdac_8bit_array_3.drv<63:0>.n452 hgu_cdac_8bit_array_3.drv<63:0>.n451 0.0419706
R4163 hgu_cdac_8bit_array_3.drv<63:0>.n447 hgu_cdac_8bit_array_3.drv<63:0>.n446 0.0419706
R4164 hgu_cdac_8bit_array_3.drv<63:0>.n443 hgu_cdac_8bit_array_3.drv<63:0>.n442 0.0419706
R4165 hgu_cdac_8bit_array_3.drv<63:0>.n438 hgu_cdac_8bit_array_3.drv<63:0>.n437 0.0419706
R4166 hgu_cdac_8bit_array_3.drv<63:0>.n434 hgu_cdac_8bit_array_3.drv<63:0>.n433 0.0419706
R4167 hgu_cdac_8bit_array_3.drv<63:0>.n429 hgu_cdac_8bit_array_3.drv<63:0>.n428 0.0419706
R4168 hgu_cdac_8bit_array_3.drv<63:0>.n425 hgu_cdac_8bit_array_3.drv<63:0>.n424 0.0419706
R4169 hgu_cdac_8bit_array_3.drv<63:0>.n420 hgu_cdac_8bit_array_3.drv<63:0>.n419 0.0419706
R4170 hgu_cdac_8bit_array_3.drv<63:0>.n416 hgu_cdac_8bit_array_3.drv<63:0>.n415 0.0419706
R4171 hgu_cdac_8bit_array_3.drv<63:0>.n411 hgu_cdac_8bit_array_3.drv<63:0>.n410 0.0419706
R4172 hgu_cdac_8bit_array_3.drv<63:0>.n407 hgu_cdac_8bit_array_3.drv<63:0>.n406 0.0419706
R4173 hgu_cdac_8bit_array_3.drv<63:0>.n402 hgu_cdac_8bit_array_3.drv<63:0>.n401 0.0419706
R4174 hgu_cdac_8bit_array_3.drv<63:0>.n398 hgu_cdac_8bit_array_3.drv<63:0>.n397 0.0419706
R4175 hgu_cdac_8bit_array_3.drv<63:0>.n393 hgu_cdac_8bit_array_3.drv<63:0>.n392 0.0419706
R4176 hgu_cdac_8bit_array_3.drv<63:0>.n389 hgu_cdac_8bit_array_3.drv<63:0>.n388 0.0419706
R4177 hgu_cdac_8bit_array_3.drv<63:0>.n384 hgu_cdac_8bit_array_3.drv<63:0>.n383 0.0419706
R4178 hgu_cdac_8bit_array_3.drv<63:0>.n380 hgu_cdac_8bit_array_3.drv<63:0>.n379 0.0419706
R4179 hgu_cdac_8bit_array_3.drv<63:0>.n375 hgu_cdac_8bit_array_3.drv<63:0>.n374 0.0419706
R4180 hgu_cdac_8bit_array_3.drv<63:0>.n316 hgu_cdac_8bit_array_3.drv<63:0>.n315 0.0278438
R4181 hgu_cdac_8bit_array_3.drv<63:0>.n366 hgu_cdac_8bit_array_3.drv<63:0>.n362 0.0180781
R4182 hgu_cdac_8bit_array_3.drv<63:0>.n368 hgu_cdac_8bit_array_3.drv<63:0>.n366 0.0180781
R4183 hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_8bit_array_3.drv<63:0>.n81 0.0157059
R4184 hgu_cdac_8bit_array_3.drv<63:0>.n40 hgu_cdac_8bit_array_3.drv<63:0>.n39 0.0143235
R4185 hgu_cdac_8bit_array_3.drv<63:0>.n42 hgu_cdac_8bit_array_3.drv<63:0>.n41 0.0143235
R4186 hgu_cdac_8bit_array_3.drv<63:0>.n49 hgu_cdac_8bit_array_3.drv<63:0>.n48 0.0143235
R4187 hgu_cdac_8bit_array_3.drv<63:0>.n51 hgu_cdac_8bit_array_3.drv<63:0>.n50 0.0143235
R4188 hgu_cdac_8bit_array_3.drv<63:0>.n58 hgu_cdac_8bit_array_3.drv<63:0>.n57 0.0143235
R4189 hgu_cdac_8bit_array_3.drv<63:0>.n60 hgu_cdac_8bit_array_3.drv<63:0>.n59 0.0143235
R4190 hgu_cdac_8bit_array_3.drv<63:0>.n67 hgu_cdac_8bit_array_3.drv<63:0>.n66 0.0143235
R4191 hgu_cdac_8bit_array_3.drv<63:0>.n69 hgu_cdac_8bit_array_3.drv<63:0>.n68 0.0143235
R4192 hgu_cdac_8bit_array_3.drv<63:0>.n76 hgu_cdac_8bit_array_3.drv<63:0>.n75 0.0143235
R4193 hgu_cdac_8bit_array_3.drv<63:0>.n78 hgu_cdac_8bit_array_3.drv<63:0>.n77 0.0143235
R4194 hgu_cdac_8bit_array_3.drv<63:0>.n600 hgu_cdac_8bit_array_3.drv<63:0>.n599 0.0143235
R4195 hgu_cdac_8bit_array_3.drv<63:0>.n598 hgu_cdac_8bit_array_3.drv<63:0>.n597 0.0143235
R4196 hgu_cdac_8bit_array_3.drv<63:0>.n591 hgu_cdac_8bit_array_3.drv<63:0>.n590 0.0143235
R4197 hgu_cdac_8bit_array_3.drv<63:0>.n589 hgu_cdac_8bit_array_3.drv<63:0>.n588 0.0143235
R4198 hgu_cdac_8bit_array_3.drv<63:0>.n582 hgu_cdac_8bit_array_3.drv<63:0>.n581 0.0143235
R4199 hgu_cdac_8bit_array_3.drv<63:0>.n580 hgu_cdac_8bit_array_3.drv<63:0>.n579 0.0143235
R4200 hgu_cdac_8bit_array_3.drv<63:0>.n573 hgu_cdac_8bit_array_3.drv<63:0>.n572 0.0143235
R4201 hgu_cdac_8bit_array_3.drv<63:0>.n571 hgu_cdac_8bit_array_3.drv<63:0>.n570 0.0143235
R4202 hgu_cdac_8bit_array_3.drv<63:0>.n564 hgu_cdac_8bit_array_3.drv<63:0>.n563 0.0143235
R4203 hgu_cdac_8bit_array_3.drv<63:0>.n562 hgu_cdac_8bit_array_3.drv<63:0>.n561 0.0143235
R4204 hgu_cdac_8bit_array_3.drv<63:0>.n555 hgu_cdac_8bit_array_3.drv<63:0>.n554 0.0143235
R4205 hgu_cdac_8bit_array_3.drv<63:0>.n553 hgu_cdac_8bit_array_3.drv<63:0>.n552 0.0143235
R4206 hgu_cdac_8bit_array_3.drv<63:0>.n546 hgu_cdac_8bit_array_3.drv<63:0>.n545 0.0143235
R4207 hgu_cdac_8bit_array_3.drv<63:0>.n544 hgu_cdac_8bit_array_3.drv<63:0>.n543 0.0143235
R4208 hgu_cdac_8bit_array_3.drv<63:0>.n537 hgu_cdac_8bit_array_3.drv<63:0>.n536 0.0143235
R4209 hgu_cdac_8bit_array_3.drv<63:0>.n535 hgu_cdac_8bit_array_3.drv<63:0>.n534 0.0143235
R4210 hgu_cdac_8bit_array_3.drv<63:0>.n528 hgu_cdac_8bit_array_3.drv<63:0>.n527 0.0143235
R4211 hgu_cdac_8bit_array_3.drv<63:0>.n526 hgu_cdac_8bit_array_3.drv<63:0>.n525 0.0143235
R4212 hgu_cdac_8bit_array_3.drv<63:0>.n519 hgu_cdac_8bit_array_3.drv<63:0>.n518 0.0143235
R4213 hgu_cdac_8bit_array_3.drv<63:0>.n517 hgu_cdac_8bit_array_3.drv<63:0>.n516 0.0143235
R4214 hgu_cdac_8bit_array_3.drv<63:0>.n510 hgu_cdac_8bit_array_3.drv<63:0>.n509 0.0143235
R4215 hgu_cdac_8bit_array_3.drv<63:0>.n508 hgu_cdac_8bit_array_3.drv<63:0>.n507 0.0143235
R4216 hgu_cdac_8bit_array_3.drv<63:0>.n503 hgu_cdac_8bit_array_3.drv<63:0>.n502 0.0143235
R4217 hgu_cdac_8bit_array_3.drv<63:0>.n500 hgu_cdac_8bit_array_3.drv<63:0>.n499 0.0143235
R4218 hgu_cdac_8bit_array_3.drv<63:0>.n498 hgu_cdac_8bit_array_3.drv<63:0>.n497 0.0143235
R4219 hgu_cdac_8bit_array_3.drv<63:0>.n491 hgu_cdac_8bit_array_3.drv<63:0>.n490 0.0143235
R4220 hgu_cdac_8bit_array_3.drv<63:0>.n489 hgu_cdac_8bit_array_3.drv<63:0>.n488 0.0143235
R4221 hgu_cdac_8bit_array_3.drv<63:0>.n482 hgu_cdac_8bit_array_3.drv<63:0>.n481 0.0143235
R4222 hgu_cdac_8bit_array_3.drv<63:0>.n480 hgu_cdac_8bit_array_3.drv<63:0>.n479 0.0143235
R4223 hgu_cdac_8bit_array_3.drv<63:0>.n473 hgu_cdac_8bit_array_3.drv<63:0>.n472 0.0143235
R4224 hgu_cdac_8bit_array_3.drv<63:0>.n471 hgu_cdac_8bit_array_3.drv<63:0>.n470 0.0143235
R4225 hgu_cdac_8bit_array_3.drv<63:0>.n464 hgu_cdac_8bit_array_3.drv<63:0>.n463 0.0143235
R4226 hgu_cdac_8bit_array_3.drv<63:0>.n462 hgu_cdac_8bit_array_3.drv<63:0>.n461 0.0143235
R4227 hgu_cdac_8bit_array_3.drv<63:0>.n455 hgu_cdac_8bit_array_3.drv<63:0>.n454 0.0143235
R4228 hgu_cdac_8bit_array_3.drv<63:0>.n453 hgu_cdac_8bit_array_3.drv<63:0>.n452 0.0143235
R4229 hgu_cdac_8bit_array_3.drv<63:0>.n446 hgu_cdac_8bit_array_3.drv<63:0>.n445 0.0143235
R4230 hgu_cdac_8bit_array_3.drv<63:0>.n444 hgu_cdac_8bit_array_3.drv<63:0>.n443 0.0143235
R4231 hgu_cdac_8bit_array_3.drv<63:0>.n437 hgu_cdac_8bit_array_3.drv<63:0>.n436 0.0143235
R4232 hgu_cdac_8bit_array_3.drv<63:0>.n435 hgu_cdac_8bit_array_3.drv<63:0>.n434 0.0143235
R4233 hgu_cdac_8bit_array_3.drv<63:0>.n428 hgu_cdac_8bit_array_3.drv<63:0>.n427 0.0143235
R4234 hgu_cdac_8bit_array_3.drv<63:0>.n426 hgu_cdac_8bit_array_3.drv<63:0>.n425 0.0143235
R4235 hgu_cdac_8bit_array_3.drv<63:0>.n419 hgu_cdac_8bit_array_3.drv<63:0>.n418 0.0143235
R4236 hgu_cdac_8bit_array_3.drv<63:0>.n417 hgu_cdac_8bit_array_3.drv<63:0>.n416 0.0143235
R4237 hgu_cdac_8bit_array_3.drv<63:0>.n410 hgu_cdac_8bit_array_3.drv<63:0>.n409 0.0143235
R4238 hgu_cdac_8bit_array_3.drv<63:0>.n408 hgu_cdac_8bit_array_3.drv<63:0>.n407 0.0143235
R4239 hgu_cdac_8bit_array_3.drv<63:0>.n401 hgu_cdac_8bit_array_3.drv<63:0>.n400 0.0143235
R4240 hgu_cdac_8bit_array_3.drv<63:0>.n399 hgu_cdac_8bit_array_3.drv<63:0>.n398 0.0143235
R4241 hgu_cdac_8bit_array_3.drv<63:0>.n392 hgu_cdac_8bit_array_3.drv<63:0>.n391 0.0143235
R4242 hgu_cdac_8bit_array_3.drv<63:0>.n390 hgu_cdac_8bit_array_3.drv<63:0>.n389 0.0143235
R4243 hgu_cdac_8bit_array_3.drv<63:0>.n383 hgu_cdac_8bit_array_3.drv<63:0>.n382 0.0143235
R4244 hgu_cdac_8bit_array_3.drv<63:0>.n381 hgu_cdac_8bit_array_3.drv<63:0>.n380 0.0143235
R4245 d<5>.n1 d<5>.n0 77.1205
R4246 d<5>.n2 d<5>.n1 77.1205
R4247 d<5>.n3 d<5>.n2 77.1205
R4248 d<5>.n4 d<5>.n3 77.1205
R4249 d<5>.n5 d<5>.n4 77.1205
R4250 d<5>.n6 d<5>.n5 77.1205
R4251 d<5>.n7 d<5>.n6 77.1205
R4252 d<5>.n8 d<5>.n7 77.1205
R4253 d<5>.n9 d<5>.n8 77.1205
R4254 d<5>.n10 d<5>.n9 77.1205
R4255 d<5>.n11 d<5>.n10 77.1205
R4256 d<5>.n12 d<5>.n11 77.1205
R4257 d<5>.n13 d<5>.n12 77.1205
R4258 d<5>.n14 d<5>.n13 77.1205
R4259 d<5>.n15 d<5>.n14 77.1205
R4260 d<5>.n16 d<5>.n15 77.1205
R4261 d<5>.n17 d<5>.n16 77.1205
R4262 d<5>.n18 d<5>.n17 77.1205
R4263 d<5>.n19 d<5>.n18 77.1205
R4264 d<5>.n20 d<5>.n19 77.1205
R4265 d<5>.n21 d<5>.n20 77.1205
R4266 d<5>.n22 d<5>.n21 77.1205
R4267 d<5>.n23 d<5>.n22 77.1205
R4268 d<5>.n24 d<5>.n23 77.1205
R4269 d<5>.n25 d<5>.n24 77.1205
R4270 d<5>.n26 d<5>.n25 77.1205
R4271 d<5>.n27 d<5>.n26 77.1205
R4272 d<5>.n28 d<5>.n27 77.1205
R4273 d<5>.n29 d<5>.n28 77.1205
R4274 d<5>.n30 d<5>.n29 77.1205
R4275 d<5>.n31 d<5>.n30 77.1205
R4276 d<5>.n0 d<5>.t17 69.5462
R4277 d<5>.n1 d<5>.t58 69.5462
R4278 d<5>.n2 d<5>.t50 69.5462
R4279 d<5>.n3 d<5>.t44 69.5462
R4280 d<5>.n4 d<5>.t19 69.5462
R4281 d<5>.n5 d<5>.t40 69.5462
R4282 d<5>.n6 d<5>.t15 69.5462
R4283 d<5>.n7 d<5>.t24 69.5462
R4284 d<5>.n8 d<5>.t61 69.5462
R4285 d<5>.n9 d<5>.t41 69.5462
R4286 d<5>.n10 d<5>.t32 69.5462
R4287 d<5>.n11 d<5>.t7 69.5462
R4288 d<5>.n12 d<5>.t0 69.5462
R4289 d<5>.n13 d<5>.t20 69.5462
R4290 d<5>.n14 d<5>.t9 69.5462
R4291 d<5>.n15 d<5>.t52 69.5462
R4292 d<5>.n16 d<5>.t29 69.5462
R4293 d<5>.n17 d<5>.t21 69.5462
R4294 d<5>.n18 d<5>.t12 69.5462
R4295 d<5>.n19 d<5>.t54 69.5462
R4296 d<5>.n20 d<5>.t30 69.5462
R4297 d<5>.n21 d<5>.t63 69.5462
R4298 d<5>.n22 d<5>.t57 69.5462
R4299 d<5>.n23 d<5>.t35 69.5462
R4300 d<5>.n24 d<5>.t8 69.5462
R4301 d<5>.n25 d<5>.t2 69.5462
R4302 d<5>.n26 d<5>.t43 69.5462
R4303 d<5>.n27 d<5>.t37 69.5462
R4304 d<5>.n28 d<5>.t4 69.5462
R4305 d<5>.n29 d<5>.t47 69.5462
R4306 d<5>.n30 d<5>.t23 69.5462
R4307 d<5>.n31 d<5>.t60 69.5462
R4308 d<5>.n0 d<5>.t31 53.0205
R4309 d<5>.n1 d<5>.t6 53.0205
R4310 d<5>.n2 d<5>.t62 53.0205
R4311 d<5>.n3 d<5>.t56 53.0205
R4312 d<5>.n4 d<5>.t33 53.0205
R4313 d<5>.n5 d<5>.t51 53.0205
R4314 d<5>.n6 d<5>.t28 53.0205
R4315 d<5>.n7 d<5>.t39 53.0205
R4316 d<5>.n8 d<5>.t11 53.0205
R4317 d<5>.n9 d<5>.t53 53.0205
R4318 d<5>.n10 d<5>.t46 53.0205
R4319 d<5>.n11 d<5>.t22 53.0205
R4320 d<5>.n12 d<5>.t14 53.0205
R4321 d<5>.n13 d<5>.t34 53.0205
R4322 d<5>.n14 d<5>.t26 53.0205
R4323 d<5>.n15 d<5>.t1 53.0205
R4324 d<5>.n16 d<5>.t42 53.0205
R4325 d<5>.n17 d<5>.t36 53.0205
R4326 d<5>.n18 d<5>.t27 53.0205
R4327 d<5>.n19 d<5>.t3 53.0205
R4328 d<5>.n20 d<5>.t45 53.0205
R4329 d<5>.n21 d<5>.t13 53.0205
R4330 d<5>.n22 d<5>.t5 53.0205
R4331 d<5>.n23 d<5>.t48 53.0205
R4332 d<5>.n24 d<5>.t25 53.0205
R4333 d<5>.n25 d<5>.t16 53.0205
R4334 d<5>.n26 d<5>.t55 53.0205
R4335 d<5>.n27 d<5>.t49 53.0205
R4336 d<5>.n28 d<5>.t18 53.0205
R4337 d<5>.n29 d<5>.t59 53.0205
R4338 d<5>.n30 d<5>.t38 53.0205
R4339 d<5>.n31 d<5>.t10 53.0205
R4340 d<5> d<5>.n31 21.088
R4341 hgu_cdac_8bit_array_3.drv<31:0>.n32 hgu_cdac_8bit_array_3.drv<31:0>.t48 41.4291
R4342 hgu_cdac_8bit_array_3.drv<31:0>.n32 hgu_cdac_8bit_array_3.drv<31:0>.t14 41.4291
R4343 hgu_cdac_8bit_array_3.drv<31:0>.n62 hgu_cdac_8bit_array_3.drv<31:0>.t56 41.4291
R4344 hgu_cdac_8bit_array_3.drv<31:0>.n62 hgu_cdac_8bit_array_3.drv<31:0>.t6 41.4291
R4345 hgu_cdac_8bit_array_3.drv<31:0>.n46 hgu_cdac_8bit_array_3.drv<31:0>.t62 41.4291
R4346 hgu_cdac_8bit_array_3.drv<31:0>.n46 hgu_cdac_8bit_array_3.drv<31:0>.t57 41.4291
R4347 hgu_cdac_8bit_array_3.drv<31:0>.n44 hgu_cdac_8bit_array_3.drv<31:0>.t55 41.4291
R4348 hgu_cdac_8bit_array_3.drv<31:0>.n44 hgu_cdac_8bit_array_3.drv<31:0>.t60 41.4291
R4349 hgu_cdac_8bit_array_3.drv<31:0>.n50 hgu_cdac_8bit_array_3.drv<31:0>.t10 41.4291
R4350 hgu_cdac_8bit_array_3.drv<31:0>.n50 hgu_cdac_8bit_array_3.drv<31:0>.t51 41.4291
R4351 hgu_cdac_8bit_array_3.drv<31:0>.n29 hgu_cdac_8bit_array_3.drv<31:0>.t4 41.4291
R4352 hgu_cdac_8bit_array_3.drv<31:0>.n29 hgu_cdac_8bit_array_3.drv<31:0>.t59 41.4291
R4353 hgu_cdac_8bit_array_3.drv<31:0>.n258 hgu_cdac_8bit_array_3.drv<31:0>.t52 41.4291
R4354 hgu_cdac_8bit_array_3.drv<31:0>.n258 hgu_cdac_8bit_array_3.drv<31:0>.t5 41.4291
R4355 hgu_cdac_8bit_array_3.drv<31:0>.n256 hgu_cdac_8bit_array_3.drv<31:0>.t0 41.4291
R4356 hgu_cdac_8bit_array_3.drv<31:0>.n256 hgu_cdac_8bit_array_3.drv<31:0>.t63 41.4291
R4357 hgu_cdac_8bit_array_3.drv<31:0>.n248 hgu_cdac_8bit_array_3.drv<31:0>.t58 41.4291
R4358 hgu_cdac_8bit_array_3.drv<31:0>.n248 hgu_cdac_8bit_array_3.drv<31:0>.t61 41.4291
R4359 hgu_cdac_8bit_array_3.drv<31:0>.n251 hgu_cdac_8bit_array_3.drv<31:0>.t13 41.4291
R4360 hgu_cdac_8bit_array_3.drv<31:0>.n251 hgu_cdac_8bit_array_3.drv<31:0>.t1 41.4291
R4361 hgu_cdac_8bit_array_3.drv<31:0>.n245 hgu_cdac_8bit_array_3.drv<31:0>.t7 41.4291
R4362 hgu_cdac_8bit_array_3.drv<31:0>.n245 hgu_cdac_8bit_array_3.drv<31:0>.t47 41.4291
R4363 hgu_cdac_8bit_array_3.drv<31:0>.n9 hgu_cdac_8bit_array_3.drv<31:0>.t49 41.4291
R4364 hgu_cdac_8bit_array_3.drv<31:0>.n9 hgu_cdac_8bit_array_3.drv<31:0>.t3 41.4291
R4365 hgu_cdac_8bit_array_3.drv<31:0>.n3 hgu_cdac_8bit_array_3.drv<31:0>.t11 41.4291
R4366 hgu_cdac_8bit_array_3.drv<31:0>.n3 hgu_cdac_8bit_array_3.drv<31:0>.t8 41.4291
R4367 hgu_cdac_8bit_array_3.drv<31:0>.n5 hgu_cdac_8bit_array_3.drv<31:0>.t50 41.4291
R4368 hgu_cdac_8bit_array_3.drv<31:0>.n5 hgu_cdac_8bit_array_3.drv<31:0>.t53 41.4291
R4369 hgu_cdac_8bit_array_3.drv<31:0>.n24 hgu_cdac_8bit_array_3.drv<31:0>.t12 41.4291
R4370 hgu_cdac_8bit_array_3.drv<31:0>.n24 hgu_cdac_8bit_array_3.drv<31:0>.t9 41.4291
R4371 hgu_cdac_8bit_array_3.drv<31:0>.n21 hgu_cdac_8bit_array_3.drv<31:0>.t2 41.4291
R4372 hgu_cdac_8bit_array_3.drv<31:0>.n21 hgu_cdac_8bit_array_3.drv<31:0>.t54 41.4291
R4373 hgu_cdac_8bit_array_3.drv<31:0>.n33 hgu_cdac_8bit_array_3.drv<31:0>.t30 34.0065
R4374 hgu_cdac_8bit_array_3.drv<31:0>.n33 hgu_cdac_8bit_array_3.drv<31:0>.t43 34.0065
R4375 hgu_cdac_8bit_array_3.drv<31:0>.n63 hgu_cdac_8bit_array_3.drv<31:0>.t38 34.0065
R4376 hgu_cdac_8bit_array_3.drv<31:0>.n63 hgu_cdac_8bit_array_3.drv<31:0>.t18 34.0065
R4377 hgu_cdac_8bit_array_3.drv<31:0>.n47 hgu_cdac_8bit_array_3.drv<31:0>.t22 34.0065
R4378 hgu_cdac_8bit_array_3.drv<31:0>.n47 hgu_cdac_8bit_array_3.drv<31:0>.t24 34.0065
R4379 hgu_cdac_8bit_array_3.drv<31:0>.n45 hgu_cdac_8bit_array_3.drv<31:0>.t37 34.0065
R4380 hgu_cdac_8bit_array_3.drv<31:0>.n45 hgu_cdac_8bit_array_3.drv<31:0>.t27 34.0065
R4381 hgu_cdac_8bit_array_3.drv<31:0>.n51 hgu_cdac_8bit_array_3.drv<31:0>.t39 34.0065
R4382 hgu_cdac_8bit_array_3.drv<31:0>.n51 hgu_cdac_8bit_array_3.drv<31:0>.t33 34.0065
R4383 hgu_cdac_8bit_array_3.drv<31:0>.n30 hgu_cdac_8bit_array_3.drv<31:0>.t16 34.0065
R4384 hgu_cdac_8bit_array_3.drv<31:0>.n30 hgu_cdac_8bit_array_3.drv<31:0>.t26 34.0065
R4385 hgu_cdac_8bit_array_3.drv<31:0>.n259 hgu_cdac_8bit_array_3.drv<31:0>.t34 34.0065
R4386 hgu_cdac_8bit_array_3.drv<31:0>.n259 hgu_cdac_8bit_array_3.drv<31:0>.t17 34.0065
R4387 hgu_cdac_8bit_array_3.drv<31:0>.n257 hgu_cdac_8bit_array_3.drv<31:0>.t44 34.0065
R4388 hgu_cdac_8bit_array_3.drv<31:0>.n257 hgu_cdac_8bit_array_3.drv<31:0>.t23 34.0065
R4389 hgu_cdac_8bit_array_3.drv<31:0>.n249 hgu_cdac_8bit_array_3.drv<31:0>.t25 34.0065
R4390 hgu_cdac_8bit_array_3.drv<31:0>.n249 hgu_cdac_8bit_array_3.drv<31:0>.t28 34.0065
R4391 hgu_cdac_8bit_array_3.drv<31:0>.n252 hgu_cdac_8bit_array_3.drv<31:0>.t42 34.0065
R4392 hgu_cdac_8bit_array_3.drv<31:0>.n252 hgu_cdac_8bit_array_3.drv<31:0>.t45 34.0065
R4393 hgu_cdac_8bit_array_3.drv<31:0>.n246 hgu_cdac_8bit_array_3.drv<31:0>.t19 34.0065
R4394 hgu_cdac_8bit_array_3.drv<31:0>.n246 hgu_cdac_8bit_array_3.drv<31:0>.t29 34.0065
R4395 hgu_cdac_8bit_array_3.drv<31:0>.n10 hgu_cdac_8bit_array_3.drv<31:0>.t31 34.0065
R4396 hgu_cdac_8bit_array_3.drv<31:0>.n10 hgu_cdac_8bit_array_3.drv<31:0>.t15 34.0065
R4397 hgu_cdac_8bit_array_3.drv<31:0>.n4 hgu_cdac_8bit_array_3.drv<31:0>.t40 34.0065
R4398 hgu_cdac_8bit_array_3.drv<31:0>.n4 hgu_cdac_8bit_array_3.drv<31:0>.t20 34.0065
R4399 hgu_cdac_8bit_array_3.drv<31:0>.n6 hgu_cdac_8bit_array_3.drv<31:0>.t32 34.0065
R4400 hgu_cdac_8bit_array_3.drv<31:0>.n6 hgu_cdac_8bit_array_3.drv<31:0>.t35 34.0065
R4401 hgu_cdac_8bit_array_3.drv<31:0>.n25 hgu_cdac_8bit_array_3.drv<31:0>.t41 34.0065
R4402 hgu_cdac_8bit_array_3.drv<31:0>.n25 hgu_cdac_8bit_array_3.drv<31:0>.t21 34.0065
R4403 hgu_cdac_8bit_array_3.drv<31:0>.n22 hgu_cdac_8bit_array_3.drv<31:0>.t46 34.0065
R4404 hgu_cdac_8bit_array_3.drv<31:0>.n22 hgu_cdac_8bit_array_3.drv<31:0>.t36 34.0065
R4405 hgu_cdac_8bit_array_3.drv<31:0>.n72 hgu_cdac_8bit_array_3.drv<31:0>.n64 10.9368
R4406 hgu_cdac_8bit_array_3.drv<31:0>.n265 hgu_cdac_8bit_array_3.drv<31:0>.n1 10.8469
R4407 hgu_cdac_8bit_array_3.drv<31:0>.n28 hgu_cdac_8bit_array_3.drv<31:0>.n27 10.8445
R4408 hgu_cdac_8bit_array_3.drv<31:0>.n255 hgu_cdac_8bit_array_3.drv<31:0>.n254 10.8414
R4409 hgu_cdac_8bit_array_3.drv<31:0>.n13 hgu_cdac_8bit_array_3.drv<31:0>.n12 10.8285
R4410 hgu_cdac_8bit_array_3.drv<31:0>.n43 hgu_cdac_8bit_array_3.drv<31:0>.n35 10.8239
R4411 hgu_cdac_8bit_array_3.drv<31:0>.n61 hgu_cdac_8bit_array_3.drv<31:0>.n53 10.8235
R4412 hgu_cdac_8bit_array_3.drv<31:0>.n8 hgu_cdac_8bit_array_3.drv<31:0>.n7 0.9906
R4413 hgu_cdac_8bit_array_3.drv<31:0>.n49 hgu_cdac_8bit_array_3.drv<31:0>.n48 0.987754
R4414 hgu_cdac_8bit_array_3.drv<31:0>.n1 hgu_cdac_8bit_array_3.drv<31:0>.n0 0.957599
R4415 hgu_cdac_8bit_array_3.drv<31:0>.n253 hgu_cdac_8bit_array_3.drv<31:0>.n250 0.957397
R4416 hgu_cdac_8bit_array_3.drv<31:0>.n27 hgu_cdac_8bit_array_3.drv<31:0>.n23 0.838862
R4417 hgu_cdac_8bit_array_3.drv<31:0>.n12 hgu_cdac_8bit_array_3.drv<31:0>.n11 0.787138
R4418 hgu_cdac_8bit_array_3.drv<31:0>.n53 hgu_cdac_8bit_array_3.drv<31:0>.n52 0.77316
R4419 hgu_cdac_8bit_array_3.drv<31:0>.n34 hgu_cdac_8bit_array_3.drv<31:0>.n33 0.558205
R4420 hgu_cdac_8bit_array_3.drv<31:0>.n48 hgu_cdac_8bit_array_3.drv<31:0>.n47 0.558205
R4421 hgu_cdac_8bit_array_3.drv<31:0>.n52 hgu_cdac_8bit_array_3.drv<31:0>.n51 0.558205
R4422 hgu_cdac_8bit_array_3.drv<31:0>.n31 hgu_cdac_8bit_array_3.drv<31:0>.n30 0.558205
R4423 hgu_cdac_8bit_array_3.drv<31:0>.n250 hgu_cdac_8bit_array_3.drv<31:0>.n249 0.558205
R4424 hgu_cdac_8bit_array_3.drv<31:0>.n253 hgu_cdac_8bit_array_3.drv<31:0>.n252 0.558205
R4425 hgu_cdac_8bit_array_3.drv<31:0>.n247 hgu_cdac_8bit_array_3.drv<31:0>.n246 0.558205
R4426 hgu_cdac_8bit_array_3.drv<31:0>.n11 hgu_cdac_8bit_array_3.drv<31:0>.n10 0.558205
R4427 hgu_cdac_8bit_array_3.drv<31:0>.n7 hgu_cdac_8bit_array_3.drv<31:0>.n6 0.558205
R4428 hgu_cdac_8bit_array_3.drv<31:0>.n23 hgu_cdac_8bit_array_3.drv<31:0>.n22 0.558205
R4429 hgu_cdac_8bit_array_3.drv<31:0>.n0 hgu_cdac_8bit_array_3.drv<31:0>.n259 0.550852
R4430 hgu_cdac_8bit_array_3.drv<31:0>.n254 hgu_cdac_8bit_array_3.drv<31:0>.n247 0.545759
R4431 hgu_cdac_8bit_array_3.drv<31:0>.n35 hgu_cdac_8bit_array_3.drv<31:0>.n31 0.428333
R4432 hgu_cdac_8bit_array_3.drv<31:0>.n1 hgu_cdac_8bit_array_3.drv<31:0>.n257 0.381734
R4433 hgu_cdac_8bit_array_3.drv<31:0>.n64 hgu_cdac_8bit_array_3.drv<31:0>.n63 0.378057
R4434 hgu_cdac_8bit_array_3.drv<31:0>.n8 hgu_cdac_8bit_array_3.drv<31:0>.n4 0.378057
R4435 hgu_cdac_8bit_array_3.drv<31:0>.n26 hgu_cdac_8bit_array_3.drv<31:0>.n25 0.378057
R4436 hgu_cdac_8bit_array_3.drv<31:0>.n35 hgu_cdac_8bit_array_3.drv<31:0>.n34 0.367988
R4437 hgu_cdac_8bit_array_3.drv<31:0>.n49 hgu_cdac_8bit_array_3.drv<31:0>.n45 0.355999
R4438 hgu_cdac_8bit_array_3.drv<31:0>.n125 hgu_cdac_8bit_array_3.drv<31:0> 0.338468
R4439 hgu_cdac_8bit_array_3.drv<31:0>.n129 hgu_cdac_8bit_array_3.drv<31:0>.n124 0.330451
R4440 hgu_cdac_8bit_array_3.drv<31:0>.n138 hgu_cdac_8bit_array_3.drv<31:0>.n121 0.330451
R4441 hgu_cdac_8bit_array_3.drv<31:0>.n147 hgu_cdac_8bit_array_3.drv<31:0>.n114 0.330451
R4442 hgu_cdac_8bit_array_3.drv<31:0>.n156 hgu_cdac_8bit_array_3.drv<31:0>.n107 0.330451
R4443 hgu_cdac_8bit_array_3.drv<31:0>.n165 hgu_cdac_8bit_array_3.drv<31:0>.n100 0.330451
R4444 hgu_cdac_8bit_array_3.drv<31:0>.n174 hgu_cdac_8bit_array_3.drv<31:0>.n93 0.330451
R4445 hgu_cdac_8bit_array_3.drv<31:0>.n183 hgu_cdac_8bit_array_3.drv<31:0>.n86 0.330451
R4446 hgu_cdac_8bit_array_3.drv<31:0>.n192 hgu_cdac_8bit_array_3.drv<31:0>.n79 0.330451
R4447 hgu_cdac_8bit_array_3.drv<31:0>.n270 hgu_cdac_8bit_array_3.drv<31:0> 0.321667
R4448 hgu_cdac_8bit_array_3.drv<31:0>.n279 hgu_cdac_8bit_array_3.drv<31:0> 0.321667
R4449 hgu_cdac_8bit_array_3.drv<31:0>.n288 hgu_cdac_8bit_array_3.drv<31:0> 0.321667
R4450 hgu_cdac_8bit_array_3.drv<31:0>.n231 hgu_cdac_8bit_array_3.drv<31:0> 0.321667
R4451 hgu_cdac_8bit_array_3.drv<31:0>.n222 hgu_cdac_8bit_array_3.drv<31:0> 0.321667
R4452 hgu_cdac_8bit_array_3.drv<31:0>.n213 hgu_cdac_8bit_array_3.drv<31:0> 0.321667
R4453 hgu_cdac_8bit_array_3.drv<31:0>.n195 hgu_cdac_8bit_array_3.drv<31:0> 0.321667
R4454 hgu_cdac_8bit_array_3.drv<31:0>.n186 hgu_cdac_8bit_array_3.drv<31:0> 0.321667
R4455 hgu_cdac_8bit_array_3.drv<31:0>.n177 hgu_cdac_8bit_array_3.drv<31:0> 0.321667
R4456 hgu_cdac_8bit_array_3.drv<31:0>.n168 hgu_cdac_8bit_array_3.drv<31:0> 0.321667
R4457 hgu_cdac_8bit_array_3.drv<31:0>.n159 hgu_cdac_8bit_array_3.drv<31:0> 0.321667
R4458 hgu_cdac_8bit_array_3.drv<31:0>.n150 hgu_cdac_8bit_array_3.drv<31:0> 0.321667
R4459 hgu_cdac_8bit_array_3.drv<31:0>.n141 hgu_cdac_8bit_array_3.drv<31:0> 0.321667
R4460 hgu_cdac_8bit_array_3.drv<31:0>.n132 hgu_cdac_8bit_array_3.drv<31:0> 0.321667
R4461 hgu_cdac_8bit_array_3.drv<31:0>.n0 hgu_cdac_8bit_array_3.drv<31:0>.n258 0.308208
R4462 hgu_cdac_8bit_array_3.drv<31:0>.n34 hgu_cdac_8bit_array_3.drv<31:0>.n32 0.300856
R4463 hgu_cdac_8bit_array_3.drv<31:0>.n48 hgu_cdac_8bit_array_3.drv<31:0>.n46 0.300856
R4464 hgu_cdac_8bit_array_3.drv<31:0>.n52 hgu_cdac_8bit_array_3.drv<31:0>.n50 0.300856
R4465 hgu_cdac_8bit_array_3.drv<31:0>.n31 hgu_cdac_8bit_array_3.drv<31:0>.n29 0.300856
R4466 hgu_cdac_8bit_array_3.drv<31:0>.n250 hgu_cdac_8bit_array_3.drv<31:0>.n248 0.300856
R4467 hgu_cdac_8bit_array_3.drv<31:0>.n253 hgu_cdac_8bit_array_3.drv<31:0>.n251 0.300856
R4468 hgu_cdac_8bit_array_3.drv<31:0>.n247 hgu_cdac_8bit_array_3.drv<31:0>.n245 0.300856
R4469 hgu_cdac_8bit_array_3.drv<31:0>.n11 hgu_cdac_8bit_array_3.drv<31:0>.n9 0.300856
R4470 hgu_cdac_8bit_array_3.drv<31:0>.n7 hgu_cdac_8bit_array_3.drv<31:0>.n5 0.300856
R4471 hgu_cdac_8bit_array_3.drv<31:0>.n23 hgu_cdac_8bit_array_3.drv<31:0>.n21 0.300856
R4472 hgu_cdac_8bit_array_3.drv<31:0>.n126 hgu_cdac_8bit_array_3.drv<31:0> 0.2966
R4473 hgu_cdac_8bit_array_3.drv<31:0>.n135 hgu_cdac_8bit_array_3.drv<31:0> 0.2966
R4474 hgu_cdac_8bit_array_3.drv<31:0>.n144 hgu_cdac_8bit_array_3.drv<31:0> 0.2966
R4475 hgu_cdac_8bit_array_3.drv<31:0>.n153 hgu_cdac_8bit_array_3.drv<31:0> 0.2966
R4476 hgu_cdac_8bit_array_3.drv<31:0>.n162 hgu_cdac_8bit_array_3.drv<31:0> 0.2966
R4477 hgu_cdac_8bit_array_3.drv<31:0>.n171 hgu_cdac_8bit_array_3.drv<31:0> 0.2966
R4478 hgu_cdac_8bit_array_3.drv<31:0>.n180 hgu_cdac_8bit_array_3.drv<31:0> 0.2966
R4479 hgu_cdac_8bit_array_3.drv<31:0>.n189 hgu_cdac_8bit_array_3.drv<31:0> 0.2966
R4480 hgu_cdac_8bit_array_3.drv<31:0>.n198 hgu_cdac_8bit_array_3.drv<31:0> 0.2966
R4481 hgu_cdac_8bit_array_3.drv<31:0>.n207 hgu_cdac_8bit_array_3.drv<31:0> 0.2966
R4482 hgu_cdac_8bit_array_3.drv<31:0>.n216 hgu_cdac_8bit_array_3.drv<31:0> 0.2966
R4483 hgu_cdac_8bit_array_3.drv<31:0>.n225 hgu_cdac_8bit_array_3.drv<31:0> 0.2966
R4484 hgu_cdac_8bit_array_3.drv<31:0>.n234 hgu_cdac_8bit_array_3.drv<31:0> 0.2966
R4485 hgu_cdac_8bit_array_3.drv<31:0>.n285 hgu_cdac_8bit_array_3.drv<31:0> 0.2966
R4486 hgu_cdac_8bit_array_3.drv<31:0>.n276 hgu_cdac_8bit_array_3.drv<31:0> 0.2966
R4487 hgu_cdac_8bit_array_3.drv<31:0>.n267 hgu_cdac_8bit_array_3.drv<31:0> 0.2966
R4488 hgu_cdac_8bit_array_3.drv<31:0>.n254 hgu_cdac_8bit_array_3.drv<31:0>.n253 0.261276
R4489 hgu_cdac_8bit_array_3.drv<31:0>.n204 hgu_cdac_8bit_array_3.drv<31:0> 0.248033
R4490 hgu_cdac_8bit_array_3.drv<31:0>.n64 hgu_cdac_8bit_array_3.drv<31:0>.n62 0.245708
R4491 hgu_cdac_8bit_array_3.drv<31:0>.n49 hgu_cdac_8bit_array_3.drv<31:0>.n44 0.245708
R4492 hgu_cdac_8bit_array_3.drv<31:0>.n8 hgu_cdac_8bit_array_3.drv<31:0>.n3 0.245708
R4493 hgu_cdac_8bit_array_3.drv<31:0>.n26 hgu_cdac_8bit_array_3.drv<31:0>.n24 0.245708
R4494 hgu_cdac_8bit_array_3.drv<31:0>.n1 hgu_cdac_8bit_array_3.drv<31:0>.n256 0.243985
R4495 hgu_cdac_8bit_array_3.drv<31:0>.n267 hgu_cdac_8bit_array_3.drv<31:0>.n266 0.240665
R4496 hgu_cdac_8bit_array_3.drv<31:0>.n273 hgu_cdac_8bit_array_3.drv<31:0>.n265 0.182836
R4497 hgu_cdac_8bit_array_3.drv<31:0>.n210 hgu_cdac_8bit_array_3.drv<31:0>.n61 0.182836
R4498 hgu_cdac_8bit_array_3.drv<31:0>.n201 hgu_cdac_8bit_array_3.drv<31:0>.n72 0.182836
R4499 hgu_cdac_8bit_array_3.drv<31:0>.n219 hgu_cdac_8bit_array_3.drv<31:0>.n43 0.182836
R4500 hgu_cdac_8bit_array_3.drv<31:0>.n228 hgu_cdac_8bit_array_3.drv<31:0>.n28 0.182836
R4501 hgu_cdac_8bit_array_3.drv<31:0>.n237 hgu_cdac_8bit_array_3.drv<31:0>.n13 0.182836
R4502 hgu_cdac_8bit_array_3.drv<31:0>.n282 hgu_cdac_8bit_array_3.drv<31:0>.n255 0.182836
R4503 hgu_cdac_8bit_array_3.drv<31:0>.n72 hgu_cdac_8bit_array_3.drv<31:0>.n71 0.149114
R4504 hgu_cdac_8bit_array_3.drv<31:0>.n61 hgu_cdac_8bit_array_3.drv<31:0>.n60 0.149114
R4505 hgu_cdac_8bit_array_3.drv<31:0>.n43 hgu_cdac_8bit_array_3.drv<31:0>.n42 0.149114
R4506 hgu_cdac_8bit_array_3.drv<31:0>.n28 hgu_cdac_8bit_array_3.drv<31:0>.n20 0.149114
R4507 hgu_cdac_8bit_array_3.drv<31:0>.n13 hgu_cdac_8bit_array_3.drv<31:0>.n2 0.149114
R4508 hgu_cdac_8bit_array_3.drv<31:0>.n255 hgu_cdac_8bit_array_3.drv<31:0>.n244 0.149114
R4509 hgu_cdac_8bit_array_3.drv<31:0>.n265 hgu_cdac_8bit_array_3.drv<31:0>.n264 0.149114
R4510 hgu_cdac_8bit_array_3.drv<31:0>.n12 hgu_cdac_8bit_array_3.drv<31:0>.n8 0.0766719
R4511 hgu_cdac_8bit_array_3.drv<31:0>.n53 hgu_cdac_8bit_array_3.drv<31:0>.n49 0.0737143
R4512 hgu_cdac_8bit_array_3.drv<31:0>.n129 hgu_cdac_8bit_array_3.drv<31:0>.n128 0.0716912
R4513 hgu_cdac_8bit_array_3.drv<31:0>.n130 hgu_cdac_8bit_array_3.drv<31:0>.n129 0.0716912
R4514 hgu_cdac_8bit_array_3.drv<31:0>.n138 hgu_cdac_8bit_array_3.drv<31:0>.n137 0.0716912
R4515 hgu_cdac_8bit_array_3.drv<31:0>.n139 hgu_cdac_8bit_array_3.drv<31:0>.n138 0.0716912
R4516 hgu_cdac_8bit_array_3.drv<31:0>.n147 hgu_cdac_8bit_array_3.drv<31:0>.n146 0.0716912
R4517 hgu_cdac_8bit_array_3.drv<31:0>.n148 hgu_cdac_8bit_array_3.drv<31:0>.n147 0.0716912
R4518 hgu_cdac_8bit_array_3.drv<31:0>.n156 hgu_cdac_8bit_array_3.drv<31:0>.n155 0.0716912
R4519 hgu_cdac_8bit_array_3.drv<31:0>.n157 hgu_cdac_8bit_array_3.drv<31:0>.n156 0.0716912
R4520 hgu_cdac_8bit_array_3.drv<31:0>.n165 hgu_cdac_8bit_array_3.drv<31:0>.n164 0.0716912
R4521 hgu_cdac_8bit_array_3.drv<31:0>.n166 hgu_cdac_8bit_array_3.drv<31:0>.n165 0.0716912
R4522 hgu_cdac_8bit_array_3.drv<31:0>.n174 hgu_cdac_8bit_array_3.drv<31:0>.n173 0.0716912
R4523 hgu_cdac_8bit_array_3.drv<31:0>.n175 hgu_cdac_8bit_array_3.drv<31:0>.n174 0.0716912
R4524 hgu_cdac_8bit_array_3.drv<31:0>.n183 hgu_cdac_8bit_array_3.drv<31:0>.n182 0.0716912
R4525 hgu_cdac_8bit_array_3.drv<31:0>.n184 hgu_cdac_8bit_array_3.drv<31:0>.n183 0.0716912
R4526 hgu_cdac_8bit_array_3.drv<31:0>.n192 hgu_cdac_8bit_array_3.drv<31:0>.n191 0.0716912
R4527 hgu_cdac_8bit_array_3.drv<31:0>.n193 hgu_cdac_8bit_array_3.drv<31:0>.n192 0.0716912
R4528 hgu_cdac_8bit_array_3.drv<31:0>.n201 hgu_cdac_8bit_array_3.drv<31:0>.n200 0.0716912
R4529 hgu_cdac_8bit_array_3.drv<31:0>.n202 hgu_cdac_8bit_array_3.drv<31:0>.n201 0.0716912
R4530 hgu_cdac_8bit_array_3.drv<31:0>.n210 hgu_cdac_8bit_array_3.drv<31:0>.n209 0.0716912
R4531 hgu_cdac_8bit_array_3.drv<31:0>.n211 hgu_cdac_8bit_array_3.drv<31:0>.n210 0.0716912
R4532 hgu_cdac_8bit_array_3.drv<31:0>.n219 hgu_cdac_8bit_array_3.drv<31:0>.n218 0.0716912
R4533 hgu_cdac_8bit_array_3.drv<31:0>.n220 hgu_cdac_8bit_array_3.drv<31:0>.n219 0.0716912
R4534 hgu_cdac_8bit_array_3.drv<31:0>.n228 hgu_cdac_8bit_array_3.drv<31:0>.n227 0.0716912
R4535 hgu_cdac_8bit_array_3.drv<31:0>.n229 hgu_cdac_8bit_array_3.drv<31:0>.n228 0.0716912
R4536 hgu_cdac_8bit_array_3.drv<31:0>.n237 hgu_cdac_8bit_array_3.drv<31:0>.n236 0.0716912
R4537 hgu_cdac_8bit_array_3.drv<31:0>.n283 hgu_cdac_8bit_array_3.drv<31:0>.n282 0.0716912
R4538 hgu_cdac_8bit_array_3.drv<31:0>.n282 hgu_cdac_8bit_array_3.drv<31:0>.n281 0.0716912
R4539 hgu_cdac_8bit_array_3.drv<31:0>.n274 hgu_cdac_8bit_array_3.drv<31:0>.n273 0.0716912
R4540 hgu_cdac_8bit_array_3.drv<31:0>.n273 hgu_cdac_8bit_array_3.drv<31:0>.n272 0.0716912
R4541 hgu_cdac_8bit_array_3.drv<31:0>.n124 hgu_cdac_8bit_array_3.drv<31:0>.n123 0.0716912
R4542 hgu_cdac_8bit_array_3.drv<31:0>.n121 hgu_cdac_8bit_array_3.drv<31:0>.n120 0.0716912
R4543 hgu_cdac_8bit_array_3.drv<31:0>.n114 hgu_cdac_8bit_array_3.drv<31:0>.n113 0.0716912
R4544 hgu_cdac_8bit_array_3.drv<31:0>.n107 hgu_cdac_8bit_array_3.drv<31:0>.n106 0.0716912
R4545 hgu_cdac_8bit_array_3.drv<31:0>.n100 hgu_cdac_8bit_array_3.drv<31:0>.n99 0.0716912
R4546 hgu_cdac_8bit_array_3.drv<31:0>.n93 hgu_cdac_8bit_array_3.drv<31:0>.n92 0.0716912
R4547 hgu_cdac_8bit_array_3.drv<31:0>.n86 hgu_cdac_8bit_array_3.drv<31:0>.n85 0.0716912
R4548 hgu_cdac_8bit_array_3.drv<31:0>.n79 hgu_cdac_8bit_array_3.drv<31:0>.n78 0.0716912
R4549 hgu_cdac_8bit_array_3.drv<31:0>.n71 hgu_cdac_8bit_array_3.drv<31:0>.n70 0.0716912
R4550 hgu_cdac_8bit_array_3.drv<31:0>.n60 hgu_cdac_8bit_array_3.drv<31:0>.n59 0.0716912
R4551 hgu_cdac_8bit_array_3.drv<31:0>.n42 hgu_cdac_8bit_array_3.drv<31:0>.n41 0.0716912
R4552 hgu_cdac_8bit_array_3.drv<31:0>.n20 hgu_cdac_8bit_array_3.drv<31:0>.n19 0.0716912
R4553 hgu_cdac_8bit_array_3.drv<31:0>.n244 hgu_cdac_8bit_array_3.drv<31:0>.n243 0.0716912
R4554 hgu_cdac_8bit_array_3.drv<31:0>.n264 hgu_cdac_8bit_array_3.drv<31:0>.n263 0.0716912
R4555 hgu_cdac_8bit_array_3.drv<31:0>.n126 hgu_cdac_8bit_array_3.drv<31:0>.n125 0.0665339
R4556 hgu_cdac_8bit_array_3.drv<31:0>.n128 hgu_cdac_8bit_array_3.drv<31:0>.n127 0.0557941
R4557 hgu_cdac_8bit_array_3.drv<31:0>.n131 hgu_cdac_8bit_array_3.drv<31:0>.n130 0.0557941
R4558 hgu_cdac_8bit_array_3.drv<31:0>.n134 hgu_cdac_8bit_array_3.drv<31:0>.n133 0.0557941
R4559 hgu_cdac_8bit_array_3.drv<31:0>.n137 hgu_cdac_8bit_array_3.drv<31:0>.n136 0.0557941
R4560 hgu_cdac_8bit_array_3.drv<31:0>.n140 hgu_cdac_8bit_array_3.drv<31:0>.n139 0.0557941
R4561 hgu_cdac_8bit_array_3.drv<31:0>.n143 hgu_cdac_8bit_array_3.drv<31:0>.n142 0.0557941
R4562 hgu_cdac_8bit_array_3.drv<31:0>.n146 hgu_cdac_8bit_array_3.drv<31:0>.n145 0.0557941
R4563 hgu_cdac_8bit_array_3.drv<31:0>.n149 hgu_cdac_8bit_array_3.drv<31:0>.n148 0.0557941
R4564 hgu_cdac_8bit_array_3.drv<31:0>.n152 hgu_cdac_8bit_array_3.drv<31:0>.n151 0.0557941
R4565 hgu_cdac_8bit_array_3.drv<31:0>.n155 hgu_cdac_8bit_array_3.drv<31:0>.n154 0.0557941
R4566 hgu_cdac_8bit_array_3.drv<31:0>.n158 hgu_cdac_8bit_array_3.drv<31:0>.n157 0.0557941
R4567 hgu_cdac_8bit_array_3.drv<31:0>.n161 hgu_cdac_8bit_array_3.drv<31:0>.n160 0.0557941
R4568 hgu_cdac_8bit_array_3.drv<31:0>.n164 hgu_cdac_8bit_array_3.drv<31:0>.n163 0.0557941
R4569 hgu_cdac_8bit_array_3.drv<31:0>.n167 hgu_cdac_8bit_array_3.drv<31:0>.n166 0.0557941
R4570 hgu_cdac_8bit_array_3.drv<31:0>.n170 hgu_cdac_8bit_array_3.drv<31:0>.n169 0.0557941
R4571 hgu_cdac_8bit_array_3.drv<31:0>.n173 hgu_cdac_8bit_array_3.drv<31:0>.n172 0.0557941
R4572 hgu_cdac_8bit_array_3.drv<31:0>.n176 hgu_cdac_8bit_array_3.drv<31:0>.n175 0.0557941
R4573 hgu_cdac_8bit_array_3.drv<31:0>.n179 hgu_cdac_8bit_array_3.drv<31:0>.n178 0.0557941
R4574 hgu_cdac_8bit_array_3.drv<31:0>.n182 hgu_cdac_8bit_array_3.drv<31:0>.n181 0.0557941
R4575 hgu_cdac_8bit_array_3.drv<31:0>.n185 hgu_cdac_8bit_array_3.drv<31:0>.n184 0.0557941
R4576 hgu_cdac_8bit_array_3.drv<31:0>.n188 hgu_cdac_8bit_array_3.drv<31:0>.n187 0.0557941
R4577 hgu_cdac_8bit_array_3.drv<31:0>.n191 hgu_cdac_8bit_array_3.drv<31:0>.n190 0.0557941
R4578 hgu_cdac_8bit_array_3.drv<31:0>.n194 hgu_cdac_8bit_array_3.drv<31:0>.n193 0.0557941
R4579 hgu_cdac_8bit_array_3.drv<31:0>.n197 hgu_cdac_8bit_array_3.drv<31:0>.n196 0.0557941
R4580 hgu_cdac_8bit_array_3.drv<31:0>.n200 hgu_cdac_8bit_array_3.drv<31:0>.n199 0.0557941
R4581 hgu_cdac_8bit_array_3.drv<31:0>.n203 hgu_cdac_8bit_array_3.drv<31:0>.n202 0.0557941
R4582 hgu_cdac_8bit_array_3.drv<31:0>.n206 hgu_cdac_8bit_array_3.drv<31:0>.n205 0.0557941
R4583 hgu_cdac_8bit_array_3.drv<31:0>.n209 hgu_cdac_8bit_array_3.drv<31:0>.n208 0.0557941
R4584 hgu_cdac_8bit_array_3.drv<31:0>.n212 hgu_cdac_8bit_array_3.drv<31:0>.n211 0.0557941
R4585 hgu_cdac_8bit_array_3.drv<31:0>.n215 hgu_cdac_8bit_array_3.drv<31:0>.n214 0.0557941
R4586 hgu_cdac_8bit_array_3.drv<31:0>.n218 hgu_cdac_8bit_array_3.drv<31:0>.n217 0.0557941
R4587 hgu_cdac_8bit_array_3.drv<31:0>.n221 hgu_cdac_8bit_array_3.drv<31:0>.n220 0.0557941
R4588 hgu_cdac_8bit_array_3.drv<31:0>.n224 hgu_cdac_8bit_array_3.drv<31:0>.n223 0.0557941
R4589 hgu_cdac_8bit_array_3.drv<31:0>.n227 hgu_cdac_8bit_array_3.drv<31:0>.n226 0.0557941
R4590 hgu_cdac_8bit_array_3.drv<31:0>.n230 hgu_cdac_8bit_array_3.drv<31:0>.n229 0.0557941
R4591 hgu_cdac_8bit_array_3.drv<31:0>.n233 hgu_cdac_8bit_array_3.drv<31:0>.n232 0.0557941
R4592 hgu_cdac_8bit_array_3.drv<31:0>.n236 hgu_cdac_8bit_array_3.drv<31:0>.n235 0.0557941
R4593 hgu_cdac_8bit_array_3.drv<31:0>.n290 hgu_cdac_8bit_array_3.drv<31:0>.n289 0.0557941
R4594 hgu_cdac_8bit_array_3.drv<31:0>.n287 hgu_cdac_8bit_array_3.drv<31:0>.n286 0.0557941
R4595 hgu_cdac_8bit_array_3.drv<31:0>.n284 hgu_cdac_8bit_array_3.drv<31:0>.n283 0.0557941
R4596 hgu_cdac_8bit_array_3.drv<31:0>.n281 hgu_cdac_8bit_array_3.drv<31:0>.n280 0.0557941
R4597 hgu_cdac_8bit_array_3.drv<31:0>.n278 hgu_cdac_8bit_array_3.drv<31:0>.n277 0.0557941
R4598 hgu_cdac_8bit_array_3.drv<31:0>.n275 hgu_cdac_8bit_array_3.drv<31:0>.n274 0.0557941
R4599 hgu_cdac_8bit_array_3.drv<31:0>.n272 hgu_cdac_8bit_array_3.drv<31:0>.n271 0.0557941
R4600 hgu_cdac_8bit_array_3.drv<31:0>.n269 hgu_cdac_8bit_array_3.drv<31:0>.n268 0.0557941
R4601 hgu_cdac_8bit_array_3.drv<31:0>.n123 hgu_cdac_8bit_array_3.drv<31:0>.n122 0.0557941
R4602 hgu_cdac_8bit_array_3.drv<31:0>.n116 hgu_cdac_8bit_array_3.drv<31:0>.n115 0.0557941
R4603 hgu_cdac_8bit_array_3.drv<31:0>.n117 hgu_cdac_8bit_array_3.drv<31:0>.n116 0.0557941
R4604 hgu_cdac_8bit_array_3.drv<31:0>.n118 hgu_cdac_8bit_array_3.drv<31:0>.n117 0.0557941
R4605 hgu_cdac_8bit_array_3.drv<31:0>.n119 hgu_cdac_8bit_array_3.drv<31:0>.n118 0.0557941
R4606 hgu_cdac_8bit_array_3.drv<31:0>.n120 hgu_cdac_8bit_array_3.drv<31:0>.n119 0.0557941
R4607 hgu_cdac_8bit_array_3.drv<31:0>.n109 hgu_cdac_8bit_array_3.drv<31:0>.n108 0.0557941
R4608 hgu_cdac_8bit_array_3.drv<31:0>.n110 hgu_cdac_8bit_array_3.drv<31:0>.n109 0.0557941
R4609 hgu_cdac_8bit_array_3.drv<31:0>.n111 hgu_cdac_8bit_array_3.drv<31:0>.n110 0.0557941
R4610 hgu_cdac_8bit_array_3.drv<31:0>.n112 hgu_cdac_8bit_array_3.drv<31:0>.n111 0.0557941
R4611 hgu_cdac_8bit_array_3.drv<31:0>.n113 hgu_cdac_8bit_array_3.drv<31:0>.n112 0.0557941
R4612 hgu_cdac_8bit_array_3.drv<31:0>.n102 hgu_cdac_8bit_array_3.drv<31:0>.n101 0.0557941
R4613 hgu_cdac_8bit_array_3.drv<31:0>.n103 hgu_cdac_8bit_array_3.drv<31:0>.n102 0.0557941
R4614 hgu_cdac_8bit_array_3.drv<31:0>.n104 hgu_cdac_8bit_array_3.drv<31:0>.n103 0.0557941
R4615 hgu_cdac_8bit_array_3.drv<31:0>.n105 hgu_cdac_8bit_array_3.drv<31:0>.n104 0.0557941
R4616 hgu_cdac_8bit_array_3.drv<31:0>.n106 hgu_cdac_8bit_array_3.drv<31:0>.n105 0.0557941
R4617 hgu_cdac_8bit_array_3.drv<31:0>.n95 hgu_cdac_8bit_array_3.drv<31:0>.n94 0.0557941
R4618 hgu_cdac_8bit_array_3.drv<31:0>.n96 hgu_cdac_8bit_array_3.drv<31:0>.n95 0.0557941
R4619 hgu_cdac_8bit_array_3.drv<31:0>.n97 hgu_cdac_8bit_array_3.drv<31:0>.n96 0.0557941
R4620 hgu_cdac_8bit_array_3.drv<31:0>.n98 hgu_cdac_8bit_array_3.drv<31:0>.n97 0.0557941
R4621 hgu_cdac_8bit_array_3.drv<31:0>.n99 hgu_cdac_8bit_array_3.drv<31:0>.n98 0.0557941
R4622 hgu_cdac_8bit_array_3.drv<31:0>.n88 hgu_cdac_8bit_array_3.drv<31:0>.n87 0.0557941
R4623 hgu_cdac_8bit_array_3.drv<31:0>.n89 hgu_cdac_8bit_array_3.drv<31:0>.n88 0.0557941
R4624 hgu_cdac_8bit_array_3.drv<31:0>.n90 hgu_cdac_8bit_array_3.drv<31:0>.n89 0.0557941
R4625 hgu_cdac_8bit_array_3.drv<31:0>.n91 hgu_cdac_8bit_array_3.drv<31:0>.n90 0.0557941
R4626 hgu_cdac_8bit_array_3.drv<31:0>.n92 hgu_cdac_8bit_array_3.drv<31:0>.n91 0.0557941
R4627 hgu_cdac_8bit_array_3.drv<31:0>.n81 hgu_cdac_8bit_array_3.drv<31:0>.n80 0.0557941
R4628 hgu_cdac_8bit_array_3.drv<31:0>.n82 hgu_cdac_8bit_array_3.drv<31:0>.n81 0.0557941
R4629 hgu_cdac_8bit_array_3.drv<31:0>.n83 hgu_cdac_8bit_array_3.drv<31:0>.n82 0.0557941
R4630 hgu_cdac_8bit_array_3.drv<31:0>.n84 hgu_cdac_8bit_array_3.drv<31:0>.n83 0.0557941
R4631 hgu_cdac_8bit_array_3.drv<31:0>.n85 hgu_cdac_8bit_array_3.drv<31:0>.n84 0.0557941
R4632 hgu_cdac_8bit_array_3.drv<31:0>.n74 hgu_cdac_8bit_array_3.drv<31:0>.n73 0.0557941
R4633 hgu_cdac_8bit_array_3.drv<31:0>.n75 hgu_cdac_8bit_array_3.drv<31:0>.n74 0.0557941
R4634 hgu_cdac_8bit_array_3.drv<31:0>.n76 hgu_cdac_8bit_array_3.drv<31:0>.n75 0.0557941
R4635 hgu_cdac_8bit_array_3.drv<31:0>.n77 hgu_cdac_8bit_array_3.drv<31:0>.n76 0.0557941
R4636 hgu_cdac_8bit_array_3.drv<31:0>.n78 hgu_cdac_8bit_array_3.drv<31:0>.n77 0.0557941
R4637 hgu_cdac_8bit_array_3.drv<31:0>.n66 hgu_cdac_8bit_array_3.drv<31:0>.n65 0.0557941
R4638 hgu_cdac_8bit_array_3.drv<31:0>.n67 hgu_cdac_8bit_array_3.drv<31:0>.n66 0.0557941
R4639 hgu_cdac_8bit_array_3.drv<31:0>.n68 hgu_cdac_8bit_array_3.drv<31:0>.n67 0.0557941
R4640 hgu_cdac_8bit_array_3.drv<31:0>.n69 hgu_cdac_8bit_array_3.drv<31:0>.n68 0.0557941
R4641 hgu_cdac_8bit_array_3.drv<31:0>.n70 hgu_cdac_8bit_array_3.drv<31:0>.n69 0.0557941
R4642 hgu_cdac_8bit_array_3.drv<31:0>.n55 hgu_cdac_8bit_array_3.drv<31:0>.n54 0.0557941
R4643 hgu_cdac_8bit_array_3.drv<31:0>.n56 hgu_cdac_8bit_array_3.drv<31:0>.n55 0.0557941
R4644 hgu_cdac_8bit_array_3.drv<31:0>.n57 hgu_cdac_8bit_array_3.drv<31:0>.n56 0.0557941
R4645 hgu_cdac_8bit_array_3.drv<31:0>.n58 hgu_cdac_8bit_array_3.drv<31:0>.n57 0.0557941
R4646 hgu_cdac_8bit_array_3.drv<31:0>.n59 hgu_cdac_8bit_array_3.drv<31:0>.n58 0.0557941
R4647 hgu_cdac_8bit_array_3.drv<31:0>.n37 hgu_cdac_8bit_array_3.drv<31:0>.n36 0.0557941
R4648 hgu_cdac_8bit_array_3.drv<31:0>.n38 hgu_cdac_8bit_array_3.drv<31:0>.n37 0.0557941
R4649 hgu_cdac_8bit_array_3.drv<31:0>.n39 hgu_cdac_8bit_array_3.drv<31:0>.n38 0.0557941
R4650 hgu_cdac_8bit_array_3.drv<31:0>.n40 hgu_cdac_8bit_array_3.drv<31:0>.n39 0.0557941
R4651 hgu_cdac_8bit_array_3.drv<31:0>.n41 hgu_cdac_8bit_array_3.drv<31:0>.n40 0.0557941
R4652 hgu_cdac_8bit_array_3.drv<31:0>.n15 hgu_cdac_8bit_array_3.drv<31:0>.n14 0.0557941
R4653 hgu_cdac_8bit_array_3.drv<31:0>.n16 hgu_cdac_8bit_array_3.drv<31:0>.n15 0.0557941
R4654 hgu_cdac_8bit_array_3.drv<31:0>.n17 hgu_cdac_8bit_array_3.drv<31:0>.n16 0.0557941
R4655 hgu_cdac_8bit_array_3.drv<31:0>.n18 hgu_cdac_8bit_array_3.drv<31:0>.n17 0.0557941
R4656 hgu_cdac_8bit_array_3.drv<31:0>.n19 hgu_cdac_8bit_array_3.drv<31:0>.n18 0.0557941
R4657 hgu_cdac_8bit_array_3.drv<31:0>.n243 hgu_cdac_8bit_array_3.drv<31:0>.n242 0.0557941
R4658 hgu_cdac_8bit_array_3.drv<31:0>.n242 hgu_cdac_8bit_array_3.drv<31:0>.n241 0.0557941
R4659 hgu_cdac_8bit_array_3.drv<31:0>.n241 hgu_cdac_8bit_array_3.drv<31:0>.n240 0.0557941
R4660 hgu_cdac_8bit_array_3.drv<31:0>.n240 hgu_cdac_8bit_array_3.drv<31:0>.n239 0.0557941
R4661 hgu_cdac_8bit_array_3.drv<31:0>.n239 hgu_cdac_8bit_array_3.drv<31:0>.n238 0.0557941
R4662 hgu_cdac_8bit_array_3.drv<31:0>.n263 hgu_cdac_8bit_array_3.drv<31:0>.n262 0.0557941
R4663 hgu_cdac_8bit_array_3.drv<31:0>.n262 hgu_cdac_8bit_array_3.drv<31:0>.n261 0.0557941
R4664 hgu_cdac_8bit_array_3.drv<31:0>.n261 hgu_cdac_8bit_array_3.drv<31:0>.n260 0.0557941
R4665 hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_8bit_array_3.drv<31:0>.n290 0.0544118
R4666 hgu_cdac_8bit_array_3.drv<31:0>.n27 hgu_cdac_8bit_array_3.drv<31:0>.n26 0.0532344
R4667 hgu_cdac_8bit_array_3.drv<31:0>.n127 hgu_cdac_8bit_array_3.drv<31:0>.n126 0.0419706
R4668 hgu_cdac_8bit_array_3.drv<31:0>.n132 hgu_cdac_8bit_array_3.drv<31:0>.n131 0.0419706
R4669 hgu_cdac_8bit_array_3.drv<31:0>.n136 hgu_cdac_8bit_array_3.drv<31:0>.n135 0.0419706
R4670 hgu_cdac_8bit_array_3.drv<31:0>.n141 hgu_cdac_8bit_array_3.drv<31:0>.n140 0.0419706
R4671 hgu_cdac_8bit_array_3.drv<31:0>.n145 hgu_cdac_8bit_array_3.drv<31:0>.n144 0.0419706
R4672 hgu_cdac_8bit_array_3.drv<31:0>.n150 hgu_cdac_8bit_array_3.drv<31:0>.n149 0.0419706
R4673 hgu_cdac_8bit_array_3.drv<31:0>.n154 hgu_cdac_8bit_array_3.drv<31:0>.n153 0.0419706
R4674 hgu_cdac_8bit_array_3.drv<31:0>.n159 hgu_cdac_8bit_array_3.drv<31:0>.n158 0.0419706
R4675 hgu_cdac_8bit_array_3.drv<31:0>.n163 hgu_cdac_8bit_array_3.drv<31:0>.n162 0.0419706
R4676 hgu_cdac_8bit_array_3.drv<31:0>.n168 hgu_cdac_8bit_array_3.drv<31:0>.n167 0.0419706
R4677 hgu_cdac_8bit_array_3.drv<31:0>.n172 hgu_cdac_8bit_array_3.drv<31:0>.n171 0.0419706
R4678 hgu_cdac_8bit_array_3.drv<31:0>.n177 hgu_cdac_8bit_array_3.drv<31:0>.n176 0.0419706
R4679 hgu_cdac_8bit_array_3.drv<31:0>.n181 hgu_cdac_8bit_array_3.drv<31:0>.n180 0.0419706
R4680 hgu_cdac_8bit_array_3.drv<31:0>.n186 hgu_cdac_8bit_array_3.drv<31:0>.n185 0.0419706
R4681 hgu_cdac_8bit_array_3.drv<31:0>.n190 hgu_cdac_8bit_array_3.drv<31:0>.n189 0.0419706
R4682 hgu_cdac_8bit_array_3.drv<31:0>.n195 hgu_cdac_8bit_array_3.drv<31:0>.n194 0.0419706
R4683 hgu_cdac_8bit_array_3.drv<31:0>.n199 hgu_cdac_8bit_array_3.drv<31:0>.n198 0.0419706
R4684 hgu_cdac_8bit_array_3.drv<31:0>.n204 hgu_cdac_8bit_array_3.drv<31:0>.n203 0.0419706
R4685 hgu_cdac_8bit_array_3.drv<31:0>.n208 hgu_cdac_8bit_array_3.drv<31:0>.n207 0.0419706
R4686 hgu_cdac_8bit_array_3.drv<31:0>.n213 hgu_cdac_8bit_array_3.drv<31:0>.n212 0.0419706
R4687 hgu_cdac_8bit_array_3.drv<31:0>.n217 hgu_cdac_8bit_array_3.drv<31:0>.n216 0.0419706
R4688 hgu_cdac_8bit_array_3.drv<31:0>.n222 hgu_cdac_8bit_array_3.drv<31:0>.n221 0.0419706
R4689 hgu_cdac_8bit_array_3.drv<31:0>.n226 hgu_cdac_8bit_array_3.drv<31:0>.n225 0.0419706
R4690 hgu_cdac_8bit_array_3.drv<31:0>.n231 hgu_cdac_8bit_array_3.drv<31:0>.n230 0.0419706
R4691 hgu_cdac_8bit_array_3.drv<31:0>.n235 hgu_cdac_8bit_array_3.drv<31:0>.n234 0.0419706
R4692 hgu_cdac_8bit_array_3.drv<31:0>.n289 hgu_cdac_8bit_array_3.drv<31:0>.n288 0.0419706
R4693 hgu_cdac_8bit_array_3.drv<31:0>.n285 hgu_cdac_8bit_array_3.drv<31:0>.n284 0.0419706
R4694 hgu_cdac_8bit_array_3.drv<31:0>.n280 hgu_cdac_8bit_array_3.drv<31:0>.n279 0.0419706
R4695 hgu_cdac_8bit_array_3.drv<31:0>.n276 hgu_cdac_8bit_array_3.drv<31:0>.n275 0.0419706
R4696 hgu_cdac_8bit_array_3.drv<31:0>.n271 hgu_cdac_8bit_array_3.drv<31:0>.n270 0.0419706
R4697 hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_8bit_array_3.drv<31:0>.n237 0.0177794
R4698 hgu_cdac_8bit_array_3.drv<31:0>.n133 hgu_cdac_8bit_array_3.drv<31:0>.n132 0.0143235
R4699 hgu_cdac_8bit_array_3.drv<31:0>.n135 hgu_cdac_8bit_array_3.drv<31:0>.n134 0.0143235
R4700 hgu_cdac_8bit_array_3.drv<31:0>.n142 hgu_cdac_8bit_array_3.drv<31:0>.n141 0.0143235
R4701 hgu_cdac_8bit_array_3.drv<31:0>.n144 hgu_cdac_8bit_array_3.drv<31:0>.n143 0.0143235
R4702 hgu_cdac_8bit_array_3.drv<31:0>.n151 hgu_cdac_8bit_array_3.drv<31:0>.n150 0.0143235
R4703 hgu_cdac_8bit_array_3.drv<31:0>.n153 hgu_cdac_8bit_array_3.drv<31:0>.n152 0.0143235
R4704 hgu_cdac_8bit_array_3.drv<31:0>.n160 hgu_cdac_8bit_array_3.drv<31:0>.n159 0.0143235
R4705 hgu_cdac_8bit_array_3.drv<31:0>.n162 hgu_cdac_8bit_array_3.drv<31:0>.n161 0.0143235
R4706 hgu_cdac_8bit_array_3.drv<31:0>.n169 hgu_cdac_8bit_array_3.drv<31:0>.n168 0.0143235
R4707 hgu_cdac_8bit_array_3.drv<31:0>.n171 hgu_cdac_8bit_array_3.drv<31:0>.n170 0.0143235
R4708 hgu_cdac_8bit_array_3.drv<31:0>.n178 hgu_cdac_8bit_array_3.drv<31:0>.n177 0.0143235
R4709 hgu_cdac_8bit_array_3.drv<31:0>.n180 hgu_cdac_8bit_array_3.drv<31:0>.n179 0.0143235
R4710 hgu_cdac_8bit_array_3.drv<31:0>.n187 hgu_cdac_8bit_array_3.drv<31:0>.n186 0.0143235
R4711 hgu_cdac_8bit_array_3.drv<31:0>.n189 hgu_cdac_8bit_array_3.drv<31:0>.n188 0.0143235
R4712 hgu_cdac_8bit_array_3.drv<31:0>.n196 hgu_cdac_8bit_array_3.drv<31:0>.n195 0.0143235
R4713 hgu_cdac_8bit_array_3.drv<31:0>.n198 hgu_cdac_8bit_array_3.drv<31:0>.n197 0.0143235
R4714 hgu_cdac_8bit_array_3.drv<31:0>.n205 hgu_cdac_8bit_array_3.drv<31:0>.n204 0.0143235
R4715 hgu_cdac_8bit_array_3.drv<31:0>.n207 hgu_cdac_8bit_array_3.drv<31:0>.n206 0.0143235
R4716 hgu_cdac_8bit_array_3.drv<31:0>.n214 hgu_cdac_8bit_array_3.drv<31:0>.n213 0.0143235
R4717 hgu_cdac_8bit_array_3.drv<31:0>.n216 hgu_cdac_8bit_array_3.drv<31:0>.n215 0.0143235
R4718 hgu_cdac_8bit_array_3.drv<31:0>.n223 hgu_cdac_8bit_array_3.drv<31:0>.n222 0.0143235
R4719 hgu_cdac_8bit_array_3.drv<31:0>.n225 hgu_cdac_8bit_array_3.drv<31:0>.n224 0.0143235
R4720 hgu_cdac_8bit_array_3.drv<31:0>.n232 hgu_cdac_8bit_array_3.drv<31:0>.n231 0.0143235
R4721 hgu_cdac_8bit_array_3.drv<31:0>.n234 hgu_cdac_8bit_array_3.drv<31:0>.n233 0.0143235
R4722 hgu_cdac_8bit_array_3.drv<31:0>.n288 hgu_cdac_8bit_array_3.drv<31:0>.n287 0.0143235
R4723 hgu_cdac_8bit_array_3.drv<31:0>.n286 hgu_cdac_8bit_array_3.drv<31:0>.n285 0.0143235
R4724 hgu_cdac_8bit_array_3.drv<31:0>.n279 hgu_cdac_8bit_array_3.drv<31:0>.n278 0.0143235
R4725 hgu_cdac_8bit_array_3.drv<31:0>.n277 hgu_cdac_8bit_array_3.drv<31:0>.n276 0.0143235
R4726 hgu_cdac_8bit_array_3.drv<31:0>.n270 hgu_cdac_8bit_array_3.drv<31:0>.n269 0.0143235
R4727 hgu_cdac_8bit_array_3.drv<31:0>.n268 hgu_cdac_8bit_array_3.drv<31:0>.n267 0.0143235
R4728 VSS.n1051 VSS.n1050 4683.73
R4729 VSS.n846 VSS.n845 4009.33
R4730 VSS.n601 VSS.n600 3413.49
R4731 VSS.n905 VSS.n904 3100.34
R4732 VSS.n811 VSS.n810 2862.07
R4733 VSS.n870 VSS.n869 2703.23
R4734 VSS.n743 VSS.n742 2639.69
R4735 VSS.n597 VSS.n3 2629.01
R4736 VSS.n971 VSS.n970 2544.38
R4737 VSS.n497 VSS.n496 2085.79
R4738 VSS.n1054 VSS.n1053 1597.5
R4739 VSS.n499 VSS.n495 1590.54
R4740 VSS.n881 VSS.n880 1527.78
R4741 VSS.n443 VSS.n442 1292.49
R4742 VSS.n445 VSS.n441 985.322
R4743 VSS.n861 VSS.t444 977.779
R4744 VSS.n898 VSS.t422 977.779
R4745 VSS.n863 VSS.t476 977.779
R4746 VSS.n865 VSS.t186 977.779
R4747 VSS.n811 VSS.t440 977.779
R4748 VSS.n964 VSS.t496 977.779
R4749 VSS.n813 VSS.t170 977.779
R4750 VSS.n815 VSS.t494 977.779
R4751 VSS.n820 VSS.t378 977.779
R4752 VSS.n956 VSS.t368 977.779
R4753 VSS.n822 VSS.t386 977.779
R4754 VSS.n950 VSS.t446 977.779
R4755 VSS.n826 VSS.t500 977.779
R4756 VSS.n828 VSS.t438 977.779
R4757 VSS.n833 VSS.t178 977.779
R4758 VSS.n942 VSS.t400 977.779
R4759 VSS.n835 VSS.t364 977.779
R4760 VSS.n936 VSS.t466 977.779
R4761 VSS.n839 VSS.t468 977.779
R4762 VSS.n841 VSS.t392 977.779
R4763 VSS.n1051 VSS.t130 977.779
R4764 VSS.n745 VSS.t154 977.779
R4765 VSS.n1044 VSS.t98 977.779
R4766 VSS.n747 VSS.t102 977.779
R4767 VSS.n1038 VSS.t128 977.779
R4768 VSS.n752 VSS.t108 977.779
R4769 VSS.n754 VSS.t132 977.779
R4770 VSS.n758 VSS.t120 977.779
R4771 VSS.n1030 VSS.t150 977.779
R4772 VSS.n760 VSS.t106 977.779
R4773 VSS.n1024 VSS.t114 977.779
R4774 VSS.n765 VSS.t140 977.779
R4775 VSS.n767 VSS.t146 977.779
R4776 VSS.n771 VSS.t126 977.779
R4777 VSS.n1016 VSS.t136 977.779
R4778 VSS.n773 VSS.t160 977.779
R4779 VSS.n1010 VSS.t118 977.779
R4780 VSS.n778 VSS.t124 977.779
R4781 VSS.n780 VSS.t134 977.779
R4782 VSS.n784 VSS.t158 977.779
R4783 VSS.n1002 VSS.t116 977.779
R4784 VSS.n786 VSS.t148 977.779
R4785 VSS.n996 VSS.t156 977.779
R4786 VSS.n791 VSS.t112 977.779
R4787 VSS.n793 VSS.t138 977.779
R4788 VSS.n797 VSS.t144 977.779
R4789 VSS.n988 VSS.t104 977.779
R4790 VSS.n799 VSS.t110 977.779
R4791 VSS.n982 VSS.t142 977.779
R4792 VSS.n804 VSS.t100 977.779
R4793 VSS.n806 VSS.t122 977.779
R4794 VSS.n975 VSS.t152 977.779
R4795 VSS.n605 VSS.t284 977.779
R4796 VSS.n610 VSS.t268 977.779
R4797 VSS.n610 VSS.t322 977.779
R4798 VSS.n1197 VSS.t244 977.779
R4799 VSS.n612 VSS.t296 977.779
R4800 VSS.n1191 VSS.t220 977.779
R4801 VSS.n616 VSS.t234 977.779
R4802 VSS.n618 VSS.t276 977.779
R4803 VSS.n623 VSS.t292 977.779
R4804 VSS.n1183 VSS.t344 977.779
R4805 VSS.n625 VSS.t262 977.779
R4806 VSS.n1177 VSS.t272 977.779
R4807 VSS.n629 VSS.t338 977.779
R4808 VSS.n631 VSS.t256 977.779
R4809 VSS.n636 VSS.t300 977.779
R4810 VSS.n1169 VSS.t318 977.779
R4811 VSS.n638 VSS.t334 977.779
R4812 VSS.n1163 VSS.t252 977.779
R4813 VSS.n642 VSS.t298 977.779
R4814 VSS.n644 VSS.t314 977.779
R4815 VSS.n649 VSS.t274 977.779
R4816 VSS.n1155 VSS.t286 977.779
R4817 VSS.n651 VSS.t306 977.779
R4818 VSS.n1149 VSS.t230 977.779
R4819 VSS.n655 VSS.t270 977.779
R4820 VSS.n657 VSS.t324 977.779
R4821 VSS.n662 VSS.t302 977.779
R4822 VSS.n1141 VSS.t226 977.779
R4823 VSS.n664 VSS.t312 977.779
R4824 VSS.n1135 VSS.t330 977.779
R4825 VSS.n668 VSS.t248 977.779
R4826 VSS.n670 VSS.t264 977.779
R4827 VSS.n675 VSS.t310 977.779
R4828 VSS.n1127 VSS.t328 977.779
R4829 VSS.n677 VSS.t246 977.779
R4830 VSS.n1121 VSS.t288 977.779
R4831 VSS.n681 VSS.t224 977.779
R4832 VSS.n683 VSS.t240 977.779
R4833 VSS.n688 VSS.t282 977.779
R4834 VSS.n1113 VSS.t336 977.779
R4835 VSS.n690 VSS.t222 977.779
R4836 VSS.n1107 VSS.t238 977.779
R4837 VSS.n694 VSS.t280 977.779
R4838 VSS.n696 VSS.t332 977.779
R4839 VSS.n701 VSS.t260 977.779
R4840 VSS.n1099 VSS.t308 977.779
R4841 VSS.n703 VSS.t326 977.779
R4842 VSS.n1093 VSS.t340 977.779
R4843 VSS.n707 VSS.t258 977.779
R4844 VSS.n709 VSS.t304 977.779
R4845 VSS.n714 VSS.t228 977.779
R4846 VSS.n1085 VSS.t250 977.779
R4847 VSS.n716 VSS.t294 977.779
R4848 VSS.n1079 VSS.t218 977.779
R4849 VSS.n720 VSS.t236 977.779
R4850 VSS.n722 VSS.t278 977.779
R4851 VSS.n727 VSS.t290 977.779
R4852 VSS.n1071 VSS.t342 977.779
R4853 VSS.n729 VSS.t232 977.779
R4854 VSS.n1065 VSS.t320 977.779
R4855 VSS.n733 VSS.t242 977.779
R4856 VSS.n735 VSS.t254 977.779
R4857 VSS.n740 VSS.t266 977.779
R4858 VSS.n1057 VSS.t316 977.779
R4859 VSS.n928 VSS.t452 977.779
R4860 VSS.n848 VSS.t456 977.779
R4861 VSS.n922 VSS.t460 977.779
R4862 VSS.n850 VSS.t462 977.779
R4863 VSS.n916 VSS.t450 977.779
R4864 VSS.n855 VSS.t454 977.779
R4865 VSS.n857 VSS.t458 977.779
R4866 VSS.n909 VSS.t448 977.779
R4867 VSS.n872 VSS.t394 977.779
R4868 VSS.n890 VSS.t388 977.779
R4869 VSS.n885 VSS.t390 977.779
R4870 VSS.n973 VSS.n969 845.635
R4871 VSS.n931 VSS.n930 408.765
R4872 VSS.n412 VSS.n411 404.312
R4873 VSS.n396 VSS.n395 367.822
R4874 VSS.n414 VSS.n410 308.036
R4875 VSS.n907 VSS.n903 308.036
R4876 VSS.n383 VSS.n382 291.923
R4877 VSS.n398 VSS.n394 280.488
R4878 VSS.n600 VSS.n599 274.284
R4879 VSS.n385 VSS.n381 222.609
R4880 VSS.n883 VSS.n879 186.992
R4881 VSS.n893 VSS.n892 173.636
R4882 VSS.n1 VSS.n0 170.837
R4883 VSS.n94 VSS.t380 46.7081
R4884 VSS.n105 VSS.t348 46.7081
R4885 VSS.n108 VSS.t176 46.7081
R4886 VSS.n90 VSS.t354 46.7081
R4887 VSS.n114 VSS.t410 46.7081
R4888 VSS.n117 VSS.t442 46.7081
R4889 VSS.n85 VSS.t188 46.7081
R4890 VSS.n123 VSS.t82 46.7081
R4891 VSS.n126 VSS.t94 46.7081
R4892 VSS.n81 VSS.t408 46.7081
R4893 VSS.n132 VSS.t398 46.7081
R4894 VSS.n135 VSS.t194 46.7081
R4895 VSS.n76 VSS.t356 46.7081
R4896 VSS.n141 VSS.t162 46.7081
R4897 VSS.n144 VSS.t404 46.7081
R4898 VSS.n72 VSS.t216 46.7081
R4899 VSS.n150 VSS.t180 46.7081
R4900 VSS.n153 VSS.t366 46.7081
R4901 VSS.n67 VSS.t426 46.7081
R4902 VSS.n159 VSS.t68 46.7081
R4903 VSS.n162 VSS.t196 46.7081
R4904 VSS.n63 VSS.t184 46.7081
R4905 VSS.n168 VSS.t472 46.7081
R4906 VSS.n171 VSS.t168 46.7081
R4907 VSS.n58 VSS.t78 46.7081
R4908 VSS.n177 VSS.t172 46.7081
R4909 VSS.n180 VSS.t370 46.7081
R4910 VSS.n54 VSS.t200 46.7081
R4911 VSS.n186 VSS.t434 46.7081
R4912 VSS.n189 VSS.t474 46.7081
R4913 VSS.n49 VSS.t80 46.7081
R4914 VSS.n195 VSS.t374 46.7081
R4915 VSS.n198 VSS.t420 46.7081
R4916 VSS.n45 VSS.t174 46.7081
R4917 VSS.n204 VSS.t498 46.7081
R4918 VSS.n207 VSS.t214 46.7081
R4919 VSS.n40 VSS.t198 46.7081
R4920 VSS.n213 VSS.t436 46.7081
R4921 VSS.n216 VSS.t182 46.7081
R4922 VSS.n36 VSS.t70 46.7081
R4923 VSS.n222 VSS.t166 46.7081
R4924 VSS.n225 VSS.t406 46.7081
R4925 VSS.n31 VSS.t432 46.7081
R4926 VSS.n231 VSS.t430 46.7081
R4927 VSS.n234 VSS.t64 46.7081
R4928 VSS.n27 VSS.t384 46.7081
R4929 VSS.n240 VSS.t86 46.7081
R4930 VSS.n243 VSS.t88 46.7081
R4931 VSS.n22 VSS.t382 46.7081
R4932 VSS.n249 VSS.t212 46.7081
R4933 VSS.n252 VSS.t418 46.7081
R4934 VSS.n18 VSS.t360 46.7081
R4935 VSS.n258 VSS.t372 46.7081
R4936 VSS.n261 VSS.t362 46.7081
R4937 VSS.n13 VSS.t396 46.7081
R4938 VSS.n267 VSS.t504 46.7081
R4939 VSS.n270 VSS.t84 46.7081
R4940 VSS.n9 VSS.t424 46.7081
R4941 VSS.n276 VSS.t192 46.7081
R4942 VSS.n279 VSS.t350 46.7081
R4943 VSS.n4 VSS.t416 46.7081
R4944 VSS.n285 VSS.t210 46.7081
R4945 VSS.n288 VSS.t164 46.7081
R4946 VSS.n599 VSS.t376 46.7081
R4947 VSS.n1 VSS.t6 46.7081
R4948 VSS.n591 VSS.t28 46.7081
R4949 VSS.n588 VSS.t20 46.7081
R4950 VSS.n292 VSS.t48 46.7081
R4951 VSS.n582 VSS.t4 46.7081
R4952 VSS.n579 VSS.t14 46.7081
R4953 VSS.n297 VSS.t38 46.7081
R4954 VSS.n573 VSS.t0 46.7081
R4955 VSS.n570 VSS.t26 46.7081
R4956 VSS.n301 VSS.t32 46.7081
R4957 VSS.n564 VSS.t58 46.7081
R4958 VSS.n561 VSS.t16 46.7081
R4959 VSS.n306 VSS.t24 46.7081
R4960 VSS.n555 VSS.t30 46.7081
R4961 VSS.n552 VSS.t56 46.7081
R4962 VSS.n310 VSS.t36 46.7081
R4963 VSS.n546 VSS.t46 46.7081
R4964 VSS.n543 VSS.t54 46.7081
R4965 VSS.n315 VSS.t12 46.7081
R4966 VSS.n537 VSS.t34 46.7081
R4967 VSS.n536 VSS.t44 46.7081
R4968 VSS.n319 VSS.t2 46.7081
R4969 VSS.n528 VSS.t8 46.7081
R4970 VSS.n525 VSS.t42 46.7081
R4971 VSS.n324 VSS.t62 46.7081
R4972 VSS.n519 VSS.t22 46.7081
R4973 VSS.n516 VSS.t50 46.7081
R4974 VSS.n328 VSS.t40 46.7081
R4975 VSS.n510 VSS.t60 46.7081
R4976 VSS.n507 VSS.t18 46.7081
R4977 VSS.n333 VSS.t52 46.7081
R4978 VSS.n501 VSS.t10 46.7081
R4979 VSS.n493 VSS.t502 46.7081
R4980 VSS.n488 VSS.t190 46.7081
R4981 VSS.n485 VSS.t208 46.7081
R4982 VSS.n337 VSS.t358 46.7081
R4983 VSS.n479 VSS.t202 46.7081
R4984 VSS.n476 VSS.t352 46.7081
R4985 VSS.n342 VSS.t204 46.7081
R4986 VSS.n470 VSS.t92 46.7081
R4987 VSS.n467 VSS.t66 46.7081
R4988 VSS.n346 VSS.t414 46.7081
R4989 VSS.n461 VSS.t96 46.7081
R4990 VSS.n458 VSS.t506 46.7081
R4991 VSS.n351 VSS.t206 46.7081
R4992 VSS.n452 VSS.t76 46.7081
R4993 VSS.n449 VSS.t74 46.7081
R4994 VSS.n355 VSS.t428 46.7081
R4995 VSS.n439 VSS.t482 46.7081
R4996 VSS.n434 VSS.t488 46.7081
R4997 VSS.n431 VSS.t484 46.7081
R4998 VSS.n359 VSS.t492 46.7081
R4999 VSS.n425 VSS.t486 46.7081
R5000 VSS.n422 VSS.t490 46.7081
R5001 VSS.n364 VSS.t478 46.7081
R5002 VSS.n416 VSS.t480 46.7081
R5003 VSS.n408 VSS.t402 46.7081
R5004 VSS.n368 VSS.t72 46.7081
R5005 VSS.n402 VSS.t412 46.7081
R5006 VSS.n370 VSS.t470 46.7081
R5007 VSS.n392 VSS.t90 46.7081
R5008 VSS.n387 VSS.t464 46.7081
R5009 VSS.n379 VSS.t346 46.7081
R5010 VSS VSS.n536 43.7889
R5011 VSS.n877 VSS.t395 41.7588
R5012 VSS.n884 VSS.t391 41.7588
R5013 VSS.n889 VSS.t389 41.7588
R5014 VSS.n894 VSS.t187 41.7588
R5015 VSS.n902 VSS.t445 41.7588
R5016 VSS.n908 VSS.t449 41.7588
R5017 VSS.n927 VSS.t453 41.7588
R5018 VSS.n932 VSS.t393 41.7588
R5019 VSS.n968 VSS.t441 41.7588
R5020 VSS.n974 VSS.t153 41.7588
R5021 VSS.n1049 VSS.t131 41.7588
R5022 VSS.n1055 VSS.t317 41.7588
R5023 VSS.n604 VSS.t285 41.7588
R5024 VSS.n415 VSS.t481 41.7588
R5025 VSS.n438 VSS.t483 41.7588
R5026 VSS.n446 VSS.t429 41.7588
R5027 VSS.n492 VSS.t503 41.7588
R5028 VSS.n500 VSS.t11 41.7588
R5029 VSS.n595 VSS.t7 41.7588
R5030 VSS.n407 VSS.t403 41.7588
R5031 VSS.n399 VSS.t471 41.7588
R5032 VSS.n391 VSS.t91 41.7588
R5033 VSS.n386 VSS.t465 41.7588
R5034 VSS.n102 VSS.t381 41.7588
R5035 VSS.n596 VSS.t377 41.7588
R5036 VSS.n377 VSS.t347 41.7588
R5037 VSS.n868 VSS.t423 41.4291
R5038 VSS.n868 VSS.t477 41.4291
R5039 VSS.n860 VSS.t455 41.4291
R5040 VSS.n860 VSS.t459 41.4291
R5041 VSS.n854 VSS.t463 41.4291
R5042 VSS.n854 VSS.t451 41.4291
R5043 VSS.n853 VSS.t457 41.4291
R5044 VSS.n853 VSS.t461 41.4291
R5045 VSS.n844 VSS.t467 41.4291
R5046 VSS.n844 VSS.t469 41.4291
R5047 VSS.n838 VSS.t401 41.4291
R5048 VSS.n838 VSS.t365 41.4291
R5049 VSS.n832 VSS.t439 41.4291
R5050 VSS.n832 VSS.t179 41.4291
R5051 VSS.n831 VSS.t447 41.4291
R5052 VSS.n831 VSS.t501 41.4291
R5053 VSS.n825 VSS.t369 41.4291
R5054 VSS.n825 VSS.t387 41.4291
R5055 VSS.n819 VSS.t495 41.4291
R5056 VSS.n819 VSS.t379 41.4291
R5057 VSS.n818 VSS.t497 41.4291
R5058 VSS.n818 VSS.t171 41.4291
R5059 VSS.n809 VSS.t101 41.4291
R5060 VSS.n809 VSS.t123 41.4291
R5061 VSS.n803 VSS.t111 41.4291
R5062 VSS.n803 VSS.t143 41.4291
R5063 VSS.n802 VSS.t145 41.4291
R5064 VSS.n802 VSS.t105 41.4291
R5065 VSS.n796 VSS.t113 41.4291
R5066 VSS.n796 VSS.t139 41.4291
R5067 VSS.n790 VSS.t149 41.4291
R5068 VSS.n790 VSS.t157 41.4291
R5069 VSS.n789 VSS.t159 41.4291
R5070 VSS.n789 VSS.t117 41.4291
R5071 VSS.n783 VSS.t125 41.4291
R5072 VSS.n783 VSS.t135 41.4291
R5073 VSS.n777 VSS.t161 41.4291
R5074 VSS.n777 VSS.t119 41.4291
R5075 VSS.n776 VSS.t127 41.4291
R5076 VSS.n776 VSS.t137 41.4291
R5077 VSS.n770 VSS.t141 41.4291
R5078 VSS.n770 VSS.t147 41.4291
R5079 VSS.n764 VSS.t107 41.4291
R5080 VSS.n764 VSS.t115 41.4291
R5081 VSS.n763 VSS.t121 41.4291
R5082 VSS.n763 VSS.t151 41.4291
R5083 VSS.n757 VSS.t109 41.4291
R5084 VSS.n757 VSS.t133 41.4291
R5085 VSS.n751 VSS.t103 41.4291
R5086 VSS.n751 VSS.t129 41.4291
R5087 VSS.n750 VSS.t155 41.4291
R5088 VSS.n750 VSS.t99 41.4291
R5089 VSS.n739 VSS.t255 41.4291
R5090 VSS.n739 VSS.t267 41.4291
R5091 VSS.n738 VSS.t321 41.4291
R5092 VSS.n738 VSS.t243 41.4291
R5093 VSS.n732 VSS.t343 41.4291
R5094 VSS.n732 VSS.t233 41.4291
R5095 VSS.n726 VSS.t279 41.4291
R5096 VSS.n726 VSS.t291 41.4291
R5097 VSS.n725 VSS.t219 41.4291
R5098 VSS.n725 VSS.t237 41.4291
R5099 VSS.n719 VSS.t251 41.4291
R5100 VSS.n719 VSS.t295 41.4291
R5101 VSS.n713 VSS.t305 41.4291
R5102 VSS.n713 VSS.t229 41.4291
R5103 VSS.n712 VSS.t341 41.4291
R5104 VSS.n712 VSS.t259 41.4291
R5105 VSS.n706 VSS.t309 41.4291
R5106 VSS.n706 VSS.t327 41.4291
R5107 VSS.n700 VSS.t333 41.4291
R5108 VSS.n700 VSS.t261 41.4291
R5109 VSS.n699 VSS.t239 41.4291
R5110 VSS.n699 VSS.t281 41.4291
R5111 VSS.n693 VSS.t337 41.4291
R5112 VSS.n693 VSS.t223 41.4291
R5113 VSS.n687 VSS.t241 41.4291
R5114 VSS.n687 VSS.t283 41.4291
R5115 VSS.n686 VSS.t289 41.4291
R5116 VSS.n686 VSS.t225 41.4291
R5117 VSS.n680 VSS.t329 41.4291
R5118 VSS.n680 VSS.t247 41.4291
R5119 VSS.n674 VSS.t265 41.4291
R5120 VSS.n674 VSS.t311 41.4291
R5121 VSS.n673 VSS.t331 41.4291
R5122 VSS.n673 VSS.t249 41.4291
R5123 VSS.n667 VSS.t227 41.4291
R5124 VSS.n667 VSS.t313 41.4291
R5125 VSS.n661 VSS.t325 41.4291
R5126 VSS.n661 VSS.t303 41.4291
R5127 VSS.n660 VSS.t231 41.4291
R5128 VSS.n660 VSS.t271 41.4291
R5129 VSS.n654 VSS.t287 41.4291
R5130 VSS.n654 VSS.t307 41.4291
R5131 VSS.n648 VSS.t315 41.4291
R5132 VSS.n648 VSS.t275 41.4291
R5133 VSS.n647 VSS.t253 41.4291
R5134 VSS.n647 VSS.t299 41.4291
R5135 VSS.n641 VSS.t319 41.4291
R5136 VSS.n641 VSS.t335 41.4291
R5137 VSS.n635 VSS.t257 41.4291
R5138 VSS.n635 VSS.t301 41.4291
R5139 VSS.n634 VSS.t273 41.4291
R5140 VSS.n634 VSS.t339 41.4291
R5141 VSS.n628 VSS.t345 41.4291
R5142 VSS.n628 VSS.t263 41.4291
R5143 VSS.n622 VSS.t277 41.4291
R5144 VSS.n622 VSS.t293 41.4291
R5145 VSS.n621 VSS.t221 41.4291
R5146 VSS.n621 VSS.t235 41.4291
R5147 VSS.n615 VSS.t245 41.4291
R5148 VSS.n615 VSS.t297 41.4291
R5149 VSS.n609 VSS.t269 41.4291
R5150 VSS.n609 VSS.t323 41.4291
R5151 VSS.n367 VSS.t491 41.4291
R5152 VSS.n367 VSS.t479 41.4291
R5153 VSS.n363 VSS.t493 41.4291
R5154 VSS.n363 VSS.t487 41.4291
R5155 VSS.n362 VSS.t489 41.4291
R5156 VSS.n362 VSS.t485 41.4291
R5157 VSS.n358 VSS.t77 41.4291
R5158 VSS.n358 VSS.t75 41.4291
R5159 VSS.n354 VSS.t507 41.4291
R5160 VSS.n354 VSS.t207 41.4291
R5161 VSS.n350 VSS.t415 41.4291
R5162 VSS.n350 VSS.t97 41.4291
R5163 VSS.n349 VSS.t93 41.4291
R5164 VSS.n349 VSS.t67 41.4291
R5165 VSS.n345 VSS.t353 41.4291
R5166 VSS.n345 VSS.t205 41.4291
R5167 VSS.n341 VSS.t359 41.4291
R5168 VSS.n341 VSS.t203 41.4291
R5169 VSS.n340 VSS.t191 41.4291
R5170 VSS.n340 VSS.t209 41.4291
R5171 VSS.n336 VSS.t19 41.4291
R5172 VSS.n336 VSS.t53 41.4291
R5173 VSS.n332 VSS.t41 41.4291
R5174 VSS.n332 VSS.t61 41.4291
R5175 VSS.n331 VSS.t23 41.4291
R5176 VSS.n331 VSS.t51 41.4291
R5177 VSS.n327 VSS.t43 41.4291
R5178 VSS.n327 VSS.t63 41.4291
R5179 VSS.n323 VSS.t3 41.4291
R5180 VSS.n323 VSS.t9 41.4291
R5181 VSS.n322 VSS.t35 41.4291
R5182 VSS.n322 VSS.t45 41.4291
R5183 VSS.n318 VSS.t55 41.4291
R5184 VSS.n318 VSS.t13 41.4291
R5185 VSS.n314 VSS.t37 41.4291
R5186 VSS.n314 VSS.t47 41.4291
R5187 VSS.n313 VSS.t31 41.4291
R5188 VSS.n313 VSS.t57 41.4291
R5189 VSS.n309 VSS.t17 41.4291
R5190 VSS.n309 VSS.t25 41.4291
R5191 VSS.n305 VSS.t33 41.4291
R5192 VSS.n305 VSS.t59 41.4291
R5193 VSS.n304 VSS.t1 41.4291
R5194 VSS.n304 VSS.t27 41.4291
R5195 VSS.n300 VSS.t15 41.4291
R5196 VSS.n300 VSS.t39 41.4291
R5197 VSS.n296 VSS.t49 41.4291
R5198 VSS.n296 VSS.t5 41.4291
R5199 VSS.n295 VSS.t29 41.4291
R5200 VSS.n295 VSS.t21 41.4291
R5201 VSS.n373 VSS.t73 41.4291
R5202 VSS.n373 VSS.t413 41.4291
R5203 VSS.n7 VSS.t211 41.4291
R5204 VSS.n7 VSS.t165 41.4291
R5205 VSS.n8 VSS.t351 41.4291
R5206 VSS.n8 VSS.t417 41.4291
R5207 VSS.n12 VSS.t425 41.4291
R5208 VSS.n12 VSS.t193 41.4291
R5209 VSS.n16 VSS.t505 41.4291
R5210 VSS.n16 VSS.t85 41.4291
R5211 VSS.n17 VSS.t363 41.4291
R5212 VSS.n17 VSS.t397 41.4291
R5213 VSS.n21 VSS.t361 41.4291
R5214 VSS.n21 VSS.t373 41.4291
R5215 VSS.n25 VSS.t213 41.4291
R5216 VSS.n25 VSS.t419 41.4291
R5217 VSS.n26 VSS.t89 41.4291
R5218 VSS.n26 VSS.t383 41.4291
R5219 VSS.n30 VSS.t385 41.4291
R5220 VSS.n30 VSS.t87 41.4291
R5221 VSS.n34 VSS.t431 41.4291
R5222 VSS.n34 VSS.t65 41.4291
R5223 VSS.n35 VSS.t407 41.4291
R5224 VSS.n35 VSS.t433 41.4291
R5225 VSS.n39 VSS.t71 41.4291
R5226 VSS.n39 VSS.t167 41.4291
R5227 VSS.n43 VSS.t437 41.4291
R5228 VSS.n43 VSS.t183 41.4291
R5229 VSS.n44 VSS.t215 41.4291
R5230 VSS.n44 VSS.t199 41.4291
R5231 VSS.n48 VSS.t175 41.4291
R5232 VSS.n48 VSS.t499 41.4291
R5233 VSS.n52 VSS.t375 41.4291
R5234 VSS.n52 VSS.t421 41.4291
R5235 VSS.n53 VSS.t475 41.4291
R5236 VSS.n53 VSS.t81 41.4291
R5237 VSS.n57 VSS.t201 41.4291
R5238 VSS.n57 VSS.t435 41.4291
R5239 VSS.n61 VSS.t173 41.4291
R5240 VSS.n61 VSS.t371 41.4291
R5241 VSS.n62 VSS.t169 41.4291
R5242 VSS.n62 VSS.t79 41.4291
R5243 VSS.n66 VSS.t185 41.4291
R5244 VSS.n66 VSS.t473 41.4291
R5245 VSS.n70 VSS.t69 41.4291
R5246 VSS.n70 VSS.t197 41.4291
R5247 VSS.n71 VSS.t367 41.4291
R5248 VSS.n71 VSS.t427 41.4291
R5249 VSS.n75 VSS.t217 41.4291
R5250 VSS.n75 VSS.t181 41.4291
R5251 VSS.n79 VSS.t163 41.4291
R5252 VSS.n79 VSS.t405 41.4291
R5253 VSS.n80 VSS.t195 41.4291
R5254 VSS.n80 VSS.t357 41.4291
R5255 VSS.n84 VSS.t409 41.4291
R5256 VSS.n84 VSS.t399 41.4291
R5257 VSS.n88 VSS.t83 41.4291
R5258 VSS.n88 VSS.t95 41.4291
R5259 VSS.n89 VSS.t443 41.4291
R5260 VSS.n89 VSS.t189 41.4291
R5261 VSS.n93 VSS.t355 41.4291
R5262 VSS.n93 VSS.t411 41.4291
R5263 VSS.n97 VSS.t349 41.4291
R5264 VSS.n97 VSS.t177 41.4291
R5265 VSS.n107 VSS.n96 35.6179
R5266 VSS.n110 VSS.n107 35.6179
R5267 VSS.n110 VSS.n92 35.6179
R5268 VSS.n116 VSS.n92 35.6179
R5269 VSS.n119 VSS.n116 35.6179
R5270 VSS.n119 VSS.n87 35.6179
R5271 VSS.n125 VSS.n87 35.6179
R5272 VSS.n128 VSS.n125 35.6179
R5273 VSS.n128 VSS.n83 35.6179
R5274 VSS.n134 VSS.n83 35.6179
R5275 VSS.n137 VSS.n134 35.6179
R5276 VSS.n137 VSS.n78 35.6179
R5277 VSS.n143 VSS.n78 35.6179
R5278 VSS.n146 VSS.n143 35.6179
R5279 VSS.n146 VSS.n74 35.6179
R5280 VSS.n152 VSS.n74 35.6179
R5281 VSS.n155 VSS.n152 35.6179
R5282 VSS.n155 VSS.n69 35.6179
R5283 VSS.n161 VSS.n69 35.6179
R5284 VSS.n164 VSS.n161 35.6179
R5285 VSS.n164 VSS.n65 35.6179
R5286 VSS.n170 VSS.n65 35.6179
R5287 VSS.n173 VSS.n170 35.6179
R5288 VSS.n173 VSS.n60 35.6179
R5289 VSS.n179 VSS.n60 35.6179
R5290 VSS.n182 VSS.n179 35.6179
R5291 VSS.n182 VSS.n56 35.6179
R5292 VSS.n188 VSS.n56 35.6179
R5293 VSS.n191 VSS.n188 35.6179
R5294 VSS.n191 VSS.n51 35.6179
R5295 VSS.n197 VSS.n51 35.6179
R5296 VSS.n200 VSS.n197 35.6179
R5297 VSS.n200 VSS.n47 35.6179
R5298 VSS.n206 VSS.n47 35.6179
R5299 VSS.n209 VSS.n206 35.6179
R5300 VSS.n209 VSS.n42 35.6179
R5301 VSS.n215 VSS.n42 35.6179
R5302 VSS.n218 VSS.n215 35.6179
R5303 VSS.n218 VSS.n38 35.6179
R5304 VSS.n224 VSS.n38 35.6179
R5305 VSS.n227 VSS.n224 35.6179
R5306 VSS.n227 VSS.n33 35.6179
R5307 VSS.n233 VSS.n33 35.6179
R5308 VSS.n236 VSS.n233 35.6179
R5309 VSS.n236 VSS.n29 35.6179
R5310 VSS.n242 VSS.n29 35.6179
R5311 VSS.n245 VSS.n242 35.6179
R5312 VSS.n245 VSS.n24 35.6179
R5313 VSS.n251 VSS.n24 35.6179
R5314 VSS.n254 VSS.n251 35.6179
R5315 VSS.n254 VSS.n20 35.6179
R5316 VSS.n260 VSS.n20 35.6179
R5317 VSS.n263 VSS.n260 35.6179
R5318 VSS.n263 VSS.n15 35.6179
R5319 VSS.n269 VSS.n15 35.6179
R5320 VSS.n272 VSS.n269 35.6179
R5321 VSS.n272 VSS.n11 35.6179
R5322 VSS.n278 VSS.n11 35.6179
R5323 VSS.n281 VSS.n278 35.6179
R5324 VSS.n281 VSS.n6 35.6179
R5325 VSS.n287 VSS.n6 35.6179
R5326 VSS.n290 VSS.n287 35.6179
R5327 VSS.n593 VSS.n590 35.6179
R5328 VSS.n590 VSS.n294 35.6179
R5329 VSS.n584 VSS.n294 35.6179
R5330 VSS.n584 VSS.n581 35.6179
R5331 VSS.n581 VSS.n299 35.6179
R5332 VSS.n575 VSS.n299 35.6179
R5333 VSS.n575 VSS.n572 35.6179
R5334 VSS.n572 VSS.n303 35.6179
R5335 VSS.n566 VSS.n303 35.6179
R5336 VSS.n566 VSS.n563 35.6179
R5337 VSS.n563 VSS.n308 35.6179
R5338 VSS.n557 VSS.n308 35.6179
R5339 VSS.n557 VSS.n554 35.6179
R5340 VSS.n554 VSS.n312 35.6179
R5341 VSS.n548 VSS.n312 35.6179
R5342 VSS.n548 VSS.n545 35.6179
R5343 VSS.n545 VSS.n317 35.6179
R5344 VSS.n539 VSS.n317 35.6179
R5345 VSS.n539 VSS.n534 35.6179
R5346 VSS.n534 VSS.n321 35.6179
R5347 VSS.n530 VSS.n321 35.6179
R5348 VSS.n530 VSS.n527 35.6179
R5349 VSS.n527 VSS.n326 35.6179
R5350 VSS.n521 VSS.n326 35.6179
R5351 VSS.n521 VSS.n518 35.6179
R5352 VSS.n518 VSS.n330 35.6179
R5353 VSS.n512 VSS.n330 35.6179
R5354 VSS.n512 VSS.n509 35.6179
R5355 VSS.n509 VSS.n335 35.6179
R5356 VSS.n503 VSS.n335 35.6179
R5357 VSS.n490 VSS.n487 35.6179
R5358 VSS.n487 VSS.n339 35.6179
R5359 VSS.n481 VSS.n339 35.6179
R5360 VSS.n481 VSS.n478 35.6179
R5361 VSS.n478 VSS.n344 35.6179
R5362 VSS.n472 VSS.n344 35.6179
R5363 VSS.n472 VSS.n469 35.6179
R5364 VSS.n469 VSS.n348 35.6179
R5365 VSS.n463 VSS.n348 35.6179
R5366 VSS.n463 VSS.n460 35.6179
R5367 VSS.n460 VSS.n353 35.6179
R5368 VSS.n454 VSS.n353 35.6179
R5369 VSS.n454 VSS.n451 35.6179
R5370 VSS.n451 VSS.n357 35.6179
R5371 VSS.n436 VSS.n433 35.6179
R5372 VSS.n433 VSS.n361 35.6179
R5373 VSS.n427 VSS.n361 35.6179
R5374 VSS.n427 VSS.n424 35.6179
R5375 VSS.n424 VSS.n366 35.6179
R5376 VSS.n418 VSS.n366 35.6179
R5377 VSS.n405 VSS.n404 35.6179
R5378 VSS.n404 VSS.n372 35.6179
R5379 VSS.n1200 VSS.n1199 35.6179
R5380 VSS.n1199 VSS.n614 35.6179
R5381 VSS.n1193 VSS.n614 35.6179
R5382 VSS.n1193 VSS.n1190 35.6179
R5383 VSS.n1190 VSS.n620 35.6179
R5384 VSS.n1186 VSS.n620 35.6179
R5385 VSS.n1186 VSS.n1185 35.6179
R5386 VSS.n1185 VSS.n627 35.6179
R5387 VSS.n1179 VSS.n627 35.6179
R5388 VSS.n1179 VSS.n1176 35.6179
R5389 VSS.n1176 VSS.n633 35.6179
R5390 VSS.n1172 VSS.n633 35.6179
R5391 VSS.n1172 VSS.n1171 35.6179
R5392 VSS.n1171 VSS.n640 35.6179
R5393 VSS.n1165 VSS.n640 35.6179
R5394 VSS.n1165 VSS.n1162 35.6179
R5395 VSS.n1162 VSS.n646 35.6179
R5396 VSS.n1158 VSS.n646 35.6179
R5397 VSS.n1158 VSS.n1157 35.6179
R5398 VSS.n1157 VSS.n653 35.6179
R5399 VSS.n1151 VSS.n653 35.6179
R5400 VSS.n1151 VSS.n1148 35.6179
R5401 VSS.n1148 VSS.n659 35.6179
R5402 VSS.n1144 VSS.n659 35.6179
R5403 VSS.n1144 VSS.n1143 35.6179
R5404 VSS.n1143 VSS.n666 35.6179
R5405 VSS.n1137 VSS.n666 35.6179
R5406 VSS.n1137 VSS.n1134 35.6179
R5407 VSS.n1134 VSS.n672 35.6179
R5408 VSS.n1130 VSS.n672 35.6179
R5409 VSS.n1130 VSS.n1129 35.6179
R5410 VSS.n1129 VSS.n679 35.6179
R5411 VSS.n1123 VSS.n679 35.6179
R5412 VSS.n1123 VSS.n1120 35.6179
R5413 VSS.n1120 VSS.n685 35.6179
R5414 VSS.n1116 VSS.n685 35.6179
R5415 VSS.n1116 VSS.n1115 35.6179
R5416 VSS.n1115 VSS.n692 35.6179
R5417 VSS.n1109 VSS.n692 35.6179
R5418 VSS.n1109 VSS.n1106 35.6179
R5419 VSS.n1106 VSS.n698 35.6179
R5420 VSS.n1102 VSS.n698 35.6179
R5421 VSS.n1102 VSS.n1101 35.6179
R5422 VSS.n1101 VSS.n705 35.6179
R5423 VSS.n1095 VSS.n705 35.6179
R5424 VSS.n1095 VSS.n1092 35.6179
R5425 VSS.n1092 VSS.n711 35.6179
R5426 VSS.n1088 VSS.n711 35.6179
R5427 VSS.n1088 VSS.n1087 35.6179
R5428 VSS.n1087 VSS.n718 35.6179
R5429 VSS.n1081 VSS.n718 35.6179
R5430 VSS.n1081 VSS.n1078 35.6179
R5431 VSS.n1078 VSS.n724 35.6179
R5432 VSS.n1074 VSS.n724 35.6179
R5433 VSS.n1074 VSS.n1073 35.6179
R5434 VSS.n1073 VSS.n731 35.6179
R5435 VSS.n1067 VSS.n731 35.6179
R5436 VSS.n1067 VSS.n1064 35.6179
R5437 VSS.n1064 VSS.n737 35.6179
R5438 VSS.n1060 VSS.n737 35.6179
R5439 VSS.n1060 VSS.n1059 35.6179
R5440 VSS.n1047 VSS.n1046 35.6179
R5441 VSS.n1046 VSS.n749 35.6179
R5442 VSS.n1040 VSS.n749 35.6179
R5443 VSS.n1040 VSS.n1037 35.6179
R5444 VSS.n1037 VSS.n756 35.6179
R5445 VSS.n1033 VSS.n756 35.6179
R5446 VSS.n1033 VSS.n1032 35.6179
R5447 VSS.n1032 VSS.n762 35.6179
R5448 VSS.n1026 VSS.n762 35.6179
R5449 VSS.n1026 VSS.n1023 35.6179
R5450 VSS.n1023 VSS.n769 35.6179
R5451 VSS.n1019 VSS.n769 35.6179
R5452 VSS.n1019 VSS.n1018 35.6179
R5453 VSS.n1018 VSS.n775 35.6179
R5454 VSS.n1012 VSS.n775 35.6179
R5455 VSS.n1012 VSS.n1009 35.6179
R5456 VSS.n1009 VSS.n782 35.6179
R5457 VSS.n1005 VSS.n782 35.6179
R5458 VSS.n1005 VSS.n1004 35.6179
R5459 VSS.n1004 VSS.n788 35.6179
R5460 VSS.n998 VSS.n788 35.6179
R5461 VSS.n998 VSS.n995 35.6179
R5462 VSS.n995 VSS.n795 35.6179
R5463 VSS.n991 VSS.n795 35.6179
R5464 VSS.n991 VSS.n990 35.6179
R5465 VSS.n990 VSS.n801 35.6179
R5466 VSS.n984 VSS.n801 35.6179
R5467 VSS.n984 VSS.n981 35.6179
R5468 VSS.n981 VSS.n808 35.6179
R5469 VSS.n977 VSS.n808 35.6179
R5470 VSS.n966 VSS.n963 35.6179
R5471 VSS.n963 VSS.n817 35.6179
R5472 VSS.n959 VSS.n817 35.6179
R5473 VSS.n959 VSS.n958 35.6179
R5474 VSS.n958 VSS.n824 35.6179
R5475 VSS.n952 VSS.n824 35.6179
R5476 VSS.n952 VSS.n949 35.6179
R5477 VSS.n949 VSS.n830 35.6179
R5478 VSS.n945 VSS.n830 35.6179
R5479 VSS.n945 VSS.n944 35.6179
R5480 VSS.n944 VSS.n837 35.6179
R5481 VSS.n938 VSS.n837 35.6179
R5482 VSS.n938 VSS.n935 35.6179
R5483 VSS.n935 VSS.n843 35.6179
R5484 VSS.n925 VSS.n924 35.6179
R5485 VSS.n924 VSS.n852 35.6179
R5486 VSS.n918 VSS.n852 35.6179
R5487 VSS.n918 VSS.n915 35.6179
R5488 VSS.n915 VSS.n859 35.6179
R5489 VSS.n911 VSS.n859 35.6179
R5490 VSS.n900 VSS.n897 35.6179
R5491 VSS.n897 VSS.n867 35.6179
R5492 VSS.n98 VSS 27.2232
R5493 VSS VSS.n98 6.40136
R5494 VSS.t34 VSS 2.91972
R5495 VSS.n98 VSS 2.50734
R5496 VSS.n378 VSS 1.858
R5497 VSS.n878 VSS 1.538
R5498 VSS.n896 VSS.n868 0.330267
R5499 VSS.n913 VSS.n860 0.330267
R5500 VSS.n919 VSS.n854 0.330267
R5501 VSS.n921 VSS.n853 0.330267
R5502 VSS.n934 VSS.n844 0.330267
R5503 VSS.n940 VSS.n838 0.330267
R5504 VSS.n946 VSS.n832 0.330267
R5505 VSS.n948 VSS.n831 0.330267
R5506 VSS.n954 VSS.n825 0.330267
R5507 VSS.n960 VSS.n819 0.330267
R5508 VSS.n962 VSS.n818 0.330267
R5509 VSS.n979 VSS.n809 0.330267
R5510 VSS.n985 VSS.n803 0.330267
R5511 VSS.n987 VSS.n802 0.330267
R5512 VSS.n993 VSS.n796 0.330267
R5513 VSS.n999 VSS.n790 0.330267
R5514 VSS.n1001 VSS.n789 0.330267
R5515 VSS.n1007 VSS.n783 0.330267
R5516 VSS.n1013 VSS.n777 0.330267
R5517 VSS.n1015 VSS.n776 0.330267
R5518 VSS.n1021 VSS.n770 0.330267
R5519 VSS.n1027 VSS.n764 0.330267
R5520 VSS.n1029 VSS.n763 0.330267
R5521 VSS.n1035 VSS.n757 0.330267
R5522 VSS.n1041 VSS.n751 0.330267
R5523 VSS.n1043 VSS.n750 0.330267
R5524 VSS.n1061 VSS.n739 0.330267
R5525 VSS.n1063 VSS.n738 0.330267
R5526 VSS.n1069 VSS.n732 0.330267
R5527 VSS.n1075 VSS.n726 0.330267
R5528 VSS.n1077 VSS.n725 0.330267
R5529 VSS.n1083 VSS.n719 0.330267
R5530 VSS.n1089 VSS.n713 0.330267
R5531 VSS.n1091 VSS.n712 0.330267
R5532 VSS.n1097 VSS.n706 0.330267
R5533 VSS.n1103 VSS.n700 0.330267
R5534 VSS.n1105 VSS.n699 0.330267
R5535 VSS.n1111 VSS.n693 0.330267
R5536 VSS.n1117 VSS.n687 0.330267
R5537 VSS.n1119 VSS.n686 0.330267
R5538 VSS.n1125 VSS.n680 0.330267
R5539 VSS.n1131 VSS.n674 0.330267
R5540 VSS.n1133 VSS.n673 0.330267
R5541 VSS.n1139 VSS.n667 0.330267
R5542 VSS.n1145 VSS.n661 0.330267
R5543 VSS.n1147 VSS.n660 0.330267
R5544 VSS.n1153 VSS.n654 0.330267
R5545 VSS.n1159 VSS.n648 0.330267
R5546 VSS.n1161 VSS.n647 0.330267
R5547 VSS.n1167 VSS.n641 0.330267
R5548 VSS.n1173 VSS.n635 0.330267
R5549 VSS.n1175 VSS.n634 0.330267
R5550 VSS.n1181 VSS.n628 0.330267
R5551 VSS.n1187 VSS.n622 0.330267
R5552 VSS.n1189 VSS.n621 0.330267
R5553 VSS.n1195 VSS.n615 0.330267
R5554 VSS.n1201 VSS.n609 0.330267
R5555 VSS.n420 VSS.n367 0.330267
R5556 VSS.n428 VSS.n363 0.330267
R5557 VSS.n430 VSS.n362 0.330267
R5558 VSS.n448 VSS.n358 0.330267
R5559 VSS.n456 VSS.n354 0.330267
R5560 VSS.n464 VSS.n350 0.330267
R5561 VSS.n466 VSS.n349 0.330267
R5562 VSS.n474 VSS.n345 0.330267
R5563 VSS.n482 VSS.n341 0.330267
R5564 VSS.n484 VSS.n340 0.330267
R5565 VSS.n505 VSS.n336 0.330267
R5566 VSS.n513 VSS.n332 0.330267
R5567 VSS.n515 VSS.n331 0.330267
R5568 VSS.n523 VSS.n327 0.330267
R5569 VSS.n531 VSS.n323 0.330267
R5570 VSS.n533 VSS.n322 0.330267
R5571 VSS.n541 VSS.n318 0.330267
R5572 VSS.n549 VSS.n314 0.330267
R5573 VSS.n551 VSS.n313 0.330267
R5574 VSS.n559 VSS.n309 0.330267
R5575 VSS.n567 VSS.n305 0.330267
R5576 VSS.n569 VSS.n304 0.330267
R5577 VSS.n577 VSS.n300 0.330267
R5578 VSS.n585 VSS.n296 0.330267
R5579 VSS.n587 VSS.n295 0.330267
R5580 VSS.n401 VSS.n373 0.330267
R5581 VSS.n284 VSS.n7 0.330267
R5582 VSS.n282 VSS.n8 0.330267
R5583 VSS.n274 VSS.n12 0.330267
R5584 VSS.n266 VSS.n16 0.330267
R5585 VSS.n264 VSS.n17 0.330267
R5586 VSS.n256 VSS.n21 0.330267
R5587 VSS.n248 VSS.n25 0.330267
R5588 VSS.n246 VSS.n26 0.330267
R5589 VSS.n238 VSS.n30 0.330267
R5590 VSS.n230 VSS.n34 0.330267
R5591 VSS.n228 VSS.n35 0.330267
R5592 VSS.n220 VSS.n39 0.330267
R5593 VSS.n212 VSS.n43 0.330267
R5594 VSS.n210 VSS.n44 0.330267
R5595 VSS.n202 VSS.n48 0.330267
R5596 VSS.n194 VSS.n52 0.330267
R5597 VSS.n192 VSS.n53 0.330267
R5598 VSS.n184 VSS.n57 0.330267
R5599 VSS.n176 VSS.n61 0.330267
R5600 VSS.n174 VSS.n62 0.330267
R5601 VSS.n166 VSS.n66 0.330267
R5602 VSS.n158 VSS.n70 0.330267
R5603 VSS.n156 VSS.n71 0.330267
R5604 VSS.n148 VSS.n75 0.330267
R5605 VSS.n140 VSS.n79 0.330267
R5606 VSS.n138 VSS.n80 0.330267
R5607 VSS.n130 VSS.n84 0.330267
R5608 VSS.n122 VSS.n88 0.330267
R5609 VSS.n120 VSS.n89 0.330267
R5610 VSS.n112 VSS.n93 0.330267
R5611 VSS.n104 VSS.n97 0.330267
R5612 VSS.n103 VSS.n102 0.3205
R5613 VSS.n596 VSS.n291 0.3205
R5614 VSS.n595 VSS.n594 0.3205
R5615 VSS.n504 VSS.n500 0.3205
R5616 VSS.n492 VSS.n491 0.3205
R5617 VSS.n447 VSS.n446 0.3205
R5618 VSS.n438 VSS.n437 0.3205
R5619 VSS.n419 VSS.n415 0.3205
R5620 VSS.n407 VSS.n406 0.3205
R5621 VSS.n400 VSS.n399 0.3205
R5622 VSS.n391 VSS.n390 0.3205
R5623 VSS.n390 VSS.n386 0.3205
R5624 VSS.n378 VSS.n377 0.3205
R5625 VSS.n608 VSS.n604 0.3205
R5626 VSS.n1056 VSS.n1055 0.3205
R5627 VSS.n1049 VSS.n1048 0.3205
R5628 VSS.n978 VSS.n974 0.3205
R5629 VSS.n968 VSS.n967 0.3205
R5630 VSS.n933 VSS.n932 0.3205
R5631 VSS.n927 VSS.n926 0.3205
R5632 VSS.n912 VSS.n908 0.3205
R5633 VSS.n902 VSS.n901 0.3205
R5634 VSS.n895 VSS.n894 0.3205
R5635 VSS.n889 VSS.n888 0.3205
R5636 VSS.n888 VSS.n884 0.3205
R5637 VSS.n878 VSS.n877 0.3205
R5638 VSS VSS.n103 0.238
R5639 VSS VSS.n111 0.238
R5640 VSS.n113 VSS 0.238
R5641 VSS VSS.n121 0.238
R5642 VSS VSS.n129 0.238
R5643 VSS.n131 VSS 0.238
R5644 VSS VSS.n139 0.238
R5645 VSS VSS.n147 0.238
R5646 VSS.n149 VSS 0.238
R5647 VSS VSS.n157 0.238
R5648 VSS VSS.n165 0.238
R5649 VSS.n167 VSS 0.238
R5650 VSS VSS.n175 0.238
R5651 VSS VSS.n183 0.238
R5652 VSS.n185 VSS 0.238
R5653 VSS VSS.n193 0.238
R5654 VSS VSS.n201 0.238
R5655 VSS.n203 VSS 0.238
R5656 VSS VSS.n211 0.238
R5657 VSS VSS.n219 0.238
R5658 VSS.n221 VSS 0.238
R5659 VSS VSS.n229 0.238
R5660 VSS VSS.n237 0.238
R5661 VSS.n239 VSS 0.238
R5662 VSS VSS.n247 0.238
R5663 VSS VSS.n255 0.238
R5664 VSS.n257 VSS 0.238
R5665 VSS VSS.n265 0.238
R5666 VSS VSS.n273 0.238
R5667 VSS.n275 VSS 0.238
R5668 VSS VSS.n283 0.238
R5669 VSS.n594 VSS 0.238
R5670 VSS.n586 VSS 0.238
R5671 VSS.n578 VSS 0.238
R5672 VSS.n576 VSS 0.238
R5673 VSS.n568 VSS 0.238
R5674 VSS.n560 VSS 0.238
R5675 VSS.n558 VSS 0.238
R5676 VSS.n550 VSS 0.238
R5677 VSS.n542 VSS 0.238
R5678 VSS.n540 VSS 0.238
R5679 VSS.n532 VSS 0.238
R5680 VSS.n524 VSS 0.238
R5681 VSS.n522 VSS 0.238
R5682 VSS.n514 VSS 0.238
R5683 VSS.n506 VSS 0.238
R5684 VSS.n491 VSS 0.238
R5685 VSS.n483 VSS 0.238
R5686 VSS.n475 VSS 0.238
R5687 VSS.n473 VSS 0.238
R5688 VSS.n465 VSS 0.238
R5689 VSS.n457 VSS 0.238
R5690 VSS.n455 VSS 0.238
R5691 VSS.n437 VSS 0.238
R5692 VSS.n429 VSS 0.238
R5693 VSS.n421 VSS 0.238
R5694 VSS.n406 VSS 0.238
R5695 VSS VSS.n608 0.238
R5696 VSS.n1196 VSS 0.238
R5697 VSS.n1194 VSS 0.238
R5698 VSS.n1188 VSS 0.238
R5699 VSS.n1182 VSS 0.238
R5700 VSS.n1180 VSS 0.238
R5701 VSS.n1174 VSS 0.238
R5702 VSS.n1168 VSS 0.238
R5703 VSS.n1166 VSS 0.238
R5704 VSS.n1160 VSS 0.238
R5705 VSS.n1154 VSS 0.238
R5706 VSS.n1152 VSS 0.238
R5707 VSS.n1146 VSS 0.238
R5708 VSS.n1140 VSS 0.238
R5709 VSS.n1138 VSS 0.238
R5710 VSS.n1132 VSS 0.238
R5711 VSS.n1126 VSS 0.238
R5712 VSS.n1124 VSS 0.238
R5713 VSS.n1118 VSS 0.238
R5714 VSS.n1112 VSS 0.238
R5715 VSS.n1110 VSS 0.238
R5716 VSS.n1104 VSS 0.238
R5717 VSS.n1098 VSS 0.238
R5718 VSS.n1096 VSS 0.238
R5719 VSS.n1090 VSS 0.238
R5720 VSS.n1084 VSS 0.238
R5721 VSS.n1082 VSS 0.238
R5722 VSS.n1076 VSS 0.238
R5723 VSS.n1070 VSS 0.238
R5724 VSS.n1068 VSS 0.238
R5725 VSS.n1062 VSS 0.238
R5726 VSS.n1048 VSS 0.238
R5727 VSS.n1042 VSS 0.238
R5728 VSS.n1036 VSS 0.238
R5729 VSS.n1034 VSS 0.238
R5730 VSS.n1028 VSS 0.238
R5731 VSS.n1022 VSS 0.238
R5732 VSS.n1020 VSS 0.238
R5733 VSS.n1014 VSS 0.238
R5734 VSS.n1008 VSS 0.238
R5735 VSS.n1006 VSS 0.238
R5736 VSS.n1000 VSS 0.238
R5737 VSS.n994 VSS 0.238
R5738 VSS.n992 VSS 0.238
R5739 VSS.n986 VSS 0.238
R5740 VSS.n980 VSS 0.238
R5741 VSS.n967 VSS 0.238
R5742 VSS.n961 VSS 0.238
R5743 VSS.n955 VSS 0.238
R5744 VSS.n953 VSS 0.238
R5745 VSS.n947 VSS 0.238
R5746 VSS.n941 VSS 0.238
R5747 VSS.n939 VSS 0.238
R5748 VSS.n926 VSS 0.238
R5749 VSS.n920 VSS 0.238
R5750 VSS.n914 VSS 0.238
R5751 VSS.n901 VSS 0.238
R5752 VSS.n111 VSS 0.178
R5753 VSS.n113 VSS 0.178
R5754 VSS.n121 VSS 0.178
R5755 VSS.n129 VSS 0.178
R5756 VSS.n131 VSS 0.178
R5757 VSS.n139 VSS 0.178
R5758 VSS.n147 VSS 0.178
R5759 VSS.n149 VSS 0.178
R5760 VSS.n157 VSS 0.178
R5761 VSS.n165 VSS 0.178
R5762 VSS.n167 VSS 0.178
R5763 VSS.n175 VSS 0.178
R5764 VSS.n183 VSS 0.178
R5765 VSS.n185 VSS 0.178
R5766 VSS.n193 VSS 0.178
R5767 VSS.n201 VSS 0.178
R5768 VSS.n203 VSS 0.178
R5769 VSS.n211 VSS 0.178
R5770 VSS.n219 VSS 0.178
R5771 VSS.n221 VSS 0.178
R5772 VSS.n229 VSS 0.178
R5773 VSS.n237 VSS 0.178
R5774 VSS.n239 VSS 0.178
R5775 VSS.n247 VSS 0.178
R5776 VSS.n255 VSS 0.178
R5777 VSS.n257 VSS 0.178
R5778 VSS.n265 VSS 0.178
R5779 VSS.n273 VSS 0.178
R5780 VSS.n275 VSS 0.178
R5781 VSS.n283 VSS 0.178
R5782 VSS.n291 VSS 0.178
R5783 VSS VSS.n586 0.178
R5784 VSS.n578 VSS 0.178
R5785 VSS VSS.n576 0.178
R5786 VSS VSS.n568 0.178
R5787 VSS.n560 VSS 0.178
R5788 VSS VSS.n558 0.178
R5789 VSS VSS.n550 0.178
R5790 VSS.n542 VSS 0.178
R5791 VSS VSS.n540 0.178
R5792 VSS VSS.n532 0.178
R5793 VSS.n524 VSS 0.178
R5794 VSS VSS.n522 0.178
R5795 VSS VSS.n514 0.178
R5796 VSS.n506 VSS 0.178
R5797 VSS VSS.n504 0.178
R5798 VSS VSS.n483 0.178
R5799 VSS.n475 VSS 0.178
R5800 VSS VSS.n473 0.178
R5801 VSS VSS.n465 0.178
R5802 VSS.n457 VSS 0.178
R5803 VSS VSS.n455 0.178
R5804 VSS VSS.n447 0.178
R5805 VSS VSS.n429 0.178
R5806 VSS.n421 VSS 0.178
R5807 VSS VSS.n419 0.178
R5808 VSS VSS.n400 0.178
R5809 VSS.n1196 VSS 0.178
R5810 VSS VSS.n1194 0.178
R5811 VSS VSS.n1188 0.178
R5812 VSS.n1182 VSS 0.178
R5813 VSS VSS.n1180 0.178
R5814 VSS VSS.n1174 0.178
R5815 VSS.n1168 VSS 0.178
R5816 VSS VSS.n1166 0.178
R5817 VSS VSS.n1160 0.178
R5818 VSS.n1154 VSS 0.178
R5819 VSS VSS.n1152 0.178
R5820 VSS VSS.n1146 0.178
R5821 VSS.n1140 VSS 0.178
R5822 VSS VSS.n1138 0.178
R5823 VSS VSS.n1132 0.178
R5824 VSS.n1126 VSS 0.178
R5825 VSS VSS.n1124 0.178
R5826 VSS VSS.n1118 0.178
R5827 VSS.n1112 VSS 0.178
R5828 VSS VSS.n1110 0.178
R5829 VSS VSS.n1104 0.178
R5830 VSS.n1098 VSS 0.178
R5831 VSS VSS.n1096 0.178
R5832 VSS VSS.n1090 0.178
R5833 VSS.n1084 VSS 0.178
R5834 VSS VSS.n1082 0.178
R5835 VSS VSS.n1076 0.178
R5836 VSS.n1070 VSS 0.178
R5837 VSS VSS.n1068 0.178
R5838 VSS VSS.n1062 0.178
R5839 VSS.n1056 VSS 0.178
R5840 VSS VSS.n1042 0.178
R5841 VSS.n1036 VSS 0.178
R5842 VSS VSS.n1034 0.178
R5843 VSS VSS.n1028 0.178
R5844 VSS.n1022 VSS 0.178
R5845 VSS VSS.n1020 0.178
R5846 VSS VSS.n1014 0.178
R5847 VSS.n1008 VSS 0.178
R5848 VSS VSS.n1006 0.178
R5849 VSS VSS.n1000 0.178
R5850 VSS.n994 VSS 0.178
R5851 VSS VSS.n992 0.178
R5852 VSS VSS.n986 0.178
R5853 VSS.n980 VSS 0.178
R5854 VSS VSS.n978 0.178
R5855 VSS VSS.n961 0.178
R5856 VSS.n955 VSS 0.178
R5857 VSS VSS.n953 0.178
R5858 VSS VSS.n947 0.178
R5859 VSS.n941 VSS 0.178
R5860 VSS VSS.n939 0.178
R5861 VSS VSS.n933 0.178
R5862 VSS VSS.n920 0.178
R5863 VSS.n914 VSS 0.178
R5864 VSS VSS.n912 0.178
R5865 VSS VSS.n895 0.178
R5866 VSS.n104 VSS 0.143
R5867 VSS VSS.n112 0.143
R5868 VSS VSS.n120 0.143
R5869 VSS.n122 VSS 0.143
R5870 VSS VSS.n130 0.143
R5871 VSS VSS.n138 0.143
R5872 VSS.n140 VSS 0.143
R5873 VSS VSS.n148 0.143
R5874 VSS VSS.n156 0.143
R5875 VSS.n158 VSS 0.143
R5876 VSS VSS.n166 0.143
R5877 VSS VSS.n174 0.143
R5878 VSS.n176 VSS 0.143
R5879 VSS VSS.n184 0.143
R5880 VSS VSS.n192 0.143
R5881 VSS.n194 VSS 0.143
R5882 VSS VSS.n202 0.143
R5883 VSS VSS.n210 0.143
R5884 VSS.n212 VSS 0.143
R5885 VSS VSS.n220 0.143
R5886 VSS VSS.n228 0.143
R5887 VSS.n230 VSS 0.143
R5888 VSS VSS.n238 0.143
R5889 VSS VSS.n246 0.143
R5890 VSS.n248 VSS 0.143
R5891 VSS VSS.n256 0.143
R5892 VSS VSS.n264 0.143
R5893 VSS.n266 VSS 0.143
R5894 VSS VSS.n274 0.143
R5895 VSS VSS.n282 0.143
R5896 VSS.n284 VSS 0.143
R5897 VSS.n596 VSS 0.143
R5898 VSS.n587 VSS 0.143
R5899 VSS.n585 VSS 0.143
R5900 VSS.n577 VSS 0.143
R5901 VSS.n569 VSS 0.143
R5902 VSS.n567 VSS 0.143
R5903 VSS.n559 VSS 0.143
R5904 VSS.n551 VSS 0.143
R5905 VSS.n549 VSS 0.143
R5906 VSS.n541 VSS 0.143
R5907 VSS.n533 VSS 0.143
R5908 VSS.n531 VSS 0.143
R5909 VSS.n523 VSS 0.143
R5910 VSS.n515 VSS 0.143
R5911 VSS.n513 VSS 0.143
R5912 VSS.n505 VSS 0.143
R5913 VSS.n500 VSS 0.143
R5914 VSS.n484 VSS 0.143
R5915 VSS.n482 VSS 0.143
R5916 VSS.n474 VSS 0.143
R5917 VSS.n466 VSS 0.143
R5918 VSS.n464 VSS 0.143
R5919 VSS.n456 VSS 0.143
R5920 VSS.n448 VSS 0.143
R5921 VSS.n446 VSS 0.143
R5922 VSS.n430 VSS 0.143
R5923 VSS.n428 VSS 0.143
R5924 VSS.n420 VSS 0.143
R5925 VSS.n415 VSS 0.143
R5926 VSS.n401 VSS 0.143
R5927 VSS.n399 VSS 0.143
R5928 VSS.n386 VSS 0.143
R5929 VSS.n377 VSS 0.143
R5930 VSS.n1201 VSS 0.143
R5931 VSS.n1195 VSS 0.143
R5932 VSS.n1189 VSS 0.143
R5933 VSS.n1187 VSS 0.143
R5934 VSS.n1181 VSS 0.143
R5935 VSS.n1175 VSS 0.143
R5936 VSS.n1173 VSS 0.143
R5937 VSS.n1167 VSS 0.143
R5938 VSS.n1161 VSS 0.143
R5939 VSS.n1159 VSS 0.143
R5940 VSS.n1153 VSS 0.143
R5941 VSS.n1147 VSS 0.143
R5942 VSS.n1145 VSS 0.143
R5943 VSS.n1139 VSS 0.143
R5944 VSS.n1133 VSS 0.143
R5945 VSS.n1131 VSS 0.143
R5946 VSS.n1125 VSS 0.143
R5947 VSS.n1119 VSS 0.143
R5948 VSS.n1117 VSS 0.143
R5949 VSS.n1111 VSS 0.143
R5950 VSS.n1105 VSS 0.143
R5951 VSS.n1103 VSS 0.143
R5952 VSS.n1097 VSS 0.143
R5953 VSS.n1091 VSS 0.143
R5954 VSS.n1089 VSS 0.143
R5955 VSS.n1083 VSS 0.143
R5956 VSS.n1077 VSS 0.143
R5957 VSS.n1075 VSS 0.143
R5958 VSS.n1069 VSS 0.143
R5959 VSS.n1063 VSS 0.143
R5960 VSS.n1061 VSS 0.143
R5961 VSS.n1055 VSS 0.143
R5962 VSS.n1043 VSS 0.143
R5963 VSS.n1041 VSS 0.143
R5964 VSS.n1035 VSS 0.143
R5965 VSS.n1029 VSS 0.143
R5966 VSS.n1027 VSS 0.143
R5967 VSS.n1021 VSS 0.143
R5968 VSS.n1015 VSS 0.143
R5969 VSS.n1013 VSS 0.143
R5970 VSS.n1007 VSS 0.143
R5971 VSS.n1001 VSS 0.143
R5972 VSS.n999 VSS 0.143
R5973 VSS.n993 VSS 0.143
R5974 VSS.n987 VSS 0.143
R5975 VSS.n985 VSS 0.143
R5976 VSS.n979 VSS 0.143
R5977 VSS.n974 VSS 0.143
R5978 VSS.n962 VSS 0.143
R5979 VSS.n960 VSS 0.143
R5980 VSS.n954 VSS 0.143
R5981 VSS.n948 VSS 0.143
R5982 VSS.n946 VSS 0.143
R5983 VSS.n940 VSS 0.143
R5984 VSS.n934 VSS 0.143
R5985 VSS.n932 VSS 0.143
R5986 VSS.n921 VSS 0.143
R5987 VSS.n919 VSS 0.143
R5988 VSS.n913 VSS 0.143
R5989 VSS.n908 VSS 0.143
R5990 VSS.n896 VSS 0.143
R5991 VSS.n894 VSS 0.143
R5992 VSS.n884 VSS 0.143
R5993 VSS.n877 VSS 0.143
R5994 VSS.n102 VSS 0.083
R5995 VSS.n104 VSS 0.083
R5996 VSS.n112 VSS 0.083
R5997 VSS.n120 VSS 0.083
R5998 VSS.n122 VSS 0.083
R5999 VSS.n130 VSS 0.083
R6000 VSS.n138 VSS 0.083
R6001 VSS.n140 VSS 0.083
R6002 VSS.n148 VSS 0.083
R6003 VSS.n156 VSS 0.083
R6004 VSS.n158 VSS 0.083
R6005 VSS.n166 VSS 0.083
R6006 VSS.n174 VSS 0.083
R6007 VSS.n176 VSS 0.083
R6008 VSS.n184 VSS 0.083
R6009 VSS.n192 VSS 0.083
R6010 VSS.n194 VSS 0.083
R6011 VSS.n202 VSS 0.083
R6012 VSS.n210 VSS 0.083
R6013 VSS.n212 VSS 0.083
R6014 VSS.n220 VSS 0.083
R6015 VSS.n228 VSS 0.083
R6016 VSS.n230 VSS 0.083
R6017 VSS.n238 VSS 0.083
R6018 VSS.n246 VSS 0.083
R6019 VSS.n248 VSS 0.083
R6020 VSS.n256 VSS 0.083
R6021 VSS.n264 VSS 0.083
R6022 VSS.n266 VSS 0.083
R6023 VSS.n274 VSS 0.083
R6024 VSS.n282 VSS 0.083
R6025 VSS.n284 VSS 0.083
R6026 VSS VSS.n595 0.083
R6027 VSS.n587 VSS 0.083
R6028 VSS VSS.n585 0.083
R6029 VSS VSS.n577 0.083
R6030 VSS.n569 VSS 0.083
R6031 VSS VSS.n567 0.083
R6032 VSS VSS.n559 0.083
R6033 VSS.n551 VSS 0.083
R6034 VSS VSS.n549 0.083
R6035 VSS VSS.n541 0.083
R6036 VSS.n533 VSS 0.083
R6037 VSS VSS.n531 0.083
R6038 VSS VSS.n523 0.083
R6039 VSS.n515 VSS 0.083
R6040 VSS VSS.n513 0.083
R6041 VSS VSS.n505 0.083
R6042 VSS.n492 VSS 0.083
R6043 VSS.n484 VSS 0.083
R6044 VSS VSS.n482 0.083
R6045 VSS VSS.n474 0.083
R6046 VSS.n466 VSS 0.083
R6047 VSS VSS.n464 0.083
R6048 VSS VSS.n456 0.083
R6049 VSS.n448 VSS 0.083
R6050 VSS.n438 VSS 0.083
R6051 VSS.n430 VSS 0.083
R6052 VSS VSS.n428 0.083
R6053 VSS VSS.n420 0.083
R6054 VSS.n407 VSS 0.083
R6055 VSS.n401 VSS 0.083
R6056 VSS.n391 VSS 0.083
R6057 VSS.n604 VSS 0.083
R6058 VSS VSS.n1201 0.083
R6059 VSS VSS.n1195 0.083
R6060 VSS.n1189 VSS 0.083
R6061 VSS VSS.n1187 0.083
R6062 VSS VSS.n1181 0.083
R6063 VSS.n1175 VSS 0.083
R6064 VSS VSS.n1173 0.083
R6065 VSS VSS.n1167 0.083
R6066 VSS.n1161 VSS 0.083
R6067 VSS VSS.n1159 0.083
R6068 VSS VSS.n1153 0.083
R6069 VSS.n1147 VSS 0.083
R6070 VSS VSS.n1145 0.083
R6071 VSS VSS.n1139 0.083
R6072 VSS.n1133 VSS 0.083
R6073 VSS VSS.n1131 0.083
R6074 VSS VSS.n1125 0.083
R6075 VSS.n1119 VSS 0.083
R6076 VSS VSS.n1117 0.083
R6077 VSS VSS.n1111 0.083
R6078 VSS.n1105 VSS 0.083
R6079 VSS VSS.n1103 0.083
R6080 VSS VSS.n1097 0.083
R6081 VSS.n1091 VSS 0.083
R6082 VSS VSS.n1089 0.083
R6083 VSS VSS.n1083 0.083
R6084 VSS.n1077 VSS 0.083
R6085 VSS VSS.n1075 0.083
R6086 VSS VSS.n1069 0.083
R6087 VSS.n1063 VSS 0.083
R6088 VSS VSS.n1061 0.083
R6089 VSS.n1049 VSS 0.083
R6090 VSS.n1043 VSS 0.083
R6091 VSS VSS.n1041 0.083
R6092 VSS VSS.n1035 0.083
R6093 VSS.n1029 VSS 0.083
R6094 VSS VSS.n1027 0.083
R6095 VSS VSS.n1021 0.083
R6096 VSS.n1015 VSS 0.083
R6097 VSS VSS.n1013 0.083
R6098 VSS VSS.n1007 0.083
R6099 VSS.n1001 VSS 0.083
R6100 VSS VSS.n999 0.083
R6101 VSS VSS.n993 0.083
R6102 VSS.n987 VSS 0.083
R6103 VSS VSS.n985 0.083
R6104 VSS VSS.n979 0.083
R6105 VSS.n968 VSS 0.083
R6106 VSS.n962 VSS 0.083
R6107 VSS VSS.n960 0.083
R6108 VSS VSS.n954 0.083
R6109 VSS.n948 VSS 0.083
R6110 VSS VSS.n946 0.083
R6111 VSS VSS.n940 0.083
R6112 VSS.n934 VSS 0.083
R6113 VSS.n927 VSS 0.083
R6114 VSS.n921 VSS 0.083
R6115 VSS VSS.n919 0.083
R6116 VSS VSS.n913 0.083
R6117 VSS.n902 VSS 0.083
R6118 VSS.n896 VSS 0.083
R6119 VSS.n889 VSS 0.083
R6120 VSS.n96 VSS.n95 0.00170947
R6121 VSS.n95 VSS.n94 0.00170947
R6122 VSS.n107 VSS.n106 0.00170947
R6123 VSS.n106 VSS.n105 0.00170947
R6124 VSS.n110 VSS.n109 0.00170947
R6125 VSS.n109 VSS.n108 0.00170947
R6126 VSS.n92 VSS.n91 0.00170947
R6127 VSS.n91 VSS.n90 0.00170947
R6128 VSS.n116 VSS.n115 0.00170947
R6129 VSS.n115 VSS.n114 0.00170947
R6130 VSS.n119 VSS.n118 0.00170947
R6131 VSS.n118 VSS.n117 0.00170947
R6132 VSS.n87 VSS.n86 0.00170947
R6133 VSS.n86 VSS.n85 0.00170947
R6134 VSS.n125 VSS.n124 0.00170947
R6135 VSS.n124 VSS.n123 0.00170947
R6136 VSS.n128 VSS.n127 0.00170947
R6137 VSS.n127 VSS.n126 0.00170947
R6138 VSS.n83 VSS.n82 0.00170947
R6139 VSS.n82 VSS.n81 0.00170947
R6140 VSS.n134 VSS.n133 0.00170947
R6141 VSS.n133 VSS.n132 0.00170947
R6142 VSS.n137 VSS.n136 0.00170947
R6143 VSS.n136 VSS.n135 0.00170947
R6144 VSS.n78 VSS.n77 0.00170947
R6145 VSS.n77 VSS.n76 0.00170947
R6146 VSS.n143 VSS.n142 0.00170947
R6147 VSS.n142 VSS.n141 0.00170947
R6148 VSS.n146 VSS.n145 0.00170947
R6149 VSS.n145 VSS.n144 0.00170947
R6150 VSS.n74 VSS.n73 0.00170947
R6151 VSS.n73 VSS.n72 0.00170947
R6152 VSS.n152 VSS.n151 0.00170947
R6153 VSS.n151 VSS.n150 0.00170947
R6154 VSS.n155 VSS.n154 0.00170947
R6155 VSS.n154 VSS.n153 0.00170947
R6156 VSS.n69 VSS.n68 0.00170947
R6157 VSS.n68 VSS.n67 0.00170947
R6158 VSS.n161 VSS.n160 0.00170947
R6159 VSS.n160 VSS.n159 0.00170947
R6160 VSS.n164 VSS.n163 0.00170947
R6161 VSS.n163 VSS.n162 0.00170947
R6162 VSS.n65 VSS.n64 0.00170947
R6163 VSS.n64 VSS.n63 0.00170947
R6164 VSS.n170 VSS.n169 0.00170947
R6165 VSS.n169 VSS.n168 0.00170947
R6166 VSS.n173 VSS.n172 0.00170947
R6167 VSS.n172 VSS.n171 0.00170947
R6168 VSS.n60 VSS.n59 0.00170947
R6169 VSS.n59 VSS.n58 0.00170947
R6170 VSS.n179 VSS.n178 0.00170947
R6171 VSS.n178 VSS.n177 0.00170947
R6172 VSS.n182 VSS.n181 0.00170947
R6173 VSS.n181 VSS.n180 0.00170947
R6174 VSS.n56 VSS.n55 0.00170947
R6175 VSS.n55 VSS.n54 0.00170947
R6176 VSS.n188 VSS.n187 0.00170947
R6177 VSS.n187 VSS.n186 0.00170947
R6178 VSS.n191 VSS.n190 0.00170947
R6179 VSS.n190 VSS.n189 0.00170947
R6180 VSS.n51 VSS.n50 0.00170947
R6181 VSS.n50 VSS.n49 0.00170947
R6182 VSS.n197 VSS.n196 0.00170947
R6183 VSS.n196 VSS.n195 0.00170947
R6184 VSS.n200 VSS.n199 0.00170947
R6185 VSS.n199 VSS.n198 0.00170947
R6186 VSS.n47 VSS.n46 0.00170947
R6187 VSS.n46 VSS.n45 0.00170947
R6188 VSS.n206 VSS.n205 0.00170947
R6189 VSS.n205 VSS.n204 0.00170947
R6190 VSS.n209 VSS.n208 0.00170947
R6191 VSS.n208 VSS.n207 0.00170947
R6192 VSS.n42 VSS.n41 0.00170947
R6193 VSS.n41 VSS.n40 0.00170947
R6194 VSS.n215 VSS.n214 0.00170947
R6195 VSS.n214 VSS.n213 0.00170947
R6196 VSS.n218 VSS.n217 0.00170947
R6197 VSS.n217 VSS.n216 0.00170947
R6198 VSS.n38 VSS.n37 0.00170947
R6199 VSS.n37 VSS.n36 0.00170947
R6200 VSS.n224 VSS.n223 0.00170947
R6201 VSS.n223 VSS.n222 0.00170947
R6202 VSS.n227 VSS.n226 0.00170947
R6203 VSS.n226 VSS.n225 0.00170947
R6204 VSS.n33 VSS.n32 0.00170947
R6205 VSS.n32 VSS.n31 0.00170947
R6206 VSS.n233 VSS.n232 0.00170947
R6207 VSS.n232 VSS.n231 0.00170947
R6208 VSS.n236 VSS.n235 0.00170947
R6209 VSS.n235 VSS.n234 0.00170947
R6210 VSS.n29 VSS.n28 0.00170947
R6211 VSS.n28 VSS.n27 0.00170947
R6212 VSS.n242 VSS.n241 0.00170947
R6213 VSS.n241 VSS.n240 0.00170947
R6214 VSS.n245 VSS.n244 0.00170947
R6215 VSS.n244 VSS.n243 0.00170947
R6216 VSS.n24 VSS.n23 0.00170947
R6217 VSS.n23 VSS.n22 0.00170947
R6218 VSS.n251 VSS.n250 0.00170947
R6219 VSS.n250 VSS.n249 0.00170947
R6220 VSS.n254 VSS.n253 0.00170947
R6221 VSS.n253 VSS.n252 0.00170947
R6222 VSS.n20 VSS.n19 0.00170947
R6223 VSS.n19 VSS.n18 0.00170947
R6224 VSS.n260 VSS.n259 0.00170947
R6225 VSS.n259 VSS.n258 0.00170947
R6226 VSS.n263 VSS.n262 0.00170947
R6227 VSS.n262 VSS.n261 0.00170947
R6228 VSS.n15 VSS.n14 0.00170947
R6229 VSS.n14 VSS.n13 0.00170947
R6230 VSS.n269 VSS.n268 0.00170947
R6231 VSS.n268 VSS.n267 0.00170947
R6232 VSS.n272 VSS.n271 0.00170947
R6233 VSS.n271 VSS.n270 0.00170947
R6234 VSS.n11 VSS.n10 0.00170947
R6235 VSS.n10 VSS.n9 0.00170947
R6236 VSS.n278 VSS.n277 0.00170947
R6237 VSS.n277 VSS.n276 0.00170947
R6238 VSS.n281 VSS.n280 0.00170947
R6239 VSS.n280 VSS.n279 0.00170947
R6240 VSS.n6 VSS.n5 0.00170947
R6241 VSS.n5 VSS.n4 0.00170947
R6242 VSS.n287 VSS.n286 0.00170947
R6243 VSS.n286 VSS.n285 0.00170947
R6244 VSS.n290 VSS.n289 0.00170947
R6245 VSS.n289 VSS.n288 0.00170947
R6246 VSS.n598 VSS.n597 0.00170947
R6247 VSS.n599 VSS.n598 0.00170947
R6248 VSS.n101 VSS.n100 0.00170947
R6249 VSS.n100 VSS.n99 0.00170947
R6250 VSS.n405 VSS.n369 0.00170947
R6251 VSS.n369 VSS.n368 0.00170947
R6252 VSS.n389 VSS.n388 0.00170947
R6253 VSS.n388 VSS.n387 0.00170947
R6254 VSS.n385 VSS.n384 0.00170947
R6255 VSS.n384 VSS.n383 0.00170947
R6256 VSS.n381 VSS.n380 0.00170947
R6257 VSS.n380 VSS.n379 0.00170947
R6258 VSS.n376 VSS.n375 0.00170947
R6259 VSS.n375 VSS.n374 0.00170947
R6260 VSS.n394 VSS.n393 0.00170947
R6261 VSS.n393 VSS.n392 0.00170947
R6262 VSS.n404 VSS.n403 0.00170947
R6263 VSS.n403 VSS.n402 0.00170947
R6264 VSS.n372 VSS.n371 0.00170947
R6265 VSS.n371 VSS.n370 0.00170947
R6266 VSS.n398 VSS.n397 0.00170947
R6267 VSS.n397 VSS.n396 0.00170947
R6268 VSS.n410 VSS.n409 0.00170947
R6269 VSS.n409 VSS.n408 0.00170947
R6270 VSS.n3 VSS.n2 0.00170947
R6271 VSS.n2 VSS.n1 0.00170947
R6272 VSS.n593 VSS.n592 0.00170947
R6273 VSS.n592 VSS.n591 0.00170947
R6274 VSS.n590 VSS.n589 0.00170947
R6275 VSS.n589 VSS.n588 0.00170947
R6276 VSS.n294 VSS.n293 0.00170947
R6277 VSS.n293 VSS.n292 0.00170947
R6278 VSS.n584 VSS.n583 0.00170947
R6279 VSS.n583 VSS.n582 0.00170947
R6280 VSS.n581 VSS.n580 0.00170947
R6281 VSS.n580 VSS.n579 0.00170947
R6282 VSS.n299 VSS.n298 0.00170947
R6283 VSS.n298 VSS.n297 0.00170947
R6284 VSS.n575 VSS.n574 0.00170947
R6285 VSS.n574 VSS.n573 0.00170947
R6286 VSS.n572 VSS.n571 0.00170947
R6287 VSS.n571 VSS.n570 0.00170947
R6288 VSS.n303 VSS.n302 0.00170947
R6289 VSS.n302 VSS.n301 0.00170947
R6290 VSS.n566 VSS.n565 0.00170947
R6291 VSS.n565 VSS.n564 0.00170947
R6292 VSS.n563 VSS.n562 0.00170947
R6293 VSS.n562 VSS.n561 0.00170947
R6294 VSS.n308 VSS.n307 0.00170947
R6295 VSS.n307 VSS.n306 0.00170947
R6296 VSS.n557 VSS.n556 0.00170947
R6297 VSS.n556 VSS.n555 0.00170947
R6298 VSS.n554 VSS.n553 0.00170947
R6299 VSS.n553 VSS.n552 0.00170947
R6300 VSS.n312 VSS.n311 0.00170947
R6301 VSS.n311 VSS.n310 0.00170947
R6302 VSS.n548 VSS.n547 0.00170947
R6303 VSS.n547 VSS.n546 0.00170947
R6304 VSS.n545 VSS.n544 0.00170947
R6305 VSS.n544 VSS.n543 0.00170947
R6306 VSS.n317 VSS.n316 0.00170947
R6307 VSS.n316 VSS.n315 0.00170947
R6308 VSS.n539 VSS.n538 0.00170947
R6309 VSS.n538 VSS.n537 0.00170947
R6310 VSS.n535 VSS.n534 0.00170947
R6311 VSS.n536 VSS.n535 0.00170947
R6312 VSS.n321 VSS.n320 0.00170947
R6313 VSS.n320 VSS.n319 0.00170947
R6314 VSS.n530 VSS.n529 0.00170947
R6315 VSS.n529 VSS.n528 0.00170947
R6316 VSS.n527 VSS.n526 0.00170947
R6317 VSS.n526 VSS.n525 0.00170947
R6318 VSS.n326 VSS.n325 0.00170947
R6319 VSS.n325 VSS.n324 0.00170947
R6320 VSS.n521 VSS.n520 0.00170947
R6321 VSS.n520 VSS.n519 0.00170947
R6322 VSS.n518 VSS.n517 0.00170947
R6323 VSS.n517 VSS.n516 0.00170947
R6324 VSS.n330 VSS.n329 0.00170947
R6325 VSS.n329 VSS.n328 0.00170947
R6326 VSS.n512 VSS.n511 0.00170947
R6327 VSS.n511 VSS.n510 0.00170947
R6328 VSS.n509 VSS.n508 0.00170947
R6329 VSS.n508 VSS.n507 0.00170947
R6330 VSS.n335 VSS.n334 0.00170947
R6331 VSS.n334 VSS.n333 0.00170947
R6332 VSS.n503 VSS.n502 0.00170947
R6333 VSS.n502 VSS.n501 0.00170947
R6334 VSS.n499 VSS.n498 0.00170947
R6335 VSS.n498 VSS.n497 0.00170947
R6336 VSS.n495 VSS.n494 0.00170947
R6337 VSS.n494 VSS.n493 0.00170947
R6338 VSS.n490 VSS.n489 0.00170947
R6339 VSS.n489 VSS.n488 0.00170947
R6340 VSS.n487 VSS.n486 0.00170947
R6341 VSS.n486 VSS.n485 0.00170947
R6342 VSS.n339 VSS.n338 0.00170947
R6343 VSS.n338 VSS.n337 0.00170947
R6344 VSS.n481 VSS.n480 0.00170947
R6345 VSS.n480 VSS.n479 0.00170947
R6346 VSS.n478 VSS.n477 0.00170947
R6347 VSS.n477 VSS.n476 0.00170947
R6348 VSS.n344 VSS.n343 0.00170947
R6349 VSS.n343 VSS.n342 0.00170947
R6350 VSS.n472 VSS.n471 0.00170947
R6351 VSS.n471 VSS.n470 0.00170947
R6352 VSS.n469 VSS.n468 0.00170947
R6353 VSS.n468 VSS.n467 0.00170947
R6354 VSS.n348 VSS.n347 0.00170947
R6355 VSS.n347 VSS.n346 0.00170947
R6356 VSS.n463 VSS.n462 0.00170947
R6357 VSS.n462 VSS.n461 0.00170947
R6358 VSS.n460 VSS.n459 0.00170947
R6359 VSS.n459 VSS.n458 0.00170947
R6360 VSS.n353 VSS.n352 0.00170947
R6361 VSS.n352 VSS.n351 0.00170947
R6362 VSS.n454 VSS.n453 0.00170947
R6363 VSS.n453 VSS.n452 0.00170947
R6364 VSS.n451 VSS.n450 0.00170947
R6365 VSS.n450 VSS.n449 0.00170947
R6366 VSS.n357 VSS.n356 0.00170947
R6367 VSS.n356 VSS.n355 0.00170947
R6368 VSS.n445 VSS.n444 0.00170947
R6369 VSS.n444 VSS.n443 0.00170947
R6370 VSS.n441 VSS.n440 0.00170947
R6371 VSS.n440 VSS.n439 0.00170947
R6372 VSS.n436 VSS.n435 0.00170947
R6373 VSS.n435 VSS.n434 0.00170947
R6374 VSS.n433 VSS.n432 0.00170947
R6375 VSS.n432 VSS.n431 0.00170947
R6376 VSS.n361 VSS.n360 0.00170947
R6377 VSS.n360 VSS.n359 0.00170947
R6378 VSS.n427 VSS.n426 0.00170947
R6379 VSS.n426 VSS.n425 0.00170947
R6380 VSS.n424 VSS.n423 0.00170947
R6381 VSS.n423 VSS.n422 0.00170947
R6382 VSS.n366 VSS.n365 0.00170947
R6383 VSS.n365 VSS.n364 0.00170947
R6384 VSS.n418 VSS.n417 0.00170947
R6385 VSS.n417 VSS.n416 0.00170947
R6386 VSS.n414 VSS.n413 0.00170947
R6387 VSS.n413 VSS.n412 0.00170947
R6388 VSS.n883 VSS.n882 0.00170947
R6389 VSS.n882 VSS.n881 0.00170947
R6390 VSS.n907 VSS.n906 0.00170947
R6391 VSS.n906 VSS.n905 0.00170947
R6392 VSS.n973 VSS.n972 0.00170947
R6393 VSS.n972 VSS.n971 0.00170947
R6394 VSS.n603 VSS.n602 0.00170947
R6395 VSS.n602 VSS.n601 0.00170947
R6396 VSS.n969 VSS.n812 0.00170947
R6397 VSS.n812 VSS.n811 0.00170947
R6398 VSS.n903 VSS.n862 0.00170947
R6399 VSS.n862 VSS.n861 0.00170947
R6400 VSS.n879 VSS.n873 0.00170947
R6401 VSS.n873 VSS.n872 0.00170947
R6402 VSS.n607 VSS.n606 0.00170947
R6403 VSS.n606 VSS.n605 0.00170947
R6404 VSS.n1200 VSS.n611 0.00170947
R6405 VSS.n611 VSS.n610 0.00170947
R6406 VSS.n1199 VSS.n1198 0.00170947
R6407 VSS.n1198 VSS.n1197 0.00170947
R6408 VSS.n614 VSS.n613 0.00170947
R6409 VSS.n613 VSS.n612 0.00170947
R6410 VSS.n1193 VSS.n1192 0.00170947
R6411 VSS.n1192 VSS.n1191 0.00170947
R6412 VSS.n1190 VSS.n617 0.00170947
R6413 VSS.n617 VSS.n616 0.00170947
R6414 VSS.n620 VSS.n619 0.00170947
R6415 VSS.n619 VSS.n618 0.00170947
R6416 VSS.n1186 VSS.n624 0.00170947
R6417 VSS.n624 VSS.n623 0.00170947
R6418 VSS.n1185 VSS.n1184 0.00170947
R6419 VSS.n1184 VSS.n1183 0.00170947
R6420 VSS.n627 VSS.n626 0.00170947
R6421 VSS.n626 VSS.n625 0.00170947
R6422 VSS.n1179 VSS.n1178 0.00170947
R6423 VSS.n1178 VSS.n1177 0.00170947
R6424 VSS.n1176 VSS.n630 0.00170947
R6425 VSS.n630 VSS.n629 0.00170947
R6426 VSS.n633 VSS.n632 0.00170947
R6427 VSS.n632 VSS.n631 0.00170947
R6428 VSS.n1172 VSS.n637 0.00170947
R6429 VSS.n637 VSS.n636 0.00170947
R6430 VSS.n1171 VSS.n1170 0.00170947
R6431 VSS.n1170 VSS.n1169 0.00170947
R6432 VSS.n640 VSS.n639 0.00170947
R6433 VSS.n639 VSS.n638 0.00170947
R6434 VSS.n1165 VSS.n1164 0.00170947
R6435 VSS.n1164 VSS.n1163 0.00170947
R6436 VSS.n1162 VSS.n643 0.00170947
R6437 VSS.n643 VSS.n642 0.00170947
R6438 VSS.n646 VSS.n645 0.00170947
R6439 VSS.n645 VSS.n644 0.00170947
R6440 VSS.n1158 VSS.n650 0.00170947
R6441 VSS.n650 VSS.n649 0.00170947
R6442 VSS.n1157 VSS.n1156 0.00170947
R6443 VSS.n1156 VSS.n1155 0.00170947
R6444 VSS.n653 VSS.n652 0.00170947
R6445 VSS.n652 VSS.n651 0.00170947
R6446 VSS.n1151 VSS.n1150 0.00170947
R6447 VSS.n1150 VSS.n1149 0.00170947
R6448 VSS.n1148 VSS.n656 0.00170947
R6449 VSS.n656 VSS.n655 0.00170947
R6450 VSS.n659 VSS.n658 0.00170947
R6451 VSS.n658 VSS.n657 0.00170947
R6452 VSS.n1144 VSS.n663 0.00170947
R6453 VSS.n663 VSS.n662 0.00170947
R6454 VSS.n1143 VSS.n1142 0.00170947
R6455 VSS.n1142 VSS.n1141 0.00170947
R6456 VSS.n666 VSS.n665 0.00170947
R6457 VSS.n665 VSS.n664 0.00170947
R6458 VSS.n1137 VSS.n1136 0.00170947
R6459 VSS.n1136 VSS.n1135 0.00170947
R6460 VSS.n1134 VSS.n669 0.00170947
R6461 VSS.n669 VSS.n668 0.00170947
R6462 VSS.n672 VSS.n671 0.00170947
R6463 VSS.n671 VSS.n670 0.00170947
R6464 VSS.n1130 VSS.n676 0.00170947
R6465 VSS.n676 VSS.n675 0.00170947
R6466 VSS.n1129 VSS.n1128 0.00170947
R6467 VSS.n1128 VSS.n1127 0.00170947
R6468 VSS.n679 VSS.n678 0.00170947
R6469 VSS.n678 VSS.n677 0.00170947
R6470 VSS.n1123 VSS.n1122 0.00170947
R6471 VSS.n1122 VSS.n1121 0.00170947
R6472 VSS.n1120 VSS.n682 0.00170947
R6473 VSS.n682 VSS.n681 0.00170947
R6474 VSS.n685 VSS.n684 0.00170947
R6475 VSS.n684 VSS.n683 0.00170947
R6476 VSS.n1116 VSS.n689 0.00170947
R6477 VSS.n689 VSS.n688 0.00170947
R6478 VSS.n1115 VSS.n1114 0.00170947
R6479 VSS.n1114 VSS.n1113 0.00170947
R6480 VSS.n692 VSS.n691 0.00170947
R6481 VSS.n691 VSS.n690 0.00170947
R6482 VSS.n1109 VSS.n1108 0.00170947
R6483 VSS.n1108 VSS.n1107 0.00170947
R6484 VSS.n1106 VSS.n695 0.00170947
R6485 VSS.n695 VSS.n694 0.00170947
R6486 VSS.n698 VSS.n697 0.00170947
R6487 VSS.n697 VSS.n696 0.00170947
R6488 VSS.n1102 VSS.n702 0.00170947
R6489 VSS.n702 VSS.n701 0.00170947
R6490 VSS.n1101 VSS.n1100 0.00170947
R6491 VSS.n1100 VSS.n1099 0.00170947
R6492 VSS.n705 VSS.n704 0.00170947
R6493 VSS.n704 VSS.n703 0.00170947
R6494 VSS.n1095 VSS.n1094 0.00170947
R6495 VSS.n1094 VSS.n1093 0.00170947
R6496 VSS.n1092 VSS.n708 0.00170947
R6497 VSS.n708 VSS.n707 0.00170947
R6498 VSS.n711 VSS.n710 0.00170947
R6499 VSS.n710 VSS.n709 0.00170947
R6500 VSS.n1088 VSS.n715 0.00170947
R6501 VSS.n715 VSS.n714 0.00170947
R6502 VSS.n1087 VSS.n1086 0.00170947
R6503 VSS.n1086 VSS.n1085 0.00170947
R6504 VSS.n718 VSS.n717 0.00170947
R6505 VSS.n717 VSS.n716 0.00170947
R6506 VSS.n1081 VSS.n1080 0.00170947
R6507 VSS.n1080 VSS.n1079 0.00170947
R6508 VSS.n1078 VSS.n721 0.00170947
R6509 VSS.n721 VSS.n720 0.00170947
R6510 VSS.n724 VSS.n723 0.00170947
R6511 VSS.n723 VSS.n722 0.00170947
R6512 VSS.n1074 VSS.n728 0.00170947
R6513 VSS.n728 VSS.n727 0.00170947
R6514 VSS.n1073 VSS.n1072 0.00170947
R6515 VSS.n1072 VSS.n1071 0.00170947
R6516 VSS.n731 VSS.n730 0.00170947
R6517 VSS.n730 VSS.n729 0.00170947
R6518 VSS.n1067 VSS.n1066 0.00170947
R6519 VSS.n1066 VSS.n1065 0.00170947
R6520 VSS.n1064 VSS.n734 0.00170947
R6521 VSS.n734 VSS.n733 0.00170947
R6522 VSS.n737 VSS.n736 0.00170947
R6523 VSS.n736 VSS.n735 0.00170947
R6524 VSS.n1060 VSS.n741 0.00170947
R6525 VSS.n741 VSS.n740 0.00170947
R6526 VSS.n1059 VSS.n1058 0.00170947
R6527 VSS.n1058 VSS.n1057 0.00170947
R6528 VSS.n1054 VSS.n744 0.00170947
R6529 VSS.n744 VSS.n743 0.00170947
R6530 VSS.n1053 VSS.n1052 0.00170947
R6531 VSS.n1052 VSS.n1051 0.00170947
R6532 VSS.n1047 VSS.n746 0.00170947
R6533 VSS.n746 VSS.n745 0.00170947
R6534 VSS.n1046 VSS.n1045 0.00170947
R6535 VSS.n1045 VSS.n1044 0.00170947
R6536 VSS.n749 VSS.n748 0.00170947
R6537 VSS.n748 VSS.n747 0.00170947
R6538 VSS.n1040 VSS.n1039 0.00170947
R6539 VSS.n1039 VSS.n1038 0.00170947
R6540 VSS.n1037 VSS.n753 0.00170947
R6541 VSS.n753 VSS.n752 0.00170947
R6542 VSS.n756 VSS.n755 0.00170947
R6543 VSS.n755 VSS.n754 0.00170947
R6544 VSS.n1033 VSS.n759 0.00170947
R6545 VSS.n759 VSS.n758 0.00170947
R6546 VSS.n1032 VSS.n1031 0.00170947
R6547 VSS.n1031 VSS.n1030 0.00170947
R6548 VSS.n762 VSS.n761 0.00170947
R6549 VSS.n761 VSS.n760 0.00170947
R6550 VSS.n1026 VSS.n1025 0.00170947
R6551 VSS.n1025 VSS.n1024 0.00170947
R6552 VSS.n1023 VSS.n766 0.00170947
R6553 VSS.n766 VSS.n765 0.00170947
R6554 VSS.n769 VSS.n768 0.00170947
R6555 VSS.n768 VSS.n767 0.00170947
R6556 VSS.n1019 VSS.n772 0.00170947
R6557 VSS.n772 VSS.n771 0.00170947
R6558 VSS.n1018 VSS.n1017 0.00170947
R6559 VSS.n1017 VSS.n1016 0.00170947
R6560 VSS.n775 VSS.n774 0.00170947
R6561 VSS.n774 VSS.n773 0.00170947
R6562 VSS.n1012 VSS.n1011 0.00170947
R6563 VSS.n1011 VSS.n1010 0.00170947
R6564 VSS.n1009 VSS.n779 0.00170947
R6565 VSS.n779 VSS.n778 0.00170947
R6566 VSS.n782 VSS.n781 0.00170947
R6567 VSS.n781 VSS.n780 0.00170947
R6568 VSS.n1005 VSS.n785 0.00170947
R6569 VSS.n785 VSS.n784 0.00170947
R6570 VSS.n1004 VSS.n1003 0.00170947
R6571 VSS.n1003 VSS.n1002 0.00170947
R6572 VSS.n788 VSS.n787 0.00170947
R6573 VSS.n787 VSS.n786 0.00170947
R6574 VSS.n998 VSS.n997 0.00170947
R6575 VSS.n997 VSS.n996 0.00170947
R6576 VSS.n995 VSS.n792 0.00170947
R6577 VSS.n792 VSS.n791 0.00170947
R6578 VSS.n795 VSS.n794 0.00170947
R6579 VSS.n794 VSS.n793 0.00170947
R6580 VSS.n991 VSS.n798 0.00170947
R6581 VSS.n798 VSS.n797 0.00170947
R6582 VSS.n990 VSS.n989 0.00170947
R6583 VSS.n989 VSS.n988 0.00170947
R6584 VSS.n801 VSS.n800 0.00170947
R6585 VSS.n800 VSS.n799 0.00170947
R6586 VSS.n984 VSS.n983 0.00170947
R6587 VSS.n983 VSS.n982 0.00170947
R6588 VSS.n981 VSS.n805 0.00170947
R6589 VSS.n805 VSS.n804 0.00170947
R6590 VSS.n808 VSS.n807 0.00170947
R6591 VSS.n807 VSS.n806 0.00170947
R6592 VSS.n977 VSS.n976 0.00170947
R6593 VSS.n976 VSS.n975 0.00170947
R6594 VSS.n966 VSS.n965 0.00170947
R6595 VSS.n965 VSS.n964 0.00170947
R6596 VSS.n963 VSS.n814 0.00170947
R6597 VSS.n814 VSS.n813 0.00170947
R6598 VSS.n817 VSS.n816 0.00170947
R6599 VSS.n816 VSS.n815 0.00170947
R6600 VSS.n959 VSS.n821 0.00170947
R6601 VSS.n821 VSS.n820 0.00170947
R6602 VSS.n958 VSS.n957 0.00170947
R6603 VSS.n957 VSS.n956 0.00170947
R6604 VSS.n824 VSS.n823 0.00170947
R6605 VSS.n823 VSS.n822 0.00170947
R6606 VSS.n952 VSS.n951 0.00170947
R6607 VSS.n951 VSS.n950 0.00170947
R6608 VSS.n949 VSS.n827 0.00170947
R6609 VSS.n827 VSS.n826 0.00170947
R6610 VSS.n830 VSS.n829 0.00170947
R6611 VSS.n829 VSS.n828 0.00170947
R6612 VSS.n945 VSS.n834 0.00170947
R6613 VSS.n834 VSS.n833 0.00170947
R6614 VSS.n944 VSS.n943 0.00170947
R6615 VSS.n943 VSS.n942 0.00170947
R6616 VSS.n837 VSS.n836 0.00170947
R6617 VSS.n836 VSS.n835 0.00170947
R6618 VSS.n938 VSS.n937 0.00170947
R6619 VSS.n937 VSS.n936 0.00170947
R6620 VSS.n935 VSS.n840 0.00170947
R6621 VSS.n840 VSS.n839 0.00170947
R6622 VSS.n843 VSS.n842 0.00170947
R6623 VSS.n842 VSS.n841 0.00170947
R6624 VSS.n931 VSS.n847 0.00170947
R6625 VSS.n847 VSS.n846 0.00170947
R6626 VSS.n930 VSS.n929 0.00170947
R6627 VSS.n929 VSS.n928 0.00170947
R6628 VSS.n925 VSS.n849 0.00170947
R6629 VSS.n849 VSS.n848 0.00170947
R6630 VSS.n924 VSS.n923 0.00170947
R6631 VSS.n923 VSS.n922 0.00170947
R6632 VSS.n852 VSS.n851 0.00170947
R6633 VSS.n851 VSS.n850 0.00170947
R6634 VSS.n918 VSS.n917 0.00170947
R6635 VSS.n917 VSS.n916 0.00170947
R6636 VSS.n915 VSS.n856 0.00170947
R6637 VSS.n856 VSS.n855 0.00170947
R6638 VSS.n859 VSS.n858 0.00170947
R6639 VSS.n858 VSS.n857 0.00170947
R6640 VSS.n911 VSS.n910 0.00170947
R6641 VSS.n910 VSS.n909 0.00170947
R6642 VSS.n900 VSS.n899 0.00170947
R6643 VSS.n899 VSS.n898 0.00170947
R6644 VSS.n897 VSS.n864 0.00170947
R6645 VSS.n864 VSS.n863 0.00170947
R6646 VSS.n867 VSS.n866 0.00170947
R6647 VSS.n866 VSS.n865 0.00170947
R6648 VSS.n893 VSS.n871 0.00170947
R6649 VSS.n871 VSS.n870 0.00170947
R6650 VSS.n892 VSS.n891 0.00170947
R6651 VSS.n891 VSS.n890 0.00170947
R6652 VSS.n887 VSS.n886 0.00170947
R6653 VSS.n886 VSS.n885 0.00170947
R6654 VSS.n876 VSS.n875 0.00170947
R6655 VSS.n875 VSS.n874 0.00170947
R6656 VSS.n377 VSS.n376 0.00118117
R6657 VSS.n103 VSS.n96 0.00118117
R6658 VSS.n107 VSS.n104 0.00118117
R6659 VSS.n111 VSS.n110 0.00118117
R6660 VSS.n112 VSS.n92 0.00118117
R6661 VSS.n116 VSS.n113 0.00118117
R6662 VSS.n120 VSS.n119 0.00118117
R6663 VSS.n121 VSS.n87 0.00118117
R6664 VSS.n125 VSS.n122 0.00118117
R6665 VSS.n129 VSS.n128 0.00118117
R6666 VSS.n130 VSS.n83 0.00118117
R6667 VSS.n134 VSS.n131 0.00118117
R6668 VSS.n138 VSS.n137 0.00118117
R6669 VSS.n139 VSS.n78 0.00118117
R6670 VSS.n143 VSS.n140 0.00118117
R6671 VSS.n147 VSS.n146 0.00118117
R6672 VSS.n148 VSS.n74 0.00118117
R6673 VSS.n152 VSS.n149 0.00118117
R6674 VSS.n156 VSS.n155 0.00118117
R6675 VSS.n157 VSS.n69 0.00118117
R6676 VSS.n161 VSS.n158 0.00118117
R6677 VSS.n165 VSS.n164 0.00118117
R6678 VSS.n166 VSS.n65 0.00118117
R6679 VSS.n170 VSS.n167 0.00118117
R6680 VSS.n174 VSS.n173 0.00118117
R6681 VSS.n175 VSS.n60 0.00118117
R6682 VSS.n179 VSS.n176 0.00118117
R6683 VSS.n183 VSS.n182 0.00118117
R6684 VSS.n184 VSS.n56 0.00118117
R6685 VSS.n188 VSS.n185 0.00118117
R6686 VSS.n192 VSS.n191 0.00118117
R6687 VSS.n193 VSS.n51 0.00118117
R6688 VSS.n197 VSS.n194 0.00118117
R6689 VSS.n201 VSS.n200 0.00118117
R6690 VSS.n202 VSS.n47 0.00118117
R6691 VSS.n206 VSS.n203 0.00118117
R6692 VSS.n210 VSS.n209 0.00118117
R6693 VSS.n211 VSS.n42 0.00118117
R6694 VSS.n215 VSS.n212 0.00118117
R6695 VSS.n219 VSS.n218 0.00118117
R6696 VSS.n220 VSS.n38 0.00118117
R6697 VSS.n224 VSS.n221 0.00118117
R6698 VSS.n228 VSS.n227 0.00118117
R6699 VSS.n229 VSS.n33 0.00118117
R6700 VSS.n233 VSS.n230 0.00118117
R6701 VSS.n237 VSS.n236 0.00118117
R6702 VSS.n238 VSS.n29 0.00118117
R6703 VSS.n242 VSS.n239 0.00118117
R6704 VSS.n246 VSS.n245 0.00118117
R6705 VSS.n247 VSS.n24 0.00118117
R6706 VSS.n251 VSS.n248 0.00118117
R6707 VSS.n255 VSS.n254 0.00118117
R6708 VSS.n256 VSS.n20 0.00118117
R6709 VSS.n260 VSS.n257 0.00118117
R6710 VSS.n264 VSS.n263 0.00118117
R6711 VSS.n265 VSS.n15 0.00118117
R6712 VSS.n269 VSS.n266 0.00118117
R6713 VSS.n273 VSS.n272 0.00118117
R6714 VSS.n274 VSS.n11 0.00118117
R6715 VSS.n278 VSS.n275 0.00118117
R6716 VSS.n282 VSS.n281 0.00118117
R6717 VSS.n283 VSS.n6 0.00118117
R6718 VSS.n287 VSS.n284 0.00118117
R6719 VSS.n291 VSS.n290 0.00118117
R6720 VSS.n597 VSS.n596 0.00118117
R6721 VSS.n102 VSS.n101 0.00118117
R6722 VSS.n390 VSS.n389 0.00118117
R6723 VSS.n386 VSS.n385 0.00118117
R6724 VSS.n381 VSS.n378 0.00118117
R6725 VSS.n394 VSS.n391 0.00118117
R6726 VSS.n406 VSS.n405 0.00118117
R6727 VSS.n404 VSS.n401 0.00118117
R6728 VSS.n400 VSS.n372 0.00118117
R6729 VSS.n399 VSS.n398 0.00118117
R6730 VSS.n410 VSS.n407 0.00118117
R6731 VSS.n595 VSS.n3 0.00118117
R6732 VSS.n594 VSS.n593 0.00118117
R6733 VSS.n590 VSS.n587 0.00118117
R6734 VSS.n586 VSS.n294 0.00118117
R6735 VSS.n585 VSS.n584 0.00118117
R6736 VSS.n581 VSS.n578 0.00118117
R6737 VSS.n577 VSS.n299 0.00118117
R6738 VSS.n576 VSS.n575 0.00118117
R6739 VSS.n572 VSS.n569 0.00118117
R6740 VSS.n568 VSS.n303 0.00118117
R6741 VSS.n567 VSS.n566 0.00118117
R6742 VSS.n563 VSS.n560 0.00118117
R6743 VSS.n559 VSS.n308 0.00118117
R6744 VSS.n558 VSS.n557 0.00118117
R6745 VSS.n554 VSS.n551 0.00118117
R6746 VSS.n550 VSS.n312 0.00118117
R6747 VSS.n549 VSS.n548 0.00118117
R6748 VSS.n545 VSS.n542 0.00118117
R6749 VSS.n541 VSS.n317 0.00118117
R6750 VSS.n540 VSS.n539 0.00118117
R6751 VSS.n534 VSS.n533 0.00118117
R6752 VSS.n532 VSS.n321 0.00118117
R6753 VSS.n531 VSS.n530 0.00118117
R6754 VSS.n527 VSS.n524 0.00118117
R6755 VSS.n523 VSS.n326 0.00118117
R6756 VSS.n522 VSS.n521 0.00118117
R6757 VSS.n518 VSS.n515 0.00118117
R6758 VSS.n514 VSS.n330 0.00118117
R6759 VSS.n513 VSS.n512 0.00118117
R6760 VSS.n509 VSS.n506 0.00118117
R6761 VSS.n505 VSS.n335 0.00118117
R6762 VSS.n504 VSS.n503 0.00118117
R6763 VSS.n500 VSS.n499 0.00118117
R6764 VSS.n495 VSS.n492 0.00118117
R6765 VSS.n491 VSS.n490 0.00118117
R6766 VSS.n487 VSS.n484 0.00118117
R6767 VSS.n483 VSS.n339 0.00118117
R6768 VSS.n482 VSS.n481 0.00118117
R6769 VSS.n478 VSS.n475 0.00118117
R6770 VSS.n474 VSS.n344 0.00118117
R6771 VSS.n473 VSS.n472 0.00118117
R6772 VSS.n469 VSS.n466 0.00118117
R6773 VSS.n465 VSS.n348 0.00118117
R6774 VSS.n464 VSS.n463 0.00118117
R6775 VSS.n460 VSS.n457 0.00118117
R6776 VSS.n456 VSS.n353 0.00118117
R6777 VSS.n455 VSS.n454 0.00118117
R6778 VSS.n451 VSS.n448 0.00118117
R6779 VSS.n447 VSS.n357 0.00118117
R6780 VSS.n446 VSS.n445 0.00118117
R6781 VSS.n441 VSS.n438 0.00118117
R6782 VSS.n437 VSS.n436 0.00118117
R6783 VSS.n433 VSS.n430 0.00118117
R6784 VSS.n429 VSS.n361 0.00118117
R6785 VSS.n428 VSS.n427 0.00118117
R6786 VSS.n424 VSS.n421 0.00118117
R6787 VSS.n420 VSS.n366 0.00118117
R6788 VSS.n419 VSS.n418 0.00118117
R6789 VSS.n415 VSS.n414 0.00118117
R6790 VSS.n604 VSS.n603 0.00118117
R6791 VSS.n608 VSS.n607 0.00118117
R6792 VSS.n1201 VSS.n1200 0.00118117
R6793 VSS.n1199 VSS.n1196 0.00118117
R6794 VSS.n1195 VSS.n614 0.00118117
R6795 VSS.n1194 VSS.n1193 0.00118117
R6796 VSS.n1190 VSS.n1189 0.00118117
R6797 VSS.n1188 VSS.n620 0.00118117
R6798 VSS.n1187 VSS.n1186 0.00118117
R6799 VSS.n1185 VSS.n1182 0.00118117
R6800 VSS.n1181 VSS.n627 0.00118117
R6801 VSS.n1180 VSS.n1179 0.00118117
R6802 VSS.n1176 VSS.n1175 0.00118117
R6803 VSS.n1174 VSS.n633 0.00118117
R6804 VSS.n1173 VSS.n1172 0.00118117
R6805 VSS.n1171 VSS.n1168 0.00118117
R6806 VSS.n1167 VSS.n640 0.00118117
R6807 VSS.n1166 VSS.n1165 0.00118117
R6808 VSS.n1162 VSS.n1161 0.00118117
R6809 VSS.n1160 VSS.n646 0.00118117
R6810 VSS.n1159 VSS.n1158 0.00118117
R6811 VSS.n1157 VSS.n1154 0.00118117
R6812 VSS.n1153 VSS.n653 0.00118117
R6813 VSS.n1152 VSS.n1151 0.00118117
R6814 VSS.n1148 VSS.n1147 0.00118117
R6815 VSS.n1146 VSS.n659 0.00118117
R6816 VSS.n1145 VSS.n1144 0.00118117
R6817 VSS.n1143 VSS.n1140 0.00118117
R6818 VSS.n1139 VSS.n666 0.00118117
R6819 VSS.n1138 VSS.n1137 0.00118117
R6820 VSS.n1134 VSS.n1133 0.00118117
R6821 VSS.n1132 VSS.n672 0.00118117
R6822 VSS.n1131 VSS.n1130 0.00118117
R6823 VSS.n1129 VSS.n1126 0.00118117
R6824 VSS.n1125 VSS.n679 0.00118117
R6825 VSS.n1124 VSS.n1123 0.00118117
R6826 VSS.n1120 VSS.n1119 0.00118117
R6827 VSS.n1118 VSS.n685 0.00118117
R6828 VSS.n1117 VSS.n1116 0.00118117
R6829 VSS.n1115 VSS.n1112 0.00118117
R6830 VSS.n1111 VSS.n692 0.00118117
R6831 VSS.n1110 VSS.n1109 0.00118117
R6832 VSS.n1106 VSS.n1105 0.00118117
R6833 VSS.n1104 VSS.n698 0.00118117
R6834 VSS.n1103 VSS.n1102 0.00118117
R6835 VSS.n1101 VSS.n1098 0.00118117
R6836 VSS.n1097 VSS.n705 0.00118117
R6837 VSS.n1096 VSS.n1095 0.00118117
R6838 VSS.n1092 VSS.n1091 0.00118117
R6839 VSS.n1090 VSS.n711 0.00118117
R6840 VSS.n1089 VSS.n1088 0.00118117
R6841 VSS.n1087 VSS.n1084 0.00118117
R6842 VSS.n1083 VSS.n718 0.00118117
R6843 VSS.n1082 VSS.n1081 0.00118117
R6844 VSS.n1078 VSS.n1077 0.00118117
R6845 VSS.n1076 VSS.n724 0.00118117
R6846 VSS.n1075 VSS.n1074 0.00118117
R6847 VSS.n1073 VSS.n1070 0.00118117
R6848 VSS.n1069 VSS.n731 0.00118117
R6849 VSS.n1068 VSS.n1067 0.00118117
R6850 VSS.n1064 VSS.n1063 0.00118117
R6851 VSS.n1062 VSS.n737 0.00118117
R6852 VSS.n1061 VSS.n1060 0.00118117
R6853 VSS.n1059 VSS.n1056 0.00118117
R6854 VSS.n1055 VSS.n1054 0.00118117
R6855 VSS.n1053 VSS.n1049 0.00118117
R6856 VSS.n1048 VSS.n1047 0.00118117
R6857 VSS.n1046 VSS.n1043 0.00118117
R6858 VSS.n1042 VSS.n749 0.00118117
R6859 VSS.n1041 VSS.n1040 0.00118117
R6860 VSS.n1037 VSS.n1036 0.00118117
R6861 VSS.n1035 VSS.n756 0.00118117
R6862 VSS.n1034 VSS.n1033 0.00118117
R6863 VSS.n1032 VSS.n1029 0.00118117
R6864 VSS.n1028 VSS.n762 0.00118117
R6865 VSS.n1027 VSS.n1026 0.00118117
R6866 VSS.n1023 VSS.n1022 0.00118117
R6867 VSS.n1021 VSS.n769 0.00118117
R6868 VSS.n1020 VSS.n1019 0.00118117
R6869 VSS.n1018 VSS.n1015 0.00118117
R6870 VSS.n1014 VSS.n775 0.00118117
R6871 VSS.n1013 VSS.n1012 0.00118117
R6872 VSS.n1009 VSS.n1008 0.00118117
R6873 VSS.n1007 VSS.n782 0.00118117
R6874 VSS.n1006 VSS.n1005 0.00118117
R6875 VSS.n1004 VSS.n1001 0.00118117
R6876 VSS.n1000 VSS.n788 0.00118117
R6877 VSS.n999 VSS.n998 0.00118117
R6878 VSS.n995 VSS.n994 0.00118117
R6879 VSS.n993 VSS.n795 0.00118117
R6880 VSS.n992 VSS.n991 0.00118117
R6881 VSS.n990 VSS.n987 0.00118117
R6882 VSS.n986 VSS.n801 0.00118117
R6883 VSS.n985 VSS.n984 0.00118117
R6884 VSS.n981 VSS.n980 0.00118117
R6885 VSS.n979 VSS.n808 0.00118117
R6886 VSS.n978 VSS.n977 0.00118117
R6887 VSS.n974 VSS.n973 0.00118117
R6888 VSS.n969 VSS.n968 0.00118117
R6889 VSS.n967 VSS.n966 0.00118117
R6890 VSS.n963 VSS.n962 0.00118117
R6891 VSS.n961 VSS.n817 0.00118117
R6892 VSS.n960 VSS.n959 0.00118117
R6893 VSS.n958 VSS.n955 0.00118117
R6894 VSS.n954 VSS.n824 0.00118117
R6895 VSS.n953 VSS.n952 0.00118117
R6896 VSS.n949 VSS.n948 0.00118117
R6897 VSS.n947 VSS.n830 0.00118117
R6898 VSS.n946 VSS.n945 0.00118117
R6899 VSS.n944 VSS.n941 0.00118117
R6900 VSS.n940 VSS.n837 0.00118117
R6901 VSS.n939 VSS.n938 0.00118117
R6902 VSS.n935 VSS.n934 0.00118117
R6903 VSS.n933 VSS.n843 0.00118117
R6904 VSS.n932 VSS.n931 0.00118117
R6905 VSS.n930 VSS.n927 0.00118117
R6906 VSS.n926 VSS.n925 0.00118117
R6907 VSS.n924 VSS.n921 0.00118117
R6908 VSS.n920 VSS.n852 0.00118117
R6909 VSS.n919 VSS.n918 0.00118117
R6910 VSS.n915 VSS.n914 0.00118117
R6911 VSS.n913 VSS.n859 0.00118117
R6912 VSS.n912 VSS.n911 0.00118117
R6913 VSS.n908 VSS.n907 0.00118117
R6914 VSS.n903 VSS.n902 0.00118117
R6915 VSS.n901 VSS.n900 0.00118117
R6916 VSS.n897 VSS.n896 0.00118117
R6917 VSS.n895 VSS.n867 0.00118117
R6918 VSS.n894 VSS.n893 0.00118117
R6919 VSS.n892 VSS.n889 0.00118117
R6920 VSS.n888 VSS.n887 0.00118117
R6921 VSS.n884 VSS.n883 0.00118117
R6922 VSS.n879 VSS.n878 0.00118117
R6923 VSS.n877 VSS.n876 0.00118117
R6924 db<6>.n1 db<6>.n0 88.1376
R6925 db<6>.n2 db<6>.n1 88.1376
R6926 db<6>.n3 db<6>.n2 88.1376
R6927 db<6>.n4 db<6>.n3 88.1376
R6928 db<6>.n5 db<6>.n4 88.1376
R6929 db<6>.n6 db<6>.n5 88.1376
R6930 db<6>.n7 db<6>.n6 88.1376
R6931 db<6>.n8 db<6>.n7 88.1376
R6932 db<6>.n9 db<6>.n8 88.1376
R6933 db<6>.n10 db<6>.n9 88.1376
R6934 db<6>.n11 db<6>.n10 88.1376
R6935 db<6>.n12 db<6>.n11 88.1376
R6936 db<6>.n13 db<6>.n12 88.1376
R6937 db<6>.n14 db<6>.n13 88.1376
R6938 db<6>.n15 db<6>.n14 88.1376
R6939 db<6>.n16 db<6>.n15 88.1376
R6940 db<6>.n17 db<6>.n16 88.1376
R6941 db<6>.n18 db<6>.n17 88.1376
R6942 db<6>.n19 db<6>.n18 88.1376
R6943 db<6>.n20 db<6>.n19 88.1376
R6944 db<6>.n21 db<6>.n20 88.1376
R6945 db<6>.n22 db<6>.n21 88.1376
R6946 db<6>.n23 db<6>.n22 88.1376
R6947 db<6>.n24 db<6>.n23 88.1376
R6948 db<6>.n25 db<6>.n24 88.1376
R6949 db<6>.n26 db<6>.n25 88.1376
R6950 db<6>.n27 db<6>.n26 88.1376
R6951 db<6>.n28 db<6>.n27 88.1376
R6952 db<6>.n29 db<6>.n28 88.1376
R6953 db<6>.n30 db<6>.n29 88.1376
R6954 db<6>.n31 db<6>.n30 88.1376
R6955 db<6>.n32 db<6>.n31 88.1376
R6956 db<6>.n33 db<6>.n32 88.1376
R6957 db<6>.n34 db<6>.n33 88.1376
R6958 db<6>.n35 db<6>.n34 88.1376
R6959 db<6>.n36 db<6>.n35 88.1376
R6960 db<6>.n37 db<6>.n36 88.1376
R6961 db<6>.n38 db<6>.n37 88.1376
R6962 db<6>.n39 db<6>.n38 88.1376
R6963 db<6>.n40 db<6>.n39 88.1376
R6964 db<6>.n41 db<6>.n40 88.1376
R6965 db<6>.n42 db<6>.n41 88.1376
R6966 db<6>.n43 db<6>.n42 88.1376
R6967 db<6>.n44 db<6>.n43 88.1376
R6968 db<6>.n45 db<6>.n44 88.1376
R6969 db<6>.n46 db<6>.n45 88.1376
R6970 db<6>.n47 db<6>.n46 88.1376
R6971 db<6>.n48 db<6>.n47 88.1376
R6972 db<6>.n49 db<6>.n48 88.1376
R6973 db<6>.n50 db<6>.n49 88.1376
R6974 db<6>.n51 db<6>.n50 88.1376
R6975 db<6>.n52 db<6>.n51 88.1376
R6976 db<6>.n53 db<6>.n52 88.1376
R6977 db<6>.n54 db<6>.n53 88.1376
R6978 db<6>.n55 db<6>.n54 88.1376
R6979 db<6>.n56 db<6>.n55 88.1376
R6980 db<6>.n57 db<6>.n56 88.1376
R6981 db<6>.n58 db<6>.n57 88.1376
R6982 db<6>.n59 db<6>.n58 88.1376
R6983 db<6>.n60 db<6>.n59 88.1376
R6984 db<6>.n61 db<6>.n60 88.1376
R6985 db<6>.n62 db<6>.n61 88.1376
R6986 db<6>.n63 db<6>.n62 88.1376
R6987 db<6>.n0 db<6>.t14 69.5462
R6988 db<6>.n1 db<6>.t96 69.5462
R6989 db<6>.n2 db<6>.t81 69.5462
R6990 db<6>.n3 db<6>.t66 69.5462
R6991 db<6>.n4 db<6>.t105 69.5462
R6992 db<6>.n5 db<6>.t55 69.5462
R6993 db<6>.n6 db<6>.t9 69.5462
R6994 db<6>.n7 db<6>.t26 69.5462
R6995 db<6>.n8 db<6>.t110 69.5462
R6996 db<6>.n9 db<6>.t58 69.5462
R6997 db<6>.n10 db<6>.t40 69.5462
R6998 db<6>.n11 db<6>.t126 69.5462
R6999 db<6>.n12 db<6>.t67 69.5462
R7000 db<6>.n13 db<6>.t18 69.5462
R7001 db<6>.n14 db<6>.t4 69.5462
R7002 db<6>.n15 db<6>.t85 69.5462
R7003 db<6>.n16 db<6>.t34 69.5462
R7004 db<6>.n17 db<6>.t21 69.5462
R7005 db<6>.n18 db<6>.t7 69.5462
R7006 db<6>.n19 db<6>.t87 69.5462
R7007 db<6>.n20 db<6>.t127 69.5462
R7008 db<6>.n21 db<6>.t112 69.5462
R7009 db<6>.n22 db<6>.t95 69.5462
R7010 db<6>.n23 db<6>.t44 69.5462
R7011 db<6>.n24 db<6>.t1 69.5462
R7012 db<6>.n25 db<6>.t115 69.5462
R7013 db<6>.n26 db<6>.t65 69.5462
R7014 db<6>.n27 db<6>.t47 69.5462
R7015 db<6>.n28 db<6>.t121 69.5462
R7016 db<6>.n29 db<6>.t70 69.5462
R7017 db<6>.n30 db<6>.t25 69.5462
R7018 db<6>.n31 db<6>.t109 69.5462
R7019 db<6>.n32 db<6>.t125 69.5462
R7020 db<6>.n33 db<6>.t73 69.5462
R7021 db<6>.n34 db<6>.t27 69.5462
R7022 db<6>.n35 db<6>.t99 69.5462
R7023 db<6>.n36 db<6>.t45 69.5462
R7024 db<6>.n37 db<6>.t32 69.5462
R7025 db<6>.n38 db<6>.t117 69.5462
R7026 db<6>.n39 db<6>.t102 69.5462
R7027 db<6>.n40 db<6>.t50 69.5462
R7028 db<6>.n41 db<6>.t6 69.5462
R7029 db<6>.n42 db<6>.t119 69.5462
R7030 db<6>.n43 db<6>.t59 69.5462
R7031 db<6>.n44 db<6>.t12 69.5462
R7032 db<6>.n45 db<6>.t93 69.5462
R7033 db<6>.n46 db<6>.t77 69.5462
R7034 db<6>.n47 db<6>.t63 69.5462
R7035 db<6>.n48 db<6>.t15 69.5462
R7036 db<6>.n49 db<6>.t98 69.5462
R7037 db<6>.n50 db<6>.t82 69.5462
R7038 db<6>.n51 db<6>.t118 69.5462
R7039 db<6>.n52 db<6>.t106 69.5462
R7040 db<6>.n53 db<6>.t88 69.5462
R7041 db<6>.n54 db<6>.t38 69.5462
R7042 db<6>.n55 db<6>.t123 69.5462
R7043 db<6>.n56 db<6>.t72 69.5462
R7044 db<6>.n57 db<6>.t91 69.5462
R7045 db<6>.n58 db<6>.t41 69.5462
R7046 db<6>.n59 db<6>.t97 69.5462
R7047 db<6>.n60 db<6>.t79 69.5462
R7048 db<6>.n61 db<6>.t30 69.5462
R7049 db<6>.n62 db<6>.t19 69.5462
R7050 db<6>.n63 db<6>.t101 69.5462
R7051 db<6>.n0 db<6>.t103 59.9062
R7052 db<6>.n1 db<6>.t51 59.9062
R7053 db<6>.n2 db<6>.t37 59.9062
R7054 db<6>.n3 db<6>.t23 59.9062
R7055 db<6>.n4 db<6>.t60 59.9062
R7056 db<6>.n5 db<6>.t13 59.9062
R7057 db<6>.n6 db<6>.t94 59.9062
R7058 db<6>.n7 db<6>.t114 59.9062
R7059 db<6>.n8 db<6>.t64 59.9062
R7060 db<6>.n9 db<6>.t16 59.9062
R7061 db<6>.n10 db<6>.t2 59.9062
R7062 db<6>.n11 db<6>.t83 59.9062
R7063 db<6>.n12 db<6>.t24 59.9062
R7064 db<6>.n13 db<6>.t107 59.9062
R7065 db<6>.n14 db<6>.t89 59.9062
R7066 db<6>.n15 db<6>.t39 59.9062
R7067 db<6>.n16 db<6>.t124 59.9062
R7068 db<6>.n17 db<6>.t111 59.9062
R7069 db<6>.n18 db<6>.t92 59.9062
R7070 db<6>.n19 db<6>.t42 59.9062
R7071 db<6>.n20 db<6>.t84 59.9062
R7072 db<6>.n21 db<6>.t68 59.9062
R7073 db<6>.n22 db<6>.t49 59.9062
R7074 db<6>.n23 db<6>.t5 59.9062
R7075 db<6>.n24 db<6>.t86 59.9062
R7076 db<6>.n25 db<6>.t69 59.9062
R7077 db<6>.n26 db<6>.t22 59.9062
R7078 db<6>.n27 db<6>.t10 59.9062
R7079 db<6>.n28 db<6>.t76 59.9062
R7080 db<6>.n29 db<6>.t28 59.9062
R7081 db<6>.n30 db<6>.t113 59.9062
R7082 db<6>.n31 db<6>.t62 59.9062
R7083 db<6>.n32 db<6>.t80 59.9062
R7084 db<6>.n33 db<6>.t31 59.9062
R7085 db<6>.n34 db<6>.t116 59.9062
R7086 db<6>.n35 db<6>.t54 59.9062
R7087 db<6>.n36 db<6>.t8 59.9062
R7088 db<6>.n37 db<6>.t122 59.9062
R7089 db<6>.n38 db<6>.t71 59.9062
R7090 db<6>.n39 db<6>.t57 59.9062
R7091 db<6>.n40 db<6>.t11 59.9062
R7092 db<6>.n41 db<6>.t90 59.9062
R7093 db<6>.n42 db<6>.t75 59.9062
R7094 db<6>.n43 db<6>.t17 59.9062
R7095 db<6>.n44 db<6>.t100 59.9062
R7096 db<6>.n45 db<6>.t48 59.9062
R7097 db<6>.n46 db<6>.t33 59.9062
R7098 db<6>.n47 db<6>.t20 59.9062
R7099 db<6>.n48 db<6>.t104 59.9062
R7100 db<6>.n49 db<6>.t53 59.9062
R7101 db<6>.n50 db<6>.t36 59.9062
R7102 db<6>.n51 db<6>.t74 59.9062
R7103 db<6>.n52 db<6>.t61 59.9062
R7104 db<6>.n53 db<6>.t43 59.9062
R7105 db<6>.n54 db<6>.t0 59.9062
R7106 db<6>.n55 db<6>.t78 59.9062
R7107 db<6>.n56 db<6>.t29 59.9062
R7108 db<6>.n57 db<6>.t46 59.9062
R7109 db<6>.n58 db<6>.t3 59.9062
R7110 db<6>.n59 db<6>.t52 59.9062
R7111 db<6>.n60 db<6>.t35 59.9062
R7112 db<6>.n61 db<6>.t120 59.9062
R7113 db<6>.n62 db<6>.t108 59.9062
R7114 db<6>.n63 db<6>.t56 59.9062
R7115 db<6> db<6>.n63 24.1005
R7116 hgu_cdac_8bit_array_2.drv<63:0>.n136 hgu_cdac_8bit_array_2.drv<63:0>.t101 41.4291
R7117 hgu_cdac_8bit_array_2.drv<63:0>.n136 hgu_cdac_8bit_array_2.drv<63:0>.t124 41.4291
R7118 hgu_cdac_8bit_array_2.drv<63:0>.n32 hgu_cdac_8bit_array_2.drv<63:0>.t74 41.4291
R7119 hgu_cdac_8bit_array_2.drv<63:0>.n32 hgu_cdac_8bit_array_2.drv<63:0>.t100 41.4291
R7120 hgu_cdac_8bit_array_2.drv<63:0>.n30 hgu_cdac_8bit_array_2.drv<63:0>.t107 41.4291
R7121 hgu_cdac_8bit_array_2.drv<63:0>.n30 hgu_cdac_8bit_array_2.drv<63:0>.t115 41.4291
R7122 hgu_cdac_8bit_array_2.drv<63:0>.n35 hgu_cdac_8bit_array_2.drv<63:0>.t94 41.4291
R7123 hgu_cdac_8bit_array_2.drv<63:0>.n35 hgu_cdac_8bit_array_2.drv<63:0>.t120 41.4291
R7124 hgu_cdac_8bit_array_2.drv<63:0>.n15 hgu_cdac_8bit_array_2.drv<63:0>.t76 41.4291
R7125 hgu_cdac_8bit_array_2.drv<63:0>.n15 hgu_cdac_8bit_array_2.drv<63:0>.t68 41.4291
R7126 hgu_cdac_8bit_array_2.drv<63:0>.n18 hgu_cdac_8bit_array_2.drv<63:0>.t91 41.4291
R7127 hgu_cdac_8bit_array_2.drv<63:0>.n18 hgu_cdac_8bit_array_2.drv<63:0>.t119 41.4291
R7128 hgu_cdac_8bit_array_2.drv<63:0>.n4 hgu_cdac_8bit_array_2.drv<63:0>.t126 41.4291
R7129 hgu_cdac_8bit_array_2.drv<63:0>.n4 hgu_cdac_8bit_array_2.drv<63:0>.t82 41.4291
R7130 hgu_cdac_8bit_array_2.drv<63:0>.n7 hgu_cdac_8bit_array_2.drv<63:0>.t114 41.4291
R7131 hgu_cdac_8bit_array_2.drv<63:0>.n7 hgu_cdac_8bit_array_2.drv<63:0>.t72 41.4291
R7132 hgu_cdac_8bit_array_2.drv<63:0>.n9 hgu_cdac_8bit_array_2.drv<63:0>.t79 41.4291
R7133 hgu_cdac_8bit_array_2.drv<63:0>.n9 hgu_cdac_8bit_array_2.drv<63:0>.t106 41.4291
R7134 hgu_cdac_8bit_array_2.drv<63:0>.n115 hgu_cdac_8bit_array_2.drv<63:0>.t64 41.4291
R7135 hgu_cdac_8bit_array_2.drv<63:0>.n115 hgu_cdac_8bit_array_2.drv<63:0>.t70 41.4291
R7136 hgu_cdac_8bit_array_2.drv<63:0>.n118 hgu_cdac_8bit_array_2.drv<63:0>.t77 41.4291
R7137 hgu_cdac_8bit_array_2.drv<63:0>.n118 hgu_cdac_8bit_array_2.drv<63:0>.t105 41.4291
R7138 hgu_cdac_8bit_array_2.drv<63:0>.n130 hgu_cdac_8bit_array_2.drv<63:0>.t81 41.4291
R7139 hgu_cdac_8bit_array_2.drv<63:0>.n130 hgu_cdac_8bit_array_2.drv<63:0>.t90 41.4291
R7140 hgu_cdac_8bit_array_2.drv<63:0>.n272 hgu_cdac_8bit_array_2.drv<63:0>.t71 41.4291
R7141 hgu_cdac_8bit_array_2.drv<63:0>.n272 hgu_cdac_8bit_array_2.drv<63:0>.t96 41.4291
R7142 hgu_cdac_8bit_array_2.drv<63:0>.n260 hgu_cdac_8bit_array_2.drv<63:0>.t109 41.4291
R7143 hgu_cdac_8bit_array_2.drv<63:0>.n260 hgu_cdac_8bit_array_2.drv<63:0>.t66 41.4291
R7144 hgu_cdac_8bit_array_2.drv<63:0>.n257 hgu_cdac_8bit_array_2.drv<63:0>.t125 41.4291
R7145 hgu_cdac_8bit_array_2.drv<63:0>.n257 hgu_cdac_8bit_array_2.drv<63:0>.t99 41.4291
R7146 hgu_cdac_8bit_array_2.drv<63:0>.n245 hgu_cdac_8bit_array_2.drv<63:0>.t112 41.4291
R7147 hgu_cdac_8bit_array_2.drv<63:0>.n245 hgu_cdac_8bit_array_2.drv<63:0>.t103 41.4291
R7148 hgu_cdac_8bit_array_2.drv<63:0>.n242 hgu_cdac_8bit_array_2.drv<63:0>.t127 41.4291
R7149 hgu_cdac_8bit_array_2.drv<63:0>.n242 hgu_cdac_8bit_array_2.drv<63:0>.t84 41.4291
R7150 hgu_cdac_8bit_array_2.drv<63:0>.n229 hgu_cdac_8bit_array_2.drv<63:0>.t93 41.4291
R7151 hgu_cdac_8bit_array_2.drv<63:0>.n229 hgu_cdac_8bit_array_2.drv<63:0>.t104 41.4291
R7152 hgu_cdac_8bit_array_2.drv<63:0>.n227 hgu_cdac_8bit_array_2.drv<63:0>.t108 41.4291
R7153 hgu_cdac_8bit_array_2.drv<63:0>.n227 hgu_cdac_8bit_array_2.drv<63:0>.t87 41.4291
R7154 hgu_cdac_8bit_array_2.drv<63:0>.n224 hgu_cdac_8bit_array_2.drv<63:0>.t73 41.4291
R7155 hgu_cdac_8bit_array_2.drv<63:0>.n224 hgu_cdac_8bit_array_2.drv<63:0>.t98 41.4291
R7156 hgu_cdac_8bit_array_2.drv<63:0>.n212 hgu_cdac_8bit_array_2.drv<63:0>.t110 41.4291
R7157 hgu_cdac_8bit_array_2.drv<63:0>.n212 hgu_cdac_8bit_array_2.drv<63:0>.t117 41.4291
R7158 hgu_cdac_8bit_array_2.drv<63:0>.n209 hgu_cdac_8bit_array_2.drv<63:0>.t75 41.4291
R7159 hgu_cdac_8bit_array_2.drv<63:0>.n209 hgu_cdac_8bit_array_2.drv<63:0>.t102 41.4291
R7160 hgu_cdac_8bit_array_2.drv<63:0>.n197 hgu_cdac_8bit_array_2.drv<63:0>.t86 41.4291
R7161 hgu_cdac_8bit_array_2.drv<63:0>.n197 hgu_cdac_8bit_array_2.drv<63:0>.t118 41.4291
R7162 hgu_cdac_8bit_array_2.drv<63:0>.n191 hgu_cdac_8bit_array_2.drv<63:0>.t121 41.4291
R7163 hgu_cdac_8bit_array_2.drv<63:0>.n191 hgu_cdac_8bit_array_2.drv<63:0>.t78 41.4291
R7164 hgu_cdac_8bit_array_2.drv<63:0>.n193 hgu_cdac_8bit_array_2.drv<63:0>.t88 41.4291
R7165 hgu_cdac_8bit_array_2.drv<63:0>.n193 hgu_cdac_8bit_array_2.drv<63:0>.t95 41.4291
R7166 hgu_cdac_8bit_array_2.drv<63:0>.n179 hgu_cdac_8bit_array_2.drv<63:0>.t123 41.4291
R7167 hgu_cdac_8bit_array_2.drv<63:0>.n179 hgu_cdac_8bit_array_2.drv<63:0>.t65 41.4291
R7168 hgu_cdac_8bit_array_2.drv<63:0>.n164 hgu_cdac_8bit_array_2.drv<63:0>.t67 41.4291
R7169 hgu_cdac_8bit_array_2.drv<63:0>.n164 hgu_cdac_8bit_array_2.drv<63:0>.t97 41.4291
R7170 hgu_cdac_8bit_array_2.drv<63:0>.n167 hgu_cdac_8bit_array_2.drv<63:0>.t83 41.4291
R7171 hgu_cdac_8bit_array_2.drv<63:0>.n167 hgu_cdac_8bit_array_2.drv<63:0>.t111 41.4291
R7172 hgu_cdac_8bit_array_2.drv<63:0>.n161 hgu_cdac_8bit_array_2.drv<63:0>.t69 41.4291
R7173 hgu_cdac_8bit_array_2.drv<63:0>.n161 hgu_cdac_8bit_array_2.drv<63:0>.t92 41.4291
R7174 hgu_cdac_8bit_array_2.drv<63:0>.n150 hgu_cdac_8bit_array_2.drv<63:0>.t85 41.4291
R7175 hgu_cdac_8bit_array_2.drv<63:0>.n150 hgu_cdac_8bit_array_2.drv<63:0>.t113 41.4291
R7176 hgu_cdac_8bit_array_2.drv<63:0>.n148 hgu_cdac_8bit_array_2.drv<63:0>.t116 41.4291
R7177 hgu_cdac_8bit_array_2.drv<63:0>.n148 hgu_cdac_8bit_array_2.drv<63:0>.t122 41.4291
R7178 hgu_cdac_8bit_array_2.drv<63:0>.n134 hgu_cdac_8bit_array_2.drv<63:0>.t80 41.4291
R7179 hgu_cdac_8bit_array_2.drv<63:0>.n134 hgu_cdac_8bit_array_2.drv<63:0>.t89 41.4291
R7180 hgu_cdac_8bit_array_2.drv<63:0>.n132 hgu_cdac_8bit_array_2.drv<63:0>.t20 34.0065
R7181 hgu_cdac_8bit_array_2.drv<63:0>.n132 hgu_cdac_8bit_array_2.drv<63:0>.t43 34.0065
R7182 hgu_cdac_8bit_array_2.drv<63:0>.n31 hgu_cdac_8bit_array_2.drv<63:0>.t57 34.0065
R7183 hgu_cdac_8bit_array_2.drv<63:0>.n31 hgu_cdac_8bit_array_2.drv<63:0>.t19 34.0065
R7184 hgu_cdac_8bit_array_2.drv<63:0>.n29 hgu_cdac_8bit_array_2.drv<63:0>.t27 34.0065
R7185 hgu_cdac_8bit_array_2.drv<63:0>.n29 hgu_cdac_8bit_array_2.drv<63:0>.t34 34.0065
R7186 hgu_cdac_8bit_array_2.drv<63:0>.n34 hgu_cdac_8bit_array_2.drv<63:0>.t13 34.0065
R7187 hgu_cdac_8bit_array_2.drv<63:0>.n34 hgu_cdac_8bit_array_2.drv<63:0>.t39 34.0065
R7188 hgu_cdac_8bit_array_2.drv<63:0>.n14 hgu_cdac_8bit_array_2.drv<63:0>.t59 34.0065
R7189 hgu_cdac_8bit_array_2.drv<63:0>.n14 hgu_cdac_8bit_array_2.drv<63:0>.t51 34.0065
R7190 hgu_cdac_8bit_array_2.drv<63:0>.n17 hgu_cdac_8bit_array_2.drv<63:0>.t10 34.0065
R7191 hgu_cdac_8bit_array_2.drv<63:0>.n17 hgu_cdac_8bit_array_2.drv<63:0>.t38 34.0065
R7192 hgu_cdac_8bit_array_2.drv<63:0>.n3 hgu_cdac_8bit_array_2.drv<63:0>.t45 34.0065
R7193 hgu_cdac_8bit_array_2.drv<63:0>.n3 hgu_cdac_8bit_array_2.drv<63:0>.t1 34.0065
R7194 hgu_cdac_8bit_array_2.drv<63:0>.n6 hgu_cdac_8bit_array_2.drv<63:0>.t33 34.0065
R7195 hgu_cdac_8bit_array_2.drv<63:0>.n6 hgu_cdac_8bit_array_2.drv<63:0>.t55 34.0065
R7196 hgu_cdac_8bit_array_2.drv<63:0>.n8 hgu_cdac_8bit_array_2.drv<63:0>.t62 34.0065
R7197 hgu_cdac_8bit_array_2.drv<63:0>.n8 hgu_cdac_8bit_array_2.drv<63:0>.t25 34.0065
R7198 hgu_cdac_8bit_array_2.drv<63:0>.n114 hgu_cdac_8bit_array_2.drv<63:0>.t47 34.0065
R7199 hgu_cdac_8bit_array_2.drv<63:0>.n114 hgu_cdac_8bit_array_2.drv<63:0>.t53 34.0065
R7200 hgu_cdac_8bit_array_2.drv<63:0>.n117 hgu_cdac_8bit_array_2.drv<63:0>.t60 34.0065
R7201 hgu_cdac_8bit_array_2.drv<63:0>.n117 hgu_cdac_8bit_array_2.drv<63:0>.t24 34.0065
R7202 hgu_cdac_8bit_array_2.drv<63:0>.n129 hgu_cdac_8bit_array_2.drv<63:0>.t0 34.0065
R7203 hgu_cdac_8bit_array_2.drv<63:0>.n129 hgu_cdac_8bit_array_2.drv<63:0>.t9 34.0065
R7204 hgu_cdac_8bit_array_2.drv<63:0>.n271 hgu_cdac_8bit_array_2.drv<63:0>.t54 34.0065
R7205 hgu_cdac_8bit_array_2.drv<63:0>.n271 hgu_cdac_8bit_array_2.drv<63:0>.t15 34.0065
R7206 hgu_cdac_8bit_array_2.drv<63:0>.n259 hgu_cdac_8bit_array_2.drv<63:0>.t28 34.0065
R7207 hgu_cdac_8bit_array_2.drv<63:0>.n259 hgu_cdac_8bit_array_2.drv<63:0>.t49 34.0065
R7208 hgu_cdac_8bit_array_2.drv<63:0>.n256 hgu_cdac_8bit_array_2.drv<63:0>.t44 34.0065
R7209 hgu_cdac_8bit_array_2.drv<63:0>.n256 hgu_cdac_8bit_array_2.drv<63:0>.t18 34.0065
R7210 hgu_cdac_8bit_array_2.drv<63:0>.n244 hgu_cdac_8bit_array_2.drv<63:0>.t31 34.0065
R7211 hgu_cdac_8bit_array_2.drv<63:0>.n244 hgu_cdac_8bit_array_2.drv<63:0>.t22 34.0065
R7212 hgu_cdac_8bit_array_2.drv<63:0>.n241 hgu_cdac_8bit_array_2.drv<63:0>.t46 34.0065
R7213 hgu_cdac_8bit_array_2.drv<63:0>.n241 hgu_cdac_8bit_array_2.drv<63:0>.t3 34.0065
R7214 hgu_cdac_8bit_array_2.drv<63:0>.n228 hgu_cdac_8bit_array_2.drv<63:0>.t12 34.0065
R7215 hgu_cdac_8bit_array_2.drv<63:0>.n228 hgu_cdac_8bit_array_2.drv<63:0>.t23 34.0065
R7216 hgu_cdac_8bit_array_2.drv<63:0>.n226 hgu_cdac_8bit_array_2.drv<63:0>.t26 34.0065
R7217 hgu_cdac_8bit_array_2.drv<63:0>.n226 hgu_cdac_8bit_array_2.drv<63:0>.t6 34.0065
R7218 hgu_cdac_8bit_array_2.drv<63:0>.n223 hgu_cdac_8bit_array_2.drv<63:0>.t56 34.0065
R7219 hgu_cdac_8bit_array_2.drv<63:0>.n223 hgu_cdac_8bit_array_2.drv<63:0>.t17 34.0065
R7220 hgu_cdac_8bit_array_2.drv<63:0>.n211 hgu_cdac_8bit_array_2.drv<63:0>.t29 34.0065
R7221 hgu_cdac_8bit_array_2.drv<63:0>.n211 hgu_cdac_8bit_array_2.drv<63:0>.t36 34.0065
R7222 hgu_cdac_8bit_array_2.drv<63:0>.n208 hgu_cdac_8bit_array_2.drv<63:0>.t58 34.0065
R7223 hgu_cdac_8bit_array_2.drv<63:0>.n208 hgu_cdac_8bit_array_2.drv<63:0>.t21 34.0065
R7224 hgu_cdac_8bit_array_2.drv<63:0>.n196 hgu_cdac_8bit_array_2.drv<63:0>.t5 34.0065
R7225 hgu_cdac_8bit_array_2.drv<63:0>.n196 hgu_cdac_8bit_array_2.drv<63:0>.t37 34.0065
R7226 hgu_cdac_8bit_array_2.drv<63:0>.n190 hgu_cdac_8bit_array_2.drv<63:0>.t40 34.0065
R7227 hgu_cdac_8bit_array_2.drv<63:0>.n190 hgu_cdac_8bit_array_2.drv<63:0>.t61 34.0065
R7228 hgu_cdac_8bit_array_2.drv<63:0>.n192 hgu_cdac_8bit_array_2.drv<63:0>.t7 34.0065
R7229 hgu_cdac_8bit_array_2.drv<63:0>.n192 hgu_cdac_8bit_array_2.drv<63:0>.t14 34.0065
R7230 hgu_cdac_8bit_array_2.drv<63:0>.n178 hgu_cdac_8bit_array_2.drv<63:0>.t42 34.0065
R7231 hgu_cdac_8bit_array_2.drv<63:0>.n178 hgu_cdac_8bit_array_2.drv<63:0>.t48 34.0065
R7232 hgu_cdac_8bit_array_2.drv<63:0>.n163 hgu_cdac_8bit_array_2.drv<63:0>.t50 34.0065
R7233 hgu_cdac_8bit_array_2.drv<63:0>.n163 hgu_cdac_8bit_array_2.drv<63:0>.t16 34.0065
R7234 hgu_cdac_8bit_array_2.drv<63:0>.n166 hgu_cdac_8bit_array_2.drv<63:0>.t2 34.0065
R7235 hgu_cdac_8bit_array_2.drv<63:0>.n166 hgu_cdac_8bit_array_2.drv<63:0>.t30 34.0065
R7236 hgu_cdac_8bit_array_2.drv<63:0>.n160 hgu_cdac_8bit_array_2.drv<63:0>.t52 34.0065
R7237 hgu_cdac_8bit_array_2.drv<63:0>.n160 hgu_cdac_8bit_array_2.drv<63:0>.t11 34.0065
R7238 hgu_cdac_8bit_array_2.drv<63:0>.n149 hgu_cdac_8bit_array_2.drv<63:0>.t4 34.0065
R7239 hgu_cdac_8bit_array_2.drv<63:0>.n149 hgu_cdac_8bit_array_2.drv<63:0>.t32 34.0065
R7240 hgu_cdac_8bit_array_2.drv<63:0>.n147 hgu_cdac_8bit_array_2.drv<63:0>.t35 34.0065
R7241 hgu_cdac_8bit_array_2.drv<63:0>.n147 hgu_cdac_8bit_array_2.drv<63:0>.t41 34.0065
R7242 hgu_cdac_8bit_array_2.drv<63:0>.n133 hgu_cdac_8bit_array_2.drv<63:0>.t63 34.0065
R7243 hgu_cdac_8bit_array_2.drv<63:0>.n133 hgu_cdac_8bit_array_2.drv<63:0>.t8 34.0065
R7244 hgu_cdac_8bit_array_2.drv<63:0>.n189 hgu_cdac_8bit_array_2.drv<63:0>.n181 12.9862
R7245 hgu_cdac_8bit_array_2.drv<63:0>.n280 hgu_cdac_8bit_array_2.drv<63:0>.n1 12.5753
R7246 hgu_cdac_8bit_array_2.drv<63:0>.n128 hgu_cdac_8bit_array_2.drv<63:0>.n120 12.2311
R7247 hgu_cdac_8bit_array_2.drv<63:0>.n270 hgu_cdac_8bit_array_2.drv<63:0>.n262 11.7398
R7248 hgu_cdac_8bit_array_2.drv<63:0>.n255 hgu_cdac_8bit_array_2.drv<63:0>.n247 11.7383
R7249 hgu_cdac_8bit_array_2.drv<63:0>.n146 hgu_cdac_8bit_array_2.drv<63:0>.n138 11.7381
R7250 hgu_cdac_8bit_array_2.drv<63:0>.n159 hgu_cdac_8bit_array_2.drv<63:0>.n2 11.7381
R7251 hgu_cdac_8bit_array_2.drv<63:0>.n177 hgu_cdac_8bit_array_2.drv<63:0>.n169 11.7381
R7252 hgu_cdac_8bit_array_2.drv<63:0>.n207 hgu_cdac_8bit_array_2.drv<63:0>.n199 11.7381
R7253 hgu_cdac_8bit_array_2.drv<63:0>.n222 hgu_cdac_8bit_array_2.drv<63:0>.n214 11.7381
R7254 hgu_cdac_8bit_array_2.drv<63:0>.n240 hgu_cdac_8bit_array_2.drv<63:0>.n232 11.7381
R7255 hgu_cdac_8bit_array_2.drv<63:0>.n28 hgu_cdac_8bit_array_2.drv<63:0>.n20 11.7374
R7256 hgu_cdac_8bit_array_2.drv<63:0>.n45 hgu_cdac_8bit_array_2.drv<63:0>.n37 11.7374
R7257 hgu_cdac_8bit_array_2.drv<63:0>.n13 hgu_cdac_8bit_array_2.drv<63:0>.n12 11.7367
R7258 hgu_cdac_8bit_array_2.drv<63:0>.n33 hgu_cdac_8bit_array_2.drv<63:0>.n0 0.9906
R7259 hgu_cdac_8bit_array_2.drv<63:0>.n11 hgu_cdac_8bit_array_2.drv<63:0>.n10 0.9906
R7260 hgu_cdac_8bit_array_2.drv<63:0>.n231 hgu_cdac_8bit_array_2.drv<63:0>.n230 0.9906
R7261 hgu_cdac_8bit_array_2.drv<63:0>.n195 hgu_cdac_8bit_array_2.drv<63:0>.n194 0.9906
R7262 hgu_cdac_8bit_array_2.drv<63:0>.n168 hgu_cdac_8bit_array_2.drv<63:0>.n165 0.957397
R7263 hgu_cdac_8bit_array_2.drv<63:0>.n137 hgu_cdac_8bit_array_2.drv<63:0>.n135 0.957397
R7264 hgu_cdac_8bit_array_2.drv<63:0>.n2 hgu_cdac_8bit_array_2.drv<63:0>.n151 0.950931
R7265 hgu_cdac_8bit_array_2.drv<63:0>.n12 hgu_cdac_8bit_array_2.drv<63:0>.n5 0.843172
R7266 hgu_cdac_8bit_array_2.drv<63:0>.n199 hgu_cdac_8bit_array_2.drv<63:0>.n198 0.838862
R7267 hgu_cdac_8bit_array_2.drv<63:0>.n232 hgu_cdac_8bit_array_2.drv<63:0>.n225 0.778517
R7268 hgu_cdac_8bit_array_2.drv<63:0>.n37 hgu_cdac_8bit_array_2.drv<63:0>.n36 0.774207
R7269 hgu_cdac_8bit_array_2.drv<63:0>.n247 hgu_cdac_8bit_array_2.drv<63:0>.n246 0.744035
R7270 hgu_cdac_8bit_array_2.drv<63:0>.n120 hgu_cdac_8bit_array_2.drv<63:0>.n119 0.623345
R7271 hgu_cdac_8bit_array_2.drv<63:0>.n137 hgu_cdac_8bit_array_2.drv<63:0>.n132 0.561881
R7272 hgu_cdac_8bit_array_2.drv<63:0>.n36 hgu_cdac_8bit_array_2.drv<63:0>.n34 0.561881
R7273 hgu_cdac_8bit_array_2.drv<63:0>.n16 hgu_cdac_8bit_array_2.drv<63:0>.n14 0.561881
R7274 hgu_cdac_8bit_array_2.drv<63:0>.n19 hgu_cdac_8bit_array_2.drv<63:0>.n17 0.561881
R7275 hgu_cdac_8bit_array_2.drv<63:0>.n5 hgu_cdac_8bit_array_2.drv<63:0>.n3 0.561881
R7276 hgu_cdac_8bit_array_2.drv<63:0>.n10 hgu_cdac_8bit_array_2.drv<63:0>.n8 0.561881
R7277 hgu_cdac_8bit_array_2.drv<63:0>.n116 hgu_cdac_8bit_array_2.drv<63:0>.n114 0.561881
R7278 hgu_cdac_8bit_array_2.drv<63:0>.n119 hgu_cdac_8bit_array_2.drv<63:0>.n117 0.561881
R7279 hgu_cdac_8bit_array_2.drv<63:0>.n131 hgu_cdac_8bit_array_2.drv<63:0>.n129 0.561881
R7280 hgu_cdac_8bit_array_2.drv<63:0>.n261 hgu_cdac_8bit_array_2.drv<63:0>.n259 0.561881
R7281 hgu_cdac_8bit_array_2.drv<63:0>.n258 hgu_cdac_8bit_array_2.drv<63:0>.n256 0.561881
R7282 hgu_cdac_8bit_array_2.drv<63:0>.n246 hgu_cdac_8bit_array_2.drv<63:0>.n244 0.561881
R7283 hgu_cdac_8bit_array_2.drv<63:0>.n230 hgu_cdac_8bit_array_2.drv<63:0>.n228 0.561881
R7284 hgu_cdac_8bit_array_2.drv<63:0>.n225 hgu_cdac_8bit_array_2.drv<63:0>.n223 0.561881
R7285 hgu_cdac_8bit_array_2.drv<63:0>.n213 hgu_cdac_8bit_array_2.drv<63:0>.n211 0.561881
R7286 hgu_cdac_8bit_array_2.drv<63:0>.n210 hgu_cdac_8bit_array_2.drv<63:0>.n208 0.561881
R7287 hgu_cdac_8bit_array_2.drv<63:0>.n198 hgu_cdac_8bit_array_2.drv<63:0>.n196 0.561881
R7288 hgu_cdac_8bit_array_2.drv<63:0>.n194 hgu_cdac_8bit_array_2.drv<63:0>.n192 0.561881
R7289 hgu_cdac_8bit_array_2.drv<63:0>.n180 hgu_cdac_8bit_array_2.drv<63:0>.n178 0.561881
R7290 hgu_cdac_8bit_array_2.drv<63:0>.n165 hgu_cdac_8bit_array_2.drv<63:0>.n163 0.561881
R7291 hgu_cdac_8bit_array_2.drv<63:0>.n168 hgu_cdac_8bit_array_2.drv<63:0>.n166 0.561881
R7292 hgu_cdac_8bit_array_2.drv<63:0>.n162 hgu_cdac_8bit_array_2.drv<63:0>.n160 0.561881
R7293 hgu_cdac_8bit_array_2.drv<63:0>.n151 hgu_cdac_8bit_array_2.drv<63:0>.n149 0.561881
R7294 hgu_cdac_8bit_array_2.drv<63:0>.n135 hgu_cdac_8bit_array_2.drv<63:0>.n133 0.561881
R7295 hgu_cdac_8bit_array_2.drv<63:0>.n0 hgu_cdac_8bit_array_2.drv<63:0>.n31 0.558205
R7296 hgu_cdac_8bit_array_2.drv<63:0>.n1 hgu_cdac_8bit_array_2.drv<63:0>.n271 0.558205
R7297 hgu_cdac_8bit_array_2.drv<63:0>.n138 hgu_cdac_8bit_array_2.drv<63:0>.n131 0.550069
R7298 hgu_cdac_8bit_array_2.drv<63:0>.n169 hgu_cdac_8bit_array_2.drv<63:0>.n168 0.545759
R7299 hgu_cdac_8bit_array_2.drv<63:0>.n262 hgu_cdac_8bit_array_2.drv<63:0>.n258 0.480142
R7300 hgu_cdac_8bit_array_2.drv<63:0>.n20 hgu_cdac_8bit_array_2.drv<63:0>.n16 0.438
R7301 hgu_cdac_8bit_array_2.drv<63:0>.n214 hgu_cdac_8bit_array_2.drv<63:0>.n213 0.43369
R7302 hgu_cdac_8bit_array_2.drv<63:0>.n11 hgu_cdac_8bit_array_2.drv<63:0>.n6 0.381734
R7303 hgu_cdac_8bit_array_2.drv<63:0>.n33 hgu_cdac_8bit_array_2.drv<63:0>.n29 0.378057
R7304 hgu_cdac_8bit_array_2.drv<63:0>.n243 hgu_cdac_8bit_array_2.drv<63:0>.n241 0.378057
R7305 hgu_cdac_8bit_array_2.drv<63:0>.n231 hgu_cdac_8bit_array_2.drv<63:0>.n226 0.378057
R7306 hgu_cdac_8bit_array_2.drv<63:0>.n195 hgu_cdac_8bit_array_2.drv<63:0>.n190 0.378057
R7307 hgu_cdac_8bit_array_2.drv<63:0>.n2 hgu_cdac_8bit_array_2.drv<63:0>.n147 0.378057
R7308 hgu_cdac_8bit_array_2.drv<63:0>.n214 hgu_cdac_8bit_array_2.drv<63:0>.n210 0.373345
R7309 hgu_cdac_8bit_array_2.drv<63:0>.n20 hgu_cdac_8bit_array_2.drv<63:0>.n19 0.369034
R7310 hgu_cdac_8bit_array_2.drv<63:0>.n64 hgu_cdac_8bit_array_2.drv<63:0> 0.338468
R7311 hgu_cdac_8bit_array_2.drv<63:0>.n68 hgu_cdac_8bit_array_2.drv<63:0>.n63 0.330451
R7312 hgu_cdac_8bit_array_2.drv<63:0>.n77 hgu_cdac_8bit_array_2.drv<63:0>.n60 0.330451
R7313 hgu_cdac_8bit_array_2.drv<63:0>.n496 hgu_cdac_8bit_array_2.drv<63:0>.n287 0.330451
R7314 hgu_cdac_8bit_array_2.drv<63:0>.n487 hgu_cdac_8bit_array_2.drv<63:0>.n294 0.330451
R7315 hgu_cdac_8bit_array_2.drv<63:0>.n478 hgu_cdac_8bit_array_2.drv<63:0>.n301 0.330451
R7316 hgu_cdac_8bit_array_2.drv<63:0>.n469 hgu_cdac_8bit_array_2.drv<63:0>.n308 0.330451
R7317 hgu_cdac_8bit_array_2.drv<63:0>.n460 hgu_cdac_8bit_array_2.drv<63:0>.n315 0.330451
R7318 hgu_cdac_8bit_array_2.drv<63:0>.n451 hgu_cdac_8bit_array_2.drv<63:0>.n322 0.330451
R7319 hgu_cdac_8bit_array_2.drv<63:0>.n442 hgu_cdac_8bit_array_2.drv<63:0>.n329 0.330451
R7320 hgu_cdac_8bit_array_2.drv<63:0>.n433 hgu_cdac_8bit_array_2.drv<63:0>.n336 0.330451
R7321 hgu_cdac_8bit_array_2.drv<63:0>.n424 hgu_cdac_8bit_array_2.drv<63:0>.n343 0.330451
R7322 hgu_cdac_8bit_array_2.drv<63:0>.n415 hgu_cdac_8bit_array_2.drv<63:0>.n350 0.330451
R7323 hgu_cdac_8bit_array_2.drv<63:0>.n406 hgu_cdac_8bit_array_2.drv<63:0>.n357 0.330451
R7324 hgu_cdac_8bit_array_2.drv<63:0>.n397 hgu_cdac_8bit_array_2.drv<63:0>.n364 0.330451
R7325 hgu_cdac_8bit_array_2.drv<63:0>.n388 hgu_cdac_8bit_array_2.drv<63:0>.n371 0.330451
R7326 hgu_cdac_8bit_array_2.drv<63:0>.n379 hgu_cdac_8bit_array_2.drv<63:0>.n374 0.330451
R7327 hgu_cdac_8bit_array_2.drv<63:0>.n262 hgu_cdac_8bit_array_2.drv<63:0>.n261 0.324969
R7328 hgu_cdac_8bit_array_2.drv<63:0>.n376 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7329 hgu_cdac_8bit_array_2.drv<63:0>.n385 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7330 hgu_cdac_8bit_array_2.drv<63:0>.n394 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7331 hgu_cdac_8bit_array_2.drv<63:0>.n403 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7332 hgu_cdac_8bit_array_2.drv<63:0>.n412 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7333 hgu_cdac_8bit_array_2.drv<63:0>.n421 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7334 hgu_cdac_8bit_array_2.drv<63:0>.n430 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7335 hgu_cdac_8bit_array_2.drv<63:0>.n439 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7336 hgu_cdac_8bit_array_2.drv<63:0>.n448 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7337 hgu_cdac_8bit_array_2.drv<63:0>.n457 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7338 hgu_cdac_8bit_array_2.drv<63:0>.n466 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7339 hgu_cdac_8bit_array_2.drv<63:0>.n475 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7340 hgu_cdac_8bit_array_2.drv<63:0>.n484 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7341 hgu_cdac_8bit_array_2.drv<63:0>.n493 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7342 hgu_cdac_8bit_array_2.drv<63:0>.n502 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7343 hgu_cdac_8bit_array_2.drv<63:0>.n512 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7344 hgu_cdac_8bit_array_2.drv<63:0>.n521 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7345 hgu_cdac_8bit_array_2.drv<63:0>.n530 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7346 hgu_cdac_8bit_array_2.drv<63:0>.n539 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7347 hgu_cdac_8bit_array_2.drv<63:0>.n548 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7348 hgu_cdac_8bit_array_2.drv<63:0>.n557 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7349 hgu_cdac_8bit_array_2.drv<63:0>.n566 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7350 hgu_cdac_8bit_array_2.drv<63:0>.n575 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7351 hgu_cdac_8bit_array_2.drv<63:0>.n584 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7352 hgu_cdac_8bit_array_2.drv<63:0>.n593 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7353 hgu_cdac_8bit_array_2.drv<63:0>.n602 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7354 hgu_cdac_8bit_array_2.drv<63:0>.n107 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7355 hgu_cdac_8bit_array_2.drv<63:0>.n98 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7356 hgu_cdac_8bit_array_2.drv<63:0>.n89 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7357 hgu_cdac_8bit_array_2.drv<63:0>.n80 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7358 hgu_cdac_8bit_array_2.drv<63:0>.n71 hgu_cdac_8bit_array_2.drv<63:0> 0.321667
R7359 hgu_cdac_8bit_array_2.drv<63:0>.n1 hgu_cdac_8bit_array_2.drv<63:0>.n272 0.317975
R7360 hgu_cdac_8bit_array_2.drv<63:0>.n375 hgu_cdac_8bit_array_2.drv<63:0> 0.313448
R7361 hgu_cdac_8bit_array_2.drv<63:0>.n0 hgu_cdac_8bit_array_2.drv<63:0>.n32 0.300856
R7362 hgu_cdac_8bit_array_2.drv<63:0>.n137 hgu_cdac_8bit_array_2.drv<63:0>.n136 0.297179
R7363 hgu_cdac_8bit_array_2.drv<63:0>.n36 hgu_cdac_8bit_array_2.drv<63:0>.n35 0.297179
R7364 hgu_cdac_8bit_array_2.drv<63:0>.n16 hgu_cdac_8bit_array_2.drv<63:0>.n15 0.297179
R7365 hgu_cdac_8bit_array_2.drv<63:0>.n19 hgu_cdac_8bit_array_2.drv<63:0>.n18 0.297179
R7366 hgu_cdac_8bit_array_2.drv<63:0>.n5 hgu_cdac_8bit_array_2.drv<63:0>.n4 0.297179
R7367 hgu_cdac_8bit_array_2.drv<63:0>.n10 hgu_cdac_8bit_array_2.drv<63:0>.n9 0.297179
R7368 hgu_cdac_8bit_array_2.drv<63:0>.n116 hgu_cdac_8bit_array_2.drv<63:0>.n115 0.297179
R7369 hgu_cdac_8bit_array_2.drv<63:0>.n119 hgu_cdac_8bit_array_2.drv<63:0>.n118 0.297179
R7370 hgu_cdac_8bit_array_2.drv<63:0>.n131 hgu_cdac_8bit_array_2.drv<63:0>.n130 0.297179
R7371 hgu_cdac_8bit_array_2.drv<63:0>.n261 hgu_cdac_8bit_array_2.drv<63:0>.n260 0.297179
R7372 hgu_cdac_8bit_array_2.drv<63:0>.n258 hgu_cdac_8bit_array_2.drv<63:0>.n257 0.297179
R7373 hgu_cdac_8bit_array_2.drv<63:0>.n246 hgu_cdac_8bit_array_2.drv<63:0>.n245 0.297179
R7374 hgu_cdac_8bit_array_2.drv<63:0>.n230 hgu_cdac_8bit_array_2.drv<63:0>.n229 0.297179
R7375 hgu_cdac_8bit_array_2.drv<63:0>.n225 hgu_cdac_8bit_array_2.drv<63:0>.n224 0.297179
R7376 hgu_cdac_8bit_array_2.drv<63:0>.n213 hgu_cdac_8bit_array_2.drv<63:0>.n212 0.297179
R7377 hgu_cdac_8bit_array_2.drv<63:0>.n210 hgu_cdac_8bit_array_2.drv<63:0>.n209 0.297179
R7378 hgu_cdac_8bit_array_2.drv<63:0>.n198 hgu_cdac_8bit_array_2.drv<63:0>.n197 0.297179
R7379 hgu_cdac_8bit_array_2.drv<63:0>.n194 hgu_cdac_8bit_array_2.drv<63:0>.n193 0.297179
R7380 hgu_cdac_8bit_array_2.drv<63:0>.n180 hgu_cdac_8bit_array_2.drv<63:0>.n179 0.297179
R7381 hgu_cdac_8bit_array_2.drv<63:0>.n165 hgu_cdac_8bit_array_2.drv<63:0>.n164 0.297179
R7382 hgu_cdac_8bit_array_2.drv<63:0>.n168 hgu_cdac_8bit_array_2.drv<63:0>.n167 0.297179
R7383 hgu_cdac_8bit_array_2.drv<63:0>.n162 hgu_cdac_8bit_array_2.drv<63:0>.n161 0.297179
R7384 hgu_cdac_8bit_array_2.drv<63:0>.n151 hgu_cdac_8bit_array_2.drv<63:0>.n150 0.297179
R7385 hgu_cdac_8bit_array_2.drv<63:0>.n135 hgu_cdac_8bit_array_2.drv<63:0>.n134 0.297179
R7386 hgu_cdac_8bit_array_2.drv<63:0>.n65 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7387 hgu_cdac_8bit_array_2.drv<63:0>.n74 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7388 hgu_cdac_8bit_array_2.drv<63:0>.n83 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7389 hgu_cdac_8bit_array_2.drv<63:0>.n92 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7390 hgu_cdac_8bit_array_2.drv<63:0>.n101 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7391 hgu_cdac_8bit_array_2.drv<63:0>.n110 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7392 hgu_cdac_8bit_array_2.drv<63:0>.n599 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7393 hgu_cdac_8bit_array_2.drv<63:0>.n590 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7394 hgu_cdac_8bit_array_2.drv<63:0>.n581 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7395 hgu_cdac_8bit_array_2.drv<63:0>.n572 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7396 hgu_cdac_8bit_array_2.drv<63:0>.n563 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7397 hgu_cdac_8bit_array_2.drv<63:0>.n554 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7398 hgu_cdac_8bit_array_2.drv<63:0>.n545 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7399 hgu_cdac_8bit_array_2.drv<63:0>.n536 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7400 hgu_cdac_8bit_array_2.drv<63:0>.n527 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7401 hgu_cdac_8bit_array_2.drv<63:0>.n518 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7402 hgu_cdac_8bit_array_2.drv<63:0>.n509 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7403 hgu_cdac_8bit_array_2.drv<63:0>.n499 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7404 hgu_cdac_8bit_array_2.drv<63:0>.n490 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7405 hgu_cdac_8bit_array_2.drv<63:0>.n481 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7406 hgu_cdac_8bit_array_2.drv<63:0>.n472 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7407 hgu_cdac_8bit_array_2.drv<63:0>.n463 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7408 hgu_cdac_8bit_array_2.drv<63:0>.n454 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7409 hgu_cdac_8bit_array_2.drv<63:0>.n445 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7410 hgu_cdac_8bit_array_2.drv<63:0>.n436 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7411 hgu_cdac_8bit_array_2.drv<63:0>.n427 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7412 hgu_cdac_8bit_array_2.drv<63:0>.n418 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7413 hgu_cdac_8bit_array_2.drv<63:0>.n409 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7414 hgu_cdac_8bit_array_2.drv<63:0>.n400 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7415 hgu_cdac_8bit_array_2.drv<63:0>.n391 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7416 hgu_cdac_8bit_array_2.drv<63:0>.n382 hgu_cdac_8bit_array_2.drv<63:0> 0.2966
R7417 hgu_cdac_8bit_array_2.drv<63:0>.n169 hgu_cdac_8bit_array_2.drv<63:0>.n162 0.261276
R7418 hgu_cdac_8bit_array_2.drv<63:0>.n138 hgu_cdac_8bit_array_2.drv<63:0>.n137 0.256966
R7419 hgu_cdac_8bit_array_2.drv<63:0>.n2 hgu_cdac_8bit_array_2.drv<63:0>.n148 0.247662
R7420 hgu_cdac_8bit_array_2.drv<63:0>.n33 hgu_cdac_8bit_array_2.drv<63:0>.n30 0.245708
R7421 hgu_cdac_8bit_array_2.drv<63:0>.n243 hgu_cdac_8bit_array_2.drv<63:0>.n242 0.245708
R7422 hgu_cdac_8bit_array_2.drv<63:0>.n231 hgu_cdac_8bit_array_2.drv<63:0>.n227 0.245708
R7423 hgu_cdac_8bit_array_2.drv<63:0>.n195 hgu_cdac_8bit_array_2.drv<63:0>.n191 0.245708
R7424 hgu_cdac_8bit_array_2.drv<63:0>.n11 hgu_cdac_8bit_array_2.drv<63:0>.n7 0.242032
R7425 hgu_cdac_8bit_array_2.drv<63:0>.n120 hgu_cdac_8bit_array_2.drv<63:0>.n116 0.18369
R7426 hgu_cdac_8bit_array_2.drv<63:0>.n181 hgu_cdac_8bit_array_2.drv<63:0>.n180 0.18369
R7427 hgu_cdac_8bit_array_2.drv<63:0>.n587 hgu_cdac_8bit_array_2.drv<63:0>.n146 0.18292
R7428 hgu_cdac_8bit_array_2.drv<63:0>.n578 hgu_cdac_8bit_array_2.drv<63:0>.n159 0.18292
R7429 hgu_cdac_8bit_array_2.drv<63:0>.n569 hgu_cdac_8bit_array_2.drv<63:0>.n177 0.18292
R7430 hgu_cdac_8bit_array_2.drv<63:0>.n560 hgu_cdac_8bit_array_2.drv<63:0>.n189 0.18292
R7431 hgu_cdac_8bit_array_2.drv<63:0>.n551 hgu_cdac_8bit_array_2.drv<63:0>.n207 0.18292
R7432 hgu_cdac_8bit_array_2.drv<63:0>.n542 hgu_cdac_8bit_array_2.drv<63:0>.n222 0.18292
R7433 hgu_cdac_8bit_array_2.drv<63:0>.n533 hgu_cdac_8bit_array_2.drv<63:0>.n240 0.18292
R7434 hgu_cdac_8bit_array_2.drv<63:0>.n596 hgu_cdac_8bit_array_2.drv<63:0>.n128 0.182836
R7435 hgu_cdac_8bit_array_2.drv<63:0>.n113 hgu_cdac_8bit_array_2.drv<63:0>.n13 0.182836
R7436 hgu_cdac_8bit_array_2.drv<63:0>.n104 hgu_cdac_8bit_array_2.drv<63:0>.n28 0.182836
R7437 hgu_cdac_8bit_array_2.drv<63:0>.n95 hgu_cdac_8bit_array_2.drv<63:0>.n45 0.182836
R7438 hgu_cdac_8bit_array_2.drv<63:0>.n86 hgu_cdac_8bit_array_2.drv<63:0>.n53 0.182836
R7439 hgu_cdac_8bit_array_2.drv<63:0>.n524 hgu_cdac_8bit_array_2.drv<63:0>.n255 0.182836
R7440 hgu_cdac_8bit_array_2.drv<63:0>.n515 hgu_cdac_8bit_array_2.drv<63:0>.n270 0.182836
R7441 hgu_cdac_8bit_array_2.drv<63:0>.n506 hgu_cdac_8bit_array_2.drv<63:0>.n280 0.182836
R7442 hgu_cdac_8bit_array_2.drv<63:0>.n146 hgu_cdac_8bit_array_2.drv<63:0>.n145 0.149226
R7443 hgu_cdac_8bit_array_2.drv<63:0>.n159 hgu_cdac_8bit_array_2.drv<63:0>.n158 0.149226
R7444 hgu_cdac_8bit_array_2.drv<63:0>.n177 hgu_cdac_8bit_array_2.drv<63:0>.n176 0.149226
R7445 hgu_cdac_8bit_array_2.drv<63:0>.n189 hgu_cdac_8bit_array_2.drv<63:0>.n188 0.149226
R7446 hgu_cdac_8bit_array_2.drv<63:0>.n207 hgu_cdac_8bit_array_2.drv<63:0>.n206 0.149226
R7447 hgu_cdac_8bit_array_2.drv<63:0>.n222 hgu_cdac_8bit_array_2.drv<63:0>.n221 0.149226
R7448 hgu_cdac_8bit_array_2.drv<63:0>.n240 hgu_cdac_8bit_array_2.drv<63:0>.n239 0.149226
R7449 hgu_cdac_8bit_array_2.drv<63:0>.n53 hgu_cdac_8bit_array_2.drv<63:0>.n52 0.149114
R7450 hgu_cdac_8bit_array_2.drv<63:0>.n45 hgu_cdac_8bit_array_2.drv<63:0>.n44 0.149114
R7451 hgu_cdac_8bit_array_2.drv<63:0>.n28 hgu_cdac_8bit_array_2.drv<63:0>.n27 0.149114
R7452 hgu_cdac_8bit_array_2.drv<63:0>.n128 hgu_cdac_8bit_array_2.drv<63:0>.n127 0.149114
R7453 hgu_cdac_8bit_array_2.drv<63:0>.n255 hgu_cdac_8bit_array_2.drv<63:0>.n254 0.149114
R7454 hgu_cdac_8bit_array_2.drv<63:0>.n270 hgu_cdac_8bit_array_2.drv<63:0>.n269 0.149114
R7455 hgu_cdac_8bit_array_2.drv<63:0>.n280 hgu_cdac_8bit_array_2.drv<63:0>.n279 0.149114
R7456 hgu_cdac_8bit_array_2.drv<63:0>.n247 hgu_cdac_8bit_array_2.drv<63:0>.n243 0.0962031
R7457 hgu_cdac_8bit_array_2.drv<63:0>.n37 hgu_cdac_8bit_array_2.drv<63:0>.n33 0.0825312
R7458 hgu_cdac_8bit_array_2.drv<63:0>.n232 hgu_cdac_8bit_array_2.drv<63:0>.n231 0.0805781
R7459 hgu_cdac_8bit_array_2.drv<63:0>.n68 hgu_cdac_8bit_array_2.drv<63:0>.n67 0.0716912
R7460 hgu_cdac_8bit_array_2.drv<63:0>.n69 hgu_cdac_8bit_array_2.drv<63:0>.n68 0.0716912
R7461 hgu_cdac_8bit_array_2.drv<63:0>.n77 hgu_cdac_8bit_array_2.drv<63:0>.n76 0.0716912
R7462 hgu_cdac_8bit_array_2.drv<63:0>.n78 hgu_cdac_8bit_array_2.drv<63:0>.n77 0.0716912
R7463 hgu_cdac_8bit_array_2.drv<63:0>.n86 hgu_cdac_8bit_array_2.drv<63:0>.n85 0.0716912
R7464 hgu_cdac_8bit_array_2.drv<63:0>.n87 hgu_cdac_8bit_array_2.drv<63:0>.n86 0.0716912
R7465 hgu_cdac_8bit_array_2.drv<63:0>.n95 hgu_cdac_8bit_array_2.drv<63:0>.n94 0.0716912
R7466 hgu_cdac_8bit_array_2.drv<63:0>.n96 hgu_cdac_8bit_array_2.drv<63:0>.n95 0.0716912
R7467 hgu_cdac_8bit_array_2.drv<63:0>.n104 hgu_cdac_8bit_array_2.drv<63:0>.n103 0.0716912
R7468 hgu_cdac_8bit_array_2.drv<63:0>.n105 hgu_cdac_8bit_array_2.drv<63:0>.n104 0.0716912
R7469 hgu_cdac_8bit_array_2.drv<63:0>.n113 hgu_cdac_8bit_array_2.drv<63:0>.n112 0.0716912
R7470 hgu_cdac_8bit_array_2.drv<63:0>.n597 hgu_cdac_8bit_array_2.drv<63:0>.n596 0.0716912
R7471 hgu_cdac_8bit_array_2.drv<63:0>.n596 hgu_cdac_8bit_array_2.drv<63:0>.n595 0.0716912
R7472 hgu_cdac_8bit_array_2.drv<63:0>.n588 hgu_cdac_8bit_array_2.drv<63:0>.n587 0.0716912
R7473 hgu_cdac_8bit_array_2.drv<63:0>.n587 hgu_cdac_8bit_array_2.drv<63:0>.n586 0.0716912
R7474 hgu_cdac_8bit_array_2.drv<63:0>.n579 hgu_cdac_8bit_array_2.drv<63:0>.n578 0.0716912
R7475 hgu_cdac_8bit_array_2.drv<63:0>.n578 hgu_cdac_8bit_array_2.drv<63:0>.n577 0.0716912
R7476 hgu_cdac_8bit_array_2.drv<63:0>.n570 hgu_cdac_8bit_array_2.drv<63:0>.n569 0.0716912
R7477 hgu_cdac_8bit_array_2.drv<63:0>.n569 hgu_cdac_8bit_array_2.drv<63:0>.n568 0.0716912
R7478 hgu_cdac_8bit_array_2.drv<63:0>.n561 hgu_cdac_8bit_array_2.drv<63:0>.n560 0.0716912
R7479 hgu_cdac_8bit_array_2.drv<63:0>.n560 hgu_cdac_8bit_array_2.drv<63:0>.n559 0.0716912
R7480 hgu_cdac_8bit_array_2.drv<63:0>.n552 hgu_cdac_8bit_array_2.drv<63:0>.n551 0.0716912
R7481 hgu_cdac_8bit_array_2.drv<63:0>.n551 hgu_cdac_8bit_array_2.drv<63:0>.n550 0.0716912
R7482 hgu_cdac_8bit_array_2.drv<63:0>.n543 hgu_cdac_8bit_array_2.drv<63:0>.n542 0.0716912
R7483 hgu_cdac_8bit_array_2.drv<63:0>.n542 hgu_cdac_8bit_array_2.drv<63:0>.n541 0.0716912
R7484 hgu_cdac_8bit_array_2.drv<63:0>.n534 hgu_cdac_8bit_array_2.drv<63:0>.n533 0.0716912
R7485 hgu_cdac_8bit_array_2.drv<63:0>.n533 hgu_cdac_8bit_array_2.drv<63:0>.n532 0.0716912
R7486 hgu_cdac_8bit_array_2.drv<63:0>.n525 hgu_cdac_8bit_array_2.drv<63:0>.n524 0.0716912
R7487 hgu_cdac_8bit_array_2.drv<63:0>.n524 hgu_cdac_8bit_array_2.drv<63:0>.n523 0.0716912
R7488 hgu_cdac_8bit_array_2.drv<63:0>.n516 hgu_cdac_8bit_array_2.drv<63:0>.n515 0.0716912
R7489 hgu_cdac_8bit_array_2.drv<63:0>.n515 hgu_cdac_8bit_array_2.drv<63:0>.n514 0.0716912
R7490 hgu_cdac_8bit_array_2.drv<63:0>.n507 hgu_cdac_8bit_array_2.drv<63:0>.n506 0.0716912
R7491 hgu_cdac_8bit_array_2.drv<63:0>.n506 hgu_cdac_8bit_array_2.drv<63:0>.n505 0.0716912
R7492 hgu_cdac_8bit_array_2.drv<63:0>.n497 hgu_cdac_8bit_array_2.drv<63:0>.n496 0.0716912
R7493 hgu_cdac_8bit_array_2.drv<63:0>.n496 hgu_cdac_8bit_array_2.drv<63:0>.n495 0.0716912
R7494 hgu_cdac_8bit_array_2.drv<63:0>.n488 hgu_cdac_8bit_array_2.drv<63:0>.n487 0.0716912
R7495 hgu_cdac_8bit_array_2.drv<63:0>.n487 hgu_cdac_8bit_array_2.drv<63:0>.n486 0.0716912
R7496 hgu_cdac_8bit_array_2.drv<63:0>.n479 hgu_cdac_8bit_array_2.drv<63:0>.n478 0.0716912
R7497 hgu_cdac_8bit_array_2.drv<63:0>.n478 hgu_cdac_8bit_array_2.drv<63:0>.n477 0.0716912
R7498 hgu_cdac_8bit_array_2.drv<63:0>.n470 hgu_cdac_8bit_array_2.drv<63:0>.n469 0.0716912
R7499 hgu_cdac_8bit_array_2.drv<63:0>.n469 hgu_cdac_8bit_array_2.drv<63:0>.n468 0.0716912
R7500 hgu_cdac_8bit_array_2.drv<63:0>.n461 hgu_cdac_8bit_array_2.drv<63:0>.n460 0.0716912
R7501 hgu_cdac_8bit_array_2.drv<63:0>.n460 hgu_cdac_8bit_array_2.drv<63:0>.n459 0.0716912
R7502 hgu_cdac_8bit_array_2.drv<63:0>.n452 hgu_cdac_8bit_array_2.drv<63:0>.n451 0.0716912
R7503 hgu_cdac_8bit_array_2.drv<63:0>.n451 hgu_cdac_8bit_array_2.drv<63:0>.n450 0.0716912
R7504 hgu_cdac_8bit_array_2.drv<63:0>.n443 hgu_cdac_8bit_array_2.drv<63:0>.n442 0.0716912
R7505 hgu_cdac_8bit_array_2.drv<63:0>.n442 hgu_cdac_8bit_array_2.drv<63:0>.n441 0.0716912
R7506 hgu_cdac_8bit_array_2.drv<63:0>.n434 hgu_cdac_8bit_array_2.drv<63:0>.n433 0.0716912
R7507 hgu_cdac_8bit_array_2.drv<63:0>.n433 hgu_cdac_8bit_array_2.drv<63:0>.n432 0.0716912
R7508 hgu_cdac_8bit_array_2.drv<63:0>.n425 hgu_cdac_8bit_array_2.drv<63:0>.n424 0.0716912
R7509 hgu_cdac_8bit_array_2.drv<63:0>.n424 hgu_cdac_8bit_array_2.drv<63:0>.n423 0.0716912
R7510 hgu_cdac_8bit_array_2.drv<63:0>.n416 hgu_cdac_8bit_array_2.drv<63:0>.n415 0.0716912
R7511 hgu_cdac_8bit_array_2.drv<63:0>.n415 hgu_cdac_8bit_array_2.drv<63:0>.n414 0.0716912
R7512 hgu_cdac_8bit_array_2.drv<63:0>.n407 hgu_cdac_8bit_array_2.drv<63:0>.n406 0.0716912
R7513 hgu_cdac_8bit_array_2.drv<63:0>.n406 hgu_cdac_8bit_array_2.drv<63:0>.n405 0.0716912
R7514 hgu_cdac_8bit_array_2.drv<63:0>.n398 hgu_cdac_8bit_array_2.drv<63:0>.n397 0.0716912
R7515 hgu_cdac_8bit_array_2.drv<63:0>.n397 hgu_cdac_8bit_array_2.drv<63:0>.n396 0.0716912
R7516 hgu_cdac_8bit_array_2.drv<63:0>.n389 hgu_cdac_8bit_array_2.drv<63:0>.n388 0.0716912
R7517 hgu_cdac_8bit_array_2.drv<63:0>.n388 hgu_cdac_8bit_array_2.drv<63:0>.n387 0.0716912
R7518 hgu_cdac_8bit_array_2.drv<63:0>.n380 hgu_cdac_8bit_array_2.drv<63:0>.n379 0.0716912
R7519 hgu_cdac_8bit_array_2.drv<63:0>.n379 hgu_cdac_8bit_array_2.drv<63:0>.n378 0.0716912
R7520 hgu_cdac_8bit_array_2.drv<63:0>.n63 hgu_cdac_8bit_array_2.drv<63:0>.n62 0.0716912
R7521 hgu_cdac_8bit_array_2.drv<63:0>.n60 hgu_cdac_8bit_array_2.drv<63:0>.n59 0.0716912
R7522 hgu_cdac_8bit_array_2.drv<63:0>.n52 hgu_cdac_8bit_array_2.drv<63:0>.n51 0.0716912
R7523 hgu_cdac_8bit_array_2.drv<63:0>.n44 hgu_cdac_8bit_array_2.drv<63:0>.n43 0.0716912
R7524 hgu_cdac_8bit_array_2.drv<63:0>.n27 hgu_cdac_8bit_array_2.drv<63:0>.n26 0.0716912
R7525 hgu_cdac_8bit_array_2.drv<63:0>.n127 hgu_cdac_8bit_array_2.drv<63:0>.n126 0.0716912
R7526 hgu_cdac_8bit_array_2.drv<63:0>.n145 hgu_cdac_8bit_array_2.drv<63:0>.n144 0.0716912
R7527 hgu_cdac_8bit_array_2.drv<63:0>.n158 hgu_cdac_8bit_array_2.drv<63:0>.n157 0.0716912
R7528 hgu_cdac_8bit_array_2.drv<63:0>.n176 hgu_cdac_8bit_array_2.drv<63:0>.n175 0.0716912
R7529 hgu_cdac_8bit_array_2.drv<63:0>.n188 hgu_cdac_8bit_array_2.drv<63:0>.n187 0.0716912
R7530 hgu_cdac_8bit_array_2.drv<63:0>.n206 hgu_cdac_8bit_array_2.drv<63:0>.n205 0.0716912
R7531 hgu_cdac_8bit_array_2.drv<63:0>.n221 hgu_cdac_8bit_array_2.drv<63:0>.n220 0.0716912
R7532 hgu_cdac_8bit_array_2.drv<63:0>.n239 hgu_cdac_8bit_array_2.drv<63:0>.n238 0.0716912
R7533 hgu_cdac_8bit_array_2.drv<63:0>.n254 hgu_cdac_8bit_array_2.drv<63:0>.n253 0.0716912
R7534 hgu_cdac_8bit_array_2.drv<63:0>.n269 hgu_cdac_8bit_array_2.drv<63:0>.n268 0.0716912
R7535 hgu_cdac_8bit_array_2.drv<63:0>.n279 hgu_cdac_8bit_array_2.drv<63:0>.n278 0.0716912
R7536 hgu_cdac_8bit_array_2.drv<63:0>.n287 hgu_cdac_8bit_array_2.drv<63:0>.n286 0.0716912
R7537 hgu_cdac_8bit_array_2.drv<63:0>.n294 hgu_cdac_8bit_array_2.drv<63:0>.n293 0.0716912
R7538 hgu_cdac_8bit_array_2.drv<63:0>.n301 hgu_cdac_8bit_array_2.drv<63:0>.n300 0.0716912
R7539 hgu_cdac_8bit_array_2.drv<63:0>.n308 hgu_cdac_8bit_array_2.drv<63:0>.n307 0.0716912
R7540 hgu_cdac_8bit_array_2.drv<63:0>.n315 hgu_cdac_8bit_array_2.drv<63:0>.n314 0.0716912
R7541 hgu_cdac_8bit_array_2.drv<63:0>.n322 hgu_cdac_8bit_array_2.drv<63:0>.n321 0.0716912
R7542 hgu_cdac_8bit_array_2.drv<63:0>.n329 hgu_cdac_8bit_array_2.drv<63:0>.n328 0.0716912
R7543 hgu_cdac_8bit_array_2.drv<63:0>.n336 hgu_cdac_8bit_array_2.drv<63:0>.n335 0.0716912
R7544 hgu_cdac_8bit_array_2.drv<63:0>.n343 hgu_cdac_8bit_array_2.drv<63:0>.n342 0.0716912
R7545 hgu_cdac_8bit_array_2.drv<63:0>.n350 hgu_cdac_8bit_array_2.drv<63:0>.n349 0.0716912
R7546 hgu_cdac_8bit_array_2.drv<63:0>.n357 hgu_cdac_8bit_array_2.drv<63:0>.n356 0.0716912
R7547 hgu_cdac_8bit_array_2.drv<63:0>.n364 hgu_cdac_8bit_array_2.drv<63:0>.n363 0.0716912
R7548 hgu_cdac_8bit_array_2.drv<63:0>.n371 hgu_cdac_8bit_array_2.drv<63:0>.n370 0.0716912
R7549 hgu_cdac_8bit_array_2.drv<63:0>.n374 hgu_cdac_8bit_array_2.drv<63:0>.n373 0.0716912
R7550 hgu_cdac_8bit_array_2.drv<63:0>.n504 hgu_cdac_8bit_array_2.drv<63:0> 0.0694333
R7551 hgu_cdac_8bit_array_2.drv<63:0>.n65 hgu_cdac_8bit_array_2.drv<63:0>.n64 0.0665339
R7552 hgu_cdac_8bit_array_2.drv<63:0>.n376 hgu_cdac_8bit_array_2.drv<63:0>.n375 0.0664894
R7553 hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_8bit_array_2.drv<63:0>.n604 0.0564853
R7554 hgu_cdac_8bit_array_2.drv<63:0>.n67 hgu_cdac_8bit_array_2.drv<63:0>.n66 0.0557941
R7555 hgu_cdac_8bit_array_2.drv<63:0>.n70 hgu_cdac_8bit_array_2.drv<63:0>.n69 0.0557941
R7556 hgu_cdac_8bit_array_2.drv<63:0>.n73 hgu_cdac_8bit_array_2.drv<63:0>.n72 0.0557941
R7557 hgu_cdac_8bit_array_2.drv<63:0>.n76 hgu_cdac_8bit_array_2.drv<63:0>.n75 0.0557941
R7558 hgu_cdac_8bit_array_2.drv<63:0>.n79 hgu_cdac_8bit_array_2.drv<63:0>.n78 0.0557941
R7559 hgu_cdac_8bit_array_2.drv<63:0>.n82 hgu_cdac_8bit_array_2.drv<63:0>.n81 0.0557941
R7560 hgu_cdac_8bit_array_2.drv<63:0>.n85 hgu_cdac_8bit_array_2.drv<63:0>.n84 0.0557941
R7561 hgu_cdac_8bit_array_2.drv<63:0>.n88 hgu_cdac_8bit_array_2.drv<63:0>.n87 0.0557941
R7562 hgu_cdac_8bit_array_2.drv<63:0>.n91 hgu_cdac_8bit_array_2.drv<63:0>.n90 0.0557941
R7563 hgu_cdac_8bit_array_2.drv<63:0>.n94 hgu_cdac_8bit_array_2.drv<63:0>.n93 0.0557941
R7564 hgu_cdac_8bit_array_2.drv<63:0>.n97 hgu_cdac_8bit_array_2.drv<63:0>.n96 0.0557941
R7565 hgu_cdac_8bit_array_2.drv<63:0>.n100 hgu_cdac_8bit_array_2.drv<63:0>.n99 0.0557941
R7566 hgu_cdac_8bit_array_2.drv<63:0>.n103 hgu_cdac_8bit_array_2.drv<63:0>.n102 0.0557941
R7567 hgu_cdac_8bit_array_2.drv<63:0>.n106 hgu_cdac_8bit_array_2.drv<63:0>.n105 0.0557941
R7568 hgu_cdac_8bit_array_2.drv<63:0>.n109 hgu_cdac_8bit_array_2.drv<63:0>.n108 0.0557941
R7569 hgu_cdac_8bit_array_2.drv<63:0>.n112 hgu_cdac_8bit_array_2.drv<63:0>.n111 0.0557941
R7570 hgu_cdac_8bit_array_2.drv<63:0>.n604 hgu_cdac_8bit_array_2.drv<63:0>.n603 0.0557941
R7571 hgu_cdac_8bit_array_2.drv<63:0>.n601 hgu_cdac_8bit_array_2.drv<63:0>.n600 0.0557941
R7572 hgu_cdac_8bit_array_2.drv<63:0>.n598 hgu_cdac_8bit_array_2.drv<63:0>.n597 0.0557941
R7573 hgu_cdac_8bit_array_2.drv<63:0>.n595 hgu_cdac_8bit_array_2.drv<63:0>.n594 0.0557941
R7574 hgu_cdac_8bit_array_2.drv<63:0>.n592 hgu_cdac_8bit_array_2.drv<63:0>.n591 0.0557941
R7575 hgu_cdac_8bit_array_2.drv<63:0>.n589 hgu_cdac_8bit_array_2.drv<63:0>.n588 0.0557941
R7576 hgu_cdac_8bit_array_2.drv<63:0>.n586 hgu_cdac_8bit_array_2.drv<63:0>.n585 0.0557941
R7577 hgu_cdac_8bit_array_2.drv<63:0>.n583 hgu_cdac_8bit_array_2.drv<63:0>.n582 0.0557941
R7578 hgu_cdac_8bit_array_2.drv<63:0>.n580 hgu_cdac_8bit_array_2.drv<63:0>.n579 0.0557941
R7579 hgu_cdac_8bit_array_2.drv<63:0>.n577 hgu_cdac_8bit_array_2.drv<63:0>.n576 0.0557941
R7580 hgu_cdac_8bit_array_2.drv<63:0>.n574 hgu_cdac_8bit_array_2.drv<63:0>.n573 0.0557941
R7581 hgu_cdac_8bit_array_2.drv<63:0>.n571 hgu_cdac_8bit_array_2.drv<63:0>.n570 0.0557941
R7582 hgu_cdac_8bit_array_2.drv<63:0>.n568 hgu_cdac_8bit_array_2.drv<63:0>.n567 0.0557941
R7583 hgu_cdac_8bit_array_2.drv<63:0>.n565 hgu_cdac_8bit_array_2.drv<63:0>.n564 0.0557941
R7584 hgu_cdac_8bit_array_2.drv<63:0>.n562 hgu_cdac_8bit_array_2.drv<63:0>.n561 0.0557941
R7585 hgu_cdac_8bit_array_2.drv<63:0>.n559 hgu_cdac_8bit_array_2.drv<63:0>.n558 0.0557941
R7586 hgu_cdac_8bit_array_2.drv<63:0>.n556 hgu_cdac_8bit_array_2.drv<63:0>.n555 0.0557941
R7587 hgu_cdac_8bit_array_2.drv<63:0>.n553 hgu_cdac_8bit_array_2.drv<63:0>.n552 0.0557941
R7588 hgu_cdac_8bit_array_2.drv<63:0>.n550 hgu_cdac_8bit_array_2.drv<63:0>.n549 0.0557941
R7589 hgu_cdac_8bit_array_2.drv<63:0>.n547 hgu_cdac_8bit_array_2.drv<63:0>.n546 0.0557941
R7590 hgu_cdac_8bit_array_2.drv<63:0>.n544 hgu_cdac_8bit_array_2.drv<63:0>.n543 0.0557941
R7591 hgu_cdac_8bit_array_2.drv<63:0>.n541 hgu_cdac_8bit_array_2.drv<63:0>.n540 0.0557941
R7592 hgu_cdac_8bit_array_2.drv<63:0>.n538 hgu_cdac_8bit_array_2.drv<63:0>.n537 0.0557941
R7593 hgu_cdac_8bit_array_2.drv<63:0>.n535 hgu_cdac_8bit_array_2.drv<63:0>.n534 0.0557941
R7594 hgu_cdac_8bit_array_2.drv<63:0>.n532 hgu_cdac_8bit_array_2.drv<63:0>.n531 0.0557941
R7595 hgu_cdac_8bit_array_2.drv<63:0>.n529 hgu_cdac_8bit_array_2.drv<63:0>.n528 0.0557941
R7596 hgu_cdac_8bit_array_2.drv<63:0>.n526 hgu_cdac_8bit_array_2.drv<63:0>.n525 0.0557941
R7597 hgu_cdac_8bit_array_2.drv<63:0>.n523 hgu_cdac_8bit_array_2.drv<63:0>.n522 0.0557941
R7598 hgu_cdac_8bit_array_2.drv<63:0>.n520 hgu_cdac_8bit_array_2.drv<63:0>.n519 0.0557941
R7599 hgu_cdac_8bit_array_2.drv<63:0>.n517 hgu_cdac_8bit_array_2.drv<63:0>.n516 0.0557941
R7600 hgu_cdac_8bit_array_2.drv<63:0>.n514 hgu_cdac_8bit_array_2.drv<63:0>.n513 0.0557941
R7601 hgu_cdac_8bit_array_2.drv<63:0>.n511 hgu_cdac_8bit_array_2.drv<63:0>.n510 0.0557941
R7602 hgu_cdac_8bit_array_2.drv<63:0>.n508 hgu_cdac_8bit_array_2.drv<63:0>.n507 0.0557941
R7603 hgu_cdac_8bit_array_2.drv<63:0>.n501 hgu_cdac_8bit_array_2.drv<63:0>.n500 0.0557941
R7604 hgu_cdac_8bit_array_2.drv<63:0>.n498 hgu_cdac_8bit_array_2.drv<63:0>.n497 0.0557941
R7605 hgu_cdac_8bit_array_2.drv<63:0>.n495 hgu_cdac_8bit_array_2.drv<63:0>.n494 0.0557941
R7606 hgu_cdac_8bit_array_2.drv<63:0>.n492 hgu_cdac_8bit_array_2.drv<63:0>.n491 0.0557941
R7607 hgu_cdac_8bit_array_2.drv<63:0>.n489 hgu_cdac_8bit_array_2.drv<63:0>.n488 0.0557941
R7608 hgu_cdac_8bit_array_2.drv<63:0>.n486 hgu_cdac_8bit_array_2.drv<63:0>.n485 0.0557941
R7609 hgu_cdac_8bit_array_2.drv<63:0>.n483 hgu_cdac_8bit_array_2.drv<63:0>.n482 0.0557941
R7610 hgu_cdac_8bit_array_2.drv<63:0>.n480 hgu_cdac_8bit_array_2.drv<63:0>.n479 0.0557941
R7611 hgu_cdac_8bit_array_2.drv<63:0>.n477 hgu_cdac_8bit_array_2.drv<63:0>.n476 0.0557941
R7612 hgu_cdac_8bit_array_2.drv<63:0>.n474 hgu_cdac_8bit_array_2.drv<63:0>.n473 0.0557941
R7613 hgu_cdac_8bit_array_2.drv<63:0>.n471 hgu_cdac_8bit_array_2.drv<63:0>.n470 0.0557941
R7614 hgu_cdac_8bit_array_2.drv<63:0>.n468 hgu_cdac_8bit_array_2.drv<63:0>.n467 0.0557941
R7615 hgu_cdac_8bit_array_2.drv<63:0>.n465 hgu_cdac_8bit_array_2.drv<63:0>.n464 0.0557941
R7616 hgu_cdac_8bit_array_2.drv<63:0>.n462 hgu_cdac_8bit_array_2.drv<63:0>.n461 0.0557941
R7617 hgu_cdac_8bit_array_2.drv<63:0>.n459 hgu_cdac_8bit_array_2.drv<63:0>.n458 0.0557941
R7618 hgu_cdac_8bit_array_2.drv<63:0>.n456 hgu_cdac_8bit_array_2.drv<63:0>.n455 0.0557941
R7619 hgu_cdac_8bit_array_2.drv<63:0>.n453 hgu_cdac_8bit_array_2.drv<63:0>.n452 0.0557941
R7620 hgu_cdac_8bit_array_2.drv<63:0>.n450 hgu_cdac_8bit_array_2.drv<63:0>.n449 0.0557941
R7621 hgu_cdac_8bit_array_2.drv<63:0>.n447 hgu_cdac_8bit_array_2.drv<63:0>.n446 0.0557941
R7622 hgu_cdac_8bit_array_2.drv<63:0>.n444 hgu_cdac_8bit_array_2.drv<63:0>.n443 0.0557941
R7623 hgu_cdac_8bit_array_2.drv<63:0>.n441 hgu_cdac_8bit_array_2.drv<63:0>.n440 0.0557941
R7624 hgu_cdac_8bit_array_2.drv<63:0>.n438 hgu_cdac_8bit_array_2.drv<63:0>.n437 0.0557941
R7625 hgu_cdac_8bit_array_2.drv<63:0>.n435 hgu_cdac_8bit_array_2.drv<63:0>.n434 0.0557941
R7626 hgu_cdac_8bit_array_2.drv<63:0>.n432 hgu_cdac_8bit_array_2.drv<63:0>.n431 0.0557941
R7627 hgu_cdac_8bit_array_2.drv<63:0>.n429 hgu_cdac_8bit_array_2.drv<63:0>.n428 0.0557941
R7628 hgu_cdac_8bit_array_2.drv<63:0>.n426 hgu_cdac_8bit_array_2.drv<63:0>.n425 0.0557941
R7629 hgu_cdac_8bit_array_2.drv<63:0>.n423 hgu_cdac_8bit_array_2.drv<63:0>.n422 0.0557941
R7630 hgu_cdac_8bit_array_2.drv<63:0>.n420 hgu_cdac_8bit_array_2.drv<63:0>.n419 0.0557941
R7631 hgu_cdac_8bit_array_2.drv<63:0>.n417 hgu_cdac_8bit_array_2.drv<63:0>.n416 0.0557941
R7632 hgu_cdac_8bit_array_2.drv<63:0>.n414 hgu_cdac_8bit_array_2.drv<63:0>.n413 0.0557941
R7633 hgu_cdac_8bit_array_2.drv<63:0>.n411 hgu_cdac_8bit_array_2.drv<63:0>.n410 0.0557941
R7634 hgu_cdac_8bit_array_2.drv<63:0>.n408 hgu_cdac_8bit_array_2.drv<63:0>.n407 0.0557941
R7635 hgu_cdac_8bit_array_2.drv<63:0>.n405 hgu_cdac_8bit_array_2.drv<63:0>.n404 0.0557941
R7636 hgu_cdac_8bit_array_2.drv<63:0>.n402 hgu_cdac_8bit_array_2.drv<63:0>.n401 0.0557941
R7637 hgu_cdac_8bit_array_2.drv<63:0>.n399 hgu_cdac_8bit_array_2.drv<63:0>.n398 0.0557941
R7638 hgu_cdac_8bit_array_2.drv<63:0>.n396 hgu_cdac_8bit_array_2.drv<63:0>.n395 0.0557941
R7639 hgu_cdac_8bit_array_2.drv<63:0>.n393 hgu_cdac_8bit_array_2.drv<63:0>.n392 0.0557941
R7640 hgu_cdac_8bit_array_2.drv<63:0>.n390 hgu_cdac_8bit_array_2.drv<63:0>.n389 0.0557941
R7641 hgu_cdac_8bit_array_2.drv<63:0>.n387 hgu_cdac_8bit_array_2.drv<63:0>.n386 0.0557941
R7642 hgu_cdac_8bit_array_2.drv<63:0>.n384 hgu_cdac_8bit_array_2.drv<63:0>.n383 0.0557941
R7643 hgu_cdac_8bit_array_2.drv<63:0>.n381 hgu_cdac_8bit_array_2.drv<63:0>.n380 0.0557941
R7644 hgu_cdac_8bit_array_2.drv<63:0>.n378 hgu_cdac_8bit_array_2.drv<63:0>.n377 0.0557941
R7645 hgu_cdac_8bit_array_2.drv<63:0>.n62 hgu_cdac_8bit_array_2.drv<63:0>.n61 0.0557941
R7646 hgu_cdac_8bit_array_2.drv<63:0>.n55 hgu_cdac_8bit_array_2.drv<63:0>.n54 0.0557941
R7647 hgu_cdac_8bit_array_2.drv<63:0>.n56 hgu_cdac_8bit_array_2.drv<63:0>.n55 0.0557941
R7648 hgu_cdac_8bit_array_2.drv<63:0>.n57 hgu_cdac_8bit_array_2.drv<63:0>.n56 0.0557941
R7649 hgu_cdac_8bit_array_2.drv<63:0>.n58 hgu_cdac_8bit_array_2.drv<63:0>.n57 0.0557941
R7650 hgu_cdac_8bit_array_2.drv<63:0>.n59 hgu_cdac_8bit_array_2.drv<63:0>.n58 0.0557941
R7651 hgu_cdac_8bit_array_2.drv<63:0>.n47 hgu_cdac_8bit_array_2.drv<63:0>.n46 0.0557941
R7652 hgu_cdac_8bit_array_2.drv<63:0>.n48 hgu_cdac_8bit_array_2.drv<63:0>.n47 0.0557941
R7653 hgu_cdac_8bit_array_2.drv<63:0>.n49 hgu_cdac_8bit_array_2.drv<63:0>.n48 0.0557941
R7654 hgu_cdac_8bit_array_2.drv<63:0>.n50 hgu_cdac_8bit_array_2.drv<63:0>.n49 0.0557941
R7655 hgu_cdac_8bit_array_2.drv<63:0>.n51 hgu_cdac_8bit_array_2.drv<63:0>.n50 0.0557941
R7656 hgu_cdac_8bit_array_2.drv<63:0>.n39 hgu_cdac_8bit_array_2.drv<63:0>.n38 0.0557941
R7657 hgu_cdac_8bit_array_2.drv<63:0>.n40 hgu_cdac_8bit_array_2.drv<63:0>.n39 0.0557941
R7658 hgu_cdac_8bit_array_2.drv<63:0>.n41 hgu_cdac_8bit_array_2.drv<63:0>.n40 0.0557941
R7659 hgu_cdac_8bit_array_2.drv<63:0>.n42 hgu_cdac_8bit_array_2.drv<63:0>.n41 0.0557941
R7660 hgu_cdac_8bit_array_2.drv<63:0>.n43 hgu_cdac_8bit_array_2.drv<63:0>.n42 0.0557941
R7661 hgu_cdac_8bit_array_2.drv<63:0>.n22 hgu_cdac_8bit_array_2.drv<63:0>.n21 0.0557941
R7662 hgu_cdac_8bit_array_2.drv<63:0>.n23 hgu_cdac_8bit_array_2.drv<63:0>.n22 0.0557941
R7663 hgu_cdac_8bit_array_2.drv<63:0>.n24 hgu_cdac_8bit_array_2.drv<63:0>.n23 0.0557941
R7664 hgu_cdac_8bit_array_2.drv<63:0>.n25 hgu_cdac_8bit_array_2.drv<63:0>.n24 0.0557941
R7665 hgu_cdac_8bit_array_2.drv<63:0>.n26 hgu_cdac_8bit_array_2.drv<63:0>.n25 0.0557941
R7666 hgu_cdac_8bit_array_2.drv<63:0>.n126 hgu_cdac_8bit_array_2.drv<63:0>.n125 0.0557941
R7667 hgu_cdac_8bit_array_2.drv<63:0>.n125 hgu_cdac_8bit_array_2.drv<63:0>.n124 0.0557941
R7668 hgu_cdac_8bit_array_2.drv<63:0>.n124 hgu_cdac_8bit_array_2.drv<63:0>.n123 0.0557941
R7669 hgu_cdac_8bit_array_2.drv<63:0>.n123 hgu_cdac_8bit_array_2.drv<63:0>.n122 0.0557941
R7670 hgu_cdac_8bit_array_2.drv<63:0>.n122 hgu_cdac_8bit_array_2.drv<63:0>.n121 0.0557941
R7671 hgu_cdac_8bit_array_2.drv<63:0>.n144 hgu_cdac_8bit_array_2.drv<63:0>.n143 0.0557941
R7672 hgu_cdac_8bit_array_2.drv<63:0>.n143 hgu_cdac_8bit_array_2.drv<63:0>.n142 0.0557941
R7673 hgu_cdac_8bit_array_2.drv<63:0>.n142 hgu_cdac_8bit_array_2.drv<63:0>.n141 0.0557941
R7674 hgu_cdac_8bit_array_2.drv<63:0>.n141 hgu_cdac_8bit_array_2.drv<63:0>.n140 0.0557941
R7675 hgu_cdac_8bit_array_2.drv<63:0>.n140 hgu_cdac_8bit_array_2.drv<63:0>.n139 0.0557941
R7676 hgu_cdac_8bit_array_2.drv<63:0>.n157 hgu_cdac_8bit_array_2.drv<63:0>.n156 0.0557941
R7677 hgu_cdac_8bit_array_2.drv<63:0>.n156 hgu_cdac_8bit_array_2.drv<63:0>.n155 0.0557941
R7678 hgu_cdac_8bit_array_2.drv<63:0>.n155 hgu_cdac_8bit_array_2.drv<63:0>.n154 0.0557941
R7679 hgu_cdac_8bit_array_2.drv<63:0>.n154 hgu_cdac_8bit_array_2.drv<63:0>.n153 0.0557941
R7680 hgu_cdac_8bit_array_2.drv<63:0>.n153 hgu_cdac_8bit_array_2.drv<63:0>.n152 0.0557941
R7681 hgu_cdac_8bit_array_2.drv<63:0>.n175 hgu_cdac_8bit_array_2.drv<63:0>.n174 0.0557941
R7682 hgu_cdac_8bit_array_2.drv<63:0>.n174 hgu_cdac_8bit_array_2.drv<63:0>.n173 0.0557941
R7683 hgu_cdac_8bit_array_2.drv<63:0>.n173 hgu_cdac_8bit_array_2.drv<63:0>.n172 0.0557941
R7684 hgu_cdac_8bit_array_2.drv<63:0>.n172 hgu_cdac_8bit_array_2.drv<63:0>.n171 0.0557941
R7685 hgu_cdac_8bit_array_2.drv<63:0>.n171 hgu_cdac_8bit_array_2.drv<63:0>.n170 0.0557941
R7686 hgu_cdac_8bit_array_2.drv<63:0>.n187 hgu_cdac_8bit_array_2.drv<63:0>.n186 0.0557941
R7687 hgu_cdac_8bit_array_2.drv<63:0>.n186 hgu_cdac_8bit_array_2.drv<63:0>.n185 0.0557941
R7688 hgu_cdac_8bit_array_2.drv<63:0>.n185 hgu_cdac_8bit_array_2.drv<63:0>.n184 0.0557941
R7689 hgu_cdac_8bit_array_2.drv<63:0>.n184 hgu_cdac_8bit_array_2.drv<63:0>.n183 0.0557941
R7690 hgu_cdac_8bit_array_2.drv<63:0>.n183 hgu_cdac_8bit_array_2.drv<63:0>.n182 0.0557941
R7691 hgu_cdac_8bit_array_2.drv<63:0>.n205 hgu_cdac_8bit_array_2.drv<63:0>.n204 0.0557941
R7692 hgu_cdac_8bit_array_2.drv<63:0>.n204 hgu_cdac_8bit_array_2.drv<63:0>.n203 0.0557941
R7693 hgu_cdac_8bit_array_2.drv<63:0>.n203 hgu_cdac_8bit_array_2.drv<63:0>.n202 0.0557941
R7694 hgu_cdac_8bit_array_2.drv<63:0>.n202 hgu_cdac_8bit_array_2.drv<63:0>.n201 0.0557941
R7695 hgu_cdac_8bit_array_2.drv<63:0>.n201 hgu_cdac_8bit_array_2.drv<63:0>.n200 0.0557941
R7696 hgu_cdac_8bit_array_2.drv<63:0>.n220 hgu_cdac_8bit_array_2.drv<63:0>.n219 0.0557941
R7697 hgu_cdac_8bit_array_2.drv<63:0>.n219 hgu_cdac_8bit_array_2.drv<63:0>.n218 0.0557941
R7698 hgu_cdac_8bit_array_2.drv<63:0>.n218 hgu_cdac_8bit_array_2.drv<63:0>.n217 0.0557941
R7699 hgu_cdac_8bit_array_2.drv<63:0>.n217 hgu_cdac_8bit_array_2.drv<63:0>.n216 0.0557941
R7700 hgu_cdac_8bit_array_2.drv<63:0>.n216 hgu_cdac_8bit_array_2.drv<63:0>.n215 0.0557941
R7701 hgu_cdac_8bit_array_2.drv<63:0>.n238 hgu_cdac_8bit_array_2.drv<63:0>.n237 0.0557941
R7702 hgu_cdac_8bit_array_2.drv<63:0>.n237 hgu_cdac_8bit_array_2.drv<63:0>.n236 0.0557941
R7703 hgu_cdac_8bit_array_2.drv<63:0>.n236 hgu_cdac_8bit_array_2.drv<63:0>.n235 0.0557941
R7704 hgu_cdac_8bit_array_2.drv<63:0>.n235 hgu_cdac_8bit_array_2.drv<63:0>.n234 0.0557941
R7705 hgu_cdac_8bit_array_2.drv<63:0>.n234 hgu_cdac_8bit_array_2.drv<63:0>.n233 0.0557941
R7706 hgu_cdac_8bit_array_2.drv<63:0>.n253 hgu_cdac_8bit_array_2.drv<63:0>.n252 0.0557941
R7707 hgu_cdac_8bit_array_2.drv<63:0>.n252 hgu_cdac_8bit_array_2.drv<63:0>.n251 0.0557941
R7708 hgu_cdac_8bit_array_2.drv<63:0>.n251 hgu_cdac_8bit_array_2.drv<63:0>.n250 0.0557941
R7709 hgu_cdac_8bit_array_2.drv<63:0>.n250 hgu_cdac_8bit_array_2.drv<63:0>.n249 0.0557941
R7710 hgu_cdac_8bit_array_2.drv<63:0>.n249 hgu_cdac_8bit_array_2.drv<63:0>.n248 0.0557941
R7711 hgu_cdac_8bit_array_2.drv<63:0>.n268 hgu_cdac_8bit_array_2.drv<63:0>.n267 0.0557941
R7712 hgu_cdac_8bit_array_2.drv<63:0>.n267 hgu_cdac_8bit_array_2.drv<63:0>.n266 0.0557941
R7713 hgu_cdac_8bit_array_2.drv<63:0>.n266 hgu_cdac_8bit_array_2.drv<63:0>.n265 0.0557941
R7714 hgu_cdac_8bit_array_2.drv<63:0>.n265 hgu_cdac_8bit_array_2.drv<63:0>.n264 0.0557941
R7715 hgu_cdac_8bit_array_2.drv<63:0>.n264 hgu_cdac_8bit_array_2.drv<63:0>.n263 0.0557941
R7716 hgu_cdac_8bit_array_2.drv<63:0>.n278 hgu_cdac_8bit_array_2.drv<63:0>.n277 0.0557941
R7717 hgu_cdac_8bit_array_2.drv<63:0>.n277 hgu_cdac_8bit_array_2.drv<63:0>.n276 0.0557941
R7718 hgu_cdac_8bit_array_2.drv<63:0>.n276 hgu_cdac_8bit_array_2.drv<63:0>.n275 0.0557941
R7719 hgu_cdac_8bit_array_2.drv<63:0>.n275 hgu_cdac_8bit_array_2.drv<63:0>.n274 0.0557941
R7720 hgu_cdac_8bit_array_2.drv<63:0>.n274 hgu_cdac_8bit_array_2.drv<63:0>.n273 0.0557941
R7721 hgu_cdac_8bit_array_2.drv<63:0>.n286 hgu_cdac_8bit_array_2.drv<63:0>.n285 0.0557941
R7722 hgu_cdac_8bit_array_2.drv<63:0>.n285 hgu_cdac_8bit_array_2.drv<63:0>.n284 0.0557941
R7723 hgu_cdac_8bit_array_2.drv<63:0>.n284 hgu_cdac_8bit_array_2.drv<63:0>.n283 0.0557941
R7724 hgu_cdac_8bit_array_2.drv<63:0>.n283 hgu_cdac_8bit_array_2.drv<63:0>.n282 0.0557941
R7725 hgu_cdac_8bit_array_2.drv<63:0>.n282 hgu_cdac_8bit_array_2.drv<63:0>.n281 0.0557941
R7726 hgu_cdac_8bit_array_2.drv<63:0>.n293 hgu_cdac_8bit_array_2.drv<63:0>.n292 0.0557941
R7727 hgu_cdac_8bit_array_2.drv<63:0>.n292 hgu_cdac_8bit_array_2.drv<63:0>.n291 0.0557941
R7728 hgu_cdac_8bit_array_2.drv<63:0>.n291 hgu_cdac_8bit_array_2.drv<63:0>.n290 0.0557941
R7729 hgu_cdac_8bit_array_2.drv<63:0>.n290 hgu_cdac_8bit_array_2.drv<63:0>.n289 0.0557941
R7730 hgu_cdac_8bit_array_2.drv<63:0>.n289 hgu_cdac_8bit_array_2.drv<63:0>.n288 0.0557941
R7731 hgu_cdac_8bit_array_2.drv<63:0>.n300 hgu_cdac_8bit_array_2.drv<63:0>.n299 0.0557941
R7732 hgu_cdac_8bit_array_2.drv<63:0>.n299 hgu_cdac_8bit_array_2.drv<63:0>.n298 0.0557941
R7733 hgu_cdac_8bit_array_2.drv<63:0>.n298 hgu_cdac_8bit_array_2.drv<63:0>.n297 0.0557941
R7734 hgu_cdac_8bit_array_2.drv<63:0>.n297 hgu_cdac_8bit_array_2.drv<63:0>.n296 0.0557941
R7735 hgu_cdac_8bit_array_2.drv<63:0>.n296 hgu_cdac_8bit_array_2.drv<63:0>.n295 0.0557941
R7736 hgu_cdac_8bit_array_2.drv<63:0>.n307 hgu_cdac_8bit_array_2.drv<63:0>.n306 0.0557941
R7737 hgu_cdac_8bit_array_2.drv<63:0>.n306 hgu_cdac_8bit_array_2.drv<63:0>.n305 0.0557941
R7738 hgu_cdac_8bit_array_2.drv<63:0>.n305 hgu_cdac_8bit_array_2.drv<63:0>.n304 0.0557941
R7739 hgu_cdac_8bit_array_2.drv<63:0>.n304 hgu_cdac_8bit_array_2.drv<63:0>.n303 0.0557941
R7740 hgu_cdac_8bit_array_2.drv<63:0>.n303 hgu_cdac_8bit_array_2.drv<63:0>.n302 0.0557941
R7741 hgu_cdac_8bit_array_2.drv<63:0>.n314 hgu_cdac_8bit_array_2.drv<63:0>.n313 0.0557941
R7742 hgu_cdac_8bit_array_2.drv<63:0>.n313 hgu_cdac_8bit_array_2.drv<63:0>.n312 0.0557941
R7743 hgu_cdac_8bit_array_2.drv<63:0>.n312 hgu_cdac_8bit_array_2.drv<63:0>.n311 0.0557941
R7744 hgu_cdac_8bit_array_2.drv<63:0>.n311 hgu_cdac_8bit_array_2.drv<63:0>.n310 0.0557941
R7745 hgu_cdac_8bit_array_2.drv<63:0>.n310 hgu_cdac_8bit_array_2.drv<63:0>.n309 0.0557941
R7746 hgu_cdac_8bit_array_2.drv<63:0>.n321 hgu_cdac_8bit_array_2.drv<63:0>.n320 0.0557941
R7747 hgu_cdac_8bit_array_2.drv<63:0>.n320 hgu_cdac_8bit_array_2.drv<63:0>.n319 0.0557941
R7748 hgu_cdac_8bit_array_2.drv<63:0>.n319 hgu_cdac_8bit_array_2.drv<63:0>.n318 0.0557941
R7749 hgu_cdac_8bit_array_2.drv<63:0>.n318 hgu_cdac_8bit_array_2.drv<63:0>.n317 0.0557941
R7750 hgu_cdac_8bit_array_2.drv<63:0>.n317 hgu_cdac_8bit_array_2.drv<63:0>.n316 0.0557941
R7751 hgu_cdac_8bit_array_2.drv<63:0>.n328 hgu_cdac_8bit_array_2.drv<63:0>.n327 0.0557941
R7752 hgu_cdac_8bit_array_2.drv<63:0>.n327 hgu_cdac_8bit_array_2.drv<63:0>.n326 0.0557941
R7753 hgu_cdac_8bit_array_2.drv<63:0>.n326 hgu_cdac_8bit_array_2.drv<63:0>.n325 0.0557941
R7754 hgu_cdac_8bit_array_2.drv<63:0>.n325 hgu_cdac_8bit_array_2.drv<63:0>.n324 0.0557941
R7755 hgu_cdac_8bit_array_2.drv<63:0>.n324 hgu_cdac_8bit_array_2.drv<63:0>.n323 0.0557941
R7756 hgu_cdac_8bit_array_2.drv<63:0>.n335 hgu_cdac_8bit_array_2.drv<63:0>.n334 0.0557941
R7757 hgu_cdac_8bit_array_2.drv<63:0>.n334 hgu_cdac_8bit_array_2.drv<63:0>.n333 0.0557941
R7758 hgu_cdac_8bit_array_2.drv<63:0>.n333 hgu_cdac_8bit_array_2.drv<63:0>.n332 0.0557941
R7759 hgu_cdac_8bit_array_2.drv<63:0>.n332 hgu_cdac_8bit_array_2.drv<63:0>.n331 0.0557941
R7760 hgu_cdac_8bit_array_2.drv<63:0>.n331 hgu_cdac_8bit_array_2.drv<63:0>.n330 0.0557941
R7761 hgu_cdac_8bit_array_2.drv<63:0>.n342 hgu_cdac_8bit_array_2.drv<63:0>.n341 0.0557941
R7762 hgu_cdac_8bit_array_2.drv<63:0>.n341 hgu_cdac_8bit_array_2.drv<63:0>.n340 0.0557941
R7763 hgu_cdac_8bit_array_2.drv<63:0>.n340 hgu_cdac_8bit_array_2.drv<63:0>.n339 0.0557941
R7764 hgu_cdac_8bit_array_2.drv<63:0>.n339 hgu_cdac_8bit_array_2.drv<63:0>.n338 0.0557941
R7765 hgu_cdac_8bit_array_2.drv<63:0>.n338 hgu_cdac_8bit_array_2.drv<63:0>.n337 0.0557941
R7766 hgu_cdac_8bit_array_2.drv<63:0>.n349 hgu_cdac_8bit_array_2.drv<63:0>.n348 0.0557941
R7767 hgu_cdac_8bit_array_2.drv<63:0>.n348 hgu_cdac_8bit_array_2.drv<63:0>.n347 0.0557941
R7768 hgu_cdac_8bit_array_2.drv<63:0>.n347 hgu_cdac_8bit_array_2.drv<63:0>.n346 0.0557941
R7769 hgu_cdac_8bit_array_2.drv<63:0>.n346 hgu_cdac_8bit_array_2.drv<63:0>.n345 0.0557941
R7770 hgu_cdac_8bit_array_2.drv<63:0>.n345 hgu_cdac_8bit_array_2.drv<63:0>.n344 0.0557941
R7771 hgu_cdac_8bit_array_2.drv<63:0>.n356 hgu_cdac_8bit_array_2.drv<63:0>.n355 0.0557941
R7772 hgu_cdac_8bit_array_2.drv<63:0>.n355 hgu_cdac_8bit_array_2.drv<63:0>.n354 0.0557941
R7773 hgu_cdac_8bit_array_2.drv<63:0>.n354 hgu_cdac_8bit_array_2.drv<63:0>.n353 0.0557941
R7774 hgu_cdac_8bit_array_2.drv<63:0>.n353 hgu_cdac_8bit_array_2.drv<63:0>.n352 0.0557941
R7775 hgu_cdac_8bit_array_2.drv<63:0>.n352 hgu_cdac_8bit_array_2.drv<63:0>.n351 0.0557941
R7776 hgu_cdac_8bit_array_2.drv<63:0>.n363 hgu_cdac_8bit_array_2.drv<63:0>.n362 0.0557941
R7777 hgu_cdac_8bit_array_2.drv<63:0>.n362 hgu_cdac_8bit_array_2.drv<63:0>.n361 0.0557941
R7778 hgu_cdac_8bit_array_2.drv<63:0>.n361 hgu_cdac_8bit_array_2.drv<63:0>.n360 0.0557941
R7779 hgu_cdac_8bit_array_2.drv<63:0>.n360 hgu_cdac_8bit_array_2.drv<63:0>.n359 0.0557941
R7780 hgu_cdac_8bit_array_2.drv<63:0>.n359 hgu_cdac_8bit_array_2.drv<63:0>.n358 0.0557941
R7781 hgu_cdac_8bit_array_2.drv<63:0>.n370 hgu_cdac_8bit_array_2.drv<63:0>.n369 0.0557941
R7782 hgu_cdac_8bit_array_2.drv<63:0>.n369 hgu_cdac_8bit_array_2.drv<63:0>.n368 0.0557941
R7783 hgu_cdac_8bit_array_2.drv<63:0>.n368 hgu_cdac_8bit_array_2.drv<63:0>.n367 0.0557941
R7784 hgu_cdac_8bit_array_2.drv<63:0>.n367 hgu_cdac_8bit_array_2.drv<63:0>.n366 0.0557941
R7785 hgu_cdac_8bit_array_2.drv<63:0>.n366 hgu_cdac_8bit_array_2.drv<63:0>.n365 0.0557941
R7786 hgu_cdac_8bit_array_2.drv<63:0>.n373 hgu_cdac_8bit_array_2.drv<63:0>.n372 0.0557941
R7787 hgu_cdac_8bit_array_2.drv<63:0>.n199 hgu_cdac_8bit_array_2.drv<63:0>.n195 0.0532344
R7788 hgu_cdac_8bit_array_2.drv<63:0>.n12 hgu_cdac_8bit_array_2.drv<63:0>.n11 0.0512812
R7789 hgu_cdac_8bit_array_2.drv<63:0>.n66 hgu_cdac_8bit_array_2.drv<63:0>.n65 0.0419706
R7790 hgu_cdac_8bit_array_2.drv<63:0>.n71 hgu_cdac_8bit_array_2.drv<63:0>.n70 0.0419706
R7791 hgu_cdac_8bit_array_2.drv<63:0>.n75 hgu_cdac_8bit_array_2.drv<63:0>.n74 0.0419706
R7792 hgu_cdac_8bit_array_2.drv<63:0>.n80 hgu_cdac_8bit_array_2.drv<63:0>.n79 0.0419706
R7793 hgu_cdac_8bit_array_2.drv<63:0>.n84 hgu_cdac_8bit_array_2.drv<63:0>.n83 0.0419706
R7794 hgu_cdac_8bit_array_2.drv<63:0>.n89 hgu_cdac_8bit_array_2.drv<63:0>.n88 0.0419706
R7795 hgu_cdac_8bit_array_2.drv<63:0>.n93 hgu_cdac_8bit_array_2.drv<63:0>.n92 0.0419706
R7796 hgu_cdac_8bit_array_2.drv<63:0>.n98 hgu_cdac_8bit_array_2.drv<63:0>.n97 0.0419706
R7797 hgu_cdac_8bit_array_2.drv<63:0>.n102 hgu_cdac_8bit_array_2.drv<63:0>.n101 0.0419706
R7798 hgu_cdac_8bit_array_2.drv<63:0>.n107 hgu_cdac_8bit_array_2.drv<63:0>.n106 0.0419706
R7799 hgu_cdac_8bit_array_2.drv<63:0>.n111 hgu_cdac_8bit_array_2.drv<63:0>.n110 0.0419706
R7800 hgu_cdac_8bit_array_2.drv<63:0>.n603 hgu_cdac_8bit_array_2.drv<63:0>.n602 0.0419706
R7801 hgu_cdac_8bit_array_2.drv<63:0>.n599 hgu_cdac_8bit_array_2.drv<63:0>.n598 0.0419706
R7802 hgu_cdac_8bit_array_2.drv<63:0>.n594 hgu_cdac_8bit_array_2.drv<63:0>.n593 0.0419706
R7803 hgu_cdac_8bit_array_2.drv<63:0>.n590 hgu_cdac_8bit_array_2.drv<63:0>.n589 0.0419706
R7804 hgu_cdac_8bit_array_2.drv<63:0>.n585 hgu_cdac_8bit_array_2.drv<63:0>.n584 0.0419706
R7805 hgu_cdac_8bit_array_2.drv<63:0>.n581 hgu_cdac_8bit_array_2.drv<63:0>.n580 0.0419706
R7806 hgu_cdac_8bit_array_2.drv<63:0>.n576 hgu_cdac_8bit_array_2.drv<63:0>.n575 0.0419706
R7807 hgu_cdac_8bit_array_2.drv<63:0>.n572 hgu_cdac_8bit_array_2.drv<63:0>.n571 0.0419706
R7808 hgu_cdac_8bit_array_2.drv<63:0>.n567 hgu_cdac_8bit_array_2.drv<63:0>.n566 0.0419706
R7809 hgu_cdac_8bit_array_2.drv<63:0>.n563 hgu_cdac_8bit_array_2.drv<63:0>.n562 0.0419706
R7810 hgu_cdac_8bit_array_2.drv<63:0>.n558 hgu_cdac_8bit_array_2.drv<63:0>.n557 0.0419706
R7811 hgu_cdac_8bit_array_2.drv<63:0>.n554 hgu_cdac_8bit_array_2.drv<63:0>.n553 0.0419706
R7812 hgu_cdac_8bit_array_2.drv<63:0>.n549 hgu_cdac_8bit_array_2.drv<63:0>.n548 0.0419706
R7813 hgu_cdac_8bit_array_2.drv<63:0>.n545 hgu_cdac_8bit_array_2.drv<63:0>.n544 0.0419706
R7814 hgu_cdac_8bit_array_2.drv<63:0>.n540 hgu_cdac_8bit_array_2.drv<63:0>.n539 0.0419706
R7815 hgu_cdac_8bit_array_2.drv<63:0>.n536 hgu_cdac_8bit_array_2.drv<63:0>.n535 0.0419706
R7816 hgu_cdac_8bit_array_2.drv<63:0>.n531 hgu_cdac_8bit_array_2.drv<63:0>.n530 0.0419706
R7817 hgu_cdac_8bit_array_2.drv<63:0>.n527 hgu_cdac_8bit_array_2.drv<63:0>.n526 0.0419706
R7818 hgu_cdac_8bit_array_2.drv<63:0>.n522 hgu_cdac_8bit_array_2.drv<63:0>.n521 0.0419706
R7819 hgu_cdac_8bit_array_2.drv<63:0>.n518 hgu_cdac_8bit_array_2.drv<63:0>.n517 0.0419706
R7820 hgu_cdac_8bit_array_2.drv<63:0>.n513 hgu_cdac_8bit_array_2.drv<63:0>.n512 0.0419706
R7821 hgu_cdac_8bit_array_2.drv<63:0>.n509 hgu_cdac_8bit_array_2.drv<63:0>.n508 0.0419706
R7822 hgu_cdac_8bit_array_2.drv<63:0>.n504 hgu_cdac_8bit_array_2.drv<63:0>.n503 0.0419706
R7823 hgu_cdac_8bit_array_2.drv<63:0>.n503 hgu_cdac_8bit_array_2.drv<63:0>.n502 0.0419706
R7824 hgu_cdac_8bit_array_2.drv<63:0>.n499 hgu_cdac_8bit_array_2.drv<63:0>.n498 0.0419706
R7825 hgu_cdac_8bit_array_2.drv<63:0>.n494 hgu_cdac_8bit_array_2.drv<63:0>.n493 0.0419706
R7826 hgu_cdac_8bit_array_2.drv<63:0>.n490 hgu_cdac_8bit_array_2.drv<63:0>.n489 0.0419706
R7827 hgu_cdac_8bit_array_2.drv<63:0>.n485 hgu_cdac_8bit_array_2.drv<63:0>.n484 0.0419706
R7828 hgu_cdac_8bit_array_2.drv<63:0>.n481 hgu_cdac_8bit_array_2.drv<63:0>.n480 0.0419706
R7829 hgu_cdac_8bit_array_2.drv<63:0>.n476 hgu_cdac_8bit_array_2.drv<63:0>.n475 0.0419706
R7830 hgu_cdac_8bit_array_2.drv<63:0>.n472 hgu_cdac_8bit_array_2.drv<63:0>.n471 0.0419706
R7831 hgu_cdac_8bit_array_2.drv<63:0>.n467 hgu_cdac_8bit_array_2.drv<63:0>.n466 0.0419706
R7832 hgu_cdac_8bit_array_2.drv<63:0>.n463 hgu_cdac_8bit_array_2.drv<63:0>.n462 0.0419706
R7833 hgu_cdac_8bit_array_2.drv<63:0>.n458 hgu_cdac_8bit_array_2.drv<63:0>.n457 0.0419706
R7834 hgu_cdac_8bit_array_2.drv<63:0>.n454 hgu_cdac_8bit_array_2.drv<63:0>.n453 0.0419706
R7835 hgu_cdac_8bit_array_2.drv<63:0>.n449 hgu_cdac_8bit_array_2.drv<63:0>.n448 0.0419706
R7836 hgu_cdac_8bit_array_2.drv<63:0>.n445 hgu_cdac_8bit_array_2.drv<63:0>.n444 0.0419706
R7837 hgu_cdac_8bit_array_2.drv<63:0>.n440 hgu_cdac_8bit_array_2.drv<63:0>.n439 0.0419706
R7838 hgu_cdac_8bit_array_2.drv<63:0>.n436 hgu_cdac_8bit_array_2.drv<63:0>.n435 0.0419706
R7839 hgu_cdac_8bit_array_2.drv<63:0>.n431 hgu_cdac_8bit_array_2.drv<63:0>.n430 0.0419706
R7840 hgu_cdac_8bit_array_2.drv<63:0>.n427 hgu_cdac_8bit_array_2.drv<63:0>.n426 0.0419706
R7841 hgu_cdac_8bit_array_2.drv<63:0>.n422 hgu_cdac_8bit_array_2.drv<63:0>.n421 0.0419706
R7842 hgu_cdac_8bit_array_2.drv<63:0>.n418 hgu_cdac_8bit_array_2.drv<63:0>.n417 0.0419706
R7843 hgu_cdac_8bit_array_2.drv<63:0>.n413 hgu_cdac_8bit_array_2.drv<63:0>.n412 0.0419706
R7844 hgu_cdac_8bit_array_2.drv<63:0>.n409 hgu_cdac_8bit_array_2.drv<63:0>.n408 0.0419706
R7845 hgu_cdac_8bit_array_2.drv<63:0>.n404 hgu_cdac_8bit_array_2.drv<63:0>.n403 0.0419706
R7846 hgu_cdac_8bit_array_2.drv<63:0>.n400 hgu_cdac_8bit_array_2.drv<63:0>.n399 0.0419706
R7847 hgu_cdac_8bit_array_2.drv<63:0>.n395 hgu_cdac_8bit_array_2.drv<63:0>.n394 0.0419706
R7848 hgu_cdac_8bit_array_2.drv<63:0>.n391 hgu_cdac_8bit_array_2.drv<63:0>.n390 0.0419706
R7849 hgu_cdac_8bit_array_2.drv<63:0>.n386 hgu_cdac_8bit_array_2.drv<63:0>.n385 0.0419706
R7850 hgu_cdac_8bit_array_2.drv<63:0>.n382 hgu_cdac_8bit_array_2.drv<63:0>.n381 0.0419706
R7851 hgu_cdac_8bit_array_2.drv<63:0>.n377 hgu_cdac_8bit_array_2.drv<63:0>.n376 0.0419706
R7852 hgu_cdac_8bit_array_2.drv<63:0> hgu_cdac_8bit_array_2.drv<63:0>.n113 0.0157059
R7853 hgu_cdac_8bit_array_2.drv<63:0>.n72 hgu_cdac_8bit_array_2.drv<63:0>.n71 0.0143235
R7854 hgu_cdac_8bit_array_2.drv<63:0>.n74 hgu_cdac_8bit_array_2.drv<63:0>.n73 0.0143235
R7855 hgu_cdac_8bit_array_2.drv<63:0>.n81 hgu_cdac_8bit_array_2.drv<63:0>.n80 0.0143235
R7856 hgu_cdac_8bit_array_2.drv<63:0>.n83 hgu_cdac_8bit_array_2.drv<63:0>.n82 0.0143235
R7857 hgu_cdac_8bit_array_2.drv<63:0>.n90 hgu_cdac_8bit_array_2.drv<63:0>.n89 0.0143235
R7858 hgu_cdac_8bit_array_2.drv<63:0>.n92 hgu_cdac_8bit_array_2.drv<63:0>.n91 0.0143235
R7859 hgu_cdac_8bit_array_2.drv<63:0>.n99 hgu_cdac_8bit_array_2.drv<63:0>.n98 0.0143235
R7860 hgu_cdac_8bit_array_2.drv<63:0>.n101 hgu_cdac_8bit_array_2.drv<63:0>.n100 0.0143235
R7861 hgu_cdac_8bit_array_2.drv<63:0>.n108 hgu_cdac_8bit_array_2.drv<63:0>.n107 0.0143235
R7862 hgu_cdac_8bit_array_2.drv<63:0>.n110 hgu_cdac_8bit_array_2.drv<63:0>.n109 0.0143235
R7863 hgu_cdac_8bit_array_2.drv<63:0>.n602 hgu_cdac_8bit_array_2.drv<63:0>.n601 0.0143235
R7864 hgu_cdac_8bit_array_2.drv<63:0>.n600 hgu_cdac_8bit_array_2.drv<63:0>.n599 0.0143235
R7865 hgu_cdac_8bit_array_2.drv<63:0>.n593 hgu_cdac_8bit_array_2.drv<63:0>.n592 0.0143235
R7866 hgu_cdac_8bit_array_2.drv<63:0>.n591 hgu_cdac_8bit_array_2.drv<63:0>.n590 0.0143235
R7867 hgu_cdac_8bit_array_2.drv<63:0>.n584 hgu_cdac_8bit_array_2.drv<63:0>.n583 0.0143235
R7868 hgu_cdac_8bit_array_2.drv<63:0>.n582 hgu_cdac_8bit_array_2.drv<63:0>.n581 0.0143235
R7869 hgu_cdac_8bit_array_2.drv<63:0>.n575 hgu_cdac_8bit_array_2.drv<63:0>.n574 0.0143235
R7870 hgu_cdac_8bit_array_2.drv<63:0>.n573 hgu_cdac_8bit_array_2.drv<63:0>.n572 0.0143235
R7871 hgu_cdac_8bit_array_2.drv<63:0>.n566 hgu_cdac_8bit_array_2.drv<63:0>.n565 0.0143235
R7872 hgu_cdac_8bit_array_2.drv<63:0>.n564 hgu_cdac_8bit_array_2.drv<63:0>.n563 0.0143235
R7873 hgu_cdac_8bit_array_2.drv<63:0>.n557 hgu_cdac_8bit_array_2.drv<63:0>.n556 0.0143235
R7874 hgu_cdac_8bit_array_2.drv<63:0>.n555 hgu_cdac_8bit_array_2.drv<63:0>.n554 0.0143235
R7875 hgu_cdac_8bit_array_2.drv<63:0>.n548 hgu_cdac_8bit_array_2.drv<63:0>.n547 0.0143235
R7876 hgu_cdac_8bit_array_2.drv<63:0>.n546 hgu_cdac_8bit_array_2.drv<63:0>.n545 0.0143235
R7877 hgu_cdac_8bit_array_2.drv<63:0>.n539 hgu_cdac_8bit_array_2.drv<63:0>.n538 0.0143235
R7878 hgu_cdac_8bit_array_2.drv<63:0>.n537 hgu_cdac_8bit_array_2.drv<63:0>.n536 0.0143235
R7879 hgu_cdac_8bit_array_2.drv<63:0>.n530 hgu_cdac_8bit_array_2.drv<63:0>.n529 0.0143235
R7880 hgu_cdac_8bit_array_2.drv<63:0>.n528 hgu_cdac_8bit_array_2.drv<63:0>.n527 0.0143235
R7881 hgu_cdac_8bit_array_2.drv<63:0>.n521 hgu_cdac_8bit_array_2.drv<63:0>.n520 0.0143235
R7882 hgu_cdac_8bit_array_2.drv<63:0>.n519 hgu_cdac_8bit_array_2.drv<63:0>.n518 0.0143235
R7883 hgu_cdac_8bit_array_2.drv<63:0>.n512 hgu_cdac_8bit_array_2.drv<63:0>.n511 0.0143235
R7884 hgu_cdac_8bit_array_2.drv<63:0>.n510 hgu_cdac_8bit_array_2.drv<63:0>.n509 0.0143235
R7885 hgu_cdac_8bit_array_2.drv<63:0>.n505 hgu_cdac_8bit_array_2.drv<63:0>.n504 0.0143235
R7886 hgu_cdac_8bit_array_2.drv<63:0>.n502 hgu_cdac_8bit_array_2.drv<63:0>.n501 0.0143235
R7887 hgu_cdac_8bit_array_2.drv<63:0>.n500 hgu_cdac_8bit_array_2.drv<63:0>.n499 0.0143235
R7888 hgu_cdac_8bit_array_2.drv<63:0>.n493 hgu_cdac_8bit_array_2.drv<63:0>.n492 0.0143235
R7889 hgu_cdac_8bit_array_2.drv<63:0>.n491 hgu_cdac_8bit_array_2.drv<63:0>.n490 0.0143235
R7890 hgu_cdac_8bit_array_2.drv<63:0>.n484 hgu_cdac_8bit_array_2.drv<63:0>.n483 0.0143235
R7891 hgu_cdac_8bit_array_2.drv<63:0>.n482 hgu_cdac_8bit_array_2.drv<63:0>.n481 0.0143235
R7892 hgu_cdac_8bit_array_2.drv<63:0>.n475 hgu_cdac_8bit_array_2.drv<63:0>.n474 0.0143235
R7893 hgu_cdac_8bit_array_2.drv<63:0>.n473 hgu_cdac_8bit_array_2.drv<63:0>.n472 0.0143235
R7894 hgu_cdac_8bit_array_2.drv<63:0>.n466 hgu_cdac_8bit_array_2.drv<63:0>.n465 0.0143235
R7895 hgu_cdac_8bit_array_2.drv<63:0>.n464 hgu_cdac_8bit_array_2.drv<63:0>.n463 0.0143235
R7896 hgu_cdac_8bit_array_2.drv<63:0>.n457 hgu_cdac_8bit_array_2.drv<63:0>.n456 0.0143235
R7897 hgu_cdac_8bit_array_2.drv<63:0>.n455 hgu_cdac_8bit_array_2.drv<63:0>.n454 0.0143235
R7898 hgu_cdac_8bit_array_2.drv<63:0>.n448 hgu_cdac_8bit_array_2.drv<63:0>.n447 0.0143235
R7899 hgu_cdac_8bit_array_2.drv<63:0>.n446 hgu_cdac_8bit_array_2.drv<63:0>.n445 0.0143235
R7900 hgu_cdac_8bit_array_2.drv<63:0>.n439 hgu_cdac_8bit_array_2.drv<63:0>.n438 0.0143235
R7901 hgu_cdac_8bit_array_2.drv<63:0>.n437 hgu_cdac_8bit_array_2.drv<63:0>.n436 0.0143235
R7902 hgu_cdac_8bit_array_2.drv<63:0>.n430 hgu_cdac_8bit_array_2.drv<63:0>.n429 0.0143235
R7903 hgu_cdac_8bit_array_2.drv<63:0>.n428 hgu_cdac_8bit_array_2.drv<63:0>.n427 0.0143235
R7904 hgu_cdac_8bit_array_2.drv<63:0>.n421 hgu_cdac_8bit_array_2.drv<63:0>.n420 0.0143235
R7905 hgu_cdac_8bit_array_2.drv<63:0>.n419 hgu_cdac_8bit_array_2.drv<63:0>.n418 0.0143235
R7906 hgu_cdac_8bit_array_2.drv<63:0>.n412 hgu_cdac_8bit_array_2.drv<63:0>.n411 0.0143235
R7907 hgu_cdac_8bit_array_2.drv<63:0>.n410 hgu_cdac_8bit_array_2.drv<63:0>.n409 0.0143235
R7908 hgu_cdac_8bit_array_2.drv<63:0>.n403 hgu_cdac_8bit_array_2.drv<63:0>.n402 0.0143235
R7909 hgu_cdac_8bit_array_2.drv<63:0>.n401 hgu_cdac_8bit_array_2.drv<63:0>.n400 0.0143235
R7910 hgu_cdac_8bit_array_2.drv<63:0>.n394 hgu_cdac_8bit_array_2.drv<63:0>.n393 0.0143235
R7911 hgu_cdac_8bit_array_2.drv<63:0>.n392 hgu_cdac_8bit_array_2.drv<63:0>.n391 0.0143235
R7912 hgu_cdac_8bit_array_2.drv<63:0>.n385 hgu_cdac_8bit_array_2.drv<63:0>.n384 0.0143235
R7913 hgu_cdac_8bit_array_2.drv<63:0>.n383 hgu_cdac_8bit_array_2.drv<63:0>.n382 0.0143235
R7914 d<4>.n1 d<4>.n0 88.1376
R7915 d<4>.n2 d<4>.n1 88.1376
R7916 d<4>.n3 d<4>.n2 88.1376
R7917 d<4>.n4 d<4>.n3 88.1376
R7918 d<4>.n5 d<4>.n4 88.1376
R7919 d<4>.n6 d<4>.n5 88.1376
R7920 d<4>.n7 d<4>.n6 88.1376
R7921 d<4>.n8 d<4>.n7 88.1376
R7922 d<4>.n9 d<4>.n8 88.1376
R7923 d<4>.n10 d<4>.n9 88.1376
R7924 d<4>.n11 d<4>.n10 88.1376
R7925 d<4>.n12 d<4>.n11 88.1376
R7926 d<4>.n13 d<4>.n12 88.1376
R7927 d<4>.n14 d<4>.n13 88.1376
R7928 d<4>.n15 d<4>.n14 88.1376
R7929 d<4>.n0 d<4>.t14 69.5462
R7930 d<4>.n1 d<4>.t4 69.5462
R7931 d<4>.n2 d<4>.t0 69.5462
R7932 d<4>.n3 d<4>.t18 69.5462
R7933 d<4>.n4 d<4>.t30 69.5462
R7934 d<4>.n5 d<4>.t24 69.5462
R7935 d<4>.n6 d<4>.t20 69.5462
R7936 d<4>.n7 d<4>.t10 69.5462
R7937 d<4>.n8 d<4>.t31 69.5462
R7938 d<4>.n9 d<4>.t25 69.5462
R7939 d<4>.n10 d<4>.t22 69.5462
R7940 d<4>.n11 d<4>.t12 69.5462
R7941 d<4>.n12 d<4>.t19 69.5462
R7942 d<4>.n13 d<4>.t15 69.5462
R7943 d<4>.n14 d<4>.t6 69.5462
R7944 d<4>.n15 d<4>.t2 69.5462
R7945 d<4>.n0 d<4>.t21 59.9062
R7946 d<4>.n1 d<4>.t11 59.9062
R7947 d<4>.n2 d<4>.t8 59.9062
R7948 d<4>.n3 d<4>.t26 59.9062
R7949 d<4>.n4 d<4>.t5 59.9062
R7950 d<4>.n5 d<4>.t1 59.9062
R7951 d<4>.n6 d<4>.t28 59.9062
R7952 d<4>.n7 d<4>.t16 59.9062
R7953 d<4>.n8 d<4>.t7 59.9062
R7954 d<4>.n9 d<4>.t3 59.9062
R7955 d<4>.n10 d<4>.t29 59.9062
R7956 d<4>.n11 d<4>.t17 59.9062
R7957 d<4>.n12 d<4>.t27 59.9062
R7958 d<4>.n13 d<4>.t23 59.9062
R7959 d<4>.n14 d<4>.t13 59.9062
R7960 d<4>.n15 d<4>.t9 59.9062
R7961 d<4> d<4>.n15 24.1005
R7962 hgu_cdac_8bit_array_3.drv<15:0>.n18 hgu_cdac_8bit_array_3.drv<15:0>.t27 41.4291
R7963 hgu_cdac_8bit_array_3.drv<15:0>.n18 hgu_cdac_8bit_array_3.drv<15:0>.t19 41.4291
R7964 hgu_cdac_8bit_array_3.drv<15:0>.n103 hgu_cdac_8bit_array_3.drv<15:0>.t24 41.4291
R7965 hgu_cdac_8bit_array_3.drv<15:0>.n103 hgu_cdac_8bit_array_3.drv<15:0>.t26 41.4291
R7966 hgu_cdac_8bit_array_3.drv<15:0>.n98 hgu_cdac_8bit_array_3.drv<15:0>.t18 41.4291
R7967 hgu_cdac_8bit_array_3.drv<15:0>.n98 hgu_cdac_8bit_array_3.drv<15:0>.t20 41.4291
R7968 hgu_cdac_8bit_array_3.drv<15:0>.n19 hgu_cdac_8bit_array_3.drv<15:0>.t29 41.4291
R7969 hgu_cdac_8bit_array_3.drv<15:0>.n19 hgu_cdac_8bit_array_3.drv<15:0>.t31 41.4291
R7970 hgu_cdac_8bit_array_3.drv<15:0>.n75 hgu_cdac_8bit_array_3.drv<15:0>.t17 41.4291
R7971 hgu_cdac_8bit_array_3.drv<15:0>.n75 hgu_cdac_8bit_array_3.drv<15:0>.t23 41.4291
R7972 hgu_cdac_8bit_array_3.drv<15:0>.n78 hgu_cdac_8bit_array_3.drv<15:0>.t28 41.4291
R7973 hgu_cdac_8bit_array_3.drv<15:0>.n78 hgu_cdac_8bit_array_3.drv<15:0>.t30 41.4291
R7974 hgu_cdac_8bit_array_3.drv<15:0>.n95 hgu_cdac_8bit_array_3.drv<15:0>.t16 41.4291
R7975 hgu_cdac_8bit_array_3.drv<15:0>.n95 hgu_cdac_8bit_array_3.drv<15:0>.t22 41.4291
R7976 hgu_cdac_8bit_array_3.drv<15:0>.n14 hgu_cdac_8bit_array_3.drv<15:0>.t21 41.4291
R7977 hgu_cdac_8bit_array_3.drv<15:0>.n14 hgu_cdac_8bit_array_3.drv<15:0>.t25 41.4291
R7978 hgu_cdac_8bit_array_3.drv<15:0>.n104 hgu_cdac_8bit_array_3.drv<15:0>.t12 34.0065
R7979 hgu_cdac_8bit_array_3.drv<15:0>.n104 hgu_cdac_8bit_array_3.drv<15:0>.t14 34.0065
R7980 hgu_cdac_8bit_array_3.drv<15:0>.n99 hgu_cdac_8bit_array_3.drv<15:0>.t6 34.0065
R7981 hgu_cdac_8bit_array_3.drv<15:0>.n99 hgu_cdac_8bit_array_3.drv<15:0>.t8 34.0065
R7982 hgu_cdac_8bit_array_3.drv<15:0>.n20 hgu_cdac_8bit_array_3.drv<15:0>.t1 34.0065
R7983 hgu_cdac_8bit_array_3.drv<15:0>.n20 hgu_cdac_8bit_array_3.drv<15:0>.t3 34.0065
R7984 hgu_cdac_8bit_array_3.drv<15:0>.n76 hgu_cdac_8bit_array_3.drv<15:0>.t5 34.0065
R7985 hgu_cdac_8bit_array_3.drv<15:0>.n76 hgu_cdac_8bit_array_3.drv<15:0>.t11 34.0065
R7986 hgu_cdac_8bit_array_3.drv<15:0>.n79 hgu_cdac_8bit_array_3.drv<15:0>.t0 34.0065
R7987 hgu_cdac_8bit_array_3.drv<15:0>.n79 hgu_cdac_8bit_array_3.drv<15:0>.t2 34.0065
R7988 hgu_cdac_8bit_array_3.drv<15:0>.n96 hgu_cdac_8bit_array_3.drv<15:0>.t4 34.0065
R7989 hgu_cdac_8bit_array_3.drv<15:0>.n96 hgu_cdac_8bit_array_3.drv<15:0>.t10 34.0065
R7990 hgu_cdac_8bit_array_3.drv<15:0>.n15 hgu_cdac_8bit_array_3.drv<15:0>.t9 34.0065
R7991 hgu_cdac_8bit_array_3.drv<15:0>.n15 hgu_cdac_8bit_array_3.drv<15:0>.t13 34.0065
R7992 hgu_cdac_8bit_array_3.drv<15:0>.n22 hgu_cdac_8bit_array_3.drv<15:0>.t15 34.0065
R7993 hgu_cdac_8bit_array_3.drv<15:0>.n22 hgu_cdac_8bit_array_3.drv<15:0>.t7 34.0065
R7994 hgu_cdac_8bit_array_3.drv<15:0>.n106 hgu_cdac_8bit_array_3.drv<15:0>.n105 11.5085
R7995 hgu_cdac_8bit_array_3.drv<15:0>.n102 hgu_cdac_8bit_array_3.drv<15:0>.n101 10.6947
R7996 hgu_cdac_8bit_array_3.drv<15:0>.n89 hgu_cdac_8bit_array_3.drv<15:0>.n81 10.6943
R7997 hgu_cdac_8bit_array_3.drv<15:0>.n25 hgu_cdac_8bit_array_3.drv<15:0>.n24 10.6923
R7998 hgu_cdac_8bit_array_3.drv<15:0>.n23 hgu_cdac_8bit_array_3.drv<15:0>.n21 0.9906
R7999 hgu_cdac_8bit_array_3.drv<15:0>.n81 hgu_cdac_8bit_array_3.drv<15:0>.n80 0.752655
R8000 hgu_cdac_8bit_array_3.drv<15:0>.n24 hgu_cdac_8bit_array_3.drv<15:0>.n17 0.752655
R8001 hgu_cdac_8bit_array_3.drv<15:0>.n100 hgu_cdac_8bit_array_3.drv<15:0>.n99 0.558205
R8002 hgu_cdac_8bit_array_3.drv<15:0>.n21 hgu_cdac_8bit_array_3.drv<15:0>.n20 0.558205
R8003 hgu_cdac_8bit_array_3.drv<15:0>.n80 hgu_cdac_8bit_array_3.drv<15:0>.n79 0.558205
R8004 hgu_cdac_8bit_array_3.drv<15:0>.n97 hgu_cdac_8bit_array_3.drv<15:0>.n96 0.558205
R8005 hgu_cdac_8bit_array_3.drv<15:0>.n16 hgu_cdac_8bit_array_3.drv<15:0>.n15 0.529944
R8006 hgu_cdac_8bit_array_3.drv<15:0>.n105 hgu_cdac_8bit_array_3.drv<15:0>.n104 0.473646
R8007 hgu_cdac_8bit_array_3.drv<15:0>.n101 hgu_cdac_8bit_array_3.drv<15:0>.n97 0.455241
R8008 hgu_cdac_8bit_array_3.drv<15:0>.n77 hgu_cdac_8bit_array_3.drv<15:0>.n76 0.381734
R8009 hgu_cdac_8bit_array_3.drv<15:0>.n23 hgu_cdac_8bit_array_3.drv<15:0>.n22 0.378057
R8010 hgu_cdac_8bit_array_3.drv<15:0>.n101 hgu_cdac_8bit_array_3.drv<15:0>.n100 0.351793
R8011 hgu_cdac_8bit_array_3.drv<15:0>.n51 hgu_cdac_8bit_array_3.drv<15:0> 0.338468
R8012 hgu_cdac_8bit_array_3.drv<15:0>.n55 hgu_cdac_8bit_array_3.drv<15:0>.n50 0.330451
R8013 hgu_cdac_8bit_array_3.drv<15:0>.n60 hgu_cdac_8bit_array_3.drv<15:0>.n47 0.330451
R8014 hgu_cdac_8bit_array_3.drv<15:0>.n65 hgu_cdac_8bit_array_3.drv<15:0>.n40 0.330451
R8015 hgu_cdac_8bit_array_3.drv<15:0>.n12 hgu_cdac_8bit_array_3.drv<15:0> 0.321667
R8016 hgu_cdac_8bit_array_3.drv<15:0>.n10 hgu_cdac_8bit_array_3.drv<15:0> 0.321667
R8017 hgu_cdac_8bit_array_3.drv<15:0>.n8 hgu_cdac_8bit_array_3.drv<15:0> 0.321667
R8018 hgu_cdac_8bit_array_3.drv<15:0>.n6 hgu_cdac_8bit_array_3.drv<15:0> 0.321667
R8019 hgu_cdac_8bit_array_3.drv<15:0>.n2 hgu_cdac_8bit_array_3.drv<15:0> 0.321667
R8020 hgu_cdac_8bit_array_3.drv<15:0>.n0 hgu_cdac_8bit_array_3.drv<15:0> 0.321667
R8021 hgu_cdac_8bit_array_3.drv<15:0>.n100 hgu_cdac_8bit_array_3.drv<15:0>.n98 0.300856
R8022 hgu_cdac_8bit_array_3.drv<15:0>.n21 hgu_cdac_8bit_array_3.drv<15:0>.n19 0.300856
R8023 hgu_cdac_8bit_array_3.drv<15:0>.n80 hgu_cdac_8bit_array_3.drv<15:0>.n78 0.300856
R8024 hgu_cdac_8bit_array_3.drv<15:0>.n97 hgu_cdac_8bit_array_3.drv<15:0>.n95 0.300856
R8025 hgu_cdac_8bit_array_3.drv<15:0>.n17 hgu_cdac_8bit_array_3.drv<15:0>.n14 0.300856
R8026 hgu_cdac_8bit_array_3.drv<15:0>.n52 hgu_cdac_8bit_array_3.drv<15:0> 0.2966
R8027 hgu_cdac_8bit_array_3.drv<15:0>.n1 hgu_cdac_8bit_array_3.drv<15:0> 0.2966
R8028 hgu_cdac_8bit_array_3.drv<15:0>.n3 hgu_cdac_8bit_array_3.drv<15:0> 0.2966
R8029 hgu_cdac_8bit_array_3.drv<15:0>.n5 hgu_cdac_8bit_array_3.drv<15:0> 0.2966
R8030 hgu_cdac_8bit_array_3.drv<15:0>.n7 hgu_cdac_8bit_array_3.drv<15:0> 0.2966
R8031 hgu_cdac_8bit_array_3.drv<15:0>.n9 hgu_cdac_8bit_array_3.drv<15:0> 0.2966
R8032 hgu_cdac_8bit_array_3.drv<15:0>.n11 hgu_cdac_8bit_array_3.drv<15:0> 0.2966
R8033 hgu_cdac_8bit_array_3.drv<15:0>.n13 hgu_cdac_8bit_array_3.drv<15:0> 0.2966
R8034 hgu_cdac_8bit_array_3.drv<15:0>.n23 hgu_cdac_8bit_array_3.drv<15:0>.n18 0.245708
R8035 hgu_cdac_8bit_array_3.drv<15:0>.n105 hgu_cdac_8bit_array_3.drv<15:0>.n103 0.245708
R8036 hgu_cdac_8bit_array_3.drv<15:0>.n77 hgu_cdac_8bit_array_3.drv<15:0>.n75 0.242032
R8037 hgu_cdac_8bit_array_3.drv<15:0>.n13 hgu_cdac_8bit_array_3.drv<15:0>.n106 0.2409
R8038 hgu_cdac_8bit_array_3.drv<15:0>.n70 hgu_cdac_8bit_array_3.drv<15:0>.n33 0.182836
R8039 hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_8bit_array_3.drv<15:0>.n25 0.182836
R8040 hgu_cdac_8bit_array_3.drv<15:0>.n114 hgu_cdac_8bit_array_3.drv<15:0>.n89 0.182836
R8041 hgu_cdac_8bit_array_3.drv<15:0>.n109 hgu_cdac_8bit_array_3.drv<15:0>.n102 0.182836
R8042 hgu_cdac_8bit_array_3.drv<15:0>.n33 hgu_cdac_8bit_array_3.drv<15:0>.n32 0.149114
R8043 hgu_cdac_8bit_array_3.drv<15:0>.n89 hgu_cdac_8bit_array_3.drv<15:0>.n88 0.149114
R8044 hgu_cdac_8bit_array_3.drv<15:0>.n102 hgu_cdac_8bit_array_3.drv<15:0>.n94 0.149114
R8045 hgu_cdac_8bit_array_3.drv<15:0>.n4 hgu_cdac_8bit_array_3.drv<15:0> 0.118
R8046 hgu_cdac_8bit_array_3.drv<15:0>.n81 hgu_cdac_8bit_array_3.drv<15:0>.n77 0.0922969
R8047 hgu_cdac_8bit_array_3.drv<15:0>.n24 hgu_cdac_8bit_array_3.drv<15:0>.n23 0.0922969
R8048 hgu_cdac_8bit_array_3.drv<15:0>.n55 hgu_cdac_8bit_array_3.drv<15:0>.n54 0.0716912
R8049 hgu_cdac_8bit_array_3.drv<15:0>.n56 hgu_cdac_8bit_array_3.drv<15:0>.n55 0.0716912
R8050 hgu_cdac_8bit_array_3.drv<15:0>.n60 hgu_cdac_8bit_array_3.drv<15:0>.n59 0.0716912
R8051 hgu_cdac_8bit_array_3.drv<15:0>.n61 hgu_cdac_8bit_array_3.drv<15:0>.n60 0.0716912
R8052 hgu_cdac_8bit_array_3.drv<15:0>.n65 hgu_cdac_8bit_array_3.drv<15:0>.n64 0.0716912
R8053 hgu_cdac_8bit_array_3.drv<15:0>.n66 hgu_cdac_8bit_array_3.drv<15:0>.n65 0.0716912
R8054 hgu_cdac_8bit_array_3.drv<15:0>.n70 hgu_cdac_8bit_array_3.drv<15:0>.n69 0.0716912
R8055 hgu_cdac_8bit_array_3.drv<15:0>.n71 hgu_cdac_8bit_array_3.drv<15:0>.n70 0.0716912
R8056 hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_8bit_array_3.drv<15:0>.n74 0.0716912
R8057 hgu_cdac_8bit_array_3.drv<15:0>.n115 hgu_cdac_8bit_array_3.drv<15:0>.n114 0.0716912
R8058 hgu_cdac_8bit_array_3.drv<15:0>.n114 hgu_cdac_8bit_array_3.drv<15:0>.n113 0.0716912
R8059 hgu_cdac_8bit_array_3.drv<15:0>.n110 hgu_cdac_8bit_array_3.drv<15:0>.n109 0.0716912
R8060 hgu_cdac_8bit_array_3.drv<15:0>.n109 hgu_cdac_8bit_array_3.drv<15:0>.n108 0.0716912
R8061 hgu_cdac_8bit_array_3.drv<15:0>.n50 hgu_cdac_8bit_array_3.drv<15:0>.n49 0.0716912
R8062 hgu_cdac_8bit_array_3.drv<15:0>.n47 hgu_cdac_8bit_array_3.drv<15:0>.n46 0.0716912
R8063 hgu_cdac_8bit_array_3.drv<15:0>.n40 hgu_cdac_8bit_array_3.drv<15:0>.n39 0.0716912
R8064 hgu_cdac_8bit_array_3.drv<15:0>.n32 hgu_cdac_8bit_array_3.drv<15:0>.n31 0.0716912
R8065 hgu_cdac_8bit_array_3.drv<15:0>.n88 hgu_cdac_8bit_array_3.drv<15:0>.n87 0.0716912
R8066 hgu_cdac_8bit_array_3.drv<15:0>.n94 hgu_cdac_8bit_array_3.drv<15:0>.n93 0.0716912
R8067 hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_8bit_array_3.drv<15:0>.n118 0.0716912
R8068 hgu_cdac_8bit_array_3.drv<15:0>.n12 hgu_cdac_8bit_array_3.drv<15:0>.n13 0.0696176
R8069 hgu_cdac_8bit_array_3.drv<15:0>.n52 hgu_cdac_8bit_array_3.drv<15:0>.n51 0.0665339
R8070 hgu_cdac_8bit_array_3.drv<15:0>.n17 hgu_cdac_8bit_array_3.drv<15:0>.n16 0.063
R8071 hgu_cdac_8bit_array_3.drv<15:0>.n54 hgu_cdac_8bit_array_3.drv<15:0>.n53 0.0557941
R8072 hgu_cdac_8bit_array_3.drv<15:0>.n57 hgu_cdac_8bit_array_3.drv<15:0>.n56 0.0557941
R8073 hgu_cdac_8bit_array_3.drv<15:0>.n1 hgu_cdac_8bit_array_3.drv<15:0>.n0 0.0557941
R8074 hgu_cdac_8bit_array_3.drv<15:0>.n59 hgu_cdac_8bit_array_3.drv<15:0>.n58 0.0557941
R8075 hgu_cdac_8bit_array_3.drv<15:0>.n62 hgu_cdac_8bit_array_3.drv<15:0>.n61 0.0557941
R8076 hgu_cdac_8bit_array_3.drv<15:0>.n3 hgu_cdac_8bit_array_3.drv<15:0>.n2 0.0557941
R8077 hgu_cdac_8bit_array_3.drv<15:0>.n64 hgu_cdac_8bit_array_3.drv<15:0>.n63 0.0557941
R8078 hgu_cdac_8bit_array_3.drv<15:0>.n67 hgu_cdac_8bit_array_3.drv<15:0>.n66 0.0557941
R8079 hgu_cdac_8bit_array_3.drv<15:0>.n5 hgu_cdac_8bit_array_3.drv<15:0>.n4 0.0557941
R8080 hgu_cdac_8bit_array_3.drv<15:0>.n69 hgu_cdac_8bit_array_3.drv<15:0>.n68 0.0557941
R8081 hgu_cdac_8bit_array_3.drv<15:0>.n72 hgu_cdac_8bit_array_3.drv<15:0>.n71 0.0557941
R8082 hgu_cdac_8bit_array_3.drv<15:0>.n7 hgu_cdac_8bit_array_3.drv<15:0>.n6 0.0557941
R8083 hgu_cdac_8bit_array_3.drv<15:0>.n74 hgu_cdac_8bit_array_3.drv<15:0>.n73 0.0557941
R8084 hgu_cdac_8bit_array_3.drv<15:0>.n118 hgu_cdac_8bit_array_3.drv<15:0>.n117 0.0557941
R8085 hgu_cdac_8bit_array_3.drv<15:0>.n8 hgu_cdac_8bit_array_3.drv<15:0>.n9 0.0557941
R8086 hgu_cdac_8bit_array_3.drv<15:0>.n116 hgu_cdac_8bit_array_3.drv<15:0>.n115 0.0557941
R8087 hgu_cdac_8bit_array_3.drv<15:0>.n113 hgu_cdac_8bit_array_3.drv<15:0>.n112 0.0557941
R8088 hgu_cdac_8bit_array_3.drv<15:0>.n10 hgu_cdac_8bit_array_3.drv<15:0>.n11 0.0557941
R8089 hgu_cdac_8bit_array_3.drv<15:0>.n111 hgu_cdac_8bit_array_3.drv<15:0>.n110 0.0557941
R8090 hgu_cdac_8bit_array_3.drv<15:0>.n108 hgu_cdac_8bit_array_3.drv<15:0>.n107 0.0557941
R8091 hgu_cdac_8bit_array_3.drv<15:0>.n49 hgu_cdac_8bit_array_3.drv<15:0>.n48 0.0557941
R8092 hgu_cdac_8bit_array_3.drv<15:0>.n42 hgu_cdac_8bit_array_3.drv<15:0>.n41 0.0557941
R8093 hgu_cdac_8bit_array_3.drv<15:0>.n43 hgu_cdac_8bit_array_3.drv<15:0>.n42 0.0557941
R8094 hgu_cdac_8bit_array_3.drv<15:0>.n44 hgu_cdac_8bit_array_3.drv<15:0>.n43 0.0557941
R8095 hgu_cdac_8bit_array_3.drv<15:0>.n45 hgu_cdac_8bit_array_3.drv<15:0>.n44 0.0557941
R8096 hgu_cdac_8bit_array_3.drv<15:0>.n46 hgu_cdac_8bit_array_3.drv<15:0>.n45 0.0557941
R8097 hgu_cdac_8bit_array_3.drv<15:0>.n35 hgu_cdac_8bit_array_3.drv<15:0>.n34 0.0557941
R8098 hgu_cdac_8bit_array_3.drv<15:0>.n36 hgu_cdac_8bit_array_3.drv<15:0>.n35 0.0557941
R8099 hgu_cdac_8bit_array_3.drv<15:0>.n37 hgu_cdac_8bit_array_3.drv<15:0>.n36 0.0557941
R8100 hgu_cdac_8bit_array_3.drv<15:0>.n38 hgu_cdac_8bit_array_3.drv<15:0>.n37 0.0557941
R8101 hgu_cdac_8bit_array_3.drv<15:0>.n39 hgu_cdac_8bit_array_3.drv<15:0>.n38 0.0557941
R8102 hgu_cdac_8bit_array_3.drv<15:0>.n27 hgu_cdac_8bit_array_3.drv<15:0>.n26 0.0557941
R8103 hgu_cdac_8bit_array_3.drv<15:0>.n28 hgu_cdac_8bit_array_3.drv<15:0>.n27 0.0557941
R8104 hgu_cdac_8bit_array_3.drv<15:0>.n29 hgu_cdac_8bit_array_3.drv<15:0>.n28 0.0557941
R8105 hgu_cdac_8bit_array_3.drv<15:0>.n30 hgu_cdac_8bit_array_3.drv<15:0>.n29 0.0557941
R8106 hgu_cdac_8bit_array_3.drv<15:0>.n31 hgu_cdac_8bit_array_3.drv<15:0>.n30 0.0557941
R8107 hgu_cdac_8bit_array_3.drv<15:0>.n87 hgu_cdac_8bit_array_3.drv<15:0>.n86 0.0557941
R8108 hgu_cdac_8bit_array_3.drv<15:0>.n86 hgu_cdac_8bit_array_3.drv<15:0>.n85 0.0557941
R8109 hgu_cdac_8bit_array_3.drv<15:0>.n85 hgu_cdac_8bit_array_3.drv<15:0>.n84 0.0557941
R8110 hgu_cdac_8bit_array_3.drv<15:0>.n84 hgu_cdac_8bit_array_3.drv<15:0>.n83 0.0557941
R8111 hgu_cdac_8bit_array_3.drv<15:0>.n83 hgu_cdac_8bit_array_3.drv<15:0>.n82 0.0557941
R8112 hgu_cdac_8bit_array_3.drv<15:0>.n93 hgu_cdac_8bit_array_3.drv<15:0>.n92 0.0557941
R8113 hgu_cdac_8bit_array_3.drv<15:0>.n92 hgu_cdac_8bit_array_3.drv<15:0>.n91 0.0557941
R8114 hgu_cdac_8bit_array_3.drv<15:0>.n91 hgu_cdac_8bit_array_3.drv<15:0>.n90 0.0557941
R8115 hgu_cdac_8bit_array_3.drv<15:0>.n107 hgu_cdac_8bit_array_3.drv<15:0>.n12 0.0557941
R8116 hgu_cdac_8bit_array_3.drv<15:0>.n11 hgu_cdac_8bit_array_3.drv<15:0>.n111 0.0557941
R8117 hgu_cdac_8bit_array_3.drv<15:0>.n112 hgu_cdac_8bit_array_3.drv<15:0>.n10 0.0557941
R8118 hgu_cdac_8bit_array_3.drv<15:0>.n9 hgu_cdac_8bit_array_3.drv<15:0>.n116 0.0557941
R8119 hgu_cdac_8bit_array_3.drv<15:0>.n117 hgu_cdac_8bit_array_3.drv<15:0>.n8 0.0557941
R8120 hgu_cdac_8bit_array_3.drv<15:0>.n73 hgu_cdac_8bit_array_3.drv<15:0>.n7 0.0557941
R8121 hgu_cdac_8bit_array_3.drv<15:0>.n6 hgu_cdac_8bit_array_3.drv<15:0>.n72 0.0557941
R8122 hgu_cdac_8bit_array_3.drv<15:0>.n68 hgu_cdac_8bit_array_3.drv<15:0>.n5 0.0557941
R8123 hgu_cdac_8bit_array_3.drv<15:0>.n4 hgu_cdac_8bit_array_3.drv<15:0>.n67 0.0557941
R8124 hgu_cdac_8bit_array_3.drv<15:0>.n63 hgu_cdac_8bit_array_3.drv<15:0>.n3 0.0557941
R8125 hgu_cdac_8bit_array_3.drv<15:0>.n2 hgu_cdac_8bit_array_3.drv<15:0>.n62 0.0557941
R8126 hgu_cdac_8bit_array_3.drv<15:0>.n58 hgu_cdac_8bit_array_3.drv<15:0>.n1 0.0557941
R8127 hgu_cdac_8bit_array_3.drv<15:0>.n0 hgu_cdac_8bit_array_3.drv<15:0>.n57 0.0557941
R8128 hgu_cdac_8bit_array_3.drv<15:0>.n53 hgu_cdac_8bit_array_3.drv<15:0>.n52 0.0419706
R8129 hgu_cdac_8bit_array_3.drv<1:0>.n1 hgu_cdac_8bit_array_3.drv<1:0>.t2 41.4291
R8130 hgu_cdac_8bit_array_3.drv<1:0>.n1 hgu_cdac_8bit_array_3.drv<1:0>.t3 41.4291
R8131 hgu_cdac_8bit_array_3.drv<1:0>.n2 hgu_cdac_8bit_array_3.drv<1:0>.t1 34.0065
R8132 hgu_cdac_8bit_array_3.drv<1:0>.n2 hgu_cdac_8bit_array_3.drv<1:0>.t0 34.0065
R8133 hgu_cdac_8bit_array_3.drv<1:0>.n4 hgu_cdac_8bit_array_3.drv<1:0>.n3 10.9504
R8134 hgu_cdac_8bit_array_3.drv<1:0>.n3 hgu_cdac_8bit_array_3.drv<1:0>.n1 0.389091
R8135 hgu_cdac_8bit_array_3.drv<1:0>.n3 hgu_cdac_8bit_array_3.drv<1:0>.n2 0.337616
R8136 hgu_cdac_8bit_array_3.drv<1:0>.n0 hgu_cdac_8bit_array_3.drv<1:0> 0.2966
R8137 hgu_cdac_8bit_array_3.drv<1:0>.n0 hgu_cdac_8bit_array_3.drv<1:0>.n4 0.238934
R8138 hgu_cdac_8bit_array_3.drv<1:0> hgu_cdac_8bit_array_3.drv<1:0>.n0 0.228564
R8139 hgu_cdac_8bit_array_3.drv<1:0>.n0 hgu_cdac_8bit_array_3.drv<1:0> 0.201033
R8140 db<4>.n1 db<4>.n0 88.1376
R8141 db<4>.n2 db<4>.n1 88.1376
R8142 db<4>.n3 db<4>.n2 88.1376
R8143 db<4>.n4 db<4>.n3 88.1376
R8144 db<4>.n5 db<4>.n4 88.1376
R8145 db<4>.n6 db<4>.n5 88.1376
R8146 db<4>.n7 db<4>.n6 88.1376
R8147 db<4>.n8 db<4>.n7 88.1376
R8148 db<4>.n9 db<4>.n8 88.1376
R8149 db<4>.n10 db<4>.n9 88.1376
R8150 db<4>.n11 db<4>.n10 88.1376
R8151 db<4>.n12 db<4>.n11 88.1376
R8152 db<4>.n13 db<4>.n12 88.1376
R8153 db<4>.n14 db<4>.n13 88.1376
R8154 db<4>.n15 db<4>.n14 88.1376
R8155 db<4>.n0 db<4>.t24 69.5462
R8156 db<4>.n1 db<4>.t17 69.5462
R8157 db<4>.n2 db<4>.t2 69.5462
R8158 db<4>.n3 db<4>.t0 69.5462
R8159 db<4>.n4 db<4>.t21 69.5462
R8160 db<4>.n5 db<4>.t19 69.5462
R8161 db<4>.n6 db<4>.t4 69.5462
R8162 db<4>.n7 db<4>.t25 69.5462
R8163 db<4>.n8 db<4>.t22 69.5462
R8164 db<4>.n9 db<4>.t8 69.5462
R8165 db<4>.n10 db<4>.t28 69.5462
R8166 db<4>.n11 db<4>.t15 69.5462
R8167 db<4>.n12 db<4>.t12 69.5462
R8168 db<4>.n13 db<4>.t9 69.5462
R8169 db<4>.n14 db<4>.t29 69.5462
R8170 db<4>.n15 db<4>.t16 69.5462
R8171 db<4>.n0 db<4>.t13 59.9062
R8172 db<4>.n1 db<4>.t6 59.9062
R8173 db<4>.n2 db<4>.t26 59.9062
R8174 db<4>.n3 db<4>.t23 59.9062
R8175 db<4>.n4 db<4>.t10 59.9062
R8176 db<4>.n5 db<4>.t7 59.9062
R8177 db<4>.n6 db<4>.t27 59.9062
R8178 db<4>.n7 db<4>.t14 59.9062
R8179 db<4>.n8 db<4>.t11 59.9062
R8180 db<4>.n9 db<4>.t30 59.9062
R8181 db<4>.n10 db<4>.t18 59.9062
R8182 db<4>.n11 db<4>.t3 59.9062
R8183 db<4>.n12 db<4>.t1 59.9062
R8184 db<4>.n13 db<4>.t31 59.9062
R8185 db<4>.n14 db<4>.t20 59.9062
R8186 db<4>.n15 db<4>.t5 59.9062
R8187 db<4> db<4>.n15 24.1005
R8188 hgu_cdac_8bit_array_2.drv<15:0>.n70 hgu_cdac_8bit_array_2.drv<15:0>.t24 41.4291
R8189 hgu_cdac_8bit_array_2.drv<15:0>.n70 hgu_cdac_8bit_array_2.drv<15:0>.t28 41.4291
R8190 hgu_cdac_8bit_array_2.drv<15:0>.n17 hgu_cdac_8bit_array_2.drv<15:0>.t21 41.4291
R8191 hgu_cdac_8bit_array_2.drv<15:0>.n17 hgu_cdac_8bit_array_2.drv<15:0>.t29 41.4291
R8192 hgu_cdac_8bit_array_2.drv<15:0>.n27 hgu_cdac_8bit_array_2.drv<15:0>.t31 41.4291
R8193 hgu_cdac_8bit_array_2.drv<15:0>.n27 hgu_cdac_8bit_array_2.drv<15:0>.t16 41.4291
R8194 hgu_cdac_8bit_array_2.drv<15:0>.n29 hgu_cdac_8bit_array_2.drv<15:0>.t22 41.4291
R8195 hgu_cdac_8bit_array_2.drv<15:0>.n29 hgu_cdac_8bit_array_2.drv<15:0>.t30 41.4291
R8196 hgu_cdac_8bit_array_2.drv<15:0>.n45 hgu_cdac_8bit_array_2.drv<15:0>.t25 41.4291
R8197 hgu_cdac_8bit_array_2.drv<15:0>.n45 hgu_cdac_8bit_array_2.drv<15:0>.t17 41.4291
R8198 hgu_cdac_8bit_array_2.drv<15:0>.n42 hgu_cdac_8bit_array_2.drv<15:0>.t18 41.4291
R8199 hgu_cdac_8bit_array_2.drv<15:0>.n42 hgu_cdac_8bit_array_2.drv<15:0>.t23 41.4291
R8200 hgu_cdac_8bit_array_2.drv<15:0>.n60 hgu_cdac_8bit_array_2.drv<15:0>.t26 41.4291
R8201 hgu_cdac_8bit_array_2.drv<15:0>.n60 hgu_cdac_8bit_array_2.drv<15:0>.t27 41.4291
R8202 hgu_cdac_8bit_array_2.drv<15:0>.n57 hgu_cdac_8bit_array_2.drv<15:0>.t19 41.4291
R8203 hgu_cdac_8bit_array_2.drv<15:0>.n57 hgu_cdac_8bit_array_2.drv<15:0>.t20 41.4291
R8204 hgu_cdac_8bit_array_2.drv<15:0>.n69 hgu_cdac_8bit_array_2.drv<15:0>.t3 34.0065
R8205 hgu_cdac_8bit_array_2.drv<15:0>.n69 hgu_cdac_8bit_array_2.drv<15:0>.t7 34.0065
R8206 hgu_cdac_8bit_array_2.drv<15:0>.n16 hgu_cdac_8bit_array_2.drv<15:0>.t0 34.0065
R8207 hgu_cdac_8bit_array_2.drv<15:0>.n16 hgu_cdac_8bit_array_2.drv<15:0>.t8 34.0065
R8208 hgu_cdac_8bit_array_2.drv<15:0>.n26 hgu_cdac_8bit_array_2.drv<15:0>.t10 34.0065
R8209 hgu_cdac_8bit_array_2.drv<15:0>.n26 hgu_cdac_8bit_array_2.drv<15:0>.t11 34.0065
R8210 hgu_cdac_8bit_array_2.drv<15:0>.n28 hgu_cdac_8bit_array_2.drv<15:0>.t1 34.0065
R8211 hgu_cdac_8bit_array_2.drv<15:0>.n28 hgu_cdac_8bit_array_2.drv<15:0>.t9 34.0065
R8212 hgu_cdac_8bit_array_2.drv<15:0>.n44 hgu_cdac_8bit_array_2.drv<15:0>.t4 34.0065
R8213 hgu_cdac_8bit_array_2.drv<15:0>.n44 hgu_cdac_8bit_array_2.drv<15:0>.t12 34.0065
R8214 hgu_cdac_8bit_array_2.drv<15:0>.n41 hgu_cdac_8bit_array_2.drv<15:0>.t13 34.0065
R8215 hgu_cdac_8bit_array_2.drv<15:0>.n41 hgu_cdac_8bit_array_2.drv<15:0>.t2 34.0065
R8216 hgu_cdac_8bit_array_2.drv<15:0>.n59 hgu_cdac_8bit_array_2.drv<15:0>.t5 34.0065
R8217 hgu_cdac_8bit_array_2.drv<15:0>.n59 hgu_cdac_8bit_array_2.drv<15:0>.t6 34.0065
R8218 hgu_cdac_8bit_array_2.drv<15:0>.n56 hgu_cdac_8bit_array_2.drv<15:0>.t14 34.0065
R8219 hgu_cdac_8bit_array_2.drv<15:0>.n56 hgu_cdac_8bit_array_2.drv<15:0>.t15 34.0065
R8220 hgu_cdac_8bit_array_2.drv<15:0>.n25 hgu_cdac_8bit_array_2.drv<15:0>.n15 12.8819
R8221 hgu_cdac_8bit_array_2.drv<15:0>.n71 hgu_cdac_8bit_array_2.drv<15:0>.n0 12.635
R8222 hgu_cdac_8bit_array_2.drv<15:0>.n40 hgu_cdac_8bit_array_2.drv<15:0>.n32 11.7313
R8223 hgu_cdac_8bit_array_2.drv<15:0>.n68 hgu_cdac_8bit_array_2.drv<15:0>.n62 11.7296
R8224 hgu_cdac_8bit_array_2.drv<15:0>.n55 hgu_cdac_8bit_array_2.drv<15:0>.n47 11.7296
R8225 hgu_cdac_8bit_array_2.drv<15:0>.n31 hgu_cdac_8bit_array_2.drv<15:0>.n30 0.990089
R8226 hgu_cdac_8bit_array_2.drv<15:0>.n47 hgu_cdac_8bit_array_2.drv<15:0>.n43 0.752655
R8227 hgu_cdac_8bit_array_2.drv<15:0>.n15 hgu_cdac_8bit_array_2.drv<15:0>.n16 0.561881
R8228 hgu_cdac_8bit_array_2.drv<15:0>.n30 hgu_cdac_8bit_array_2.drv<15:0>.n28 0.561881
R8229 hgu_cdac_8bit_array_2.drv<15:0>.n43 hgu_cdac_8bit_array_2.drv<15:0>.n41 0.561881
R8230 hgu_cdac_8bit_array_2.drv<15:0>.n61 hgu_cdac_8bit_array_2.drv<15:0>.n59 0.561881
R8231 hgu_cdac_8bit_array_2.drv<15:0>.n58 hgu_cdac_8bit_array_2.drv<15:0>.n56 0.561881
R8232 hgu_cdac_8bit_array_2.drv<15:0>.n0 hgu_cdac_8bit_array_2.drv<15:0>.n69 0.543499
R8233 hgu_cdac_8bit_array_2.drv<15:0>.n62 hgu_cdac_8bit_array_2.drv<15:0>.n61 0.459552
R8234 hgu_cdac_8bit_array_2.drv<15:0>.n46 hgu_cdac_8bit_array_2.drv<15:0>.n44 0.378057
R8235 hgu_cdac_8bit_array_2.drv<15:0>.n31 hgu_cdac_8bit_array_2.drv<15:0>.n26 0.374381
R8236 hgu_cdac_8bit_array_2.drv<15:0>.n62 hgu_cdac_8bit_array_2.drv<15:0>.n58 0.347483
R8237 hgu_cdac_8bit_array_2.drv<15:0>.n113 hgu_cdac_8bit_array_2.drv<15:0>.n100 0.330451
R8238 hgu_cdac_8bit_array_2.drv<15:0>.n108 hgu_cdac_8bit_array_2.drv<15:0>.n103 0.330451
R8239 hgu_cdac_8bit_array_2.drv<15:0>.n105 hgu_cdac_8bit_array_2.drv<15:0> 0.321667
R8240 hgu_cdac_8bit_array_2.drv<15:0>.n13 hgu_cdac_8bit_array_2.drv<15:0> 0.321667
R8241 hgu_cdac_8bit_array_2.drv<15:0>.n11 hgu_cdac_8bit_array_2.drv<15:0> 0.321667
R8242 hgu_cdac_8bit_array_2.drv<15:0>.n9 hgu_cdac_8bit_array_2.drv<15:0> 0.321667
R8243 hgu_cdac_8bit_array_2.drv<15:0>.n5 hgu_cdac_8bit_array_2.drv<15:0> 0.321667
R8244 hgu_cdac_8bit_array_2.drv<15:0>.n3 hgu_cdac_8bit_array_2.drv<15:0> 0.321667
R8245 hgu_cdac_8bit_array_2.drv<15:0>.n1 hgu_cdac_8bit_array_2.drv<15:0> 0.321667
R8246 hgu_cdac_8bit_array_2.drv<15:0>.n0 hgu_cdac_8bit_array_2.drv<15:0>.n70 0.315561
R8247 hgu_cdac_8bit_array_2.drv<15:0>.n104 hgu_cdac_8bit_array_2.drv<15:0> 0.313448
R8248 hgu_cdac_8bit_array_2.drv<15:0>.n30 hgu_cdac_8bit_array_2.drv<15:0>.n29 0.297179
R8249 hgu_cdac_8bit_array_2.drv<15:0>.n43 hgu_cdac_8bit_array_2.drv<15:0>.n42 0.297179
R8250 hgu_cdac_8bit_array_2.drv<15:0>.n61 hgu_cdac_8bit_array_2.drv<15:0>.n60 0.297179
R8251 hgu_cdac_8bit_array_2.drv<15:0>.n58 hgu_cdac_8bit_array_2.drv<15:0>.n57 0.297179
R8252 hgu_cdac_8bit_array_2.drv<15:0>.n15 hgu_cdac_8bit_array_2.drv<15:0>.n17 0.297179
R8253 hgu_cdac_8bit_array_2.drv<15:0>.n2 hgu_cdac_8bit_array_2.drv<15:0> 0.2966
R8254 hgu_cdac_8bit_array_2.drv<15:0>.n4 hgu_cdac_8bit_array_2.drv<15:0> 0.2966
R8255 hgu_cdac_8bit_array_2.drv<15:0>.n6 hgu_cdac_8bit_array_2.drv<15:0> 0.2966
R8256 hgu_cdac_8bit_array_2.drv<15:0>.n8 hgu_cdac_8bit_array_2.drv<15:0> 0.2966
R8257 hgu_cdac_8bit_array_2.drv<15:0>.n10 hgu_cdac_8bit_array_2.drv<15:0> 0.2966
R8258 hgu_cdac_8bit_array_2.drv<15:0>.n12 hgu_cdac_8bit_array_2.drv<15:0> 0.2966
R8259 hgu_cdac_8bit_array_2.drv<15:0>.n14 hgu_cdac_8bit_array_2.drv<15:0> 0.2966
R8260 hgu_cdac_8bit_array_2.drv<15:0>.n31 hgu_cdac_8bit_array_2.drv<15:0>.n27 0.245708
R8261 hgu_cdac_8bit_array_2.drv<15:0>.n46 hgu_cdac_8bit_array_2.drv<15:0>.n45 0.245708
R8262 hgu_cdac_8bit_array_2.drv<15:0>.n1 hgu_cdac_8bit_array_2.drv<15:0>.n71 0.241319
R8263 hgu_cdac_8bit_array_2.drv<15:0>.n74 hgu_cdac_8bit_array_2.drv<15:0>.n68 0.18292
R8264 hgu_cdac_8bit_array_2.drv<15:0>.n79 hgu_cdac_8bit_array_2.drv<15:0>.n55 0.18292
R8265 hgu_cdac_8bit_array_2.drv<15:0>.n84 hgu_cdac_8bit_array_2.drv<15:0>.n40 0.182836
R8266 hgu_cdac_8bit_array_2.drv<15:0>.n89 hgu_cdac_8bit_array_2.drv<15:0>.n25 0.182836
R8267 hgu_cdac_8bit_array_2.drv<15:0>.n68 hgu_cdac_8bit_array_2.drv<15:0>.n67 0.149226
R8268 hgu_cdac_8bit_array_2.drv<15:0>.n55 hgu_cdac_8bit_array_2.drv<15:0>.n54 0.149226
R8269 hgu_cdac_8bit_array_2.drv<15:0>.n40 hgu_cdac_8bit_array_2.drv<15:0>.n39 0.149114
R8270 hgu_cdac_8bit_array_2.drv<15:0>.n25 hgu_cdac_8bit_array_2.drv<15:0>.n24 0.149114
R8271 hgu_cdac_8bit_array_2.drv<15:0>.n7 hgu_cdac_8bit_array_2.drv<15:0> 0.118
R8272 hgu_cdac_8bit_array_2.drv<15:0>.n47 hgu_cdac_8bit_array_2.drv<15:0>.n46 0.0922969
R8273 hgu_cdac_8bit_array_2.drv<15:0>.n32 hgu_cdac_8bit_array_2.drv<15:0>.n31 0.0908846
R8274 hgu_cdac_8bit_array_2.drv<15:0>.n74 hgu_cdac_8bit_array_2.drv<15:0>.n73 0.0716912
R8275 hgu_cdac_8bit_array_2.drv<15:0>.n75 hgu_cdac_8bit_array_2.drv<15:0>.n74 0.0716912
R8276 hgu_cdac_8bit_array_2.drv<15:0>.n79 hgu_cdac_8bit_array_2.drv<15:0>.n78 0.0716912
R8277 hgu_cdac_8bit_array_2.drv<15:0>.n80 hgu_cdac_8bit_array_2.drv<15:0>.n79 0.0716912
R8278 hgu_cdac_8bit_array_2.drv<15:0>.n84 hgu_cdac_8bit_array_2.drv<15:0>.n83 0.0716912
R8279 hgu_cdac_8bit_array_2.drv<15:0>.n85 hgu_cdac_8bit_array_2.drv<15:0>.n84 0.0716912
R8280 hgu_cdac_8bit_array_2.drv<15:0>.n89 hgu_cdac_8bit_array_2.drv<15:0>.n88 0.0716912
R8281 hgu_cdac_8bit_array_2.drv<15:0>.n90 hgu_cdac_8bit_array_2.drv<15:0>.n89 0.0716912
R8282 hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_8bit_array_2.drv<15:0>.n93 0.0716912
R8283 hgu_cdac_8bit_array_2.drv<15:0>.n114 hgu_cdac_8bit_array_2.drv<15:0>.n113 0.0716912
R8284 hgu_cdac_8bit_array_2.drv<15:0>.n113 hgu_cdac_8bit_array_2.drv<15:0>.n112 0.0716912
R8285 hgu_cdac_8bit_array_2.drv<15:0>.n109 hgu_cdac_8bit_array_2.drv<15:0>.n108 0.0716912
R8286 hgu_cdac_8bit_array_2.drv<15:0>.n108 hgu_cdac_8bit_array_2.drv<15:0>.n107 0.0716912
R8287 hgu_cdac_8bit_array_2.drv<15:0>.n67 hgu_cdac_8bit_array_2.drv<15:0>.n66 0.0716912
R8288 hgu_cdac_8bit_array_2.drv<15:0>.n54 hgu_cdac_8bit_array_2.drv<15:0>.n53 0.0716912
R8289 hgu_cdac_8bit_array_2.drv<15:0>.n39 hgu_cdac_8bit_array_2.drv<15:0>.n38 0.0716912
R8290 hgu_cdac_8bit_array_2.drv<15:0>.n24 hgu_cdac_8bit_array_2.drv<15:0>.n23 0.0716912
R8291 hgu_cdac_8bit_array_2.drv<15:0>.n100 hgu_cdac_8bit_array_2.drv<15:0>.n99 0.0716912
R8292 hgu_cdac_8bit_array_2.drv<15:0>.n103 hgu_cdac_8bit_array_2.drv<15:0>.n102 0.0716912
R8293 hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_8bit_array_2.drv<15:0>.n117 0.0716912
R8294 hgu_cdac_8bit_array_2.drv<15:0>.n2 hgu_cdac_8bit_array_2.drv<15:0>.n1 0.0696176
R8295 hgu_cdac_8bit_array_2.drv<15:0>.n105 hgu_cdac_8bit_array_2.drv<15:0>.n104 0.0664894
R8296 hgu_cdac_8bit_array_2.drv<15:0>.n73 hgu_cdac_8bit_array_2.drv<15:0>.n72 0.0557941
R8297 hgu_cdac_8bit_array_2.drv<15:0>.n76 hgu_cdac_8bit_array_2.drv<15:0>.n75 0.0557941
R8298 hgu_cdac_8bit_array_2.drv<15:0>.n4 hgu_cdac_8bit_array_2.drv<15:0>.n3 0.0557941
R8299 hgu_cdac_8bit_array_2.drv<15:0>.n78 hgu_cdac_8bit_array_2.drv<15:0>.n77 0.0557941
R8300 hgu_cdac_8bit_array_2.drv<15:0>.n81 hgu_cdac_8bit_array_2.drv<15:0>.n80 0.0557941
R8301 hgu_cdac_8bit_array_2.drv<15:0>.n6 hgu_cdac_8bit_array_2.drv<15:0>.n5 0.0557941
R8302 hgu_cdac_8bit_array_2.drv<15:0>.n83 hgu_cdac_8bit_array_2.drv<15:0>.n82 0.0557941
R8303 hgu_cdac_8bit_array_2.drv<15:0>.n86 hgu_cdac_8bit_array_2.drv<15:0>.n85 0.0557941
R8304 hgu_cdac_8bit_array_2.drv<15:0>.n8 hgu_cdac_8bit_array_2.drv<15:0>.n7 0.0557941
R8305 hgu_cdac_8bit_array_2.drv<15:0>.n88 hgu_cdac_8bit_array_2.drv<15:0>.n87 0.0557941
R8306 hgu_cdac_8bit_array_2.drv<15:0>.n91 hgu_cdac_8bit_array_2.drv<15:0>.n90 0.0557941
R8307 hgu_cdac_8bit_array_2.drv<15:0>.n10 hgu_cdac_8bit_array_2.drv<15:0>.n9 0.0557941
R8308 hgu_cdac_8bit_array_2.drv<15:0>.n93 hgu_cdac_8bit_array_2.drv<15:0>.n92 0.0557941
R8309 hgu_cdac_8bit_array_2.drv<15:0>.n117 hgu_cdac_8bit_array_2.drv<15:0>.n116 0.0557941
R8310 hgu_cdac_8bit_array_2.drv<15:0>.n11 hgu_cdac_8bit_array_2.drv<15:0>.n12 0.0557941
R8311 hgu_cdac_8bit_array_2.drv<15:0>.n115 hgu_cdac_8bit_array_2.drv<15:0>.n114 0.0557941
R8312 hgu_cdac_8bit_array_2.drv<15:0>.n112 hgu_cdac_8bit_array_2.drv<15:0>.n111 0.0557941
R8313 hgu_cdac_8bit_array_2.drv<15:0>.n13 hgu_cdac_8bit_array_2.drv<15:0>.n14 0.0557941
R8314 hgu_cdac_8bit_array_2.drv<15:0>.n110 hgu_cdac_8bit_array_2.drv<15:0>.n109 0.0557941
R8315 hgu_cdac_8bit_array_2.drv<15:0>.n107 hgu_cdac_8bit_array_2.drv<15:0>.n106 0.0557941
R8316 hgu_cdac_8bit_array_2.drv<15:0>.n64 hgu_cdac_8bit_array_2.drv<15:0>.n63 0.0557941
R8317 hgu_cdac_8bit_array_2.drv<15:0>.n65 hgu_cdac_8bit_array_2.drv<15:0>.n64 0.0557941
R8318 hgu_cdac_8bit_array_2.drv<15:0>.n66 hgu_cdac_8bit_array_2.drv<15:0>.n65 0.0557941
R8319 hgu_cdac_8bit_array_2.drv<15:0>.n49 hgu_cdac_8bit_array_2.drv<15:0>.n48 0.0557941
R8320 hgu_cdac_8bit_array_2.drv<15:0>.n50 hgu_cdac_8bit_array_2.drv<15:0>.n49 0.0557941
R8321 hgu_cdac_8bit_array_2.drv<15:0>.n51 hgu_cdac_8bit_array_2.drv<15:0>.n50 0.0557941
R8322 hgu_cdac_8bit_array_2.drv<15:0>.n52 hgu_cdac_8bit_array_2.drv<15:0>.n51 0.0557941
R8323 hgu_cdac_8bit_array_2.drv<15:0>.n53 hgu_cdac_8bit_array_2.drv<15:0>.n52 0.0557941
R8324 hgu_cdac_8bit_array_2.drv<15:0>.n34 hgu_cdac_8bit_array_2.drv<15:0>.n33 0.0557941
R8325 hgu_cdac_8bit_array_2.drv<15:0>.n35 hgu_cdac_8bit_array_2.drv<15:0>.n34 0.0557941
R8326 hgu_cdac_8bit_array_2.drv<15:0>.n36 hgu_cdac_8bit_array_2.drv<15:0>.n35 0.0557941
R8327 hgu_cdac_8bit_array_2.drv<15:0>.n37 hgu_cdac_8bit_array_2.drv<15:0>.n36 0.0557941
R8328 hgu_cdac_8bit_array_2.drv<15:0>.n38 hgu_cdac_8bit_array_2.drv<15:0>.n37 0.0557941
R8329 hgu_cdac_8bit_array_2.drv<15:0>.n19 hgu_cdac_8bit_array_2.drv<15:0>.n18 0.0557941
R8330 hgu_cdac_8bit_array_2.drv<15:0>.n20 hgu_cdac_8bit_array_2.drv<15:0>.n19 0.0557941
R8331 hgu_cdac_8bit_array_2.drv<15:0>.n21 hgu_cdac_8bit_array_2.drv<15:0>.n20 0.0557941
R8332 hgu_cdac_8bit_array_2.drv<15:0>.n22 hgu_cdac_8bit_array_2.drv<15:0>.n21 0.0557941
R8333 hgu_cdac_8bit_array_2.drv<15:0>.n23 hgu_cdac_8bit_array_2.drv<15:0>.n22 0.0557941
R8334 hgu_cdac_8bit_array_2.drv<15:0>.n99 hgu_cdac_8bit_array_2.drv<15:0>.n98 0.0557941
R8335 hgu_cdac_8bit_array_2.drv<15:0>.n98 hgu_cdac_8bit_array_2.drv<15:0>.n97 0.0557941
R8336 hgu_cdac_8bit_array_2.drv<15:0>.n97 hgu_cdac_8bit_array_2.drv<15:0>.n96 0.0557941
R8337 hgu_cdac_8bit_array_2.drv<15:0>.n96 hgu_cdac_8bit_array_2.drv<15:0>.n95 0.0557941
R8338 hgu_cdac_8bit_array_2.drv<15:0>.n95 hgu_cdac_8bit_array_2.drv<15:0>.n94 0.0557941
R8339 hgu_cdac_8bit_array_2.drv<15:0>.n102 hgu_cdac_8bit_array_2.drv<15:0>.n101 0.0557941
R8340 hgu_cdac_8bit_array_2.drv<15:0>.n14 hgu_cdac_8bit_array_2.drv<15:0>.n110 0.0557941
R8341 hgu_cdac_8bit_array_2.drv<15:0>.n111 hgu_cdac_8bit_array_2.drv<15:0>.n13 0.0557941
R8342 hgu_cdac_8bit_array_2.drv<15:0>.n12 hgu_cdac_8bit_array_2.drv<15:0>.n115 0.0557941
R8343 hgu_cdac_8bit_array_2.drv<15:0>.n116 hgu_cdac_8bit_array_2.drv<15:0>.n11 0.0557941
R8344 hgu_cdac_8bit_array_2.drv<15:0>.n92 hgu_cdac_8bit_array_2.drv<15:0>.n10 0.0557941
R8345 hgu_cdac_8bit_array_2.drv<15:0>.n9 hgu_cdac_8bit_array_2.drv<15:0>.n91 0.0557941
R8346 hgu_cdac_8bit_array_2.drv<15:0>.n87 hgu_cdac_8bit_array_2.drv<15:0>.n8 0.0557941
R8347 hgu_cdac_8bit_array_2.drv<15:0>.n7 hgu_cdac_8bit_array_2.drv<15:0>.n86 0.0557941
R8348 hgu_cdac_8bit_array_2.drv<15:0>.n82 hgu_cdac_8bit_array_2.drv<15:0>.n6 0.0557941
R8349 hgu_cdac_8bit_array_2.drv<15:0>.n5 hgu_cdac_8bit_array_2.drv<15:0>.n81 0.0557941
R8350 hgu_cdac_8bit_array_2.drv<15:0>.n77 hgu_cdac_8bit_array_2.drv<15:0>.n4 0.0557941
R8351 hgu_cdac_8bit_array_2.drv<15:0>.n3 hgu_cdac_8bit_array_2.drv<15:0>.n76 0.0557941
R8352 hgu_cdac_8bit_array_2.drv<15:0>.n72 hgu_cdac_8bit_array_2.drv<15:0>.n2 0.0557941
R8353 hgu_cdac_8bit_array_2.drv<15:0>.n106 hgu_cdac_8bit_array_2.drv<15:0>.n105 0.0419706
R8354 db<1>.n1 db<1>.n0 88.1376
R8355 db<1>.n1 db<1> 79.1862
R8356 db<1>.n1 db<1>.t1 69.5462
R8357 db<1>.n0 db<1>.t3 69.5462
R8358 db<1>.n0 db<1>.t2 59.9062
R8359 db<1>.n1 db<1> 30.9862
R8360 db<1> db<1>.t0 28.9205
R8361 db<1> db<1>.n1 24.1005
R8362 hgu_cdac_8bit_array_2.drv<1:0>.n0 hgu_cdac_8bit_array_2.drv<1:0>.t2 41.4291
R8363 hgu_cdac_8bit_array_2.drv<1:0>.n0 hgu_cdac_8bit_array_2.drv<1:0>.t3 41.4291
R8364 hgu_cdac_8bit_array_2.drv<1:0>.n1 hgu_cdac_8bit_array_2.drv<1:0>.t0 34.0065
R8365 hgu_cdac_8bit_array_2.drv<1:0>.n1 hgu_cdac_8bit_array_2.drv<1:0>.t1 34.0065
R8366 hgu_cdac_8bit_array_2.drv<1:0> hgu_cdac_8bit_array_2.drv<1:0>.n2 13.3608
R8367 hgu_cdac_8bit_array_2.drv<1:0>.n2 hgu_cdac_8bit_array_2.drv<1:0>.n0 0.389091
R8368 hgu_cdac_8bit_array_2.drv<1:0>.n2 hgu_cdac_8bit_array_2.drv<1:0>.n1 0.337616
R8369 db<2>.n1 db<2>.n0 88.1376
R8370 db<2>.n2 db<2>.n1 88.1376
R8371 db<2>.n3 db<2>.n2 88.1376
R8372 db<2>.n0 db<2>.t5 69.5462
R8373 db<2>.n1 db<2>.t4 69.5462
R8374 db<2>.n2 db<2>.t0 69.5462
R8375 db<2>.n3 db<2>.t6 69.5462
R8376 db<2>.n0 db<2>.t2 59.9062
R8377 db<2>.n1 db<2>.t1 59.9062
R8378 db<2>.n2 db<2>.t7 59.9062
R8379 db<2>.n3 db<2>.t3 59.9062
R8380 db<2> db<2>.n3 24.1005
R8381 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n6 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t6 41.4291
R8382 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n6 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t7 41.4291
R8383 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n8 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t4 41.4291
R8384 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n8 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t5 41.4291
R8385 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n5 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t1 34.0065
R8386 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n5 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t2 34.0065
R8387 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n7 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t3 34.0065
R8388 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n7 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t0 34.0065
R8389 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n11 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n9 12.7104
R8390 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n9 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n7 0.561881
R8391 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n4 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n5 0.543499
R8392 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n2 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT 0.321667
R8393 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n4 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n6 0.315561
R8394 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n1 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT 0.313448
R8395 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n9 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n8 0.297179
R8396 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n3 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT 0.2966
R8397 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n11 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n10 0.282934
R8398 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n4 12.7579
R8399 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n11 0.174435
R8400 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n3 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n0 0.168456
R8401 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n0 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n2 0.126985
R8402 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n3 0.124175
R8403 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n2 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n1 0.10796
R8404 db<0> db<0>.t1 148.732
R8405 db<0> db<0>.t0 28.9205
R8406 hgu_cdac_8bit_array_2.drv<0>.n0 hgu_cdac_8bit_array_2.drv<0>.t1 41.6853
R8407 hgu_cdac_8bit_array_2.drv<0>.n0 hgu_cdac_8bit_array_2.drv<0>.t0 34.4833
R8408 hgu_cdac_8bit_array_2.drv<0> hgu_cdac_8bit_array_2.drv<0>.n0 10.7727
R8409 d<2>.n1 d<2>.n0 88.1376
R8410 d<2>.n2 d<2>.n1 88.1376
R8411 d<2>.n3 d<2>.n2 88.1376
R8412 d<2>.n0 d<2>.t2 69.5462
R8413 d<2>.n1 d<2>.t7 69.5462
R8414 d<2>.n2 d<2>.t5 69.5462
R8415 d<2>.n3 d<2>.t1 69.5462
R8416 d<2>.n0 d<2>.t4 59.9062
R8417 d<2>.n1 d<2>.t0 59.9062
R8418 d<2>.n2 d<2>.t6 59.9062
R8419 d<2>.n3 d<2>.t3 59.9062
R8420 d<2> d<2>.n3 24.1005
R8421 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n5 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t5 41.4291
R8422 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n5 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t7 41.4291
R8423 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n8 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t4 41.4291
R8424 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n8 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t6 41.4291
R8425 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n6 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t2 34.0065
R8426 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n6 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t0 34.0065
R8427 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n9 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t1 34.0065
R8428 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n9 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t3 34.0065
R8429 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n11 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n10 11.6043
R8430 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n7 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n1 11.2783
R8431 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n10 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n9 0.554528
R8432 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n1 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n6 0.53362
R8433 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n1 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n5 0.359679
R8434 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n3 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT 0.321667
R8435 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n10 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n8 0.304532
R8436 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n4 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT 0.2966
R8437 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n2 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT 0.2966
R8438 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n2 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n11 0.240665
R8439 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n7 0.182836
R8440 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n4 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n0 0.168456
R8441 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n0 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n3 0.126985
R8442 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n3 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n2 0.124912
R8443 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n4 0.124069
R8444 d<0> d<0>.t1 119.124
R8445 d<0> d<0>.t0 58.5291
R8446 hgu_cdac_8bit_array_3.drv<0>.n0 hgu_cdac_8bit_array_3.drv<0>.t1 41.8324
R8447 hgu_cdac_8bit_array_3.drv<0>.n0 hgu_cdac_8bit_array_3.drv<0>.t0 34.4955
R8448 hgu_cdac_8bit_array_3.drv<0> hgu_cdac_8bit_array_3.drv<0>.n0 9.32419
R8449 tb<2>.n5 tb<2>.n4 0.243676
R8450 tb<2>.n9 tb<2>.n8 0.204769
R8451 tb<2>.n0 tb<2> 0.170237
R8452 tb<2>.n2 tb<2>.n0 0.156119
R8453 tb<2>.n14 tb<2> 0.15456
R8454 tb<2>.n7 tb<2>.n2 0.128732
R8455 tb<2>.n7 tb<2>.n6 0.124872
R8456 tb<2>.n16 tb<2>.n15 0.124872
R8457 tb<2>.n5 tb<2> 0.124715
R8458 tb<2>.n11 tb<2>.n10 0.11555
R8459 tb<2>.n10 tb<2> 0.102244
R8460 tb<2>.n15 tb<2>.n14 0.0420764
R8461 tb<2>.n6 tb<2>.n5 0.0226851
R8462 tb<2>.n12 tb<2>.n11 0.01225
R8463 tb<2>.n17 tb<2>.n16 0.0101019
R8464 tb<2>.n15 tb<2>.n13 0.00864247
R8465 tb<2>.n6 tb<2>.n3 0.00864247
R8466 tb<2>.n13 tb<2>.n12 0.00687288
R8467 tb<2>.n2 tb<2>.n1 0.00494962
R8468 tb<2> tb<2>.n17 0.0041207
R8469 tb<2>.n8 tb<2>.n7 0.00349062
R8470 tb<2>.n16 tb<2>.n9 0.00349062
R8471 t<4>.n86 t<4>.n3 3.4105
R8472 t<4>.n88 t<4>.n87 3.4105
R8473 t<4>.n25 t<4>.n22 1.7055
R8474 t<4>.n27 t<4>.n26 1.7055
R8475 t<4>.n28 t<4>.n21 1.7055
R8476 t<4>.n30 t<4>.n29 1.7055
R8477 t<4>.n31 t<4>.n20 1.7055
R8478 t<4>.n34 t<4>.n33 1.7055
R8479 t<4>.n35 t<4>.n19 1.7055
R8480 t<4>.n37 t<4>.n36 1.7055
R8481 t<4>.n38 t<4>.n18 1.7055
R8482 t<4>.n40 t<4>.n39 1.7055
R8483 t<4>.n41 t<4>.n17 1.7055
R8484 t<4>.n43 t<4>.n42 1.7055
R8485 t<4>.n45 t<4>.n16 1.7055
R8486 t<4>.n47 t<4>.n46 1.7055
R8487 t<4>.n48 t<4>.n15 1.7055
R8488 t<4>.n50 t<4>.n49 1.7055
R8489 t<4>.n51 t<4>.n14 1.7055
R8490 t<4>.n54 t<4>.n53 1.7055
R8491 t<4>.n55 t<4>.n13 1.7055
R8492 t<4>.n57 t<4>.n56 1.7055
R8493 t<4>.n58 t<4>.n12 1.7055
R8494 t<4>.n60 t<4>.n59 1.7055
R8495 t<4>.n61 t<4>.n11 1.7055
R8496 t<4>.n63 t<4>.n62 1.7055
R8497 t<4>.n65 t<4>.n10 1.7055
R8498 t<4>.n67 t<4>.n66 1.7055
R8499 t<4>.n68 t<4>.n9 1.7055
R8500 t<4>.n70 t<4>.n69 1.7055
R8501 t<4>.n71 t<4>.n8 1.7055
R8502 t<4>.n73 t<4>.n72 1.7055
R8503 t<4>.n75 t<4>.n74 1.7055
R8504 t<4>.n76 t<4>.n6 1.7055
R8505 t<4>.n78 t<4>.n77 1.7055
R8506 t<4>.n79 t<4>.n5 1.7055
R8507 t<4>.n81 t<4>.n80 1.7055
R8508 t<4>.n82 t<4>.n4 1.7055
R8509 t<4>.n85 t<4>.n84 1.7055
R8510 t<4>.n93 t<4>.n92 0.397694
R8511 t<4>.n95 t<4>.n94 0.3805
R8512 t<4>.n89 t<4>.n2 0.3805
R8513 t<4>.n180 t<4>.n179 0.3805
R8514 t<4>.n23 t<4>.n22 0.342446
R8515 t<4>.n92 t<4>.n91 0.3424
R8516 t<4>.n185 t<4>.n184 0.3424
R8517 t<4>.n23 t<4> 0.255933
R8518 t<4>.n97 t<4> 0.24623
R8519 t<4>.n24 t<4>.n23 0.207891
R8520 t<4>.n93 t<4>.n0 0.193586
R8521 t<4>.n98 t<4>.n97 0.17426
R8522 t<4>.n144 t<4>.n143 0.142882
R8523 t<4>.n150 t<4>.n149 0.142882
R8524 t<4>.n156 t<4>.n155 0.142882
R8525 t<4>.n162 t<4>.n161 0.142882
R8526 t<4>.n168 t<4>.n167 0.142882
R8527 t<4>.n174 t<4>.n173 0.142882
R8528 t<4>.n101 t<4>.n100 0.142882
R8529 t<4>.n108 t<4>.n107 0.142882
R8530 t<4>.n115 t<4>.n114 0.142882
R8531 t<4>.n122 t<4>.n121 0.142882
R8532 t<4>.n129 t<4>.n128 0.142882
R8533 t<4>.n136 t<4>.n135 0.142882
R8534 t<4>.n29 t<4>.n20 0.142882
R8535 t<4>.n41 t<4>.n40 0.142882
R8536 t<4>.n49 t<4>.n14 0.142882
R8537 t<4>.n61 t<4>.n60 0.142882
R8538 t<4>.n69 t<4>.n8 0.142882
R8539 t<4>.n80 t<4>.n79 0.142882
R8540 t<4>.n31 t<4>.n30 0.142882
R8541 t<4>.n39 t<4>.n17 0.142882
R8542 t<4>.n51 t<4>.n50 0.142882
R8543 t<4>.n59 t<4>.n11 0.142882
R8544 t<4>.n71 t<4>.n70 0.142882
R8545 t<4>.n81 t<4>.n5 0.142882
R8546 t<4>.n1 t<4>.n0 0.130613
R8547 t<4>.n90 t<4>.n0 0.125385
R8548 t<4>.n96 t<4> 0.124566
R8549 t<4>.n187 t<4>.n186 0.119792
R8550 t<4>.n83 t<4> 0.0976333
R8551 t<4>.n7 t<4> 0.0976333
R8552 t<4>.n64 t<4> 0.0976333
R8553 t<4>.n52 t<4> 0.0976333
R8554 t<4>.n44 t<4> 0.0976333
R8555 t<4>.n32 t<4> 0.0976333
R8556 t<4>.n24 t<4> 0.0976333
R8557 t<4> t<4>.n95 0.0807031
R8558 t<4>.n98 t<4> 0.0725667
R8559 t<4>.n105 t<4> 0.0725667
R8560 t<4>.n112 t<4> 0.0725667
R8561 t<4>.n119 t<4> 0.0725667
R8562 t<4>.n126 t<4> 0.0725667
R8563 t<4>.n133 t<4> 0.0725667
R8564 t<4>.n141 t<4> 0.0725667
R8565 t<4>.n143 t<4>.n142 0.0557941
R8566 t<4>.n145 t<4>.n144 0.0557941
R8567 t<4>.n146 t<4>.n145 0.0557941
R8568 t<4>.n147 t<4>.n146 0.0557941
R8569 t<4>.n148 t<4>.n147 0.0557941
R8570 t<4>.n149 t<4>.n148 0.0557941
R8571 t<4>.n151 t<4>.n150 0.0557941
R8572 t<4>.n152 t<4>.n151 0.0557941
R8573 t<4>.n153 t<4>.n152 0.0557941
R8574 t<4>.n154 t<4>.n153 0.0557941
R8575 t<4>.n155 t<4>.n154 0.0557941
R8576 t<4>.n157 t<4>.n156 0.0557941
R8577 t<4>.n158 t<4>.n157 0.0557941
R8578 t<4>.n159 t<4>.n158 0.0557941
R8579 t<4>.n160 t<4>.n159 0.0557941
R8580 t<4>.n161 t<4>.n160 0.0557941
R8581 t<4>.n163 t<4>.n162 0.0557941
R8582 t<4>.n164 t<4>.n163 0.0557941
R8583 t<4>.n165 t<4>.n164 0.0557941
R8584 t<4>.n166 t<4>.n165 0.0557941
R8585 t<4>.n167 t<4>.n166 0.0557941
R8586 t<4>.n169 t<4>.n168 0.0557941
R8587 t<4>.n170 t<4>.n169 0.0557941
R8588 t<4>.n171 t<4>.n170 0.0557941
R8589 t<4>.n172 t<4>.n171 0.0557941
R8590 t<4>.n173 t<4>.n172 0.0557941
R8591 t<4>.n175 t<4>.n174 0.0557941
R8592 t<4>.n176 t<4>.n175 0.0557941
R8593 t<4>.n100 t<4>.n99 0.0557941
R8594 t<4>.n102 t<4>.n101 0.0557941
R8595 t<4>.n103 t<4>.n102 0.0557941
R8596 t<4>.n104 t<4>.n103 0.0557941
R8597 t<4>.n107 t<4>.n106 0.0557941
R8598 t<4>.n109 t<4>.n108 0.0557941
R8599 t<4>.n110 t<4>.n109 0.0557941
R8600 t<4>.n111 t<4>.n110 0.0557941
R8601 t<4>.n114 t<4>.n113 0.0557941
R8602 t<4>.n116 t<4>.n115 0.0557941
R8603 t<4>.n117 t<4>.n116 0.0557941
R8604 t<4>.n118 t<4>.n117 0.0557941
R8605 t<4>.n121 t<4>.n120 0.0557941
R8606 t<4>.n123 t<4>.n122 0.0557941
R8607 t<4>.n124 t<4>.n123 0.0557941
R8608 t<4>.n125 t<4>.n124 0.0557941
R8609 t<4>.n128 t<4>.n127 0.0557941
R8610 t<4>.n130 t<4>.n129 0.0557941
R8611 t<4>.n131 t<4>.n130 0.0557941
R8612 t<4>.n132 t<4>.n131 0.0557941
R8613 t<4>.n135 t<4>.n134 0.0557941
R8614 t<4>.n137 t<4>.n136 0.0557941
R8615 t<4>.n138 t<4>.n137 0.0557941
R8616 t<4>.n27 t<4>.n22 0.0557941
R8617 t<4>.n28 t<4>.n27 0.0557941
R8618 t<4>.n29 t<4>.n28 0.0557941
R8619 t<4>.n34 t<4>.n20 0.0557941
R8620 t<4>.n35 t<4>.n34 0.0557941
R8621 t<4>.n36 t<4>.n35 0.0557941
R8622 t<4>.n36 t<4>.n18 0.0557941
R8623 t<4>.n40 t<4>.n18 0.0557941
R8624 t<4>.n42 t<4>.n41 0.0557941
R8625 t<4>.n42 t<4>.n16 0.0557941
R8626 t<4>.n47 t<4>.n16 0.0557941
R8627 t<4>.n48 t<4>.n47 0.0557941
R8628 t<4>.n49 t<4>.n48 0.0557941
R8629 t<4>.n54 t<4>.n14 0.0557941
R8630 t<4>.n55 t<4>.n54 0.0557941
R8631 t<4>.n56 t<4>.n55 0.0557941
R8632 t<4>.n56 t<4>.n12 0.0557941
R8633 t<4>.n60 t<4>.n12 0.0557941
R8634 t<4>.n62 t<4>.n61 0.0557941
R8635 t<4>.n62 t<4>.n10 0.0557941
R8636 t<4>.n67 t<4>.n10 0.0557941
R8637 t<4>.n68 t<4>.n67 0.0557941
R8638 t<4>.n69 t<4>.n68 0.0557941
R8639 t<4>.n73 t<4>.n8 0.0557941
R8640 t<4>.n74 t<4>.n73 0.0557941
R8641 t<4>.n74 t<4>.n6 0.0557941
R8642 t<4>.n78 t<4>.n6 0.0557941
R8643 t<4>.n79 t<4>.n78 0.0557941
R8644 t<4>.n80 t<4>.n4 0.0557941
R8645 t<4>.n85 t<4>.n4 0.0557941
R8646 t<4>.n26 t<4>.n25 0.0557941
R8647 t<4>.n26 t<4>.n21 0.0557941
R8648 t<4>.n30 t<4>.n21 0.0557941
R8649 t<4>.n33 t<4>.n31 0.0557941
R8650 t<4>.n37 t<4>.n19 0.0557941
R8651 t<4>.n38 t<4>.n37 0.0557941
R8652 t<4>.n39 t<4>.n38 0.0557941
R8653 t<4>.n43 t<4>.n17 0.0557941
R8654 t<4>.n46 t<4>.n45 0.0557941
R8655 t<4>.n46 t<4>.n15 0.0557941
R8656 t<4>.n50 t<4>.n15 0.0557941
R8657 t<4>.n53 t<4>.n51 0.0557941
R8658 t<4>.n57 t<4>.n13 0.0557941
R8659 t<4>.n58 t<4>.n57 0.0557941
R8660 t<4>.n59 t<4>.n58 0.0557941
R8661 t<4>.n63 t<4>.n11 0.0557941
R8662 t<4>.n66 t<4>.n65 0.0557941
R8663 t<4>.n66 t<4>.n9 0.0557941
R8664 t<4>.n70 t<4>.n9 0.0557941
R8665 t<4>.n72 t<4>.n71 0.0557941
R8666 t<4>.n76 t<4>.n75 0.0557941
R8667 t<4>.n77 t<4>.n76 0.0557941
R8668 t<4>.n77 t<4>.n5 0.0557941
R8669 t<4>.n82 t<4>.n81 0.0557941
R8670 t<4>.n177 t<4>.n176 0.0509559
R8671 t<4>.n139 t<4>.n138 0.0509559
R8672 t<4>.n86 t<4>.n85 0.0509559
R8673 t<4>.n84 t<4>.n3 0.0509559
R8674 t<4>.n99 t<4>.n98 0.0419706
R8675 t<4>.n106 t<4>.n105 0.0419706
R8676 t<4>.n113 t<4>.n112 0.0419706
R8677 t<4>.n120 t<4>.n119 0.0419706
R8678 t<4>.n127 t<4>.n126 0.0419706
R8679 t<4>.n134 t<4>.n133 0.0419706
R8680 t<4>.n33 t<4>.n32 0.0419706
R8681 t<4>.n44 t<4>.n43 0.0419706
R8682 t<4>.n53 t<4>.n52 0.0419706
R8683 t<4>.n64 t<4>.n63 0.0419706
R8684 t<4>.n72 t<4>.n7 0.0419706
R8685 t<4>.n83 t<4>.n82 0.0419706
R8686 t<4>.n92 t<4>.n2 0.0385147
R8687 t<4>.n185 t<4>.n183 0.0281471
R8688 t<4>.n186 t<4>.n185 0.0220232
R8689 t<4>.n179 t<4>.n178 0.0177794
R8690 t<4>.n87 t<4>.n2 0.0177794
R8691 t<4>.n182 t<4>.n181 0.0170882
R8692 t<4>.n186 t<4>.n180 0.0170118
R8693 t<4>.n105 t<4>.n104 0.0143235
R8694 t<4>.n112 t<4>.n111 0.0143235
R8695 t<4>.n119 t<4>.n118 0.0143235
R8696 t<4>.n126 t<4>.n125 0.0143235
R8697 t<4>.n133 t<4>.n132 0.0143235
R8698 t<4>.n141 t<4>.n140 0.0143235
R8699 t<4>.n25 t<4>.n24 0.0143235
R8700 t<4>.n32 t<4>.n19 0.0143235
R8701 t<4>.n45 t<4>.n44 0.0143235
R8702 t<4>.n52 t<4>.n13 0.0143235
R8703 t<4>.n65 t<4>.n64 0.0143235
R8704 t<4>.n75 t<4>.n7 0.0143235
R8705 t<4>.n84 t<4>.n83 0.0143235
R8706 t<4>.n89 t<4>.n88 0.0138432
R8707 t<4>.n183 t<4>.n182 0.0115588
R8708 t<4>.n91 t<4>.n1 0.0110482
R8709 t<4>.n188 t<4>.n187 0.0100893
R8710 t<4>.n91 t<4>.n90 0.00752478
R8711 t<4>.n90 t<4>.n89 0.006246
R8712 t<4>.n178 t<4>.n177 0.00533824
R8713 t<4>.n140 t<4>.n139 0.00533824
R8714 t<4>.n87 t<4>.n86 0.00533824
R8715 t<4>.n88 t<4>.n3 0.00533824
R8716 t<4>.n94 t<4>.n93 0.00527966
R8717 t<4>.n180 t<4>.n141 0.00395588
R8718 t<4>.n95 t<4>.n0 0.00349062
R8719 t<4>.n187 t<4>.n96 0.00349062
R8720 t<4> t<4>.n188 0.00331784
R8721 t<4>.n94 t<4>.n1 0.00208685
R8722 t<2>.n5 t<2>.n3 0.473358
R8723 t<2>.n8 t<2>.n7 0.3805
R8724 t<2>.n6 t<2>.n5 0.3424
R8725 t<2>.n5 t<2>.n4 0.243676
R8726 t<2>.n3 t<2> 0.170237
R8727 t<2>.n3 t<2>.n1 0.156119
R8728 t<2>.n14 t<2> 0.15456
R8729 t<2>.n1 t<2>.n0 0.128732
R8730 t<2>.n2 t<2>.n0 0.124872
R8731 t<2>.n16 t<2>.n15 0.124872
R8732 t<2>.n4 t<2> 0.124715
R8733 t<2>.n9 t<2> 0.120759
R8734 t<2>.n11 t<2>.n10 0.11555
R8735 t<2>.n10 t<2> 0.102244
R8736 t<2> t<2>.n8 0.0845094
R8737 t<2>.n15 t<2>.n14 0.0420764
R8738 t<2>.n4 t<2>.n2 0.0226851
R8739 t<2>.n12 t<2>.n11 0.01225
R8740 t<2>.n17 t<2>.n16 0.0101019
R8741 t<2>.n15 t<2>.n13 0.00864247
R8742 t<2>.n6 t<2>.n2 0.00864247
R8743 t<2>.n13 t<2>.n12 0.00687288
R8744 t<2>.n7 t<2>.n6 0.00687288
R8745 t<2>.n7 t<2>.n1 0.00494962
R8746 t<2> t<2>.n17 0.0041207
R8747 t<2>.n8 t<2>.n0 0.00349062
R8748 t<2>.n16 t<2>.n9 0.00349062
R8749 tb<6>.n597 tb<6>.n596 0.3805
R8750 tb<6>.n398 tb<6>.n397 0.3424
R8751 tb<6>.n407 tb<6>.n406 0.3424
R8752 tb<6>.n0 tb<6> 0.271393
R8753 tb<6>.n403 tb<6>.n402 0.204749
R8754 tb<6>.n1 tb<6>.n0 0.174213
R8755 tb<6>.n591 tb<6>.n590 0.142882
R8756 tb<6>.n585 tb<6>.n584 0.142882
R8757 tb<6>.n579 tb<6>.n578 0.142882
R8758 tb<6>.n573 tb<6>.n572 0.142882
R8759 tb<6>.n567 tb<6>.n566 0.142882
R8760 tb<6>.n561 tb<6>.n560 0.142882
R8761 tb<6>.n555 tb<6>.n554 0.142882
R8762 tb<6>.n549 tb<6>.n548 0.142882
R8763 tb<6>.n543 tb<6>.n542 0.142882
R8764 tb<6>.n537 tb<6>.n536 0.142882
R8765 tb<6>.n531 tb<6>.n530 0.142882
R8766 tb<6>.n525 tb<6>.n524 0.142882
R8767 tb<6>.n519 tb<6>.n518 0.142882
R8768 tb<6>.n513 tb<6>.n512 0.142882
R8769 tb<6>.n507 tb<6>.n506 0.142882
R8770 tb<6>.n501 tb<6>.n500 0.142882
R8771 tb<6>.n495 tb<6>.n494 0.142882
R8772 tb<6>.n489 tb<6>.n488 0.142882
R8773 tb<6>.n483 tb<6>.n482 0.142882
R8774 tb<6>.n477 tb<6>.n476 0.142882
R8775 tb<6>.n471 tb<6>.n470 0.142882
R8776 tb<6>.n465 tb<6>.n464 0.142882
R8777 tb<6>.n459 tb<6>.n458 0.142882
R8778 tb<6>.n453 tb<6>.n452 0.142882
R8779 tb<6>.n447 tb<6>.n446 0.142882
R8780 tb<6>.n441 tb<6>.n440 0.142882
R8781 tb<6>.n435 tb<6>.n434 0.142882
R8782 tb<6>.n429 tb<6>.n428 0.142882
R8783 tb<6>.n423 tb<6>.n422 0.142882
R8784 tb<6>.n417 tb<6>.n416 0.142882
R8785 tb<6>.n391 tb<6>.n390 0.142882
R8786 tb<6>.n385 tb<6>.n384 0.142882
R8787 tb<6>.n379 tb<6>.n378 0.142882
R8788 tb<6>.n373 tb<6>.n372 0.142882
R8789 tb<6>.n367 tb<6>.n366 0.142882
R8790 tb<6>.n361 tb<6>.n360 0.142882
R8791 tb<6>.n355 tb<6>.n354 0.142882
R8792 tb<6>.n349 tb<6>.n348 0.142882
R8793 tb<6>.n343 tb<6>.n342 0.142882
R8794 tb<6>.n337 tb<6>.n336 0.142882
R8795 tb<6>.n331 tb<6>.n330 0.142882
R8796 tb<6>.n325 tb<6>.n324 0.142882
R8797 tb<6>.n319 tb<6>.n318 0.142882
R8798 tb<6>.n313 tb<6>.n312 0.142882
R8799 tb<6>.n307 tb<6>.n306 0.142882
R8800 tb<6>.n301 tb<6>.n300 0.142882
R8801 tb<6>.n295 tb<6>.n294 0.142882
R8802 tb<6>.n289 tb<6>.n288 0.142882
R8803 tb<6>.n283 tb<6>.n282 0.142882
R8804 tb<6>.n277 tb<6>.n276 0.142882
R8805 tb<6>.n271 tb<6>.n270 0.142882
R8806 tb<6>.n265 tb<6>.n264 0.142882
R8807 tb<6>.n259 tb<6>.n258 0.142882
R8808 tb<6>.n253 tb<6>.n252 0.142882
R8809 tb<6>.n247 tb<6>.n246 0.142882
R8810 tb<6>.n241 tb<6>.n240 0.142882
R8811 tb<6>.n235 tb<6>.n234 0.142882
R8812 tb<6>.n229 tb<6>.n228 0.142882
R8813 tb<6>.n223 tb<6>.n222 0.142882
R8814 tb<6>.n217 tb<6>.n216 0.142882
R8815 tb<6>.n207 tb<6>.n206 0.142882
R8816 tb<6>.n200 tb<6>.n199 0.142882
R8817 tb<6>.n193 tb<6>.n192 0.142882
R8818 tb<6>.n186 tb<6>.n185 0.142882
R8819 tb<6>.n179 tb<6>.n178 0.142882
R8820 tb<6>.n172 tb<6>.n171 0.142882
R8821 tb<6>.n165 tb<6>.n164 0.142882
R8822 tb<6>.n158 tb<6>.n157 0.142882
R8823 tb<6>.n151 tb<6>.n150 0.142882
R8824 tb<6>.n144 tb<6>.n143 0.142882
R8825 tb<6>.n137 tb<6>.n136 0.142882
R8826 tb<6>.n130 tb<6>.n129 0.142882
R8827 tb<6>.n123 tb<6>.n122 0.142882
R8828 tb<6>.n116 tb<6>.n115 0.142882
R8829 tb<6>.n109 tb<6>.n108 0.142882
R8830 tb<6>.n102 tb<6>.n101 0.142882
R8831 tb<6>.n95 tb<6>.n94 0.142882
R8832 tb<6>.n88 tb<6>.n87 0.142882
R8833 tb<6>.n81 tb<6>.n80 0.142882
R8834 tb<6>.n74 tb<6>.n73 0.142882
R8835 tb<6>.n67 tb<6>.n66 0.142882
R8836 tb<6>.n60 tb<6>.n59 0.142882
R8837 tb<6>.n53 tb<6>.n52 0.142882
R8838 tb<6>.n46 tb<6>.n45 0.142882
R8839 tb<6>.n39 tb<6>.n38 0.142882
R8840 tb<6>.n32 tb<6>.n31 0.142882
R8841 tb<6>.n25 tb<6>.n24 0.142882
R8842 tb<6>.n18 tb<6>.n17 0.142882
R8843 tb<6>.n11 tb<6>.n10 0.142882
R8844 tb<6>.n4 tb<6>.n3 0.142882
R8845 tb<6>.n599 tb<6>.n405 0.127395
R8846 tb<6>.n599 tb<6>.n598 0.124744
R8847 tb<6>.n1 tb<6> 0.0976333
R8848 tb<6>.n8 tb<6> 0.0976333
R8849 tb<6>.n15 tb<6> 0.0976333
R8850 tb<6>.n22 tb<6> 0.0976333
R8851 tb<6>.n29 tb<6> 0.0976333
R8852 tb<6>.n36 tb<6> 0.0976333
R8853 tb<6>.n43 tb<6> 0.0976333
R8854 tb<6>.n50 tb<6> 0.0976333
R8855 tb<6>.n57 tb<6> 0.0976333
R8856 tb<6>.n64 tb<6> 0.0976333
R8857 tb<6>.n71 tb<6> 0.0976333
R8858 tb<6>.n78 tb<6> 0.0976333
R8859 tb<6>.n85 tb<6> 0.0976333
R8860 tb<6>.n92 tb<6> 0.0976333
R8861 tb<6>.n99 tb<6> 0.0976333
R8862 tb<6>.n106 tb<6> 0.0976333
R8863 tb<6>.n113 tb<6> 0.0976333
R8864 tb<6>.n120 tb<6> 0.0976333
R8865 tb<6>.n127 tb<6> 0.0976333
R8866 tb<6>.n134 tb<6> 0.0976333
R8867 tb<6>.n141 tb<6> 0.0976333
R8868 tb<6>.n148 tb<6> 0.0976333
R8869 tb<6>.n155 tb<6> 0.0976333
R8870 tb<6>.n162 tb<6> 0.0976333
R8871 tb<6>.n169 tb<6> 0.0976333
R8872 tb<6>.n176 tb<6> 0.0976333
R8873 tb<6>.n183 tb<6> 0.0976333
R8874 tb<6>.n190 tb<6> 0.0976333
R8875 tb<6>.n197 tb<6> 0.0976333
R8876 tb<6>.n204 tb<6> 0.0976333
R8877 tb<6>.n213 tb<6> 0.0976333
R8878 tb<6>.n401 tb<6>.n400 0.0762548
R8879 tb<6>.n409 tb<6> 0.0725667
R8880 tb<6>.n593 tb<6>.n592 0.0557941
R8881 tb<6>.n592 tb<6>.n591 0.0557941
R8882 tb<6>.n590 tb<6>.n589 0.0557941
R8883 tb<6>.n589 tb<6>.n588 0.0557941
R8884 tb<6>.n588 tb<6>.n587 0.0557941
R8885 tb<6>.n587 tb<6>.n586 0.0557941
R8886 tb<6>.n586 tb<6>.n585 0.0557941
R8887 tb<6>.n584 tb<6>.n583 0.0557941
R8888 tb<6>.n583 tb<6>.n582 0.0557941
R8889 tb<6>.n582 tb<6>.n581 0.0557941
R8890 tb<6>.n581 tb<6>.n580 0.0557941
R8891 tb<6>.n580 tb<6>.n579 0.0557941
R8892 tb<6>.n578 tb<6>.n577 0.0557941
R8893 tb<6>.n577 tb<6>.n576 0.0557941
R8894 tb<6>.n576 tb<6>.n575 0.0557941
R8895 tb<6>.n575 tb<6>.n574 0.0557941
R8896 tb<6>.n574 tb<6>.n573 0.0557941
R8897 tb<6>.n572 tb<6>.n571 0.0557941
R8898 tb<6>.n571 tb<6>.n570 0.0557941
R8899 tb<6>.n570 tb<6>.n569 0.0557941
R8900 tb<6>.n569 tb<6>.n568 0.0557941
R8901 tb<6>.n568 tb<6>.n567 0.0557941
R8902 tb<6>.n566 tb<6>.n565 0.0557941
R8903 tb<6>.n565 tb<6>.n564 0.0557941
R8904 tb<6>.n564 tb<6>.n563 0.0557941
R8905 tb<6>.n563 tb<6>.n562 0.0557941
R8906 tb<6>.n562 tb<6>.n561 0.0557941
R8907 tb<6>.n560 tb<6>.n559 0.0557941
R8908 tb<6>.n559 tb<6>.n558 0.0557941
R8909 tb<6>.n558 tb<6>.n557 0.0557941
R8910 tb<6>.n557 tb<6>.n556 0.0557941
R8911 tb<6>.n556 tb<6>.n555 0.0557941
R8912 tb<6>.n554 tb<6>.n553 0.0557941
R8913 tb<6>.n553 tb<6>.n552 0.0557941
R8914 tb<6>.n552 tb<6>.n551 0.0557941
R8915 tb<6>.n551 tb<6>.n550 0.0557941
R8916 tb<6>.n550 tb<6>.n549 0.0557941
R8917 tb<6>.n548 tb<6>.n547 0.0557941
R8918 tb<6>.n547 tb<6>.n546 0.0557941
R8919 tb<6>.n546 tb<6>.n545 0.0557941
R8920 tb<6>.n545 tb<6>.n544 0.0557941
R8921 tb<6>.n544 tb<6>.n543 0.0557941
R8922 tb<6>.n542 tb<6>.n541 0.0557941
R8923 tb<6>.n541 tb<6>.n540 0.0557941
R8924 tb<6>.n540 tb<6>.n539 0.0557941
R8925 tb<6>.n539 tb<6>.n538 0.0557941
R8926 tb<6>.n538 tb<6>.n537 0.0557941
R8927 tb<6>.n536 tb<6>.n535 0.0557941
R8928 tb<6>.n535 tb<6>.n534 0.0557941
R8929 tb<6>.n534 tb<6>.n533 0.0557941
R8930 tb<6>.n533 tb<6>.n532 0.0557941
R8931 tb<6>.n532 tb<6>.n531 0.0557941
R8932 tb<6>.n530 tb<6>.n529 0.0557941
R8933 tb<6>.n529 tb<6>.n528 0.0557941
R8934 tb<6>.n528 tb<6>.n527 0.0557941
R8935 tb<6>.n527 tb<6>.n526 0.0557941
R8936 tb<6>.n526 tb<6>.n525 0.0557941
R8937 tb<6>.n524 tb<6>.n523 0.0557941
R8938 tb<6>.n523 tb<6>.n522 0.0557941
R8939 tb<6>.n522 tb<6>.n521 0.0557941
R8940 tb<6>.n521 tb<6>.n520 0.0557941
R8941 tb<6>.n520 tb<6>.n519 0.0557941
R8942 tb<6>.n518 tb<6>.n517 0.0557941
R8943 tb<6>.n517 tb<6>.n516 0.0557941
R8944 tb<6>.n516 tb<6>.n515 0.0557941
R8945 tb<6>.n515 tb<6>.n514 0.0557941
R8946 tb<6>.n514 tb<6>.n513 0.0557941
R8947 tb<6>.n512 tb<6>.n511 0.0557941
R8948 tb<6>.n511 tb<6>.n510 0.0557941
R8949 tb<6>.n510 tb<6>.n509 0.0557941
R8950 tb<6>.n509 tb<6>.n508 0.0557941
R8951 tb<6>.n508 tb<6>.n507 0.0557941
R8952 tb<6>.n506 tb<6>.n505 0.0557941
R8953 tb<6>.n505 tb<6>.n504 0.0557941
R8954 tb<6>.n504 tb<6>.n503 0.0557941
R8955 tb<6>.n503 tb<6>.n502 0.0557941
R8956 tb<6>.n502 tb<6>.n501 0.0557941
R8957 tb<6>.n500 tb<6>.n499 0.0557941
R8958 tb<6>.n499 tb<6>.n498 0.0557941
R8959 tb<6>.n498 tb<6>.n497 0.0557941
R8960 tb<6>.n497 tb<6>.n496 0.0557941
R8961 tb<6>.n496 tb<6>.n495 0.0557941
R8962 tb<6>.n494 tb<6>.n493 0.0557941
R8963 tb<6>.n493 tb<6>.n492 0.0557941
R8964 tb<6>.n492 tb<6>.n491 0.0557941
R8965 tb<6>.n491 tb<6>.n490 0.0557941
R8966 tb<6>.n490 tb<6>.n489 0.0557941
R8967 tb<6>.n488 tb<6>.n487 0.0557941
R8968 tb<6>.n487 tb<6>.n486 0.0557941
R8969 tb<6>.n486 tb<6>.n485 0.0557941
R8970 tb<6>.n485 tb<6>.n484 0.0557941
R8971 tb<6>.n484 tb<6>.n483 0.0557941
R8972 tb<6>.n482 tb<6>.n481 0.0557941
R8973 tb<6>.n481 tb<6>.n480 0.0557941
R8974 tb<6>.n480 tb<6>.n479 0.0557941
R8975 tb<6>.n479 tb<6>.n478 0.0557941
R8976 tb<6>.n478 tb<6>.n477 0.0557941
R8977 tb<6>.n476 tb<6>.n475 0.0557941
R8978 tb<6>.n475 tb<6>.n474 0.0557941
R8979 tb<6>.n474 tb<6>.n473 0.0557941
R8980 tb<6>.n473 tb<6>.n472 0.0557941
R8981 tb<6>.n472 tb<6>.n471 0.0557941
R8982 tb<6>.n470 tb<6>.n469 0.0557941
R8983 tb<6>.n469 tb<6>.n468 0.0557941
R8984 tb<6>.n468 tb<6>.n467 0.0557941
R8985 tb<6>.n467 tb<6>.n466 0.0557941
R8986 tb<6>.n466 tb<6>.n465 0.0557941
R8987 tb<6>.n464 tb<6>.n463 0.0557941
R8988 tb<6>.n463 tb<6>.n462 0.0557941
R8989 tb<6>.n462 tb<6>.n461 0.0557941
R8990 tb<6>.n461 tb<6>.n460 0.0557941
R8991 tb<6>.n460 tb<6>.n459 0.0557941
R8992 tb<6>.n458 tb<6>.n457 0.0557941
R8993 tb<6>.n457 tb<6>.n456 0.0557941
R8994 tb<6>.n456 tb<6>.n455 0.0557941
R8995 tb<6>.n455 tb<6>.n454 0.0557941
R8996 tb<6>.n454 tb<6>.n453 0.0557941
R8997 tb<6>.n452 tb<6>.n451 0.0557941
R8998 tb<6>.n451 tb<6>.n450 0.0557941
R8999 tb<6>.n450 tb<6>.n449 0.0557941
R9000 tb<6>.n449 tb<6>.n448 0.0557941
R9001 tb<6>.n448 tb<6>.n447 0.0557941
R9002 tb<6>.n446 tb<6>.n445 0.0557941
R9003 tb<6>.n445 tb<6>.n444 0.0557941
R9004 tb<6>.n444 tb<6>.n443 0.0557941
R9005 tb<6>.n443 tb<6>.n442 0.0557941
R9006 tb<6>.n442 tb<6>.n441 0.0557941
R9007 tb<6>.n440 tb<6>.n439 0.0557941
R9008 tb<6>.n439 tb<6>.n438 0.0557941
R9009 tb<6>.n438 tb<6>.n437 0.0557941
R9010 tb<6>.n437 tb<6>.n436 0.0557941
R9011 tb<6>.n436 tb<6>.n435 0.0557941
R9012 tb<6>.n434 tb<6>.n433 0.0557941
R9013 tb<6>.n433 tb<6>.n432 0.0557941
R9014 tb<6>.n432 tb<6>.n431 0.0557941
R9015 tb<6>.n431 tb<6>.n430 0.0557941
R9016 tb<6>.n430 tb<6>.n429 0.0557941
R9017 tb<6>.n428 tb<6>.n427 0.0557941
R9018 tb<6>.n427 tb<6>.n426 0.0557941
R9019 tb<6>.n426 tb<6>.n425 0.0557941
R9020 tb<6>.n425 tb<6>.n424 0.0557941
R9021 tb<6>.n424 tb<6>.n423 0.0557941
R9022 tb<6>.n422 tb<6>.n421 0.0557941
R9023 tb<6>.n421 tb<6>.n420 0.0557941
R9024 tb<6>.n420 tb<6>.n419 0.0557941
R9025 tb<6>.n419 tb<6>.n418 0.0557941
R9026 tb<6>.n418 tb<6>.n417 0.0557941
R9027 tb<6>.n416 tb<6>.n415 0.0557941
R9028 tb<6>.n415 tb<6>.n414 0.0557941
R9029 tb<6>.n414 tb<6>.n413 0.0557941
R9030 tb<6>.n408 tb<6> 0.0557941
R9031 tb<6>.n393 tb<6>.n392 0.0557941
R9032 tb<6>.n392 tb<6>.n391 0.0557941
R9033 tb<6>.n390 tb<6>.n389 0.0557941
R9034 tb<6>.n389 tb<6>.n388 0.0557941
R9035 tb<6>.n388 tb<6>.n387 0.0557941
R9036 tb<6>.n387 tb<6>.n386 0.0557941
R9037 tb<6>.n386 tb<6>.n385 0.0557941
R9038 tb<6>.n384 tb<6>.n383 0.0557941
R9039 tb<6>.n383 tb<6>.n382 0.0557941
R9040 tb<6>.n382 tb<6>.n381 0.0557941
R9041 tb<6>.n381 tb<6>.n380 0.0557941
R9042 tb<6>.n380 tb<6>.n379 0.0557941
R9043 tb<6>.n378 tb<6>.n377 0.0557941
R9044 tb<6>.n377 tb<6>.n376 0.0557941
R9045 tb<6>.n376 tb<6>.n375 0.0557941
R9046 tb<6>.n375 tb<6>.n374 0.0557941
R9047 tb<6>.n374 tb<6>.n373 0.0557941
R9048 tb<6>.n372 tb<6>.n371 0.0557941
R9049 tb<6>.n371 tb<6>.n370 0.0557941
R9050 tb<6>.n370 tb<6>.n369 0.0557941
R9051 tb<6>.n369 tb<6>.n368 0.0557941
R9052 tb<6>.n368 tb<6>.n367 0.0557941
R9053 tb<6>.n366 tb<6>.n365 0.0557941
R9054 tb<6>.n365 tb<6>.n364 0.0557941
R9055 tb<6>.n364 tb<6>.n363 0.0557941
R9056 tb<6>.n363 tb<6>.n362 0.0557941
R9057 tb<6>.n362 tb<6>.n361 0.0557941
R9058 tb<6>.n360 tb<6>.n359 0.0557941
R9059 tb<6>.n359 tb<6>.n358 0.0557941
R9060 tb<6>.n358 tb<6>.n357 0.0557941
R9061 tb<6>.n357 tb<6>.n356 0.0557941
R9062 tb<6>.n356 tb<6>.n355 0.0557941
R9063 tb<6>.n354 tb<6>.n353 0.0557941
R9064 tb<6>.n353 tb<6>.n352 0.0557941
R9065 tb<6>.n352 tb<6>.n351 0.0557941
R9066 tb<6>.n351 tb<6>.n350 0.0557941
R9067 tb<6>.n350 tb<6>.n349 0.0557941
R9068 tb<6>.n348 tb<6>.n347 0.0557941
R9069 tb<6>.n347 tb<6>.n346 0.0557941
R9070 tb<6>.n346 tb<6>.n345 0.0557941
R9071 tb<6>.n345 tb<6>.n344 0.0557941
R9072 tb<6>.n344 tb<6>.n343 0.0557941
R9073 tb<6>.n342 tb<6>.n341 0.0557941
R9074 tb<6>.n341 tb<6>.n340 0.0557941
R9075 tb<6>.n340 tb<6>.n339 0.0557941
R9076 tb<6>.n339 tb<6>.n338 0.0557941
R9077 tb<6>.n338 tb<6>.n337 0.0557941
R9078 tb<6>.n336 tb<6>.n335 0.0557941
R9079 tb<6>.n335 tb<6>.n334 0.0557941
R9080 tb<6>.n334 tb<6>.n333 0.0557941
R9081 tb<6>.n333 tb<6>.n332 0.0557941
R9082 tb<6>.n332 tb<6>.n331 0.0557941
R9083 tb<6>.n330 tb<6>.n329 0.0557941
R9084 tb<6>.n329 tb<6>.n328 0.0557941
R9085 tb<6>.n328 tb<6>.n327 0.0557941
R9086 tb<6>.n327 tb<6>.n326 0.0557941
R9087 tb<6>.n326 tb<6>.n325 0.0557941
R9088 tb<6>.n324 tb<6>.n323 0.0557941
R9089 tb<6>.n323 tb<6>.n322 0.0557941
R9090 tb<6>.n322 tb<6>.n321 0.0557941
R9091 tb<6>.n321 tb<6>.n320 0.0557941
R9092 tb<6>.n320 tb<6>.n319 0.0557941
R9093 tb<6>.n318 tb<6>.n317 0.0557941
R9094 tb<6>.n317 tb<6>.n316 0.0557941
R9095 tb<6>.n316 tb<6>.n315 0.0557941
R9096 tb<6>.n315 tb<6>.n314 0.0557941
R9097 tb<6>.n314 tb<6>.n313 0.0557941
R9098 tb<6>.n312 tb<6>.n311 0.0557941
R9099 tb<6>.n311 tb<6>.n310 0.0557941
R9100 tb<6>.n310 tb<6>.n309 0.0557941
R9101 tb<6>.n309 tb<6>.n308 0.0557941
R9102 tb<6>.n308 tb<6>.n307 0.0557941
R9103 tb<6>.n306 tb<6>.n305 0.0557941
R9104 tb<6>.n305 tb<6>.n304 0.0557941
R9105 tb<6>.n304 tb<6>.n303 0.0557941
R9106 tb<6>.n303 tb<6>.n302 0.0557941
R9107 tb<6>.n302 tb<6>.n301 0.0557941
R9108 tb<6>.n300 tb<6>.n299 0.0557941
R9109 tb<6>.n299 tb<6>.n298 0.0557941
R9110 tb<6>.n298 tb<6>.n297 0.0557941
R9111 tb<6>.n297 tb<6>.n296 0.0557941
R9112 tb<6>.n296 tb<6>.n295 0.0557941
R9113 tb<6>.n294 tb<6>.n293 0.0557941
R9114 tb<6>.n293 tb<6>.n292 0.0557941
R9115 tb<6>.n292 tb<6>.n291 0.0557941
R9116 tb<6>.n291 tb<6>.n290 0.0557941
R9117 tb<6>.n290 tb<6>.n289 0.0557941
R9118 tb<6>.n288 tb<6>.n287 0.0557941
R9119 tb<6>.n287 tb<6>.n286 0.0557941
R9120 tb<6>.n286 tb<6>.n285 0.0557941
R9121 tb<6>.n285 tb<6>.n284 0.0557941
R9122 tb<6>.n284 tb<6>.n283 0.0557941
R9123 tb<6>.n282 tb<6>.n281 0.0557941
R9124 tb<6>.n281 tb<6>.n280 0.0557941
R9125 tb<6>.n280 tb<6>.n279 0.0557941
R9126 tb<6>.n279 tb<6>.n278 0.0557941
R9127 tb<6>.n278 tb<6>.n277 0.0557941
R9128 tb<6>.n276 tb<6>.n275 0.0557941
R9129 tb<6>.n275 tb<6>.n274 0.0557941
R9130 tb<6>.n274 tb<6>.n273 0.0557941
R9131 tb<6>.n273 tb<6>.n272 0.0557941
R9132 tb<6>.n272 tb<6>.n271 0.0557941
R9133 tb<6>.n270 tb<6>.n269 0.0557941
R9134 tb<6>.n269 tb<6>.n268 0.0557941
R9135 tb<6>.n268 tb<6>.n267 0.0557941
R9136 tb<6>.n267 tb<6>.n266 0.0557941
R9137 tb<6>.n266 tb<6>.n265 0.0557941
R9138 tb<6>.n264 tb<6>.n263 0.0557941
R9139 tb<6>.n263 tb<6>.n262 0.0557941
R9140 tb<6>.n262 tb<6>.n261 0.0557941
R9141 tb<6>.n261 tb<6>.n260 0.0557941
R9142 tb<6>.n260 tb<6>.n259 0.0557941
R9143 tb<6>.n258 tb<6>.n257 0.0557941
R9144 tb<6>.n257 tb<6>.n256 0.0557941
R9145 tb<6>.n256 tb<6>.n255 0.0557941
R9146 tb<6>.n255 tb<6>.n254 0.0557941
R9147 tb<6>.n254 tb<6>.n253 0.0557941
R9148 tb<6>.n252 tb<6>.n251 0.0557941
R9149 tb<6>.n251 tb<6>.n250 0.0557941
R9150 tb<6>.n250 tb<6>.n249 0.0557941
R9151 tb<6>.n249 tb<6>.n248 0.0557941
R9152 tb<6>.n248 tb<6>.n247 0.0557941
R9153 tb<6>.n246 tb<6>.n245 0.0557941
R9154 tb<6>.n245 tb<6>.n244 0.0557941
R9155 tb<6>.n244 tb<6>.n243 0.0557941
R9156 tb<6>.n243 tb<6>.n242 0.0557941
R9157 tb<6>.n242 tb<6>.n241 0.0557941
R9158 tb<6>.n240 tb<6>.n239 0.0557941
R9159 tb<6>.n239 tb<6>.n238 0.0557941
R9160 tb<6>.n238 tb<6>.n237 0.0557941
R9161 tb<6>.n237 tb<6>.n236 0.0557941
R9162 tb<6>.n236 tb<6>.n235 0.0557941
R9163 tb<6>.n234 tb<6>.n233 0.0557941
R9164 tb<6>.n233 tb<6>.n232 0.0557941
R9165 tb<6>.n232 tb<6>.n231 0.0557941
R9166 tb<6>.n231 tb<6>.n230 0.0557941
R9167 tb<6>.n230 tb<6>.n229 0.0557941
R9168 tb<6>.n228 tb<6>.n227 0.0557941
R9169 tb<6>.n227 tb<6>.n226 0.0557941
R9170 tb<6>.n226 tb<6>.n225 0.0557941
R9171 tb<6>.n225 tb<6>.n224 0.0557941
R9172 tb<6>.n224 tb<6>.n223 0.0557941
R9173 tb<6>.n222 tb<6>.n221 0.0557941
R9174 tb<6>.n221 tb<6>.n220 0.0557941
R9175 tb<6>.n220 tb<6>.n219 0.0557941
R9176 tb<6>.n219 tb<6>.n218 0.0557941
R9177 tb<6>.n218 tb<6>.n217 0.0557941
R9178 tb<6>.n216 tb<6>.n215 0.0557941
R9179 tb<6>.n209 tb<6>.n208 0.0557941
R9180 tb<6>.n208 tb<6>.n207 0.0557941
R9181 tb<6>.n206 tb<6>.n205 0.0557941
R9182 tb<6>.n203 tb<6>.n202 0.0557941
R9183 tb<6>.n202 tb<6>.n201 0.0557941
R9184 tb<6>.n201 tb<6>.n200 0.0557941
R9185 tb<6>.n199 tb<6>.n198 0.0557941
R9186 tb<6>.n196 tb<6>.n195 0.0557941
R9187 tb<6>.n195 tb<6>.n194 0.0557941
R9188 tb<6>.n194 tb<6>.n193 0.0557941
R9189 tb<6>.n192 tb<6>.n191 0.0557941
R9190 tb<6>.n189 tb<6>.n188 0.0557941
R9191 tb<6>.n188 tb<6>.n187 0.0557941
R9192 tb<6>.n187 tb<6>.n186 0.0557941
R9193 tb<6>.n185 tb<6>.n184 0.0557941
R9194 tb<6>.n182 tb<6>.n181 0.0557941
R9195 tb<6>.n181 tb<6>.n180 0.0557941
R9196 tb<6>.n180 tb<6>.n179 0.0557941
R9197 tb<6>.n178 tb<6>.n177 0.0557941
R9198 tb<6>.n175 tb<6>.n174 0.0557941
R9199 tb<6>.n174 tb<6>.n173 0.0557941
R9200 tb<6>.n173 tb<6>.n172 0.0557941
R9201 tb<6>.n171 tb<6>.n170 0.0557941
R9202 tb<6>.n168 tb<6>.n167 0.0557941
R9203 tb<6>.n167 tb<6>.n166 0.0557941
R9204 tb<6>.n166 tb<6>.n165 0.0557941
R9205 tb<6>.n164 tb<6>.n163 0.0557941
R9206 tb<6>.n161 tb<6>.n160 0.0557941
R9207 tb<6>.n160 tb<6>.n159 0.0557941
R9208 tb<6>.n159 tb<6>.n158 0.0557941
R9209 tb<6>.n157 tb<6>.n156 0.0557941
R9210 tb<6>.n154 tb<6>.n153 0.0557941
R9211 tb<6>.n153 tb<6>.n152 0.0557941
R9212 tb<6>.n152 tb<6>.n151 0.0557941
R9213 tb<6>.n150 tb<6>.n149 0.0557941
R9214 tb<6>.n147 tb<6>.n146 0.0557941
R9215 tb<6>.n146 tb<6>.n145 0.0557941
R9216 tb<6>.n145 tb<6>.n144 0.0557941
R9217 tb<6>.n143 tb<6>.n142 0.0557941
R9218 tb<6>.n140 tb<6>.n139 0.0557941
R9219 tb<6>.n139 tb<6>.n138 0.0557941
R9220 tb<6>.n138 tb<6>.n137 0.0557941
R9221 tb<6>.n136 tb<6>.n135 0.0557941
R9222 tb<6>.n133 tb<6>.n132 0.0557941
R9223 tb<6>.n132 tb<6>.n131 0.0557941
R9224 tb<6>.n131 tb<6>.n130 0.0557941
R9225 tb<6>.n129 tb<6>.n128 0.0557941
R9226 tb<6>.n126 tb<6>.n125 0.0557941
R9227 tb<6>.n125 tb<6>.n124 0.0557941
R9228 tb<6>.n124 tb<6>.n123 0.0557941
R9229 tb<6>.n122 tb<6>.n121 0.0557941
R9230 tb<6>.n119 tb<6>.n118 0.0557941
R9231 tb<6>.n118 tb<6>.n117 0.0557941
R9232 tb<6>.n117 tb<6>.n116 0.0557941
R9233 tb<6>.n115 tb<6>.n114 0.0557941
R9234 tb<6>.n112 tb<6>.n111 0.0557941
R9235 tb<6>.n111 tb<6>.n110 0.0557941
R9236 tb<6>.n110 tb<6>.n109 0.0557941
R9237 tb<6>.n108 tb<6>.n107 0.0557941
R9238 tb<6>.n105 tb<6>.n104 0.0557941
R9239 tb<6>.n104 tb<6>.n103 0.0557941
R9240 tb<6>.n103 tb<6>.n102 0.0557941
R9241 tb<6>.n101 tb<6>.n100 0.0557941
R9242 tb<6>.n98 tb<6>.n97 0.0557941
R9243 tb<6>.n97 tb<6>.n96 0.0557941
R9244 tb<6>.n96 tb<6>.n95 0.0557941
R9245 tb<6>.n94 tb<6>.n93 0.0557941
R9246 tb<6>.n91 tb<6>.n90 0.0557941
R9247 tb<6>.n90 tb<6>.n89 0.0557941
R9248 tb<6>.n89 tb<6>.n88 0.0557941
R9249 tb<6>.n87 tb<6>.n86 0.0557941
R9250 tb<6>.n84 tb<6>.n83 0.0557941
R9251 tb<6>.n83 tb<6>.n82 0.0557941
R9252 tb<6>.n82 tb<6>.n81 0.0557941
R9253 tb<6>.n80 tb<6>.n79 0.0557941
R9254 tb<6>.n77 tb<6>.n76 0.0557941
R9255 tb<6>.n76 tb<6>.n75 0.0557941
R9256 tb<6>.n75 tb<6>.n74 0.0557941
R9257 tb<6>.n73 tb<6>.n72 0.0557941
R9258 tb<6>.n70 tb<6>.n69 0.0557941
R9259 tb<6>.n69 tb<6>.n68 0.0557941
R9260 tb<6>.n68 tb<6>.n67 0.0557941
R9261 tb<6>.n66 tb<6>.n65 0.0557941
R9262 tb<6>.n63 tb<6>.n62 0.0557941
R9263 tb<6>.n62 tb<6>.n61 0.0557941
R9264 tb<6>.n61 tb<6>.n60 0.0557941
R9265 tb<6>.n59 tb<6>.n58 0.0557941
R9266 tb<6>.n56 tb<6>.n55 0.0557941
R9267 tb<6>.n55 tb<6>.n54 0.0557941
R9268 tb<6>.n54 tb<6>.n53 0.0557941
R9269 tb<6>.n52 tb<6>.n51 0.0557941
R9270 tb<6>.n49 tb<6>.n48 0.0557941
R9271 tb<6>.n48 tb<6>.n47 0.0557941
R9272 tb<6>.n47 tb<6>.n46 0.0557941
R9273 tb<6>.n45 tb<6>.n44 0.0557941
R9274 tb<6>.n42 tb<6>.n41 0.0557941
R9275 tb<6>.n41 tb<6>.n40 0.0557941
R9276 tb<6>.n40 tb<6>.n39 0.0557941
R9277 tb<6>.n38 tb<6>.n37 0.0557941
R9278 tb<6>.n35 tb<6>.n34 0.0557941
R9279 tb<6>.n34 tb<6>.n33 0.0557941
R9280 tb<6>.n33 tb<6>.n32 0.0557941
R9281 tb<6>.n31 tb<6>.n30 0.0557941
R9282 tb<6>.n28 tb<6>.n27 0.0557941
R9283 tb<6>.n27 tb<6>.n26 0.0557941
R9284 tb<6>.n26 tb<6>.n25 0.0557941
R9285 tb<6>.n24 tb<6>.n23 0.0557941
R9286 tb<6>.n21 tb<6>.n20 0.0557941
R9287 tb<6>.n20 tb<6>.n19 0.0557941
R9288 tb<6>.n19 tb<6>.n18 0.0557941
R9289 tb<6>.n17 tb<6>.n16 0.0557941
R9290 tb<6>.n14 tb<6>.n13 0.0557941
R9291 tb<6>.n13 tb<6>.n12 0.0557941
R9292 tb<6>.n12 tb<6>.n11 0.0557941
R9293 tb<6>.n10 tb<6>.n9 0.0557941
R9294 tb<6>.n7 tb<6>.n6 0.0557941
R9295 tb<6>.n6 tb<6>.n5 0.0557941
R9296 tb<6>.n5 tb<6>.n4 0.0557941
R9297 tb<6>.n3 tb<6>.n2 0.0557941
R9298 tb<6>.n397 tb<6>.n396 0.0488824
R9299 tb<6>.n409 tb<6>.n408 0.0419706
R9300 tb<6>.n205 tb<6>.n204 0.0419706
R9301 tb<6>.n198 tb<6>.n197 0.0419706
R9302 tb<6>.n191 tb<6>.n190 0.0419706
R9303 tb<6>.n184 tb<6>.n183 0.0419706
R9304 tb<6>.n177 tb<6>.n176 0.0419706
R9305 tb<6>.n170 tb<6>.n169 0.0419706
R9306 tb<6>.n163 tb<6>.n162 0.0419706
R9307 tb<6>.n156 tb<6>.n155 0.0419706
R9308 tb<6>.n149 tb<6>.n148 0.0419706
R9309 tb<6>.n142 tb<6>.n141 0.0419706
R9310 tb<6>.n135 tb<6>.n134 0.0419706
R9311 tb<6>.n128 tb<6>.n127 0.0419706
R9312 tb<6>.n121 tb<6>.n120 0.0419706
R9313 tb<6>.n114 tb<6>.n113 0.0419706
R9314 tb<6>.n107 tb<6>.n106 0.0419706
R9315 tb<6>.n100 tb<6>.n99 0.0419706
R9316 tb<6>.n93 tb<6>.n92 0.0419706
R9317 tb<6>.n86 tb<6>.n85 0.0419706
R9318 tb<6>.n79 tb<6>.n78 0.0419706
R9319 tb<6>.n72 tb<6>.n71 0.0419706
R9320 tb<6>.n65 tb<6>.n64 0.0419706
R9321 tb<6>.n58 tb<6>.n57 0.0419706
R9322 tb<6>.n51 tb<6>.n50 0.0419706
R9323 tb<6>.n44 tb<6>.n43 0.0419706
R9324 tb<6>.n37 tb<6>.n36 0.0419706
R9325 tb<6>.n30 tb<6>.n29 0.0419706
R9326 tb<6>.n23 tb<6>.n22 0.0419706
R9327 tb<6>.n16 tb<6>.n15 0.0419706
R9328 tb<6>.n9 tb<6>.n8 0.0419706
R9329 tb<6>.n2 tb<6>.n1 0.0419706
R9330 tb<6>.n594 tb<6>.n593 0.0405882
R9331 tb<6>.n411 tb<6>.n410 0.0405882
R9332 tb<6>.n394 tb<6>.n393 0.0405882
R9333 tb<6>.n210 tb<6>.n209 0.0405882
R9334 tb<6>.n595 tb<6>.n594 0.0157059
R9335 tb<6>.n395 tb<6>.n394 0.0157059
R9336 tb<6>.n410 tb<6>.n409 0.0143235
R9337 tb<6>.n204 tb<6>.n203 0.0143235
R9338 tb<6>.n197 tb<6>.n196 0.0143235
R9339 tb<6>.n190 tb<6>.n189 0.0143235
R9340 tb<6>.n183 tb<6>.n182 0.0143235
R9341 tb<6>.n176 tb<6>.n175 0.0143235
R9342 tb<6>.n169 tb<6>.n168 0.0143235
R9343 tb<6>.n162 tb<6>.n161 0.0143235
R9344 tb<6>.n155 tb<6>.n154 0.0143235
R9345 tb<6>.n148 tb<6>.n147 0.0143235
R9346 tb<6>.n141 tb<6>.n140 0.0143235
R9347 tb<6>.n134 tb<6>.n133 0.0143235
R9348 tb<6>.n127 tb<6>.n126 0.0143235
R9349 tb<6>.n120 tb<6>.n119 0.0143235
R9350 tb<6>.n113 tb<6>.n112 0.0143235
R9351 tb<6>.n106 tb<6>.n105 0.0143235
R9352 tb<6>.n99 tb<6>.n98 0.0143235
R9353 tb<6>.n92 tb<6>.n91 0.0143235
R9354 tb<6>.n85 tb<6>.n84 0.0143235
R9355 tb<6>.n78 tb<6>.n77 0.0143235
R9356 tb<6>.n71 tb<6>.n70 0.0143235
R9357 tb<6>.n64 tb<6>.n63 0.0143235
R9358 tb<6>.n57 tb<6>.n56 0.0143235
R9359 tb<6>.n50 tb<6>.n49 0.0143235
R9360 tb<6>.n43 tb<6>.n42 0.0143235
R9361 tb<6>.n36 tb<6>.n35 0.0143235
R9362 tb<6>.n29 tb<6>.n28 0.0143235
R9363 tb<6>.n22 tb<6>.n21 0.0143235
R9364 tb<6>.n15 tb<6>.n14 0.0143235
R9365 tb<6>.n8 tb<6>.n7 0.0143235
R9366 tb<6>.n600 tb<6>.n599 0.0100455
R9367 tb<6>.n412 tb<6>.n411 0.0098016
R9368 tb<6>.n211 tb<6>.n210 0.0098016
R9369 tb<6>.n405 tb<6>.n404 0.0089954
R9370 tb<6>.n214 tb<6>.n213 0.00892479
R9371 tb<6>.n598 tb<6>.n407 0.00883373
R9372 tb<6>.n598 tb<6>.n597 0.00783691
R9373 tb<6>.n596 tb<6>.n595 0.00741176
R9374 tb<6>.n396 tb<6>.n395 0.00741176
R9375 tb<6>.n400 tb<6>.n399 0.00606092
R9376 tb<6>.n399 tb<6>.n398 0.00567797
R9377 tb<6>.n398 tb<6>.n214 0.00494174
R9378 tb<6> tb<6>.n600 0.00455166
R9379 tb<6>.n402 tb<6>.n401 0.00349062
R9380 tb<6>.n599 tb<6>.n403 0.00347205
R9381 tb<6>.n597 tb<6>.n412 0.00249153
R9382 tb<6>.n213 tb<6>.n212 0.00249153
R9383 tb<6>.n212 tb<6>.n211 0.00249153
R9384 t<6>.n395 t<6>.n394 3.4105
R9385 t<6>.n396 t<6>.n3 3.4105
R9386 t<6>.n393 t<6>.n5 1.7055
R9387 t<6>.n392 t<6>.n391 1.7055
R9388 t<6>.n390 t<6>.n6 1.7055
R9389 t<6>.n389 t<6>.n388 1.7055
R9390 t<6>.n387 t<6>.n7 1.7055
R9391 t<6>.n386 t<6>.n385 1.7055
R9392 t<6>.n384 t<6>.n8 1.7055
R9393 t<6>.n383 t<6>.n382 1.7055
R9394 t<6>.n381 t<6>.n10 1.7055
R9395 t<6>.n380 t<6>.n379 1.7055
R9396 t<6>.n378 t<6>.n11 1.7055
R9397 t<6>.n376 t<6>.n375 1.7055
R9398 t<6>.n374 t<6>.n12 1.7055
R9399 t<6>.n373 t<6>.n372 1.7055
R9400 t<6>.n371 t<6>.n13 1.7055
R9401 t<6>.n370 t<6>.n369 1.7055
R9402 t<6>.n368 t<6>.n14 1.7055
R9403 t<6>.n367 t<6>.n366 1.7055
R9404 t<6>.n365 t<6>.n15 1.7055
R9405 t<6>.n364 t<6>.n363 1.7055
R9406 t<6>.n362 t<6>.n17 1.7055
R9407 t<6>.n361 t<6>.n360 1.7055
R9408 t<6>.n359 t<6>.n18 1.7055
R9409 t<6>.n357 t<6>.n356 1.7055
R9410 t<6>.n355 t<6>.n19 1.7055
R9411 t<6>.n354 t<6>.n353 1.7055
R9412 t<6>.n352 t<6>.n20 1.7055
R9413 t<6>.n351 t<6>.n350 1.7055
R9414 t<6>.n349 t<6>.n21 1.7055
R9415 t<6>.n348 t<6>.n347 1.7055
R9416 t<6>.n346 t<6>.n22 1.7055
R9417 t<6>.n345 t<6>.n344 1.7055
R9418 t<6>.n343 t<6>.n24 1.7055
R9419 t<6>.n342 t<6>.n341 1.7055
R9420 t<6>.n340 t<6>.n25 1.7055
R9421 t<6>.n338 t<6>.n337 1.7055
R9422 t<6>.n336 t<6>.n26 1.7055
R9423 t<6>.n335 t<6>.n334 1.7055
R9424 t<6>.n333 t<6>.n27 1.7055
R9425 t<6>.n332 t<6>.n331 1.7055
R9426 t<6>.n330 t<6>.n28 1.7055
R9427 t<6>.n329 t<6>.n328 1.7055
R9428 t<6>.n327 t<6>.n29 1.7055
R9429 t<6>.n326 t<6>.n325 1.7055
R9430 t<6>.n324 t<6>.n31 1.7055
R9431 t<6>.n323 t<6>.n322 1.7055
R9432 t<6>.n321 t<6>.n32 1.7055
R9433 t<6>.n319 t<6>.n318 1.7055
R9434 t<6>.n317 t<6>.n33 1.7055
R9435 t<6>.n316 t<6>.n315 1.7055
R9436 t<6>.n314 t<6>.n34 1.7055
R9437 t<6>.n313 t<6>.n312 1.7055
R9438 t<6>.n311 t<6>.n35 1.7055
R9439 t<6>.n310 t<6>.n309 1.7055
R9440 t<6>.n308 t<6>.n36 1.7055
R9441 t<6>.n307 t<6>.n306 1.7055
R9442 t<6>.n305 t<6>.n38 1.7055
R9443 t<6>.n304 t<6>.n303 1.7055
R9444 t<6>.n302 t<6>.n39 1.7055
R9445 t<6>.n300 t<6>.n299 1.7055
R9446 t<6>.n298 t<6>.n40 1.7055
R9447 t<6>.n297 t<6>.n296 1.7055
R9448 t<6>.n295 t<6>.n41 1.7055
R9449 t<6>.n294 t<6>.n293 1.7055
R9450 t<6>.n292 t<6>.n42 1.7055
R9451 t<6>.n291 t<6>.n290 1.7055
R9452 t<6>.n289 t<6>.n43 1.7055
R9453 t<6>.n288 t<6>.n287 1.7055
R9454 t<6>.n286 t<6>.n45 1.7055
R9455 t<6>.n285 t<6>.n284 1.7055
R9456 t<6>.n283 t<6>.n46 1.7055
R9457 t<6>.n281 t<6>.n280 1.7055
R9458 t<6>.n279 t<6>.n47 1.7055
R9459 t<6>.n278 t<6>.n277 1.7055
R9460 t<6>.n276 t<6>.n48 1.7055
R9461 t<6>.n275 t<6>.n274 1.7055
R9462 t<6>.n273 t<6>.n49 1.7055
R9463 t<6>.n272 t<6>.n271 1.7055
R9464 t<6>.n270 t<6>.n50 1.7055
R9465 t<6>.n269 t<6>.n268 1.7055
R9466 t<6>.n267 t<6>.n52 1.7055
R9467 t<6>.n266 t<6>.n265 1.7055
R9468 t<6>.n264 t<6>.n53 1.7055
R9469 t<6>.n262 t<6>.n261 1.7055
R9470 t<6>.n260 t<6>.n54 1.7055
R9471 t<6>.n259 t<6>.n258 1.7055
R9472 t<6>.n257 t<6>.n55 1.7055
R9473 t<6>.n256 t<6>.n255 1.7055
R9474 t<6>.n254 t<6>.n56 1.7055
R9475 t<6>.n253 t<6>.n252 1.7055
R9476 t<6>.n251 t<6>.n57 1.7055
R9477 t<6>.n250 t<6>.n249 1.7055
R9478 t<6>.n248 t<6>.n59 1.7055
R9479 t<6>.n247 t<6>.n246 1.7055
R9480 t<6>.n245 t<6>.n60 1.7055
R9481 t<6>.n243 t<6>.n242 1.7055
R9482 t<6>.n241 t<6>.n61 1.7055
R9483 t<6>.n240 t<6>.n239 1.7055
R9484 t<6>.n238 t<6>.n62 1.7055
R9485 t<6>.n237 t<6>.n236 1.7055
R9486 t<6>.n235 t<6>.n63 1.7055
R9487 t<6>.n234 t<6>.n233 1.7055
R9488 t<6>.n232 t<6>.n64 1.7055
R9489 t<6>.n231 t<6>.n230 1.7055
R9490 t<6>.n229 t<6>.n66 1.7055
R9491 t<6>.n228 t<6>.n227 1.7055
R9492 t<6>.n226 t<6>.n67 1.7055
R9493 t<6>.n224 t<6>.n223 1.7055
R9494 t<6>.n222 t<6>.n68 1.7055
R9495 t<6>.n221 t<6>.n220 1.7055
R9496 t<6>.n219 t<6>.n69 1.7055
R9497 t<6>.n218 t<6>.n217 1.7055
R9498 t<6>.n216 t<6>.n70 1.7055
R9499 t<6>.n215 t<6>.n214 1.7055
R9500 t<6>.n213 t<6>.n71 1.7055
R9501 t<6>.n212 t<6>.n211 1.7055
R9502 t<6>.n210 t<6>.n73 1.7055
R9503 t<6>.n209 t<6>.n208 1.7055
R9504 t<6>.n207 t<6>.n74 1.7055
R9505 t<6>.n205 t<6>.n204 1.7055
R9506 t<6>.n203 t<6>.n75 1.7055
R9507 t<6>.n202 t<6>.n201 1.7055
R9508 t<6>.n200 t<6>.n76 1.7055
R9509 t<6>.n199 t<6>.n198 1.7055
R9510 t<6>.n197 t<6>.n77 1.7055
R9511 t<6>.n196 t<6>.n195 1.7055
R9512 t<6>.n194 t<6>.n78 1.7055
R9513 t<6>.n193 t<6>.n192 1.7055
R9514 t<6>.n191 t<6>.n80 1.7055
R9515 t<6>.n190 t<6>.n189 1.7055
R9516 t<6>.n188 t<6>.n81 1.7055
R9517 t<6>.n186 t<6>.n185 1.7055
R9518 t<6>.n184 t<6>.n82 1.7055
R9519 t<6>.n183 t<6>.n182 1.7055
R9520 t<6>.n181 t<6>.n83 1.7055
R9521 t<6>.n180 t<6>.n179 1.7055
R9522 t<6>.n178 t<6>.n84 1.7055
R9523 t<6>.n177 t<6>.n176 1.7055
R9524 t<6>.n175 t<6>.n85 1.7055
R9525 t<6>.n174 t<6>.n173 1.7055
R9526 t<6>.n172 t<6>.n87 1.7055
R9527 t<6>.n171 t<6>.n170 1.7055
R9528 t<6>.n169 t<6>.n88 1.7055
R9529 t<6>.n167 t<6>.n166 1.7055
R9530 t<6>.n165 t<6>.n89 1.7055
R9531 t<6>.n164 t<6>.n163 1.7055
R9532 t<6>.n162 t<6>.n90 1.7055
R9533 t<6>.n161 t<6>.n160 1.7055
R9534 t<6>.n159 t<6>.n91 1.7055
R9535 t<6>.n158 t<6>.n157 1.7055
R9536 t<6>.n156 t<6>.n92 1.7055
R9537 t<6>.n155 t<6>.n154 1.7055
R9538 t<6>.n153 t<6>.n94 1.7055
R9539 t<6>.n152 t<6>.n151 1.7055
R9540 t<6>.n150 t<6>.n95 1.7055
R9541 t<6>.n148 t<6>.n147 1.7055
R9542 t<6>.n146 t<6>.n96 1.7055
R9543 t<6>.n145 t<6>.n144 1.7055
R9544 t<6>.n143 t<6>.n97 1.7055
R9545 t<6>.n142 t<6>.n141 1.7055
R9546 t<6>.n140 t<6>.n98 1.7055
R9547 t<6>.n139 t<6>.n138 1.7055
R9548 t<6>.n137 t<6>.n99 1.7055
R9549 t<6>.n136 t<6>.n135 1.7055
R9550 t<6>.n134 t<6>.n101 1.7055
R9551 t<6>.n133 t<6>.n132 1.7055
R9552 t<6>.n131 t<6>.n102 1.7055
R9553 t<6>.n129 t<6>.n128 1.7055
R9554 t<6>.n127 t<6>.n103 1.7055
R9555 t<6>.n126 t<6>.n125 1.7055
R9556 t<6>.n124 t<6>.n104 1.7055
R9557 t<6>.n123 t<6>.n122 1.7055
R9558 t<6>.n121 t<6>.n105 1.7055
R9559 t<6>.n120 t<6>.n119 1.7055
R9560 t<6>.n118 t<6>.n106 1.7055
R9561 t<6>.n117 t<6>.n116 1.7055
R9562 t<6>.n115 t<6>.n108 1.7055
R9563 t<6>.n114 t<6>.n113 1.7055
R9564 t<6>.n112 t<6>.n109 1.7055
R9565 t<6>.n399 t<6>.n1 0.404561
R9566 t<6>.n596 t<6>.n595 0.3805
R9567 t<6>.n397 t<6>.n0 0.3805
R9568 t<6>.n398 t<6>.n397 0.3805
R9569 t<6>.n402 t<6>.n401 0.3805
R9570 t<6>.n407 t<6>.n406 0.3424
R9571 t<6>.n400 t<6>.n399 0.3424
R9572 t<6>.n110 t<6>.n109 0.304086
R9573 t<6>.n110 t<6> 0.271393
R9574 t<6>.n2 t<6>.n0 0.189029
R9575 t<6>.n111 t<6>.n110 0.174213
R9576 t<6>.n388 t<6>.n6 0.142882
R9577 t<6>.n381 t<6>.n380 0.142882
R9578 t<6>.n369 t<6>.n13 0.142882
R9579 t<6>.n362 t<6>.n361 0.142882
R9580 t<6>.n350 t<6>.n20 0.142882
R9581 t<6>.n343 t<6>.n342 0.142882
R9582 t<6>.n331 t<6>.n27 0.142882
R9583 t<6>.n324 t<6>.n323 0.142882
R9584 t<6>.n312 t<6>.n34 0.142882
R9585 t<6>.n305 t<6>.n304 0.142882
R9586 t<6>.n293 t<6>.n41 0.142882
R9587 t<6>.n286 t<6>.n285 0.142882
R9588 t<6>.n274 t<6>.n48 0.142882
R9589 t<6>.n267 t<6>.n266 0.142882
R9590 t<6>.n255 t<6>.n55 0.142882
R9591 t<6>.n248 t<6>.n247 0.142882
R9592 t<6>.n236 t<6>.n62 0.142882
R9593 t<6>.n229 t<6>.n228 0.142882
R9594 t<6>.n217 t<6>.n69 0.142882
R9595 t<6>.n210 t<6>.n209 0.142882
R9596 t<6>.n198 t<6>.n76 0.142882
R9597 t<6>.n191 t<6>.n190 0.142882
R9598 t<6>.n179 t<6>.n83 0.142882
R9599 t<6>.n172 t<6>.n171 0.142882
R9600 t<6>.n160 t<6>.n90 0.142882
R9601 t<6>.n153 t<6>.n152 0.142882
R9602 t<6>.n141 t<6>.n97 0.142882
R9603 t<6>.n134 t<6>.n133 0.142882
R9604 t<6>.n122 t<6>.n104 0.142882
R9605 t<6>.n115 t<6>.n114 0.142882
R9606 t<6>.n390 t<6>.n389 0.142882
R9607 t<6>.n379 t<6>.n10 0.142882
R9608 t<6>.n371 t<6>.n370 0.142882
R9609 t<6>.n360 t<6>.n17 0.142882
R9610 t<6>.n352 t<6>.n351 0.142882
R9611 t<6>.n341 t<6>.n24 0.142882
R9612 t<6>.n333 t<6>.n332 0.142882
R9613 t<6>.n322 t<6>.n31 0.142882
R9614 t<6>.n314 t<6>.n313 0.142882
R9615 t<6>.n303 t<6>.n38 0.142882
R9616 t<6>.n295 t<6>.n294 0.142882
R9617 t<6>.n284 t<6>.n45 0.142882
R9618 t<6>.n276 t<6>.n275 0.142882
R9619 t<6>.n265 t<6>.n52 0.142882
R9620 t<6>.n257 t<6>.n256 0.142882
R9621 t<6>.n246 t<6>.n59 0.142882
R9622 t<6>.n238 t<6>.n237 0.142882
R9623 t<6>.n227 t<6>.n66 0.142882
R9624 t<6>.n219 t<6>.n218 0.142882
R9625 t<6>.n208 t<6>.n73 0.142882
R9626 t<6>.n200 t<6>.n199 0.142882
R9627 t<6>.n189 t<6>.n80 0.142882
R9628 t<6>.n181 t<6>.n180 0.142882
R9629 t<6>.n170 t<6>.n87 0.142882
R9630 t<6>.n162 t<6>.n161 0.142882
R9631 t<6>.n151 t<6>.n94 0.142882
R9632 t<6>.n143 t<6>.n142 0.142882
R9633 t<6>.n132 t<6>.n101 0.142882
R9634 t<6>.n124 t<6>.n123 0.142882
R9635 t<6>.n113 t<6>.n108 0.142882
R9636 t<6>.n590 t<6>.n589 0.142882
R9637 t<6>.n584 t<6>.n583 0.142882
R9638 t<6>.n578 t<6>.n577 0.142882
R9639 t<6>.n572 t<6>.n571 0.142882
R9640 t<6>.n566 t<6>.n565 0.142882
R9641 t<6>.n560 t<6>.n559 0.142882
R9642 t<6>.n554 t<6>.n553 0.142882
R9643 t<6>.n548 t<6>.n547 0.142882
R9644 t<6>.n542 t<6>.n541 0.142882
R9645 t<6>.n536 t<6>.n535 0.142882
R9646 t<6>.n530 t<6>.n529 0.142882
R9647 t<6>.n524 t<6>.n523 0.142882
R9648 t<6>.n518 t<6>.n517 0.142882
R9649 t<6>.n512 t<6>.n511 0.142882
R9650 t<6>.n506 t<6>.n505 0.142882
R9651 t<6>.n500 t<6>.n499 0.142882
R9652 t<6>.n494 t<6>.n493 0.142882
R9653 t<6>.n488 t<6>.n487 0.142882
R9654 t<6>.n482 t<6>.n481 0.142882
R9655 t<6>.n476 t<6>.n475 0.142882
R9656 t<6>.n470 t<6>.n469 0.142882
R9657 t<6>.n464 t<6>.n463 0.142882
R9658 t<6>.n458 t<6>.n457 0.142882
R9659 t<6>.n452 t<6>.n451 0.142882
R9660 t<6>.n446 t<6>.n445 0.142882
R9661 t<6>.n440 t<6>.n439 0.142882
R9662 t<6>.n434 t<6>.n433 0.142882
R9663 t<6>.n428 t<6>.n427 0.142882
R9664 t<6>.n422 t<6>.n421 0.142882
R9665 t<6>.n416 t<6>.n415 0.142882
R9666 t<6>.n598 t<6>.n405 0.127395
R9667 t<6>.n403 t<6> 0.125633
R9668 t<6>.n598 t<6>.n597 0.124744
R9669 t<6>.n111 t<6> 0.0976333
R9670 t<6>.n107 t<6> 0.0976333
R9671 t<6>.n130 t<6> 0.0976333
R9672 t<6>.n100 t<6> 0.0976333
R9673 t<6>.n149 t<6> 0.0976333
R9674 t<6>.n93 t<6> 0.0976333
R9675 t<6>.n168 t<6> 0.0976333
R9676 t<6>.n86 t<6> 0.0976333
R9677 t<6>.n187 t<6> 0.0976333
R9678 t<6>.n79 t<6> 0.0976333
R9679 t<6>.n206 t<6> 0.0976333
R9680 t<6>.n72 t<6> 0.0976333
R9681 t<6>.n225 t<6> 0.0976333
R9682 t<6>.n65 t<6> 0.0976333
R9683 t<6>.n244 t<6> 0.0976333
R9684 t<6>.n58 t<6> 0.0976333
R9685 t<6>.n263 t<6> 0.0976333
R9686 t<6>.n51 t<6> 0.0976333
R9687 t<6>.n282 t<6> 0.0976333
R9688 t<6>.n44 t<6> 0.0976333
R9689 t<6>.n301 t<6> 0.0976333
R9690 t<6>.n37 t<6> 0.0976333
R9691 t<6>.n320 t<6> 0.0976333
R9692 t<6>.n30 t<6> 0.0976333
R9693 t<6>.n339 t<6> 0.0976333
R9694 t<6>.n23 t<6> 0.0976333
R9695 t<6>.n358 t<6> 0.0976333
R9696 t<6>.n16 t<6> 0.0976333
R9697 t<6>.n377 t<6> 0.0976333
R9698 t<6>.n9 t<6> 0.0976333
R9699 t<6>.n4 t<6> 0.0976333
R9700 t<6> t<6>.n402 0.0796156
R9701 t<6>.n1 t<6>.n0 0.0762548
R9702 t<6>.n408 t<6> 0.0725667
R9703 t<6>.n393 t<6>.n392 0.0557941
R9704 t<6>.n392 t<6>.n6 0.0557941
R9705 t<6>.n388 t<6>.n387 0.0557941
R9706 t<6>.n387 t<6>.n386 0.0557941
R9707 t<6>.n386 t<6>.n8 0.0557941
R9708 t<6>.n382 t<6>.n8 0.0557941
R9709 t<6>.n382 t<6>.n381 0.0557941
R9710 t<6>.n380 t<6>.n11 0.0557941
R9711 t<6>.n375 t<6>.n11 0.0557941
R9712 t<6>.n375 t<6>.n374 0.0557941
R9713 t<6>.n374 t<6>.n373 0.0557941
R9714 t<6>.n373 t<6>.n13 0.0557941
R9715 t<6>.n369 t<6>.n368 0.0557941
R9716 t<6>.n368 t<6>.n367 0.0557941
R9717 t<6>.n367 t<6>.n15 0.0557941
R9718 t<6>.n363 t<6>.n15 0.0557941
R9719 t<6>.n363 t<6>.n362 0.0557941
R9720 t<6>.n361 t<6>.n18 0.0557941
R9721 t<6>.n356 t<6>.n18 0.0557941
R9722 t<6>.n356 t<6>.n355 0.0557941
R9723 t<6>.n355 t<6>.n354 0.0557941
R9724 t<6>.n354 t<6>.n20 0.0557941
R9725 t<6>.n350 t<6>.n349 0.0557941
R9726 t<6>.n349 t<6>.n348 0.0557941
R9727 t<6>.n348 t<6>.n22 0.0557941
R9728 t<6>.n344 t<6>.n22 0.0557941
R9729 t<6>.n344 t<6>.n343 0.0557941
R9730 t<6>.n342 t<6>.n25 0.0557941
R9731 t<6>.n337 t<6>.n25 0.0557941
R9732 t<6>.n337 t<6>.n336 0.0557941
R9733 t<6>.n336 t<6>.n335 0.0557941
R9734 t<6>.n335 t<6>.n27 0.0557941
R9735 t<6>.n331 t<6>.n330 0.0557941
R9736 t<6>.n330 t<6>.n329 0.0557941
R9737 t<6>.n329 t<6>.n29 0.0557941
R9738 t<6>.n325 t<6>.n29 0.0557941
R9739 t<6>.n325 t<6>.n324 0.0557941
R9740 t<6>.n323 t<6>.n32 0.0557941
R9741 t<6>.n318 t<6>.n32 0.0557941
R9742 t<6>.n318 t<6>.n317 0.0557941
R9743 t<6>.n317 t<6>.n316 0.0557941
R9744 t<6>.n316 t<6>.n34 0.0557941
R9745 t<6>.n312 t<6>.n311 0.0557941
R9746 t<6>.n311 t<6>.n310 0.0557941
R9747 t<6>.n310 t<6>.n36 0.0557941
R9748 t<6>.n306 t<6>.n36 0.0557941
R9749 t<6>.n306 t<6>.n305 0.0557941
R9750 t<6>.n304 t<6>.n39 0.0557941
R9751 t<6>.n299 t<6>.n39 0.0557941
R9752 t<6>.n299 t<6>.n298 0.0557941
R9753 t<6>.n298 t<6>.n297 0.0557941
R9754 t<6>.n297 t<6>.n41 0.0557941
R9755 t<6>.n293 t<6>.n292 0.0557941
R9756 t<6>.n292 t<6>.n291 0.0557941
R9757 t<6>.n291 t<6>.n43 0.0557941
R9758 t<6>.n287 t<6>.n43 0.0557941
R9759 t<6>.n287 t<6>.n286 0.0557941
R9760 t<6>.n285 t<6>.n46 0.0557941
R9761 t<6>.n280 t<6>.n46 0.0557941
R9762 t<6>.n280 t<6>.n279 0.0557941
R9763 t<6>.n279 t<6>.n278 0.0557941
R9764 t<6>.n278 t<6>.n48 0.0557941
R9765 t<6>.n274 t<6>.n273 0.0557941
R9766 t<6>.n273 t<6>.n272 0.0557941
R9767 t<6>.n272 t<6>.n50 0.0557941
R9768 t<6>.n268 t<6>.n50 0.0557941
R9769 t<6>.n268 t<6>.n267 0.0557941
R9770 t<6>.n266 t<6>.n53 0.0557941
R9771 t<6>.n261 t<6>.n53 0.0557941
R9772 t<6>.n261 t<6>.n260 0.0557941
R9773 t<6>.n260 t<6>.n259 0.0557941
R9774 t<6>.n259 t<6>.n55 0.0557941
R9775 t<6>.n255 t<6>.n254 0.0557941
R9776 t<6>.n254 t<6>.n253 0.0557941
R9777 t<6>.n253 t<6>.n57 0.0557941
R9778 t<6>.n249 t<6>.n57 0.0557941
R9779 t<6>.n249 t<6>.n248 0.0557941
R9780 t<6>.n247 t<6>.n60 0.0557941
R9781 t<6>.n242 t<6>.n60 0.0557941
R9782 t<6>.n242 t<6>.n241 0.0557941
R9783 t<6>.n241 t<6>.n240 0.0557941
R9784 t<6>.n240 t<6>.n62 0.0557941
R9785 t<6>.n236 t<6>.n235 0.0557941
R9786 t<6>.n235 t<6>.n234 0.0557941
R9787 t<6>.n234 t<6>.n64 0.0557941
R9788 t<6>.n230 t<6>.n64 0.0557941
R9789 t<6>.n230 t<6>.n229 0.0557941
R9790 t<6>.n228 t<6>.n67 0.0557941
R9791 t<6>.n223 t<6>.n67 0.0557941
R9792 t<6>.n223 t<6>.n222 0.0557941
R9793 t<6>.n222 t<6>.n221 0.0557941
R9794 t<6>.n221 t<6>.n69 0.0557941
R9795 t<6>.n217 t<6>.n216 0.0557941
R9796 t<6>.n216 t<6>.n215 0.0557941
R9797 t<6>.n215 t<6>.n71 0.0557941
R9798 t<6>.n211 t<6>.n71 0.0557941
R9799 t<6>.n211 t<6>.n210 0.0557941
R9800 t<6>.n209 t<6>.n74 0.0557941
R9801 t<6>.n204 t<6>.n74 0.0557941
R9802 t<6>.n204 t<6>.n203 0.0557941
R9803 t<6>.n203 t<6>.n202 0.0557941
R9804 t<6>.n202 t<6>.n76 0.0557941
R9805 t<6>.n198 t<6>.n197 0.0557941
R9806 t<6>.n197 t<6>.n196 0.0557941
R9807 t<6>.n196 t<6>.n78 0.0557941
R9808 t<6>.n192 t<6>.n78 0.0557941
R9809 t<6>.n192 t<6>.n191 0.0557941
R9810 t<6>.n190 t<6>.n81 0.0557941
R9811 t<6>.n185 t<6>.n81 0.0557941
R9812 t<6>.n185 t<6>.n184 0.0557941
R9813 t<6>.n184 t<6>.n183 0.0557941
R9814 t<6>.n183 t<6>.n83 0.0557941
R9815 t<6>.n179 t<6>.n178 0.0557941
R9816 t<6>.n178 t<6>.n177 0.0557941
R9817 t<6>.n177 t<6>.n85 0.0557941
R9818 t<6>.n173 t<6>.n85 0.0557941
R9819 t<6>.n173 t<6>.n172 0.0557941
R9820 t<6>.n171 t<6>.n88 0.0557941
R9821 t<6>.n166 t<6>.n88 0.0557941
R9822 t<6>.n166 t<6>.n165 0.0557941
R9823 t<6>.n165 t<6>.n164 0.0557941
R9824 t<6>.n164 t<6>.n90 0.0557941
R9825 t<6>.n160 t<6>.n159 0.0557941
R9826 t<6>.n159 t<6>.n158 0.0557941
R9827 t<6>.n158 t<6>.n92 0.0557941
R9828 t<6>.n154 t<6>.n92 0.0557941
R9829 t<6>.n154 t<6>.n153 0.0557941
R9830 t<6>.n152 t<6>.n95 0.0557941
R9831 t<6>.n147 t<6>.n95 0.0557941
R9832 t<6>.n147 t<6>.n146 0.0557941
R9833 t<6>.n146 t<6>.n145 0.0557941
R9834 t<6>.n145 t<6>.n97 0.0557941
R9835 t<6>.n141 t<6>.n140 0.0557941
R9836 t<6>.n140 t<6>.n139 0.0557941
R9837 t<6>.n139 t<6>.n99 0.0557941
R9838 t<6>.n135 t<6>.n99 0.0557941
R9839 t<6>.n135 t<6>.n134 0.0557941
R9840 t<6>.n133 t<6>.n102 0.0557941
R9841 t<6>.n128 t<6>.n102 0.0557941
R9842 t<6>.n128 t<6>.n127 0.0557941
R9843 t<6>.n127 t<6>.n126 0.0557941
R9844 t<6>.n126 t<6>.n104 0.0557941
R9845 t<6>.n122 t<6>.n121 0.0557941
R9846 t<6>.n121 t<6>.n120 0.0557941
R9847 t<6>.n120 t<6>.n106 0.0557941
R9848 t<6>.n116 t<6>.n106 0.0557941
R9849 t<6>.n116 t<6>.n115 0.0557941
R9850 t<6>.n114 t<6>.n109 0.0557941
R9851 t<6>.n391 t<6>.n5 0.0557941
R9852 t<6>.n391 t<6>.n390 0.0557941
R9853 t<6>.n389 t<6>.n7 0.0557941
R9854 t<6>.n385 t<6>.n384 0.0557941
R9855 t<6>.n384 t<6>.n383 0.0557941
R9856 t<6>.n383 t<6>.n10 0.0557941
R9857 t<6>.n379 t<6>.n378 0.0557941
R9858 t<6>.n376 t<6>.n12 0.0557941
R9859 t<6>.n372 t<6>.n12 0.0557941
R9860 t<6>.n372 t<6>.n371 0.0557941
R9861 t<6>.n370 t<6>.n14 0.0557941
R9862 t<6>.n366 t<6>.n365 0.0557941
R9863 t<6>.n365 t<6>.n364 0.0557941
R9864 t<6>.n364 t<6>.n17 0.0557941
R9865 t<6>.n360 t<6>.n359 0.0557941
R9866 t<6>.n357 t<6>.n19 0.0557941
R9867 t<6>.n353 t<6>.n19 0.0557941
R9868 t<6>.n353 t<6>.n352 0.0557941
R9869 t<6>.n351 t<6>.n21 0.0557941
R9870 t<6>.n347 t<6>.n346 0.0557941
R9871 t<6>.n346 t<6>.n345 0.0557941
R9872 t<6>.n345 t<6>.n24 0.0557941
R9873 t<6>.n341 t<6>.n340 0.0557941
R9874 t<6>.n338 t<6>.n26 0.0557941
R9875 t<6>.n334 t<6>.n26 0.0557941
R9876 t<6>.n334 t<6>.n333 0.0557941
R9877 t<6>.n332 t<6>.n28 0.0557941
R9878 t<6>.n328 t<6>.n327 0.0557941
R9879 t<6>.n327 t<6>.n326 0.0557941
R9880 t<6>.n326 t<6>.n31 0.0557941
R9881 t<6>.n322 t<6>.n321 0.0557941
R9882 t<6>.n319 t<6>.n33 0.0557941
R9883 t<6>.n315 t<6>.n33 0.0557941
R9884 t<6>.n315 t<6>.n314 0.0557941
R9885 t<6>.n313 t<6>.n35 0.0557941
R9886 t<6>.n309 t<6>.n308 0.0557941
R9887 t<6>.n308 t<6>.n307 0.0557941
R9888 t<6>.n307 t<6>.n38 0.0557941
R9889 t<6>.n303 t<6>.n302 0.0557941
R9890 t<6>.n300 t<6>.n40 0.0557941
R9891 t<6>.n296 t<6>.n40 0.0557941
R9892 t<6>.n296 t<6>.n295 0.0557941
R9893 t<6>.n294 t<6>.n42 0.0557941
R9894 t<6>.n290 t<6>.n289 0.0557941
R9895 t<6>.n289 t<6>.n288 0.0557941
R9896 t<6>.n288 t<6>.n45 0.0557941
R9897 t<6>.n284 t<6>.n283 0.0557941
R9898 t<6>.n281 t<6>.n47 0.0557941
R9899 t<6>.n277 t<6>.n47 0.0557941
R9900 t<6>.n277 t<6>.n276 0.0557941
R9901 t<6>.n275 t<6>.n49 0.0557941
R9902 t<6>.n271 t<6>.n270 0.0557941
R9903 t<6>.n270 t<6>.n269 0.0557941
R9904 t<6>.n269 t<6>.n52 0.0557941
R9905 t<6>.n265 t<6>.n264 0.0557941
R9906 t<6>.n262 t<6>.n54 0.0557941
R9907 t<6>.n258 t<6>.n54 0.0557941
R9908 t<6>.n258 t<6>.n257 0.0557941
R9909 t<6>.n256 t<6>.n56 0.0557941
R9910 t<6>.n252 t<6>.n251 0.0557941
R9911 t<6>.n251 t<6>.n250 0.0557941
R9912 t<6>.n250 t<6>.n59 0.0557941
R9913 t<6>.n246 t<6>.n245 0.0557941
R9914 t<6>.n243 t<6>.n61 0.0557941
R9915 t<6>.n239 t<6>.n61 0.0557941
R9916 t<6>.n239 t<6>.n238 0.0557941
R9917 t<6>.n237 t<6>.n63 0.0557941
R9918 t<6>.n233 t<6>.n232 0.0557941
R9919 t<6>.n232 t<6>.n231 0.0557941
R9920 t<6>.n231 t<6>.n66 0.0557941
R9921 t<6>.n227 t<6>.n226 0.0557941
R9922 t<6>.n224 t<6>.n68 0.0557941
R9923 t<6>.n220 t<6>.n68 0.0557941
R9924 t<6>.n220 t<6>.n219 0.0557941
R9925 t<6>.n218 t<6>.n70 0.0557941
R9926 t<6>.n214 t<6>.n213 0.0557941
R9927 t<6>.n213 t<6>.n212 0.0557941
R9928 t<6>.n212 t<6>.n73 0.0557941
R9929 t<6>.n208 t<6>.n207 0.0557941
R9930 t<6>.n205 t<6>.n75 0.0557941
R9931 t<6>.n201 t<6>.n75 0.0557941
R9932 t<6>.n201 t<6>.n200 0.0557941
R9933 t<6>.n199 t<6>.n77 0.0557941
R9934 t<6>.n195 t<6>.n194 0.0557941
R9935 t<6>.n194 t<6>.n193 0.0557941
R9936 t<6>.n193 t<6>.n80 0.0557941
R9937 t<6>.n189 t<6>.n188 0.0557941
R9938 t<6>.n186 t<6>.n82 0.0557941
R9939 t<6>.n182 t<6>.n82 0.0557941
R9940 t<6>.n182 t<6>.n181 0.0557941
R9941 t<6>.n180 t<6>.n84 0.0557941
R9942 t<6>.n176 t<6>.n175 0.0557941
R9943 t<6>.n175 t<6>.n174 0.0557941
R9944 t<6>.n174 t<6>.n87 0.0557941
R9945 t<6>.n170 t<6>.n169 0.0557941
R9946 t<6>.n167 t<6>.n89 0.0557941
R9947 t<6>.n163 t<6>.n89 0.0557941
R9948 t<6>.n163 t<6>.n162 0.0557941
R9949 t<6>.n161 t<6>.n91 0.0557941
R9950 t<6>.n157 t<6>.n156 0.0557941
R9951 t<6>.n156 t<6>.n155 0.0557941
R9952 t<6>.n155 t<6>.n94 0.0557941
R9953 t<6>.n151 t<6>.n150 0.0557941
R9954 t<6>.n148 t<6>.n96 0.0557941
R9955 t<6>.n144 t<6>.n96 0.0557941
R9956 t<6>.n144 t<6>.n143 0.0557941
R9957 t<6>.n142 t<6>.n98 0.0557941
R9958 t<6>.n138 t<6>.n137 0.0557941
R9959 t<6>.n137 t<6>.n136 0.0557941
R9960 t<6>.n136 t<6>.n101 0.0557941
R9961 t<6>.n132 t<6>.n131 0.0557941
R9962 t<6>.n129 t<6>.n103 0.0557941
R9963 t<6>.n125 t<6>.n103 0.0557941
R9964 t<6>.n125 t<6>.n124 0.0557941
R9965 t<6>.n123 t<6>.n105 0.0557941
R9966 t<6>.n119 t<6>.n118 0.0557941
R9967 t<6>.n118 t<6>.n117 0.0557941
R9968 t<6>.n117 t<6>.n108 0.0557941
R9969 t<6>.n113 t<6>.n112 0.0557941
R9970 t<6>.n592 t<6>.n591 0.0557941
R9971 t<6>.n591 t<6>.n590 0.0557941
R9972 t<6>.n589 t<6>.n588 0.0557941
R9973 t<6>.n588 t<6>.n587 0.0557941
R9974 t<6>.n587 t<6>.n586 0.0557941
R9975 t<6>.n586 t<6>.n585 0.0557941
R9976 t<6>.n585 t<6>.n584 0.0557941
R9977 t<6>.n583 t<6>.n582 0.0557941
R9978 t<6>.n582 t<6>.n581 0.0557941
R9979 t<6>.n581 t<6>.n580 0.0557941
R9980 t<6>.n580 t<6>.n579 0.0557941
R9981 t<6>.n579 t<6>.n578 0.0557941
R9982 t<6>.n577 t<6>.n576 0.0557941
R9983 t<6>.n576 t<6>.n575 0.0557941
R9984 t<6>.n575 t<6>.n574 0.0557941
R9985 t<6>.n574 t<6>.n573 0.0557941
R9986 t<6>.n573 t<6>.n572 0.0557941
R9987 t<6>.n571 t<6>.n570 0.0557941
R9988 t<6>.n570 t<6>.n569 0.0557941
R9989 t<6>.n569 t<6>.n568 0.0557941
R9990 t<6>.n568 t<6>.n567 0.0557941
R9991 t<6>.n567 t<6>.n566 0.0557941
R9992 t<6>.n565 t<6>.n564 0.0557941
R9993 t<6>.n564 t<6>.n563 0.0557941
R9994 t<6>.n563 t<6>.n562 0.0557941
R9995 t<6>.n562 t<6>.n561 0.0557941
R9996 t<6>.n561 t<6>.n560 0.0557941
R9997 t<6>.n559 t<6>.n558 0.0557941
R9998 t<6>.n558 t<6>.n557 0.0557941
R9999 t<6>.n557 t<6>.n556 0.0557941
R10000 t<6>.n556 t<6>.n555 0.0557941
R10001 t<6>.n555 t<6>.n554 0.0557941
R10002 t<6>.n553 t<6>.n552 0.0557941
R10003 t<6>.n552 t<6>.n551 0.0557941
R10004 t<6>.n551 t<6>.n550 0.0557941
R10005 t<6>.n550 t<6>.n549 0.0557941
R10006 t<6>.n549 t<6>.n548 0.0557941
R10007 t<6>.n547 t<6>.n546 0.0557941
R10008 t<6>.n546 t<6>.n545 0.0557941
R10009 t<6>.n545 t<6>.n544 0.0557941
R10010 t<6>.n544 t<6>.n543 0.0557941
R10011 t<6>.n543 t<6>.n542 0.0557941
R10012 t<6>.n541 t<6>.n540 0.0557941
R10013 t<6>.n540 t<6>.n539 0.0557941
R10014 t<6>.n539 t<6>.n538 0.0557941
R10015 t<6>.n538 t<6>.n537 0.0557941
R10016 t<6>.n537 t<6>.n536 0.0557941
R10017 t<6>.n535 t<6>.n534 0.0557941
R10018 t<6>.n534 t<6>.n533 0.0557941
R10019 t<6>.n533 t<6>.n532 0.0557941
R10020 t<6>.n532 t<6>.n531 0.0557941
R10021 t<6>.n531 t<6>.n530 0.0557941
R10022 t<6>.n529 t<6>.n528 0.0557941
R10023 t<6>.n528 t<6>.n527 0.0557941
R10024 t<6>.n527 t<6>.n526 0.0557941
R10025 t<6>.n526 t<6>.n525 0.0557941
R10026 t<6>.n525 t<6>.n524 0.0557941
R10027 t<6>.n523 t<6>.n522 0.0557941
R10028 t<6>.n522 t<6>.n521 0.0557941
R10029 t<6>.n521 t<6>.n520 0.0557941
R10030 t<6>.n520 t<6>.n519 0.0557941
R10031 t<6>.n519 t<6>.n518 0.0557941
R10032 t<6>.n517 t<6>.n516 0.0557941
R10033 t<6>.n516 t<6>.n515 0.0557941
R10034 t<6>.n515 t<6>.n514 0.0557941
R10035 t<6>.n514 t<6>.n513 0.0557941
R10036 t<6>.n513 t<6>.n512 0.0557941
R10037 t<6>.n511 t<6>.n510 0.0557941
R10038 t<6>.n510 t<6>.n509 0.0557941
R10039 t<6>.n509 t<6>.n508 0.0557941
R10040 t<6>.n508 t<6>.n507 0.0557941
R10041 t<6>.n507 t<6>.n506 0.0557941
R10042 t<6>.n505 t<6>.n504 0.0557941
R10043 t<6>.n504 t<6>.n503 0.0557941
R10044 t<6>.n503 t<6>.n502 0.0557941
R10045 t<6>.n502 t<6>.n501 0.0557941
R10046 t<6>.n501 t<6>.n500 0.0557941
R10047 t<6>.n499 t<6>.n498 0.0557941
R10048 t<6>.n498 t<6>.n497 0.0557941
R10049 t<6>.n497 t<6>.n496 0.0557941
R10050 t<6>.n496 t<6>.n495 0.0557941
R10051 t<6>.n495 t<6>.n494 0.0557941
R10052 t<6>.n493 t<6>.n492 0.0557941
R10053 t<6>.n492 t<6>.n491 0.0557941
R10054 t<6>.n491 t<6>.n490 0.0557941
R10055 t<6>.n490 t<6>.n489 0.0557941
R10056 t<6>.n489 t<6>.n488 0.0557941
R10057 t<6>.n487 t<6>.n486 0.0557941
R10058 t<6>.n486 t<6>.n485 0.0557941
R10059 t<6>.n485 t<6>.n484 0.0557941
R10060 t<6>.n484 t<6>.n483 0.0557941
R10061 t<6>.n483 t<6>.n482 0.0557941
R10062 t<6>.n481 t<6>.n480 0.0557941
R10063 t<6>.n480 t<6>.n479 0.0557941
R10064 t<6>.n479 t<6>.n478 0.0557941
R10065 t<6>.n478 t<6>.n477 0.0557941
R10066 t<6>.n477 t<6>.n476 0.0557941
R10067 t<6>.n475 t<6>.n474 0.0557941
R10068 t<6>.n474 t<6>.n473 0.0557941
R10069 t<6>.n473 t<6>.n472 0.0557941
R10070 t<6>.n472 t<6>.n471 0.0557941
R10071 t<6>.n471 t<6>.n470 0.0557941
R10072 t<6>.n469 t<6>.n468 0.0557941
R10073 t<6>.n468 t<6>.n467 0.0557941
R10074 t<6>.n467 t<6>.n466 0.0557941
R10075 t<6>.n466 t<6>.n465 0.0557941
R10076 t<6>.n465 t<6>.n464 0.0557941
R10077 t<6>.n463 t<6>.n462 0.0557941
R10078 t<6>.n462 t<6>.n461 0.0557941
R10079 t<6>.n461 t<6>.n460 0.0557941
R10080 t<6>.n460 t<6>.n459 0.0557941
R10081 t<6>.n459 t<6>.n458 0.0557941
R10082 t<6>.n457 t<6>.n456 0.0557941
R10083 t<6>.n456 t<6>.n455 0.0557941
R10084 t<6>.n455 t<6>.n454 0.0557941
R10085 t<6>.n454 t<6>.n453 0.0557941
R10086 t<6>.n453 t<6>.n452 0.0557941
R10087 t<6>.n451 t<6>.n450 0.0557941
R10088 t<6>.n450 t<6>.n449 0.0557941
R10089 t<6>.n449 t<6>.n448 0.0557941
R10090 t<6>.n448 t<6>.n447 0.0557941
R10091 t<6>.n447 t<6>.n446 0.0557941
R10092 t<6>.n445 t<6>.n444 0.0557941
R10093 t<6>.n444 t<6>.n443 0.0557941
R10094 t<6>.n443 t<6>.n442 0.0557941
R10095 t<6>.n442 t<6>.n441 0.0557941
R10096 t<6>.n441 t<6>.n440 0.0557941
R10097 t<6>.n439 t<6>.n438 0.0557941
R10098 t<6>.n438 t<6>.n437 0.0557941
R10099 t<6>.n437 t<6>.n436 0.0557941
R10100 t<6>.n436 t<6>.n435 0.0557941
R10101 t<6>.n435 t<6>.n434 0.0557941
R10102 t<6>.n433 t<6>.n432 0.0557941
R10103 t<6>.n432 t<6>.n431 0.0557941
R10104 t<6>.n431 t<6>.n430 0.0557941
R10105 t<6>.n430 t<6>.n429 0.0557941
R10106 t<6>.n429 t<6>.n428 0.0557941
R10107 t<6>.n427 t<6>.n426 0.0557941
R10108 t<6>.n426 t<6>.n425 0.0557941
R10109 t<6>.n425 t<6>.n424 0.0557941
R10110 t<6>.n424 t<6>.n423 0.0557941
R10111 t<6>.n423 t<6>.n422 0.0557941
R10112 t<6>.n421 t<6>.n420 0.0557941
R10113 t<6>.n420 t<6>.n419 0.0557941
R10114 t<6>.n419 t<6>.n418 0.0557941
R10115 t<6>.n418 t<6>.n417 0.0557941
R10116 t<6>.n417 t<6>.n416 0.0557941
R10117 t<6>.n415 t<6>.n414 0.0557941
R10118 t<6>.n414 t<6>.n413 0.0557941
R10119 t<6>.n413 t<6>.n412 0.0557941
R10120 t<6>.n399 t<6>.n398 0.0488824
R10121 t<6>.n9 t<6>.n7 0.0419706
R10122 t<6>.n378 t<6>.n377 0.0419706
R10123 t<6>.n16 t<6>.n14 0.0419706
R10124 t<6>.n359 t<6>.n358 0.0419706
R10125 t<6>.n23 t<6>.n21 0.0419706
R10126 t<6>.n340 t<6>.n339 0.0419706
R10127 t<6>.n30 t<6>.n28 0.0419706
R10128 t<6>.n321 t<6>.n320 0.0419706
R10129 t<6>.n37 t<6>.n35 0.0419706
R10130 t<6>.n302 t<6>.n301 0.0419706
R10131 t<6>.n44 t<6>.n42 0.0419706
R10132 t<6>.n283 t<6>.n282 0.0419706
R10133 t<6>.n51 t<6>.n49 0.0419706
R10134 t<6>.n264 t<6>.n263 0.0419706
R10135 t<6>.n58 t<6>.n56 0.0419706
R10136 t<6>.n245 t<6>.n244 0.0419706
R10137 t<6>.n65 t<6>.n63 0.0419706
R10138 t<6>.n226 t<6>.n225 0.0419706
R10139 t<6>.n72 t<6>.n70 0.0419706
R10140 t<6>.n207 t<6>.n206 0.0419706
R10141 t<6>.n79 t<6>.n77 0.0419706
R10142 t<6>.n188 t<6>.n187 0.0419706
R10143 t<6>.n86 t<6>.n84 0.0419706
R10144 t<6>.n169 t<6>.n168 0.0419706
R10145 t<6>.n93 t<6>.n91 0.0419706
R10146 t<6>.n150 t<6>.n149 0.0419706
R10147 t<6>.n100 t<6>.n98 0.0419706
R10148 t<6>.n131 t<6>.n130 0.0419706
R10149 t<6>.n107 t<6>.n105 0.0419706
R10150 t<6>.n112 t<6>.n111 0.0419706
R10151 t<6>.n408 t<6> 0.0419706
R10152 t<6>.n394 t<6>.n393 0.0405882
R10153 t<6>.n395 t<6>.n5 0.0405882
R10154 t<6>.n593 t<6>.n592 0.0405882
R10155 t<6>.n410 t<6>.n409 0.0405882
R10156 t<6>.n394 t<6>.n3 0.0157059
R10157 t<6>.n594 t<6>.n593 0.0157059
R10158 t<6>.n385 t<6>.n9 0.0143235
R10159 t<6>.n377 t<6>.n376 0.0143235
R10160 t<6>.n366 t<6>.n16 0.0143235
R10161 t<6>.n358 t<6>.n357 0.0143235
R10162 t<6>.n347 t<6>.n23 0.0143235
R10163 t<6>.n339 t<6>.n338 0.0143235
R10164 t<6>.n328 t<6>.n30 0.0143235
R10165 t<6>.n320 t<6>.n319 0.0143235
R10166 t<6>.n309 t<6>.n37 0.0143235
R10167 t<6>.n301 t<6>.n300 0.0143235
R10168 t<6>.n290 t<6>.n44 0.0143235
R10169 t<6>.n282 t<6>.n281 0.0143235
R10170 t<6>.n271 t<6>.n51 0.0143235
R10171 t<6>.n263 t<6>.n262 0.0143235
R10172 t<6>.n252 t<6>.n58 0.0143235
R10173 t<6>.n244 t<6>.n243 0.0143235
R10174 t<6>.n233 t<6>.n65 0.0143235
R10175 t<6>.n225 t<6>.n224 0.0143235
R10176 t<6>.n214 t<6>.n72 0.0143235
R10177 t<6>.n206 t<6>.n205 0.0143235
R10178 t<6>.n195 t<6>.n79 0.0143235
R10179 t<6>.n187 t<6>.n186 0.0143235
R10180 t<6>.n176 t<6>.n86 0.0143235
R10181 t<6>.n168 t<6>.n167 0.0143235
R10182 t<6>.n157 t<6>.n93 0.0143235
R10183 t<6>.n149 t<6>.n148 0.0143235
R10184 t<6>.n138 t<6>.n100 0.0143235
R10185 t<6>.n130 t<6>.n129 0.0143235
R10186 t<6>.n119 t<6>.n107 0.0143235
R10187 t<6>.n409 t<6>.n408 0.0143235
R10188 t<6>.n599 t<6>.n598 0.0100455
R10189 t<6>.n396 t<6>.n395 0.0098016
R10190 t<6>.n411 t<6>.n410 0.0098016
R10191 t<6>.n405 t<6>.n404 0.0089954
R10192 t<6>.n4 t<6>.n2 0.00892479
R10193 t<6>.n597 t<6>.n407 0.00883373
R10194 t<6>.n597 t<6>.n596 0.00783691
R10195 t<6>.n398 t<6>.n3 0.00741176
R10196 t<6>.n595 t<6>.n594 0.00741176
R10197 t<6>.n401 t<6>.n1 0.00606092
R10198 t<6>.n401 t<6>.n400 0.00567797
R10199 t<6>.n400 t<6>.n2 0.00494174
R10200 t<6> t<6>.n599 0.00455166
R10201 t<6>.n402 t<6>.n0 0.00349062
R10202 t<6>.n598 t<6>.n403 0.00347205
R10203 t<6>.n397 t<6>.n4 0.00249153
R10204 t<6>.n397 t<6>.n396 0.00249153
R10205 t<6>.n596 t<6>.n411 0.00249153
R10206 tb<3>.n1 tb<3> 0.255933
R10207 tb<3>.n2 tb<3>.n1 0.207891
R10208 tb<3>.n23 tb<3>.n22 0.204769
R10209 tb<3>.n32 tb<3>.n0 0.201793
R10210 tb<3>.n31 tb<3>.n25 0.185301
R10211 tb<3>.n31 tb<3>.n30 0.177515
R10212 tb<3>.n7 tb<3>.n6 0.142882
R10213 tb<3>.n24 tb<3> 0.119615
R10214 tb<3>.n25 tb<3>.n24 0.118419
R10215 tb<3>.n16 tb<3> 0.108543
R10216 tb<3>.n9 tb<3> 0.0976333
R10217 tb<3>.n2 tb<3> 0.0976333
R10218 tb<3>.n21 tb<3>.n20 0.0876263
R10219 tb<3>.n17 tb<3>.n16 0.0750151
R10220 tb<3>.n19 tb<3>.n18 0.0571765
R10221 tb<3>.n4 tb<3>.n3 0.0557941
R10222 tb<3>.n5 tb<3>.n4 0.0557941
R10223 tb<3>.n6 tb<3>.n5 0.0557941
R10224 tb<3>.n8 tb<3>.n7 0.0557941
R10225 tb<3>.n11 tb<3>.n10 0.0557941
R10226 tb<3>.n12 tb<3>.n11 0.0557941
R10227 tb<3>.n27 tb<3>.n26 0.0468088
R10228 tb<3>.n13 tb<3>.n12 0.0468088
R10229 tb<3>.n20 tb<3>.n15 0.0457975
R10230 tb<3>.n26 tb<3> 0.0419706
R10231 tb<3>.n9 tb<3>.n8 0.0419706
R10232 tb<3>.n30 tb<3>.n29 0.0279692
R10233 tb<3>.n20 tb<3>.n19 0.0215457
R10234 tb<3>.n3 tb<3>.n2 0.0143235
R10235 tb<3>.n10 tb<3>.n9 0.0143235
R10236 tb<3>.n29 tb<3>.n28 0.0136324
R10237 tb<3>.n15 tb<3>.n14 0.0136324
R10238 tb<3>.n18 tb<3>.n17 0.0123976
R10239 tb<3>.n32 tb<3>.n31 0.0100893
R10240 tb<3>.n28 tb<3>.n27 0.00948529
R10241 tb<3>.n14 tb<3>.n13 0.00948529
R10242 tb<3> tb<3>.n32 0.00449597
R10243 tb<3>.n22 tb<3>.n21 0.00349062
R10244 tb<3>.n31 tb<3>.n23 0.00349062
R10245 t<3>.n27 t<3>.n26 3.4105
R10246 t<3>.n28 t<3>.n4 3.4105
R10247 t<3>.n12 t<3>.n9 1.7055
R10248 t<3>.n14 t<3>.n13 1.7055
R10249 t<3>.n15 t<3>.n8 1.7055
R10250 t<3>.n17 t<3>.n16 1.7055
R10251 t<3>.n18 t<3>.n7 1.7055
R10252 t<3>.n20 t<3>.n19 1.7055
R10253 t<3>.n22 t<3>.n6 1.7055
R10254 t<3>.n24 t<3>.n23 1.7055
R10255 t<3>.n25 t<3>.n5 1.7055
R10256 t<3>.n32 t<3>.n31 0.48427
R10257 t<3>.n35 t<3>.n34 0.3805
R10258 t<3>.n30 t<3>.n29 0.3805
R10259 t<3>.n12 t<3>.n11 0.342446
R10260 t<3>.n33 t<3>.n32 0.3424
R10261 t<3>.n11 t<3> 0.255933
R10262 t<3>.n11 t<3>.n10 0.207891
R10263 t<3>.n46 t<3>.n0 0.201793
R10264 t<3>.n3 t<3>.n1 0.185301
R10265 t<3>.n45 t<3>.n39 0.185301
R10266 t<3>.n45 t<3>.n44 0.177515
R10267 t<3>.n18 t<3>.n17 0.142882
R10268 t<3>.n16 t<3>.n7 0.142882
R10269 t<3>.n32 t<3>.n30 0.12975
R10270 t<3>.n36 t<3> 0.123659
R10271 t<3>.n37 t<3> 0.119615
R10272 t<3>.n39 t<3>.n37 0.118419
R10273 t<3>.n31 t<3> 0.108543
R10274 t<3>.n21 t<3> 0.0976333
R10275 t<3>.n10 t<3> 0.0976333
R10276 t<3>.n2 t<3>.n1 0.0876263
R10277 t<3> t<3>.n35 0.0816094
R10278 t<3>.n31 t<3>.n3 0.0750151
R10279 t<3>.n34 t<3>.n33 0.0571765
R10280 t<3>.n13 t<3>.n12 0.0557941
R10281 t<3>.n13 t<3>.n8 0.0557941
R10282 t<3>.n17 t<3>.n8 0.0557941
R10283 t<3>.n19 t<3>.n18 0.0557941
R10284 t<3>.n19 t<3>.n6 0.0557941
R10285 t<3>.n24 t<3>.n6 0.0557941
R10286 t<3>.n25 t<3>.n24 0.0557941
R10287 t<3>.n14 t<3>.n9 0.0557941
R10288 t<3>.n15 t<3>.n14 0.0557941
R10289 t<3>.n16 t<3>.n15 0.0557941
R10290 t<3>.n20 t<3>.n7 0.0557941
R10291 t<3>.n23 t<3>.n22 0.0557941
R10292 t<3>.n23 t<3>.n5 0.0557941
R10293 t<3>.n41 t<3>.n40 0.0468088
R10294 t<3>.n26 t<3>.n25 0.0468088
R10295 t<3>.n27 t<3>.n5 0.0468088
R10296 t<3>.n29 t<3>.n2 0.0457975
R10297 t<3>.n40 t<3> 0.0419706
R10298 t<3>.n21 t<3>.n20 0.0419706
R10299 t<3>.n44 t<3>.n43 0.0279692
R10300 t<3>.n34 t<3>.n2 0.0215457
R10301 t<3>.n10 t<3>.n9 0.0143235
R10302 t<3>.n22 t<3>.n21 0.0143235
R10303 t<3>.n43 t<3>.n42 0.0136324
R10304 t<3>.n30 t<3>.n4 0.0136324
R10305 t<3>.n29 t<3>.n28 0.0136324
R10306 t<3>.n39 t<3>.n38 0.0123976
R10307 t<3>.n33 t<3>.n3 0.0123976
R10308 t<3>.n46 t<3>.n45 0.0100893
R10309 t<3>.n42 t<3>.n41 0.00948529
R10310 t<3>.n26 t<3>.n4 0.00948529
R10311 t<3>.n28 t<3>.n27 0.00948529
R10312 t<3> t<3>.n46 0.00449597
R10313 t<3>.n35 t<3>.n1 0.00349062
R10314 t<3>.n45 t<3>.n36 0.00349062
R10315 t<5>.n191 t<5>.n3 3.4105
R10316 t<5>.n193 t<5>.n192 3.4105
R10317 t<5>.n49 t<5>.n46 1.7055
R10318 t<5>.n51 t<5>.n50 1.7055
R10319 t<5>.n52 t<5>.n45 1.7055
R10320 t<5>.n54 t<5>.n53 1.7055
R10321 t<5>.n55 t<5>.n44 1.7055
R10322 t<5>.n58 t<5>.n57 1.7055
R10323 t<5>.n59 t<5>.n43 1.7055
R10324 t<5>.n61 t<5>.n60 1.7055
R10325 t<5>.n62 t<5>.n42 1.7055
R10326 t<5>.n64 t<5>.n63 1.7055
R10327 t<5>.n65 t<5>.n41 1.7055
R10328 t<5>.n67 t<5>.n66 1.7055
R10329 t<5>.n69 t<5>.n40 1.7055
R10330 t<5>.n71 t<5>.n70 1.7055
R10331 t<5>.n72 t<5>.n39 1.7055
R10332 t<5>.n74 t<5>.n73 1.7055
R10333 t<5>.n75 t<5>.n38 1.7055
R10334 t<5>.n78 t<5>.n77 1.7055
R10335 t<5>.n79 t<5>.n37 1.7055
R10336 t<5>.n81 t<5>.n80 1.7055
R10337 t<5>.n82 t<5>.n36 1.7055
R10338 t<5>.n84 t<5>.n83 1.7055
R10339 t<5>.n85 t<5>.n35 1.7055
R10340 t<5>.n87 t<5>.n86 1.7055
R10341 t<5>.n89 t<5>.n34 1.7055
R10342 t<5>.n91 t<5>.n90 1.7055
R10343 t<5>.n92 t<5>.n33 1.7055
R10344 t<5>.n94 t<5>.n93 1.7055
R10345 t<5>.n95 t<5>.n32 1.7055
R10346 t<5>.n98 t<5>.n97 1.7055
R10347 t<5>.n99 t<5>.n31 1.7055
R10348 t<5>.n101 t<5>.n100 1.7055
R10349 t<5>.n102 t<5>.n30 1.7055
R10350 t<5>.n104 t<5>.n103 1.7055
R10351 t<5>.n105 t<5>.n29 1.7055
R10352 t<5>.n107 t<5>.n106 1.7055
R10353 t<5>.n109 t<5>.n28 1.7055
R10354 t<5>.n111 t<5>.n110 1.7055
R10355 t<5>.n112 t<5>.n27 1.7055
R10356 t<5>.n114 t<5>.n113 1.7055
R10357 t<5>.n115 t<5>.n26 1.7055
R10358 t<5>.n118 t<5>.n117 1.7055
R10359 t<5>.n119 t<5>.n25 1.7055
R10360 t<5>.n121 t<5>.n120 1.7055
R10361 t<5>.n122 t<5>.n24 1.7055
R10362 t<5>.n125 t<5>.n124 1.7055
R10363 t<5>.n126 t<5>.n23 1.7055
R10364 t<5>.n128 t<5>.n127 1.7055
R10365 t<5>.n130 t<5>.n22 1.7055
R10366 t<5>.n132 t<5>.n131 1.7055
R10367 t<5>.n133 t<5>.n21 1.7055
R10368 t<5>.n135 t<5>.n134 1.7055
R10369 t<5>.n136 t<5>.n20 1.7055
R10370 t<5>.n139 t<5>.n138 1.7055
R10371 t<5>.n140 t<5>.n19 1.7055
R10372 t<5>.n142 t<5>.n141 1.7055
R10373 t<5>.n143 t<5>.n18 1.7055
R10374 t<5>.n145 t<5>.n144 1.7055
R10375 t<5>.n146 t<5>.n17 1.7055
R10376 t<5>.n148 t<5>.n147 1.7055
R10377 t<5>.n150 t<5>.n16 1.7055
R10378 t<5>.n152 t<5>.n151 1.7055
R10379 t<5>.n153 t<5>.n15 1.7055
R10380 t<5>.n155 t<5>.n154 1.7055
R10381 t<5>.n156 t<5>.n14 1.7055
R10382 t<5>.n159 t<5>.n158 1.7055
R10383 t<5>.n160 t<5>.n13 1.7055
R10384 t<5>.n162 t<5>.n161 1.7055
R10385 t<5>.n163 t<5>.n12 1.7055
R10386 t<5>.n165 t<5>.n164 1.7055
R10387 t<5>.n166 t<5>.n11 1.7055
R10388 t<5>.n168 t<5>.n167 1.7055
R10389 t<5>.n170 t<5>.n10 1.7055
R10390 t<5>.n172 t<5>.n171 1.7055
R10391 t<5>.n173 t<5>.n9 1.7055
R10392 t<5>.n175 t<5>.n174 1.7055
R10393 t<5>.n176 t<5>.n8 1.7055
R10394 t<5>.n178 t<5>.n177 1.7055
R10395 t<5>.n180 t<5>.n179 1.7055
R10396 t<5>.n181 t<5>.n6 1.7055
R10397 t<5>.n183 t<5>.n182 1.7055
R10398 t<5>.n184 t<5>.n5 1.7055
R10399 t<5>.n186 t<5>.n185 1.7055
R10400 t<5>.n187 t<5>.n4 1.7055
R10401 t<5>.n190 t<5>.n189 1.7055
R10402 t<5>.n123 t<5> 0.746233
R10403 t<5>.n198 t<5>.n197 0.397694
R10404 t<5>.n200 t<5>.n199 0.3805
R10405 t<5>.n194 t<5>.n2 0.3805
R10406 t<5>.n389 t<5>.n388 0.3805
R10407 t<5>.n47 t<5>.n46 0.342446
R10408 t<5>.n197 t<5>.n196 0.3424
R10409 t<5>.n394 t<5>.n393 0.3424
R10410 t<5>.n47 t<5> 0.255933
R10411 t<5>.n202 t<5> 0.24623
R10412 t<5>.n48 t<5>.n47 0.207891
R10413 t<5>.n198 t<5>.n0 0.193586
R10414 t<5>.n203 t<5>.n202 0.17426
R10415 t<5>.n305 t<5>.n304 0.142882
R10416 t<5>.n311 t<5>.n310 0.142882
R10417 t<5>.n317 t<5>.n316 0.142882
R10418 t<5>.n323 t<5>.n322 0.142882
R10419 t<5>.n329 t<5>.n328 0.142882
R10420 t<5>.n335 t<5>.n334 0.142882
R10421 t<5>.n341 t<5>.n340 0.142882
R10422 t<5>.n347 t<5>.n346 0.142882
R10423 t<5>.n353 t<5>.n352 0.142882
R10424 t<5>.n359 t<5>.n358 0.142882
R10425 t<5>.n365 t<5>.n364 0.142882
R10426 t<5>.n371 t<5>.n370 0.142882
R10427 t<5>.n377 t<5>.n376 0.142882
R10428 t<5>.n383 t<5>.n382 0.142882
R10429 t<5>.n206 t<5>.n205 0.142882
R10430 t<5>.n213 t<5>.n212 0.142882
R10431 t<5>.n220 t<5>.n219 0.142882
R10432 t<5>.n227 t<5>.n226 0.142882
R10433 t<5>.n234 t<5>.n233 0.142882
R10434 t<5>.n241 t<5>.n240 0.142882
R10435 t<5>.n248 t<5>.n247 0.142882
R10436 t<5>.n255 t<5>.n254 0.142882
R10437 t<5>.n262 t<5>.n261 0.142882
R10438 t<5>.n269 t<5>.n268 0.142882
R10439 t<5>.n276 t<5>.n275 0.142882
R10440 t<5>.n283 t<5>.n282 0.142882
R10441 t<5>.n290 t<5>.n289 0.142882
R10442 t<5>.n297 t<5>.n296 0.142882
R10443 t<5>.n53 t<5>.n44 0.142882
R10444 t<5>.n65 t<5>.n64 0.142882
R10445 t<5>.n73 t<5>.n38 0.142882
R10446 t<5>.n85 t<5>.n84 0.142882
R10447 t<5>.n93 t<5>.n32 0.142882
R10448 t<5>.n105 t<5>.n104 0.142882
R10449 t<5>.n113 t<5>.n26 0.142882
R10450 t<5>.n126 t<5>.n125 0.142882
R10451 t<5>.n134 t<5>.n20 0.142882
R10452 t<5>.n146 t<5>.n145 0.142882
R10453 t<5>.n154 t<5>.n14 0.142882
R10454 t<5>.n166 t<5>.n165 0.142882
R10455 t<5>.n174 t<5>.n8 0.142882
R10456 t<5>.n185 t<5>.n184 0.142882
R10457 t<5>.n55 t<5>.n54 0.142882
R10458 t<5>.n63 t<5>.n41 0.142882
R10459 t<5>.n75 t<5>.n74 0.142882
R10460 t<5>.n83 t<5>.n35 0.142882
R10461 t<5>.n95 t<5>.n94 0.142882
R10462 t<5>.n103 t<5>.n29 0.142882
R10463 t<5>.n115 t<5>.n114 0.142882
R10464 t<5>.n124 t<5>.n23 0.142882
R10465 t<5>.n136 t<5>.n135 0.142882
R10466 t<5>.n144 t<5>.n17 0.142882
R10467 t<5>.n156 t<5>.n155 0.142882
R10468 t<5>.n164 t<5>.n11 0.142882
R10469 t<5>.n176 t<5>.n175 0.142882
R10470 t<5>.n186 t<5>.n5 0.142882
R10471 t<5>.n1 t<5>.n0 0.130613
R10472 t<5>.n201 t<5> 0.125653
R10473 t<5>.n195 t<5>.n0 0.125385
R10474 t<5>.n396 t<5>.n395 0.119792
R10475 t<5>.n188 t<5> 0.0976333
R10476 t<5>.n7 t<5> 0.0976333
R10477 t<5>.n169 t<5> 0.0976333
R10478 t<5>.n157 t<5> 0.0976333
R10479 t<5>.n149 t<5> 0.0976333
R10480 t<5>.n137 t<5> 0.0976333
R10481 t<5>.n129 t<5> 0.0976333
R10482 t<5>.n116 t<5> 0.0976333
R10483 t<5>.n108 t<5> 0.0976333
R10484 t<5>.n96 t<5> 0.0976333
R10485 t<5>.n88 t<5> 0.0976333
R10486 t<5>.n76 t<5> 0.0976333
R10487 t<5>.n68 t<5> 0.0976333
R10488 t<5>.n56 t<5> 0.0976333
R10489 t<5>.n48 t<5> 0.0976333
R10490 t<5> t<5>.n200 0.0796156
R10491 t<5>.n203 t<5> 0.0725667
R10492 t<5>.n210 t<5> 0.0725667
R10493 t<5>.n217 t<5> 0.0725667
R10494 t<5>.n224 t<5> 0.0725667
R10495 t<5>.n231 t<5> 0.0725667
R10496 t<5>.n238 t<5> 0.0725667
R10497 t<5>.n245 t<5> 0.0725667
R10498 t<5>.n252 t<5> 0.0725667
R10499 t<5>.n259 t<5> 0.0725667
R10500 t<5>.n266 t<5> 0.0725667
R10501 t<5>.n273 t<5> 0.0725667
R10502 t<5>.n280 t<5> 0.0725667
R10503 t<5>.n287 t<5> 0.0725667
R10504 t<5>.n294 t<5> 0.0725667
R10505 t<5>.n302 t<5> 0.0725667
R10506 t<5>.n304 t<5>.n303 0.0557941
R10507 t<5>.n306 t<5>.n305 0.0557941
R10508 t<5>.n307 t<5>.n306 0.0557941
R10509 t<5>.n308 t<5>.n307 0.0557941
R10510 t<5>.n309 t<5>.n308 0.0557941
R10511 t<5>.n310 t<5>.n309 0.0557941
R10512 t<5>.n312 t<5>.n311 0.0557941
R10513 t<5>.n313 t<5>.n312 0.0557941
R10514 t<5>.n314 t<5>.n313 0.0557941
R10515 t<5>.n315 t<5>.n314 0.0557941
R10516 t<5>.n316 t<5>.n315 0.0557941
R10517 t<5>.n318 t<5>.n317 0.0557941
R10518 t<5>.n319 t<5>.n318 0.0557941
R10519 t<5>.n320 t<5>.n319 0.0557941
R10520 t<5>.n321 t<5>.n320 0.0557941
R10521 t<5>.n322 t<5>.n321 0.0557941
R10522 t<5>.n324 t<5>.n323 0.0557941
R10523 t<5>.n325 t<5>.n324 0.0557941
R10524 t<5>.n326 t<5>.n325 0.0557941
R10525 t<5>.n327 t<5>.n326 0.0557941
R10526 t<5>.n328 t<5>.n327 0.0557941
R10527 t<5>.n330 t<5>.n329 0.0557941
R10528 t<5>.n331 t<5>.n330 0.0557941
R10529 t<5>.n332 t<5>.n331 0.0557941
R10530 t<5>.n333 t<5>.n332 0.0557941
R10531 t<5>.n334 t<5>.n333 0.0557941
R10532 t<5>.n336 t<5>.n335 0.0557941
R10533 t<5>.n337 t<5>.n336 0.0557941
R10534 t<5>.n338 t<5>.n337 0.0557941
R10535 t<5>.n339 t<5>.n338 0.0557941
R10536 t<5>.n340 t<5>.n339 0.0557941
R10537 t<5>.n342 t<5>.n341 0.0557941
R10538 t<5>.n343 t<5>.n342 0.0557941
R10539 t<5>.n344 t<5>.n343 0.0557941
R10540 t<5>.n345 t<5>.n344 0.0557941
R10541 t<5>.n346 t<5>.n345 0.0557941
R10542 t<5>.n348 t<5>.n347 0.0557941
R10543 t<5>.n349 t<5>.n348 0.0557941
R10544 t<5>.n350 t<5>.n349 0.0557941
R10545 t<5>.n351 t<5>.n350 0.0557941
R10546 t<5>.n352 t<5>.n351 0.0557941
R10547 t<5>.n354 t<5>.n353 0.0557941
R10548 t<5>.n355 t<5>.n354 0.0557941
R10549 t<5>.n356 t<5>.n355 0.0557941
R10550 t<5>.n357 t<5>.n356 0.0557941
R10551 t<5>.n358 t<5>.n357 0.0557941
R10552 t<5>.n360 t<5>.n359 0.0557941
R10553 t<5>.n361 t<5>.n360 0.0557941
R10554 t<5>.n362 t<5>.n361 0.0557941
R10555 t<5>.n363 t<5>.n362 0.0557941
R10556 t<5>.n364 t<5>.n363 0.0557941
R10557 t<5>.n366 t<5>.n365 0.0557941
R10558 t<5>.n367 t<5>.n366 0.0557941
R10559 t<5>.n368 t<5>.n367 0.0557941
R10560 t<5>.n369 t<5>.n368 0.0557941
R10561 t<5>.n370 t<5>.n369 0.0557941
R10562 t<5>.n372 t<5>.n371 0.0557941
R10563 t<5>.n373 t<5>.n372 0.0557941
R10564 t<5>.n374 t<5>.n373 0.0557941
R10565 t<5>.n375 t<5>.n374 0.0557941
R10566 t<5>.n376 t<5>.n375 0.0557941
R10567 t<5>.n378 t<5>.n377 0.0557941
R10568 t<5>.n379 t<5>.n378 0.0557941
R10569 t<5>.n380 t<5>.n379 0.0557941
R10570 t<5>.n381 t<5>.n380 0.0557941
R10571 t<5>.n382 t<5>.n381 0.0557941
R10572 t<5>.n384 t<5>.n383 0.0557941
R10573 t<5>.n385 t<5>.n384 0.0557941
R10574 t<5>.n205 t<5>.n204 0.0557941
R10575 t<5>.n207 t<5>.n206 0.0557941
R10576 t<5>.n208 t<5>.n207 0.0557941
R10577 t<5>.n209 t<5>.n208 0.0557941
R10578 t<5>.n212 t<5>.n211 0.0557941
R10579 t<5>.n214 t<5>.n213 0.0557941
R10580 t<5>.n215 t<5>.n214 0.0557941
R10581 t<5>.n216 t<5>.n215 0.0557941
R10582 t<5>.n219 t<5>.n218 0.0557941
R10583 t<5>.n221 t<5>.n220 0.0557941
R10584 t<5>.n222 t<5>.n221 0.0557941
R10585 t<5>.n223 t<5>.n222 0.0557941
R10586 t<5>.n226 t<5>.n225 0.0557941
R10587 t<5>.n228 t<5>.n227 0.0557941
R10588 t<5>.n229 t<5>.n228 0.0557941
R10589 t<5>.n230 t<5>.n229 0.0557941
R10590 t<5>.n233 t<5>.n232 0.0557941
R10591 t<5>.n235 t<5>.n234 0.0557941
R10592 t<5>.n236 t<5>.n235 0.0557941
R10593 t<5>.n237 t<5>.n236 0.0557941
R10594 t<5>.n240 t<5>.n239 0.0557941
R10595 t<5>.n242 t<5>.n241 0.0557941
R10596 t<5>.n243 t<5>.n242 0.0557941
R10597 t<5>.n244 t<5>.n243 0.0557941
R10598 t<5>.n247 t<5>.n246 0.0557941
R10599 t<5>.n249 t<5>.n248 0.0557941
R10600 t<5>.n250 t<5>.n249 0.0557941
R10601 t<5>.n251 t<5>.n250 0.0557941
R10602 t<5>.n254 t<5>.n253 0.0557941
R10603 t<5>.n256 t<5>.n255 0.0557941
R10604 t<5>.n257 t<5>.n256 0.0557941
R10605 t<5>.n258 t<5>.n257 0.0557941
R10606 t<5>.n261 t<5>.n260 0.0557941
R10607 t<5>.n263 t<5>.n262 0.0557941
R10608 t<5>.n264 t<5>.n263 0.0557941
R10609 t<5>.n265 t<5>.n264 0.0557941
R10610 t<5>.n268 t<5>.n267 0.0557941
R10611 t<5>.n270 t<5>.n269 0.0557941
R10612 t<5>.n271 t<5>.n270 0.0557941
R10613 t<5>.n272 t<5>.n271 0.0557941
R10614 t<5>.n275 t<5>.n274 0.0557941
R10615 t<5>.n277 t<5>.n276 0.0557941
R10616 t<5>.n278 t<5>.n277 0.0557941
R10617 t<5>.n279 t<5>.n278 0.0557941
R10618 t<5>.n282 t<5>.n281 0.0557941
R10619 t<5>.n284 t<5>.n283 0.0557941
R10620 t<5>.n285 t<5>.n284 0.0557941
R10621 t<5>.n286 t<5>.n285 0.0557941
R10622 t<5>.n289 t<5>.n288 0.0557941
R10623 t<5>.n291 t<5>.n290 0.0557941
R10624 t<5>.n292 t<5>.n291 0.0557941
R10625 t<5>.n293 t<5>.n292 0.0557941
R10626 t<5>.n296 t<5>.n295 0.0557941
R10627 t<5>.n298 t<5>.n297 0.0557941
R10628 t<5>.n299 t<5>.n298 0.0557941
R10629 t<5>.n51 t<5>.n46 0.0557941
R10630 t<5>.n52 t<5>.n51 0.0557941
R10631 t<5>.n53 t<5>.n52 0.0557941
R10632 t<5>.n58 t<5>.n44 0.0557941
R10633 t<5>.n59 t<5>.n58 0.0557941
R10634 t<5>.n60 t<5>.n59 0.0557941
R10635 t<5>.n60 t<5>.n42 0.0557941
R10636 t<5>.n64 t<5>.n42 0.0557941
R10637 t<5>.n66 t<5>.n65 0.0557941
R10638 t<5>.n66 t<5>.n40 0.0557941
R10639 t<5>.n71 t<5>.n40 0.0557941
R10640 t<5>.n72 t<5>.n71 0.0557941
R10641 t<5>.n73 t<5>.n72 0.0557941
R10642 t<5>.n78 t<5>.n38 0.0557941
R10643 t<5>.n79 t<5>.n78 0.0557941
R10644 t<5>.n80 t<5>.n79 0.0557941
R10645 t<5>.n80 t<5>.n36 0.0557941
R10646 t<5>.n84 t<5>.n36 0.0557941
R10647 t<5>.n86 t<5>.n85 0.0557941
R10648 t<5>.n86 t<5>.n34 0.0557941
R10649 t<5>.n91 t<5>.n34 0.0557941
R10650 t<5>.n92 t<5>.n91 0.0557941
R10651 t<5>.n93 t<5>.n92 0.0557941
R10652 t<5>.n98 t<5>.n32 0.0557941
R10653 t<5>.n99 t<5>.n98 0.0557941
R10654 t<5>.n100 t<5>.n99 0.0557941
R10655 t<5>.n100 t<5>.n30 0.0557941
R10656 t<5>.n104 t<5>.n30 0.0557941
R10657 t<5>.n106 t<5>.n105 0.0557941
R10658 t<5>.n106 t<5>.n28 0.0557941
R10659 t<5>.n111 t<5>.n28 0.0557941
R10660 t<5>.n112 t<5>.n111 0.0557941
R10661 t<5>.n113 t<5>.n112 0.0557941
R10662 t<5>.n118 t<5>.n26 0.0557941
R10663 t<5>.n119 t<5>.n118 0.0557941
R10664 t<5>.n120 t<5>.n119 0.0557941
R10665 t<5>.n120 t<5>.n24 0.0557941
R10666 t<5>.n125 t<5>.n24 0.0557941
R10667 t<5>.n127 t<5>.n126 0.0557941
R10668 t<5>.n127 t<5>.n22 0.0557941
R10669 t<5>.n132 t<5>.n22 0.0557941
R10670 t<5>.n133 t<5>.n132 0.0557941
R10671 t<5>.n134 t<5>.n133 0.0557941
R10672 t<5>.n139 t<5>.n20 0.0557941
R10673 t<5>.n140 t<5>.n139 0.0557941
R10674 t<5>.n141 t<5>.n140 0.0557941
R10675 t<5>.n141 t<5>.n18 0.0557941
R10676 t<5>.n145 t<5>.n18 0.0557941
R10677 t<5>.n147 t<5>.n146 0.0557941
R10678 t<5>.n147 t<5>.n16 0.0557941
R10679 t<5>.n152 t<5>.n16 0.0557941
R10680 t<5>.n153 t<5>.n152 0.0557941
R10681 t<5>.n154 t<5>.n153 0.0557941
R10682 t<5>.n159 t<5>.n14 0.0557941
R10683 t<5>.n160 t<5>.n159 0.0557941
R10684 t<5>.n161 t<5>.n160 0.0557941
R10685 t<5>.n161 t<5>.n12 0.0557941
R10686 t<5>.n165 t<5>.n12 0.0557941
R10687 t<5>.n167 t<5>.n166 0.0557941
R10688 t<5>.n167 t<5>.n10 0.0557941
R10689 t<5>.n172 t<5>.n10 0.0557941
R10690 t<5>.n173 t<5>.n172 0.0557941
R10691 t<5>.n174 t<5>.n173 0.0557941
R10692 t<5>.n178 t<5>.n8 0.0557941
R10693 t<5>.n179 t<5>.n178 0.0557941
R10694 t<5>.n179 t<5>.n6 0.0557941
R10695 t<5>.n183 t<5>.n6 0.0557941
R10696 t<5>.n184 t<5>.n183 0.0557941
R10697 t<5>.n185 t<5>.n4 0.0557941
R10698 t<5>.n190 t<5>.n4 0.0557941
R10699 t<5>.n50 t<5>.n49 0.0557941
R10700 t<5>.n50 t<5>.n45 0.0557941
R10701 t<5>.n54 t<5>.n45 0.0557941
R10702 t<5>.n57 t<5>.n55 0.0557941
R10703 t<5>.n61 t<5>.n43 0.0557941
R10704 t<5>.n62 t<5>.n61 0.0557941
R10705 t<5>.n63 t<5>.n62 0.0557941
R10706 t<5>.n67 t<5>.n41 0.0557941
R10707 t<5>.n70 t<5>.n69 0.0557941
R10708 t<5>.n70 t<5>.n39 0.0557941
R10709 t<5>.n74 t<5>.n39 0.0557941
R10710 t<5>.n77 t<5>.n75 0.0557941
R10711 t<5>.n81 t<5>.n37 0.0557941
R10712 t<5>.n82 t<5>.n81 0.0557941
R10713 t<5>.n83 t<5>.n82 0.0557941
R10714 t<5>.n87 t<5>.n35 0.0557941
R10715 t<5>.n90 t<5>.n89 0.0557941
R10716 t<5>.n90 t<5>.n33 0.0557941
R10717 t<5>.n94 t<5>.n33 0.0557941
R10718 t<5>.n97 t<5>.n95 0.0557941
R10719 t<5>.n101 t<5>.n31 0.0557941
R10720 t<5>.n102 t<5>.n101 0.0557941
R10721 t<5>.n103 t<5>.n102 0.0557941
R10722 t<5>.n107 t<5>.n29 0.0557941
R10723 t<5>.n110 t<5>.n109 0.0557941
R10724 t<5>.n110 t<5>.n27 0.0557941
R10725 t<5>.n114 t<5>.n27 0.0557941
R10726 t<5>.n117 t<5>.n115 0.0557941
R10727 t<5>.n121 t<5>.n25 0.0557941
R10728 t<5>.n122 t<5>.n121 0.0557941
R10729 t<5>.n128 t<5>.n23 0.0557941
R10730 t<5>.n131 t<5>.n130 0.0557941
R10731 t<5>.n131 t<5>.n21 0.0557941
R10732 t<5>.n135 t<5>.n21 0.0557941
R10733 t<5>.n138 t<5>.n136 0.0557941
R10734 t<5>.n142 t<5>.n19 0.0557941
R10735 t<5>.n143 t<5>.n142 0.0557941
R10736 t<5>.n144 t<5>.n143 0.0557941
R10737 t<5>.n148 t<5>.n17 0.0557941
R10738 t<5>.n151 t<5>.n150 0.0557941
R10739 t<5>.n151 t<5>.n15 0.0557941
R10740 t<5>.n155 t<5>.n15 0.0557941
R10741 t<5>.n158 t<5>.n156 0.0557941
R10742 t<5>.n162 t<5>.n13 0.0557941
R10743 t<5>.n163 t<5>.n162 0.0557941
R10744 t<5>.n164 t<5>.n163 0.0557941
R10745 t<5>.n168 t<5>.n11 0.0557941
R10746 t<5>.n171 t<5>.n170 0.0557941
R10747 t<5>.n171 t<5>.n9 0.0557941
R10748 t<5>.n175 t<5>.n9 0.0557941
R10749 t<5>.n177 t<5>.n176 0.0557941
R10750 t<5>.n181 t<5>.n180 0.0557941
R10751 t<5>.n182 t<5>.n181 0.0557941
R10752 t<5>.n182 t<5>.n5 0.0557941
R10753 t<5>.n187 t<5>.n186 0.0557941
R10754 t<5>.n386 t<5>.n385 0.0509559
R10755 t<5>.n300 t<5>.n299 0.0509559
R10756 t<5>.n191 t<5>.n190 0.0509559
R10757 t<5>.n189 t<5>.n3 0.0509559
R10758 t<5>.n204 t<5>.n203 0.0419706
R10759 t<5>.n211 t<5>.n210 0.0419706
R10760 t<5>.n218 t<5>.n217 0.0419706
R10761 t<5>.n225 t<5>.n224 0.0419706
R10762 t<5>.n232 t<5>.n231 0.0419706
R10763 t<5>.n239 t<5>.n238 0.0419706
R10764 t<5>.n246 t<5>.n245 0.0419706
R10765 t<5>.n253 t<5>.n252 0.0419706
R10766 t<5>.n260 t<5>.n259 0.0419706
R10767 t<5>.n267 t<5>.n266 0.0419706
R10768 t<5>.n274 t<5>.n273 0.0419706
R10769 t<5>.n281 t<5>.n280 0.0419706
R10770 t<5>.n288 t<5>.n287 0.0419706
R10771 t<5>.n295 t<5>.n294 0.0419706
R10772 t<5>.n57 t<5>.n56 0.0419706
R10773 t<5>.n68 t<5>.n67 0.0419706
R10774 t<5>.n77 t<5>.n76 0.0419706
R10775 t<5>.n88 t<5>.n87 0.0419706
R10776 t<5>.n97 t<5>.n96 0.0419706
R10777 t<5>.n108 t<5>.n107 0.0419706
R10778 t<5>.n117 t<5>.n116 0.0419706
R10779 t<5>.n123 t<5>.n122 0.0419706
R10780 t<5>.n129 t<5>.n128 0.0419706
R10781 t<5>.n138 t<5>.n137 0.0419706
R10782 t<5>.n149 t<5>.n148 0.0419706
R10783 t<5>.n158 t<5>.n157 0.0419706
R10784 t<5>.n169 t<5>.n168 0.0419706
R10785 t<5>.n177 t<5>.n7 0.0419706
R10786 t<5>.n188 t<5>.n187 0.0419706
R10787 t<5>.n197 t<5>.n2 0.0385147
R10788 t<5>.n394 t<5>.n392 0.0281471
R10789 t<5>.n395 t<5>.n394 0.0220232
R10790 t<5>.n388 t<5>.n387 0.0177794
R10791 t<5>.n192 t<5>.n2 0.0177794
R10792 t<5>.n391 t<5>.n390 0.0170882
R10793 t<5>.n395 t<5>.n389 0.0170118
R10794 t<5>.n210 t<5>.n209 0.0143235
R10795 t<5>.n217 t<5>.n216 0.0143235
R10796 t<5>.n224 t<5>.n223 0.0143235
R10797 t<5>.n231 t<5>.n230 0.0143235
R10798 t<5>.n238 t<5>.n237 0.0143235
R10799 t<5>.n245 t<5>.n244 0.0143235
R10800 t<5>.n252 t<5>.n251 0.0143235
R10801 t<5>.n259 t<5>.n258 0.0143235
R10802 t<5>.n266 t<5>.n265 0.0143235
R10803 t<5>.n273 t<5>.n272 0.0143235
R10804 t<5>.n280 t<5>.n279 0.0143235
R10805 t<5>.n287 t<5>.n286 0.0143235
R10806 t<5>.n294 t<5>.n293 0.0143235
R10807 t<5>.n302 t<5>.n301 0.0143235
R10808 t<5>.n49 t<5>.n48 0.0143235
R10809 t<5>.n56 t<5>.n43 0.0143235
R10810 t<5>.n69 t<5>.n68 0.0143235
R10811 t<5>.n76 t<5>.n37 0.0143235
R10812 t<5>.n89 t<5>.n88 0.0143235
R10813 t<5>.n96 t<5>.n31 0.0143235
R10814 t<5>.n109 t<5>.n108 0.0143235
R10815 t<5>.n116 t<5>.n25 0.0143235
R10816 t<5>.n124 t<5>.n123 0.0143235
R10817 t<5>.n130 t<5>.n129 0.0143235
R10818 t<5>.n137 t<5>.n19 0.0143235
R10819 t<5>.n150 t<5>.n149 0.0143235
R10820 t<5>.n157 t<5>.n13 0.0143235
R10821 t<5>.n170 t<5>.n169 0.0143235
R10822 t<5>.n180 t<5>.n7 0.0143235
R10823 t<5>.n189 t<5>.n188 0.0143235
R10824 t<5>.n194 t<5>.n193 0.0138432
R10825 t<5>.n392 t<5>.n391 0.0115588
R10826 t<5>.n196 t<5>.n1 0.0110482
R10827 t<5>.n397 t<5>.n396 0.0100893
R10828 t<5>.n196 t<5>.n195 0.00752478
R10829 t<5>.n195 t<5>.n194 0.006246
R10830 t<5>.n387 t<5>.n386 0.00533824
R10831 t<5>.n301 t<5>.n300 0.00533824
R10832 t<5>.n192 t<5>.n191 0.00533824
R10833 t<5>.n193 t<5>.n3 0.00533824
R10834 t<5>.n199 t<5>.n198 0.00527966
R10835 t<5> t<5>.n397 0.00503972
R10836 t<5>.n389 t<5>.n302 0.00395588
R10837 t<5>.n200 t<5>.n0 0.00349062
R10838 t<5>.n396 t<5>.n201 0.00349062
R10839 t<5>.n199 t<5>.n1 0.00208685
R10840 tb<1> tb<1>.n4 0.546915
R10841 tb<1>.n4 tb<1>.n3 0.191835
R10842 tb<1>.n3 tb<1>.n2 0.190255
R10843 tb<1>.n1 tb<1>.n0 0.190195
R10844 tb<1>.n1 tb<1> 0.145828
R10845 tb<1>.n3 tb<1>.n1 0.0214975
R10846 tb<1>.n2 tb<1> 0.0101926
R10847 tb<1>.n2 tb<1>.n0 0.0101019
R10848 tb<1>.n4 tb<1>.n0 0.00250189
R10849 t<1>.n4 t<1>.n3 0.190255
R10850 t<1>.n2 t<1>.n0 0.190195
R10851 t<1>.n0 t<1> 0.145828
R10852 t<1>.n1 t<1> 0.122193
R10853 t<1> t<1>.n4 0.0101926
R10854 t<1>.n4 t<1>.n2 0.0101019
R10855 t<1>.n2 t<1>.n1 0.00250189
R10856 tb<4>.n0 tb<4> 0.255933
R10857 tb<4>.n52 tb<4> 0.24623
R10858 tb<4>.n1 tb<4>.n0 0.207891
R10859 tb<4>.n51 tb<4>.n50 0.204769
R10860 tb<4>.n53 tb<4>.n52 0.17426
R10861 tb<4>.n56 tb<4>.n55 0.142882
R10862 tb<4>.n63 tb<4>.n62 0.142882
R10863 tb<4>.n70 tb<4>.n69 0.142882
R10864 tb<4>.n77 tb<4>.n76 0.142882
R10865 tb<4>.n84 tb<4>.n83 0.142882
R10866 tb<4>.n91 tb<4>.n90 0.142882
R10867 tb<4>.n6 tb<4>.n5 0.142882
R10868 tb<4>.n13 tb<4>.n12 0.142882
R10869 tb<4>.n20 tb<4>.n19 0.142882
R10870 tb<4>.n27 tb<4>.n26 0.142882
R10871 tb<4>.n34 tb<4>.n33 0.142882
R10872 tb<4>.n41 tb<4>.n40 0.142882
R10873 tb<4>.n49 tb<4>.n48 0.125385
R10874 tb<4>.n98 tb<4>.n97 0.119792
R10875 tb<4>.n43 tb<4> 0.0976333
R10876 tb<4>.n36 tb<4> 0.0976333
R10877 tb<4>.n29 tb<4> 0.0976333
R10878 tb<4>.n22 tb<4> 0.0976333
R10879 tb<4>.n15 tb<4> 0.0976333
R10880 tb<4>.n8 tb<4> 0.0976333
R10881 tb<4>.n1 tb<4> 0.0976333
R10882 tb<4>.n53 tb<4> 0.0725667
R10883 tb<4>.n60 tb<4> 0.0725667
R10884 tb<4>.n67 tb<4> 0.0725667
R10885 tb<4>.n74 tb<4> 0.0725667
R10886 tb<4>.n81 tb<4> 0.0725667
R10887 tb<4>.n88 tb<4> 0.0725667
R10888 tb<4>.n55 tb<4>.n54 0.0557941
R10889 tb<4>.n57 tb<4>.n56 0.0557941
R10890 tb<4>.n58 tb<4>.n57 0.0557941
R10891 tb<4>.n59 tb<4>.n58 0.0557941
R10892 tb<4>.n62 tb<4>.n61 0.0557941
R10893 tb<4>.n64 tb<4>.n63 0.0557941
R10894 tb<4>.n65 tb<4>.n64 0.0557941
R10895 tb<4>.n66 tb<4>.n65 0.0557941
R10896 tb<4>.n69 tb<4>.n68 0.0557941
R10897 tb<4>.n71 tb<4>.n70 0.0557941
R10898 tb<4>.n72 tb<4>.n71 0.0557941
R10899 tb<4>.n73 tb<4>.n72 0.0557941
R10900 tb<4>.n76 tb<4>.n75 0.0557941
R10901 tb<4>.n78 tb<4>.n77 0.0557941
R10902 tb<4>.n79 tb<4>.n78 0.0557941
R10903 tb<4>.n80 tb<4>.n79 0.0557941
R10904 tb<4>.n83 tb<4>.n82 0.0557941
R10905 tb<4>.n85 tb<4>.n84 0.0557941
R10906 tb<4>.n86 tb<4>.n85 0.0557941
R10907 tb<4>.n87 tb<4>.n86 0.0557941
R10908 tb<4>.n90 tb<4>.n89 0.0557941
R10909 tb<4>.n92 tb<4>.n91 0.0557941
R10910 tb<4>.n93 tb<4>.n92 0.0557941
R10911 tb<4>.n3 tb<4>.n2 0.0557941
R10912 tb<4>.n4 tb<4>.n3 0.0557941
R10913 tb<4>.n5 tb<4>.n4 0.0557941
R10914 tb<4>.n7 tb<4>.n6 0.0557941
R10915 tb<4>.n10 tb<4>.n9 0.0557941
R10916 tb<4>.n11 tb<4>.n10 0.0557941
R10917 tb<4>.n12 tb<4>.n11 0.0557941
R10918 tb<4>.n14 tb<4>.n13 0.0557941
R10919 tb<4>.n17 tb<4>.n16 0.0557941
R10920 tb<4>.n18 tb<4>.n17 0.0557941
R10921 tb<4>.n19 tb<4>.n18 0.0557941
R10922 tb<4>.n21 tb<4>.n20 0.0557941
R10923 tb<4>.n24 tb<4>.n23 0.0557941
R10924 tb<4>.n25 tb<4>.n24 0.0557941
R10925 tb<4>.n26 tb<4>.n25 0.0557941
R10926 tb<4>.n28 tb<4>.n27 0.0557941
R10927 tb<4>.n31 tb<4>.n30 0.0557941
R10928 tb<4>.n32 tb<4>.n31 0.0557941
R10929 tb<4>.n33 tb<4>.n32 0.0557941
R10930 tb<4>.n35 tb<4>.n34 0.0557941
R10931 tb<4>.n38 tb<4>.n37 0.0557941
R10932 tb<4>.n39 tb<4>.n38 0.0557941
R10933 tb<4>.n40 tb<4>.n39 0.0557941
R10934 tb<4>.n42 tb<4>.n41 0.0557941
R10935 tb<4>.n94 tb<4>.n93 0.0509559
R10936 tb<4>.n45 tb<4>.n44 0.0509559
R10937 tb<4>.n54 tb<4>.n53 0.0419706
R10938 tb<4>.n61 tb<4>.n60 0.0419706
R10939 tb<4>.n68 tb<4>.n67 0.0419706
R10940 tb<4>.n75 tb<4>.n74 0.0419706
R10941 tb<4>.n82 tb<4>.n81 0.0419706
R10942 tb<4>.n89 tb<4>.n88 0.0419706
R10943 tb<4>.n8 tb<4>.n7 0.0419706
R10944 tb<4>.n15 tb<4>.n14 0.0419706
R10945 tb<4>.n22 tb<4>.n21 0.0419706
R10946 tb<4>.n29 tb<4>.n28 0.0419706
R10947 tb<4>.n36 tb<4>.n35 0.0419706
R10948 tb<4>.n43 tb<4>.n42 0.0419706
R10949 tb<4>.n97 tb<4>.n96 0.0170118
R10950 tb<4>.n60 tb<4>.n59 0.0143235
R10951 tb<4>.n67 tb<4>.n66 0.0143235
R10952 tb<4>.n74 tb<4>.n73 0.0143235
R10953 tb<4>.n81 tb<4>.n80 0.0143235
R10954 tb<4>.n88 tb<4>.n87 0.0143235
R10955 tb<4> tb<4>.n95 0.0143235
R10956 tb<4>.n2 tb<4>.n1 0.0143235
R10957 tb<4>.n9 tb<4>.n8 0.0143235
R10958 tb<4>.n16 tb<4>.n15 0.0143235
R10959 tb<4>.n23 tb<4>.n22 0.0143235
R10960 tb<4>.n30 tb<4>.n29 0.0143235
R10961 tb<4>.n37 tb<4>.n36 0.0143235
R10962 tb<4>.n44 tb<4>.n43 0.0143235
R10963 tb<4>.n47 tb<4>.n46 0.0138432
R10964 tb<4>.n99 tb<4>.n98 0.0100893
R10965 tb<4>.n48 tb<4>.n47 0.006246
R10966 tb<4>.n95 tb<4>.n94 0.00533824
R10967 tb<4>.n46 tb<4>.n45 0.00533824
R10968 tb<4>.n96 tb<4> 0.00395588
R10969 tb<4>.n50 tb<4>.n49 0.00349062
R10970 tb<4>.n98 tb<4>.n51 0.00349062
R10971 tb<4> tb<4>.n99 0.00331784
R10972 tb<5>.n59 tb<5> 0.746233
R10973 tb<5>.n197 tb<5>.n196 0.3805
R10974 tb<5>.n293 tb<5>.n292 0.3805
R10975 tb<5>.n4 tb<5>.n3 0.3424
R10976 tb<5>.n298 tb<5>.n297 0.3424
R10977 tb<5>.n5 tb<5> 0.255933
R10978 tb<5>.n6 tb<5>.n5 0.207891
R10979 tb<5>.n201 tb<5>.n200 0.204769
R10980 tb<5>.n209 tb<5>.n208 0.142882
R10981 tb<5>.n215 tb<5>.n214 0.142882
R10982 tb<5>.n221 tb<5>.n220 0.142882
R10983 tb<5>.n227 tb<5>.n226 0.142882
R10984 tb<5>.n233 tb<5>.n232 0.142882
R10985 tb<5>.n239 tb<5>.n238 0.142882
R10986 tb<5>.n245 tb<5>.n244 0.142882
R10987 tb<5>.n251 tb<5>.n250 0.142882
R10988 tb<5>.n257 tb<5>.n256 0.142882
R10989 tb<5>.n263 tb<5>.n262 0.142882
R10990 tb<5>.n269 tb<5>.n268 0.142882
R10991 tb<5>.n275 tb<5>.n274 0.142882
R10992 tb<5>.n281 tb<5>.n280 0.142882
R10993 tb<5>.n287 tb<5>.n286 0.142882
R10994 tb<5>.n113 tb<5>.n112 0.142882
R10995 tb<5>.n119 tb<5>.n118 0.142882
R10996 tb<5>.n125 tb<5>.n124 0.142882
R10997 tb<5>.n131 tb<5>.n130 0.142882
R10998 tb<5>.n137 tb<5>.n136 0.142882
R10999 tb<5>.n143 tb<5>.n142 0.142882
R11000 tb<5>.n149 tb<5>.n148 0.142882
R11001 tb<5>.n155 tb<5>.n154 0.142882
R11002 tb<5>.n161 tb<5>.n160 0.142882
R11003 tb<5>.n167 tb<5>.n166 0.142882
R11004 tb<5>.n173 tb<5>.n172 0.142882
R11005 tb<5>.n179 tb<5>.n178 0.142882
R11006 tb<5>.n185 tb<5>.n184 0.142882
R11007 tb<5>.n191 tb<5>.n190 0.142882
R11008 tb<5>.n11 tb<5>.n10 0.142882
R11009 tb<5>.n18 tb<5>.n17 0.142882
R11010 tb<5>.n25 tb<5>.n24 0.142882
R11011 tb<5>.n32 tb<5>.n31 0.142882
R11012 tb<5>.n39 tb<5>.n38 0.142882
R11013 tb<5>.n46 tb<5>.n45 0.142882
R11014 tb<5>.n53 tb<5>.n52 0.142882
R11015 tb<5>.n61 tb<5>.n60 0.142882
R11016 tb<5>.n68 tb<5>.n67 0.142882
R11017 tb<5>.n75 tb<5>.n74 0.142882
R11018 tb<5>.n82 tb<5>.n81 0.142882
R11019 tb<5>.n89 tb<5>.n88 0.142882
R11020 tb<5>.n96 tb<5>.n95 0.142882
R11021 tb<5>.n103 tb<5>.n102 0.142882
R11022 tb<5>.n199 tb<5>.n2 0.130613
R11023 tb<5>.n199 tb<5>.n198 0.125385
R11024 tb<5>.n300 tb<5>.n299 0.119792
R11025 tb<5>.n105 tb<5> 0.0976333
R11026 tb<5>.n98 tb<5> 0.0976333
R11027 tb<5>.n91 tb<5> 0.0976333
R11028 tb<5>.n84 tb<5> 0.0976333
R11029 tb<5>.n77 tb<5> 0.0976333
R11030 tb<5>.n70 tb<5> 0.0976333
R11031 tb<5>.n63 tb<5> 0.0976333
R11032 tb<5>.n55 tb<5> 0.0976333
R11033 tb<5>.n48 tb<5> 0.0976333
R11034 tb<5>.n41 tb<5> 0.0976333
R11035 tb<5>.n34 tb<5> 0.0976333
R11036 tb<5>.n27 tb<5> 0.0976333
R11037 tb<5>.n20 tb<5> 0.0976333
R11038 tb<5>.n13 tb<5> 0.0976333
R11039 tb<5>.n6 tb<5> 0.0976333
R11040 tb<5>.n206 tb<5> 0.0725667
R11041 tb<5>.n208 tb<5>.n207 0.0557941
R11042 tb<5>.n210 tb<5>.n209 0.0557941
R11043 tb<5>.n211 tb<5>.n210 0.0557941
R11044 tb<5>.n212 tb<5>.n211 0.0557941
R11045 tb<5>.n213 tb<5>.n212 0.0557941
R11046 tb<5>.n214 tb<5>.n213 0.0557941
R11047 tb<5>.n216 tb<5>.n215 0.0557941
R11048 tb<5>.n217 tb<5>.n216 0.0557941
R11049 tb<5>.n218 tb<5>.n217 0.0557941
R11050 tb<5>.n219 tb<5>.n218 0.0557941
R11051 tb<5>.n220 tb<5>.n219 0.0557941
R11052 tb<5>.n222 tb<5>.n221 0.0557941
R11053 tb<5>.n223 tb<5>.n222 0.0557941
R11054 tb<5>.n224 tb<5>.n223 0.0557941
R11055 tb<5>.n225 tb<5>.n224 0.0557941
R11056 tb<5>.n226 tb<5>.n225 0.0557941
R11057 tb<5>.n228 tb<5>.n227 0.0557941
R11058 tb<5>.n229 tb<5>.n228 0.0557941
R11059 tb<5>.n230 tb<5>.n229 0.0557941
R11060 tb<5>.n231 tb<5>.n230 0.0557941
R11061 tb<5>.n232 tb<5>.n231 0.0557941
R11062 tb<5>.n234 tb<5>.n233 0.0557941
R11063 tb<5>.n235 tb<5>.n234 0.0557941
R11064 tb<5>.n236 tb<5>.n235 0.0557941
R11065 tb<5>.n237 tb<5>.n236 0.0557941
R11066 tb<5>.n238 tb<5>.n237 0.0557941
R11067 tb<5>.n240 tb<5>.n239 0.0557941
R11068 tb<5>.n241 tb<5>.n240 0.0557941
R11069 tb<5>.n242 tb<5>.n241 0.0557941
R11070 tb<5>.n243 tb<5>.n242 0.0557941
R11071 tb<5>.n244 tb<5>.n243 0.0557941
R11072 tb<5>.n246 tb<5>.n245 0.0557941
R11073 tb<5>.n247 tb<5>.n246 0.0557941
R11074 tb<5>.n248 tb<5>.n247 0.0557941
R11075 tb<5>.n249 tb<5>.n248 0.0557941
R11076 tb<5>.n250 tb<5>.n249 0.0557941
R11077 tb<5>.n252 tb<5>.n251 0.0557941
R11078 tb<5>.n253 tb<5>.n252 0.0557941
R11079 tb<5>.n254 tb<5>.n253 0.0557941
R11080 tb<5>.n255 tb<5>.n254 0.0557941
R11081 tb<5>.n256 tb<5>.n255 0.0557941
R11082 tb<5>.n258 tb<5>.n257 0.0557941
R11083 tb<5>.n259 tb<5>.n258 0.0557941
R11084 tb<5>.n260 tb<5>.n259 0.0557941
R11085 tb<5>.n261 tb<5>.n260 0.0557941
R11086 tb<5>.n262 tb<5>.n261 0.0557941
R11087 tb<5>.n264 tb<5>.n263 0.0557941
R11088 tb<5>.n265 tb<5>.n264 0.0557941
R11089 tb<5>.n266 tb<5>.n265 0.0557941
R11090 tb<5>.n267 tb<5>.n266 0.0557941
R11091 tb<5>.n268 tb<5>.n267 0.0557941
R11092 tb<5>.n270 tb<5>.n269 0.0557941
R11093 tb<5>.n271 tb<5>.n270 0.0557941
R11094 tb<5>.n272 tb<5>.n271 0.0557941
R11095 tb<5>.n273 tb<5>.n272 0.0557941
R11096 tb<5>.n274 tb<5>.n273 0.0557941
R11097 tb<5>.n276 tb<5>.n275 0.0557941
R11098 tb<5>.n277 tb<5>.n276 0.0557941
R11099 tb<5>.n278 tb<5>.n277 0.0557941
R11100 tb<5>.n279 tb<5>.n278 0.0557941
R11101 tb<5>.n280 tb<5>.n279 0.0557941
R11102 tb<5>.n282 tb<5>.n281 0.0557941
R11103 tb<5>.n283 tb<5>.n282 0.0557941
R11104 tb<5>.n284 tb<5>.n283 0.0557941
R11105 tb<5>.n285 tb<5>.n284 0.0557941
R11106 tb<5>.n286 tb<5>.n285 0.0557941
R11107 tb<5>.n288 tb<5>.n287 0.0557941
R11108 tb<5>.n289 tb<5>.n288 0.0557941
R11109 tb<5>.n202 tb<5> 0.0557941
R11110 tb<5>.n203 tb<5>.n202 0.0557941
R11111 tb<5>.n110 tb<5>.n109 0.0557941
R11112 tb<5>.n111 tb<5>.n110 0.0557941
R11113 tb<5>.n112 tb<5>.n111 0.0557941
R11114 tb<5>.n114 tb<5>.n113 0.0557941
R11115 tb<5>.n115 tb<5>.n114 0.0557941
R11116 tb<5>.n116 tb<5>.n115 0.0557941
R11117 tb<5>.n117 tb<5>.n116 0.0557941
R11118 tb<5>.n118 tb<5>.n117 0.0557941
R11119 tb<5>.n120 tb<5>.n119 0.0557941
R11120 tb<5>.n121 tb<5>.n120 0.0557941
R11121 tb<5>.n122 tb<5>.n121 0.0557941
R11122 tb<5>.n123 tb<5>.n122 0.0557941
R11123 tb<5>.n124 tb<5>.n123 0.0557941
R11124 tb<5>.n126 tb<5>.n125 0.0557941
R11125 tb<5>.n127 tb<5>.n126 0.0557941
R11126 tb<5>.n128 tb<5>.n127 0.0557941
R11127 tb<5>.n129 tb<5>.n128 0.0557941
R11128 tb<5>.n130 tb<5>.n129 0.0557941
R11129 tb<5>.n132 tb<5>.n131 0.0557941
R11130 tb<5>.n133 tb<5>.n132 0.0557941
R11131 tb<5>.n134 tb<5>.n133 0.0557941
R11132 tb<5>.n135 tb<5>.n134 0.0557941
R11133 tb<5>.n136 tb<5>.n135 0.0557941
R11134 tb<5>.n138 tb<5>.n137 0.0557941
R11135 tb<5>.n139 tb<5>.n138 0.0557941
R11136 tb<5>.n140 tb<5>.n139 0.0557941
R11137 tb<5>.n141 tb<5>.n140 0.0557941
R11138 tb<5>.n142 tb<5>.n141 0.0557941
R11139 tb<5>.n144 tb<5>.n143 0.0557941
R11140 tb<5>.n145 tb<5>.n144 0.0557941
R11141 tb<5>.n146 tb<5>.n145 0.0557941
R11142 tb<5>.n147 tb<5>.n146 0.0557941
R11143 tb<5>.n148 tb<5>.n147 0.0557941
R11144 tb<5>.n150 tb<5>.n149 0.0557941
R11145 tb<5>.n151 tb<5>.n150 0.0557941
R11146 tb<5>.n152 tb<5>.n151 0.0557941
R11147 tb<5>.n153 tb<5>.n152 0.0557941
R11148 tb<5>.n154 tb<5>.n153 0.0557941
R11149 tb<5>.n156 tb<5>.n155 0.0557941
R11150 tb<5>.n157 tb<5>.n156 0.0557941
R11151 tb<5>.n158 tb<5>.n157 0.0557941
R11152 tb<5>.n159 tb<5>.n158 0.0557941
R11153 tb<5>.n160 tb<5>.n159 0.0557941
R11154 tb<5>.n162 tb<5>.n161 0.0557941
R11155 tb<5>.n163 tb<5>.n162 0.0557941
R11156 tb<5>.n164 tb<5>.n163 0.0557941
R11157 tb<5>.n165 tb<5>.n164 0.0557941
R11158 tb<5>.n166 tb<5>.n165 0.0557941
R11159 tb<5>.n168 tb<5>.n167 0.0557941
R11160 tb<5>.n169 tb<5>.n168 0.0557941
R11161 tb<5>.n170 tb<5>.n169 0.0557941
R11162 tb<5>.n171 tb<5>.n170 0.0557941
R11163 tb<5>.n172 tb<5>.n171 0.0557941
R11164 tb<5>.n174 tb<5>.n173 0.0557941
R11165 tb<5>.n175 tb<5>.n174 0.0557941
R11166 tb<5>.n176 tb<5>.n175 0.0557941
R11167 tb<5>.n177 tb<5>.n176 0.0557941
R11168 tb<5>.n178 tb<5>.n177 0.0557941
R11169 tb<5>.n180 tb<5>.n179 0.0557941
R11170 tb<5>.n181 tb<5>.n180 0.0557941
R11171 tb<5>.n182 tb<5>.n181 0.0557941
R11172 tb<5>.n183 tb<5>.n182 0.0557941
R11173 tb<5>.n184 tb<5>.n183 0.0557941
R11174 tb<5>.n186 tb<5>.n185 0.0557941
R11175 tb<5>.n187 tb<5>.n186 0.0557941
R11176 tb<5>.n188 tb<5>.n187 0.0557941
R11177 tb<5>.n189 tb<5>.n188 0.0557941
R11178 tb<5>.n190 tb<5>.n189 0.0557941
R11179 tb<5>.n192 tb<5>.n191 0.0557941
R11180 tb<5>.n193 tb<5>.n192 0.0557941
R11181 tb<5>.n8 tb<5>.n7 0.0557941
R11182 tb<5>.n9 tb<5>.n8 0.0557941
R11183 tb<5>.n10 tb<5>.n9 0.0557941
R11184 tb<5>.n12 tb<5>.n11 0.0557941
R11185 tb<5>.n15 tb<5>.n14 0.0557941
R11186 tb<5>.n16 tb<5>.n15 0.0557941
R11187 tb<5>.n17 tb<5>.n16 0.0557941
R11188 tb<5>.n19 tb<5>.n18 0.0557941
R11189 tb<5>.n22 tb<5>.n21 0.0557941
R11190 tb<5>.n23 tb<5>.n22 0.0557941
R11191 tb<5>.n24 tb<5>.n23 0.0557941
R11192 tb<5>.n26 tb<5>.n25 0.0557941
R11193 tb<5>.n29 tb<5>.n28 0.0557941
R11194 tb<5>.n30 tb<5>.n29 0.0557941
R11195 tb<5>.n31 tb<5>.n30 0.0557941
R11196 tb<5>.n33 tb<5>.n32 0.0557941
R11197 tb<5>.n36 tb<5>.n35 0.0557941
R11198 tb<5>.n37 tb<5>.n36 0.0557941
R11199 tb<5>.n38 tb<5>.n37 0.0557941
R11200 tb<5>.n40 tb<5>.n39 0.0557941
R11201 tb<5>.n43 tb<5>.n42 0.0557941
R11202 tb<5>.n44 tb<5>.n43 0.0557941
R11203 tb<5>.n45 tb<5>.n44 0.0557941
R11204 tb<5>.n47 tb<5>.n46 0.0557941
R11205 tb<5>.n50 tb<5>.n49 0.0557941
R11206 tb<5>.n51 tb<5>.n50 0.0557941
R11207 tb<5>.n52 tb<5>.n51 0.0557941
R11208 tb<5>.n54 tb<5>.n53 0.0557941
R11209 tb<5>.n57 tb<5>.n56 0.0557941
R11210 tb<5>.n58 tb<5>.n57 0.0557941
R11211 tb<5>.n62 tb<5>.n61 0.0557941
R11212 tb<5>.n65 tb<5>.n64 0.0557941
R11213 tb<5>.n66 tb<5>.n65 0.0557941
R11214 tb<5>.n67 tb<5>.n66 0.0557941
R11215 tb<5>.n69 tb<5>.n68 0.0557941
R11216 tb<5>.n72 tb<5>.n71 0.0557941
R11217 tb<5>.n73 tb<5>.n72 0.0557941
R11218 tb<5>.n74 tb<5>.n73 0.0557941
R11219 tb<5>.n76 tb<5>.n75 0.0557941
R11220 tb<5>.n79 tb<5>.n78 0.0557941
R11221 tb<5>.n80 tb<5>.n79 0.0557941
R11222 tb<5>.n81 tb<5>.n80 0.0557941
R11223 tb<5>.n83 tb<5>.n82 0.0557941
R11224 tb<5>.n86 tb<5>.n85 0.0557941
R11225 tb<5>.n87 tb<5>.n86 0.0557941
R11226 tb<5>.n88 tb<5>.n87 0.0557941
R11227 tb<5>.n90 tb<5>.n89 0.0557941
R11228 tb<5>.n93 tb<5>.n92 0.0557941
R11229 tb<5>.n94 tb<5>.n93 0.0557941
R11230 tb<5>.n95 tb<5>.n94 0.0557941
R11231 tb<5>.n97 tb<5>.n96 0.0557941
R11232 tb<5>.n100 tb<5>.n99 0.0557941
R11233 tb<5>.n101 tb<5>.n100 0.0557941
R11234 tb<5>.n102 tb<5>.n101 0.0557941
R11235 tb<5>.n104 tb<5>.n103 0.0557941
R11236 tb<5>.n290 tb<5>.n289 0.0509559
R11237 tb<5>.n204 tb<5>.n203 0.0509559
R11238 tb<5>.n194 tb<5>.n193 0.0509559
R11239 tb<5>.n107 tb<5>.n106 0.0509559
R11240 tb<5>.n13 tb<5>.n12 0.0419706
R11241 tb<5>.n20 tb<5>.n19 0.0419706
R11242 tb<5>.n27 tb<5>.n26 0.0419706
R11243 tb<5>.n34 tb<5>.n33 0.0419706
R11244 tb<5>.n41 tb<5>.n40 0.0419706
R11245 tb<5>.n48 tb<5>.n47 0.0419706
R11246 tb<5>.n55 tb<5>.n54 0.0419706
R11247 tb<5>.n59 tb<5>.n58 0.0419706
R11248 tb<5>.n63 tb<5>.n62 0.0419706
R11249 tb<5>.n70 tb<5>.n69 0.0419706
R11250 tb<5>.n77 tb<5>.n76 0.0419706
R11251 tb<5>.n84 tb<5>.n83 0.0419706
R11252 tb<5>.n91 tb<5>.n90 0.0419706
R11253 tb<5>.n98 tb<5>.n97 0.0419706
R11254 tb<5>.n105 tb<5>.n104 0.0419706
R11255 tb<5>.n298 tb<5>.n296 0.0281471
R11256 tb<5>.n299 tb<5>.n298 0.0220232
R11257 tb<5>.n292 tb<5>.n291 0.0177794
R11258 tb<5>.n196 tb<5>.n195 0.0177794
R11259 tb<5>.n295 tb<5>.n294 0.0170882
R11260 tb<5>.n299 tb<5>.n293 0.0170118
R11261 tb<5>.n206 tb<5>.n205 0.0143235
R11262 tb<5>.n7 tb<5>.n6 0.0143235
R11263 tb<5>.n14 tb<5>.n13 0.0143235
R11264 tb<5>.n21 tb<5>.n20 0.0143235
R11265 tb<5>.n28 tb<5>.n27 0.0143235
R11266 tb<5>.n35 tb<5>.n34 0.0143235
R11267 tb<5>.n42 tb<5>.n41 0.0143235
R11268 tb<5>.n49 tb<5>.n48 0.0143235
R11269 tb<5>.n56 tb<5>.n55 0.0143235
R11270 tb<5>.n60 tb<5>.n59 0.0143235
R11271 tb<5>.n64 tb<5>.n63 0.0143235
R11272 tb<5>.n71 tb<5>.n70 0.0143235
R11273 tb<5>.n78 tb<5>.n77 0.0143235
R11274 tb<5>.n85 tb<5>.n84 0.0143235
R11275 tb<5>.n92 tb<5>.n91 0.0143235
R11276 tb<5>.n99 tb<5>.n98 0.0143235
R11277 tb<5>.n106 tb<5>.n105 0.0143235
R11278 tb<5>.n197 tb<5>.n108 0.0138432
R11279 tb<5>.n296 tb<5>.n295 0.0115588
R11280 tb<5>.n301 tb<5>.n300 0.0100893
R11281 tb<5>.n198 tb<5>.n4 0.00752478
R11282 tb<5>.n198 tb<5>.n197 0.006246
R11283 tb<5>.n291 tb<5>.n290 0.00533824
R11284 tb<5>.n205 tb<5>.n204 0.00533824
R11285 tb<5>.n195 tb<5>.n194 0.00533824
R11286 tb<5>.n108 tb<5>.n107 0.00533824
R11287 tb<5>.n1 tb<5>.n0 0.00527966
R11288 tb<5> tb<5>.n301 0.00503972
R11289 tb<5>.n293 tb<5>.n206 0.00395588
R11290 tb<5>.n200 tb<5>.n199 0.00349062
R11291 tb<5>.n300 tb<5>.n201 0.00349062
R11292 tb<5>.n2 tb<5>.n1 0.00208685
C0 hgu_cdac_8bit_array_2.drv<0> t<1> 0.0206f
C1 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT d<2> 0.249f
C2 hgu_cdac_8bit_array_3.drv<0> d<0> 0.0391f
C3 VDD hgu_cdac_8bit_array_3.drv<63:0> 1.5f
C4 t<2> tb<2> 0.394f
C5 hgu_cdac_8bit_array_3.drv<15:0> db<4> 0.0274f
C6 hgu_cdac_8bit_array_3.drv<0> t<2> 1.24e-19
C7 t<5> db<5> 0.387f
C8 VDD hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT 0.197f
C9 hgu_cdac_8bit_array_3.drv<1:0> t<1> 11.6f
C10 hgu_cdac_8bit_array_2.drv<31:0> hgu_cdac_8bit_array_2.drv<63:0> 2.28f
C11 VDD db<2> 0.251f
C12 hgu_cdac_8bit_array_3.drv<1:0> d<1> 0.0914f
C13 VREF db<3> 0.213f
C14 VDD t<3> 0.0631f
C15 VREF hgu_cdac_8bit_array_2.drv<0> 0.153f
C16 hgu_cdac_8bit_array_3.drv<0> t<1> 0.369f
C17 VREF t<5> 0.222f
C18 VREF hgu_cdac_8bit_array_2.drv<15:0> 2.12f
C19 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT d<3> 1.78e-19
C20 hgu_cdac_8bit_array_3.drv<0> d<1> 0.00519f
C21 t<1> t<2> 0.503f
C22 hgu_cdac_8bit_array_2.drv<63:0> tb<6> 0.325p
C23 d<0> d<1> 0.00414f
C24 hgu_cdac_8bit_array_3.drv<1:0> VREF 0.378f
C25 hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_8bit_array_2.drv<31:0> 0.967f
C26 t<3> d<3> 0.0494f
C27 hgu_cdac_8bit_array_2.drv<63:0> t<6> 4.72f
C28 VDD db<3> 0.509f
C29 VDD hgu_cdac_8bit_array_2.drv<0> 0.0314f
C30 VDD t<5> 0.226f
C31 hgu_cdac_8bit_array_3.drv<0> VREF 0.257f
C32 VDD hgu_cdac_8bit_array_2.drv<15:0> 0.14f
C33 hgu_cdac_8bit_array_3.drv<15:0> VREF 2.69f
C34 VREF d<0> 0.0246f
C35 hgu_cdac_8bit_array_3.drv<1:0> d<2> 2.5e-19
C36 VREF db<4> 0.43f
C37 VREF t<2> 0.0296f
C38 t<1> d<1> 0.0127f
C39 hgu_cdac_8bit_array_3.drv<63:0> tb<6> 0.00302f
C40 hgu_cdac_8bit_array_3.drv<0> d<2> 7.36e-19
C41 VDD hgu_cdac_8bit_array_3.drv<1:0> 0.0923f
C42 hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_8bit_array_3.drv<63:0> 2.29f
C43 tb<3> tb<4> 0.316f
C44 d<3> db<3> 0.03f
C45 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT hgu_cdac_8bit_array_2.drv<7:0> 1.08f
C46 hgu_cdac_8bit_array_3.drv<63:0> t<6> 0.328p
C47 t<2> d<2> 0.0256f
C48 VDD hgu_cdac_8bit_array_3.drv<0> 0.124f
C49 hgu_cdac_8bit_array_2.drv<31:0> tb<5> 0.163p
C50 VREF t<1> 0.0223f
C51 VDD hgu_cdac_8bit_array_3.drv<15:0> 0.471f
C52 VDD d<0> 0.0602f
C53 VDD db<4> 0.997f
C54 VREF d<1> 0.0484f
C55 VDD t<2> 0.0406f
C56 VREF db<5> 0.876f
C57 hgu_cdac_8bit_array_2.drv<31:0> t<5> 2.38f
C58 hgu_cdac_8bit_array_2.drv<15:0> hgu_cdac_8bit_array_2.drv<31:0> 2.28f
C59 t<3> t<4> 0.316f
C60 tb<5> tb<6> 0.186f
C61 tb<4> tb<5> 0.318f
C62 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT hgu_cdac_8bit_array_2.drv<7:0> 1.89e-21
C63 hgu_cdac_8bit_array_2.drv<7:0> tb<3> 42.3f
C64 hgu_cdac_8bit_array_3.drv<15:0> d<3> 1.49e-19
C65 d<1> d<2> 0.00443f
C66 hgu_cdac_8bit_array_2.drv<7:0> db<2> 1.93e-19
C67 hgu_cdac_8bit_array_3.drv<31:0> tb<5> 0.00263f
C68 VDD t<1> 0.0297f
C69 hgu_cdac_8bit_array_2.drv<7:0> t<3> 0.671f
C70 hgu_cdac_8bit_array_2.drv<15:0> tb<4> 82.5f
C71 VDD d<1> 0.128f
C72 VDD db<5> 2f
C73 hgu_cdac_8bit_array_3.drv<31:0> t<5> 0.165p
C74 hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_8bit_array_2.drv<15:0> 0.966f
C75 VREF d<2> 0.102f
C76 t<4> db<3> 0.00263f
C77 t<5> t<6> 0.186f
C78 t<4> t<5> 0.318f
C79 VREF db<6> 1.76f
C80 hgu_cdac_8bit_array_3.drv<63:0> d<6> 4.14f
C81 hgu_cdac_8bit_array_2.drv<15:0> t<4> 1.55f
C82 VDD VREF 49.1f
C83 hgu_cdac_8bit_array_3.drv<15:0> d<4> 1.03f
C84 db<0> db<1> 0.00352f
C85 hgu_cdac_8bit_array_2.drv<7:0> db<3> 0.448f
C86 t<5> d<5> 0.18f
C87 hgu_cdac_8bit_array_3.drv<15:0> tb<4> 0.00202f
C88 hgu_cdac_8bit_array_2.drv<7:0> hgu_cdac_8bit_array_2.drv<15:0> 2.27f
C89 hgu_cdac_8bit_array_2.drv<0> hgu_cdac_unit_0.CBOT 4.71e-19
C90 hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_8bit_array_3.drv<31:0> 2.29f
C91 VDD d<2> 0.251f
C92 VDD db<6> 4f
C93 hgu_cdac_8bit_array_3.drv<31:0> db<4> 0.0168f
C94 hgu_cdac_8bit_array_3.drv<15:0> t<4> 83.1f
C95 hgu_cdac_8bit_array_2.drv<0> hgu_cdac_unit_1.CBOT 0.387f
C96 VREF d<3> 0.212f
C97 t<4> db<4> 0.189f
C98 hgu_cdac_8bit_array_2.drv<31:0> db<5> 1.88f
C99 hgu_cdac_8bit_array_2.drv<7:0> tb<2> 0.016f
C100 hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_8bit_array_2.drv<7:0> 0.0699f
C101 d<2> d<3> 0.0026f
C102 hgu_cdac_8bit_array_3.drv<1:0> hgu_cdac_unit_1.CBOT 0.703f
C103 VREF hgu_cdac_8bit_array_2.drv<31:0> 4.1f
C104 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT db<1> 2.67e-19
C105 hgu_cdac_8bit_array_2.drv<7:0> t<2> 1.01e-20
C106 VDD d<3> 0.509f
C107 hgu_cdac_8bit_array_3.drv<0> hgu_cdac_unit_1.CBOT 0.00742f
C108 hgu_cdac_8bit_array_3.drv<63:0> hgu_cdac_8bit_array_2.drv<63:0> 7.25f
C109 hgu_cdac_8bit_array_3.drv<31:0> db<5> 0.0251f
C110 VREF d<4> 0.43f
C111 VDD hgu_cdac_8bit_array_2.drv<31:0> 0.252f
C112 hgu_cdac_8bit_array_3.drv<31:0> VREF 5.04f
C113 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT db<1> 0.00419f
C114 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT 2.13f
C115 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT tb<3> 0.03f
C116 VREF t<6> 0.525f
C117 VREF t<4> 0.114f
C118 db<1> db<2> 0.00284f
C119 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT db<2> 0.219f
C120 hgu_cdac_8bit_array_2.drv<0> db<0> 0.0294f
C121 t<1> hgu_cdac_unit_1.CBOT 0.381f
C122 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT t<3> 0.0103f
C123 VDD d<4> 0.997f
C124 hgu_cdac_8bit_array_2.drv<63:0> tb<5> 0.00164f
C125 t<6> db<6> 0.764f
C126 VREF d<5> 0.874f
C127 VREF hgu_cdac_8bit_array_2.drv<7:0> 1.07f
C128 hgu_cdac_8bit_array_3.drv<1:0> db<0> 2.72e-19
C129 VDD hgu_cdac_8bit_array_3.drv<31:0> 0.785f
C130 VDD t<6> 0.655f
C131 VDD t<4> 0.122f
C132 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT db<2> 0.0356f
C133 hgu_cdac_8bit_array_3.drv<0> db<0> 0.0154f
C134 d<3> d<4> 0.00198f
C135 d<0> db<0> 0.00636f
C136 hgu_cdac_8bit_array_2.drv<0> db<1> 7.56e-19
C137 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT t<3> 0.0216f
C138 t<3> tb<3> 0.636f
C139 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT db<3> 2.04e-19
C140 t<3> db<2> 0.00154f
C141 VDD d<5> 2f
C142 VDD hgu_cdac_8bit_array_2.drv<7:0> 0.0789f
C143 VREF d<6> 1.75f
C144 hgu_cdac_8bit_array_3.drv<1:0> db<1> 0.0135f
C145 hgu_cdac_8bit_array_3.drv<1:0> hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT 2.6e-20
C146 hgu_cdac_8bit_array_2.drv<31:0> tb<6> 0.0162f
C147 hgu_cdac_8bit_array_2.drv<31:0> tb<4> 0.00164f
C148 hgu_cdac_8bit_array_3.drv<63:0> t<5> 0.00511f
C149 t<1> db<0> 8.18e-19
C150 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT tb<2> 22.1f
C151 hgu_cdac_8bit_array_3.drv<31:0> hgu_cdac_8bit_array_2.drv<31:0> 3.77f
C152 hgu_cdac_8bit_array_3.drv<0> db<1> 4.18e-19
C153 hgu_cdac_8bit_array_3.drv<0> hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT 1.87e-20
C154 hgu_cdac_8bit_array_2.drv<15:0> tb<3> 0.00163f
C155 hgu_cdac_8bit_array_2.drv<7:0> d<3> 0.00405f
C156 hgu_cdac_8bit_array_2.drv<31:0> t<6> 0.0156f
C157 db<2> db<3> 0.0026f
C158 t<2> db<1> 0.00113f
C159 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT t<2> 0.571f
C160 t<3> db<3> 0.101f
C161 VDD d<6> 4f
C162 hgu_cdac_8bit_array_3.drv<1:0> hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT 1.11f
C163 t<4> d<4> 0.0905f
C164 VREF db<0> 0.0246f
C165 t<6> tb<6> 4.02f
C166 t<4> tb<4> 1.12f
C167 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT tb<2> 0.0014f
C168 tb<2> tb<3> 0.455f
C169 t<1> db<1> 0.0252f
C170 hgu_cdac_8bit_array_3.drv<0> hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT 0.00224f
C171 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT t<1> 6.12e-21
C172 t<5> tb<5> 2.08f
C173 hgu_cdac_8bit_array_3.drv<31:0> t<6> 0.00164f
C174 hgu_cdac_8bit_array_2.drv<15:0> tb<5> 0.323f
C175 hgu_cdac_8bit_array_3.drv<31:0> t<4> 0.0053f
C176 d<1> db<1> 0.00636f
C177 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT t<2> 22.2f
C178 hgu_cdac_8bit_array_2.drv<7:0> tb<4> 0.321f
C179 hgu_cdac_8bit_array_3.drv<15:0> t<3> 0.0213f
C180 t<2> db<2> 0.0514f
C181 hgu_cdac_8bit_array_2.drv<15:0> t<5> 0.0336f
C182 VREF hgu_cdac_8bit_array_2.drv<63:0> 8.33f
C183 VDD db<0> 0.0601f
C184 hgu_cdac_8bit_array_3.drv<31:0> d<5> 2.09f
C185 t<2> t<3> 0.455f
C186 hgu_cdac_8bit_array_2.drv<7:0> t<4> 0.00788f
C187 VREF db<1> 0.0484f
C188 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT t<1> 0.0226f
C189 VREF hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT 0.564f
C190 hgu_cdac_8bit_array_3.drv<1:0> hgu_cdac_8bit_array_2.drv<0> 0.13f
C191 hgu_cdac_8bit_array_3.drv<63:0> db<5> 0.0173f
C192 hgu_cdac_8bit_array_2.drv<63:0> db<6> 3.93f
C193 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT d<1> 0.00506f
C194 hgu_cdac_8bit_array_2.drv<0> tb<2> 2.41e-19
C195 hgu_cdac_8bit_array_3.drv<0> hgu_cdac_8bit_array_2.drv<0> 0.483f
C196 hgu_cdac_8bit_array_3.drv<15:0> db<3> 2.16e-19
C197 hgu_cdac_8bit_array_3.drv<15:0> t<5> 0.296f
C198 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT d<2> 0.0016f
C199 hgu_cdac_8bit_array_3.drv<15:0> hgu_cdac_8bit_array_2.drv<15:0> 2.96f
C200 t<5> db<4> 0.00575f
C201 hgu_cdac_8bit_array_3.drv<63:0> VREF 9.96f
C202 VDD hgu_cdac_8bit_array_2.drv<63:0> 0.509f
C203 hgu_cdac_8bit_array_2.drv<15:0> db<4> 0.976f
C204 VDD db<1> 0.128f
C205 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT VREF 0.826f
C206 VDD hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT 0.0484f
C207 hgu_cdac_8bit_array_3.drv<0> hgu_cdac_8bit_array_3.drv<1:0> 1.19f
C208 t<6> d<6> 0.36f
C209 hgu_cdac_8bit_array_3.drv<1:0> d<0> 2.76e-19
C210 VREF db<2> 0.102f
C211 hgu_cdac_8bit_array_3.drv<63:0> db<6> 0.0514f
C212 hgu_cdac_8bit_array_3.drv<1:0> t<2> 0.0233f
C213 VREF t<3> 0.0584f
C214 db<6> VSS 12.7f
C215 db<5> VSS 6.38f
C216 db<4> VSS 3.21f
C217 db<3> VSS 1.58f
C218 db<2> VSS 0.819f
C219 db<1> VSS 0.42f
C220 db<0> VSS 0.23f
C221 d<6> VSS 12.7f
C222 d<5> VSS 6.38f
C223 d<4> VSS 3.21f
C224 d<3> VSS 1.58f
C225 d<2> VSS 0.818f
C226 d<1> VSS 0.417f
C227 d<0> VSS 0.229f
C228 hgu_cdac_unit_0.CBOT VSS 0.995f $ **FLOATING
C229 tb<6> VSS -0.602p
C230 tb<5> VSS -1.21p
C231 tb<4> VSS 0.244p
C232 tb<3> VSS 27.2f
C233 tb<2> VSS 9.17f
C234 hgu_cdac_unit_1.CBOT VSS 0.812f $ **FLOATING
C235 t<6> VSS -0.689p
C236 t<5> VSS -1.79p
C237 t<4> VSS 0.337p
C238 t<3> VSS 50.4f
C239 t<2> VSS 18.8f
C240 t<1> VSS 10.1f
C241 hgu_cdac_8bit_array_2.drv<63:0> VSS 0.177p
C242 hgu_cdac_8bit_array_2.drv<31:0> VSS 0.186p
C243 hgu_cdac_8bit_array_2.drv<15:0> VSS 34.7f
C244 hgu_cdac_8bit_array_2.drv<7:0> VSS 14.4f
C245 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT VSS 12f
C246 hgu_cdac_8bit_array_2.drv<0> VSS 5.76f
C247 VREF VSS 34.9f
C248 hgu_cdac_8bit_array_3.drv<63:0> VSS 0.184p
C249 hgu_cdac_8bit_array_3.drv<31:0> VSS 86.7f
C250 hgu_cdac_8bit_array_3.drv<15:0> VSS 44.6f
C251 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT VSS 8.11f
C252 hgu_cdac_8bit_array_3.drv<1:0> VSS 5.58f
C253 hgu_cdac_8bit_array_3.drv<0> VSS 5.48f
C254 VDD VSS 53.3f
C255 tb<5>.n0 VSS -10.3f
C256 tb<5>.n1 VSS 34.4f
C257 tb<5>.n2 VSS -3.9f
C258 tb<5>.n3 VSS -11.6f
C259 tb<5>.n4 VSS -9.65f
C260 tb<5>.n5 VSS 40.7f
C261 tb<5>.n6 VSS -4.76f
C262 tb<5>.n7 VSS -2.66f
C263 tb<5>.n8 VSS -4.25f
C264 tb<5>.n9 VSS 7.82f
C265 tb<5>.n10 VSS 28.6f
C266 tb<5>.n11 VSS -7.6f
C267 tb<5>.n12 VSS -3.72f
C268 tb<5>.n13 VSS -5.03f
C269 tb<5>.n14 VSS -2.66f
C270 tb<5>.n15 VSS -4.25f
C271 tb<5>.n16 VSS 7.82f
C272 tb<5>.n17 VSS 28.6f
C273 tb<5>.n18 VSS -7.6f
C274 tb<5>.n19 VSS -3.72f
C275 tb<5>.n20 VSS -5.03f
C276 tb<5>.n21 VSS -2.66f
C277 tb<5>.n22 VSS -4.25f
C278 tb<5>.n23 VSS 7.82f
C279 tb<5>.n24 VSS 28.6f
C280 tb<5>.n25 VSS -7.6f
C281 tb<5>.n26 VSS -3.72f
C282 tb<5>.n27 VSS -5.03f
C283 tb<5>.n28 VSS -2.66f
C284 tb<5>.n29 VSS -4.25f
C285 tb<5>.n30 VSS 7.82f
C286 tb<5>.n31 VSS 28.6f
C287 tb<5>.n32 VSS -7.6f
C288 tb<5>.n33 VSS -3.72f
C289 tb<5>.n34 VSS -5.03f
C290 tb<5>.n35 VSS -2.66f
C291 tb<5>.n36 VSS -4.25f
C292 tb<5>.n37 VSS 7.82f
C293 tb<5>.n38 VSS 28.6f
C294 tb<5>.n39 VSS -7.6f
C295 tb<5>.n40 VSS -3.72f
C296 tb<5>.n41 VSS -5.03f
C297 tb<5>.n42 VSS -2.66f
C298 tb<5>.n43 VSS -4.25f
C299 tb<5>.n44 VSS 7.82f
C300 tb<5>.n45 VSS 28.6f
C301 tb<5>.n46 VSS -7.6f
C302 tb<5>.n47 VSS -3.72f
C303 tb<5>.n48 VSS -5.03f
C304 tb<5>.n49 VSS -2.66f
C305 tb<5>.n50 VSS -4.25f
C306 tb<5>.n51 VSS 7.82f
C307 tb<5>.n52 VSS 28.6f
C308 tb<5>.n53 VSS -7.6f
C309 tb<5>.n54 VSS -3.72f
C310 tb<5>.n55 VSS -5.03f
C311 tb<5>.n56 VSS -2.66f
C312 tb<5>.n57 VSS -4.25f
C313 tb<5>.n58 VSS -3.72f
C314 tb<5>.n59 VSS -24.4f
C315 tb<5>.n60 VSS -6f
C316 tb<5>.n61 VSS -7.6f
C317 tb<5>.n62 VSS -3.72f
C318 tb<5>.n63 VSS -5.03f
C319 tb<5>.n64 VSS -2.66f
C320 tb<5>.n65 VSS -4.25f
C321 tb<5>.n66 VSS 7.82f
C322 tb<5>.n67 VSS 28.6f
C323 tb<5>.n68 VSS -7.6f
C324 tb<5>.n69 VSS -3.72f
C325 tb<5>.n70 VSS -5.03f
C326 tb<5>.n71 VSS -2.66f
C327 tb<5>.n72 VSS -4.25f
C328 tb<5>.n73 VSS 7.82f
C329 tb<5>.n74 VSS 28.6f
C330 tb<5>.n75 VSS -7.6f
C331 tb<5>.n76 VSS -3.72f
C332 tb<5>.n77 VSS -5.03f
C333 tb<5>.n78 VSS -2.66f
C334 tb<5>.n79 VSS -4.25f
C335 tb<5>.n80 VSS 7.82f
C336 tb<5>.n81 VSS 28.6f
C337 tb<5>.n82 VSS -7.6f
C338 tb<5>.n83 VSS -3.72f
C339 tb<5>.n84 VSS -5.03f
C340 tb<5>.n85 VSS -2.66f
C341 tb<5>.n86 VSS -4.25f
C342 tb<5>.n87 VSS 7.82f
C343 tb<5>.n88 VSS 28.6f
C344 tb<5>.n89 VSS -7.6f
C345 tb<5>.n90 VSS -3.72f
C346 tb<5>.n91 VSS -5.03f
C347 tb<5>.n92 VSS -2.66f
C348 tb<5>.n93 VSS -4.25f
C349 tb<5>.n94 VSS 7.82f
C350 tb<5>.n95 VSS 28.6f
C351 tb<5>.n96 VSS -7.6f
C352 tb<5>.n97 VSS -3.72f
C353 tb<5>.n98 VSS -5.03f
C354 tb<5>.n99 VSS -2.66f
C355 tb<5>.n100 VSS -4.25f
C356 tb<5>.n101 VSS 7.82f
C357 tb<5>.n102 VSS 28.6f
C358 tb<5>.n103 VSS -7.6f
C359 tb<5>.n104 VSS -3.72f
C360 tb<5>.n105 VSS -5.03f
C361 tb<5>.n106 VSS -2.47f
C362 tb<5>.n107 VSS -2.13f
C363 tb<5>.n108 VSS -0.78f
C364 tb<5>.n109 VSS 44.8f
C365 tb<5>.n110 VSS 32f
C366 tb<5>.n111 VSS 7.82f
C367 tb<5>.n112 VSS -7.6f
C368 tb<5>.n113 VSS 28.6f
C369 tb<5>.n114 VSS 7.82f
C370 tb<5>.n115 VSS -4.25f
C371 tb<5>.n116 VSS 32f
C372 tb<5>.n117 VSS 7.82f
C373 tb<5>.n118 VSS -7.6f
C374 tb<5>.n119 VSS 28.6f
C375 tb<5>.n120 VSS 7.82f
C376 tb<5>.n121 VSS -4.25f
C377 tb<5>.n122 VSS 32f
C378 tb<5>.n123 VSS 7.82f
C379 tb<5>.n124 VSS -7.6f
C380 tb<5>.n125 VSS 28.6f
C381 tb<5>.n126 VSS 7.82f
C382 tb<5>.n127 VSS -4.25f
C383 tb<5>.n128 VSS 32f
C384 tb<5>.n129 VSS 7.82f
C385 tb<5>.n130 VSS -7.6f
C386 tb<5>.n131 VSS 28.6f
C387 tb<5>.n132 VSS 7.82f
C388 tb<5>.n133 VSS -4.25f
C389 tb<5>.n134 VSS 32f
C390 tb<5>.n135 VSS 7.82f
C391 tb<5>.n136 VSS -7.6f
C392 tb<5>.n137 VSS 28.6f
C393 tb<5>.n138 VSS 7.82f
C394 tb<5>.n139 VSS -4.25f
C395 tb<5>.n140 VSS 32f
C396 tb<5>.n141 VSS 7.82f
C397 tb<5>.n142 VSS -7.6f
C398 tb<5>.n143 VSS 28.6f
C399 tb<5>.n144 VSS 7.82f
C400 tb<5>.n145 VSS -4.25f
C401 tb<5>.n146 VSS 32f
C402 tb<5>.n147 VSS 7.82f
C403 tb<5>.n148 VSS -7.6f
C404 tb<5>.n149 VSS 28.6f
C405 tb<5>.n150 VSS 7.82f
C406 tb<5>.n151 VSS -4.25f
C407 tb<5>.n152 VSS 32f
C408 tb<5>.n153 VSS 7.82f
C409 tb<5>.n154 VSS -7.6f
C410 tb<5>.n155 VSS 28.6f
C411 tb<5>.n156 VSS 7.82f
C412 tb<5>.n157 VSS -4.25f
C413 tb<5>.n158 VSS 32f
C414 tb<5>.n159 VSS 7.82f
C415 tb<5>.n160 VSS -7.6f
C416 tb<5>.n161 VSS 28.6f
C417 tb<5>.n162 VSS 7.82f
C418 tb<5>.n163 VSS -4.25f
C419 tb<5>.n164 VSS 32f
C420 tb<5>.n165 VSS 7.82f
C421 tb<5>.n166 VSS -7.6f
C422 tb<5>.n167 VSS 28.6f
C423 tb<5>.n168 VSS 7.82f
C424 tb<5>.n169 VSS -4.25f
C425 tb<5>.n170 VSS 32f
C426 tb<5>.n171 VSS 7.82f
C427 tb<5>.n172 VSS -7.6f
C428 tb<5>.n173 VSS 28.6f
C429 tb<5>.n174 VSS 7.82f
C430 tb<5>.n175 VSS -4.25f
C431 tb<5>.n176 VSS 32f
C432 tb<5>.n177 VSS 7.82f
C433 tb<5>.n178 VSS -7.6f
C434 tb<5>.n179 VSS 28.6f
C435 tb<5>.n180 VSS 7.82f
C436 tb<5>.n181 VSS -4.25f
C437 tb<5>.n182 VSS 32f
C438 tb<5>.n183 VSS 7.82f
C439 tb<5>.n184 VSS -7.6f
C440 tb<5>.n185 VSS 28.6f
C441 tb<5>.n186 VSS 7.82f
C442 tb<5>.n187 VSS -4.25f
C443 tb<5>.n188 VSS 32f
C444 tb<5>.n189 VSS 7.82f
C445 tb<5>.n190 VSS -7.6f
C446 tb<5>.n191 VSS 28.6f
C447 tb<5>.n192 VSS 7.82f
C448 tb<5>.n193 VSS -4.06f
C449 tb<5>.n194 VSS -2.13f
C450 tb<5>.n195 VSS 8.81f
C451 tb<5>.n196 VSS 36.5f
C452 tb<5>.n197 VSS -5.82f
C453 tb<5>.n198 VSS -1.4f
C454 tb<5>.n199 VSS -62.3f
C455 tb<5>.n200 VSS -0.286p
C456 tb<5>.n201 VSS -0.286p
C457 tb<5>.n202 VSS 7.82f
C458 tb<5>.n203 VSS -4.06f
C459 tb<5>.n204 VSS -2.13f
C460 tb<5>.n205 VSS -0.717f
C461 tb<5>.n206 VSS -2.82f
C462 tb<5>.n207 VSS 47.9f
C463 tb<5>.n208 VSS 28.6f
C464 tb<5>.n209 VSS -7.6f
C465 tb<5>.n210 VSS 7.82f
C466 tb<5>.n211 VSS 32f
C467 tb<5>.n212 VSS -4.25f
C468 tb<5>.n213 VSS 7.82f
C469 tb<5>.n214 VSS 28.6f
C470 tb<5>.n215 VSS -7.6f
C471 tb<5>.n216 VSS 7.82f
C472 tb<5>.n217 VSS 32f
C473 tb<5>.n218 VSS -4.25f
C474 tb<5>.n219 VSS 7.82f
C475 tb<5>.n220 VSS 28.6f
C476 tb<5>.n221 VSS -7.6f
C477 tb<5>.n222 VSS 7.82f
C478 tb<5>.n223 VSS 32f
C479 tb<5>.n224 VSS -4.25f
C480 tb<5>.n225 VSS 7.82f
C481 tb<5>.n226 VSS 28.6f
C482 tb<5>.n227 VSS -7.6f
C483 tb<5>.n228 VSS 7.82f
C484 tb<5>.n229 VSS 32f
C485 tb<5>.n230 VSS -4.25f
C486 tb<5>.n231 VSS 7.82f
C487 tb<5>.n232 VSS 28.6f
C488 tb<5>.n233 VSS -7.6f
C489 tb<5>.n234 VSS 7.82f
C490 tb<5>.n235 VSS 32f
C491 tb<5>.n236 VSS -4.25f
C492 tb<5>.n237 VSS 7.82f
C493 tb<5>.n238 VSS 28.6f
C494 tb<5>.n239 VSS -7.6f
C495 tb<5>.n240 VSS 7.82f
C496 tb<5>.n241 VSS 32f
C497 tb<5>.n242 VSS -4.25f
C498 tb<5>.n243 VSS 7.82f
C499 tb<5>.n244 VSS 28.6f
C500 tb<5>.n245 VSS -7.6f
C501 tb<5>.n246 VSS 7.82f
C502 tb<5>.n247 VSS 32f
C503 tb<5>.n248 VSS -4.25f
C504 tb<5>.n249 VSS 7.82f
C505 tb<5>.n250 VSS 28.6f
C506 tb<5>.n251 VSS -7.6f
C507 tb<5>.n252 VSS 7.82f
C508 tb<5>.n253 VSS 32f
C509 tb<5>.n254 VSS -4.25f
C510 tb<5>.n255 VSS 7.82f
C511 tb<5>.n256 VSS 28.6f
C512 tb<5>.n257 VSS -7.6f
C513 tb<5>.n258 VSS 7.82f
C514 tb<5>.n259 VSS 32f
C515 tb<5>.n260 VSS -4.25f
C516 tb<5>.n261 VSS 7.82f
C517 tb<5>.n262 VSS 28.6f
C518 tb<5>.n263 VSS -7.6f
C519 tb<5>.n264 VSS 7.82f
C520 tb<5>.n265 VSS 32f
C521 tb<5>.n266 VSS -4.25f
C522 tb<5>.n267 VSS 7.82f
C523 tb<5>.n268 VSS 28.6f
C524 tb<5>.n269 VSS -7.6f
C525 tb<5>.n270 VSS 7.82f
C526 tb<5>.n271 VSS 32f
C527 tb<5>.n272 VSS -4.25f
C528 tb<5>.n273 VSS 7.82f
C529 tb<5>.n274 VSS 28.6f
C530 tb<5>.n275 VSS -7.6f
C531 tb<5>.n276 VSS 7.82f
C532 tb<5>.n277 VSS 32f
C533 tb<5>.n278 VSS -4.25f
C534 tb<5>.n279 VSS 7.82f
C535 tb<5>.n280 VSS 28.6f
C536 tb<5>.n281 VSS -7.6f
C537 tb<5>.n282 VSS 7.82f
C538 tb<5>.n283 VSS 32f
C539 tb<5>.n284 VSS -4.25f
C540 tb<5>.n285 VSS 7.82f
C541 tb<5>.n286 VSS 28.6f
C542 tb<5>.n287 VSS -7.6f
C543 tb<5>.n288 VSS 7.82f
C544 tb<5>.n289 VSS 32.2f
C545 tb<5>.n290 VSS -2.13f
C546 tb<5>.n291 VSS -0.85f
C547 tb<5>.n292 VSS -2.13f
C548 tb<5>.n293 VSS -1.33f
C549 tb<5>.n294 VSS 0.454f
C550 tb<5>.n295 VSS -30.6f
C551 tb<5>.n296 VSS -1.49f
C552 tb<5>.n297 VSS 31.6f
C553 tb<5>.n298 VSS -2.37f
C554 tb<5>.n299 VSS -0.413f
C555 tb<5>.n300 VSS -17.8f
C556 tb<5>.n301 VSS -17.3f
C557 tb<4>.n0 VSS -13.3f
C558 tb<4>.n1 VSS 1.55f
C559 tb<4>.n2 VSS 0.867f
C560 tb<4>.n3 VSS 1.39f
C561 tb<4>.n4 VSS -2.55f
C562 tb<4>.n5 VSS -9.34f
C563 tb<4>.n6 VSS 2.48f
C564 tb<4>.n7 VSS 1.21f
C565 tb<4>.n8 VSS 1.64f
C566 tb<4>.n9 VSS 0.867f
C567 tb<4>.n10 VSS 1.39f
C568 tb<4>.n11 VSS -2.55f
C569 tb<4>.n12 VSS -9.34f
C570 tb<4>.n13 VSS 2.48f
C571 tb<4>.n14 VSS 1.21f
C572 tb<4>.n15 VSS 1.64f
C573 tb<4>.n16 VSS 0.867f
C574 tb<4>.n17 VSS 1.39f
C575 tb<4>.n18 VSS -2.55f
C576 tb<4>.n19 VSS -9.34f
C577 tb<4>.n20 VSS 2.48f
C578 tb<4>.n21 VSS 1.21f
C579 tb<4>.n22 VSS 1.64f
C580 tb<4>.n23 VSS 0.867f
C581 tb<4>.n24 VSS 1.39f
C582 tb<4>.n25 VSS -2.55f
C583 tb<4>.n26 VSS -9.34f
C584 tb<4>.n27 VSS 2.48f
C585 tb<4>.n28 VSS 1.21f
C586 tb<4>.n29 VSS 1.64f
C587 tb<4>.n30 VSS 0.867f
C588 tb<4>.n31 VSS 1.39f
C589 tb<4>.n32 VSS -2.55f
C590 tb<4>.n33 VSS -9.34f
C591 tb<4>.n34 VSS 2.48f
C592 tb<4>.n35 VSS 1.21f
C593 tb<4>.n36 VSS 1.64f
C594 tb<4>.n37 VSS 0.867f
C595 tb<4>.n38 VSS 1.39f
C596 tb<4>.n39 VSS -2.55f
C597 tb<4>.n40 VSS -9.34f
C598 tb<4>.n41 VSS 2.48f
C599 tb<4>.n42 VSS 1.21f
C600 tb<4>.n43 VSS 1.64f
C601 tb<4>.n44 VSS 0.806f
C602 tb<4>.n45 VSS 0.694f
C603 tb<4>.n46 VSS 0.254f
C604 tb<4>.n47 VSS -0.153p
C605 tb<4>.n48 VSS 7.41f
C606 tb<4>.n49 VSS 13.7f
C607 tb<4>.n50 VSS 93.3f
C608 tb<4>.n51 VSS 93.3f
C609 tb<4>.n52 VSS -16.6f
C610 tb<4>.n53 VSS -1.15f
C611 tb<4>.n54 VSS 1.21f
C612 tb<4>.n55 VSS 2.48f
C613 tb<4>.n56 VSS -9.34f
C614 tb<4>.n57 VSS -2.55f
C615 tb<4>.n58 VSS 1.39f
C616 tb<4>.n59 VSS 0.867f
C617 tb<4>.n60 VSS 1.4f
C618 tb<4>.n61 VSS 1.21f
C619 tb<4>.n62 VSS 2.48f
C620 tb<4>.n63 VSS -9.34f
C621 tb<4>.n64 VSS -2.55f
C622 tb<4>.n65 VSS 1.39f
C623 tb<4>.n66 VSS 0.867f
C624 tb<4>.n67 VSS 1.4f
C625 tb<4>.n68 VSS 1.21f
C626 tb<4>.n69 VSS 2.48f
C627 tb<4>.n70 VSS -9.34f
C628 tb<4>.n71 VSS -2.55f
C629 tb<4>.n72 VSS 1.39f
C630 tb<4>.n73 VSS 0.867f
C631 tb<4>.n74 VSS 1.4f
C632 tb<4>.n75 VSS 1.21f
C633 tb<4>.n76 VSS 2.48f
C634 tb<4>.n77 VSS -9.34f
C635 tb<4>.n78 VSS -2.55f
C636 tb<4>.n79 VSS 1.39f
C637 tb<4>.n80 VSS 0.867f
C638 tb<4>.n81 VSS 1.4f
C639 tb<4>.n82 VSS 1.21f
C640 tb<4>.n83 VSS 2.48f
C641 tb<4>.n84 VSS -9.34f
C642 tb<4>.n85 VSS -2.55f
C643 tb<4>.n86 VSS 1.39f
C644 tb<4>.n87 VSS 0.867f
C645 tb<4>.n88 VSS 1.4f
C646 tb<4>.n89 VSS 1.21f
C647 tb<4>.n90 VSS 2.48f
C648 tb<4>.n91 VSS -9.34f
C649 tb<4>.n92 VSS -2.55f
C650 tb<4>.n93 VSS 1.33f
C651 tb<4>.n94 VSS 0.694f
C652 tb<4>.n95 VSS 0.234f
C653 tb<4>.n96 VSS -0.138p
C654 tb<4>.n97 VSS 0.905f
C655 tb<4>.n98 VSS 5.79f
C656 tb<4>.n99 VSS 4.74f
C657 t<1>.n0 VSS -0.634f
C658 t<1>.n1 VSS 2.68f
C659 t<1>.n2 VSS 0.29f
C660 t<1>.n3 VSS 0.406f
C661 t<1>.n4 VSS 0.376f
C662 tb<1>.n0 VSS 0.288f
C663 tb<1>.n1 VSS -0.629f
C664 tb<1>.n2 VSS 0.373f
C665 tb<1>.n3 VSS 0.403f
C666 tb<1>.n4 VSS 7.84f
C667 t<5>.n0 VSS -63.6f
C668 t<5>.n1 VSS -3.98f
C669 t<5>.n2 VSS 37.3f
C670 t<5>.n3 VSS -2.17f
C671 t<5>.n4 VSS 7.99f
C672 t<5>.n5 VSS 29.2f
C673 t<5>.n6 VSS 32.6f
C674 t<5>.n7 VSS -5.14f
C675 t<5>.n8 VSS 29.2f
C676 t<5>.n9 VSS 7.99f
C677 t<5>.n10 VSS -4.34f
C678 t<5>.n11 VSS -7.76f
C679 t<5>.n12 VSS 7.99f
C680 t<5>.n13 VSS -2.71f
C681 t<5>.n14 VSS 29.2f
C682 t<5>.n15 VSS 7.99f
C683 t<5>.n16 VSS -4.34f
C684 t<5>.n17 VSS -7.76f
C685 t<5>.n18 VSS 7.99f
C686 t<5>.n19 VSS -2.71f
C687 t<5>.n20 VSS 29.2f
C688 t<5>.n21 VSS 7.99f
C689 t<5>.n22 VSS -4.34f
C690 t<5>.n23 VSS -7.76f
C691 t<5>.n24 VSS 7.99f
C692 t<5>.n25 VSS -2.71f
C693 t<5>.n26 VSS 29.2f
C694 t<5>.n27 VSS 7.99f
C695 t<5>.n28 VSS -4.34f
C696 t<5>.n29 VSS -7.76f
C697 t<5>.n30 VSS 7.99f
C698 t<5>.n31 VSS -2.71f
C699 t<5>.n32 VSS 29.2f
C700 t<5>.n33 VSS 7.99f
C701 t<5>.n34 VSS -4.34f
C702 t<5>.n35 VSS -7.76f
C703 t<5>.n36 VSS 7.99f
C704 t<5>.n37 VSS -2.71f
C705 t<5>.n38 VSS 29.2f
C706 t<5>.n39 VSS 7.99f
C707 t<5>.n40 VSS -4.34f
C708 t<5>.n41 VSS -7.76f
C709 t<5>.n42 VSS 7.99f
C710 t<5>.n43 VSS -2.71f
C711 t<5>.n44 VSS 29.2f
C712 t<5>.n45 VSS 7.99f
C713 t<5>.n46 VSS 45.7f
C714 t<5>.n47 VSS 41.5f
C715 t<5>.n48 VSS -4.86f
C716 t<5>.n49 VSS -2.71f
C717 t<5>.n50 VSS -4.34f
C718 t<5>.n51 VSS 32.6f
C719 t<5>.n52 VSS 7.99f
C720 t<5>.n53 VSS -7.76f
C721 t<5>.n54 VSS 29.2f
C722 t<5>.n55 VSS -7.76f
C723 t<5>.n56 VSS -5.14f
C724 t<5>.n57 VSS -3.8f
C725 t<5>.n58 VSS 7.99f
C726 t<5>.n59 VSS -4.34f
C727 t<5>.n60 VSS 32.6f
C728 t<5>.n61 VSS -4.34f
C729 t<5>.n62 VSS 7.99f
C730 t<5>.n63 VSS 29.2f
C731 t<5>.n64 VSS -7.76f
C732 t<5>.n65 VSS 29.2f
C733 t<5>.n66 VSS 7.99f
C734 t<5>.n67 VSS -3.8f
C735 t<5>.n68 VSS -5.14f
C736 t<5>.n69 VSS -2.71f
C737 t<5>.n70 VSS -4.34f
C738 t<5>.n71 VSS 32.6f
C739 t<5>.n72 VSS 7.99f
C740 t<5>.n73 VSS -7.76f
C741 t<5>.n74 VSS 29.2f
C742 t<5>.n75 VSS -7.76f
C743 t<5>.n76 VSS -5.14f
C744 t<5>.n77 VSS -3.8f
C745 t<5>.n78 VSS 7.99f
C746 t<5>.n79 VSS -4.34f
C747 t<5>.n80 VSS 32.6f
C748 t<5>.n81 VSS -4.34f
C749 t<5>.n82 VSS 7.99f
C750 t<5>.n83 VSS 29.2f
C751 t<5>.n84 VSS -7.76f
C752 t<5>.n85 VSS 29.2f
C753 t<5>.n86 VSS 7.99f
C754 t<5>.n87 VSS -3.8f
C755 t<5>.n88 VSS -5.14f
C756 t<5>.n89 VSS -2.71f
C757 t<5>.n90 VSS -4.34f
C758 t<5>.n91 VSS 32.6f
C759 t<5>.n92 VSS 7.99f
C760 t<5>.n93 VSS -7.76f
C761 t<5>.n94 VSS 29.2f
C762 t<5>.n95 VSS -7.76f
C763 t<5>.n96 VSS -5.14f
C764 t<5>.n97 VSS -3.8f
C765 t<5>.n98 VSS 7.99f
C766 t<5>.n99 VSS -4.34f
C767 t<5>.n100 VSS 32.6f
C768 t<5>.n101 VSS -4.34f
C769 t<5>.n102 VSS 7.99f
C770 t<5>.n103 VSS 29.2f
C771 t<5>.n104 VSS -7.76f
C772 t<5>.n105 VSS 29.2f
C773 t<5>.n106 VSS 7.99f
C774 t<5>.n107 VSS -3.8f
C775 t<5>.n108 VSS -5.14f
C776 t<5>.n109 VSS -2.71f
C777 t<5>.n110 VSS -4.34f
C778 t<5>.n111 VSS 32.6f
C779 t<5>.n112 VSS 7.99f
C780 t<5>.n113 VSS -7.76f
C781 t<5>.n114 VSS 29.2f
C782 t<5>.n115 VSS -7.76f
C783 t<5>.n116 VSS -5.14f
C784 t<5>.n117 VSS -3.8f
C785 t<5>.n118 VSS 7.99f
C786 t<5>.n119 VSS -4.34f
C787 t<5>.n120 VSS 32.6f
C788 t<5>.n121 VSS -4.34f
C789 t<5>.n122 VSS -3.8f
C790 t<5>.n123 VSS -25f
C791 t<5>.n124 VSS -6.13f
C792 t<5>.n125 VSS -7.76f
C793 t<5>.n126 VSS 29.2f
C794 t<5>.n127 VSS 7.99f
C795 t<5>.n128 VSS -3.8f
C796 t<5>.n129 VSS -5.14f
C797 t<5>.n130 VSS -2.71f
C798 t<5>.n131 VSS -4.34f
C799 t<5>.n132 VSS 32.6f
C800 t<5>.n133 VSS 7.99f
C801 t<5>.n134 VSS -7.76f
C802 t<5>.n135 VSS 29.2f
C803 t<5>.n136 VSS -7.76f
C804 t<5>.n137 VSS -5.14f
C805 t<5>.n138 VSS -3.8f
C806 t<5>.n139 VSS 7.99f
C807 t<5>.n140 VSS -4.34f
C808 t<5>.n141 VSS 32.6f
C809 t<5>.n142 VSS -4.34f
C810 t<5>.n143 VSS 7.99f
C811 t<5>.n144 VSS 29.2f
C812 t<5>.n145 VSS -7.76f
C813 t<5>.n146 VSS 29.2f
C814 t<5>.n147 VSS 7.99f
C815 t<5>.n148 VSS -3.8f
C816 t<5>.n149 VSS -5.14f
C817 t<5>.n150 VSS -2.71f
C818 t<5>.n151 VSS -4.34f
C819 t<5>.n152 VSS 32.6f
C820 t<5>.n153 VSS 7.99f
C821 t<5>.n154 VSS -7.76f
C822 t<5>.n155 VSS 29.2f
C823 t<5>.n156 VSS -7.76f
C824 t<5>.n157 VSS -5.14f
C825 t<5>.n158 VSS -3.8f
C826 t<5>.n159 VSS 7.99f
C827 t<5>.n160 VSS -4.34f
C828 t<5>.n161 VSS 32.6f
C829 t<5>.n162 VSS -4.34f
C830 t<5>.n163 VSS 7.99f
C831 t<5>.n164 VSS 29.2f
C832 t<5>.n165 VSS -7.76f
C833 t<5>.n166 VSS 29.2f
C834 t<5>.n167 VSS 7.99f
C835 t<5>.n168 VSS -3.8f
C836 t<5>.n169 VSS -5.14f
C837 t<5>.n170 VSS -2.71f
C838 t<5>.n171 VSS -4.34f
C839 t<5>.n172 VSS 32.6f
C840 t<5>.n173 VSS 7.99f
C841 t<5>.n174 VSS -7.76f
C842 t<5>.n175 VSS 29.2f
C843 t<5>.n176 VSS -7.76f
C844 t<5>.n177 VSS -3.8f
C845 t<5>.n178 VSS 7.99f
C846 t<5>.n179 VSS -4.34f
C847 t<5>.n180 VSS -2.71f
C848 t<5>.n181 VSS -4.34f
C849 t<5>.n182 VSS 7.99f
C850 t<5>.n183 VSS 7.99f
C851 t<5>.n184 VSS -7.76f
C852 t<5>.n185 VSS 29.2f
C853 t<5>.n186 VSS -7.76f
C854 t<5>.n187 VSS -3.8f
C855 t<5>.n188 VSS -5.14f
C856 t<5>.n189 VSS -2.52f
C857 t<5>.n190 VSS -4.15f
C858 t<5>.n191 VSS -2.17f
C859 t<5>.n192 VSS 8.99f
C860 t<5>.n193 VSS -0.796f
C861 t<5>.n194 VSS -5.95f
C862 t<5>.n195 VSS -1.43f
C863 t<5>.n196 VSS -9.86f
C864 t<5>.n197 VSS -11.9f
C865 t<5>.n198 VSS -10.5f
C866 t<5>.n199 VSS 35.1f
C867 t<5>.n200 VSS -0.116p
C868 t<5>.n201 VSS -0.181p
C869 t<5>.n202 VSS 52f
C870 t<5>.n203 VSS 3.6f
C871 t<5>.n204 VSS -3.8f
C872 t<5>.n205 VSS -7.76f
C873 t<5>.n206 VSS 29.2f
C874 t<5>.n207 VSS 7.99f
C875 t<5>.n208 VSS -4.34f
C876 t<5>.n209 VSS -2.71f
C877 t<5>.n210 VSS -4.37f
C878 t<5>.n211 VSS -3.8f
C879 t<5>.n212 VSS -7.76f
C880 t<5>.n213 VSS 29.2f
C881 t<5>.n214 VSS 7.99f
C882 t<5>.n215 VSS -4.34f
C883 t<5>.n216 VSS -2.71f
C884 t<5>.n217 VSS -4.37f
C885 t<5>.n218 VSS -3.8f
C886 t<5>.n219 VSS -7.76f
C887 t<5>.n220 VSS 29.2f
C888 t<5>.n221 VSS 7.99f
C889 t<5>.n222 VSS -4.34f
C890 t<5>.n223 VSS -2.71f
C891 t<5>.n224 VSS -4.37f
C892 t<5>.n225 VSS -3.8f
C893 t<5>.n226 VSS -7.76f
C894 t<5>.n227 VSS 29.2f
C895 t<5>.n228 VSS 7.99f
C896 t<5>.n229 VSS -4.34f
C897 t<5>.n230 VSS -2.71f
C898 t<5>.n231 VSS -4.37f
C899 t<5>.n232 VSS -3.8f
C900 t<5>.n233 VSS -7.76f
C901 t<5>.n234 VSS 29.2f
C902 t<5>.n235 VSS 7.99f
C903 t<5>.n236 VSS -4.34f
C904 t<5>.n237 VSS -2.71f
C905 t<5>.n238 VSS -4.37f
C906 t<5>.n239 VSS -3.8f
C907 t<5>.n240 VSS -7.76f
C908 t<5>.n241 VSS 29.2f
C909 t<5>.n242 VSS 7.99f
C910 t<5>.n243 VSS -4.34f
C911 t<5>.n244 VSS -2.71f
C912 t<5>.n245 VSS -4.37f
C913 t<5>.n246 VSS -3.8f
C914 t<5>.n247 VSS -7.76f
C915 t<5>.n248 VSS 29.2f
C916 t<5>.n249 VSS 7.99f
C917 t<5>.n250 VSS -4.34f
C918 t<5>.n251 VSS -2.71f
C919 t<5>.n252 VSS -4.37f
C920 t<5>.n253 VSS -3.8f
C921 t<5>.n254 VSS -7.76f
C922 t<5>.n255 VSS 29.2f
C923 t<5>.n256 VSS 7.99f
C924 t<5>.n257 VSS -4.34f
C925 t<5>.n258 VSS -2.71f
C926 t<5>.n259 VSS -4.37f
C927 t<5>.n260 VSS -3.8f
C928 t<5>.n261 VSS -7.76f
C929 t<5>.n262 VSS 29.2f
C930 t<5>.n263 VSS 7.99f
C931 t<5>.n264 VSS -4.34f
C932 t<5>.n265 VSS -2.71f
C933 t<5>.n266 VSS -4.37f
C934 t<5>.n267 VSS -3.8f
C935 t<5>.n268 VSS -7.76f
C936 t<5>.n269 VSS 29.2f
C937 t<5>.n270 VSS 7.99f
C938 t<5>.n271 VSS -4.34f
C939 t<5>.n272 VSS -2.71f
C940 t<5>.n273 VSS -4.37f
C941 t<5>.n274 VSS -3.8f
C942 t<5>.n275 VSS -7.76f
C943 t<5>.n276 VSS 29.2f
C944 t<5>.n277 VSS 7.99f
C945 t<5>.n278 VSS -4.34f
C946 t<5>.n279 VSS -2.71f
C947 t<5>.n280 VSS -4.37f
C948 t<5>.n281 VSS -3.8f
C949 t<5>.n282 VSS -7.76f
C950 t<5>.n283 VSS 29.2f
C951 t<5>.n284 VSS 7.99f
C952 t<5>.n285 VSS -4.34f
C953 t<5>.n286 VSS -2.71f
C954 t<5>.n287 VSS -4.37f
C955 t<5>.n288 VSS -3.8f
C956 t<5>.n289 VSS -7.76f
C957 t<5>.n290 VSS 29.2f
C958 t<5>.n291 VSS 7.99f
C959 t<5>.n292 VSS -4.34f
C960 t<5>.n293 VSS -2.71f
C961 t<5>.n294 VSS -4.37f
C962 t<5>.n295 VSS -3.8f
C963 t<5>.n296 VSS -7.76f
C964 t<5>.n297 VSS 29.2f
C965 t<5>.n298 VSS 7.99f
C966 t<5>.n299 VSS -4.15f
C967 t<5>.n300 VSS -2.17f
C968 t<5>.n301 VSS -0.732f
C969 t<5>.n302 VSS -2.88f
C970 t<5>.n303 VSS 48.9f
C971 t<5>.n304 VSS 29.2f
C972 t<5>.n305 VSS -7.76f
C973 t<5>.n306 VSS 7.99f
C974 t<5>.n307 VSS 32.6f
C975 t<5>.n308 VSS -4.34f
C976 t<5>.n309 VSS 7.99f
C977 t<5>.n310 VSS 29.2f
C978 t<5>.n311 VSS -7.76f
C979 t<5>.n312 VSS 7.99f
C980 t<5>.n313 VSS 32.6f
C981 t<5>.n314 VSS -4.34f
C982 t<5>.n315 VSS 7.99f
C983 t<5>.n316 VSS 29.2f
C984 t<5>.n317 VSS -7.76f
C985 t<5>.n318 VSS 7.99f
C986 t<5>.n319 VSS 32.6f
C987 t<5>.n320 VSS -4.34f
C988 t<5>.n321 VSS 7.99f
C989 t<5>.n322 VSS 29.2f
C990 t<5>.n323 VSS -7.76f
C991 t<5>.n324 VSS 7.99f
C992 t<5>.n325 VSS 32.6f
C993 t<5>.n326 VSS -4.34f
C994 t<5>.n327 VSS 7.99f
C995 t<5>.n328 VSS 29.2f
C996 t<5>.n329 VSS -7.76f
C997 t<5>.n330 VSS 7.99f
C998 t<5>.n331 VSS 32.6f
C999 t<5>.n332 VSS -4.34f
C1000 t<5>.n333 VSS 7.99f
C1001 t<5>.n334 VSS 29.2f
C1002 t<5>.n335 VSS -7.76f
C1003 t<5>.n336 VSS 7.99f
C1004 t<5>.n337 VSS 32.6f
C1005 t<5>.n338 VSS -4.34f
C1006 t<5>.n339 VSS 7.99f
C1007 t<5>.n340 VSS 29.2f
C1008 t<5>.n341 VSS -7.76f
C1009 t<5>.n342 VSS 7.99f
C1010 t<5>.n343 VSS 32.6f
C1011 t<5>.n344 VSS -4.34f
C1012 t<5>.n345 VSS 7.99f
C1013 t<5>.n346 VSS 29.2f
C1014 t<5>.n347 VSS -7.76f
C1015 t<5>.n348 VSS 7.99f
C1016 t<5>.n349 VSS 32.6f
C1017 t<5>.n350 VSS -4.34f
C1018 t<5>.n351 VSS 7.99f
C1019 t<5>.n352 VSS 29.2f
C1020 t<5>.n353 VSS -7.76f
C1021 t<5>.n354 VSS 7.99f
C1022 t<5>.n355 VSS 32.6f
C1023 t<5>.n356 VSS -4.34f
C1024 t<5>.n357 VSS 7.99f
C1025 t<5>.n358 VSS 29.2f
C1026 t<5>.n359 VSS -7.76f
C1027 t<5>.n360 VSS 7.99f
C1028 t<5>.n361 VSS 32.6f
C1029 t<5>.n362 VSS -4.34f
C1030 t<5>.n363 VSS 7.99f
C1031 t<5>.n364 VSS 29.2f
C1032 t<5>.n365 VSS -7.76f
C1033 t<5>.n366 VSS 7.99f
C1034 t<5>.n367 VSS 32.6f
C1035 t<5>.n368 VSS -4.34f
C1036 t<5>.n369 VSS 7.99f
C1037 t<5>.n370 VSS 29.2f
C1038 t<5>.n371 VSS -7.76f
C1039 t<5>.n372 VSS 7.99f
C1040 t<5>.n373 VSS 32.6f
C1041 t<5>.n374 VSS -4.34f
C1042 t<5>.n375 VSS 7.99f
C1043 t<5>.n376 VSS 29.2f
C1044 t<5>.n377 VSS -7.76f
C1045 t<5>.n378 VSS 7.99f
C1046 t<5>.n379 VSS 32.6f
C1047 t<5>.n380 VSS -4.34f
C1048 t<5>.n381 VSS 7.99f
C1049 t<5>.n382 VSS 29.2f
C1050 t<5>.n383 VSS -7.76f
C1051 t<5>.n384 VSS 7.99f
C1052 t<5>.n385 VSS 32.8f
C1053 t<5>.n386 VSS -2.17f
C1054 t<5>.n387 VSS -0.868f
C1055 t<5>.n388 VSS -2.17f
C1056 t<5>.n389 VSS -1.36f
C1057 t<5>.n390 VSS 0.463f
C1058 t<5>.n391 VSS -31.2f
C1059 t<5>.n392 VSS -1.52f
C1060 t<5>.n393 VSS 32.3f
C1061 t<5>.n394 VSS -2.42f
C1062 t<5>.n395 VSS -0.422f
C1063 t<5>.n396 VSS -18.1f
C1064 t<5>.n397 VSS -17.7f
C1065 t<3>.n0 VSS 2.8f
C1066 t<3>.n1 VSS 5.22f
C1067 t<3>.n2 VSS 0.048f
C1068 t<3>.n3 VSS 0.242f
C1069 t<3>.n4 VSS 0.0698f
C1070 t<3>.n5 VSS -0.0935f
C1071 t<3>.n6 VSS 0.349f
C1072 t<3>.n7 VSS 0.623f
C1073 t<3>.n8 VSS -0.642f
C1074 t<3>.n9 VSS 0.218f
C1075 t<3>.n10 VSS 0.391f
C1076 t<3>.n11 VSS -3.34f
C1077 t<3>.n12 VSS -3.68f
C1078 t<3>.n13 VSS -2.62f
C1079 t<3>.n14 VSS 0.349f
C1080 t<3>.n15 VSS -0.642f
C1081 t<3>.n16 VSS -2.35f
C1082 t<3>.n17 VSS 0.623f
C1083 t<3>.n18 VSS -2.35f
C1084 t<3>.n19 VSS -0.642f
C1085 t<3>.n20 VSS 0.305f
C1086 t<3>.n21 VSS 0.413f
C1087 t<3>.n22 VSS 0.218f
C1088 t<3>.n23 VSS 0.349f
C1089 t<3>.n24 VSS -2.62f
C1090 t<3>.n25 VSS -0.67f
C1091 t<3>.n26 VSS 0.174f
C1092 t<3>.n27 VSS -3.37f
C1093 t<3>.n28 VSS 0.0698f
C1094 t<3>.n29 VSS 0.256f
C1095 t<3>.n30 VSS 0.449f
C1096 t<3>.n31 VSS -1.81f
C1097 t<3>.n32 VSS -4.89f
C1098 t<3>.n33 VSS 0.253f
C1099 t<3>.n34 VSS 2.97f
C1100 t<3>.n35 VSS 9.52f
C1101 t<3>.n36 VSS 14.3f
C1102 t<3>.n37 VSS -0.191f
C1103 t<3>.n38 VSS -5f
C1104 t<3>.n39 VSS -1.66f
C1105 t<3>.n40 VSS 0.277f
C1106 t<3>.n41 VSS 0.174f
C1107 t<3>.n42 VSS 0.0698f
C1108 t<3>.n43 VSS -11.3f
C1109 t<3>.n44 VSS 0.0791f
C1110 t<3>.n45 VSS 1.45f
C1111 t<3>.n46 VSS 1.35f
C1112 tb<3>.n0 VSS 2.78f
C1113 tb<3>.n1 VSS -3.31f
C1114 tb<3>.n2 VSS 0.388f
C1115 tb<3>.n3 VSS 0.216f
C1116 tb<3>.n4 VSS 0.346f
C1117 tb<3>.n5 VSS -0.637f
C1118 tb<3>.n6 VSS -2.33f
C1119 tb<3>.n7 VSS 0.619f
C1120 tb<3>.n8 VSS 0.303f
C1121 tb<3>.n9 VSS 0.41f
C1122 tb<3>.n10 VSS 0.216f
C1123 tb<3>.n11 VSS 0.346f
C1124 tb<3>.n12 VSS -0.0929f
C1125 tb<3>.n13 VSS -3.35f
C1126 tb<3>.n14 VSS 0.0693f
C1127 tb<3>.n15 VSS -11.2f
C1128 tb<3>.n16 VSS -1.79f
C1129 tb<3>.n17 VSS 0.24f
C1130 tb<3>.n18 VSS -4.61f
C1131 tb<3>.n19 VSS 2.95f
C1132 tb<3>.n20 VSS 0.0476f
C1133 tb<3>.n21 VSS 5.18f
C1134 tb<3>.n22 VSS 23.3f
C1135 tb<3>.n23 VSS 23.3f
C1136 tb<3>.n24 VSS -0.19f
C1137 tb<3>.n25 VSS -6.61f
C1138 tb<3>.n26 VSS 0.275f
C1139 tb<3>.n27 VSS 0.173f
C1140 tb<3>.n28 VSS 0.0693f
C1141 tb<3>.n29 VSS -11.2f
C1142 tb<3>.n30 VSS 0.0786f
C1143 tb<3>.n31 VSS 1.44f
C1144 tb<3>.n32 VSS 1.34f
C1145 t<6>.n0 VSS -16.1f
C1146 t<6>.n1 VSS -2.42f
C1147 t<6>.n2 VSS -0.679f
C1148 t<6>.n3 VSS -0.221f
C1149 t<6>.n4 VSS -2.23f
C1150 t<6>.n5 VSS -0.952f
C1151 t<6>.n6 VSS -1.97f
C1152 t<6>.n7 VSS -0.965f
C1153 t<6>.n8 VSS 8.3f
C1154 t<6>.n9 VSS -1.31f
C1155 t<6>.n10 VSS 7.43f
C1156 t<6>.n11 VSS 2.03f
C1157 t<6>.n12 VSS -1.1f
C1158 t<6>.n13 VSS -1.97f
C1159 t<6>.n14 VSS -0.965f
C1160 t<6>.n15 VSS 8.3f
C1161 t<6>.n16 VSS -1.31f
C1162 t<6>.n17 VSS 7.43f
C1163 t<6>.n18 VSS 2.03f
C1164 t<6>.n19 VSS -1.1f
C1165 t<6>.n20 VSS -1.97f
C1166 t<6>.n21 VSS -0.965f
C1167 t<6>.n22 VSS 8.3f
C1168 t<6>.n23 VSS -1.31f
C1169 t<6>.n24 VSS 7.43f
C1170 t<6>.n25 VSS 2.03f
C1171 t<6>.n26 VSS -1.1f
C1172 t<6>.n27 VSS -1.97f
C1173 t<6>.n28 VSS -0.965f
C1174 t<6>.n29 VSS 8.3f
C1175 t<6>.n30 VSS -1.31f
C1176 t<6>.n31 VSS 7.43f
C1177 t<6>.n32 VSS 2.03f
C1178 t<6>.n33 VSS -1.1f
C1179 t<6>.n34 VSS -1.97f
C1180 t<6>.n35 VSS -0.965f
C1181 t<6>.n36 VSS 8.3f
C1182 t<6>.n37 VSS -1.31f
C1183 t<6>.n38 VSS 7.43f
C1184 t<6>.n39 VSS 2.03f
C1185 t<6>.n40 VSS -1.1f
C1186 t<6>.n41 VSS -1.97f
C1187 t<6>.n42 VSS -0.965f
C1188 t<6>.n43 VSS 8.3f
C1189 t<6>.n44 VSS -1.31f
C1190 t<6>.n45 VSS 7.43f
C1191 t<6>.n46 VSS 2.03f
C1192 t<6>.n47 VSS -1.1f
C1193 t<6>.n48 VSS -1.97f
C1194 t<6>.n49 VSS -0.965f
C1195 t<6>.n50 VSS 8.3f
C1196 t<6>.n51 VSS -1.31f
C1197 t<6>.n52 VSS 7.43f
C1198 t<6>.n53 VSS 2.03f
C1199 t<6>.n54 VSS -1.1f
C1200 t<6>.n55 VSS -1.97f
C1201 t<6>.n56 VSS -0.965f
C1202 t<6>.n57 VSS 8.3f
C1203 t<6>.n58 VSS -1.31f
C1204 t<6>.n59 VSS 7.43f
C1205 t<6>.n60 VSS 2.03f
C1206 t<6>.n61 VSS -1.1f
C1207 t<6>.n62 VSS -1.97f
C1208 t<6>.n63 VSS -0.965f
C1209 t<6>.n64 VSS 8.3f
C1210 t<6>.n65 VSS -1.31f
C1211 t<6>.n66 VSS 7.43f
C1212 t<6>.n67 VSS 2.03f
C1213 t<6>.n68 VSS -1.1f
C1214 t<6>.n69 VSS -1.97f
C1215 t<6>.n70 VSS -0.965f
C1216 t<6>.n71 VSS 8.3f
C1217 t<6>.n72 VSS -1.31f
C1218 t<6>.n73 VSS 7.43f
C1219 t<6>.n74 VSS 2.03f
C1220 t<6>.n75 VSS -1.1f
C1221 t<6>.n76 VSS -1.97f
C1222 t<6>.n77 VSS -0.965f
C1223 t<6>.n78 VSS 8.3f
C1224 t<6>.n79 VSS -1.31f
C1225 t<6>.n80 VSS 7.43f
C1226 t<6>.n81 VSS 2.03f
C1227 t<6>.n82 VSS -1.1f
C1228 t<6>.n83 VSS -1.97f
C1229 t<6>.n84 VSS -0.965f
C1230 t<6>.n85 VSS 8.3f
C1231 t<6>.n86 VSS -1.31f
C1232 t<6>.n87 VSS 7.43f
C1233 t<6>.n88 VSS 2.03f
C1234 t<6>.n89 VSS -1.1f
C1235 t<6>.n90 VSS -1.97f
C1236 t<6>.n91 VSS -0.965f
C1237 t<6>.n92 VSS 8.3f
C1238 t<6>.n93 VSS -1.31f
C1239 t<6>.n94 VSS 7.43f
C1240 t<6>.n95 VSS 2.03f
C1241 t<6>.n96 VSS -1.1f
C1242 t<6>.n97 VSS -1.97f
C1243 t<6>.n98 VSS -0.965f
C1244 t<6>.n99 VSS 8.3f
C1245 t<6>.n100 VSS -1.31f
C1246 t<6>.n101 VSS 7.43f
C1247 t<6>.n102 VSS 2.03f
C1248 t<6>.n103 VSS -1.1f
C1249 t<6>.n104 VSS -1.97f
C1250 t<6>.n105 VSS -0.965f
C1251 t<6>.n106 VSS 8.3f
C1252 t<6>.n107 VSS -1.31f
C1253 t<6>.n108 VSS 7.43f
C1254 t<6>.n109 VSS 12.4f
C1255 t<6>.n110 VSS 13.9f
C1256 t<6>.n111 VSS 0.72f
C1257 t<6>.n112 VSS -0.965f
C1258 t<6>.n113 VSS -1.97f
C1259 t<6>.n114 VSS 7.43f
C1260 t<6>.n115 VSS -1.97f
C1261 t<6>.n116 VSS 2.03f
C1262 t<6>.n117 VSS 2.03f
C1263 t<6>.n118 VSS -1.1f
C1264 t<6>.n119 VSS -0.69f
C1265 t<6>.n120 VSS -1.1f
C1266 t<6>.n121 VSS 2.03f
C1267 t<6>.n122 VSS 7.43f
C1268 t<6>.n123 VSS -1.97f
C1269 t<6>.n124 VSS 7.43f
C1270 t<6>.n125 VSS 2.03f
C1271 t<6>.n126 VSS 2.03f
C1272 t<6>.n127 VSS 8.3f
C1273 t<6>.n128 VSS -1.1f
C1274 t<6>.n129 VSS -0.69f
C1275 t<6>.n130 VSS -1.31f
C1276 t<6>.n131 VSS -0.965f
C1277 t<6>.n132 VSS -1.97f
C1278 t<6>.n133 VSS 7.43f
C1279 t<6>.n134 VSS -1.97f
C1280 t<6>.n135 VSS 2.03f
C1281 t<6>.n136 VSS 2.03f
C1282 t<6>.n137 VSS -1.1f
C1283 t<6>.n138 VSS -0.69f
C1284 t<6>.n139 VSS -1.1f
C1285 t<6>.n140 VSS 2.03f
C1286 t<6>.n141 VSS 7.43f
C1287 t<6>.n142 VSS -1.97f
C1288 t<6>.n143 VSS 7.43f
C1289 t<6>.n144 VSS 2.03f
C1290 t<6>.n145 VSS 2.03f
C1291 t<6>.n146 VSS 8.3f
C1292 t<6>.n147 VSS -1.1f
C1293 t<6>.n148 VSS -0.69f
C1294 t<6>.n149 VSS -1.31f
C1295 t<6>.n150 VSS -0.965f
C1296 t<6>.n151 VSS -1.97f
C1297 t<6>.n152 VSS 7.43f
C1298 t<6>.n153 VSS -1.97f
C1299 t<6>.n154 VSS 2.03f
C1300 t<6>.n155 VSS 2.03f
C1301 t<6>.n156 VSS -1.1f
C1302 t<6>.n157 VSS -0.69f
C1303 t<6>.n158 VSS -1.1f
C1304 t<6>.n159 VSS 2.03f
C1305 t<6>.n160 VSS 7.43f
C1306 t<6>.n161 VSS -1.97f
C1307 t<6>.n162 VSS 7.43f
C1308 t<6>.n163 VSS 2.03f
C1309 t<6>.n164 VSS 2.03f
C1310 t<6>.n165 VSS 8.3f
C1311 t<6>.n166 VSS -1.1f
C1312 t<6>.n167 VSS -0.69f
C1313 t<6>.n168 VSS -1.31f
C1314 t<6>.n169 VSS -0.965f
C1315 t<6>.n170 VSS -1.97f
C1316 t<6>.n171 VSS 7.43f
C1317 t<6>.n172 VSS -1.97f
C1318 t<6>.n173 VSS 2.03f
C1319 t<6>.n174 VSS 2.03f
C1320 t<6>.n175 VSS -1.1f
C1321 t<6>.n176 VSS -0.69f
C1322 t<6>.n177 VSS -1.1f
C1323 t<6>.n178 VSS 2.03f
C1324 t<6>.n179 VSS 7.43f
C1325 t<6>.n180 VSS -1.97f
C1326 t<6>.n181 VSS 7.43f
C1327 t<6>.n182 VSS 2.03f
C1328 t<6>.n183 VSS 2.03f
C1329 t<6>.n184 VSS 8.3f
C1330 t<6>.n185 VSS -1.1f
C1331 t<6>.n186 VSS -0.69f
C1332 t<6>.n187 VSS -1.31f
C1333 t<6>.n188 VSS -0.965f
C1334 t<6>.n189 VSS -1.97f
C1335 t<6>.n190 VSS 7.43f
C1336 t<6>.n191 VSS -1.97f
C1337 t<6>.n192 VSS 2.03f
C1338 t<6>.n193 VSS 2.03f
C1339 t<6>.n194 VSS -1.1f
C1340 t<6>.n195 VSS -0.69f
C1341 t<6>.n196 VSS -1.1f
C1342 t<6>.n197 VSS 2.03f
C1343 t<6>.n198 VSS 7.43f
C1344 t<6>.n199 VSS -1.97f
C1345 t<6>.n200 VSS 7.43f
C1346 t<6>.n201 VSS 2.03f
C1347 t<6>.n202 VSS 2.03f
C1348 t<6>.n203 VSS 8.3f
C1349 t<6>.n204 VSS -1.1f
C1350 t<6>.n205 VSS -0.69f
C1351 t<6>.n206 VSS -1.31f
C1352 t<6>.n207 VSS -0.965f
C1353 t<6>.n208 VSS -1.97f
C1354 t<6>.n209 VSS 7.43f
C1355 t<6>.n210 VSS -1.97f
C1356 t<6>.n211 VSS 2.03f
C1357 t<6>.n212 VSS 2.03f
C1358 t<6>.n213 VSS -1.1f
C1359 t<6>.n214 VSS -0.69f
C1360 t<6>.n215 VSS -1.1f
C1361 t<6>.n216 VSS 2.03f
C1362 t<6>.n217 VSS 7.43f
C1363 t<6>.n218 VSS -1.97f
C1364 t<6>.n219 VSS 7.43f
C1365 t<6>.n220 VSS 2.03f
C1366 t<6>.n221 VSS 2.03f
C1367 t<6>.n222 VSS 8.3f
C1368 t<6>.n223 VSS -1.1f
C1369 t<6>.n224 VSS -0.69f
C1370 t<6>.n225 VSS -1.31f
C1371 t<6>.n226 VSS -0.965f
C1372 t<6>.n227 VSS -1.97f
C1373 t<6>.n228 VSS 7.43f
C1374 t<6>.n229 VSS -1.97f
C1375 t<6>.n230 VSS 2.03f
C1376 t<6>.n231 VSS 2.03f
C1377 t<6>.n232 VSS -1.1f
C1378 t<6>.n233 VSS -0.69f
C1379 t<6>.n234 VSS -1.1f
C1380 t<6>.n235 VSS 2.03f
C1381 t<6>.n236 VSS 7.43f
C1382 t<6>.n237 VSS -1.97f
C1383 t<6>.n238 VSS 7.43f
C1384 t<6>.n239 VSS 2.03f
C1385 t<6>.n240 VSS 2.03f
C1386 t<6>.n241 VSS 8.3f
C1387 t<6>.n242 VSS -1.1f
C1388 t<6>.n243 VSS -0.69f
C1389 t<6>.n244 VSS -1.31f
C1390 t<6>.n245 VSS -0.965f
C1391 t<6>.n246 VSS -1.97f
C1392 t<6>.n247 VSS 7.43f
C1393 t<6>.n248 VSS -1.97f
C1394 t<6>.n249 VSS 2.03f
C1395 t<6>.n250 VSS 2.03f
C1396 t<6>.n251 VSS -1.1f
C1397 t<6>.n252 VSS -0.69f
C1398 t<6>.n253 VSS -1.1f
C1399 t<6>.n254 VSS 2.03f
C1400 t<6>.n255 VSS 7.43f
C1401 t<6>.n256 VSS -1.97f
C1402 t<6>.n257 VSS 7.43f
C1403 t<6>.n258 VSS 2.03f
C1404 t<6>.n259 VSS 2.03f
C1405 t<6>.n260 VSS 8.3f
C1406 t<6>.n261 VSS -1.1f
C1407 t<6>.n262 VSS -0.69f
C1408 t<6>.n263 VSS -1.31f
C1409 t<6>.n264 VSS -0.965f
C1410 t<6>.n265 VSS -1.97f
C1411 t<6>.n266 VSS 7.43f
C1412 t<6>.n267 VSS -1.97f
C1413 t<6>.n268 VSS 2.03f
C1414 t<6>.n269 VSS 2.03f
C1415 t<6>.n270 VSS -1.1f
C1416 t<6>.n271 VSS -0.69f
C1417 t<6>.n272 VSS -1.1f
C1418 t<6>.n273 VSS 2.03f
C1419 t<6>.n274 VSS 7.43f
C1420 t<6>.n275 VSS -1.97f
C1421 t<6>.n276 VSS 7.43f
C1422 t<6>.n277 VSS 2.03f
C1423 t<6>.n278 VSS 2.03f
C1424 t<6>.n279 VSS 8.3f
C1425 t<6>.n280 VSS -1.1f
C1426 t<6>.n281 VSS -0.69f
C1427 t<6>.n282 VSS -1.31f
C1428 t<6>.n283 VSS -0.965f
C1429 t<6>.n284 VSS -1.97f
C1430 t<6>.n285 VSS 7.43f
C1431 t<6>.n286 VSS -1.97f
C1432 t<6>.n287 VSS 2.03f
C1433 t<6>.n288 VSS 2.03f
C1434 t<6>.n289 VSS -1.1f
C1435 t<6>.n290 VSS -0.69f
C1436 t<6>.n291 VSS -1.1f
C1437 t<6>.n292 VSS 2.03f
C1438 t<6>.n293 VSS 7.43f
C1439 t<6>.n294 VSS -1.97f
C1440 t<6>.n295 VSS 7.43f
C1441 t<6>.n296 VSS 2.03f
C1442 t<6>.n297 VSS 2.03f
C1443 t<6>.n298 VSS 8.3f
C1444 t<6>.n299 VSS -1.1f
C1445 t<6>.n300 VSS -0.69f
C1446 t<6>.n301 VSS -1.31f
C1447 t<6>.n302 VSS -0.965f
C1448 t<6>.n303 VSS -1.97f
C1449 t<6>.n304 VSS 7.43f
C1450 t<6>.n305 VSS -1.97f
C1451 t<6>.n306 VSS 2.03f
C1452 t<6>.n307 VSS 2.03f
C1453 t<6>.n308 VSS -1.1f
C1454 t<6>.n309 VSS -0.69f
C1455 t<6>.n310 VSS -1.1f
C1456 t<6>.n311 VSS 2.03f
C1457 t<6>.n312 VSS 7.43f
C1458 t<6>.n313 VSS -1.97f
C1459 t<6>.n314 VSS 7.43f
C1460 t<6>.n315 VSS 2.03f
C1461 t<6>.n316 VSS 2.03f
C1462 t<6>.n317 VSS 8.3f
C1463 t<6>.n318 VSS -1.1f
C1464 t<6>.n319 VSS -0.69f
C1465 t<6>.n320 VSS -1.31f
C1466 t<6>.n321 VSS -0.965f
C1467 t<6>.n322 VSS -1.97f
C1468 t<6>.n323 VSS 7.43f
C1469 t<6>.n324 VSS -1.97f
C1470 t<6>.n325 VSS 2.03f
C1471 t<6>.n326 VSS 2.03f
C1472 t<6>.n327 VSS -1.1f
C1473 t<6>.n328 VSS -0.69f
C1474 t<6>.n329 VSS -1.1f
C1475 t<6>.n330 VSS 2.03f
C1476 t<6>.n331 VSS 7.43f
C1477 t<6>.n332 VSS -1.97f
C1478 t<6>.n333 VSS 7.43f
C1479 t<6>.n334 VSS 2.03f
C1480 t<6>.n335 VSS 2.03f
C1481 t<6>.n336 VSS 8.3f
C1482 t<6>.n337 VSS -1.1f
C1483 t<6>.n338 VSS -0.69f
C1484 t<6>.n339 VSS -1.31f
C1485 t<6>.n340 VSS -0.965f
C1486 t<6>.n341 VSS -1.97f
C1487 t<6>.n342 VSS 7.43f
C1488 t<6>.n343 VSS -1.97f
C1489 t<6>.n344 VSS 2.03f
C1490 t<6>.n345 VSS 2.03f
C1491 t<6>.n346 VSS -1.1f
C1492 t<6>.n347 VSS -0.69f
C1493 t<6>.n348 VSS -1.1f
C1494 t<6>.n349 VSS 2.03f
C1495 t<6>.n350 VSS 7.43f
C1496 t<6>.n351 VSS -1.97f
C1497 t<6>.n352 VSS 7.43f
C1498 t<6>.n353 VSS 2.03f
C1499 t<6>.n354 VSS 2.03f
C1500 t<6>.n355 VSS 8.3f
C1501 t<6>.n356 VSS -1.1f
C1502 t<6>.n357 VSS -0.69f
C1503 t<6>.n358 VSS -1.31f
C1504 t<6>.n359 VSS -0.965f
C1505 t<6>.n360 VSS -1.97f
C1506 t<6>.n361 VSS 7.43f
C1507 t<6>.n362 VSS -1.97f
C1508 t<6>.n363 VSS 2.03f
C1509 t<6>.n364 VSS 2.03f
C1510 t<6>.n365 VSS -1.1f
C1511 t<6>.n366 VSS -0.69f
C1512 t<6>.n367 VSS -1.1f
C1513 t<6>.n368 VSS 2.03f
C1514 t<6>.n369 VSS 7.43f
C1515 t<6>.n370 VSS -1.97f
C1516 t<6>.n371 VSS 7.43f
C1517 t<6>.n372 VSS 2.03f
C1518 t<6>.n373 VSS 2.03f
C1519 t<6>.n374 VSS 8.3f
C1520 t<6>.n375 VSS -1.1f
C1521 t<6>.n376 VSS -0.69f
C1522 t<6>.n377 VSS -1.31f
C1523 t<6>.n378 VSS -0.965f
C1524 t<6>.n379 VSS -1.97f
C1525 t<6>.n380 VSS 7.43f
C1526 t<6>.n381 VSS -1.97f
C1527 t<6>.n382 VSS 2.03f
C1528 t<6>.n383 VSS 2.03f
C1529 t<6>.n384 VSS -1.1f
C1530 t<6>.n385 VSS -0.69f
C1531 t<6>.n386 VSS -1.1f
C1532 t<6>.n387 VSS 2.03f
C1533 t<6>.n388 VSS 7.43f
C1534 t<6>.n389 VSS -1.97f
C1535 t<6>.n390 VSS 7.43f
C1536 t<6>.n391 VSS 2.03f
C1537 t<6>.n392 VSS 2.03f
C1538 t<6>.n393 VSS 8.45f
C1539 t<6>.n394 VSS -0.552f
C1540 t<6>.n395 VSS -0.56f
C1541 t<6>.n396 VSS -0.791f
C1542 t<6>.n397 VSS -0.479f
C1543 t<6>.n398 VSS -0.552f
C1544 t<6>.n399 VSS 8.06f
C1545 t<6>.n400 VSS -1.58f
C1546 t<6>.n401 VSS -2.39f
C1547 t<6>.n402 VSS -29.4f
C1548 t<6>.n403 VSS -45.9f
C1549 t<6>.n404 VSS 2.38f
C1550 t<6>.n405 VSS 4.54f
C1551 t<6>.n406 VSS -1.31f
C1552 t<6>.n407 VSS -2.03f
C1553 t<6>.n408 VSS -1.11f
C1554 t<6>.n409 VSS -0.538f
C1555 t<6>.n410 VSS -0.56f
C1556 t<6>.n411 VSS -0.791f
C1557 t<6>.n412 VSS 11.6f
C1558 t<6>.n413 VSS 8.3f
C1559 t<6>.n414 VSS 2.03f
C1560 t<6>.n415 VSS -1.97f
C1561 t<6>.n416 VSS 7.43f
C1562 t<6>.n417 VSS 2.03f
C1563 t<6>.n418 VSS -1.1f
C1564 t<6>.n419 VSS 8.3f
C1565 t<6>.n420 VSS 2.03f
C1566 t<6>.n421 VSS -1.97f
C1567 t<6>.n422 VSS 7.43f
C1568 t<6>.n423 VSS 2.03f
C1569 t<6>.n424 VSS -1.1f
C1570 t<6>.n425 VSS 8.3f
C1571 t<6>.n426 VSS 2.03f
C1572 t<6>.n427 VSS -1.97f
C1573 t<6>.n428 VSS 7.43f
C1574 t<6>.n429 VSS 2.03f
C1575 t<6>.n430 VSS -1.1f
C1576 t<6>.n431 VSS 8.3f
C1577 t<6>.n432 VSS 2.03f
C1578 t<6>.n433 VSS -1.97f
C1579 t<6>.n434 VSS 7.43f
C1580 t<6>.n435 VSS 2.03f
C1581 t<6>.n436 VSS -1.1f
C1582 t<6>.n437 VSS 8.3f
C1583 t<6>.n438 VSS 2.03f
C1584 t<6>.n439 VSS -1.97f
C1585 t<6>.n440 VSS 7.43f
C1586 t<6>.n441 VSS 2.03f
C1587 t<6>.n442 VSS -1.1f
C1588 t<6>.n443 VSS 8.3f
C1589 t<6>.n444 VSS 2.03f
C1590 t<6>.n445 VSS -1.97f
C1591 t<6>.n446 VSS 7.43f
C1592 t<6>.n447 VSS 2.03f
C1593 t<6>.n448 VSS -1.1f
C1594 t<6>.n449 VSS 8.3f
C1595 t<6>.n450 VSS 2.03f
C1596 t<6>.n451 VSS -1.97f
C1597 t<6>.n452 VSS 7.43f
C1598 t<6>.n453 VSS 2.03f
C1599 t<6>.n454 VSS -1.1f
C1600 t<6>.n455 VSS 8.3f
C1601 t<6>.n456 VSS 2.03f
C1602 t<6>.n457 VSS -1.97f
C1603 t<6>.n458 VSS 7.43f
C1604 t<6>.n459 VSS 2.03f
C1605 t<6>.n460 VSS -1.1f
C1606 t<6>.n461 VSS 8.3f
C1607 t<6>.n462 VSS 2.03f
C1608 t<6>.n463 VSS -1.97f
C1609 t<6>.n464 VSS 7.43f
C1610 t<6>.n465 VSS 2.03f
C1611 t<6>.n466 VSS -1.1f
C1612 t<6>.n467 VSS 8.3f
C1613 t<6>.n468 VSS 2.03f
C1614 t<6>.n469 VSS -1.97f
C1615 t<6>.n470 VSS 7.43f
C1616 t<6>.n471 VSS 2.03f
C1617 t<6>.n472 VSS -1.1f
C1618 t<6>.n473 VSS 8.3f
C1619 t<6>.n474 VSS 2.03f
C1620 t<6>.n475 VSS -1.97f
C1621 t<6>.n476 VSS 7.43f
C1622 t<6>.n477 VSS 2.03f
C1623 t<6>.n478 VSS -1.1f
C1624 t<6>.n479 VSS 8.3f
C1625 t<6>.n480 VSS 2.03f
C1626 t<6>.n481 VSS -1.97f
C1627 t<6>.n482 VSS 7.43f
C1628 t<6>.n483 VSS 2.03f
C1629 t<6>.n484 VSS -1.1f
C1630 t<6>.n485 VSS 8.3f
C1631 t<6>.n486 VSS 2.03f
C1632 t<6>.n487 VSS -1.97f
C1633 t<6>.n488 VSS 7.43f
C1634 t<6>.n489 VSS 2.03f
C1635 t<6>.n490 VSS -1.1f
C1636 t<6>.n491 VSS 8.3f
C1637 t<6>.n492 VSS 2.03f
C1638 t<6>.n493 VSS -1.97f
C1639 t<6>.n494 VSS 7.43f
C1640 t<6>.n495 VSS 2.03f
C1641 t<6>.n496 VSS -1.1f
C1642 t<6>.n497 VSS 8.3f
C1643 t<6>.n498 VSS 2.03f
C1644 t<6>.n499 VSS -1.97f
C1645 t<6>.n500 VSS 7.43f
C1646 t<6>.n501 VSS 2.03f
C1647 t<6>.n502 VSS -1.1f
C1648 t<6>.n503 VSS 8.3f
C1649 t<6>.n504 VSS 2.03f
C1650 t<6>.n505 VSS -1.97f
C1651 t<6>.n506 VSS 7.43f
C1652 t<6>.n507 VSS 2.03f
C1653 t<6>.n508 VSS -1.1f
C1654 t<6>.n509 VSS 8.3f
C1655 t<6>.n510 VSS 2.03f
C1656 t<6>.n511 VSS -1.97f
C1657 t<6>.n512 VSS 7.43f
C1658 t<6>.n513 VSS 2.03f
C1659 t<6>.n514 VSS -1.1f
C1660 t<6>.n515 VSS 8.3f
C1661 t<6>.n516 VSS 2.03f
C1662 t<6>.n517 VSS -1.97f
C1663 t<6>.n518 VSS 7.43f
C1664 t<6>.n519 VSS 2.03f
C1665 t<6>.n520 VSS -1.1f
C1666 t<6>.n521 VSS 8.3f
C1667 t<6>.n522 VSS 2.03f
C1668 t<6>.n523 VSS -1.97f
C1669 t<6>.n524 VSS 7.43f
C1670 t<6>.n525 VSS 2.03f
C1671 t<6>.n526 VSS -1.1f
C1672 t<6>.n527 VSS 8.3f
C1673 t<6>.n528 VSS 2.03f
C1674 t<6>.n529 VSS -1.97f
C1675 t<6>.n530 VSS 7.43f
C1676 t<6>.n531 VSS 2.03f
C1677 t<6>.n532 VSS -1.1f
C1678 t<6>.n533 VSS 8.3f
C1679 t<6>.n534 VSS 2.03f
C1680 t<6>.n535 VSS -1.97f
C1681 t<6>.n536 VSS 7.43f
C1682 t<6>.n537 VSS 2.03f
C1683 t<6>.n538 VSS -1.1f
C1684 t<6>.n539 VSS 8.3f
C1685 t<6>.n540 VSS 2.03f
C1686 t<6>.n541 VSS -1.97f
C1687 t<6>.n542 VSS 7.43f
C1688 t<6>.n543 VSS 2.03f
C1689 t<6>.n544 VSS -1.1f
C1690 t<6>.n545 VSS 8.3f
C1691 t<6>.n546 VSS 2.03f
C1692 t<6>.n547 VSS -1.97f
C1693 t<6>.n548 VSS 7.43f
C1694 t<6>.n549 VSS 2.03f
C1695 t<6>.n550 VSS -1.1f
C1696 t<6>.n551 VSS 8.3f
C1697 t<6>.n552 VSS 2.03f
C1698 t<6>.n553 VSS -1.97f
C1699 t<6>.n554 VSS 7.43f
C1700 t<6>.n555 VSS 2.03f
C1701 t<6>.n556 VSS -1.1f
C1702 t<6>.n557 VSS 8.3f
C1703 t<6>.n558 VSS 2.03f
C1704 t<6>.n559 VSS -1.97f
C1705 t<6>.n560 VSS 7.43f
C1706 t<6>.n561 VSS 2.03f
C1707 t<6>.n562 VSS -1.1f
C1708 t<6>.n563 VSS 8.3f
C1709 t<6>.n564 VSS 2.03f
C1710 t<6>.n565 VSS -1.97f
C1711 t<6>.n566 VSS 7.43f
C1712 t<6>.n567 VSS 2.03f
C1713 t<6>.n568 VSS -1.1f
C1714 t<6>.n569 VSS 8.3f
C1715 t<6>.n570 VSS 2.03f
C1716 t<6>.n571 VSS -1.97f
C1717 t<6>.n572 VSS 7.43f
C1718 t<6>.n573 VSS 2.03f
C1719 t<6>.n574 VSS -1.1f
C1720 t<6>.n575 VSS 8.3f
C1721 t<6>.n576 VSS 2.03f
C1722 t<6>.n577 VSS -1.97f
C1723 t<6>.n578 VSS 7.43f
C1724 t<6>.n579 VSS 2.03f
C1725 t<6>.n580 VSS -1.1f
C1726 t<6>.n581 VSS 8.3f
C1727 t<6>.n582 VSS 2.03f
C1728 t<6>.n583 VSS -1.97f
C1729 t<6>.n584 VSS 7.43f
C1730 t<6>.n585 VSS 2.03f
C1731 t<6>.n586 VSS -1.1f
C1732 t<6>.n587 VSS 8.3f
C1733 t<6>.n588 VSS 2.03f
C1734 t<6>.n589 VSS -1.97f
C1735 t<6>.n590 VSS 7.43f
C1736 t<6>.n591 VSS 2.03f
C1737 t<6>.n592 VSS -0.952f
C1738 t<6>.n593 VSS -0.552f
C1739 t<6>.n594 VSS -0.221f
C1740 t<6>.n595 VSS 10.2f
C1741 t<6>.n596 VSS -1.67f
C1742 t<6>.n597 VSS -0.512f
C1743 t<6>.n598 VSS -4.64f
C1744 t<6>.n599 VSS -3.96f
C1745 tb<6>.n0 VSS 13.7f
C1746 tb<6>.n1 VSS 0.705f
C1747 tb<6>.n2 VSS -0.946f
C1748 tb<6>.n3 VSS -1.93f
C1749 tb<6>.n4 VSS 7.28f
C1750 tb<6>.n5 VSS 1.99f
C1751 tb<6>.n6 VSS -1.08f
C1752 tb<6>.n7 VSS -0.676f
C1753 tb<6>.n8 VSS -1.28f
C1754 tb<6>.n9 VSS -0.946f
C1755 tb<6>.n10 VSS -1.93f
C1756 tb<6>.n11 VSS 7.28f
C1757 tb<6>.n12 VSS 1.99f
C1758 tb<6>.n13 VSS -1.08f
C1759 tb<6>.n14 VSS -0.676f
C1760 tb<6>.n15 VSS -1.28f
C1761 tb<6>.n16 VSS -0.946f
C1762 tb<6>.n17 VSS -1.93f
C1763 tb<6>.n18 VSS 7.28f
C1764 tb<6>.n19 VSS 1.99f
C1765 tb<6>.n20 VSS -1.08f
C1766 tb<6>.n21 VSS -0.676f
C1767 tb<6>.n22 VSS -1.28f
C1768 tb<6>.n23 VSS -0.946f
C1769 tb<6>.n24 VSS -1.93f
C1770 tb<6>.n25 VSS 7.28f
C1771 tb<6>.n26 VSS 1.99f
C1772 tb<6>.n27 VSS -1.08f
C1773 tb<6>.n28 VSS -0.676f
C1774 tb<6>.n29 VSS -1.28f
C1775 tb<6>.n30 VSS -0.946f
C1776 tb<6>.n31 VSS -1.93f
C1777 tb<6>.n32 VSS 7.28f
C1778 tb<6>.n33 VSS 1.99f
C1779 tb<6>.n34 VSS -1.08f
C1780 tb<6>.n35 VSS -0.676f
C1781 tb<6>.n36 VSS -1.28f
C1782 tb<6>.n37 VSS -0.946f
C1783 tb<6>.n38 VSS -1.93f
C1784 tb<6>.n39 VSS 7.28f
C1785 tb<6>.n40 VSS 1.99f
C1786 tb<6>.n41 VSS -1.08f
C1787 tb<6>.n42 VSS -0.676f
C1788 tb<6>.n43 VSS -1.28f
C1789 tb<6>.n44 VSS -0.946f
C1790 tb<6>.n45 VSS -1.93f
C1791 tb<6>.n46 VSS 7.28f
C1792 tb<6>.n47 VSS 1.99f
C1793 tb<6>.n48 VSS -1.08f
C1794 tb<6>.n49 VSS -0.676f
C1795 tb<6>.n50 VSS -1.28f
C1796 tb<6>.n51 VSS -0.946f
C1797 tb<6>.n52 VSS -1.93f
C1798 tb<6>.n53 VSS 7.28f
C1799 tb<6>.n54 VSS 1.99f
C1800 tb<6>.n55 VSS -1.08f
C1801 tb<6>.n56 VSS -0.676f
C1802 tb<6>.n57 VSS -1.28f
C1803 tb<6>.n58 VSS -0.946f
C1804 tb<6>.n59 VSS -1.93f
C1805 tb<6>.n60 VSS 7.28f
C1806 tb<6>.n61 VSS 1.99f
C1807 tb<6>.n62 VSS -1.08f
C1808 tb<6>.n63 VSS -0.676f
C1809 tb<6>.n64 VSS -1.28f
C1810 tb<6>.n65 VSS -0.946f
C1811 tb<6>.n66 VSS -1.93f
C1812 tb<6>.n67 VSS 7.28f
C1813 tb<6>.n68 VSS 1.99f
C1814 tb<6>.n69 VSS -1.08f
C1815 tb<6>.n70 VSS -0.676f
C1816 tb<6>.n71 VSS -1.28f
C1817 tb<6>.n72 VSS -0.946f
C1818 tb<6>.n73 VSS -1.93f
C1819 tb<6>.n74 VSS 7.28f
C1820 tb<6>.n75 VSS 1.99f
C1821 tb<6>.n76 VSS -1.08f
C1822 tb<6>.n77 VSS -0.676f
C1823 tb<6>.n78 VSS -1.28f
C1824 tb<6>.n79 VSS -0.946f
C1825 tb<6>.n80 VSS -1.93f
C1826 tb<6>.n81 VSS 7.28f
C1827 tb<6>.n82 VSS 1.99f
C1828 tb<6>.n83 VSS -1.08f
C1829 tb<6>.n84 VSS -0.676f
C1830 tb<6>.n85 VSS -1.28f
C1831 tb<6>.n86 VSS -0.946f
C1832 tb<6>.n87 VSS -1.93f
C1833 tb<6>.n88 VSS 7.28f
C1834 tb<6>.n89 VSS 1.99f
C1835 tb<6>.n90 VSS -1.08f
C1836 tb<6>.n91 VSS -0.676f
C1837 tb<6>.n92 VSS -1.28f
C1838 tb<6>.n93 VSS -0.946f
C1839 tb<6>.n94 VSS -1.93f
C1840 tb<6>.n95 VSS 7.28f
C1841 tb<6>.n96 VSS 1.99f
C1842 tb<6>.n97 VSS -1.08f
C1843 tb<6>.n98 VSS -0.676f
C1844 tb<6>.n99 VSS -1.28f
C1845 tb<6>.n100 VSS -0.946f
C1846 tb<6>.n101 VSS -1.93f
C1847 tb<6>.n102 VSS 7.28f
C1848 tb<6>.n103 VSS 1.99f
C1849 tb<6>.n104 VSS -1.08f
C1850 tb<6>.n105 VSS -0.676f
C1851 tb<6>.n106 VSS -1.28f
C1852 tb<6>.n107 VSS -0.946f
C1853 tb<6>.n108 VSS -1.93f
C1854 tb<6>.n109 VSS 7.28f
C1855 tb<6>.n110 VSS 1.99f
C1856 tb<6>.n111 VSS -1.08f
C1857 tb<6>.n112 VSS -0.676f
C1858 tb<6>.n113 VSS -1.28f
C1859 tb<6>.n114 VSS -0.946f
C1860 tb<6>.n115 VSS -1.93f
C1861 tb<6>.n116 VSS 7.28f
C1862 tb<6>.n117 VSS 1.99f
C1863 tb<6>.n118 VSS -1.08f
C1864 tb<6>.n119 VSS -0.676f
C1865 tb<6>.n120 VSS -1.28f
C1866 tb<6>.n121 VSS -0.946f
C1867 tb<6>.n122 VSS -1.93f
C1868 tb<6>.n123 VSS 7.28f
C1869 tb<6>.n124 VSS 1.99f
C1870 tb<6>.n125 VSS -1.08f
C1871 tb<6>.n126 VSS -0.676f
C1872 tb<6>.n127 VSS -1.28f
C1873 tb<6>.n128 VSS -0.946f
C1874 tb<6>.n129 VSS -1.93f
C1875 tb<6>.n130 VSS 7.28f
C1876 tb<6>.n131 VSS 1.99f
C1877 tb<6>.n132 VSS -1.08f
C1878 tb<6>.n133 VSS -0.676f
C1879 tb<6>.n134 VSS -1.28f
C1880 tb<6>.n135 VSS -0.946f
C1881 tb<6>.n136 VSS -1.93f
C1882 tb<6>.n137 VSS 7.28f
C1883 tb<6>.n138 VSS 1.99f
C1884 tb<6>.n139 VSS -1.08f
C1885 tb<6>.n140 VSS -0.676f
C1886 tb<6>.n141 VSS -1.28f
C1887 tb<6>.n142 VSS -0.946f
C1888 tb<6>.n143 VSS -1.93f
C1889 tb<6>.n144 VSS 7.28f
C1890 tb<6>.n145 VSS 1.99f
C1891 tb<6>.n146 VSS -1.08f
C1892 tb<6>.n147 VSS -0.676f
C1893 tb<6>.n148 VSS -1.28f
C1894 tb<6>.n149 VSS -0.946f
C1895 tb<6>.n150 VSS -1.93f
C1896 tb<6>.n151 VSS 7.28f
C1897 tb<6>.n152 VSS 1.99f
C1898 tb<6>.n153 VSS -1.08f
C1899 tb<6>.n154 VSS -0.676f
C1900 tb<6>.n155 VSS -1.28f
C1901 tb<6>.n156 VSS -0.946f
C1902 tb<6>.n157 VSS -1.93f
C1903 tb<6>.n158 VSS 7.28f
C1904 tb<6>.n159 VSS 1.99f
C1905 tb<6>.n160 VSS -1.08f
C1906 tb<6>.n161 VSS -0.676f
C1907 tb<6>.n162 VSS -1.28f
C1908 tb<6>.n163 VSS -0.946f
C1909 tb<6>.n164 VSS -1.93f
C1910 tb<6>.n165 VSS 7.28f
C1911 tb<6>.n166 VSS 1.99f
C1912 tb<6>.n167 VSS -1.08f
C1913 tb<6>.n168 VSS -0.676f
C1914 tb<6>.n169 VSS -1.28f
C1915 tb<6>.n170 VSS -0.946f
C1916 tb<6>.n171 VSS -1.93f
C1917 tb<6>.n172 VSS 7.28f
C1918 tb<6>.n173 VSS 1.99f
C1919 tb<6>.n174 VSS -1.08f
C1920 tb<6>.n175 VSS -0.676f
C1921 tb<6>.n176 VSS -1.28f
C1922 tb<6>.n177 VSS -0.946f
C1923 tb<6>.n178 VSS -1.93f
C1924 tb<6>.n179 VSS 7.28f
C1925 tb<6>.n180 VSS 1.99f
C1926 tb<6>.n181 VSS -1.08f
C1927 tb<6>.n182 VSS -0.676f
C1928 tb<6>.n183 VSS -1.28f
C1929 tb<6>.n184 VSS -0.946f
C1930 tb<6>.n185 VSS -1.93f
C1931 tb<6>.n186 VSS 7.28f
C1932 tb<6>.n187 VSS 1.99f
C1933 tb<6>.n188 VSS -1.08f
C1934 tb<6>.n189 VSS -0.676f
C1935 tb<6>.n190 VSS -1.28f
C1936 tb<6>.n191 VSS -0.946f
C1937 tb<6>.n192 VSS -1.93f
C1938 tb<6>.n193 VSS 7.28f
C1939 tb<6>.n194 VSS 1.99f
C1940 tb<6>.n195 VSS -1.08f
C1941 tb<6>.n196 VSS -0.676f
C1942 tb<6>.n197 VSS -1.28f
C1943 tb<6>.n198 VSS -0.946f
C1944 tb<6>.n199 VSS -1.93f
C1945 tb<6>.n200 VSS 7.28f
C1946 tb<6>.n201 VSS 1.99f
C1947 tb<6>.n202 VSS -1.08f
C1948 tb<6>.n203 VSS -0.676f
C1949 tb<6>.n204 VSS -1.28f
C1950 tb<6>.n205 VSS -0.946f
C1951 tb<6>.n206 VSS -1.93f
C1952 tb<6>.n207 VSS 7.28f
C1953 tb<6>.n208 VSS 1.99f
C1954 tb<6>.n209 VSS -0.932f
C1955 tb<6>.n210 VSS -0.549f
C1956 tb<6>.n211 VSS -0.775f
C1957 tb<6>.n212 VSS -0.469f
C1958 tb<6>.n213 VSS -2.18f
C1959 tb<6>.n214 VSS -0.665f
C1960 tb<6>.n215 VSS 12.2f
C1961 tb<6>.n216 VSS 7.28f
C1962 tb<6>.n217 VSS -1.93f
C1963 tb<6>.n218 VSS 1.99f
C1964 tb<6>.n219 VSS 8.13f
C1965 tb<6>.n220 VSS -1.08f
C1966 tb<6>.n221 VSS 1.99f
C1967 tb<6>.n222 VSS 7.28f
C1968 tb<6>.n223 VSS -1.93f
C1969 tb<6>.n224 VSS 1.99f
C1970 tb<6>.n225 VSS 8.13f
C1971 tb<6>.n226 VSS -1.08f
C1972 tb<6>.n227 VSS 1.99f
C1973 tb<6>.n228 VSS 7.28f
C1974 tb<6>.n229 VSS -1.93f
C1975 tb<6>.n230 VSS 1.99f
C1976 tb<6>.n231 VSS 8.13f
C1977 tb<6>.n232 VSS -1.08f
C1978 tb<6>.n233 VSS 1.99f
C1979 tb<6>.n234 VSS 7.28f
C1980 tb<6>.n235 VSS -1.93f
C1981 tb<6>.n236 VSS 1.99f
C1982 tb<6>.n237 VSS 8.13f
C1983 tb<6>.n238 VSS -1.08f
C1984 tb<6>.n239 VSS 1.99f
C1985 tb<6>.n240 VSS 7.28f
C1986 tb<6>.n241 VSS -1.93f
C1987 tb<6>.n242 VSS 1.99f
C1988 tb<6>.n243 VSS 8.13f
C1989 tb<6>.n244 VSS -1.08f
C1990 tb<6>.n245 VSS 1.99f
C1991 tb<6>.n246 VSS 7.28f
C1992 tb<6>.n247 VSS -1.93f
C1993 tb<6>.n248 VSS 1.99f
C1994 tb<6>.n249 VSS 8.13f
C1995 tb<6>.n250 VSS -1.08f
C1996 tb<6>.n251 VSS 1.99f
C1997 tb<6>.n252 VSS 7.28f
C1998 tb<6>.n253 VSS -1.93f
C1999 tb<6>.n254 VSS 1.99f
C2000 tb<6>.n255 VSS 8.13f
C2001 tb<6>.n256 VSS -1.08f
C2002 tb<6>.n257 VSS 1.99f
C2003 tb<6>.n258 VSS 7.28f
C2004 tb<6>.n259 VSS -1.93f
C2005 tb<6>.n260 VSS 1.99f
C2006 tb<6>.n261 VSS 8.13f
C2007 tb<6>.n262 VSS -1.08f
C2008 tb<6>.n263 VSS 1.99f
C2009 tb<6>.n264 VSS 7.28f
C2010 tb<6>.n265 VSS -1.93f
C2011 tb<6>.n266 VSS 1.99f
C2012 tb<6>.n267 VSS 8.13f
C2013 tb<6>.n268 VSS -1.08f
C2014 tb<6>.n269 VSS 1.99f
C2015 tb<6>.n270 VSS 7.28f
C2016 tb<6>.n271 VSS -1.93f
C2017 tb<6>.n272 VSS 1.99f
C2018 tb<6>.n273 VSS 8.13f
C2019 tb<6>.n274 VSS -1.08f
C2020 tb<6>.n275 VSS 1.99f
C2021 tb<6>.n276 VSS 7.28f
C2022 tb<6>.n277 VSS -1.93f
C2023 tb<6>.n278 VSS 1.99f
C2024 tb<6>.n279 VSS 8.13f
C2025 tb<6>.n280 VSS -1.08f
C2026 tb<6>.n281 VSS 1.99f
C2027 tb<6>.n282 VSS 7.28f
C2028 tb<6>.n283 VSS -1.93f
C2029 tb<6>.n284 VSS 1.99f
C2030 tb<6>.n285 VSS 8.13f
C2031 tb<6>.n286 VSS -1.08f
C2032 tb<6>.n287 VSS 1.99f
C2033 tb<6>.n288 VSS 7.28f
C2034 tb<6>.n289 VSS -1.93f
C2035 tb<6>.n290 VSS 1.99f
C2036 tb<6>.n291 VSS 8.13f
C2037 tb<6>.n292 VSS -1.08f
C2038 tb<6>.n293 VSS 1.99f
C2039 tb<6>.n294 VSS 7.28f
C2040 tb<6>.n295 VSS -1.93f
C2041 tb<6>.n296 VSS 1.99f
C2042 tb<6>.n297 VSS 8.13f
C2043 tb<6>.n298 VSS -1.08f
C2044 tb<6>.n299 VSS 1.99f
C2045 tb<6>.n300 VSS 7.28f
C2046 tb<6>.n301 VSS -1.93f
C2047 tb<6>.n302 VSS 1.99f
C2048 tb<6>.n303 VSS 8.13f
C2049 tb<6>.n304 VSS -1.08f
C2050 tb<6>.n305 VSS 1.99f
C2051 tb<6>.n306 VSS 7.28f
C2052 tb<6>.n307 VSS -1.93f
C2053 tb<6>.n308 VSS 1.99f
C2054 tb<6>.n309 VSS 8.13f
C2055 tb<6>.n310 VSS -1.08f
C2056 tb<6>.n311 VSS 1.99f
C2057 tb<6>.n312 VSS 7.28f
C2058 tb<6>.n313 VSS -1.93f
C2059 tb<6>.n314 VSS 1.99f
C2060 tb<6>.n315 VSS 8.13f
C2061 tb<6>.n316 VSS -1.08f
C2062 tb<6>.n317 VSS 1.99f
C2063 tb<6>.n318 VSS 7.28f
C2064 tb<6>.n319 VSS -1.93f
C2065 tb<6>.n320 VSS 1.99f
C2066 tb<6>.n321 VSS 8.13f
C2067 tb<6>.n322 VSS -1.08f
C2068 tb<6>.n323 VSS 1.99f
C2069 tb<6>.n324 VSS 7.28f
C2070 tb<6>.n325 VSS -1.93f
C2071 tb<6>.n326 VSS 1.99f
C2072 tb<6>.n327 VSS 8.13f
C2073 tb<6>.n328 VSS -1.08f
C2074 tb<6>.n329 VSS 1.99f
C2075 tb<6>.n330 VSS 7.28f
C2076 tb<6>.n331 VSS -1.93f
C2077 tb<6>.n332 VSS 1.99f
C2078 tb<6>.n333 VSS 8.13f
C2079 tb<6>.n334 VSS -1.08f
C2080 tb<6>.n335 VSS 1.99f
C2081 tb<6>.n336 VSS 7.28f
C2082 tb<6>.n337 VSS -1.93f
C2083 tb<6>.n338 VSS 1.99f
C2084 tb<6>.n339 VSS 8.13f
C2085 tb<6>.n340 VSS -1.08f
C2086 tb<6>.n341 VSS 1.99f
C2087 tb<6>.n342 VSS 7.28f
C2088 tb<6>.n343 VSS -1.93f
C2089 tb<6>.n344 VSS 1.99f
C2090 tb<6>.n345 VSS 8.13f
C2091 tb<6>.n346 VSS -1.08f
C2092 tb<6>.n347 VSS 1.99f
C2093 tb<6>.n348 VSS 7.28f
C2094 tb<6>.n349 VSS -1.93f
C2095 tb<6>.n350 VSS 1.99f
C2096 tb<6>.n351 VSS 8.13f
C2097 tb<6>.n352 VSS -1.08f
C2098 tb<6>.n353 VSS 1.99f
C2099 tb<6>.n354 VSS 7.28f
C2100 tb<6>.n355 VSS -1.93f
C2101 tb<6>.n356 VSS 1.99f
C2102 tb<6>.n357 VSS 8.13f
C2103 tb<6>.n358 VSS -1.08f
C2104 tb<6>.n359 VSS 1.99f
C2105 tb<6>.n360 VSS 7.28f
C2106 tb<6>.n361 VSS -1.93f
C2107 tb<6>.n362 VSS 1.99f
C2108 tb<6>.n363 VSS 8.13f
C2109 tb<6>.n364 VSS -1.08f
C2110 tb<6>.n365 VSS 1.99f
C2111 tb<6>.n366 VSS 7.28f
C2112 tb<6>.n367 VSS -1.93f
C2113 tb<6>.n368 VSS 1.99f
C2114 tb<6>.n369 VSS 8.13f
C2115 tb<6>.n370 VSS -1.08f
C2116 tb<6>.n371 VSS 1.99f
C2117 tb<6>.n372 VSS 7.28f
C2118 tb<6>.n373 VSS -1.93f
C2119 tb<6>.n374 VSS 1.99f
C2120 tb<6>.n375 VSS 8.13f
C2121 tb<6>.n376 VSS -1.08f
C2122 tb<6>.n377 VSS 1.99f
C2123 tb<6>.n378 VSS 7.28f
C2124 tb<6>.n379 VSS -1.93f
C2125 tb<6>.n380 VSS 1.99f
C2126 tb<6>.n381 VSS 8.13f
C2127 tb<6>.n382 VSS -1.08f
C2128 tb<6>.n383 VSS 1.99f
C2129 tb<6>.n384 VSS 7.28f
C2130 tb<6>.n385 VSS -1.93f
C2131 tb<6>.n386 VSS 1.99f
C2132 tb<6>.n387 VSS 8.13f
C2133 tb<6>.n388 VSS -1.08f
C2134 tb<6>.n389 VSS 1.99f
C2135 tb<6>.n390 VSS 7.28f
C2136 tb<6>.n391 VSS -1.93f
C2137 tb<6>.n392 VSS 1.99f
C2138 tb<6>.n393 VSS 8.28f
C2139 tb<6>.n394 VSS -0.541f
C2140 tb<6>.n395 VSS -0.216f
C2141 tb<6>.n396 VSS -0.541f
C2142 tb<6>.n397 VSS 7.9f
C2143 tb<6>.n398 VSS -1.55f
C2144 tb<6>.n399 VSS -2.34f
C2145 tb<6>.n400 VSS -2.37f
C2146 tb<6>.n401 VSS -15.8f
C2147 tb<6>.n402 VSS -72.7f
C2148 tb<6>.n403 VSS -72.7f
C2149 tb<6>.n404 VSS 2.34f
C2150 tb<6>.n405 VSS 4.44f
C2151 tb<6>.n406 VSS -1.28f
C2152 tb<6>.n407 VSS -1.99f
C2153 tb<6>.n408 VSS -0.946f
C2154 tb<6>.n409 VSS -1.09f
C2155 tb<6>.n410 VSS -0.527f
C2156 tb<6>.n411 VSS -0.549f
C2157 tb<6>.n412 VSS -0.775f
C2158 tb<6>.n413 VSS 11.4f
C2159 tb<6>.n414 VSS 8.13f
C2160 tb<6>.n415 VSS 1.99f
C2161 tb<6>.n416 VSS -1.93f
C2162 tb<6>.n417 VSS 7.28f
C2163 tb<6>.n418 VSS 1.99f
C2164 tb<6>.n419 VSS -1.08f
C2165 tb<6>.n420 VSS 8.13f
C2166 tb<6>.n421 VSS 1.99f
C2167 tb<6>.n422 VSS -1.93f
C2168 tb<6>.n423 VSS 7.28f
C2169 tb<6>.n424 VSS 1.99f
C2170 tb<6>.n425 VSS -1.08f
C2171 tb<6>.n426 VSS 8.13f
C2172 tb<6>.n427 VSS 1.99f
C2173 tb<6>.n428 VSS -1.93f
C2174 tb<6>.n429 VSS 7.28f
C2175 tb<6>.n430 VSS 1.99f
C2176 tb<6>.n431 VSS -1.08f
C2177 tb<6>.n432 VSS 8.13f
C2178 tb<6>.n433 VSS 1.99f
C2179 tb<6>.n434 VSS -1.93f
C2180 tb<6>.n435 VSS 7.28f
C2181 tb<6>.n436 VSS 1.99f
C2182 tb<6>.n437 VSS -1.08f
C2183 tb<6>.n438 VSS 8.13f
C2184 tb<6>.n439 VSS 1.99f
C2185 tb<6>.n440 VSS -1.93f
C2186 tb<6>.n441 VSS 7.28f
C2187 tb<6>.n442 VSS 1.99f
C2188 tb<6>.n443 VSS -1.08f
C2189 tb<6>.n444 VSS 8.13f
C2190 tb<6>.n445 VSS 1.99f
C2191 tb<6>.n446 VSS -1.93f
C2192 tb<6>.n447 VSS 7.28f
C2193 tb<6>.n448 VSS 1.99f
C2194 tb<6>.n449 VSS -1.08f
C2195 tb<6>.n450 VSS 8.13f
C2196 tb<6>.n451 VSS 1.99f
C2197 tb<6>.n452 VSS -1.93f
C2198 tb<6>.n453 VSS 7.28f
C2199 tb<6>.n454 VSS 1.99f
C2200 tb<6>.n455 VSS -1.08f
C2201 tb<6>.n456 VSS 8.13f
C2202 tb<6>.n457 VSS 1.99f
C2203 tb<6>.n458 VSS -1.93f
C2204 tb<6>.n459 VSS 7.28f
C2205 tb<6>.n460 VSS 1.99f
C2206 tb<6>.n461 VSS -1.08f
C2207 tb<6>.n462 VSS 8.13f
C2208 tb<6>.n463 VSS 1.99f
C2209 tb<6>.n464 VSS -1.93f
C2210 tb<6>.n465 VSS 7.28f
C2211 tb<6>.n466 VSS 1.99f
C2212 tb<6>.n467 VSS -1.08f
C2213 tb<6>.n468 VSS 8.13f
C2214 tb<6>.n469 VSS 1.99f
C2215 tb<6>.n470 VSS -1.93f
C2216 tb<6>.n471 VSS 7.28f
C2217 tb<6>.n472 VSS 1.99f
C2218 tb<6>.n473 VSS -1.08f
C2219 tb<6>.n474 VSS 8.13f
C2220 tb<6>.n475 VSS 1.99f
C2221 tb<6>.n476 VSS -1.93f
C2222 tb<6>.n477 VSS 7.28f
C2223 tb<6>.n478 VSS 1.99f
C2224 tb<6>.n479 VSS -1.08f
C2225 tb<6>.n480 VSS 8.13f
C2226 tb<6>.n481 VSS 1.99f
C2227 tb<6>.n482 VSS -1.93f
C2228 tb<6>.n483 VSS 7.28f
C2229 tb<6>.n484 VSS 1.99f
C2230 tb<6>.n485 VSS -1.08f
C2231 tb<6>.n486 VSS 8.13f
C2232 tb<6>.n487 VSS 1.99f
C2233 tb<6>.n488 VSS -1.93f
C2234 tb<6>.n489 VSS 7.28f
C2235 tb<6>.n490 VSS 1.99f
C2236 tb<6>.n491 VSS -1.08f
C2237 tb<6>.n492 VSS 8.13f
C2238 tb<6>.n493 VSS 1.99f
C2239 tb<6>.n494 VSS -1.93f
C2240 tb<6>.n495 VSS 7.28f
C2241 tb<6>.n496 VSS 1.99f
C2242 tb<6>.n497 VSS -1.08f
C2243 tb<6>.n498 VSS 8.13f
C2244 tb<6>.n499 VSS 1.99f
C2245 tb<6>.n500 VSS -1.93f
C2246 tb<6>.n501 VSS 7.28f
C2247 tb<6>.n502 VSS 1.99f
C2248 tb<6>.n503 VSS -1.08f
C2249 tb<6>.n504 VSS 8.13f
C2250 tb<6>.n505 VSS 1.99f
C2251 tb<6>.n506 VSS -1.93f
C2252 tb<6>.n507 VSS 7.28f
C2253 tb<6>.n508 VSS 1.99f
C2254 tb<6>.n509 VSS -1.08f
C2255 tb<6>.n510 VSS 8.13f
C2256 tb<6>.n511 VSS 1.99f
C2257 tb<6>.n512 VSS -1.93f
C2258 tb<6>.n513 VSS 7.28f
C2259 tb<6>.n514 VSS 1.99f
C2260 tb<6>.n515 VSS -1.08f
C2261 tb<6>.n516 VSS 8.13f
C2262 tb<6>.n517 VSS 1.99f
C2263 tb<6>.n518 VSS -1.93f
C2264 tb<6>.n519 VSS 7.28f
C2265 tb<6>.n520 VSS 1.99f
C2266 tb<6>.n521 VSS -1.08f
C2267 tb<6>.n522 VSS 8.13f
C2268 tb<6>.n523 VSS 1.99f
C2269 tb<6>.n524 VSS -1.93f
C2270 tb<6>.n525 VSS 7.28f
C2271 tb<6>.n526 VSS 1.99f
C2272 tb<6>.n527 VSS -1.08f
C2273 tb<6>.n528 VSS 8.13f
C2274 tb<6>.n529 VSS 1.99f
C2275 tb<6>.n530 VSS -1.93f
C2276 tb<6>.n531 VSS 7.28f
C2277 tb<6>.n532 VSS 1.99f
C2278 tb<6>.n533 VSS -1.08f
C2279 tb<6>.n534 VSS 8.13f
C2280 tb<6>.n535 VSS 1.99f
C2281 tb<6>.n536 VSS -1.93f
C2282 tb<6>.n537 VSS 7.28f
C2283 tb<6>.n538 VSS 1.99f
C2284 tb<6>.n539 VSS -1.08f
C2285 tb<6>.n540 VSS 8.13f
C2286 tb<6>.n541 VSS 1.99f
C2287 tb<6>.n542 VSS -1.93f
C2288 tb<6>.n543 VSS 7.28f
C2289 tb<6>.n544 VSS 1.99f
C2290 tb<6>.n545 VSS -1.08f
C2291 tb<6>.n546 VSS 8.13f
C2292 tb<6>.n547 VSS 1.99f
C2293 tb<6>.n548 VSS -1.93f
C2294 tb<6>.n549 VSS 7.28f
C2295 tb<6>.n550 VSS 1.99f
C2296 tb<6>.n551 VSS -1.08f
C2297 tb<6>.n552 VSS 8.13f
C2298 tb<6>.n553 VSS 1.99f
C2299 tb<6>.n554 VSS -1.93f
C2300 tb<6>.n555 VSS 7.28f
C2301 tb<6>.n556 VSS 1.99f
C2302 tb<6>.n557 VSS -1.08f
C2303 tb<6>.n558 VSS 8.13f
C2304 tb<6>.n559 VSS 1.99f
C2305 tb<6>.n560 VSS -1.93f
C2306 tb<6>.n561 VSS 7.28f
C2307 tb<6>.n562 VSS 1.99f
C2308 tb<6>.n563 VSS -1.08f
C2309 tb<6>.n564 VSS 8.13f
C2310 tb<6>.n565 VSS 1.99f
C2311 tb<6>.n566 VSS -1.93f
C2312 tb<6>.n567 VSS 7.28f
C2313 tb<6>.n568 VSS 1.99f
C2314 tb<6>.n569 VSS -1.08f
C2315 tb<6>.n570 VSS 8.13f
C2316 tb<6>.n571 VSS 1.99f
C2317 tb<6>.n572 VSS -1.93f
C2318 tb<6>.n573 VSS 7.28f
C2319 tb<6>.n574 VSS 1.99f
C2320 tb<6>.n575 VSS -1.08f
C2321 tb<6>.n576 VSS 8.13f
C2322 tb<6>.n577 VSS 1.99f
C2323 tb<6>.n578 VSS -1.93f
C2324 tb<6>.n579 VSS 7.28f
C2325 tb<6>.n580 VSS 1.99f
C2326 tb<6>.n581 VSS -1.08f
C2327 tb<6>.n582 VSS 8.13f
C2328 tb<6>.n583 VSS 1.99f
C2329 tb<6>.n584 VSS -1.93f
C2330 tb<6>.n585 VSS 7.28f
C2331 tb<6>.n586 VSS 1.99f
C2332 tb<6>.n587 VSS -1.08f
C2333 tb<6>.n588 VSS 8.13f
C2334 tb<6>.n589 VSS 1.99f
C2335 tb<6>.n590 VSS -1.93f
C2336 tb<6>.n591 VSS 7.28f
C2337 tb<6>.n592 VSS 1.99f
C2338 tb<6>.n593 VSS -0.932f
C2339 tb<6>.n594 VSS -0.541f
C2340 tb<6>.n595 VSS -0.216f
C2341 tb<6>.n596 VSS 9.99f
C2342 tb<6>.n597 VSS -1.64f
C2343 tb<6>.n598 VSS -0.502f
C2344 tb<6>.n599 VSS -4.54f
C2345 tb<6>.n600 VSS -3.88f
C2346 t<2>.n0 VSS 2.12f
C2347 t<2>.n1 VSS -0.206f
C2348 t<2>.n2 VSS 0.295f
C2349 t<2>.n3 VSS -0.94f
C2350 t<2>.n4 VSS -0.737f
C2351 t<2>.n5 VSS -2.95f
C2352 t<2>.n6 VSS 0.28f
C2353 t<2>.n7 VSS 0.362f
C2354 t<2>.n8 VSS 4.11f
C2355 t<2>.n9 VSS 5.83f
C2356 t<2>.n10 VSS -1.08f
C2357 t<2>.n11 VSS 0.686f
C2358 t<2>.n12 VSS 0.287f
C2359 t<2>.n13 VSS -0.753f
C2360 t<2>.n14 VSS -3.03f
C2361 t<2>.n15 VSS -0.138f
C2362 t<2>.n16 VSS 0.605f
C2363 t<2>.n17 VSS 0.496f
C2364 t<4>.n0 VSS 20.5f
C2365 t<4>.n1 VSS 1.28f
C2366 t<4>.n2 VSS -12f
C2367 t<4>.n3 VSS 0.699f
C2368 t<4>.n4 VSS -2.57f
C2369 t<4>.n5 VSS -9.41f
C2370 t<4>.n6 VSS -10.5f
C2371 t<4>.n7 VSS 1.65f
C2372 t<4>.n8 VSS -9.41f
C2373 t<4>.n9 VSS -2.57f
C2374 t<4>.n10 VSS 1.4f
C2375 t<4>.n11 VSS 2.5f
C2376 t<4>.n12 VSS -2.57f
C2377 t<4>.n13 VSS 0.873f
C2378 t<4>.n14 VSS -9.41f
C2379 t<4>.n15 VSS -2.57f
C2380 t<4>.n16 VSS 1.4f
C2381 t<4>.n17 VSS 2.5f
C2382 t<4>.n18 VSS -2.57f
C2383 t<4>.n19 VSS 0.873f
C2384 t<4>.n20 VSS -9.41f
C2385 t<4>.n21 VSS -2.57f
C2386 t<4>.n22 VSS -14.7f
C2387 t<4>.n23 VSS -13.4f
C2388 t<4>.n24 VSS 1.57f
C2389 t<4>.n25 VSS 0.873f
C2390 t<4>.n26 VSS 1.4f
C2391 t<4>.n27 VSS -10.5f
C2392 t<4>.n28 VSS -2.57f
C2393 t<4>.n29 VSS 2.5f
C2394 t<4>.n30 VSS -9.41f
C2395 t<4>.n31 VSS 2.5f
C2396 t<4>.n32 VSS 1.65f
C2397 t<4>.n33 VSS 1.22f
C2398 t<4>.n34 VSS -2.57f
C2399 t<4>.n35 VSS 1.4f
C2400 t<4>.n36 VSS -10.5f
C2401 t<4>.n37 VSS 1.4f
C2402 t<4>.n38 VSS -2.57f
C2403 t<4>.n39 VSS -9.41f
C2404 t<4>.n40 VSS 2.5f
C2405 t<4>.n41 VSS -9.41f
C2406 t<4>.n42 VSS -2.57f
C2407 t<4>.n43 VSS 1.22f
C2408 t<4>.n44 VSS 1.65f
C2409 t<4>.n45 VSS 0.873f
C2410 t<4>.n46 VSS 1.4f
C2411 t<4>.n47 VSS -10.5f
C2412 t<4>.n48 VSS -2.57f
C2413 t<4>.n49 VSS 2.5f
C2414 t<4>.n50 VSS -9.41f
C2415 t<4>.n51 VSS 2.5f
C2416 t<4>.n52 VSS 1.65f
C2417 t<4>.n53 VSS 1.22f
C2418 t<4>.n54 VSS -2.57f
C2419 t<4>.n55 VSS 1.4f
C2420 t<4>.n56 VSS -10.5f
C2421 t<4>.n57 VSS 1.4f
C2422 t<4>.n58 VSS -2.57f
C2423 t<4>.n59 VSS -9.41f
C2424 t<4>.n60 VSS 2.5f
C2425 t<4>.n61 VSS -9.41f
C2426 t<4>.n62 VSS -2.57f
C2427 t<4>.n63 VSS 1.22f
C2428 t<4>.n64 VSS 1.65f
C2429 t<4>.n65 VSS 0.873f
C2430 t<4>.n66 VSS 1.4f
C2431 t<4>.n67 VSS -10.5f
C2432 t<4>.n68 VSS -2.57f
C2433 t<4>.n69 VSS 2.5f
C2434 t<4>.n70 VSS -9.41f
C2435 t<4>.n71 VSS 2.5f
C2436 t<4>.n72 VSS 1.22f
C2437 t<4>.n73 VSS -2.57f
C2438 t<4>.n74 VSS 1.4f
C2439 t<4>.n75 VSS 0.873f
C2440 t<4>.n76 VSS 1.4f
C2441 t<4>.n77 VSS -2.57f
C2442 t<4>.n78 VSS -2.57f
C2443 t<4>.n79 VSS 2.5f
C2444 t<4>.n80 VSS -9.41f
C2445 t<4>.n81 VSS 2.5f
C2446 t<4>.n82 VSS 1.22f
C2447 t<4>.n83 VSS 1.65f
C2448 t<4>.n84 VSS 0.812f
C2449 t<4>.n85 VSS 1.34f
C2450 t<4>.n86 VSS 0.699f
C2451 t<4>.n87 VSS -2.9f
C2452 t<4>.n88 VSS 0.256f
C2453 t<4>.n89 VSS 1.91f
C2454 t<4>.n90 VSS 0.462f
C2455 t<4>.n91 VSS 3.17f
C2456 t<4>.n92 VSS 3.82f
C2457 t<4>.n93 VSS 3.38f
C2458 t<4>.n94 VSS -11.3f
C2459 t<4>.n95 VSS 37.7f
C2460 t<4>.n96 VSS 57.6f
C2461 t<4>.n97 VSS -16.7f
C2462 t<4>.n98 VSS -1.16f
C2463 t<4>.n99 VSS 1.22f
C2464 t<4>.n100 VSS 2.5f
C2465 t<4>.n101 VSS -9.41f
C2466 t<4>.n102 VSS -2.57f
C2467 t<4>.n103 VSS 1.4f
C2468 t<4>.n104 VSS 0.873f
C2469 t<4>.n105 VSS 1.41f
C2470 t<4>.n106 VSS 1.22f
C2471 t<4>.n107 VSS 2.5f
C2472 t<4>.n108 VSS -9.41f
C2473 t<4>.n109 VSS -2.57f
C2474 t<4>.n110 VSS 1.4f
C2475 t<4>.n111 VSS 0.873f
C2476 t<4>.n112 VSS 1.41f
C2477 t<4>.n113 VSS 1.22f
C2478 t<4>.n114 VSS 2.5f
C2479 t<4>.n115 VSS -9.41f
C2480 t<4>.n116 VSS -2.57f
C2481 t<4>.n117 VSS 1.4f
C2482 t<4>.n118 VSS 0.873f
C2483 t<4>.n119 VSS 1.41f
C2484 t<4>.n120 VSS 1.22f
C2485 t<4>.n121 VSS 2.5f
C2486 t<4>.n122 VSS -9.41f
C2487 t<4>.n123 VSS -2.57f
C2488 t<4>.n124 VSS 1.4f
C2489 t<4>.n125 VSS 0.873f
C2490 t<4>.n126 VSS 1.41f
C2491 t<4>.n127 VSS 1.22f
C2492 t<4>.n128 VSS 2.5f
C2493 t<4>.n129 VSS -9.41f
C2494 t<4>.n130 VSS -2.57f
C2495 t<4>.n131 VSS 1.4f
C2496 t<4>.n132 VSS 0.873f
C2497 t<4>.n133 VSS 1.41f
C2498 t<4>.n134 VSS 1.22f
C2499 t<4>.n135 VSS 2.5f
C2500 t<4>.n136 VSS -9.41f
C2501 t<4>.n137 VSS -2.57f
C2502 t<4>.n138 VSS 1.34f
C2503 t<4>.n139 VSS 0.699f
C2504 t<4>.n140 VSS 0.236f
C2505 t<4>.n141 VSS 0.927f
C2506 t<4>.n142 VSS -15.7f
C2507 t<4>.n143 VSS -9.41f
C2508 t<4>.n144 VSS 2.5f
C2509 t<4>.n145 VSS -2.57f
C2510 t<4>.n146 VSS -10.5f
C2511 t<4>.n147 VSS 1.4f
C2512 t<4>.n148 VSS -2.57f
C2513 t<4>.n149 VSS -9.41f
C2514 t<4>.n150 VSS 2.5f
C2515 t<4>.n151 VSS -2.57f
C2516 t<4>.n152 VSS -10.5f
C2517 t<4>.n153 VSS 1.4f
C2518 t<4>.n154 VSS -2.57f
C2519 t<4>.n155 VSS -9.41f
C2520 t<4>.n156 VSS 2.5f
C2521 t<4>.n157 VSS -2.57f
C2522 t<4>.n158 VSS -10.5f
C2523 t<4>.n159 VSS 1.4f
C2524 t<4>.n160 VSS -2.57f
C2525 t<4>.n161 VSS -9.41f
C2526 t<4>.n162 VSS 2.5f
C2527 t<4>.n163 VSS -2.57f
C2528 t<4>.n164 VSS -10.5f
C2529 t<4>.n165 VSS 1.4f
C2530 t<4>.n166 VSS -2.57f
C2531 t<4>.n167 VSS -9.41f
C2532 t<4>.n168 VSS 2.5f
C2533 t<4>.n169 VSS -2.57f
C2534 t<4>.n170 VSS -10.5f
C2535 t<4>.n171 VSS 1.4f
C2536 t<4>.n172 VSS -2.57f
C2537 t<4>.n173 VSS -9.41f
C2538 t<4>.n174 VSS 2.5f
C2539 t<4>.n175 VSS -2.57f
C2540 t<4>.n176 VSS -10.6f
C2541 t<4>.n177 VSS 0.699f
C2542 t<4>.n178 VSS 0.279f
C2543 t<4>.n179 VSS 0.699f
C2544 t<4>.n180 VSS 0.438f
C2545 t<4>.n181 VSS -0.149f
C2546 t<4>.n182 VSS 10f
C2547 t<4>.n183 VSS 0.489f
C2548 t<4>.n184 VSS -10.4f
C2549 t<4>.n185 VSS 0.78f
C2550 t<4>.n186 VSS 0.136f
C2551 t<4>.n187 VSS 5.84f
C2552 t<4>.n188 VSS 4.77f
C2553 tb<2>.n0 VSS -0.935f
C2554 tb<2>.n1 VSS 0.36f
C2555 tb<2>.n2 VSS -0.206f
C2556 tb<2>.n3 VSS 0.279f
C2557 tb<2>.n4 VSS -2.94f
C2558 tb<2>.n5 VSS -0.733f
C2559 tb<2>.n6 VSS 0.293f
C2560 tb<2>.n7 VSS 2.11f
C2561 tb<2>.n8 VSS 9.75f
C2562 tb<2>.n9 VSS 9.75f
C2563 tb<2>.n10 VSS -1.07f
C2564 tb<2>.n11 VSS 0.683f
C2565 tb<2>.n12 VSS 0.286f
C2566 tb<2>.n13 VSS -0.75f
C2567 tb<2>.n14 VSS -3.01f
C2568 tb<2>.n15 VSS -0.137f
C2569 tb<2>.n16 VSS 0.602f
C2570 tb<2>.n17 VSS 0.494f
C2571 hgu_cdac_8bit_array_3.drv<0>.t1 VSS 0.0151f
C2572 hgu_cdac_8bit_array_3.drv<0>.t0 VSS 0.0308f
C2573 hgu_cdac_8bit_array_3.drv<0>.n0 VSS 1.41f
C2574 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n0 VSS 1.01f
C2575 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n1 VSS 2.29f
C2576 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n2 VSS 0.757f
C2577 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n3 VSS -0.386f
C2578 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n4 VSS -0.507f
C2579 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t5 VSS 0.0314f
C2580 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t7 VSS 0.0314f
C2581 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n5 VSS 0.232f
C2582 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t2 VSS 0.0629f
C2583 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t0 VSS 0.0629f
C2584 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n6 VSS 0.419f
C2585 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n7 VSS 4.96f
C2586 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t4 VSS 0.0314f
C2587 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t6 VSS 0.0314f
C2588 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n8 VSS 0.233f
C2589 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t1 VSS 0.0629f
C2590 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.t3 VSS 0.0629f
C2591 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n9 VSS 0.478f
C2592 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n10 VSS 2.34f
C2593 hgu_cdac_8bit_array_3.hgu_cdac_cap_4_0.CBOT.n11 VSS 6.79f
C2594 hgu_cdac_8bit_array_2.drv<0>.t1 VSS 0.0129f
C2595 hgu_cdac_8bit_array_2.drv<0>.t0 VSS 0.0275f
C2596 hgu_cdac_8bit_array_2.drv<0>.n0 VSS 1.52f
C2597 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n0 VSS 0.89f
C2598 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n1 VSS 2.59f
C2599 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n2 VSS -0.371f
C2600 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n3 VSS 0.277f
C2601 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n4 VSS 2.47f
C2602 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t1 VSS 0.0595f
C2603 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t2 VSS 0.0595f
C2604 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n5 VSS 0.451f
C2605 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t6 VSS 0.0297f
C2606 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t7 VSS 0.0297f
C2607 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n6 VSS 0.219f
C2608 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t3 VSS 0.0595f
C2609 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t0 VSS 0.0595f
C2610 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n7 VSS 0.453f
C2611 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t4 VSS 0.0297f
C2612 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.t5 VSS 0.0297f
C2613 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n8 VSS 0.219f
C2614 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n9 VSS 2.42f
C2615 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n10 VSS -0.397f
C2616 hgu_cdac_8bit_array_2.hgu_cdac_cap_4_0.CBOT.n11 VSS 5.99f
C2617 hgu_cdac_8bit_array_2.drv<1:0>.t2 VSS 0.0213f
C2618 hgu_cdac_8bit_array_2.drv<1:0>.t3 VSS 0.0213f
C2619 hgu_cdac_8bit_array_2.drv<1:0>.n0 VSS 0.166f
C2620 hgu_cdac_8bit_array_2.drv<1:0>.t0 VSS 0.0426f
C2621 hgu_cdac_8bit_array_2.drv<1:0>.t1 VSS 0.0426f
C2622 hgu_cdac_8bit_array_2.drv<1:0>.n1 VSS 0.301f
C2623 hgu_cdac_8bit_array_2.drv<1:0>.n2 VSS 2.22f
C2624 hgu_cdac_8bit_array_2.drv<15:0>.n0 VSS 3.64f
C2625 hgu_cdac_8bit_array_2.drv<15:0>.n1 VSS 1.12f
C2626 hgu_cdac_8bit_array_2.drv<15:0>.n2 VSS 0.643f
C2627 hgu_cdac_8bit_array_2.drv<15:0>.n3 VSS 0.679f
C2628 hgu_cdac_8bit_array_2.drv<15:0>.n4 VSS 0.643f
C2629 hgu_cdac_8bit_array_2.drv<15:0>.n5 VSS 0.679f
C2630 hgu_cdac_8bit_array_2.drv<15:0>.n6 VSS 0.643f
C2631 hgu_cdac_8bit_array_2.drv<15:0>.n7 VSS 0.391f
C2632 hgu_cdac_8bit_array_2.drv<15:0>.n8 VSS 0.643f
C2633 hgu_cdac_8bit_array_2.drv<15:0>.n9 VSS 0.679f
C2634 hgu_cdac_8bit_array_2.drv<15:0>.n10 VSS 0.643f
C2635 hgu_cdac_8bit_array_2.drv<15:0>.n11 VSS 0.679f
C2636 hgu_cdac_8bit_array_2.drv<15:0>.n12 VSS 0.643f
C2637 hgu_cdac_8bit_array_2.drv<15:0>.n13 VSS 0.679f
C2638 hgu_cdac_8bit_array_2.drv<15:0>.n14 VSS 0.643f
C2639 hgu_cdac_8bit_array_2.drv<15:0>.n15 VSS 3.67f
C2640 hgu_cdac_8bit_array_2.drv<15:0>.t0 VSS 0.0898f
C2641 hgu_cdac_8bit_array_2.drv<15:0>.t8 VSS 0.0898f
C2642 hgu_cdac_8bit_array_2.drv<15:0>.n16 VSS 0.684f
C2643 hgu_cdac_8bit_array_2.drv<15:0>.t21 VSS 0.0449f
C2644 hgu_cdac_8bit_array_2.drv<15:0>.t29 VSS 0.0449f
C2645 hgu_cdac_8bit_array_2.drv<15:0>.n17 VSS 0.329f
C2646 hgu_cdac_8bit_array_2.drv<15:0>.n18 VSS -1.48f
C2647 hgu_cdac_8bit_array_2.drv<15:0>.n19 VSS -0.941f
C2648 hgu_cdac_8bit_array_2.drv<15:0>.n20 VSS -1.51f
C2649 hgu_cdac_8bit_array_2.drv<15:0>.n21 VSS -1.51f
C2650 hgu_cdac_8bit_array_2.drv<15:0>.n22 VSS -0.941f
C2651 hgu_cdac_8bit_array_2.drv<15:0>.n23 VSS -1.48f
C2652 hgu_cdac_8bit_array_2.drv<15:0>.n24 VSS 3.4f
C2653 hgu_cdac_8bit_array_2.drv<15:0>.n25 VSS 7.79f
C2654 hgu_cdac_8bit_array_2.drv<15:0>.t10 VSS 0.0898f
C2655 hgu_cdac_8bit_array_2.drv<15:0>.t11 VSS 0.0898f
C2656 hgu_cdac_8bit_array_2.drv<15:0>.n26 VSS 0.644f
C2657 hgu_cdac_8bit_array_2.drv<15:0>.t31 VSS 0.0449f
C2658 hgu_cdac_8bit_array_2.drv<15:0>.t16 VSS 0.0449f
C2659 hgu_cdac_8bit_array_2.drv<15:0>.n27 VSS 0.317f
C2660 hgu_cdac_8bit_array_2.drv<15:0>.t1 VSS 0.0898f
C2661 hgu_cdac_8bit_array_2.drv<15:0>.t9 VSS 0.0898f
C2662 hgu_cdac_8bit_array_2.drv<15:0>.n28 VSS 0.684f
C2663 hgu_cdac_8bit_array_2.drv<15:0>.t22 VSS 0.0449f
C2664 hgu_cdac_8bit_array_2.drv<15:0>.t30 VSS 0.0449f
C2665 hgu_cdac_8bit_array_2.drv<15:0>.n29 VSS 0.33f
C2666 hgu_cdac_8bit_array_2.drv<15:0>.n30 VSS 0.43f
C2667 hgu_cdac_8bit_array_2.drv<15:0>.n31 VSS 0.367f
C2668 hgu_cdac_8bit_array_2.drv<15:0>.n32 VSS 3.39f
C2669 hgu_cdac_8bit_array_2.drv<15:0>.n33 VSS -1.48f
C2670 hgu_cdac_8bit_array_2.drv<15:0>.n34 VSS -0.941f
C2671 hgu_cdac_8bit_array_2.drv<15:0>.n35 VSS -1.51f
C2672 hgu_cdac_8bit_array_2.drv<15:0>.n36 VSS -1.51f
C2673 hgu_cdac_8bit_array_2.drv<15:0>.n37 VSS -0.941f
C2674 hgu_cdac_8bit_array_2.drv<15:0>.n38 VSS -1.48f
C2675 hgu_cdac_8bit_array_2.drv<15:0>.n39 VSS 3.4f
C2676 hgu_cdac_8bit_array_2.drv<15:0>.n40 VSS 7.39f
C2677 hgu_cdac_8bit_array_2.drv<15:0>.t13 VSS 0.0898f
C2678 hgu_cdac_8bit_array_2.drv<15:0>.t2 VSS 0.0898f
C2679 hgu_cdac_8bit_array_2.drv<15:0>.n41 VSS 0.684f
C2680 hgu_cdac_8bit_array_2.drv<15:0>.t18 VSS 0.0449f
C2681 hgu_cdac_8bit_array_2.drv<15:0>.t23 VSS 0.0449f
C2682 hgu_cdac_8bit_array_2.drv<15:0>.n42 VSS 0.33f
C2683 hgu_cdac_8bit_array_2.drv<15:0>.n43 VSS 0.398f
C2684 hgu_cdac_8bit_array_2.drv<15:0>.t4 VSS 0.0898f
C2685 hgu_cdac_8bit_array_2.drv<15:0>.t12 VSS 0.0898f
C2686 hgu_cdac_8bit_array_2.drv<15:0>.n44 VSS 0.644f
C2687 hgu_cdac_8bit_array_2.drv<15:0>.t25 VSS 0.0449f
C2688 hgu_cdac_8bit_array_2.drv<15:0>.t17 VSS 0.0449f
C2689 hgu_cdac_8bit_array_2.drv<15:0>.n45 VSS 0.317f
C2690 hgu_cdac_8bit_array_2.drv<15:0>.n46 VSS 0.365f
C2691 hgu_cdac_8bit_array_2.drv<15:0>.n47 VSS 3.39f
C2692 hgu_cdac_8bit_array_2.drv<15:0>.n48 VSS -1.48f
C2693 hgu_cdac_8bit_array_2.drv<15:0>.n49 VSS -0.941f
C2694 hgu_cdac_8bit_array_2.drv<15:0>.n50 VSS -1.51f
C2695 hgu_cdac_8bit_array_2.drv<15:0>.n51 VSS -1.51f
C2696 hgu_cdac_8bit_array_2.drv<15:0>.n52 VSS -0.941f
C2697 hgu_cdac_8bit_array_2.drv<15:0>.n53 VSS -1.48f
C2698 hgu_cdac_8bit_array_2.drv<15:0>.n54 VSS 3.4f
C2699 hgu_cdac_8bit_array_2.drv<15:0>.n55 VSS 7.39f
C2700 hgu_cdac_8bit_array_2.drv<15:0>.t14 VSS 0.0898f
C2701 hgu_cdac_8bit_array_2.drv<15:0>.t15 VSS 0.0898f
C2702 hgu_cdac_8bit_array_2.drv<15:0>.n56 VSS 0.684f
C2703 hgu_cdac_8bit_array_2.drv<15:0>.t19 VSS 0.0449f
C2704 hgu_cdac_8bit_array_2.drv<15:0>.t20 VSS 0.0449f
C2705 hgu_cdac_8bit_array_2.drv<15:0>.n57 VSS 0.33f
C2706 hgu_cdac_8bit_array_2.drv<15:0>.n58 VSS 0.351f
C2707 hgu_cdac_8bit_array_2.drv<15:0>.t5 VSS 0.0898f
C2708 hgu_cdac_8bit_array_2.drv<15:0>.t6 VSS 0.0898f
C2709 hgu_cdac_8bit_array_2.drv<15:0>.n59 VSS 0.684f
C2710 hgu_cdac_8bit_array_2.drv<15:0>.t26 VSS 0.0449f
C2711 hgu_cdac_8bit_array_2.drv<15:0>.t27 VSS 0.0449f
C2712 hgu_cdac_8bit_array_2.drv<15:0>.n60 VSS 0.33f
C2713 hgu_cdac_8bit_array_2.drv<15:0>.n61 VSS 0.363f
C2714 hgu_cdac_8bit_array_2.drv<15:0>.n62 VSS 3.4f
C2715 hgu_cdac_8bit_array_2.drv<15:0>.n63 VSS -1.78f
C2716 hgu_cdac_8bit_array_2.drv<15:0>.n64 VSS -1.51f
C2717 hgu_cdac_8bit_array_2.drv<15:0>.n65 VSS -0.941f
C2718 hgu_cdac_8bit_array_2.drv<15:0>.n66 VSS -1.48f
C2719 hgu_cdac_8bit_array_2.drv<15:0>.n67 VSS 3.4f
C2720 hgu_cdac_8bit_array_2.drv<15:0>.n68 VSS 7.39f
C2721 hgu_cdac_8bit_array_2.drv<15:0>.t3 VSS 0.0898f
C2722 hgu_cdac_8bit_array_2.drv<15:0>.t7 VSS 0.0898f
C2723 hgu_cdac_8bit_array_2.drv<15:0>.n69 VSS 0.68f
C2724 hgu_cdac_8bit_array_2.drv<15:0>.t24 VSS 0.0449f
C2725 hgu_cdac_8bit_array_2.drv<15:0>.t28 VSS 0.0449f
C2726 hgu_cdac_8bit_array_2.drv<15:0>.n70 VSS 0.33f
C2727 hgu_cdac_8bit_array_2.drv<15:0>.n71 VSS 10.1f
C2728 hgu_cdac_8bit_array_2.drv<15:0>.n72 VSS -0.395f
C2729 hgu_cdac_8bit_array_2.drv<15:0>.n73 VSS -1.48f
C2730 hgu_cdac_8bit_array_2.drv<15:0>.n74 VSS 3.75f
C2731 hgu_cdac_8bit_array_2.drv<15:0>.n75 VSS -1.48f
C2732 hgu_cdac_8bit_array_2.drv<15:0>.n76 VSS -0.395f
C2733 hgu_cdac_8bit_array_2.drv<15:0>.n77 VSS -0.395f
C2734 hgu_cdac_8bit_array_2.drv<15:0>.n78 VSS -1.48f
C2735 hgu_cdac_8bit_array_2.drv<15:0>.n79 VSS 3.75f
C2736 hgu_cdac_8bit_array_2.drv<15:0>.n80 VSS -1.48f
C2737 hgu_cdac_8bit_array_2.drv<15:0>.n81 VSS -0.395f
C2738 hgu_cdac_8bit_array_2.drv<15:0>.n82 VSS -0.395f
C2739 hgu_cdac_8bit_array_2.drv<15:0>.n83 VSS -1.48f
C2740 hgu_cdac_8bit_array_2.drv<15:0>.n84 VSS 3.75f
C2741 hgu_cdac_8bit_array_2.drv<15:0>.n85 VSS -1.48f
C2742 hgu_cdac_8bit_array_2.drv<15:0>.n86 VSS -0.395f
C2743 hgu_cdac_8bit_array_2.drv<15:0>.n87 VSS -0.395f
C2744 hgu_cdac_8bit_array_2.drv<15:0>.n88 VSS -1.48f
C2745 hgu_cdac_8bit_array_2.drv<15:0>.n89 VSS 3.75f
C2746 hgu_cdac_8bit_array_2.drv<15:0>.n90 VSS -1.48f
C2747 hgu_cdac_8bit_array_2.drv<15:0>.n91 VSS -0.395f
C2748 hgu_cdac_8bit_array_2.drv<15:0>.n92 VSS -0.395f
C2749 hgu_cdac_8bit_array_2.drv<15:0>.n93 VSS -1.48f
C2750 hgu_cdac_8bit_array_2.drv<15:0>.n94 VSS -1.48f
C2751 hgu_cdac_8bit_array_2.drv<15:0>.n95 VSS -0.941f
C2752 hgu_cdac_8bit_array_2.drv<15:0>.n96 VSS -1.51f
C2753 hgu_cdac_8bit_array_2.drv<15:0>.n97 VSS -1.51f
C2754 hgu_cdac_8bit_array_2.drv<15:0>.n98 VSS -0.941f
C2755 hgu_cdac_8bit_array_2.drv<15:0>.n99 VSS -1.48f
C2756 hgu_cdac_8bit_array_2.drv<15:0>.n100 VSS 5.26f
C2757 hgu_cdac_8bit_array_2.drv<15:0>.n101 VSS -1.31f
C2758 hgu_cdac_8bit_array_2.drv<15:0>.n102 VSS -1.48f
C2759 hgu_cdac_8bit_array_2.drv<15:0>.n103 VSS 5.26f
C2760 hgu_cdac_8bit_array_2.drv<15:0>.n104 VSS 3.91f
C2761 hgu_cdac_8bit_array_2.drv<15:0>.n105 VSS 0.669f
C2762 hgu_cdac_8bit_array_2.drv<15:0>.n106 VSS -0.395f
C2763 hgu_cdac_8bit_array_2.drv<15:0>.n107 VSS -1.48f
C2764 hgu_cdac_8bit_array_2.drv<15:0>.n108 VSS 5.26f
C2765 hgu_cdac_8bit_array_2.drv<15:0>.n109 VSS -1.48f
C2766 hgu_cdac_8bit_array_2.drv<15:0>.n110 VSS -0.395f
C2767 hgu_cdac_8bit_array_2.drv<15:0>.n111 VSS -0.395f
C2768 hgu_cdac_8bit_array_2.drv<15:0>.n112 VSS -1.48f
C2769 hgu_cdac_8bit_array_2.drv<15:0>.n113 VSS 5.26f
C2770 hgu_cdac_8bit_array_2.drv<15:0>.n114 VSS -1.48f
C2771 hgu_cdac_8bit_array_2.drv<15:0>.n115 VSS -0.395f
C2772 hgu_cdac_8bit_array_2.drv<15:0>.n116 VSS -0.395f
C2773 hgu_cdac_8bit_array_2.drv<15:0>.n117 VSS -1.51f
C2774 hgu_cdac_8bit_array_3.drv<1:0>.n0 VSS 0.247f
C2775 hgu_cdac_8bit_array_3.drv<1:0>.t2 VSS 0.0231f
C2776 hgu_cdac_8bit_array_3.drv<1:0>.t3 VSS 0.0231f
C2777 hgu_cdac_8bit_array_3.drv<1:0>.n1 VSS 0.181f
C2778 hgu_cdac_8bit_array_3.drv<1:0>.t1 VSS 0.0463f
C2779 hgu_cdac_8bit_array_3.drv<1:0>.t0 VSS 0.0463f
C2780 hgu_cdac_8bit_array_3.drv<1:0>.n2 VSS 0.327f
C2781 hgu_cdac_8bit_array_3.drv<1:0>.n3 VSS 1.53f
C2782 hgu_cdac_8bit_array_3.drv<1:0>.n4 VSS 5.16f
C2783 hgu_cdac_8bit_array_3.drv<15:0>.n0 VSS 0.714f
C2784 hgu_cdac_8bit_array_3.drv<15:0>.n1 VSS 0.677f
C2785 hgu_cdac_8bit_array_3.drv<15:0>.n2 VSS 0.714f
C2786 hgu_cdac_8bit_array_3.drv<15:0>.n3 VSS 0.677f
C2787 hgu_cdac_8bit_array_3.drv<15:0>.n4 VSS 0.412f
C2788 hgu_cdac_8bit_array_3.drv<15:0>.n5 VSS 0.677f
C2789 hgu_cdac_8bit_array_3.drv<15:0>.n6 VSS 0.714f
C2790 hgu_cdac_8bit_array_3.drv<15:0>.n7 VSS 0.677f
C2791 hgu_cdac_8bit_array_3.drv<15:0>.n8 VSS 0.714f
C2792 hgu_cdac_8bit_array_3.drv<15:0>.n9 VSS 0.677f
C2793 hgu_cdac_8bit_array_3.drv<15:0>.n10 VSS 0.714f
C2794 hgu_cdac_8bit_array_3.drv<15:0>.n11 VSS 0.677f
C2795 hgu_cdac_8bit_array_3.drv<15:0>.n12 VSS 0.714f
C2796 hgu_cdac_8bit_array_3.drv<15:0>.n13 VSS 1.14f
C2797 hgu_cdac_8bit_array_3.drv<15:0>.t21 VSS 0.0472f
C2798 hgu_cdac_8bit_array_3.drv<15:0>.t25 VSS 0.0472f
C2799 hgu_cdac_8bit_array_3.drv<15:0>.n14 VSS 0.349f
C2800 hgu_cdac_8bit_array_3.drv<15:0>.t9 VSS 0.0945f
C2801 hgu_cdac_8bit_array_3.drv<15:0>.t13 VSS 0.0945f
C2802 hgu_cdac_8bit_array_3.drv<15:0>.n15 VSS 0.629f
C2803 hgu_cdac_8bit_array_3.drv<15:0>.n16 VSS 3.65f
C2804 hgu_cdac_8bit_array_3.drv<15:0>.n17 VSS 0.187f
C2805 hgu_cdac_8bit_array_3.drv<15:0>.t27 VSS 0.0472f
C2806 hgu_cdac_8bit_array_3.drv<15:0>.t19 VSS 0.0472f
C2807 hgu_cdac_8bit_array_3.drv<15:0>.n18 VSS 0.334f
C2808 hgu_cdac_8bit_array_3.drv<15:0>.t29 VSS 0.0472f
C2809 hgu_cdac_8bit_array_3.drv<15:0>.t31 VSS 0.0472f
C2810 hgu_cdac_8bit_array_3.drv<15:0>.n19 VSS 0.349f
C2811 hgu_cdac_8bit_array_3.drv<15:0>.t1 VSS 0.0945f
C2812 hgu_cdac_8bit_array_3.drv<15:0>.t3 VSS 0.0945f
C2813 hgu_cdac_8bit_array_3.drv<15:0>.n20 VSS 0.719f
C2814 hgu_cdac_8bit_array_3.drv<15:0>.n21 VSS 0.453f
C2815 hgu_cdac_8bit_array_3.drv<15:0>.t15 VSS 0.0945f
C2816 hgu_cdac_8bit_array_3.drv<15:0>.t7 VSS 0.0945f
C2817 hgu_cdac_8bit_array_3.drv<15:0>.n22 VSS 0.678f
C2818 hgu_cdac_8bit_array_3.drv<15:0>.n23 VSS 0.385f
C2819 hgu_cdac_8bit_array_3.drv<15:0>.n24 VSS 3.26f
C2820 hgu_cdac_8bit_array_3.drv<15:0>.n25 VSS -5.57f
C2821 hgu_cdac_8bit_array_3.drv<15:0>.n26 VSS -1.56f
C2822 hgu_cdac_8bit_array_3.drv<15:0>.n27 VSS -0.99f
C2823 hgu_cdac_8bit_array_3.drv<15:0>.n28 VSS -1.59f
C2824 hgu_cdac_8bit_array_3.drv<15:0>.n29 VSS -1.59f
C2825 hgu_cdac_8bit_array_3.drv<15:0>.n30 VSS -0.99f
C2826 hgu_cdac_8bit_array_3.drv<15:0>.n31 VSS -1.56f
C2827 hgu_cdac_8bit_array_3.drv<15:0>.n32 VSS 3.57f
C2828 hgu_cdac_8bit_array_3.drv<15:0>.n33 VSS 7.71f
C2829 hgu_cdac_8bit_array_3.drv<15:0>.n34 VSS -1.56f
C2830 hgu_cdac_8bit_array_3.drv<15:0>.n35 VSS -0.99f
C2831 hgu_cdac_8bit_array_3.drv<15:0>.n36 VSS -1.59f
C2832 hgu_cdac_8bit_array_3.drv<15:0>.n37 VSS -1.59f
C2833 hgu_cdac_8bit_array_3.drv<15:0>.n38 VSS -0.99f
C2834 hgu_cdac_8bit_array_3.drv<15:0>.n39 VSS -1.56f
C2835 hgu_cdac_8bit_array_3.drv<15:0>.n40 VSS 5.53f
C2836 hgu_cdac_8bit_array_3.drv<15:0>.n41 VSS -1.56f
C2837 hgu_cdac_8bit_array_3.drv<15:0>.n42 VSS -0.99f
C2838 hgu_cdac_8bit_array_3.drv<15:0>.n43 VSS -1.59f
C2839 hgu_cdac_8bit_array_3.drv<15:0>.n44 VSS -1.59f
C2840 hgu_cdac_8bit_array_3.drv<15:0>.n45 VSS -0.99f
C2841 hgu_cdac_8bit_array_3.drv<15:0>.n46 VSS -1.56f
C2842 hgu_cdac_8bit_array_3.drv<15:0>.n47 VSS 5.53f
C2843 hgu_cdac_8bit_array_3.drv<15:0>.n48 VSS -1.38f
C2844 hgu_cdac_8bit_array_3.drv<15:0>.n49 VSS -1.56f
C2845 hgu_cdac_8bit_array_3.drv<15:0>.n50 VSS 5.53f
C2846 hgu_cdac_8bit_array_3.drv<15:0>.n51 VSS 4.16f
C2847 hgu_cdac_8bit_array_3.drv<15:0>.n52 VSS 0.667f
C2848 hgu_cdac_8bit_array_3.drv<15:0>.n53 VSS -0.416f
C2849 hgu_cdac_8bit_array_3.drv<15:0>.n54 VSS -1.56f
C2850 hgu_cdac_8bit_array_3.drv<15:0>.n55 VSS 5.54f
C2851 hgu_cdac_8bit_array_3.drv<15:0>.n56 VSS -1.56f
C2852 hgu_cdac_8bit_array_3.drv<15:0>.n57 VSS -0.416f
C2853 hgu_cdac_8bit_array_3.drv<15:0>.n58 VSS -0.416f
C2854 hgu_cdac_8bit_array_3.drv<15:0>.n59 VSS -1.56f
C2855 hgu_cdac_8bit_array_3.drv<15:0>.n60 VSS 5.54f
C2856 hgu_cdac_8bit_array_3.drv<15:0>.n61 VSS -1.56f
C2857 hgu_cdac_8bit_array_3.drv<15:0>.n62 VSS -0.416f
C2858 hgu_cdac_8bit_array_3.drv<15:0>.n63 VSS -0.416f
C2859 hgu_cdac_8bit_array_3.drv<15:0>.n64 VSS -1.56f
C2860 hgu_cdac_8bit_array_3.drv<15:0>.n65 VSS 5.54f
C2861 hgu_cdac_8bit_array_3.drv<15:0>.n66 VSS -1.56f
C2862 hgu_cdac_8bit_array_3.drv<15:0>.n67 VSS -0.416f
C2863 hgu_cdac_8bit_array_3.drv<15:0>.n68 VSS -0.416f
C2864 hgu_cdac_8bit_array_3.drv<15:0>.n69 VSS -1.56f
C2865 hgu_cdac_8bit_array_3.drv<15:0>.n70 VSS 3.94f
C2866 hgu_cdac_8bit_array_3.drv<15:0>.n71 VSS -1.56f
C2867 hgu_cdac_8bit_array_3.drv<15:0>.n72 VSS -0.416f
C2868 hgu_cdac_8bit_array_3.drv<15:0>.n73 VSS -0.416f
C2869 hgu_cdac_8bit_array_3.drv<15:0>.n74 VSS -1.56f
C2870 hgu_cdac_8bit_array_3.drv<15:0>.t17 VSS 0.0472f
C2871 hgu_cdac_8bit_array_3.drv<15:0>.t23 VSS 0.0472f
C2872 hgu_cdac_8bit_array_3.drv<15:0>.n75 VSS 0.333f
C2873 hgu_cdac_8bit_array_3.drv<15:0>.t5 VSS 0.0945f
C2874 hgu_cdac_8bit_array_3.drv<15:0>.t11 VSS 0.0945f
C2875 hgu_cdac_8bit_array_3.drv<15:0>.n76 VSS 0.679f
C2876 hgu_cdac_8bit_array_3.drv<15:0>.n77 VSS 0.385f
C2877 hgu_cdac_8bit_array_3.drv<15:0>.t28 VSS 0.0472f
C2878 hgu_cdac_8bit_array_3.drv<15:0>.t30 VSS 0.0472f
C2879 hgu_cdac_8bit_array_3.drv<15:0>.n78 VSS 0.349f
C2880 hgu_cdac_8bit_array_3.drv<15:0>.t0 VSS 0.0945f
C2881 hgu_cdac_8bit_array_3.drv<15:0>.t2 VSS 0.0945f
C2882 hgu_cdac_8bit_array_3.drv<15:0>.n79 VSS 0.719f
C2883 hgu_cdac_8bit_array_3.drv<15:0>.n80 VSS 0.419f
C2884 hgu_cdac_8bit_array_3.drv<15:0>.n81 VSS 3.26f
C2885 hgu_cdac_8bit_array_3.drv<15:0>.n82 VSS -1.56f
C2886 hgu_cdac_8bit_array_3.drv<15:0>.n83 VSS -0.99f
C2887 hgu_cdac_8bit_array_3.drv<15:0>.n84 VSS -1.59f
C2888 hgu_cdac_8bit_array_3.drv<15:0>.n85 VSS -1.59f
C2889 hgu_cdac_8bit_array_3.drv<15:0>.n86 VSS -0.99f
C2890 hgu_cdac_8bit_array_3.drv<15:0>.n87 VSS -1.56f
C2891 hgu_cdac_8bit_array_3.drv<15:0>.n88 VSS 3.57f
C2892 hgu_cdac_8bit_array_3.drv<15:0>.n89 VSS 7.42f
C2893 hgu_cdac_8bit_array_3.drv<15:0>.n90 VSS -1.87f
C2894 hgu_cdac_8bit_array_3.drv<15:0>.n91 VSS -1.59f
C2895 hgu_cdac_8bit_array_3.drv<15:0>.n92 VSS -0.99f
C2896 hgu_cdac_8bit_array_3.drv<15:0>.n93 VSS -1.56f
C2897 hgu_cdac_8bit_array_3.drv<15:0>.n94 VSS 3.57f
C2898 hgu_cdac_8bit_array_3.drv<15:0>.t16 VSS 0.0472f
C2899 hgu_cdac_8bit_array_3.drv<15:0>.t22 VSS 0.0472f
C2900 hgu_cdac_8bit_array_3.drv<15:0>.n95 VSS 0.349f
C2901 hgu_cdac_8bit_array_3.drv<15:0>.t4 VSS 0.0945f
C2902 hgu_cdac_8bit_array_3.drv<15:0>.t10 VSS 0.0945f
C2903 hgu_cdac_8bit_array_3.drv<15:0>.n96 VSS 0.719f
C2904 hgu_cdac_8bit_array_3.drv<15:0>.n97 VSS 0.382f
C2905 hgu_cdac_8bit_array_3.drv<15:0>.t18 VSS 0.0472f
C2906 hgu_cdac_8bit_array_3.drv<15:0>.t20 VSS 0.0472f
C2907 hgu_cdac_8bit_array_3.drv<15:0>.n98 VSS 0.349f
C2908 hgu_cdac_8bit_array_3.drv<15:0>.t6 VSS 0.0945f
C2909 hgu_cdac_8bit_array_3.drv<15:0>.t8 VSS 0.0945f
C2910 hgu_cdac_8bit_array_3.drv<15:0>.n99 VSS 0.719f
C2911 hgu_cdac_8bit_array_3.drv<15:0>.n100 VSS 0.377f
C2912 hgu_cdac_8bit_array_3.drv<15:0>.n101 VSS 3.26f
C2913 hgu_cdac_8bit_array_3.drv<15:0>.n102 VSS 7.42f
C2914 hgu_cdac_8bit_array_3.drv<15:0>.t24 VSS 0.0472f
C2915 hgu_cdac_8bit_array_3.drv<15:0>.t26 VSS 0.0472f
C2916 hgu_cdac_8bit_array_3.drv<15:0>.n103 VSS 0.334f
C2917 hgu_cdac_8bit_array_3.drv<15:0>.t12 VSS 0.0945f
C2918 hgu_cdac_8bit_array_3.drv<15:0>.t14 VSS 0.0945f
C2919 hgu_cdac_8bit_array_3.drv<15:0>.n104 VSS 0.701f
C2920 hgu_cdac_8bit_array_3.drv<15:0>.n105 VSS 3.67f
C2921 hgu_cdac_8bit_array_3.drv<15:0>.n106 VSS 10.4f
C2922 hgu_cdac_8bit_array_3.drv<15:0>.n107 VSS -0.416f
C2923 hgu_cdac_8bit_array_3.drv<15:0>.n108 VSS -1.56f
C2924 hgu_cdac_8bit_array_3.drv<15:0>.n109 VSS 3.94f
C2925 hgu_cdac_8bit_array_3.drv<15:0>.n110 VSS -1.56f
C2926 hgu_cdac_8bit_array_3.drv<15:0>.n111 VSS -0.416f
C2927 hgu_cdac_8bit_array_3.drv<15:0>.n112 VSS -0.416f
C2928 hgu_cdac_8bit_array_3.drv<15:0>.n113 VSS -1.56f
C2929 hgu_cdac_8bit_array_3.drv<15:0>.n114 VSS 3.94f
C2930 hgu_cdac_8bit_array_3.drv<15:0>.n115 VSS -1.56f
C2931 hgu_cdac_8bit_array_3.drv<15:0>.n116 VSS -0.416f
C2932 hgu_cdac_8bit_array_3.drv<15:0>.n117 VSS -0.416f
C2933 hgu_cdac_8bit_array_3.drv<15:0>.n118 VSS -1.59f
C2934 hgu_cdac_8bit_array_2.drv<63:0>.n0 VSS 4.16f
C2935 hgu_cdac_8bit_array_2.drv<63:0>.n1 VSS 4.15f
C2936 hgu_cdac_8bit_array_2.drv<63:0>.n2 VSS 4.28f
C2937 hgu_cdac_8bit_array_2.drv<63:0>.t45 VSS 0.104f
C2938 hgu_cdac_8bit_array_2.drv<63:0>.t1 VSS 0.104f
C2939 hgu_cdac_8bit_array_2.drv<63:0>.n3 VSS 0.793f
C2940 hgu_cdac_8bit_array_2.drv<63:0>.t126 VSS 0.0521f
C2941 hgu_cdac_8bit_array_2.drv<63:0>.t82 VSS 0.0521f
C2942 hgu_cdac_8bit_array_2.drv<63:0>.n4 VSS 0.383f
C2943 hgu_cdac_8bit_array_2.drv<63:0>.n5 VSS 0.474f
C2944 hgu_cdac_8bit_array_2.drv<63:0>.t33 VSS 0.104f
C2945 hgu_cdac_8bit_array_2.drv<63:0>.t55 VSS 0.104f
C2946 hgu_cdac_8bit_array_2.drv<63:0>.n6 VSS 0.748f
C2947 hgu_cdac_8bit_array_2.drv<63:0>.t114 VSS 0.0521f
C2948 hgu_cdac_8bit_array_2.drv<63:0>.t72 VSS 0.0521f
C2949 hgu_cdac_8bit_array_2.drv<63:0>.n7 VSS 0.367f
C2950 hgu_cdac_8bit_array_2.drv<63:0>.t62 VSS 0.104f
C2951 hgu_cdac_8bit_array_2.drv<63:0>.t25 VSS 0.104f
C2952 hgu_cdac_8bit_array_2.drv<63:0>.n8 VSS 0.793f
C2953 hgu_cdac_8bit_array_2.drv<63:0>.t79 VSS 0.0521f
C2954 hgu_cdac_8bit_array_2.drv<63:0>.t106 VSS 0.0521f
C2955 hgu_cdac_8bit_array_2.drv<63:0>.n9 VSS 0.383f
C2956 hgu_cdac_8bit_array_2.drv<63:0>.n10 VSS 0.493f
C2957 hgu_cdac_8bit_array_2.drv<63:0>.n11 VSS 0.395f
C2958 hgu_cdac_8bit_array_2.drv<63:0>.n12 VSS 3.92f
C2959 hgu_cdac_8bit_array_2.drv<63:0>.n13 VSS -5.78f
C2960 hgu_cdac_8bit_array_2.drv<63:0>.t59 VSS 0.104f
C2961 hgu_cdac_8bit_array_2.drv<63:0>.t51 VSS 0.104f
C2962 hgu_cdac_8bit_array_2.drv<63:0>.n14 VSS 0.793f
C2963 hgu_cdac_8bit_array_2.drv<63:0>.t76 VSS 0.0521f
C2964 hgu_cdac_8bit_array_2.drv<63:0>.t68 VSS 0.0521f
C2965 hgu_cdac_8bit_array_2.drv<63:0>.n15 VSS 0.383f
C2966 hgu_cdac_8bit_array_2.drv<63:0>.n16 VSS 0.418f
C2967 hgu_cdac_8bit_array_2.drv<63:0>.t10 VSS 0.104f
C2968 hgu_cdac_8bit_array_2.drv<63:0>.t38 VSS 0.104f
C2969 hgu_cdac_8bit_array_2.drv<63:0>.n17 VSS 0.793f
C2970 hgu_cdac_8bit_array_2.drv<63:0>.t91 VSS 0.0521f
C2971 hgu_cdac_8bit_array_2.drv<63:0>.t119 VSS 0.0521f
C2972 hgu_cdac_8bit_array_2.drv<63:0>.n18 VSS 0.383f
C2973 hgu_cdac_8bit_array_2.drv<63:0>.n19 VSS 0.409f
C2974 hgu_cdac_8bit_array_2.drv<63:0>.n20 VSS 3.94f
C2975 hgu_cdac_8bit_array_2.drv<63:0>.n21 VSS -1.72f
C2976 hgu_cdac_8bit_array_2.drv<63:0>.n22 VSS -1.09f
C2977 hgu_cdac_8bit_array_2.drv<63:0>.n23 VSS -1.75f
C2978 hgu_cdac_8bit_array_2.drv<63:0>.n24 VSS -1.75f
C2979 hgu_cdac_8bit_array_2.drv<63:0>.n25 VSS -1.09f
C2980 hgu_cdac_8bit_array_2.drv<63:0>.n26 VSS -1.72f
C2981 hgu_cdac_8bit_array_2.drv<63:0>.n27 VSS 3.94f
C2982 hgu_cdac_8bit_array_2.drv<63:0>.n28 VSS 8.53f
C2983 hgu_cdac_8bit_array_2.drv<63:0>.t27 VSS 0.104f
C2984 hgu_cdac_8bit_array_2.drv<63:0>.t34 VSS 0.104f
C2985 hgu_cdac_8bit_array_2.drv<63:0>.n29 VSS 0.747f
C2986 hgu_cdac_8bit_array_2.drv<63:0>.t107 VSS 0.0521f
C2987 hgu_cdac_8bit_array_2.drv<63:0>.t115 VSS 0.0521f
C2988 hgu_cdac_8bit_array_2.drv<63:0>.n30 VSS 0.368f
C2989 hgu_cdac_8bit_array_2.drv<63:0>.t57 VSS 0.104f
C2990 hgu_cdac_8bit_array_2.drv<63:0>.t19 VSS 0.104f
C2991 hgu_cdac_8bit_array_2.drv<63:0>.n31 VSS 0.792f
C2992 hgu_cdac_8bit_array_2.drv<63:0>.t74 VSS 0.0521f
C2993 hgu_cdac_8bit_array_2.drv<63:0>.t100 VSS 0.0521f
C2994 hgu_cdac_8bit_array_2.drv<63:0>.n32 VSS 0.383f
C2995 hgu_cdac_8bit_array_2.drv<63:0>.n33 VSS 0.417f
C2996 hgu_cdac_8bit_array_2.drv<63:0>.t13 VSS 0.104f
C2997 hgu_cdac_8bit_array_2.drv<63:0>.t39 VSS 0.104f
C2998 hgu_cdac_8bit_array_2.drv<63:0>.n34 VSS 0.793f
C2999 hgu_cdac_8bit_array_2.drv<63:0>.t94 VSS 0.0521f
C3000 hgu_cdac_8bit_array_2.drv<63:0>.t120 VSS 0.0521f
C3001 hgu_cdac_8bit_array_2.drv<63:0>.n35 VSS 0.383f
C3002 hgu_cdac_8bit_array_2.drv<63:0>.n36 VSS 0.464f
C3003 hgu_cdac_8bit_array_2.drv<63:0>.n37 VSS 3.93f
C3004 hgu_cdac_8bit_array_2.drv<63:0>.n38 VSS -1.72f
C3005 hgu_cdac_8bit_array_2.drv<63:0>.n39 VSS -1.09f
C3006 hgu_cdac_8bit_array_2.drv<63:0>.n40 VSS -1.75f
C3007 hgu_cdac_8bit_array_2.drv<63:0>.n41 VSS -1.75f
C3008 hgu_cdac_8bit_array_2.drv<63:0>.n42 VSS -1.09f
C3009 hgu_cdac_8bit_array_2.drv<63:0>.n43 VSS -1.72f
C3010 hgu_cdac_8bit_array_2.drv<63:0>.n44 VSS 3.94f
C3011 hgu_cdac_8bit_array_2.drv<63:0>.n45 VSS 8.53f
C3012 hgu_cdac_8bit_array_2.drv<63:0>.n46 VSS -1.72f
C3013 hgu_cdac_8bit_array_2.drv<63:0>.n47 VSS -1.09f
C3014 hgu_cdac_8bit_array_2.drv<63:0>.n48 VSS -1.75f
C3015 hgu_cdac_8bit_array_2.drv<63:0>.n49 VSS -1.75f
C3016 hgu_cdac_8bit_array_2.drv<63:0>.n50 VSS -1.09f
C3017 hgu_cdac_8bit_array_2.drv<63:0>.n51 VSS -1.72f
C3018 hgu_cdac_8bit_array_2.drv<63:0>.n52 VSS 3.94f
C3019 hgu_cdac_8bit_array_2.drv<63:0>.n53 VSS 8.87f
C3020 hgu_cdac_8bit_array_2.drv<63:0>.n54 VSS -1.72f
C3021 hgu_cdac_8bit_array_2.drv<63:0>.n55 VSS -1.09f
C3022 hgu_cdac_8bit_array_2.drv<63:0>.n56 VSS -1.75f
C3023 hgu_cdac_8bit_array_2.drv<63:0>.n57 VSS -1.75f
C3024 hgu_cdac_8bit_array_2.drv<63:0>.n58 VSS -1.09f
C3025 hgu_cdac_8bit_array_2.drv<63:0>.n59 VSS -1.72f
C3026 hgu_cdac_8bit_array_2.drv<63:0>.n60 VSS 6.09f
C3027 hgu_cdac_8bit_array_2.drv<63:0>.n61 VSS -1.52f
C3028 hgu_cdac_8bit_array_2.drv<63:0>.n62 VSS -1.72f
C3029 hgu_cdac_8bit_array_2.drv<63:0>.n63 VSS 6.09f
C3030 hgu_cdac_8bit_array_2.drv<63:0>.n64 VSS 4.59f
C3031 hgu_cdac_8bit_array_2.drv<63:0>.n65 VSS 0.735f
C3032 hgu_cdac_8bit_array_2.drv<63:0>.n66 VSS -0.458f
C3033 hgu_cdac_8bit_array_2.drv<63:0>.n67 VSS -1.72f
C3034 hgu_cdac_8bit_array_2.drv<63:0>.n68 VSS 6.1f
C3035 hgu_cdac_8bit_array_2.drv<63:0>.n69 VSS -1.72f
C3036 hgu_cdac_8bit_array_2.drv<63:0>.n70 VSS -0.458f
C3037 hgu_cdac_8bit_array_2.drv<63:0>.n71 VSS 0.642f
C3038 hgu_cdac_8bit_array_2.drv<63:0>.n72 VSS 0.145f
C3039 hgu_cdac_8bit_array_2.drv<63:0>.n73 VSS 0.145f
C3040 hgu_cdac_8bit_array_2.drv<63:0>.n74 VSS 0.601f
C3041 hgu_cdac_8bit_array_2.drv<63:0>.n75 VSS -0.458f
C3042 hgu_cdac_8bit_array_2.drv<63:0>.n76 VSS -1.72f
C3043 hgu_cdac_8bit_array_2.drv<63:0>.n77 VSS 6.1f
C3044 hgu_cdac_8bit_array_2.drv<63:0>.n78 VSS -1.72f
C3045 hgu_cdac_8bit_array_2.drv<63:0>.n79 VSS -0.458f
C3046 hgu_cdac_8bit_array_2.drv<63:0>.n80 VSS 0.642f
C3047 hgu_cdac_8bit_array_2.drv<63:0>.n81 VSS 0.145f
C3048 hgu_cdac_8bit_array_2.drv<63:0>.n82 VSS 0.145f
C3049 hgu_cdac_8bit_array_2.drv<63:0>.n83 VSS 0.601f
C3050 hgu_cdac_8bit_array_2.drv<63:0>.n84 VSS -0.458f
C3051 hgu_cdac_8bit_array_2.drv<63:0>.n85 VSS -1.72f
C3052 hgu_cdac_8bit_array_2.drv<63:0>.n86 VSS 4.35f
C3053 hgu_cdac_8bit_array_2.drv<63:0>.n87 VSS -1.72f
C3054 hgu_cdac_8bit_array_2.drv<63:0>.n88 VSS -0.458f
C3055 hgu_cdac_8bit_array_2.drv<63:0>.n89 VSS 0.642f
C3056 hgu_cdac_8bit_array_2.drv<63:0>.n90 VSS 0.145f
C3057 hgu_cdac_8bit_array_2.drv<63:0>.n91 VSS 0.145f
C3058 hgu_cdac_8bit_array_2.drv<63:0>.n92 VSS 0.601f
C3059 hgu_cdac_8bit_array_2.drv<63:0>.n93 VSS -0.458f
C3060 hgu_cdac_8bit_array_2.drv<63:0>.n94 VSS -1.72f
C3061 hgu_cdac_8bit_array_2.drv<63:0>.n95 VSS 4.35f
C3062 hgu_cdac_8bit_array_2.drv<63:0>.n96 VSS -1.72f
C3063 hgu_cdac_8bit_array_2.drv<63:0>.n97 VSS -0.458f
C3064 hgu_cdac_8bit_array_2.drv<63:0>.n98 VSS 0.642f
C3065 hgu_cdac_8bit_array_2.drv<63:0>.n99 VSS 0.145f
C3066 hgu_cdac_8bit_array_2.drv<63:0>.n100 VSS 0.145f
C3067 hgu_cdac_8bit_array_2.drv<63:0>.n101 VSS 0.601f
C3068 hgu_cdac_8bit_array_2.drv<63:0>.n102 VSS -0.458f
C3069 hgu_cdac_8bit_array_2.drv<63:0>.n103 VSS -1.72f
C3070 hgu_cdac_8bit_array_2.drv<63:0>.n104 VSS 4.35f
C3071 hgu_cdac_8bit_array_2.drv<63:0>.n105 VSS -1.72f
C3072 hgu_cdac_8bit_array_2.drv<63:0>.n106 VSS -0.458f
C3073 hgu_cdac_8bit_array_2.drv<63:0>.n107 VSS 0.642f
C3074 hgu_cdac_8bit_array_2.drv<63:0>.n108 VSS 0.145f
C3075 hgu_cdac_8bit_array_2.drv<63:0>.n109 VSS 0.145f
C3076 hgu_cdac_8bit_array_2.drv<63:0>.n110 VSS 0.601f
C3077 hgu_cdac_8bit_array_2.drv<63:0>.n111 VSS -0.458f
C3078 hgu_cdac_8bit_array_2.drv<63:0>.n112 VSS -1.72f
C3079 hgu_cdac_8bit_array_2.drv<63:0>.n113 VSS 4.23f
C3080 hgu_cdac_8bit_array_2.drv<63:0>.t47 VSS 0.104f
C3081 hgu_cdac_8bit_array_2.drv<63:0>.t53 VSS 0.104f
C3082 hgu_cdac_8bit_array_2.drv<63:0>.n114 VSS 0.793f
C3083 hgu_cdac_8bit_array_2.drv<63:0>.t64 VSS 0.0521f
C3084 hgu_cdac_8bit_array_2.drv<63:0>.t70 VSS 0.0521f
C3085 hgu_cdac_8bit_array_2.drv<63:0>.n115 VSS 0.383f
C3086 hgu_cdac_8bit_array_2.drv<63:0>.n116 VSS 0.389f
C3087 hgu_cdac_8bit_array_2.drv<63:0>.t60 VSS 0.104f
C3088 hgu_cdac_8bit_array_2.drv<63:0>.t24 VSS 0.104f
C3089 hgu_cdac_8bit_array_2.drv<63:0>.n117 VSS 0.793f
C3090 hgu_cdac_8bit_array_2.drv<63:0>.t77 VSS 0.0521f
C3091 hgu_cdac_8bit_array_2.drv<63:0>.t105 VSS 0.0521f
C3092 hgu_cdac_8bit_array_2.drv<63:0>.n118 VSS 0.383f
C3093 hgu_cdac_8bit_array_2.drv<63:0>.n119 VSS 0.443f
C3094 hgu_cdac_8bit_array_2.drv<63:0>.n120 VSS 3.79f
C3095 hgu_cdac_8bit_array_2.drv<63:0>.n121 VSS -1.72f
C3096 hgu_cdac_8bit_array_2.drv<63:0>.n122 VSS -1.09f
C3097 hgu_cdac_8bit_array_2.drv<63:0>.n123 VSS -1.75f
C3098 hgu_cdac_8bit_array_2.drv<63:0>.n124 VSS -1.75f
C3099 hgu_cdac_8bit_array_2.drv<63:0>.n125 VSS -1.09f
C3100 hgu_cdac_8bit_array_2.drv<63:0>.n126 VSS -1.72f
C3101 hgu_cdac_8bit_array_2.drv<63:0>.n127 VSS 3.94f
C3102 hgu_cdac_8bit_array_2.drv<63:0>.n128 VSS 8.67f
C3103 hgu_cdac_8bit_array_2.drv<63:0>.t0 VSS 0.104f
C3104 hgu_cdac_8bit_array_2.drv<63:0>.t9 VSS 0.104f
C3105 hgu_cdac_8bit_array_2.drv<63:0>.n129 VSS 0.793f
C3106 hgu_cdac_8bit_array_2.drv<63:0>.t81 VSS 0.0521f
C3107 hgu_cdac_8bit_array_2.drv<63:0>.t90 VSS 0.0521f
C3108 hgu_cdac_8bit_array_2.drv<63:0>.n130 VSS 0.383f
C3109 hgu_cdac_8bit_array_2.drv<63:0>.n131 VSS 0.433f
C3110 hgu_cdac_8bit_array_2.drv<63:0>.t20 VSS 0.104f
C3111 hgu_cdac_8bit_array_2.drv<63:0>.t43 VSS 0.104f
C3112 hgu_cdac_8bit_array_2.drv<63:0>.n132 VSS 0.793f
C3113 hgu_cdac_8bit_array_2.drv<63:0>.t63 VSS 0.104f
C3114 hgu_cdac_8bit_array_2.drv<63:0>.t8 VSS 0.104f
C3115 hgu_cdac_8bit_array_2.drv<63:0>.n133 VSS 0.793f
C3116 hgu_cdac_8bit_array_2.drv<63:0>.t80 VSS 0.0521f
C3117 hgu_cdac_8bit_array_2.drv<63:0>.t89 VSS 0.0521f
C3118 hgu_cdac_8bit_array_2.drv<63:0>.n134 VSS 0.383f
C3119 hgu_cdac_8bit_array_2.drv<63:0>.n135 VSS 0.49f
C3120 hgu_cdac_8bit_array_2.drv<63:0>.t101 VSS 0.0521f
C3121 hgu_cdac_8bit_array_2.drv<63:0>.t124 VSS 0.0521f
C3122 hgu_cdac_8bit_array_2.drv<63:0>.n136 VSS 0.383f
C3123 hgu_cdac_8bit_array_2.drv<63:0>.n137 VSS 0.396f
C3124 hgu_cdac_8bit_array_2.drv<63:0>.n138 VSS 3.94f
C3125 hgu_cdac_8bit_array_2.drv<63:0>.n139 VSS -1.72f
C3126 hgu_cdac_8bit_array_2.drv<63:0>.n140 VSS -1.09f
C3127 hgu_cdac_8bit_array_2.drv<63:0>.n141 VSS -1.75f
C3128 hgu_cdac_8bit_array_2.drv<63:0>.n142 VSS -1.75f
C3129 hgu_cdac_8bit_array_2.drv<63:0>.n143 VSS -1.09f
C3130 hgu_cdac_8bit_array_2.drv<63:0>.n144 VSS -1.72f
C3131 hgu_cdac_8bit_array_2.drv<63:0>.n145 VSS 3.94f
C3132 hgu_cdac_8bit_array_2.drv<63:0>.n146 VSS 8.53f
C3133 hgu_cdac_8bit_array_2.drv<63:0>.t35 VSS 0.104f
C3134 hgu_cdac_8bit_array_2.drv<63:0>.t41 VSS 0.104f
C3135 hgu_cdac_8bit_array_2.drv<63:0>.n147 VSS 0.747f
C3136 hgu_cdac_8bit_array_2.drv<63:0>.t116 VSS 0.0521f
C3137 hgu_cdac_8bit_array_2.drv<63:0>.t122 VSS 0.0521f
C3138 hgu_cdac_8bit_array_2.drv<63:0>.n148 VSS 0.368f
C3139 hgu_cdac_8bit_array_2.drv<63:0>.t4 VSS 0.104f
C3140 hgu_cdac_8bit_array_2.drv<63:0>.t32 VSS 0.104f
C3141 hgu_cdac_8bit_array_2.drv<63:0>.n149 VSS 0.793f
C3142 hgu_cdac_8bit_array_2.drv<63:0>.t85 VSS 0.0521f
C3143 hgu_cdac_8bit_array_2.drv<63:0>.t113 VSS 0.0521f
C3144 hgu_cdac_8bit_array_2.drv<63:0>.n150 VSS 0.383f
C3145 hgu_cdac_8bit_array_2.drv<63:0>.n151 VSS 0.489f
C3146 hgu_cdac_8bit_array_2.drv<63:0>.n152 VSS -1.72f
C3147 hgu_cdac_8bit_array_2.drv<63:0>.n153 VSS -1.09f
C3148 hgu_cdac_8bit_array_2.drv<63:0>.n154 VSS -1.75f
C3149 hgu_cdac_8bit_array_2.drv<63:0>.n155 VSS -1.75f
C3150 hgu_cdac_8bit_array_2.drv<63:0>.n156 VSS -1.09f
C3151 hgu_cdac_8bit_array_2.drv<63:0>.n157 VSS -1.72f
C3152 hgu_cdac_8bit_array_2.drv<63:0>.n158 VSS 3.94f
C3153 hgu_cdac_8bit_array_2.drv<63:0>.n159 VSS 8.53f
C3154 hgu_cdac_8bit_array_2.drv<63:0>.t52 VSS 0.104f
C3155 hgu_cdac_8bit_array_2.drv<63:0>.t11 VSS 0.104f
C3156 hgu_cdac_8bit_array_2.drv<63:0>.n160 VSS 0.793f
C3157 hgu_cdac_8bit_array_2.drv<63:0>.t69 VSS 0.0521f
C3158 hgu_cdac_8bit_array_2.drv<63:0>.t92 VSS 0.0521f
C3159 hgu_cdac_8bit_array_2.drv<63:0>.n161 VSS 0.383f
C3160 hgu_cdac_8bit_array_2.drv<63:0>.n162 VSS 0.396f
C3161 hgu_cdac_8bit_array_2.drv<63:0>.t50 VSS 0.104f
C3162 hgu_cdac_8bit_array_2.drv<63:0>.t16 VSS 0.104f
C3163 hgu_cdac_8bit_array_2.drv<63:0>.n163 VSS 0.793f
C3164 hgu_cdac_8bit_array_2.drv<63:0>.t67 VSS 0.0521f
C3165 hgu_cdac_8bit_array_2.drv<63:0>.t97 VSS 0.0521f
C3166 hgu_cdac_8bit_array_2.drv<63:0>.n164 VSS 0.383f
C3167 hgu_cdac_8bit_array_2.drv<63:0>.n165 VSS 0.443f
C3168 hgu_cdac_8bit_array_2.drv<63:0>.t2 VSS 0.104f
C3169 hgu_cdac_8bit_array_2.drv<63:0>.t30 VSS 0.104f
C3170 hgu_cdac_8bit_array_2.drv<63:0>.n166 VSS 0.793f
C3171 hgu_cdac_8bit_array_2.drv<63:0>.t83 VSS 0.0521f
C3172 hgu_cdac_8bit_array_2.drv<63:0>.t111 VSS 0.0521f
C3173 hgu_cdac_8bit_array_2.drv<63:0>.n167 VSS 0.383f
C3174 hgu_cdac_8bit_array_2.drv<63:0>.n168 VSS 0.433f
C3175 hgu_cdac_8bit_array_2.drv<63:0>.n169 VSS 3.94f
C3176 hgu_cdac_8bit_array_2.drv<63:0>.n170 VSS -1.72f
C3177 hgu_cdac_8bit_array_2.drv<63:0>.n171 VSS -1.09f
C3178 hgu_cdac_8bit_array_2.drv<63:0>.n172 VSS -1.75f
C3179 hgu_cdac_8bit_array_2.drv<63:0>.n173 VSS -1.75f
C3180 hgu_cdac_8bit_array_2.drv<63:0>.n174 VSS -1.09f
C3181 hgu_cdac_8bit_array_2.drv<63:0>.n175 VSS -1.72f
C3182 hgu_cdac_8bit_array_2.drv<63:0>.n176 VSS 3.94f
C3183 hgu_cdac_8bit_array_2.drv<63:0>.n177 VSS 8.53f
C3184 hgu_cdac_8bit_array_2.drv<63:0>.t42 VSS 0.104f
C3185 hgu_cdac_8bit_array_2.drv<63:0>.t48 VSS 0.104f
C3186 hgu_cdac_8bit_array_2.drv<63:0>.n178 VSS 0.793f
C3187 hgu_cdac_8bit_array_2.drv<63:0>.t123 VSS 0.0521f
C3188 hgu_cdac_8bit_array_2.drv<63:0>.t65 VSS 0.0521f
C3189 hgu_cdac_8bit_array_2.drv<63:0>.n179 VSS 0.383f
C3190 hgu_cdac_8bit_array_2.drv<63:0>.n180 VSS 0.389f
C3191 hgu_cdac_8bit_array_2.drv<63:0>.n181 VSS 3.59f
C3192 hgu_cdac_8bit_array_2.drv<63:0>.n182 VSS -1.72f
C3193 hgu_cdac_8bit_array_2.drv<63:0>.n183 VSS -1.09f
C3194 hgu_cdac_8bit_array_2.drv<63:0>.n184 VSS -1.75f
C3195 hgu_cdac_8bit_array_2.drv<63:0>.n185 VSS -1.75f
C3196 hgu_cdac_8bit_array_2.drv<63:0>.n186 VSS -1.09f
C3197 hgu_cdac_8bit_array_2.drv<63:0>.n187 VSS -1.72f
C3198 hgu_cdac_8bit_array_2.drv<63:0>.n188 VSS 3.94f
C3199 hgu_cdac_8bit_array_2.drv<63:0>.n189 VSS 8.87f
C3200 hgu_cdac_8bit_array_2.drv<63:0>.t40 VSS 0.104f
C3201 hgu_cdac_8bit_array_2.drv<63:0>.t61 VSS 0.104f
C3202 hgu_cdac_8bit_array_2.drv<63:0>.n190 VSS 0.747f
C3203 hgu_cdac_8bit_array_2.drv<63:0>.t121 VSS 0.0521f
C3204 hgu_cdac_8bit_array_2.drv<63:0>.t78 VSS 0.0521f
C3205 hgu_cdac_8bit_array_2.drv<63:0>.n191 VSS 0.368f
C3206 hgu_cdac_8bit_array_2.drv<63:0>.t7 VSS 0.104f
C3207 hgu_cdac_8bit_array_2.drv<63:0>.t14 VSS 0.104f
C3208 hgu_cdac_8bit_array_2.drv<63:0>.n192 VSS 0.793f
C3209 hgu_cdac_8bit_array_2.drv<63:0>.t88 VSS 0.0521f
C3210 hgu_cdac_8bit_array_2.drv<63:0>.t95 VSS 0.0521f
C3211 hgu_cdac_8bit_array_2.drv<63:0>.n193 VSS 0.383f
C3212 hgu_cdac_8bit_array_2.drv<63:0>.n194 VSS 0.493f
C3213 hgu_cdac_8bit_array_2.drv<63:0>.n195 VSS 0.396f
C3214 hgu_cdac_8bit_array_2.drv<63:0>.t5 VSS 0.104f
C3215 hgu_cdac_8bit_array_2.drv<63:0>.t37 VSS 0.104f
C3216 hgu_cdac_8bit_array_2.drv<63:0>.n196 VSS 0.793f
C3217 hgu_cdac_8bit_array_2.drv<63:0>.t86 VSS 0.0521f
C3218 hgu_cdac_8bit_array_2.drv<63:0>.t118 VSS 0.0521f
C3219 hgu_cdac_8bit_array_2.drv<63:0>.n197 VSS 0.383f
C3220 hgu_cdac_8bit_array_2.drv<63:0>.n198 VSS 0.474f
C3221 hgu_cdac_8bit_array_2.drv<63:0>.n199 VSS 3.92f
C3222 hgu_cdac_8bit_array_2.drv<63:0>.n200 VSS -1.72f
C3223 hgu_cdac_8bit_array_2.drv<63:0>.n201 VSS -1.09f
C3224 hgu_cdac_8bit_array_2.drv<63:0>.n202 VSS -1.75f
C3225 hgu_cdac_8bit_array_2.drv<63:0>.n203 VSS -1.75f
C3226 hgu_cdac_8bit_array_2.drv<63:0>.n204 VSS -1.09f
C3227 hgu_cdac_8bit_array_2.drv<63:0>.n205 VSS -1.72f
C3228 hgu_cdac_8bit_array_2.drv<63:0>.n206 VSS 3.94f
C3229 hgu_cdac_8bit_array_2.drv<63:0>.n207 VSS 8.53f
C3230 hgu_cdac_8bit_array_2.drv<63:0>.t58 VSS 0.104f
C3231 hgu_cdac_8bit_array_2.drv<63:0>.t21 VSS 0.104f
C3232 hgu_cdac_8bit_array_2.drv<63:0>.n208 VSS 0.793f
C3233 hgu_cdac_8bit_array_2.drv<63:0>.t75 VSS 0.0521f
C3234 hgu_cdac_8bit_array_2.drv<63:0>.t102 VSS 0.0521f
C3235 hgu_cdac_8bit_array_2.drv<63:0>.n209 VSS 0.383f
C3236 hgu_cdac_8bit_array_2.drv<63:0>.n210 VSS 0.41f
C3237 hgu_cdac_8bit_array_2.drv<63:0>.t29 VSS 0.104f
C3238 hgu_cdac_8bit_array_2.drv<63:0>.t36 VSS 0.104f
C3239 hgu_cdac_8bit_array_2.drv<63:0>.n211 VSS 0.793f
C3240 hgu_cdac_8bit_array_2.drv<63:0>.t110 VSS 0.0521f
C3241 hgu_cdac_8bit_array_2.drv<63:0>.t117 VSS 0.0521f
C3242 hgu_cdac_8bit_array_2.drv<63:0>.n212 VSS 0.383f
C3243 hgu_cdac_8bit_array_2.drv<63:0>.n213 VSS 0.418f
C3244 hgu_cdac_8bit_array_2.drv<63:0>.n214 VSS 3.94f
C3245 hgu_cdac_8bit_array_2.drv<63:0>.n215 VSS -1.72f
C3246 hgu_cdac_8bit_array_2.drv<63:0>.n216 VSS -1.09f
C3247 hgu_cdac_8bit_array_2.drv<63:0>.n217 VSS -1.75f
C3248 hgu_cdac_8bit_array_2.drv<63:0>.n218 VSS -1.75f
C3249 hgu_cdac_8bit_array_2.drv<63:0>.n219 VSS -1.09f
C3250 hgu_cdac_8bit_array_2.drv<63:0>.n220 VSS -1.72f
C3251 hgu_cdac_8bit_array_2.drv<63:0>.n221 VSS 3.94f
C3252 hgu_cdac_8bit_array_2.drv<63:0>.n222 VSS 8.53f
C3253 hgu_cdac_8bit_array_2.drv<63:0>.t56 VSS 0.104f
C3254 hgu_cdac_8bit_array_2.drv<63:0>.t17 VSS 0.104f
C3255 hgu_cdac_8bit_array_2.drv<63:0>.n223 VSS 0.793f
C3256 hgu_cdac_8bit_array_2.drv<63:0>.t73 VSS 0.0521f
C3257 hgu_cdac_8bit_array_2.drv<63:0>.t98 VSS 0.0521f
C3258 hgu_cdac_8bit_array_2.drv<63:0>.n224 VSS 0.383f
C3259 hgu_cdac_8bit_array_2.drv<63:0>.n225 VSS 0.465f
C3260 hgu_cdac_8bit_array_2.drv<63:0>.t26 VSS 0.104f
C3261 hgu_cdac_8bit_array_2.drv<63:0>.t6 VSS 0.104f
C3262 hgu_cdac_8bit_array_2.drv<63:0>.n226 VSS 0.747f
C3263 hgu_cdac_8bit_array_2.drv<63:0>.t108 VSS 0.0521f
C3264 hgu_cdac_8bit_array_2.drv<63:0>.t87 VSS 0.0521f
C3265 hgu_cdac_8bit_array_2.drv<63:0>.n227 VSS 0.368f
C3266 hgu_cdac_8bit_array_2.drv<63:0>.t12 VSS 0.104f
C3267 hgu_cdac_8bit_array_2.drv<63:0>.t23 VSS 0.104f
C3268 hgu_cdac_8bit_array_2.drv<63:0>.n228 VSS 0.793f
C3269 hgu_cdac_8bit_array_2.drv<63:0>.t93 VSS 0.0521f
C3270 hgu_cdac_8bit_array_2.drv<63:0>.t104 VSS 0.0521f
C3271 hgu_cdac_8bit_array_2.drv<63:0>.n229 VSS 0.383f
C3272 hgu_cdac_8bit_array_2.drv<63:0>.n230 VSS 0.499f
C3273 hgu_cdac_8bit_array_2.drv<63:0>.n231 VSS 0.416f
C3274 hgu_cdac_8bit_array_2.drv<63:0>.n232 VSS 3.93f
C3275 hgu_cdac_8bit_array_2.drv<63:0>.n233 VSS -1.72f
C3276 hgu_cdac_8bit_array_2.drv<63:0>.n234 VSS -1.09f
C3277 hgu_cdac_8bit_array_2.drv<63:0>.n235 VSS -1.75f
C3278 hgu_cdac_8bit_array_2.drv<63:0>.n236 VSS -1.75f
C3279 hgu_cdac_8bit_array_2.drv<63:0>.n237 VSS -1.09f
C3280 hgu_cdac_8bit_array_2.drv<63:0>.n238 VSS -1.72f
C3281 hgu_cdac_8bit_array_2.drv<63:0>.n239 VSS 3.94f
C3282 hgu_cdac_8bit_array_2.drv<63:0>.n240 VSS 8.53f
C3283 hgu_cdac_8bit_array_2.drv<63:0>.t46 VSS 0.104f
C3284 hgu_cdac_8bit_array_2.drv<63:0>.t3 VSS 0.104f
C3285 hgu_cdac_8bit_array_2.drv<63:0>.n241 VSS 0.747f
C3286 hgu_cdac_8bit_array_2.drv<63:0>.t127 VSS 0.0521f
C3287 hgu_cdac_8bit_array_2.drv<63:0>.t84 VSS 0.0521f
C3288 hgu_cdac_8bit_array_2.drv<63:0>.n242 VSS 0.368f
C3289 hgu_cdac_8bit_array_2.drv<63:0>.n243 VSS 0.427f
C3290 hgu_cdac_8bit_array_2.drv<63:0>.t31 VSS 0.104f
C3291 hgu_cdac_8bit_array_2.drv<63:0>.t22 VSS 0.104f
C3292 hgu_cdac_8bit_array_2.drv<63:0>.n244 VSS 0.793f
C3293 hgu_cdac_8bit_array_2.drv<63:0>.t112 VSS 0.0521f
C3294 hgu_cdac_8bit_array_2.drv<63:0>.t103 VSS 0.0521f
C3295 hgu_cdac_8bit_array_2.drv<63:0>.n245 VSS 0.383f
C3296 hgu_cdac_8bit_array_2.drv<63:0>.n246 VSS 0.46f
C3297 hgu_cdac_8bit_array_2.drv<63:0>.n247 VSS 3.93f
C3298 hgu_cdac_8bit_array_2.drv<63:0>.n248 VSS -1.72f
C3299 hgu_cdac_8bit_array_2.drv<63:0>.n249 VSS -1.09f
C3300 hgu_cdac_8bit_array_2.drv<63:0>.n250 VSS -1.75f
C3301 hgu_cdac_8bit_array_2.drv<63:0>.n251 VSS -1.75f
C3302 hgu_cdac_8bit_array_2.drv<63:0>.n252 VSS -1.09f
C3303 hgu_cdac_8bit_array_2.drv<63:0>.n253 VSS -1.72f
C3304 hgu_cdac_8bit_array_2.drv<63:0>.n254 VSS 3.94f
C3305 hgu_cdac_8bit_array_2.drv<63:0>.n255 VSS 8.53f
C3306 hgu_cdac_8bit_array_2.drv<63:0>.t44 VSS 0.104f
C3307 hgu_cdac_8bit_array_2.drv<63:0>.t18 VSS 0.104f
C3308 hgu_cdac_8bit_array_2.drv<63:0>.n256 VSS 0.793f
C3309 hgu_cdac_8bit_array_2.drv<63:0>.t125 VSS 0.0521f
C3310 hgu_cdac_8bit_array_2.drv<63:0>.t99 VSS 0.0521f
C3311 hgu_cdac_8bit_array_2.drv<63:0>.n257 VSS 0.383f
C3312 hgu_cdac_8bit_array_2.drv<63:0>.n258 VSS 0.424f
C3313 hgu_cdac_8bit_array_2.drv<63:0>.t28 VSS 0.104f
C3314 hgu_cdac_8bit_array_2.drv<63:0>.t49 VSS 0.104f
C3315 hgu_cdac_8bit_array_2.drv<63:0>.n259 VSS 0.793f
C3316 hgu_cdac_8bit_array_2.drv<63:0>.t109 VSS 0.0521f
C3317 hgu_cdac_8bit_array_2.drv<63:0>.t66 VSS 0.0521f
C3318 hgu_cdac_8bit_array_2.drv<63:0>.n260 VSS 0.383f
C3319 hgu_cdac_8bit_array_2.drv<63:0>.n261 VSS 0.404f
C3320 hgu_cdac_8bit_array_2.drv<63:0>.n262 VSS 3.94f
C3321 hgu_cdac_8bit_array_2.drv<63:0>.n263 VSS -1.72f
C3322 hgu_cdac_8bit_array_2.drv<63:0>.n264 VSS -1.09f
C3323 hgu_cdac_8bit_array_2.drv<63:0>.n265 VSS -1.75f
C3324 hgu_cdac_8bit_array_2.drv<63:0>.n266 VSS -1.75f
C3325 hgu_cdac_8bit_array_2.drv<63:0>.n267 VSS -1.09f
C3326 hgu_cdac_8bit_array_2.drv<63:0>.n268 VSS -1.72f
C3327 hgu_cdac_8bit_array_2.drv<63:0>.n269 VSS 3.94f
C3328 hgu_cdac_8bit_array_2.drv<63:0>.n270 VSS 8.53f
C3329 hgu_cdac_8bit_array_2.drv<63:0>.t54 VSS 0.104f
C3330 hgu_cdac_8bit_array_2.drv<63:0>.t15 VSS 0.104f
C3331 hgu_cdac_8bit_array_2.drv<63:0>.n271 VSS 0.792f
C3332 hgu_cdac_8bit_array_2.drv<63:0>.t71 VSS 0.0521f
C3333 hgu_cdac_8bit_array_2.drv<63:0>.t96 VSS 0.0521f
C3334 hgu_cdac_8bit_array_2.drv<63:0>.n272 VSS 0.344f
C3335 hgu_cdac_8bit_array_2.drv<63:0>.n273 VSS -1.72f
C3336 hgu_cdac_8bit_array_2.drv<63:0>.n274 VSS -1.09f
C3337 hgu_cdac_8bit_array_2.drv<63:0>.n275 VSS -1.75f
C3338 hgu_cdac_8bit_array_2.drv<63:0>.n276 VSS -1.75f
C3339 hgu_cdac_8bit_array_2.drv<63:0>.n277 VSS -1.09f
C3340 hgu_cdac_8bit_array_2.drv<63:0>.n278 VSS -1.72f
C3341 hgu_cdac_8bit_array_2.drv<63:0>.n279 VSS 3.94f
C3342 hgu_cdac_8bit_array_2.drv<63:0>.n280 VSS 8.79f
C3343 hgu_cdac_8bit_array_2.drv<63:0>.n281 VSS -1.72f
C3344 hgu_cdac_8bit_array_2.drv<63:0>.n282 VSS -1.09f
C3345 hgu_cdac_8bit_array_2.drv<63:0>.n283 VSS -1.75f
C3346 hgu_cdac_8bit_array_2.drv<63:0>.n284 VSS -1.75f
C3347 hgu_cdac_8bit_array_2.drv<63:0>.n285 VSS -1.09f
C3348 hgu_cdac_8bit_array_2.drv<63:0>.n286 VSS -1.72f
C3349 hgu_cdac_8bit_array_2.drv<63:0>.n287 VSS 6.09f
C3350 hgu_cdac_8bit_array_2.drv<63:0>.n288 VSS -1.72f
C3351 hgu_cdac_8bit_array_2.drv<63:0>.n289 VSS -1.09f
C3352 hgu_cdac_8bit_array_2.drv<63:0>.n290 VSS -1.75f
C3353 hgu_cdac_8bit_array_2.drv<63:0>.n291 VSS -1.75f
C3354 hgu_cdac_8bit_array_2.drv<63:0>.n292 VSS -1.09f
C3355 hgu_cdac_8bit_array_2.drv<63:0>.n293 VSS -1.72f
C3356 hgu_cdac_8bit_array_2.drv<63:0>.n294 VSS 6.09f
C3357 hgu_cdac_8bit_array_2.drv<63:0>.n295 VSS -1.72f
C3358 hgu_cdac_8bit_array_2.drv<63:0>.n296 VSS -1.09f
C3359 hgu_cdac_8bit_array_2.drv<63:0>.n297 VSS -1.75f
C3360 hgu_cdac_8bit_array_2.drv<63:0>.n298 VSS -1.75f
C3361 hgu_cdac_8bit_array_2.drv<63:0>.n299 VSS -1.09f
C3362 hgu_cdac_8bit_array_2.drv<63:0>.n300 VSS -1.72f
C3363 hgu_cdac_8bit_array_2.drv<63:0>.n301 VSS 6.09f
C3364 hgu_cdac_8bit_array_2.drv<63:0>.n302 VSS -1.72f
C3365 hgu_cdac_8bit_array_2.drv<63:0>.n303 VSS -1.09f
C3366 hgu_cdac_8bit_array_2.drv<63:0>.n304 VSS -1.75f
C3367 hgu_cdac_8bit_array_2.drv<63:0>.n305 VSS -1.75f
C3368 hgu_cdac_8bit_array_2.drv<63:0>.n306 VSS -1.09f
C3369 hgu_cdac_8bit_array_2.drv<63:0>.n307 VSS -1.72f
C3370 hgu_cdac_8bit_array_2.drv<63:0>.n308 VSS 6.09f
C3371 hgu_cdac_8bit_array_2.drv<63:0>.n309 VSS -1.72f
C3372 hgu_cdac_8bit_array_2.drv<63:0>.n310 VSS -1.09f
C3373 hgu_cdac_8bit_array_2.drv<63:0>.n311 VSS -1.75f
C3374 hgu_cdac_8bit_array_2.drv<63:0>.n312 VSS -1.75f
C3375 hgu_cdac_8bit_array_2.drv<63:0>.n313 VSS -1.09f
C3376 hgu_cdac_8bit_array_2.drv<63:0>.n314 VSS -1.72f
C3377 hgu_cdac_8bit_array_2.drv<63:0>.n315 VSS 6.09f
C3378 hgu_cdac_8bit_array_2.drv<63:0>.n316 VSS -1.72f
C3379 hgu_cdac_8bit_array_2.drv<63:0>.n317 VSS -1.09f
C3380 hgu_cdac_8bit_array_2.drv<63:0>.n318 VSS -1.75f
C3381 hgu_cdac_8bit_array_2.drv<63:0>.n319 VSS -1.75f
C3382 hgu_cdac_8bit_array_2.drv<63:0>.n320 VSS -1.09f
C3383 hgu_cdac_8bit_array_2.drv<63:0>.n321 VSS -1.72f
C3384 hgu_cdac_8bit_array_2.drv<63:0>.n322 VSS 6.09f
C3385 hgu_cdac_8bit_array_2.drv<63:0>.n323 VSS -1.72f
C3386 hgu_cdac_8bit_array_2.drv<63:0>.n324 VSS -1.09f
C3387 hgu_cdac_8bit_array_2.drv<63:0>.n325 VSS -1.75f
C3388 hgu_cdac_8bit_array_2.drv<63:0>.n326 VSS -1.75f
C3389 hgu_cdac_8bit_array_2.drv<63:0>.n327 VSS -1.09f
C3390 hgu_cdac_8bit_array_2.drv<63:0>.n328 VSS -1.72f
C3391 hgu_cdac_8bit_array_2.drv<63:0>.n329 VSS 6.09f
C3392 hgu_cdac_8bit_array_2.drv<63:0>.n330 VSS -1.72f
C3393 hgu_cdac_8bit_array_2.drv<63:0>.n331 VSS -1.09f
C3394 hgu_cdac_8bit_array_2.drv<63:0>.n332 VSS -1.75f
C3395 hgu_cdac_8bit_array_2.drv<63:0>.n333 VSS -1.75f
C3396 hgu_cdac_8bit_array_2.drv<63:0>.n334 VSS -1.09f
C3397 hgu_cdac_8bit_array_2.drv<63:0>.n335 VSS -1.72f
C3398 hgu_cdac_8bit_array_2.drv<63:0>.n336 VSS 6.09f
C3399 hgu_cdac_8bit_array_2.drv<63:0>.n337 VSS -1.72f
C3400 hgu_cdac_8bit_array_2.drv<63:0>.n338 VSS -1.09f
C3401 hgu_cdac_8bit_array_2.drv<63:0>.n339 VSS -1.75f
C3402 hgu_cdac_8bit_array_2.drv<63:0>.n340 VSS -1.75f
C3403 hgu_cdac_8bit_array_2.drv<63:0>.n341 VSS -1.09f
C3404 hgu_cdac_8bit_array_2.drv<63:0>.n342 VSS -1.72f
C3405 hgu_cdac_8bit_array_2.drv<63:0>.n343 VSS 6.09f
C3406 hgu_cdac_8bit_array_2.drv<63:0>.n344 VSS -1.72f
C3407 hgu_cdac_8bit_array_2.drv<63:0>.n345 VSS -1.09f
C3408 hgu_cdac_8bit_array_2.drv<63:0>.n346 VSS -1.75f
C3409 hgu_cdac_8bit_array_2.drv<63:0>.n347 VSS -1.75f
C3410 hgu_cdac_8bit_array_2.drv<63:0>.n348 VSS -1.09f
C3411 hgu_cdac_8bit_array_2.drv<63:0>.n349 VSS -1.72f
C3412 hgu_cdac_8bit_array_2.drv<63:0>.n350 VSS 6.09f
C3413 hgu_cdac_8bit_array_2.drv<63:0>.n351 VSS -1.72f
C3414 hgu_cdac_8bit_array_2.drv<63:0>.n352 VSS -1.09f
C3415 hgu_cdac_8bit_array_2.drv<63:0>.n353 VSS -1.75f
C3416 hgu_cdac_8bit_array_2.drv<63:0>.n354 VSS -1.75f
C3417 hgu_cdac_8bit_array_2.drv<63:0>.n355 VSS -1.09f
C3418 hgu_cdac_8bit_array_2.drv<63:0>.n356 VSS -1.72f
C3419 hgu_cdac_8bit_array_2.drv<63:0>.n357 VSS 6.09f
C3420 hgu_cdac_8bit_array_2.drv<63:0>.n358 VSS -1.72f
C3421 hgu_cdac_8bit_array_2.drv<63:0>.n359 VSS -1.09f
C3422 hgu_cdac_8bit_array_2.drv<63:0>.n360 VSS -1.75f
C3423 hgu_cdac_8bit_array_2.drv<63:0>.n361 VSS -1.75f
C3424 hgu_cdac_8bit_array_2.drv<63:0>.n362 VSS -1.09f
C3425 hgu_cdac_8bit_array_2.drv<63:0>.n363 VSS -1.72f
C3426 hgu_cdac_8bit_array_2.drv<63:0>.n364 VSS 6.09f
C3427 hgu_cdac_8bit_array_2.drv<63:0>.n365 VSS -1.72f
C3428 hgu_cdac_8bit_array_2.drv<63:0>.n366 VSS -1.09f
C3429 hgu_cdac_8bit_array_2.drv<63:0>.n367 VSS -1.75f
C3430 hgu_cdac_8bit_array_2.drv<63:0>.n368 VSS -1.75f
C3431 hgu_cdac_8bit_array_2.drv<63:0>.n369 VSS -1.09f
C3432 hgu_cdac_8bit_array_2.drv<63:0>.n370 VSS -1.72f
C3433 hgu_cdac_8bit_array_2.drv<63:0>.n371 VSS 6.09f
C3434 hgu_cdac_8bit_array_2.drv<63:0>.n372 VSS -1.52f
C3435 hgu_cdac_8bit_array_2.drv<63:0>.n373 VSS -1.72f
C3436 hgu_cdac_8bit_array_2.drv<63:0>.n374 VSS 6.09f
C3437 hgu_cdac_8bit_array_2.drv<63:0>.n375 VSS 4.53f
C3438 hgu_cdac_8bit_array_2.drv<63:0>.n376 VSS 0.776f
C3439 hgu_cdac_8bit_array_2.drv<63:0>.n377 VSS -0.458f
C3440 hgu_cdac_8bit_array_2.drv<63:0>.n378 VSS -1.72f
C3441 hgu_cdac_8bit_array_2.drv<63:0>.n379 VSS 6.1f
C3442 hgu_cdac_8bit_array_2.drv<63:0>.n380 VSS -1.72f
C3443 hgu_cdac_8bit_array_2.drv<63:0>.n381 VSS -0.458f
C3444 hgu_cdac_8bit_array_2.drv<63:0>.n382 VSS 0.601f
C3445 hgu_cdac_8bit_array_2.drv<63:0>.n383 VSS 0.145f
C3446 hgu_cdac_8bit_array_2.drv<63:0>.n384 VSS 0.145f
C3447 hgu_cdac_8bit_array_2.drv<63:0>.n385 VSS 0.642f
C3448 hgu_cdac_8bit_array_2.drv<63:0>.n386 VSS -0.458f
C3449 hgu_cdac_8bit_array_2.drv<63:0>.n387 VSS -1.72f
C3450 hgu_cdac_8bit_array_2.drv<63:0>.n388 VSS 6.1f
C3451 hgu_cdac_8bit_array_2.drv<63:0>.n389 VSS -1.72f
C3452 hgu_cdac_8bit_array_2.drv<63:0>.n390 VSS -0.458f
C3453 hgu_cdac_8bit_array_2.drv<63:0>.n391 VSS 0.601f
C3454 hgu_cdac_8bit_array_2.drv<63:0>.n392 VSS 0.145f
C3455 hgu_cdac_8bit_array_2.drv<63:0>.n393 VSS 0.145f
C3456 hgu_cdac_8bit_array_2.drv<63:0>.n394 VSS 0.642f
C3457 hgu_cdac_8bit_array_2.drv<63:0>.n395 VSS -0.458f
C3458 hgu_cdac_8bit_array_2.drv<63:0>.n396 VSS -1.72f
C3459 hgu_cdac_8bit_array_2.drv<63:0>.n397 VSS 6.1f
C3460 hgu_cdac_8bit_array_2.drv<63:0>.n398 VSS -1.72f
C3461 hgu_cdac_8bit_array_2.drv<63:0>.n399 VSS -0.458f
C3462 hgu_cdac_8bit_array_2.drv<63:0>.n400 VSS 0.601f
C3463 hgu_cdac_8bit_array_2.drv<63:0>.n401 VSS 0.145f
C3464 hgu_cdac_8bit_array_2.drv<63:0>.n402 VSS 0.145f
C3465 hgu_cdac_8bit_array_2.drv<63:0>.n403 VSS 0.642f
C3466 hgu_cdac_8bit_array_2.drv<63:0>.n404 VSS -0.458f
C3467 hgu_cdac_8bit_array_2.drv<63:0>.n405 VSS -1.72f
C3468 hgu_cdac_8bit_array_2.drv<63:0>.n406 VSS 6.1f
C3469 hgu_cdac_8bit_array_2.drv<63:0>.n407 VSS -1.72f
C3470 hgu_cdac_8bit_array_2.drv<63:0>.n408 VSS -0.458f
C3471 hgu_cdac_8bit_array_2.drv<63:0>.n409 VSS 0.601f
C3472 hgu_cdac_8bit_array_2.drv<63:0>.n410 VSS 0.145f
C3473 hgu_cdac_8bit_array_2.drv<63:0>.n411 VSS 0.145f
C3474 hgu_cdac_8bit_array_2.drv<63:0>.n412 VSS 0.642f
C3475 hgu_cdac_8bit_array_2.drv<63:0>.n413 VSS -0.458f
C3476 hgu_cdac_8bit_array_2.drv<63:0>.n414 VSS -1.72f
C3477 hgu_cdac_8bit_array_2.drv<63:0>.n415 VSS 6.1f
C3478 hgu_cdac_8bit_array_2.drv<63:0>.n416 VSS -1.72f
C3479 hgu_cdac_8bit_array_2.drv<63:0>.n417 VSS -0.458f
C3480 hgu_cdac_8bit_array_2.drv<63:0>.n418 VSS 0.601f
C3481 hgu_cdac_8bit_array_2.drv<63:0>.n419 VSS 0.145f
C3482 hgu_cdac_8bit_array_2.drv<63:0>.n420 VSS 0.145f
C3483 hgu_cdac_8bit_array_2.drv<63:0>.n421 VSS 0.642f
C3484 hgu_cdac_8bit_array_2.drv<63:0>.n422 VSS -0.458f
C3485 hgu_cdac_8bit_array_2.drv<63:0>.n423 VSS -1.72f
C3486 hgu_cdac_8bit_array_2.drv<63:0>.n424 VSS 6.1f
C3487 hgu_cdac_8bit_array_2.drv<63:0>.n425 VSS -1.72f
C3488 hgu_cdac_8bit_array_2.drv<63:0>.n426 VSS -0.458f
C3489 hgu_cdac_8bit_array_2.drv<63:0>.n427 VSS 0.601f
C3490 hgu_cdac_8bit_array_2.drv<63:0>.n428 VSS 0.145f
C3491 hgu_cdac_8bit_array_2.drv<63:0>.n429 VSS 0.145f
C3492 hgu_cdac_8bit_array_2.drv<63:0>.n430 VSS 0.642f
C3493 hgu_cdac_8bit_array_2.drv<63:0>.n431 VSS -0.458f
C3494 hgu_cdac_8bit_array_2.drv<63:0>.n432 VSS -1.72f
C3495 hgu_cdac_8bit_array_2.drv<63:0>.n433 VSS 6.1f
C3496 hgu_cdac_8bit_array_2.drv<63:0>.n434 VSS -1.72f
C3497 hgu_cdac_8bit_array_2.drv<63:0>.n435 VSS -0.458f
C3498 hgu_cdac_8bit_array_2.drv<63:0>.n436 VSS 0.601f
C3499 hgu_cdac_8bit_array_2.drv<63:0>.n437 VSS 0.145f
C3500 hgu_cdac_8bit_array_2.drv<63:0>.n438 VSS 0.145f
C3501 hgu_cdac_8bit_array_2.drv<63:0>.n439 VSS 0.642f
C3502 hgu_cdac_8bit_array_2.drv<63:0>.n440 VSS -0.458f
C3503 hgu_cdac_8bit_array_2.drv<63:0>.n441 VSS -1.72f
C3504 hgu_cdac_8bit_array_2.drv<63:0>.n442 VSS 6.1f
C3505 hgu_cdac_8bit_array_2.drv<63:0>.n443 VSS -1.72f
C3506 hgu_cdac_8bit_array_2.drv<63:0>.n444 VSS -0.458f
C3507 hgu_cdac_8bit_array_2.drv<63:0>.n445 VSS 0.601f
C3508 hgu_cdac_8bit_array_2.drv<63:0>.n446 VSS 0.145f
C3509 hgu_cdac_8bit_array_2.drv<63:0>.n447 VSS 0.145f
C3510 hgu_cdac_8bit_array_2.drv<63:0>.n448 VSS 0.642f
C3511 hgu_cdac_8bit_array_2.drv<63:0>.n449 VSS -0.458f
C3512 hgu_cdac_8bit_array_2.drv<63:0>.n450 VSS -1.72f
C3513 hgu_cdac_8bit_array_2.drv<63:0>.n451 VSS 6.1f
C3514 hgu_cdac_8bit_array_2.drv<63:0>.n452 VSS -1.72f
C3515 hgu_cdac_8bit_array_2.drv<63:0>.n453 VSS -0.458f
C3516 hgu_cdac_8bit_array_2.drv<63:0>.n454 VSS 0.601f
C3517 hgu_cdac_8bit_array_2.drv<63:0>.n455 VSS 0.145f
C3518 hgu_cdac_8bit_array_2.drv<63:0>.n456 VSS 0.145f
C3519 hgu_cdac_8bit_array_2.drv<63:0>.n457 VSS 0.642f
C3520 hgu_cdac_8bit_array_2.drv<63:0>.n458 VSS -0.458f
C3521 hgu_cdac_8bit_array_2.drv<63:0>.n459 VSS -1.72f
C3522 hgu_cdac_8bit_array_2.drv<63:0>.n460 VSS 6.1f
C3523 hgu_cdac_8bit_array_2.drv<63:0>.n461 VSS -1.72f
C3524 hgu_cdac_8bit_array_2.drv<63:0>.n462 VSS -0.458f
C3525 hgu_cdac_8bit_array_2.drv<63:0>.n463 VSS 0.601f
C3526 hgu_cdac_8bit_array_2.drv<63:0>.n464 VSS 0.145f
C3527 hgu_cdac_8bit_array_2.drv<63:0>.n465 VSS 0.145f
C3528 hgu_cdac_8bit_array_2.drv<63:0>.n466 VSS 0.642f
C3529 hgu_cdac_8bit_array_2.drv<63:0>.n467 VSS -0.458f
C3530 hgu_cdac_8bit_array_2.drv<63:0>.n468 VSS -1.72f
C3531 hgu_cdac_8bit_array_2.drv<63:0>.n469 VSS 6.1f
C3532 hgu_cdac_8bit_array_2.drv<63:0>.n470 VSS -1.72f
C3533 hgu_cdac_8bit_array_2.drv<63:0>.n471 VSS -0.458f
C3534 hgu_cdac_8bit_array_2.drv<63:0>.n472 VSS 0.601f
C3535 hgu_cdac_8bit_array_2.drv<63:0>.n473 VSS 0.145f
C3536 hgu_cdac_8bit_array_2.drv<63:0>.n474 VSS 0.145f
C3537 hgu_cdac_8bit_array_2.drv<63:0>.n475 VSS 0.642f
C3538 hgu_cdac_8bit_array_2.drv<63:0>.n476 VSS -0.458f
C3539 hgu_cdac_8bit_array_2.drv<63:0>.n477 VSS -1.72f
C3540 hgu_cdac_8bit_array_2.drv<63:0>.n478 VSS 6.1f
C3541 hgu_cdac_8bit_array_2.drv<63:0>.n479 VSS -1.72f
C3542 hgu_cdac_8bit_array_2.drv<63:0>.n480 VSS -0.458f
C3543 hgu_cdac_8bit_array_2.drv<63:0>.n481 VSS 0.601f
C3544 hgu_cdac_8bit_array_2.drv<63:0>.n482 VSS 0.145f
C3545 hgu_cdac_8bit_array_2.drv<63:0>.n483 VSS 0.145f
C3546 hgu_cdac_8bit_array_2.drv<63:0>.n484 VSS 0.642f
C3547 hgu_cdac_8bit_array_2.drv<63:0>.n485 VSS -0.458f
C3548 hgu_cdac_8bit_array_2.drv<63:0>.n486 VSS -1.72f
C3549 hgu_cdac_8bit_array_2.drv<63:0>.n487 VSS 6.1f
C3550 hgu_cdac_8bit_array_2.drv<63:0>.n488 VSS -1.72f
C3551 hgu_cdac_8bit_array_2.drv<63:0>.n489 VSS -0.458f
C3552 hgu_cdac_8bit_array_2.drv<63:0>.n490 VSS 0.601f
C3553 hgu_cdac_8bit_array_2.drv<63:0>.n491 VSS 0.145f
C3554 hgu_cdac_8bit_array_2.drv<63:0>.n492 VSS 0.145f
C3555 hgu_cdac_8bit_array_2.drv<63:0>.n493 VSS 0.642f
C3556 hgu_cdac_8bit_array_2.drv<63:0>.n494 VSS -0.458f
C3557 hgu_cdac_8bit_array_2.drv<63:0>.n495 VSS -1.72f
C3558 hgu_cdac_8bit_array_2.drv<63:0>.n496 VSS 6.1f
C3559 hgu_cdac_8bit_array_2.drv<63:0>.n497 VSS -1.72f
C3560 hgu_cdac_8bit_array_2.drv<63:0>.n498 VSS -0.458f
C3561 hgu_cdac_8bit_array_2.drv<63:0>.n499 VSS 0.601f
C3562 hgu_cdac_8bit_array_2.drv<63:0>.n500 VSS 0.145f
C3563 hgu_cdac_8bit_array_2.drv<63:0>.n501 VSS 0.145f
C3564 hgu_cdac_8bit_array_2.drv<63:0>.n502 VSS 0.642f
C3565 hgu_cdac_8bit_array_2.drv<63:0>.n503 VSS 0.174f
C3566 hgu_cdac_8bit_array_2.drv<63:0>.n504 VSS 0.229f
C3567 hgu_cdac_8bit_array_2.drv<63:0>.n505 VSS 0.179f
C3568 hgu_cdac_8bit_array_2.drv<63:0>.n506 VSS 4.35f
C3569 hgu_cdac_8bit_array_2.drv<63:0>.n507 VSS -1.72f
C3570 hgu_cdac_8bit_array_2.drv<63:0>.n508 VSS -0.458f
C3571 hgu_cdac_8bit_array_2.drv<63:0>.n509 VSS 0.601f
C3572 hgu_cdac_8bit_array_2.drv<63:0>.n510 VSS 0.145f
C3573 hgu_cdac_8bit_array_2.drv<63:0>.n511 VSS 0.145f
C3574 hgu_cdac_8bit_array_2.drv<63:0>.n512 VSS 0.642f
C3575 hgu_cdac_8bit_array_2.drv<63:0>.n513 VSS -0.458f
C3576 hgu_cdac_8bit_array_2.drv<63:0>.n514 VSS -1.72f
C3577 hgu_cdac_8bit_array_2.drv<63:0>.n515 VSS 4.35f
C3578 hgu_cdac_8bit_array_2.drv<63:0>.n516 VSS -1.72f
C3579 hgu_cdac_8bit_array_2.drv<63:0>.n517 VSS -0.458f
C3580 hgu_cdac_8bit_array_2.drv<63:0>.n518 VSS 0.601f
C3581 hgu_cdac_8bit_array_2.drv<63:0>.n519 VSS 0.145f
C3582 hgu_cdac_8bit_array_2.drv<63:0>.n520 VSS 0.145f
C3583 hgu_cdac_8bit_array_2.drv<63:0>.n521 VSS 0.642f
C3584 hgu_cdac_8bit_array_2.drv<63:0>.n522 VSS -0.458f
C3585 hgu_cdac_8bit_array_2.drv<63:0>.n523 VSS -1.72f
C3586 hgu_cdac_8bit_array_2.drv<63:0>.n524 VSS 4.35f
C3587 hgu_cdac_8bit_array_2.drv<63:0>.n525 VSS -1.72f
C3588 hgu_cdac_8bit_array_2.drv<63:0>.n526 VSS -0.458f
C3589 hgu_cdac_8bit_array_2.drv<63:0>.n527 VSS 0.601f
C3590 hgu_cdac_8bit_array_2.drv<63:0>.n528 VSS 0.145f
C3591 hgu_cdac_8bit_array_2.drv<63:0>.n529 VSS 0.145f
C3592 hgu_cdac_8bit_array_2.drv<63:0>.n530 VSS 0.642f
C3593 hgu_cdac_8bit_array_2.drv<63:0>.n531 VSS -0.458f
C3594 hgu_cdac_8bit_array_2.drv<63:0>.n532 VSS -1.72f
C3595 hgu_cdac_8bit_array_2.drv<63:0>.n533 VSS 4.35f
C3596 hgu_cdac_8bit_array_2.drv<63:0>.n534 VSS -1.72f
C3597 hgu_cdac_8bit_array_2.drv<63:0>.n535 VSS -0.458f
C3598 hgu_cdac_8bit_array_2.drv<63:0>.n536 VSS 0.601f
C3599 hgu_cdac_8bit_array_2.drv<63:0>.n537 VSS 0.145f
C3600 hgu_cdac_8bit_array_2.drv<63:0>.n538 VSS 0.145f
C3601 hgu_cdac_8bit_array_2.drv<63:0>.n539 VSS 0.642f
C3602 hgu_cdac_8bit_array_2.drv<63:0>.n540 VSS -0.458f
C3603 hgu_cdac_8bit_array_2.drv<63:0>.n541 VSS -1.72f
C3604 hgu_cdac_8bit_array_2.drv<63:0>.n542 VSS 4.35f
C3605 hgu_cdac_8bit_array_2.drv<63:0>.n543 VSS -1.72f
C3606 hgu_cdac_8bit_array_2.drv<63:0>.n544 VSS -0.458f
C3607 hgu_cdac_8bit_array_2.drv<63:0>.n545 VSS 0.601f
C3608 hgu_cdac_8bit_array_2.drv<63:0>.n546 VSS 0.145f
C3609 hgu_cdac_8bit_array_2.drv<63:0>.n547 VSS 0.145f
C3610 hgu_cdac_8bit_array_2.drv<63:0>.n548 VSS 0.642f
C3611 hgu_cdac_8bit_array_2.drv<63:0>.n549 VSS -0.458f
C3612 hgu_cdac_8bit_array_2.drv<63:0>.n550 VSS -1.72f
C3613 hgu_cdac_8bit_array_2.drv<63:0>.n551 VSS 4.35f
C3614 hgu_cdac_8bit_array_2.drv<63:0>.n552 VSS -1.72f
C3615 hgu_cdac_8bit_array_2.drv<63:0>.n553 VSS -0.458f
C3616 hgu_cdac_8bit_array_2.drv<63:0>.n554 VSS 0.601f
C3617 hgu_cdac_8bit_array_2.drv<63:0>.n555 VSS 0.145f
C3618 hgu_cdac_8bit_array_2.drv<63:0>.n556 VSS 0.145f
C3619 hgu_cdac_8bit_array_2.drv<63:0>.n557 VSS 0.642f
C3620 hgu_cdac_8bit_array_2.drv<63:0>.n558 VSS -0.458f
C3621 hgu_cdac_8bit_array_2.drv<63:0>.n559 VSS -1.72f
C3622 hgu_cdac_8bit_array_2.drv<63:0>.n560 VSS 4.35f
C3623 hgu_cdac_8bit_array_2.drv<63:0>.n561 VSS -1.72f
C3624 hgu_cdac_8bit_array_2.drv<63:0>.n562 VSS -0.458f
C3625 hgu_cdac_8bit_array_2.drv<63:0>.n563 VSS 0.601f
C3626 hgu_cdac_8bit_array_2.drv<63:0>.n564 VSS 0.145f
C3627 hgu_cdac_8bit_array_2.drv<63:0>.n565 VSS 0.145f
C3628 hgu_cdac_8bit_array_2.drv<63:0>.n566 VSS 0.642f
C3629 hgu_cdac_8bit_array_2.drv<63:0>.n567 VSS -0.458f
C3630 hgu_cdac_8bit_array_2.drv<63:0>.n568 VSS -1.72f
C3631 hgu_cdac_8bit_array_2.drv<63:0>.n569 VSS 4.35f
C3632 hgu_cdac_8bit_array_2.drv<63:0>.n570 VSS -1.72f
C3633 hgu_cdac_8bit_array_2.drv<63:0>.n571 VSS -0.458f
C3634 hgu_cdac_8bit_array_2.drv<63:0>.n572 VSS 0.601f
C3635 hgu_cdac_8bit_array_2.drv<63:0>.n573 VSS 0.145f
C3636 hgu_cdac_8bit_array_2.drv<63:0>.n574 VSS 0.145f
C3637 hgu_cdac_8bit_array_2.drv<63:0>.n575 VSS 0.642f
C3638 hgu_cdac_8bit_array_2.drv<63:0>.n576 VSS -0.458f
C3639 hgu_cdac_8bit_array_2.drv<63:0>.n577 VSS -1.72f
C3640 hgu_cdac_8bit_array_2.drv<63:0>.n578 VSS 4.35f
C3641 hgu_cdac_8bit_array_2.drv<63:0>.n579 VSS -1.72f
C3642 hgu_cdac_8bit_array_2.drv<63:0>.n580 VSS -0.458f
C3643 hgu_cdac_8bit_array_2.drv<63:0>.n581 VSS 0.601f
C3644 hgu_cdac_8bit_array_2.drv<63:0>.n582 VSS 0.145f
C3645 hgu_cdac_8bit_array_2.drv<63:0>.n583 VSS 0.145f
C3646 hgu_cdac_8bit_array_2.drv<63:0>.n584 VSS 0.642f
C3647 hgu_cdac_8bit_array_2.drv<63:0>.n585 VSS -0.458f
C3648 hgu_cdac_8bit_array_2.drv<63:0>.n586 VSS -1.72f
C3649 hgu_cdac_8bit_array_2.drv<63:0>.n587 VSS 4.35f
C3650 hgu_cdac_8bit_array_2.drv<63:0>.n588 VSS -1.72f
C3651 hgu_cdac_8bit_array_2.drv<63:0>.n589 VSS -0.458f
C3652 hgu_cdac_8bit_array_2.drv<63:0>.n590 VSS 0.601f
C3653 hgu_cdac_8bit_array_2.drv<63:0>.n591 VSS 0.145f
C3654 hgu_cdac_8bit_array_2.drv<63:0>.n592 VSS 0.145f
C3655 hgu_cdac_8bit_array_2.drv<63:0>.n593 VSS 0.642f
C3656 hgu_cdac_8bit_array_2.drv<63:0>.n594 VSS -0.458f
C3657 hgu_cdac_8bit_array_2.drv<63:0>.n595 VSS -1.72f
C3658 hgu_cdac_8bit_array_2.drv<63:0>.n596 VSS 4.35f
C3659 hgu_cdac_8bit_array_2.drv<63:0>.n597 VSS -1.72f
C3660 hgu_cdac_8bit_array_2.drv<63:0>.n598 VSS -0.458f
C3661 hgu_cdac_8bit_array_2.drv<63:0>.n599 VSS 0.601f
C3662 hgu_cdac_8bit_array_2.drv<63:0>.n600 VSS 0.145f
C3663 hgu_cdac_8bit_array_2.drv<63:0>.n601 VSS 0.145f
C3664 hgu_cdac_8bit_array_2.drv<63:0>.n602 VSS 0.642f
C3665 hgu_cdac_8bit_array_2.drv<63:0>.n603 VSS -0.458f
C3666 hgu_cdac_8bit_array_2.drv<63:0>.n604 VSS -1.75f
C3667 db<6>.t101 VSS 0.0333f
C3668 db<6>.t56 VSS 0.0191f
C3669 db<6>.t19 VSS 0.0333f
C3670 db<6>.t108 VSS 0.0191f
C3671 db<6>.t30 VSS 0.0333f
C3672 db<6>.t120 VSS 0.0191f
C3673 db<6>.t79 VSS 0.0333f
C3674 db<6>.t35 VSS 0.0191f
C3675 db<6>.t97 VSS 0.0333f
C3676 db<6>.t52 VSS 0.0191f
C3677 db<6>.t41 VSS 0.0333f
C3678 db<6>.t3 VSS 0.0191f
C3679 db<6>.t91 VSS 0.0333f
C3680 db<6>.t46 VSS 0.0191f
C3681 db<6>.t72 VSS 0.0333f
C3682 db<6>.t29 VSS 0.0191f
C3683 db<6>.t123 VSS 0.0333f
C3684 db<6>.t78 VSS 0.0191f
C3685 db<6>.t38 VSS 0.0333f
C3686 db<6>.t0 VSS 0.0191f
C3687 db<6>.t88 VSS 0.0333f
C3688 db<6>.t43 VSS 0.0191f
C3689 db<6>.t106 VSS 0.0333f
C3690 db<6>.t61 VSS 0.0191f
C3691 db<6>.t118 VSS 0.0333f
C3692 db<6>.t74 VSS 0.0191f
C3693 db<6>.t82 VSS 0.0333f
C3694 db<6>.t36 VSS 0.0191f
C3695 db<6>.t98 VSS 0.0333f
C3696 db<6>.t53 VSS 0.0191f
C3697 db<6>.t15 VSS 0.0333f
C3698 db<6>.t104 VSS 0.0191f
C3699 db<6>.t63 VSS 0.0333f
C3700 db<6>.t20 VSS 0.0191f
C3701 db<6>.t77 VSS 0.0333f
C3702 db<6>.t33 VSS 0.0191f
C3703 db<6>.t93 VSS 0.0333f
C3704 db<6>.t48 VSS 0.0191f
C3705 db<6>.t12 VSS 0.0333f
C3706 db<6>.t100 VSS 0.0191f
C3707 db<6>.t59 VSS 0.0333f
C3708 db<6>.t17 VSS 0.0191f
C3709 db<6>.t119 VSS 0.0333f
C3710 db<6>.t75 VSS 0.0191f
C3711 db<6>.t6 VSS 0.0333f
C3712 db<6>.t90 VSS 0.0191f
C3713 db<6>.t50 VSS 0.0333f
C3714 db<6>.t11 VSS 0.0191f
C3715 db<6>.t102 VSS 0.0333f
C3716 db<6>.t57 VSS 0.0191f
C3717 db<6>.t117 VSS 0.0333f
C3718 db<6>.t71 VSS 0.0191f
C3719 db<6>.t32 VSS 0.0333f
C3720 db<6>.t122 VSS 0.0191f
C3721 db<6>.t45 VSS 0.0333f
C3722 db<6>.t8 VSS 0.0191f
C3723 db<6>.t99 VSS 0.0333f
C3724 db<6>.t54 VSS 0.0191f
C3725 db<6>.t27 VSS 0.0333f
C3726 db<6>.t116 VSS 0.0191f
C3727 db<6>.t73 VSS 0.0333f
C3728 db<6>.t31 VSS 0.0191f
C3729 db<6>.t125 VSS 0.0333f
C3730 db<6>.t80 VSS 0.0191f
C3731 db<6>.t109 VSS 0.0333f
C3732 db<6>.t62 VSS 0.0191f
C3733 db<6>.t25 VSS 0.0333f
C3734 db<6>.t113 VSS 0.0191f
C3735 db<6>.t70 VSS 0.0333f
C3736 db<6>.t28 VSS 0.0191f
C3737 db<6>.t121 VSS 0.0333f
C3738 db<6>.t76 VSS 0.0191f
C3739 db<6>.t47 VSS 0.0333f
C3740 db<6>.t10 VSS 0.0191f
C3741 db<6>.t65 VSS 0.0333f
C3742 db<6>.t22 VSS 0.0191f
C3743 db<6>.t115 VSS 0.0333f
C3744 db<6>.t69 VSS 0.0191f
C3745 db<6>.t1 VSS 0.0333f
C3746 db<6>.t86 VSS 0.0191f
C3747 db<6>.t44 VSS 0.0333f
C3748 db<6>.t5 VSS 0.0191f
C3749 db<6>.t95 VSS 0.0333f
C3750 db<6>.t49 VSS 0.0191f
C3751 db<6>.t112 VSS 0.0333f
C3752 db<6>.t68 VSS 0.0191f
C3753 db<6>.t127 VSS 0.0333f
C3754 db<6>.t84 VSS 0.0191f
C3755 db<6>.t87 VSS 0.0333f
C3756 db<6>.t42 VSS 0.0191f
C3757 db<6>.t7 VSS 0.0333f
C3758 db<6>.t92 VSS 0.0191f
C3759 db<6>.t21 VSS 0.0333f
C3760 db<6>.t111 VSS 0.0191f
C3761 db<6>.t34 VSS 0.0333f
C3762 db<6>.t124 VSS 0.0191f
C3763 db<6>.t85 VSS 0.0333f
C3764 db<6>.t39 VSS 0.0191f
C3765 db<6>.t4 VSS 0.0333f
C3766 db<6>.t89 VSS 0.0191f
C3767 db<6>.t18 VSS 0.0333f
C3768 db<6>.t107 VSS 0.0191f
C3769 db<6>.t67 VSS 0.0333f
C3770 db<6>.t24 VSS 0.0191f
C3771 db<6>.t126 VSS 0.0333f
C3772 db<6>.t83 VSS 0.0191f
C3773 db<6>.t40 VSS 0.0333f
C3774 db<6>.t2 VSS 0.0191f
C3775 db<6>.t58 VSS 0.0333f
C3776 db<6>.t16 VSS 0.0191f
C3777 db<6>.t110 VSS 0.0333f
C3778 db<6>.t64 VSS 0.0191f
C3779 db<6>.t26 VSS 0.0333f
C3780 db<6>.t114 VSS 0.0191f
C3781 db<6>.t9 VSS 0.0333f
C3782 db<6>.t94 VSS 0.0191f
C3783 db<6>.t55 VSS 0.0333f
C3784 db<6>.t13 VSS 0.0191f
C3785 db<6>.t105 VSS 0.0333f
C3786 db<6>.t60 VSS 0.0191f
C3787 db<6>.t66 VSS 0.0333f
C3788 db<6>.t23 VSS 0.0191f
C3789 db<6>.t81 VSS 0.0333f
C3790 db<6>.t37 VSS 0.0191f
C3791 db<6>.t96 VSS 0.0333f
C3792 db<6>.t51 VSS 0.0191f
C3793 db<6>.t14 VSS 0.0333f
C3794 db<6>.t103 VSS 0.0191f
C3795 db<6>.n0 VSS 0.062f
C3796 db<6>.n1 VSS 0.0713f
C3797 db<6>.n2 VSS 0.0713f
C3798 db<6>.n3 VSS 0.0713f
C3799 db<6>.n4 VSS 0.0713f
C3800 db<6>.n5 VSS 0.0713f
C3801 db<6>.n6 VSS 0.0713f
C3802 db<6>.n7 VSS 0.0713f
C3803 db<6>.n8 VSS 0.0713f
C3804 db<6>.n9 VSS 0.0713f
C3805 db<6>.n10 VSS 0.0713f
C3806 db<6>.n11 VSS 0.0713f
C3807 db<6>.n12 VSS 0.0713f
C3808 db<6>.n13 VSS 0.0713f
C3809 db<6>.n14 VSS 0.0713f
C3810 db<6>.n15 VSS 0.0713f
C3811 db<6>.n16 VSS 0.0713f
C3812 db<6>.n17 VSS 0.0713f
C3813 db<6>.n18 VSS 0.0713f
C3814 db<6>.n19 VSS 0.0713f
C3815 db<6>.n20 VSS 0.0713f
C3816 db<6>.n21 VSS 0.0713f
C3817 db<6>.n22 VSS 0.0713f
C3818 db<6>.n23 VSS 0.0713f
C3819 db<6>.n24 VSS 0.0713f
C3820 db<6>.n25 VSS 0.0713f
C3821 db<6>.n26 VSS 0.0713f
C3822 db<6>.n27 VSS 0.0713f
C3823 db<6>.n28 VSS 0.0713f
C3824 db<6>.n29 VSS 0.0713f
C3825 db<6>.n30 VSS 0.0713f
C3826 db<6>.n31 VSS 0.0713f
C3827 db<6>.n32 VSS 0.0713f
C3828 db<6>.n33 VSS 0.0713f
C3829 db<6>.n34 VSS 0.0713f
C3830 db<6>.n35 VSS 0.0713f
C3831 db<6>.n36 VSS 0.0713f
C3832 db<6>.n37 VSS 0.0713f
C3833 db<6>.n38 VSS 0.0713f
C3834 db<6>.n39 VSS 0.0713f
C3835 db<6>.n40 VSS 0.0713f
C3836 db<6>.n41 VSS 0.0713f
C3837 db<6>.n42 VSS 0.0713f
C3838 db<6>.n43 VSS 0.0713f
C3839 db<6>.n44 VSS 0.0713f
C3840 db<6>.n45 VSS 0.0713f
C3841 db<6>.n46 VSS 0.0713f
C3842 db<6>.n47 VSS 0.0713f
C3843 db<6>.n48 VSS 0.0713f
C3844 db<6>.n49 VSS 0.0713f
C3845 db<6>.n50 VSS 0.0713f
C3846 db<6>.n51 VSS 0.0713f
C3847 db<6>.n52 VSS 0.0713f
C3848 db<6>.n53 VSS 0.0713f
C3849 db<6>.n54 VSS 0.0713f
C3850 db<6>.n55 VSS 0.0713f
C3851 db<6>.n56 VSS 0.0713f
C3852 db<6>.n57 VSS 0.0713f
C3853 db<6>.n58 VSS 0.0713f
C3854 db<6>.n59 VSS 0.0713f
C3855 db<6>.n60 VSS 0.0713f
C3856 db<6>.n61 VSS 0.0713f
C3857 db<6>.n62 VSS 0.0713f
C3858 db<6>.n63 VSS 0.0564f
C3859 hgu_cdac_8bit_array_3.drv<31:0>.n0 VSS 3.93f
C3860 hgu_cdac_8bit_array_3.drv<31:0>.n1 VSS 3.95f
C3861 hgu_cdac_8bit_array_3.drv<31:0>.n2 VSS -14.5f
C3862 hgu_cdac_8bit_array_3.drv<31:0>.t11 VSS 0.0528f
C3863 hgu_cdac_8bit_array_3.drv<31:0>.t8 VSS 0.0528f
C3864 hgu_cdac_8bit_array_3.drv<31:0>.n3 VSS 0.373f
C3865 hgu_cdac_8bit_array_3.drv<31:0>.t40 VSS 0.106f
C3866 hgu_cdac_8bit_array_3.drv<31:0>.t20 VSS 0.106f
C3867 hgu_cdac_8bit_array_3.drv<31:0>.n4 VSS 0.758f
C3868 hgu_cdac_8bit_array_3.drv<31:0>.t50 VSS 0.0528f
C3869 hgu_cdac_8bit_array_3.drv<31:0>.t53 VSS 0.0528f
C3870 hgu_cdac_8bit_array_3.drv<31:0>.n5 VSS 0.39f
C3871 hgu_cdac_8bit_array_3.drv<31:0>.t32 VSS 0.106f
C3872 hgu_cdac_8bit_array_3.drv<31:0>.t35 VSS 0.106f
C3873 hgu_cdac_8bit_array_3.drv<31:0>.n6 VSS 0.804f
C3874 hgu_cdac_8bit_array_3.drv<31:0>.n7 VSS 0.506f
C3875 hgu_cdac_8bit_array_3.drv<31:0>.n8 VSS 0.419f
C3876 hgu_cdac_8bit_array_3.drv<31:0>.t49 VSS 0.0528f
C3877 hgu_cdac_8bit_array_3.drv<31:0>.t3 VSS 0.0528f
C3878 hgu_cdac_8bit_array_3.drv<31:0>.n9 VSS 0.39f
C3879 hgu_cdac_8bit_array_3.drv<31:0>.t31 VSS 0.106f
C3880 hgu_cdac_8bit_array_3.drv<31:0>.t15 VSS 0.106f
C3881 hgu_cdac_8bit_array_3.drv<31:0>.n10 VSS 0.804f
C3882 hgu_cdac_8bit_array_3.drv<31:0>.n11 VSS 0.473f
C3883 hgu_cdac_8bit_array_3.drv<31:0>.n12 VSS 3.64f
C3884 hgu_cdac_8bit_array_3.drv<31:0>.n13 VSS 8.27f
C3885 hgu_cdac_8bit_array_3.drv<31:0>.n14 VSS -1.74f
C3886 hgu_cdac_8bit_array_3.drv<31:0>.n15 VSS -1.11f
C3887 hgu_cdac_8bit_array_3.drv<31:0>.n16 VSS -1.78f
C3888 hgu_cdac_8bit_array_3.drv<31:0>.n17 VSS -1.78f
C3889 hgu_cdac_8bit_array_3.drv<31:0>.n18 VSS -1.11f
C3890 hgu_cdac_8bit_array_3.drv<31:0>.n19 VSS -1.74f
C3891 hgu_cdac_8bit_array_3.drv<31:0>.n20 VSS 4f
C3892 hgu_cdac_8bit_array_3.drv<31:0>.t2 VSS 0.0528f
C3893 hgu_cdac_8bit_array_3.drv<31:0>.t54 VSS 0.0528f
C3894 hgu_cdac_8bit_array_3.drv<31:0>.n21 VSS 0.39f
C3895 hgu_cdac_8bit_array_3.drv<31:0>.t46 VSS 0.106f
C3896 hgu_cdac_8bit_array_3.drv<31:0>.t36 VSS 0.106f
C3897 hgu_cdac_8bit_array_3.drv<31:0>.n22 VSS 0.804f
C3898 hgu_cdac_8bit_array_3.drv<31:0>.n23 VSS 0.48f
C3899 hgu_cdac_8bit_array_3.drv<31:0>.t12 VSS 0.0528f
C3900 hgu_cdac_8bit_array_3.drv<31:0>.t9 VSS 0.0528f
C3901 hgu_cdac_8bit_array_3.drv<31:0>.n24 VSS 0.373f
C3902 hgu_cdac_8bit_array_3.drv<31:0>.t41 VSS 0.106f
C3903 hgu_cdac_8bit_array_3.drv<31:0>.t21 VSS 0.106f
C3904 hgu_cdac_8bit_array_3.drv<31:0>.n25 VSS 0.758f
C3905 hgu_cdac_8bit_array_3.drv<31:0>.n26 VSS 0.402f
C3906 hgu_cdac_8bit_array_3.drv<31:0>.n27 VSS 3.58f
C3907 hgu_cdac_8bit_array_3.drv<31:0>.n28 VSS 8.26f
C3908 hgu_cdac_8bit_array_3.drv<31:0>.t4 VSS 0.0528f
C3909 hgu_cdac_8bit_array_3.drv<31:0>.t59 VSS 0.0528f
C3910 hgu_cdac_8bit_array_3.drv<31:0>.n29 VSS 0.39f
C3911 hgu_cdac_8bit_array_3.drv<31:0>.t16 VSS 0.106f
C3912 hgu_cdac_8bit_array_3.drv<31:0>.t26 VSS 0.106f
C3913 hgu_cdac_8bit_array_3.drv<31:0>.n30 VSS 0.804f
C3914 hgu_cdac_8bit_array_3.drv<31:0>.n31 VSS 0.423f
C3915 hgu_cdac_8bit_array_3.drv<31:0>.t48 VSS 0.0528f
C3916 hgu_cdac_8bit_array_3.drv<31:0>.t14 VSS 0.0528f
C3917 hgu_cdac_8bit_array_3.drv<31:0>.n32 VSS 0.39f
C3918 hgu_cdac_8bit_array_3.drv<31:0>.t30 VSS 0.106f
C3919 hgu_cdac_8bit_array_3.drv<31:0>.t43 VSS 0.106f
C3920 hgu_cdac_8bit_array_3.drv<31:0>.n33 VSS 0.804f
C3921 hgu_cdac_8bit_array_3.drv<31:0>.n34 VSS 0.415f
C3922 hgu_cdac_8bit_array_3.drv<31:0>.n35 VSS 3.61f
C3923 hgu_cdac_8bit_array_3.drv<31:0>.n36 VSS -1.74f
C3924 hgu_cdac_8bit_array_3.drv<31:0>.n37 VSS -1.11f
C3925 hgu_cdac_8bit_array_3.drv<31:0>.n38 VSS -1.78f
C3926 hgu_cdac_8bit_array_3.drv<31:0>.n39 VSS -1.78f
C3927 hgu_cdac_8bit_array_3.drv<31:0>.n40 VSS -1.11f
C3928 hgu_cdac_8bit_array_3.drv<31:0>.n41 VSS -1.74f
C3929 hgu_cdac_8bit_array_3.drv<31:0>.n42 VSS 4f
C3930 hgu_cdac_8bit_array_3.drv<31:0>.n43 VSS 8.25f
C3931 hgu_cdac_8bit_array_3.drv<31:0>.t55 VSS 0.0528f
C3932 hgu_cdac_8bit_array_3.drv<31:0>.t60 VSS 0.0528f
C3933 hgu_cdac_8bit_array_3.drv<31:0>.n44 VSS 0.373f
C3934 hgu_cdac_8bit_array_3.drv<31:0>.t37 VSS 0.106f
C3935 hgu_cdac_8bit_array_3.drv<31:0>.t27 VSS 0.106f
C3936 hgu_cdac_8bit_array_3.drv<31:0>.n45 VSS 0.752f
C3937 hgu_cdac_8bit_array_3.drv<31:0>.t62 VSS 0.0528f
C3938 hgu_cdac_8bit_array_3.drv<31:0>.t57 VSS 0.0528f
C3939 hgu_cdac_8bit_array_3.drv<31:0>.n46 VSS 0.39f
C3940 hgu_cdac_8bit_array_3.drv<31:0>.t22 VSS 0.106f
C3941 hgu_cdac_8bit_array_3.drv<31:0>.t24 VSS 0.106f
C3942 hgu_cdac_8bit_array_3.drv<31:0>.n47 VSS 0.804f
C3943 hgu_cdac_8bit_array_3.drv<31:0>.n48 VSS 0.506f
C3944 hgu_cdac_8bit_array_3.drv<31:0>.n49 VSS 0.429f
C3945 hgu_cdac_8bit_array_3.drv<31:0>.t10 VSS 0.0528f
C3946 hgu_cdac_8bit_array_3.drv<31:0>.t51 VSS 0.0528f
C3947 hgu_cdac_8bit_array_3.drv<31:0>.n50 VSS 0.39f
C3948 hgu_cdac_8bit_array_3.drv<31:0>.t39 VSS 0.106f
C3949 hgu_cdac_8bit_array_3.drv<31:0>.t33 VSS 0.106f
C3950 hgu_cdac_8bit_array_3.drv<31:0>.n51 VSS 0.804f
C3951 hgu_cdac_8bit_array_3.drv<31:0>.n52 VSS 0.471f
C3952 hgu_cdac_8bit_array_3.drv<31:0>.n53 VSS 3.59f
C3953 hgu_cdac_8bit_array_3.drv<31:0>.n54 VSS -1.74f
C3954 hgu_cdac_8bit_array_3.drv<31:0>.n55 VSS -1.11f
C3955 hgu_cdac_8bit_array_3.drv<31:0>.n56 VSS -1.78f
C3956 hgu_cdac_8bit_array_3.drv<31:0>.n57 VSS -1.78f
C3957 hgu_cdac_8bit_array_3.drv<31:0>.n58 VSS -1.11f
C3958 hgu_cdac_8bit_array_3.drv<31:0>.n59 VSS -1.74f
C3959 hgu_cdac_8bit_array_3.drv<31:0>.n60 VSS 4f
C3960 hgu_cdac_8bit_array_3.drv<31:0>.n61 VSS 8.25f
C3961 hgu_cdac_8bit_array_3.drv<31:0>.t56 VSS 0.0528f
C3962 hgu_cdac_8bit_array_3.drv<31:0>.t6 VSS 0.0528f
C3963 hgu_cdac_8bit_array_3.drv<31:0>.n62 VSS 0.373f
C3964 hgu_cdac_8bit_array_3.drv<31:0>.t38 VSS 0.106f
C3965 hgu_cdac_8bit_array_3.drv<31:0>.t18 VSS 0.106f
C3966 hgu_cdac_8bit_array_3.drv<31:0>.n63 VSS 0.758f
C3967 hgu_cdac_8bit_array_3.drv<31:0>.n64 VSS 3.91f
C3968 hgu_cdac_8bit_array_3.drv<31:0>.n65 VSS -1.74f
C3969 hgu_cdac_8bit_array_3.drv<31:0>.n66 VSS -1.11f
C3970 hgu_cdac_8bit_array_3.drv<31:0>.n67 VSS -1.78f
C3971 hgu_cdac_8bit_array_3.drv<31:0>.n68 VSS -1.78f
C3972 hgu_cdac_8bit_array_3.drv<31:0>.n69 VSS -1.11f
C3973 hgu_cdac_8bit_array_3.drv<31:0>.n70 VSS -1.74f
C3974 hgu_cdac_8bit_array_3.drv<31:0>.n71 VSS 4f
C3975 hgu_cdac_8bit_array_3.drv<31:0>.n72 VSS 8.29f
C3976 hgu_cdac_8bit_array_3.drv<31:0>.n73 VSS -1.74f
C3977 hgu_cdac_8bit_array_3.drv<31:0>.n74 VSS -1.11f
C3978 hgu_cdac_8bit_array_3.drv<31:0>.n75 VSS -1.78f
C3979 hgu_cdac_8bit_array_3.drv<31:0>.n76 VSS -1.78f
C3980 hgu_cdac_8bit_array_3.drv<31:0>.n77 VSS -1.11f
C3981 hgu_cdac_8bit_array_3.drv<31:0>.n78 VSS -1.74f
C3982 hgu_cdac_8bit_array_3.drv<31:0>.n79 VSS 6.18f
C3983 hgu_cdac_8bit_array_3.drv<31:0>.n80 VSS -1.74f
C3984 hgu_cdac_8bit_array_3.drv<31:0>.n81 VSS -1.11f
C3985 hgu_cdac_8bit_array_3.drv<31:0>.n82 VSS -1.78f
C3986 hgu_cdac_8bit_array_3.drv<31:0>.n83 VSS -1.78f
C3987 hgu_cdac_8bit_array_3.drv<31:0>.n84 VSS -1.11f
C3988 hgu_cdac_8bit_array_3.drv<31:0>.n85 VSS -1.74f
C3989 hgu_cdac_8bit_array_3.drv<31:0>.n86 VSS 6.18f
C3990 hgu_cdac_8bit_array_3.drv<31:0>.n87 VSS -1.74f
C3991 hgu_cdac_8bit_array_3.drv<31:0>.n88 VSS -1.11f
C3992 hgu_cdac_8bit_array_3.drv<31:0>.n89 VSS -1.78f
C3993 hgu_cdac_8bit_array_3.drv<31:0>.n90 VSS -1.78f
C3994 hgu_cdac_8bit_array_3.drv<31:0>.n91 VSS -1.11f
C3995 hgu_cdac_8bit_array_3.drv<31:0>.n92 VSS -1.74f
C3996 hgu_cdac_8bit_array_3.drv<31:0>.n93 VSS 6.18f
C3997 hgu_cdac_8bit_array_3.drv<31:0>.n94 VSS -1.74f
C3998 hgu_cdac_8bit_array_3.drv<31:0>.n95 VSS -1.11f
C3999 hgu_cdac_8bit_array_3.drv<31:0>.n96 VSS -1.78f
C4000 hgu_cdac_8bit_array_3.drv<31:0>.n97 VSS -1.78f
C4001 hgu_cdac_8bit_array_3.drv<31:0>.n98 VSS -1.11f
C4002 hgu_cdac_8bit_array_3.drv<31:0>.n99 VSS -1.74f
C4003 hgu_cdac_8bit_array_3.drv<31:0>.n100 VSS 6.18f
C4004 hgu_cdac_8bit_array_3.drv<31:0>.n101 VSS -1.74f
C4005 hgu_cdac_8bit_array_3.drv<31:0>.n102 VSS -1.11f
C4006 hgu_cdac_8bit_array_3.drv<31:0>.n103 VSS -1.78f
C4007 hgu_cdac_8bit_array_3.drv<31:0>.n104 VSS -1.78f
C4008 hgu_cdac_8bit_array_3.drv<31:0>.n105 VSS -1.11f
C4009 hgu_cdac_8bit_array_3.drv<31:0>.n106 VSS -1.74f
C4010 hgu_cdac_8bit_array_3.drv<31:0>.n107 VSS 6.18f
C4011 hgu_cdac_8bit_array_3.drv<31:0>.n108 VSS -1.74f
C4012 hgu_cdac_8bit_array_3.drv<31:0>.n109 VSS -1.11f
C4013 hgu_cdac_8bit_array_3.drv<31:0>.n110 VSS -1.78f
C4014 hgu_cdac_8bit_array_3.drv<31:0>.n111 VSS -1.78f
C4015 hgu_cdac_8bit_array_3.drv<31:0>.n112 VSS -1.11f
C4016 hgu_cdac_8bit_array_3.drv<31:0>.n113 VSS -1.74f
C4017 hgu_cdac_8bit_array_3.drv<31:0>.n114 VSS 6.18f
C4018 hgu_cdac_8bit_array_3.drv<31:0>.n115 VSS -1.74f
C4019 hgu_cdac_8bit_array_3.drv<31:0>.n116 VSS -1.11f
C4020 hgu_cdac_8bit_array_3.drv<31:0>.n117 VSS -1.78f
C4021 hgu_cdac_8bit_array_3.drv<31:0>.n118 VSS -1.78f
C4022 hgu_cdac_8bit_array_3.drv<31:0>.n119 VSS -1.11f
C4023 hgu_cdac_8bit_array_3.drv<31:0>.n120 VSS -1.74f
C4024 hgu_cdac_8bit_array_3.drv<31:0>.n121 VSS 6.18f
C4025 hgu_cdac_8bit_array_3.drv<31:0>.n122 VSS -1.54f
C4026 hgu_cdac_8bit_array_3.drv<31:0>.n123 VSS -1.74f
C4027 hgu_cdac_8bit_array_3.drv<31:0>.n124 VSS 6.18f
C4028 hgu_cdac_8bit_array_3.drv<31:0>.n125 VSS 4.65f
C4029 hgu_cdac_8bit_array_3.drv<31:0>.n126 VSS 0.746f
C4030 hgu_cdac_8bit_array_3.drv<31:0>.n127 VSS -0.465f
C4031 hgu_cdac_8bit_array_3.drv<31:0>.n128 VSS -1.74f
C4032 hgu_cdac_8bit_array_3.drv<31:0>.n129 VSS 6.19f
C4033 hgu_cdac_8bit_array_3.drv<31:0>.n130 VSS -1.74f
C4034 hgu_cdac_8bit_array_3.drv<31:0>.n131 VSS -0.465f
C4035 hgu_cdac_8bit_array_3.drv<31:0>.n132 VSS 0.651f
C4036 hgu_cdac_8bit_array_3.drv<31:0>.n133 VSS 0.147f
C4037 hgu_cdac_8bit_array_3.drv<31:0>.n134 VSS 0.147f
C4038 hgu_cdac_8bit_array_3.drv<31:0>.n135 VSS 0.61f
C4039 hgu_cdac_8bit_array_3.drv<31:0>.n136 VSS -0.465f
C4040 hgu_cdac_8bit_array_3.drv<31:0>.n137 VSS -1.74f
C4041 hgu_cdac_8bit_array_3.drv<31:0>.n138 VSS 6.19f
C4042 hgu_cdac_8bit_array_3.drv<31:0>.n139 VSS -1.74f
C4043 hgu_cdac_8bit_array_3.drv<31:0>.n140 VSS -0.465f
C4044 hgu_cdac_8bit_array_3.drv<31:0>.n141 VSS 0.651f
C4045 hgu_cdac_8bit_array_3.drv<31:0>.n142 VSS 0.147f
C4046 hgu_cdac_8bit_array_3.drv<31:0>.n143 VSS 0.147f
C4047 hgu_cdac_8bit_array_3.drv<31:0>.n144 VSS 0.61f
C4048 hgu_cdac_8bit_array_3.drv<31:0>.n145 VSS -0.465f
C4049 hgu_cdac_8bit_array_3.drv<31:0>.n146 VSS -1.74f
C4050 hgu_cdac_8bit_array_3.drv<31:0>.n147 VSS 6.19f
C4051 hgu_cdac_8bit_array_3.drv<31:0>.n148 VSS -1.74f
C4052 hgu_cdac_8bit_array_3.drv<31:0>.n149 VSS -0.465f
C4053 hgu_cdac_8bit_array_3.drv<31:0>.n150 VSS 0.651f
C4054 hgu_cdac_8bit_array_3.drv<31:0>.n151 VSS 0.147f
C4055 hgu_cdac_8bit_array_3.drv<31:0>.n152 VSS 0.147f
C4056 hgu_cdac_8bit_array_3.drv<31:0>.n153 VSS 0.61f
C4057 hgu_cdac_8bit_array_3.drv<31:0>.n154 VSS -0.465f
C4058 hgu_cdac_8bit_array_3.drv<31:0>.n155 VSS -1.74f
C4059 hgu_cdac_8bit_array_3.drv<31:0>.n156 VSS 6.19f
C4060 hgu_cdac_8bit_array_3.drv<31:0>.n157 VSS -1.74f
C4061 hgu_cdac_8bit_array_3.drv<31:0>.n158 VSS -0.465f
C4062 hgu_cdac_8bit_array_3.drv<31:0>.n159 VSS 0.651f
C4063 hgu_cdac_8bit_array_3.drv<31:0>.n160 VSS 0.147f
C4064 hgu_cdac_8bit_array_3.drv<31:0>.n161 VSS 0.147f
C4065 hgu_cdac_8bit_array_3.drv<31:0>.n162 VSS 0.61f
C4066 hgu_cdac_8bit_array_3.drv<31:0>.n163 VSS -0.465f
C4067 hgu_cdac_8bit_array_3.drv<31:0>.n164 VSS -1.74f
C4068 hgu_cdac_8bit_array_3.drv<31:0>.n165 VSS 6.19f
C4069 hgu_cdac_8bit_array_3.drv<31:0>.n166 VSS -1.74f
C4070 hgu_cdac_8bit_array_3.drv<31:0>.n167 VSS -0.465f
C4071 hgu_cdac_8bit_array_3.drv<31:0>.n168 VSS 0.651f
C4072 hgu_cdac_8bit_array_3.drv<31:0>.n169 VSS 0.147f
C4073 hgu_cdac_8bit_array_3.drv<31:0>.n170 VSS 0.147f
C4074 hgu_cdac_8bit_array_3.drv<31:0>.n171 VSS 0.61f
C4075 hgu_cdac_8bit_array_3.drv<31:0>.n172 VSS -0.465f
C4076 hgu_cdac_8bit_array_3.drv<31:0>.n173 VSS -1.74f
C4077 hgu_cdac_8bit_array_3.drv<31:0>.n174 VSS 6.19f
C4078 hgu_cdac_8bit_array_3.drv<31:0>.n175 VSS -1.74f
C4079 hgu_cdac_8bit_array_3.drv<31:0>.n176 VSS -0.465f
C4080 hgu_cdac_8bit_array_3.drv<31:0>.n177 VSS 0.651f
C4081 hgu_cdac_8bit_array_3.drv<31:0>.n178 VSS 0.147f
C4082 hgu_cdac_8bit_array_3.drv<31:0>.n179 VSS 0.147f
C4083 hgu_cdac_8bit_array_3.drv<31:0>.n180 VSS 0.61f
C4084 hgu_cdac_8bit_array_3.drv<31:0>.n181 VSS -0.465f
C4085 hgu_cdac_8bit_array_3.drv<31:0>.n182 VSS -1.74f
C4086 hgu_cdac_8bit_array_3.drv<31:0>.n183 VSS 6.19f
C4087 hgu_cdac_8bit_array_3.drv<31:0>.n184 VSS -1.74f
C4088 hgu_cdac_8bit_array_3.drv<31:0>.n185 VSS -0.465f
C4089 hgu_cdac_8bit_array_3.drv<31:0>.n186 VSS 0.651f
C4090 hgu_cdac_8bit_array_3.drv<31:0>.n187 VSS 0.147f
C4091 hgu_cdac_8bit_array_3.drv<31:0>.n188 VSS 0.147f
C4092 hgu_cdac_8bit_array_3.drv<31:0>.n189 VSS 0.61f
C4093 hgu_cdac_8bit_array_3.drv<31:0>.n190 VSS -0.465f
C4094 hgu_cdac_8bit_array_3.drv<31:0>.n191 VSS -1.74f
C4095 hgu_cdac_8bit_array_3.drv<31:0>.n192 VSS 6.19f
C4096 hgu_cdac_8bit_array_3.drv<31:0>.n193 VSS -1.74f
C4097 hgu_cdac_8bit_array_3.drv<31:0>.n194 VSS -0.465f
C4098 hgu_cdac_8bit_array_3.drv<31:0>.n195 VSS 0.651f
C4099 hgu_cdac_8bit_array_3.drv<31:0>.n196 VSS 0.147f
C4100 hgu_cdac_8bit_array_3.drv<31:0>.n197 VSS 0.147f
C4101 hgu_cdac_8bit_array_3.drv<31:0>.n198 VSS 0.61f
C4102 hgu_cdac_8bit_array_3.drv<31:0>.n199 VSS -0.465f
C4103 hgu_cdac_8bit_array_3.drv<31:0>.n200 VSS -1.74f
C4104 hgu_cdac_8bit_array_3.drv<31:0>.n201 VSS 4.41f
C4105 hgu_cdac_8bit_array_3.drv<31:0>.n202 VSS -1.74f
C4106 hgu_cdac_8bit_array_3.drv<31:0>.n203 VSS -0.465f
C4107 hgu_cdac_8bit_array_3.drv<31:0>.n204 VSS 0.529f
C4108 hgu_cdac_8bit_array_3.drv<31:0>.n205 VSS 0.147f
C4109 hgu_cdac_8bit_array_3.drv<31:0>.n206 VSS 0.147f
C4110 hgu_cdac_8bit_array_3.drv<31:0>.n207 VSS 0.61f
C4111 hgu_cdac_8bit_array_3.drv<31:0>.n208 VSS -0.465f
C4112 hgu_cdac_8bit_array_3.drv<31:0>.n209 VSS -1.74f
C4113 hgu_cdac_8bit_array_3.drv<31:0>.n210 VSS 4.41f
C4114 hgu_cdac_8bit_array_3.drv<31:0>.n211 VSS -1.74f
C4115 hgu_cdac_8bit_array_3.drv<31:0>.n212 VSS -0.465f
C4116 hgu_cdac_8bit_array_3.drv<31:0>.n213 VSS 0.651f
C4117 hgu_cdac_8bit_array_3.drv<31:0>.n214 VSS 0.147f
C4118 hgu_cdac_8bit_array_3.drv<31:0>.n215 VSS 0.147f
C4119 hgu_cdac_8bit_array_3.drv<31:0>.n216 VSS 0.61f
C4120 hgu_cdac_8bit_array_3.drv<31:0>.n217 VSS -0.465f
C4121 hgu_cdac_8bit_array_3.drv<31:0>.n218 VSS -1.74f
C4122 hgu_cdac_8bit_array_3.drv<31:0>.n219 VSS 4.41f
C4123 hgu_cdac_8bit_array_3.drv<31:0>.n220 VSS -1.74f
C4124 hgu_cdac_8bit_array_3.drv<31:0>.n221 VSS -0.465f
C4125 hgu_cdac_8bit_array_3.drv<31:0>.n222 VSS 0.651f
C4126 hgu_cdac_8bit_array_3.drv<31:0>.n223 VSS 0.147f
C4127 hgu_cdac_8bit_array_3.drv<31:0>.n224 VSS 0.147f
C4128 hgu_cdac_8bit_array_3.drv<31:0>.n225 VSS 0.61f
C4129 hgu_cdac_8bit_array_3.drv<31:0>.n226 VSS -0.465f
C4130 hgu_cdac_8bit_array_3.drv<31:0>.n227 VSS -1.74f
C4131 hgu_cdac_8bit_array_3.drv<31:0>.n228 VSS 4.41f
C4132 hgu_cdac_8bit_array_3.drv<31:0>.n229 VSS -1.74f
C4133 hgu_cdac_8bit_array_3.drv<31:0>.n230 VSS -0.465f
C4134 hgu_cdac_8bit_array_3.drv<31:0>.n231 VSS 0.651f
C4135 hgu_cdac_8bit_array_3.drv<31:0>.n232 VSS 0.147f
C4136 hgu_cdac_8bit_array_3.drv<31:0>.n233 VSS 0.147f
C4137 hgu_cdac_8bit_array_3.drv<31:0>.n234 VSS 0.61f
C4138 hgu_cdac_8bit_array_3.drv<31:0>.n235 VSS -0.465f
C4139 hgu_cdac_8bit_array_3.drv<31:0>.n236 VSS -1.74f
C4140 hgu_cdac_8bit_array_3.drv<31:0>.n237 VSS 4.29f
C4141 hgu_cdac_8bit_array_3.drv<31:0>.n238 VSS -1.74f
C4142 hgu_cdac_8bit_array_3.drv<31:0>.n239 VSS -1.11f
C4143 hgu_cdac_8bit_array_3.drv<31:0>.n240 VSS -1.78f
C4144 hgu_cdac_8bit_array_3.drv<31:0>.n241 VSS -1.78f
C4145 hgu_cdac_8bit_array_3.drv<31:0>.n242 VSS -1.11f
C4146 hgu_cdac_8bit_array_3.drv<31:0>.n243 VSS -1.74f
C4147 hgu_cdac_8bit_array_3.drv<31:0>.n244 VSS 4f
C4148 hgu_cdac_8bit_array_3.drv<31:0>.t7 VSS 0.0528f
C4149 hgu_cdac_8bit_array_3.drv<31:0>.t47 VSS 0.0528f
C4150 hgu_cdac_8bit_array_3.drv<31:0>.n245 VSS 0.39f
C4151 hgu_cdac_8bit_array_3.drv<31:0>.t19 VSS 0.106f
C4152 hgu_cdac_8bit_array_3.drv<31:0>.t29 VSS 0.106f
C4153 hgu_cdac_8bit_array_3.drv<31:0>.n246 VSS 0.804f
C4154 hgu_cdac_8bit_array_3.drv<31:0>.n247 VSS 0.439f
C4155 hgu_cdac_8bit_array_3.drv<31:0>.t58 VSS 0.0528f
C4156 hgu_cdac_8bit_array_3.drv<31:0>.t61 VSS 0.0528f
C4157 hgu_cdac_8bit_array_3.drv<31:0>.n248 VSS 0.39f
C4158 hgu_cdac_8bit_array_3.drv<31:0>.t25 VSS 0.106f
C4159 hgu_cdac_8bit_array_3.drv<31:0>.t28 VSS 0.106f
C4160 hgu_cdac_8bit_array_3.drv<31:0>.n249 VSS 0.804f
C4161 hgu_cdac_8bit_array_3.drv<31:0>.n250 VSS 0.496f
C4162 hgu_cdac_8bit_array_3.drv<31:0>.t13 VSS 0.0528f
C4163 hgu_cdac_8bit_array_3.drv<31:0>.t1 VSS 0.0528f
C4164 hgu_cdac_8bit_array_3.drv<31:0>.n251 VSS 0.39f
C4165 hgu_cdac_8bit_array_3.drv<31:0>.t42 VSS 0.106f
C4166 hgu_cdac_8bit_array_3.drv<31:0>.t45 VSS 0.106f
C4167 hgu_cdac_8bit_array_3.drv<31:0>.n252 VSS 0.804f
C4168 hgu_cdac_8bit_array_3.drv<31:0>.n253 VSS 0.402f
C4169 hgu_cdac_8bit_array_3.drv<31:0>.n254 VSS 3.6f
C4170 hgu_cdac_8bit_array_3.drv<31:0>.n255 VSS 8.26f
C4171 hgu_cdac_8bit_array_3.drv<31:0>.t0 VSS 0.0528f
C4172 hgu_cdac_8bit_array_3.drv<31:0>.t63 VSS 0.0528f
C4173 hgu_cdac_8bit_array_3.drv<31:0>.n256 VSS 0.372f
C4174 hgu_cdac_8bit_array_3.drv<31:0>.t44 VSS 0.106f
C4175 hgu_cdac_8bit_array_3.drv<31:0>.t23 VSS 0.106f
C4176 hgu_cdac_8bit_array_3.drv<31:0>.n257 VSS 0.759f
C4177 hgu_cdac_8bit_array_3.drv<31:0>.t52 VSS 0.0528f
C4178 hgu_cdac_8bit_array_3.drv<31:0>.t5 VSS 0.0528f
C4179 hgu_cdac_8bit_array_3.drv<31:0>.n258 VSS 0.39f
C4180 hgu_cdac_8bit_array_3.drv<31:0>.t34 VSS 0.106f
C4181 hgu_cdac_8bit_array_3.drv<31:0>.t17 VSS 0.106f
C4182 hgu_cdac_8bit_array_3.drv<31:0>.n259 VSS 0.802f
C4183 hgu_cdac_8bit_array_3.drv<31:0>.n260 VSS -2.09f
C4184 hgu_cdac_8bit_array_3.drv<31:0>.n261 VSS -1.78f
C4185 hgu_cdac_8bit_array_3.drv<31:0>.n262 VSS -1.11f
C4186 hgu_cdac_8bit_array_3.drv<31:0>.n263 VSS -1.74f
C4187 hgu_cdac_8bit_array_3.drv<31:0>.n264 VSS 4f
C4188 hgu_cdac_8bit_array_3.drv<31:0>.n265 VSS 8.26f
C4189 hgu_cdac_8bit_array_3.drv<31:0>.n266 VSS 11.6f
C4190 hgu_cdac_8bit_array_3.drv<31:0>.n267 VSS 1.12f
C4191 hgu_cdac_8bit_array_3.drv<31:0>.n268 VSS 0.147f
C4192 hgu_cdac_8bit_array_3.drv<31:0>.n269 VSS 0.147f
C4193 hgu_cdac_8bit_array_3.drv<31:0>.n270 VSS 0.651f
C4194 hgu_cdac_8bit_array_3.drv<31:0>.n271 VSS -0.465f
C4195 hgu_cdac_8bit_array_3.drv<31:0>.n272 VSS -1.74f
C4196 hgu_cdac_8bit_array_3.drv<31:0>.n273 VSS 4.41f
C4197 hgu_cdac_8bit_array_3.drv<31:0>.n274 VSS -1.74f
C4198 hgu_cdac_8bit_array_3.drv<31:0>.n275 VSS -0.465f
C4199 hgu_cdac_8bit_array_3.drv<31:0>.n276 VSS 0.61f
C4200 hgu_cdac_8bit_array_3.drv<31:0>.n277 VSS 0.147f
C4201 hgu_cdac_8bit_array_3.drv<31:0>.n278 VSS 0.147f
C4202 hgu_cdac_8bit_array_3.drv<31:0>.n279 VSS 0.651f
C4203 hgu_cdac_8bit_array_3.drv<31:0>.n280 VSS -0.465f
C4204 hgu_cdac_8bit_array_3.drv<31:0>.n281 VSS -1.74f
C4205 hgu_cdac_8bit_array_3.drv<31:0>.n282 VSS 4.41f
C4206 hgu_cdac_8bit_array_3.drv<31:0>.n283 VSS -1.74f
C4207 hgu_cdac_8bit_array_3.drv<31:0>.n284 VSS -0.465f
C4208 hgu_cdac_8bit_array_3.drv<31:0>.n285 VSS 0.61f
C4209 hgu_cdac_8bit_array_3.drv<31:0>.n286 VSS 0.147f
C4210 hgu_cdac_8bit_array_3.drv<31:0>.n287 VSS 0.147f
C4211 hgu_cdac_8bit_array_3.drv<31:0>.n288 VSS 0.651f
C4212 hgu_cdac_8bit_array_3.drv<31:0>.n289 VSS -0.465f
C4213 hgu_cdac_8bit_array_3.drv<31:0>.n290 VSS -1.78f
C4214 d<5>.t10 VSS 0.00914f
C4215 d<5>.t60 VSS 0.0174f
C4216 d<5>.t38 VSS 0.00914f
C4217 d<5>.t23 VSS 0.0174f
C4218 d<5>.t59 VSS 0.00914f
C4219 d<5>.t47 VSS 0.0174f
C4220 d<5>.t18 VSS 0.00914f
C4221 d<5>.t4 VSS 0.0174f
C4222 d<5>.t49 VSS 0.00914f
C4223 d<5>.t37 VSS 0.0174f
C4224 d<5>.t55 VSS 0.00914f
C4225 d<5>.t43 VSS 0.0174f
C4226 d<5>.t16 VSS 0.00914f
C4227 d<5>.t2 VSS 0.0174f
C4228 d<5>.t25 VSS 0.00914f
C4229 d<5>.t8 VSS 0.0174f
C4230 d<5>.t48 VSS 0.00914f
C4231 d<5>.t35 VSS 0.0174f
C4232 d<5>.t5 VSS 0.00914f
C4233 d<5>.t57 VSS 0.0174f
C4234 d<5>.t13 VSS 0.00914f
C4235 d<5>.t63 VSS 0.0174f
C4236 d<5>.t45 VSS 0.00914f
C4237 d<5>.t30 VSS 0.0174f
C4238 d<5>.t3 VSS 0.00914f
C4239 d<5>.t54 VSS 0.0174f
C4240 d<5>.t27 VSS 0.00914f
C4241 d<5>.t12 VSS 0.0174f
C4242 d<5>.t36 VSS 0.00914f
C4243 d<5>.t21 VSS 0.0174f
C4244 d<5>.t42 VSS 0.00914f
C4245 d<5>.t29 VSS 0.0174f
C4246 d<5>.t1 VSS 0.00914f
C4247 d<5>.t52 VSS 0.0174f
C4248 d<5>.t26 VSS 0.00914f
C4249 d<5>.t9 VSS 0.0174f
C4250 d<5>.t34 VSS 0.00914f
C4251 d<5>.t20 VSS 0.0174f
C4252 d<5>.t14 VSS 0.00914f
C4253 d<5>.t0 VSS 0.0174f
C4254 d<5>.t22 VSS 0.00914f
C4255 d<5>.t7 VSS 0.0174f
C4256 d<5>.t46 VSS 0.00914f
C4257 d<5>.t32 VSS 0.0174f
C4258 d<5>.t53 VSS 0.00914f
C4259 d<5>.t41 VSS 0.0174f
C4260 d<5>.t11 VSS 0.00914f
C4261 d<5>.t61 VSS 0.0174f
C4262 d<5>.t39 VSS 0.00914f
C4263 d<5>.t24 VSS 0.0174f
C4264 d<5>.t28 VSS 0.00914f
C4265 d<5>.t15 VSS 0.0174f
C4266 d<5>.t51 VSS 0.00914f
C4267 d<5>.t40 VSS 0.0174f
C4268 d<5>.t33 VSS 0.00914f
C4269 d<5>.t19 VSS 0.0174f
C4270 d<5>.t56 VSS 0.00914f
C4271 d<5>.t44 VSS 0.0174f
C4272 d<5>.t62 VSS 0.00914f
C4273 d<5>.t50 VSS 0.0174f
C4274 d<5>.t6 VSS 0.00914f
C4275 d<5>.t58 VSS 0.0174f
C4276 d<5>.t31 VSS 0.00914f
C4277 d<5>.t17 VSS 0.0174f
C4278 d<5>.n0 VSS 0.0339f
C4279 d<5>.n1 VSS 0.0395f
C4280 d<5>.n2 VSS 0.0395f
C4281 d<5>.n3 VSS 0.0395f
C4282 d<5>.n4 VSS 0.0395f
C4283 d<5>.n5 VSS 0.0395f
C4284 d<5>.n6 VSS 0.0395f
C4285 d<5>.n7 VSS 0.0395f
C4286 d<5>.n8 VSS 0.0395f
C4287 d<5>.n9 VSS 0.0395f
C4288 d<5>.n10 VSS 0.0395f
C4289 d<5>.n11 VSS 0.0395f
C4290 d<5>.n12 VSS 0.0395f
C4291 d<5>.n13 VSS 0.0395f
C4292 d<5>.n14 VSS 0.0395f
C4293 d<5>.n15 VSS 0.0395f
C4294 d<5>.n16 VSS 0.0395f
C4295 d<5>.n17 VSS 0.0395f
C4296 d<5>.n18 VSS 0.0395f
C4297 d<5>.n19 VSS 0.0395f
C4298 d<5>.n20 VSS 0.0395f
C4299 d<5>.n21 VSS 0.0395f
C4300 d<5>.n22 VSS 0.0395f
C4301 d<5>.n23 VSS 0.0395f
C4302 d<5>.n24 VSS 0.0395f
C4303 d<5>.n25 VSS 0.0395f
C4304 d<5>.n26 VSS 0.0395f
C4305 d<5>.n27 VSS 0.0395f
C4306 d<5>.n28 VSS 0.0395f
C4307 d<5>.n29 VSS 0.0395f
C4308 d<5>.n30 VSS 0.0395f
C4309 d<5>.n31 VSS 0.0306f
C4310 hgu_cdac_8bit_array_3.drv<63:0>.n0 VSS 4.24f
C4311 hgu_cdac_8bit_array_3.drv<63:0>.n1 VSS -1.85f
C4312 hgu_cdac_8bit_array_3.drv<63:0>.n2 VSS -1.17f
C4313 hgu_cdac_8bit_array_3.drv<63:0>.n3 VSS -1.88f
C4314 hgu_cdac_8bit_array_3.drv<63:0>.n4 VSS -1.88f
C4315 hgu_cdac_8bit_array_3.drv<63:0>.n5 VSS -1.17f
C4316 hgu_cdac_8bit_array_3.drv<63:0>.n6 VSS -1.85f
C4317 hgu_cdac_8bit_array_3.drv<63:0>.n7 VSS 6.55f
C4318 hgu_cdac_8bit_array_3.drv<63:0>.n8 VSS -1.85f
C4319 hgu_cdac_8bit_array_3.drv<63:0>.n9 VSS -1.17f
C4320 hgu_cdac_8bit_array_3.drv<63:0>.n10 VSS -1.88f
C4321 hgu_cdac_8bit_array_3.drv<63:0>.n11 VSS -1.88f
C4322 hgu_cdac_8bit_array_3.drv<63:0>.n12 VSS -1.17f
C4323 hgu_cdac_8bit_array_3.drv<63:0>.n13 VSS -1.85f
C4324 hgu_cdac_8bit_array_3.drv<63:0>.n14 VSS 6.55f
C4325 hgu_cdac_8bit_array_3.drv<63:0>.n15 VSS -1.85f
C4326 hgu_cdac_8bit_array_3.drv<63:0>.n16 VSS -1.17f
C4327 hgu_cdac_8bit_array_3.drv<63:0>.n17 VSS -1.88f
C4328 hgu_cdac_8bit_array_3.drv<63:0>.n18 VSS -1.88f
C4329 hgu_cdac_8bit_array_3.drv<63:0>.n19 VSS -1.17f
C4330 hgu_cdac_8bit_array_3.drv<63:0>.n20 VSS -1.85f
C4331 hgu_cdac_8bit_array_3.drv<63:0>.n21 VSS 6.55f
C4332 hgu_cdac_8bit_array_3.drv<63:0>.n22 VSS -1.85f
C4333 hgu_cdac_8bit_array_3.drv<63:0>.n23 VSS -1.17f
C4334 hgu_cdac_8bit_array_3.drv<63:0>.n24 VSS -1.88f
C4335 hgu_cdac_8bit_array_3.drv<63:0>.n25 VSS -1.88f
C4336 hgu_cdac_8bit_array_3.drv<63:0>.n26 VSS -1.17f
C4337 hgu_cdac_8bit_array_3.drv<63:0>.n27 VSS -1.85f
C4338 hgu_cdac_8bit_array_3.drv<63:0>.n28 VSS 6.55f
C4339 hgu_cdac_8bit_array_3.drv<63:0>.n29 VSS -1.63f
C4340 hgu_cdac_8bit_array_3.drv<63:0>.n30 VSS -1.85f
C4341 hgu_cdac_8bit_array_3.drv<63:0>.n31 VSS 6.55f
C4342 hgu_cdac_8bit_array_3.drv<63:0>.n32 VSS 4.93f
C4343 hgu_cdac_8bit_array_3.drv<63:0>.n33 VSS 0.79f
C4344 hgu_cdac_8bit_array_3.drv<63:0>.n34 VSS -0.492f
C4345 hgu_cdac_8bit_array_3.drv<63:0>.n35 VSS -1.85f
C4346 hgu_cdac_8bit_array_3.drv<63:0>.n36 VSS 6.56f
C4347 hgu_cdac_8bit_array_3.drv<63:0>.n37 VSS -1.85f
C4348 hgu_cdac_8bit_array_3.drv<63:0>.n38 VSS -0.492f
C4349 hgu_cdac_8bit_array_3.drv<63:0>.n39 VSS 0.69f
C4350 hgu_cdac_8bit_array_3.drv<63:0>.n40 VSS 0.156f
C4351 hgu_cdac_8bit_array_3.drv<63:0>.n41 VSS 0.156f
C4352 hgu_cdac_8bit_array_3.drv<63:0>.n42 VSS 0.646f
C4353 hgu_cdac_8bit_array_3.drv<63:0>.n43 VSS -0.492f
C4354 hgu_cdac_8bit_array_3.drv<63:0>.n44 VSS -1.85f
C4355 hgu_cdac_8bit_array_3.drv<63:0>.n45 VSS 6.56f
C4356 hgu_cdac_8bit_array_3.drv<63:0>.n46 VSS -1.85f
C4357 hgu_cdac_8bit_array_3.drv<63:0>.n47 VSS -0.492f
C4358 hgu_cdac_8bit_array_3.drv<63:0>.n48 VSS 0.69f
C4359 hgu_cdac_8bit_array_3.drv<63:0>.n49 VSS 0.156f
C4360 hgu_cdac_8bit_array_3.drv<63:0>.n50 VSS 0.156f
C4361 hgu_cdac_8bit_array_3.drv<63:0>.n51 VSS 0.646f
C4362 hgu_cdac_8bit_array_3.drv<63:0>.n52 VSS -0.492f
C4363 hgu_cdac_8bit_array_3.drv<63:0>.n53 VSS -1.85f
C4364 hgu_cdac_8bit_array_3.drv<63:0>.n54 VSS 6.56f
C4365 hgu_cdac_8bit_array_3.drv<63:0>.n55 VSS -1.85f
C4366 hgu_cdac_8bit_array_3.drv<63:0>.n56 VSS -0.492f
C4367 hgu_cdac_8bit_array_3.drv<63:0>.n57 VSS 0.69f
C4368 hgu_cdac_8bit_array_3.drv<63:0>.n58 VSS 0.156f
C4369 hgu_cdac_8bit_array_3.drv<63:0>.n59 VSS 0.156f
C4370 hgu_cdac_8bit_array_3.drv<63:0>.n60 VSS 0.646f
C4371 hgu_cdac_8bit_array_3.drv<63:0>.n61 VSS -0.492f
C4372 hgu_cdac_8bit_array_3.drv<63:0>.n62 VSS -1.85f
C4373 hgu_cdac_8bit_array_3.drv<63:0>.n63 VSS 6.56f
C4374 hgu_cdac_8bit_array_3.drv<63:0>.n64 VSS -1.85f
C4375 hgu_cdac_8bit_array_3.drv<63:0>.n65 VSS -0.492f
C4376 hgu_cdac_8bit_array_3.drv<63:0>.n66 VSS 0.69f
C4377 hgu_cdac_8bit_array_3.drv<63:0>.n67 VSS 0.156f
C4378 hgu_cdac_8bit_array_3.drv<63:0>.n68 VSS 0.156f
C4379 hgu_cdac_8bit_array_3.drv<63:0>.n69 VSS 0.646f
C4380 hgu_cdac_8bit_array_3.drv<63:0>.n70 VSS -0.492f
C4381 hgu_cdac_8bit_array_3.drv<63:0>.n71 VSS -1.85f
C4382 hgu_cdac_8bit_array_3.drv<63:0>.n72 VSS 6.56f
C4383 hgu_cdac_8bit_array_3.drv<63:0>.n73 VSS -1.85f
C4384 hgu_cdac_8bit_array_3.drv<63:0>.n74 VSS -0.492f
C4385 hgu_cdac_8bit_array_3.drv<63:0>.n75 VSS 0.69f
C4386 hgu_cdac_8bit_array_3.drv<63:0>.n76 VSS 0.156f
C4387 hgu_cdac_8bit_array_3.drv<63:0>.n77 VSS 0.156f
C4388 hgu_cdac_8bit_array_3.drv<63:0>.n78 VSS 0.646f
C4389 hgu_cdac_8bit_array_3.drv<63:0>.n79 VSS -0.492f
C4390 hgu_cdac_8bit_array_3.drv<63:0>.n80 VSS -1.85f
C4391 hgu_cdac_8bit_array_3.drv<63:0>.n81 VSS -6.63f
C4392 hgu_cdac_8bit_array_3.drv<63:0>.n82 VSS -1.85f
C4393 hgu_cdac_8bit_array_3.drv<63:0>.n83 VSS -1.17f
C4394 hgu_cdac_8bit_array_3.drv<63:0>.n84 VSS -1.88f
C4395 hgu_cdac_8bit_array_3.drv<63:0>.n85 VSS -1.88f
C4396 hgu_cdac_8bit_array_3.drv<63:0>.n86 VSS -1.17f
C4397 hgu_cdac_8bit_array_3.drv<63:0>.n87 VSS -1.85f
C4398 hgu_cdac_8bit_array_3.drv<63:0>.n88 VSS 6.55f
C4399 hgu_cdac_8bit_array_3.drv<63:0>.n89 VSS -1.85f
C4400 hgu_cdac_8bit_array_3.drv<63:0>.n90 VSS -1.17f
C4401 hgu_cdac_8bit_array_3.drv<63:0>.n91 VSS -1.88f
C4402 hgu_cdac_8bit_array_3.drv<63:0>.n92 VSS -1.88f
C4403 hgu_cdac_8bit_array_3.drv<63:0>.n93 VSS -1.17f
C4404 hgu_cdac_8bit_array_3.drv<63:0>.n94 VSS -1.85f
C4405 hgu_cdac_8bit_array_3.drv<63:0>.n95 VSS 6.55f
C4406 hgu_cdac_8bit_array_3.drv<63:0>.n96 VSS -1.85f
C4407 hgu_cdac_8bit_array_3.drv<63:0>.n97 VSS -1.17f
C4408 hgu_cdac_8bit_array_3.drv<63:0>.n98 VSS -1.88f
C4409 hgu_cdac_8bit_array_3.drv<63:0>.n99 VSS -1.88f
C4410 hgu_cdac_8bit_array_3.drv<63:0>.n100 VSS -1.17f
C4411 hgu_cdac_8bit_array_3.drv<63:0>.n101 VSS -1.85f
C4412 hgu_cdac_8bit_array_3.drv<63:0>.n102 VSS 6.55f
C4413 hgu_cdac_8bit_array_3.drv<63:0>.n103 VSS -1.85f
C4414 hgu_cdac_8bit_array_3.drv<63:0>.n104 VSS -1.17f
C4415 hgu_cdac_8bit_array_3.drv<63:0>.n105 VSS -1.88f
C4416 hgu_cdac_8bit_array_3.drv<63:0>.n106 VSS -1.88f
C4417 hgu_cdac_8bit_array_3.drv<63:0>.n107 VSS -1.17f
C4418 hgu_cdac_8bit_array_3.drv<63:0>.n108 VSS -1.85f
C4419 hgu_cdac_8bit_array_3.drv<63:0>.n109 VSS 6.55f
C4420 hgu_cdac_8bit_array_3.drv<63:0>.n110 VSS -1.85f
C4421 hgu_cdac_8bit_array_3.drv<63:0>.n111 VSS -1.17f
C4422 hgu_cdac_8bit_array_3.drv<63:0>.n112 VSS -1.88f
C4423 hgu_cdac_8bit_array_3.drv<63:0>.n113 VSS -1.88f
C4424 hgu_cdac_8bit_array_3.drv<63:0>.n114 VSS -1.17f
C4425 hgu_cdac_8bit_array_3.drv<63:0>.n115 VSS -1.85f
C4426 hgu_cdac_8bit_array_3.drv<63:0>.n116 VSS 6.55f
C4427 hgu_cdac_8bit_array_3.drv<63:0>.n117 VSS -1.85f
C4428 hgu_cdac_8bit_array_3.drv<63:0>.n118 VSS -1.17f
C4429 hgu_cdac_8bit_array_3.drv<63:0>.n119 VSS -1.88f
C4430 hgu_cdac_8bit_array_3.drv<63:0>.n120 VSS -1.88f
C4431 hgu_cdac_8bit_array_3.drv<63:0>.n121 VSS -1.17f
C4432 hgu_cdac_8bit_array_3.drv<63:0>.n122 VSS -1.85f
C4433 hgu_cdac_8bit_array_3.drv<63:0>.n123 VSS 6.55f
C4434 hgu_cdac_8bit_array_3.drv<63:0>.n124 VSS -1.85f
C4435 hgu_cdac_8bit_array_3.drv<63:0>.n125 VSS -1.17f
C4436 hgu_cdac_8bit_array_3.drv<63:0>.n126 VSS -1.88f
C4437 hgu_cdac_8bit_array_3.drv<63:0>.n127 VSS -1.88f
C4438 hgu_cdac_8bit_array_3.drv<63:0>.n128 VSS -1.17f
C4439 hgu_cdac_8bit_array_3.drv<63:0>.n129 VSS -1.85f
C4440 hgu_cdac_8bit_array_3.drv<63:0>.n130 VSS 6.55f
C4441 hgu_cdac_8bit_array_3.drv<63:0>.n131 VSS -1.85f
C4442 hgu_cdac_8bit_array_3.drv<63:0>.n132 VSS -1.17f
C4443 hgu_cdac_8bit_array_3.drv<63:0>.n133 VSS -1.88f
C4444 hgu_cdac_8bit_array_3.drv<63:0>.n134 VSS -1.88f
C4445 hgu_cdac_8bit_array_3.drv<63:0>.n135 VSS -1.17f
C4446 hgu_cdac_8bit_array_3.drv<63:0>.n136 VSS -1.85f
C4447 hgu_cdac_8bit_array_3.drv<63:0>.n137 VSS 6.55f
C4448 hgu_cdac_8bit_array_3.drv<63:0>.n138 VSS -1.85f
C4449 hgu_cdac_8bit_array_3.drv<63:0>.n139 VSS -1.17f
C4450 hgu_cdac_8bit_array_3.drv<63:0>.n140 VSS -1.88f
C4451 hgu_cdac_8bit_array_3.drv<63:0>.n141 VSS -1.88f
C4452 hgu_cdac_8bit_array_3.drv<63:0>.n142 VSS -1.17f
C4453 hgu_cdac_8bit_array_3.drv<63:0>.n143 VSS -1.85f
C4454 hgu_cdac_8bit_array_3.drv<63:0>.n144 VSS 6.55f
C4455 hgu_cdac_8bit_array_3.drv<63:0>.n145 VSS -1.85f
C4456 hgu_cdac_8bit_array_3.drv<63:0>.n146 VSS -1.17f
C4457 hgu_cdac_8bit_array_3.drv<63:0>.n147 VSS -1.88f
C4458 hgu_cdac_8bit_array_3.drv<63:0>.n148 VSS -1.88f
C4459 hgu_cdac_8bit_array_3.drv<63:0>.n149 VSS -1.17f
C4460 hgu_cdac_8bit_array_3.drv<63:0>.n150 VSS -1.85f
C4461 hgu_cdac_8bit_array_3.drv<63:0>.n151 VSS 6.55f
C4462 hgu_cdac_8bit_array_3.drv<63:0>.n152 VSS -1.85f
C4463 hgu_cdac_8bit_array_3.drv<63:0>.n153 VSS -1.17f
C4464 hgu_cdac_8bit_array_3.drv<63:0>.n154 VSS -1.88f
C4465 hgu_cdac_8bit_array_3.drv<63:0>.n155 VSS -1.88f
C4466 hgu_cdac_8bit_array_3.drv<63:0>.n156 VSS -1.17f
C4467 hgu_cdac_8bit_array_3.drv<63:0>.n157 VSS -1.85f
C4468 hgu_cdac_8bit_array_3.drv<63:0>.n158 VSS 6.55f
C4469 hgu_cdac_8bit_array_3.drv<63:0>.t101 VSS 0.0559f
C4470 hgu_cdac_8bit_array_3.drv<63:0>.t98 VSS 0.0559f
C4471 hgu_cdac_8bit_array_3.drv<63:0>.n159 VSS 0.413f
C4472 hgu_cdac_8bit_array_3.drv<63:0>.t73 VSS 0.112f
C4473 hgu_cdac_8bit_array_3.drv<63:0>.t65 VSS 0.112f
C4474 hgu_cdac_8bit_array_3.drv<63:0>.n160 VSS 0.852f
C4475 hgu_cdac_8bit_array_3.drv<63:0>.n161 VSS 4.13f
C4476 hgu_cdac_8bit_array_3.drv<63:0>.n162 VSS -1.85f
C4477 hgu_cdac_8bit_array_3.drv<63:0>.n163 VSS -1.17f
C4478 hgu_cdac_8bit_array_3.drv<63:0>.n164 VSS -1.88f
C4479 hgu_cdac_8bit_array_3.drv<63:0>.n165 VSS -1.88f
C4480 hgu_cdac_8bit_array_3.drv<63:0>.n166 VSS -1.17f
C4481 hgu_cdac_8bit_array_3.drv<63:0>.n167 VSS -1.85f
C4482 hgu_cdac_8bit_array_3.drv<63:0>.n168 VSS 4.23f
C4483 hgu_cdac_8bit_array_3.drv<63:0>.n169 VSS 9.01f
C4484 hgu_cdac_8bit_array_3.drv<63:0>.n170 VSS -1.85f
C4485 hgu_cdac_8bit_array_3.drv<63:0>.n171 VSS -1.17f
C4486 hgu_cdac_8bit_array_3.drv<63:0>.n172 VSS -1.88f
C4487 hgu_cdac_8bit_array_3.drv<63:0>.n173 VSS -1.88f
C4488 hgu_cdac_8bit_array_3.drv<63:0>.n174 VSS -1.17f
C4489 hgu_cdac_8bit_array_3.drv<63:0>.n175 VSS -1.85f
C4490 hgu_cdac_8bit_array_3.drv<63:0>.n176 VSS 4.23f
C4491 hgu_cdac_8bit_array_3.drv<63:0>.t112 VSS 0.0559f
C4492 hgu_cdac_8bit_array_3.drv<63:0>.t118 VSS 0.0559f
C4493 hgu_cdac_8bit_array_3.drv<63:0>.n177 VSS 0.413f
C4494 hgu_cdac_8bit_array_3.drv<63:0>.t28 VSS 0.112f
C4495 hgu_cdac_8bit_array_3.drv<63:0>.t53 VSS 0.112f
C4496 hgu_cdac_8bit_array_3.drv<63:0>.n178 VSS 0.852f
C4497 hgu_cdac_8bit_array_3.drv<63:0>.n179 VSS 0.467f
C4498 hgu_cdac_8bit_array_3.drv<63:0>.t7 VSS 0.0559f
C4499 hgu_cdac_8bit_array_3.drv<63:0>.t111 VSS 0.0559f
C4500 hgu_cdac_8bit_array_3.drv<63:0>.n180 VSS 0.413f
C4501 hgu_cdac_8bit_array_3.drv<63:0>.t79 VSS 0.112f
C4502 hgu_cdac_8bit_array_3.drv<63:0>.t41 VSS 0.112f
C4503 hgu_cdac_8bit_array_3.drv<63:0>.n181 VSS 0.852f
C4504 hgu_cdac_8bit_array_3.drv<63:0>.t1 VSS 0.0559f
C4505 hgu_cdac_8bit_array_3.drv<63:0>.t23 VSS 0.0559f
C4506 hgu_cdac_8bit_array_3.drv<63:0>.n182 VSS 0.413f
C4507 hgu_cdac_8bit_array_3.drv<63:0>.t49 VSS 0.112f
C4508 hgu_cdac_8bit_array_3.drv<63:0>.t70 VSS 0.112f
C4509 hgu_cdac_8bit_array_3.drv<63:0>.n183 VSS 0.852f
C4510 hgu_cdac_8bit_array_3.drv<63:0>.n184 VSS 0.527f
C4511 hgu_cdac_8bit_array_3.drv<63:0>.n185 VSS 0.424f
C4512 hgu_cdac_8bit_array_3.drv<63:0>.n186 VSS 3.86f
C4513 hgu_cdac_8bit_array_3.drv<63:0>.n187 VSS 8.79f
C4514 hgu_cdac_8bit_array_3.drv<63:0>.n188 VSS -1.85f
C4515 hgu_cdac_8bit_array_3.drv<63:0>.n189 VSS -1.17f
C4516 hgu_cdac_8bit_array_3.drv<63:0>.n190 VSS -1.88f
C4517 hgu_cdac_8bit_array_3.drv<63:0>.n191 VSS -1.88f
C4518 hgu_cdac_8bit_array_3.drv<63:0>.n192 VSS -1.17f
C4519 hgu_cdac_8bit_array_3.drv<63:0>.n193 VSS -1.85f
C4520 hgu_cdac_8bit_array_3.drv<63:0>.n194 VSS 4.23f
C4521 hgu_cdac_8bit_array_3.drv<63:0>.t5 VSS 0.0559f
C4522 hgu_cdac_8bit_array_3.drv<63:0>.t20 VSS 0.0559f
C4523 hgu_cdac_8bit_array_3.drv<63:0>.n195 VSS 0.395f
C4524 hgu_cdac_8bit_array_3.drv<63:0>.t77 VSS 0.112f
C4525 hgu_cdac_8bit_array_3.drv<63:0>.t39 VSS 0.112f
C4526 hgu_cdac_8bit_array_3.drv<63:0>.n196 VSS 0.803f
C4527 hgu_cdac_8bit_array_3.drv<63:0>.t95 VSS 0.0559f
C4528 hgu_cdac_8bit_array_3.drv<63:0>.t21 VSS 0.0559f
C4529 hgu_cdac_8bit_array_3.drv<63:0>.n197 VSS 0.413f
C4530 hgu_cdac_8bit_array_3.drv<63:0>.t62 VSS 0.112f
C4531 hgu_cdac_8bit_array_3.drv<63:0>.t67 VSS 0.112f
C4532 hgu_cdac_8bit_array_3.drv<63:0>.n198 VSS 0.852f
C4533 hgu_cdac_8bit_array_3.drv<63:0>.n199 VSS 0.526f
C4534 hgu_cdac_8bit_array_3.drv<63:0>.n200 VSS 8.79f
C4535 hgu_cdac_8bit_array_3.drv<63:0>.t125 VSS 0.0559f
C4536 hgu_cdac_8bit_array_3.drv<63:0>.t12 VSS 0.0559f
C4537 hgu_cdac_8bit_array_3.drv<63:0>.n201 VSS 0.413f
C4538 hgu_cdac_8bit_array_3.drv<63:0>.t36 VSS 0.112f
C4539 hgu_cdac_8bit_array_3.drv<63:0>.t59 VSS 0.112f
C4540 hgu_cdac_8bit_array_3.drv<63:0>.n202 VSS 0.852f
C4541 hgu_cdac_8bit_array_3.drv<63:0>.n203 VSS 0.426f
C4542 hgu_cdac_8bit_array_3.drv<63:0>.t9 VSS 0.0559f
C4543 hgu_cdac_8bit_array_3.drv<63:0>.t93 VSS 0.0559f
C4544 hgu_cdac_8bit_array_3.drv<63:0>.n204 VSS 0.413f
C4545 hgu_cdac_8bit_array_3.drv<63:0>.t81 VSS 0.112f
C4546 hgu_cdac_8bit_array_3.drv<63:0>.t26 VSS 0.112f
C4547 hgu_cdac_8bit_array_3.drv<63:0>.n205 VSS 0.852f
C4548 hgu_cdac_8bit_array_3.drv<63:0>.n206 VSS 0.464f
C4549 hgu_cdac_8bit_array_3.drv<63:0>.n207 VSS 3.86f
C4550 hgu_cdac_8bit_array_3.drv<63:0>.n208 VSS -1.85f
C4551 hgu_cdac_8bit_array_3.drv<63:0>.n209 VSS -1.17f
C4552 hgu_cdac_8bit_array_3.drv<63:0>.n210 VSS -1.88f
C4553 hgu_cdac_8bit_array_3.drv<63:0>.n211 VSS -1.88f
C4554 hgu_cdac_8bit_array_3.drv<63:0>.n212 VSS -1.17f
C4555 hgu_cdac_8bit_array_3.drv<63:0>.n213 VSS -1.85f
C4556 hgu_cdac_8bit_array_3.drv<63:0>.n214 VSS 4.23f
C4557 hgu_cdac_8bit_array_3.drv<63:0>.n215 VSS 8.79f
C4558 hgu_cdac_8bit_array_3.drv<63:0>.t123 VSS 0.0559f
C4559 hgu_cdac_8bit_array_3.drv<63:0>.t10 VSS 0.0559f
C4560 hgu_cdac_8bit_array_3.drv<63:0>.n216 VSS 0.413f
C4561 hgu_cdac_8bit_array_3.drv<63:0>.t34 VSS 0.112f
C4562 hgu_cdac_8bit_array_3.drv<63:0>.t57 VSS 0.112f
C4563 hgu_cdac_8bit_array_3.drv<63:0>.n217 VSS 0.852f
C4564 hgu_cdac_8bit_array_3.drv<63:0>.n218 VSS 0.496f
C4565 hgu_cdac_8bit_array_3.drv<63:0>.t8 VSS 0.0559f
C4566 hgu_cdac_8bit_array_3.drv<63:0>.t91 VSS 0.0559f
C4567 hgu_cdac_8bit_array_3.drv<63:0>.n219 VSS 0.395f
C4568 hgu_cdac_8bit_array_3.drv<63:0>.t80 VSS 0.112f
C4569 hgu_cdac_8bit_array_3.drv<63:0>.t88 VSS 0.112f
C4570 hgu_cdac_8bit_array_3.drv<63:0>.n220 VSS 0.802f
C4571 hgu_cdac_8bit_array_3.drv<63:0>.t22 VSS 0.0559f
C4572 hgu_cdac_8bit_array_3.drv<63:0>.t102 VSS 0.0559f
C4573 hgu_cdac_8bit_array_3.drv<63:0>.n221 VSS 0.413f
C4574 hgu_cdac_8bit_array_3.drv<63:0>.t68 VSS 0.112f
C4575 hgu_cdac_8bit_array_3.drv<63:0>.t74 VSS 0.112f
C4576 hgu_cdac_8bit_array_3.drv<63:0>.n222 VSS 0.852f
C4577 hgu_cdac_8bit_array_3.drv<63:0>.n223 VSS 0.536f
C4578 hgu_cdac_8bit_array_3.drv<63:0>.n224 VSS 0.457f
C4579 hgu_cdac_8bit_array_3.drv<63:0>.n225 VSS 3.9f
C4580 hgu_cdac_8bit_array_3.drv<63:0>.n226 VSS -1.85f
C4581 hgu_cdac_8bit_array_3.drv<63:0>.n227 VSS -1.17f
C4582 hgu_cdac_8bit_array_3.drv<63:0>.n228 VSS -1.88f
C4583 hgu_cdac_8bit_array_3.drv<63:0>.n229 VSS -1.88f
C4584 hgu_cdac_8bit_array_3.drv<63:0>.n230 VSS -1.17f
C4585 hgu_cdac_8bit_array_3.drv<63:0>.n231 VSS -1.85f
C4586 hgu_cdac_8bit_array_3.drv<63:0>.n232 VSS 4.23f
C4587 hgu_cdac_8bit_array_3.drv<63:0>.n233 VSS 8.79f
C4588 hgu_cdac_8bit_array_3.drv<63:0>.t107 VSS 0.0559f
C4589 hgu_cdac_8bit_array_3.drv<63:0>.t19 VSS 0.0559f
C4590 hgu_cdac_8bit_array_3.drv<63:0>.n234 VSS 0.395f
C4591 hgu_cdac_8bit_array_3.drv<63:0>.t84 VSS 0.112f
C4592 hgu_cdac_8bit_array_3.drv<63:0>.t46 VSS 0.112f
C4593 hgu_cdac_8bit_array_3.drv<63:0>.n235 VSS 0.803f
C4594 hgu_cdac_8bit_array_3.drv<63:0>.n236 VSS 0.429f
C4595 hgu_cdac_8bit_array_3.drv<63:0>.t99 VSS 0.0559f
C4596 hgu_cdac_8bit_array_3.drv<63:0>.t113 VSS 0.0559f
C4597 hgu_cdac_8bit_array_3.drv<63:0>.n237 VSS 0.413f
C4598 hgu_cdac_8bit_array_3.drv<63:0>.t66 VSS 0.112f
C4599 hgu_cdac_8bit_array_3.drv<63:0>.t29 VSS 0.112f
C4600 hgu_cdac_8bit_array_3.drv<63:0>.n238 VSS 0.852f
C4601 hgu_cdac_8bit_array_3.drv<63:0>.n239 VSS 0.508f
C4602 hgu_cdac_8bit_array_3.drv<63:0>.n240 VSS 3.85f
C4603 hgu_cdac_8bit_array_3.drv<63:0>.n241 VSS -1.85f
C4604 hgu_cdac_8bit_array_3.drv<63:0>.n242 VSS -1.17f
C4605 hgu_cdac_8bit_array_3.drv<63:0>.n243 VSS -1.88f
C4606 hgu_cdac_8bit_array_3.drv<63:0>.n244 VSS -1.88f
C4607 hgu_cdac_8bit_array_3.drv<63:0>.n245 VSS -1.17f
C4608 hgu_cdac_8bit_array_3.drv<63:0>.n246 VSS -1.85f
C4609 hgu_cdac_8bit_array_3.drv<63:0>.n247 VSS 4.23f
C4610 hgu_cdac_8bit_array_3.drv<63:0>.n248 VSS 8.79f
C4611 hgu_cdac_8bit_array_3.drv<63:0>.t105 VSS 0.0559f
C4612 hgu_cdac_8bit_array_3.drv<63:0>.t17 VSS 0.0559f
C4613 hgu_cdac_8bit_array_3.drv<63:0>.n249 VSS 0.413f
C4614 hgu_cdac_8bit_array_3.drv<63:0>.t82 VSS 0.112f
C4615 hgu_cdac_8bit_array_3.drv<63:0>.t44 VSS 0.112f
C4616 hgu_cdac_8bit_array_3.drv<63:0>.n250 VSS 0.852f
C4617 hgu_cdac_8bit_array_3.drv<63:0>.n251 VSS 0.442f
C4618 hgu_cdac_8bit_array_3.drv<63:0>.t90 VSS 0.0559f
C4619 hgu_cdac_8bit_array_3.drv<63:0>.t116 VSS 0.0559f
C4620 hgu_cdac_8bit_array_3.drv<63:0>.n252 VSS 0.413f
C4621 hgu_cdac_8bit_array_3.drv<63:0>.t87 VSS 0.112f
C4622 hgu_cdac_8bit_array_3.drv<63:0>.t32 VSS 0.112f
C4623 hgu_cdac_8bit_array_3.drv<63:0>.n253 VSS 0.852f
C4624 hgu_cdac_8bit_array_3.drv<63:0>.t120 VSS 0.0559f
C4625 hgu_cdac_8bit_array_3.drv<63:0>.t96 VSS 0.0559f
C4626 hgu_cdac_8bit_array_3.drv<63:0>.n254 VSS 0.413f
C4627 hgu_cdac_8bit_array_3.drv<63:0>.t55 VSS 0.112f
C4628 hgu_cdac_8bit_array_3.drv<63:0>.t63 VSS 0.112f
C4629 hgu_cdac_8bit_array_3.drv<63:0>.n255 VSS 0.852f
C4630 hgu_cdac_8bit_array_3.drv<63:0>.t109 VSS 0.0559f
C4631 hgu_cdac_8bit_array_3.drv<63:0>.t115 VSS 0.0559f
C4632 hgu_cdac_8bit_array_3.drv<63:0>.n256 VSS 0.413f
C4633 hgu_cdac_8bit_array_3.drv<63:0>.t86 VSS 0.112f
C4634 hgu_cdac_8bit_array_3.drv<63:0>.t31 VSS 0.112f
C4635 hgu_cdac_8bit_array_3.drv<63:0>.n257 VSS 0.852f
C4636 hgu_cdac_8bit_array_3.drv<63:0>.n258 VSS 0.524f
C4637 hgu_cdac_8bit_array_3.drv<63:0>.n259 VSS 0.524f
C4638 hgu_cdac_8bit_array_3.drv<63:0>.n260 VSS 0.448f
C4639 hgu_cdac_8bit_array_3.drv<63:0>.n261 VSS 3.87f
C4640 hgu_cdac_8bit_array_3.drv<63:0>.n262 VSS -1.85f
C4641 hgu_cdac_8bit_array_3.drv<63:0>.n263 VSS -1.17f
C4642 hgu_cdac_8bit_array_3.drv<63:0>.n264 VSS -1.88f
C4643 hgu_cdac_8bit_array_3.drv<63:0>.n265 VSS -1.88f
C4644 hgu_cdac_8bit_array_3.drv<63:0>.n266 VSS -1.17f
C4645 hgu_cdac_8bit_array_3.drv<63:0>.n267 VSS -1.85f
C4646 hgu_cdac_8bit_array_3.drv<63:0>.n268 VSS 4.23f
C4647 hgu_cdac_8bit_array_3.drv<63:0>.n269 VSS 8.79f
C4648 hgu_cdac_8bit_array_3.drv<63:0>.n270 VSS -1.85f
C4649 hgu_cdac_8bit_array_3.drv<63:0>.n271 VSS -1.17f
C4650 hgu_cdac_8bit_array_3.drv<63:0>.n272 VSS -1.88f
C4651 hgu_cdac_8bit_array_3.drv<63:0>.n273 VSS -1.88f
C4652 hgu_cdac_8bit_array_3.drv<63:0>.n274 VSS -1.17f
C4653 hgu_cdac_8bit_array_3.drv<63:0>.n275 VSS -1.85f
C4654 hgu_cdac_8bit_array_3.drv<63:0>.n276 VSS 2.58f
C4655 hgu_cdac_8bit_array_3.drv<63:0>.t16 VSS 0.0559f
C4656 hgu_cdac_8bit_array_3.drv<63:0>.t4 VSS 0.0559f
C4657 hgu_cdac_8bit_array_3.drv<63:0>.n277 VSS 0.395f
C4658 hgu_cdac_8bit_array_3.drv<63:0>.t43 VSS 0.112f
C4659 hgu_cdac_8bit_array_3.drv<63:0>.t51 VSS 0.112f
C4660 hgu_cdac_8bit_array_3.drv<63:0>.n278 VSS 0.803f
C4661 hgu_cdac_8bit_array_3.drv<63:0>.t119 VSS 0.0559f
C4662 hgu_cdac_8bit_array_3.drv<63:0>.t103 VSS 0.0559f
C4663 hgu_cdac_8bit_array_3.drv<63:0>.n279 VSS 0.413f
C4664 hgu_cdac_8bit_array_3.drv<63:0>.t54 VSS 0.112f
C4665 hgu_cdac_8bit_array_3.drv<63:0>.t75 VSS 0.112f
C4666 hgu_cdac_8bit_array_3.drv<63:0>.n280 VSS 0.852f
C4667 hgu_cdac_8bit_array_3.drv<63:0>.n281 VSS 0.53f
C4668 hgu_cdac_8bit_array_3.drv<63:0>.n282 VSS 0.457f
C4669 hgu_cdac_8bit_array_3.drv<63:0>.n283 VSS 3.7f
C4670 hgu_cdac_8bit_array_3.drv<63:0>.n284 VSS -1.85f
C4671 hgu_cdac_8bit_array_3.drv<63:0>.n285 VSS -1.17f
C4672 hgu_cdac_8bit_array_3.drv<63:0>.n286 VSS -1.88f
C4673 hgu_cdac_8bit_array_3.drv<63:0>.n287 VSS -1.88f
C4674 hgu_cdac_8bit_array_3.drv<63:0>.n288 VSS -1.17f
C4675 hgu_cdac_8bit_array_3.drv<63:0>.n289 VSS -1.85f
C4676 hgu_cdac_8bit_array_3.drv<63:0>.n290 VSS 4.23f
C4677 hgu_cdac_8bit_array_3.drv<63:0>.n291 VSS 8.9f
C4678 hgu_cdac_8bit_array_3.drv<63:0>.n292 VSS -1.85f
C4679 hgu_cdac_8bit_array_3.drv<63:0>.n293 VSS -1.17f
C4680 hgu_cdac_8bit_array_3.drv<63:0>.n294 VSS -1.88f
C4681 hgu_cdac_8bit_array_3.drv<63:0>.n295 VSS -1.88f
C4682 hgu_cdac_8bit_array_3.drv<63:0>.n296 VSS -1.17f
C4683 hgu_cdac_8bit_array_3.drv<63:0>.n297 VSS -1.85f
C4684 hgu_cdac_8bit_array_3.drv<63:0>.n298 VSS 4.23f
C4685 hgu_cdac_8bit_array_3.drv<63:0>.t100 VSS 0.0559f
C4686 hgu_cdac_8bit_array_3.drv<63:0>.t124 VSS 0.0559f
C4687 hgu_cdac_8bit_array_3.drv<63:0>.n299 VSS 0.413f
C4688 hgu_cdac_8bit_array_3.drv<63:0>.t72 VSS 0.112f
C4689 hgu_cdac_8bit_array_3.drv<63:0>.t35 VSS 0.112f
C4690 hgu_cdac_8bit_array_3.drv<63:0>.n300 VSS 0.852f
C4691 hgu_cdac_8bit_array_3.drv<63:0>.n301 VSS 0.548f
C4692 hgu_cdac_8bit_array_3.drv<63:0>.t15 VSS 0.0559f
C4693 hgu_cdac_8bit_array_3.drv<63:0>.t3 VSS 0.0559f
C4694 hgu_cdac_8bit_array_3.drv<63:0>.n302 VSS 0.413f
C4695 hgu_cdac_8bit_array_3.drv<63:0>.t42 VSS 0.112f
C4696 hgu_cdac_8bit_array_3.drv<63:0>.t50 VSS 0.112f
C4697 hgu_cdac_8bit_array_3.drv<63:0>.n303 VSS 0.852f
C4698 hgu_cdac_8bit_array_3.drv<63:0>.n304 VSS 0.457f
C4699 hgu_cdac_8bit_array_3.drv<63:0>.t25 VSS 0.0559f
C4700 hgu_cdac_8bit_array_3.drv<63:0>.t122 VSS 0.0559f
C4701 hgu_cdac_8bit_array_3.drv<63:0>.n305 VSS 0.413f
C4702 hgu_cdac_8bit_array_3.drv<63:0>.t71 VSS 0.112f
C4703 hgu_cdac_8bit_array_3.drv<63:0>.t33 VSS 0.112f
C4704 hgu_cdac_8bit_array_3.drv<63:0>.n306 VSS 0.852f
C4705 hgu_cdac_8bit_array_3.drv<63:0>.n307 VSS 0.449f
C4706 hgu_cdac_8bit_array_3.drv<63:0>.n308 VSS 3.85f
C4707 hgu_cdac_8bit_array_3.drv<63:0>.n309 VSS 8.79f
C4708 hgu_cdac_8bit_array_3.drv<63:0>.t14 VSS 0.0559f
C4709 hgu_cdac_8bit_array_3.drv<63:0>.t108 VSS 0.0559f
C4710 hgu_cdac_8bit_array_3.drv<63:0>.n310 VSS 0.413f
C4711 hgu_cdac_8bit_array_3.drv<63:0>.t61 VSS 0.112f
C4712 hgu_cdac_8bit_array_3.drv<63:0>.t85 VSS 0.112f
C4713 hgu_cdac_8bit_array_3.drv<63:0>.n311 VSS 0.852f
C4714 hgu_cdac_8bit_array_3.drv<63:0>.n312 VSS 0.517f
C4715 hgu_cdac_8bit_array_3.drv<63:0>.t114 VSS 0.0559f
C4716 hgu_cdac_8bit_array_3.drv<63:0>.t126 VSS 0.0559f
C4717 hgu_cdac_8bit_array_3.drv<63:0>.n313 VSS 0.395f
C4718 hgu_cdac_8bit_array_3.drv<63:0>.t30 VSS 0.112f
C4719 hgu_cdac_8bit_array_3.drv<63:0>.t37 VSS 0.112f
C4720 hgu_cdac_8bit_array_3.drv<63:0>.n314 VSS 0.803f
C4721 hgu_cdac_8bit_array_3.drv<63:0>.n315 VSS 0.339f
C4722 hgu_cdac_8bit_array_3.drv<63:0>.n316 VSS 3.83f
C4723 hgu_cdac_8bit_array_3.drv<63:0>.n317 VSS -1.85f
C4724 hgu_cdac_8bit_array_3.drv<63:0>.n318 VSS -1.17f
C4725 hgu_cdac_8bit_array_3.drv<63:0>.n319 VSS -1.88f
C4726 hgu_cdac_8bit_array_3.drv<63:0>.n320 VSS -1.88f
C4727 hgu_cdac_8bit_array_3.drv<63:0>.n321 VSS -1.17f
C4728 hgu_cdac_8bit_array_3.drv<63:0>.n322 VSS -1.85f
C4729 hgu_cdac_8bit_array_3.drv<63:0>.n323 VSS 4.23f
C4730 hgu_cdac_8bit_array_3.drv<63:0>.n324 VSS 8.79f
C4731 hgu_cdac_8bit_array_3.drv<63:0>.t13 VSS 0.0559f
C4732 hgu_cdac_8bit_array_3.drv<63:0>.t106 VSS 0.0559f
C4733 hgu_cdac_8bit_array_3.drv<63:0>.n325 VSS 0.413f
C4734 hgu_cdac_8bit_array_3.drv<63:0>.t60 VSS 0.112f
C4735 hgu_cdac_8bit_array_3.drv<63:0>.t83 VSS 0.112f
C4736 hgu_cdac_8bit_array_3.drv<63:0>.n326 VSS 0.852f
C4737 hgu_cdac_8bit_array_3.drv<63:0>.n327 VSS 0.6f
C4738 hgu_cdac_8bit_array_3.drv<63:0>.t18 VSS 0.0559f
C4739 hgu_cdac_8bit_array_3.drv<63:0>.t121 VSS 0.0559f
C4740 hgu_cdac_8bit_array_3.drv<63:0>.n328 VSS 0.413f
C4741 hgu_cdac_8bit_array_3.drv<63:0>.t45 VSS 0.112f
C4742 hgu_cdac_8bit_array_3.drv<63:0>.t56 VSS 0.112f
C4743 hgu_cdac_8bit_array_3.drv<63:0>.n329 VSS 0.852f
C4744 hgu_cdac_8bit_array_3.drv<63:0>.n330 VSS 0.419f
C4745 hgu_cdac_8bit_array_3.drv<63:0>.t6 VSS 0.0559f
C4746 hgu_cdac_8bit_array_3.drv<63:0>.t110 VSS 0.0559f
C4747 hgu_cdac_8bit_array_3.drv<63:0>.n331 VSS 0.413f
C4748 hgu_cdac_8bit_array_3.drv<63:0>.t78 VSS 0.112f
C4749 hgu_cdac_8bit_array_3.drv<63:0>.t40 VSS 0.112f
C4750 hgu_cdac_8bit_array_3.drv<63:0>.n332 VSS 0.852f
C4751 hgu_cdac_8bit_array_3.drv<63:0>.n333 VSS 0.518f
C4752 hgu_cdac_8bit_array_3.drv<63:0>.n334 VSS 3.82f
C4753 hgu_cdac_8bit_array_3.drv<63:0>.n335 VSS -1.85f
C4754 hgu_cdac_8bit_array_3.drv<63:0>.n336 VSS -1.17f
C4755 hgu_cdac_8bit_array_3.drv<63:0>.n337 VSS -1.88f
C4756 hgu_cdac_8bit_array_3.drv<63:0>.n338 VSS -1.88f
C4757 hgu_cdac_8bit_array_3.drv<63:0>.n339 VSS -1.17f
C4758 hgu_cdac_8bit_array_3.drv<63:0>.n340 VSS -1.85f
C4759 hgu_cdac_8bit_array_3.drv<63:0>.n341 VSS 4.23f
C4760 hgu_cdac_8bit_array_3.drv<63:0>.n342 VSS 8.79f
C4761 hgu_cdac_8bit_array_3.drv<63:0>.t2 VSS 0.0559f
C4762 hgu_cdac_8bit_array_3.drv<63:0>.t24 VSS 0.0559f
C4763 hgu_cdac_8bit_array_3.drv<63:0>.n343 VSS 0.413f
C4764 hgu_cdac_8bit_array_3.drv<63:0>.t48 VSS 0.112f
C4765 hgu_cdac_8bit_array_3.drv<63:0>.t69 VSS 0.112f
C4766 hgu_cdac_8bit_array_3.drv<63:0>.n344 VSS 0.852f
C4767 hgu_cdac_8bit_array_3.drv<63:0>.n345 VSS 0.474f
C4768 hgu_cdac_8bit_array_3.drv<63:0>.t104 VSS 0.0559f
C4769 hgu_cdac_8bit_array_3.drv<63:0>.t127 VSS 0.0559f
C4770 hgu_cdac_8bit_array_3.drv<63:0>.n346 VSS 0.413f
C4771 hgu_cdac_8bit_array_3.drv<63:0>.t76 VSS 0.112f
C4772 hgu_cdac_8bit_array_3.drv<63:0>.t38 VSS 0.112f
C4773 hgu_cdac_8bit_array_3.drv<63:0>.n347 VSS 0.852f
C4774 hgu_cdac_8bit_array_3.drv<63:0>.n348 VSS 0.419f
C4775 hgu_cdac_8bit_array_3.drv<63:0>.n349 VSS 3.86f
C4776 hgu_cdac_8bit_array_3.drv<63:0>.n350 VSS -1.85f
C4777 hgu_cdac_8bit_array_3.drv<63:0>.n351 VSS -1.17f
C4778 hgu_cdac_8bit_array_3.drv<63:0>.n352 VSS -1.88f
C4779 hgu_cdac_8bit_array_3.drv<63:0>.n353 VSS -1.88f
C4780 hgu_cdac_8bit_array_3.drv<63:0>.n354 VSS -1.17f
C4781 hgu_cdac_8bit_array_3.drv<63:0>.n355 VSS -1.85f
C4782 hgu_cdac_8bit_array_3.drv<63:0>.n356 VSS 4.23f
C4783 hgu_cdac_8bit_array_3.drv<63:0>.n357 VSS 8.79f
C4784 hgu_cdac_8bit_array_3.drv<63:0>.t0 VSS 0.0559f
C4785 hgu_cdac_8bit_array_3.drv<63:0>.t94 VSS 0.0559f
C4786 hgu_cdac_8bit_array_3.drv<63:0>.n358 VSS 0.413f
C4787 hgu_cdac_8bit_array_3.drv<63:0>.t47 VSS 0.112f
C4788 hgu_cdac_8bit_array_3.drv<63:0>.t27 VSS 0.112f
C4789 hgu_cdac_8bit_array_3.drv<63:0>.n359 VSS 0.852f
C4790 hgu_cdac_8bit_array_3.drv<63:0>.n360 VSS 0.522f
C4791 hgu_cdac_8bit_array_3.drv<63:0>.t117 VSS 0.0559f
C4792 hgu_cdac_8bit_array_3.drv<63:0>.t11 VSS 0.0559f
C4793 hgu_cdac_8bit_array_3.drv<63:0>.n361 VSS 0.407f
C4794 hgu_cdac_8bit_array_3.drv<63:0>.n362 VSS 0.275f
C4795 hgu_cdac_8bit_array_3.drv<63:0>.t97 VSS 0.0559f
C4796 hgu_cdac_8bit_array_3.drv<63:0>.t92 VSS 0.0559f
C4797 hgu_cdac_8bit_array_3.drv<63:0>.n363 VSS 0.413f
C4798 hgu_cdac_8bit_array_3.drv<63:0>.t64 VSS 0.112f
C4799 hgu_cdac_8bit_array_3.drv<63:0>.t89 VSS 0.112f
C4800 hgu_cdac_8bit_array_3.drv<63:0>.n364 VSS 0.76f
C4801 hgu_cdac_8bit_array_3.drv<63:0>.n365 VSS 0.431f
C4802 hgu_cdac_8bit_array_3.drv<63:0>.n366 VSS 0.0832f
C4803 hgu_cdac_8bit_array_3.drv<63:0>.t52 VSS 0.112f
C4804 hgu_cdac_8bit_array_3.drv<63:0>.t58 VSS 0.112f
C4805 hgu_cdac_8bit_array_3.drv<63:0>.n367 VSS 0.825f
C4806 hgu_cdac_8bit_array_3.drv<63:0>.n368 VSS 3.8f
C4807 hgu_cdac_8bit_array_3.drv<63:0>.n369 VSS 1.53f
C4808 hgu_cdac_8bit_array_3.drv<63:0>.n370 VSS -1.85f
C4809 hgu_cdac_8bit_array_3.drv<63:0>.n371 VSS 4.23f
C4810 hgu_cdac_8bit_array_3.drv<63:0>.n372 VSS 8.79f
C4811 hgu_cdac_8bit_array_3.drv<63:0>.n373 VSS 9.84f
C4812 hgu_cdac_8bit_array_3.drv<63:0>.n374 VSS 0.834f
C4813 hgu_cdac_8bit_array_3.drv<63:0>.n375 VSS -0.492f
C4814 hgu_cdac_8bit_array_3.drv<63:0>.n376 VSS -1.85f
C4815 hgu_cdac_8bit_array_3.drv<63:0>.n377 VSS 4.67f
C4816 hgu_cdac_8bit_array_3.drv<63:0>.n378 VSS -1.85f
C4817 hgu_cdac_8bit_array_3.drv<63:0>.n379 VSS -0.492f
C4818 hgu_cdac_8bit_array_3.drv<63:0>.n380 VSS 0.646f
C4819 hgu_cdac_8bit_array_3.drv<63:0>.n381 VSS 0.156f
C4820 hgu_cdac_8bit_array_3.drv<63:0>.n382 VSS 0.156f
C4821 hgu_cdac_8bit_array_3.drv<63:0>.n383 VSS 0.69f
C4822 hgu_cdac_8bit_array_3.drv<63:0>.n384 VSS -0.492f
C4823 hgu_cdac_8bit_array_3.drv<63:0>.n385 VSS -1.85f
C4824 hgu_cdac_8bit_array_3.drv<63:0>.n386 VSS 4.67f
C4825 hgu_cdac_8bit_array_3.drv<63:0>.n387 VSS -1.85f
C4826 hgu_cdac_8bit_array_3.drv<63:0>.n388 VSS -0.492f
C4827 hgu_cdac_8bit_array_3.drv<63:0>.n389 VSS 0.646f
C4828 hgu_cdac_8bit_array_3.drv<63:0>.n390 VSS 0.156f
C4829 hgu_cdac_8bit_array_3.drv<63:0>.n391 VSS 0.156f
C4830 hgu_cdac_8bit_array_3.drv<63:0>.n392 VSS 0.69f
C4831 hgu_cdac_8bit_array_3.drv<63:0>.n393 VSS -0.492f
C4832 hgu_cdac_8bit_array_3.drv<63:0>.n394 VSS -1.85f
C4833 hgu_cdac_8bit_array_3.drv<63:0>.n395 VSS 4.67f
C4834 hgu_cdac_8bit_array_3.drv<63:0>.n396 VSS -1.85f
C4835 hgu_cdac_8bit_array_3.drv<63:0>.n397 VSS -0.492f
C4836 hgu_cdac_8bit_array_3.drv<63:0>.n398 VSS 0.646f
C4837 hgu_cdac_8bit_array_3.drv<63:0>.n399 VSS 0.156f
C4838 hgu_cdac_8bit_array_3.drv<63:0>.n400 VSS 0.156f
C4839 hgu_cdac_8bit_array_3.drv<63:0>.n401 VSS 0.69f
C4840 hgu_cdac_8bit_array_3.drv<63:0>.n402 VSS -0.492f
C4841 hgu_cdac_8bit_array_3.drv<63:0>.n403 VSS -1.85f
C4842 hgu_cdac_8bit_array_3.drv<63:0>.n404 VSS 4.67f
C4843 hgu_cdac_8bit_array_3.drv<63:0>.n405 VSS -1.85f
C4844 hgu_cdac_8bit_array_3.drv<63:0>.n406 VSS -0.492f
C4845 hgu_cdac_8bit_array_3.drv<63:0>.n407 VSS 0.646f
C4846 hgu_cdac_8bit_array_3.drv<63:0>.n408 VSS 0.156f
C4847 hgu_cdac_8bit_array_3.drv<63:0>.n409 VSS 0.156f
C4848 hgu_cdac_8bit_array_3.drv<63:0>.n410 VSS 0.69f
C4849 hgu_cdac_8bit_array_3.drv<63:0>.n411 VSS -0.492f
C4850 hgu_cdac_8bit_array_3.drv<63:0>.n412 VSS -1.85f
C4851 hgu_cdac_8bit_array_3.drv<63:0>.n413 VSS 4.67f
C4852 hgu_cdac_8bit_array_3.drv<63:0>.n414 VSS -1.85f
C4853 hgu_cdac_8bit_array_3.drv<63:0>.n415 VSS -0.492f
C4854 hgu_cdac_8bit_array_3.drv<63:0>.n416 VSS 0.646f
C4855 hgu_cdac_8bit_array_3.drv<63:0>.n417 VSS 0.156f
C4856 hgu_cdac_8bit_array_3.drv<63:0>.n418 VSS 0.156f
C4857 hgu_cdac_8bit_array_3.drv<63:0>.n419 VSS 0.69f
C4858 hgu_cdac_8bit_array_3.drv<63:0>.n420 VSS -0.492f
C4859 hgu_cdac_8bit_array_3.drv<63:0>.n421 VSS -1.85f
C4860 hgu_cdac_8bit_array_3.drv<63:0>.n422 VSS 4.67f
C4861 hgu_cdac_8bit_array_3.drv<63:0>.n423 VSS -1.85f
C4862 hgu_cdac_8bit_array_3.drv<63:0>.n424 VSS -0.492f
C4863 hgu_cdac_8bit_array_3.drv<63:0>.n425 VSS 0.646f
C4864 hgu_cdac_8bit_array_3.drv<63:0>.n426 VSS 0.156f
C4865 hgu_cdac_8bit_array_3.drv<63:0>.n427 VSS 0.156f
C4866 hgu_cdac_8bit_array_3.drv<63:0>.n428 VSS 0.69f
C4867 hgu_cdac_8bit_array_3.drv<63:0>.n429 VSS -0.492f
C4868 hgu_cdac_8bit_array_3.drv<63:0>.n430 VSS -1.85f
C4869 hgu_cdac_8bit_array_3.drv<63:0>.n431 VSS 3.32f
C4870 hgu_cdac_8bit_array_3.drv<63:0>.n432 VSS -1.85f
C4871 hgu_cdac_8bit_array_3.drv<63:0>.n433 VSS -0.492f
C4872 hgu_cdac_8bit_array_3.drv<63:0>.n434 VSS 0.646f
C4873 hgu_cdac_8bit_array_3.drv<63:0>.n435 VSS 0.156f
C4874 hgu_cdac_8bit_array_3.drv<63:0>.n436 VSS 0.156f
C4875 hgu_cdac_8bit_array_3.drv<63:0>.n437 VSS 0.69f
C4876 hgu_cdac_8bit_array_3.drv<63:0>.n438 VSS -0.492f
C4877 hgu_cdac_8bit_array_3.drv<63:0>.n439 VSS -1.85f
C4878 hgu_cdac_8bit_array_3.drv<63:0>.n440 VSS 4.67f
C4879 hgu_cdac_8bit_array_3.drv<63:0>.n441 VSS -1.85f
C4880 hgu_cdac_8bit_array_3.drv<63:0>.n442 VSS -0.492f
C4881 hgu_cdac_8bit_array_3.drv<63:0>.n443 VSS 0.646f
C4882 hgu_cdac_8bit_array_3.drv<63:0>.n444 VSS 0.156f
C4883 hgu_cdac_8bit_array_3.drv<63:0>.n445 VSS 0.156f
C4884 hgu_cdac_8bit_array_3.drv<63:0>.n446 VSS 0.69f
C4885 hgu_cdac_8bit_array_3.drv<63:0>.n447 VSS -0.492f
C4886 hgu_cdac_8bit_array_3.drv<63:0>.n448 VSS -1.85f
C4887 hgu_cdac_8bit_array_3.drv<63:0>.n449 VSS 4.67f
C4888 hgu_cdac_8bit_array_3.drv<63:0>.n450 VSS -1.85f
C4889 hgu_cdac_8bit_array_3.drv<63:0>.n451 VSS -0.492f
C4890 hgu_cdac_8bit_array_3.drv<63:0>.n452 VSS 0.646f
C4891 hgu_cdac_8bit_array_3.drv<63:0>.n453 VSS 0.156f
C4892 hgu_cdac_8bit_array_3.drv<63:0>.n454 VSS 0.156f
C4893 hgu_cdac_8bit_array_3.drv<63:0>.n455 VSS 0.69f
C4894 hgu_cdac_8bit_array_3.drv<63:0>.n456 VSS -0.492f
C4895 hgu_cdac_8bit_array_3.drv<63:0>.n457 VSS -1.85f
C4896 hgu_cdac_8bit_array_3.drv<63:0>.n458 VSS 4.67f
C4897 hgu_cdac_8bit_array_3.drv<63:0>.n459 VSS -1.85f
C4898 hgu_cdac_8bit_array_3.drv<63:0>.n460 VSS -0.492f
C4899 hgu_cdac_8bit_array_3.drv<63:0>.n461 VSS 0.646f
C4900 hgu_cdac_8bit_array_3.drv<63:0>.n462 VSS 0.156f
C4901 hgu_cdac_8bit_array_3.drv<63:0>.n463 VSS 0.156f
C4902 hgu_cdac_8bit_array_3.drv<63:0>.n464 VSS 0.69f
C4903 hgu_cdac_8bit_array_3.drv<63:0>.n465 VSS -0.492f
C4904 hgu_cdac_8bit_array_3.drv<63:0>.n466 VSS -1.85f
C4905 hgu_cdac_8bit_array_3.drv<63:0>.n467 VSS 4.67f
C4906 hgu_cdac_8bit_array_3.drv<63:0>.n468 VSS -1.85f
C4907 hgu_cdac_8bit_array_3.drv<63:0>.n469 VSS -0.492f
C4908 hgu_cdac_8bit_array_3.drv<63:0>.n470 VSS 0.646f
C4909 hgu_cdac_8bit_array_3.drv<63:0>.n471 VSS 0.156f
C4910 hgu_cdac_8bit_array_3.drv<63:0>.n472 VSS 0.156f
C4911 hgu_cdac_8bit_array_3.drv<63:0>.n473 VSS 0.69f
C4912 hgu_cdac_8bit_array_3.drv<63:0>.n474 VSS -0.492f
C4913 hgu_cdac_8bit_array_3.drv<63:0>.n475 VSS -1.85f
C4914 hgu_cdac_8bit_array_3.drv<63:0>.n476 VSS 4.67f
C4915 hgu_cdac_8bit_array_3.drv<63:0>.n477 VSS -1.85f
C4916 hgu_cdac_8bit_array_3.drv<63:0>.n478 VSS -0.492f
C4917 hgu_cdac_8bit_array_3.drv<63:0>.n479 VSS 0.646f
C4918 hgu_cdac_8bit_array_3.drv<63:0>.n480 VSS 0.156f
C4919 hgu_cdac_8bit_array_3.drv<63:0>.n481 VSS 0.156f
C4920 hgu_cdac_8bit_array_3.drv<63:0>.n482 VSS 0.69f
C4921 hgu_cdac_8bit_array_3.drv<63:0>.n483 VSS -0.492f
C4922 hgu_cdac_8bit_array_3.drv<63:0>.n484 VSS -1.85f
C4923 hgu_cdac_8bit_array_3.drv<63:0>.n485 VSS 4.67f
C4924 hgu_cdac_8bit_array_3.drv<63:0>.n486 VSS -1.85f
C4925 hgu_cdac_8bit_array_3.drv<63:0>.n487 VSS -0.492f
C4926 hgu_cdac_8bit_array_3.drv<63:0>.n488 VSS 0.646f
C4927 hgu_cdac_8bit_array_3.drv<63:0>.n489 VSS 0.156f
C4928 hgu_cdac_8bit_array_3.drv<63:0>.n490 VSS 0.156f
C4929 hgu_cdac_8bit_array_3.drv<63:0>.n491 VSS 0.69f
C4930 hgu_cdac_8bit_array_3.drv<63:0>.n492 VSS -0.492f
C4931 hgu_cdac_8bit_array_3.drv<63:0>.n493 VSS -1.85f
C4932 hgu_cdac_8bit_array_3.drv<63:0>.n494 VSS 4.67f
C4933 hgu_cdac_8bit_array_3.drv<63:0>.n495 VSS -1.85f
C4934 hgu_cdac_8bit_array_3.drv<63:0>.n496 VSS -0.492f
C4935 hgu_cdac_8bit_array_3.drv<63:0>.n497 VSS 0.646f
C4936 hgu_cdac_8bit_array_3.drv<63:0>.n498 VSS 0.156f
C4937 hgu_cdac_8bit_array_3.drv<63:0>.n499 VSS 0.156f
C4938 hgu_cdac_8bit_array_3.drv<63:0>.n500 VSS 0.69f
C4939 hgu_cdac_8bit_array_3.drv<63:0>.n501 VSS 0.187f
C4940 hgu_cdac_8bit_array_3.drv<63:0>.n502 VSS 0.246f
C4941 hgu_cdac_8bit_array_3.drv<63:0>.n503 VSS 0.192f
C4942 hgu_cdac_8bit_array_3.drv<63:0>.n504 VSS 6.56f
C4943 hgu_cdac_8bit_array_3.drv<63:0>.n505 VSS -1.85f
C4944 hgu_cdac_8bit_array_3.drv<63:0>.n506 VSS -0.492f
C4945 hgu_cdac_8bit_array_3.drv<63:0>.n507 VSS 0.646f
C4946 hgu_cdac_8bit_array_3.drv<63:0>.n508 VSS 0.156f
C4947 hgu_cdac_8bit_array_3.drv<63:0>.n509 VSS 0.156f
C4948 hgu_cdac_8bit_array_3.drv<63:0>.n510 VSS 0.69f
C4949 hgu_cdac_8bit_array_3.drv<63:0>.n511 VSS -0.492f
C4950 hgu_cdac_8bit_array_3.drv<63:0>.n512 VSS -1.85f
C4951 hgu_cdac_8bit_array_3.drv<63:0>.n513 VSS 6.56f
C4952 hgu_cdac_8bit_array_3.drv<63:0>.n514 VSS -1.85f
C4953 hgu_cdac_8bit_array_3.drv<63:0>.n515 VSS -0.492f
C4954 hgu_cdac_8bit_array_3.drv<63:0>.n516 VSS 0.646f
C4955 hgu_cdac_8bit_array_3.drv<63:0>.n517 VSS 0.156f
C4956 hgu_cdac_8bit_array_3.drv<63:0>.n518 VSS 0.156f
C4957 hgu_cdac_8bit_array_3.drv<63:0>.n519 VSS 0.69f
C4958 hgu_cdac_8bit_array_3.drv<63:0>.n520 VSS -0.492f
C4959 hgu_cdac_8bit_array_3.drv<63:0>.n521 VSS -1.85f
C4960 hgu_cdac_8bit_array_3.drv<63:0>.n522 VSS 6.56f
C4961 hgu_cdac_8bit_array_3.drv<63:0>.n523 VSS -1.85f
C4962 hgu_cdac_8bit_array_3.drv<63:0>.n524 VSS -0.492f
C4963 hgu_cdac_8bit_array_3.drv<63:0>.n525 VSS 0.646f
C4964 hgu_cdac_8bit_array_3.drv<63:0>.n526 VSS 0.156f
C4965 hgu_cdac_8bit_array_3.drv<63:0>.n527 VSS 0.156f
C4966 hgu_cdac_8bit_array_3.drv<63:0>.n528 VSS 0.69f
C4967 hgu_cdac_8bit_array_3.drv<63:0>.n529 VSS -0.492f
C4968 hgu_cdac_8bit_array_3.drv<63:0>.n530 VSS -1.85f
C4969 hgu_cdac_8bit_array_3.drv<63:0>.n531 VSS 6.56f
C4970 hgu_cdac_8bit_array_3.drv<63:0>.n532 VSS -1.85f
C4971 hgu_cdac_8bit_array_3.drv<63:0>.n533 VSS -0.492f
C4972 hgu_cdac_8bit_array_3.drv<63:0>.n534 VSS 0.646f
C4973 hgu_cdac_8bit_array_3.drv<63:0>.n535 VSS 0.156f
C4974 hgu_cdac_8bit_array_3.drv<63:0>.n536 VSS 0.156f
C4975 hgu_cdac_8bit_array_3.drv<63:0>.n537 VSS 0.69f
C4976 hgu_cdac_8bit_array_3.drv<63:0>.n538 VSS -0.492f
C4977 hgu_cdac_8bit_array_3.drv<63:0>.n539 VSS -1.85f
C4978 hgu_cdac_8bit_array_3.drv<63:0>.n540 VSS 6.56f
C4979 hgu_cdac_8bit_array_3.drv<63:0>.n541 VSS -1.85f
C4980 hgu_cdac_8bit_array_3.drv<63:0>.n542 VSS -0.492f
C4981 hgu_cdac_8bit_array_3.drv<63:0>.n543 VSS 0.646f
C4982 hgu_cdac_8bit_array_3.drv<63:0>.n544 VSS 0.156f
C4983 hgu_cdac_8bit_array_3.drv<63:0>.n545 VSS 0.156f
C4984 hgu_cdac_8bit_array_3.drv<63:0>.n546 VSS 0.69f
C4985 hgu_cdac_8bit_array_3.drv<63:0>.n547 VSS -0.492f
C4986 hgu_cdac_8bit_array_3.drv<63:0>.n548 VSS -1.85f
C4987 hgu_cdac_8bit_array_3.drv<63:0>.n549 VSS 6.56f
C4988 hgu_cdac_8bit_array_3.drv<63:0>.n550 VSS -1.85f
C4989 hgu_cdac_8bit_array_3.drv<63:0>.n551 VSS -0.492f
C4990 hgu_cdac_8bit_array_3.drv<63:0>.n552 VSS 0.646f
C4991 hgu_cdac_8bit_array_3.drv<63:0>.n553 VSS 0.156f
C4992 hgu_cdac_8bit_array_3.drv<63:0>.n554 VSS 0.156f
C4993 hgu_cdac_8bit_array_3.drv<63:0>.n555 VSS 0.69f
C4994 hgu_cdac_8bit_array_3.drv<63:0>.n556 VSS -0.492f
C4995 hgu_cdac_8bit_array_3.drv<63:0>.n557 VSS -1.85f
C4996 hgu_cdac_8bit_array_3.drv<63:0>.n558 VSS 6.56f
C4997 hgu_cdac_8bit_array_3.drv<63:0>.n559 VSS -1.85f
C4998 hgu_cdac_8bit_array_3.drv<63:0>.n560 VSS -0.492f
C4999 hgu_cdac_8bit_array_3.drv<63:0>.n561 VSS 0.646f
C5000 hgu_cdac_8bit_array_3.drv<63:0>.n562 VSS 0.156f
C5001 hgu_cdac_8bit_array_3.drv<63:0>.n563 VSS 0.156f
C5002 hgu_cdac_8bit_array_3.drv<63:0>.n564 VSS 0.69f
C5003 hgu_cdac_8bit_array_3.drv<63:0>.n565 VSS -0.492f
C5004 hgu_cdac_8bit_array_3.drv<63:0>.n566 VSS -1.85f
C5005 hgu_cdac_8bit_array_3.drv<63:0>.n567 VSS 6.56f
C5006 hgu_cdac_8bit_array_3.drv<63:0>.n568 VSS -1.85f
C5007 hgu_cdac_8bit_array_3.drv<63:0>.n569 VSS -0.492f
C5008 hgu_cdac_8bit_array_3.drv<63:0>.n570 VSS 0.646f
C5009 hgu_cdac_8bit_array_3.drv<63:0>.n571 VSS 0.156f
C5010 hgu_cdac_8bit_array_3.drv<63:0>.n572 VSS 0.156f
C5011 hgu_cdac_8bit_array_3.drv<63:0>.n573 VSS 0.69f
C5012 hgu_cdac_8bit_array_3.drv<63:0>.n574 VSS -0.492f
C5013 hgu_cdac_8bit_array_3.drv<63:0>.n575 VSS -1.85f
C5014 hgu_cdac_8bit_array_3.drv<63:0>.n576 VSS 6.56f
C5015 hgu_cdac_8bit_array_3.drv<63:0>.n577 VSS -1.85f
C5016 hgu_cdac_8bit_array_3.drv<63:0>.n578 VSS -0.492f
C5017 hgu_cdac_8bit_array_3.drv<63:0>.n579 VSS 0.646f
C5018 hgu_cdac_8bit_array_3.drv<63:0>.n580 VSS 0.156f
C5019 hgu_cdac_8bit_array_3.drv<63:0>.n581 VSS 0.156f
C5020 hgu_cdac_8bit_array_3.drv<63:0>.n582 VSS 0.69f
C5021 hgu_cdac_8bit_array_3.drv<63:0>.n583 VSS -0.492f
C5022 hgu_cdac_8bit_array_3.drv<63:0>.n584 VSS -1.85f
C5023 hgu_cdac_8bit_array_3.drv<63:0>.n585 VSS 6.56f
C5024 hgu_cdac_8bit_array_3.drv<63:0>.n586 VSS -1.85f
C5025 hgu_cdac_8bit_array_3.drv<63:0>.n587 VSS -0.492f
C5026 hgu_cdac_8bit_array_3.drv<63:0>.n588 VSS 0.646f
C5027 hgu_cdac_8bit_array_3.drv<63:0>.n589 VSS 0.156f
C5028 hgu_cdac_8bit_array_3.drv<63:0>.n590 VSS 0.156f
C5029 hgu_cdac_8bit_array_3.drv<63:0>.n591 VSS 0.69f
C5030 hgu_cdac_8bit_array_3.drv<63:0>.n592 VSS -0.492f
C5031 hgu_cdac_8bit_array_3.drv<63:0>.n593 VSS -1.85f
C5032 hgu_cdac_8bit_array_3.drv<63:0>.n594 VSS 6.56f
C5033 hgu_cdac_8bit_array_3.drv<63:0>.n595 VSS -1.85f
C5034 hgu_cdac_8bit_array_3.drv<63:0>.n596 VSS -0.492f
C5035 hgu_cdac_8bit_array_3.drv<63:0>.n597 VSS 0.646f
C5036 hgu_cdac_8bit_array_3.drv<63:0>.n598 VSS 0.156f
C5037 hgu_cdac_8bit_array_3.drv<63:0>.n599 VSS 0.156f
C5038 hgu_cdac_8bit_array_3.drv<63:0>.n600 VSS 0.69f
C5039 hgu_cdac_8bit_array_3.drv<63:0>.n601 VSS -0.492f
C5040 hgu_cdac_8bit_array_3.drv<63:0>.n602 VSS -1.88f
C5041 d<6>.t31 VSS 0.0196f
C5042 d<6>.t0 VSS 0.0341f
C5043 d<6>.t75 VSS 0.0196f
C5044 d<6>.t51 VSS 0.0341f
C5045 d<6>.t88 VSS 0.0196f
C5046 d<6>.t64 VSS 0.0341f
C5047 d<6>.t103 VSS 0.0196f
C5048 d<6>.t77 VSS 0.0341f
C5049 d<6>.t26 VSS 0.0196f
C5050 d<6>.t124 VSS 0.0341f
C5051 d<6>.t112 VSS 0.0196f
C5052 d<6>.t86 VSS 0.0341f
C5053 d<6>.t2 VSS 0.0196f
C5054 d<6>.t101 VSS 0.0341f
C5055 d<6>.t53 VSS 0.0196f
C5056 d<6>.t24 VSS 0.0341f
C5057 d<6>.t65 VSS 0.0196f
C5058 d<6>.t40 VSS 0.0341f
C5059 d<6>.t108 VSS 0.0196f
C5060 d<6>.t84 VSS 0.0341f
C5061 d<6>.t126 VSS 0.0196f
C5062 d<6>.t99 VSS 0.0341f
C5063 d<6>.t50 VSS 0.0196f
C5064 d<6>.t20 VSS 0.0341f
C5065 d<6>.t92 VSS 0.0196f
C5066 d<6>.t70 VSS 0.0341f
C5067 d<6>.t117 VSS 0.0196f
C5068 d<6>.t91 VSS 0.0341f
C5069 d<6>.t41 VSS 0.0196f
C5070 d<6>.t12 VSS 0.0341f
C5071 d<6>.t85 VSS 0.0196f
C5072 d<6>.t61 VSS 0.0341f
C5073 d<6>.t5 VSS 0.0196f
C5074 d<6>.t105 VSS 0.0341f
C5075 d<6>.t21 VSS 0.0196f
C5076 d<6>.t120 VSS 0.0341f
C5077 d<6>.t37 VSS 0.0196f
C5078 d<6>.t8 VSS 0.0341f
C5079 d<6>.t82 VSS 0.0196f
C5080 d<6>.t59 VSS 0.0341f
C5081 d<6>.t14 VSS 0.0196f
C5082 d<6>.t113 VSS 0.0341f
C5083 d<6>.t62 VSS 0.0196f
C5084 d<6>.t36 VSS 0.0341f
C5085 d<6>.t106 VSS 0.0196f
C5086 d<6>.t81 VSS 0.0341f
C5087 d<6>.t121 VSS 0.0196f
C5088 d<6>.t96 VSS 0.0341f
C5089 d<6>.t10 VSS 0.0196f
C5090 d<6>.t110 VSS 0.0341f
C5091 d<6>.t60 VSS 0.0196f
C5092 d<6>.t34 VSS 0.0341f
C5093 d<6>.t104 VSS 0.0196f
C5094 d<6>.t78 VSS 0.0341f
C5095 d<6>.t119 VSS 0.0196f
C5096 d<6>.t94 VSS 0.0341f
C5097 d<6>.t54 VSS 0.0196f
C5098 d<6>.t27 VSS 0.0341f
C5099 d<6>.t97 VSS 0.0196f
C5100 d<6>.t74 VSS 0.0341f
C5101 d<6>.t17 VSS 0.0196f
C5102 d<6>.t116 VSS 0.0341f
C5103 d<6>.t35 VSS 0.0196f
C5104 d<6>.t6 VSS 0.0341f
C5105 d<6>.t79 VSS 0.0196f
C5106 d<6>.t57 VSS 0.0341f
C5107 d<6>.t95 VSS 0.0196f
C5108 d<6>.t71 VSS 0.0341f
C5109 d<6>.t15 VSS 0.0196f
C5110 d<6>.t114 VSS 0.0341f
C5111 d<6>.t33 VSS 0.0196f
C5112 d<6>.t4 VSS 0.0341f
C5113 d<6>.t118 VSS 0.0196f
C5114 d<6>.t93 VSS 0.0341f
C5115 d<6>.t43 VSS 0.0196f
C5116 d<6>.t13 VSS 0.0341f
C5117 d<6>.t23 VSS 0.0196f
C5118 d<6>.t122 VSS 0.0341f
C5119 d<6>.t72 VSS 0.0196f
C5120 d<6>.t46 VSS 0.0341f
C5121 d<6>.t115 VSS 0.0196f
C5122 d<6>.t89 VSS 0.0341f
C5123 d<6>.t38 VSS 0.0196f
C5124 d<6>.t9 VSS 0.0341f
C5125 d<6>.t55 VSS 0.0196f
C5126 d<6>.t28 VSS 0.0341f
C5127 d<6>.t68 VSS 0.0196f
C5128 d<6>.t42 VSS 0.0341f
C5129 d<6>.t32 VSS 0.0196f
C5130 d<6>.t3 VSS 0.0341f
C5131 d<6>.t48 VSS 0.0196f
C5132 d<6>.t18 VSS 0.0341f
C5133 d<6>.t90 VSS 0.0196f
C5134 d<6>.t67 VSS 0.0341f
C5135 d<6>.t11 VSS 0.0196f
C5136 d<6>.t111 VSS 0.0341f
C5137 d<6>.t29 VSS 0.0196f
C5138 d<6>.t127 VSS 0.0341f
C5139 d<6>.t45 VSS 0.0196f
C5140 d<6>.t16 VSS 0.0341f
C5141 d<6>.t87 VSS 0.0196f
C5142 d<6>.t63 VSS 0.0341f
C5143 d<6>.t7 VSS 0.0196f
C5144 d<6>.t107 VSS 0.0341f
C5145 d<6>.t69 VSS 0.0196f
C5146 d<6>.t44 VSS 0.0341f
C5147 d<6>.t80 VSS 0.0196f
C5148 d<6>.t58 VSS 0.0341f
C5149 d<6>.t1 VSS 0.0196f
C5150 d<6>.t100 VSS 0.0341f
C5151 d<6>.t52 VSS 0.0196f
C5152 d<6>.t22 VSS 0.0341f
C5153 d<6>.t66 VSS 0.0196f
C5154 d<6>.t39 VSS 0.0341f
C5155 d<6>.t109 VSS 0.0196f
C5156 d<6>.t83 VSS 0.0341f
C5157 d<6>.t125 VSS 0.0196f
C5158 d<6>.t98 VSS 0.0341f
C5159 d<6>.t49 VSS 0.0196f
C5160 d<6>.t19 VSS 0.0341f
C5161 d<6>.t102 VSS 0.0196f
C5162 d<6>.t76 VSS 0.0341f
C5163 d<6>.t25 VSS 0.0196f
C5164 d<6>.t123 VSS 0.0341f
C5165 d<6>.t73 VSS 0.0196f
C5166 d<6>.t47 VSS 0.0341f
C5167 d<6>.t56 VSS 0.0196f
C5168 d<6>.t30 VSS 0.0341f
C5169 d<6>.n0 VSS 0.0636f
C5170 d<6>.n1 VSS 0.0732f
C5171 d<6>.n2 VSS 0.0732f
C5172 d<6>.n3 VSS 0.0732f
C5173 d<6>.n4 VSS 0.0732f
C5174 d<6>.n5 VSS 0.0732f
C5175 d<6>.n6 VSS 0.0732f
C5176 d<6>.n7 VSS 0.0732f
C5177 d<6>.n8 VSS 0.0732f
C5178 d<6>.n9 VSS 0.0732f
C5179 d<6>.n10 VSS 0.0732f
C5180 d<6>.n11 VSS 0.0732f
C5181 d<6>.n12 VSS 0.0732f
C5182 d<6>.n13 VSS 0.0732f
C5183 d<6>.n14 VSS 0.0732f
C5184 d<6>.n15 VSS 0.0732f
C5185 d<6>.n16 VSS 0.0732f
C5186 d<6>.n17 VSS 0.0732f
C5187 d<6>.n18 VSS 0.0732f
C5188 d<6>.n19 VSS 0.0732f
C5189 d<6>.n20 VSS 0.0732f
C5190 d<6>.n21 VSS 0.0732f
C5191 d<6>.n22 VSS 0.0732f
C5192 d<6>.n23 VSS 0.0732f
C5193 d<6>.n24 VSS 0.0732f
C5194 d<6>.n25 VSS 0.0732f
C5195 d<6>.n26 VSS 0.0732f
C5196 d<6>.n27 VSS 0.0732f
C5197 d<6>.n28 VSS 0.0732f
C5198 d<6>.n29 VSS 0.0732f
C5199 d<6>.n30 VSS 0.0732f
C5200 d<6>.n31 VSS 0.0732f
C5201 d<6>.n32 VSS 0.0732f
C5202 d<6>.n33 VSS 0.0732f
C5203 d<6>.n34 VSS 0.0732f
C5204 d<6>.n35 VSS 0.0732f
C5205 d<6>.n36 VSS 0.0732f
C5206 d<6>.n37 VSS 0.0732f
C5207 d<6>.n38 VSS 0.0732f
C5208 d<6>.n39 VSS 0.0732f
C5209 d<6>.n40 VSS 0.0732f
C5210 d<6>.n41 VSS 0.0732f
C5211 d<6>.n42 VSS 0.0732f
C5212 d<6>.n43 VSS 0.0732f
C5213 d<6>.n44 VSS 0.0732f
C5214 d<6>.n45 VSS 0.0732f
C5215 d<6>.n46 VSS 0.0732f
C5216 d<6>.n47 VSS 0.0732f
C5217 d<6>.n48 VSS 0.0732f
C5218 d<6>.n49 VSS 0.0732f
C5219 d<6>.n50 VSS 0.0732f
C5220 d<6>.n51 VSS 0.0732f
C5221 d<6>.n52 VSS 0.0732f
C5222 d<6>.n53 VSS 0.0732f
C5223 d<6>.n54 VSS 0.0732f
C5224 d<6>.n55 VSS 0.0732f
C5225 d<6>.n56 VSS 0.0732f
C5226 d<6>.n57 VSS 0.0732f
C5227 d<6>.n58 VSS 0.0732f
C5228 d<6>.n59 VSS 0.0732f
C5229 d<6>.n60 VSS 0.0732f
C5230 d<6>.n61 VSS 0.0732f
C5231 d<6>.n62 VSS 0.0732f
C5232 d<6>.n63 VSS 0.0578f
C5233 hgu_cdac_8bit_array_2.drv<31:0>.n0 VSS 10.2f
C5234 hgu_cdac_8bit_array_2.drv<31:0>.n1 VSS -4.18f
C5235 hgu_cdac_8bit_array_2.drv<31:0>.n2 VSS -2.65f
C5236 hgu_cdac_8bit_array_2.drv<31:0>.n3 VSS -4.26f
C5237 hgu_cdac_8bit_array_2.drv<31:0>.n4 VSS -4.26f
C5238 hgu_cdac_8bit_array_2.drv<31:0>.n5 VSS -2.65f
C5239 hgu_cdac_8bit_array_2.drv<31:0>.n6 VSS -4.18f
C5240 hgu_cdac_8bit_array_2.drv<31:0>.n7 VSS 14.8f
C5241 hgu_cdac_8bit_array_2.drv<31:0>.n8 VSS -4.18f
C5242 hgu_cdac_8bit_array_2.drv<31:0>.n9 VSS -2.65f
C5243 hgu_cdac_8bit_array_2.drv<31:0>.n10 VSS -4.26f
C5244 hgu_cdac_8bit_array_2.drv<31:0>.n11 VSS -4.26f
C5245 hgu_cdac_8bit_array_2.drv<31:0>.n12 VSS -2.65f
C5246 hgu_cdac_8bit_array_2.drv<31:0>.n13 VSS -4.18f
C5247 hgu_cdac_8bit_array_2.drv<31:0>.n14 VSS 14.8f
C5248 hgu_cdac_8bit_array_2.drv<31:0>.n15 VSS -4.18f
C5249 hgu_cdac_8bit_array_2.drv<31:0>.n16 VSS -2.65f
C5250 hgu_cdac_8bit_array_2.drv<31:0>.n17 VSS -4.26f
C5251 hgu_cdac_8bit_array_2.drv<31:0>.n18 VSS -4.26f
C5252 hgu_cdac_8bit_array_2.drv<31:0>.n19 VSS -2.65f
C5253 hgu_cdac_8bit_array_2.drv<31:0>.n20 VSS -4.18f
C5254 hgu_cdac_8bit_array_2.drv<31:0>.n21 VSS 14.8f
C5255 hgu_cdac_8bit_array_2.drv<31:0>.n22 VSS -4.18f
C5256 hgu_cdac_8bit_array_2.drv<31:0>.n23 VSS -2.65f
C5257 hgu_cdac_8bit_array_2.drv<31:0>.n24 VSS -4.26f
C5258 hgu_cdac_8bit_array_2.drv<31:0>.n25 VSS -4.26f
C5259 hgu_cdac_8bit_array_2.drv<31:0>.n26 VSS -2.65f
C5260 hgu_cdac_8bit_array_2.drv<31:0>.n27 VSS -4.18f
C5261 hgu_cdac_8bit_array_2.drv<31:0>.n28 VSS 14.8f
C5262 hgu_cdac_8bit_array_2.drv<31:0>.n29 VSS -4.18f
C5263 hgu_cdac_8bit_array_2.drv<31:0>.n30 VSS -2.65f
C5264 hgu_cdac_8bit_array_2.drv<31:0>.n31 VSS -4.26f
C5265 hgu_cdac_8bit_array_2.drv<31:0>.n32 VSS -4.26f
C5266 hgu_cdac_8bit_array_2.drv<31:0>.n33 VSS -2.65f
C5267 hgu_cdac_8bit_array_2.drv<31:0>.n34 VSS -4.18f
C5268 hgu_cdac_8bit_array_2.drv<31:0>.n35 VSS 14.8f
C5269 hgu_cdac_8bit_array_2.drv<31:0>.n36 VSS -4.18f
C5270 hgu_cdac_8bit_array_2.drv<31:0>.n37 VSS -2.65f
C5271 hgu_cdac_8bit_array_2.drv<31:0>.n38 VSS -4.26f
C5272 hgu_cdac_8bit_array_2.drv<31:0>.n39 VSS -4.26f
C5273 hgu_cdac_8bit_array_2.drv<31:0>.n40 VSS -2.65f
C5274 hgu_cdac_8bit_array_2.drv<31:0>.n41 VSS -4.18f
C5275 hgu_cdac_8bit_array_2.drv<31:0>.n42 VSS 5.02f
C5276 hgu_cdac_8bit_array_2.drv<31:0>.n43 VSS -4.18f
C5277 hgu_cdac_8bit_array_2.drv<31:0>.n44 VSS -2.65f
C5278 hgu_cdac_8bit_array_2.drv<31:0>.n45 VSS -4.26f
C5279 hgu_cdac_8bit_array_2.drv<31:0>.n46 VSS -4.26f
C5280 hgu_cdac_8bit_array_2.drv<31:0>.n47 VSS -2.65f
C5281 hgu_cdac_8bit_array_2.drv<31:0>.n48 VSS -4.18f
C5282 hgu_cdac_8bit_array_2.drv<31:0>.n49 VSS 5.02f
C5283 hgu_cdac_8bit_array_2.drv<31:0>.n50 VSS -4.18f
C5284 hgu_cdac_8bit_array_2.drv<31:0>.n51 VSS -2.65f
C5285 hgu_cdac_8bit_array_2.drv<31:0>.n52 VSS -4.26f
C5286 hgu_cdac_8bit_array_2.drv<31:0>.n53 VSS -4.26f
C5287 hgu_cdac_8bit_array_2.drv<31:0>.n54 VSS -2.65f
C5288 hgu_cdac_8bit_array_2.drv<31:0>.n55 VSS -4.18f
C5289 hgu_cdac_8bit_array_2.drv<31:0>.n56 VSS 5.02f
C5290 hgu_cdac_8bit_array_2.drv<31:0>.n57 VSS -4.18f
C5291 hgu_cdac_8bit_array_2.drv<31:0>.n58 VSS -2.65f
C5292 hgu_cdac_8bit_array_2.drv<31:0>.n59 VSS -4.26f
C5293 hgu_cdac_8bit_array_2.drv<31:0>.n60 VSS -4.26f
C5294 hgu_cdac_8bit_array_2.drv<31:0>.n61 VSS -2.65f
C5295 hgu_cdac_8bit_array_2.drv<31:0>.n62 VSS -4.18f
C5296 hgu_cdac_8bit_array_2.drv<31:0>.n63 VSS 5.02f
C5297 hgu_cdac_8bit_array_2.drv<31:0>.n64 VSS -4.18f
C5298 hgu_cdac_8bit_array_2.drv<31:0>.n65 VSS -2.65f
C5299 hgu_cdac_8bit_array_2.drv<31:0>.n66 VSS -4.26f
C5300 hgu_cdac_8bit_array_2.drv<31:0>.n67 VSS -4.26f
C5301 hgu_cdac_8bit_array_2.drv<31:0>.n68 VSS -2.65f
C5302 hgu_cdac_8bit_array_2.drv<31:0>.n69 VSS -4.18f
C5303 hgu_cdac_8bit_array_2.drv<31:0>.n70 VSS 5.02f
C5304 hgu_cdac_8bit_array_2.drv<31:0>.n71 VSS -4.18f
C5305 hgu_cdac_8bit_array_2.drv<31:0>.n72 VSS -2.65f
C5306 hgu_cdac_8bit_array_2.drv<31:0>.n73 VSS -4.26f
C5307 hgu_cdac_8bit_array_2.drv<31:0>.n74 VSS -4.26f
C5308 hgu_cdac_8bit_array_2.drv<31:0>.n75 VSS -2.65f
C5309 hgu_cdac_8bit_array_2.drv<31:0>.n76 VSS -4.18f
C5310 hgu_cdac_8bit_array_2.drv<31:0>.n77 VSS 5.02f
C5311 hgu_cdac_8bit_array_2.drv<31:0>.n78 VSS -5.01f
C5312 hgu_cdac_8bit_array_2.drv<31:0>.n79 VSS -4.26f
C5313 hgu_cdac_8bit_array_2.drv<31:0>.n80 VSS -2.65f
C5314 hgu_cdac_8bit_array_2.drv<31:0>.n81 VSS -4.18f
C5315 hgu_cdac_8bit_array_2.drv<31:0>.n82 VSS 5.02f
C5316 hgu_cdac_8bit_array_2.drv<31:0>.t37 VSS 0.253f
C5317 hgu_cdac_8bit_array_2.drv<31:0>.t16 VSS 0.253f
C5318 hgu_cdac_8bit_array_2.drv<31:0>.n83 VSS 1.93f
C5319 hgu_cdac_8bit_array_2.drv<31:0>.t12 VSS 0.253f
C5320 hgu_cdac_8bit_array_2.drv<31:0>.t26 VSS 0.253f
C5321 hgu_cdac_8bit_array_2.drv<31:0>.n84 VSS 1.93f
C5322 hgu_cdac_8bit_array_2.drv<31:0>.t63 VSS 0.127f
C5323 hgu_cdac_8bit_array_2.drv<31:0>.t57 VSS 0.127f
C5324 hgu_cdac_8bit_array_2.drv<31:0>.n85 VSS 0.931f
C5325 hgu_cdac_8bit_array_2.drv<31:0>.t36 VSS 0.253f
C5326 hgu_cdac_8bit_array_2.drv<31:0>.t41 VSS 0.253f
C5327 hgu_cdac_8bit_array_2.drv<31:0>.n86 VSS 1.93f
C5328 hgu_cdac_8bit_array_2.drv<31:0>.t50 VSS 0.127f
C5329 hgu_cdac_8bit_array_2.drv<31:0>.t60 VSS 0.127f
C5330 hgu_cdac_8bit_array_2.drv<31:0>.n87 VSS 0.931f
C5331 hgu_cdac_8bit_array_2.drv<31:0>.t21 VSS 0.253f
C5332 hgu_cdac_8bit_array_2.drv<31:0>.t34 VSS 0.253f
C5333 hgu_cdac_8bit_array_2.drv<31:0>.n88 VSS 1.93f
C5334 hgu_cdac_8bit_array_2.drv<31:0>.t4 VSS 0.127f
C5335 hgu_cdac_8bit_array_2.drv<31:0>.t11 VSS 0.127f
C5336 hgu_cdac_8bit_array_2.drv<31:0>.n89 VSS 0.931f
C5337 hgu_cdac_8bit_array_2.drv<31:0>.t15 VSS 0.253f
C5338 hgu_cdac_8bit_array_2.drv<31:0>.t18 VSS 0.253f
C5339 hgu_cdac_8bit_array_2.drv<31:0>.n90 VSS 1.93f
C5340 hgu_cdac_8bit_array_2.drv<31:0>.t46 VSS 0.127f
C5341 hgu_cdac_8bit_array_2.drv<31:0>.t1 VSS 0.127f
C5342 hgu_cdac_8bit_array_2.drv<31:0>.n91 VSS 0.931f
C5343 hgu_cdac_8bit_array_2.drv<31:0>.t31 VSS 0.253f
C5344 hgu_cdac_8bit_array_2.drv<31:0>.t42 VSS 0.253f
C5345 hgu_cdac_8bit_array_2.drv<31:0>.n92 VSS 1.93f
C5346 hgu_cdac_8bit_array_2.drv<31:0>.t9 VSS 0.127f
C5347 hgu_cdac_8bit_array_2.drv<31:0>.t61 VSS 0.127f
C5348 hgu_cdac_8bit_array_2.drv<31:0>.n93 VSS 0.931f
C5349 hgu_cdac_8bit_array_2.drv<31:0>.t14 VSS 0.253f
C5350 hgu_cdac_8bit_array_2.drv<31:0>.t17 VSS 0.253f
C5351 hgu_cdac_8bit_array_2.drv<31:0>.n94 VSS 1.93f
C5352 hgu_cdac_8bit_array_2.drv<31:0>.t45 VSS 0.127f
C5353 hgu_cdac_8bit_array_2.drv<31:0>.t48 VSS 0.127f
C5354 hgu_cdac_8bit_array_2.drv<31:0>.n95 VSS 0.931f
C5355 hgu_cdac_8bit_array_2.drv<31:0>.t30 VSS 0.253f
C5356 hgu_cdac_8bit_array_2.drv<31:0>.t20 VSS 0.253f
C5357 hgu_cdac_8bit_array_2.drv<31:0>.n96 VSS 1.93f
C5358 hgu_cdac_8bit_array_2.drv<31:0>.t8 VSS 0.127f
C5359 hgu_cdac_8bit_array_2.drv<31:0>.t3 VSS 0.127f
C5360 hgu_cdac_8bit_array_2.drv<31:0>.n97 VSS 0.931f
C5361 hgu_cdac_8bit_array_2.drv<31:0>.t25 VSS 0.253f
C5362 hgu_cdac_8bit_array_2.drv<31:0>.t29 VSS 0.253f
C5363 hgu_cdac_8bit_array_2.drv<31:0>.n98 VSS 1.93f
C5364 hgu_cdac_8bit_array_2.drv<31:0>.t56 VSS 0.127f
C5365 hgu_cdac_8bit_array_2.drv<31:0>.t7 VSS 0.127f
C5366 hgu_cdac_8bit_array_2.drv<31:0>.n99 VSS 0.931f
C5367 hgu_cdac_8bit_array_2.drv<31:0>.t40 VSS 0.253f
C5368 hgu_cdac_8bit_array_2.drv<31:0>.t19 VSS 0.253f
C5369 hgu_cdac_8bit_array_2.drv<31:0>.n100 VSS 1.93f
C5370 hgu_cdac_8bit_array_2.drv<31:0>.t59 VSS 0.127f
C5371 hgu_cdac_8bit_array_2.drv<31:0>.t2 VSS 0.127f
C5372 hgu_cdac_8bit_array_2.drv<31:0>.n101 VSS 0.931f
C5373 hgu_cdac_8bit_array_2.drv<31:0>.t24 VSS 0.253f
C5374 hgu_cdac_8bit_array_2.drv<31:0>.t35 VSS 0.253f
C5375 hgu_cdac_8bit_array_2.drv<31:0>.n102 VSS 1.93f
C5376 hgu_cdac_8bit_array_2.drv<31:0>.t55 VSS 0.127f
C5377 hgu_cdac_8bit_array_2.drv<31:0>.t49 VSS 0.127f
C5378 hgu_cdac_8bit_array_2.drv<31:0>.n103 VSS 0.931f
C5379 hgu_cdac_8bit_array_2.drv<31:0>.t38 VSS 0.253f
C5380 hgu_cdac_8bit_array_2.drv<31:0>.t23 VSS 0.253f
C5381 hgu_cdac_8bit_array_2.drv<31:0>.n104 VSS 1.93f
C5382 hgu_cdac_8bit_array_2.drv<31:0>.t52 VSS 0.127f
C5383 hgu_cdac_8bit_array_2.drv<31:0>.t54 VSS 0.127f
C5384 hgu_cdac_8bit_array_2.drv<31:0>.n105 VSS 0.931f
C5385 hgu_cdac_8bit_array_2.drv<31:0>.t33 VSS 0.253f
C5386 hgu_cdac_8bit_array_2.drv<31:0>.t13 VSS 0.253f
C5387 hgu_cdac_8bit_array_2.drv<31:0>.n106 VSS 1.93f
C5388 hgu_cdac_8bit_array_2.drv<31:0>.t0 VSS 0.127f
C5389 hgu_cdac_8bit_array_2.drv<31:0>.t44 VSS 0.127f
C5390 hgu_cdac_8bit_array_2.drv<31:0>.n107 VSS 0.931f
C5391 hgu_cdac_8bit_array_2.drv<31:0>.t27 VSS 0.253f
C5392 hgu_cdac_8bit_array_2.drv<31:0>.t22 VSS 0.253f
C5393 hgu_cdac_8bit_array_2.drv<31:0>.n108 VSS 1.93f
C5394 hgu_cdac_8bit_array_2.drv<31:0>.t58 VSS 0.127f
C5395 hgu_cdac_8bit_array_2.drv<31:0>.t5 VSS 0.127f
C5396 hgu_cdac_8bit_array_2.drv<31:0>.n109 VSS 0.931f
C5397 hgu_cdac_8bit_array_2.drv<31:0>.t28 VSS 0.253f
C5398 hgu_cdac_8bit_array_2.drv<31:0>.t39 VSS 0.253f
C5399 hgu_cdac_8bit_array_2.drv<31:0>.n110 VSS 1.93f
C5400 hgu_cdac_8bit_array_2.drv<31:0>.t6 VSS 0.127f
C5401 hgu_cdac_8bit_array_2.drv<31:0>.t53 VSS 0.127f
C5402 hgu_cdac_8bit_array_2.drv<31:0>.n111 VSS 0.837f
C5403 hgu_cdac_8bit_array_2.drv<31:0>.n112 VSS 0.841f
C5404 hgu_cdac_8bit_array_2.drv<31:0>.t32 VSS 0.253f
C5405 hgu_cdac_8bit_array_2.drv<31:0>.t43 VSS 0.253f
C5406 hgu_cdac_8bit_array_2.drv<31:0>.n113 VSS 1.93f
C5407 hgu_cdac_8bit_array_2.drv<31:0>.t10 VSS 0.127f
C5408 hgu_cdac_8bit_array_2.drv<31:0>.t62 VSS 0.127f
C5409 hgu_cdac_8bit_array_2.drv<31:0>.n114 VSS 0.931f
C5410 hgu_cdac_8bit_array_2.drv<31:0>.n115 VSS 1.19f
C5411 hgu_cdac_8bit_array_2.drv<31:0>.n116 VSS 1.19f
C5412 hgu_cdac_8bit_array_2.drv<31:0>.n117 VSS 1.19f
C5413 hgu_cdac_8bit_array_2.drv<31:0>.n118 VSS 1.19f
C5414 hgu_cdac_8bit_array_2.drv<31:0>.n119 VSS 1.19f
C5415 hgu_cdac_8bit_array_2.drv<31:0>.n120 VSS 1.19f
C5416 hgu_cdac_8bit_array_2.drv<31:0>.n121 VSS 1.19f
C5417 hgu_cdac_8bit_array_2.drv<31:0>.n122 VSS 1.19f
C5418 hgu_cdac_8bit_array_2.drv<31:0>.n123 VSS 1.19f
C5419 hgu_cdac_8bit_array_2.drv<31:0>.n124 VSS 1.19f
C5420 hgu_cdac_8bit_array_2.drv<31:0>.n125 VSS 1.19f
C5421 hgu_cdac_8bit_array_2.drv<31:0>.n126 VSS 1.19f
C5422 hgu_cdac_8bit_array_2.drv<31:0>.n127 VSS 1.19f
C5423 hgu_cdac_8bit_array_2.drv<31:0>.n128 VSS 1.19f
C5424 hgu_cdac_8bit_array_2.drv<31:0>.t51 VSS 0.127f
C5425 hgu_cdac_8bit_array_2.drv<31:0>.t47 VSS 0.127f
C5426 hgu_cdac_8bit_array_2.drv<31:0>.n129 VSS 0.835f
C5427 hgu_cdac_8bit_array_2.drv<31:0>.n130 VSS 28.5f
C5428 hgu_cdac_8bit_array_2.drv<31:0>.n131 VSS 2.79f
C5429 hgu_cdac_8bit_array_2.drv<31:0>.n132 VSS 0.353f
C5430 hgu_cdac_8bit_array_2.drv<31:0>.n133 VSS 0.353f
C5431 hgu_cdac_8bit_array_2.drv<31:0>.n134 VSS 1.46f
C5432 hgu_cdac_8bit_array_2.drv<31:0>.n135 VSS -1.11f
C5433 hgu_cdac_8bit_array_2.drv<31:0>.n136 VSS -4.18f
C5434 hgu_cdac_8bit_array_2.drv<31:0>.n137 VSS 6.86f
C5435 hgu_cdac_8bit_array_2.drv<31:0>.n138 VSS -4.18f
C5436 hgu_cdac_8bit_array_2.drv<31:0>.n139 VSS -1.11f
C5437 hgu_cdac_8bit_array_2.drv<31:0>.n140 VSS 1.56f
C5438 hgu_cdac_8bit_array_2.drv<31:0>.n141 VSS 0.353f
C5439 hgu_cdac_8bit_array_2.drv<31:0>.n142 VSS 0.353f
C5440 hgu_cdac_8bit_array_2.drv<31:0>.n143 VSS 1.46f
C5441 hgu_cdac_8bit_array_2.drv<31:0>.n144 VSS -1.11f
C5442 hgu_cdac_8bit_array_2.drv<31:0>.n145 VSS -4.18f
C5443 hgu_cdac_8bit_array_2.drv<31:0>.n146 VSS 6.86f
C5444 hgu_cdac_8bit_array_2.drv<31:0>.n147 VSS -4.18f
C5445 hgu_cdac_8bit_array_2.drv<31:0>.n148 VSS -1.11f
C5446 hgu_cdac_8bit_array_2.drv<31:0>.n149 VSS 1.56f
C5447 hgu_cdac_8bit_array_2.drv<31:0>.n150 VSS 0.353f
C5448 hgu_cdac_8bit_array_2.drv<31:0>.n151 VSS 0.353f
C5449 hgu_cdac_8bit_array_2.drv<31:0>.n152 VSS 1.46f
C5450 hgu_cdac_8bit_array_2.drv<31:0>.n153 VSS -1.11f
C5451 hgu_cdac_8bit_array_2.drv<31:0>.n154 VSS -4.18f
C5452 hgu_cdac_8bit_array_2.drv<31:0>.n155 VSS 6.86f
C5453 hgu_cdac_8bit_array_2.drv<31:0>.n156 VSS -4.18f
C5454 hgu_cdac_8bit_array_2.drv<31:0>.n157 VSS -1.11f
C5455 hgu_cdac_8bit_array_2.drv<31:0>.n158 VSS 1.56f
C5456 hgu_cdac_8bit_array_2.drv<31:0>.n159 VSS 0.353f
C5457 hgu_cdac_8bit_array_2.drv<31:0>.n160 VSS 0.353f
C5458 hgu_cdac_8bit_array_2.drv<31:0>.n161 VSS 1.46f
C5459 hgu_cdac_8bit_array_2.drv<31:0>.n162 VSS -1.11f
C5460 hgu_cdac_8bit_array_2.drv<31:0>.n163 VSS -4.18f
C5461 hgu_cdac_8bit_array_2.drv<31:0>.n164 VSS 6.86f
C5462 hgu_cdac_8bit_array_2.drv<31:0>.n165 VSS -4.18f
C5463 hgu_cdac_8bit_array_2.drv<31:0>.n166 VSS -1.11f
C5464 hgu_cdac_8bit_array_2.drv<31:0>.n167 VSS 1.56f
C5465 hgu_cdac_8bit_array_2.drv<31:0>.n168 VSS 0.353f
C5466 hgu_cdac_8bit_array_2.drv<31:0>.n169 VSS 0.353f
C5467 hgu_cdac_8bit_array_2.drv<31:0>.n170 VSS 1.46f
C5468 hgu_cdac_8bit_array_2.drv<31:0>.n171 VSS -1.11f
C5469 hgu_cdac_8bit_array_2.drv<31:0>.n172 VSS -4.18f
C5470 hgu_cdac_8bit_array_2.drv<31:0>.n173 VSS 6.86f
C5471 hgu_cdac_8bit_array_2.drv<31:0>.n174 VSS -4.18f
C5472 hgu_cdac_8bit_array_2.drv<31:0>.n175 VSS -1.11f
C5473 hgu_cdac_8bit_array_2.drv<31:0>.n176 VSS 1.56f
C5474 hgu_cdac_8bit_array_2.drv<31:0>.n177 VSS 0.353f
C5475 hgu_cdac_8bit_array_2.drv<31:0>.n178 VSS 0.353f
C5476 hgu_cdac_8bit_array_2.drv<31:0>.n179 VSS 1.46f
C5477 hgu_cdac_8bit_array_2.drv<31:0>.n180 VSS -1.11f
C5478 hgu_cdac_8bit_array_2.drv<31:0>.n181 VSS -4.18f
C5479 hgu_cdac_8bit_array_2.drv<31:0>.n182 VSS 6.86f
C5480 hgu_cdac_8bit_array_2.drv<31:0>.n183 VSS -4.18f
C5481 hgu_cdac_8bit_array_2.drv<31:0>.n184 VSS -1.11f
C5482 hgu_cdac_8bit_array_2.drv<31:0>.n185 VSS 1.56f
C5483 hgu_cdac_8bit_array_2.drv<31:0>.n186 VSS 0.353f
C5484 hgu_cdac_8bit_array_2.drv<31:0>.n187 VSS 0.353f
C5485 hgu_cdac_8bit_array_2.drv<31:0>.n188 VSS 1.46f
C5486 hgu_cdac_8bit_array_2.drv<31:0>.n189 VSS -1.11f
C5487 hgu_cdac_8bit_array_2.drv<31:0>.n190 VSS -4.18f
C5488 hgu_cdac_8bit_array_2.drv<31:0>.n191 VSS 6.86f
C5489 hgu_cdac_8bit_array_2.drv<31:0>.n192 VSS -4.18f
C5490 hgu_cdac_8bit_array_2.drv<31:0>.n193 VSS -1.11f
C5491 hgu_cdac_8bit_array_2.drv<31:0>.n194 VSS 1.56f
C5492 hgu_cdac_8bit_array_2.drv<31:0>.n195 VSS 0.353f
C5493 hgu_cdac_8bit_array_2.drv<31:0>.n196 VSS 0.353f
C5494 hgu_cdac_8bit_array_2.drv<31:0>.n197 VSS 1.46f
C5495 hgu_cdac_8bit_array_2.drv<31:0>.n198 VSS -1.11f
C5496 hgu_cdac_8bit_array_2.drv<31:0>.n199 VSS -4.18f
C5497 hgu_cdac_8bit_array_2.drv<31:0>.n200 VSS 14.8f
C5498 hgu_cdac_8bit_array_2.drv<31:0>.n201 VSS -4.18f
C5499 hgu_cdac_8bit_array_2.drv<31:0>.n202 VSS -1.11f
C5500 hgu_cdac_8bit_array_2.drv<31:0>.n203 VSS 1.56f
C5501 hgu_cdac_8bit_array_2.drv<31:0>.n204 VSS 0.353f
C5502 hgu_cdac_8bit_array_2.drv<31:0>.n205 VSS 0.353f
C5503 hgu_cdac_8bit_array_2.drv<31:0>.n206 VSS 1.46f
C5504 hgu_cdac_8bit_array_2.drv<31:0>.n207 VSS -1.11f
C5505 hgu_cdac_8bit_array_2.drv<31:0>.n208 VSS -4.18f
C5506 hgu_cdac_8bit_array_2.drv<31:0>.n209 VSS 14.8f
C5507 hgu_cdac_8bit_array_2.drv<31:0>.n210 VSS -4.18f
C5508 hgu_cdac_8bit_array_2.drv<31:0>.n211 VSS -1.11f
C5509 hgu_cdac_8bit_array_2.drv<31:0>.n212 VSS 1.27f
C5510 hgu_cdac_8bit_array_2.drv<31:0>.n213 VSS 0.353f
C5511 hgu_cdac_8bit_array_2.drv<31:0>.n214 VSS 0.353f
C5512 hgu_cdac_8bit_array_2.drv<31:0>.n215 VSS 1.46f
C5513 hgu_cdac_8bit_array_2.drv<31:0>.n216 VSS -1.11f
C5514 hgu_cdac_8bit_array_2.drv<31:0>.n217 VSS -4.18f
C5515 hgu_cdac_8bit_array_2.drv<31:0>.n218 VSS 14.8f
C5516 hgu_cdac_8bit_array_2.drv<31:0>.n219 VSS -4.18f
C5517 hgu_cdac_8bit_array_2.drv<31:0>.n220 VSS -1.11f
C5518 hgu_cdac_8bit_array_2.drv<31:0>.n221 VSS 1.56f
C5519 hgu_cdac_8bit_array_2.drv<31:0>.n222 VSS 0.353f
C5520 hgu_cdac_8bit_array_2.drv<31:0>.n223 VSS 0.353f
C5521 hgu_cdac_8bit_array_2.drv<31:0>.n224 VSS 1.46f
C5522 hgu_cdac_8bit_array_2.drv<31:0>.n225 VSS -1.11f
C5523 hgu_cdac_8bit_array_2.drv<31:0>.n226 VSS -4.18f
C5524 hgu_cdac_8bit_array_2.drv<31:0>.n227 VSS 14.8f
C5525 hgu_cdac_8bit_array_2.drv<31:0>.n228 VSS -4.18f
C5526 hgu_cdac_8bit_array_2.drv<31:0>.n229 VSS -1.11f
C5527 hgu_cdac_8bit_array_2.drv<31:0>.n230 VSS 1.56f
C5528 hgu_cdac_8bit_array_2.drv<31:0>.n231 VSS 0.353f
C5529 hgu_cdac_8bit_array_2.drv<31:0>.n232 VSS 0.353f
C5530 hgu_cdac_8bit_array_2.drv<31:0>.n233 VSS 1.46f
C5531 hgu_cdac_8bit_array_2.drv<31:0>.n234 VSS -1.11f
C5532 hgu_cdac_8bit_array_2.drv<31:0>.n235 VSS -4.18f
C5533 hgu_cdac_8bit_array_2.drv<31:0>.n236 VSS 14.8f
C5534 hgu_cdac_8bit_array_2.drv<31:0>.n237 VSS -4.18f
C5535 hgu_cdac_8bit_array_2.drv<31:0>.n238 VSS -1.11f
C5536 hgu_cdac_8bit_array_2.drv<31:0>.n239 VSS 1.56f
C5537 hgu_cdac_8bit_array_2.drv<31:0>.n240 VSS 0.353f
C5538 hgu_cdac_8bit_array_2.drv<31:0>.n241 VSS 0.353f
C5539 hgu_cdac_8bit_array_2.drv<31:0>.n242 VSS 1.46f
C5540 hgu_cdac_8bit_array_2.drv<31:0>.n243 VSS -1.11f
C5541 hgu_cdac_8bit_array_2.drv<31:0>.n244 VSS -4.18f
C5542 hgu_cdac_8bit_array_2.drv<31:0>.n245 VSS -15f
C5543 hgu_cdac_8bit_array_2.drv<31:0>.n246 VSS -4.18f
C5544 hgu_cdac_8bit_array_2.drv<31:0>.n247 VSS -2.65f
C5545 hgu_cdac_8bit_array_2.drv<31:0>.n248 VSS -4.26f
C5546 hgu_cdac_8bit_array_2.drv<31:0>.n249 VSS -4.26f
C5547 hgu_cdac_8bit_array_2.drv<31:0>.n250 VSS -2.65f
C5548 hgu_cdac_8bit_array_2.drv<31:0>.n251 VSS -4.18f
C5549 hgu_cdac_8bit_array_2.drv<31:0>.n252 VSS 14.8f
C5550 hgu_cdac_8bit_array_2.drv<31:0>.n253 VSS -3.7f
C5551 hgu_cdac_8bit_array_2.drv<31:0>.n254 VSS -4.18f
C5552 hgu_cdac_8bit_array_2.drv<31:0>.n255 VSS 14.8f
C5553 hgu_cdac_8bit_array_2.drv<31:0>.n256 VSS 11f
C5554 hgu_cdac_8bit_array_2.drv<31:0>.n257 VSS 1.89f
C5555 hgu_cdac_8bit_array_2.drv<31:0>.n258 VSS -1.11f
C5556 hgu_cdac_8bit_array_2.drv<31:0>.n259 VSS -4.18f
C5557 hgu_cdac_8bit_array_2.drv<31:0>.n260 VSS 14.8f
C5558 hgu_cdac_8bit_array_2.drv<31:0>.n261 VSS -4.18f
C5559 hgu_cdac_8bit_array_2.drv<31:0>.n262 VSS -1.11f
C5560 hgu_cdac_8bit_array_2.drv<31:0>.n263 VSS 1.46f
C5561 hgu_cdac_8bit_array_2.drv<31:0>.n264 VSS 0.353f
C5562 hgu_cdac_8bit_array_2.drv<31:0>.n265 VSS 0.353f
C5563 hgu_cdac_8bit_array_2.drv<31:0>.n266 VSS 1.56f
C5564 hgu_cdac_8bit_array_2.drv<31:0>.n267 VSS -1.11f
C5565 hgu_cdac_8bit_array_2.drv<31:0>.n268 VSS -4.18f
C5566 hgu_cdac_8bit_array_2.drv<31:0>.n269 VSS 14.8f
C5567 hgu_cdac_8bit_array_2.drv<31:0>.n270 VSS -4.18f
C5568 hgu_cdac_8bit_array_2.drv<31:0>.n271 VSS -1.11f
C5569 hgu_cdac_8bit_array_2.drv<31:0>.n272 VSS 1.46f
C5570 hgu_cdac_8bit_array_2.drv<31:0>.n273 VSS 0.353f
C5571 hgu_cdac_8bit_array_2.drv<31:0>.n274 VSS 0.353f
C5572 hgu_cdac_8bit_array_2.drv<31:0>.n275 VSS 1.56f
C5573 hgu_cdac_8bit_array_2.drv<31:0>.n276 VSS -1.11f
C5574 hgu_cdac_8bit_array_2.drv<31:0>.n277 VSS -4.27f
C5575 hgu_cdac_8bit_array_2.drv<7:0>.n0 VSS 0.248f
C5576 hgu_cdac_8bit_array_2.drv<7:0>.n1 VSS 1.01f
C5577 hgu_cdac_8bit_array_2.drv<7:0>.n2 VSS 0.582f
C5578 hgu_cdac_8bit_array_2.drv<7:0>.n3 VSS -0.357f
C5579 hgu_cdac_8bit_array_2.drv<7:0>.n4 VSS 0.484f
C5580 hgu_cdac_8bit_array_2.drv<7:0>.n5 VSS 0.582f
C5581 hgu_cdac_8bit_array_2.drv<7:0>.n6 VSS 0.614f
C5582 hgu_cdac_8bit_array_2.drv<7:0>.n7 VSS -0.357f
C5583 hgu_cdac_8bit_array_2.drv<7:0>.n8 VSS 0.582f
C5584 hgu_cdac_8bit_array_2.drv<7:0>.t8 VSS 0.0812f
C5585 hgu_cdac_8bit_array_2.drv<7:0>.t12 VSS 0.0812f
C5586 hgu_cdac_8bit_array_2.drv<7:0>.n9 VSS 0.619f
C5587 hgu_cdac_8bit_array_2.drv<7:0>.t7 VSS 0.0406f
C5588 hgu_cdac_8bit_array_2.drv<7:0>.t3 VSS 0.0406f
C5589 hgu_cdac_8bit_array_2.drv<7:0>.n10 VSS 0.299f
C5590 hgu_cdac_8bit_array_2.drv<7:0>.n11 VSS 0.381f
C5591 hgu_cdac_8bit_array_2.drv<7:0>.t15 VSS 0.0812f
C5592 hgu_cdac_8bit_array_2.drv<7:0>.t10 VSS 0.0812f
C5593 hgu_cdac_8bit_array_2.drv<7:0>.n12 VSS 0.619f
C5594 hgu_cdac_8bit_array_2.drv<7:0>.t6 VSS 0.0406f
C5595 hgu_cdac_8bit_array_2.drv<7:0>.t1 VSS 0.0406f
C5596 hgu_cdac_8bit_array_2.drv<7:0>.n13 VSS 0.299f
C5597 hgu_cdac_8bit_array_2.drv<7:0>.n14 VSS 2.7f
C5598 hgu_cdac_8bit_array_2.drv<7:0>.n15 VSS 5.94f
C5599 hgu_cdac_8bit_array_2.drv<7:0>.n16 VSS -1.61f
C5600 hgu_cdac_8bit_array_2.drv<7:0>.n17 VSS -1.37f
C5601 hgu_cdac_8bit_array_2.drv<7:0>.n18 VSS -0.851f
C5602 hgu_cdac_8bit_array_2.drv<7:0>.n19 VSS -1.34f
C5603 hgu_cdac_8bit_array_2.drv<7:0>.n20 VSS 3.07f
C5604 hgu_cdac_8bit_array_2.drv<7:0>.n21 VSS 2.74f
C5605 hgu_cdac_8bit_array_2.drv<7:0>.n22 VSS 5.7f
C5606 hgu_cdac_8bit_array_2.drv<7:0>.n23 VSS -0.357f
C5607 hgu_cdac_8bit_array_2.drv<7:0>.n24 VSS -1.34f
C5608 hgu_cdac_8bit_array_2.drv<7:0>.n25 VSS 3.39f
C5609 hgu_cdac_8bit_array_2.drv<7:0>.n26 VSS -1.34f
C5610 hgu_cdac_8bit_array_2.drv<7:0>.n27 VSS -0.357f
C5611 hgu_cdac_8bit_array_2.drv<7:0>.n28 VSS -1.34f
C5612 hgu_cdac_8bit_array_2.drv<7:0>.t9 VSS 0.0812f
C5613 hgu_cdac_8bit_array_2.drv<7:0>.t11 VSS 0.0812f
C5614 hgu_cdac_8bit_array_2.drv<7:0>.n29 VSS 0.619f
C5615 hgu_cdac_8bit_array_2.drv<7:0>.t0 VSS 0.0406f
C5616 hgu_cdac_8bit_array_2.drv<7:0>.t2 VSS 0.0406f
C5617 hgu_cdac_8bit_array_2.drv<7:0>.n30 VSS 0.299f
C5618 hgu_cdac_8bit_array_2.drv<7:0>.n31 VSS 0.381f
C5619 hgu_cdac_8bit_array_2.drv<7:0>.t13 VSS 0.0812f
C5620 hgu_cdac_8bit_array_2.drv<7:0>.t14 VSS 0.0812f
C5621 hgu_cdac_8bit_array_2.drv<7:0>.n32 VSS 0.619f
C5622 hgu_cdac_8bit_array_2.drv<7:0>.t4 VSS 0.0406f
C5623 hgu_cdac_8bit_array_2.drv<7:0>.t5 VSS 0.0406f
C5624 hgu_cdac_8bit_array_2.drv<7:0>.n33 VSS 0.299f
C5625 hgu_cdac_8bit_array_2.drv<7:0>.n34 VSS 3.26f
C5626 hgu_cdac_8bit_array_2.drv<7:0>.n35 VSS -1.19f
C5627 hgu_cdac_8bit_array_2.drv<7:0>.n36 VSS -1.34f
C5628 hgu_cdac_8bit_array_2.drv<7:0>.n37 VSS 3.07f
C5629 hgu_cdac_8bit_array_2.drv<7:0>.n38 VSS 6.83f
C5630 hgu_cdac_8bit_array_2.drv<7:0>.n39 VSS 3.53f
C5631 hgu_cdac_8bit_array_2.drv<7:0>.n40 VSS -1.34f
C5632 hgu_cdac_8bit_array_2.drv<7:0>.n41 VSS 3.39f
C5633 hgu_cdac_8bit_array_2.drv<7:0>.n42 VSS -1.34f
C5634 hgu_cdac_8bit_array_2.drv<7:0>.n43 VSS -0.357f
C5635 hgu_cdac_8bit_array_2.drv<7:0>.n44 VSS -1.37f
C5636 VDD.n0 VSS 0.17f
C5637 VDD.n1 VSS 0.0176f
C5638 VDD.n2 VSS 0.0118f
C5639 VDD.t106 VSS 0.0741f
C5640 VDD.n3 VSS 0.0741f
C5641 VDD.n4 VSS 0.0177f
C5642 VDD.n5 VSS 0.0177f
C5643 VDD.n6 VSS 0.0171f
C5644 VDD.t110 VSS 0.0741f
C5645 VDD.t195 VSS 0.0741f
C5646 VDD.n7 VSS 0.0741f
C5647 VDD.n8 VSS 0.0177f
C5648 VDD.t58 VSS 0.0741f
C5649 VDD.n9 VSS 0.0741f
C5650 VDD.n10 VSS 0.0177f
C5651 VDD.n11 VSS 0.0177f
C5652 VDD.t175 VSS 0.0741f
C5653 VDD.n12 VSS 0.0741f
C5654 VDD.n13 VSS 0.0177f
C5655 VDD.t83 VSS 0.0741f
C5656 VDD.n14 VSS 0.0741f
C5657 VDD.n15 VSS 0.0177f
C5658 VDD.n16 VSS 0.0177f
C5659 VDD.t214 VSS 0.0741f
C5660 VDD.n17 VSS 0.0741f
C5661 VDD.n18 VSS 0.0177f
C5662 VDD.t119 VSS 0.0741f
C5663 VDD.n19 VSS 0.0741f
C5664 VDD.n20 VSS 0.0177f
C5665 VDD.n21 VSS 0.0177f
C5666 VDD.t76 VSS 0.0741f
C5667 VDD.n22 VSS 0.0741f
C5668 VDD.n23 VSS 0.0177f
C5669 VDD.t210 VSS 0.0741f
C5670 VDD.n24 VSS 0.0741f
C5671 VDD.n25 VSS 0.0177f
C5672 VDD.n26 VSS 0.0177f
C5673 VDD.t86 VSS 0.0741f
C5674 VDD.n27 VSS 0.0741f
C5675 VDD.n28 VSS 0.0177f
C5676 VDD.t34 VSS 0.0741f
C5677 VDD.n29 VSS 0.0741f
C5678 VDD.n30 VSS 0.0177f
C5679 VDD.n31 VSS 0.0177f
C5680 VDD.t156 VSS 0.0741f
C5681 VDD.n32 VSS 0.0741f
C5682 VDD.n33 VSS 0.0177f
C5683 VDD.t124 VSS 0.0741f
C5684 VDD.n34 VSS 0.0741f
C5685 VDD.n35 VSS 0.0177f
C5686 VDD.n36 VSS 0.0177f
C5687 VDD.t141 VSS 0.0741f
C5688 VDD.n37 VSS 0.0741f
C5689 VDD.n38 VSS 0.0177f
C5690 VDD.t109 VSS 0.0741f
C5691 VDD.n39 VSS 0.0741f
C5692 VDD.n40 VSS 0.0177f
C5693 VDD.n41 VSS 0.0177f
C5694 VDD.t189 VSS 0.0741f
C5695 VDD.n42 VSS 0.0741f
C5696 VDD.n43 VSS 0.0177f
C5697 VDD.t242 VSS 0.0741f
C5698 VDD.n44 VSS 0.0741f
C5699 VDD.n45 VSS 0.0177f
C5700 VDD.n46 VSS 0.0177f
C5701 VDD.t235 VSS 0.0741f
C5702 VDD.n47 VSS 0.0741f
C5703 VDD.n48 VSS 0.0177f
C5704 VDD.t215 VSS 0.0741f
C5705 VDD.n49 VSS 0.0741f
C5706 VDD.n50 VSS 0.0177f
C5707 VDD.n51 VSS 0.0177f
C5708 VDD.t82 VSS 0.0741f
C5709 VDD.n52 VSS 0.0741f
C5710 VDD.n53 VSS 0.0177f
C5711 VDD.t213 VSS 0.0741f
C5712 VDD.n54 VSS 0.0741f
C5713 VDD.n55 VSS 0.0177f
C5714 VDD.n56 VSS 0.0177f
C5715 VDD.t237 VSS 0.0741f
C5716 VDD.n57 VSS 0.0741f
C5717 VDD.n58 VSS 0.0177f
C5718 VDD.t234 VSS 0.0741f
C5719 VDD.n59 VSS 0.0741f
C5720 VDD.n60 VSS 0.0177f
C5721 VDD.n61 VSS 0.0177f
C5722 VDD.t207 VSS 0.0741f
C5723 VDD.n62 VSS 0.0741f
C5724 VDD.n63 VSS 0.0177f
C5725 VDD.t62 VSS 0.0741f
C5726 VDD.n64 VSS 0.0741f
C5727 VDD.n65 VSS 0.0177f
C5728 VDD.n66 VSS 0.0177f
C5729 VDD.t15 VSS 0.0741f
C5730 VDD.n67 VSS 0.0741f
C5731 VDD.n68 VSS 0.0177f
C5732 VDD.t233 VSS 0.0741f
C5733 VDD.n69 VSS 0.0741f
C5734 VDD.n70 VSS 0.0177f
C5735 VDD.n71 VSS 0.0177f
C5736 VDD.t114 VSS 0.0741f
C5737 VDD.n72 VSS 0.0741f
C5738 VDD.n73 VSS 0.0177f
C5739 VDD.t197 VSS 0.0741f
C5740 VDD.n74 VSS 0.0741f
C5741 VDD.n75 VSS 0.0177f
C5742 VDD.n76 VSS 0.0177f
C5743 VDD.t85 VSS 0.0741f
C5744 VDD.n77 VSS 0.0741f
C5745 VDD.n78 VSS 0.0177f
C5746 VDD.t246 VSS 0.0741f
C5747 VDD.n79 VSS 0.0741f
C5748 VDD.n80 VSS 0.0177f
C5749 VDD.n81 VSS 0.0177f
C5750 VDD.t194 VSS 0.0741f
C5751 VDD.n82 VSS 0.0741f
C5752 VDD.n83 VSS 0.0177f
C5753 VDD.t212 VSS 0.0741f
C5754 VDD.n84 VSS 0.0741f
C5755 VDD.n85 VSS 0.0177f
C5756 VDD.n86 VSS 0.0177f
C5757 VDD.t196 VSS 0.0741f
C5758 VDD.n87 VSS 0.0741f
C5759 VDD.n88 VSS 0.0177f
C5760 VDD.t59 VSS 0.0741f
C5761 VDD.n89 VSS 0.0741f
C5762 VDD.n90 VSS 0.0177f
C5763 VDD.n91 VSS 0.0177f
C5764 VDD.t66 VSS 0.0741f
C5765 VDD.n92 VSS 0.0741f
C5766 VDD.n93 VSS 0.0177f
C5767 VDD.t72 VSS 0.0741f
C5768 VDD.n94 VSS 0.0741f
C5769 VDD.n95 VSS 0.0177f
C5770 VDD.n96 VSS 0.0177f
C5771 VDD.t73 VSS 0.0741f
C5772 VDD.n97 VSS 0.0741f
C5773 VDD.n98 VSS 0.0177f
C5774 VDD.t22 VSS 0.0741f
C5775 VDD.n99 VSS 0.0741f
C5776 VDD.n100 VSS 0.0177f
C5777 VDD.n101 VSS 0.0177f
C5778 VDD.t203 VSS 0.0741f
C5779 VDD.n102 VSS 0.0741f
C5780 VDD.n103 VSS 0.0177f
C5781 VDD.t31 VSS 0.0741f
C5782 VDD.n104 VSS 0.0741f
C5783 VDD.n105 VSS 0.0177f
C5784 VDD.n106 VSS 0.0177f
C5785 VDD.t38 VSS 0.0741f
C5786 VDD.n107 VSS 0.0741f
C5787 VDD.n108 VSS 0.0177f
C5788 VDD.n109 VSS 0.17f
C5789 VDD.t93 VSS 0.0741f
C5790 VDD.n110 VSS 0.0741f
C5791 VDD.n111 VSS 0.0177f
C5792 VDD.t71 VSS 0.0741f
C5793 VDD.n112 VSS 0.0741f
C5794 VDD.n113 VSS 0.0177f
C5795 VDD.n114 VSS 0.0177f
C5796 VDD.t226 VSS 0.0741f
C5797 VDD.n115 VSS 0.0741f
C5798 VDD.n116 VSS 0.0177f
C5799 VDD.t75 VSS 0.0741f
C5800 VDD.n117 VSS 0.0741f
C5801 VDD.n118 VSS 0.0177f
C5802 VDD.n119 VSS 0.0177f
C5803 VDD.t224 VSS 0.0741f
C5804 VDD.n120 VSS 0.0741f
C5805 VDD.n121 VSS 0.0177f
C5806 VDD.t167 VSS 0.0741f
C5807 VDD.n122 VSS 0.0741f
C5808 VDD.n123 VSS 0.0177f
C5809 VDD.n124 VSS 0.0177f
C5810 VDD.t32 VSS 0.0741f
C5811 VDD.n125 VSS 0.0741f
C5812 VDD.n126 VSS 0.0177f
C5813 VDD.t79 VSS 0.0741f
C5814 VDD.n127 VSS 0.0741f
C5815 VDD.n128 VSS 0.0177f
C5816 VDD.n129 VSS 0.0177f
C5817 VDD.t13 VSS 0.0741f
C5818 VDD.n130 VSS 0.0741f
C5819 VDD.n131 VSS 0.0177f
C5820 VDD.t165 VSS 0.0741f
C5821 VDD.n132 VSS 0.0741f
C5822 VDD.n133 VSS 0.0177f
C5823 VDD.n134 VSS 0.0177f
C5824 VDD.t128 VSS 0.0741f
C5825 VDD.n135 VSS 0.0741f
C5826 VDD.n136 VSS 0.0177f
C5827 VDD.t177 VSS 0.0741f
C5828 VDD.n137 VSS 0.0741f
C5829 VDD.n138 VSS 0.0177f
C5830 VDD.n139 VSS 0.0177f
C5831 VDD.t121 VSS 0.0741f
C5832 VDD.n140 VSS 0.0741f
C5833 VDD.n141 VSS 0.0177f
C5834 VDD.t45 VSS 0.0741f
C5835 VDD.n142 VSS 0.0741f
C5836 VDD.n143 VSS 0.0177f
C5837 VDD.n144 VSS 0.0177f
C5838 VDD.t225 VSS 0.0741f
C5839 VDD.n145 VSS 0.0741f
C5840 VDD.n146 VSS 0.0177f
C5841 VDD.t64 VSS 0.0741f
C5842 VDD.n147 VSS 0.0741f
C5843 VDD.n148 VSS 0.0177f
C5844 VDD.n149 VSS 0.0177f
C5845 VDD.t3 VSS 0.0741f
C5846 VDD.n150 VSS 0.0741f
C5847 VDD.n151 VSS 0.0177f
C5848 VDD.t99 VSS 0.0741f
C5849 VDD.n152 VSS 0.0741f
C5850 VDD.n153 VSS 0.0177f
C5851 VDD.n154 VSS 0.0177f
C5852 VDD.t134 VSS 0.0741f
C5853 VDD.n155 VSS 0.0741f
C5854 VDD.n156 VSS 0.0177f
C5855 VDD.t191 VSS 0.0741f
C5856 VDD.n157 VSS 0.0741f
C5857 VDD.n158 VSS 0.0177f
C5858 VDD.n159 VSS 0.0177f
C5859 VDD.t23 VSS 0.0741f
C5860 VDD.n160 VSS 0.0741f
C5861 VDD.n161 VSS 0.0177f
C5862 VDD.t89 VSS 0.0741f
C5863 VDD.n162 VSS 0.0741f
C5864 VDD.n163 VSS 0.0177f
C5865 VDD.n164 VSS 0.0177f
C5866 VDD.t140 VSS 0.0741f
C5867 VDD.n165 VSS 0.0741f
C5868 VDD.n166 VSS 0.0177f
C5869 VDD.t132 VSS 0.0741f
C5870 VDD.n167 VSS 0.0741f
C5871 VDD.n168 VSS 0.0177f
C5872 VDD.n169 VSS 0.0177f
C5873 VDD.t100 VSS 0.0741f
C5874 VDD.n170 VSS 0.0741f
C5875 VDD.n171 VSS 0.0177f
C5876 VDD.t102 VSS 0.0741f
C5877 VDD.n172 VSS 0.0741f
C5878 VDD.n173 VSS 0.0177f
C5879 VDD.n174 VSS 0.0177f
C5880 VDD.t20 VSS 0.0741f
C5881 VDD.n175 VSS 0.0741f
C5882 VDD.n176 VSS 0.0177f
C5883 VDD.t152 VSS 0.0741f
C5884 VDD.n177 VSS 0.0741f
C5885 VDD.n178 VSS 0.0177f
C5886 VDD.n179 VSS 0.0177f
C5887 VDD.t231 VSS 0.0741f
C5888 VDD.n180 VSS 0.0741f
C5889 VDD.n181 VSS 0.0177f
C5890 VDD.t9 VSS 0.0741f
C5891 VDD.n182 VSS 0.0741f
C5892 VDD.n183 VSS 0.0177f
C5893 VDD.n184 VSS 0.0177f
C5894 VDD.t69 VSS 0.0741f
C5895 VDD.n185 VSS 0.0741f
C5896 VDD.n186 VSS 0.0177f
C5897 VDD.t96 VSS 0.0741f
C5898 VDD.n187 VSS 0.0741f
C5899 VDD.n188 VSS 0.0177f
C5900 VDD.n189 VSS 0.0177f
C5901 VDD.t143 VSS 0.0741f
C5902 VDD.n190 VSS 0.0741f
C5903 VDD.n191 VSS 0.0177f
C5904 VDD.t169 VSS 0.0741f
C5905 VDD.n192 VSS 0.0741f
C5906 VDD.n193 VSS 0.0177f
C5907 VDD.n194 VSS 0.0177f
C5908 VDD.t154 VSS 0.0741f
C5909 VDD.n195 VSS 0.0741f
C5910 VDD.n196 VSS 0.0177f
C5911 VDD.t137 VSS 0.0741f
C5912 VDD.n197 VSS 0.0741f
C5913 VDD.n198 VSS 0.0177f
C5914 VDD.n199 VSS 0.0177f
C5915 VDD.t0 VSS 0.0741f
C5916 VDD.n200 VSS 0.0741f
C5917 VDD.n201 VSS 0.0177f
C5918 VDD.t11 VSS 0.0741f
C5919 VDD.n202 VSS 0.0741f
C5920 VDD.n203 VSS 0.0177f
C5921 VDD.n204 VSS 0.0177f
C5922 VDD.t24 VSS 0.0741f
C5923 VDD.n205 VSS 0.0741f
C5924 VDD.n206 VSS 0.0177f
C5925 VDD.t50 VSS 0.0741f
C5926 VDD.n207 VSS 0.0741f
C5927 VDD.n208 VSS 0.0177f
C5928 VDD.n209 VSS 0.0177f
C5929 VDD.t5 VSS 0.0741f
C5930 VDD.n210 VSS 0.0741f
C5931 VDD.n211 VSS 0.0177f
C5932 VDD.t216 VSS 0.0741f
C5933 VDD.n212 VSS 0.0741f
C5934 VDD.n213 VSS 0.0177f
C5935 VDD.n214 VSS 0.0177f
C5936 VDD.t168 VSS 0.0741f
C5937 VDD.n215 VSS 0.17f
C5938 VDD.t118 VSS 0.0741f
C5939 VDD.n216 VSS 0.0741f
C5940 VDD.n217 VSS 0.0177f
C5941 VDD.t95 VSS 0.0741f
C5942 VDD.n218 VSS 0.0741f
C5943 VDD.n219 VSS 0.0177f
C5944 VDD.n220 VSS 0.0177f
C5945 VDD.t98 VSS 0.0741f
C5946 VDD.n221 VSS 0.0741f
C5947 VDD.n222 VSS 0.0177f
C5948 VDD.t4 VSS 0.0741f
C5949 VDD.n223 VSS 0.0741f
C5950 VDD.n224 VSS 0.0177f
C5951 VDD.n225 VSS 0.0177f
C5952 VDD.t200 VSS 0.0741f
C5953 VDD.n226 VSS 0.0741f
C5954 VDD.n227 VSS 0.0177f
C5955 VDD.t223 VSS 0.0741f
C5956 VDD.n228 VSS 0.0741f
C5957 VDD.n229 VSS 0.0177f
C5958 VDD.n230 VSS 0.0177f
C5959 VDD.t92 VSS 0.0741f
C5960 VDD.n231 VSS 0.0741f
C5961 VDD.n232 VSS 0.0177f
C5962 VDD.t151 VSS 0.0741f
C5963 VDD.n233 VSS 0.0741f
C5964 VDD.n234 VSS 0.0177f
C5965 VDD.n235 VSS 0.0177f
C5966 VDD.t14 VSS 0.0741f
C5967 VDD.n236 VSS 0.0741f
C5968 VDD.n237 VSS 0.0177f
C5969 VDD.t133 VSS 0.0741f
C5970 VDD.n238 VSS 0.0741f
C5971 VDD.n239 VSS 0.0177f
C5972 VDD.n240 VSS 0.0177f
C5973 VDD.t198 VSS 0.0741f
C5974 VDD.n241 VSS 0.0741f
C5975 VDD.n242 VSS 0.0177f
C5976 VDD.t161 VSS 0.0741f
C5977 VDD.n243 VSS 0.0741f
C5978 VDD.n244 VSS 0.0177f
C5979 VDD.n245 VSS 0.0177f
C5980 VDD.t171 VSS 0.0741f
C5981 VDD.n246 VSS 0.0741f
C5982 VDD.n247 VSS 0.0177f
C5983 VDD.t142 VSS 0.0741f
C5984 VDD.n248 VSS 0.0741f
C5985 VDD.n249 VSS 0.0177f
C5986 VDD.n250 VSS 0.0177f
C5987 VDD.t91 VSS 0.0741f
C5988 VDD.n251 VSS 0.0741f
C5989 VDD.n252 VSS 0.0177f
C5990 VDD.t97 VSS 0.0741f
C5991 VDD.n253 VSS 0.0741f
C5992 VDD.n254 VSS 0.0177f
C5993 VDD.n255 VSS 0.0177f
C5994 VDD.t94 VSS 0.0741f
C5995 VDD.n256 VSS 0.0741f
C5996 VDD.n257 VSS 0.0177f
C5997 VDD.t173 VSS 0.0741f
C5998 VDD.n258 VSS 0.0741f
C5999 VDD.n259 VSS 0.0177f
C6000 VDD.n260 VSS 0.0177f
C6001 VDD.t138 VSS 0.0741f
C6002 VDD.n261 VSS 0.0741f
C6003 VDD.n262 VSS 0.0177f
C6004 VDD.t46 VSS 0.0741f
C6005 VDD.n263 VSS 0.0741f
C6006 VDD.n264 VSS 0.0177f
C6007 VDD.n265 VSS 0.0177f
C6008 VDD.n266 VSS 0.17f
C6009 VDD.t166 VSS 0.0741f
C6010 VDD.n267 VSS 0.0741f
C6011 VDD.n268 VSS 0.0177f
C6012 VDD.t170 VSS 0.0741f
C6013 VDD.n269 VSS 0.0741f
C6014 VDD.n270 VSS 0.0177f
C6015 VDD.n271 VSS 0.0177f
C6016 VDD.t21 VSS 0.0741f
C6017 VDD.n272 VSS 0.0741f
C6018 VDD.n273 VSS 0.0177f
C6019 VDD.t146 VSS 0.0741f
C6020 VDD.n274 VSS 0.0741f
C6021 VDD.n275 VSS 0.0177f
C6022 VDD.n276 VSS 0.0177f
C6023 VDD.t116 VSS 0.0741f
C6024 VDD.n277 VSS 0.0741f
C6025 VDD.n278 VSS 0.0177f
C6026 VDD.t101 VSS 0.0741f
C6027 VDD.n279 VSS 0.0741f
C6028 VDD.n280 VSS 0.0177f
C6029 VDD.n281 VSS 0.0177f
C6030 VDD.t149 VSS 0.0741f
C6031 VDD.n282 VSS 0.0741f
C6032 VDD.n283 VSS 0.0177f
C6033 VDD.t63 VSS 0.0741f
C6034 VDD.n284 VSS 0.0741f
C6035 VDD.n285 VSS 0.0177f
C6036 VDD.n286 VSS 0.0177f
C6037 VDD.t127 VSS 0.0741f
C6038 VDD.n287 VSS 0.0741f
C6039 VDD.n288 VSS 0.0177f
C6040 VDD.t74 VSS 0.0741f
C6041 VDD.n289 VSS 0.0741f
C6042 VDD.n290 VSS 0.0177f
C6043 VDD.n291 VSS 0.0177f
C6044 VDD.t61 VSS 0.0741f
C6045 VDD.n292 VSS 0.0741f
C6046 VDD.n293 VSS 0.0177f
C6047 VDD.t55 VSS 0.0741f
C6048 VDD.n294 VSS 0.0741f
C6049 VDD.n295 VSS 0.0177f
C6050 VDD.n296 VSS 0.0177f
C6051 VDD.t219 VSS 0.0741f
C6052 VDD.n297 VSS 0.0741f
C6053 VDD.n298 VSS 0.0177f
C6054 VDD.t239 VSS 0.0741f
C6055 VDD.n299 VSS 0.0741f
C6056 VDD.n300 VSS 0.0177f
C6057 VDD.n301 VSS 0.0177f
C6058 VDD.t28 VSS 0.0741f
C6059 VDD.n302 VSS 0.0741f
C6060 VDD.n303 VSS 0.0177f
C6061 VDD.t205 VSS 0.0741f
C6062 VDD.n304 VSS 0.0741f
C6063 VDD.n305 VSS 0.0177f
C6064 VDD.n306 VSS 0.0177f
C6065 VDD.t42 VSS 0.0741f
C6066 VDD.n307 VSS 0.0741f
C6067 VDD.n308 VSS 0.0177f
C6068 VDD.t6 VSS 0.0741f
C6069 VDD.n309 VSS 0.0741f
C6070 VDD.n310 VSS 0.0177f
C6071 VDD.n311 VSS 0.0177f
C6072 VDD.t54 VSS 0.0741f
C6073 VDD.n312 VSS 0.0741f
C6074 VDD.n313 VSS 0.0177f
C6075 VDD.t19 VSS 0.0741f
C6076 VDD.n314 VSS 0.0741f
C6077 VDD.n315 VSS 0.0177f
C6078 VDD.n316 VSS 0.0177f
C6079 VDD.t209 VSS 0.0741f
C6080 VDD.n317 VSS 0.17f
C6081 VDD.t248 VSS 0.0741f
C6082 VDD.n318 VSS 0.0741f
C6083 VDD.n319 VSS 0.0177f
C6084 VDD.t112 VSS 0.0741f
C6085 VDD.n320 VSS 0.0741f
C6086 VDD.n321 VSS 0.0177f
C6087 VDD.n322 VSS 0.0177f
C6088 VDD.t117 VSS 0.0741f
C6089 VDD.n323 VSS 0.0741f
C6090 VDD.n324 VSS 0.0177f
C6091 VDD.t1 VSS 0.0741f
C6092 VDD.n325 VSS 0.0741f
C6093 VDD.n326 VSS 0.0177f
C6094 VDD.n327 VSS 0.0177f
C6095 VDD.t131 VSS 0.0741f
C6096 VDD.n328 VSS 0.0741f
C6097 VDD.n329 VSS 0.0177f
C6098 VDD.t243 VSS 0.0741f
C6099 VDD.n330 VSS 0.0741f
C6100 VDD.n331 VSS 0.0177f
C6101 VDD.n332 VSS 0.0177f
C6102 VDD.t113 VSS 0.0741f
C6103 VDD.n333 VSS 0.0741f
C6104 VDD.n334 VSS 0.0177f
C6105 VDD.t178 VSS 0.0741f
C6106 VDD.n335 VSS 0.0741f
C6107 VDD.n336 VSS 0.0177f
C6108 VDD.n337 VSS 0.0177f
C6109 VDD.t81 VSS 0.0741f
C6110 VDD.n338 VSS 0.0741f
C6111 VDD.n339 VSS 0.0177f
C6112 VDD.t218 VSS 0.0741f
C6113 VDD.n340 VSS 0.0741f
C6114 VDD.n341 VSS 0.0177f
C6115 VDD.n342 VSS 0.0177f
C6116 VDD.n343 VSS 0.17f
C6117 VDD.t2 VSS 0.0741f
C6118 VDD.n344 VSS 0.0741f
C6119 VDD.n345 VSS 0.0177f
C6120 VDD.t29 VSS 0.0741f
C6121 VDD.n346 VSS 0.0741f
C6122 VDD.n347 VSS 0.0177f
C6123 VDD.n348 VSS 0.0177f
C6124 VDD.t105 VSS 0.0741f
C6125 VDD.n349 VSS 0.0741f
C6126 VDD.n350 VSS 0.0177f
C6127 VDD.t115 VSS 0.0741f
C6128 VDD.n351 VSS 0.0741f
C6129 VDD.n352 VSS 0.0177f
C6130 VDD.n353 VSS 0.0177f
C6131 VDD.t57 VSS 0.0741f
C6132 VDD.n354 VSS 0.0741f
C6133 VDD.n355 VSS 0.0177f
C6134 VDD.t49 VSS 0.0741f
C6135 VDD.n356 VSS 0.0741f
C6136 VDD.n357 VSS 0.0177f
C6137 VDD.n358 VSS 0.0177f
C6138 VDD.t180 VSS 0.0741f
C6139 VDD.n359 VSS 0.0741f
C6140 VDD.n360 VSS 0.0177f
C6141 VDD.t120 VSS 0.0741f
C6142 VDD.n361 VSS 0.0741f
C6143 VDD.n362 VSS 0.0177f
C6144 VDD.n363 VSS 0.0177f
C6145 VDD.t183 VSS 0.0741f
C6146 VDD.n364 VSS 0.0741f
C6147 VDD.n365 VSS 0.0177f
C6148 VDD.t217 VSS 0.0741f
C6149 VDD.n366 VSS 0.0741f
C6150 VDD.n367 VSS 0.0177f
C6151 VDD.n368 VSS 0.0177f
C6152 VDD.t35 VSS 0.0741f
C6153 VDD.n369 VSS 0.17f
C6154 VDD.t221 VSS 0.0741f
C6155 VDD.n370 VSS 0.0741f
C6156 VDD.n371 VSS 0.0177f
C6157 VDD.t153 VSS 0.127f
C6158 VDD.n372 VSS 0.0754f
C6159 VDD.n373 VSS 0.0177f
C6160 VDD.n374 VSS 0.0177f
C6161 VDD.t172 VSS 0.125f
C6162 VDD.n375 VSS 0.125f
C6163 VDD.n376 VSS 0.0177f
C6164 VDD.t147 VSS 0.125f
C6165 VDD.n377 VSS 0.125f
C6166 VDD.n378 VSS 0.0177f
C6167 VDD.n379 VSS 0.0177f
C6168 VDD.t228 VSS 0.127f
C6169 VDD.n380 VSS 0.125f
C6170 VDD.n381 VSS 0.0177f
C6171 VDD.t229 VSS 0.0741f
C6172 VDD.n382 VSS 0.0754f
C6173 VDD.n383 VSS 0.0177f
C6174 VDD.n384 VSS 0.0177f
C6175 VDD.t230 VSS 0.0741f
C6176 VDD.n385 VSS 0.0741f
C6177 VDD.n386 VSS 0.0177f
C6178 VDD.n387 VSS 0.17f
C6179 VDD.t181 VSS 0.0741f
C6180 VDD.n388 VSS 0.0741f
C6181 VDD.n389 VSS 0.0177f
C6182 VDD.t87 VSS 0.0946f
C6183 VDD.n390 VSS 0.0774f
C6184 VDD.n391 VSS 0.0532f
C6185 VDD.n392 VSS 0.0177f
C6186 VDD.n393 VSS 0.0177f
C6187 VDD.t222 VSS 0.0946f
C6188 VDD.n394 VSS 0.0774f
C6189 VDD.t185 VSS 0.0741f
C6190 VDD.n395 VSS 0.0532f
C6191 VDD.n396 VSS 0.0177f
C6192 VDD.t145 VSS 0.0741f
C6193 VDD.n397 VSS 0.0741f
C6194 VDD.n398 VSS 0.0177f
C6195 VDD.n399 VSS 0.0177f
C6196 VDD.n400 VSS 0.0728f
C6197 VDD.t240 VSS 0.226f
C6198 VDD.t155 VSS 0.125f
C6199 VDD.n401 VSS 0.125f
C6200 VDD.n402 VSS 0.0177f
C6201 VDD.n403 VSS 0.0177f
C6202 VDD.t184 VSS 0.226f
C6203 VDD.n404 VSS 0.125f
C6204 VDD.n405 VSS 0.0177f
C6205 VDD.n406 VSS 0.037f
C6206 VDD.t244 VSS 0.221f
C6207 VDD.t108 VSS 0.221f
C6208 VDD.n407 VSS 0.208f
C6209 VDD.n408 VSS 0.012f
C6210 VDD.n409 VSS 0.0658f
C6211 VDD.n410 VSS 0.0728f
C6212 VDD.n411 VSS 0.0561f
C6213 VDD.n412 VSS 0.00964f
C6214 VDD.n413 VSS 0.0554f
C6215 VDD.n414 VSS 0.0177f
C6216 VDD.n415 VSS 0.0138f
C6217 VDD.n416 VSS 0.0118f
C6218 VDD.n417 VSS 0.00964f
C6219 VDD.n418 VSS 0.0432f
C6220 VDD.n419 VSS 0.17f
C6221 VDD.n420 VSS 0.0432f
C6222 VDD.n421 VSS 0.0138f
C6223 VDD.t30 VSS 0.0741f
C6224 VDD.n422 VSS 0.0741f
C6225 VDD.n423 VSS 0.0177f
C6226 VDD.n424 VSS 0.0177f
C6227 VDD.n425 VSS 0.0151f
C6228 VDD.n426 VSS 0.00633f
C6229 VDD.n427 VSS 0.013f
C6230 VDD.n428 VSS 0.0177f
C6231 VDD.n429 VSS 0.0802f
C6232 VDD.n430 VSS 0.0177f
C6233 VDD.n431 VSS 0.0177f
C6234 VDD.n432 VSS 0.00633f
C6235 VDD.n433 VSS 0.013f
C6236 VDD.n434 VSS 0.00633f
C6237 VDD.t245 VSS 0.0741f
C6238 VDD.n435 VSS 0.0741f
C6239 VDD.n436 VSS 0.0177f
C6240 VDD.n437 VSS 0.0177f
C6241 VDD.n438 VSS 0.0177f
C6242 VDD.n439 VSS 0.0171f
C6243 VDD.n440 VSS 0.0118f
C6244 VDD.t192 VSS 0.0741f
C6245 VDD.n441 VSS 0.17f
C6246 VDD.n442 VSS 0.0501f
C6247 VDD.n443 VSS 0.0501f
C6248 VDD.n444 VSS 0.0138f
C6249 VDD.n445 VSS 0.0151f
C6250 VDD.t227 VSS 0.0741f
C6251 VDD.n446 VSS 0.0741f
C6252 VDD.n447 VSS 0.0177f
C6253 VDD.n448 VSS 0.0177f
C6254 VDD.n449 VSS 0.0177f
C6255 VDD.n450 VSS 0.00633f
C6256 VDD.n451 VSS 0.013f
C6257 VDD.n452 VSS 0.00633f
C6258 VDD.n453 VSS 0.0177f
C6259 VDD.t88 VSS 0.125f
C6260 VDD.n454 VSS 0.125f
C6261 VDD.n455 VSS 0.0177f
C6262 VDD.n456 VSS 0.0177f
C6263 VDD.n457 VSS 0.013f
C6264 VDD.n458 VSS 0.00633f
C6265 VDD.n459 VSS 0.013f
C6266 VDD.t80 VSS 0.125f
C6267 VDD.n460 VSS 0.125f
C6268 VDD.n461 VSS 0.0177f
C6269 VDD.n462 VSS 0.0177f
C6270 VDD.n463 VSS 0.0177f
C6271 VDD.n464 VSS 0.00633f
C6272 VDD.n465 VSS 0.013f
C6273 VDD.n466 VSS 0.00633f
C6274 VDD.n467 VSS 0.0177f
C6275 VDD.t158 VSS 0.0741f
C6276 VDD.n468 VSS 0.0741f
C6277 VDD.n469 VSS 0.0177f
C6278 VDD.n470 VSS 0.0177f
C6279 VDD.n471 VSS 0.0171f
C6280 VDD.n472 VSS 0.0118f
C6281 VDD.n473 VSS 0.0752f
C6282 VDD.n474 VSS 0.17f
C6283 VDD.n475 VSS 0.0752f
C6284 VDD.n476 VSS 0.0138f
C6285 VDD.n477 VSS 0.0151f
C6286 VDD.n478 VSS 0.00633f
C6287 VDD.t201 VSS 0.0741f
C6288 VDD.n479 VSS 0.0741f
C6289 VDD.n480 VSS 0.0177f
C6290 VDD.n481 VSS 0.0177f
C6291 VDD.n482 VSS 0.0177f
C6292 VDD.n483 VSS 0.013f
C6293 VDD.n484 VSS 0.00633f
C6294 VDD.n485 VSS 0.013f
C6295 VDD.n486 VSS 0.0177f
C6296 VDD.t10 VSS 0.0741f
C6297 VDD.n487 VSS 0.0741f
C6298 VDD.n488 VSS 0.0177f
C6299 VDD.n489 VSS 0.0177f
C6300 VDD.n490 VSS 0.00633f
C6301 VDD.n491 VSS 0.013f
C6302 VDD.n492 VSS 0.00633f
C6303 VDD.t206 VSS 0.0741f
C6304 VDD.n493 VSS 0.0741f
C6305 VDD.n494 VSS 0.0177f
C6306 VDD.n495 VSS 0.0177f
C6307 VDD.n496 VSS 0.0177f
C6308 VDD.n497 VSS 0.013f
C6309 VDD.n498 VSS 0.00633f
C6310 VDD.n499 VSS 0.013f
C6311 VDD.n500 VSS 0.0177f
C6312 VDD.t26 VSS 0.0741f
C6313 VDD.n501 VSS 0.0741f
C6314 VDD.n502 VSS 0.0177f
C6315 VDD.n503 VSS 0.0177f
C6316 VDD.n504 VSS 0.00633f
C6317 VDD.n505 VSS 0.013f
C6318 VDD.n506 VSS 0.00633f
C6319 VDD.t144 VSS 0.0741f
C6320 VDD.n507 VSS 0.0741f
C6321 VDD.n508 VSS 0.0177f
C6322 VDD.n509 VSS 0.0177f
C6323 VDD.n510 VSS 0.0177f
C6324 VDD.n511 VSS 0.0171f
C6325 VDD.n512 VSS 0.0118f
C6326 VDD.t70 VSS 0.0741f
C6327 VDD.n513 VSS 0.17f
C6328 VDD.n514 VSS 0.046f
C6329 VDD.n515 VSS 0.046f
C6330 VDD.n516 VSS 0.0138f
C6331 VDD.n517 VSS 0.0151f
C6332 VDD.n518 VSS 0.00633f
C6333 VDD.n519 VSS 0.0177f
C6334 VDD.t160 VSS 0.0741f
C6335 VDD.n520 VSS 0.0741f
C6336 VDD.n521 VSS 0.0177f
C6337 VDD.n522 VSS 0.0177f
C6338 VDD.n523 VSS 0.013f
C6339 VDD.n524 VSS 0.00633f
C6340 VDD.n525 VSS 0.013f
C6341 VDD.t67 VSS 0.0741f
C6342 VDD.n526 VSS 0.0741f
C6343 VDD.n527 VSS 0.0177f
C6344 VDD.n528 VSS 0.0177f
C6345 VDD.n529 VSS 0.0177f
C6346 VDD.n530 VSS 0.00633f
C6347 VDD.n531 VSS 0.013f
C6348 VDD.n532 VSS 0.00633f
C6349 VDD.n533 VSS 0.0177f
C6350 VDD.t232 VSS 0.0741f
C6351 VDD.n534 VSS 0.0741f
C6352 VDD.n535 VSS 0.0177f
C6353 VDD.n536 VSS 0.0177f
C6354 VDD.n537 VSS 0.013f
C6355 VDD.n538 VSS 0.00633f
C6356 VDD.n539 VSS 0.013f
C6357 VDD.t159 VSS 0.0741f
C6358 VDD.n540 VSS 0.0741f
C6359 VDD.n541 VSS 0.0177f
C6360 VDD.n542 VSS 0.0177f
C6361 VDD.n543 VSS 0.0177f
C6362 VDD.n544 VSS 0.00633f
C6363 VDD.n545 VSS 0.013f
C6364 VDD.n546 VSS 0.00633f
C6365 VDD.n547 VSS 0.0177f
C6366 VDD.t41 VSS 0.0741f
C6367 VDD.n548 VSS 0.0741f
C6368 VDD.n549 VSS 0.0177f
C6369 VDD.n550 VSS 0.0177f
C6370 VDD.n551 VSS 0.0171f
C6371 VDD.n552 VSS 0.0118f
C6372 VDD.n553 VSS 0.0404f
C6373 VDD.n554 VSS 0.17f
C6374 VDD.n555 VSS 0.0404f
C6375 VDD.n556 VSS 0.0138f
C6376 VDD.t36 VSS 0.0741f
C6377 VDD.n557 VSS 0.0741f
C6378 VDD.n558 VSS 0.0177f
C6379 VDD.n559 VSS 0.0177f
C6380 VDD.n560 VSS 0.0151f
C6381 VDD.n561 VSS 0.00633f
C6382 VDD.n562 VSS 0.013f
C6383 VDD.n563 VSS 0.0177f
C6384 VDD.t17 VSS 0.0741f
C6385 VDD.n564 VSS 0.0741f
C6386 VDD.n565 VSS 0.0177f
C6387 VDD.n566 VSS 0.0177f
C6388 VDD.n567 VSS 0.00633f
C6389 VDD.n568 VSS 0.013f
C6390 VDD.n569 VSS 0.00633f
C6391 VDD.t37 VSS 0.0741f
C6392 VDD.n570 VSS 0.0741f
C6393 VDD.n571 VSS 0.0177f
C6394 VDD.n572 VSS 0.0177f
C6395 VDD.n573 VSS 0.0177f
C6396 VDD.n574 VSS 0.013f
C6397 VDD.n575 VSS 0.00633f
C6398 VDD.n576 VSS 0.013f
C6399 VDD.n577 VSS 0.0177f
C6400 VDD.t182 VSS 0.0741f
C6401 VDD.n578 VSS 0.0741f
C6402 VDD.n579 VSS 0.0177f
C6403 VDD.n580 VSS 0.0177f
C6404 VDD.n581 VSS 0.00633f
C6405 VDD.n582 VSS 0.013f
C6406 VDD.n583 VSS 0.00633f
C6407 VDD.t136 VSS 0.0741f
C6408 VDD.n584 VSS 0.0741f
C6409 VDD.n585 VSS 0.0177f
C6410 VDD.n586 VSS 0.0177f
C6411 VDD.n587 VSS 0.0177f
C6412 VDD.n588 VSS 0.013f
C6413 VDD.n589 VSS 0.00633f
C6414 VDD.n590 VSS 0.013f
C6415 VDD.n591 VSS 0.0177f
C6416 VDD.t164 VSS 0.0741f
C6417 VDD.n592 VSS 0.0741f
C6418 VDD.n593 VSS 0.0177f
C6419 VDD.n594 VSS 0.0177f
C6420 VDD.n595 VSS 0.00633f
C6421 VDD.n596 VSS 0.013f
C6422 VDD.n597 VSS 0.00633f
C6423 VDD.t53 VSS 0.0741f
C6424 VDD.n598 VSS 0.0741f
C6425 VDD.n599 VSS 0.0177f
C6426 VDD.n600 VSS 0.0177f
C6427 VDD.n601 VSS 0.0177f
C6428 VDD.n602 VSS 0.013f
C6429 VDD.n603 VSS 0.00633f
C6430 VDD.n604 VSS 0.013f
C6431 VDD.n605 VSS 0.0177f
C6432 VDD.t78 VSS 0.0741f
C6433 VDD.n606 VSS 0.0741f
C6434 VDD.n607 VSS 0.0177f
C6435 VDD.n608 VSS 0.0177f
C6436 VDD.n609 VSS 0.00633f
C6437 VDD.n610 VSS 0.013f
C6438 VDD.n611 VSS 0.00633f
C6439 VDD.t68 VSS 0.0741f
C6440 VDD.n612 VSS 0.0741f
C6441 VDD.n613 VSS 0.0177f
C6442 VDD.n614 VSS 0.0177f
C6443 VDD.n615 VSS 0.0177f
C6444 VDD.n616 VSS 0.013f
C6445 VDD.n617 VSS 0.00633f
C6446 VDD.n618 VSS 0.013f
C6447 VDD.n619 VSS 0.0177f
C6448 VDD.t247 VSS 0.0741f
C6449 VDD.n620 VSS 0.0741f
C6450 VDD.n621 VSS 0.0177f
C6451 VDD.n622 VSS 0.0177f
C6452 VDD.n623 VSS 0.00633f
C6453 VDD.n624 VSS 0.013f
C6454 VDD.n625 VSS 0.00633f
C6455 VDD.t90 VSS 0.0741f
C6456 VDD.n626 VSS 0.0741f
C6457 VDD.n627 VSS 0.0177f
C6458 VDD.n628 VSS 0.0177f
C6459 VDD.n629 VSS 0.0177f
C6460 VDD.n630 VSS 0.0171f
C6461 VDD.n631 VSS 0.0118f
C6462 VDD.t176 VSS 0.0741f
C6463 VDD.n632 VSS 0.17f
C6464 VDD.n633 VSS 0.0896f
C6465 VDD.n634 VSS 0.0896f
C6466 VDD.n635 VSS 0.0138f
C6467 VDD.t162 VSS 0.0741f
C6468 VDD.n636 VSS 0.0741f
C6469 VDD.n637 VSS 0.0177f
C6470 VDD.n638 VSS 0.0177f
C6471 VDD.n639 VSS 0.0151f
C6472 VDD.n640 VSS 0.00633f
C6473 VDD.n641 VSS 0.013f
C6474 VDD.t56 VSS 0.0741f
C6475 VDD.n642 VSS 0.0741f
C6476 VDD.n643 VSS 0.0177f
C6477 VDD.n644 VSS 0.0177f
C6478 VDD.n645 VSS 0.0177f
C6479 VDD.n646 VSS 0.00633f
C6480 VDD.n647 VSS 0.013f
C6481 VDD.n648 VSS 0.00633f
C6482 VDD.n649 VSS 0.0177f
C6483 VDD.t107 VSS 0.0741f
C6484 VDD.n650 VSS 0.0741f
C6485 VDD.n651 VSS 0.0177f
C6486 VDD.n652 VSS 0.0177f
C6487 VDD.n653 VSS 0.013f
C6488 VDD.n654 VSS 0.00633f
C6489 VDD.n655 VSS 0.013f
C6490 VDD.t241 VSS 0.0741f
C6491 VDD.n656 VSS 0.0741f
C6492 VDD.n657 VSS 0.0177f
C6493 VDD.n658 VSS 0.0177f
C6494 VDD.n659 VSS 0.0177f
C6495 VDD.n660 VSS 0.00633f
C6496 VDD.n661 VSS 0.013f
C6497 VDD.n662 VSS 0.00633f
C6498 VDD.n663 VSS 0.0177f
C6499 VDD.t51 VSS 0.0741f
C6500 VDD.n664 VSS 0.0741f
C6501 VDD.n665 VSS 0.0177f
C6502 VDD.n666 VSS 0.0177f
C6503 VDD.n667 VSS 0.013f
C6504 VDD.n668 VSS 0.00633f
C6505 VDD.n669 VSS 0.013f
C6506 VDD.t65 VSS 0.0741f
C6507 VDD.n670 VSS 0.0741f
C6508 VDD.n671 VSS 0.0177f
C6509 VDD.n672 VSS 0.0177f
C6510 VDD.n673 VSS 0.0177f
C6511 VDD.n674 VSS 0.00633f
C6512 VDD.n675 VSS 0.013f
C6513 VDD.n676 VSS 0.00633f
C6514 VDD.n677 VSS 0.0177f
C6515 VDD.t199 VSS 0.0741f
C6516 VDD.n678 VSS 0.0741f
C6517 VDD.n679 VSS 0.0177f
C6518 VDD.n680 VSS 0.0177f
C6519 VDD.n681 VSS 0.013f
C6520 VDD.n682 VSS 0.00633f
C6521 VDD.n683 VSS 0.013f
C6522 VDD.t174 VSS 0.0741f
C6523 VDD.n684 VSS 0.0741f
C6524 VDD.n685 VSS 0.0177f
C6525 VDD.n686 VSS 0.0177f
C6526 VDD.n687 VSS 0.0177f
C6527 VDD.n688 VSS 0.00633f
C6528 VDD.n689 VSS 0.013f
C6529 VDD.n690 VSS 0.00633f
C6530 VDD.n691 VSS 0.0177f
C6531 VDD.t163 VSS 0.0741f
C6532 VDD.n692 VSS 0.0741f
C6533 VDD.n693 VSS 0.0177f
C6534 VDD.n694 VSS 0.0177f
C6535 VDD.n695 VSS 0.013f
C6536 VDD.n696 VSS 0.00633f
C6537 VDD.n697 VSS 0.013f
C6538 VDD.t104 VSS 0.0741f
C6539 VDD.n698 VSS 0.0741f
C6540 VDD.n699 VSS 0.0177f
C6541 VDD.n700 VSS 0.0177f
C6542 VDD.n701 VSS 0.0177f
C6543 VDD.n702 VSS 0.00633f
C6544 VDD.n703 VSS 0.013f
C6545 VDD.n704 VSS 0.00633f
C6546 VDD.n705 VSS 0.0177f
C6547 VDD.t193 VSS 0.0741f
C6548 VDD.n706 VSS 0.0741f
C6549 VDD.n707 VSS 0.0177f
C6550 VDD.n708 VSS 0.0177f
C6551 VDD.n709 VSS 0.0171f
C6552 VDD.n710 VSS 0.0118f
C6553 VDD.n711 VSS 0.0421f
C6554 VDD.n712 VSS 0.17f
C6555 VDD.n713 VSS 0.0421f
C6556 VDD.n714 VSS 0.0138f
C6557 VDD.n715 VSS 0.0151f
C6558 VDD.n716 VSS 0.00633f
C6559 VDD.t52 VSS 0.0741f
C6560 VDD.n717 VSS 0.0741f
C6561 VDD.n718 VSS 0.0177f
C6562 VDD.n719 VSS 0.0177f
C6563 VDD.n720 VSS 0.0177f
C6564 VDD.n721 VSS 0.013f
C6565 VDD.n722 VSS 0.00633f
C6566 VDD.n723 VSS 0.013f
C6567 VDD.n724 VSS 0.0177f
C6568 VDD.t186 VSS 0.0741f
C6569 VDD.n725 VSS 0.0741f
C6570 VDD.n726 VSS 0.0177f
C6571 VDD.n727 VSS 0.0177f
C6572 VDD.n728 VSS 0.00633f
C6573 VDD.n729 VSS 0.013f
C6574 VDD.n730 VSS 0.00633f
C6575 VDD.t43 VSS 0.0741f
C6576 VDD.n731 VSS 0.0741f
C6577 VDD.n732 VSS 0.0177f
C6578 VDD.n733 VSS 0.0177f
C6579 VDD.n734 VSS 0.0177f
C6580 VDD.n735 VSS 0.013f
C6581 VDD.n736 VSS 0.00633f
C6582 VDD.n737 VSS 0.013f
C6583 VDD.n738 VSS 0.0177f
C6584 VDD.t47 VSS 0.0741f
C6585 VDD.n739 VSS 0.0741f
C6586 VDD.n740 VSS 0.0177f
C6587 VDD.n741 VSS 0.0177f
C6588 VDD.n742 VSS 0.00633f
C6589 VDD.n743 VSS 0.013f
C6590 VDD.n744 VSS 0.00633f
C6591 VDD.t12 VSS 0.0741f
C6592 VDD.n745 VSS 0.0741f
C6593 VDD.n746 VSS 0.0177f
C6594 VDD.n747 VSS 0.0177f
C6595 VDD.n748 VSS 0.0177f
C6596 VDD.n749 VSS 0.013f
C6597 VDD.n750 VSS 0.00633f
C6598 VDD.n751 VSS 0.013f
C6599 VDD.n752 VSS 0.0177f
C6600 VDD.t39 VSS 0.0741f
C6601 VDD.n753 VSS 0.0741f
C6602 VDD.n754 VSS 0.0177f
C6603 VDD.n755 VSS 0.0177f
C6604 VDD.n756 VSS 0.00633f
C6605 VDD.n757 VSS 0.013f
C6606 VDD.n758 VSS 0.00633f
C6607 VDD.t129 VSS 0.0741f
C6608 VDD.n759 VSS 0.0741f
C6609 VDD.n760 VSS 0.0177f
C6610 VDD.n761 VSS 0.0177f
C6611 VDD.n762 VSS 0.0177f
C6612 VDD.n763 VSS 0.013f
C6613 VDD.n764 VSS 0.00633f
C6614 VDD.n765 VSS 0.013f
C6615 VDD.n766 VSS 0.0177f
C6616 VDD.t111 VSS 0.0741f
C6617 VDD.n767 VSS 0.0741f
C6618 VDD.n768 VSS 0.0177f
C6619 VDD.n769 VSS 0.0177f
C6620 VDD.n770 VSS 0.00633f
C6621 VDD.n771 VSS 0.013f
C6622 VDD.n772 VSS 0.00633f
C6623 VDD.t187 VSS 0.0741f
C6624 VDD.n773 VSS 0.0741f
C6625 VDD.n774 VSS 0.0177f
C6626 VDD.n775 VSS 0.0177f
C6627 VDD.n776 VSS 0.0177f
C6628 VDD.n777 VSS 0.013f
C6629 VDD.n778 VSS 0.00633f
C6630 VDD.n779 VSS 0.013f
C6631 VDD.n780 VSS 0.0177f
C6632 VDD.t190 VSS 0.0741f
C6633 VDD.n781 VSS 0.0741f
C6634 VDD.n782 VSS 0.0177f
C6635 VDD.n783 VSS 0.0177f
C6636 VDD.n784 VSS 0.00633f
C6637 VDD.n785 VSS 0.013f
C6638 VDD.n786 VSS 0.00633f
C6639 VDD.t44 VSS 0.0741f
C6640 VDD.n787 VSS 0.0741f
C6641 VDD.n788 VSS 0.0177f
C6642 VDD.n789 VSS 0.0177f
C6643 VDD.n790 VSS 0.0177f
C6644 VDD.n791 VSS 0.013f
C6645 VDD.n792 VSS 0.00633f
C6646 VDD.n793 VSS 0.013f
C6647 VDD.n794 VSS 0.0177f
C6648 VDD.t122 VSS 0.0741f
C6649 VDD.n795 VSS 0.0741f
C6650 VDD.n796 VSS 0.0177f
C6651 VDD.n797 VSS 0.0177f
C6652 VDD.n798 VSS 0.00633f
C6653 VDD.n799 VSS 0.013f
C6654 VDD.n800 VSS 0.00633f
C6655 VDD.t220 VSS 0.0741f
C6656 VDD.n801 VSS 0.0741f
C6657 VDD.n802 VSS 0.0177f
C6658 VDD.n803 VSS 0.0177f
C6659 VDD.n804 VSS 0.0177f
C6660 VDD.n805 VSS 0.013f
C6661 VDD.n806 VSS 0.00633f
C6662 VDD.n807 VSS 0.013f
C6663 VDD.n808 VSS 0.0177f
C6664 VDD.t48 VSS 0.0741f
C6665 VDD.n809 VSS 0.0741f
C6666 VDD.n810 VSS 0.0177f
C6667 VDD.n811 VSS 0.0177f
C6668 VDD.n812 VSS 0.00633f
C6669 VDD.n813 VSS 0.013f
C6670 VDD.n814 VSS 0.00633f
C6671 VDD.t33 VSS 0.0741f
C6672 VDD.n815 VSS 0.0741f
C6673 VDD.n816 VSS 0.0177f
C6674 VDD.n817 VSS 0.0177f
C6675 VDD.n818 VSS 0.0177f
C6676 VDD.n819 VSS 0.013f
C6677 VDD.n820 VSS 0.00633f
C6678 VDD.n821 VSS 0.013f
C6679 VDD.n822 VSS 0.0177f
C6680 VDD.t139 VSS 0.0741f
C6681 VDD.n823 VSS 0.0741f
C6682 VDD.n824 VSS 0.0177f
C6683 VDD.n825 VSS 0.0177f
C6684 VDD.n826 VSS 0.00633f
C6685 VDD.n827 VSS 0.013f
C6686 VDD.n828 VSS 0.00633f
C6687 VDD.t188 VSS 0.0741f
C6688 VDD.n829 VSS 0.0741f
C6689 VDD.n830 VSS 0.0177f
C6690 VDD.n831 VSS 0.0177f
C6691 VDD.n832 VSS 0.0177f
C6692 VDD.n833 VSS 0.013f
C6693 VDD.n834 VSS 0.00633f
C6694 VDD.n835 VSS 0.013f
C6695 VDD.n836 VSS 0.0177f
C6696 VDD.t77 VSS 0.0741f
C6697 VDD.n837 VSS 0.0741f
C6698 VDD.n838 VSS 0.0177f
C6699 VDD.n839 VSS 0.0177f
C6700 VDD.n840 VSS 0.00633f
C6701 VDD.n841 VSS 0.013f
C6702 VDD.n842 VSS 0.00633f
C6703 VDD.t135 VSS 0.0741f
C6704 VDD.n843 VSS 0.0741f
C6705 VDD.n844 VSS 0.0177f
C6706 VDD.n845 VSS 0.0177f
C6707 VDD.n846 VSS 0.0177f
C6708 VDD.n847 VSS 0.013f
C6709 VDD.n848 VSS 0.00633f
C6710 VDD.n849 VSS 0.013f
C6711 VDD.n850 VSS 0.0177f
C6712 VDD.t204 VSS 0.0741f
C6713 VDD.n851 VSS 0.0741f
C6714 VDD.n852 VSS 0.0177f
C6715 VDD.n853 VSS 0.0177f
C6716 VDD.n854 VSS 0.00633f
C6717 VDD.n855 VSS 0.013f
C6718 VDD.n856 VSS 0.00633f
C6719 VDD.t150 VSS 0.0741f
C6720 VDD.n857 VSS 0.0741f
C6721 VDD.n858 VSS 0.0177f
C6722 VDD.n859 VSS 0.0177f
C6723 VDD.n860 VSS 0.0177f
C6724 VDD.n861 VSS 0.0171f
C6725 VDD.n862 VSS 0.0118f
C6726 VDD.t103 VSS 0.0741f
C6727 VDD.n863 VSS 0.17f
C6728 VDD.n864 VSS 0.0627f
C6729 VDD.n865 VSS 0.0627f
C6730 VDD.n866 VSS 0.0138f
C6731 VDD.n867 VSS 0.0151f
C6732 VDD.t7 VSS 0.0741f
C6733 VDD.n868 VSS 0.0741f
C6734 VDD.n869 VSS 0.0177f
C6735 VDD.n870 VSS 0.0177f
C6736 VDD.n871 VSS 0.0177f
C6737 VDD.n872 VSS 0.00633f
C6738 VDD.n873 VSS 0.013f
C6739 VDD.n874 VSS 0.00633f
C6740 VDD.n875 VSS 0.0177f
C6741 VDD.t211 VSS 0.0741f
C6742 VDD.n876 VSS 0.0741f
C6743 VDD.n877 VSS 0.0177f
C6744 VDD.n878 VSS 0.0177f
C6745 VDD.n879 VSS 0.013f
C6746 VDD.n880 VSS 0.00633f
C6747 VDD.n881 VSS 0.013f
C6748 VDD.t208 VSS 0.0741f
C6749 VDD.n882 VSS 0.0741f
C6750 VDD.n883 VSS 0.0177f
C6751 VDD.n884 VSS 0.0177f
C6752 VDD.n885 VSS 0.0177f
C6753 VDD.n886 VSS 0.00633f
C6754 VDD.n887 VSS 0.013f
C6755 VDD.n888 VSS 0.00633f
C6756 VDD.n889 VSS 0.0177f
C6757 VDD.t125 VSS 0.0741f
C6758 VDD.n890 VSS 0.0741f
C6759 VDD.n891 VSS 0.0177f
C6760 VDD.n892 VSS 0.0177f
C6761 VDD.n893 VSS 0.013f
C6762 VDD.n894 VSS 0.00633f
C6763 VDD.n895 VSS 0.013f
C6764 VDD.t16 VSS 0.0741f
C6765 VDD.n896 VSS 0.0741f
C6766 VDD.n897 VSS 0.0177f
C6767 VDD.n898 VSS 0.0177f
C6768 VDD.n899 VSS 0.0177f
C6769 VDD.n900 VSS 0.00633f
C6770 VDD.n901 VSS 0.013f
C6771 VDD.n902 VSS 0.00633f
C6772 VDD.n903 VSS 0.0177f
C6773 VDD.t40 VSS 0.0741f
C6774 VDD.n904 VSS 0.0741f
C6775 VDD.n905 VSS 0.0177f
C6776 VDD.n906 VSS 0.0177f
C6777 VDD.n907 VSS 0.013f
C6778 VDD.n908 VSS 0.00633f
C6779 VDD.n909 VSS 0.013f
C6780 VDD.t84 VSS 0.0741f
C6781 VDD.n910 VSS 0.0741f
C6782 VDD.n911 VSS 0.0177f
C6783 VDD.n912 VSS 0.0177f
C6784 VDD.n913 VSS 0.0177f
C6785 VDD.n914 VSS 0.00633f
C6786 VDD.n915 VSS 0.013f
C6787 VDD.n916 VSS 0.00633f
C6788 VDD.n917 VSS 0.0177f
C6789 VDD.t202 VSS 0.0741f
C6790 VDD.n918 VSS 0.0741f
C6791 VDD.n919 VSS 0.0177f
C6792 VDD.n920 VSS 0.0177f
C6793 VDD.n921 VSS 0.013f
C6794 VDD.n922 VSS 0.00633f
C6795 VDD.n923 VSS 0.013f
C6796 VDD.t8 VSS 0.0741f
C6797 VDD.n924 VSS 0.0741f
C6798 VDD.n925 VSS 0.0177f
C6799 VDD.n926 VSS 0.0177f
C6800 VDD.n927 VSS 0.0177f
C6801 VDD.n928 VSS 0.00633f
C6802 VDD.n929 VSS 0.013f
C6803 VDD.n930 VSS 0.00633f
C6804 VDD.n931 VSS 0.0177f
C6805 VDD.t18 VSS 0.0741f
C6806 VDD.n932 VSS 0.0741f
C6807 VDD.n933 VSS 0.0177f
C6808 VDD.n934 VSS 0.0177f
C6809 VDD.n935 VSS 0.013f
C6810 VDD.n936 VSS 0.00633f
C6811 VDD.n937 VSS 0.013f
C6812 VDD.t123 VSS 0.0741f
C6813 VDD.n938 VSS 0.0741f
C6814 VDD.n939 VSS 0.0177f
C6815 VDD.n940 VSS 0.0177f
C6816 VDD.n941 VSS 0.0177f
C6817 VDD.n942 VSS 0.00633f
C6818 VDD.n943 VSS 0.013f
C6819 VDD.n944 VSS 0.00633f
C6820 VDD.n945 VSS 0.0177f
C6821 VDD.t60 VSS 0.0741f
C6822 VDD.n946 VSS 0.0741f
C6823 VDD.n947 VSS 0.0177f
C6824 VDD.n948 VSS 0.0177f
C6825 VDD.n949 VSS 0.013f
C6826 VDD.n950 VSS 0.00633f
C6827 VDD.n951 VSS 0.013f
C6828 VDD.t179 VSS 0.0741f
C6829 VDD.n952 VSS 0.0741f
C6830 VDD.n953 VSS 0.0177f
C6831 VDD.n954 VSS 0.0177f
C6832 VDD.n955 VSS 0.0177f
C6833 VDD.n956 VSS 0.00633f
C6834 VDD.n957 VSS 0.013f
C6835 VDD.n958 VSS 0.00633f
C6836 VDD.n959 VSS 0.0177f
C6837 VDD.t126 VSS 0.0741f
C6838 VDD.n960 VSS 0.0741f
C6839 VDD.n961 VSS 0.0177f
C6840 VDD.n962 VSS 0.0177f
C6841 VDD.n963 VSS 0.013f
C6842 VDD.n964 VSS 0.00633f
C6843 VDD.n965 VSS 0.013f
C6844 VDD.t130 VSS 0.0741f
C6845 VDD.n966 VSS 0.0741f
C6846 VDD.n967 VSS 0.0177f
C6847 VDD.n968 VSS 0.0177f
C6848 VDD.n969 VSS 0.0177f
C6849 VDD.n970 VSS 0.00633f
C6850 VDD.n971 VSS 0.013f
C6851 VDD.n972 VSS 0.00633f
C6852 VDD.n973 VSS 0.0177f
C6853 VDD.t148 VSS 0.0741f
C6854 VDD.n974 VSS 0.0741f
C6855 VDD.n975 VSS 0.0177f
C6856 VDD.n976 VSS 0.0177f
C6857 VDD.n977 VSS 0.013f
C6858 VDD.n978 VSS 0.00633f
C6859 VDD.n979 VSS 0.013f
C6860 VDD.t27 VSS 0.0741f
C6861 VDD.n980 VSS 0.0741f
C6862 VDD.n981 VSS 0.0177f
C6863 VDD.n982 VSS 0.0177f
C6864 VDD.n983 VSS 0.0177f
C6865 VDD.n984 VSS 0.00633f
C6866 VDD.n985 VSS 0.013f
C6867 VDD.n986 VSS 0.00633f
C6868 VDD.n987 VSS 0.0177f
C6869 VDD.t238 VSS 0.0741f
C6870 VDD.n988 VSS 0.0741f
C6871 VDD.n989 VSS 0.0177f
C6872 VDD.n990 VSS 0.0177f
C6873 VDD.n991 VSS 0.013f
C6874 VDD.n992 VSS 0.00633f
C6875 VDD.n993 VSS 0.013f
C6876 VDD.t25 VSS 0.0741f
C6877 VDD.n994 VSS 0.0741f
C6878 VDD.n995 VSS 0.0177f
C6879 VDD.n996 VSS 0.0177f
C6880 VDD.n997 VSS 0.0177f
C6881 VDD.n998 VSS 0.00633f
C6882 VDD.n999 VSS 0.013f
C6883 VDD.n1000 VSS 0.00633f
C6884 VDD.n1001 VSS 0.0177f
C6885 VDD.t157 VSS 0.0741f
C6886 VDD.n1002 VSS 0.0741f
C6887 VDD.n1003 VSS 0.0177f
C6888 VDD.n1004 VSS 0.0177f
C6889 VDD.n1005 VSS 0.013f
C6890 VDD.n1006 VSS 0.00633f
C6891 VDD.n1007 VSS 0.013f
C6892 VDD.t236 VSS 0.0741f
C6893 VDD.n1008 VSS 0.0741f
C6894 VDD.n1009 VSS 0.0177f
C6895 VDD.n1010 VSS 0.0177f
C6896 VDD.n1011 VSS 0.0177f
C6897 VDD.n1012 VSS 0.00633f
C6898 VREF.t249 VSS 0.0352f
C6899 VREF.n0 VSS 0.471f
C6900 VREF.t185 VSS 0.0352f
C6901 VREF.n1 VSS 0.344f
C6902 VREF.t184 VSS 0.0352f
C6903 VREF.n2 VSS 0.474f
C6904 VREF.t30 VSS 0.0352f
C6905 VREF.n3 VSS 0.344f
C6906 VREF.t186 VSS 0.0321f
C6907 VREF.t145 VSS 0.0321f
C6908 VREF.n4 VSS 0.233f
C6909 VREF.n5 VSS 0.0878f
C6910 VREF.t223 VSS 0.0352f
C6911 VREF.n6 VSS 0.575f
C6912 VREF.t229 VSS 0.0352f
C6913 VREF.n7 VSS 0.344f
C6914 VREF.t232 VSS 0.0321f
C6915 VREF.t234 VSS 0.0321f
C6916 VREF.n8 VSS 0.233f
C6917 VREF.n9 VSS 0.0876f
C6918 VREF.t228 VSS 0.0321f
C6919 VREF.t230 VSS 0.0321f
C6920 VREF.n10 VSS 0.233f
C6921 VREF.n11 VSS 0.0876f
C6922 VREF.t233 VSS 0.0321f
C6923 VREF.t235 VSS 0.0321f
C6924 VREF.n12 VSS 0.233f
C6925 VREF.n13 VSS 0.0878f
C6926 VREF.t231 VSS 0.0352f
C6927 VREF.n14 VSS 0.651f
C6928 VREF.t218 VSS 0.0352f
C6929 VREF.n15 VSS 0.344f
C6930 VREF.t183 VSS 0.0321f
C6931 VREF.t202 VSS 0.0321f
C6932 VREF.n16 VSS 0.233f
C6933 VREF.n17 VSS 0.0876f
C6934 VREF.t180 VSS 0.0321f
C6935 VREF.t120 VSS 0.0321f
C6936 VREF.n18 VSS 0.233f
C6937 VREF.n19 VSS 0.0876f
C6938 VREF.t49 VSS 0.0321f
C6939 VREF.t10 VSS 0.0321f
C6940 VREF.n20 VSS 0.233f
C6941 VREF.n21 VSS 0.0876f
C6942 VREF.t57 VSS 0.0321f
C6943 VREF.t207 VSS 0.0321f
C6944 VREF.n22 VSS 0.233f
C6945 VREF.n23 VSS 0.0876f
C6946 VREF.t105 VSS 0.0321f
C6947 VREF.t115 VSS 0.0321f
C6948 VREF.n24 VSS 0.233f
C6949 VREF.n25 VSS 0.0876f
C6950 VREF.t29 VSS 0.0321f
C6951 VREF.t26 VSS 0.0321f
C6952 VREF.n26 VSS 0.233f
C6953 VREF.n27 VSS 0.0876f
C6954 VREF.t2 VSS 0.0321f
C6955 VREF.t144 VSS 0.0321f
C6956 VREF.n28 VSS 0.233f
C6957 VREF.n29 VSS 0.0878f
C6958 VREF.t70 VSS 0.0352f
C6959 VREF.n30 VSS 0.982f
C6960 VREF.t36 VSS 0.0352f
C6961 VREF.n31 VSS 0.344f
C6962 VREF.t54 VSS 0.0321f
C6963 VREF.t19 VSS 0.0321f
C6964 VREF.n32 VSS 0.233f
C6965 VREF.n33 VSS 0.0876f
C6966 VREF.t6 VSS 0.0321f
C6967 VREF.t17 VSS 0.0321f
C6968 VREF.n34 VSS 0.233f
C6969 VREF.n35 VSS 0.0876f
C6970 VREF.t42 VSS 0.0321f
C6971 VREF.t37 VSS 0.0321f
C6972 VREF.n36 VSS 0.233f
C6973 VREF.n37 VSS 0.0876f
C6974 VREF.t28 VSS 0.0321f
C6975 VREF.t206 VSS 0.0321f
C6976 VREF.n38 VSS 0.233f
C6977 VREF.n39 VSS 0.0876f
C6978 VREF.t244 VSS 0.0321f
C6979 VREF.t182 VSS 0.0321f
C6980 VREF.n40 VSS 0.233f
C6981 VREF.n41 VSS 0.0876f
C6982 VREF.t220 VSS 0.0321f
C6983 VREF.t136 VSS 0.0321f
C6984 VREF.n42 VSS 0.233f
C6985 VREF.n43 VSS 0.0876f
C6986 VREF.t61 VSS 0.0321f
C6987 VREF.t55 VSS 0.0321f
C6988 VREF.n44 VSS 0.233f
C6989 VREF.n45 VSS 0.0876f
C6990 VREF.t74 VSS 0.0321f
C6991 VREF.t164 VSS 0.0321f
C6992 VREF.n46 VSS 0.233f
C6993 VREF.n47 VSS 0.0876f
C6994 VREF.t127 VSS 0.0321f
C6995 VREF.t53 VSS 0.0321f
C6996 VREF.n48 VSS 0.233f
C6997 VREF.n49 VSS 0.0876f
C6998 VREF.t149 VSS 0.0321f
C6999 VREF.t63 VSS 0.0321f
C7000 VREF.n50 VSS 0.233f
C7001 VREF.n51 VSS 0.0876f
C7002 VREF.t101 VSS 0.0321f
C7003 VREF.t78 VSS 0.0321f
C7004 VREF.n52 VSS 0.233f
C7005 VREF.n53 VSS 0.0876f
C7006 VREF.t116 VSS 0.0321f
C7007 VREF.t68 VSS 0.0321f
C7008 VREF.n54 VSS 0.233f
C7009 VREF.n55 VSS 0.0876f
C7010 VREF.t21 VSS 0.0321f
C7011 VREF.t146 VSS 0.0321f
C7012 VREF.n56 VSS 0.233f
C7013 VREF.n57 VSS 0.0876f
C7014 VREF.t170 VSS 0.0321f
C7015 VREF.t252 VSS 0.0321f
C7016 VREF.n58 VSS 0.233f
C7017 VREF.n59 VSS 0.0876f
C7018 VREF.t166 VSS 0.0321f
C7019 VREF.t90 VSS 0.0321f
C7020 VREF.n60 VSS 0.233f
C7021 VREF.n61 VSS 0.0878f
C7022 VREF.t176 VSS 0.0352f
C7023 VREF.n62 VSS 1.55f
C7024 VREF.t217 VSS 0.0352f
C7025 VREF.n63 VSS 0.344f
C7026 VREF.t5 VSS 0.0321f
C7027 VREF.t52 VSS 0.0321f
C7028 VREF.n64 VSS 0.233f
C7029 VREF.n65 VSS 0.0876f
C7030 VREF.t24 VSS 0.0321f
C7031 VREF.t50 VSS 0.0321f
C7032 VREF.n66 VSS 0.233f
C7033 VREF.n67 VSS 0.0876f
C7034 VREF.t11 VSS 0.0321f
C7035 VREF.t187 VSS 0.0321f
C7036 VREF.n68 VSS 0.233f
C7037 VREF.n69 VSS 0.0876f
C7038 VREF.t0 VSS 0.0321f
C7039 VREF.t43 VSS 0.0321f
C7040 VREF.n70 VSS 0.233f
C7041 VREF.n71 VSS 0.0876f
C7042 VREF.t154 VSS 0.0321f
C7043 VREF.t137 VSS 0.0321f
C7044 VREF.n72 VSS 0.233f
C7045 VREF.n73 VSS 0.0876f
C7046 VREF.t169 VSS 0.0321f
C7047 VREF.t47 VSS 0.0321f
C7048 VREF.n74 VSS 0.233f
C7049 VREF.n75 VSS 0.0876f
C7050 VREF.t143 VSS 0.0321f
C7051 VREF.t12 VSS 0.0321f
C7052 VREF.n76 VSS 0.233f
C7053 VREF.n77 VSS 0.0876f
C7054 VREF.t69 VSS 0.0321f
C7055 VREF.t96 VSS 0.0321f
C7056 VREF.n78 VSS 0.233f
C7057 VREF.n79 VSS 0.0876f
C7058 VREF.t9 VSS 0.0321f
C7059 VREF.t39 VSS 0.0321f
C7060 VREF.n80 VSS 0.233f
C7061 VREF.n81 VSS 0.0876f
C7062 VREF.t236 VSS 0.0321f
C7063 VREF.t129 VSS 0.0321f
C7064 VREF.n82 VSS 0.233f
C7065 VREF.n83 VSS 0.0876f
C7066 VREF.t20 VSS 0.0321f
C7067 VREF.t152 VSS 0.0321f
C7068 VREF.n84 VSS 0.233f
C7069 VREF.n85 VSS 0.0876f
C7070 VREF.t102 VSS 0.0321f
C7071 VREF.t111 VSS 0.0321f
C7072 VREF.n86 VSS 0.233f
C7073 VREF.n87 VSS 0.0876f
C7074 VREF.t100 VSS 0.0321f
C7075 VREF.t188 VSS 0.0321f
C7076 VREF.n88 VSS 0.233f
C7077 VREF.n89 VSS 0.0876f
C7078 VREF.t140 VSS 0.0321f
C7079 VREF.t132 VSS 0.0321f
C7080 VREF.n90 VSS 0.233f
C7081 VREF.n91 VSS 0.0876f
C7082 VREF.t89 VSS 0.0321f
C7083 VREF.t191 VSS 0.0321f
C7084 VREF.n92 VSS 0.233f
C7085 VREF.n93 VSS 0.0876f
C7086 VREF.t23 VSS 0.0321f
C7087 VREF.t44 VSS 0.0321f
C7088 VREF.n94 VSS 0.233f
C7089 VREF.n95 VSS 0.0876f
C7090 VREF.t134 VSS 0.0321f
C7091 VREF.t192 VSS 0.0321f
C7092 VREF.n96 VSS 0.233f
C7093 VREF.n97 VSS 0.0876f
C7094 VREF.t99 VSS 0.0321f
C7095 VREF.t122 VSS 0.0321f
C7096 VREF.n98 VSS 0.233f
C7097 VREF.n99 VSS 0.0876f
C7098 VREF.t3 VSS 0.0321f
C7099 VREF.t221 VSS 0.0321f
C7100 VREF.n100 VSS 0.233f
C7101 VREF.n101 VSS 0.0876f
C7102 VREF.t226 VSS 0.0321f
C7103 VREF.t64 VSS 0.0321f
C7104 VREF.n102 VSS 0.233f
C7105 VREF.n103 VSS 0.0876f
C7106 VREF.t45 VSS 0.0321f
C7107 VREF.t48 VSS 0.0321f
C7108 VREF.n104 VSS 0.233f
C7109 VREF.n105 VSS 0.0876f
C7110 VREF.t121 VSS 0.0321f
C7111 VREF.t33 VSS 0.0321f
C7112 VREF.n106 VSS 0.233f
C7113 VREF.n107 VSS 0.0876f
C7114 VREF.t128 VSS 0.0321f
C7115 VREF.t177 VSS 0.0321f
C7116 VREF.n108 VSS 0.233f
C7117 VREF.n109 VSS 0.0876f
C7118 VREF.t165 VSS 0.0321f
C7119 VREF.t139 VSS 0.0321f
C7120 VREF.n110 VSS 0.233f
C7121 VREF.n111 VSS 0.0876f
C7122 VREF.t13 VSS 0.0321f
C7123 VREF.t189 VSS 0.0321f
C7124 VREF.n112 VSS 0.233f
C7125 VREF.n113 VSS 0.0876f
C7126 VREF.t32 VSS 0.0321f
C7127 VREF.t79 VSS 0.0321f
C7128 VREF.n114 VSS 0.233f
C7129 VREF.n115 VSS 0.0876f
C7130 VREF.t167 VSS 0.0321f
C7131 VREF.t77 VSS 0.0321f
C7132 VREF.n116 VSS 0.233f
C7133 VREF.n117 VSS 0.0876f
C7134 VREF.t225 VSS 0.0321f
C7135 VREF.t135 VSS 0.0321f
C7136 VREF.n118 VSS 0.233f
C7137 VREF.n119 VSS 0.0876f
C7138 VREF.t227 VSS 0.0321f
C7139 VREF.t75 VSS 0.0321f
C7140 VREF.n120 VSS 0.233f
C7141 VREF.n121 VSS 0.0876f
C7142 VREF.t71 VSS 0.0321f
C7143 VREF.t205 VSS 0.0321f
C7144 VREF.n122 VSS 0.233f
C7145 VREF.n123 VSS 0.0876f
C7146 VREF.t93 VSS 0.0321f
C7147 VREF.t150 VSS 0.0321f
C7148 VREF.n124 VSS 0.233f
C7149 VREF.n125 VSS 0.0878f
C7150 VREF.t103 VSS 0.0352f
C7151 VREF.t108 VSS 0.0351f
C7152 VREF.n126 VSS 0.208f
C7153 VREF.t155 VSS 0.0351f
C7154 VREF.n127 VSS 0.0555f
C7155 VREF.t245 VSS 0.0351f
C7156 VREF.n128 VSS 0.266f
C7157 VREF.t87 VSS 0.0351f
C7158 VREF.n129 VSS 0.0552f
C7159 VREF.t181 VSS 0.0321f
C7160 VREF.t250 VSS 0.0321f
C7161 VREF.n130 VSS 0.231f
C7162 VREF.n131 VSS 0.0609f
C7163 VREF.t193 VSS 0.0351f
C7164 VREF.n132 VSS 0.286f
C7165 VREF.t88 VSS 0.0351f
C7166 VREF.n133 VSS 0.0552f
C7167 VREF.t80 VSS 0.0321f
C7168 VREF.t147 VSS 0.0321f
C7169 VREF.n134 VSS 0.231f
C7170 VREF.n135 VSS 0.0607f
C7171 VREF.t153 VSS 0.0321f
C7172 VREF.t172 VSS 0.0321f
C7173 VREF.n136 VSS 0.231f
C7174 VREF.n137 VSS 0.0607f
C7175 VREF.t158 VSS 0.0321f
C7176 VREF.t222 VSS 0.0321f
C7177 VREF.n138 VSS 0.231f
C7178 VREF.n139 VSS 0.0609f
C7179 VREF.t35 VSS 0.0351f
C7180 VREF.n140 VSS 0.799f
C7181 VREF.t219 VSS 0.0351f
C7182 VREF.n141 VSS 0.0552f
C7183 VREF.t160 VSS 0.0321f
C7184 VREF.t81 VSS 0.0321f
C7185 VREF.n142 VSS 0.231f
C7186 VREF.n143 VSS 0.0607f
C7187 VREF.t67 VSS 0.0321f
C7188 VREF.t178 VSS 0.0321f
C7189 VREF.n144 VSS 0.231f
C7190 VREF.n145 VSS 0.0607f
C7191 VREF.t248 VSS 0.0321f
C7192 VREF.t113 VSS 0.0321f
C7193 VREF.n146 VSS 0.231f
C7194 VREF.n147 VSS 0.0607f
C7195 VREF.t237 VSS 0.0321f
C7196 VREF.t131 VSS 0.0321f
C7197 VREF.n148 VSS 0.231f
C7198 VREF.n149 VSS 0.0607f
C7199 VREF.t159 VSS 0.0321f
C7200 VREF.t1 VSS 0.0321f
C7201 VREF.n150 VSS 0.231f
C7202 VREF.n151 VSS 0.0607f
C7203 VREF.t112 VSS 0.0321f
C7204 VREF.t117 VSS 0.0321f
C7205 VREF.n152 VSS 0.231f
C7206 VREF.n153 VSS 0.0607f
C7207 VREF.t41 VSS 0.0321f
C7208 VREF.t253 VSS 0.0321f
C7209 VREF.n154 VSS 0.231f
C7210 VREF.n155 VSS 0.0609f
C7211 VREF.t210 VSS 0.0351f
C7212 VREF.n156 VSS 1.26f
C7213 VREF.t162 VSS 0.0351f
C7214 VREF.n157 VSS 0.0552f
C7215 VREF.t56 VSS 0.0321f
C7216 VREF.t46 VSS 0.0321f
C7217 VREF.n158 VSS 0.231f
C7218 VREF.n159 VSS 0.0607f
C7219 VREF.t173 VSS 0.0321f
C7220 VREF.t138 VSS 0.0321f
C7221 VREF.n160 VSS 0.231f
C7222 VREF.n161 VSS 0.0607f
C7223 VREF.t107 VSS 0.0321f
C7224 VREF.t94 VSS 0.0321f
C7225 VREF.n162 VSS 0.231f
C7226 VREF.n163 VSS 0.0607f
C7227 VREF.t246 VSS 0.0321f
C7228 VREF.t97 VSS 0.0321f
C7229 VREF.n164 VSS 0.231f
C7230 VREF.n165 VSS 0.0607f
C7231 VREF.t142 VSS 0.0321f
C7232 VREF.t91 VSS 0.0321f
C7233 VREF.n166 VSS 0.231f
C7234 VREF.n167 VSS 0.0607f
C7235 VREF.t51 VSS 0.0321f
C7236 VREF.t171 VSS 0.0321f
C7237 VREF.n168 VSS 0.231f
C7238 VREF.n169 VSS 0.0607f
C7239 VREF.t65 VSS 0.0321f
C7240 VREF.t161 VSS 0.0321f
C7241 VREF.n170 VSS 0.231f
C7242 VREF.n171 VSS 0.0607f
C7243 VREF.t133 VSS 0.0321f
C7244 VREF.t199 VSS 0.0321f
C7245 VREF.n172 VSS 0.231f
C7246 VREF.n173 VSS 0.0607f
C7247 VREF.t200 VSS 0.0321f
C7248 VREF.t14 VSS 0.0321f
C7249 VREF.n174 VSS 0.231f
C7250 VREF.n175 VSS 0.0607f
C7251 VREF.t174 VSS 0.0321f
C7252 VREF.t151 VSS 0.0321f
C7253 VREF.n176 VSS 0.231f
C7254 VREF.n177 VSS 0.0607f
C7255 VREF.t224 VSS 0.0321f
C7256 VREF.t92 VSS 0.0321f
C7257 VREF.n178 VSS 0.231f
C7258 VREF.n179 VSS 0.0607f
C7259 VREF.t163 VSS 0.0321f
C7260 VREF.t201 VSS 0.0321f
C7261 VREF.n180 VSS 0.231f
C7262 VREF.n181 VSS 0.0607f
C7263 VREF.t104 VSS 0.0321f
C7264 VREF.t4 VSS 0.0321f
C7265 VREF.n182 VSS 0.231f
C7266 VREF.n183 VSS 0.0607f
C7267 VREF.t95 VSS 0.0321f
C7268 VREF.t98 VSS 0.0321f
C7269 VREF.n184 VSS 0.231f
C7270 VREF.n185 VSS 0.0607f
C7271 VREF.t194 VSS 0.0321f
C7272 VREF.t118 VSS 0.0321f
C7273 VREF.n186 VSS 0.231f
C7274 VREF.n187 VSS 0.0609f
C7275 VREF.t168 VSS 0.0351f
C7276 VREF.n188 VSS 2.04f
C7277 VREF.t7 VSS 0.0351f
C7278 VREF.n189 VSS 0.0552f
C7279 VREF.t31 VSS 0.0321f
C7280 VREF.t38 VSS 0.0321f
C7281 VREF.n190 VSS 0.231f
C7282 VREF.n191 VSS 0.0607f
C7283 VREF.t212 VSS 0.0321f
C7284 VREF.t204 VSS 0.0321f
C7285 VREF.n192 VSS 0.231f
C7286 VREF.n193 VSS 0.0607f
C7287 VREF.t209 VSS 0.0321f
C7288 VREF.t22 VSS 0.0321f
C7289 VREF.n194 VSS 0.231f
C7290 VREF.n195 VSS 0.0607f
C7291 VREF.t72 VSS 0.0321f
C7292 VREF.t73 VSS 0.0321f
C7293 VREF.n196 VSS 0.231f
C7294 VREF.n197 VSS 0.0607f
C7295 VREF.t125 VSS 0.0321f
C7296 VREF.t66 VSS 0.0321f
C7297 VREF.n198 VSS 0.231f
C7298 VREF.n199 VSS 0.0607f
C7299 VREF.t16 VSS 0.0321f
C7300 VREF.t59 VSS 0.0321f
C7301 VREF.n200 VSS 0.231f
C7302 VREF.n201 VSS 0.0607f
C7303 VREF.t213 VSS 0.0321f
C7304 VREF.t197 VSS 0.0321f
C7305 VREF.n202 VSS 0.231f
C7306 VREF.n203 VSS 0.0607f
C7307 VREF.t40 VSS 0.0321f
C7308 VREF.t195 VSS 0.0321f
C7309 VREF.n204 VSS 0.231f
C7310 VREF.n205 VSS 0.0607f
C7311 VREF.t84 VSS 0.0321f
C7312 VREF.t251 VSS 0.0321f
C7313 VREF.n206 VSS 0.231f
C7314 VREF.n207 VSS 0.0607f
C7315 VREF.t198 VSS 0.0321f
C7316 VREF.t85 VSS 0.0321f
C7317 VREF.n208 VSS 0.231f
C7318 VREF.n209 VSS 0.0607f
C7319 VREF.t203 VSS 0.0321f
C7320 VREF.t114 VSS 0.0321f
C7321 VREF.n210 VSS 0.231f
C7322 VREF.n211 VSS 0.0607f
C7323 VREF.t8 VSS 0.0321f
C7324 VREF.t238 VSS 0.0321f
C7325 VREF.n212 VSS 0.231f
C7326 VREF.n213 VSS 0.0607f
C7327 VREF.t62 VSS 0.0321f
C7328 VREF.t15 VSS 0.0321f
C7329 VREF.n214 VSS 0.231f
C7330 VREF.n215 VSS 0.0607f
C7331 VREF.t18 VSS 0.0321f
C7332 VREF.t208 VSS 0.0321f
C7333 VREF.n216 VSS 0.231f
C7334 VREF.n217 VSS 0.0607f
C7335 VREF.t123 VSS 0.0321f
C7336 VREF.t239 VSS 0.0321f
C7337 VREF.n218 VSS 0.231f
C7338 VREF.n219 VSS 0.0607f
C7339 VREF.t214 VSS 0.0321f
C7340 VREF.t242 VSS 0.0321f
C7341 VREF.n220 VSS 0.231f
C7342 VREF.n221 VSS 0.0607f
C7343 VREF.t60 VSS 0.0321f
C7344 VREF.t82 VSS 0.0321f
C7345 VREF.n222 VSS 0.231f
C7346 VREF.n223 VSS 0.0607f
C7347 VREF.t179 VSS 0.0321f
C7348 VREF.t216 VSS 0.0321f
C7349 VREF.n224 VSS 0.231f
C7350 VREF.n225 VSS 0.0607f
C7351 VREF.t247 VSS 0.0321f
C7352 VREF.t240 VSS 0.0321f
C7353 VREF.n226 VSS 0.231f
C7354 VREF.n227 VSS 0.0607f
C7355 VREF.t126 VSS 0.0321f
C7356 VREF.t190 VSS 0.0321f
C7357 VREF.n228 VSS 0.231f
C7358 VREF.n229 VSS 0.0607f
C7359 VREF.t130 VSS 0.0321f
C7360 VREF.t109 VSS 0.0321f
C7361 VREF.n230 VSS 0.231f
C7362 VREF.n231 VSS 0.0607f
C7363 VREF.t124 VSS 0.0321f
C7364 VREF.t141 VSS 0.0321f
C7365 VREF.n232 VSS 0.231f
C7366 VREF.n233 VSS 0.0607f
C7367 VREF.t148 VSS 0.0321f
C7368 VREF.t156 VSS 0.0321f
C7369 VREF.n234 VSS 0.231f
C7370 VREF.n235 VSS 0.0607f
C7371 VREF.t27 VSS 0.0321f
C7372 VREF.t34 VSS 0.0321f
C7373 VREF.n236 VSS 0.231f
C7374 VREF.n237 VSS 0.0607f
C7375 VREF.t211 VSS 0.0321f
C7376 VREF.t86 VSS 0.0321f
C7377 VREF.n238 VSS 0.231f
C7378 VREF.n239 VSS 0.0607f
C7379 VREF.t243 VSS 0.0321f
C7380 VREF.t76 VSS 0.0321f
C7381 VREF.n240 VSS 0.231f
C7382 VREF.n241 VSS 0.0607f
C7383 VREF.t25 VSS 0.0321f
C7384 VREF.t119 VSS 0.0321f
C7385 VREF.n242 VSS 0.231f
C7386 VREF.n243 VSS 0.0607f
C7387 VREF.t83 VSS 0.0321f
C7388 VREF.t215 VSS 0.0321f
C7389 VREF.n244 VSS 0.231f
C7390 VREF.n245 VSS 0.0607f
C7391 VREF.t157 VSS 0.0321f
C7392 VREF.t175 VSS 0.0321f
C7393 VREF.n246 VSS 0.231f
C7394 VREF.n247 VSS 0.0607f
C7395 VREF.t241 VSS 0.0321f
C7396 VREF.t58 VSS 0.0321f
C7397 VREF.n248 VSS 0.231f
C7398 VREF.n249 VSS 0.0607f
C7399 VREF.t110 VSS 0.0321f
C7400 VREF.t196 VSS 0.0321f
C7401 VREF.n250 VSS 0.231f
C7402 VREF.n251 VSS 0.0609f
C7403 VREF.t106 VSS 0.0351f
C7404 VREF.n252 VSS 0.15f
C7405 VREF.n253 VSS 2.19f
C7406 VREF.n254 VSS 2.39f
C7407 hgu_cdac_8bit_array_3.drv<7:0>.n0 VSS 0.771f
C7408 hgu_cdac_8bit_array_3.drv<7:0>.n1 VSS 12.7f
C7409 hgu_cdac_8bit_array_3.drv<7:0>.n2 VSS 0.648f
C7410 hgu_cdac_8bit_array_3.drv<7:0>.n3 VSS 0.648f
C7411 hgu_cdac_8bit_array_3.drv<7:0>.n4 VSS 3.18f
C7412 hgu_cdac_8bit_array_3.drv<7:0>.t9 VSS 0.0387f
C7413 hgu_cdac_8bit_array_3.drv<7:0>.t10 VSS 0.0387f
C7414 hgu_cdac_8bit_array_3.drv<7:0>.t5 VSS 0.0773f
C7415 hgu_cdac_8bit_array_3.drv<7:0>.t11 VSS 0.0773f
C7416 hgu_cdac_8bit_array_3.drv<7:0>.n5 VSS 0.589f
C7417 hgu_cdac_8bit_array_3.drv<7:0>.t1 VSS 0.0387f
C7418 hgu_cdac_8bit_array_3.drv<7:0>.t6 VSS 0.0387f
C7419 hgu_cdac_8bit_array_3.drv<7:0>.t13 VSS 0.0773f
C7420 hgu_cdac_8bit_array_3.drv<7:0>.t15 VSS 0.0773f
C7421 hgu_cdac_8bit_array_3.drv<7:0>.n6 VSS 0.589f
C7422 hgu_cdac_8bit_array_3.drv<7:0>.t2 VSS 0.0387f
C7423 hgu_cdac_8bit_array_3.drv<7:0>.t7 VSS 0.0387f
C7424 hgu_cdac_8bit_array_3.drv<7:0>.t14 VSS 0.0773f
C7425 hgu_cdac_8bit_array_3.drv<7:0>.t3 VSS 0.0773f
C7426 hgu_cdac_8bit_array_3.drv<7:0>.n7 VSS 0.516f
C7427 hgu_cdac_8bit_array_3.drv<7:0>.n8 VSS 5.98f
C7428 hgu_cdac_8bit_array_3.drv<7:0>.t8 VSS 0.0387f
C7429 hgu_cdac_8bit_array_3.drv<7:0>.t0 VSS 0.0387f
C7430 hgu_cdac_8bit_array_3.drv<7:0>.t4 VSS 0.0773f
C7431 hgu_cdac_8bit_array_3.drv<7:0>.t12 VSS 0.0773f
C7432 hgu_cdac_8bit_array_3.drv<7:0>.n9 VSS 0.589f
.ends

