magic
tech sky130A
magscale 1 2
timestamp 1699112127
<< pwell >>
rect 1924 1412 1950 1444
rect 2530 1412 2556 1444
rect 3136 1412 3162 1444
rect 3742 1412 3768 1444
rect 4348 1412 4374 1444
rect 4954 1412 4980 1444
rect 5560 1412 5586 1444
rect 6166 1412 6192 1444
rect 1918 -112 1944 -80
rect 2524 -112 2550 -80
rect 3130 -112 3156 -80
rect 3736 -112 3762 -80
rect 4342 -112 4368 -80
rect 4948 -112 4974 -80
rect 5554 -112 5580 -80
rect 6160 -112 6186 -80
<< psubdiff >>
rect 4096 526 4140 608
<< metal3 >>
rect 1598 1858 6512 1860
rect 1598 1794 1702 1858
rect 1766 1794 1782 1858
rect 1846 1794 1862 1858
rect 1926 1794 1942 1858
rect 2006 1794 2022 1858
rect 2086 1794 2102 1858
rect 2166 1794 2308 1858
rect 2372 1794 2388 1858
rect 2452 1794 2468 1858
rect 2532 1794 2548 1858
rect 2612 1794 2628 1858
rect 2692 1794 2708 1858
rect 2772 1794 2914 1858
rect 2978 1794 2994 1858
rect 3058 1794 3074 1858
rect 3138 1794 3154 1858
rect 3218 1794 3234 1858
rect 3298 1794 3314 1858
rect 3378 1794 3520 1858
rect 3584 1794 3600 1858
rect 3664 1794 3680 1858
rect 3744 1794 3760 1858
rect 3824 1794 3840 1858
rect 3904 1794 3920 1858
rect 3984 1794 4126 1858
rect 4190 1794 4206 1858
rect 4270 1794 4286 1858
rect 4350 1794 4366 1858
rect 4430 1794 4446 1858
rect 4510 1794 4526 1858
rect 4590 1794 4732 1858
rect 4796 1794 4812 1858
rect 4876 1794 4892 1858
rect 4956 1794 4972 1858
rect 5036 1794 5052 1858
rect 5116 1794 5132 1858
rect 5196 1794 5338 1858
rect 5402 1794 5418 1858
rect 5482 1794 5498 1858
rect 5562 1794 5578 1858
rect 5642 1794 5658 1858
rect 5722 1794 5738 1858
rect 5802 1794 5944 1858
rect 6008 1794 6024 1858
rect 6088 1794 6104 1858
rect 6168 1794 6184 1858
rect 6248 1794 6264 1858
rect 6328 1794 6344 1858
rect 6408 1794 6512 1858
rect 1598 1792 6512 1794
rect 1598 1638 1664 1728
rect 1598 1574 1599 1638
rect 1663 1574 1664 1638
rect 1598 1558 1664 1574
rect 1598 1494 1599 1558
rect 1663 1494 1664 1558
rect 1598 1478 1664 1494
rect 1598 1414 1599 1478
rect 1663 1414 1664 1478
rect 1598 1398 1664 1414
rect 1598 1334 1599 1398
rect 1663 1334 1664 1398
rect 1598 1318 1664 1334
rect 1598 1254 1599 1318
rect 1663 1254 1664 1318
rect 1598 1238 1664 1254
rect 1598 1174 1599 1238
rect 1663 1174 1664 1238
rect 1598 1158 1664 1174
rect 1598 1094 1599 1158
rect 1663 1094 1664 1158
rect 1598 1078 1664 1094
rect 1598 1014 1599 1078
rect 1663 1014 1664 1078
rect 1598 998 1664 1014
rect 1598 934 1599 998
rect 1663 934 1664 998
rect 1598 918 1664 934
rect 1598 854 1599 918
rect 1663 854 1664 918
rect 1598 700 1664 854
rect 1724 762 1784 1792
rect 1844 700 1904 1732
rect 1964 762 2024 1792
rect 2084 700 2144 1732
rect 2204 1638 2270 1728
rect 2204 1574 2205 1638
rect 2269 1574 2270 1638
rect 2204 1558 2270 1574
rect 2204 1494 2205 1558
rect 2269 1494 2270 1558
rect 2204 1478 2270 1494
rect 2204 1414 2205 1478
rect 2269 1414 2270 1478
rect 2204 1398 2270 1414
rect 2204 1334 2205 1398
rect 2269 1334 2270 1398
rect 2204 1318 2270 1334
rect 2204 1254 2205 1318
rect 2269 1254 2270 1318
rect 2204 1238 2270 1254
rect 2204 1174 2205 1238
rect 2269 1174 2270 1238
rect 2204 1158 2270 1174
rect 2204 1094 2205 1158
rect 2269 1094 2270 1158
rect 2204 1078 2270 1094
rect 2204 1014 2205 1078
rect 2269 1014 2270 1078
rect 2204 998 2270 1014
rect 2204 934 2205 998
rect 2269 934 2270 998
rect 2204 918 2270 934
rect 2204 854 2205 918
rect 2269 854 2270 918
rect 2204 700 2270 854
rect 2330 762 2390 1792
rect 2450 700 2510 1732
rect 2570 762 2630 1792
rect 2690 700 2750 1732
rect 2810 1638 2876 1728
rect 2810 1574 2811 1638
rect 2875 1574 2876 1638
rect 2810 1558 2876 1574
rect 2810 1494 2811 1558
rect 2875 1494 2876 1558
rect 2810 1478 2876 1494
rect 2810 1414 2811 1478
rect 2875 1414 2876 1478
rect 2810 1398 2876 1414
rect 2810 1334 2811 1398
rect 2875 1334 2876 1398
rect 2810 1318 2876 1334
rect 2810 1254 2811 1318
rect 2875 1254 2876 1318
rect 2810 1238 2876 1254
rect 2810 1174 2811 1238
rect 2875 1174 2876 1238
rect 2810 1158 2876 1174
rect 2810 1094 2811 1158
rect 2875 1094 2876 1158
rect 2810 1078 2876 1094
rect 2810 1014 2811 1078
rect 2875 1014 2876 1078
rect 2810 998 2876 1014
rect 2810 934 2811 998
rect 2875 934 2876 998
rect 2810 918 2876 934
rect 2810 854 2811 918
rect 2875 854 2876 918
rect 2810 700 2876 854
rect 2936 762 2996 1792
rect 3056 700 3116 1732
rect 3176 762 3236 1792
rect 3296 700 3356 1732
rect 3416 1638 3482 1728
rect 3416 1574 3417 1638
rect 3481 1574 3482 1638
rect 3416 1558 3482 1574
rect 3416 1494 3417 1558
rect 3481 1494 3482 1558
rect 3416 1478 3482 1494
rect 3416 1414 3417 1478
rect 3481 1414 3482 1478
rect 3416 1398 3482 1414
rect 3416 1334 3417 1398
rect 3481 1334 3482 1398
rect 3416 1318 3482 1334
rect 3416 1254 3417 1318
rect 3481 1254 3482 1318
rect 3416 1238 3482 1254
rect 3416 1174 3417 1238
rect 3481 1174 3482 1238
rect 3416 1158 3482 1174
rect 3416 1094 3417 1158
rect 3481 1094 3482 1158
rect 3416 1078 3482 1094
rect 3416 1014 3417 1078
rect 3481 1014 3482 1078
rect 3416 998 3482 1014
rect 3416 934 3417 998
rect 3481 934 3482 998
rect 3416 918 3482 934
rect 3416 854 3417 918
rect 3481 854 3482 918
rect 3416 700 3482 854
rect 3542 762 3602 1792
rect 3662 700 3722 1732
rect 3782 762 3842 1792
rect 3902 700 3962 1732
rect 4022 1638 4088 1728
rect 4022 1574 4023 1638
rect 4087 1574 4088 1638
rect 4022 1558 4088 1574
rect 4022 1494 4023 1558
rect 4087 1494 4088 1558
rect 4022 1478 4088 1494
rect 4022 1414 4023 1478
rect 4087 1414 4088 1478
rect 4022 1398 4088 1414
rect 4022 1334 4023 1398
rect 4087 1334 4088 1398
rect 4022 1318 4088 1334
rect 4022 1254 4023 1318
rect 4087 1254 4088 1318
rect 4022 1238 4088 1254
rect 4022 1174 4023 1238
rect 4087 1174 4088 1238
rect 4022 1158 4088 1174
rect 4022 1094 4023 1158
rect 4087 1094 4088 1158
rect 4022 1078 4088 1094
rect 4022 1014 4023 1078
rect 4087 1014 4088 1078
rect 4022 998 4088 1014
rect 4022 934 4023 998
rect 4087 934 4088 998
rect 4022 918 4088 934
rect 4022 854 4023 918
rect 4087 854 4088 918
rect 4022 700 4088 854
rect 4148 762 4208 1792
rect 4268 700 4328 1732
rect 4388 762 4448 1792
rect 4508 700 4568 1732
rect 4628 1638 4694 1728
rect 4628 1574 4629 1638
rect 4693 1574 4694 1638
rect 4628 1558 4694 1574
rect 4628 1494 4629 1558
rect 4693 1494 4694 1558
rect 4628 1478 4694 1494
rect 4628 1414 4629 1478
rect 4693 1414 4694 1478
rect 4628 1398 4694 1414
rect 4628 1334 4629 1398
rect 4693 1334 4694 1398
rect 4628 1318 4694 1334
rect 4628 1254 4629 1318
rect 4693 1254 4694 1318
rect 4628 1238 4694 1254
rect 4628 1174 4629 1238
rect 4693 1174 4694 1238
rect 4628 1158 4694 1174
rect 4628 1094 4629 1158
rect 4693 1094 4694 1158
rect 4628 1078 4694 1094
rect 4628 1014 4629 1078
rect 4693 1014 4694 1078
rect 4628 998 4694 1014
rect 4628 934 4629 998
rect 4693 934 4694 998
rect 4628 918 4694 934
rect 4628 854 4629 918
rect 4693 854 4694 918
rect 4628 700 4694 854
rect 4754 762 4814 1792
rect 4874 700 4934 1732
rect 4994 762 5054 1792
rect 5114 700 5174 1732
rect 5234 1638 5300 1728
rect 5234 1574 5235 1638
rect 5299 1574 5300 1638
rect 5234 1558 5300 1574
rect 5234 1494 5235 1558
rect 5299 1494 5300 1558
rect 5234 1478 5300 1494
rect 5234 1414 5235 1478
rect 5299 1414 5300 1478
rect 5234 1398 5300 1414
rect 5234 1334 5235 1398
rect 5299 1334 5300 1398
rect 5234 1318 5300 1334
rect 5234 1254 5235 1318
rect 5299 1254 5300 1318
rect 5234 1238 5300 1254
rect 5234 1174 5235 1238
rect 5299 1174 5300 1238
rect 5234 1158 5300 1174
rect 5234 1094 5235 1158
rect 5299 1094 5300 1158
rect 5234 1078 5300 1094
rect 5234 1014 5235 1078
rect 5299 1014 5300 1078
rect 5234 998 5300 1014
rect 5234 934 5235 998
rect 5299 934 5300 998
rect 5234 918 5300 934
rect 5234 854 5235 918
rect 5299 854 5300 918
rect 5234 700 5300 854
rect 5360 762 5420 1792
rect 5480 700 5540 1732
rect 5600 762 5660 1792
rect 5720 700 5780 1732
rect 5840 1638 5906 1728
rect 5840 1574 5841 1638
rect 5905 1574 5906 1638
rect 5840 1558 5906 1574
rect 5840 1494 5841 1558
rect 5905 1494 5906 1558
rect 5840 1478 5906 1494
rect 5840 1414 5841 1478
rect 5905 1414 5906 1478
rect 5840 1398 5906 1414
rect 5840 1334 5841 1398
rect 5905 1334 5906 1398
rect 5840 1318 5906 1334
rect 5840 1254 5841 1318
rect 5905 1254 5906 1318
rect 5840 1238 5906 1254
rect 5840 1174 5841 1238
rect 5905 1174 5906 1238
rect 5840 1158 5906 1174
rect 5840 1094 5841 1158
rect 5905 1094 5906 1158
rect 5840 1078 5906 1094
rect 5840 1014 5841 1078
rect 5905 1014 5906 1078
rect 5840 998 5906 1014
rect 5840 934 5841 998
rect 5905 934 5906 998
rect 5840 918 5906 934
rect 5840 854 5841 918
rect 5905 854 5906 918
rect 5840 700 5906 854
rect 5966 762 6026 1792
rect 6086 700 6146 1732
rect 6206 762 6266 1792
rect 6326 700 6386 1732
rect 6446 1638 6512 1728
rect 6446 1574 6447 1638
rect 6511 1574 6512 1638
rect 6446 1558 6512 1574
rect 6446 1494 6447 1558
rect 6511 1494 6512 1558
rect 6446 1478 6512 1494
rect 6446 1414 6447 1478
rect 6511 1414 6512 1478
rect 6446 1398 6512 1414
rect 6446 1334 6447 1398
rect 6511 1334 6512 1398
rect 6446 1318 6512 1334
rect 6446 1254 6447 1318
rect 6511 1254 6512 1318
rect 6446 1238 6512 1254
rect 6446 1174 6447 1238
rect 6511 1174 6512 1238
rect 6446 1158 6512 1174
rect 6446 1094 6447 1158
rect 6511 1094 6512 1158
rect 6446 1078 6512 1094
rect 6446 1014 6447 1078
rect 6511 1014 6512 1078
rect 6446 998 6512 1014
rect 6446 934 6447 998
rect 6511 934 6512 998
rect 6446 918 6512 934
rect 6446 854 6447 918
rect 6511 854 6512 918
rect 6446 700 6512 854
rect 1598 698 6512 700
rect 1598 634 1702 698
rect 1766 634 1782 698
rect 1846 634 1862 698
rect 1926 634 1942 698
rect 2006 634 2022 698
rect 2086 634 2102 698
rect 2166 634 2308 698
rect 2372 634 2388 698
rect 2452 634 2468 698
rect 2532 634 2548 698
rect 2612 634 2628 698
rect 2692 634 2708 698
rect 2772 634 2914 698
rect 2978 634 2994 698
rect 3058 634 3074 698
rect 3138 634 3154 698
rect 3218 634 3234 698
rect 3298 634 3314 698
rect 3378 634 3520 698
rect 3584 634 3600 698
rect 3664 634 3680 698
rect 3744 634 3760 698
rect 3824 634 3840 698
rect 3904 634 3920 698
rect 3984 634 4126 698
rect 4190 634 4206 698
rect 4270 634 4286 698
rect 4350 634 4366 698
rect 4430 634 4446 698
rect 4510 634 4526 698
rect 4590 634 4732 698
rect 4796 634 4812 698
rect 4876 634 4892 698
rect 4956 634 4972 698
rect 5036 634 5052 698
rect 5116 634 5132 698
rect 5196 634 5338 698
rect 5402 634 5418 698
rect 5482 634 5498 698
rect 5562 634 5578 698
rect 5642 634 5658 698
rect 5722 634 5738 698
rect 5802 634 5944 698
rect 6008 634 6024 698
rect 6088 634 6104 698
rect 6168 634 6184 698
rect 6248 634 6264 698
rect 6328 634 6344 698
rect 6408 634 6512 698
rect 1598 632 6512 634
rect 1598 478 1664 632
rect 1598 414 1599 478
rect 1663 414 1664 478
rect 1598 398 1664 414
rect 1598 334 1599 398
rect 1663 334 1664 398
rect 1598 318 1664 334
rect 1598 254 1599 318
rect 1663 254 1664 318
rect 1598 238 1664 254
rect 1598 174 1599 238
rect 1663 174 1664 238
rect 1598 158 1664 174
rect 1598 94 1599 158
rect 1663 94 1664 158
rect 1598 78 1664 94
rect 1598 14 1599 78
rect 1663 14 1664 78
rect 1598 -2 1664 14
rect 1598 -66 1599 -2
rect 1663 -66 1664 -2
rect 1598 -82 1664 -66
rect 1598 -146 1599 -82
rect 1663 -146 1664 -82
rect 1598 -162 1664 -146
rect 1598 -226 1599 -162
rect 1663 -226 1664 -162
rect 1598 -242 1664 -226
rect 1598 -306 1599 -242
rect 1663 -306 1664 -242
rect 1598 -396 1664 -306
rect 1724 -400 1784 632
rect 1844 -460 1904 570
rect 1964 -400 2024 632
rect 2084 -460 2144 570
rect 2204 478 2270 632
rect 2204 414 2205 478
rect 2269 414 2270 478
rect 2204 398 2270 414
rect 2204 334 2205 398
rect 2269 334 2270 398
rect 2204 318 2270 334
rect 2204 254 2205 318
rect 2269 254 2270 318
rect 2204 238 2270 254
rect 2204 174 2205 238
rect 2269 174 2270 238
rect 2204 158 2270 174
rect 2204 94 2205 158
rect 2269 94 2270 158
rect 2204 78 2270 94
rect 2204 14 2205 78
rect 2269 14 2270 78
rect 2204 -2 2270 14
rect 2204 -66 2205 -2
rect 2269 -66 2270 -2
rect 2204 -82 2270 -66
rect 2204 -146 2205 -82
rect 2269 -146 2270 -82
rect 2204 -162 2270 -146
rect 2204 -226 2205 -162
rect 2269 -226 2270 -162
rect 2204 -242 2270 -226
rect 2204 -306 2205 -242
rect 2269 -306 2270 -242
rect 2204 -396 2270 -306
rect 2330 -400 2390 632
rect 2450 -460 2510 570
rect 2570 -400 2630 632
rect 2690 -460 2750 570
rect 2810 478 2876 632
rect 2810 414 2811 478
rect 2875 414 2876 478
rect 2810 398 2876 414
rect 2810 334 2811 398
rect 2875 334 2876 398
rect 2810 318 2876 334
rect 2810 254 2811 318
rect 2875 254 2876 318
rect 2810 238 2876 254
rect 2810 174 2811 238
rect 2875 174 2876 238
rect 2810 158 2876 174
rect 2810 94 2811 158
rect 2875 94 2876 158
rect 2810 78 2876 94
rect 2810 14 2811 78
rect 2875 14 2876 78
rect 2810 -2 2876 14
rect 2810 -66 2811 -2
rect 2875 -66 2876 -2
rect 2810 -82 2876 -66
rect 2810 -146 2811 -82
rect 2875 -146 2876 -82
rect 2810 -162 2876 -146
rect 2810 -226 2811 -162
rect 2875 -226 2876 -162
rect 2810 -242 2876 -226
rect 2810 -306 2811 -242
rect 2875 -306 2876 -242
rect 2810 -396 2876 -306
rect 2936 -400 2996 632
rect 3056 -460 3116 570
rect 3176 -400 3236 632
rect 3296 -460 3356 570
rect 3416 478 3482 632
rect 3416 414 3417 478
rect 3481 414 3482 478
rect 3416 398 3482 414
rect 3416 334 3417 398
rect 3481 334 3482 398
rect 3416 318 3482 334
rect 3416 254 3417 318
rect 3481 254 3482 318
rect 3416 238 3482 254
rect 3416 174 3417 238
rect 3481 174 3482 238
rect 3416 158 3482 174
rect 3416 94 3417 158
rect 3481 94 3482 158
rect 3416 78 3482 94
rect 3416 14 3417 78
rect 3481 14 3482 78
rect 3416 -2 3482 14
rect 3416 -66 3417 -2
rect 3481 -66 3482 -2
rect 3416 -82 3482 -66
rect 3416 -146 3417 -82
rect 3481 -146 3482 -82
rect 3416 -162 3482 -146
rect 3416 -226 3417 -162
rect 3481 -226 3482 -162
rect 3416 -242 3482 -226
rect 3416 -306 3417 -242
rect 3481 -306 3482 -242
rect 3416 -396 3482 -306
rect 3542 -400 3602 632
rect 3662 -460 3722 570
rect 3782 -400 3842 632
rect 3902 -460 3962 570
rect 4022 478 4088 632
rect 4022 414 4023 478
rect 4087 414 4088 478
rect 4022 398 4088 414
rect 4022 334 4023 398
rect 4087 334 4088 398
rect 4022 318 4088 334
rect 4022 254 4023 318
rect 4087 254 4088 318
rect 4022 238 4088 254
rect 4022 174 4023 238
rect 4087 174 4088 238
rect 4022 158 4088 174
rect 4022 94 4023 158
rect 4087 94 4088 158
rect 4022 78 4088 94
rect 4022 14 4023 78
rect 4087 14 4088 78
rect 4022 -2 4088 14
rect 4022 -66 4023 -2
rect 4087 -66 4088 -2
rect 4022 -82 4088 -66
rect 4022 -146 4023 -82
rect 4087 -146 4088 -82
rect 4022 -162 4088 -146
rect 4022 -226 4023 -162
rect 4087 -226 4088 -162
rect 4022 -242 4088 -226
rect 4022 -306 4023 -242
rect 4087 -306 4088 -242
rect 4022 -396 4088 -306
rect 4148 -400 4208 632
rect 4268 -460 4328 570
rect 4388 -400 4448 632
rect 4508 -460 4568 570
rect 4628 478 4694 632
rect 4628 414 4629 478
rect 4693 414 4694 478
rect 4628 398 4694 414
rect 4628 334 4629 398
rect 4693 334 4694 398
rect 4628 318 4694 334
rect 4628 254 4629 318
rect 4693 254 4694 318
rect 4628 238 4694 254
rect 4628 174 4629 238
rect 4693 174 4694 238
rect 4628 158 4694 174
rect 4628 94 4629 158
rect 4693 94 4694 158
rect 4628 78 4694 94
rect 4628 14 4629 78
rect 4693 14 4694 78
rect 4628 -2 4694 14
rect 4628 -66 4629 -2
rect 4693 -66 4694 -2
rect 4628 -82 4694 -66
rect 4628 -146 4629 -82
rect 4693 -146 4694 -82
rect 4628 -162 4694 -146
rect 4628 -226 4629 -162
rect 4693 -226 4694 -162
rect 4628 -242 4694 -226
rect 4628 -306 4629 -242
rect 4693 -306 4694 -242
rect 4628 -396 4694 -306
rect 4754 -400 4814 632
rect 4874 -460 4934 570
rect 4994 -400 5054 632
rect 5114 -460 5174 570
rect 5234 478 5300 632
rect 5234 414 5235 478
rect 5299 414 5300 478
rect 5234 398 5300 414
rect 5234 334 5235 398
rect 5299 334 5300 398
rect 5234 318 5300 334
rect 5234 254 5235 318
rect 5299 254 5300 318
rect 5234 238 5300 254
rect 5234 174 5235 238
rect 5299 174 5300 238
rect 5234 158 5300 174
rect 5234 94 5235 158
rect 5299 94 5300 158
rect 5234 78 5300 94
rect 5234 14 5235 78
rect 5299 14 5300 78
rect 5234 -2 5300 14
rect 5234 -66 5235 -2
rect 5299 -66 5300 -2
rect 5234 -82 5300 -66
rect 5234 -146 5235 -82
rect 5299 -146 5300 -82
rect 5234 -162 5300 -146
rect 5234 -226 5235 -162
rect 5299 -226 5300 -162
rect 5234 -242 5300 -226
rect 5234 -306 5235 -242
rect 5299 -306 5300 -242
rect 5234 -396 5300 -306
rect 5360 -400 5420 632
rect 5480 -460 5540 570
rect 5600 -400 5660 632
rect 5720 -460 5780 570
rect 5840 478 5906 632
rect 5840 414 5841 478
rect 5905 414 5906 478
rect 5840 398 5906 414
rect 5840 334 5841 398
rect 5905 334 5906 398
rect 5840 318 5906 334
rect 5840 254 5841 318
rect 5905 254 5906 318
rect 5840 238 5906 254
rect 5840 174 5841 238
rect 5905 174 5906 238
rect 5840 158 5906 174
rect 5840 94 5841 158
rect 5905 94 5906 158
rect 5840 78 5906 94
rect 5840 14 5841 78
rect 5905 14 5906 78
rect 5840 -2 5906 14
rect 5840 -66 5841 -2
rect 5905 -66 5906 -2
rect 5840 -82 5906 -66
rect 5840 -146 5841 -82
rect 5905 -146 5906 -82
rect 5840 -162 5906 -146
rect 5840 -226 5841 -162
rect 5905 -226 5906 -162
rect 5840 -242 5906 -226
rect 5840 -306 5841 -242
rect 5905 -306 5906 -242
rect 5840 -396 5906 -306
rect 5966 -400 6026 632
rect 6086 -460 6146 570
rect 6206 -400 6266 632
rect 6326 -460 6386 570
rect 6446 478 6512 632
rect 6446 414 6447 478
rect 6511 414 6512 478
rect 6446 398 6512 414
rect 6446 334 6447 398
rect 6511 334 6512 398
rect 6446 318 6512 334
rect 6446 254 6447 318
rect 6511 254 6512 318
rect 6446 238 6512 254
rect 6446 174 6447 238
rect 6511 174 6512 238
rect 6446 158 6512 174
rect 6446 94 6447 158
rect 6511 94 6512 158
rect 6446 78 6512 94
rect 6446 14 6447 78
rect 6511 14 6512 78
rect 6446 -2 6512 14
rect 6446 -66 6447 -2
rect 6511 -66 6512 -2
rect 6446 -82 6512 -66
rect 6446 -146 6447 -82
rect 6511 -146 6512 -82
rect 6446 -162 6512 -146
rect 6446 -226 6447 -162
rect 6511 -226 6512 -162
rect 6446 -242 6512 -226
rect 6446 -306 6447 -242
rect 6511 -306 6512 -242
rect 6446 -396 6512 -306
rect 1598 -462 6512 -460
rect 1598 -526 1702 -462
rect 1766 -526 1782 -462
rect 1846 -526 1862 -462
rect 1926 -526 1942 -462
rect 2006 -526 2022 -462
rect 2086 -526 2102 -462
rect 2166 -526 2308 -462
rect 2372 -526 2388 -462
rect 2452 -526 2468 -462
rect 2532 -526 2548 -462
rect 2612 -526 2628 -462
rect 2692 -526 2708 -462
rect 2772 -526 2914 -462
rect 2978 -526 2994 -462
rect 3058 -526 3074 -462
rect 3138 -526 3154 -462
rect 3218 -526 3234 -462
rect 3298 -526 3314 -462
rect 3378 -526 3520 -462
rect 3584 -526 3600 -462
rect 3664 -526 3680 -462
rect 3744 -526 3760 -462
rect 3824 -526 3840 -462
rect 3904 -526 3920 -462
rect 3984 -526 4126 -462
rect 4190 -526 4206 -462
rect 4270 -526 4286 -462
rect 4350 -526 4366 -462
rect 4430 -526 4446 -462
rect 4510 -526 4526 -462
rect 4590 -526 4732 -462
rect 4796 -526 4812 -462
rect 4876 -526 4892 -462
rect 4956 -526 4972 -462
rect 5036 -526 5052 -462
rect 5116 -526 5132 -462
rect 5196 -526 5338 -462
rect 5402 -526 5418 -462
rect 5482 -526 5498 -462
rect 5562 -526 5578 -462
rect 5642 -526 5658 -462
rect 5722 -526 5738 -462
rect 5802 -526 5944 -462
rect 6008 -526 6024 -462
rect 6088 -526 6104 -462
rect 6168 -526 6184 -462
rect 6248 -526 6264 -462
rect 6328 -526 6344 -462
rect 6408 -526 6512 -462
rect 1598 -528 6512 -526
<< via3 >>
rect 1702 1794 1766 1858
rect 1782 1794 1846 1858
rect 1862 1794 1926 1858
rect 1942 1794 2006 1858
rect 2022 1794 2086 1858
rect 2102 1794 2166 1858
rect 2308 1794 2372 1858
rect 2388 1794 2452 1858
rect 2468 1794 2532 1858
rect 2548 1794 2612 1858
rect 2628 1794 2692 1858
rect 2708 1794 2772 1858
rect 2914 1794 2978 1858
rect 2994 1794 3058 1858
rect 3074 1794 3138 1858
rect 3154 1794 3218 1858
rect 3234 1794 3298 1858
rect 3314 1794 3378 1858
rect 3520 1794 3584 1858
rect 3600 1794 3664 1858
rect 3680 1794 3744 1858
rect 3760 1794 3824 1858
rect 3840 1794 3904 1858
rect 3920 1794 3984 1858
rect 4126 1794 4190 1858
rect 4206 1794 4270 1858
rect 4286 1794 4350 1858
rect 4366 1794 4430 1858
rect 4446 1794 4510 1858
rect 4526 1794 4590 1858
rect 4732 1794 4796 1858
rect 4812 1794 4876 1858
rect 4892 1794 4956 1858
rect 4972 1794 5036 1858
rect 5052 1794 5116 1858
rect 5132 1794 5196 1858
rect 5338 1794 5402 1858
rect 5418 1794 5482 1858
rect 5498 1794 5562 1858
rect 5578 1794 5642 1858
rect 5658 1794 5722 1858
rect 5738 1794 5802 1858
rect 5944 1794 6008 1858
rect 6024 1794 6088 1858
rect 6104 1794 6168 1858
rect 6184 1794 6248 1858
rect 6264 1794 6328 1858
rect 6344 1794 6408 1858
rect 1599 1574 1663 1638
rect 1599 1494 1663 1558
rect 1599 1414 1663 1478
rect 1599 1334 1663 1398
rect 1599 1254 1663 1318
rect 1599 1174 1663 1238
rect 1599 1094 1663 1158
rect 1599 1014 1663 1078
rect 1599 934 1663 998
rect 1599 854 1663 918
rect 2205 1574 2269 1638
rect 2205 1494 2269 1558
rect 2205 1414 2269 1478
rect 2205 1334 2269 1398
rect 2205 1254 2269 1318
rect 2205 1174 2269 1238
rect 2205 1094 2269 1158
rect 2205 1014 2269 1078
rect 2205 934 2269 998
rect 2205 854 2269 918
rect 2811 1574 2875 1638
rect 2811 1494 2875 1558
rect 2811 1414 2875 1478
rect 2811 1334 2875 1398
rect 2811 1254 2875 1318
rect 2811 1174 2875 1238
rect 2811 1094 2875 1158
rect 2811 1014 2875 1078
rect 2811 934 2875 998
rect 2811 854 2875 918
rect 3417 1574 3481 1638
rect 3417 1494 3481 1558
rect 3417 1414 3481 1478
rect 3417 1334 3481 1398
rect 3417 1254 3481 1318
rect 3417 1174 3481 1238
rect 3417 1094 3481 1158
rect 3417 1014 3481 1078
rect 3417 934 3481 998
rect 3417 854 3481 918
rect 4023 1574 4087 1638
rect 4023 1494 4087 1558
rect 4023 1414 4087 1478
rect 4023 1334 4087 1398
rect 4023 1254 4087 1318
rect 4023 1174 4087 1238
rect 4023 1094 4087 1158
rect 4023 1014 4087 1078
rect 4023 934 4087 998
rect 4023 854 4087 918
rect 4629 1574 4693 1638
rect 4629 1494 4693 1558
rect 4629 1414 4693 1478
rect 4629 1334 4693 1398
rect 4629 1254 4693 1318
rect 4629 1174 4693 1238
rect 4629 1094 4693 1158
rect 4629 1014 4693 1078
rect 4629 934 4693 998
rect 4629 854 4693 918
rect 5235 1574 5299 1638
rect 5235 1494 5299 1558
rect 5235 1414 5299 1478
rect 5235 1334 5299 1398
rect 5235 1254 5299 1318
rect 5235 1174 5299 1238
rect 5235 1094 5299 1158
rect 5235 1014 5299 1078
rect 5235 934 5299 998
rect 5235 854 5299 918
rect 5841 1574 5905 1638
rect 5841 1494 5905 1558
rect 5841 1414 5905 1478
rect 5841 1334 5905 1398
rect 5841 1254 5905 1318
rect 5841 1174 5905 1238
rect 5841 1094 5905 1158
rect 5841 1014 5905 1078
rect 5841 934 5905 998
rect 5841 854 5905 918
rect 6447 1574 6511 1638
rect 6447 1494 6511 1558
rect 6447 1414 6511 1478
rect 6447 1334 6511 1398
rect 6447 1254 6511 1318
rect 6447 1174 6511 1238
rect 6447 1094 6511 1158
rect 6447 1014 6511 1078
rect 6447 934 6511 998
rect 6447 854 6511 918
rect 1702 634 1766 698
rect 1782 634 1846 698
rect 1862 634 1926 698
rect 1942 634 2006 698
rect 2022 634 2086 698
rect 2102 634 2166 698
rect 2308 634 2372 698
rect 2388 634 2452 698
rect 2468 634 2532 698
rect 2548 634 2612 698
rect 2628 634 2692 698
rect 2708 634 2772 698
rect 2914 634 2978 698
rect 2994 634 3058 698
rect 3074 634 3138 698
rect 3154 634 3218 698
rect 3234 634 3298 698
rect 3314 634 3378 698
rect 3520 634 3584 698
rect 3600 634 3664 698
rect 3680 634 3744 698
rect 3760 634 3824 698
rect 3840 634 3904 698
rect 3920 634 3984 698
rect 4126 634 4190 698
rect 4206 634 4270 698
rect 4286 634 4350 698
rect 4366 634 4430 698
rect 4446 634 4510 698
rect 4526 634 4590 698
rect 4732 634 4796 698
rect 4812 634 4876 698
rect 4892 634 4956 698
rect 4972 634 5036 698
rect 5052 634 5116 698
rect 5132 634 5196 698
rect 5338 634 5402 698
rect 5418 634 5482 698
rect 5498 634 5562 698
rect 5578 634 5642 698
rect 5658 634 5722 698
rect 5738 634 5802 698
rect 5944 634 6008 698
rect 6024 634 6088 698
rect 6104 634 6168 698
rect 6184 634 6248 698
rect 6264 634 6328 698
rect 6344 634 6408 698
rect 1599 414 1663 478
rect 1599 334 1663 398
rect 1599 254 1663 318
rect 1599 174 1663 238
rect 1599 94 1663 158
rect 1599 14 1663 78
rect 1599 -66 1663 -2
rect 1599 -146 1663 -82
rect 1599 -226 1663 -162
rect 1599 -306 1663 -242
rect 2205 414 2269 478
rect 2205 334 2269 398
rect 2205 254 2269 318
rect 2205 174 2269 238
rect 2205 94 2269 158
rect 2205 14 2269 78
rect 2205 -66 2269 -2
rect 2205 -146 2269 -82
rect 2205 -226 2269 -162
rect 2205 -306 2269 -242
rect 2811 414 2875 478
rect 2811 334 2875 398
rect 2811 254 2875 318
rect 2811 174 2875 238
rect 2811 94 2875 158
rect 2811 14 2875 78
rect 2811 -66 2875 -2
rect 2811 -146 2875 -82
rect 2811 -226 2875 -162
rect 2811 -306 2875 -242
rect 3417 414 3481 478
rect 3417 334 3481 398
rect 3417 254 3481 318
rect 3417 174 3481 238
rect 3417 94 3481 158
rect 3417 14 3481 78
rect 3417 -66 3481 -2
rect 3417 -146 3481 -82
rect 3417 -226 3481 -162
rect 3417 -306 3481 -242
rect 4023 414 4087 478
rect 4023 334 4087 398
rect 4023 254 4087 318
rect 4023 174 4087 238
rect 4023 94 4087 158
rect 4023 14 4087 78
rect 4023 -66 4087 -2
rect 4023 -146 4087 -82
rect 4023 -226 4087 -162
rect 4023 -306 4087 -242
rect 4629 414 4693 478
rect 4629 334 4693 398
rect 4629 254 4693 318
rect 4629 174 4693 238
rect 4629 94 4693 158
rect 4629 14 4693 78
rect 4629 -66 4693 -2
rect 4629 -146 4693 -82
rect 4629 -226 4693 -162
rect 4629 -306 4693 -242
rect 5235 414 5299 478
rect 5235 334 5299 398
rect 5235 254 5299 318
rect 5235 174 5299 238
rect 5235 94 5299 158
rect 5235 14 5299 78
rect 5235 -66 5299 -2
rect 5235 -146 5299 -82
rect 5235 -226 5299 -162
rect 5235 -306 5299 -242
rect 5841 414 5905 478
rect 5841 334 5905 398
rect 5841 254 5905 318
rect 5841 174 5905 238
rect 5841 94 5905 158
rect 5841 14 5905 78
rect 5841 -66 5905 -2
rect 5841 -146 5905 -82
rect 5841 -226 5905 -162
rect 5841 -306 5905 -242
rect 6447 414 6511 478
rect 6447 334 6511 398
rect 6447 254 6511 318
rect 6447 174 6511 238
rect 6447 94 6511 158
rect 6447 14 6511 78
rect 6447 -66 6511 -2
rect 6447 -146 6511 -82
rect 6447 -226 6511 -162
rect 6447 -306 6511 -242
rect 1702 -526 1766 -462
rect 1782 -526 1846 -462
rect 1862 -526 1926 -462
rect 1942 -526 2006 -462
rect 2022 -526 2086 -462
rect 2102 -526 2166 -462
rect 2308 -526 2372 -462
rect 2388 -526 2452 -462
rect 2468 -526 2532 -462
rect 2548 -526 2612 -462
rect 2628 -526 2692 -462
rect 2708 -526 2772 -462
rect 2914 -526 2978 -462
rect 2994 -526 3058 -462
rect 3074 -526 3138 -462
rect 3154 -526 3218 -462
rect 3234 -526 3298 -462
rect 3314 -526 3378 -462
rect 3520 -526 3584 -462
rect 3600 -526 3664 -462
rect 3680 -526 3744 -462
rect 3760 -526 3824 -462
rect 3840 -526 3904 -462
rect 3920 -526 3984 -462
rect 4126 -526 4190 -462
rect 4206 -526 4270 -462
rect 4286 -526 4350 -462
rect 4366 -526 4430 -462
rect 4446 -526 4510 -462
rect 4526 -526 4590 -462
rect 4732 -526 4796 -462
rect 4812 -526 4876 -462
rect 4892 -526 4956 -462
rect 4972 -526 5036 -462
rect 5052 -526 5116 -462
rect 5132 -526 5196 -462
rect 5338 -526 5402 -462
rect 5418 -526 5482 -462
rect 5498 -526 5562 -462
rect 5578 -526 5642 -462
rect 5658 -526 5722 -462
rect 5738 -526 5802 -462
rect 5944 -526 6008 -462
rect 6024 -526 6088 -462
rect 6104 -526 6168 -462
rect 6184 -526 6248 -462
rect 6264 -526 6328 -462
rect 6344 -526 6408 -462
<< metal4 >>
rect 1598 1858 6512 1860
rect 1598 1794 1702 1858
rect 1766 1794 1782 1858
rect 1846 1794 1862 1858
rect 1926 1794 1942 1858
rect 2006 1794 2022 1858
rect 2086 1794 2102 1858
rect 2166 1794 2308 1858
rect 2372 1794 2388 1858
rect 2452 1794 2468 1858
rect 2532 1794 2548 1858
rect 2612 1794 2628 1858
rect 2692 1794 2708 1858
rect 2772 1794 2914 1858
rect 2978 1794 2994 1858
rect 3058 1794 3074 1858
rect 3138 1794 3154 1858
rect 3218 1794 3234 1858
rect 3298 1794 3314 1858
rect 3378 1794 3520 1858
rect 3584 1794 3600 1858
rect 3664 1794 3680 1858
rect 3744 1794 3760 1858
rect 3824 1794 3840 1858
rect 3904 1794 3920 1858
rect 3984 1794 4126 1858
rect 4190 1794 4206 1858
rect 4270 1794 4286 1858
rect 4350 1794 4366 1858
rect 4430 1794 4446 1858
rect 4510 1794 4526 1858
rect 4590 1794 4732 1858
rect 4796 1794 4812 1858
rect 4876 1794 4892 1858
rect 4956 1794 4972 1858
rect 5036 1794 5052 1858
rect 5116 1794 5132 1858
rect 5196 1794 5338 1858
rect 5402 1794 5418 1858
rect 5482 1794 5498 1858
rect 5562 1794 5578 1858
rect 5642 1794 5658 1858
rect 5722 1794 5738 1858
rect 5802 1794 5944 1858
rect 6008 1794 6024 1858
rect 6088 1794 6104 1858
rect 6168 1794 6184 1858
rect 6248 1794 6264 1858
rect 6328 1794 6344 1858
rect 6408 1794 6512 1858
rect 1598 1792 6512 1794
rect 1598 1638 1664 1728
rect 1598 1574 1599 1638
rect 1663 1574 1664 1638
rect 1598 1558 1664 1574
rect 1598 1494 1599 1558
rect 1663 1494 1664 1558
rect 1598 1478 1664 1494
rect 1598 1414 1599 1478
rect 1663 1414 1664 1478
rect 1598 1398 1664 1414
rect 1598 1334 1599 1398
rect 1663 1334 1664 1398
rect 1598 1318 1664 1334
rect 1598 1254 1599 1318
rect 1663 1254 1664 1318
rect 1598 1238 1664 1254
rect 1598 1174 1599 1238
rect 1663 1174 1664 1238
rect 1598 1158 1664 1174
rect 1598 1094 1599 1158
rect 1663 1094 1664 1158
rect 1598 1078 1664 1094
rect 1598 1014 1599 1078
rect 1663 1014 1664 1078
rect 1598 998 1664 1014
rect 1598 934 1599 998
rect 1663 934 1664 998
rect 1598 918 1664 934
rect 1598 854 1599 918
rect 1663 854 1664 918
rect 1598 700 1664 854
rect 1724 700 1784 1732
rect 1844 762 1904 1792
rect 1964 700 2024 1732
rect 2084 762 2144 1792
rect 2204 1638 2270 1728
rect 2204 1574 2205 1638
rect 2269 1574 2270 1638
rect 2204 1558 2270 1574
rect 2204 1494 2205 1558
rect 2269 1494 2270 1558
rect 2204 1478 2270 1494
rect 2204 1414 2205 1478
rect 2269 1414 2270 1478
rect 2204 1398 2270 1414
rect 2204 1334 2205 1398
rect 2269 1334 2270 1398
rect 2204 1318 2270 1334
rect 2204 1254 2205 1318
rect 2269 1254 2270 1318
rect 2204 1238 2270 1254
rect 2204 1174 2205 1238
rect 2269 1174 2270 1238
rect 2204 1158 2270 1174
rect 2204 1094 2205 1158
rect 2269 1094 2270 1158
rect 2204 1078 2270 1094
rect 2204 1014 2205 1078
rect 2269 1014 2270 1078
rect 2204 998 2270 1014
rect 2204 934 2205 998
rect 2269 934 2270 998
rect 2204 918 2270 934
rect 2204 854 2205 918
rect 2269 854 2270 918
rect 2204 700 2270 854
rect 2330 700 2390 1732
rect 2450 762 2510 1792
rect 2570 700 2630 1732
rect 2690 762 2750 1792
rect 2810 1638 2876 1728
rect 2810 1574 2811 1638
rect 2875 1574 2876 1638
rect 2810 1558 2876 1574
rect 2810 1494 2811 1558
rect 2875 1494 2876 1558
rect 2810 1478 2876 1494
rect 2810 1414 2811 1478
rect 2875 1414 2876 1478
rect 2810 1398 2876 1414
rect 2810 1334 2811 1398
rect 2875 1334 2876 1398
rect 2810 1318 2876 1334
rect 2810 1254 2811 1318
rect 2875 1254 2876 1318
rect 2810 1238 2876 1254
rect 2810 1174 2811 1238
rect 2875 1174 2876 1238
rect 2810 1158 2876 1174
rect 2810 1094 2811 1158
rect 2875 1094 2876 1158
rect 2810 1078 2876 1094
rect 2810 1014 2811 1078
rect 2875 1014 2876 1078
rect 2810 998 2876 1014
rect 2810 934 2811 998
rect 2875 934 2876 998
rect 2810 918 2876 934
rect 2810 854 2811 918
rect 2875 854 2876 918
rect 2810 700 2876 854
rect 2936 700 2996 1732
rect 3056 762 3116 1792
rect 3176 700 3236 1732
rect 3296 762 3356 1792
rect 3416 1638 3482 1728
rect 3416 1574 3417 1638
rect 3481 1574 3482 1638
rect 3416 1558 3482 1574
rect 3416 1494 3417 1558
rect 3481 1494 3482 1558
rect 3416 1478 3482 1494
rect 3416 1414 3417 1478
rect 3481 1414 3482 1478
rect 3416 1398 3482 1414
rect 3416 1334 3417 1398
rect 3481 1334 3482 1398
rect 3416 1318 3482 1334
rect 3416 1254 3417 1318
rect 3481 1254 3482 1318
rect 3416 1238 3482 1254
rect 3416 1174 3417 1238
rect 3481 1174 3482 1238
rect 3416 1158 3482 1174
rect 3416 1094 3417 1158
rect 3481 1094 3482 1158
rect 3416 1078 3482 1094
rect 3416 1014 3417 1078
rect 3481 1014 3482 1078
rect 3416 998 3482 1014
rect 3416 934 3417 998
rect 3481 934 3482 998
rect 3416 918 3482 934
rect 3416 854 3417 918
rect 3481 854 3482 918
rect 3416 700 3482 854
rect 3542 700 3602 1732
rect 3662 762 3722 1792
rect 3782 700 3842 1732
rect 3902 762 3962 1792
rect 4022 1638 4088 1728
rect 4022 1574 4023 1638
rect 4087 1574 4088 1638
rect 4022 1558 4088 1574
rect 4022 1494 4023 1558
rect 4087 1494 4088 1558
rect 4022 1478 4088 1494
rect 4022 1414 4023 1478
rect 4087 1414 4088 1478
rect 4022 1398 4088 1414
rect 4022 1334 4023 1398
rect 4087 1334 4088 1398
rect 4022 1318 4088 1334
rect 4022 1254 4023 1318
rect 4087 1254 4088 1318
rect 4022 1238 4088 1254
rect 4022 1174 4023 1238
rect 4087 1174 4088 1238
rect 4022 1158 4088 1174
rect 4022 1094 4023 1158
rect 4087 1094 4088 1158
rect 4022 1078 4088 1094
rect 4022 1014 4023 1078
rect 4087 1014 4088 1078
rect 4022 998 4088 1014
rect 4022 934 4023 998
rect 4087 934 4088 998
rect 4022 918 4088 934
rect 4022 854 4023 918
rect 4087 854 4088 918
rect 4022 700 4088 854
rect 4148 700 4208 1732
rect 4268 762 4328 1792
rect 4388 700 4448 1732
rect 4508 762 4568 1792
rect 4628 1638 4694 1728
rect 4628 1574 4629 1638
rect 4693 1574 4694 1638
rect 4628 1558 4694 1574
rect 4628 1494 4629 1558
rect 4693 1494 4694 1558
rect 4628 1478 4694 1494
rect 4628 1414 4629 1478
rect 4693 1414 4694 1478
rect 4628 1398 4694 1414
rect 4628 1334 4629 1398
rect 4693 1334 4694 1398
rect 4628 1318 4694 1334
rect 4628 1254 4629 1318
rect 4693 1254 4694 1318
rect 4628 1238 4694 1254
rect 4628 1174 4629 1238
rect 4693 1174 4694 1238
rect 4628 1158 4694 1174
rect 4628 1094 4629 1158
rect 4693 1094 4694 1158
rect 4628 1078 4694 1094
rect 4628 1014 4629 1078
rect 4693 1014 4694 1078
rect 4628 998 4694 1014
rect 4628 934 4629 998
rect 4693 934 4694 998
rect 4628 918 4694 934
rect 4628 854 4629 918
rect 4693 854 4694 918
rect 4628 700 4694 854
rect 4754 700 4814 1732
rect 4874 762 4934 1792
rect 4994 700 5054 1732
rect 5114 762 5174 1792
rect 5234 1638 5300 1728
rect 5234 1574 5235 1638
rect 5299 1574 5300 1638
rect 5234 1558 5300 1574
rect 5234 1494 5235 1558
rect 5299 1494 5300 1558
rect 5234 1478 5300 1494
rect 5234 1414 5235 1478
rect 5299 1414 5300 1478
rect 5234 1398 5300 1414
rect 5234 1334 5235 1398
rect 5299 1334 5300 1398
rect 5234 1318 5300 1334
rect 5234 1254 5235 1318
rect 5299 1254 5300 1318
rect 5234 1238 5300 1254
rect 5234 1174 5235 1238
rect 5299 1174 5300 1238
rect 5234 1158 5300 1174
rect 5234 1094 5235 1158
rect 5299 1094 5300 1158
rect 5234 1078 5300 1094
rect 5234 1014 5235 1078
rect 5299 1014 5300 1078
rect 5234 998 5300 1014
rect 5234 934 5235 998
rect 5299 934 5300 998
rect 5234 918 5300 934
rect 5234 854 5235 918
rect 5299 854 5300 918
rect 5234 700 5300 854
rect 5360 700 5420 1732
rect 5480 762 5540 1792
rect 5600 700 5660 1732
rect 5720 762 5780 1792
rect 5840 1638 5906 1728
rect 5840 1574 5841 1638
rect 5905 1574 5906 1638
rect 5840 1558 5906 1574
rect 5840 1494 5841 1558
rect 5905 1494 5906 1558
rect 5840 1478 5906 1494
rect 5840 1414 5841 1478
rect 5905 1414 5906 1478
rect 5840 1398 5906 1414
rect 5840 1334 5841 1398
rect 5905 1334 5906 1398
rect 5840 1318 5906 1334
rect 5840 1254 5841 1318
rect 5905 1254 5906 1318
rect 5840 1238 5906 1254
rect 5840 1174 5841 1238
rect 5905 1174 5906 1238
rect 5840 1158 5906 1174
rect 5840 1094 5841 1158
rect 5905 1094 5906 1158
rect 5840 1078 5906 1094
rect 5840 1014 5841 1078
rect 5905 1014 5906 1078
rect 5840 998 5906 1014
rect 5840 934 5841 998
rect 5905 934 5906 998
rect 5840 918 5906 934
rect 5840 854 5841 918
rect 5905 854 5906 918
rect 5840 700 5906 854
rect 5966 700 6026 1732
rect 6086 762 6146 1792
rect 6206 700 6266 1732
rect 6326 762 6386 1792
rect 6446 1638 6512 1728
rect 6446 1574 6447 1638
rect 6511 1574 6512 1638
rect 6446 1558 6512 1574
rect 6446 1494 6447 1558
rect 6511 1494 6512 1558
rect 6446 1478 6512 1494
rect 6446 1414 6447 1478
rect 6511 1414 6512 1478
rect 6446 1398 6512 1414
rect 6446 1334 6447 1398
rect 6511 1334 6512 1398
rect 6446 1318 6512 1334
rect 6446 1254 6447 1318
rect 6511 1254 6512 1318
rect 6446 1238 6512 1254
rect 6446 1174 6447 1238
rect 6511 1174 6512 1238
rect 6446 1158 6512 1174
rect 6446 1094 6447 1158
rect 6511 1094 6512 1158
rect 6446 1078 6512 1094
rect 6446 1014 6447 1078
rect 6511 1014 6512 1078
rect 6446 998 6512 1014
rect 6446 934 6447 998
rect 6511 934 6512 998
rect 6446 918 6512 934
rect 6446 854 6447 918
rect 6511 854 6512 918
rect 6446 700 6512 854
rect 1598 698 6512 700
rect 1598 634 1702 698
rect 1766 634 1782 698
rect 1846 634 1862 698
rect 1926 634 1942 698
rect 2006 634 2022 698
rect 2086 634 2102 698
rect 2166 634 2308 698
rect 2372 634 2388 698
rect 2452 634 2468 698
rect 2532 634 2548 698
rect 2612 634 2628 698
rect 2692 634 2708 698
rect 2772 634 2914 698
rect 2978 634 2994 698
rect 3058 634 3074 698
rect 3138 634 3154 698
rect 3218 634 3234 698
rect 3298 634 3314 698
rect 3378 634 3520 698
rect 3584 634 3600 698
rect 3664 634 3680 698
rect 3744 634 3760 698
rect 3824 634 3840 698
rect 3904 634 3920 698
rect 3984 634 4126 698
rect 4190 634 4206 698
rect 4270 634 4286 698
rect 4350 634 4366 698
rect 4430 634 4446 698
rect 4510 634 4526 698
rect 4590 634 4732 698
rect 4796 634 4812 698
rect 4876 634 4892 698
rect 4956 634 4972 698
rect 5036 634 5052 698
rect 5116 634 5132 698
rect 5196 634 5338 698
rect 5402 634 5418 698
rect 5482 634 5498 698
rect 5562 634 5578 698
rect 5642 634 5658 698
rect 5722 634 5738 698
rect 5802 634 5944 698
rect 6008 634 6024 698
rect 6088 634 6104 698
rect 6168 634 6184 698
rect 6248 634 6264 698
rect 6328 634 6344 698
rect 6408 634 6512 698
rect 1598 632 6512 634
rect 1598 478 1664 632
rect 1598 414 1599 478
rect 1663 414 1664 478
rect 1598 398 1664 414
rect 1598 334 1599 398
rect 1663 334 1664 398
rect 1598 318 1664 334
rect 1598 254 1599 318
rect 1663 254 1664 318
rect 1598 238 1664 254
rect 1598 174 1599 238
rect 1663 174 1664 238
rect 1598 158 1664 174
rect 1598 94 1599 158
rect 1663 94 1664 158
rect 1598 78 1664 94
rect 1598 14 1599 78
rect 1663 14 1664 78
rect 1598 -2 1664 14
rect 1598 -66 1599 -2
rect 1663 -66 1664 -2
rect 1598 -82 1664 -66
rect 1598 -146 1599 -82
rect 1663 -146 1664 -82
rect 1598 -162 1664 -146
rect 1598 -226 1599 -162
rect 1663 -226 1664 -162
rect 1598 -242 1664 -226
rect 1598 -306 1599 -242
rect 1663 -306 1664 -242
rect 1598 -396 1664 -306
rect 1724 -460 1784 570
rect 1844 -400 1904 632
rect 1964 -460 2024 570
rect 2084 -400 2144 632
rect 2204 478 2270 632
rect 2204 414 2205 478
rect 2269 414 2270 478
rect 2204 398 2270 414
rect 2204 334 2205 398
rect 2269 334 2270 398
rect 2204 318 2270 334
rect 2204 254 2205 318
rect 2269 254 2270 318
rect 2204 238 2270 254
rect 2204 174 2205 238
rect 2269 174 2270 238
rect 2204 158 2270 174
rect 2204 94 2205 158
rect 2269 94 2270 158
rect 2204 78 2270 94
rect 2204 14 2205 78
rect 2269 14 2270 78
rect 2204 -2 2270 14
rect 2204 -66 2205 -2
rect 2269 -66 2270 -2
rect 2204 -82 2270 -66
rect 2204 -146 2205 -82
rect 2269 -146 2270 -82
rect 2204 -162 2270 -146
rect 2204 -226 2205 -162
rect 2269 -226 2270 -162
rect 2204 -242 2270 -226
rect 2204 -306 2205 -242
rect 2269 -306 2270 -242
rect 2204 -396 2270 -306
rect 2330 -460 2390 570
rect 2450 -400 2510 632
rect 2570 -460 2630 570
rect 2690 -400 2750 632
rect 2810 478 2876 632
rect 2810 414 2811 478
rect 2875 414 2876 478
rect 2810 398 2876 414
rect 2810 334 2811 398
rect 2875 334 2876 398
rect 2810 318 2876 334
rect 2810 254 2811 318
rect 2875 254 2876 318
rect 2810 238 2876 254
rect 2810 174 2811 238
rect 2875 174 2876 238
rect 2810 158 2876 174
rect 2810 94 2811 158
rect 2875 94 2876 158
rect 2810 78 2876 94
rect 2810 14 2811 78
rect 2875 14 2876 78
rect 2810 -2 2876 14
rect 2810 -66 2811 -2
rect 2875 -66 2876 -2
rect 2810 -82 2876 -66
rect 2810 -146 2811 -82
rect 2875 -146 2876 -82
rect 2810 -162 2876 -146
rect 2810 -226 2811 -162
rect 2875 -226 2876 -162
rect 2810 -242 2876 -226
rect 2810 -306 2811 -242
rect 2875 -306 2876 -242
rect 2810 -396 2876 -306
rect 2936 -460 2996 570
rect 3056 -400 3116 632
rect 3176 -460 3236 570
rect 3296 -400 3356 632
rect 3416 478 3482 632
rect 3416 414 3417 478
rect 3481 414 3482 478
rect 3416 398 3482 414
rect 3416 334 3417 398
rect 3481 334 3482 398
rect 3416 318 3482 334
rect 3416 254 3417 318
rect 3481 254 3482 318
rect 3416 238 3482 254
rect 3416 174 3417 238
rect 3481 174 3482 238
rect 3416 158 3482 174
rect 3416 94 3417 158
rect 3481 94 3482 158
rect 3416 78 3482 94
rect 3416 14 3417 78
rect 3481 14 3482 78
rect 3416 -2 3482 14
rect 3416 -66 3417 -2
rect 3481 -66 3482 -2
rect 3416 -82 3482 -66
rect 3416 -146 3417 -82
rect 3481 -146 3482 -82
rect 3416 -162 3482 -146
rect 3416 -226 3417 -162
rect 3481 -226 3482 -162
rect 3416 -242 3482 -226
rect 3416 -306 3417 -242
rect 3481 -306 3482 -242
rect 3416 -396 3482 -306
rect 3542 -460 3602 570
rect 3662 -400 3722 632
rect 3782 -460 3842 570
rect 3902 -400 3962 632
rect 4022 478 4088 632
rect 4022 414 4023 478
rect 4087 414 4088 478
rect 4022 398 4088 414
rect 4022 334 4023 398
rect 4087 334 4088 398
rect 4022 318 4088 334
rect 4022 254 4023 318
rect 4087 254 4088 318
rect 4022 238 4088 254
rect 4022 174 4023 238
rect 4087 174 4088 238
rect 4022 158 4088 174
rect 4022 94 4023 158
rect 4087 94 4088 158
rect 4022 78 4088 94
rect 4022 14 4023 78
rect 4087 14 4088 78
rect 4022 -2 4088 14
rect 4022 -66 4023 -2
rect 4087 -66 4088 -2
rect 4022 -82 4088 -66
rect 4022 -146 4023 -82
rect 4087 -146 4088 -82
rect 4022 -162 4088 -146
rect 4022 -226 4023 -162
rect 4087 -226 4088 -162
rect 4022 -242 4088 -226
rect 4022 -306 4023 -242
rect 4087 -306 4088 -242
rect 4022 -396 4088 -306
rect 4148 -460 4208 570
rect 4268 -400 4328 632
rect 4388 -460 4448 570
rect 4508 -400 4568 632
rect 4628 478 4694 632
rect 4628 414 4629 478
rect 4693 414 4694 478
rect 4628 398 4694 414
rect 4628 334 4629 398
rect 4693 334 4694 398
rect 4628 318 4694 334
rect 4628 254 4629 318
rect 4693 254 4694 318
rect 4628 238 4694 254
rect 4628 174 4629 238
rect 4693 174 4694 238
rect 4628 158 4694 174
rect 4628 94 4629 158
rect 4693 94 4694 158
rect 4628 78 4694 94
rect 4628 14 4629 78
rect 4693 14 4694 78
rect 4628 -2 4694 14
rect 4628 -66 4629 -2
rect 4693 -66 4694 -2
rect 4628 -82 4694 -66
rect 4628 -146 4629 -82
rect 4693 -146 4694 -82
rect 4628 -162 4694 -146
rect 4628 -226 4629 -162
rect 4693 -226 4694 -162
rect 4628 -242 4694 -226
rect 4628 -306 4629 -242
rect 4693 -306 4694 -242
rect 4628 -396 4694 -306
rect 4754 -460 4814 570
rect 4874 -400 4934 632
rect 4994 -460 5054 570
rect 5114 -400 5174 632
rect 5234 478 5300 632
rect 5234 414 5235 478
rect 5299 414 5300 478
rect 5234 398 5300 414
rect 5234 334 5235 398
rect 5299 334 5300 398
rect 5234 318 5300 334
rect 5234 254 5235 318
rect 5299 254 5300 318
rect 5234 238 5300 254
rect 5234 174 5235 238
rect 5299 174 5300 238
rect 5234 158 5300 174
rect 5234 94 5235 158
rect 5299 94 5300 158
rect 5234 78 5300 94
rect 5234 14 5235 78
rect 5299 14 5300 78
rect 5234 -2 5300 14
rect 5234 -66 5235 -2
rect 5299 -66 5300 -2
rect 5234 -82 5300 -66
rect 5234 -146 5235 -82
rect 5299 -146 5300 -82
rect 5234 -162 5300 -146
rect 5234 -226 5235 -162
rect 5299 -226 5300 -162
rect 5234 -242 5300 -226
rect 5234 -306 5235 -242
rect 5299 -306 5300 -242
rect 5234 -396 5300 -306
rect 5360 -460 5420 570
rect 5480 -400 5540 632
rect 5600 -460 5660 570
rect 5720 -400 5780 632
rect 5840 478 5906 632
rect 5840 414 5841 478
rect 5905 414 5906 478
rect 5840 398 5906 414
rect 5840 334 5841 398
rect 5905 334 5906 398
rect 5840 318 5906 334
rect 5840 254 5841 318
rect 5905 254 5906 318
rect 5840 238 5906 254
rect 5840 174 5841 238
rect 5905 174 5906 238
rect 5840 158 5906 174
rect 5840 94 5841 158
rect 5905 94 5906 158
rect 5840 78 5906 94
rect 5840 14 5841 78
rect 5905 14 5906 78
rect 5840 -2 5906 14
rect 5840 -66 5841 -2
rect 5905 -66 5906 -2
rect 5840 -82 5906 -66
rect 5840 -146 5841 -82
rect 5905 -146 5906 -82
rect 5840 -162 5906 -146
rect 5840 -226 5841 -162
rect 5905 -226 5906 -162
rect 5840 -242 5906 -226
rect 5840 -306 5841 -242
rect 5905 -306 5906 -242
rect 5840 -396 5906 -306
rect 5966 -460 6026 570
rect 6086 -400 6146 632
rect 6206 -460 6266 570
rect 6326 -400 6386 632
rect 6446 478 6512 632
rect 6446 414 6447 478
rect 6511 414 6512 478
rect 6446 398 6512 414
rect 6446 334 6447 398
rect 6511 334 6512 398
rect 6446 318 6512 334
rect 6446 254 6447 318
rect 6511 254 6512 318
rect 6446 238 6512 254
rect 6446 174 6447 238
rect 6511 174 6512 238
rect 6446 158 6512 174
rect 6446 94 6447 158
rect 6511 94 6512 158
rect 6446 78 6512 94
rect 6446 14 6447 78
rect 6511 14 6512 78
rect 6446 -2 6512 14
rect 6446 -66 6447 -2
rect 6511 -66 6512 -2
rect 6446 -82 6512 -66
rect 6446 -146 6447 -82
rect 6511 -146 6512 -82
rect 6446 -162 6512 -146
rect 6446 -226 6447 -162
rect 6511 -226 6512 -162
rect 6446 -242 6512 -226
rect 6446 -306 6447 -242
rect 6511 -306 6512 -242
rect 6446 -396 6512 -306
rect 1598 -462 6512 -460
rect 1598 -526 1702 -462
rect 1766 -526 1782 -462
rect 1846 -526 1862 -462
rect 1926 -526 1942 -462
rect 2006 -526 2022 -462
rect 2086 -526 2102 -462
rect 2166 -526 2308 -462
rect 2372 -526 2388 -462
rect 2452 -526 2468 -462
rect 2532 -526 2548 -462
rect 2612 -526 2628 -462
rect 2692 -526 2708 -462
rect 2772 -526 2914 -462
rect 2978 -526 2994 -462
rect 3058 -526 3074 -462
rect 3138 -526 3154 -462
rect 3218 -526 3234 -462
rect 3298 -526 3314 -462
rect 3378 -526 3520 -462
rect 3584 -526 3600 -462
rect 3664 -526 3680 -462
rect 3744 -526 3760 -462
rect 3824 -526 3840 -462
rect 3904 -526 3920 -462
rect 3984 -526 4126 -462
rect 4190 -526 4206 -462
rect 4270 -526 4286 -462
rect 4350 -526 4366 -462
rect 4430 -526 4446 -462
rect 4510 -526 4526 -462
rect 4590 -526 4732 -462
rect 4796 -526 4812 -462
rect 4876 -526 4892 -462
rect 4956 -526 4972 -462
rect 5036 -526 5052 -462
rect 5116 -526 5132 -462
rect 5196 -526 5338 -462
rect 5402 -526 5418 -462
rect 5482 -526 5498 -462
rect 5562 -526 5578 -462
rect 5642 -526 5658 -462
rect 5722 -526 5738 -462
rect 5802 -526 5944 -462
rect 6008 -526 6024 -462
rect 6088 -526 6104 -462
rect 6168 -526 6184 -462
rect 6248 -526 6264 -462
rect 6328 -526 6344 -462
rect 6408 -526 6512 -462
rect 1598 -528 6512 -526
<< labels >>
flabel metal4 4402 770 4438 850 0 FreeSans 320 0 0 0 CBOT
port 2 nsew
flabel metal4 3678 800 3714 880 0 FreeSans 320 0 0 0 CTOP
port 4 nsew
flabel metal4 3792 426 3836 508 0 FreeSans 320 0 0 0 CTOP
port 8 nsew
flabel psubdiff 4096 526 4140 608 0 FreeSans 320 0 0 0 SUB
port 10 nsew
flabel pwell 2530 1412 2556 1444 0 FreeSans 160 0 0 0 x1[3].SUB
flabel metal4 2588 1078 2614 1110 0 FreeSans 320 0 0 0 x1[3].CBOT
flabel metal4 2470 1668 2496 1700 0 FreeSans 320 0 0 0 x1[3].CTOP
flabel pwell 1924 1412 1950 1444 0 FreeSans 160 0 0 0 x1[1].SUB
flabel metal4 1982 1078 2008 1110 0 FreeSans 320 0 0 0 x1[1].CBOT
flabel metal4 1864 1668 1890 1700 0 FreeSans 320 0 0 0 x1[1].CTOP
flabel pwell 4348 1412 4374 1444 0 FreeSans 160 0 0 0 x1[9].SUB
flabel metal4 4406 1078 4432 1110 0 FreeSans 320 0 0 0 x1[9].CBOT
flabel metal4 4288 1668 4314 1700 0 FreeSans 320 0 0 0 x1[9].CTOP
flabel pwell 3742 1412 3768 1444 0 FreeSans 160 0 0 0 x1[7].SUB
flabel metal4 3800 1078 3826 1110 0 FreeSans 320 0 0 0 x1[7].CBOT
flabel metal4 3682 1668 3708 1700 0 FreeSans 320 0 0 0 x1[7].CTOP
flabel pwell 3136 1412 3162 1444 0 FreeSans 160 0 0 0 x1[5].SUB
flabel metal4 3194 1078 3220 1110 0 FreeSans 320 0 0 0 x1[5].CBOT
flabel metal4 3076 1668 3102 1700 0 FreeSans 320 0 0 0 x1[5].CTOP
flabel pwell 5560 1412 5586 1444 0 FreeSans 160 0 0 0 x1[13].SUB
flabel metal4 5618 1078 5644 1110 0 FreeSans 320 0 0 0 x1[13].CBOT
flabel metal4 5500 1668 5526 1700 0 FreeSans 320 0 0 0 x1[13].CTOP
flabel pwell 4954 1412 4980 1444 0 FreeSans 160 0 0 0 x1[11].SUB
flabel metal4 5012 1078 5038 1110 0 FreeSans 320 0 0 0 x1[11].CBOT
flabel metal4 4894 1668 4920 1700 0 FreeSans 320 0 0 0 x1[11].CTOP
flabel pwell 6166 1412 6192 1444 0 FreeSans 160 0 0 0 x1[15].SUB
flabel metal4 6224 1078 6250 1110 0 FreeSans 320 0 0 0 x1[15].CBOT
flabel metal4 6106 1668 6132 1700 0 FreeSans 320 0 0 0 x1[15].CTOP
flabel pwell 6160 -112 6186 -80 0 FreeSans 160 0 0 0 x1[14].SUB
flabel metal4 6102 222 6128 254 0 FreeSans 320 0 0 0 x1[14].CBOT
flabel metal4 6220 -368 6246 -336 0 FreeSans 320 0 0 0 x1[14].CTOP
flabel pwell 5554 -112 5580 -80 0 FreeSans 160 0 0 0 x1[12].SUB
flabel metal4 5496 222 5522 254 0 FreeSans 320 0 0 0 x1[12].CBOT
flabel metal4 5614 -368 5640 -336 0 FreeSans 320 0 0 0 x1[12].CTOP
flabel pwell 4948 -112 4974 -80 0 FreeSans 160 0 0 0 x1[10].SUB
flabel metal4 4890 222 4916 254 0 FreeSans 320 0 0 0 x1[10].CBOT
flabel metal4 5008 -368 5034 -336 0 FreeSans 320 0 0 0 x1[10].CTOP
flabel pwell 4342 -112 4368 -80 0 FreeSans 160 0 0 0 x1[8].SUB
flabel metal4 4284 222 4310 254 0 FreeSans 320 0 0 0 x1[8].CBOT
flabel metal4 4402 -368 4428 -336 0 FreeSans 320 0 0 0 x1[8].CTOP
flabel pwell 3736 -112 3762 -80 0 FreeSans 160 0 0 0 x1[6].SUB
flabel metal4 3678 222 3704 254 0 FreeSans 320 0 0 0 x1[6].CBOT
flabel metal4 3796 -368 3822 -336 0 FreeSans 320 0 0 0 x1[6].CTOP
flabel pwell 3130 -112 3156 -80 0 FreeSans 160 0 0 0 x1[4].SUB
flabel metal4 3072 222 3098 254 0 FreeSans 320 0 0 0 x1[4].CBOT
flabel metal4 3190 -368 3216 -336 0 FreeSans 320 0 0 0 x1[4].CTOP
flabel pwell 2524 -112 2550 -80 0 FreeSans 160 0 0 0 x1[2].SUB
flabel metal4 2466 222 2492 254 0 FreeSans 320 0 0 0 x1[2].CBOT
flabel metal4 2584 -368 2610 -336 0 FreeSans 320 0 0 0 x1[2].CTOP
flabel pwell 1918 -112 1944 -80 0 FreeSans 160 0 0 0 x1[0].SUB
flabel metal4 1860 222 1886 254 0 FreeSans 320 0 0 0 x1[0].CBOT
flabel metal4 1978 -368 2004 -336 0 FreeSans 320 0 0 0 x1[0].CTOP
<< end >>
