* NGSPICE file created from hgu_cdac_cap_2.ext - technology: sky130A

.subckt hgu_cdac_cap_2 SUB
C0 x1.CBOT x2.CTOP 5.11f
C1 x2.CTOP x2.CBOT 5.11f
C2 x1.CBOT SUB 1.38f $ **FLOATING
C3 x2.CBOT SUB 1.38f $ **FLOATING
.ends

