* NGSPICE file created from hgu_cdac_cap_2.ext - technology: sky130A

.subckt hgu_cdac_cap_2 SUB CBOT CTOP
C0 CTOP CBOT 10.2f
C1 CTOP SUB 1.1f
C2 CBOT SUB 2.17f
.ends

