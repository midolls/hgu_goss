magic
tech sky130A
magscale 1 2
timestamp 1697718446
<< nwell >>
rect 1419 162 4041 469
rect 1987 156 2086 162
rect 3434 160 3704 162
<< pdiff >>
rect 3549 338 3595 339
rect 3549 281 3555 338
rect 3589 281 3595 338
rect 3948 316 3987 339
<< ndiffc >>
rect 3467 0 3501 34
rect 3555 0 3589 34
rect 3643 0 3677 34
rect 1468 -46 1502 -12
rect 3354 -41 3388 -7
<< pdiffc >>
rect 1468 200 1502 234
rect 1925 194 1959 228
rect 3467 224 3501 337
rect 3555 224 3589 338
rect 3643 224 3677 337
<< poly >>
rect 1513 127 1912 157
rect 3513 155 3631 172
rect 1749 116 1815 127
rect 1749 82 1765 116
rect 1799 82 1815 116
rect 1749 63 1815 82
rect 3513 121 3541 155
rect 3575 121 3631 155
rect 3513 75 3631 121
rect 1513 33 3343 63
<< polycont >>
rect 1765 82 1799 116
rect 3541 121 3575 155
<< locali >>
rect 1444 401 1468 435
rect 1502 401 1540 435
rect 1574 401 1612 435
rect 1646 401 1684 435
rect 1718 401 1756 435
rect 1790 401 1828 435
rect 1862 401 1900 435
rect 1934 401 1972 435
rect 2006 401 3412 435
rect 3446 401 3484 435
rect 3518 401 3556 435
rect 3590 401 3628 435
rect 3662 401 3700 435
rect 3734 401 3772 435
rect 3806 401 3844 435
rect 3878 401 3916 435
rect 3950 401 3988 435
rect 4022 401 4060 435
rect 4094 401 4104 435
rect 1468 234 1502 401
rect 1468 172 1502 200
rect 1925 228 1959 401
rect 3467 337 3501 401
rect 3467 202 3501 224
rect 3555 338 3589 363
rect 3555 201 3589 224
rect 3643 337 3677 362
rect 1925 155 1959 194
rect 3643 155 3677 224
rect 1749 116 1815 132
rect 1924 121 2402 155
rect 2809 121 3541 155
rect 3575 121 3597 155
rect 3643 121 4104 155
rect 1455 82 1765 116
rect 1799 82 1815 116
rect 1455 81 1815 82
rect 1749 66 1815 81
rect 1468 -12 1502 18
rect 1468 -100 1502 -46
rect 3354 -7 3388 121
rect 3354 -66 3388 -41
rect 3467 34 3501 60
rect 3467 -100 3501 0
rect 3555 34 3589 60
rect 3555 -24 3589 0
rect 3643 34 3677 121
rect 3643 -24 3677 0
rect 1433 -134 1468 -100
rect 1502 -134 1540 -100
rect 1574 -134 1612 -100
rect 1646 -134 1684 -100
rect 1718 -134 1756 -100
rect 1790 -134 1828 -100
rect 1862 -134 1900 -100
rect 1934 -134 1972 -100
rect 2006 -134 2044 -100
rect 2078 -134 2116 -100
rect 2150 -134 2188 -100
rect 2222 -134 2260 -100
rect 2294 -134 2332 -100
rect 2366 -134 2404 -100
rect 2438 -134 2476 -100
rect 2510 -134 2548 -100
rect 2582 -134 2620 -100
rect 2654 -134 2692 -100
rect 2726 -134 2764 -100
rect 2798 -134 2836 -100
rect 2870 -134 2908 -100
rect 2942 -134 2980 -100
rect 3014 -134 3052 -100
rect 3086 -134 3124 -100
rect 3158 -134 3196 -100
rect 3230 -134 3268 -100
rect 3302 -134 3340 -100
rect 3374 -134 3412 -100
rect 3446 -134 3484 -100
rect 3518 -134 3556 -100
rect 3590 -134 3628 -100
rect 3662 -134 3700 -100
rect 3734 -134 3772 -100
rect 3806 -134 3844 -100
rect 3878 -134 3916 -100
rect 3950 -134 3988 -100
rect 4022 -134 4060 -100
rect 4094 -134 4104 -100
<< viali >>
rect 1468 401 1502 435
rect 1540 401 1574 435
rect 1612 401 1646 435
rect 1684 401 1718 435
rect 1756 401 1790 435
rect 1828 401 1862 435
rect 1900 401 1934 435
rect 1972 401 2006 435
rect 3412 401 3446 435
rect 3484 401 3518 435
rect 3556 401 3590 435
rect 3628 401 3662 435
rect 3700 401 3734 435
rect 3772 401 3806 435
rect 3844 401 3878 435
rect 3916 401 3950 435
rect 3988 401 4022 435
rect 4060 401 4094 435
rect 3555 293 3589 327
rect 3555 0 3589 34
rect 1468 -134 1502 -100
rect 1540 -134 1574 -100
rect 1612 -134 1646 -100
rect 1684 -134 1718 -100
rect 1756 -134 1790 -100
rect 1828 -134 1862 -100
rect 1900 -134 1934 -100
rect 1972 -134 2006 -100
rect 2044 -134 2078 -100
rect 2116 -134 2150 -100
rect 2188 -134 2222 -100
rect 2260 -134 2294 -100
rect 2332 -134 2366 -100
rect 2404 -134 2438 -100
rect 2476 -134 2510 -100
rect 2548 -134 2582 -100
rect 2620 -134 2654 -100
rect 2692 -134 2726 -100
rect 2764 -134 2798 -100
rect 2836 -134 2870 -100
rect 2908 -134 2942 -100
rect 2980 -134 3014 -100
rect 3052 -134 3086 -100
rect 3124 -134 3158 -100
rect 3196 -134 3230 -100
rect 3268 -134 3302 -100
rect 3340 -134 3374 -100
rect 3412 -134 3446 -100
rect 3484 -134 3518 -100
rect 3556 -134 3590 -100
rect 3628 -134 3662 -100
rect 3700 -134 3734 -100
rect 3772 -134 3806 -100
rect 3844 -134 3878 -100
rect 3916 -134 3950 -100
rect 3988 -134 4022 -100
rect 4060 -134 4094 -100
<< metal1 >>
rect 1444 435 4104 469
rect 1444 401 1468 435
rect 1502 401 1540 435
rect 1574 401 1612 435
rect 1646 401 1684 435
rect 1718 401 1756 435
rect 1790 401 1828 435
rect 1862 401 1900 435
rect 1934 401 1972 435
rect 2006 401 3412 435
rect 3446 401 3484 435
rect 3518 401 3556 435
rect 3590 401 3628 435
rect 3662 401 3700 435
rect 3734 401 3772 435
rect 3806 401 3844 435
rect 3878 401 3916 435
rect 3950 401 3988 435
rect 4022 401 4060 435
rect 4094 401 4104 435
rect 1444 367 4104 401
rect 3549 327 3987 339
rect 3549 293 3555 327
rect 3589 316 3987 327
rect 3589 307 3980 316
rect 3589 293 3595 307
rect 3549 281 3595 293
rect 3852 174 3885 208
rect 3489 141 3885 174
rect 3489 -66 3521 141
rect 4015 113 4047 367
rect 3845 81 4047 113
rect 3845 75 3891 81
rect 3549 34 3596 60
rect 3549 0 3555 34
rect 3589 0 3596 34
rect 3549 -5 3596 0
rect 3941 -5 3987 1
rect 3549 -38 3987 -5
rect 1433 -100 4104 -66
rect 1433 -134 1468 -100
rect 1502 -134 1540 -100
rect 1574 -134 1612 -100
rect 1646 -134 1684 -100
rect 1718 -134 1756 -100
rect 1790 -134 1828 -100
rect 1862 -134 1900 -100
rect 1934 -134 1972 -100
rect 2006 -134 2044 -100
rect 2078 -134 2116 -100
rect 2150 -134 2188 -100
rect 2222 -134 2260 -100
rect 2294 -134 2332 -100
rect 2366 -134 2404 -100
rect 2438 -134 2476 -100
rect 2510 -134 2548 -100
rect 2582 -134 2620 -100
rect 2654 -134 2692 -100
rect 2726 -134 2764 -100
rect 2798 -134 2836 -100
rect 2870 -134 2908 -100
rect 2942 -134 2980 -100
rect 3014 -134 3052 -100
rect 3086 -134 3124 -100
rect 3158 -134 3196 -100
rect 3230 -134 3268 -100
rect 3302 -134 3340 -100
rect 3374 -134 3412 -100
rect 3446 -134 3484 -100
rect 3518 -134 3556 -100
rect 3590 -134 3628 -100
rect 3662 -134 3700 -100
rect 3734 -134 3772 -100
rect 3806 -134 3844 -100
rect 3878 -134 3916 -100
rect 3950 -134 3988 -100
rect 4022 -134 4060 -100
rect 4094 -134 4104 -100
rect 1433 -168 4104 -134
use sky130_fd_pr__nfet_01v8_MVW3GX  XM1
timestamp 1697717772
transform 1 0 3868 0 -1 41
box -125 -130 125 68
use sky130_fd_pr__pfet_01v8_XYYHBL  XM2
timestamp 1697716041
transform 1 0 3868 0 1 282
box -162 -177 162 118
use sky130_fd_pr__pfet_01v8_NSZ2Q7  XM3
timestamp 1697716041
transform 1 0 2710 0 1 261
box -727 -156 725 156
use sky130_fd_pr__nfet_01v8_L7T3GD  XM4
timestamp 1697704885
transform -1 0 3328 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__pfet_01v8_M479BZ  XM5
timestamp 1697713470
transform -1 0 1897 0 1 214
box -109 -83 109 90
use sky130_fd_pr__nfet_01v8_L7T3GD  XM6
timestamp 1697704885
transform -1 0 3256 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__pfet_01v8_M479BZ  XM7
timestamp 1697713470
transform -1 0 1825 0 1 214
box -109 -83 109 90
use sky130_fd_pr__pfet_01v8_M479BZ  XM8
timestamp 1697713470
transform -1 0 1744 0 1 214
box -109 -83 109 90
use sky130_fd_pr__pfet_01v8_M479BZ  XM9
timestamp 1697713470
transform -1 0 1672 0 1 214
box -109 -83 109 90
use sky130_fd_pr__pfet_01v8_M479BZ  XM10
timestamp 1697713470
transform -1 0 1600 0 1 214
box -109 -83 109 90
use sky130_fd_pr__pfet_01v8_M479BZ  XM11
timestamp 1697713470
transform -1 0 1528 0 1 214
box -109 -83 109 90
use sky130_fd_pr__nfet_01v8_L7T3GD  XM12
timestamp 1697704885
transform -1 0 1888 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM13
timestamp 1697704885
transform 1 0 3616 0 1 18
box -73 -69 73 68
use sky130_fd_pr__pfet_01v8_XYUFBL  XM14
timestamp 1697713470
transform 1 0 3528 0 1 282
box -109 -127 110 116
use sky130_fd_pr__nfet_01v8_L7T3GD  XM15
timestamp 1697704885
transform 1 0 3528 0 1 18
box -73 -69 73 68
use sky130_fd_pr__pfet_01v8_XYUFBL  XM16
timestamp 1697713470
transform 1 0 3616 0 1 282
box -109 -127 110 116
use sky130_fd_pr__nfet_01v8_L7T3GD  XM17
timestamp 1697704885
transform -1 0 2608 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM18
timestamp 1697704885
transform -1 0 2536 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM19
timestamp 1697704885
transform -1 0 2464 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM20
timestamp 1697704885
transform -1 0 2392 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM21
timestamp 1697704885
transform -1 0 3184 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM22
timestamp 1697704885
transform -1 0 3112 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM23
timestamp 1697704885
transform -1 0 3040 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM24
timestamp 1697704885
transform -1 0 2968 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM25
timestamp 1697704885
transform -1 0 2896 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM26
timestamp 1697704885
transform -1 0 2824 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM27
timestamp 1697704885
transform -1 0 2752 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM28
timestamp 1697704885
transform -1 0 2680 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM29
timestamp 1697704885
transform -1 0 2320 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM30
timestamp 1697704885
transform -1 0 2248 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM31
timestamp 1697704885
transform -1 0 2176 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM32
timestamp 1697704885
transform -1 0 2104 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM33
timestamp 1697704885
transform -1 0 2032 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM34
timestamp 1697704885
transform -1 0 1960 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM36
timestamp 1697704885
transform -1 0 1816 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM37
timestamp 1697704885
transform -1 0 1744 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM38
timestamp 1697704885
transform -1 0 1672 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM39
timestamp 1697704885
transform -1 0 1600 0 1 -24
box -73 -69 73 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM40
timestamp 1697704885
transform -1 0 1528 0 1 -24
box -73 -69 73 68
<< end >>
