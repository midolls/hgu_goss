magic
tech sky130A
magscale 1 2
timestamp 1697441537
<< error_s >>
rect 476 -710 6752 -674
rect 476 -852 512 -710
rect 1634 -778 2656 -776
rect 1232 -812 2656 -778
rect 1232 -814 1670 -812
rect 1232 -852 1268 -814
rect 2620 -852 2656 -812
rect 4322 -828 4832 -792
rect 4322 -852 4358 -828
rect 4796 -852 4832 -828
rect 5128 -852 5550 -844
rect 6716 -852 6752 -710
rect 476 -888 1232 -852
rect 2656 -888 4322 -852
rect 4832 -888 5128 -852
rect 5550 -878 6752 -852
rect 6028 -888 6752 -878
rect 4496 -1834 4554 -1828
rect 4716 -1834 4774 -1828
rect 4496 -1868 4508 -1834
rect 4716 -1868 4728 -1834
rect 4496 -1874 4554 -1868
rect 4716 -1874 4774 -1868
rect 4562 -2074 4620 -2068
rect 4762 -2074 4820 -2068
rect 4562 -2108 4574 -2074
rect 4762 -2108 4774 -2074
rect 4562 -2114 4620 -2108
rect 4762 -2114 4820 -2108
rect 5064 -2566 5204 -2474
rect 5318 -3080 5458 -2566
rect 1866 -3614 1924 -3608
rect 1866 -3648 1878 -3614
rect 1866 -3654 1924 -3648
<< nwell >>
rect 4728 -1280 4794 -1210
rect 1244 -1518 1310 -1516
rect 1244 -1582 1314 -1518
rect 2012 -1528 2076 -1520
rect 2574 -1614 2638 -1606
<< nsubdiff >>
rect 512 -852 6716 -710
<< poly >>
rect 4728 -1226 4794 -1210
rect 4728 -1260 4744 -1226
rect 4778 -1260 4794 -1226
rect 4728 -1280 4794 -1260
rect 1226 -1516 1256 -1414
rect 1226 -1532 1310 -1516
rect 1226 -1566 1260 -1532
rect 1294 -1566 1310 -1532
rect 1226 -1582 1310 -1566
rect 1226 -1829 1256 -1582
rect 2630 -1608 2660 -1412
rect 2574 -1624 2660 -1608
rect 5324 -1622 5354 -1231
rect 2574 -1658 2590 -1624
rect 2624 -1658 2660 -1624
rect 2574 -1674 2660 -1658
rect 2630 -1784 2660 -1674
rect 4576 -2682 4606 -2344
rect 4776 -2682 4806 -2305
rect 4978 -2394 5008 -2296
rect 4942 -2410 5008 -2394
rect 4942 -2444 4958 -2410
rect 4992 -2444 5008 -2410
rect 4942 -2460 5008 -2444
rect 4978 -2682 5008 -2460
rect 5514 -2785 5544 -2337
<< polycont >>
rect 4744 -1260 4778 -1226
rect 1260 -1566 1294 -1532
rect 2590 -1658 2624 -1624
rect 4958 -2444 4992 -2410
<< locali >>
rect 508 -730 6712 -710
rect 508 -732 3130 -730
rect 508 -836 538 -732
rect 646 -836 754 -732
rect 862 -836 970 -732
rect 1078 -836 1186 -732
rect 1294 -836 1402 -732
rect 1510 -836 1618 -732
rect 1726 -836 1834 -732
rect 1942 -836 2050 -732
rect 2158 -836 2266 -732
rect 2374 -836 2482 -732
rect 2590 -836 2698 -732
rect 2806 -836 2914 -732
rect 3022 -834 3130 -732
rect 3238 -834 3346 -730
rect 3454 -834 3562 -730
rect 3670 -834 3778 -730
rect 3886 -834 3994 -730
rect 4102 -834 4210 -730
rect 4318 -834 4426 -730
rect 4534 -834 4642 -730
rect 4750 -834 4858 -730
rect 4966 -834 5074 -730
rect 5182 -834 5290 -730
rect 5398 -834 5506 -730
rect 5614 -834 5722 -730
rect 5830 -834 5938 -730
rect 6046 -834 6154 -730
rect 6262 -834 6370 -730
rect 6478 -834 6586 -730
rect 6694 -834 6712 -730
rect 3022 -836 6712 -834
rect 508 -852 6712 -836
rect 1578 -1066 1624 -852
rect 1866 -1050 1912 -852
rect 1978 -1032 2024 -852
rect 2266 -1030 2312 -852
rect 4728 -1260 4744 -1226
rect 4778 -1260 4794 -1226
rect 1244 -1566 1260 -1532
rect 1294 -1566 1310 -1532
rect 2574 -1658 2590 -1624
rect 2624 -1658 2640 -1624
rect 4942 -2444 4958 -2410
rect 4992 -2444 5008 -2410
rect 1322 -4632 2964 -4614
rect 1322 -4634 1468 -4632
rect 1322 -4692 1360 -4634
rect 1414 -4690 1468 -4634
rect 1522 -4690 1574 -4632
rect 1628 -4690 1682 -4632
rect 1736 -4634 2094 -4632
rect 1736 -4690 1792 -4634
rect 1414 -4692 1792 -4690
rect 1846 -4692 1894 -4634
rect 1948 -4692 1994 -4634
rect 2048 -4690 2094 -4634
rect 2148 -4690 2194 -4632
rect 2248 -4634 2494 -4632
rect 2248 -4690 2292 -4634
rect 2048 -4692 2292 -4690
rect 2346 -4692 2394 -4634
rect 2448 -4690 2494 -4634
rect 2548 -4634 2692 -4632
rect 2548 -4690 2594 -4634
rect 2448 -4692 2594 -4690
rect 2648 -4690 2692 -4634
rect 2746 -4690 2792 -4632
rect 2846 -4690 2892 -4632
rect 2946 -4690 2964 -4632
rect 2648 -4692 2964 -4690
rect 1322 -4712 2964 -4692
<< viali >>
rect 538 -836 646 -732
rect 754 -836 862 -732
rect 970 -836 1078 -732
rect 1186 -836 1294 -732
rect 1402 -836 1510 -732
rect 1618 -836 1726 -732
rect 1834 -836 1942 -732
rect 2050 -836 2158 -732
rect 2266 -836 2374 -732
rect 2482 -836 2590 -732
rect 2698 -836 2806 -732
rect 2914 -836 3022 -732
rect 3130 -834 3238 -730
rect 3346 -834 3454 -730
rect 3562 -834 3670 -730
rect 3778 -834 3886 -730
rect 3994 -834 4102 -730
rect 4210 -834 4318 -730
rect 4426 -834 4534 -730
rect 4642 -834 4750 -730
rect 4858 -834 4966 -730
rect 5074 -834 5182 -730
rect 5290 -834 5398 -730
rect 5506 -834 5614 -730
rect 5722 -834 5830 -730
rect 5938 -834 6046 -730
rect 6154 -834 6262 -730
rect 6370 -834 6478 -730
rect 6586 -834 6694 -730
rect 4744 -1260 4778 -1226
rect 1260 -1566 1294 -1532
rect 2590 -1658 2624 -1624
rect 4958 -2444 4992 -2410
rect 1360 -4692 1414 -4634
rect 1468 -4690 1522 -4632
rect 1574 -4690 1628 -4632
rect 1682 -4690 1736 -4632
rect 1792 -4692 1846 -4634
rect 1894 -4692 1948 -4634
rect 1994 -4692 2048 -4634
rect 2094 -4690 2148 -4632
rect 2194 -4690 2248 -4632
rect 2292 -4692 2346 -4634
rect 2394 -4692 2448 -4634
rect 2494 -4690 2548 -4632
rect 2594 -4692 2648 -4634
rect 2692 -4690 2746 -4632
rect 2792 -4690 2846 -4632
rect 2892 -4690 2946 -4632
<< metal1 >>
rect -870 112 -670 312
rect -870 -288 -670 -88
rect -870 -688 -670 -488
rect 508 -710 708 -652
rect 2188 -710 2440 -708
rect 508 -730 6716 -710
rect 508 -732 3130 -730
rect 508 -836 538 -732
rect 646 -836 754 -732
rect 862 -836 970 -732
rect 1078 -836 1186 -732
rect 1294 -836 1402 -732
rect 1510 -836 1618 -732
rect 1726 -836 1834 -732
rect 1942 -836 2050 -732
rect 2158 -836 2266 -732
rect 2374 -836 2482 -732
rect 2590 -836 2698 -732
rect 2806 -836 2914 -732
rect 3022 -834 3130 -732
rect 3238 -834 3346 -730
rect 3454 -834 3562 -730
rect 3670 -834 3778 -730
rect 3886 -834 3994 -730
rect 4102 -834 4210 -730
rect 4318 -834 4426 -730
rect 4534 -834 4642 -730
rect 4750 -834 4858 -730
rect 4966 -834 5074 -730
rect 5182 -834 5290 -730
rect 5398 -834 5506 -730
rect 5614 -834 5722 -730
rect 5830 -834 5938 -730
rect 6046 -834 6154 -730
rect 6262 -834 6370 -730
rect 6478 -834 6586 -730
rect 6694 -834 6716 -730
rect 3022 -836 6716 -834
rect 508 -852 6716 -836
rect 1536 -854 1578 -852
rect 2518 -856 2670 -852
rect 4732 -1226 4790 -1220
rect 4732 -1260 4744 -1226
rect 4778 -1260 4790 -1226
rect -870 -1488 -670 -1288
rect -870 -1888 -670 -1688
rect 748 -1776 794 -1330
rect 1174 -1440 1220 -1350
rect 1702 -1364 1788 -1346
rect 1696 -1392 1800 -1364
rect 2096 -1366 2182 -1344
rect 1702 -1396 1788 -1392
rect 2096 -1394 2206 -1366
rect 982 -1486 1220 -1440
rect 982 -1744 1040 -1486
rect 748 -1822 990 -1776
rect 1174 -1878 1220 -1486
rect 1414 -1498 1472 -1438
rect 1616 -1496 1674 -1448
rect 1250 -1524 1314 -1518
rect 1740 -1520 1786 -1396
rect 1250 -1526 1256 -1524
rect 1248 -1576 1256 -1526
rect 1308 -1576 1314 -1524
rect 1248 -1582 1314 -1576
rect 1724 -1526 1788 -1520
rect 1724 -1578 1730 -1526
rect 1782 -1578 1788 -1526
rect 1724 -1584 1788 -1578
rect 1732 -1784 1778 -1584
rect 1816 -1606 1874 -1442
rect 2016 -1520 2074 -1444
rect 2012 -1526 2076 -1520
rect 2012 -1578 2018 -1526
rect 2070 -1578 2076 -1526
rect 2012 -1584 2076 -1578
rect 1812 -1612 1876 -1606
rect 1812 -1664 1818 -1612
rect 1870 -1664 1876 -1612
rect 1812 -1670 1876 -1664
rect 1816 -1740 1874 -1670
rect 2016 -1724 2074 -1584
rect 2104 -1606 2150 -1394
rect 2216 -1494 2274 -1436
rect 2416 -1494 2474 -1436
rect 2666 -1438 2712 -1342
rect 2666 -1484 2904 -1438
rect 2104 -1612 2168 -1606
rect 2104 -1664 2110 -1612
rect 2162 -1664 2168 -1612
rect 2104 -1670 2168 -1664
rect 2574 -1612 2638 -1606
rect 2574 -1664 2580 -1612
rect 2632 -1664 2638 -1612
rect 2574 -1670 2638 -1664
rect 2112 -1784 2158 -1670
rect 1732 -1786 1818 -1784
rect 1732 -1832 1824 -1786
rect 1732 -1834 1818 -1832
rect 2072 -1834 2158 -1784
rect 2666 -1870 2712 -1484
rect 2846 -1742 2904 -1484
rect 3092 -1772 3138 -1326
rect 4732 -1410 4790 -1260
rect 4458 -1454 4790 -1410
rect 4458 -1670 4504 -1454
rect 4732 -1456 4790 -1454
rect 5364 -1272 5410 -1172
rect 5364 -1318 5650 -1272
rect 4760 -1494 4826 -1488
rect 4760 -1546 4768 -1494
rect 4820 -1546 4826 -1494
rect 4760 -1552 4826 -1546
rect 4766 -1656 4812 -1552
rect 5364 -1700 5410 -1318
rect 5592 -1576 5650 -1318
rect 2896 -1818 3138 -1772
rect -870 -2288 -670 -2088
rect 1472 -2156 1530 -2098
rect 1664 -2222 1710 -2014
rect 2370 -2158 2428 -2100
rect 4616 -2228 4764 -2156
rect 4612 -2302 4764 -2228
rect 4612 -2410 4658 -2302
rect 4946 -2410 5004 -2404
rect 4612 -2444 4958 -2410
rect 4992 -2444 5006 -2410
rect 4612 -2446 5006 -2444
rect -870 -2688 -670 -2488
rect 1278 -2702 1328 -2574
rect 1664 -2628 1710 -2578
rect 1866 -2628 1912 -2574
rect 1664 -2674 1912 -2628
rect 1978 -2628 2024 -2576
rect 2178 -2628 2224 -2578
rect 1978 -2674 2224 -2628
rect 2560 -2702 2610 -2560
rect 4672 -2662 4712 -2446
rect 4946 -2450 5004 -2446
rect 1278 -2748 2610 -2702
rect -870 -3088 -670 -2888
rect 1916 -2922 1962 -2748
rect 4612 -2858 4770 -2662
rect 5550 -2700 5596 -2306
rect 5778 -2700 5836 -2442
rect 5550 -2746 5836 -2700
rect 5550 -2834 5596 -2746
rect -870 -3488 -670 -3288
rect -870 -3888 -670 -3688
rect -870 -4288 -670 -4088
rect -870 -4688 -670 -4488
rect 1320 -4632 2962 -4612
rect 1320 -4634 1468 -4632
rect 1320 -4692 1360 -4634
rect 1414 -4690 1468 -4634
rect 1522 -4690 1574 -4632
rect 1628 -4690 1682 -4632
rect 1736 -4634 2094 -4632
rect 1736 -4690 1792 -4634
rect 1414 -4692 1792 -4690
rect 1846 -4692 1894 -4634
rect 1948 -4692 1994 -4634
rect 2048 -4690 2094 -4634
rect 2148 -4690 2194 -4632
rect 2248 -4634 2494 -4632
rect 2248 -4690 2292 -4634
rect 2048 -4692 2292 -4690
rect 2346 -4692 2394 -4634
rect 2448 -4690 2494 -4634
rect 2548 -4634 2692 -4632
rect 2548 -4690 2594 -4634
rect 2448 -4692 2594 -4690
rect 2648 -4690 2692 -4634
rect 2746 -4690 2792 -4632
rect 2846 -4690 2892 -4632
rect 2946 -4690 2962 -4632
rect 2648 -4692 2962 -4690
rect 1320 -4710 2962 -4692
rect -870 -5088 -670 -4888
<< via1 >>
rect 1256 -1532 1308 -1524
rect 1256 -1566 1260 -1532
rect 1260 -1566 1294 -1532
rect 1294 -1566 1308 -1532
rect 1256 -1576 1308 -1566
rect 1730 -1578 1782 -1526
rect 2018 -1578 2070 -1526
rect 1818 -1664 1870 -1612
rect 2110 -1664 2162 -1612
rect 2580 -1624 2632 -1612
rect 2580 -1658 2590 -1624
rect 2590 -1658 2624 -1624
rect 2624 -1658 2632 -1624
rect 2580 -1664 2632 -1658
rect 4768 -1546 4820 -1494
<< metal2 >>
rect 1250 -1524 1314 -1518
rect 1724 -1524 1788 -1520
rect 1250 -1576 1256 -1524
rect 1308 -1526 1788 -1524
rect 2012 -1526 2076 -1520
rect 1308 -1576 1730 -1526
rect 1250 -1582 1314 -1576
rect 1724 -1578 1730 -1576
rect 1782 -1578 2018 -1526
rect 2070 -1578 2076 -1526
rect 4532 -1548 4598 -1502
rect 1724 -1584 1788 -1578
rect 2012 -1584 2076 -1578
rect 1812 -1612 1876 -1606
rect 1812 -1664 1818 -1612
rect 1870 -1614 1876 -1612
rect 2104 -1612 2168 -1606
rect 2574 -1612 2638 -1606
rect 2104 -1614 2110 -1612
rect 1870 -1664 2110 -1614
rect 2162 -1664 2580 -1612
rect 2632 -1664 2638 -1612
rect 1812 -1670 1876 -1664
rect 2104 -1670 2168 -1664
rect 2574 -1670 2638 -1664
<< rmetal2 >>
rect 4506 -1502 4558 -1268
rect 4760 -1494 4826 -1488
rect 4760 -1502 4768 -1494
rect 4506 -1548 4532 -1502
rect 4598 -1546 4768 -1502
rect 4820 -1546 4826 -1494
rect 4598 -1548 4826 -1546
rect 4760 -1552 4826 -1548
use sky130_fd_pr__nfet_01v8_PWNS5P  XM1
timestamp 1697007148
transform 1 0 1895 0 -1 -3176
box -73 -430 73 488
use sky130_fd_pr__nfet_01v8_lvt_F5PS5H  XM2
timestamp 1697420474
transform 1 0 2393 0 1 -2392
box -221 -226 221 290
use sky130_fd_pr__nfet_01v8_lvt_F5PS5H  XM3
timestamp 1697420474
transform 1 0 1495 0 1 -2390
box -221 -226 221 290
use sky130_fd_pr__nfet_01v8_PWNS5P  XM4
timestamp 1697007148
transform 1 0 1845 0 1 -2186
box -73 -430 73 488
use sky130_fd_pr__nfet_01v8_PWNS5P  XM5
timestamp 1697007148
transform 1 0 2045 0 1 -2188
box -73 -430 73 488
use sky130_fd_pr__pfet_01v8_XGAKDL  XM6
timestamp 1697360394
transform 1 0 1845 0 1 -1195
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XGAKDL  XM7
timestamp 1697360394
transform 1 0 2045 0 1 -1195
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XGAKDL  XM8
timestamp 1697360394
transform 1 0 1645 0 1 -1197
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XGAKDL  XM9
timestamp 1697360394
transform 1 0 1443 0 1 -1197
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XGAKDL  XM10
timestamp 1697360394
transform 1 0 2245 0 1 -1195
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XGAKDL  XM11
timestamp 1697360394
transform 1 0 2445 0 1 -1195
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_MQX2PY  XM12
timestamp 1697008372
transform 1 0 2645 0 1 -1311
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_L7T3GD  XM13
timestamp 1697008372
transform 1 0 2645 0 1 -1852
box -73 -80 73 80
use sky130_fd_pr__pfet_01v8_HFBCFR  XM14
timestamp 1697012471
transform 1 0 2971 0 1 -1330
box -311 -286 311 286
use sky130_fd_pr__nfet_01v8_648S5X  XM15
timestamp 1697012471
transform 1 0 2875 0 1 -1872
box -73 -138 73 188
use sky130_fd_pr__pfet_01v8_MQX2PY  XM16
timestamp 1697008372
transform 1 0 4533 0 1 -1095
box -211 -303 211 303
use sky130_fd_pr__pfet_01v8_MQX2PY  XM17
timestamp 1697008372
transform 1 0 4621 0 1 -1095
box -211 -303 211 303
use sky130_fd_pr__pfet_01v8_MQX2PY  XM18
timestamp 1697008372
transform -1 0 1241 0 1 -1313
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_9NW3WL  XM19
timestamp 1697022684
transform 1 0 4745 0 -1 -1712
box -73 -122 73 172
use sky130_fd_pr__nfet_01v8_L7T3GD  XM20
timestamp 1697008372
transform -1 0 1239 0 1 -1890
box -73 -80 73 80
use sky130_fd_pr__pfet_01v8_HFBCFR  XM21
timestamp 1697012471
transform -1 0 915 0 1 -1332
box -311 -286 311 286
use sky130_fd_pr__nfet_01v8_648S5X  XM22
timestamp 1697012471
transform -1 0 1011 0 1 -1876
box -73 -138 73 188
use sky130_fd_pr__nfet_01v8_9NW3WL  XM23
timestamp 1697022684
transform 1 0 4525 0 -1 -1712
box -73 -122 73 172
use sky130_fd_pr__pfet_01v8_MQX2PY  XM24
timestamp 1697008372
transform 1 0 4591 0 1 -2775
box -211 -303 211 303
use sky130_fd_pr__pfet_01v8_MQX2PY  XM25
timestamp 1697008372
transform 1 0 4791 0 1 -2775
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_9NW3WL  XM26
timestamp 1697022684
transform 1 0 4591 0 1 -2230
box -73 -122 73 172
use sky130_fd_pr__nfet_01v8_9NW3WL  XM27
timestamp 1697022684
transform 1 0 4791 0 1 -2230
box -73 -122 73 172
use sky130_fd_pr__pfet_01v8_MQX2PY  XM28
timestamp 1697008372
transform 1 0 4993 0 1 -2777
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_L7T3GD  XM29
timestamp 1697008372
transform 1 0 4993 0 1 -2238
box -73 -80 73 80
use sky130_fd_pr__pfet_01v8_MQX2PY  XM30
timestamp 1697008372
transform 1 0 5339 0 1 -1147
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_L7T3GD  XM31
timestamp 1697008372
transform 1 0 5339 0 1 -1698
box -73 -80 73 80
use sky130_fd_pr__pfet_01v8_HFBCFR  XM32
timestamp 1697012471
transform 1 0 5717 0 1 -1164
box -311 -286 311 286
use sky130_fd_pr__nfet_01v8_648S5X  XM33
timestamp 1697012471
transform 1 0 5623 0 1 -1708
box -73 -138 73 188
use sky130_fd_pr__pfet_01v8_MQX2PY  XM34
timestamp 1697008372
transform 1 0 5529 0 -1 -2869
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_L7T3GD  XM35
timestamp 1697008372
transform 1 0 5529 0 -1 -2276
box -73 -80 73 80
use sky130_fd_pr__pfet_01v8_HFBCFR  XM36
timestamp 1697012471
transform 1 0 5903 0 -1 -2854
box -311 -286 311 286
use sky130_fd_pr__nfet_01v8_648S5X  XM37
timestamp 1697012471
transform 1 0 5807 0 -1 -2312
box -73 -138 73 188
<< labels >>
flabel metal1 508 -852 708 -652 0 FreeSans 256 0 0 0 VDD
port 3 nsew
flabel metal1 -870 112 -670 312 0 FreeSans 256 0 0 0 cdac_vn
port 0 nsew
flabel metal1 -870 -288 -670 -88 0 FreeSans 256 0 0 0 cdac_vp
port 1 nsew
flabel metal1 -870 -688 -670 -488 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 -870 -1488 -670 -1288 0 FreeSans 256 0 0 0 clk
port 4 nsew
flabel metal1 -870 -1888 -670 -1688 0 FreeSans 256 0 0 0 X
port 5 nsew
flabel metal1 -870 -2288 -670 -2088 0 FreeSans 256 0 0 0 Y
port 6 nsew
flabel metal1 -870 -2688 -670 -2488 0 FreeSans 256 0 0 0 P
port 7 nsew
flabel metal1 -870 -3088 -670 -2888 0 FreeSans 256 0 0 0 Q
port 8 nsew
flabel metal1 -870 -3488 -670 -3288 0 FreeSans 256 0 0 0 ready
port 9 nsew
flabel metal1 -870 -3888 -670 -3688 0 FreeSans 256 0 0 0 X_drive
port 10 nsew
flabel metal1 -870 -4288 -670 -4088 0 FreeSans 256 0 0 0 Y_drive
port 11 nsew
flabel metal1 -870 -4688 -670 -4488 0 FreeSans 256 0 0 0 comp_outp
port 12 nsew
flabel metal1 -870 -5088 -670 -4888 0 FreeSans 256 0 0 0 comp_outn
port 13 nsew
<< end >>
