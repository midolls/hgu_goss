magic
tech sky130A
magscale 1 2
timestamp 1699867178
<< nwell >>
rect -3292 7457 -3185 7829
rect -3397 6176 -3134 6839
<< metal1 >>
rect -8566 13489 -8560 13541
rect -8508 13539 -8502 13541
rect -8508 13492 -8447 13539
rect -8508 13489 -8502 13492
rect -6358 9032 -6352 9084
rect -6300 9032 -6294 9084
rect -6058 8808 -878 8838
rect -6058 8739 -878 8769
rect -6058 8669 -878 8699
rect -6058 8599 -878 8629
rect -6058 8530 -878 8560
rect -6058 8460 -878 8490
rect -6058 8390 -878 8420
rect -6058 8320 -878 8350
rect -6058 8251 -878 8281
rect -6058 8181 -878 8211
rect -6058 8112 -878 8142
rect -6058 8042 -878 8072
rect -6058 7972 -878 8002
rect -8565 7652 -8559 7704
rect -8507 7690 -8501 7704
rect -3334 7692 -3158 7788
rect -8507 7662 -5970 7690
rect -8507 7652 -8501 7662
rect -5998 5600 -5970 7662
rect -3447 7052 -3150 7244
rect -3443 6412 -3146 6604
rect -3421 5868 -3160 5964
rect -5397 5659 -5391 5675
rect -5422 5624 -5391 5659
rect -5397 5623 -5391 5624
rect -5339 5659 -5333 5675
rect -5339 5624 164 5659
rect -5339 5623 -5333 5624
rect -6011 5548 -6005 5600
rect -5953 5548 -5947 5600
rect -1314 5466 -1308 5518
rect -1256 5507 -1250 5518
rect -1128 5507 -1122 5517
rect -1256 5477 -1122 5507
rect -1256 5466 -1250 5477
rect -1128 5465 -1122 5477
rect -1070 5465 -1064 5517
rect -1589 5397 -1583 5449
rect -1531 5437 -1525 5449
rect -1214 5437 -1208 5447
rect -1531 5407 -1208 5437
rect -1531 5397 -1525 5407
rect -1214 5395 -1208 5407
rect -1156 5395 -1150 5447
rect -1864 5327 -1858 5379
rect -1806 5367 -1800 5379
rect -1301 5367 -1295 5378
rect -1806 5337 -1295 5367
rect -1806 5327 -1800 5337
rect -1301 5326 -1295 5337
rect -1243 5326 -1237 5378
rect -2406 5257 -2400 5309
rect -2348 5298 -2342 5309
rect -1387 5298 -1381 5308
rect -2348 5268 -1381 5298
rect -2348 5257 -2342 5268
rect -1387 5256 -1381 5268
rect -1329 5256 -1323 5308
rect -2971 5188 -2965 5240
rect -2913 5228 -2907 5240
rect -1474 5228 -1468 5239
rect -2913 5198 -1468 5228
rect -2913 5188 -2907 5198
rect -1474 5187 -1468 5198
rect -1416 5187 -1410 5239
rect -3264 5118 -3258 5170
rect -3206 5159 -3200 5170
rect -1560 5159 -1554 5169
rect -3206 5129 -1554 5159
rect -3206 5118 -3200 5129
rect -1560 5117 -1554 5129
rect -1502 5117 -1496 5169
rect -3350 5048 -3344 5100
rect -3292 5089 -3286 5100
rect -1646 5089 -1640 5099
rect -3292 5059 -1640 5089
rect -3292 5048 -3286 5059
rect -1646 5047 -1640 5059
rect -1588 5047 -1582 5099
rect -3497 4978 -3491 5030
rect -3439 5019 -3433 5030
rect -1732 5019 -1726 5029
rect -3439 4989 -1726 5019
rect -3439 4978 -3433 4989
rect -1732 4977 -1726 4989
rect -1674 4977 -1668 5029
rect -3770 4909 -3764 4961
rect -3712 4949 -3706 4961
rect -1819 4949 -1813 4960
rect -3712 4919 -1813 4949
rect -3712 4909 -3706 4919
rect -1819 4908 -1813 4919
rect -1761 4908 -1755 4960
rect -4049 4839 -4043 4891
rect -3991 4880 -3985 4891
rect -1905 4880 -1899 4890
rect -3991 4850 -1899 4880
rect -3991 4839 -3985 4850
rect -1905 4838 -1899 4850
rect -1847 4838 -1841 4890
rect -4596 4770 -4590 4822
rect -4538 4810 -4532 4822
rect -1991 4810 -1985 4820
rect -4538 4780 -1985 4810
rect -4538 4770 -4532 4780
rect -1991 4768 -1985 4780
rect -1933 4768 -1927 4820
rect -5147 4700 -5141 4752
rect -5089 4740 -5083 4752
rect -2078 4740 -2072 4751
rect -5089 4710 -2072 4740
rect -5089 4700 -5083 4710
rect -2078 4699 -2072 4710
rect -2020 4699 -2014 4751
rect -1352 -152 -1346 -100
rect -1294 -110 -1288 -100
rect -1294 -140 14484 -110
rect -1294 -152 -1288 -140
rect -804 -222 -798 -170
rect -746 -180 -740 -170
rect -746 -210 14484 -180
rect -746 -222 -740 -210
rect -537 -291 -531 -239
rect -479 -250 -473 -239
rect -479 -280 14484 -250
rect -479 -291 -473 -280
rect -251 -361 -245 -309
rect -193 -319 -187 -309
rect -193 -349 14484 -319
rect -193 -361 -187 -349
rect -24 -430 -18 -378
rect 34 -389 40 -378
rect 34 -419 14484 -389
rect 34 -430 40 -419
rect 62 -500 68 -448
rect 120 -458 126 -448
rect 120 -488 14484 -458
rect 120 -500 126 -488
rect 448 -570 454 -518
rect 506 -528 512 -518
rect 506 -558 14484 -528
rect 506 -570 512 -558
rect 994 -640 1000 -588
rect 1052 -598 1058 -588
rect 1052 -628 14484 -598
rect 1052 -640 1058 -628
rect 1541 -709 1547 -657
rect 1599 -668 1605 -657
rect 1599 -698 14484 -668
rect 1599 -709 1605 -698
rect 1827 -779 1833 -727
rect 1885 -737 1891 -727
rect 1885 -767 14484 -737
rect 1885 -779 1891 -767
rect 2093 -849 2099 -797
rect 2151 -807 2157 -797
rect 2151 -837 14484 -807
rect 2151 -849 2157 -837
rect 2240 -918 2246 -866
rect 2298 -877 2304 -866
rect 2298 -907 14484 -877
rect 2298 -918 2304 -907
rect 2327 -987 2333 -935
rect 2385 -946 2391 -935
rect 2385 -976 14484 -946
rect 2385 -987 2391 -976
rect -2409 -3092 2642 -3062
rect -2409 -3161 2642 -3131
rect -2409 -3231 2642 -3201
rect -2409 -3301 2642 -3271
rect -2409 -3370 2642 -3340
rect -2409 -3440 2642 -3410
rect -2409 -3510 2642 -3480
rect -2409 -3580 2642 -3550
rect -2409 -3649 2642 -3619
rect -2409 -3719 2642 -3689
rect -2409 -3788 2642 -3758
rect -2409 -3858 2642 -3828
rect -2409 -3928 2642 -3898
<< via1 >>
rect -8560 13489 -8508 13541
rect -6352 9032 -6300 9084
rect -8559 7652 -8507 7704
rect -5391 5623 -5339 5675
rect -6005 5548 -5953 5600
rect -1308 5466 -1256 5518
rect -1122 5465 -1070 5517
rect -1583 5397 -1531 5449
rect -1208 5395 -1156 5447
rect -1858 5327 -1806 5379
rect -1295 5326 -1243 5378
rect -2400 5257 -2348 5309
rect -1381 5256 -1329 5308
rect -2965 5188 -2913 5240
rect -1468 5187 -1416 5239
rect -3258 5118 -3206 5170
rect -1554 5117 -1502 5169
rect -3344 5048 -3292 5100
rect -1640 5047 -1588 5099
rect -3491 4978 -3439 5030
rect -1726 4977 -1674 5029
rect -3764 4909 -3712 4961
rect -1813 4908 -1761 4960
rect -4043 4839 -3991 4891
rect -1899 4838 -1847 4890
rect -4590 4770 -4538 4822
rect -1985 4768 -1933 4820
rect -5141 4700 -5089 4752
rect -2072 4699 -2020 4751
rect -1346 -152 -1294 -100
rect -798 -222 -746 -170
rect -531 -291 -479 -239
rect -245 -361 -193 -309
rect -18 -430 34 -378
rect 68 -500 120 -448
rect 454 -570 506 -518
rect 1000 -640 1052 -588
rect 1547 -709 1599 -657
rect 1833 -779 1885 -727
rect 2099 -849 2151 -797
rect 2246 -918 2298 -866
rect 2333 -987 2385 -935
<< metal2 >>
rect -8566 13489 -8560 13541
rect -8508 13489 -8502 13541
rect -8552 7704 -8524 13489
rect -6358 9032 -6352 9084
rect -6300 9032 -6294 9084
rect -8565 7652 -8559 7704
rect -8507 7652 -8501 7704
rect -6338 7615 -6310 9032
rect -5397 5623 -5391 5675
rect -5339 5623 -5333 5675
rect -6011 5548 -6005 5600
rect -5953 5548 -5947 5600
rect -5135 4752 -5093 5532
rect -4586 4822 -4544 5532
rect -4038 4891 -3996 5532
rect -3758 4961 -3716 5532
rect -3486 5030 -3444 5532
rect -3339 5100 -3297 5532
rect -3252 5170 -3210 5532
rect -2959 5240 -2917 5532
rect -2395 5309 -2353 5532
rect -1852 5379 -1810 5532
rect -1578 5449 -1536 5532
rect -1303 5518 -1261 5532
rect -1314 5466 -1308 5518
rect -1256 5466 -1250 5518
rect -1128 5465 -1122 5517
rect -1070 5465 -1064 5517
rect -1589 5397 -1583 5449
rect -1531 5397 -1525 5449
rect -1214 5395 -1208 5447
rect -1156 5395 -1150 5447
rect -1864 5327 -1858 5379
rect -1806 5327 -1800 5379
rect -1301 5326 -1295 5378
rect -1243 5326 -1237 5378
rect -2406 5257 -2400 5309
rect -2348 5257 -2342 5309
rect -1387 5256 -1381 5308
rect -1329 5256 -1323 5308
rect -2971 5188 -2965 5240
rect -2913 5188 -2907 5240
rect -1474 5187 -1468 5239
rect -1416 5187 -1410 5239
rect -3264 5118 -3258 5170
rect -3206 5118 -3200 5170
rect -1560 5117 -1554 5169
rect -1502 5117 -1496 5169
rect -3350 5048 -3344 5100
rect -3292 5048 -3286 5100
rect -1646 5047 -1640 5099
rect -1588 5047 -1582 5099
rect -3497 4978 -3491 5030
rect -3439 4978 -3433 5030
rect -1732 4977 -1726 5029
rect -1674 4977 -1668 5029
rect -3770 4909 -3764 4961
rect -3712 4909 -3706 4961
rect -1819 4908 -1813 4960
rect -1761 4908 -1755 4960
rect -4049 4839 -4043 4891
rect -3991 4839 -3985 4891
rect -1905 4838 -1899 4890
rect -1847 4838 -1841 4890
rect -4596 4770 -4590 4822
rect -4538 4770 -4532 4822
rect -1991 4768 -1985 4820
rect -1933 4768 -1927 4820
rect -5147 4700 -5141 4752
rect -5089 4700 -5083 4752
rect -2078 4699 -2072 4751
rect -2020 4699 -2014 4751
rect -2062 4591 -2020 4699
rect -1980 4591 -1938 4768
rect -1896 4591 -1854 4838
rect -1808 4591 -1766 4908
rect -1721 4591 -1679 4977
rect -1635 4591 -1593 5047
rect -1549 4591 -1507 5117
rect -1462 4591 -1420 5187
rect -1376 4591 -1334 5256
rect -1290 4591 -1248 5326
rect -1203 4591 -1161 5395
rect -1118 4591 -1076 5465
rect -1031 4592 -989 8902
rect -944 4592 -902 8902
rect -1352 -152 -1346 -100
rect -1294 -152 -1288 -100
rect -1340 -1031 -1298 -152
rect -804 -222 -798 -170
rect -746 -222 -740 -170
rect -794 -1031 -752 -222
rect -537 -291 -531 -239
rect -479 -291 -473 -239
rect -526 -1031 -484 -291
rect -251 -361 -245 -309
rect -193 -361 -187 -309
rect -239 -1031 -197 -361
rect -24 -430 -18 -378
rect 34 -430 40 -378
rect -13 -1031 29 -430
rect 62 -500 68 -448
rect 120 -500 126 -448
rect 73 -1031 115 -500
rect 448 -570 454 -518
rect 506 -570 512 -518
rect 460 -1031 502 -570
rect 994 -640 1000 -588
rect 1052 -640 1058 -588
rect 1006 -1031 1048 -640
rect 1541 -709 1547 -657
rect 1599 -709 1605 -657
rect 1552 -1031 1594 -709
rect 1827 -779 1833 -727
rect 1885 -779 1891 -727
rect 1839 -1031 1881 -779
rect 2093 -849 2099 -797
rect 2151 -849 2157 -797
rect 2104 -1031 2146 -849
rect 2240 -918 2246 -866
rect 2298 -918 2304 -866
rect 2251 -1031 2293 -918
rect 2327 -987 2333 -935
rect 2385 -987 2391 -935
rect 2338 -1031 2380 -987
<< metal4 >>
rect -5346 9209 -4382 9215
rect -5756 9030 -4382 9209
rect -5756 8938 -5568 9030
rect -5378 9028 -4382 9030
rect -5378 8938 -5174 9028
rect -5756 8936 -5174 8938
rect -4984 9026 -4382 9028
rect -4984 8936 -4767 9026
rect -5756 8934 -4767 8936
rect -4577 8934 -4382 9026
rect -5756 7770 -4382 8934
rect -3171 9018 -2207 9177
rect -3171 8926 -3042 9018
rect -2852 9014 -2207 9018
rect -2852 8926 -2616 9014
rect -3171 8922 -2616 8926
rect -2426 8922 -2207 9014
rect -5756 7764 -4792 7770
rect -5756 5870 -5344 7764
rect -3171 7733 -2207 8922
rect -6144 4549 -5862 5189
rect -4300 4549 -3323 5974
rect -1171 5863 -699 7792
rect -6144 4255 -2585 4549
rect -6144 4251 -5862 4255
use hgu_cdac_half  hgu_cdac_half_0
timestamp 1699830634
transform 1 0 -49110 0 -1 6793
box -314 0 39606 5813
use hgu_cdac_half  hgu_cdac_half_1
timestamp 1699830634
transform 1 0 -49110 0 1 7572
box -314 0 39606 5813
use hgu_cdac_sw_buffer  hgu_cdac_sw_buffer_0
timestamp 1699539897
transform -1 0 -315 0 -1 -3771
box -270 -2798 1830 -714
use hgu_cdac_sw_buffer  hgu_cdac_sw_buffer_1
timestamp 1699539897
transform -1 0 2039 0 -1 -3767
box -270 -2798 1830 -714
use hgu_cdac_sw_buffer  hgu_cdac_sw_buffer_2
timestamp 1699539897
transform -1 0 -1376 0 1 8596
box -270 -2798 1830 -714
use hgu_cdac_sw_buffer  hgu_cdac_sw_buffer_3
timestamp 1699539897
transform -1 0 -3554 0 1 8596
box -270 -2798 1830 -714
use hgu_comp_flat  hgu_comp_flat_0
timestamp 1698719859
transform 1 0 -9082 0 1 7042
box 338 -1940 3788 618
use hgu_sarlogic_flat  hgu_sarlogic_flat_0
timestamp 1699766314
transform 1 0 -10778 0 1 1682
box 2064 -1908 31250 13749
use hgu_tah  hgu_tah_0
timestamp 1699832401
transform 1 0 -51339 0 1 3641
box 711 297 1858 5355
use hgu_vgen_vref  hgu_vgen_vref_0
timestamp 1699832401
transform -1 0 -50750 0 1 -30367
box 0 0 22370 76000
<< end >>
