magic
tech sky130A
magscale 1 2
timestamp 1698592390
<< nwell >>
rect 10320 2357 15469 3189
rect 10320 2218 15615 2357
rect 10320 2027 15919 2218
rect 10320 2007 15469 2027
rect 10320 1999 10488 2007
<< pwell >>
rect 10828 1117 10854 1149
rect 11434 1117 11460 1149
rect 12040 1117 12066 1149
rect 12646 1117 12672 1149
rect 13378 1117 13404 1149
rect 13984 1117 14010 1149
rect 14716 1117 14742 1149
<< nmos >>
rect 10352 1843 10438 1873
rect 10822 1855 10852 1939
rect 11428 1855 11458 1939
rect 12034 1855 12064 1939
rect 12640 1855 12670 1939
rect 13372 1855 13402 1939
rect 13978 1855 14008 1939
rect 14710 1855 14740 1939
rect 10352 1771 10438 1801
rect 10352 1699 10438 1729
rect 10352 1627 10438 1657
rect 10352 1555 10438 1585
rect 10352 1483 10438 1513
rect 10354 1380 10438 1410
rect 10354 1308 10438 1338
rect 10354 1236 10438 1266
rect 15160 681 15244 1881
rect 15419 1821 15579 1851
rect 15695 1847 15725 1931
rect 15791 1847 15821 1931
rect 15419 1733 15579 1763
<< pmos >>
rect 10823 2055 10853 2139
rect 11429 2055 11459 2139
rect 12035 2055 12065 2139
rect 12641 2055 12671 2139
rect 13247 2055 13277 2139
rect 13853 2055 13883 2139
rect 14459 2055 14489 2139
rect 15065 2055 15095 2139
<< pmoshvt >>
rect 10357 2268 10443 2298
rect 10357 2196 10443 2226
rect 15495 2232 15579 2262
rect 15495 2144 15579 2174
rect 10357 2093 10441 2123
rect 15695 2064 15725 2148
rect 15791 2064 15821 2148
<< ndiff >>
rect 10352 1918 10438 1931
rect 10352 1884 10368 1918
rect 10424 1884 10438 1918
rect 10352 1873 10438 1884
rect 10764 1927 10822 1939
rect 10764 1867 10776 1927
rect 10810 1867 10822 1927
rect 10764 1855 10822 1867
rect 10852 1927 10910 1939
rect 10852 1867 10864 1927
rect 10898 1867 10910 1927
rect 10852 1855 10910 1867
rect 11370 1927 11428 1939
rect 11370 1867 11382 1927
rect 11416 1867 11428 1927
rect 11370 1855 11428 1867
rect 11458 1927 11516 1939
rect 11458 1867 11470 1927
rect 11504 1867 11516 1927
rect 11458 1855 11516 1867
rect 11976 1927 12034 1939
rect 11976 1867 11988 1927
rect 12022 1867 12034 1927
rect 11976 1855 12034 1867
rect 12064 1927 12122 1939
rect 12064 1867 12076 1927
rect 12110 1867 12122 1927
rect 12064 1855 12122 1867
rect 12582 1927 12640 1939
rect 12582 1867 12594 1927
rect 12628 1867 12640 1927
rect 12582 1855 12640 1867
rect 12670 1927 12728 1939
rect 12670 1867 12682 1927
rect 12716 1867 12728 1927
rect 12670 1855 12728 1867
rect 13314 1927 13372 1939
rect 13314 1867 13326 1927
rect 13360 1867 13372 1927
rect 13314 1855 13372 1867
rect 13402 1927 13460 1939
rect 13402 1867 13414 1927
rect 13448 1867 13460 1927
rect 13402 1855 13460 1867
rect 13920 1927 13978 1939
rect 13920 1867 13932 1927
rect 13966 1867 13978 1927
rect 13920 1855 13978 1867
rect 14008 1927 14066 1939
rect 14008 1867 14020 1927
rect 14054 1867 14066 1927
rect 14008 1855 14066 1867
rect 14652 1927 14710 1939
rect 14652 1867 14664 1927
rect 14698 1867 14710 1927
rect 14652 1855 14710 1867
rect 14740 1927 14798 1939
rect 14740 1867 14752 1927
rect 14786 1867 14798 1927
rect 15160 1927 15244 1939
rect 15160 1893 15172 1927
rect 15232 1893 15244 1927
rect 15633 1919 15695 1931
rect 15160 1881 15244 1893
rect 15419 1897 15579 1909
rect 14740 1855 14798 1867
rect 10352 1801 10438 1843
rect 10352 1729 10438 1771
rect 10352 1657 10438 1699
rect 10352 1585 10438 1627
rect 10352 1513 10438 1555
rect 10352 1425 10438 1483
rect 10354 1410 10438 1425
rect 10354 1338 10438 1380
rect 10354 1266 10438 1308
rect 10354 1221 10438 1236
rect 10354 1187 10368 1221
rect 10424 1187 10438 1221
rect 10354 1178 10438 1187
rect 15419 1863 15431 1897
rect 15567 1863 15579 1897
rect 15419 1851 15579 1863
rect 15633 1859 15645 1919
rect 15679 1859 15695 1919
rect 15633 1847 15695 1859
rect 15725 1919 15791 1931
rect 15725 1859 15741 1919
rect 15775 1859 15791 1919
rect 15725 1847 15791 1859
rect 15821 1919 15883 1931
rect 15821 1859 15837 1919
rect 15871 1859 15883 1919
rect 15821 1847 15883 1859
rect 15419 1809 15579 1821
rect 15419 1775 15431 1809
rect 15567 1775 15579 1809
rect 15419 1763 15579 1775
rect 15419 1721 15579 1733
rect 15419 1687 15431 1721
rect 15567 1687 15579 1721
rect 15419 1675 15579 1687
rect 15160 669 15244 681
rect 15160 635 15172 669
rect 15232 635 15244 669
rect 15160 623 15244 635
<< pdiff >>
rect 10357 2345 10443 2356
rect 10357 2311 10370 2345
rect 10430 2311 10443 2345
rect 10357 2298 10443 2311
rect 15495 2308 15579 2320
rect 15495 2274 15507 2308
rect 15567 2274 15579 2308
rect 10357 2226 10443 2268
rect 15495 2262 15579 2274
rect 10357 2138 10443 2196
rect 15495 2220 15579 2232
rect 15495 2186 15507 2220
rect 15567 2186 15579 2220
rect 15495 2174 15579 2186
rect 10357 2123 10441 2138
rect 10765 2127 10823 2139
rect 10357 2081 10441 2093
rect 10357 2047 10369 2081
rect 10429 2047 10441 2081
rect 10765 2067 10777 2127
rect 10811 2067 10823 2127
rect 10765 2055 10823 2067
rect 10853 2127 10911 2139
rect 10853 2067 10865 2127
rect 10899 2067 10911 2127
rect 10853 2055 10911 2067
rect 11371 2127 11429 2139
rect 11371 2067 11383 2127
rect 11417 2067 11429 2127
rect 11371 2055 11429 2067
rect 11459 2127 11517 2139
rect 11459 2067 11471 2127
rect 11505 2067 11517 2127
rect 11459 2055 11517 2067
rect 11977 2127 12035 2139
rect 11977 2067 11989 2127
rect 12023 2067 12035 2127
rect 11977 2055 12035 2067
rect 12065 2127 12123 2139
rect 12065 2067 12077 2127
rect 12111 2067 12123 2127
rect 12065 2055 12123 2067
rect 12583 2127 12641 2139
rect 12583 2067 12595 2127
rect 12629 2067 12641 2127
rect 12583 2055 12641 2067
rect 12671 2127 12729 2139
rect 12671 2067 12683 2127
rect 12717 2067 12729 2127
rect 12671 2055 12729 2067
rect 13189 2127 13247 2139
rect 13189 2067 13201 2127
rect 13235 2067 13247 2127
rect 13189 2055 13247 2067
rect 13277 2127 13335 2139
rect 13277 2067 13289 2127
rect 13323 2067 13335 2127
rect 13277 2055 13335 2067
rect 13795 2127 13853 2139
rect 13795 2067 13807 2127
rect 13841 2067 13853 2127
rect 13795 2055 13853 2067
rect 13883 2127 13941 2139
rect 13883 2067 13895 2127
rect 13929 2067 13941 2127
rect 13883 2055 13941 2067
rect 14401 2127 14459 2139
rect 14401 2067 14413 2127
rect 14447 2067 14459 2127
rect 14401 2055 14459 2067
rect 14489 2127 14547 2139
rect 14489 2067 14501 2127
rect 14535 2067 14547 2127
rect 14489 2055 14547 2067
rect 15007 2127 15065 2139
rect 15007 2067 15019 2127
rect 15053 2067 15065 2127
rect 15007 2055 15065 2067
rect 15095 2127 15153 2139
rect 15095 2067 15107 2127
rect 15141 2067 15153 2127
rect 15495 2132 15579 2144
rect 15495 2098 15507 2132
rect 15567 2098 15579 2132
rect 15495 2086 15579 2098
rect 15633 2136 15695 2148
rect 15095 2055 15153 2067
rect 15633 2076 15645 2136
rect 15679 2076 15695 2136
rect 15633 2064 15695 2076
rect 15725 2136 15791 2148
rect 15725 2076 15741 2136
rect 15775 2076 15791 2136
rect 15725 2064 15791 2076
rect 15821 2136 15883 2148
rect 15821 2076 15837 2136
rect 15871 2076 15883 2136
rect 15821 2064 15883 2076
rect 10357 2035 10441 2047
<< ndiffc >>
rect 10368 1884 10424 1918
rect 10776 1867 10810 1927
rect 10864 1867 10898 1927
rect 11382 1867 11416 1927
rect 11470 1867 11504 1927
rect 11988 1867 12022 1927
rect 12076 1867 12110 1927
rect 12594 1867 12628 1927
rect 12682 1867 12716 1927
rect 13326 1867 13360 1927
rect 13414 1867 13448 1927
rect 13932 1867 13966 1927
rect 14020 1867 14054 1927
rect 14664 1867 14698 1927
rect 14752 1867 14786 1927
rect 15172 1893 15232 1927
rect 10368 1187 10424 1221
rect 15431 1863 15567 1897
rect 15645 1859 15679 1919
rect 15741 1859 15775 1919
rect 15837 1859 15871 1919
rect 15431 1775 15567 1809
rect 15431 1687 15567 1721
rect 15172 635 15232 669
<< pdiffc >>
rect 10370 2311 10430 2345
rect 15507 2274 15567 2308
rect 15507 2186 15567 2220
rect 10369 2047 10429 2081
rect 10777 2067 10811 2127
rect 10865 2067 10899 2127
rect 11383 2067 11417 2127
rect 11471 2067 11505 2127
rect 11989 2067 12023 2127
rect 12077 2067 12111 2127
rect 12595 2067 12629 2127
rect 12683 2067 12717 2127
rect 13201 2067 13235 2127
rect 13289 2067 13323 2127
rect 13807 2067 13841 2127
rect 13895 2067 13929 2127
rect 14413 2067 14447 2127
rect 14501 2067 14535 2127
rect 15019 2067 15053 2127
rect 15107 2067 15141 2127
rect 15507 2098 15567 2132
rect 15645 2076 15679 2136
rect 15741 2076 15775 2136
rect 15837 2076 15871 2136
<< poly >>
rect 10312 2268 10357 2298
rect 10443 2268 10474 2298
rect 10312 2226 10342 2268
rect 10312 2196 10357 2226
rect 10443 2196 10474 2226
rect 10805 2220 10871 2236
rect 10312 2141 10342 2196
rect 10260 2125 10342 2141
rect 10260 2091 10276 2125
rect 10310 2123 10342 2125
rect 10805 2186 10821 2220
rect 10855 2186 10871 2220
rect 10805 2170 10871 2186
rect 11411 2220 11477 2236
rect 11411 2186 11427 2220
rect 11461 2186 11477 2220
rect 11411 2170 11477 2186
rect 12017 2220 12083 2236
rect 12017 2186 12033 2220
rect 12067 2186 12083 2220
rect 12017 2170 12083 2186
rect 12623 2220 12689 2236
rect 12623 2186 12639 2220
rect 12673 2186 12689 2220
rect 12623 2170 12689 2186
rect 13229 2220 13295 2236
rect 13229 2186 13245 2220
rect 13279 2186 13295 2220
rect 13229 2170 13295 2186
rect 13835 2220 13901 2236
rect 13835 2186 13851 2220
rect 13885 2186 13901 2220
rect 13835 2170 13901 2186
rect 14441 2220 14507 2236
rect 14441 2186 14457 2220
rect 14491 2186 14507 2220
rect 14441 2170 14507 2186
rect 15047 2220 15113 2236
rect 15047 2186 15063 2220
rect 15097 2186 15113 2220
rect 15446 2232 15495 2262
rect 15579 2232 15610 2262
rect 15446 2211 15480 2232
rect 15047 2170 15113 2186
rect 15404 2195 15480 2211
rect 10823 2139 10853 2170
rect 11429 2139 11459 2170
rect 12035 2139 12065 2170
rect 12641 2139 12671 2170
rect 13247 2139 13277 2170
rect 13853 2139 13883 2170
rect 14459 2139 14489 2170
rect 15065 2139 15095 2170
rect 15404 2161 15414 2195
rect 15448 2174 15480 2195
rect 15448 2161 15495 2174
rect 15404 2145 15495 2161
rect 15464 2144 15495 2145
rect 15579 2144 15610 2174
rect 15695 2148 15725 2178
rect 15791 2148 15821 2174
rect 10310 2093 10357 2123
rect 10441 2093 10471 2123
rect 10310 2091 10326 2093
rect 10260 2075 10326 2091
rect 10823 2025 10853 2055
rect 11429 2025 11459 2055
rect 12035 2025 12065 2055
rect 12641 2025 12671 2055
rect 13247 2025 13277 2055
rect 13853 2025 13883 2055
rect 14459 2025 14489 2055
rect 15065 2025 15095 2055
rect 15695 2049 15725 2064
rect 15791 2049 15821 2064
rect 15695 2033 15821 2049
rect 15695 2019 15839 2033
rect 15773 2017 15839 2019
rect 15773 1983 15789 2017
rect 15823 1983 15839 2017
rect 15773 1976 15839 1983
rect 10822 1939 10852 1965
rect 11428 1939 11458 1965
rect 12034 1939 12064 1965
rect 12640 1939 12670 1965
rect 13372 1939 13402 1965
rect 13978 1939 14008 1965
rect 14710 1939 14740 1965
rect 15695 1953 15839 1976
rect 15695 1946 15821 1953
rect 10292 1873 10337 1879
rect 10292 1843 10352 1873
rect 10438 1843 10464 1873
rect 15695 1931 15725 1946
rect 15791 1931 15821 1946
rect 10292 1835 10337 1843
rect 10307 1801 10337 1835
rect 10822 1833 10852 1855
rect 11428 1833 11458 1855
rect 12034 1833 12064 1855
rect 12640 1833 12670 1855
rect 13372 1833 13402 1855
rect 13978 1833 14008 1855
rect 14710 1833 14740 1855
rect 10804 1817 10870 1833
rect 10307 1771 10352 1801
rect 10438 1771 10464 1801
rect 10804 1783 10820 1817
rect 10854 1783 10870 1817
rect 10307 1729 10337 1771
rect 10804 1767 10870 1783
rect 11410 1817 11476 1833
rect 11410 1783 11426 1817
rect 11460 1783 11476 1817
rect 11410 1767 11476 1783
rect 12016 1817 12082 1833
rect 12016 1783 12032 1817
rect 12066 1783 12082 1817
rect 12016 1767 12082 1783
rect 12622 1817 12688 1833
rect 12622 1783 12638 1817
rect 12672 1783 12688 1817
rect 12622 1767 12688 1783
rect 13354 1817 13420 1833
rect 13354 1783 13370 1817
rect 13404 1783 13420 1817
rect 13354 1767 13420 1783
rect 13960 1817 14026 1833
rect 13960 1783 13976 1817
rect 14010 1783 14026 1817
rect 13960 1767 14026 1783
rect 14692 1817 14758 1833
rect 14692 1783 14708 1817
rect 14742 1783 14758 1817
rect 14692 1767 14758 1783
rect 10307 1699 10352 1729
rect 10438 1699 10464 1729
rect 10307 1657 10337 1699
rect 10307 1627 10352 1657
rect 10438 1627 10464 1657
rect 10307 1585 10337 1627
rect 10307 1555 10352 1585
rect 10438 1555 10464 1585
rect 10307 1513 10337 1555
rect 10307 1483 10352 1513
rect 10438 1483 10464 1513
rect 10307 1410 10337 1483
rect 10307 1380 10354 1410
rect 10438 1380 10464 1410
rect 10307 1338 10337 1380
rect 10307 1308 10354 1338
rect 10438 1308 10464 1338
rect 10307 1266 10337 1308
rect 10307 1236 10354 1266
rect 10438 1236 10464 1266
rect 15134 681 15160 1881
rect 15244 1865 15332 1881
rect 15244 697 15282 1865
rect 15316 1851 15332 1865
rect 15316 1821 15419 1851
rect 15579 1821 15605 1851
rect 15695 1821 15725 1847
rect 15791 1821 15821 1847
rect 15316 1763 15404 1821
rect 15316 1733 15419 1763
rect 15579 1733 15605 1763
rect 15316 697 15332 1733
rect 15244 681 15332 697
<< polycont >>
rect 10276 2091 10310 2125
rect 10821 2186 10855 2220
rect 11427 2186 11461 2220
rect 12033 2186 12067 2220
rect 12639 2186 12673 2220
rect 13245 2186 13279 2220
rect 13851 2186 13885 2220
rect 14457 2186 14491 2220
rect 15063 2186 15097 2220
rect 15414 2161 15448 2195
rect 15789 1983 15823 2017
rect 10820 1783 10854 1817
rect 11426 1783 11460 1817
rect 12032 1783 12066 1817
rect 12638 1783 12672 1817
rect 13370 1783 13404 1817
rect 13976 1783 14010 1817
rect 14708 1783 14742 1817
rect 15282 697 15316 1865
<< locali >>
rect 10354 2311 10370 2345
rect 10430 2311 10447 2345
rect 15491 2274 15507 2308
rect 15567 2274 15583 2308
rect 10805 2186 10821 2220
rect 10855 2186 10871 2220
rect 11411 2186 11427 2220
rect 11461 2186 11477 2220
rect 12017 2186 12033 2220
rect 12067 2186 12083 2220
rect 12623 2186 12639 2220
rect 12673 2186 12689 2220
rect 13229 2186 13245 2220
rect 13279 2186 13295 2220
rect 13835 2186 13851 2220
rect 13885 2186 13901 2220
rect 14441 2186 14457 2220
rect 14491 2186 14507 2220
rect 15047 2186 15063 2220
rect 15097 2186 15113 2220
rect 15414 2195 15448 2212
rect 15491 2186 15507 2220
rect 15567 2186 15775 2220
rect 15414 2145 15448 2161
rect 10276 2125 10310 2141
rect 10276 2075 10310 2091
rect 10777 2127 10811 2143
rect 10352 2081 10444 2082
rect 10352 2047 10369 2081
rect 10429 2047 10445 2081
rect 10777 2051 10811 2067
rect 10865 2127 10899 2143
rect 10865 2051 10899 2067
rect 11383 2127 11417 2143
rect 11383 2051 11417 2067
rect 11471 2127 11505 2143
rect 11471 2051 11505 2067
rect 11989 2127 12023 2143
rect 11989 2051 12023 2067
rect 12077 2127 12111 2143
rect 12077 2051 12111 2067
rect 12595 2127 12629 2143
rect 12595 2051 12629 2067
rect 12683 2127 12717 2143
rect 12683 2051 12717 2067
rect 13201 2127 13235 2143
rect 13201 2051 13235 2067
rect 13289 2127 13323 2143
rect 13289 2051 13323 2067
rect 13807 2127 13841 2143
rect 13807 2051 13841 2067
rect 13895 2127 13929 2143
rect 13895 2051 13929 2067
rect 14413 2127 14447 2143
rect 14413 2051 14447 2067
rect 14501 2127 14535 2143
rect 14501 2051 14535 2067
rect 15019 2127 15053 2143
rect 15019 2051 15053 2067
rect 15107 2127 15141 2143
rect 15645 2136 15679 2152
rect 15491 2098 15507 2132
rect 15567 2098 15583 2132
rect 15107 2051 15141 2067
rect 15645 2060 15679 2076
rect 15741 2136 15775 2186
rect 15741 2060 15775 2076
rect 15837 2136 15871 2152
rect 15837 2060 15871 2076
rect 10352 1918 10444 2047
rect 15773 1983 15789 2017
rect 15823 1983 15839 2017
rect 10352 1884 10368 1918
rect 10424 1884 10444 1918
rect 10776 1927 10810 1943
rect 10776 1851 10810 1867
rect 10864 1927 10898 1943
rect 10864 1851 10898 1867
rect 11382 1927 11416 1943
rect 11382 1851 11416 1867
rect 11470 1927 11504 1943
rect 11470 1851 11504 1867
rect 11988 1927 12022 1943
rect 11988 1851 12022 1867
rect 12076 1927 12110 1943
rect 12076 1851 12110 1867
rect 12594 1927 12628 1943
rect 12594 1851 12628 1867
rect 12682 1927 12716 1943
rect 12682 1851 12716 1867
rect 13326 1927 13360 1943
rect 13326 1851 13360 1867
rect 13414 1927 13448 1943
rect 13414 1851 13448 1867
rect 13932 1927 13966 1943
rect 13932 1851 13966 1867
rect 14020 1927 14054 1943
rect 14020 1851 14054 1867
rect 14664 1927 14698 1943
rect 14664 1851 14698 1867
rect 14752 1927 14786 1943
rect 15156 1893 15172 1927
rect 15232 1893 15248 1927
rect 15645 1919 15679 1935
rect 14752 1851 14786 1867
rect 15282 1865 15316 1881
rect 10804 1783 10820 1817
rect 10854 1783 10870 1817
rect 11410 1783 11426 1817
rect 11460 1783 11476 1817
rect 12016 1783 12032 1817
rect 12066 1783 12082 1817
rect 12622 1783 12638 1817
rect 12672 1783 12688 1817
rect 13354 1783 13370 1817
rect 13404 1783 13420 1817
rect 13960 1783 13976 1817
rect 14010 1783 14026 1817
rect 14692 1783 14708 1817
rect 14742 1783 14758 1817
rect 10352 1187 10368 1221
rect 10424 1187 10440 1221
rect 15415 1863 15431 1897
rect 15567 1863 15583 1897
rect 15645 1843 15679 1859
rect 15741 1919 15775 1935
rect 15741 1809 15775 1859
rect 15837 1919 15871 1935
rect 15837 1843 15871 1859
rect 15415 1775 15431 1809
rect 15567 1775 15775 1809
rect 15415 1687 15431 1721
rect 15567 1687 15583 1721
rect 15282 681 15316 697
rect 15156 635 15172 669
rect 15232 635 15248 669
<< viali >>
rect 10821 2186 10855 2220
rect 11427 2186 11461 2220
rect 12033 2186 12067 2220
rect 12639 2186 12673 2220
rect 13245 2186 13279 2220
rect 13851 2186 13885 2220
rect 14457 2186 14491 2220
rect 15063 2186 15097 2220
rect 15414 2161 15448 2195
rect 10276 2091 10310 2125
rect 10369 2047 10429 2081
rect 10777 2067 10811 2127
rect 10865 2067 10899 2127
rect 11383 2067 11417 2127
rect 11471 2067 11505 2127
rect 11989 2067 12023 2127
rect 12077 2067 12111 2127
rect 12595 2067 12629 2127
rect 12683 2067 12717 2127
rect 13201 2067 13235 2127
rect 13289 2067 13323 2127
rect 13807 2067 13841 2127
rect 13895 2067 13929 2127
rect 14413 2067 14447 2127
rect 14501 2067 14535 2127
rect 15019 2067 15053 2127
rect 15107 2067 15141 2127
rect 15645 2076 15679 2136
rect 15837 2076 15871 2136
rect 15789 1983 15823 2017
rect 10776 1867 10810 1927
rect 10864 1867 10898 1927
rect 11382 1867 11416 1927
rect 11470 1867 11504 1927
rect 11988 1867 12022 1927
rect 12076 1867 12110 1927
rect 12594 1867 12628 1927
rect 12682 1867 12716 1927
rect 13326 1867 13360 1927
rect 13414 1867 13448 1927
rect 13932 1867 13966 1927
rect 14020 1867 14054 1927
rect 14664 1867 14698 1927
rect 14752 1867 14786 1927
rect 15172 1893 15232 1927
rect 10820 1783 10854 1817
rect 11426 1783 11460 1817
rect 12032 1783 12066 1817
rect 12638 1783 12672 1817
rect 13370 1783 13404 1817
rect 13976 1783 14010 1817
rect 14708 1783 14742 1817
rect 15282 697 15316 1865
rect 15645 1859 15679 1919
rect 15837 1859 15871 1919
rect 15172 635 15232 669
<< metal1 >>
rect 10809 2220 10867 3320
rect 10809 2186 10821 2220
rect 10855 2186 10867 2220
rect 10809 2180 10867 2186
rect 11415 2220 11473 3320
rect 11415 2186 11427 2220
rect 11461 2186 11473 2220
rect 11415 2180 11473 2186
rect 12021 2220 12079 3320
rect 12021 2186 12033 2220
rect 12067 2186 12079 2220
rect 12021 2180 12079 2186
rect 12627 2220 12685 3320
rect 12627 2186 12639 2220
rect 12673 2186 12685 2220
rect 12627 2180 12685 2186
rect 13233 2220 13291 3320
rect 13233 2186 13245 2220
rect 13279 2186 13291 2220
rect 13233 2180 13291 2186
rect 13839 2220 13897 3320
rect 13839 2186 13851 2220
rect 13885 2186 13897 2220
rect 13839 2180 13897 2186
rect 14445 2220 14503 3320
rect 14445 2186 14457 2220
rect 14491 2186 14503 2220
rect 14445 2180 14503 2186
rect 15051 2220 15109 3320
rect 15051 2186 15063 2220
rect 15097 2186 15109 2220
rect 15051 2180 15109 2186
rect 15408 2195 15454 2211
rect 15408 2161 15414 2195
rect 15448 2161 15454 2195
rect 15408 2149 15454 2161
rect 10258 2125 10316 2137
rect 10258 2091 10276 2125
rect 10310 2091 10316 2125
rect 10771 2127 10817 2139
rect 10771 2110 10777 2127
rect 10258 2079 10316 2091
rect 10741 2109 10777 2110
rect 10357 2081 10441 2087
rect 10357 2047 10369 2081
rect 10429 2047 10441 2081
rect 10357 2015 10441 2047
rect 10741 2045 10747 2109
rect 10811 2045 10817 2127
rect 10859 2127 10905 2139
rect 10859 2067 10865 2127
rect 10899 2067 10905 2127
rect 11377 2127 11423 2139
rect 11377 2110 11383 2127
rect 10859 2015 10905 2067
rect 11347 2109 11383 2110
rect 11347 2045 11353 2109
rect 11417 2045 11423 2127
rect 11465 2127 11511 2139
rect 11465 2067 11471 2127
rect 11505 2067 11511 2127
rect 11983 2127 12029 2139
rect 11983 2110 11989 2127
rect 11465 2015 11511 2067
rect 11953 2109 11989 2110
rect 11953 2045 11959 2109
rect 12023 2045 12029 2127
rect 12071 2127 12117 2139
rect 12071 2067 12077 2127
rect 12111 2067 12117 2127
rect 12589 2127 12635 2139
rect 12589 2110 12595 2127
rect 12071 2015 12117 2067
rect 12559 2109 12595 2110
rect 12559 2045 12565 2109
rect 12629 2045 12635 2127
rect 12677 2127 12723 2139
rect 12677 2067 12683 2127
rect 12717 2067 12723 2127
rect 13195 2127 13241 2139
rect 13195 2110 13201 2127
rect 12677 2015 12723 2067
rect 13165 2109 13201 2110
rect 13165 2045 13171 2109
rect 13235 2045 13241 2127
rect 13283 2127 13329 2139
rect 13283 2067 13289 2127
rect 13323 2067 13329 2127
rect 13801 2127 13847 2139
rect 13801 2110 13807 2127
rect 13283 2015 13329 2067
rect 13771 2109 13807 2110
rect 13771 2045 13777 2109
rect 13841 2045 13847 2127
rect 13889 2127 13935 2139
rect 13889 2067 13895 2127
rect 13929 2067 13935 2127
rect 14407 2127 14453 2139
rect 14407 2110 14413 2127
rect 13889 2015 13935 2067
rect 14377 2109 14413 2110
rect 14377 2045 14383 2109
rect 14447 2045 14453 2127
rect 14495 2127 14541 2139
rect 14495 2067 14501 2127
rect 14535 2067 14541 2127
rect 15013 2127 15059 2139
rect 15013 2110 15019 2127
rect 14495 2015 14541 2067
rect 14983 2109 15019 2110
rect 14983 2045 14989 2109
rect 15053 2045 15059 2127
rect 15101 2127 15147 2139
rect 15101 2067 15107 2127
rect 15141 2067 15147 2127
rect 15101 2015 15147 2067
rect 15414 2015 15448 2149
rect 15639 2136 15877 2148
rect 15639 2076 15645 2136
rect 15679 2076 15837 2136
rect 15871 2076 15877 2136
rect 15639 2064 15877 2076
rect 10357 1974 15448 2015
rect 15777 2017 15854 2023
rect 15777 1983 15789 2017
rect 15823 1983 15854 2017
rect 15777 1977 15854 1983
rect 10770 1927 10816 1974
rect 10770 1867 10776 1927
rect 10810 1867 10816 1927
rect 10849 1877 10856 1941
rect 10920 1877 10926 1941
rect 11376 1927 11422 1974
rect 10770 1855 10816 1867
rect 10858 1867 10864 1877
rect 10898 1867 10904 1877
rect 10858 1855 10904 1867
rect 11376 1867 11382 1927
rect 11416 1867 11422 1927
rect 11455 1877 11462 1941
rect 11526 1877 11532 1941
rect 11982 1927 12028 1974
rect 11376 1855 11422 1867
rect 11464 1867 11470 1877
rect 11504 1867 11510 1877
rect 11464 1855 11510 1867
rect 11982 1867 11988 1927
rect 12022 1867 12028 1927
rect 12061 1877 12068 1941
rect 12132 1877 12138 1941
rect 12588 1927 12634 1974
rect 11982 1855 12028 1867
rect 12070 1867 12076 1877
rect 12110 1867 12116 1877
rect 12070 1855 12116 1867
rect 12588 1867 12594 1927
rect 12628 1867 12634 1927
rect 12667 1877 12674 1941
rect 12738 1877 12744 1941
rect 13320 1927 13366 1974
rect 12588 1855 12634 1867
rect 12676 1867 12682 1877
rect 12716 1867 12722 1877
rect 12676 1855 12722 1867
rect 13320 1867 13326 1927
rect 13360 1867 13366 1927
rect 13399 1877 13406 1941
rect 13470 1877 13476 1941
rect 13926 1927 13972 1974
rect 13320 1855 13366 1867
rect 13408 1867 13414 1877
rect 13448 1867 13454 1877
rect 13408 1855 13454 1867
rect 13926 1867 13932 1927
rect 13966 1867 13972 1927
rect 14005 1877 14012 1941
rect 14076 1877 14082 1941
rect 14658 1927 14704 1974
rect 13926 1855 13972 1867
rect 14014 1867 14020 1877
rect 14054 1867 14060 1877
rect 14014 1855 14060 1867
rect 14658 1867 14664 1927
rect 14698 1867 14704 1927
rect 14737 1877 14744 1941
rect 14808 1877 14814 1941
rect 15160 1927 15244 1933
rect 15160 1893 15172 1927
rect 15232 1893 15244 1927
rect 14658 1855 14704 1867
rect 14746 1867 14752 1877
rect 14786 1867 14792 1877
rect 14746 1855 14792 1867
rect 10807 1817 10866 1823
rect 10807 1783 10820 1817
rect 10854 1783 10866 1817
rect 10807 694 10866 1783
rect 11413 1817 11472 1823
rect 11413 1783 11426 1817
rect 11460 1783 11472 1817
rect 11413 694 11472 1783
rect 12019 1817 12078 1823
rect 12019 1783 12032 1817
rect 12066 1783 12078 1817
rect 12019 694 12078 1783
rect 12625 1817 12684 1823
rect 12625 1783 12638 1817
rect 12672 1783 12684 1817
rect 12625 694 12684 1783
rect 13357 1817 13416 1823
rect 13357 1783 13370 1817
rect 13404 1783 13416 1817
rect 13357 694 13416 1783
rect 13963 1817 14022 1823
rect 13963 1783 13976 1817
rect 14010 1783 14022 1817
rect 13963 694 14022 1783
rect 14695 1817 14754 1823
rect 14695 1783 14708 1817
rect 14742 1783 14754 1817
rect 14695 694 14754 1783
rect 15160 669 15244 1893
rect 15276 1865 15322 1974
rect 15276 697 15282 1865
rect 15316 697 15322 1865
rect 15639 1919 15877 1932
rect 15639 1859 15645 1919
rect 15679 1859 15837 1919
rect 15871 1859 15877 1919
rect 15639 1847 15877 1859
rect 15276 685 15322 697
rect 15160 635 15172 669
rect 15232 635 15244 669
rect 15160 629 15244 635
<< via1 >>
rect 10747 2067 10777 2109
rect 10777 2067 10811 2109
rect 10747 2045 10811 2067
rect 11353 2067 11383 2109
rect 11383 2067 11417 2109
rect 11353 2045 11417 2067
rect 11959 2067 11989 2109
rect 11989 2067 12023 2109
rect 11959 2045 12023 2067
rect 12565 2067 12595 2109
rect 12595 2067 12629 2109
rect 12565 2045 12629 2067
rect 13171 2067 13201 2109
rect 13201 2067 13235 2109
rect 13171 2045 13235 2067
rect 13777 2067 13807 2109
rect 13807 2067 13841 2109
rect 13777 2045 13841 2067
rect 14383 2067 14413 2109
rect 14413 2067 14447 2109
rect 14383 2045 14447 2067
rect 14989 2067 15019 2109
rect 15019 2067 15053 2109
rect 14989 2045 15053 2067
rect 10856 1927 10920 1941
rect 10856 1877 10864 1927
rect 10864 1877 10898 1927
rect 10898 1877 10920 1927
rect 11462 1927 11526 1941
rect 11462 1877 11470 1927
rect 11470 1877 11504 1927
rect 11504 1877 11526 1927
rect 12068 1927 12132 1941
rect 12068 1877 12076 1927
rect 12076 1877 12110 1927
rect 12110 1877 12132 1927
rect 12674 1927 12738 1941
rect 12674 1877 12682 1927
rect 12682 1877 12716 1927
rect 12716 1877 12738 1927
rect 13406 1927 13470 1941
rect 13406 1877 13414 1927
rect 13414 1877 13448 1927
rect 13448 1877 13470 1927
rect 14012 1927 14076 1941
rect 14012 1877 14020 1927
rect 14020 1877 14054 1927
rect 14054 1877 14076 1927
rect 14744 1927 14808 1941
rect 14744 1877 14752 1927
rect 14752 1877 14786 1927
rect 14786 1877 14808 1927
<< metal2 >>
rect 10741 2109 10817 2110
rect 11347 2109 11423 2110
rect 11953 2109 12029 2110
rect 12559 2109 12635 2110
rect 13165 2109 13241 2110
rect 13771 2109 13847 2110
rect 14377 2109 14453 2110
rect 14983 2109 15059 2110
rect 10738 2045 10747 2109
rect 10811 2045 10820 2109
rect 10738 2036 10820 2045
rect 11344 2045 11353 2109
rect 11417 2045 11426 2109
rect 11344 2036 11426 2045
rect 11950 2045 11959 2109
rect 12023 2045 12032 2109
rect 11950 2036 12032 2045
rect 12556 2045 12565 2109
rect 12629 2045 12638 2109
rect 12556 2036 12638 2045
rect 13162 2045 13171 2109
rect 13235 2045 13244 2109
rect 13162 2036 13244 2045
rect 13768 2045 13777 2109
rect 13841 2045 13850 2109
rect 13768 2036 13850 2045
rect 14374 2045 14383 2109
rect 14447 2045 14456 2109
rect 14374 2036 14456 2045
rect 14980 2045 14989 2109
rect 15053 2045 15062 2109
rect 14980 2036 15062 2045
rect 10847 1877 10856 1941
rect 10920 1877 10929 1941
rect 10847 1876 10929 1877
rect 11453 1877 11462 1941
rect 11526 1877 11535 1941
rect 11453 1876 11535 1877
rect 12059 1877 12068 1941
rect 12132 1877 12141 1941
rect 12059 1876 12141 1877
rect 12665 1877 12674 1941
rect 12738 1877 12747 1941
rect 12665 1876 12747 1877
rect 13397 1877 13406 1941
rect 13470 1877 13479 1941
rect 13397 1876 13479 1877
rect 14003 1877 14012 1941
rect 14076 1877 14085 1941
rect 14003 1876 14085 1877
rect 14735 1877 14744 1941
rect 14808 1877 14817 1941
rect 14735 1876 14817 1877
<< via2 >>
rect 10747 2045 10811 2109
rect 11353 2045 11417 2109
rect 11959 2045 12023 2109
rect 12565 2045 12629 2109
rect 13171 2045 13235 2109
rect 13777 2045 13841 2109
rect 14383 2045 14447 2109
rect 14989 2045 15053 2109
rect 10856 1877 10920 1941
rect 11462 1877 11526 1941
rect 12068 1877 12132 1941
rect 12674 1877 12738 1941
rect 13406 1877 13470 1941
rect 14012 1877 14076 1941
rect 14744 1877 14808 1941
<< metal3 >>
rect 10502 3289 15416 3291
rect 10502 3225 10606 3289
rect 10670 3225 10686 3289
rect 10750 3225 10766 3289
rect 10830 3225 10846 3289
rect 10910 3225 10926 3289
rect 10990 3225 11006 3289
rect 11070 3225 11212 3289
rect 11276 3225 11292 3289
rect 11356 3225 11372 3289
rect 11436 3225 11452 3289
rect 11516 3225 11532 3289
rect 11596 3225 11612 3289
rect 11676 3225 11818 3289
rect 11882 3225 11898 3289
rect 11962 3225 11978 3289
rect 12042 3225 12058 3289
rect 12122 3225 12138 3289
rect 12202 3225 12218 3289
rect 12282 3225 12424 3289
rect 12488 3225 12504 3289
rect 12568 3225 12584 3289
rect 12648 3225 12664 3289
rect 12728 3225 12744 3289
rect 12808 3225 12824 3289
rect 12888 3225 13030 3289
rect 13094 3225 13110 3289
rect 13174 3225 13190 3289
rect 13254 3225 13270 3289
rect 13334 3225 13350 3289
rect 13414 3225 13430 3289
rect 13494 3225 13636 3289
rect 13700 3225 13716 3289
rect 13780 3225 13796 3289
rect 13860 3225 13876 3289
rect 13940 3225 13956 3289
rect 14020 3225 14036 3289
rect 14100 3225 14242 3289
rect 14306 3225 14322 3289
rect 14386 3225 14402 3289
rect 14466 3225 14482 3289
rect 14546 3225 14562 3289
rect 14626 3225 14642 3289
rect 14706 3225 14848 3289
rect 14912 3225 14928 3289
rect 14992 3225 15008 3289
rect 15072 3225 15088 3289
rect 15152 3225 15168 3289
rect 15232 3225 15248 3289
rect 15312 3225 15416 3289
rect 10502 3223 15416 3225
rect 10502 3069 10568 3159
rect 10502 3005 10503 3069
rect 10567 3005 10568 3069
rect 10502 2989 10568 3005
rect 10502 2925 10503 2989
rect 10567 2925 10568 2989
rect 10502 2909 10568 2925
rect 10502 2845 10503 2909
rect 10567 2845 10568 2909
rect 10502 2829 10568 2845
rect 10502 2765 10503 2829
rect 10567 2765 10568 2829
rect 10502 2749 10568 2765
rect 10502 2685 10503 2749
rect 10567 2685 10568 2749
rect 10502 2669 10568 2685
rect 10502 2605 10503 2669
rect 10567 2605 10568 2669
rect 10502 2589 10568 2605
rect 10502 2525 10503 2589
rect 10567 2525 10568 2589
rect 10502 2509 10568 2525
rect 10502 2445 10503 2509
rect 10567 2445 10568 2509
rect 10502 2429 10568 2445
rect 10502 2365 10503 2429
rect 10567 2365 10568 2429
rect 10502 2349 10568 2365
rect 10502 2285 10503 2349
rect 10567 2285 10568 2349
rect 10502 2131 10568 2285
rect 10628 2131 10688 3163
rect 10748 2193 10808 3223
rect 10868 2131 10928 3163
rect 10988 2193 11048 3223
rect 11108 3069 11174 3159
rect 11108 3005 11109 3069
rect 11173 3005 11174 3069
rect 11108 2989 11174 3005
rect 11108 2925 11109 2989
rect 11173 2925 11174 2989
rect 11108 2909 11174 2925
rect 11108 2845 11109 2909
rect 11173 2845 11174 2909
rect 11108 2829 11174 2845
rect 11108 2765 11109 2829
rect 11173 2765 11174 2829
rect 11108 2749 11174 2765
rect 11108 2685 11109 2749
rect 11173 2685 11174 2749
rect 11108 2669 11174 2685
rect 11108 2605 11109 2669
rect 11173 2605 11174 2669
rect 11108 2589 11174 2605
rect 11108 2525 11109 2589
rect 11173 2525 11174 2589
rect 11108 2509 11174 2525
rect 11108 2445 11109 2509
rect 11173 2445 11174 2509
rect 11108 2429 11174 2445
rect 11108 2365 11109 2429
rect 11173 2365 11174 2429
rect 11108 2349 11174 2365
rect 11108 2285 11109 2349
rect 11173 2285 11174 2349
rect 11108 2131 11174 2285
rect 11234 2131 11294 3163
rect 11354 2193 11414 3223
rect 11474 2131 11534 3163
rect 11594 2193 11654 3223
rect 11714 3069 11780 3159
rect 11714 3005 11715 3069
rect 11779 3005 11780 3069
rect 11714 2989 11780 3005
rect 11714 2925 11715 2989
rect 11779 2925 11780 2989
rect 11714 2909 11780 2925
rect 11714 2845 11715 2909
rect 11779 2845 11780 2909
rect 11714 2829 11780 2845
rect 11714 2765 11715 2829
rect 11779 2765 11780 2829
rect 11714 2749 11780 2765
rect 11714 2685 11715 2749
rect 11779 2685 11780 2749
rect 11714 2669 11780 2685
rect 11714 2605 11715 2669
rect 11779 2605 11780 2669
rect 11714 2589 11780 2605
rect 11714 2525 11715 2589
rect 11779 2525 11780 2589
rect 11714 2509 11780 2525
rect 11714 2445 11715 2509
rect 11779 2445 11780 2509
rect 11714 2429 11780 2445
rect 11714 2365 11715 2429
rect 11779 2365 11780 2429
rect 11714 2349 11780 2365
rect 11714 2285 11715 2349
rect 11779 2285 11780 2349
rect 11714 2131 11780 2285
rect 11840 2131 11900 3163
rect 11960 2193 12020 3223
rect 12080 2131 12140 3163
rect 12200 2193 12260 3223
rect 12320 3069 12386 3159
rect 12320 3005 12321 3069
rect 12385 3005 12386 3069
rect 12320 2989 12386 3005
rect 12320 2925 12321 2989
rect 12385 2925 12386 2989
rect 12320 2909 12386 2925
rect 12320 2845 12321 2909
rect 12385 2845 12386 2909
rect 12320 2829 12386 2845
rect 12320 2765 12321 2829
rect 12385 2765 12386 2829
rect 12320 2749 12386 2765
rect 12320 2685 12321 2749
rect 12385 2685 12386 2749
rect 12320 2669 12386 2685
rect 12320 2605 12321 2669
rect 12385 2605 12386 2669
rect 12320 2589 12386 2605
rect 12320 2525 12321 2589
rect 12385 2525 12386 2589
rect 12320 2509 12386 2525
rect 12320 2445 12321 2509
rect 12385 2445 12386 2509
rect 12320 2429 12386 2445
rect 12320 2365 12321 2429
rect 12385 2365 12386 2429
rect 12320 2349 12386 2365
rect 12320 2285 12321 2349
rect 12385 2285 12386 2349
rect 12320 2131 12386 2285
rect 12446 2131 12506 3163
rect 12566 2193 12626 3223
rect 12686 2131 12746 3163
rect 12806 2193 12866 3223
rect 12926 3069 12992 3159
rect 12926 3005 12927 3069
rect 12991 3005 12992 3069
rect 12926 2989 12992 3005
rect 12926 2925 12927 2989
rect 12991 2925 12992 2989
rect 12926 2909 12992 2925
rect 12926 2845 12927 2909
rect 12991 2845 12992 2909
rect 12926 2829 12992 2845
rect 12926 2765 12927 2829
rect 12991 2765 12992 2829
rect 12926 2749 12992 2765
rect 12926 2685 12927 2749
rect 12991 2685 12992 2749
rect 12926 2669 12992 2685
rect 12926 2605 12927 2669
rect 12991 2605 12992 2669
rect 12926 2589 12992 2605
rect 12926 2525 12927 2589
rect 12991 2525 12992 2589
rect 12926 2509 12992 2525
rect 12926 2445 12927 2509
rect 12991 2445 12992 2509
rect 12926 2429 12992 2445
rect 12926 2365 12927 2429
rect 12991 2365 12992 2429
rect 12926 2349 12992 2365
rect 12926 2285 12927 2349
rect 12991 2285 12992 2349
rect 12926 2131 12992 2285
rect 13052 2131 13112 3163
rect 13172 2193 13232 3223
rect 13292 2131 13352 3163
rect 13412 2193 13472 3223
rect 13532 3069 13598 3159
rect 13532 3005 13533 3069
rect 13597 3005 13598 3069
rect 13532 2989 13598 3005
rect 13532 2925 13533 2989
rect 13597 2925 13598 2989
rect 13532 2909 13598 2925
rect 13532 2845 13533 2909
rect 13597 2845 13598 2909
rect 13532 2829 13598 2845
rect 13532 2765 13533 2829
rect 13597 2765 13598 2829
rect 13532 2749 13598 2765
rect 13532 2685 13533 2749
rect 13597 2685 13598 2749
rect 13532 2669 13598 2685
rect 13532 2605 13533 2669
rect 13597 2605 13598 2669
rect 13532 2589 13598 2605
rect 13532 2525 13533 2589
rect 13597 2525 13598 2589
rect 13532 2509 13598 2525
rect 13532 2445 13533 2509
rect 13597 2445 13598 2509
rect 13532 2429 13598 2445
rect 13532 2365 13533 2429
rect 13597 2365 13598 2429
rect 13532 2349 13598 2365
rect 13532 2285 13533 2349
rect 13597 2285 13598 2349
rect 13532 2131 13598 2285
rect 13658 2131 13718 3163
rect 13778 2193 13838 3223
rect 13898 2131 13958 3163
rect 14018 2193 14078 3223
rect 14138 3069 14204 3159
rect 14138 3005 14139 3069
rect 14203 3005 14204 3069
rect 14138 2989 14204 3005
rect 14138 2925 14139 2989
rect 14203 2925 14204 2989
rect 14138 2909 14204 2925
rect 14138 2845 14139 2909
rect 14203 2845 14204 2909
rect 14138 2829 14204 2845
rect 14138 2765 14139 2829
rect 14203 2765 14204 2829
rect 14138 2749 14204 2765
rect 14138 2685 14139 2749
rect 14203 2685 14204 2749
rect 14138 2669 14204 2685
rect 14138 2605 14139 2669
rect 14203 2605 14204 2669
rect 14138 2589 14204 2605
rect 14138 2525 14139 2589
rect 14203 2525 14204 2589
rect 14138 2509 14204 2525
rect 14138 2445 14139 2509
rect 14203 2445 14204 2509
rect 14138 2429 14204 2445
rect 14138 2365 14139 2429
rect 14203 2365 14204 2429
rect 14138 2349 14204 2365
rect 14138 2285 14139 2349
rect 14203 2285 14204 2349
rect 14138 2131 14204 2285
rect 14264 2131 14324 3163
rect 14384 2193 14444 3223
rect 14504 2131 14564 3163
rect 14624 2193 14684 3223
rect 14744 3069 14810 3159
rect 14744 3005 14745 3069
rect 14809 3005 14810 3069
rect 14744 2989 14810 3005
rect 14744 2925 14745 2989
rect 14809 2925 14810 2989
rect 14744 2909 14810 2925
rect 14744 2845 14745 2909
rect 14809 2845 14810 2909
rect 14744 2829 14810 2845
rect 14744 2765 14745 2829
rect 14809 2765 14810 2829
rect 14744 2749 14810 2765
rect 14744 2685 14745 2749
rect 14809 2685 14810 2749
rect 14744 2669 14810 2685
rect 14744 2605 14745 2669
rect 14809 2605 14810 2669
rect 14744 2589 14810 2605
rect 14744 2525 14745 2589
rect 14809 2525 14810 2589
rect 14744 2509 14810 2525
rect 14744 2445 14745 2509
rect 14809 2445 14810 2509
rect 14744 2429 14810 2445
rect 14744 2365 14745 2429
rect 14809 2365 14810 2429
rect 14744 2349 14810 2365
rect 14744 2285 14745 2349
rect 14809 2285 14810 2349
rect 14744 2131 14810 2285
rect 14870 2131 14930 3163
rect 14990 2193 15050 3223
rect 15110 2131 15170 3163
rect 15230 2193 15290 3223
rect 15350 3069 15416 3159
rect 15350 3005 15351 3069
rect 15415 3005 15416 3069
rect 15350 2989 15416 3005
rect 15350 2925 15351 2989
rect 15415 2925 15416 2989
rect 15350 2909 15416 2925
rect 15350 2845 15351 2909
rect 15415 2845 15416 2909
rect 15350 2829 15416 2845
rect 15350 2765 15351 2829
rect 15415 2765 15416 2829
rect 15350 2749 15416 2765
rect 15350 2685 15351 2749
rect 15415 2685 15416 2749
rect 15350 2669 15416 2685
rect 15350 2605 15351 2669
rect 15415 2605 15416 2669
rect 15350 2589 15416 2605
rect 15350 2525 15351 2589
rect 15415 2525 15416 2589
rect 15350 2509 15416 2525
rect 15350 2445 15351 2509
rect 15415 2445 15416 2509
rect 15350 2429 15416 2445
rect 15350 2365 15351 2429
rect 15415 2365 15416 2429
rect 15350 2349 15416 2365
rect 15350 2285 15351 2349
rect 15415 2285 15416 2349
rect 15350 2131 15416 2285
rect 10502 2129 15416 2131
rect 10502 2065 10606 2129
rect 10670 2065 10686 2129
rect 10750 2109 10766 2129
rect 10830 2065 10846 2129
rect 10910 2065 10926 2129
rect 10990 2065 11006 2129
rect 11070 2065 11212 2129
rect 11276 2065 11292 2129
rect 11356 2109 11372 2129
rect 11436 2065 11452 2129
rect 11516 2065 11532 2129
rect 11596 2065 11612 2129
rect 11676 2065 11818 2129
rect 11882 2065 11898 2129
rect 11962 2109 11978 2129
rect 12042 2065 12058 2129
rect 12122 2065 12138 2129
rect 12202 2065 12218 2129
rect 12282 2065 12424 2129
rect 12488 2065 12504 2129
rect 12568 2109 12584 2129
rect 12648 2065 12664 2129
rect 12728 2065 12744 2129
rect 12808 2065 12824 2129
rect 12888 2065 13030 2129
rect 13094 2065 13110 2129
rect 13174 2109 13190 2129
rect 13254 2065 13270 2129
rect 13334 2065 13350 2129
rect 13414 2065 13430 2129
rect 13494 2065 13636 2129
rect 13700 2065 13716 2129
rect 13780 2109 13796 2129
rect 13860 2065 13876 2129
rect 13940 2065 13956 2129
rect 14020 2065 14036 2129
rect 14100 2065 14242 2129
rect 14306 2065 14322 2129
rect 14386 2109 14402 2129
rect 14466 2065 14482 2129
rect 14546 2065 14562 2129
rect 14626 2065 14642 2129
rect 14706 2065 14848 2129
rect 14912 2065 14928 2129
rect 14992 2109 15008 2129
rect 15072 2065 15088 2129
rect 15152 2065 15168 2129
rect 15232 2065 15248 2129
rect 15312 2065 15416 2129
rect 10502 2063 10747 2065
rect 10738 2045 10747 2063
rect 10811 2063 11353 2065
rect 10811 2045 10820 2063
rect 10738 2036 10820 2045
rect 11344 2045 11353 2063
rect 11417 2063 11959 2065
rect 11417 2045 11426 2063
rect 11344 2036 11426 2045
rect 11950 2045 11959 2063
rect 12023 2063 12565 2065
rect 12023 2045 12032 2063
rect 11950 2036 12032 2045
rect 12556 2045 12565 2063
rect 12629 2063 13171 2065
rect 12629 2045 12638 2063
rect 12556 2036 12638 2045
rect 13162 2045 13171 2063
rect 13235 2063 13777 2065
rect 13235 2045 13244 2063
rect 13162 2036 13244 2045
rect 13768 2045 13777 2063
rect 13841 2063 14383 2065
rect 13841 2045 13850 2063
rect 13768 2036 13850 2045
rect 14374 2045 14383 2063
rect 14447 2063 14989 2065
rect 14447 2045 14456 2063
rect 14374 2036 14456 2045
rect 14980 2045 14989 2063
rect 15053 2063 15416 2065
rect 15053 2045 15062 2063
rect 14980 2036 15062 2045
rect 10847 1941 10929 1948
rect 10847 1929 10856 1941
rect 10502 1927 10856 1929
rect 10920 1929 10929 1941
rect 11453 1941 11535 1948
rect 11453 1929 11462 1941
rect 10920 1927 11462 1929
rect 11526 1929 11535 1941
rect 12059 1941 12141 1948
rect 12059 1929 12068 1941
rect 11526 1927 12068 1929
rect 12132 1929 12141 1941
rect 12665 1941 12747 1948
rect 12665 1929 12674 1941
rect 12132 1927 12674 1929
rect 12738 1929 12747 1941
rect 13397 1941 13479 1948
rect 13397 1929 13406 1941
rect 12738 1927 12992 1929
rect 10502 1863 10606 1927
rect 10670 1863 10686 1927
rect 10750 1863 10766 1927
rect 10830 1863 10846 1927
rect 10920 1877 10926 1927
rect 10910 1863 10926 1877
rect 10990 1863 11006 1927
rect 11070 1863 11212 1927
rect 11276 1863 11292 1927
rect 11356 1863 11372 1927
rect 11436 1863 11452 1927
rect 11526 1877 11532 1927
rect 11516 1863 11532 1877
rect 11596 1863 11612 1927
rect 11676 1863 11818 1927
rect 11882 1863 11898 1927
rect 11962 1863 11978 1927
rect 12042 1863 12058 1927
rect 12132 1877 12138 1927
rect 12122 1863 12138 1877
rect 12202 1863 12218 1927
rect 12282 1863 12424 1927
rect 12488 1863 12504 1927
rect 12568 1863 12584 1927
rect 12648 1863 12664 1927
rect 12738 1877 12744 1927
rect 12728 1863 12744 1877
rect 12808 1863 12824 1927
rect 12888 1863 12992 1927
rect 10502 1861 12992 1863
rect 10502 1707 10568 1861
rect 10502 1643 10503 1707
rect 10567 1643 10568 1707
rect 10502 1627 10568 1643
rect 10502 1563 10503 1627
rect 10567 1563 10568 1627
rect 10502 1547 10568 1563
rect 10502 1483 10503 1547
rect 10567 1483 10568 1547
rect 10502 1467 10568 1483
rect 10502 1403 10503 1467
rect 10567 1403 10568 1467
rect 10502 1387 10568 1403
rect 10502 1323 10503 1387
rect 10567 1323 10568 1387
rect 10502 1307 10568 1323
rect 10502 1243 10503 1307
rect 10567 1243 10568 1307
rect 10502 1227 10568 1243
rect 10502 1163 10503 1227
rect 10567 1163 10568 1227
rect 10502 1147 10568 1163
rect 10502 1083 10503 1147
rect 10567 1083 10568 1147
rect 10502 1067 10568 1083
rect 10502 1003 10503 1067
rect 10567 1003 10568 1067
rect 10502 987 10568 1003
rect 10502 923 10503 987
rect 10567 923 10568 987
rect 10502 833 10568 923
rect 10628 769 10688 1799
rect 10748 829 10808 1861
rect 10868 769 10928 1799
rect 10988 829 11048 1861
rect 11108 1707 11174 1861
rect 11108 1643 11109 1707
rect 11173 1643 11174 1707
rect 11108 1627 11174 1643
rect 11108 1563 11109 1627
rect 11173 1563 11174 1627
rect 11108 1547 11174 1563
rect 11108 1483 11109 1547
rect 11173 1483 11174 1547
rect 11108 1467 11174 1483
rect 11108 1403 11109 1467
rect 11173 1403 11174 1467
rect 11108 1387 11174 1403
rect 11108 1323 11109 1387
rect 11173 1323 11174 1387
rect 11108 1307 11174 1323
rect 11108 1243 11109 1307
rect 11173 1243 11174 1307
rect 11108 1227 11174 1243
rect 11108 1163 11109 1227
rect 11173 1163 11174 1227
rect 11108 1147 11174 1163
rect 11108 1083 11109 1147
rect 11173 1083 11174 1147
rect 11108 1067 11174 1083
rect 11108 1003 11109 1067
rect 11173 1003 11174 1067
rect 11108 987 11174 1003
rect 11108 923 11109 987
rect 11173 923 11174 987
rect 11108 833 11174 923
rect 11234 769 11294 1799
rect 11354 829 11414 1861
rect 11474 769 11534 1799
rect 11594 829 11654 1861
rect 11714 1707 11780 1861
rect 11714 1643 11715 1707
rect 11779 1643 11780 1707
rect 11714 1627 11780 1643
rect 11714 1563 11715 1627
rect 11779 1563 11780 1627
rect 11714 1547 11780 1563
rect 11714 1483 11715 1547
rect 11779 1483 11780 1547
rect 11714 1467 11780 1483
rect 11714 1403 11715 1467
rect 11779 1403 11780 1467
rect 11714 1387 11780 1403
rect 11714 1323 11715 1387
rect 11779 1323 11780 1387
rect 11714 1307 11780 1323
rect 11714 1243 11715 1307
rect 11779 1243 11780 1307
rect 11714 1227 11780 1243
rect 11714 1163 11715 1227
rect 11779 1163 11780 1227
rect 11714 1147 11780 1163
rect 11714 1083 11715 1147
rect 11779 1083 11780 1147
rect 11714 1067 11780 1083
rect 11714 1003 11715 1067
rect 11779 1003 11780 1067
rect 11714 987 11780 1003
rect 11714 923 11715 987
rect 11779 923 11780 987
rect 11714 833 11780 923
rect 11840 769 11900 1799
rect 11960 829 12020 1861
rect 12080 769 12140 1799
rect 12200 829 12260 1861
rect 12320 1707 12386 1861
rect 12320 1643 12321 1707
rect 12385 1643 12386 1707
rect 12320 1627 12386 1643
rect 12320 1563 12321 1627
rect 12385 1563 12386 1627
rect 12320 1547 12386 1563
rect 12320 1483 12321 1547
rect 12385 1483 12386 1547
rect 12320 1467 12386 1483
rect 12320 1403 12321 1467
rect 12385 1403 12386 1467
rect 12320 1387 12386 1403
rect 12320 1323 12321 1387
rect 12385 1323 12386 1387
rect 12320 1307 12386 1323
rect 12320 1243 12321 1307
rect 12385 1243 12386 1307
rect 12320 1227 12386 1243
rect 12320 1163 12321 1227
rect 12385 1163 12386 1227
rect 12320 1147 12386 1163
rect 12320 1083 12321 1147
rect 12385 1083 12386 1147
rect 12320 1067 12386 1083
rect 12320 1003 12321 1067
rect 12385 1003 12386 1067
rect 12320 987 12386 1003
rect 12320 923 12321 987
rect 12385 923 12386 987
rect 12320 833 12386 923
rect 12446 769 12506 1799
rect 12566 829 12626 1861
rect 12686 769 12746 1799
rect 12806 829 12866 1861
rect 12926 1707 12992 1861
rect 12926 1643 12927 1707
rect 12991 1643 12992 1707
rect 12926 1627 12992 1643
rect 12926 1563 12927 1627
rect 12991 1563 12992 1627
rect 12926 1547 12992 1563
rect 12926 1483 12927 1547
rect 12991 1483 12992 1547
rect 12926 1467 12992 1483
rect 12926 1403 12927 1467
rect 12991 1403 12992 1467
rect 12926 1387 12992 1403
rect 12926 1323 12927 1387
rect 12991 1323 12992 1387
rect 12926 1307 12992 1323
rect 12926 1243 12927 1307
rect 12991 1243 12992 1307
rect 12926 1227 12992 1243
rect 12926 1163 12927 1227
rect 12991 1163 12992 1227
rect 12926 1147 12992 1163
rect 12926 1083 12927 1147
rect 12991 1083 12992 1147
rect 12926 1067 12992 1083
rect 12926 1003 12927 1067
rect 12991 1003 12992 1067
rect 12926 987 12992 1003
rect 12926 923 12927 987
rect 12991 923 12992 987
rect 12926 833 12992 923
rect 13052 1927 13406 1929
rect 13470 1929 13479 1941
rect 14003 1941 14085 1948
rect 14003 1929 14012 1941
rect 13470 1927 14012 1929
rect 14076 1929 14085 1941
rect 14735 1941 14817 1948
rect 14735 1929 14744 1941
rect 14076 1927 14330 1929
rect 13052 1863 13156 1927
rect 13220 1863 13236 1927
rect 13300 1863 13316 1927
rect 13380 1863 13396 1927
rect 13470 1877 13476 1927
rect 13460 1863 13476 1877
rect 13540 1863 13556 1927
rect 13620 1863 13762 1927
rect 13826 1863 13842 1927
rect 13906 1863 13922 1927
rect 13986 1863 14002 1927
rect 14076 1877 14082 1927
rect 14066 1863 14082 1877
rect 14146 1863 14162 1927
rect 14226 1863 14330 1927
rect 13052 1861 14330 1863
rect 13052 1707 13118 1861
rect 13052 1643 13053 1707
rect 13117 1643 13118 1707
rect 13052 1627 13118 1643
rect 13052 1563 13053 1627
rect 13117 1563 13118 1627
rect 13052 1547 13118 1563
rect 13052 1483 13053 1547
rect 13117 1483 13118 1547
rect 13052 1467 13118 1483
rect 13052 1403 13053 1467
rect 13117 1403 13118 1467
rect 13052 1387 13118 1403
rect 13052 1323 13053 1387
rect 13117 1323 13118 1387
rect 13052 1307 13118 1323
rect 13052 1243 13053 1307
rect 13117 1243 13118 1307
rect 13052 1227 13118 1243
rect 13052 1163 13053 1227
rect 13117 1163 13118 1227
rect 13052 1147 13118 1163
rect 13052 1083 13053 1147
rect 13117 1083 13118 1147
rect 13052 1067 13118 1083
rect 13052 1003 13053 1067
rect 13117 1003 13118 1067
rect 13052 987 13118 1003
rect 13052 923 13053 987
rect 13117 923 13118 987
rect 13052 833 13118 923
rect 13178 769 13238 1799
rect 13298 829 13358 1861
rect 13418 769 13478 1799
rect 13538 829 13598 1861
rect 13658 1707 13724 1861
rect 13658 1643 13659 1707
rect 13723 1643 13724 1707
rect 13658 1627 13724 1643
rect 13658 1563 13659 1627
rect 13723 1563 13724 1627
rect 13658 1547 13724 1563
rect 13658 1483 13659 1547
rect 13723 1483 13724 1547
rect 13658 1467 13724 1483
rect 13658 1403 13659 1467
rect 13723 1403 13724 1467
rect 13658 1387 13724 1403
rect 13658 1323 13659 1387
rect 13723 1323 13724 1387
rect 13658 1307 13724 1323
rect 13658 1243 13659 1307
rect 13723 1243 13724 1307
rect 13658 1227 13724 1243
rect 13658 1163 13659 1227
rect 13723 1163 13724 1227
rect 13658 1147 13724 1163
rect 13658 1083 13659 1147
rect 13723 1083 13724 1147
rect 13658 1067 13724 1083
rect 13658 1003 13659 1067
rect 13723 1003 13724 1067
rect 13658 987 13724 1003
rect 13658 923 13659 987
rect 13723 923 13724 987
rect 13658 833 13724 923
rect 13784 769 13844 1799
rect 13904 829 13964 1861
rect 14024 769 14084 1799
rect 14144 829 14204 1861
rect 14264 1707 14330 1861
rect 14264 1643 14265 1707
rect 14329 1643 14330 1707
rect 14264 1627 14330 1643
rect 14264 1563 14265 1627
rect 14329 1563 14330 1627
rect 14264 1547 14330 1563
rect 14264 1483 14265 1547
rect 14329 1483 14330 1547
rect 14264 1467 14330 1483
rect 14264 1403 14265 1467
rect 14329 1403 14330 1467
rect 14264 1387 14330 1403
rect 14264 1323 14265 1387
rect 14329 1323 14330 1387
rect 14264 1307 14330 1323
rect 14264 1243 14265 1307
rect 14329 1243 14330 1307
rect 14264 1227 14330 1243
rect 14264 1163 14265 1227
rect 14329 1163 14330 1227
rect 14264 1147 14330 1163
rect 14264 1083 14265 1147
rect 14329 1083 14330 1147
rect 14264 1067 14330 1083
rect 14264 1003 14265 1067
rect 14329 1003 14330 1067
rect 14264 987 14330 1003
rect 14264 923 14265 987
rect 14329 923 14330 987
rect 14264 833 14330 923
rect 14390 1927 14744 1929
rect 14808 1929 14817 1941
rect 14808 1927 15062 1929
rect 14390 1863 14494 1927
rect 14558 1863 14574 1927
rect 14638 1863 14654 1927
rect 14718 1863 14734 1927
rect 14808 1877 14814 1927
rect 14798 1863 14814 1877
rect 14878 1863 14894 1927
rect 14958 1863 15062 1927
rect 14390 1861 15062 1863
rect 14390 1707 14456 1861
rect 14390 1643 14391 1707
rect 14455 1643 14456 1707
rect 14390 1627 14456 1643
rect 14390 1563 14391 1627
rect 14455 1563 14456 1627
rect 14390 1547 14456 1563
rect 14390 1483 14391 1547
rect 14455 1483 14456 1547
rect 14390 1467 14456 1483
rect 14390 1403 14391 1467
rect 14455 1403 14456 1467
rect 14390 1387 14456 1403
rect 14390 1323 14391 1387
rect 14455 1323 14456 1387
rect 14390 1307 14456 1323
rect 14390 1243 14391 1307
rect 14455 1243 14456 1307
rect 14390 1227 14456 1243
rect 14390 1163 14391 1227
rect 14455 1163 14456 1227
rect 14390 1147 14456 1163
rect 14390 1083 14391 1147
rect 14455 1083 14456 1147
rect 14390 1067 14456 1083
rect 14390 1003 14391 1067
rect 14455 1003 14456 1067
rect 14390 987 14456 1003
rect 14390 923 14391 987
rect 14455 923 14456 987
rect 14390 833 14456 923
rect 14516 769 14576 1799
rect 14636 829 14696 1861
rect 14756 769 14816 1799
rect 14876 829 14936 1861
rect 14996 1707 15062 1861
rect 14996 1643 14997 1707
rect 15061 1643 15062 1707
rect 14996 1627 15062 1643
rect 14996 1563 14997 1627
rect 15061 1563 15062 1627
rect 14996 1547 15062 1563
rect 14996 1483 14997 1547
rect 15061 1483 15062 1547
rect 14996 1467 15062 1483
rect 14996 1403 14997 1467
rect 15061 1403 15062 1467
rect 14996 1387 15062 1403
rect 14996 1323 14997 1387
rect 15061 1323 15062 1387
rect 14996 1307 15062 1323
rect 14996 1243 14997 1307
rect 15061 1243 15062 1307
rect 14996 1227 15062 1243
rect 14996 1163 14997 1227
rect 15061 1163 15062 1227
rect 14996 1147 15062 1163
rect 14996 1083 14997 1147
rect 15061 1083 15062 1147
rect 14996 1067 15062 1083
rect 14996 1003 14997 1067
rect 15061 1003 15062 1067
rect 14996 987 15062 1003
rect 14996 923 14997 987
rect 15061 923 15062 987
rect 14996 833 15062 923
rect 10502 767 12992 769
rect 10502 703 10606 767
rect 10670 703 10686 767
rect 10750 703 10766 767
rect 10830 703 10846 767
rect 10910 703 10926 767
rect 10990 703 11006 767
rect 11070 703 11212 767
rect 11276 703 11292 767
rect 11356 703 11372 767
rect 11436 703 11452 767
rect 11516 703 11532 767
rect 11596 703 11612 767
rect 11676 703 11818 767
rect 11882 703 11898 767
rect 11962 703 11978 767
rect 12042 703 12058 767
rect 12122 703 12138 767
rect 12202 703 12218 767
rect 12282 703 12424 767
rect 12488 703 12504 767
rect 12568 703 12584 767
rect 12648 703 12664 767
rect 12728 703 12744 767
rect 12808 703 12824 767
rect 12888 703 12992 767
rect 10502 701 12992 703
rect 13052 767 14330 769
rect 13052 703 13156 767
rect 13220 703 13236 767
rect 13300 703 13316 767
rect 13380 703 13396 767
rect 13460 703 13476 767
rect 13540 703 13556 767
rect 13620 703 13762 767
rect 13826 703 13842 767
rect 13906 703 13922 767
rect 13986 703 14002 767
rect 14066 703 14082 767
rect 14146 703 14162 767
rect 14226 703 14330 767
rect 13052 701 14330 703
rect 14390 767 15062 769
rect 14390 703 14494 767
rect 14558 703 14574 767
rect 14638 703 14654 767
rect 14718 703 14734 767
rect 14798 703 14814 767
rect 14878 703 14894 767
rect 14958 703 15062 767
rect 14390 701 15062 703
<< via3 >>
rect 10606 3225 10670 3289
rect 10686 3225 10750 3289
rect 10766 3225 10830 3289
rect 10846 3225 10910 3289
rect 10926 3225 10990 3289
rect 11006 3225 11070 3289
rect 11212 3225 11276 3289
rect 11292 3225 11356 3289
rect 11372 3225 11436 3289
rect 11452 3225 11516 3289
rect 11532 3225 11596 3289
rect 11612 3225 11676 3289
rect 11818 3225 11882 3289
rect 11898 3225 11962 3289
rect 11978 3225 12042 3289
rect 12058 3225 12122 3289
rect 12138 3225 12202 3289
rect 12218 3225 12282 3289
rect 12424 3225 12488 3289
rect 12504 3225 12568 3289
rect 12584 3225 12648 3289
rect 12664 3225 12728 3289
rect 12744 3225 12808 3289
rect 12824 3225 12888 3289
rect 13030 3225 13094 3289
rect 13110 3225 13174 3289
rect 13190 3225 13254 3289
rect 13270 3225 13334 3289
rect 13350 3225 13414 3289
rect 13430 3225 13494 3289
rect 13636 3225 13700 3289
rect 13716 3225 13780 3289
rect 13796 3225 13860 3289
rect 13876 3225 13940 3289
rect 13956 3225 14020 3289
rect 14036 3225 14100 3289
rect 14242 3225 14306 3289
rect 14322 3225 14386 3289
rect 14402 3225 14466 3289
rect 14482 3225 14546 3289
rect 14562 3225 14626 3289
rect 14642 3225 14706 3289
rect 14848 3225 14912 3289
rect 14928 3225 14992 3289
rect 15008 3225 15072 3289
rect 15088 3225 15152 3289
rect 15168 3225 15232 3289
rect 15248 3225 15312 3289
rect 10503 3005 10567 3069
rect 10503 2925 10567 2989
rect 10503 2845 10567 2909
rect 10503 2765 10567 2829
rect 10503 2685 10567 2749
rect 10503 2605 10567 2669
rect 10503 2525 10567 2589
rect 10503 2445 10567 2509
rect 10503 2365 10567 2429
rect 10503 2285 10567 2349
rect 11109 3005 11173 3069
rect 11109 2925 11173 2989
rect 11109 2845 11173 2909
rect 11109 2765 11173 2829
rect 11109 2685 11173 2749
rect 11109 2605 11173 2669
rect 11109 2525 11173 2589
rect 11109 2445 11173 2509
rect 11109 2365 11173 2429
rect 11109 2285 11173 2349
rect 11715 3005 11779 3069
rect 11715 2925 11779 2989
rect 11715 2845 11779 2909
rect 11715 2765 11779 2829
rect 11715 2685 11779 2749
rect 11715 2605 11779 2669
rect 11715 2525 11779 2589
rect 11715 2445 11779 2509
rect 11715 2365 11779 2429
rect 11715 2285 11779 2349
rect 12321 3005 12385 3069
rect 12321 2925 12385 2989
rect 12321 2845 12385 2909
rect 12321 2765 12385 2829
rect 12321 2685 12385 2749
rect 12321 2605 12385 2669
rect 12321 2525 12385 2589
rect 12321 2445 12385 2509
rect 12321 2365 12385 2429
rect 12321 2285 12385 2349
rect 12927 3005 12991 3069
rect 12927 2925 12991 2989
rect 12927 2845 12991 2909
rect 12927 2765 12991 2829
rect 12927 2685 12991 2749
rect 12927 2605 12991 2669
rect 12927 2525 12991 2589
rect 12927 2445 12991 2509
rect 12927 2365 12991 2429
rect 12927 2285 12991 2349
rect 13533 3005 13597 3069
rect 13533 2925 13597 2989
rect 13533 2845 13597 2909
rect 13533 2765 13597 2829
rect 13533 2685 13597 2749
rect 13533 2605 13597 2669
rect 13533 2525 13597 2589
rect 13533 2445 13597 2509
rect 13533 2365 13597 2429
rect 13533 2285 13597 2349
rect 14139 3005 14203 3069
rect 14139 2925 14203 2989
rect 14139 2845 14203 2909
rect 14139 2765 14203 2829
rect 14139 2685 14203 2749
rect 14139 2605 14203 2669
rect 14139 2525 14203 2589
rect 14139 2445 14203 2509
rect 14139 2365 14203 2429
rect 14139 2285 14203 2349
rect 14745 3005 14809 3069
rect 14745 2925 14809 2989
rect 14745 2845 14809 2909
rect 14745 2765 14809 2829
rect 14745 2685 14809 2749
rect 14745 2605 14809 2669
rect 14745 2525 14809 2589
rect 14745 2445 14809 2509
rect 14745 2365 14809 2429
rect 14745 2285 14809 2349
rect 15351 3005 15415 3069
rect 15351 2925 15415 2989
rect 15351 2845 15415 2909
rect 15351 2765 15415 2829
rect 15351 2685 15415 2749
rect 15351 2605 15415 2669
rect 15351 2525 15415 2589
rect 15351 2445 15415 2509
rect 15351 2365 15415 2429
rect 15351 2285 15415 2349
rect 10606 2065 10670 2129
rect 10686 2109 10750 2129
rect 10766 2109 10830 2129
rect 10686 2065 10747 2109
rect 10747 2065 10750 2109
rect 10766 2065 10811 2109
rect 10811 2065 10830 2109
rect 10846 2065 10910 2129
rect 10926 2065 10990 2129
rect 11006 2065 11070 2129
rect 11212 2065 11276 2129
rect 11292 2109 11356 2129
rect 11372 2109 11436 2129
rect 11292 2065 11353 2109
rect 11353 2065 11356 2109
rect 11372 2065 11417 2109
rect 11417 2065 11436 2109
rect 11452 2065 11516 2129
rect 11532 2065 11596 2129
rect 11612 2065 11676 2129
rect 11818 2065 11882 2129
rect 11898 2109 11962 2129
rect 11978 2109 12042 2129
rect 11898 2065 11959 2109
rect 11959 2065 11962 2109
rect 11978 2065 12023 2109
rect 12023 2065 12042 2109
rect 12058 2065 12122 2129
rect 12138 2065 12202 2129
rect 12218 2065 12282 2129
rect 12424 2065 12488 2129
rect 12504 2109 12568 2129
rect 12584 2109 12648 2129
rect 12504 2065 12565 2109
rect 12565 2065 12568 2109
rect 12584 2065 12629 2109
rect 12629 2065 12648 2109
rect 12664 2065 12728 2129
rect 12744 2065 12808 2129
rect 12824 2065 12888 2129
rect 13030 2065 13094 2129
rect 13110 2109 13174 2129
rect 13190 2109 13254 2129
rect 13110 2065 13171 2109
rect 13171 2065 13174 2109
rect 13190 2065 13235 2109
rect 13235 2065 13254 2109
rect 13270 2065 13334 2129
rect 13350 2065 13414 2129
rect 13430 2065 13494 2129
rect 13636 2065 13700 2129
rect 13716 2109 13780 2129
rect 13796 2109 13860 2129
rect 13716 2065 13777 2109
rect 13777 2065 13780 2109
rect 13796 2065 13841 2109
rect 13841 2065 13860 2109
rect 13876 2065 13940 2129
rect 13956 2065 14020 2129
rect 14036 2065 14100 2129
rect 14242 2065 14306 2129
rect 14322 2109 14386 2129
rect 14402 2109 14466 2129
rect 14322 2065 14383 2109
rect 14383 2065 14386 2109
rect 14402 2065 14447 2109
rect 14447 2065 14466 2109
rect 14482 2065 14546 2129
rect 14562 2065 14626 2129
rect 14642 2065 14706 2129
rect 14848 2065 14912 2129
rect 14928 2109 14992 2129
rect 15008 2109 15072 2129
rect 14928 2065 14989 2109
rect 14989 2065 14992 2109
rect 15008 2065 15053 2109
rect 15053 2065 15072 2109
rect 15088 2065 15152 2129
rect 15168 2065 15232 2129
rect 15248 2065 15312 2129
rect 10606 1863 10670 1927
rect 10686 1863 10750 1927
rect 10766 1863 10830 1927
rect 10846 1877 10856 1927
rect 10856 1877 10910 1927
rect 10846 1863 10910 1877
rect 10926 1863 10990 1927
rect 11006 1863 11070 1927
rect 11212 1863 11276 1927
rect 11292 1863 11356 1927
rect 11372 1863 11436 1927
rect 11452 1877 11462 1927
rect 11462 1877 11516 1927
rect 11452 1863 11516 1877
rect 11532 1863 11596 1927
rect 11612 1863 11676 1927
rect 11818 1863 11882 1927
rect 11898 1863 11962 1927
rect 11978 1863 12042 1927
rect 12058 1877 12068 1927
rect 12068 1877 12122 1927
rect 12058 1863 12122 1877
rect 12138 1863 12202 1927
rect 12218 1863 12282 1927
rect 12424 1863 12488 1927
rect 12504 1863 12568 1927
rect 12584 1863 12648 1927
rect 12664 1877 12674 1927
rect 12674 1877 12728 1927
rect 12664 1863 12728 1877
rect 12744 1863 12808 1927
rect 12824 1863 12888 1927
rect 10503 1643 10567 1707
rect 10503 1563 10567 1627
rect 10503 1483 10567 1547
rect 10503 1403 10567 1467
rect 10503 1323 10567 1387
rect 10503 1243 10567 1307
rect 10503 1163 10567 1227
rect 10503 1083 10567 1147
rect 10503 1003 10567 1067
rect 10503 923 10567 987
rect 11109 1643 11173 1707
rect 11109 1563 11173 1627
rect 11109 1483 11173 1547
rect 11109 1403 11173 1467
rect 11109 1323 11173 1387
rect 11109 1243 11173 1307
rect 11109 1163 11173 1227
rect 11109 1083 11173 1147
rect 11109 1003 11173 1067
rect 11109 923 11173 987
rect 11715 1643 11779 1707
rect 11715 1563 11779 1627
rect 11715 1483 11779 1547
rect 11715 1403 11779 1467
rect 11715 1323 11779 1387
rect 11715 1243 11779 1307
rect 11715 1163 11779 1227
rect 11715 1083 11779 1147
rect 11715 1003 11779 1067
rect 11715 923 11779 987
rect 12321 1643 12385 1707
rect 12321 1563 12385 1627
rect 12321 1483 12385 1547
rect 12321 1403 12385 1467
rect 12321 1323 12385 1387
rect 12321 1243 12385 1307
rect 12321 1163 12385 1227
rect 12321 1083 12385 1147
rect 12321 1003 12385 1067
rect 12321 923 12385 987
rect 12927 1643 12991 1707
rect 12927 1563 12991 1627
rect 12927 1483 12991 1547
rect 12927 1403 12991 1467
rect 12927 1323 12991 1387
rect 12927 1243 12991 1307
rect 12927 1163 12991 1227
rect 12927 1083 12991 1147
rect 12927 1003 12991 1067
rect 12927 923 12991 987
rect 13156 1863 13220 1927
rect 13236 1863 13300 1927
rect 13316 1863 13380 1927
rect 13396 1877 13406 1927
rect 13406 1877 13460 1927
rect 13396 1863 13460 1877
rect 13476 1863 13540 1927
rect 13556 1863 13620 1927
rect 13762 1863 13826 1927
rect 13842 1863 13906 1927
rect 13922 1863 13986 1927
rect 14002 1877 14012 1927
rect 14012 1877 14066 1927
rect 14002 1863 14066 1877
rect 14082 1863 14146 1927
rect 14162 1863 14226 1927
rect 13053 1643 13117 1707
rect 13053 1563 13117 1627
rect 13053 1483 13117 1547
rect 13053 1403 13117 1467
rect 13053 1323 13117 1387
rect 13053 1243 13117 1307
rect 13053 1163 13117 1227
rect 13053 1083 13117 1147
rect 13053 1003 13117 1067
rect 13053 923 13117 987
rect 13659 1643 13723 1707
rect 13659 1563 13723 1627
rect 13659 1483 13723 1547
rect 13659 1403 13723 1467
rect 13659 1323 13723 1387
rect 13659 1243 13723 1307
rect 13659 1163 13723 1227
rect 13659 1083 13723 1147
rect 13659 1003 13723 1067
rect 13659 923 13723 987
rect 14265 1643 14329 1707
rect 14265 1563 14329 1627
rect 14265 1483 14329 1547
rect 14265 1403 14329 1467
rect 14265 1323 14329 1387
rect 14265 1243 14329 1307
rect 14265 1163 14329 1227
rect 14265 1083 14329 1147
rect 14265 1003 14329 1067
rect 14265 923 14329 987
rect 14494 1863 14558 1927
rect 14574 1863 14638 1927
rect 14654 1863 14718 1927
rect 14734 1877 14744 1927
rect 14744 1877 14798 1927
rect 14734 1863 14798 1877
rect 14814 1863 14878 1927
rect 14894 1863 14958 1927
rect 14391 1643 14455 1707
rect 14391 1563 14455 1627
rect 14391 1483 14455 1547
rect 14391 1403 14455 1467
rect 14391 1323 14455 1387
rect 14391 1243 14455 1307
rect 14391 1163 14455 1227
rect 14391 1083 14455 1147
rect 14391 1003 14455 1067
rect 14391 923 14455 987
rect 14997 1643 15061 1707
rect 14997 1563 15061 1627
rect 14997 1483 15061 1547
rect 14997 1403 15061 1467
rect 14997 1323 15061 1387
rect 14997 1243 15061 1307
rect 14997 1163 15061 1227
rect 14997 1083 15061 1147
rect 14997 1003 15061 1067
rect 14997 923 15061 987
rect 10606 703 10670 767
rect 10686 703 10750 767
rect 10766 703 10830 767
rect 10846 703 10910 767
rect 10926 703 10990 767
rect 11006 703 11070 767
rect 11212 703 11276 767
rect 11292 703 11356 767
rect 11372 703 11436 767
rect 11452 703 11516 767
rect 11532 703 11596 767
rect 11612 703 11676 767
rect 11818 703 11882 767
rect 11898 703 11962 767
rect 11978 703 12042 767
rect 12058 703 12122 767
rect 12138 703 12202 767
rect 12218 703 12282 767
rect 12424 703 12488 767
rect 12504 703 12568 767
rect 12584 703 12648 767
rect 12664 703 12728 767
rect 12744 703 12808 767
rect 12824 703 12888 767
rect 13156 703 13220 767
rect 13236 703 13300 767
rect 13316 703 13380 767
rect 13396 703 13460 767
rect 13476 703 13540 767
rect 13556 703 13620 767
rect 13762 703 13826 767
rect 13842 703 13906 767
rect 13922 703 13986 767
rect 14002 703 14066 767
rect 14082 703 14146 767
rect 14162 703 14226 767
rect 14494 703 14558 767
rect 14574 703 14638 767
rect 14654 703 14718 767
rect 14734 703 14798 767
rect 14814 703 14878 767
rect 14894 703 14958 767
<< metal4 >>
rect 10231 3351 15964 3486
rect 10231 2312 10442 3351
rect 10502 3289 15416 3291
rect 10502 3225 10606 3289
rect 10670 3225 10686 3289
rect 10750 3225 10766 3289
rect 10830 3225 10846 3289
rect 10910 3225 10926 3289
rect 10990 3225 11006 3289
rect 11070 3225 11212 3289
rect 11276 3225 11292 3289
rect 11356 3225 11372 3289
rect 11436 3225 11452 3289
rect 11516 3225 11532 3289
rect 11596 3225 11612 3289
rect 11676 3225 11818 3289
rect 11882 3225 11898 3289
rect 11962 3225 11978 3289
rect 12042 3225 12058 3289
rect 12122 3225 12138 3289
rect 12202 3225 12218 3289
rect 12282 3225 12424 3289
rect 12488 3225 12504 3289
rect 12568 3225 12584 3289
rect 12648 3225 12664 3289
rect 12728 3225 12744 3289
rect 12808 3225 12824 3289
rect 12888 3225 13030 3289
rect 13094 3225 13110 3289
rect 13174 3225 13190 3289
rect 13254 3225 13270 3289
rect 13334 3225 13350 3289
rect 13414 3225 13430 3289
rect 13494 3225 13636 3289
rect 13700 3225 13716 3289
rect 13780 3225 13796 3289
rect 13860 3225 13876 3289
rect 13940 3225 13956 3289
rect 14020 3225 14036 3289
rect 14100 3225 14242 3289
rect 14306 3225 14322 3289
rect 14386 3225 14402 3289
rect 14466 3225 14482 3289
rect 14546 3225 14562 3289
rect 14626 3225 14642 3289
rect 14706 3225 14848 3289
rect 14912 3225 14928 3289
rect 14992 3225 15008 3289
rect 15072 3225 15088 3289
rect 15152 3225 15168 3289
rect 15232 3225 15248 3289
rect 15312 3225 15416 3289
rect 10502 3223 15416 3225
rect 10502 3069 10568 3159
rect 10502 3005 10503 3069
rect 10567 3005 10568 3069
rect 10502 2989 10568 3005
rect 10502 2925 10503 2989
rect 10567 2925 10568 2989
rect 10502 2909 10568 2925
rect 10502 2845 10503 2909
rect 10567 2845 10568 2909
rect 10502 2829 10568 2845
rect 10502 2765 10503 2829
rect 10567 2765 10568 2829
rect 10502 2749 10568 2765
rect 10502 2685 10503 2749
rect 10567 2685 10568 2749
rect 10502 2669 10568 2685
rect 10502 2605 10503 2669
rect 10567 2605 10568 2669
rect 10502 2589 10568 2605
rect 10502 2525 10503 2589
rect 10567 2525 10568 2589
rect 10502 2509 10568 2525
rect 10502 2445 10503 2509
rect 10567 2445 10568 2509
rect 10502 2429 10568 2445
rect 10502 2365 10503 2429
rect 10567 2365 10568 2429
rect 10502 2349 10568 2365
rect 10502 2285 10503 2349
rect 10567 2285 10568 2349
rect 10502 2131 10568 2285
rect 10628 2193 10688 3223
rect 10748 2131 10808 3163
rect 10868 2193 10928 3223
rect 10988 2131 11048 3163
rect 11108 3069 11174 3159
rect 11108 3005 11109 3069
rect 11173 3005 11174 3069
rect 11108 2989 11174 3005
rect 11108 2925 11109 2989
rect 11173 2925 11174 2989
rect 11108 2909 11174 2925
rect 11108 2845 11109 2909
rect 11173 2845 11174 2909
rect 11108 2829 11174 2845
rect 11108 2765 11109 2829
rect 11173 2765 11174 2829
rect 11108 2749 11174 2765
rect 11108 2685 11109 2749
rect 11173 2685 11174 2749
rect 11108 2669 11174 2685
rect 11108 2605 11109 2669
rect 11173 2605 11174 2669
rect 11108 2589 11174 2605
rect 11108 2525 11109 2589
rect 11173 2525 11174 2589
rect 11108 2509 11174 2525
rect 11108 2445 11109 2509
rect 11173 2445 11174 2509
rect 11108 2429 11174 2445
rect 11108 2365 11109 2429
rect 11173 2365 11174 2429
rect 11108 2349 11174 2365
rect 11108 2285 11109 2349
rect 11173 2285 11174 2349
rect 11108 2131 11174 2285
rect 11234 2193 11294 3223
rect 11354 2131 11414 3163
rect 11474 2193 11534 3223
rect 11594 2131 11654 3163
rect 11714 3069 11780 3159
rect 11714 3005 11715 3069
rect 11779 3005 11780 3069
rect 11714 2989 11780 3005
rect 11714 2925 11715 2989
rect 11779 2925 11780 2989
rect 11714 2909 11780 2925
rect 11714 2845 11715 2909
rect 11779 2845 11780 2909
rect 11714 2829 11780 2845
rect 11714 2765 11715 2829
rect 11779 2765 11780 2829
rect 11714 2749 11780 2765
rect 11714 2685 11715 2749
rect 11779 2685 11780 2749
rect 11714 2669 11780 2685
rect 11714 2605 11715 2669
rect 11779 2605 11780 2669
rect 11714 2589 11780 2605
rect 11714 2525 11715 2589
rect 11779 2525 11780 2589
rect 11714 2509 11780 2525
rect 11714 2445 11715 2509
rect 11779 2445 11780 2509
rect 11714 2429 11780 2445
rect 11714 2365 11715 2429
rect 11779 2365 11780 2429
rect 11714 2349 11780 2365
rect 11714 2285 11715 2349
rect 11779 2285 11780 2349
rect 11714 2131 11780 2285
rect 11840 2193 11900 3223
rect 11960 2131 12020 3163
rect 12080 2193 12140 3223
rect 12200 2131 12260 3163
rect 12320 3069 12386 3159
rect 12320 3005 12321 3069
rect 12385 3005 12386 3069
rect 12320 2989 12386 3005
rect 12320 2925 12321 2989
rect 12385 2925 12386 2989
rect 12320 2909 12386 2925
rect 12320 2845 12321 2909
rect 12385 2845 12386 2909
rect 12320 2829 12386 2845
rect 12320 2765 12321 2829
rect 12385 2765 12386 2829
rect 12320 2749 12386 2765
rect 12320 2685 12321 2749
rect 12385 2685 12386 2749
rect 12320 2669 12386 2685
rect 12320 2605 12321 2669
rect 12385 2605 12386 2669
rect 12320 2589 12386 2605
rect 12320 2525 12321 2589
rect 12385 2525 12386 2589
rect 12320 2509 12386 2525
rect 12320 2445 12321 2509
rect 12385 2445 12386 2509
rect 12320 2429 12386 2445
rect 12320 2365 12321 2429
rect 12385 2365 12386 2429
rect 12320 2349 12386 2365
rect 12320 2285 12321 2349
rect 12385 2285 12386 2349
rect 12320 2131 12386 2285
rect 12446 2193 12506 3223
rect 12566 2131 12626 3163
rect 12686 2193 12746 3223
rect 12806 2131 12866 3163
rect 12926 3069 12992 3159
rect 12926 3005 12927 3069
rect 12991 3005 12992 3069
rect 12926 2989 12992 3005
rect 12926 2925 12927 2989
rect 12991 2925 12992 2989
rect 12926 2909 12992 2925
rect 12926 2845 12927 2909
rect 12991 2845 12992 2909
rect 12926 2829 12992 2845
rect 12926 2765 12927 2829
rect 12991 2765 12992 2829
rect 12926 2749 12992 2765
rect 12926 2685 12927 2749
rect 12991 2685 12992 2749
rect 12926 2669 12992 2685
rect 12926 2605 12927 2669
rect 12991 2605 12992 2669
rect 12926 2589 12992 2605
rect 12926 2525 12927 2589
rect 12991 2525 12992 2589
rect 12926 2509 12992 2525
rect 12926 2445 12927 2509
rect 12991 2445 12992 2509
rect 12926 2429 12992 2445
rect 12926 2365 12927 2429
rect 12991 2365 12992 2429
rect 12926 2349 12992 2365
rect 12926 2285 12927 2349
rect 12991 2285 12992 2349
rect 12926 2131 12992 2285
rect 13052 2193 13112 3223
rect 13172 2131 13232 3163
rect 13292 2193 13352 3223
rect 13412 2131 13472 3163
rect 13532 3069 13598 3159
rect 13532 3005 13533 3069
rect 13597 3005 13598 3069
rect 13532 2989 13598 3005
rect 13532 2925 13533 2989
rect 13597 2925 13598 2989
rect 13532 2909 13598 2925
rect 13532 2845 13533 2909
rect 13597 2845 13598 2909
rect 13532 2829 13598 2845
rect 13532 2765 13533 2829
rect 13597 2765 13598 2829
rect 13532 2749 13598 2765
rect 13532 2685 13533 2749
rect 13597 2685 13598 2749
rect 13532 2669 13598 2685
rect 13532 2605 13533 2669
rect 13597 2605 13598 2669
rect 13532 2589 13598 2605
rect 13532 2525 13533 2589
rect 13597 2525 13598 2589
rect 13532 2509 13598 2525
rect 13532 2445 13533 2509
rect 13597 2445 13598 2509
rect 13532 2429 13598 2445
rect 13532 2365 13533 2429
rect 13597 2365 13598 2429
rect 13532 2349 13598 2365
rect 13532 2285 13533 2349
rect 13597 2285 13598 2349
rect 13532 2131 13598 2285
rect 13658 2193 13718 3223
rect 13778 2131 13838 3163
rect 13898 2193 13958 3223
rect 14018 2131 14078 3163
rect 14138 3069 14204 3159
rect 14138 3005 14139 3069
rect 14203 3005 14204 3069
rect 14138 2989 14204 3005
rect 14138 2925 14139 2989
rect 14203 2925 14204 2989
rect 14138 2909 14204 2925
rect 14138 2845 14139 2909
rect 14203 2845 14204 2909
rect 14138 2829 14204 2845
rect 14138 2765 14139 2829
rect 14203 2765 14204 2829
rect 14138 2749 14204 2765
rect 14138 2685 14139 2749
rect 14203 2685 14204 2749
rect 14138 2669 14204 2685
rect 14138 2605 14139 2669
rect 14203 2605 14204 2669
rect 14138 2589 14204 2605
rect 14138 2525 14139 2589
rect 14203 2525 14204 2589
rect 14138 2509 14204 2525
rect 14138 2445 14139 2509
rect 14203 2445 14204 2509
rect 14138 2429 14204 2445
rect 14138 2365 14139 2429
rect 14203 2365 14204 2429
rect 14138 2349 14204 2365
rect 14138 2285 14139 2349
rect 14203 2285 14204 2349
rect 14138 2131 14204 2285
rect 14264 2193 14324 3223
rect 14384 2131 14444 3163
rect 14504 2193 14564 3223
rect 14624 2131 14684 3163
rect 14744 3069 14810 3159
rect 14744 3005 14745 3069
rect 14809 3005 14810 3069
rect 14744 2989 14810 3005
rect 14744 2925 14745 2989
rect 14809 2925 14810 2989
rect 14744 2909 14810 2925
rect 14744 2845 14745 2909
rect 14809 2845 14810 2909
rect 14744 2829 14810 2845
rect 14744 2765 14745 2829
rect 14809 2765 14810 2829
rect 14744 2749 14810 2765
rect 14744 2685 14745 2749
rect 14809 2685 14810 2749
rect 14744 2669 14810 2685
rect 14744 2605 14745 2669
rect 14809 2605 14810 2669
rect 14744 2589 14810 2605
rect 14744 2525 14745 2589
rect 14809 2525 14810 2589
rect 14744 2509 14810 2525
rect 14744 2445 14745 2509
rect 14809 2445 14810 2509
rect 14744 2429 14810 2445
rect 14744 2365 14745 2429
rect 14809 2365 14810 2429
rect 14744 2349 14810 2365
rect 14744 2285 14745 2349
rect 14809 2285 14810 2349
rect 14744 2131 14810 2285
rect 14870 2193 14930 3223
rect 14990 2131 15050 3163
rect 15110 2193 15170 3223
rect 15230 2131 15290 3163
rect 15350 3069 15416 3159
rect 15350 3005 15351 3069
rect 15415 3005 15416 3069
rect 15350 2989 15416 3005
rect 15350 2925 15351 2989
rect 15415 2925 15416 2989
rect 15350 2909 15416 2925
rect 15350 2845 15351 2909
rect 15415 2845 15416 2909
rect 15350 2829 15416 2845
rect 15350 2765 15351 2829
rect 15415 2765 15416 2829
rect 15350 2749 15416 2765
rect 15350 2685 15351 2749
rect 15415 2685 15416 2749
rect 15350 2669 15416 2685
rect 15350 2605 15351 2669
rect 15415 2605 15416 2669
rect 15350 2589 15416 2605
rect 15350 2525 15351 2589
rect 15415 2525 15416 2589
rect 15350 2509 15416 2525
rect 15350 2445 15351 2509
rect 15415 2445 15416 2509
rect 15350 2429 15416 2445
rect 15350 2365 15351 2429
rect 15415 2365 15416 2429
rect 15536 2393 15964 3351
rect 15350 2349 15416 2365
rect 15350 2285 15351 2349
rect 15415 2285 15416 2349
rect 15350 2131 15416 2285
rect 10502 2129 15416 2131
rect 10502 2065 10606 2129
rect 10670 2065 10686 2129
rect 10750 2065 10766 2129
rect 10830 2065 10846 2129
rect 10910 2065 10926 2129
rect 10990 2065 11006 2129
rect 11070 2065 11212 2129
rect 11276 2065 11292 2129
rect 11356 2065 11372 2129
rect 11436 2065 11452 2129
rect 11516 2065 11532 2129
rect 11596 2065 11612 2129
rect 11676 2065 11818 2129
rect 11882 2065 11898 2129
rect 11962 2065 11978 2129
rect 12042 2065 12058 2129
rect 12122 2065 12138 2129
rect 12202 2065 12218 2129
rect 12282 2065 12424 2129
rect 12488 2065 12504 2129
rect 12568 2065 12584 2129
rect 12648 2065 12664 2129
rect 12728 2065 12744 2129
rect 12808 2065 12824 2129
rect 12888 2065 13030 2129
rect 13094 2065 13110 2129
rect 13174 2065 13190 2129
rect 13254 2065 13270 2129
rect 13334 2065 13350 2129
rect 13414 2065 13430 2129
rect 13494 2065 13636 2129
rect 13700 2065 13716 2129
rect 13780 2065 13796 2129
rect 13860 2065 13876 2129
rect 13940 2065 13956 2129
rect 14020 2065 14036 2129
rect 14100 2065 14242 2129
rect 14306 2065 14322 2129
rect 14386 2065 14402 2129
rect 14466 2065 14482 2129
rect 14546 2065 14562 2129
rect 14626 2065 14642 2129
rect 14706 2065 14848 2129
rect 14912 2065 14928 2129
rect 14992 2065 15008 2129
rect 15072 2065 15088 2129
rect 15152 2065 15168 2129
rect 15232 2065 15248 2129
rect 15312 2065 15416 2129
rect 10502 2063 15416 2065
rect 10502 1927 12992 1929
rect 10502 1863 10606 1927
rect 10670 1863 10686 1927
rect 10750 1863 10766 1927
rect 10830 1863 10846 1927
rect 10910 1863 10926 1927
rect 10990 1863 11006 1927
rect 11070 1863 11212 1927
rect 11276 1863 11292 1927
rect 11356 1863 11372 1927
rect 11436 1863 11452 1927
rect 11516 1863 11532 1927
rect 11596 1863 11612 1927
rect 11676 1863 11818 1927
rect 11882 1863 11898 1927
rect 11962 1863 11978 1927
rect 12042 1863 12058 1927
rect 12122 1863 12138 1927
rect 12202 1863 12218 1927
rect 12282 1863 12424 1927
rect 12488 1863 12504 1927
rect 12568 1863 12584 1927
rect 12648 1863 12664 1927
rect 12728 1863 12744 1927
rect 12808 1863 12824 1927
rect 12888 1863 12992 1927
rect 10502 1861 12992 1863
rect 10502 1707 10568 1861
rect 10502 1643 10503 1707
rect 10567 1643 10568 1707
rect 10502 1627 10568 1643
rect 10502 1563 10503 1627
rect 10567 1563 10568 1627
rect 10502 1547 10568 1563
rect 10502 1483 10503 1547
rect 10567 1483 10568 1547
rect 10502 1467 10568 1483
rect 10502 1403 10503 1467
rect 10567 1403 10568 1467
rect 10502 1387 10568 1403
rect 10502 1323 10503 1387
rect 10567 1323 10568 1387
rect 10502 1307 10568 1323
rect 10502 1243 10503 1307
rect 10567 1243 10568 1307
rect 10502 1227 10568 1243
rect 10230 641 10442 1224
rect 10502 1163 10503 1227
rect 10567 1163 10568 1227
rect 10502 1147 10568 1163
rect 10502 1083 10503 1147
rect 10567 1083 10568 1147
rect 10502 1067 10568 1083
rect 10502 1003 10503 1067
rect 10567 1003 10568 1067
rect 10502 987 10568 1003
rect 10502 923 10503 987
rect 10567 923 10568 987
rect 10502 833 10568 923
rect 10628 829 10688 1861
rect 10748 769 10808 1799
rect 10868 829 10928 1861
rect 10988 769 11048 1799
rect 11108 1707 11174 1861
rect 11108 1643 11109 1707
rect 11173 1643 11174 1707
rect 11108 1627 11174 1643
rect 11108 1563 11109 1627
rect 11173 1563 11174 1627
rect 11108 1547 11174 1563
rect 11108 1483 11109 1547
rect 11173 1483 11174 1547
rect 11108 1467 11174 1483
rect 11108 1403 11109 1467
rect 11173 1403 11174 1467
rect 11108 1387 11174 1403
rect 11108 1323 11109 1387
rect 11173 1323 11174 1387
rect 11108 1307 11174 1323
rect 11108 1243 11109 1307
rect 11173 1243 11174 1307
rect 11108 1227 11174 1243
rect 11108 1163 11109 1227
rect 11173 1163 11174 1227
rect 11108 1147 11174 1163
rect 11108 1083 11109 1147
rect 11173 1083 11174 1147
rect 11108 1067 11174 1083
rect 11108 1003 11109 1067
rect 11173 1003 11174 1067
rect 11108 987 11174 1003
rect 11108 923 11109 987
rect 11173 923 11174 987
rect 11108 833 11174 923
rect 11234 829 11294 1861
rect 11354 769 11414 1799
rect 11474 829 11534 1861
rect 11594 769 11654 1799
rect 11714 1707 11780 1861
rect 11714 1643 11715 1707
rect 11779 1643 11780 1707
rect 11714 1627 11780 1643
rect 11714 1563 11715 1627
rect 11779 1563 11780 1627
rect 11714 1547 11780 1563
rect 11714 1483 11715 1547
rect 11779 1483 11780 1547
rect 11714 1467 11780 1483
rect 11714 1403 11715 1467
rect 11779 1403 11780 1467
rect 11714 1387 11780 1403
rect 11714 1323 11715 1387
rect 11779 1323 11780 1387
rect 11714 1307 11780 1323
rect 11714 1243 11715 1307
rect 11779 1243 11780 1307
rect 11714 1227 11780 1243
rect 11714 1163 11715 1227
rect 11779 1163 11780 1227
rect 11714 1147 11780 1163
rect 11714 1083 11715 1147
rect 11779 1083 11780 1147
rect 11714 1067 11780 1083
rect 11714 1003 11715 1067
rect 11779 1003 11780 1067
rect 11714 987 11780 1003
rect 11714 923 11715 987
rect 11779 923 11780 987
rect 11714 833 11780 923
rect 11840 829 11900 1861
rect 11960 769 12020 1799
rect 12080 829 12140 1861
rect 12200 769 12260 1799
rect 12320 1707 12386 1861
rect 12320 1643 12321 1707
rect 12385 1643 12386 1707
rect 12320 1627 12386 1643
rect 12320 1563 12321 1627
rect 12385 1563 12386 1627
rect 12320 1547 12386 1563
rect 12320 1483 12321 1547
rect 12385 1483 12386 1547
rect 12320 1467 12386 1483
rect 12320 1403 12321 1467
rect 12385 1403 12386 1467
rect 12320 1387 12386 1403
rect 12320 1323 12321 1387
rect 12385 1323 12386 1387
rect 12320 1307 12386 1323
rect 12320 1243 12321 1307
rect 12385 1243 12386 1307
rect 12320 1227 12386 1243
rect 12320 1163 12321 1227
rect 12385 1163 12386 1227
rect 12320 1147 12386 1163
rect 12320 1083 12321 1147
rect 12385 1083 12386 1147
rect 12320 1067 12386 1083
rect 12320 1003 12321 1067
rect 12385 1003 12386 1067
rect 12320 987 12386 1003
rect 12320 923 12321 987
rect 12385 923 12386 987
rect 12320 833 12386 923
rect 12446 829 12506 1861
rect 12566 769 12626 1799
rect 12686 829 12746 1861
rect 12806 769 12866 1799
rect 12926 1707 12992 1861
rect 12926 1643 12927 1707
rect 12991 1643 12992 1707
rect 12926 1627 12992 1643
rect 12926 1563 12927 1627
rect 12991 1563 12992 1627
rect 12926 1547 12992 1563
rect 12926 1483 12927 1547
rect 12991 1483 12992 1547
rect 12926 1467 12992 1483
rect 12926 1403 12927 1467
rect 12991 1403 12992 1467
rect 12926 1387 12992 1403
rect 12926 1323 12927 1387
rect 12991 1323 12992 1387
rect 12926 1307 12992 1323
rect 12926 1243 12927 1307
rect 12991 1243 12992 1307
rect 12926 1227 12992 1243
rect 12926 1163 12927 1227
rect 12991 1163 12992 1227
rect 12926 1147 12992 1163
rect 12926 1083 12927 1147
rect 12991 1083 12992 1147
rect 12926 1067 12992 1083
rect 12926 1003 12927 1067
rect 12991 1003 12992 1067
rect 12926 987 12992 1003
rect 12926 923 12927 987
rect 12991 923 12992 987
rect 12926 833 12992 923
rect 13052 1927 14330 1929
rect 13052 1863 13156 1927
rect 13220 1863 13236 1927
rect 13300 1863 13316 1927
rect 13380 1863 13396 1927
rect 13460 1863 13476 1927
rect 13540 1863 13556 1927
rect 13620 1863 13762 1927
rect 13826 1863 13842 1927
rect 13906 1863 13922 1927
rect 13986 1863 14002 1927
rect 14066 1863 14082 1927
rect 14146 1863 14162 1927
rect 14226 1863 14330 1927
rect 13052 1861 14330 1863
rect 13052 1707 13118 1861
rect 13052 1643 13053 1707
rect 13117 1643 13118 1707
rect 13052 1627 13118 1643
rect 13052 1563 13053 1627
rect 13117 1563 13118 1627
rect 13052 1547 13118 1563
rect 13052 1483 13053 1547
rect 13117 1483 13118 1547
rect 13052 1467 13118 1483
rect 13052 1403 13053 1467
rect 13117 1403 13118 1467
rect 13052 1387 13118 1403
rect 13052 1323 13053 1387
rect 13117 1323 13118 1387
rect 13052 1307 13118 1323
rect 13052 1243 13053 1307
rect 13117 1243 13118 1307
rect 13052 1227 13118 1243
rect 13052 1163 13053 1227
rect 13117 1163 13118 1227
rect 13052 1147 13118 1163
rect 13052 1083 13053 1147
rect 13117 1083 13118 1147
rect 13052 1067 13118 1083
rect 13052 1003 13053 1067
rect 13117 1003 13118 1067
rect 13052 987 13118 1003
rect 13052 923 13053 987
rect 13117 923 13118 987
rect 13052 833 13118 923
rect 13178 829 13238 1861
rect 13298 769 13358 1799
rect 13418 829 13478 1861
rect 13538 769 13598 1799
rect 13658 1707 13724 1861
rect 13658 1643 13659 1707
rect 13723 1643 13724 1707
rect 13658 1627 13724 1643
rect 13658 1563 13659 1627
rect 13723 1563 13724 1627
rect 13658 1547 13724 1563
rect 13658 1483 13659 1547
rect 13723 1483 13724 1547
rect 13658 1467 13724 1483
rect 13658 1403 13659 1467
rect 13723 1403 13724 1467
rect 13658 1387 13724 1403
rect 13658 1323 13659 1387
rect 13723 1323 13724 1387
rect 13658 1307 13724 1323
rect 13658 1243 13659 1307
rect 13723 1243 13724 1307
rect 13658 1227 13724 1243
rect 13658 1163 13659 1227
rect 13723 1163 13724 1227
rect 13658 1147 13724 1163
rect 13658 1083 13659 1147
rect 13723 1083 13724 1147
rect 13658 1067 13724 1083
rect 13658 1003 13659 1067
rect 13723 1003 13724 1067
rect 13658 987 13724 1003
rect 13658 923 13659 987
rect 13723 923 13724 987
rect 13658 833 13724 923
rect 13784 829 13844 1861
rect 13904 769 13964 1799
rect 14024 829 14084 1861
rect 14144 769 14204 1799
rect 14264 1707 14330 1861
rect 14264 1643 14265 1707
rect 14329 1643 14330 1707
rect 14264 1627 14330 1643
rect 14264 1563 14265 1627
rect 14329 1563 14330 1627
rect 14264 1547 14330 1563
rect 14264 1483 14265 1547
rect 14329 1483 14330 1547
rect 14264 1467 14330 1483
rect 14264 1403 14265 1467
rect 14329 1403 14330 1467
rect 14264 1387 14330 1403
rect 14264 1323 14265 1387
rect 14329 1323 14330 1387
rect 14264 1307 14330 1323
rect 14264 1243 14265 1307
rect 14329 1243 14330 1307
rect 14264 1227 14330 1243
rect 14264 1163 14265 1227
rect 14329 1163 14330 1227
rect 14264 1147 14330 1163
rect 14264 1083 14265 1147
rect 14329 1083 14330 1147
rect 14264 1067 14330 1083
rect 14264 1003 14265 1067
rect 14329 1003 14330 1067
rect 14264 987 14330 1003
rect 14264 923 14265 987
rect 14329 923 14330 987
rect 14264 833 14330 923
rect 14390 1927 15062 1929
rect 14390 1863 14494 1927
rect 14558 1863 14574 1927
rect 14638 1863 14654 1927
rect 14718 1863 14734 1927
rect 14798 1863 14814 1927
rect 14878 1863 14894 1927
rect 14958 1863 15062 1927
rect 14390 1861 15062 1863
rect 14390 1707 14456 1861
rect 14390 1643 14391 1707
rect 14455 1643 14456 1707
rect 14390 1627 14456 1643
rect 14390 1563 14391 1627
rect 14455 1563 14456 1627
rect 14390 1547 14456 1563
rect 14390 1483 14391 1547
rect 14455 1483 14456 1547
rect 14390 1467 14456 1483
rect 14390 1403 14391 1467
rect 14455 1403 14456 1467
rect 14390 1387 14456 1403
rect 14390 1323 14391 1387
rect 14455 1323 14456 1387
rect 14390 1307 14456 1323
rect 14390 1243 14391 1307
rect 14455 1243 14456 1307
rect 14390 1227 14456 1243
rect 14390 1163 14391 1227
rect 14455 1163 14456 1227
rect 14390 1147 14456 1163
rect 14390 1083 14391 1147
rect 14455 1083 14456 1147
rect 14390 1067 14456 1083
rect 14390 1003 14391 1067
rect 14455 1003 14456 1067
rect 14390 987 14456 1003
rect 14390 923 14391 987
rect 14455 923 14456 987
rect 14390 833 14456 923
rect 14516 829 14576 1861
rect 14636 769 14696 1799
rect 14756 829 14816 1861
rect 14876 769 14936 1799
rect 14996 1707 15062 1861
rect 14996 1643 14997 1707
rect 15061 1643 15062 1707
rect 14996 1627 15062 1643
rect 14996 1563 14997 1627
rect 15061 1563 15062 1627
rect 14996 1547 15062 1563
rect 14996 1483 14997 1547
rect 15061 1483 15062 1547
rect 14996 1467 15062 1483
rect 14996 1403 14997 1467
rect 15061 1403 15062 1467
rect 14996 1387 15062 1403
rect 14996 1323 14997 1387
rect 15061 1323 15062 1387
rect 14996 1307 15062 1323
rect 14996 1243 14997 1307
rect 15061 1243 15062 1307
rect 14996 1227 15062 1243
rect 14996 1163 14997 1227
rect 15061 1163 15062 1227
rect 14996 1147 15062 1163
rect 14996 1083 14997 1147
rect 15061 1083 15062 1147
rect 14996 1067 15062 1083
rect 14996 1003 14997 1067
rect 15061 1003 15062 1067
rect 14996 987 15062 1003
rect 14996 923 14997 987
rect 15061 923 15062 987
rect 14996 833 15062 923
rect 10502 767 12992 769
rect 10502 703 10606 767
rect 10670 703 10686 767
rect 10750 703 10766 767
rect 10830 703 10846 767
rect 10910 703 10926 767
rect 10990 703 11006 767
rect 11070 703 11212 767
rect 11276 703 11292 767
rect 11356 703 11372 767
rect 11436 703 11452 767
rect 11516 703 11532 767
rect 11596 703 11612 767
rect 11676 703 11818 767
rect 11882 703 11898 767
rect 11962 703 11978 767
rect 12042 703 12058 767
rect 12122 703 12138 767
rect 12202 703 12218 767
rect 12282 703 12424 767
rect 12488 703 12504 767
rect 12568 703 12584 767
rect 12648 703 12664 767
rect 12728 703 12744 767
rect 12808 703 12824 767
rect 12888 703 12992 767
rect 10502 701 12992 703
rect 13052 767 14330 769
rect 13052 703 13156 767
rect 13220 703 13236 767
rect 13300 703 13316 767
rect 13380 703 13396 767
rect 13460 703 13476 767
rect 13540 703 13556 767
rect 13620 703 13762 767
rect 13826 703 13842 767
rect 13906 703 13922 767
rect 13986 703 14002 767
rect 14066 703 14082 767
rect 14146 703 14162 767
rect 14226 703 14330 767
rect 13052 701 14330 703
rect 14390 767 15062 769
rect 14390 703 14494 767
rect 14558 703 14574 767
rect 14638 703 14654 767
rect 14718 703 14734 767
rect 14798 703 14814 767
rect 14878 703 14894 767
rect 14958 703 15062 767
rect 14390 701 15062 703
rect 15409 641 15965 1639
rect 10230 506 15965 641
<< labels >>
flabel pwell 10828 1117 10854 1149 0 FreeSans 160 0 0 0 x2.x2.SUB
flabel metal4 10886 1451 10912 1483 0 FreeSans 320 0 0 0 x2.x2.CBOT
flabel metal4 10768 861 10794 893 0 FreeSans 320 0 0 0 x2.x2.CTOP
flabel pwell 11434 1117 11460 1149 0 FreeSans 160 0 0 0 x3[1].x2.SUB
flabel metal4 11492 1451 11518 1483 0 FreeSans 320 0 0 0 x3[1].x2.CBOT
flabel metal4 11374 861 11400 893 0 FreeSans 320 0 0 0 x3[1].x2.CTOP
flabel pwell 12040 1117 12066 1149 0 FreeSans 160 0 0 0 x3[0].x2.SUB
flabel metal4 12098 1451 12124 1483 0 FreeSans 320 0 0 0 x3[0].x2.CBOT
flabel metal4 11980 861 12006 893 0 FreeSans 320 0 0 0 x3[0].x2.CTOP
flabel pwell 12646 1117 12672 1149 0 FreeSans 160 0 0 0 x4[3].x2.SUB
flabel metal4 12704 1451 12730 1483 0 FreeSans 320 0 0 0 x4[3].x2.CBOT
flabel metal4 12586 861 12612 893 0 FreeSans 320 0 0 0 x4[3].x2.CTOP
flabel pwell 13378 1117 13404 1149 0 FreeSans 160 0 0 0 x4[2].x2.SUB
flabel metal4 13436 1451 13462 1483 0 FreeSans 320 0 0 0 x4[2].x2.CBOT
flabel metal4 13318 861 13344 893 0 FreeSans 320 0 0 0 x4[2].x2.CTOP
flabel pwell 13984 1117 14010 1149 0 FreeSans 160 0 0 0 x4[1].x2.SUB
flabel metal4 14042 1451 14068 1483 0 FreeSans 320 0 0 0 x4[1].x2.CBOT
flabel metal4 13924 861 13950 893 0 FreeSans 320 0 0 0 x4[1].x2.CTOP
flabel pwell 14716 1117 14742 1149 0 FreeSans 160 0 0 0 x4[0].x2.SUB
flabel metal4 14774 1451 14800 1483 0 FreeSans 320 0 0 0 x4[0].x2.CBOT
flabel metal4 14656 861 14682 893 0 FreeSans 320 0 0 0 x4[0].x2.CTOP
flabel metal4 10764 2509 10790 2541 0 FreeSans 320 0 0 0 x5[7].x1.CBOT
flabel metal4 10882 3099 10908 3131 0 FreeSans 320 0 0 0 x5[7].x1.CTOP
flabel nwell 10757 2763 10925 2931 0 FreeSans 320 0 0 0 x5[7].x1.SUB
flabel metal4 11370 2509 11396 2541 0 FreeSans 320 0 0 0 x5[6].x1.CBOT
flabel metal4 11488 3099 11514 3131 0 FreeSans 320 0 0 0 x5[6].x1.CTOP
flabel nwell 11363 2763 11531 2931 0 FreeSans 320 0 0 0 x5[6].x1.SUB
flabel metal4 12582 2509 12608 2541 0 FreeSans 320 0 0 0 x5[4].x1.CBOT
flabel metal4 12700 3099 12726 3131 0 FreeSans 320 0 0 0 x5[4].x1.CTOP
flabel nwell 12575 2763 12743 2931 0 FreeSans 320 0 0 0 x5[4].x1.SUB
flabel metal4 11976 2509 12002 2541 0 FreeSans 320 0 0 0 x5[5].x1.CBOT
flabel metal4 12094 3099 12120 3131 0 FreeSans 320 0 0 0 x5[5].x1.CTOP
flabel nwell 11969 2763 12137 2931 0 FreeSans 320 0 0 0 x5[5].x1.SUB
flabel metal4 13188 2509 13214 2541 0 FreeSans 320 0 0 0 x5[3].x1.CBOT
flabel metal4 13306 3099 13332 3131 0 FreeSans 320 0 0 0 x5[3].x1.CTOP
flabel nwell 13181 2763 13349 2931 0 FreeSans 320 0 0 0 x5[3].x1.SUB
flabel metal4 13794 2509 13820 2541 0 FreeSans 320 0 0 0 x5[2].x1.CBOT
flabel metal4 13912 3099 13938 3131 0 FreeSans 320 0 0 0 x5[2].x1.CTOP
flabel nwell 13787 2763 13955 2931 0 FreeSans 320 0 0 0 x5[2].x1.SUB
flabel metal4 14400 2509 14426 2541 0 FreeSans 320 0 0 0 x5[1].x1.CBOT
flabel metal4 14518 3099 14544 3131 0 FreeSans 320 0 0 0 x5[1].x1.CTOP
flabel nwell 14393 2763 14561 2931 0 FreeSans 320 0 0 0 x5[1].x1.SUB
flabel metal4 15006 2509 15032 2541 0 FreeSans 320 0 0 0 x5[0].x1.CBOT
flabel metal4 15124 3099 15150 3131 0 FreeSans 320 0 0 0 x5[0].x1.CTOP
flabel nwell 14999 2763 15167 2931 0 FreeSans 320 0 0 0 x5[0].x1.SUB
<< end >>
