magic
tech sky130A
magscale 1 2
timestamp 1697025759
<< pwell >>
rect -401 -348 401 348
<< nmos >>
rect -205 -138 205 138
<< ndiff >>
rect -263 126 -205 138
rect -263 -126 -251 126
rect -217 -126 -205 126
rect -263 -138 -205 -126
rect 205 126 263 138
rect 205 -126 217 126
rect 251 -126 263 126
rect 205 -138 263 -126
<< ndiffc >>
rect -251 -126 -217 126
rect 217 -126 251 126
<< psubdiff >>
rect -365 278 -269 312
rect 269 278 365 312
rect -365 216 -331 278
rect 331 216 365 278
rect -365 -278 -331 -216
rect 331 -278 365 -216
rect -365 -312 -269 -278
rect 269 -312 365 -278
<< psubdiffcont >>
rect -269 278 269 312
rect -365 -216 -331 216
rect 331 -216 365 216
rect -269 -312 269 -278
<< poly >>
rect -205 210 205 226
rect -205 176 -189 210
rect 189 176 205 210
rect -205 138 205 176
rect -205 -176 205 -138
rect -205 -210 -189 -176
rect 189 -210 205 -176
rect -205 -226 205 -210
<< polycont >>
rect -189 176 189 210
rect -189 -210 189 -176
<< locali >>
rect -365 278 -269 312
rect 269 278 365 312
rect -365 216 -331 278
rect 331 216 365 278
rect -205 176 -189 210
rect 189 176 205 210
rect -251 126 -217 142
rect -251 -142 -217 -126
rect 217 126 251 142
rect 217 -142 251 -126
rect -205 -210 -189 -176
rect 189 -210 205 -176
rect -365 -278 -331 -216
rect 331 -278 365 -216
rect -365 -312 -269 -278
rect 269 -312 365 -278
<< viali >>
rect -189 176 189 210
rect -251 -126 -217 126
rect 217 -126 251 126
rect -189 -210 189 -176
<< metal1 >>
rect -201 210 201 216
rect -201 176 -189 210
rect 189 176 201 210
rect -201 170 201 176
rect -257 126 -211 138
rect -257 -126 -251 126
rect -217 -126 -211 126
rect -257 -138 -211 -126
rect 211 126 257 138
rect 211 -126 217 126
rect 251 -126 257 126
rect 211 -138 257 -126
rect -201 -176 201 -170
rect -201 -210 -189 -176
rect 189 -210 201 -176
rect -201 -216 201 -210
<< properties >>
string FIXED_BBOX -348 -295 348 295
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.375 l 2.045 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
