magic
tech sky130A
timestamp 1706708090
<< nwell >>
rect 58 937 510 997
rect 230 339 247 340
rect 276 339 293 340
rect 322 339 339 340
rect 196 303 510 339
<< psubdiff >>
rect 77 655 491 663
rect 77 654 322 655
rect 77 653 277 654
rect 77 652 137 653
rect 77 635 93 652
rect 110 636 137 652
rect 154 651 229 653
rect 154 636 184 651
rect 110 635 184 636
rect 77 634 184 635
rect 201 636 229 651
rect 246 637 277 653
rect 294 638 322 654
rect 339 654 491 655
rect 339 638 370 654
rect 294 637 370 638
rect 387 653 491 654
rect 387 637 416 653
rect 246 636 416 637
rect 433 652 491 653
rect 433 636 460 652
rect 201 635 460 636
rect 477 635 491 652
rect 201 634 491 635
rect 77 623 491 634
<< nsubdiff >>
rect 77 970 491 975
rect 77 969 278 970
rect 77 952 92 969
rect 109 968 231 969
rect 109 952 138 968
rect 77 951 138 952
rect 155 951 183 968
rect 200 952 231 968
rect 248 953 278 969
rect 295 969 413 970
rect 295 953 323 969
rect 248 952 323 953
rect 340 952 368 969
rect 385 953 413 969
rect 430 969 491 970
rect 430 953 459 969
rect 385 952 459 953
rect 476 952 491 969
rect 200 951 491 952
rect 77 948 491 951
rect 215 323 230 340
rect 247 323 276 340
rect 293 323 322 340
rect 339 339 491 340
rect 339 323 367 339
rect 215 322 367 323
rect 384 322 413 339
rect 430 322 459 339
rect 476 322 491 339
<< psubdiffcont >>
rect 93 635 110 652
rect 137 636 154 653
rect 184 634 201 651
rect 229 636 246 653
rect 277 637 294 654
rect 322 638 339 655
rect 370 637 387 654
rect 416 636 433 653
rect 460 635 477 652
<< nsubdiffcont >>
rect 92 952 109 969
rect 138 951 155 968
rect 183 951 200 968
rect 231 952 248 969
rect 278 953 295 970
rect 323 952 340 969
rect 368 952 385 969
rect 413 953 430 970
rect 459 952 476 969
rect 230 323 247 340
rect 276 323 293 340
rect 322 323 339 340
rect 367 322 384 339
rect 413 322 430 339
rect 459 322 476 339
<< locali >>
rect 77 970 491 975
rect 77 969 278 970
rect 77 952 92 969
rect 109 968 231 969
rect 109 952 138 968
rect 77 951 138 952
rect 155 951 183 968
rect 200 952 231 968
rect 248 953 278 969
rect 295 969 413 970
rect 295 953 323 969
rect 248 952 323 953
rect 340 952 368 969
rect 385 953 413 969
rect 430 969 491 970
rect 430 953 459 969
rect 385 952 459 953
rect 476 952 491 969
rect 200 951 491 952
rect 77 947 491 951
rect 304 776 395 796
rect 77 655 491 663
rect 77 654 322 655
rect 77 653 277 654
rect 77 652 137 653
rect 77 635 93 652
rect 110 636 137 652
rect 154 651 229 653
rect 154 636 184 651
rect 110 635 184 636
rect 77 634 184 635
rect 201 636 229 651
rect 246 637 277 653
rect 294 638 322 654
rect 339 654 491 655
rect 339 638 370 654
rect 294 637 370 638
rect 387 653 491 654
rect 387 637 416 653
rect 246 636 416 637
rect 433 652 491 653
rect 433 636 460 652
rect 201 635 460 636
rect 477 635 491 652
rect 201 634 491 635
rect 77 623 491 634
rect 299 489 403 509
rect 215 323 230 340
rect 247 323 276 340
rect 293 323 322 340
rect 339 339 491 340
rect 339 323 367 339
rect 215 322 367 323
rect 384 322 413 339
rect 430 322 459 339
rect 476 322 491 339
<< viali >>
rect 138 848 155 865
rect 92 776 109 793
rect 180 780 197 797
rect 254 779 271 796
rect 438 778 455 795
rect 248 490 265 507
rect 436 490 453 507
<< metal1 >>
rect 487 916 639 973
rect 129 870 164 878
rect 129 865 276 870
rect 129 848 138 865
rect 155 848 276 865
rect 129 845 276 848
rect 129 841 164 845
rect 33 793 119 801
rect 33 776 92 793
rect 109 776 119 793
rect 33 768 119 776
rect 171 799 204 803
rect 250 799 276 845
rect 171 773 174 799
rect 200 773 204 799
rect 247 796 279 799
rect 247 779 254 796
rect 271 779 279 796
rect 247 773 279 779
rect 427 796 466 801
rect 171 771 204 773
rect 427 770 434 796
rect 460 770 466 796
rect 427 768 466 770
rect 53 653 230 692
rect 53 636 246 653
rect 277 637 294 654
rect 322 638 339 655
rect 370 637 387 654
rect 416 636 433 653
rect 53 595 230 636
rect 427 513 461 515
rect 72 512 271 513
rect 72 486 176 512
rect 202 507 271 512
rect 202 490 248 507
rect 265 490 271 507
rect 202 486 271 490
rect 72 484 271 486
rect 427 487 430 513
rect 457 487 461 513
rect 427 484 461 487
rect 72 483 216 484
rect 538 371 639 916
rect 230 323 247 340
rect 276 323 293 340
rect 322 323 339 340
rect 367 322 384 339
rect 486 322 639 371
<< via1 >>
rect 174 797 200 799
rect 174 780 180 797
rect 180 780 197 797
rect 197 780 200 797
rect 174 773 200 780
rect 434 795 460 796
rect 434 778 438 795
rect 438 778 455 795
rect 455 778 460 795
rect 434 770 460 778
rect 176 486 202 512
rect 430 507 457 513
rect 430 490 436 507
rect 436 490 453 507
rect 453 490 457 507
rect 430 487 457 490
<< metal2 >>
rect 171 799 204 803
rect 171 773 174 799
rect 200 783 204 799
rect 427 796 464 801
rect 200 773 207 783
rect 171 512 207 773
rect 171 486 176 512
rect 202 486 207 512
rect 171 484 207 486
rect 427 770 434 796
rect 460 770 464 796
rect 427 513 464 770
rect 427 487 430 513
rect 457 487 464 513
rect 427 484 464 487
use sky130_fd_sc_hd__inv_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 215 0 1 667
box -19 -24 157 296
use sky130_fd_sc_hd__inv_1  x2
timestamp 1701704242
transform 1 0 353 0 1 667
box -19 -24 157 296
use sky130_fd_sc_hd__inv_1  x3
timestamp 1701704242
transform -1 0 491 0 -1 619
box -19 -24 157 296
use sky130_fd_sc_hd__inv_1  x4
timestamp 1701704242
transform -1 0 353 0 -1 619
box -19 -24 157 296
use sky130_fd_sc_hd__nand2_1  x5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 215 0 1 667
box -19 -24 157 296
<< labels >>
flabel metal1 72 483 176 513 0 FreeSans 160 0 0 0 ring_osil
port 1 nsew
flabel metal1 538 322 639 973 0 FreeSans 160 0 0 0 vdd
port 2 nsew
flabel metal1 33 768 92 801 0 FreeSans 160 0 0 0 en
port 0 nsew
flabel metal1 53 595 230 692 0 FreeSans 160 0 0 0 gnd
port 5 nsew
<< end >>
