magic
tech sky130A
magscale 1 2
timestamp 1698845081
<< nwell >>
rect 9760 2342 15943 2993
rect 9262 2021 15943 2342
rect 9760 1813 15943 2021
rect 9760 1662 15989 1813
rect 10436 1629 10654 1662
rect 11168 1629 11512 1662
rect 12380 1629 12724 1662
rect 13592 1629 13936 1662
rect 14804 1629 15148 1662
rect 15578 1644 15989 1662
rect 15578 1643 15797 1644
<< pwell >>
rect 9342 1781 9528 1963
rect 9532 1781 9718 1963
rect 9342 1777 9363 1781
rect 9329 1743 9363 1777
rect 9697 1777 9718 1781
rect 9697 1743 9731 1777
rect 10575 669 10745 839
rect 11307 669 11477 839
rect 11911 669 12081 839
rect 12519 669 12689 839
rect 13123 669 13293 839
rect 13857 669 14027 839
rect 14461 669 14631 839
rect 15193 669 15363 839
<< nmos >>
rect 10885 1477 10915 1561
rect 11617 1477 11647 1561
rect 11741 1477 11771 1561
rect 12829 1477 12859 1561
rect 12953 1477 12983 1561
rect 14167 1477 14197 1561
rect 14291 1477 14321 1561
rect 15023 1477 15053 1561
rect 15673 1478 15703 1562
rect 15765 1478 15795 1562
rect 15861 1478 15891 1562
rect 9863 1293 9893 1377
rect 9935 1293 9965 1377
rect 15673 1340 15703 1424
rect 9863 1155 9893 1239
rect 9935 1155 9965 1239
rect 9863 1017 9893 1101
rect 9935 1017 9965 1101
rect 9863 879 9893 963
rect 9935 879 9965 963
rect 9863 741 9893 825
rect 9935 741 9965 825
rect 9863 603 9893 687
rect 9935 603 9965 687
rect 9863 465 9893 549
rect 9935 465 9965 549
rect 9863 327 9893 411
rect 9935 327 9965 411
<< scnmos >>
rect 9420 1807 9450 1937
rect 9610 1807 9640 1937
<< pmos >>
rect 10530 1678 10560 1762
rect 11262 1678 11292 1762
rect 11388 1678 11418 1762
rect 12474 1678 12504 1762
rect 12600 1678 12630 1762
rect 13686 1678 13716 1762
rect 13812 1678 13842 1762
rect 14898 1678 14928 1762
rect 15024 1678 15054 1762
<< scpmoshvt >>
rect 9420 2057 9450 2257
rect 9610 2057 9640 2257
<< pmoshvt >>
rect 9909 2820 9939 2904
rect 9909 2682 9939 2766
rect 9909 2544 9939 2628
rect 9909 2406 9939 2490
rect 9909 2268 9939 2352
rect 9909 2130 9939 2214
rect 15673 1819 15703 1903
rect 15673 1681 15703 1765
rect 15765 1681 15795 1765
rect 15861 1681 15891 1765
<< ndiff >>
rect 9368 1925 9420 1937
rect 9368 1891 9376 1925
rect 9410 1891 9420 1925
rect 9368 1857 9420 1891
rect 9368 1823 9376 1857
rect 9410 1823 9420 1857
rect 9368 1807 9420 1823
rect 9450 1925 9502 1937
rect 9450 1891 9460 1925
rect 9494 1891 9502 1925
rect 9450 1857 9502 1891
rect 9450 1823 9460 1857
rect 9494 1823 9502 1857
rect 9450 1807 9502 1823
rect 9558 1925 9610 1937
rect 9558 1891 9566 1925
rect 9600 1891 9610 1925
rect 9558 1857 9610 1891
rect 9558 1823 9566 1857
rect 9600 1823 9610 1857
rect 9558 1807 9610 1823
rect 9640 1925 9692 1937
rect 9640 1891 9650 1925
rect 9684 1891 9692 1925
rect 9640 1857 9692 1891
rect 9640 1823 9650 1857
rect 9684 1823 9692 1857
rect 9640 1807 9692 1823
rect 10827 1549 10885 1561
rect 10827 1489 10839 1549
rect 10873 1489 10885 1549
rect 10827 1477 10885 1489
rect 10915 1549 10973 1561
rect 10915 1489 10927 1549
rect 10961 1489 10973 1549
rect 10915 1477 10973 1489
rect 11559 1549 11617 1561
rect 11559 1489 11571 1549
rect 11605 1489 11617 1549
rect 11559 1477 11617 1489
rect 11647 1549 11741 1561
rect 11647 1489 11676 1549
rect 11710 1489 11741 1549
rect 11647 1477 11741 1489
rect 11771 1549 11829 1561
rect 11771 1489 11783 1549
rect 11817 1489 11829 1549
rect 11771 1477 11829 1489
rect 12771 1549 12829 1561
rect 12771 1489 12783 1549
rect 12817 1489 12829 1549
rect 12771 1477 12829 1489
rect 12859 1549 12953 1561
rect 12859 1489 12887 1549
rect 12921 1489 12953 1549
rect 12859 1477 12953 1489
rect 12983 1549 13041 1561
rect 12983 1489 12995 1549
rect 13029 1489 13041 1549
rect 12983 1477 13041 1489
rect 14109 1549 14167 1561
rect 14109 1489 14121 1549
rect 14155 1489 14167 1549
rect 14109 1477 14167 1489
rect 14197 1549 14291 1561
rect 14197 1489 14227 1549
rect 14261 1489 14291 1549
rect 14197 1477 14291 1489
rect 14321 1549 14379 1561
rect 14321 1489 14333 1549
rect 14367 1489 14379 1549
rect 14321 1477 14379 1489
rect 14964 1549 15023 1561
rect 14964 1489 14976 1549
rect 15010 1489 15023 1549
rect 14964 1477 15023 1489
rect 15053 1549 15111 1561
rect 15053 1489 15065 1549
rect 15099 1489 15111 1549
rect 15053 1477 15111 1489
rect 15615 1550 15673 1562
rect 15615 1490 15627 1550
rect 15661 1490 15673 1550
rect 15615 1478 15673 1490
rect 15703 1550 15765 1562
rect 15703 1490 15715 1550
rect 15749 1490 15765 1550
rect 15703 1478 15765 1490
rect 15795 1550 15861 1562
rect 15795 1490 15811 1550
rect 15845 1490 15861 1550
rect 15795 1478 15861 1490
rect 15891 1550 15953 1562
rect 15891 1490 15907 1550
rect 15941 1490 15953 1550
rect 15891 1478 15953 1490
rect 15615 1412 15673 1424
rect 9805 1365 9863 1377
rect 9805 1305 9817 1365
rect 9851 1305 9863 1365
rect 9805 1293 9863 1305
rect 9893 1293 9935 1377
rect 9965 1365 10023 1377
rect 9965 1305 9977 1365
rect 10011 1305 10023 1365
rect 15615 1352 15627 1412
rect 15661 1352 15673 1412
rect 15615 1340 15673 1352
rect 15703 1412 15761 1424
rect 15703 1352 15715 1412
rect 15749 1352 15761 1412
rect 15703 1340 15761 1352
rect 9965 1293 10023 1305
rect 9805 1227 9863 1239
rect 9805 1167 9817 1227
rect 9851 1167 9863 1227
rect 9805 1155 9863 1167
rect 9893 1155 9935 1239
rect 9965 1227 10023 1239
rect 9965 1167 9977 1227
rect 10011 1167 10023 1227
rect 9965 1155 10023 1167
rect 9805 1089 9863 1101
rect 9805 1029 9817 1089
rect 9851 1029 9863 1089
rect 9805 1017 9863 1029
rect 9893 1017 9935 1101
rect 9965 1089 10023 1101
rect 9965 1029 9977 1089
rect 10011 1029 10023 1089
rect 9965 1017 10023 1029
rect 9805 951 9863 963
rect 9805 891 9817 951
rect 9851 891 9863 951
rect 9805 879 9863 891
rect 9893 879 9935 963
rect 9965 951 10023 963
rect 9965 891 9977 951
rect 10011 891 10023 951
rect 9965 879 10023 891
rect 9805 813 9863 825
rect 9805 753 9817 813
rect 9851 753 9863 813
rect 9805 741 9863 753
rect 9893 741 9935 825
rect 9965 813 10023 825
rect 9965 753 9977 813
rect 10011 753 10023 813
rect 9965 741 10023 753
rect 9805 675 9863 687
rect 9805 615 9817 675
rect 9851 615 9863 675
rect 9805 603 9863 615
rect 9893 603 9935 687
rect 9965 675 10023 687
rect 9965 615 9977 675
rect 10011 615 10023 675
rect 9965 603 10023 615
rect 9805 537 9863 549
rect 9805 477 9817 537
rect 9851 477 9863 537
rect 9805 465 9863 477
rect 9893 465 9935 549
rect 9965 537 10023 549
rect 9965 477 9977 537
rect 10011 477 10023 537
rect 9965 465 10023 477
rect 9805 399 9863 411
rect 9805 339 9817 399
rect 9851 339 9863 399
rect 9805 327 9863 339
rect 9893 327 9935 411
rect 9965 399 10023 411
rect 9965 339 9977 399
rect 10011 339 10023 399
rect 9965 327 10023 339
<< pdiff >>
rect 9851 2892 9909 2904
rect 9851 2832 9863 2892
rect 9897 2832 9909 2892
rect 9851 2820 9909 2832
rect 9939 2892 9997 2904
rect 9939 2832 9951 2892
rect 9985 2832 9997 2892
rect 9939 2820 9997 2832
rect 9851 2754 9909 2766
rect 9851 2694 9863 2754
rect 9897 2694 9909 2754
rect 9851 2682 9909 2694
rect 9939 2754 9997 2766
rect 9939 2694 9951 2754
rect 9985 2694 9997 2754
rect 9939 2682 9997 2694
rect 9851 2616 9909 2628
rect 9851 2556 9863 2616
rect 9897 2556 9909 2616
rect 9851 2544 9909 2556
rect 9939 2616 9997 2628
rect 9939 2556 9951 2616
rect 9985 2556 9997 2616
rect 9939 2544 9997 2556
rect 9851 2478 9909 2490
rect 9851 2418 9863 2478
rect 9897 2418 9909 2478
rect 9851 2406 9909 2418
rect 9939 2478 9997 2490
rect 9939 2418 9951 2478
rect 9985 2418 9997 2478
rect 9939 2406 9997 2418
rect 9851 2340 9909 2352
rect 9851 2280 9863 2340
rect 9897 2280 9909 2340
rect 9851 2268 9909 2280
rect 9939 2340 9997 2352
rect 9939 2280 9951 2340
rect 9985 2280 9997 2340
rect 9939 2268 9997 2280
rect 9368 2245 9420 2257
rect 9368 2211 9376 2245
rect 9410 2211 9420 2245
rect 9368 2177 9420 2211
rect 9368 2143 9376 2177
rect 9410 2143 9420 2177
rect 9368 2109 9420 2143
rect 9368 2075 9376 2109
rect 9410 2075 9420 2109
rect 9368 2057 9420 2075
rect 9450 2245 9502 2257
rect 9450 2211 9460 2245
rect 9494 2211 9502 2245
rect 9450 2177 9502 2211
rect 9450 2143 9460 2177
rect 9494 2143 9502 2177
rect 9450 2109 9502 2143
rect 9450 2075 9460 2109
rect 9494 2075 9502 2109
rect 9450 2057 9502 2075
rect 9558 2245 9610 2257
rect 9558 2211 9566 2245
rect 9600 2211 9610 2245
rect 9558 2177 9610 2211
rect 9558 2143 9566 2177
rect 9600 2143 9610 2177
rect 9558 2109 9610 2143
rect 9558 2075 9566 2109
rect 9600 2075 9610 2109
rect 9558 2057 9610 2075
rect 9640 2245 9692 2257
rect 9640 2211 9650 2245
rect 9684 2211 9692 2245
rect 9640 2177 9692 2211
rect 9640 2143 9650 2177
rect 9684 2143 9692 2177
rect 9640 2109 9692 2143
rect 9851 2202 9909 2214
rect 9851 2142 9863 2202
rect 9897 2142 9909 2202
rect 9851 2130 9909 2142
rect 9939 2202 9997 2214
rect 9939 2142 9951 2202
rect 9985 2142 9997 2202
rect 9939 2130 9997 2142
rect 9640 2075 9650 2109
rect 9684 2075 9692 2109
rect 9640 2057 9692 2075
rect 15615 1891 15673 1903
rect 15615 1831 15627 1891
rect 15661 1831 15673 1891
rect 15615 1819 15673 1831
rect 15703 1891 15761 1903
rect 15703 1831 15715 1891
rect 15749 1831 15761 1891
rect 15703 1819 15761 1831
rect 10472 1750 10530 1762
rect 10472 1690 10484 1750
rect 10518 1690 10530 1750
rect 10472 1678 10530 1690
rect 10560 1750 10618 1762
rect 10560 1690 10572 1750
rect 10606 1690 10618 1750
rect 10560 1678 10618 1690
rect 11204 1750 11262 1762
rect 11204 1690 11216 1750
rect 11250 1690 11262 1750
rect 11204 1678 11262 1690
rect 11292 1750 11388 1762
rect 11292 1690 11321 1750
rect 11355 1690 11388 1750
rect 11292 1678 11388 1690
rect 11418 1750 11476 1762
rect 11418 1690 11430 1750
rect 11464 1690 11476 1750
rect 11418 1678 11476 1690
rect 12416 1750 12474 1762
rect 12416 1690 12428 1750
rect 12462 1690 12474 1750
rect 12416 1678 12474 1690
rect 12504 1750 12600 1762
rect 12504 1690 12532 1750
rect 12566 1690 12600 1750
rect 12504 1678 12600 1690
rect 12630 1750 12688 1762
rect 12630 1690 12642 1750
rect 12676 1690 12688 1750
rect 12630 1678 12688 1690
rect 13628 1750 13686 1762
rect 13628 1690 13640 1750
rect 13674 1690 13686 1750
rect 13628 1678 13686 1690
rect 13716 1750 13812 1762
rect 13716 1690 13745 1750
rect 13779 1690 13812 1750
rect 13716 1678 13812 1690
rect 13842 1750 13900 1762
rect 13842 1690 13854 1750
rect 13888 1690 13900 1750
rect 13842 1678 13900 1690
rect 14840 1750 14898 1762
rect 14840 1690 14852 1750
rect 14886 1690 14898 1750
rect 14840 1678 14898 1690
rect 14928 1750 15024 1762
rect 14928 1690 14959 1750
rect 14993 1690 15024 1750
rect 14928 1678 15024 1690
rect 15054 1750 15112 1762
rect 15054 1690 15066 1750
rect 15100 1690 15112 1750
rect 15054 1678 15112 1690
rect 15615 1753 15673 1765
rect 15615 1693 15627 1753
rect 15661 1693 15673 1753
rect 15615 1681 15673 1693
rect 15703 1753 15765 1765
rect 15703 1693 15715 1753
rect 15749 1693 15765 1753
rect 15703 1681 15765 1693
rect 15795 1753 15861 1765
rect 15795 1693 15811 1753
rect 15845 1693 15861 1753
rect 15795 1681 15861 1693
rect 15891 1753 15953 1765
rect 15891 1693 15907 1753
rect 15941 1693 15953 1753
rect 15891 1681 15953 1693
<< ndiffc >>
rect 9376 1891 9410 1925
rect 9376 1823 9410 1857
rect 9460 1891 9494 1925
rect 9460 1823 9494 1857
rect 9566 1891 9600 1925
rect 9566 1823 9600 1857
rect 9650 1891 9684 1925
rect 9650 1823 9684 1857
rect 10839 1489 10873 1549
rect 10927 1489 10961 1549
rect 11571 1489 11605 1549
rect 11676 1489 11710 1549
rect 11783 1489 11817 1549
rect 12783 1489 12817 1549
rect 12887 1489 12921 1549
rect 12995 1489 13029 1549
rect 14121 1489 14155 1549
rect 14227 1489 14261 1549
rect 14333 1489 14367 1549
rect 14976 1489 15010 1549
rect 15065 1489 15099 1549
rect 15627 1490 15661 1550
rect 15715 1490 15749 1550
rect 15811 1490 15845 1550
rect 15907 1490 15941 1550
rect 9817 1305 9851 1365
rect 9977 1305 10011 1365
rect 15627 1352 15661 1412
rect 15715 1352 15749 1412
rect 9817 1167 9851 1227
rect 9977 1167 10011 1227
rect 9817 1029 9851 1089
rect 9977 1029 10011 1089
rect 9817 891 9851 951
rect 9977 891 10011 951
rect 9817 753 9851 813
rect 9977 753 10011 813
rect 9817 615 9851 675
rect 9977 615 10011 675
rect 9817 477 9851 537
rect 9977 477 10011 537
rect 9817 339 9851 399
rect 9977 339 10011 399
<< pdiffc >>
rect 9863 2832 9897 2892
rect 9951 2832 9985 2892
rect 9863 2694 9897 2754
rect 9951 2694 9985 2754
rect 9863 2556 9897 2616
rect 9951 2556 9985 2616
rect 9863 2418 9897 2478
rect 9951 2418 9985 2478
rect 9863 2280 9897 2340
rect 9951 2280 9985 2340
rect 9376 2211 9410 2245
rect 9376 2143 9410 2177
rect 9376 2075 9410 2109
rect 9460 2211 9494 2245
rect 9460 2143 9494 2177
rect 9460 2075 9494 2109
rect 9566 2211 9600 2245
rect 9566 2143 9600 2177
rect 9566 2075 9600 2109
rect 9650 2211 9684 2245
rect 9650 2143 9684 2177
rect 9863 2142 9897 2202
rect 9951 2142 9985 2202
rect 9650 2075 9684 2109
rect 15627 1831 15661 1891
rect 15715 1831 15749 1891
rect 10484 1690 10518 1750
rect 10572 1690 10606 1750
rect 11216 1690 11250 1750
rect 11321 1690 11355 1750
rect 11430 1690 11464 1750
rect 12428 1690 12462 1750
rect 12532 1690 12566 1750
rect 12642 1690 12676 1750
rect 13640 1690 13674 1750
rect 13745 1690 13779 1750
rect 13854 1690 13888 1750
rect 14852 1690 14886 1750
rect 14959 1690 14993 1750
rect 15066 1690 15100 1750
rect 15627 1693 15661 1753
rect 15715 1693 15749 1753
rect 15811 1693 15845 1753
rect 15907 1693 15941 1753
<< poly >>
rect 9909 2904 9939 2934
rect 9909 2766 9939 2820
rect 9909 2628 9939 2682
rect 9909 2490 9939 2544
rect 9909 2352 9939 2406
rect 9420 2257 9450 2283
rect 9610 2257 9640 2283
rect 9909 2214 9939 2268
rect 9909 2099 9939 2130
rect 9891 2083 9957 2099
rect 9420 2025 9450 2057
rect 9364 2009 9450 2025
rect 9364 1975 9380 2009
rect 9414 1975 9450 2009
rect 9364 1959 9450 1975
rect 9420 1937 9450 1959
rect 9610 2025 9640 2057
rect 9891 2049 9907 2083
rect 9941 2049 9957 2083
rect 9891 2033 9957 2049
rect 9610 2009 9696 2025
rect 9610 1975 9646 2009
rect 9680 1975 9696 2009
rect 9610 1959 9696 1975
rect 9610 1937 9640 1959
rect 15673 1903 15703 1934
rect 10512 1843 10578 1859
rect 10512 1809 10528 1843
rect 10562 1809 10578 1843
rect 9420 1781 9450 1807
rect 9610 1781 9640 1807
rect 10512 1793 10578 1809
rect 11244 1843 11310 1859
rect 11244 1809 11260 1843
rect 11294 1809 11310 1843
rect 11244 1793 11310 1809
rect 11370 1843 11436 1859
rect 11370 1809 11386 1843
rect 11420 1809 11436 1843
rect 11370 1793 11436 1809
rect 12456 1843 12522 1859
rect 12456 1809 12472 1843
rect 12506 1809 12522 1843
rect 12456 1793 12522 1809
rect 12582 1843 12648 1859
rect 12582 1809 12598 1843
rect 12632 1809 12648 1843
rect 12582 1793 12648 1809
rect 13668 1843 13734 1859
rect 13668 1809 13684 1843
rect 13718 1809 13734 1843
rect 13668 1793 13734 1809
rect 13794 1843 13860 1859
rect 13794 1809 13810 1843
rect 13844 1809 13860 1843
rect 13794 1793 13860 1809
rect 14880 1843 14946 1859
rect 14880 1809 14896 1843
rect 14930 1809 14946 1843
rect 14880 1793 14946 1809
rect 15006 1843 15072 1859
rect 15006 1809 15022 1843
rect 15056 1809 15072 1843
rect 15006 1793 15072 1809
rect 10530 1762 10560 1793
rect 11262 1762 11292 1793
rect 11388 1762 11418 1793
rect 12474 1762 12504 1793
rect 12600 1762 12630 1793
rect 13686 1762 13716 1793
rect 13812 1762 13842 1793
rect 14898 1762 14928 1793
rect 15024 1762 15054 1793
rect 15673 1765 15703 1819
rect 15765 1765 15795 1791
rect 15861 1765 15891 1796
rect 10530 1650 10560 1678
rect 11262 1650 11292 1678
rect 11388 1650 11418 1678
rect 12474 1650 12504 1678
rect 12600 1650 12630 1678
rect 13686 1650 13716 1678
rect 13812 1650 13842 1678
rect 14898 1650 14928 1678
rect 15024 1650 15054 1678
rect 15673 1656 15703 1681
rect 15544 1636 15703 1656
rect 15765 1656 15795 1681
rect 15861 1656 15891 1681
rect 15765 1650 15891 1656
rect 15544 1602 15556 1636
rect 15590 1602 15703 1636
rect 10885 1561 10915 1587
rect 11617 1561 11647 1587
rect 11741 1561 11771 1587
rect 12829 1561 12859 1587
rect 12953 1561 12983 1587
rect 14167 1561 14197 1587
rect 14291 1561 14321 1587
rect 15023 1561 15053 1587
rect 15544 1583 15703 1602
rect 15747 1634 15891 1650
rect 15747 1600 15763 1634
rect 15797 1600 15891 1634
rect 15747 1584 15891 1600
rect 15673 1562 15703 1583
rect 15765 1577 15891 1584
rect 15765 1562 15795 1577
rect 15861 1562 15891 1577
rect 9881 1449 9947 1465
rect 10885 1455 10915 1477
rect 11617 1455 11647 1477
rect 11741 1455 11771 1477
rect 12829 1455 12859 1477
rect 12953 1455 12983 1477
rect 14167 1455 14197 1477
rect 14291 1455 14321 1477
rect 15023 1455 15053 1477
rect 9881 1422 9897 1449
rect 9863 1415 9897 1422
rect 9931 1422 9947 1449
rect 10867 1439 10933 1455
rect 9931 1415 9965 1422
rect 9863 1392 9965 1415
rect 9863 1377 9893 1392
rect 9935 1377 9965 1392
rect 10867 1405 10883 1439
rect 10917 1405 10933 1439
rect 10867 1389 10933 1405
rect 11599 1439 11665 1455
rect 11599 1405 11615 1439
rect 11649 1405 11665 1439
rect 11599 1389 11665 1405
rect 11723 1439 11789 1455
rect 11723 1405 11739 1439
rect 11773 1405 11789 1439
rect 11723 1389 11789 1405
rect 12811 1439 12877 1455
rect 12811 1405 12827 1439
rect 12861 1405 12877 1439
rect 12811 1389 12877 1405
rect 12935 1439 13001 1455
rect 12935 1405 12951 1439
rect 12985 1405 13001 1439
rect 12935 1389 13001 1405
rect 14149 1439 14215 1455
rect 14149 1405 14165 1439
rect 14199 1405 14215 1439
rect 14149 1389 14215 1405
rect 14273 1439 14339 1455
rect 14273 1405 14289 1439
rect 14323 1405 14339 1439
rect 14273 1389 14339 1405
rect 15005 1439 15071 1455
rect 15005 1405 15021 1439
rect 15055 1405 15071 1439
rect 15673 1424 15703 1478
rect 15765 1452 15795 1478
rect 15861 1452 15891 1478
rect 15005 1389 15071 1405
rect 15673 1313 15703 1340
rect 9863 1239 9893 1293
rect 9935 1239 9965 1293
rect 9863 1101 9893 1155
rect 9935 1101 9965 1155
rect 9863 963 9893 1017
rect 9935 963 9965 1017
rect 9863 825 9893 879
rect 9935 825 9965 879
rect 9863 687 9893 741
rect 9935 687 9965 741
rect 9863 549 9893 603
rect 9935 549 9965 603
rect 9863 411 9893 465
rect 9935 411 9965 465
rect 9863 301 9893 327
rect 9935 301 9965 327
<< polycont >>
rect 9380 1975 9414 2009
rect 9907 2049 9941 2083
rect 9646 1975 9680 2009
rect 10528 1809 10562 1843
rect 11260 1809 11294 1843
rect 11386 1809 11420 1843
rect 12472 1809 12506 1843
rect 12598 1809 12632 1843
rect 13684 1809 13718 1843
rect 13810 1809 13844 1843
rect 14896 1809 14930 1843
rect 15022 1809 15056 1843
rect 15556 1602 15590 1636
rect 15763 1600 15797 1634
rect 9897 1415 9931 1449
rect 10883 1405 10917 1439
rect 11615 1405 11649 1439
rect 11739 1405 11773 1439
rect 12827 1405 12861 1439
rect 12951 1405 12985 1439
rect 14165 1405 14199 1439
rect 14289 1405 14323 1439
rect 15021 1405 15055 1439
<< locali >>
rect 9863 2892 9897 2908
rect 9863 2816 9897 2832
rect 9951 2892 9985 2908
rect 9951 2816 9985 2832
rect 9863 2754 9897 2770
rect 9863 2678 9897 2694
rect 9951 2754 9985 2770
rect 9951 2678 9985 2694
rect 9863 2616 9897 2632
rect 9863 2540 9897 2556
rect 9951 2616 9985 2632
rect 9951 2540 9985 2556
rect 9863 2478 9897 2494
rect 9863 2402 9897 2418
rect 9951 2478 9985 2494
rect 9951 2402 9985 2418
rect 9863 2340 9897 2356
rect 9300 2287 9329 2321
rect 9363 2287 9421 2321
rect 9455 2287 9513 2321
rect 9547 2287 9605 2321
rect 9639 2287 9697 2321
rect 9731 2287 9760 2321
rect 9368 2245 9410 2287
rect 9368 2211 9376 2245
rect 9368 2177 9410 2211
rect 9368 2143 9376 2177
rect 9368 2109 9410 2143
rect 9368 2075 9376 2109
rect 9368 2059 9410 2075
rect 9444 2245 9510 2253
rect 9444 2211 9460 2245
rect 9494 2211 9510 2245
rect 9444 2178 9510 2211
rect 9444 2144 9457 2178
rect 9491 2177 9510 2178
rect 9444 2143 9460 2144
rect 9494 2143 9510 2177
rect 9444 2109 9510 2143
rect 9444 2075 9460 2109
rect 9494 2075 9510 2109
rect 9444 2057 9510 2075
rect 9364 2013 9430 2023
rect 9364 1979 9376 2013
rect 9410 2009 9430 2013
rect 9364 1975 9380 1979
rect 9414 1975 9430 2009
rect 9364 1925 9410 1941
rect 9464 1937 9510 2057
rect 9364 1891 9376 1925
rect 9364 1857 9410 1891
rect 9364 1823 9376 1857
rect 9364 1777 9410 1823
rect 9444 1925 9510 1937
rect 9444 1891 9460 1925
rect 9494 1891 9510 1925
rect 9444 1857 9510 1891
rect 9444 1823 9460 1857
rect 9494 1823 9510 1857
rect 9444 1811 9510 1823
rect 9550 2245 9616 2253
rect 9550 2211 9566 2245
rect 9600 2211 9616 2245
rect 9550 2177 9616 2211
rect 9550 2143 9566 2177
rect 9600 2143 9616 2177
rect 9550 2123 9616 2143
rect 9550 2075 9566 2123
rect 9600 2075 9616 2123
rect 9550 2057 9616 2075
rect 9650 2245 9692 2287
rect 9863 2264 9897 2280
rect 9951 2340 9985 2356
rect 9951 2264 9985 2280
rect 9684 2211 9692 2245
rect 9650 2177 9692 2211
rect 9684 2143 9692 2177
rect 9650 2109 9692 2143
rect 9863 2202 9897 2218
rect 9863 2126 9897 2142
rect 9951 2202 9985 2218
rect 9951 2126 9985 2142
rect 9684 2075 9692 2109
rect 9650 2059 9692 2075
rect 9550 1937 9596 2057
rect 9891 2049 9907 2083
rect 9941 2049 9957 2083
rect 9630 2012 9696 2023
rect 9630 2009 9650 2012
rect 9630 1975 9646 2009
rect 9684 1978 9696 2012
rect 9680 1975 9696 1978
rect 9817 2013 9866 2025
rect 9817 1979 9826 2013
rect 9860 2008 9866 2013
rect 9860 1979 10112 2008
rect 9817 1973 10112 1979
rect 9817 1966 9866 1973
rect 10077 1950 10112 1973
rect 9550 1925 9616 1937
rect 9550 1891 9566 1925
rect 9600 1891 9616 1925
rect 9550 1857 9616 1891
rect 9550 1823 9566 1857
rect 9600 1823 9616 1857
rect 9550 1811 9616 1823
rect 9650 1925 9696 1941
rect 10077 1938 10126 1950
rect 9684 1891 9696 1925
rect 9650 1857 9696 1891
rect 9818 1920 9867 1932
rect 9818 1886 9827 1920
rect 9861 1886 10028 1920
rect 10077 1904 10086 1938
rect 10120 1904 10126 1938
rect 10077 1891 10126 1904
rect 15627 1891 15661 1907
rect 9818 1873 9867 1886
rect 9684 1823 9696 1857
rect 9650 1777 9696 1823
rect 9987 1844 10028 1886
rect 10078 1845 10127 1857
rect 10078 1844 10087 1845
rect 9987 1811 10087 1844
rect 10121 1811 10127 1845
rect 9987 1810 10127 1811
rect 10078 1798 10127 1810
rect 10512 1809 10528 1843
rect 10562 1809 10578 1843
rect 11244 1809 11260 1843
rect 11294 1809 11310 1843
rect 11370 1809 11386 1843
rect 11420 1809 11436 1843
rect 12456 1809 12472 1843
rect 12506 1809 12522 1843
rect 12582 1809 12598 1843
rect 12632 1809 12648 1843
rect 13668 1809 13684 1843
rect 13718 1809 13734 1843
rect 13794 1809 13810 1843
rect 13844 1809 13860 1843
rect 14880 1809 14896 1843
rect 14930 1809 14946 1843
rect 15006 1809 15022 1843
rect 15056 1809 15072 1843
rect 15627 1815 15661 1831
rect 15715 1891 15749 1907
rect 15715 1815 15749 1831
rect 9300 1743 9329 1777
rect 9363 1743 9421 1777
rect 9455 1743 9513 1777
rect 9547 1743 9605 1777
rect 9639 1743 9697 1777
rect 9731 1743 9760 1777
rect 10484 1750 10518 1766
rect 10484 1674 10518 1690
rect 10572 1750 10606 1766
rect 10572 1674 10606 1690
rect 11216 1750 11250 1766
rect 11216 1674 11250 1690
rect 11321 1750 11355 1766
rect 11321 1674 11355 1690
rect 11430 1750 11464 1766
rect 11430 1674 11464 1690
rect 12428 1750 12462 1766
rect 12428 1674 12462 1690
rect 12532 1750 12566 1766
rect 12532 1674 12566 1690
rect 12642 1750 12676 1766
rect 12642 1674 12676 1690
rect 13640 1750 13674 1766
rect 13640 1674 13674 1690
rect 13745 1750 13779 1766
rect 13745 1674 13779 1690
rect 13854 1750 13888 1766
rect 13854 1674 13888 1690
rect 14852 1750 14886 1766
rect 14852 1674 14886 1690
rect 14959 1750 14993 1766
rect 14959 1674 14993 1690
rect 15066 1750 15100 1766
rect 15066 1674 15100 1690
rect 15627 1753 15661 1769
rect 15627 1677 15661 1693
rect 15715 1753 15749 1769
rect 15715 1677 15749 1693
rect 15811 1753 15845 1769
rect 15811 1677 15845 1693
rect 15907 1753 15941 1769
rect 15907 1677 15941 1693
rect 15540 1602 15556 1636
rect 15590 1602 15606 1636
rect 15747 1600 15763 1634
rect 15797 1600 15813 1634
rect 10839 1549 10873 1565
rect 10839 1473 10873 1489
rect 10927 1549 10961 1565
rect 10927 1473 10961 1489
rect 11571 1549 11605 1565
rect 11571 1473 11605 1489
rect 11676 1549 11710 1565
rect 11676 1473 11710 1489
rect 11783 1549 11817 1565
rect 11783 1473 11817 1489
rect 12783 1549 12817 1565
rect 12783 1473 12817 1489
rect 12887 1549 12921 1565
rect 12887 1473 12921 1489
rect 12995 1549 13029 1565
rect 12995 1473 13029 1489
rect 14121 1549 14155 1565
rect 14121 1473 14155 1489
rect 14227 1549 14261 1565
rect 14227 1473 14261 1489
rect 14333 1549 14367 1565
rect 14333 1473 14367 1489
rect 14976 1549 15010 1565
rect 14976 1473 15010 1489
rect 15065 1549 15099 1565
rect 15065 1473 15099 1489
rect 15627 1550 15661 1566
rect 15627 1474 15661 1490
rect 15715 1550 15749 1566
rect 15715 1474 15749 1490
rect 15811 1550 15845 1566
rect 15811 1474 15845 1490
rect 15907 1550 15941 1566
rect 15907 1474 15941 1490
rect 9881 1415 9897 1449
rect 9931 1415 9947 1449
rect 10867 1405 10883 1439
rect 10917 1405 10933 1439
rect 11599 1405 11615 1439
rect 11649 1405 11665 1439
rect 11723 1405 11739 1439
rect 11773 1405 11789 1439
rect 12811 1405 12827 1439
rect 12861 1405 12877 1439
rect 12935 1405 12951 1439
rect 12985 1405 13001 1439
rect 14149 1405 14165 1439
rect 14199 1405 14215 1439
rect 14273 1405 14289 1439
rect 14323 1405 14339 1439
rect 15005 1405 15021 1439
rect 15055 1405 15071 1439
rect 15627 1412 15661 1428
rect 9817 1365 9851 1381
rect 9817 1289 9851 1305
rect 9977 1365 10011 1381
rect 15627 1336 15661 1352
rect 15715 1412 15749 1428
rect 15715 1336 15749 1352
rect 9977 1289 10011 1305
rect 9817 1227 9851 1243
rect 9817 1151 9851 1167
rect 9977 1227 10011 1243
rect 9977 1151 10011 1167
rect 9817 1089 9851 1105
rect 9817 1013 9851 1029
rect 9977 1089 10011 1105
rect 9977 1013 10011 1029
rect 9817 951 9851 967
rect 9817 875 9851 891
rect 9977 951 10011 967
rect 9977 875 10011 891
rect 9817 813 9851 829
rect 9817 737 9851 753
rect 9977 813 10011 829
rect 9977 737 10011 753
rect 9817 675 9851 691
rect 9817 599 9851 615
rect 9977 675 10011 691
rect 9977 599 10011 615
rect 9817 537 9851 553
rect 9817 461 9851 477
rect 9977 537 10011 553
rect 9977 461 10011 477
rect 9817 399 9851 415
rect 9817 323 9851 339
rect 9977 399 10011 415
rect 9977 323 10011 339
<< viali >>
rect 9863 2832 9897 2892
rect 9951 2832 9985 2892
rect 9863 2694 9897 2754
rect 9951 2694 9985 2754
rect 9863 2556 9897 2616
rect 9951 2556 9985 2616
rect 9863 2418 9897 2478
rect 9951 2418 9985 2478
rect 9329 2287 9363 2321
rect 9421 2287 9455 2321
rect 9513 2287 9547 2321
rect 9605 2287 9639 2321
rect 9697 2287 9731 2321
rect 9457 2177 9491 2178
rect 9457 2144 9460 2177
rect 9460 2144 9491 2177
rect 9376 2009 9410 2013
rect 9376 1979 9380 2009
rect 9380 1979 9410 2009
rect 9566 2109 9600 2123
rect 9566 2089 9600 2109
rect 9863 2280 9897 2340
rect 9951 2280 9985 2340
rect 9863 2142 9897 2202
rect 9951 2142 9985 2202
rect 9907 2049 9941 2083
rect 9650 2009 9684 2012
rect 9650 1978 9680 2009
rect 9680 1978 9684 2009
rect 9826 1979 9860 2013
rect 9827 1886 9861 1920
rect 10086 1904 10120 1938
rect 10087 1811 10121 1845
rect 10528 1809 10562 1843
rect 11260 1809 11294 1843
rect 11386 1809 11420 1843
rect 12472 1809 12506 1843
rect 12598 1809 12632 1843
rect 13684 1809 13718 1843
rect 13810 1809 13844 1843
rect 14896 1809 14930 1843
rect 15022 1809 15056 1843
rect 15627 1831 15661 1891
rect 15715 1831 15749 1891
rect 9329 1743 9363 1777
rect 9421 1743 9455 1777
rect 9513 1743 9547 1777
rect 9605 1743 9639 1777
rect 9697 1743 9731 1777
rect 10484 1690 10518 1750
rect 10572 1690 10606 1750
rect 11216 1690 11250 1750
rect 11321 1690 11355 1750
rect 11430 1690 11464 1750
rect 12428 1690 12462 1750
rect 12532 1690 12566 1750
rect 12642 1690 12676 1750
rect 13640 1690 13674 1750
rect 13745 1690 13779 1750
rect 13854 1690 13888 1750
rect 14852 1690 14886 1750
rect 14959 1690 14993 1750
rect 15066 1690 15100 1750
rect 15627 1693 15661 1753
rect 15715 1693 15749 1753
rect 15811 1693 15845 1753
rect 15907 1693 15941 1753
rect 15556 1602 15590 1636
rect 15763 1600 15797 1634
rect 10839 1489 10873 1549
rect 10927 1489 10961 1549
rect 11571 1489 11605 1549
rect 11676 1489 11710 1549
rect 11783 1489 11817 1549
rect 12783 1489 12817 1549
rect 12887 1489 12921 1549
rect 12995 1489 13029 1549
rect 14121 1489 14155 1549
rect 14227 1489 14261 1549
rect 14333 1489 14367 1549
rect 14976 1489 15010 1549
rect 15065 1489 15099 1549
rect 15627 1490 15661 1550
rect 15715 1490 15749 1550
rect 15811 1490 15845 1550
rect 15907 1490 15941 1550
rect 9897 1415 9931 1449
rect 10883 1405 10917 1439
rect 11615 1405 11649 1439
rect 11739 1405 11773 1439
rect 12827 1405 12861 1439
rect 12951 1405 12985 1439
rect 14165 1405 14199 1439
rect 14289 1405 14323 1439
rect 15021 1405 15055 1439
rect 9817 1305 9851 1365
rect 9977 1305 10011 1365
rect 15627 1352 15661 1412
rect 15715 1352 15749 1412
rect 9817 1167 9851 1227
rect 9977 1167 10011 1227
rect 9817 1029 9851 1089
rect 9977 1029 10011 1089
rect 9817 891 9851 951
rect 9977 891 10011 951
rect 9817 753 9851 813
rect 9977 753 10011 813
rect 9817 615 9851 675
rect 9977 615 10011 675
rect 9817 477 9851 537
rect 9977 477 10011 537
rect 9817 339 9851 399
rect 9977 339 10011 399
<< metal1 >>
rect 9963 2937 10053 2953
rect 9963 2926 9982 2937
rect 9857 2892 9903 2904
rect 9857 2832 9863 2892
rect 9897 2832 9903 2892
rect 9857 2754 9903 2832
rect 9945 2892 9982 2926
rect 9945 2832 9951 2892
rect 10034 2885 10053 2937
rect 9985 2870 10053 2885
rect 9985 2832 9991 2870
rect 9945 2820 9991 2832
rect 9857 2694 9863 2754
rect 9897 2694 9903 2754
rect 9857 2682 9903 2694
rect 9945 2754 9991 2766
rect 9945 2694 9951 2754
rect 9985 2694 9991 2754
rect 9857 2616 9903 2628
rect 9857 2556 9863 2616
rect 9897 2556 9903 2616
rect 9857 2478 9903 2556
rect 9945 2616 9991 2694
rect 9945 2556 9951 2616
rect 9985 2556 9991 2616
rect 9945 2544 9991 2556
rect 9857 2418 9863 2478
rect 9897 2418 9903 2478
rect 9857 2406 9903 2418
rect 9945 2478 9991 2490
rect 9945 2418 9951 2478
rect 9985 2418 9991 2478
rect 9300 2332 9760 2352
rect 9300 2321 9365 2332
rect 9300 2287 9329 2321
rect 9363 2287 9365 2321
rect 9300 2280 9365 2287
rect 9417 2331 9640 2332
rect 9417 2321 9496 2331
rect 9548 2321 9640 2331
rect 9417 2287 9421 2321
rect 9455 2287 9496 2321
rect 9548 2287 9605 2321
rect 9639 2287 9640 2321
rect 9417 2280 9496 2287
rect 9300 2279 9496 2280
rect 9548 2280 9640 2287
rect 9692 2321 9760 2332
rect 9692 2287 9697 2321
rect 9731 2287 9760 2321
rect 9692 2280 9760 2287
rect 9548 2279 9760 2280
rect 9300 2256 9760 2279
rect 9857 2340 9903 2352
rect 9857 2280 9863 2340
rect 9897 2280 9903 2340
rect 9857 2202 9903 2280
rect 9945 2340 9991 2418
rect 9945 2280 9951 2340
rect 9985 2280 9991 2340
rect 9945 2268 9991 2280
rect 9445 2178 9817 2185
rect 9445 2144 9457 2178
rect 9491 2157 9817 2178
rect 9491 2144 9503 2157
rect 9445 2137 9503 2144
rect 9550 2123 9617 2129
rect 9550 2089 9566 2123
rect 9600 2110 9617 2123
rect 9600 2089 9761 2110
rect 9550 2082 9761 2089
rect 9630 2021 9696 2023
rect 9368 2016 9422 2020
rect 9367 2013 9422 2016
rect 9238 1979 9376 2013
rect 9410 1979 9422 2013
rect 9367 1976 9422 1979
rect 9367 1972 9421 1976
rect 9630 1969 9638 2021
rect 9690 1969 9696 2021
rect 9630 1968 9696 1969
rect 9733 1938 9761 2082
rect 9789 2025 9817 2157
rect 9857 2142 9863 2202
rect 9897 2142 9903 2202
rect 9857 2130 9903 2142
rect 9945 2202 10027 2214
rect 9945 2142 9951 2202
rect 9985 2142 10027 2202
rect 9945 2130 10027 2142
rect 9895 2083 9953 2089
rect 9895 2049 9907 2083
rect 9941 2049 9953 2083
rect 9895 2043 9953 2049
rect 9789 2013 9866 2025
rect 9789 1979 9826 2013
rect 9860 1979 9866 2013
rect 9817 1966 9866 1979
rect 9733 1920 9867 1938
rect 9733 1910 9827 1920
rect 9818 1886 9827 1910
rect 9861 1886 9867 1920
rect 9818 1873 9867 1886
rect 9300 1786 9760 1808
rect 9300 1777 9383 1786
rect 9435 1777 9503 1786
rect 9555 1777 9646 1786
rect 9698 1777 9760 1786
rect 9300 1743 9329 1777
rect 9363 1743 9383 1777
rect 9455 1743 9503 1777
rect 9555 1743 9605 1777
rect 9639 1743 9646 1777
rect 9731 1743 9760 1777
rect 9300 1734 9383 1743
rect 9435 1734 9503 1743
rect 9555 1734 9646 1743
rect 9698 1734 9760 1743
rect 9300 1712 9760 1734
rect 9895 1643 9943 2043
rect 9275 1596 9943 1643
rect 9895 1455 9943 1596
rect 9885 1449 9943 1455
rect 9644 1443 9709 1444
rect 9644 1440 9650 1443
rect 9256 1393 9650 1440
rect 9644 1391 9650 1393
rect 9702 1391 9709 1443
rect 9885 1415 9897 1449
rect 9931 1415 9943 1449
rect 9885 1409 9943 1415
rect 9981 1640 10027 2130
rect 15695 2010 15785 2026
rect 15695 1999 15714 2010
rect 15620 1958 15714 1999
rect 15766 1958 15785 2010
rect 10077 1943 10126 1950
rect 10077 1938 10696 1943
rect 10077 1904 10086 1938
rect 10120 1904 10696 1938
rect 10077 1896 10696 1904
rect 10077 1891 10126 1896
rect 10078 1849 10127 1857
rect 10647 1849 10696 1896
rect 15620 1940 15785 1958
rect 15620 1894 15667 1940
rect 15621 1891 15667 1894
rect 10078 1845 10579 1849
rect 10078 1811 10087 1845
rect 10121 1843 10579 1845
rect 10121 1811 10528 1843
rect 10078 1809 10528 1811
rect 10562 1809 10579 1843
rect 10078 1803 10579 1809
rect 10647 1843 15068 1849
rect 10647 1809 11260 1843
rect 11294 1809 11386 1843
rect 11420 1809 12472 1843
rect 12506 1809 12598 1843
rect 12632 1809 13684 1843
rect 13718 1809 13810 1843
rect 13844 1809 14896 1843
rect 14930 1809 15022 1843
rect 15056 1809 15068 1843
rect 15621 1831 15627 1891
rect 15661 1831 15667 1891
rect 15621 1819 15667 1831
rect 15709 1891 15755 1903
rect 15709 1831 15715 1891
rect 15749 1831 15755 1891
rect 15709 1822 15755 1831
rect 10647 1803 15068 1809
rect 10078 1802 10567 1803
rect 10647 1802 11093 1803
rect 10078 1798 10127 1802
rect 15709 1793 15947 1822
rect 10478 1754 10524 1762
rect 10455 1753 10534 1754
rect 10455 1689 10462 1753
rect 10526 1689 10534 1753
rect 10566 1750 10612 1762
rect 11210 1754 11256 1762
rect 10566 1690 10572 1750
rect 10606 1690 10612 1750
rect 10478 1678 10524 1689
rect 10566 1640 10612 1690
rect 11187 1753 11266 1754
rect 11187 1689 11194 1753
rect 11258 1689 11266 1753
rect 11315 1750 11361 1762
rect 11424 1754 11470 1762
rect 12422 1754 12468 1762
rect 11315 1690 11321 1750
rect 11355 1690 11361 1750
rect 11210 1678 11256 1689
rect 11315 1640 11361 1690
rect 11414 1753 11493 1754
rect 11414 1689 11422 1753
rect 11486 1689 11493 1753
rect 12399 1753 12478 1754
rect 12399 1689 12406 1753
rect 12470 1689 12478 1753
rect 12526 1750 12572 1762
rect 12636 1754 12682 1762
rect 13634 1754 13680 1762
rect 12526 1690 12532 1750
rect 12566 1690 12572 1750
rect 11424 1678 11470 1689
rect 12422 1678 12468 1689
rect 12526 1640 12572 1690
rect 12626 1753 12705 1754
rect 12626 1689 12634 1753
rect 12698 1689 12705 1753
rect 13611 1753 13690 1754
rect 13611 1689 13618 1753
rect 13682 1689 13690 1753
rect 13739 1750 13785 1762
rect 13848 1754 13894 1762
rect 14846 1754 14892 1762
rect 13739 1690 13745 1750
rect 13779 1690 13785 1750
rect 12636 1678 12682 1689
rect 13634 1678 13680 1689
rect 13739 1640 13785 1690
rect 13838 1753 13917 1754
rect 13838 1689 13846 1753
rect 13910 1689 13917 1753
rect 14823 1753 14902 1754
rect 14823 1689 14830 1753
rect 14894 1689 14902 1753
rect 14953 1750 14999 1762
rect 15060 1754 15106 1762
rect 14953 1690 14959 1750
rect 14993 1690 14999 1750
rect 13848 1678 13894 1689
rect 14846 1678 14892 1689
rect 14953 1640 14999 1690
rect 15050 1753 15129 1754
rect 15050 1689 15058 1753
rect 15122 1689 15129 1753
rect 15621 1753 15667 1765
rect 15621 1693 15627 1753
rect 15661 1693 15667 1753
rect 15060 1678 15106 1689
rect 15621 1681 15667 1693
rect 15709 1753 15755 1793
rect 15709 1693 15715 1753
rect 15749 1693 15755 1753
rect 15709 1681 15755 1693
rect 15783 1753 15873 1765
rect 15783 1749 15811 1753
rect 15845 1749 15873 1753
rect 15783 1697 15802 1749
rect 15854 1697 15873 1749
rect 15783 1693 15811 1697
rect 15845 1693 15873 1697
rect 15783 1681 15873 1693
rect 15901 1753 15947 1793
rect 15901 1693 15907 1753
rect 15941 1693 15947 1753
rect 15901 1681 15947 1693
rect 15540 1640 15606 1642
rect 9981 1636 15606 1640
rect 9981 1602 15556 1636
rect 15590 1602 15606 1636
rect 9981 1598 15606 1602
rect 9981 1377 10027 1598
rect 10833 1551 10879 1561
rect 10811 1487 10820 1551
rect 10884 1487 10893 1551
rect 10811 1486 10893 1487
rect 10921 1549 10967 1598
rect 11565 1551 11611 1561
rect 10921 1489 10927 1549
rect 10961 1489 10967 1549
rect 10833 1477 10879 1486
rect 10921 1477 10967 1489
rect 11543 1487 11552 1551
rect 11616 1487 11625 1551
rect 11543 1486 11625 1487
rect 11670 1549 11716 1598
rect 11777 1551 11823 1561
rect 12777 1551 12823 1561
rect 11670 1489 11676 1549
rect 11710 1489 11716 1549
rect 11565 1477 11611 1486
rect 11670 1477 11716 1489
rect 11763 1487 11772 1551
rect 11836 1487 11845 1551
rect 11763 1486 11845 1487
rect 12755 1487 12764 1551
rect 12828 1487 12837 1551
rect 12755 1486 12837 1487
rect 12881 1549 12927 1598
rect 12989 1551 13035 1561
rect 14115 1551 14161 1561
rect 12881 1489 12887 1549
rect 12921 1489 12927 1549
rect 11777 1477 11823 1486
rect 12777 1477 12823 1486
rect 12881 1477 12927 1489
rect 12975 1487 12984 1551
rect 13048 1487 13057 1551
rect 12975 1486 13057 1487
rect 14093 1487 14102 1551
rect 14166 1487 14175 1551
rect 14093 1486 14175 1487
rect 14221 1549 14267 1598
rect 14327 1551 14373 1561
rect 14221 1489 14227 1549
rect 14261 1489 14267 1549
rect 12989 1477 13035 1486
rect 14115 1477 14161 1486
rect 14221 1477 14267 1489
rect 14313 1487 14322 1551
rect 14386 1487 14395 1551
rect 14313 1486 14395 1487
rect 14970 1549 15016 1598
rect 15544 1596 15606 1598
rect 15639 1633 15667 1681
rect 15751 1634 15933 1640
rect 15751 1633 15763 1634
rect 15639 1604 15763 1633
rect 15639 1562 15667 1604
rect 15751 1600 15763 1604
rect 15797 1600 15933 1634
rect 15751 1594 15933 1600
rect 15059 1551 15105 1561
rect 14970 1489 14976 1549
rect 15010 1489 15016 1549
rect 14327 1477 14373 1486
rect 14970 1477 15016 1489
rect 15045 1487 15054 1551
rect 15118 1487 15127 1551
rect 15045 1486 15127 1487
rect 15621 1550 15667 1562
rect 15621 1490 15627 1550
rect 15661 1490 15667 1550
rect 15059 1477 15105 1486
rect 15621 1478 15667 1490
rect 15709 1550 15755 1562
rect 15709 1490 15715 1550
rect 15749 1490 15755 1550
rect 15709 1450 15755 1490
rect 15783 1550 15873 1562
rect 15783 1546 15811 1550
rect 15845 1546 15873 1550
rect 15783 1494 15802 1546
rect 15854 1494 15873 1546
rect 15783 1490 15811 1494
rect 15845 1490 15873 1494
rect 15783 1478 15873 1490
rect 15901 1550 15947 1562
rect 15901 1490 15907 1550
rect 15941 1490 15947 1550
rect 15901 1450 15947 1490
rect 10131 1391 10138 1443
rect 10190 1441 10196 1443
rect 10871 1441 10929 1445
rect 10190 1439 10929 1441
rect 10190 1405 10883 1439
rect 10917 1405 10929 1439
rect 10190 1394 10929 1405
rect 11603 1439 12997 1445
rect 11603 1405 11615 1439
rect 11649 1405 11739 1439
rect 11773 1405 12827 1439
rect 12861 1405 12951 1439
rect 12985 1405 12997 1439
rect 11603 1399 12997 1405
rect 14153 1439 14335 1445
rect 14153 1405 14165 1439
rect 14199 1405 14289 1439
rect 14323 1405 14335 1439
rect 14153 1399 14335 1405
rect 15009 1439 15067 1445
rect 15009 1405 15021 1439
rect 15055 1405 15067 1439
rect 10190 1391 10196 1394
rect 10131 1390 10196 1391
rect 10871 1389 10929 1394
rect 9811 1365 9857 1377
rect 9811 1305 9817 1365
rect 9851 1305 9857 1365
rect 9811 1227 9857 1305
rect 9971 1365 10027 1377
rect 9971 1305 9977 1365
rect 10011 1305 10027 1365
rect 9971 1293 10027 1305
rect 9811 1167 9817 1227
rect 9851 1167 9857 1227
rect 9811 1155 9857 1167
rect 9971 1227 10017 1239
rect 9971 1167 9977 1227
rect 10011 1167 10017 1227
rect 9811 1089 9857 1101
rect 9811 1029 9817 1089
rect 9851 1029 9857 1089
rect 9811 951 9857 1029
rect 9971 1089 10017 1167
rect 9971 1029 9977 1089
rect 10011 1029 10017 1089
rect 9971 1017 10017 1029
rect 9811 891 9817 951
rect 9851 891 9857 951
rect 9811 879 9857 891
rect 9971 951 10017 963
rect 9971 891 9977 951
rect 10011 891 10017 951
rect 9811 813 9857 825
rect 9811 753 9817 813
rect 9851 753 9857 813
rect 9811 675 9857 753
rect 9971 813 10017 891
rect 9971 753 9977 813
rect 10011 753 10017 813
rect 9971 741 10017 753
rect 9811 615 9817 675
rect 9851 615 9857 675
rect 9811 603 9857 615
rect 9971 675 10017 687
rect 9971 615 9977 675
rect 10011 615 10017 675
rect 9811 537 9857 549
rect 9811 477 9817 537
rect 9851 477 9857 537
rect 9811 399 9857 477
rect 9971 537 10017 615
rect 9971 477 9977 537
rect 10011 477 10017 537
rect 9971 465 10017 477
rect 9811 339 9817 399
rect 9851 339 9857 399
rect 9971 399 10017 411
rect 9971 375 9977 399
rect 9811 327 9857 339
rect 9932 359 9977 375
rect 10011 375 10017 399
rect 10011 359 10039 375
rect 9932 307 9968 359
rect 10020 307 10039 359
rect 9932 291 10039 307
rect 11727 268 11785 1399
rect 14153 268 14211 1399
rect 15009 267 15067 1405
rect 15621 1412 15667 1424
rect 15621 1352 15627 1412
rect 15661 1352 15667 1412
rect 15621 1300 15667 1352
rect 15709 1421 15947 1450
rect 15709 1412 15755 1421
rect 15709 1352 15715 1412
rect 15749 1352 15755 1412
rect 15709 1340 15755 1352
rect 15621 1284 15782 1300
rect 15621 1232 15711 1284
rect 15763 1232 15782 1284
rect 15621 1216 15782 1232
<< via1 >>
rect 9982 2892 10034 2937
rect 9982 2885 9985 2892
rect 9985 2885 10034 2892
rect 9365 2280 9417 2332
rect 9496 2321 9548 2331
rect 9496 2287 9513 2321
rect 9513 2287 9547 2321
rect 9547 2287 9548 2321
rect 9496 2279 9548 2287
rect 9640 2280 9692 2332
rect 9638 2012 9690 2021
rect 9638 1978 9650 2012
rect 9650 1978 9684 2012
rect 9684 1978 9690 2012
rect 9638 1969 9690 1978
rect 9383 1777 9435 1786
rect 9503 1777 9555 1786
rect 9646 1777 9698 1786
rect 9383 1743 9421 1777
rect 9421 1743 9435 1777
rect 9503 1743 9513 1777
rect 9513 1743 9547 1777
rect 9547 1743 9555 1777
rect 9646 1743 9697 1777
rect 9697 1743 9698 1777
rect 9383 1734 9435 1743
rect 9503 1734 9555 1743
rect 9646 1734 9698 1743
rect 9650 1391 9702 1443
rect 15714 1958 15766 2010
rect 10462 1750 10526 1753
rect 10462 1690 10484 1750
rect 10484 1690 10518 1750
rect 10518 1690 10526 1750
rect 10462 1689 10526 1690
rect 11194 1750 11258 1753
rect 11194 1690 11216 1750
rect 11216 1690 11250 1750
rect 11250 1690 11258 1750
rect 11194 1689 11258 1690
rect 11422 1750 11486 1753
rect 11422 1690 11430 1750
rect 11430 1690 11464 1750
rect 11464 1690 11486 1750
rect 11422 1689 11486 1690
rect 12406 1750 12470 1753
rect 12406 1690 12428 1750
rect 12428 1690 12462 1750
rect 12462 1690 12470 1750
rect 12406 1689 12470 1690
rect 12634 1750 12698 1753
rect 12634 1690 12642 1750
rect 12642 1690 12676 1750
rect 12676 1690 12698 1750
rect 12634 1689 12698 1690
rect 13618 1750 13682 1753
rect 13618 1690 13640 1750
rect 13640 1690 13674 1750
rect 13674 1690 13682 1750
rect 13618 1689 13682 1690
rect 13846 1750 13910 1753
rect 13846 1690 13854 1750
rect 13854 1690 13888 1750
rect 13888 1690 13910 1750
rect 13846 1689 13910 1690
rect 14830 1750 14894 1753
rect 14830 1690 14852 1750
rect 14852 1690 14886 1750
rect 14886 1690 14894 1750
rect 14830 1689 14894 1690
rect 15058 1750 15122 1753
rect 15058 1690 15066 1750
rect 15066 1690 15100 1750
rect 15100 1690 15122 1750
rect 15058 1689 15122 1690
rect 15802 1697 15811 1749
rect 15811 1697 15845 1749
rect 15845 1697 15854 1749
rect 10820 1549 10884 1551
rect 10820 1489 10839 1549
rect 10839 1489 10873 1549
rect 10873 1489 10884 1549
rect 10820 1487 10884 1489
rect 11552 1549 11616 1551
rect 11552 1489 11571 1549
rect 11571 1489 11605 1549
rect 11605 1489 11616 1549
rect 11552 1487 11616 1489
rect 11772 1549 11836 1551
rect 11772 1489 11783 1549
rect 11783 1489 11817 1549
rect 11817 1489 11836 1549
rect 11772 1487 11836 1489
rect 12764 1549 12828 1551
rect 12764 1489 12783 1549
rect 12783 1489 12817 1549
rect 12817 1489 12828 1549
rect 12764 1487 12828 1489
rect 12984 1549 13048 1551
rect 12984 1489 12995 1549
rect 12995 1489 13029 1549
rect 13029 1489 13048 1549
rect 12984 1487 13048 1489
rect 14102 1549 14166 1551
rect 14102 1489 14121 1549
rect 14121 1489 14155 1549
rect 14155 1489 14166 1549
rect 14102 1487 14166 1489
rect 14322 1549 14386 1551
rect 14322 1489 14333 1549
rect 14333 1489 14367 1549
rect 14367 1489 14386 1549
rect 14322 1487 14386 1489
rect 15054 1549 15118 1551
rect 15054 1489 15065 1549
rect 15065 1489 15099 1549
rect 15099 1489 15118 1549
rect 15054 1487 15118 1489
rect 15802 1494 15811 1546
rect 15811 1494 15845 1546
rect 15845 1494 15854 1546
rect 10138 1391 10190 1443
rect 9968 339 9977 359
rect 9977 339 10011 359
rect 10011 339 10020 359
rect 9968 307 10020 339
rect 15711 1232 15763 1284
<< metal2 >>
rect 9971 2939 10045 2943
rect 9971 2883 9980 2939
rect 10036 2883 10045 2939
rect 9971 2879 10045 2883
rect 9363 2334 9419 2343
rect 9363 2269 9419 2278
rect 9494 2333 9550 2342
rect 9494 2268 9550 2277
rect 9638 2334 9694 2343
rect 9638 2269 9694 2278
rect 9630 1969 9638 2021
rect 9690 1969 9696 2021
rect 9630 1968 9696 1969
rect 15703 2012 15777 2016
rect 9648 1892 9694 1968
rect 15703 1956 15712 2012
rect 15768 1956 15777 2012
rect 15703 1952 15777 1956
rect 9648 1846 9887 1892
rect 9381 1788 9437 1797
rect 9381 1723 9437 1732
rect 9501 1788 9557 1797
rect 9501 1723 9557 1732
rect 9644 1788 9700 1797
rect 9644 1723 9700 1732
rect 9644 1443 9709 1444
rect 9644 1391 9650 1443
rect 9702 1440 9709 1443
rect 9841 1440 9887 1846
rect 10455 1753 10534 1754
rect 11187 1753 11266 1754
rect 11414 1753 11493 1754
rect 12399 1753 12478 1754
rect 12626 1753 12705 1754
rect 13611 1753 13690 1754
rect 13838 1753 13917 1754
rect 14823 1753 14902 1754
rect 15050 1753 15129 1754
rect 10452 1689 10462 1753
rect 10526 1689 10535 1753
rect 11184 1689 11194 1753
rect 11258 1689 11267 1753
rect 11413 1689 11422 1753
rect 11486 1689 11496 1753
rect 12396 1689 12406 1753
rect 12470 1689 12479 1753
rect 12625 1689 12634 1753
rect 12698 1689 12708 1753
rect 13608 1689 13618 1753
rect 13682 1689 13691 1753
rect 13837 1689 13846 1753
rect 13910 1689 13920 1753
rect 14820 1689 14830 1753
rect 14894 1689 14903 1753
rect 15049 1689 15058 1753
rect 15122 1689 15132 1753
rect 15791 1751 15865 1755
rect 15791 1695 15800 1751
rect 15856 1695 15865 1751
rect 15791 1691 15865 1695
rect 10811 1487 10820 1551
rect 10884 1487 10893 1551
rect 10811 1486 10893 1487
rect 11543 1487 11552 1551
rect 11616 1487 11625 1551
rect 11543 1486 11625 1487
rect 11763 1487 11772 1551
rect 11836 1487 11845 1551
rect 11763 1486 11845 1487
rect 12755 1487 12764 1551
rect 12828 1487 12837 1551
rect 12755 1486 12837 1487
rect 12975 1487 12984 1551
rect 13048 1487 13057 1551
rect 12975 1486 13057 1487
rect 14093 1487 14102 1551
rect 14166 1487 14175 1551
rect 14093 1486 14175 1487
rect 14313 1487 14322 1551
rect 14386 1487 14395 1551
rect 14313 1486 14395 1487
rect 15045 1487 15054 1551
rect 15118 1487 15127 1551
rect 15791 1548 15865 1552
rect 15791 1492 15800 1548
rect 15856 1492 15865 1548
rect 15791 1488 15865 1492
rect 15045 1486 15127 1487
rect 10131 1440 10138 1443
rect 9702 1394 10138 1440
rect 9702 1391 9709 1394
rect 10131 1391 10138 1394
rect 10190 1391 10196 1443
rect 10131 1390 10196 1391
rect 15700 1286 15774 1290
rect 15700 1230 15709 1286
rect 15765 1230 15774 1286
rect 15700 1226 15774 1230
rect 9957 361 10031 365
rect 9957 305 9966 361
rect 10022 305 10031 361
rect 9957 301 10031 305
<< via2 >>
rect 9980 2937 10036 2939
rect 9980 2885 9982 2937
rect 9982 2885 10034 2937
rect 10034 2885 10036 2937
rect 9980 2883 10036 2885
rect 9363 2332 9419 2334
rect 9363 2280 9365 2332
rect 9365 2280 9417 2332
rect 9417 2280 9419 2332
rect 9363 2278 9419 2280
rect 9494 2331 9550 2333
rect 9494 2279 9496 2331
rect 9496 2279 9548 2331
rect 9548 2279 9550 2331
rect 9494 2277 9550 2279
rect 9638 2332 9694 2334
rect 9638 2280 9640 2332
rect 9640 2280 9692 2332
rect 9692 2280 9694 2332
rect 9638 2278 9694 2280
rect 15712 2010 15768 2012
rect 15712 1958 15714 2010
rect 15714 1958 15766 2010
rect 15766 1958 15768 2010
rect 15712 1956 15768 1958
rect 9381 1786 9437 1788
rect 9381 1734 9383 1786
rect 9383 1734 9435 1786
rect 9435 1734 9437 1786
rect 9381 1732 9437 1734
rect 9501 1786 9557 1788
rect 9501 1734 9503 1786
rect 9503 1734 9555 1786
rect 9555 1734 9557 1786
rect 9501 1732 9557 1734
rect 9644 1786 9700 1788
rect 9644 1734 9646 1786
rect 9646 1734 9698 1786
rect 9698 1734 9700 1786
rect 9644 1732 9700 1734
rect 10462 1689 10526 1753
rect 11194 1689 11258 1753
rect 11422 1689 11486 1753
rect 12406 1689 12470 1753
rect 12634 1689 12698 1753
rect 13618 1689 13682 1753
rect 13846 1689 13910 1753
rect 14830 1689 14894 1753
rect 15058 1689 15122 1753
rect 15800 1749 15856 1751
rect 15800 1697 15802 1749
rect 15802 1697 15854 1749
rect 15854 1697 15856 1749
rect 15800 1695 15856 1697
rect 10820 1487 10884 1551
rect 11552 1487 11616 1551
rect 11772 1487 11836 1551
rect 12764 1487 12828 1551
rect 12984 1487 13048 1551
rect 14102 1487 14166 1551
rect 14322 1487 14386 1551
rect 15054 1487 15118 1551
rect 15800 1546 15856 1548
rect 15800 1494 15802 1546
rect 15802 1494 15854 1546
rect 15854 1494 15856 1546
rect 15800 1492 15856 1494
rect 15709 1284 15765 1286
rect 15709 1232 15711 1284
rect 15711 1232 15763 1284
rect 15763 1232 15765 1284
rect 15709 1230 15765 1232
rect 9966 359 10022 361
rect 9966 307 9968 359
rect 9968 307 10020 359
rect 10020 307 10022 359
rect 9966 305 10022 307
<< metal3 >>
rect 9945 2943 10071 2953
rect 9945 2879 9976 2943
rect 10040 2938 10071 2943
rect 10040 2936 10641 2938
rect 10040 2879 10073 2936
rect 9945 2872 10073 2879
rect 10137 2872 10153 2936
rect 10217 2872 10233 2936
rect 10297 2872 10313 2936
rect 10377 2872 10393 2936
rect 10457 2872 10473 2936
rect 10537 2872 10641 2936
rect 9945 2870 10641 2872
rect 10701 2936 15615 2938
rect 10701 2872 10805 2936
rect 10869 2872 10885 2936
rect 10949 2872 10965 2936
rect 11029 2872 11045 2936
rect 11109 2872 11125 2936
rect 11189 2872 11205 2936
rect 11269 2872 11411 2936
rect 11475 2872 11491 2936
rect 11555 2872 11571 2936
rect 11635 2872 11651 2936
rect 11715 2872 11731 2936
rect 11795 2872 11811 2936
rect 11875 2872 12017 2936
rect 12081 2872 12097 2936
rect 12161 2872 12177 2936
rect 12241 2872 12257 2936
rect 12321 2872 12337 2936
rect 12401 2872 12417 2936
rect 12481 2872 12623 2936
rect 12687 2872 12703 2936
rect 12767 2872 12783 2936
rect 12847 2872 12863 2936
rect 12927 2872 12943 2936
rect 13007 2872 13023 2936
rect 13087 2872 13229 2936
rect 13293 2872 13309 2936
rect 13373 2872 13389 2936
rect 13453 2872 13469 2936
rect 13533 2872 13549 2936
rect 13613 2872 13629 2936
rect 13693 2872 13835 2936
rect 13899 2872 13915 2936
rect 13979 2872 13995 2936
rect 14059 2872 14075 2936
rect 14139 2872 14155 2936
rect 14219 2872 14235 2936
rect 14299 2872 14441 2936
rect 14505 2872 14521 2936
rect 14585 2872 14601 2936
rect 14665 2872 14681 2936
rect 14745 2872 14761 2936
rect 14825 2872 14841 2936
rect 14905 2872 15047 2936
rect 15111 2872 15127 2936
rect 15191 2872 15207 2936
rect 15271 2872 15287 2936
rect 15351 2872 15367 2936
rect 15431 2872 15447 2936
rect 15511 2872 15615 2936
rect 10701 2870 15615 2872
rect 9969 2716 10035 2806
rect 9969 2652 9970 2716
rect 10034 2652 10035 2716
rect 9969 2636 10035 2652
rect 9969 2572 9970 2636
rect 10034 2572 10035 2636
rect 9969 2556 10035 2572
rect 9969 2492 9970 2556
rect 10034 2492 10035 2556
rect 9969 2476 10035 2492
rect 9969 2412 9970 2476
rect 10034 2412 10035 2476
rect 9969 2396 10035 2412
rect 9318 2352 9462 2353
rect 9593 2352 9737 2353
rect 9318 2338 9737 2352
rect 9318 2274 9359 2338
rect 9423 2337 9634 2338
rect 9423 2274 9490 2337
rect 9318 2273 9490 2274
rect 9554 2274 9634 2337
rect 9698 2274 9737 2338
rect 9554 2273 9737 2274
rect 9318 2257 9737 2273
rect 9969 2332 9970 2396
rect 10034 2332 10035 2396
rect 9969 2316 10035 2332
rect 9449 2256 9593 2257
rect 9969 2252 9970 2316
rect 10034 2252 10035 2316
rect 9969 2236 10035 2252
rect 9969 2172 9970 2236
rect 10034 2172 10035 2236
rect 9969 2156 10035 2172
rect 9969 2092 9970 2156
rect 10034 2092 10035 2156
rect 9969 2076 10035 2092
rect 9969 2012 9970 2076
rect 10034 2012 10035 2076
rect 9969 1996 10035 2012
rect 9969 1932 9970 1996
rect 10034 1932 10035 1996
rect 9484 1807 9576 1808
rect 9336 1792 9743 1807
rect 9336 1728 9377 1792
rect 9441 1728 9497 1792
rect 9561 1728 9640 1792
rect 9704 1728 9743 1792
rect 9336 1711 9743 1728
rect 9969 1778 10035 1932
rect 10095 1778 10155 2810
rect 10215 1840 10275 2870
rect 10335 1778 10395 2810
rect 10455 1840 10515 2870
rect 10575 2716 10641 2806
rect 10575 2652 10576 2716
rect 10640 2652 10641 2716
rect 10575 2636 10641 2652
rect 10575 2572 10576 2636
rect 10640 2572 10641 2636
rect 10575 2556 10641 2572
rect 10575 2492 10576 2556
rect 10640 2492 10641 2556
rect 10575 2476 10641 2492
rect 10575 2412 10576 2476
rect 10640 2412 10641 2476
rect 10575 2396 10641 2412
rect 10575 2332 10576 2396
rect 10640 2332 10641 2396
rect 10575 2316 10641 2332
rect 10575 2252 10576 2316
rect 10640 2252 10641 2316
rect 10575 2236 10641 2252
rect 10575 2172 10576 2236
rect 10640 2172 10641 2236
rect 10575 2156 10641 2172
rect 10575 2092 10576 2156
rect 10640 2092 10641 2156
rect 10575 2076 10641 2092
rect 10575 2012 10576 2076
rect 10640 2012 10641 2076
rect 10575 1996 10641 2012
rect 10575 1932 10576 1996
rect 10640 1932 10641 1996
rect 10575 1778 10641 1932
rect 9969 1776 10641 1778
rect 9969 1712 10073 1776
rect 10137 1712 10153 1776
rect 10217 1712 10233 1776
rect 10297 1712 10313 1776
rect 10377 1712 10393 1776
rect 10457 1753 10473 1776
rect 10457 1712 10462 1753
rect 10537 1712 10641 1776
rect 9969 1710 10462 1712
rect 10452 1689 10462 1710
rect 10526 1710 10641 1712
rect 10701 2716 10767 2806
rect 10701 2652 10702 2716
rect 10766 2652 10767 2716
rect 10701 2636 10767 2652
rect 10701 2572 10702 2636
rect 10766 2572 10767 2636
rect 10701 2556 10767 2572
rect 10701 2492 10702 2556
rect 10766 2492 10767 2556
rect 10701 2476 10767 2492
rect 10701 2412 10702 2476
rect 10766 2412 10767 2476
rect 10701 2396 10767 2412
rect 10701 2332 10702 2396
rect 10766 2332 10767 2396
rect 10701 2316 10767 2332
rect 10701 2252 10702 2316
rect 10766 2252 10767 2316
rect 10701 2236 10767 2252
rect 10701 2172 10702 2236
rect 10766 2172 10767 2236
rect 10701 2156 10767 2172
rect 10701 2092 10702 2156
rect 10766 2092 10767 2156
rect 10701 2076 10767 2092
rect 10701 2012 10702 2076
rect 10766 2012 10767 2076
rect 10701 1996 10767 2012
rect 10701 1932 10702 1996
rect 10766 1932 10767 1996
rect 10701 1778 10767 1932
rect 10827 1778 10887 2810
rect 10947 1840 11007 2870
rect 11067 1778 11127 2810
rect 11187 1840 11247 2870
rect 11307 2716 11373 2806
rect 11307 2652 11308 2716
rect 11372 2652 11373 2716
rect 11307 2636 11373 2652
rect 11307 2572 11308 2636
rect 11372 2572 11373 2636
rect 11307 2556 11373 2572
rect 11307 2492 11308 2556
rect 11372 2492 11373 2556
rect 11307 2476 11373 2492
rect 11307 2412 11308 2476
rect 11372 2412 11373 2476
rect 11307 2396 11373 2412
rect 11307 2332 11308 2396
rect 11372 2332 11373 2396
rect 11307 2316 11373 2332
rect 11307 2252 11308 2316
rect 11372 2252 11373 2316
rect 11307 2236 11373 2252
rect 11307 2172 11308 2236
rect 11372 2172 11373 2236
rect 11307 2156 11373 2172
rect 11307 2092 11308 2156
rect 11372 2092 11373 2156
rect 11307 2076 11373 2092
rect 11307 2012 11308 2076
rect 11372 2012 11373 2076
rect 11307 1996 11373 2012
rect 11307 1932 11308 1996
rect 11372 1932 11373 1996
rect 11307 1778 11373 1932
rect 11433 1840 11493 2870
rect 11553 1778 11613 2810
rect 11673 1840 11733 2870
rect 11793 1778 11853 2810
rect 11913 2716 11979 2806
rect 11913 2652 11914 2716
rect 11978 2652 11979 2716
rect 11913 2636 11979 2652
rect 11913 2572 11914 2636
rect 11978 2572 11979 2636
rect 11913 2556 11979 2572
rect 11913 2492 11914 2556
rect 11978 2492 11979 2556
rect 11913 2476 11979 2492
rect 11913 2412 11914 2476
rect 11978 2412 11979 2476
rect 11913 2396 11979 2412
rect 11913 2332 11914 2396
rect 11978 2332 11979 2396
rect 11913 2316 11979 2332
rect 11913 2252 11914 2316
rect 11978 2252 11979 2316
rect 11913 2236 11979 2252
rect 11913 2172 11914 2236
rect 11978 2172 11979 2236
rect 11913 2156 11979 2172
rect 11913 2092 11914 2156
rect 11978 2092 11979 2156
rect 11913 2076 11979 2092
rect 11913 2012 11914 2076
rect 11978 2012 11979 2076
rect 11913 1996 11979 2012
rect 11913 1932 11914 1996
rect 11978 1932 11979 1996
rect 11913 1778 11979 1932
rect 12039 1778 12099 2810
rect 12159 1840 12219 2870
rect 12279 1778 12339 2810
rect 12399 1840 12459 2870
rect 12519 2716 12585 2806
rect 12519 2652 12520 2716
rect 12584 2652 12585 2716
rect 12519 2636 12585 2652
rect 12519 2572 12520 2636
rect 12584 2572 12585 2636
rect 12519 2556 12585 2572
rect 12519 2492 12520 2556
rect 12584 2492 12585 2556
rect 12519 2476 12585 2492
rect 12519 2412 12520 2476
rect 12584 2412 12585 2476
rect 12519 2396 12585 2412
rect 12519 2332 12520 2396
rect 12584 2332 12585 2396
rect 12519 2316 12585 2332
rect 12519 2252 12520 2316
rect 12584 2252 12585 2316
rect 12519 2236 12585 2252
rect 12519 2172 12520 2236
rect 12584 2172 12585 2236
rect 12519 2156 12585 2172
rect 12519 2092 12520 2156
rect 12584 2092 12585 2156
rect 12519 2076 12585 2092
rect 12519 2012 12520 2076
rect 12584 2012 12585 2076
rect 12519 1996 12585 2012
rect 12519 1932 12520 1996
rect 12584 1932 12585 1996
rect 12519 1778 12585 1932
rect 12645 1840 12705 2870
rect 12765 1778 12825 2810
rect 12885 1840 12945 2870
rect 13005 1778 13065 2810
rect 13125 2716 13191 2806
rect 13125 2652 13126 2716
rect 13190 2652 13191 2716
rect 13125 2636 13191 2652
rect 13125 2572 13126 2636
rect 13190 2572 13191 2636
rect 13125 2556 13191 2572
rect 13125 2492 13126 2556
rect 13190 2492 13191 2556
rect 13125 2476 13191 2492
rect 13125 2412 13126 2476
rect 13190 2412 13191 2476
rect 13125 2396 13191 2412
rect 13125 2332 13126 2396
rect 13190 2332 13191 2396
rect 13125 2316 13191 2332
rect 13125 2252 13126 2316
rect 13190 2252 13191 2316
rect 13125 2236 13191 2252
rect 13125 2172 13126 2236
rect 13190 2172 13191 2236
rect 13125 2156 13191 2172
rect 13125 2092 13126 2156
rect 13190 2092 13191 2156
rect 13125 2076 13191 2092
rect 13125 2012 13126 2076
rect 13190 2012 13191 2076
rect 13125 1996 13191 2012
rect 13125 1932 13126 1996
rect 13190 1932 13191 1996
rect 13125 1778 13191 1932
rect 13251 1778 13311 2810
rect 13371 1840 13431 2870
rect 13491 1778 13551 2810
rect 13611 1840 13671 2870
rect 13731 2716 13797 2806
rect 13731 2652 13732 2716
rect 13796 2652 13797 2716
rect 13731 2636 13797 2652
rect 13731 2572 13732 2636
rect 13796 2572 13797 2636
rect 13731 2556 13797 2572
rect 13731 2492 13732 2556
rect 13796 2492 13797 2556
rect 13731 2476 13797 2492
rect 13731 2412 13732 2476
rect 13796 2412 13797 2476
rect 13731 2396 13797 2412
rect 13731 2332 13732 2396
rect 13796 2332 13797 2396
rect 13731 2316 13797 2332
rect 13731 2252 13732 2316
rect 13796 2252 13797 2316
rect 13731 2236 13797 2252
rect 13731 2172 13732 2236
rect 13796 2172 13797 2236
rect 13731 2156 13797 2172
rect 13731 2092 13732 2156
rect 13796 2092 13797 2156
rect 13731 2076 13797 2092
rect 13731 2012 13732 2076
rect 13796 2012 13797 2076
rect 13731 1996 13797 2012
rect 13731 1932 13732 1996
rect 13796 1932 13797 1996
rect 13731 1778 13797 1932
rect 13857 1840 13917 2870
rect 13977 1778 14037 2810
rect 14097 1840 14157 2870
rect 14217 1778 14277 2810
rect 14337 2716 14403 2806
rect 14337 2652 14338 2716
rect 14402 2652 14403 2716
rect 14337 2636 14403 2652
rect 14337 2572 14338 2636
rect 14402 2572 14403 2636
rect 14337 2556 14403 2572
rect 14337 2492 14338 2556
rect 14402 2492 14403 2556
rect 14337 2476 14403 2492
rect 14337 2412 14338 2476
rect 14402 2412 14403 2476
rect 14337 2396 14403 2412
rect 14337 2332 14338 2396
rect 14402 2332 14403 2396
rect 14337 2316 14403 2332
rect 14337 2252 14338 2316
rect 14402 2252 14403 2316
rect 14337 2236 14403 2252
rect 14337 2172 14338 2236
rect 14402 2172 14403 2236
rect 14337 2156 14403 2172
rect 14337 2092 14338 2156
rect 14402 2092 14403 2156
rect 14337 2076 14403 2092
rect 14337 2012 14338 2076
rect 14402 2012 14403 2076
rect 14337 1996 14403 2012
rect 14337 1932 14338 1996
rect 14402 1932 14403 1996
rect 14337 1778 14403 1932
rect 14463 1778 14523 2810
rect 14583 1840 14643 2870
rect 14703 1778 14763 2810
rect 14823 1840 14883 2870
rect 14943 2716 15009 2806
rect 14943 2652 14944 2716
rect 15008 2652 15009 2716
rect 14943 2636 15009 2652
rect 14943 2572 14944 2636
rect 15008 2572 15009 2636
rect 14943 2556 15009 2572
rect 14943 2492 14944 2556
rect 15008 2492 15009 2556
rect 14943 2476 15009 2492
rect 14943 2412 14944 2476
rect 15008 2412 15009 2476
rect 14943 2396 15009 2412
rect 14943 2332 14944 2396
rect 15008 2332 15009 2396
rect 14943 2316 15009 2332
rect 14943 2252 14944 2316
rect 15008 2252 15009 2316
rect 14943 2236 15009 2252
rect 14943 2172 14944 2236
rect 15008 2172 15009 2236
rect 14943 2156 15009 2172
rect 14943 2092 14944 2156
rect 15008 2092 15009 2156
rect 14943 2076 15009 2092
rect 14943 2012 14944 2076
rect 15008 2012 15009 2076
rect 14943 1996 15009 2012
rect 14943 1932 14944 1996
rect 15008 1932 15009 1996
rect 14943 1778 15009 1932
rect 15069 1840 15129 2870
rect 15189 1778 15249 2810
rect 15309 1840 15369 2870
rect 15429 1778 15489 2810
rect 15549 2716 15615 2806
rect 15549 2652 15550 2716
rect 15614 2652 15615 2716
rect 15549 2636 15615 2652
rect 15549 2572 15550 2636
rect 15614 2572 15615 2636
rect 15549 2556 15615 2572
rect 15549 2492 15550 2556
rect 15614 2492 15615 2556
rect 15549 2476 15615 2492
rect 15549 2412 15550 2476
rect 15614 2412 15615 2476
rect 15549 2396 15615 2412
rect 15549 2332 15550 2396
rect 15614 2332 15615 2396
rect 15549 2316 15615 2332
rect 15549 2252 15550 2316
rect 15614 2252 15615 2316
rect 15549 2236 15615 2252
rect 15549 2172 15550 2236
rect 15614 2172 15615 2236
rect 15549 2156 15615 2172
rect 15549 2092 15550 2156
rect 15614 2092 15615 2156
rect 15549 2076 15615 2092
rect 15549 2012 15550 2076
rect 15614 2012 15615 2076
rect 15549 1996 15615 2012
rect 15549 1932 15550 1996
rect 15614 1932 15615 1996
rect 15677 2016 15803 2026
rect 15677 1952 15708 2016
rect 15772 1952 15803 2016
rect 15677 1942 15803 1952
rect 15549 1778 15615 1932
rect 10701 1776 15615 1778
rect 10701 1712 10805 1776
rect 10869 1712 10885 1776
rect 10949 1712 10965 1776
rect 11029 1712 11045 1776
rect 11109 1712 11125 1776
rect 11189 1753 11205 1776
rect 11189 1712 11194 1753
rect 11269 1712 11411 1776
rect 11475 1753 11491 1776
rect 11486 1712 11491 1753
rect 11555 1712 11571 1776
rect 11635 1712 11651 1776
rect 11715 1712 11731 1776
rect 11795 1712 11811 1776
rect 11875 1712 12017 1776
rect 12081 1712 12097 1776
rect 12161 1712 12177 1776
rect 12241 1712 12257 1776
rect 12321 1712 12337 1776
rect 12401 1753 12417 1776
rect 12401 1712 12406 1753
rect 12481 1712 12623 1776
rect 12687 1753 12703 1776
rect 12698 1712 12703 1753
rect 12767 1712 12783 1776
rect 12847 1712 12863 1776
rect 12927 1712 12943 1776
rect 13007 1712 13023 1776
rect 13087 1712 13229 1776
rect 13293 1712 13309 1776
rect 13373 1712 13389 1776
rect 13453 1712 13469 1776
rect 13533 1712 13549 1776
rect 13613 1753 13629 1776
rect 13613 1712 13618 1753
rect 13693 1712 13835 1776
rect 13899 1753 13915 1776
rect 13910 1712 13915 1753
rect 13979 1712 13995 1776
rect 14059 1712 14075 1776
rect 14139 1712 14155 1776
rect 14219 1712 14235 1776
rect 14299 1712 14441 1776
rect 14505 1712 14521 1776
rect 14585 1712 14601 1776
rect 14665 1712 14681 1776
rect 14745 1712 14761 1776
rect 14825 1753 14841 1776
rect 14825 1712 14830 1753
rect 14905 1712 15047 1776
rect 15111 1753 15127 1776
rect 15122 1712 15127 1753
rect 15191 1712 15207 1776
rect 15271 1712 15287 1776
rect 15351 1712 15367 1776
rect 15431 1712 15447 1776
rect 15511 1712 15615 1776
rect 10701 1710 11194 1712
rect 10526 1689 10535 1710
rect 10452 1684 10535 1689
rect 11184 1689 11194 1710
rect 11258 1710 11422 1712
rect 11258 1689 11267 1710
rect 11184 1684 11267 1689
rect 11413 1689 11422 1710
rect 11486 1710 12406 1712
rect 11486 1689 11496 1710
rect 11413 1684 11496 1689
rect 12396 1689 12406 1710
rect 12470 1710 12634 1712
rect 12470 1689 12479 1710
rect 12396 1684 12479 1689
rect 12625 1689 12634 1710
rect 12698 1710 13618 1712
rect 12698 1689 12708 1710
rect 12625 1684 12708 1689
rect 13608 1689 13618 1710
rect 13682 1710 13846 1712
rect 13682 1689 13691 1710
rect 13608 1684 13691 1689
rect 13837 1689 13846 1710
rect 13910 1710 14830 1712
rect 13910 1689 13920 1710
rect 13837 1684 13920 1689
rect 14820 1689 14830 1710
rect 14894 1710 15058 1712
rect 14894 1689 14903 1710
rect 14820 1684 14903 1689
rect 15049 1689 15058 1710
rect 15122 1710 15615 1712
rect 15765 1755 15891 1765
rect 15122 1689 15132 1710
rect 15049 1684 15132 1689
rect 15765 1691 15796 1755
rect 15860 1691 15891 1755
rect 15765 1681 15891 1691
rect 10811 1551 10893 1557
rect 10811 1529 10820 1551
rect 10323 1527 10820 1529
rect 10884 1529 10893 1551
rect 11543 1551 11625 1557
rect 11543 1529 11552 1551
rect 10884 1527 10995 1529
rect 10323 1463 10427 1527
rect 10491 1463 10507 1527
rect 10571 1463 10587 1527
rect 10651 1463 10667 1527
rect 10731 1463 10747 1527
rect 10811 1487 10820 1527
rect 10811 1463 10827 1487
rect 10891 1463 10995 1527
rect 10323 1461 10995 1463
rect 10323 1307 10389 1461
rect 10323 1243 10324 1307
rect 10388 1243 10389 1307
rect 10323 1227 10389 1243
rect 10323 1163 10324 1227
rect 10388 1163 10389 1227
rect 10323 1147 10389 1163
rect 10323 1083 10324 1147
rect 10388 1083 10389 1147
rect 10323 1067 10389 1083
rect 10323 1003 10324 1067
rect 10388 1003 10389 1067
rect 10323 987 10389 1003
rect 10323 923 10324 987
rect 10388 923 10389 987
rect 10323 907 10389 923
rect 10323 843 10324 907
rect 10388 843 10389 907
rect 10323 827 10389 843
rect 10323 763 10324 827
rect 10388 763 10389 827
rect 10323 747 10389 763
rect 10323 683 10324 747
rect 10388 683 10389 747
rect 10323 667 10389 683
rect 10323 603 10324 667
rect 10388 603 10389 667
rect 10323 587 10389 603
rect 10323 523 10324 587
rect 10388 523 10389 587
rect 10323 433 10389 523
rect 10449 429 10509 1461
rect 9932 365 10057 375
rect 10569 369 10629 1399
rect 10689 429 10749 1461
rect 10809 369 10869 1399
rect 10929 1307 10995 1461
rect 10929 1243 10930 1307
rect 10994 1243 10995 1307
rect 10929 1227 10995 1243
rect 10929 1163 10930 1227
rect 10994 1163 10995 1227
rect 10929 1147 10995 1163
rect 10929 1083 10930 1147
rect 10994 1083 10995 1147
rect 10929 1067 10995 1083
rect 10929 1003 10930 1067
rect 10994 1003 10995 1067
rect 10929 987 10995 1003
rect 10929 923 10930 987
rect 10994 923 10995 987
rect 10929 907 10995 923
rect 10929 843 10930 907
rect 10994 843 10995 907
rect 10929 827 10995 843
rect 10929 763 10930 827
rect 10994 763 10995 827
rect 10929 747 10995 763
rect 10929 683 10930 747
rect 10994 683 10995 747
rect 10929 667 10995 683
rect 10929 603 10930 667
rect 10994 603 10995 667
rect 10929 587 10995 603
rect 10929 523 10930 587
rect 10994 523 10995 587
rect 10929 433 10995 523
rect 11055 1527 11552 1529
rect 11616 1529 11625 1551
rect 11763 1551 11845 1557
rect 11763 1529 11772 1551
rect 11616 1527 11772 1529
rect 11836 1529 11845 1551
rect 12755 1551 12837 1557
rect 12755 1529 12764 1551
rect 11836 1527 12764 1529
rect 12828 1529 12837 1551
rect 12975 1551 13057 1557
rect 12975 1529 12984 1551
rect 12828 1527 12984 1529
rect 13048 1529 13057 1551
rect 14093 1551 14175 1557
rect 14093 1529 14102 1551
rect 13048 1527 13545 1529
rect 11055 1463 11159 1527
rect 11223 1463 11239 1527
rect 11303 1463 11319 1527
rect 11383 1463 11399 1527
rect 11463 1463 11479 1527
rect 11543 1487 11552 1527
rect 11543 1463 11559 1487
rect 11623 1463 11765 1527
rect 11836 1487 11845 1527
rect 11829 1463 11845 1487
rect 11909 1463 11925 1527
rect 11989 1463 12005 1527
rect 12069 1463 12085 1527
rect 12149 1463 12165 1527
rect 12229 1463 12371 1527
rect 12435 1463 12451 1527
rect 12515 1463 12531 1527
rect 12595 1463 12611 1527
rect 12675 1463 12691 1527
rect 12755 1487 12764 1527
rect 12755 1463 12771 1487
rect 12835 1463 12977 1527
rect 13048 1487 13057 1527
rect 13041 1463 13057 1487
rect 13121 1463 13137 1527
rect 13201 1463 13217 1527
rect 13281 1463 13297 1527
rect 13361 1463 13377 1527
rect 13441 1463 13545 1527
rect 11055 1461 13545 1463
rect 11055 1307 11121 1461
rect 11055 1243 11056 1307
rect 11120 1243 11121 1307
rect 11055 1227 11121 1243
rect 11055 1163 11056 1227
rect 11120 1163 11121 1227
rect 11055 1147 11121 1163
rect 11055 1083 11056 1147
rect 11120 1083 11121 1147
rect 11055 1067 11121 1083
rect 11055 1003 11056 1067
rect 11120 1003 11121 1067
rect 11055 987 11121 1003
rect 11055 923 11056 987
rect 11120 923 11121 987
rect 11055 907 11121 923
rect 11055 843 11056 907
rect 11120 843 11121 907
rect 11055 827 11121 843
rect 11055 763 11056 827
rect 11120 763 11121 827
rect 11055 747 11121 763
rect 11055 683 11056 747
rect 11120 683 11121 747
rect 11055 667 11121 683
rect 11055 603 11056 667
rect 11120 603 11121 667
rect 11055 587 11121 603
rect 11055 523 11056 587
rect 11120 523 11121 587
rect 11055 433 11121 523
rect 11181 429 11241 1461
rect 11301 369 11361 1399
rect 11421 429 11481 1461
rect 11541 369 11601 1399
rect 11661 1307 11727 1461
rect 11661 1243 11662 1307
rect 11726 1243 11727 1307
rect 11661 1227 11727 1243
rect 11661 1163 11662 1227
rect 11726 1163 11727 1227
rect 11661 1147 11727 1163
rect 11661 1083 11662 1147
rect 11726 1083 11727 1147
rect 11661 1067 11727 1083
rect 11661 1003 11662 1067
rect 11726 1003 11727 1067
rect 11661 987 11727 1003
rect 11661 923 11662 987
rect 11726 923 11727 987
rect 11661 907 11727 923
rect 11661 843 11662 907
rect 11726 843 11727 907
rect 11661 827 11727 843
rect 11661 763 11662 827
rect 11726 763 11727 827
rect 11661 747 11727 763
rect 11661 683 11662 747
rect 11726 683 11727 747
rect 11661 667 11727 683
rect 11661 603 11662 667
rect 11726 603 11727 667
rect 11661 587 11727 603
rect 11661 523 11662 587
rect 11726 523 11727 587
rect 11661 433 11727 523
rect 11787 369 11847 1399
rect 11907 429 11967 1461
rect 12027 369 12087 1399
rect 12147 429 12207 1461
rect 12267 1307 12333 1461
rect 12267 1243 12268 1307
rect 12332 1243 12333 1307
rect 12267 1227 12333 1243
rect 12267 1163 12268 1227
rect 12332 1163 12333 1227
rect 12267 1147 12333 1163
rect 12267 1083 12268 1147
rect 12332 1083 12333 1147
rect 12267 1067 12333 1083
rect 12267 1003 12268 1067
rect 12332 1003 12333 1067
rect 12267 987 12333 1003
rect 12267 923 12268 987
rect 12332 923 12333 987
rect 12267 907 12333 923
rect 12267 843 12268 907
rect 12332 843 12333 907
rect 12267 827 12333 843
rect 12267 763 12268 827
rect 12332 763 12333 827
rect 12267 747 12333 763
rect 12267 683 12268 747
rect 12332 683 12333 747
rect 12267 667 12333 683
rect 12267 603 12268 667
rect 12332 603 12333 667
rect 12267 587 12333 603
rect 12267 523 12268 587
rect 12332 523 12333 587
rect 12267 433 12333 523
rect 12393 429 12453 1461
rect 12513 369 12573 1399
rect 12633 429 12693 1461
rect 12753 369 12813 1399
rect 12873 1307 12939 1461
rect 12873 1243 12874 1307
rect 12938 1243 12939 1307
rect 12873 1227 12939 1243
rect 12873 1163 12874 1227
rect 12938 1163 12939 1227
rect 12873 1147 12939 1163
rect 12873 1083 12874 1147
rect 12938 1083 12939 1147
rect 12873 1067 12939 1083
rect 12873 1003 12874 1067
rect 12938 1003 12939 1067
rect 12873 987 12939 1003
rect 12873 923 12874 987
rect 12938 923 12939 987
rect 12873 907 12939 923
rect 12873 843 12874 907
rect 12938 843 12939 907
rect 12873 827 12939 843
rect 12873 763 12874 827
rect 12938 763 12939 827
rect 12873 747 12939 763
rect 12873 683 12874 747
rect 12938 683 12939 747
rect 12873 667 12939 683
rect 12873 603 12874 667
rect 12938 603 12939 667
rect 12873 587 12939 603
rect 12873 523 12874 587
rect 12938 523 12939 587
rect 12873 433 12939 523
rect 12999 369 13059 1399
rect 13119 429 13179 1461
rect 13239 369 13299 1399
rect 13359 429 13419 1461
rect 13479 1307 13545 1461
rect 13479 1243 13480 1307
rect 13544 1243 13545 1307
rect 13479 1227 13545 1243
rect 13479 1163 13480 1227
rect 13544 1163 13545 1227
rect 13479 1147 13545 1163
rect 13479 1083 13480 1147
rect 13544 1083 13545 1147
rect 13479 1067 13545 1083
rect 13479 1003 13480 1067
rect 13544 1003 13545 1067
rect 13479 987 13545 1003
rect 13479 923 13480 987
rect 13544 923 13545 987
rect 13479 907 13545 923
rect 13479 843 13480 907
rect 13544 843 13545 907
rect 13479 827 13545 843
rect 13479 763 13480 827
rect 13544 763 13545 827
rect 13479 747 13545 763
rect 13479 683 13480 747
rect 13544 683 13545 747
rect 13479 667 13545 683
rect 13479 603 13480 667
rect 13544 603 13545 667
rect 13479 587 13545 603
rect 13479 523 13480 587
rect 13544 523 13545 587
rect 13479 433 13545 523
rect 13605 1527 14102 1529
rect 14166 1529 14175 1551
rect 14313 1551 14395 1557
rect 14313 1529 14322 1551
rect 14166 1527 14322 1529
rect 14386 1529 14395 1551
rect 15045 1551 15127 1557
rect 15045 1529 15054 1551
rect 14386 1527 14883 1529
rect 13605 1463 13709 1527
rect 13773 1463 13789 1527
rect 13853 1463 13869 1527
rect 13933 1463 13949 1527
rect 14013 1463 14029 1527
rect 14093 1487 14102 1527
rect 14093 1463 14109 1487
rect 14173 1463 14315 1527
rect 14386 1487 14395 1527
rect 14379 1463 14395 1487
rect 14459 1463 14475 1527
rect 14539 1463 14555 1527
rect 14619 1463 14635 1527
rect 14699 1463 14715 1527
rect 14779 1463 14883 1527
rect 13605 1461 14883 1463
rect 13605 1307 13671 1461
rect 13605 1243 13606 1307
rect 13670 1243 13671 1307
rect 13605 1227 13671 1243
rect 13605 1163 13606 1227
rect 13670 1163 13671 1227
rect 13605 1147 13671 1163
rect 13605 1083 13606 1147
rect 13670 1083 13671 1147
rect 13605 1067 13671 1083
rect 13605 1003 13606 1067
rect 13670 1003 13671 1067
rect 13605 987 13671 1003
rect 13605 923 13606 987
rect 13670 923 13671 987
rect 13605 907 13671 923
rect 13605 843 13606 907
rect 13670 843 13671 907
rect 13605 827 13671 843
rect 13605 763 13606 827
rect 13670 763 13671 827
rect 13605 747 13671 763
rect 13605 683 13606 747
rect 13670 683 13671 747
rect 13605 667 13671 683
rect 13605 603 13606 667
rect 13670 603 13671 667
rect 13605 587 13671 603
rect 13605 523 13606 587
rect 13670 523 13671 587
rect 13605 433 13671 523
rect 13731 429 13791 1461
rect 13851 369 13911 1399
rect 13971 429 14031 1461
rect 14091 369 14151 1399
rect 14211 1307 14277 1461
rect 14211 1243 14212 1307
rect 14276 1243 14277 1307
rect 14211 1227 14277 1243
rect 14211 1163 14212 1227
rect 14276 1163 14277 1227
rect 14211 1147 14277 1163
rect 14211 1083 14212 1147
rect 14276 1083 14277 1147
rect 14211 1067 14277 1083
rect 14211 1003 14212 1067
rect 14276 1003 14277 1067
rect 14211 987 14277 1003
rect 14211 923 14212 987
rect 14276 923 14277 987
rect 14211 907 14277 923
rect 14211 843 14212 907
rect 14276 843 14277 907
rect 14211 827 14277 843
rect 14211 763 14212 827
rect 14276 763 14277 827
rect 14211 747 14277 763
rect 14211 683 14212 747
rect 14276 683 14277 747
rect 14211 667 14277 683
rect 14211 603 14212 667
rect 14276 603 14277 667
rect 14211 587 14277 603
rect 14211 523 14212 587
rect 14276 523 14277 587
rect 14211 433 14277 523
rect 14337 369 14397 1399
rect 14457 429 14517 1461
rect 14577 369 14637 1399
rect 14697 429 14757 1461
rect 14817 1307 14883 1461
rect 14817 1243 14818 1307
rect 14882 1243 14883 1307
rect 14817 1227 14883 1243
rect 14817 1163 14818 1227
rect 14882 1163 14883 1227
rect 14817 1147 14883 1163
rect 14817 1083 14818 1147
rect 14882 1083 14883 1147
rect 14817 1067 14883 1083
rect 14817 1003 14818 1067
rect 14882 1003 14883 1067
rect 14817 987 14883 1003
rect 14817 923 14818 987
rect 14882 923 14883 987
rect 14817 907 14883 923
rect 14817 843 14818 907
rect 14882 843 14883 907
rect 14817 827 14883 843
rect 14817 763 14818 827
rect 14882 763 14883 827
rect 14817 747 14883 763
rect 14817 683 14818 747
rect 14882 683 14883 747
rect 14817 667 14883 683
rect 14817 603 14818 667
rect 14882 603 14883 667
rect 14817 587 14883 603
rect 14817 523 14818 587
rect 14882 523 14883 587
rect 14817 433 14883 523
rect 14943 1527 15054 1529
rect 15118 1529 15127 1551
rect 15765 1552 15891 1562
rect 15118 1527 15615 1529
rect 14943 1463 15047 1527
rect 15118 1487 15127 1527
rect 15111 1463 15127 1487
rect 15191 1463 15207 1527
rect 15271 1463 15287 1527
rect 15351 1463 15367 1527
rect 15431 1463 15447 1527
rect 15511 1463 15615 1527
rect 15765 1488 15796 1552
rect 15860 1488 15891 1552
rect 15765 1478 15891 1488
rect 15791 1477 15865 1478
rect 14943 1461 15615 1463
rect 14943 1307 15009 1461
rect 14943 1243 14944 1307
rect 15008 1243 15009 1307
rect 14943 1227 15009 1243
rect 14943 1163 14944 1227
rect 15008 1163 15009 1227
rect 14943 1147 15009 1163
rect 14943 1083 14944 1147
rect 15008 1083 15009 1147
rect 14943 1067 15009 1083
rect 14943 1003 14944 1067
rect 15008 1003 15009 1067
rect 14943 987 15009 1003
rect 14943 923 14944 987
rect 15008 923 15009 987
rect 14943 907 15009 923
rect 14943 843 14944 907
rect 15008 843 15009 907
rect 14943 827 15009 843
rect 14943 763 14944 827
rect 15008 763 15009 827
rect 14943 747 15009 763
rect 14943 683 14944 747
rect 15008 683 15009 747
rect 14943 667 15009 683
rect 14943 603 14944 667
rect 15008 603 15009 667
rect 14943 587 15009 603
rect 14943 523 14944 587
rect 15008 523 15009 587
rect 14943 433 15009 523
rect 15069 369 15129 1399
rect 15189 429 15249 1461
rect 15309 369 15369 1399
rect 15429 429 15489 1461
rect 15549 1307 15615 1461
rect 15549 1243 15550 1307
rect 15614 1243 15615 1307
rect 15549 1227 15615 1243
rect 15549 1163 15550 1227
rect 15614 1163 15615 1227
rect 15675 1290 15800 1300
rect 15675 1226 15705 1290
rect 15769 1226 15800 1290
rect 15675 1216 15800 1226
rect 15549 1147 15615 1163
rect 15549 1083 15550 1147
rect 15614 1083 15615 1147
rect 15549 1067 15615 1083
rect 15549 1003 15550 1067
rect 15614 1003 15615 1067
rect 15549 987 15615 1003
rect 15549 923 15550 987
rect 15614 923 15615 987
rect 15549 907 15615 923
rect 15549 843 15550 907
rect 15614 843 15615 907
rect 15549 827 15615 843
rect 15549 763 15550 827
rect 15614 763 15615 827
rect 15549 747 15615 763
rect 15549 683 15550 747
rect 15614 683 15615 747
rect 15549 667 15615 683
rect 15549 603 15550 667
rect 15614 603 15615 667
rect 15549 587 15615 603
rect 15549 523 15550 587
rect 15614 523 15615 587
rect 15549 433 15615 523
rect 9932 301 9962 365
rect 10026 301 10057 365
rect 10323 367 10995 369
rect 10323 303 10427 367
rect 10491 303 10507 367
rect 10571 303 10587 367
rect 10651 303 10667 367
rect 10731 303 10747 367
rect 10811 303 10827 367
rect 10891 303 10995 367
rect 10323 301 10995 303
rect 11055 367 13545 369
rect 11055 303 11159 367
rect 11223 303 11239 367
rect 11303 303 11319 367
rect 11383 303 11399 367
rect 11463 303 11479 367
rect 11543 303 11559 367
rect 11623 303 11765 367
rect 11829 303 11845 367
rect 11909 303 11925 367
rect 11989 303 12005 367
rect 12069 303 12085 367
rect 12149 303 12165 367
rect 12229 303 12371 367
rect 12435 303 12451 367
rect 12515 303 12531 367
rect 12595 303 12611 367
rect 12675 303 12691 367
rect 12755 303 12771 367
rect 12835 303 12977 367
rect 13041 303 13057 367
rect 13121 303 13137 367
rect 13201 303 13217 367
rect 13281 303 13297 367
rect 13361 303 13377 367
rect 13441 303 13545 367
rect 11055 301 13545 303
rect 13605 367 14883 369
rect 13605 303 13709 367
rect 13773 303 13789 367
rect 13853 303 13869 367
rect 13933 303 13949 367
rect 14013 303 14029 367
rect 14093 303 14109 367
rect 14173 303 14315 367
rect 14379 303 14395 367
rect 14459 303 14475 367
rect 14539 303 14555 367
rect 14619 303 14635 367
rect 14699 303 14715 367
rect 14779 303 14883 367
rect 13605 301 14883 303
rect 14943 367 15615 369
rect 14943 303 15047 367
rect 15111 303 15127 367
rect 15191 303 15207 367
rect 15271 303 15287 367
rect 15351 303 15367 367
rect 15431 303 15447 367
rect 15511 303 15615 367
rect 14943 301 15615 303
rect 9932 291 10057 301
<< via3 >>
rect 9976 2939 10040 2943
rect 9976 2883 9980 2939
rect 9980 2883 10036 2939
rect 10036 2883 10040 2939
rect 9976 2879 10040 2883
rect 10073 2872 10137 2936
rect 10153 2872 10217 2936
rect 10233 2872 10297 2936
rect 10313 2872 10377 2936
rect 10393 2872 10457 2936
rect 10473 2872 10537 2936
rect 10805 2872 10869 2936
rect 10885 2872 10949 2936
rect 10965 2872 11029 2936
rect 11045 2872 11109 2936
rect 11125 2872 11189 2936
rect 11205 2872 11269 2936
rect 11411 2872 11475 2936
rect 11491 2872 11555 2936
rect 11571 2872 11635 2936
rect 11651 2872 11715 2936
rect 11731 2872 11795 2936
rect 11811 2872 11875 2936
rect 12017 2872 12081 2936
rect 12097 2872 12161 2936
rect 12177 2872 12241 2936
rect 12257 2872 12321 2936
rect 12337 2872 12401 2936
rect 12417 2872 12481 2936
rect 12623 2872 12687 2936
rect 12703 2872 12767 2936
rect 12783 2872 12847 2936
rect 12863 2872 12927 2936
rect 12943 2872 13007 2936
rect 13023 2872 13087 2936
rect 13229 2872 13293 2936
rect 13309 2872 13373 2936
rect 13389 2872 13453 2936
rect 13469 2872 13533 2936
rect 13549 2872 13613 2936
rect 13629 2872 13693 2936
rect 13835 2872 13899 2936
rect 13915 2872 13979 2936
rect 13995 2872 14059 2936
rect 14075 2872 14139 2936
rect 14155 2872 14219 2936
rect 14235 2872 14299 2936
rect 14441 2872 14505 2936
rect 14521 2872 14585 2936
rect 14601 2872 14665 2936
rect 14681 2872 14745 2936
rect 14761 2872 14825 2936
rect 14841 2872 14905 2936
rect 15047 2872 15111 2936
rect 15127 2872 15191 2936
rect 15207 2872 15271 2936
rect 15287 2872 15351 2936
rect 15367 2872 15431 2936
rect 15447 2872 15511 2936
rect 9970 2652 10034 2716
rect 9970 2572 10034 2636
rect 9970 2492 10034 2556
rect 9970 2412 10034 2476
rect 9359 2334 9423 2338
rect 9359 2278 9363 2334
rect 9363 2278 9419 2334
rect 9419 2278 9423 2334
rect 9359 2274 9423 2278
rect 9490 2333 9554 2337
rect 9490 2277 9494 2333
rect 9494 2277 9550 2333
rect 9550 2277 9554 2333
rect 9490 2273 9554 2277
rect 9634 2334 9698 2338
rect 9634 2278 9638 2334
rect 9638 2278 9694 2334
rect 9694 2278 9698 2334
rect 9634 2274 9698 2278
rect 9970 2332 10034 2396
rect 9970 2252 10034 2316
rect 9970 2172 10034 2236
rect 9970 2092 10034 2156
rect 9970 2012 10034 2076
rect 9970 1932 10034 1996
rect 9377 1788 9441 1792
rect 9377 1732 9381 1788
rect 9381 1732 9437 1788
rect 9437 1732 9441 1788
rect 9377 1728 9441 1732
rect 9497 1788 9561 1792
rect 9497 1732 9501 1788
rect 9501 1732 9557 1788
rect 9557 1732 9561 1788
rect 9497 1728 9561 1732
rect 9640 1788 9704 1792
rect 9640 1732 9644 1788
rect 9644 1732 9700 1788
rect 9700 1732 9704 1788
rect 9640 1728 9704 1732
rect 10576 2652 10640 2716
rect 10576 2572 10640 2636
rect 10576 2492 10640 2556
rect 10576 2412 10640 2476
rect 10576 2332 10640 2396
rect 10576 2252 10640 2316
rect 10576 2172 10640 2236
rect 10576 2092 10640 2156
rect 10576 2012 10640 2076
rect 10576 1932 10640 1996
rect 10073 1712 10137 1776
rect 10153 1712 10217 1776
rect 10233 1712 10297 1776
rect 10313 1712 10377 1776
rect 10393 1712 10457 1776
rect 10473 1753 10537 1776
rect 10473 1712 10526 1753
rect 10526 1712 10537 1753
rect 10702 2652 10766 2716
rect 10702 2572 10766 2636
rect 10702 2492 10766 2556
rect 10702 2412 10766 2476
rect 10702 2332 10766 2396
rect 10702 2252 10766 2316
rect 10702 2172 10766 2236
rect 10702 2092 10766 2156
rect 10702 2012 10766 2076
rect 10702 1932 10766 1996
rect 11308 2652 11372 2716
rect 11308 2572 11372 2636
rect 11308 2492 11372 2556
rect 11308 2412 11372 2476
rect 11308 2332 11372 2396
rect 11308 2252 11372 2316
rect 11308 2172 11372 2236
rect 11308 2092 11372 2156
rect 11308 2012 11372 2076
rect 11308 1932 11372 1996
rect 11914 2652 11978 2716
rect 11914 2572 11978 2636
rect 11914 2492 11978 2556
rect 11914 2412 11978 2476
rect 11914 2332 11978 2396
rect 11914 2252 11978 2316
rect 11914 2172 11978 2236
rect 11914 2092 11978 2156
rect 11914 2012 11978 2076
rect 11914 1932 11978 1996
rect 12520 2652 12584 2716
rect 12520 2572 12584 2636
rect 12520 2492 12584 2556
rect 12520 2412 12584 2476
rect 12520 2332 12584 2396
rect 12520 2252 12584 2316
rect 12520 2172 12584 2236
rect 12520 2092 12584 2156
rect 12520 2012 12584 2076
rect 12520 1932 12584 1996
rect 13126 2652 13190 2716
rect 13126 2572 13190 2636
rect 13126 2492 13190 2556
rect 13126 2412 13190 2476
rect 13126 2332 13190 2396
rect 13126 2252 13190 2316
rect 13126 2172 13190 2236
rect 13126 2092 13190 2156
rect 13126 2012 13190 2076
rect 13126 1932 13190 1996
rect 13732 2652 13796 2716
rect 13732 2572 13796 2636
rect 13732 2492 13796 2556
rect 13732 2412 13796 2476
rect 13732 2332 13796 2396
rect 13732 2252 13796 2316
rect 13732 2172 13796 2236
rect 13732 2092 13796 2156
rect 13732 2012 13796 2076
rect 13732 1932 13796 1996
rect 14338 2652 14402 2716
rect 14338 2572 14402 2636
rect 14338 2492 14402 2556
rect 14338 2412 14402 2476
rect 14338 2332 14402 2396
rect 14338 2252 14402 2316
rect 14338 2172 14402 2236
rect 14338 2092 14402 2156
rect 14338 2012 14402 2076
rect 14338 1932 14402 1996
rect 14944 2652 15008 2716
rect 14944 2572 15008 2636
rect 14944 2492 15008 2556
rect 14944 2412 15008 2476
rect 14944 2332 15008 2396
rect 14944 2252 15008 2316
rect 14944 2172 15008 2236
rect 14944 2092 15008 2156
rect 14944 2012 15008 2076
rect 14944 1932 15008 1996
rect 15550 2652 15614 2716
rect 15550 2572 15614 2636
rect 15550 2492 15614 2556
rect 15550 2412 15614 2476
rect 15550 2332 15614 2396
rect 15550 2252 15614 2316
rect 15550 2172 15614 2236
rect 15550 2092 15614 2156
rect 15550 2012 15614 2076
rect 15550 1932 15614 1996
rect 15708 2012 15772 2016
rect 15708 1956 15712 2012
rect 15712 1956 15768 2012
rect 15768 1956 15772 2012
rect 15708 1952 15772 1956
rect 10805 1712 10869 1776
rect 10885 1712 10949 1776
rect 10965 1712 11029 1776
rect 11045 1712 11109 1776
rect 11125 1712 11189 1776
rect 11205 1753 11269 1776
rect 11205 1712 11258 1753
rect 11258 1712 11269 1753
rect 11411 1753 11475 1776
rect 11411 1712 11422 1753
rect 11422 1712 11475 1753
rect 11491 1712 11555 1776
rect 11571 1712 11635 1776
rect 11651 1712 11715 1776
rect 11731 1712 11795 1776
rect 11811 1712 11875 1776
rect 12017 1712 12081 1776
rect 12097 1712 12161 1776
rect 12177 1712 12241 1776
rect 12257 1712 12321 1776
rect 12337 1712 12401 1776
rect 12417 1753 12481 1776
rect 12417 1712 12470 1753
rect 12470 1712 12481 1753
rect 12623 1753 12687 1776
rect 12623 1712 12634 1753
rect 12634 1712 12687 1753
rect 12703 1712 12767 1776
rect 12783 1712 12847 1776
rect 12863 1712 12927 1776
rect 12943 1712 13007 1776
rect 13023 1712 13087 1776
rect 13229 1712 13293 1776
rect 13309 1712 13373 1776
rect 13389 1712 13453 1776
rect 13469 1712 13533 1776
rect 13549 1712 13613 1776
rect 13629 1753 13693 1776
rect 13629 1712 13682 1753
rect 13682 1712 13693 1753
rect 13835 1753 13899 1776
rect 13835 1712 13846 1753
rect 13846 1712 13899 1753
rect 13915 1712 13979 1776
rect 13995 1712 14059 1776
rect 14075 1712 14139 1776
rect 14155 1712 14219 1776
rect 14235 1712 14299 1776
rect 14441 1712 14505 1776
rect 14521 1712 14585 1776
rect 14601 1712 14665 1776
rect 14681 1712 14745 1776
rect 14761 1712 14825 1776
rect 14841 1753 14905 1776
rect 14841 1712 14894 1753
rect 14894 1712 14905 1753
rect 15047 1753 15111 1776
rect 15047 1712 15058 1753
rect 15058 1712 15111 1753
rect 15127 1712 15191 1776
rect 15207 1712 15271 1776
rect 15287 1712 15351 1776
rect 15367 1712 15431 1776
rect 15447 1712 15511 1776
rect 15796 1751 15860 1755
rect 15796 1695 15800 1751
rect 15800 1695 15856 1751
rect 15856 1695 15860 1751
rect 15796 1691 15860 1695
rect 10427 1463 10491 1527
rect 10507 1463 10571 1527
rect 10587 1463 10651 1527
rect 10667 1463 10731 1527
rect 10747 1463 10811 1527
rect 10827 1487 10884 1527
rect 10884 1487 10891 1527
rect 10827 1463 10891 1487
rect 10324 1243 10388 1307
rect 10324 1163 10388 1227
rect 10324 1083 10388 1147
rect 10324 1003 10388 1067
rect 10324 923 10388 987
rect 10324 843 10388 907
rect 10324 763 10388 827
rect 10324 683 10388 747
rect 10324 603 10388 667
rect 10324 523 10388 587
rect 10930 1243 10994 1307
rect 10930 1163 10994 1227
rect 10930 1083 10994 1147
rect 10930 1003 10994 1067
rect 10930 923 10994 987
rect 10930 843 10994 907
rect 10930 763 10994 827
rect 10930 683 10994 747
rect 10930 603 10994 667
rect 10930 523 10994 587
rect 11159 1463 11223 1527
rect 11239 1463 11303 1527
rect 11319 1463 11383 1527
rect 11399 1463 11463 1527
rect 11479 1463 11543 1527
rect 11559 1487 11616 1527
rect 11616 1487 11623 1527
rect 11559 1463 11623 1487
rect 11765 1487 11772 1527
rect 11772 1487 11829 1527
rect 11765 1463 11829 1487
rect 11845 1463 11909 1527
rect 11925 1463 11989 1527
rect 12005 1463 12069 1527
rect 12085 1463 12149 1527
rect 12165 1463 12229 1527
rect 12371 1463 12435 1527
rect 12451 1463 12515 1527
rect 12531 1463 12595 1527
rect 12611 1463 12675 1527
rect 12691 1463 12755 1527
rect 12771 1487 12828 1527
rect 12828 1487 12835 1527
rect 12771 1463 12835 1487
rect 12977 1487 12984 1527
rect 12984 1487 13041 1527
rect 12977 1463 13041 1487
rect 13057 1463 13121 1527
rect 13137 1463 13201 1527
rect 13217 1463 13281 1527
rect 13297 1463 13361 1527
rect 13377 1463 13441 1527
rect 11056 1243 11120 1307
rect 11056 1163 11120 1227
rect 11056 1083 11120 1147
rect 11056 1003 11120 1067
rect 11056 923 11120 987
rect 11056 843 11120 907
rect 11056 763 11120 827
rect 11056 683 11120 747
rect 11056 603 11120 667
rect 11056 523 11120 587
rect 11662 1243 11726 1307
rect 11662 1163 11726 1227
rect 11662 1083 11726 1147
rect 11662 1003 11726 1067
rect 11662 923 11726 987
rect 11662 843 11726 907
rect 11662 763 11726 827
rect 11662 683 11726 747
rect 11662 603 11726 667
rect 11662 523 11726 587
rect 12268 1243 12332 1307
rect 12268 1163 12332 1227
rect 12268 1083 12332 1147
rect 12268 1003 12332 1067
rect 12268 923 12332 987
rect 12268 843 12332 907
rect 12268 763 12332 827
rect 12268 683 12332 747
rect 12268 603 12332 667
rect 12268 523 12332 587
rect 12874 1243 12938 1307
rect 12874 1163 12938 1227
rect 12874 1083 12938 1147
rect 12874 1003 12938 1067
rect 12874 923 12938 987
rect 12874 843 12938 907
rect 12874 763 12938 827
rect 12874 683 12938 747
rect 12874 603 12938 667
rect 12874 523 12938 587
rect 13480 1243 13544 1307
rect 13480 1163 13544 1227
rect 13480 1083 13544 1147
rect 13480 1003 13544 1067
rect 13480 923 13544 987
rect 13480 843 13544 907
rect 13480 763 13544 827
rect 13480 683 13544 747
rect 13480 603 13544 667
rect 13480 523 13544 587
rect 13709 1463 13773 1527
rect 13789 1463 13853 1527
rect 13869 1463 13933 1527
rect 13949 1463 14013 1527
rect 14029 1463 14093 1527
rect 14109 1487 14166 1527
rect 14166 1487 14173 1527
rect 14109 1463 14173 1487
rect 14315 1487 14322 1527
rect 14322 1487 14379 1527
rect 14315 1463 14379 1487
rect 14395 1463 14459 1527
rect 14475 1463 14539 1527
rect 14555 1463 14619 1527
rect 14635 1463 14699 1527
rect 14715 1463 14779 1527
rect 13606 1243 13670 1307
rect 13606 1163 13670 1227
rect 13606 1083 13670 1147
rect 13606 1003 13670 1067
rect 13606 923 13670 987
rect 13606 843 13670 907
rect 13606 763 13670 827
rect 13606 683 13670 747
rect 13606 603 13670 667
rect 13606 523 13670 587
rect 14212 1243 14276 1307
rect 14212 1163 14276 1227
rect 14212 1083 14276 1147
rect 14212 1003 14276 1067
rect 14212 923 14276 987
rect 14212 843 14276 907
rect 14212 763 14276 827
rect 14212 683 14276 747
rect 14212 603 14276 667
rect 14212 523 14276 587
rect 14818 1243 14882 1307
rect 14818 1163 14882 1227
rect 14818 1083 14882 1147
rect 14818 1003 14882 1067
rect 14818 923 14882 987
rect 14818 843 14882 907
rect 14818 763 14882 827
rect 14818 683 14882 747
rect 14818 603 14882 667
rect 14818 523 14882 587
rect 15047 1487 15054 1527
rect 15054 1487 15111 1527
rect 15047 1463 15111 1487
rect 15127 1463 15191 1527
rect 15207 1463 15271 1527
rect 15287 1463 15351 1527
rect 15367 1463 15431 1527
rect 15447 1463 15511 1527
rect 15796 1548 15860 1552
rect 15796 1492 15800 1548
rect 15800 1492 15856 1548
rect 15856 1492 15860 1548
rect 15796 1488 15860 1492
rect 14944 1243 15008 1307
rect 14944 1163 15008 1227
rect 14944 1083 15008 1147
rect 14944 1003 15008 1067
rect 14944 923 15008 987
rect 14944 843 15008 907
rect 14944 763 15008 827
rect 14944 683 15008 747
rect 14944 603 15008 667
rect 14944 523 15008 587
rect 15550 1243 15614 1307
rect 15550 1163 15614 1227
rect 15705 1286 15769 1290
rect 15705 1230 15709 1286
rect 15709 1230 15765 1286
rect 15765 1230 15769 1286
rect 15705 1226 15769 1230
rect 15550 1083 15614 1147
rect 15550 1003 15614 1067
rect 15550 923 15614 987
rect 15550 843 15614 907
rect 15550 763 15614 827
rect 15550 683 15614 747
rect 15550 603 15614 667
rect 15550 523 15614 587
rect 9962 361 10026 365
rect 9962 305 9966 361
rect 9966 305 10022 361
rect 10022 305 10026 361
rect 9962 301 10026 305
rect 10427 303 10491 367
rect 10507 303 10571 367
rect 10587 303 10651 367
rect 10667 303 10731 367
rect 10747 303 10811 367
rect 10827 303 10891 367
rect 11159 303 11223 367
rect 11239 303 11303 367
rect 11319 303 11383 367
rect 11399 303 11463 367
rect 11479 303 11543 367
rect 11559 303 11623 367
rect 11765 303 11829 367
rect 11845 303 11909 367
rect 11925 303 11989 367
rect 12005 303 12069 367
rect 12085 303 12149 367
rect 12165 303 12229 367
rect 12371 303 12435 367
rect 12451 303 12515 367
rect 12531 303 12595 367
rect 12611 303 12675 367
rect 12691 303 12755 367
rect 12771 303 12835 367
rect 12977 303 13041 367
rect 13057 303 13121 367
rect 13137 303 13201 367
rect 13217 303 13281 367
rect 13297 303 13361 367
rect 13377 303 13441 367
rect 13709 303 13773 367
rect 13789 303 13853 367
rect 13869 303 13933 367
rect 13949 303 14013 367
rect 14029 303 14093 367
rect 14109 303 14173 367
rect 14315 303 14379 367
rect 14395 303 14459 367
rect 14475 303 14539 367
rect 14555 303 14619 367
rect 14635 303 14699 367
rect 14715 303 14779 367
rect 15047 303 15111 367
rect 15127 303 15191 367
rect 15207 303 15271 367
rect 15287 303 15351 367
rect 15367 303 15431 367
rect 15447 303 15511 367
<< metal4 >>
rect 9945 2948 10071 2953
rect 9299 2943 15993 2948
rect 9299 2879 9976 2943
rect 10040 2936 15993 2943
rect 10040 2879 10073 2936
rect 9299 2872 10073 2879
rect 10137 2872 10153 2936
rect 10217 2872 10233 2936
rect 10297 2872 10313 2936
rect 10377 2872 10393 2936
rect 10457 2872 10473 2936
rect 10537 2872 10805 2936
rect 10869 2872 10885 2936
rect 10949 2872 10965 2936
rect 11029 2872 11045 2936
rect 11109 2872 11125 2936
rect 11189 2872 11205 2936
rect 11269 2872 11411 2936
rect 11475 2872 11491 2936
rect 11555 2872 11571 2936
rect 11635 2872 11651 2936
rect 11715 2872 11731 2936
rect 11795 2872 11811 2936
rect 11875 2872 12017 2936
rect 12081 2872 12097 2936
rect 12161 2872 12177 2936
rect 12241 2872 12257 2936
rect 12321 2872 12337 2936
rect 12401 2872 12417 2936
rect 12481 2872 12623 2936
rect 12687 2872 12703 2936
rect 12767 2872 12783 2936
rect 12847 2872 12863 2936
rect 12927 2872 12943 2936
rect 13007 2872 13023 2936
rect 13087 2872 13229 2936
rect 13293 2872 13309 2936
rect 13373 2872 13389 2936
rect 13453 2872 13469 2936
rect 13533 2872 13549 2936
rect 13613 2872 13629 2936
rect 13693 2872 13835 2936
rect 13899 2872 13915 2936
rect 13979 2872 13995 2936
rect 14059 2872 14075 2936
rect 14139 2872 14155 2936
rect 14219 2872 14235 2936
rect 14299 2872 14441 2936
rect 14505 2872 14521 2936
rect 14585 2872 14601 2936
rect 14665 2872 14681 2936
rect 14745 2872 14761 2936
rect 14825 2872 14841 2936
rect 14905 2872 15047 2936
rect 15111 2872 15127 2936
rect 15191 2872 15207 2936
rect 15271 2872 15287 2936
rect 15351 2872 15367 2936
rect 15431 2872 15447 2936
rect 15511 2872 15993 2936
rect 9299 2870 15993 2872
rect 9299 2338 9761 2870
rect 9299 2274 9359 2338
rect 9423 2337 9634 2338
rect 9423 2274 9490 2337
rect 9299 2273 9490 2274
rect 9554 2274 9634 2337
rect 9698 2274 9761 2338
rect 9554 2273 9761 2274
rect 9299 2255 9761 2273
rect 9969 2716 10035 2806
rect 9969 2652 9970 2716
rect 10034 2652 10035 2716
rect 9969 2636 10035 2652
rect 9969 2572 9970 2636
rect 10034 2572 10035 2636
rect 9969 2556 10035 2572
rect 9969 2492 9970 2556
rect 10034 2492 10035 2556
rect 9969 2476 10035 2492
rect 9969 2412 9970 2476
rect 10034 2412 10035 2476
rect 9969 2396 10035 2412
rect 9969 2332 9970 2396
rect 10034 2332 10035 2396
rect 9969 2316 10035 2332
rect 9969 2252 9970 2316
rect 10034 2252 10035 2316
rect 9969 2236 10035 2252
rect 9969 2172 9970 2236
rect 10034 2172 10035 2236
rect 9969 2156 10035 2172
rect 9969 2092 9970 2156
rect 10034 2092 10035 2156
rect 9969 2076 10035 2092
rect 9969 2012 9970 2076
rect 10034 2012 10035 2076
rect 9969 1996 10035 2012
rect 9969 1932 9970 1996
rect 10034 1932 10035 1996
rect 9316 1792 9747 1807
rect 9316 1728 9377 1792
rect 9441 1728 9497 1792
rect 9561 1728 9640 1792
rect 9704 1728 9747 1792
rect 9316 1713 9747 1728
rect 9317 369 9747 1713
rect 9969 1778 10035 1932
rect 10095 1840 10155 2870
rect 10215 1778 10275 2810
rect 10335 1840 10395 2870
rect 10455 1778 10515 2810
rect 10575 2716 10641 2806
rect 10575 2652 10576 2716
rect 10640 2652 10641 2716
rect 10575 2636 10641 2652
rect 10575 2572 10576 2636
rect 10640 2572 10641 2636
rect 10575 2556 10641 2572
rect 10575 2492 10576 2556
rect 10640 2492 10641 2556
rect 10575 2476 10641 2492
rect 10575 2412 10576 2476
rect 10640 2412 10641 2476
rect 10575 2396 10641 2412
rect 10575 2332 10576 2396
rect 10640 2332 10641 2396
rect 10575 2316 10641 2332
rect 10575 2252 10576 2316
rect 10640 2252 10641 2316
rect 10575 2236 10641 2252
rect 10575 2172 10576 2236
rect 10640 2172 10641 2236
rect 10575 2156 10641 2172
rect 10575 2092 10576 2156
rect 10640 2092 10641 2156
rect 10575 2076 10641 2092
rect 10575 2012 10576 2076
rect 10640 2012 10641 2076
rect 10575 1996 10641 2012
rect 10575 1932 10576 1996
rect 10640 1932 10641 1996
rect 10575 1778 10641 1932
rect 9969 1776 10641 1778
rect 9969 1712 10073 1776
rect 10137 1712 10153 1776
rect 10217 1712 10233 1776
rect 10297 1712 10313 1776
rect 10377 1712 10393 1776
rect 10457 1712 10473 1776
rect 10537 1712 10641 1776
rect 9969 1710 10641 1712
rect 10701 2716 10767 2806
rect 10701 2652 10702 2716
rect 10766 2652 10767 2716
rect 10701 2636 10767 2652
rect 10701 2572 10702 2636
rect 10766 2572 10767 2636
rect 10701 2556 10767 2572
rect 10701 2492 10702 2556
rect 10766 2492 10767 2556
rect 10701 2476 10767 2492
rect 10701 2412 10702 2476
rect 10766 2412 10767 2476
rect 10701 2396 10767 2412
rect 10701 2332 10702 2396
rect 10766 2332 10767 2396
rect 10701 2316 10767 2332
rect 10701 2252 10702 2316
rect 10766 2252 10767 2316
rect 10701 2236 10767 2252
rect 10701 2172 10702 2236
rect 10766 2172 10767 2236
rect 10701 2156 10767 2172
rect 10701 2092 10702 2156
rect 10766 2092 10767 2156
rect 10701 2076 10767 2092
rect 10701 2012 10702 2076
rect 10766 2012 10767 2076
rect 10701 1996 10767 2012
rect 10701 1932 10702 1996
rect 10766 1932 10767 1996
rect 10701 1778 10767 1932
rect 10827 1840 10887 2870
rect 10947 1778 11007 2810
rect 11067 1840 11127 2870
rect 11187 1778 11247 2810
rect 11307 2716 11373 2806
rect 11307 2652 11308 2716
rect 11372 2652 11373 2716
rect 11307 2636 11373 2652
rect 11307 2572 11308 2636
rect 11372 2572 11373 2636
rect 11307 2556 11373 2572
rect 11307 2492 11308 2556
rect 11372 2492 11373 2556
rect 11307 2476 11373 2492
rect 11307 2412 11308 2476
rect 11372 2412 11373 2476
rect 11307 2396 11373 2412
rect 11307 2332 11308 2396
rect 11372 2332 11373 2396
rect 11307 2316 11373 2332
rect 11307 2252 11308 2316
rect 11372 2252 11373 2316
rect 11307 2236 11373 2252
rect 11307 2172 11308 2236
rect 11372 2172 11373 2236
rect 11307 2156 11373 2172
rect 11307 2092 11308 2156
rect 11372 2092 11373 2156
rect 11307 2076 11373 2092
rect 11307 2012 11308 2076
rect 11372 2012 11373 2076
rect 11307 1996 11373 2012
rect 11307 1932 11308 1996
rect 11372 1932 11373 1996
rect 11307 1778 11373 1932
rect 11433 1778 11493 2810
rect 11553 1840 11613 2870
rect 11673 1778 11733 2810
rect 11793 1840 11853 2870
rect 11913 2716 11979 2806
rect 11913 2652 11914 2716
rect 11978 2652 11979 2716
rect 11913 2636 11979 2652
rect 11913 2572 11914 2636
rect 11978 2572 11979 2636
rect 11913 2556 11979 2572
rect 11913 2492 11914 2556
rect 11978 2492 11979 2556
rect 11913 2476 11979 2492
rect 11913 2412 11914 2476
rect 11978 2412 11979 2476
rect 11913 2396 11979 2412
rect 11913 2332 11914 2396
rect 11978 2332 11979 2396
rect 11913 2316 11979 2332
rect 11913 2252 11914 2316
rect 11978 2252 11979 2316
rect 11913 2236 11979 2252
rect 11913 2172 11914 2236
rect 11978 2172 11979 2236
rect 11913 2156 11979 2172
rect 11913 2092 11914 2156
rect 11978 2092 11979 2156
rect 11913 2076 11979 2092
rect 11913 2012 11914 2076
rect 11978 2012 11979 2076
rect 11913 1996 11979 2012
rect 11913 1932 11914 1996
rect 11978 1932 11979 1996
rect 11913 1778 11979 1932
rect 12039 1840 12099 2870
rect 12159 1778 12219 2810
rect 12279 1840 12339 2870
rect 12399 1778 12459 2810
rect 12519 2716 12585 2806
rect 12519 2652 12520 2716
rect 12584 2652 12585 2716
rect 12519 2636 12585 2652
rect 12519 2572 12520 2636
rect 12584 2572 12585 2636
rect 12519 2556 12585 2572
rect 12519 2492 12520 2556
rect 12584 2492 12585 2556
rect 12519 2476 12585 2492
rect 12519 2412 12520 2476
rect 12584 2412 12585 2476
rect 12519 2396 12585 2412
rect 12519 2332 12520 2396
rect 12584 2332 12585 2396
rect 12519 2316 12585 2332
rect 12519 2252 12520 2316
rect 12584 2252 12585 2316
rect 12519 2236 12585 2252
rect 12519 2172 12520 2236
rect 12584 2172 12585 2236
rect 12519 2156 12585 2172
rect 12519 2092 12520 2156
rect 12584 2092 12585 2156
rect 12519 2076 12585 2092
rect 12519 2012 12520 2076
rect 12584 2012 12585 2076
rect 12519 1996 12585 2012
rect 12519 1932 12520 1996
rect 12584 1932 12585 1996
rect 12519 1778 12585 1932
rect 12645 1778 12705 2810
rect 12765 1840 12825 2870
rect 12885 1778 12945 2810
rect 13005 1840 13065 2870
rect 13125 2716 13191 2806
rect 13125 2652 13126 2716
rect 13190 2652 13191 2716
rect 13125 2636 13191 2652
rect 13125 2572 13126 2636
rect 13190 2572 13191 2636
rect 13125 2556 13191 2572
rect 13125 2492 13126 2556
rect 13190 2492 13191 2556
rect 13125 2476 13191 2492
rect 13125 2412 13126 2476
rect 13190 2412 13191 2476
rect 13125 2396 13191 2412
rect 13125 2332 13126 2396
rect 13190 2332 13191 2396
rect 13125 2316 13191 2332
rect 13125 2252 13126 2316
rect 13190 2252 13191 2316
rect 13125 2236 13191 2252
rect 13125 2172 13126 2236
rect 13190 2172 13191 2236
rect 13125 2156 13191 2172
rect 13125 2092 13126 2156
rect 13190 2092 13191 2156
rect 13125 2076 13191 2092
rect 13125 2012 13126 2076
rect 13190 2012 13191 2076
rect 13125 1996 13191 2012
rect 13125 1932 13126 1996
rect 13190 1932 13191 1996
rect 13125 1778 13191 1932
rect 13251 1840 13311 2870
rect 13371 1778 13431 2810
rect 13491 1840 13551 2870
rect 13611 1778 13671 2810
rect 13731 2716 13797 2806
rect 13731 2652 13732 2716
rect 13796 2652 13797 2716
rect 13731 2636 13797 2652
rect 13731 2572 13732 2636
rect 13796 2572 13797 2636
rect 13731 2556 13797 2572
rect 13731 2492 13732 2556
rect 13796 2492 13797 2556
rect 13731 2476 13797 2492
rect 13731 2412 13732 2476
rect 13796 2412 13797 2476
rect 13731 2396 13797 2412
rect 13731 2332 13732 2396
rect 13796 2332 13797 2396
rect 13731 2316 13797 2332
rect 13731 2252 13732 2316
rect 13796 2252 13797 2316
rect 13731 2236 13797 2252
rect 13731 2172 13732 2236
rect 13796 2172 13797 2236
rect 13731 2156 13797 2172
rect 13731 2092 13732 2156
rect 13796 2092 13797 2156
rect 13731 2076 13797 2092
rect 13731 2012 13732 2076
rect 13796 2012 13797 2076
rect 13731 1996 13797 2012
rect 13731 1932 13732 1996
rect 13796 1932 13797 1996
rect 13731 1778 13797 1932
rect 13857 1778 13917 2810
rect 13977 1840 14037 2870
rect 14097 1778 14157 2810
rect 14217 1840 14277 2870
rect 14337 2716 14403 2806
rect 14337 2652 14338 2716
rect 14402 2652 14403 2716
rect 14337 2636 14403 2652
rect 14337 2572 14338 2636
rect 14402 2572 14403 2636
rect 14337 2556 14403 2572
rect 14337 2492 14338 2556
rect 14402 2492 14403 2556
rect 14337 2476 14403 2492
rect 14337 2412 14338 2476
rect 14402 2412 14403 2476
rect 14337 2396 14403 2412
rect 14337 2332 14338 2396
rect 14402 2332 14403 2396
rect 14337 2316 14403 2332
rect 14337 2252 14338 2316
rect 14402 2252 14403 2316
rect 14337 2236 14403 2252
rect 14337 2172 14338 2236
rect 14402 2172 14403 2236
rect 14337 2156 14403 2172
rect 14337 2092 14338 2156
rect 14402 2092 14403 2156
rect 14337 2076 14403 2092
rect 14337 2012 14338 2076
rect 14402 2012 14403 2076
rect 14337 1996 14403 2012
rect 14337 1932 14338 1996
rect 14402 1932 14403 1996
rect 14337 1778 14403 1932
rect 14463 1840 14523 2870
rect 14583 1778 14643 2810
rect 14703 1840 14763 2870
rect 14823 1778 14883 2810
rect 14943 2716 15009 2806
rect 14943 2652 14944 2716
rect 15008 2652 15009 2716
rect 14943 2636 15009 2652
rect 14943 2572 14944 2636
rect 15008 2572 15009 2636
rect 14943 2556 15009 2572
rect 14943 2492 14944 2556
rect 15008 2492 15009 2556
rect 14943 2476 15009 2492
rect 14943 2412 14944 2476
rect 15008 2412 15009 2476
rect 14943 2396 15009 2412
rect 14943 2332 14944 2396
rect 15008 2332 15009 2396
rect 14943 2316 15009 2332
rect 14943 2252 14944 2316
rect 15008 2252 15009 2316
rect 14943 2236 15009 2252
rect 14943 2172 14944 2236
rect 15008 2172 15009 2236
rect 14943 2156 15009 2172
rect 14943 2092 14944 2156
rect 15008 2092 15009 2156
rect 14943 2076 15009 2092
rect 14943 2012 14944 2076
rect 15008 2012 15009 2076
rect 14943 1996 15009 2012
rect 14943 1932 14944 1996
rect 15008 1932 15009 1996
rect 14943 1778 15009 1932
rect 15069 1778 15129 2810
rect 15189 1840 15249 2870
rect 15309 1778 15369 2810
rect 15429 1840 15489 2870
rect 15549 2716 15615 2806
rect 15549 2652 15550 2716
rect 15614 2652 15615 2716
rect 15549 2636 15615 2652
rect 15549 2572 15550 2636
rect 15614 2572 15615 2636
rect 15549 2556 15615 2572
rect 15549 2492 15550 2556
rect 15614 2492 15615 2556
rect 15549 2476 15615 2492
rect 15549 2412 15550 2476
rect 15614 2412 15615 2476
rect 15549 2396 15615 2412
rect 15549 2332 15550 2396
rect 15614 2332 15615 2396
rect 15549 2316 15615 2332
rect 15549 2252 15550 2316
rect 15614 2252 15615 2316
rect 15549 2236 15615 2252
rect 15549 2172 15550 2236
rect 15614 2172 15615 2236
rect 15549 2156 15615 2172
rect 15549 2092 15550 2156
rect 15614 2092 15615 2156
rect 15549 2076 15615 2092
rect 15549 2012 15550 2076
rect 15614 2012 15615 2076
rect 15549 1996 15615 2012
rect 15549 1932 15550 1996
rect 15614 1932 15615 1996
rect 15675 2016 15993 2870
rect 15675 1952 15708 2016
rect 15772 1952 15993 2016
rect 15675 1940 15993 1952
rect 15549 1778 15615 1932
rect 10701 1776 15615 1778
rect 10701 1712 10805 1776
rect 10869 1712 10885 1776
rect 10949 1712 10965 1776
rect 11029 1712 11045 1776
rect 11109 1712 11125 1776
rect 11189 1712 11205 1776
rect 11269 1712 11411 1776
rect 11475 1712 11491 1776
rect 11555 1712 11571 1776
rect 11635 1712 11651 1776
rect 11715 1712 11731 1776
rect 11795 1712 11811 1776
rect 11875 1712 12017 1776
rect 12081 1712 12097 1776
rect 12161 1712 12177 1776
rect 12241 1712 12257 1776
rect 12321 1712 12337 1776
rect 12401 1712 12417 1776
rect 12481 1712 12623 1776
rect 12687 1712 12703 1776
rect 12767 1712 12783 1776
rect 12847 1712 12863 1776
rect 12927 1712 12943 1776
rect 13007 1712 13023 1776
rect 13087 1712 13229 1776
rect 13293 1712 13309 1776
rect 13373 1712 13389 1776
rect 13453 1712 13469 1776
rect 13533 1712 13549 1776
rect 13613 1712 13629 1776
rect 13693 1712 13835 1776
rect 13899 1712 13915 1776
rect 13979 1712 13995 1776
rect 14059 1712 14075 1776
rect 14139 1712 14155 1776
rect 14219 1712 14235 1776
rect 14299 1712 14441 1776
rect 14505 1712 14521 1776
rect 14585 1712 14601 1776
rect 14665 1712 14681 1776
rect 14745 1712 14761 1776
rect 14825 1712 14841 1776
rect 14905 1712 15047 1776
rect 15111 1712 15127 1776
rect 15191 1712 15207 1776
rect 15271 1712 15287 1776
rect 15351 1712 15367 1776
rect 15431 1712 15447 1776
rect 15511 1712 15615 1776
rect 10701 1710 15615 1712
rect 15675 1755 15873 1765
rect 15675 1691 15796 1755
rect 15860 1691 15873 1755
rect 15675 1681 15873 1691
rect 10323 1527 10995 1529
rect 10323 1463 10427 1527
rect 10491 1463 10507 1527
rect 10571 1463 10587 1527
rect 10651 1463 10667 1527
rect 10731 1463 10747 1527
rect 10811 1463 10827 1527
rect 10891 1463 10995 1527
rect 10323 1461 10995 1463
rect 10323 1307 10389 1461
rect 10323 1243 10324 1307
rect 10388 1243 10389 1307
rect 10323 1227 10389 1243
rect 10323 1163 10324 1227
rect 10388 1163 10389 1227
rect 10323 1147 10389 1163
rect 10323 1083 10324 1147
rect 10388 1083 10389 1147
rect 10323 1067 10389 1083
rect 10323 1003 10324 1067
rect 10388 1003 10389 1067
rect 10323 987 10389 1003
rect 10323 923 10324 987
rect 10388 923 10389 987
rect 10323 907 10389 923
rect 10323 843 10324 907
rect 10388 843 10389 907
rect 10323 827 10389 843
rect 10323 763 10324 827
rect 10388 763 10389 827
rect 10323 747 10389 763
rect 10323 683 10324 747
rect 10388 683 10389 747
rect 10323 667 10389 683
rect 10323 603 10324 667
rect 10388 603 10389 667
rect 10323 587 10389 603
rect 10323 523 10324 587
rect 10388 523 10389 587
rect 10323 433 10389 523
rect 9932 369 10057 375
rect 10449 369 10509 1399
rect 10569 429 10629 1461
rect 10689 369 10749 1399
rect 10809 429 10869 1461
rect 10929 1307 10995 1461
rect 10929 1243 10930 1307
rect 10994 1243 10995 1307
rect 10929 1227 10995 1243
rect 10929 1163 10930 1227
rect 10994 1163 10995 1227
rect 10929 1147 10995 1163
rect 10929 1083 10930 1147
rect 10994 1083 10995 1147
rect 10929 1067 10995 1083
rect 10929 1003 10930 1067
rect 10994 1003 10995 1067
rect 10929 987 10995 1003
rect 10929 923 10930 987
rect 10994 923 10995 987
rect 10929 907 10995 923
rect 10929 843 10930 907
rect 10994 843 10995 907
rect 10929 827 10995 843
rect 10929 763 10930 827
rect 10994 763 10995 827
rect 10929 747 10995 763
rect 10929 683 10930 747
rect 10994 683 10995 747
rect 10929 667 10995 683
rect 10929 603 10930 667
rect 10994 603 10995 667
rect 10929 587 10995 603
rect 10929 523 10930 587
rect 10994 523 10995 587
rect 10929 433 10995 523
rect 11055 1527 13545 1529
rect 11055 1463 11159 1527
rect 11223 1463 11239 1527
rect 11303 1463 11319 1527
rect 11383 1463 11399 1527
rect 11463 1463 11479 1527
rect 11543 1463 11559 1527
rect 11623 1463 11765 1527
rect 11829 1463 11845 1527
rect 11909 1463 11925 1527
rect 11989 1463 12005 1527
rect 12069 1463 12085 1527
rect 12149 1463 12165 1527
rect 12229 1463 12371 1527
rect 12435 1463 12451 1527
rect 12515 1463 12531 1527
rect 12595 1463 12611 1527
rect 12675 1463 12691 1527
rect 12755 1463 12771 1527
rect 12835 1463 12977 1527
rect 13041 1463 13057 1527
rect 13121 1463 13137 1527
rect 13201 1463 13217 1527
rect 13281 1463 13297 1527
rect 13361 1463 13377 1527
rect 13441 1463 13545 1527
rect 11055 1461 13545 1463
rect 11055 1307 11121 1461
rect 11055 1243 11056 1307
rect 11120 1243 11121 1307
rect 11055 1227 11121 1243
rect 11055 1163 11056 1227
rect 11120 1163 11121 1227
rect 11055 1147 11121 1163
rect 11055 1083 11056 1147
rect 11120 1083 11121 1147
rect 11055 1067 11121 1083
rect 11055 1003 11056 1067
rect 11120 1003 11121 1067
rect 11055 987 11121 1003
rect 11055 923 11056 987
rect 11120 923 11121 987
rect 11055 907 11121 923
rect 11055 843 11056 907
rect 11120 843 11121 907
rect 11055 827 11121 843
rect 11055 763 11056 827
rect 11120 763 11121 827
rect 11055 747 11121 763
rect 11055 683 11056 747
rect 11120 683 11121 747
rect 11055 667 11121 683
rect 11055 603 11056 667
rect 11120 603 11121 667
rect 11055 587 11121 603
rect 11055 523 11056 587
rect 11120 523 11121 587
rect 11055 433 11121 523
rect 11181 369 11241 1399
rect 11301 429 11361 1461
rect 11421 369 11481 1399
rect 11541 429 11601 1461
rect 11661 1307 11727 1461
rect 11661 1243 11662 1307
rect 11726 1243 11727 1307
rect 11661 1227 11727 1243
rect 11661 1163 11662 1227
rect 11726 1163 11727 1227
rect 11661 1147 11727 1163
rect 11661 1083 11662 1147
rect 11726 1083 11727 1147
rect 11661 1067 11727 1083
rect 11661 1003 11662 1067
rect 11726 1003 11727 1067
rect 11661 987 11727 1003
rect 11661 923 11662 987
rect 11726 923 11727 987
rect 11661 907 11727 923
rect 11661 843 11662 907
rect 11726 843 11727 907
rect 11661 827 11727 843
rect 11661 763 11662 827
rect 11726 763 11727 827
rect 11661 747 11727 763
rect 11661 683 11662 747
rect 11726 683 11727 747
rect 11661 667 11727 683
rect 11661 603 11662 667
rect 11726 603 11727 667
rect 11661 587 11727 603
rect 11661 523 11662 587
rect 11726 523 11727 587
rect 11661 433 11727 523
rect 11787 429 11847 1461
rect 11907 369 11967 1399
rect 12027 429 12087 1461
rect 12147 369 12207 1399
rect 12267 1307 12333 1461
rect 12267 1243 12268 1307
rect 12332 1243 12333 1307
rect 12267 1227 12333 1243
rect 12267 1163 12268 1227
rect 12332 1163 12333 1227
rect 12267 1147 12333 1163
rect 12267 1083 12268 1147
rect 12332 1083 12333 1147
rect 12267 1067 12333 1083
rect 12267 1003 12268 1067
rect 12332 1003 12333 1067
rect 12267 987 12333 1003
rect 12267 923 12268 987
rect 12332 923 12333 987
rect 12267 907 12333 923
rect 12267 843 12268 907
rect 12332 843 12333 907
rect 12267 827 12333 843
rect 12267 763 12268 827
rect 12332 763 12333 827
rect 12267 747 12333 763
rect 12267 683 12268 747
rect 12332 683 12333 747
rect 12267 667 12333 683
rect 12267 603 12268 667
rect 12332 603 12333 667
rect 12267 587 12333 603
rect 12267 523 12268 587
rect 12332 523 12333 587
rect 12267 433 12333 523
rect 12393 369 12453 1399
rect 12513 429 12573 1461
rect 12633 369 12693 1399
rect 12753 429 12813 1461
rect 12873 1307 12939 1461
rect 12873 1243 12874 1307
rect 12938 1243 12939 1307
rect 12873 1227 12939 1243
rect 12873 1163 12874 1227
rect 12938 1163 12939 1227
rect 12873 1147 12939 1163
rect 12873 1083 12874 1147
rect 12938 1083 12939 1147
rect 12873 1067 12939 1083
rect 12873 1003 12874 1067
rect 12938 1003 12939 1067
rect 12873 987 12939 1003
rect 12873 923 12874 987
rect 12938 923 12939 987
rect 12873 907 12939 923
rect 12873 843 12874 907
rect 12938 843 12939 907
rect 12873 827 12939 843
rect 12873 763 12874 827
rect 12938 763 12939 827
rect 12873 747 12939 763
rect 12873 683 12874 747
rect 12938 683 12939 747
rect 12873 667 12939 683
rect 12873 603 12874 667
rect 12938 603 12939 667
rect 12873 587 12939 603
rect 12873 523 12874 587
rect 12938 523 12939 587
rect 12873 433 12939 523
rect 12999 429 13059 1461
rect 13119 369 13179 1399
rect 13239 429 13299 1461
rect 13359 369 13419 1399
rect 13479 1307 13545 1461
rect 13479 1243 13480 1307
rect 13544 1243 13545 1307
rect 13479 1227 13545 1243
rect 13479 1163 13480 1227
rect 13544 1163 13545 1227
rect 13479 1147 13545 1163
rect 13479 1083 13480 1147
rect 13544 1083 13545 1147
rect 13479 1067 13545 1083
rect 13479 1003 13480 1067
rect 13544 1003 13545 1067
rect 13479 987 13545 1003
rect 13479 923 13480 987
rect 13544 923 13545 987
rect 13479 907 13545 923
rect 13479 843 13480 907
rect 13544 843 13545 907
rect 13479 827 13545 843
rect 13479 763 13480 827
rect 13544 763 13545 827
rect 13479 747 13545 763
rect 13479 683 13480 747
rect 13544 683 13545 747
rect 13479 667 13545 683
rect 13479 603 13480 667
rect 13544 603 13545 667
rect 13479 587 13545 603
rect 13479 523 13480 587
rect 13544 523 13545 587
rect 13479 433 13545 523
rect 13605 1527 14883 1529
rect 13605 1463 13709 1527
rect 13773 1463 13789 1527
rect 13853 1463 13869 1527
rect 13933 1463 13949 1527
rect 14013 1463 14029 1527
rect 14093 1463 14109 1527
rect 14173 1463 14315 1527
rect 14379 1463 14395 1527
rect 14459 1463 14475 1527
rect 14539 1463 14555 1527
rect 14619 1463 14635 1527
rect 14699 1463 14715 1527
rect 14779 1463 14883 1527
rect 13605 1461 14883 1463
rect 13605 1307 13671 1461
rect 13605 1243 13606 1307
rect 13670 1243 13671 1307
rect 13605 1227 13671 1243
rect 13605 1163 13606 1227
rect 13670 1163 13671 1227
rect 13605 1147 13671 1163
rect 13605 1083 13606 1147
rect 13670 1083 13671 1147
rect 13605 1067 13671 1083
rect 13605 1003 13606 1067
rect 13670 1003 13671 1067
rect 13605 987 13671 1003
rect 13605 923 13606 987
rect 13670 923 13671 987
rect 13605 907 13671 923
rect 13605 843 13606 907
rect 13670 843 13671 907
rect 13605 827 13671 843
rect 13605 763 13606 827
rect 13670 763 13671 827
rect 13605 747 13671 763
rect 13605 683 13606 747
rect 13670 683 13671 747
rect 13605 667 13671 683
rect 13605 603 13606 667
rect 13670 603 13671 667
rect 13605 587 13671 603
rect 13605 523 13606 587
rect 13670 523 13671 587
rect 13605 433 13671 523
rect 13731 369 13791 1399
rect 13851 429 13911 1461
rect 13971 369 14031 1399
rect 14091 429 14151 1461
rect 14211 1307 14277 1461
rect 14211 1243 14212 1307
rect 14276 1243 14277 1307
rect 14211 1227 14277 1243
rect 14211 1163 14212 1227
rect 14276 1163 14277 1227
rect 14211 1147 14277 1163
rect 14211 1083 14212 1147
rect 14276 1083 14277 1147
rect 14211 1067 14277 1083
rect 14211 1003 14212 1067
rect 14276 1003 14277 1067
rect 14211 987 14277 1003
rect 14211 923 14212 987
rect 14276 923 14277 987
rect 14211 907 14277 923
rect 14211 843 14212 907
rect 14276 843 14277 907
rect 14211 827 14277 843
rect 14211 763 14212 827
rect 14276 763 14277 827
rect 14211 747 14277 763
rect 14211 683 14212 747
rect 14276 683 14277 747
rect 14211 667 14277 683
rect 14211 603 14212 667
rect 14276 603 14277 667
rect 14211 587 14277 603
rect 14211 523 14212 587
rect 14276 523 14277 587
rect 14211 433 14277 523
rect 14337 429 14397 1461
rect 14457 369 14517 1399
rect 14577 429 14637 1461
rect 14697 369 14757 1399
rect 14817 1307 14883 1461
rect 14817 1243 14818 1307
rect 14882 1243 14883 1307
rect 14817 1227 14883 1243
rect 14817 1163 14818 1227
rect 14882 1163 14883 1227
rect 14817 1147 14883 1163
rect 14817 1083 14818 1147
rect 14882 1083 14883 1147
rect 14817 1067 14883 1083
rect 14817 1003 14818 1067
rect 14882 1003 14883 1067
rect 14817 987 14883 1003
rect 14817 923 14818 987
rect 14882 923 14883 987
rect 14817 907 14883 923
rect 14817 843 14818 907
rect 14882 843 14883 907
rect 14817 827 14883 843
rect 14817 763 14818 827
rect 14882 763 14883 827
rect 14817 747 14883 763
rect 14817 683 14818 747
rect 14882 683 14883 747
rect 14817 667 14883 683
rect 14817 603 14818 667
rect 14882 603 14883 667
rect 14817 587 14883 603
rect 14817 523 14818 587
rect 14882 523 14883 587
rect 14817 433 14883 523
rect 14943 1527 15615 1529
rect 14943 1463 15047 1527
rect 15111 1463 15127 1527
rect 15191 1463 15207 1527
rect 15271 1463 15287 1527
rect 15351 1463 15367 1527
rect 15431 1463 15447 1527
rect 15511 1463 15615 1527
rect 14943 1461 15615 1463
rect 14943 1307 15009 1461
rect 14943 1243 14944 1307
rect 15008 1243 15009 1307
rect 14943 1227 15009 1243
rect 14943 1163 14944 1227
rect 15008 1163 15009 1227
rect 14943 1147 15009 1163
rect 14943 1083 14944 1147
rect 15008 1083 15009 1147
rect 14943 1067 15009 1083
rect 14943 1003 14944 1067
rect 15008 1003 15009 1067
rect 14943 987 15009 1003
rect 14943 923 14944 987
rect 15008 923 15009 987
rect 14943 907 15009 923
rect 14943 843 14944 907
rect 15008 843 15009 907
rect 14943 827 15009 843
rect 14943 763 14944 827
rect 15008 763 15009 827
rect 14943 747 15009 763
rect 14943 683 14944 747
rect 15008 683 15009 747
rect 14943 667 15009 683
rect 14943 603 14944 667
rect 15008 603 15009 667
rect 14943 587 15009 603
rect 14943 523 14944 587
rect 15008 523 15009 587
rect 14943 433 15009 523
rect 15069 429 15129 1461
rect 15189 369 15249 1399
rect 15309 429 15369 1461
rect 15429 369 15489 1399
rect 15549 1307 15615 1461
rect 15549 1243 15550 1307
rect 15614 1243 15615 1307
rect 15549 1227 15615 1243
rect 15549 1163 15550 1227
rect 15614 1163 15615 1227
rect 15549 1147 15615 1163
rect 15549 1083 15550 1147
rect 15614 1083 15615 1147
rect 15549 1067 15615 1083
rect 15549 1003 15550 1067
rect 15614 1003 15615 1067
rect 15549 987 15615 1003
rect 15549 923 15550 987
rect 15614 923 15615 987
rect 15549 907 15615 923
rect 15549 843 15550 907
rect 15614 843 15615 907
rect 15549 827 15615 843
rect 15549 763 15550 827
rect 15614 763 15615 827
rect 15549 747 15615 763
rect 15549 683 15550 747
rect 15614 683 15615 747
rect 15549 667 15615 683
rect 15549 603 15550 667
rect 15614 603 15615 667
rect 15549 587 15615 603
rect 15549 523 15550 587
rect 15614 523 15615 587
rect 15549 433 15615 523
rect 15675 1300 15735 1681
rect 15933 1562 15993 1940
rect 15795 1552 15993 1562
rect 15795 1488 15796 1552
rect 15860 1488 15993 1552
rect 15795 1478 15993 1488
rect 15675 1290 15993 1300
rect 15675 1226 15705 1290
rect 15769 1226 15993 1290
rect 15675 369 15993 1226
rect 9316 367 15993 369
rect 9316 365 10427 367
rect 9316 301 9962 365
rect 10026 303 10427 365
rect 10491 303 10507 367
rect 10571 303 10587 367
rect 10651 303 10667 367
rect 10731 303 10747 367
rect 10811 303 10827 367
rect 10891 303 11159 367
rect 11223 303 11239 367
rect 11303 303 11319 367
rect 11383 303 11399 367
rect 11463 303 11479 367
rect 11543 303 11559 367
rect 11623 303 11765 367
rect 11829 303 11845 367
rect 11909 303 11925 367
rect 11989 303 12005 367
rect 12069 303 12085 367
rect 12149 303 12165 367
rect 12229 303 12371 367
rect 12435 303 12451 367
rect 12515 303 12531 367
rect 12595 303 12611 367
rect 12675 303 12691 367
rect 12755 303 12771 367
rect 12835 303 12977 367
rect 13041 303 13057 367
rect 13121 303 13137 367
rect 13201 303 13217 367
rect 13281 303 13297 367
rect 13361 303 13377 367
rect 13441 303 13709 367
rect 13773 303 13789 367
rect 13853 303 13869 367
rect 13933 303 13949 367
rect 14013 303 14029 367
rect 14093 303 14109 367
rect 14173 303 14315 367
rect 14379 303 14395 367
rect 14459 303 14475 367
rect 14539 303 14555 367
rect 14619 303 14635 367
rect 14699 303 14715 367
rect 14779 303 15047 367
rect 15111 303 15127 367
rect 15191 303 15207 367
rect 15271 303 15287 367
rect 15351 303 15367 367
rect 15431 303 15447 367
rect 15511 303 15993 367
rect 10026 301 15993 303
rect 9316 291 15993 301
rect 9316 289 9812 291
<< labels >>
flabel metal1 9275 1596 9943 1643 0 FreeSans 320 0 0 0 IN
port 1 nsew
flabel metal1 15751 1594 15933 1640 0 FreeSans 320 0 0 0 OUT
port 2 nsew
flabel metal4 9299 2338 9761 2948 0 FreeSans 320 0 0 0 VDD
port 3 nsew
flabel metal4 9317 289 9747 1728 0 FreeSans 320 0 0 0 VSS
port 4 nsew
flabel metal1 9238 1979 9376 2013 0 FreeSans 320 0 0 0 code[3]
port 5 nsew
flabel metal1 9256 1393 9650 1440 0 FreeSans 320 0 0 0 code_offset
port 6 nsew
flabel metal1 15009 267 15067 1423 0 FreeSans 320 0 0 0 code[0]
port 7 nsew
flabel metal1 14153 268 14211 1445 0 FreeSans 320 0 0 0 code[1]
port 8 nsew
flabel metal1 11727 268 11785 1445 0 FreeSans 320 0 0 0 code[2]
port 10 nsew
flabel poly 9863 1392 9965 1422 0 FreeSans 320 0 0 0 x9.input_stack
flabel space 9977 1305 10011 1365 0 FreeSans 320 0 0 0 x9.output_stack
flabel space 9977 339 10011 399 0 FreeSans 320 0 0 0 x9.vss
flabel space 10569 429 10629 1463 0 FreeSans 320 0 0 0 x7.CBOT
flabel space 10689 367 10749 1399 0 FreeSans 320 0 0 0 x7.CTOP
flabel space 10575 669 10745 839 0 FreeSans 320 0 0 0 x7.SUB
flabel space 10883 1405 10917 1439 0 FreeSans 320 0 0 0 x7.SW
flabel metal4 10585 1051 10611 1083 0 FreeSans 320 0 0 0 x7.x2.CBOT
flabel metal4 10703 461 10729 493 0 FreeSans 320 0 0 0 x7.x2.CTOP
flabel pwell 10575 669 10745 839 0 FreeSans 320 0 0 0 x7.x2.SUB
flabel space 11301 429 11361 1463 0 FreeSans 320 0 0 0 x4[3].CBOT
flabel space 11421 367 11481 1399 0 FreeSans 320 0 0 0 x4[3].CTOP
flabel space 11307 669 11477 839 0 FreeSans 320 0 0 0 x4[3].SUB
flabel space 11615 1405 11649 1439 0 FreeSans 320 0 0 0 x4[3].SW
flabel metal4 11317 1051 11343 1083 0 FreeSans 320 0 0 0 x4[3].x2.CBOT
flabel metal4 11435 461 11461 493 0 FreeSans 320 0 0 0 x4[3].x2.CTOP
flabel pwell 11307 669 11477 839 0 FreeSans 320 0 0 0 x4[3].x2.SUB
flabel space 12027 429 12087 1463 0 FreeSans 320 0 0 0 x4[2].CBOT
flabel space 11907 367 11967 1399 0 FreeSans 320 0 0 0 x4[2].CTOP
flabel space 11911 669 12081 839 0 FreeSans 320 0 0 0 x4[2].SUB
flabel space 11739 1405 11773 1439 0 FreeSans 320 0 0 0 x4[2].SW
flabel metal4 12045 1051 12071 1083 0 FreeSans 320 0 0 0 x4[2].x2.CBOT
flabel metal4 11927 461 11953 493 0 FreeSans 320 0 0 0 x4[2].x2.CTOP
flabel pwell 11911 669 12081 839 0 FreeSans 320 0 0 0 x4[2].x2.SUB
flabel space 12513 429 12573 1463 0 FreeSans 320 0 0 0 x4[1].CBOT
flabel space 12633 367 12693 1399 0 FreeSans 320 0 0 0 x4[1].CTOP
flabel space 12519 669 12689 839 0 FreeSans 320 0 0 0 x4[1].SUB
flabel space 12827 1405 12861 1439 0 FreeSans 320 0 0 0 x4[1].SW
flabel metal4 12529 1051 12555 1083 0 FreeSans 320 0 0 0 x4[1].x2.CBOT
flabel metal4 12647 461 12673 493 0 FreeSans 320 0 0 0 x4[1].x2.CTOP
flabel pwell 12519 669 12689 839 0 FreeSans 320 0 0 0 x4[1].x2.SUB
flabel space 13239 429 13299 1463 0 FreeSans 320 0 0 0 x4[0].CBOT
flabel space 13119 367 13179 1399 0 FreeSans 320 0 0 0 x4[0].CTOP
flabel space 13123 669 13293 839 0 FreeSans 320 0 0 0 x4[0].SUB
flabel space 12951 1405 12985 1439 0 FreeSans 320 0 0 0 x4[0].SW
flabel metal4 13257 1051 13283 1083 0 FreeSans 320 0 0 0 x4[0].x2.CBOT
flabel metal4 13139 461 13165 493 0 FreeSans 320 0 0 0 x4[0].x2.CTOP
flabel pwell 13123 669 13293 839 0 FreeSans 320 0 0 0 x4[0].x2.SUB
flabel space 13851 429 13911 1463 0 FreeSans 320 0 0 0 x3[1].CBOT
flabel space 13971 367 14031 1399 0 FreeSans 320 0 0 0 x3[1].CTOP
flabel space 13857 669 14027 839 0 FreeSans 320 0 0 0 x3[1].SUB
flabel space 14165 1405 14199 1439 0 FreeSans 320 0 0 0 x3[1].SW
flabel metal4 13867 1051 13893 1083 0 FreeSans 320 0 0 0 x3[1].x2.CBOT
flabel metal4 13985 461 14011 493 0 FreeSans 320 0 0 0 x3[1].x2.CTOP
flabel pwell 13857 669 14027 839 0 FreeSans 320 0 0 0 x3[1].x2.SUB
flabel space 14577 429 14637 1463 0 FreeSans 320 0 0 0 x3[0].CBOT
flabel space 14457 367 14517 1399 0 FreeSans 320 0 0 0 x3[0].CTOP
flabel space 14461 669 14631 839 0 FreeSans 320 0 0 0 x3[0].SUB
flabel space 14289 1405 14323 1439 0 FreeSans 320 0 0 0 x3[0].SW
flabel metal4 14595 1051 14621 1083 0 FreeSans 320 0 0 0 x3[0].x2.CBOT
flabel metal4 14477 461 14503 493 0 FreeSans 320 0 0 0 x3[0].x2.CTOP
flabel pwell 14461 669 14631 839 0 FreeSans 320 0 0 0 x3[0].x2.SUB
flabel space 15309 429 15369 1463 0 FreeSans 320 0 0 0 x2.CBOT
flabel space 15189 367 15249 1399 0 FreeSans 320 0 0 0 x2.CTOP
flabel space 15193 669 15363 839 0 FreeSans 320 0 0 0 x2.SUB
flabel space 15021 1405 15055 1439 0 FreeSans 320 0 0 0 x2.SW
flabel metal4 15327 1051 15353 1083 0 FreeSans 320 0 0 0 x2.x2.CBOT
flabel metal4 15209 461 15235 493 0 FreeSans 320 0 0 0 x2.x2.CTOP
flabel pwell 15193 669 15363 839 0 FreeSans 320 0 0 0 x2.x2.SUB
flabel locali 9464 2049 9498 2083 0 FreeSans 340 0 0 0 x1.Y
flabel locali 9464 1981 9498 2015 0 FreeSans 340 0 0 0 x1.Y
flabel locali 9372 1981 9406 2015 0 FreeSans 340 0 0 0 x1.A
flabel metal1 9329 1743 9363 1777 0 FreeSans 200 0 0 0 x1.VGND
flabel metal1 9329 2287 9363 2321 0 FreeSans 200 0 0 0 x1.VPWR
rlabel comment 9300 1760 9300 1760 4 x1.inv_1
rlabel metal1 9300 1712 9576 1808 1 x1.VGND
rlabel metal1 9300 2256 9576 2352 1 x1.VPWR
flabel pwell 9329 1743 9363 1777 0 FreeSans 200 0 0 0 x1.VNB
flabel nwell 9329 2287 9363 2321 0 FreeSans 200 0 0 0 x1.VPB
flabel locali 9562 2049 9596 2083 0 FreeSans 340 0 0 0 x5.Y
flabel locali 9562 1981 9596 2015 0 FreeSans 340 0 0 0 x5.Y
flabel locali 9654 1981 9688 2015 0 FreeSans 340 0 0 0 x5.A
flabel metal1 9697 1743 9731 1777 0 FreeSans 200 0 0 0 x5.VGND
flabel metal1 9697 2287 9731 2321 0 FreeSans 200 0 0 0 x5.VPWR
rlabel comment 9760 1760 9760 1760 6 x5.inv_1
rlabel metal1 9484 1712 9760 1808 1 x5.VGND
rlabel metal1 9484 2256 9760 2352 1 x5.VPWR
flabel pwell 9697 1743 9731 1777 0 FreeSans 200 0 0 0 x5.VNB
flabel nwell 9697 2287 9731 2321 0 FreeSans 200 0 0 0 x5.VPB
flabel metal1 9907 2049 9941 2083 0 FreeSans 320 0 0 0 x8.input_stack
flabel space 9951 2832 9985 2892 0 FreeSans 320 0 0 0 x8.vdd
flabel space 9951 2142 9985 2202 0 FreeSans 320 0 0 0 x8.output_stack
flabel space 10221 2400 10391 2570 0 FreeSans 320 0 0 0 x6.SUB
flabel space 10215 1776 10275 2810 0 FreeSans 320 0 0 0 x6.CBOT
flabel space 10335 1840 10395 2872 0 FreeSans 320 0 0 0 x6.CTOP
flabel space 10528 1809 10562 1843 0 FreeSans 320 0 0 0 x6.SW
flabel metal4 10231 2156 10257 2188 0 FreeSans 320 0 0 0 x6.x1.CBOT
flabel metal4 10349 2746 10375 2778 0 FreeSans 320 0 0 0 x6.x1.CTOP
flabel nwell 10221 2400 10391 2570 0 FreeSans 320 0 0 0 x6.x1.SUB
flabel space 10953 2400 11123 2570 0 FreeSans 320 0 0 0 x5[7].SUB
flabel space 10947 1776 11007 2810 0 FreeSans 320 0 0 0 x5[7].CBOT
flabel space 11067 1840 11127 2872 0 FreeSans 320 0 0 0 x5[7].CTOP
flabel space 11260 1809 11294 1843 0 FreeSans 320 0 0 0 x5[7].SW
flabel metal4 10963 2156 10989 2188 0 FreeSans 320 0 0 0 x5[7].x1.CBOT
flabel metal4 11081 2746 11107 2778 0 FreeSans 320 0 0 0 x5[7].x1.CTOP
flabel nwell 10953 2400 11123 2570 0 FreeSans 320 0 0 0 x5[7].x1.SUB
flabel space 11557 2400 11727 2570 0 FreeSans 320 0 0 0 x5[6].SUB
flabel space 11673 1776 11733 2810 0 FreeSans 320 0 0 0 x5[6].CBOT
flabel space 11553 1840 11613 2872 0 FreeSans 320 0 0 0 x5[6].CTOP
flabel space 11386 1809 11420 1843 0 FreeSans 320 0 0 0 x5[6].SW
flabel metal4 11691 2156 11717 2188 0 FreeSans 320 0 0 0 x5[6].x1.CBOT
flabel metal4 11573 2746 11599 2778 0 FreeSans 320 0 0 0 x5[6].x1.CTOP
flabel nwell 11557 2400 11727 2570 0 FreeSans 320 0 0 0 x5[6].x1.SUB
flabel space 12165 2400 12335 2570 0 FreeSans 320 0 0 0 x5[5].SUB
flabel space 12159 1776 12219 2810 0 FreeSans 320 0 0 0 x5[5].CBOT
flabel space 12279 1840 12339 2872 0 FreeSans 320 0 0 0 x5[5].CTOP
flabel space 12472 1809 12506 1843 0 FreeSans 320 0 0 0 x5[5].SW
flabel metal4 12175 2156 12201 2188 0 FreeSans 320 0 0 0 x5[5].x1.CBOT
flabel metal4 12293 2746 12319 2778 0 FreeSans 320 0 0 0 x5[5].x1.CTOP
flabel nwell 12165 2400 12335 2570 0 FreeSans 320 0 0 0 x5[5].x1.SUB
flabel space 12769 2400 12939 2570 0 FreeSans 320 0 0 0 x5[4].SUB
flabel space 12885 1776 12945 2810 0 FreeSans 320 0 0 0 x5[4].CBOT
flabel space 12765 1840 12825 2872 0 FreeSans 320 0 0 0 x5[4].CTOP
flabel space 12598 1809 12632 1843 0 FreeSans 320 0 0 0 x5[4].SW
flabel metal4 12903 2156 12929 2188 0 FreeSans 320 0 0 0 x5[4].x1.CBOT
flabel metal4 12785 2746 12811 2778 0 FreeSans 320 0 0 0 x5[4].x1.CTOP
flabel nwell 12769 2400 12939 2570 0 FreeSans 320 0 0 0 x5[4].x1.SUB
flabel space 13377 2400 13547 2570 0 FreeSans 320 0 0 0 x5[3].SUB
flabel space 13371 1776 13431 2810 0 FreeSans 320 0 0 0 x5[3].CBOT
flabel space 13491 1840 13551 2872 0 FreeSans 320 0 0 0 x5[3].CTOP
flabel space 13684 1809 13718 1843 0 FreeSans 320 0 0 0 x5[3].SW
flabel metal4 13387 2156 13413 2188 0 FreeSans 320 0 0 0 x5[3].x1.CBOT
flabel metal4 13505 2746 13531 2778 0 FreeSans 320 0 0 0 x5[3].x1.CTOP
flabel nwell 13377 2400 13547 2570 0 FreeSans 320 0 0 0 x5[3].x1.SUB
flabel space 13981 2400 14151 2570 0 FreeSans 320 0 0 0 x5[2].SUB
flabel space 14097 1776 14157 2810 0 FreeSans 320 0 0 0 x5[2].CBOT
flabel space 13977 1840 14037 2872 0 FreeSans 320 0 0 0 x5[2].CTOP
flabel space 13810 1809 13844 1843 0 FreeSans 320 0 0 0 x5[2].SW
flabel metal4 14115 2156 14141 2188 0 FreeSans 320 0 0 0 x5[2].x1.CBOT
flabel metal4 13997 2746 14023 2778 0 FreeSans 320 0 0 0 x5[2].x1.CTOP
flabel nwell 13981 2400 14151 2570 0 FreeSans 320 0 0 0 x5[2].x1.SUB
flabel space 14589 2400 14759 2570 0 FreeSans 320 0 0 0 x5[1].SUB
flabel space 14583 1776 14643 2810 0 FreeSans 320 0 0 0 x5[1].CBOT
flabel space 14703 1840 14763 2872 0 FreeSans 320 0 0 0 x5[1].CTOP
flabel space 14896 1809 14930 1843 0 FreeSans 320 0 0 0 x5[1].SW
flabel metal4 14599 2156 14625 2188 0 FreeSans 320 0 0 0 x5[1].x1.CBOT
flabel metal4 14717 2746 14743 2778 0 FreeSans 320 0 0 0 x5[1].x1.CTOP
flabel nwell 14589 2400 14759 2570 0 FreeSans 320 0 0 0 x5[1].x1.SUB
flabel space 15193 2400 15363 2570 0 FreeSans 320 0 0 0 x5[0].SUB
flabel space 15309 1776 15369 2810 0 FreeSans 320 0 0 0 x5[0].CBOT
flabel space 15189 1840 15249 2872 0 FreeSans 320 0 0 0 x5[0].CTOP
flabel space 15022 1809 15056 1843 0 FreeSans 320 0 0 0 x5[0].SW
flabel metal4 15327 2156 15353 2188 0 FreeSans 320 0 0 0 x5[0].x1.CBOT
flabel metal4 15209 2746 15235 2778 0 FreeSans 320 0 0 0 x5[0].x1.CTOP
flabel nwell 15193 2400 15363 2570 0 FreeSans 320 0 0 0 x5[0].x1.SUB
<< end >>
