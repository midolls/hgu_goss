magic
tech sky130A
magscale 1 2
timestamp 1698839504
<< nmos >>
rect 143 757 173 841
rect 215 757 245 841
rect 143 619 173 703
rect 215 619 245 703
rect 143 481 173 565
rect 215 481 245 565
rect 143 343 173 427
rect 215 343 245 427
rect 143 205 173 289
rect 215 205 245 289
rect 143 67 173 151
rect 215 67 245 151
rect 143 -71 173 13
rect 215 -71 245 13
rect 143 -209 173 -125
rect 215 -209 245 -125
<< ndiff >>
rect 85 829 143 841
rect 85 769 97 829
rect 131 769 143 829
rect 85 757 143 769
rect 173 757 215 841
rect 245 829 303 841
rect 245 769 257 829
rect 291 769 303 829
rect 245 757 303 769
rect 85 691 143 703
rect 85 631 97 691
rect 131 631 143 691
rect 85 619 143 631
rect 173 619 215 703
rect 245 691 303 703
rect 245 631 257 691
rect 291 631 303 691
rect 245 619 303 631
rect 85 553 143 565
rect 85 493 97 553
rect 131 493 143 553
rect 85 481 143 493
rect 173 481 215 565
rect 245 553 303 565
rect 245 493 257 553
rect 291 493 303 553
rect 245 481 303 493
rect 85 415 143 427
rect 85 355 97 415
rect 131 355 143 415
rect 85 343 143 355
rect 173 343 215 427
rect 245 415 303 427
rect 245 355 257 415
rect 291 355 303 415
rect 245 343 303 355
rect 85 277 143 289
rect 85 217 97 277
rect 131 217 143 277
rect 85 205 143 217
rect 173 205 215 289
rect 245 277 303 289
rect 245 217 257 277
rect 291 217 303 277
rect 245 205 303 217
rect 85 139 143 151
rect 85 79 97 139
rect 131 79 143 139
rect 85 67 143 79
rect 173 67 215 151
rect 245 139 303 151
rect 245 79 257 139
rect 291 79 303 139
rect 245 67 303 79
rect 85 1 143 13
rect 85 -59 97 1
rect 131 -59 143 1
rect 85 -71 143 -59
rect 173 -71 215 13
rect 245 1 303 13
rect 245 -59 257 1
rect 291 -59 303 1
rect 245 -71 303 -59
rect 85 -137 143 -125
rect 85 -197 97 -137
rect 131 -197 143 -137
rect 85 -209 143 -197
rect 173 -209 215 -125
rect 245 -137 303 -125
rect 245 -197 257 -137
rect 291 -197 303 -137
rect 245 -209 303 -197
<< ndiffc >>
rect 97 769 131 829
rect 257 769 291 829
rect 97 631 131 691
rect 257 631 291 691
rect 97 493 131 553
rect 257 493 291 553
rect 97 355 131 415
rect 257 355 291 415
rect 97 217 131 277
rect 257 217 291 277
rect 97 79 131 139
rect 257 79 291 139
rect 97 -59 131 1
rect 257 -59 291 1
rect 97 -197 131 -137
rect 257 -197 291 -137
<< poly >>
rect 143 856 245 886
rect 143 841 173 856
rect 215 841 245 856
rect 143 703 173 757
rect 215 703 245 757
rect 143 565 173 619
rect 215 565 245 619
rect 143 427 173 481
rect 215 427 245 481
rect 143 289 173 343
rect 215 289 245 343
rect 143 151 173 205
rect 215 151 245 205
rect 143 13 173 67
rect 215 13 245 67
rect 143 -125 173 -71
rect 215 -125 245 -71
rect 143 -235 173 -209
rect 215 -235 245 -209
<< locali >>
rect 97 829 131 845
rect 97 753 131 769
rect 257 829 291 845
rect 257 753 291 769
rect 97 691 131 707
rect 97 615 131 631
rect 257 691 291 707
rect 257 615 291 631
rect 97 553 131 569
rect 97 477 131 493
rect 257 553 291 569
rect 257 477 291 493
rect 97 415 131 431
rect 97 339 131 355
rect 257 415 291 431
rect 257 339 291 355
rect 97 277 131 293
rect 97 201 131 217
rect 257 277 291 293
rect 257 201 291 217
rect 97 139 131 155
rect 97 63 131 79
rect 257 139 291 155
rect 257 63 291 79
rect 97 1 131 17
rect 97 -75 131 -59
rect 257 1 291 17
rect 257 -75 291 -59
rect 97 -137 131 -121
rect 97 -213 131 -197
rect 257 -137 291 -121
rect 257 -213 291 -197
<< viali >>
rect 97 769 131 829
rect 257 769 291 829
rect 97 631 131 691
rect 257 631 291 691
rect 97 493 131 553
rect 257 493 291 553
rect 97 355 131 415
rect 257 355 291 415
rect 97 217 131 277
rect 257 217 291 277
rect 97 79 131 139
rect 257 79 291 139
rect 97 -59 131 1
rect 257 -59 291 1
rect 97 -197 131 -137
rect 257 -197 291 -137
<< metal1 >>
rect 91 829 137 841
rect 91 769 97 829
rect 131 769 137 829
rect 91 757 137 769
rect 251 829 297 841
rect 251 769 257 829
rect 291 769 297 829
rect 91 691 137 703
rect 91 631 97 691
rect 131 631 137 691
rect 91 553 137 631
rect 251 691 297 769
rect 251 631 257 691
rect 291 631 297 691
rect 251 619 297 631
rect 91 493 97 553
rect 131 493 137 553
rect 91 481 137 493
rect 251 553 297 565
rect 251 493 257 553
rect 291 493 297 553
rect 91 415 137 427
rect 91 355 97 415
rect 131 355 137 415
rect 91 277 137 355
rect 251 415 297 493
rect 251 355 257 415
rect 291 355 297 415
rect 251 343 297 355
rect 91 217 97 277
rect 131 217 137 277
rect 91 205 137 217
rect 251 277 297 289
rect 251 217 257 277
rect 291 217 297 277
rect 91 139 137 151
rect 91 79 97 139
rect 131 79 137 139
rect 91 1 137 79
rect 251 139 297 217
rect 251 79 257 139
rect 291 79 297 139
rect 251 67 297 79
rect 91 -59 97 1
rect 131 -59 137 1
rect 91 -71 137 -59
rect 251 1 297 13
rect 251 -59 257 1
rect 291 -59 297 1
rect 91 -137 137 -125
rect 91 -197 97 -137
rect 131 -197 137 -137
rect 91 -209 137 -197
rect 251 -137 297 -59
rect 251 -197 257 -137
rect 291 -197 297 -137
rect 251 -209 297 -197
<< labels >>
flabel poly 143 856 245 886 0 FreeSans 320 0 0 0 input_stack
port 0 nsew
flabel space 97 769 131 829 0 FreeSans 320 0 0 0 output_stack
port 1 nsew
flabel space 97 -197 131 -137 0 FreeSans 320 0 0 0 vss
port 3 nsew
<< end >>
