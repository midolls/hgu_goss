../mag/hgu_sarlogic_flat.spice