magic
tech sky130A
magscale 1 2
timestamp 1699180127
<< psubdiff >>
rect 300 2029 348 2143
<< metal4 >>
rect 244 2488 280 2590
rect 364 2058 400 2148
rect 362 928 402 1006
use hgu_cdac_unit  x1
timestamp 1699173900
transform 1 0 -700 0 1 66
box 686 598 1358 1826
use hgu_cdac_unit  x2
timestamp 1699173900
transform -1 0 1344 0 -1 3650
box 686 598 1358 1826
<< labels >>
flabel psubdiff 300 2029 348 2143 0 FreeSans 160 0 0 0 SUB
port 1 nsew
flabel metal4 364 2058 400 2148 0 FreeSans 320 0 0 0 CBOT
port 4 nsew
flabel metal4 244 2488 280 2590 0 FreeSans 320 0 0 0 CTOP
port 6 nsew
flabel metal4 362 928 402 1006 0 FreeSans 320 0 0 0 CTOP
port 8 nsew
<< end >>
