magic
tech sky130A
magscale 1 2
timestamp 1699184006
<< error_p >>
rect 129 931 187 937
rect 129 897 141 931
rect 129 891 187 897
<< nwell >>
rect 48 349 268 898
rect -98 181 268 349
rect 48 40 268 181
<< pmoshvt >>
rect 143 766 173 850
rect 143 628 173 712
rect 143 490 173 574
rect 143 352 173 436
rect 143 214 173 298
rect 143 76 173 160
<< pdiff >>
rect 85 838 143 850
rect 85 778 97 838
rect 131 778 143 838
rect 85 766 143 778
rect 173 838 231 850
rect 173 778 185 838
rect 219 778 231 838
rect 173 766 231 778
rect 85 700 143 712
rect 85 640 97 700
rect 131 640 143 700
rect 85 628 143 640
rect 173 700 231 712
rect 173 640 185 700
rect 219 640 231 700
rect 173 628 231 640
rect 85 562 143 574
rect 85 502 97 562
rect 131 502 143 562
rect 85 490 143 502
rect 173 562 231 574
rect 173 502 185 562
rect 219 502 231 562
rect 173 490 231 502
rect 85 424 143 436
rect 85 364 97 424
rect 131 364 143 424
rect 85 352 143 364
rect 173 424 231 436
rect 173 364 185 424
rect 219 364 231 424
rect 173 352 231 364
rect 85 286 143 298
rect 85 226 97 286
rect 131 226 143 286
rect 85 214 143 226
rect 173 286 231 298
rect 173 226 185 286
rect 219 226 231 286
rect 173 214 231 226
rect 85 148 143 160
rect 85 88 97 148
rect 131 88 143 148
rect 85 76 143 88
rect 173 148 231 160
rect 173 88 185 148
rect 219 88 231 148
rect 173 76 231 88
<< pdiffc >>
rect 97 778 131 838
rect 185 778 219 838
rect 97 640 131 700
rect 185 640 219 700
rect 97 502 131 562
rect 185 502 219 562
rect 97 364 131 424
rect 185 364 219 424
rect 97 226 131 286
rect 185 226 219 286
rect 97 88 131 148
rect 185 88 219 148
<< nsubdiff >>
rect -52 277 31 301
rect -52 242 -28 277
rect 6 242 31 277
rect -52 217 31 242
<< nsubdiffcont >>
rect -28 242 6 277
<< poly >>
rect 125 931 191 947
rect 125 897 141 931
rect 175 897 191 931
rect 125 881 191 897
rect 143 850 173 881
rect 143 712 173 766
rect 143 574 173 628
rect 143 436 173 490
rect 143 298 173 352
rect 143 160 173 214
rect 143 46 173 76
<< polycont >>
rect 141 897 175 931
<< locali >>
rect 125 897 141 931
rect 175 897 191 931
rect 97 838 131 854
rect 97 762 131 778
rect 185 838 219 854
rect 185 762 219 778
rect 97 700 131 716
rect 97 624 131 640
rect 185 700 219 716
rect 185 624 219 640
rect 97 562 131 578
rect 97 486 131 502
rect 185 562 219 578
rect 185 486 219 502
rect 97 424 131 440
rect 97 348 131 364
rect 185 424 219 440
rect 185 348 219 364
rect -52 277 31 301
rect -52 242 -28 277
rect 6 242 31 277
rect -52 217 31 242
rect 97 286 131 302
rect -39 153 18 217
rect 97 210 131 226
rect 185 286 219 302
rect 185 210 219 226
rect 97 153 131 164
rect -39 148 131 153
rect -39 88 97 148
rect -39 82 131 88
rect -39 81 62 82
rect 97 72 131 82
rect 185 148 219 164
rect 185 72 219 88
<< viali >>
rect 141 897 175 931
rect 97 778 131 838
rect 185 778 219 838
rect 97 640 131 700
rect 185 640 219 700
rect 97 502 131 562
rect 185 502 219 562
rect 97 364 131 424
rect 185 364 219 424
rect 97 226 131 286
rect 185 226 219 286
rect 97 88 131 148
rect 185 88 219 148
<< metal1 >>
rect 129 931 187 937
rect 129 897 141 931
rect 175 897 187 931
rect 129 891 187 897
rect 91 838 137 850
rect 91 778 97 838
rect 131 778 137 838
rect 91 766 137 778
rect 179 838 225 850
rect 179 778 185 838
rect 219 778 225 838
rect 91 700 137 712
rect 91 640 97 700
rect 131 640 137 700
rect 91 562 137 640
rect 179 700 225 778
rect 179 640 185 700
rect 219 640 225 700
rect 179 628 225 640
rect 91 502 97 562
rect 131 502 137 562
rect 91 490 137 502
rect 179 562 225 574
rect 179 502 185 562
rect 219 502 225 562
rect 91 424 137 436
rect 91 364 97 424
rect 131 364 137 424
rect 91 286 137 364
rect 179 424 225 502
rect 179 364 185 424
rect 219 364 225 424
rect 179 352 225 364
rect 91 226 97 286
rect 131 226 137 286
rect 91 214 137 226
rect 179 286 225 298
rect 179 226 185 286
rect 219 226 225 286
rect 91 148 137 160
rect 91 88 97 148
rect 131 88 137 148
rect 91 76 137 88
rect 179 148 225 226
rect 179 88 185 148
rect 219 88 225 148
rect 179 76 225 88
<< labels >>
flabel metal1 141 897 175 931 0 FreeSans 320 0 0 0 input_stack
port 0 nsew
flabel nwell 97 88 131 148 0 FreeSans 320 0 0 0 vdd
port 1 nsew
flabel metal1 91 838 137 850 0 FreeSans 320 0 0 0 output_stack
port 6 nsew
<< end >>
