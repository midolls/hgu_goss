magic
tech sky130A
magscale 1 2
timestamp 1698626624
<< pwell >>
rect 1006 4374 1032 4406
rect 1612 4374 1638 4406
rect 686 4046 738 4070
rect 1602 3874 1654 3898
rect 1006 3214 1032 3246
rect 1612 3214 1638 3246
<< metal3 >>
rect 686 5184 1964 5186
rect 686 5120 790 5184
rect 854 5120 870 5184
rect 934 5120 950 5184
rect 1014 5120 1030 5184
rect 1094 5120 1110 5184
rect 1174 5120 1190 5184
rect 1254 5120 1396 5184
rect 1460 5120 1476 5184
rect 1540 5120 1556 5184
rect 1620 5120 1636 5184
rect 1700 5120 1716 5184
rect 1780 5120 1796 5184
rect 1860 5120 1964 5184
rect 686 5118 1964 5120
rect 686 4964 752 5118
rect 686 4900 687 4964
rect 751 4900 752 4964
rect 686 4884 752 4900
rect 686 4820 687 4884
rect 751 4820 752 4884
rect 686 4804 752 4820
rect 686 4740 687 4804
rect 751 4740 752 4804
rect 686 4724 752 4740
rect 686 4660 687 4724
rect 751 4660 752 4724
rect 686 4644 752 4660
rect 686 4580 687 4644
rect 751 4580 752 4644
rect 686 4564 752 4580
rect 686 4500 687 4564
rect 751 4500 752 4564
rect 686 4484 752 4500
rect 686 4420 687 4484
rect 751 4420 752 4484
rect 686 4404 752 4420
rect 686 4340 687 4404
rect 751 4340 752 4404
rect 686 4324 752 4340
rect 686 4260 687 4324
rect 751 4260 752 4324
rect 686 4244 752 4260
rect 686 4180 687 4244
rect 751 4180 752 4244
rect 686 4090 752 4180
rect 812 4086 872 5118
rect 932 4026 992 5056
rect 1052 4086 1112 5118
rect 1172 4026 1232 5056
rect 1292 4964 1358 5118
rect 1292 4900 1293 4964
rect 1357 4900 1358 4964
rect 1292 4884 1358 4900
rect 1292 4820 1293 4884
rect 1357 4820 1358 4884
rect 1292 4804 1358 4820
rect 1292 4740 1293 4804
rect 1357 4740 1358 4804
rect 1292 4724 1358 4740
rect 1292 4660 1293 4724
rect 1357 4660 1358 4724
rect 1292 4644 1358 4660
rect 1292 4580 1293 4644
rect 1357 4580 1358 4644
rect 1292 4564 1358 4580
rect 1292 4500 1293 4564
rect 1357 4500 1358 4564
rect 1292 4484 1358 4500
rect 1292 4420 1293 4484
rect 1357 4420 1358 4484
rect 1292 4404 1358 4420
rect 1292 4340 1293 4404
rect 1357 4340 1358 4404
rect 1292 4324 1358 4340
rect 1292 4260 1293 4324
rect 1357 4260 1358 4324
rect 1292 4244 1358 4260
rect 1292 4180 1293 4244
rect 1357 4180 1358 4244
rect 1292 4090 1358 4180
rect 1418 4086 1478 5118
rect 1538 4026 1598 5056
rect 1658 4086 1718 5118
rect 1778 4026 1838 5056
rect 1898 4964 1964 5118
rect 1898 4900 1899 4964
rect 1963 4900 1964 4964
rect 1898 4884 1964 4900
rect 1898 4820 1899 4884
rect 1963 4820 1964 4884
rect 1898 4804 1964 4820
rect 1898 4740 1899 4804
rect 1963 4740 1964 4804
rect 1898 4724 1964 4740
rect 1898 4660 1899 4724
rect 1963 4660 1964 4724
rect 1898 4644 1964 4660
rect 1898 4580 1899 4644
rect 1963 4580 1964 4644
rect 1898 4564 1964 4580
rect 1898 4500 1899 4564
rect 1963 4500 1964 4564
rect 1898 4484 1964 4500
rect 1898 4420 1899 4484
rect 1963 4420 1964 4484
rect 1898 4404 1964 4420
rect 1898 4340 1899 4404
rect 1963 4340 1964 4404
rect 1898 4324 1964 4340
rect 1898 4260 1899 4324
rect 1963 4260 1964 4324
rect 1898 4244 1964 4260
rect 1898 4180 1899 4244
rect 1963 4180 1964 4244
rect 1898 4090 1964 4180
rect 686 4024 1964 4026
rect 686 3960 790 4024
rect 854 3960 870 4024
rect 934 3960 950 4024
rect 1014 3960 1030 4024
rect 1094 3960 1110 4024
rect 1174 3960 1190 4024
rect 1254 3960 1396 4024
rect 1460 3960 1476 4024
rect 1540 3960 1556 4024
rect 1620 3960 1636 4024
rect 1700 3960 1716 4024
rect 1780 3960 1796 4024
rect 1860 3960 1964 4024
rect 686 3958 1964 3960
rect 686 3804 752 3958
rect 686 3740 687 3804
rect 751 3740 752 3804
rect 686 3724 752 3740
rect 686 3660 687 3724
rect 751 3660 752 3724
rect 686 3644 752 3660
rect 686 3580 687 3644
rect 751 3580 752 3644
rect 686 3564 752 3580
rect 686 3500 687 3564
rect 751 3500 752 3564
rect 686 3484 752 3500
rect 686 3420 687 3484
rect 751 3420 752 3484
rect 686 3404 752 3420
rect 686 3340 687 3404
rect 751 3340 752 3404
rect 686 3324 752 3340
rect 686 3260 687 3324
rect 751 3260 752 3324
rect 686 3244 752 3260
rect 686 3180 687 3244
rect 751 3180 752 3244
rect 686 3164 752 3180
rect 686 3100 687 3164
rect 751 3100 752 3164
rect 686 3084 752 3100
rect 686 3020 687 3084
rect 751 3020 752 3084
rect 686 2930 752 3020
rect 812 2926 872 3958
rect 932 2866 992 3896
rect 1052 2926 1112 3958
rect 1172 2866 1232 3896
rect 1292 3804 1358 3958
rect 1292 3740 1293 3804
rect 1357 3740 1358 3804
rect 1292 3724 1358 3740
rect 1292 3660 1293 3724
rect 1357 3660 1358 3724
rect 1292 3644 1358 3660
rect 1292 3580 1293 3644
rect 1357 3580 1358 3644
rect 1292 3564 1358 3580
rect 1292 3500 1293 3564
rect 1357 3500 1358 3564
rect 1292 3484 1358 3500
rect 1292 3420 1293 3484
rect 1357 3420 1358 3484
rect 1292 3404 1358 3420
rect 1292 3340 1293 3404
rect 1357 3340 1358 3404
rect 1292 3324 1358 3340
rect 1292 3260 1293 3324
rect 1357 3260 1358 3324
rect 1292 3244 1358 3260
rect 1292 3180 1293 3244
rect 1357 3180 1358 3244
rect 1292 3164 1358 3180
rect 1292 3100 1293 3164
rect 1357 3100 1358 3164
rect 1292 3084 1358 3100
rect 1292 3020 1293 3084
rect 1357 3020 1358 3084
rect 1292 2930 1358 3020
rect 1418 2926 1478 3958
rect 1538 2866 1598 3896
rect 1658 2926 1718 3958
rect 1778 2866 1838 3896
rect 1898 3804 1964 3958
rect 1898 3740 1899 3804
rect 1963 3740 1964 3804
rect 1898 3724 1964 3740
rect 1898 3660 1899 3724
rect 1963 3660 1964 3724
rect 1898 3644 1964 3660
rect 1898 3580 1899 3644
rect 1963 3580 1964 3644
rect 1898 3564 1964 3580
rect 1898 3500 1899 3564
rect 1963 3500 1964 3564
rect 1898 3484 1964 3500
rect 1898 3420 1899 3484
rect 1963 3420 1964 3484
rect 1898 3404 1964 3420
rect 1898 3340 1899 3404
rect 1963 3340 1964 3404
rect 1898 3324 1964 3340
rect 1898 3260 1899 3324
rect 1963 3260 1964 3324
rect 1898 3244 1964 3260
rect 1898 3180 1899 3244
rect 1963 3180 1964 3244
rect 1898 3164 1964 3180
rect 1898 3100 1899 3164
rect 1963 3100 1964 3164
rect 1898 3084 1964 3100
rect 1898 3020 1899 3084
rect 1963 3020 1964 3084
rect 1898 2930 1964 3020
rect 686 2864 1964 2866
rect 686 2800 790 2864
rect 854 2800 870 2864
rect 934 2800 950 2864
rect 1014 2800 1030 2864
rect 1094 2800 1110 2864
rect 1174 2800 1190 2864
rect 1254 2800 1396 2864
rect 1460 2800 1476 2864
rect 1540 2800 1556 2864
rect 1620 2800 1636 2864
rect 1700 2800 1716 2864
rect 1780 2800 1796 2864
rect 1860 2800 1964 2864
rect 686 2798 1964 2800
<< via3 >>
rect 790 5120 854 5184
rect 870 5120 934 5184
rect 950 5120 1014 5184
rect 1030 5120 1094 5184
rect 1110 5120 1174 5184
rect 1190 5120 1254 5184
rect 1396 5120 1460 5184
rect 1476 5120 1540 5184
rect 1556 5120 1620 5184
rect 1636 5120 1700 5184
rect 1716 5120 1780 5184
rect 1796 5120 1860 5184
rect 687 4900 751 4964
rect 687 4820 751 4884
rect 687 4740 751 4804
rect 687 4660 751 4724
rect 687 4580 751 4644
rect 687 4500 751 4564
rect 687 4420 751 4484
rect 687 4340 751 4404
rect 687 4260 751 4324
rect 687 4180 751 4244
rect 1293 4900 1357 4964
rect 1293 4820 1357 4884
rect 1293 4740 1357 4804
rect 1293 4660 1357 4724
rect 1293 4580 1357 4644
rect 1293 4500 1357 4564
rect 1293 4420 1357 4484
rect 1293 4340 1357 4404
rect 1293 4260 1357 4324
rect 1293 4180 1357 4244
rect 1899 4900 1963 4964
rect 1899 4820 1963 4884
rect 1899 4740 1963 4804
rect 1899 4660 1963 4724
rect 1899 4580 1963 4644
rect 1899 4500 1963 4564
rect 1899 4420 1963 4484
rect 1899 4340 1963 4404
rect 1899 4260 1963 4324
rect 1899 4180 1963 4244
rect 790 3960 854 4024
rect 870 3960 934 4024
rect 950 3960 1014 4024
rect 1030 3960 1094 4024
rect 1110 3960 1174 4024
rect 1190 3960 1254 4024
rect 1396 3960 1460 4024
rect 1476 3960 1540 4024
rect 1556 3960 1620 4024
rect 1636 3960 1700 4024
rect 1716 3960 1780 4024
rect 1796 3960 1860 4024
rect 687 3740 751 3804
rect 687 3660 751 3724
rect 687 3580 751 3644
rect 687 3500 751 3564
rect 687 3420 751 3484
rect 687 3340 751 3404
rect 687 3260 751 3324
rect 687 3180 751 3244
rect 687 3100 751 3164
rect 687 3020 751 3084
rect 1293 3740 1357 3804
rect 1293 3660 1357 3724
rect 1293 3580 1357 3644
rect 1293 3500 1357 3564
rect 1293 3420 1357 3484
rect 1293 3340 1357 3404
rect 1293 3260 1357 3324
rect 1293 3180 1357 3244
rect 1293 3100 1357 3164
rect 1293 3020 1357 3084
rect 1899 3740 1963 3804
rect 1899 3660 1963 3724
rect 1899 3580 1963 3644
rect 1899 3500 1963 3564
rect 1899 3420 1963 3484
rect 1899 3340 1963 3404
rect 1899 3260 1963 3324
rect 1899 3180 1963 3244
rect 1899 3100 1963 3164
rect 1899 3020 1963 3084
rect 790 2800 854 2864
rect 870 2800 934 2864
rect 950 2800 1014 2864
rect 1030 2800 1094 2864
rect 1110 2800 1174 2864
rect 1190 2800 1254 2864
rect 1396 2800 1460 2864
rect 1476 2800 1540 2864
rect 1556 2800 1620 2864
rect 1636 2800 1700 2864
rect 1716 2800 1780 2864
rect 1796 2800 1860 2864
<< metal4 >>
rect 686 5184 1964 5186
rect 686 5120 790 5184
rect 854 5120 870 5184
rect 934 5120 950 5184
rect 1014 5120 1030 5184
rect 1094 5120 1110 5184
rect 1174 5120 1190 5184
rect 1254 5120 1396 5184
rect 1460 5120 1476 5184
rect 1540 5120 1556 5184
rect 1620 5120 1636 5184
rect 1700 5120 1716 5184
rect 1780 5120 1796 5184
rect 1860 5120 1964 5184
rect 686 5118 1964 5120
rect 686 4964 752 5118
rect 686 4900 687 4964
rect 751 4900 752 4964
rect 686 4884 752 4900
rect 686 4820 687 4884
rect 751 4820 752 4884
rect 686 4804 752 4820
rect 686 4740 687 4804
rect 751 4740 752 4804
rect 686 4724 752 4740
rect 686 4660 687 4724
rect 751 4660 752 4724
rect 686 4644 752 4660
rect 686 4580 687 4644
rect 751 4580 752 4644
rect 686 4564 752 4580
rect 686 4500 687 4564
rect 751 4500 752 4564
rect 686 4484 752 4500
rect 686 4420 687 4484
rect 751 4420 752 4484
rect 686 4404 752 4420
rect 686 4340 687 4404
rect 751 4340 752 4404
rect 686 4324 752 4340
rect 686 4260 687 4324
rect 751 4260 752 4324
rect 686 4244 752 4260
rect 686 4180 687 4244
rect 751 4180 752 4244
rect 686 4090 752 4180
rect 812 4026 872 5056
rect 932 4086 992 5118
rect 1052 4026 1112 5056
rect 1172 4086 1232 5118
rect 1292 4964 1358 5118
rect 1292 4900 1293 4964
rect 1357 4900 1358 4964
rect 1292 4884 1358 4900
rect 1292 4820 1293 4884
rect 1357 4820 1358 4884
rect 1292 4804 1358 4820
rect 1292 4740 1293 4804
rect 1357 4740 1358 4804
rect 1292 4724 1358 4740
rect 1292 4660 1293 4724
rect 1357 4660 1358 4724
rect 1292 4644 1358 4660
rect 1292 4580 1293 4644
rect 1357 4580 1358 4644
rect 1292 4564 1358 4580
rect 1292 4500 1293 4564
rect 1357 4500 1358 4564
rect 1292 4484 1358 4500
rect 1292 4420 1293 4484
rect 1357 4420 1358 4484
rect 1292 4404 1358 4420
rect 1292 4340 1293 4404
rect 1357 4340 1358 4404
rect 1292 4324 1358 4340
rect 1292 4260 1293 4324
rect 1357 4260 1358 4324
rect 1292 4244 1358 4260
rect 1292 4180 1293 4244
rect 1357 4180 1358 4244
rect 1292 4090 1358 4180
rect 1418 4026 1478 5056
rect 1538 4086 1598 5118
rect 1658 4026 1718 5056
rect 1778 4086 1838 5118
rect 1898 4964 1964 5118
rect 1898 4900 1899 4964
rect 1963 4900 1964 4964
rect 1898 4884 1964 4900
rect 1898 4820 1899 4884
rect 1963 4820 1964 4884
rect 1898 4804 1964 4820
rect 1898 4740 1899 4804
rect 1963 4740 1964 4804
rect 1898 4724 1964 4740
rect 1898 4660 1899 4724
rect 1963 4660 1964 4724
rect 1898 4644 1964 4660
rect 1898 4580 1899 4644
rect 1963 4580 1964 4644
rect 1898 4564 1964 4580
rect 1898 4500 1899 4564
rect 1963 4500 1964 4564
rect 1898 4484 1964 4500
rect 1898 4420 1899 4484
rect 1963 4420 1964 4484
rect 1898 4404 1964 4420
rect 1898 4340 1899 4404
rect 1963 4340 1964 4404
rect 1898 4324 1964 4340
rect 1898 4260 1899 4324
rect 1963 4260 1964 4324
rect 1898 4244 1964 4260
rect 1898 4180 1899 4244
rect 1963 4180 1964 4244
rect 1898 4090 1964 4180
rect 686 4024 1964 4026
rect 686 3960 790 4024
rect 854 3960 870 4024
rect 934 3960 950 4024
rect 1014 3960 1030 4024
rect 1094 3960 1110 4024
rect 1174 3960 1190 4024
rect 1254 3960 1396 4024
rect 1460 3960 1476 4024
rect 1540 3960 1556 4024
rect 1620 3960 1636 4024
rect 1700 3960 1716 4024
rect 1780 3960 1796 4024
rect 1860 3960 1964 4024
rect 686 3958 1964 3960
rect 686 3804 752 3958
rect 686 3740 687 3804
rect 751 3740 752 3804
rect 686 3724 752 3740
rect 686 3660 687 3724
rect 751 3660 752 3724
rect 686 3644 752 3660
rect 686 3580 687 3644
rect 751 3580 752 3644
rect 686 3564 752 3580
rect 686 3500 687 3564
rect 751 3500 752 3564
rect 686 3484 752 3500
rect 686 3420 687 3484
rect 751 3420 752 3484
rect 686 3404 752 3420
rect 686 3340 687 3404
rect 751 3340 752 3404
rect 686 3324 752 3340
rect 686 3260 687 3324
rect 751 3260 752 3324
rect 686 3244 752 3260
rect 686 3180 687 3244
rect 751 3180 752 3244
rect 686 3164 752 3180
rect 686 3100 687 3164
rect 751 3100 752 3164
rect 686 3084 752 3100
rect 686 3020 687 3084
rect 751 3020 752 3084
rect 686 2930 752 3020
rect 812 2866 872 3896
rect 932 2926 992 3958
rect 1052 2866 1112 3896
rect 1172 2926 1232 3958
rect 1292 3804 1358 3958
rect 1292 3740 1293 3804
rect 1357 3740 1358 3804
rect 1292 3724 1358 3740
rect 1292 3660 1293 3724
rect 1357 3660 1358 3724
rect 1292 3644 1358 3660
rect 1292 3580 1293 3644
rect 1357 3580 1358 3644
rect 1292 3564 1358 3580
rect 1292 3500 1293 3564
rect 1357 3500 1358 3564
rect 1292 3484 1358 3500
rect 1292 3420 1293 3484
rect 1357 3420 1358 3484
rect 1292 3404 1358 3420
rect 1292 3340 1293 3404
rect 1357 3340 1358 3404
rect 1292 3324 1358 3340
rect 1292 3260 1293 3324
rect 1357 3260 1358 3324
rect 1292 3244 1358 3260
rect 1292 3180 1293 3244
rect 1357 3180 1358 3244
rect 1292 3164 1358 3180
rect 1292 3100 1293 3164
rect 1357 3100 1358 3164
rect 1292 3084 1358 3100
rect 1292 3020 1293 3084
rect 1357 3020 1358 3084
rect 1292 2930 1358 3020
rect 1418 2866 1478 3896
rect 1538 2926 1598 3958
rect 1658 2866 1718 3896
rect 1778 2926 1838 3958
rect 1898 3804 1964 3958
rect 1898 3740 1899 3804
rect 1963 3740 1964 3804
rect 1898 3724 1964 3740
rect 1898 3660 1899 3724
rect 1963 3660 1964 3724
rect 1898 3644 1964 3660
rect 1898 3580 1899 3644
rect 1963 3580 1964 3644
rect 1898 3564 1964 3580
rect 1898 3500 1899 3564
rect 1963 3500 1964 3564
rect 1898 3484 1964 3500
rect 1898 3420 1899 3484
rect 1963 3420 1964 3484
rect 1898 3404 1964 3420
rect 1898 3340 1899 3404
rect 1963 3340 1964 3404
rect 1898 3324 1964 3340
rect 1898 3260 1899 3324
rect 1963 3260 1964 3324
rect 1898 3244 1964 3260
rect 1898 3180 1899 3244
rect 1963 3180 1964 3244
rect 1898 3164 1964 3180
rect 1898 3100 1899 3164
rect 1963 3100 1964 3164
rect 1898 3084 1964 3100
rect 1898 3020 1899 3084
rect 1963 3020 1964 3084
rect 1898 2930 1964 3020
rect 686 2864 1964 2866
rect 686 2800 790 2864
rect 854 2800 870 2864
rect 934 2800 950 2864
rect 1014 2800 1030 2864
rect 1094 2800 1110 2864
rect 1174 2800 1190 2864
rect 1254 2800 1396 2864
rect 1460 2800 1476 2864
rect 1540 2800 1556 2864
rect 1620 2800 1636 2864
rect 1700 2800 1716 2864
rect 1780 2800 1796 2864
rect 1860 2800 1964 2864
rect 686 2798 1964 2800
<< labels >>
flabel pwell 686 4046 738 4070 0 FreeSans 160 0 0 0 SUB
port 1 nsew
flabel pwell 1612 4374 1638 4406 0 FreeSans 160 0 0 0 x1[3].SUB
flabel metal4 1554 4708 1580 4740 0 FreeSans 320 0 0 0 x1[3].CBOT
flabel metal4 1672 4118 1698 4150 0 FreeSans 320 0 0 0 x1[3].CTOP
flabel pwell 1612 3214 1638 3246 0 FreeSans 160 0 0 0 x1[2].SUB
flabel metal4 1554 3548 1580 3580 0 FreeSans 320 0 0 0 x1[2].CBOT
flabel metal4 1672 2958 1698 2990 0 FreeSans 320 0 0 0 x1[2].CTOP
flabel pwell 1006 4374 1032 4406 0 FreeSans 160 0 0 0 x1[1].SUB
flabel metal4 948 4708 974 4740 0 FreeSans 320 0 0 0 x1[1].CBOT
flabel metal4 1066 4118 1092 4150 0 FreeSans 320 0 0 0 x1[1].CTOP
flabel pwell 1006 3214 1032 3246 0 FreeSans 160 0 0 0 x1[0].SUB
flabel metal4 948 3548 974 3580 0 FreeSans 320 0 0 0 x1[0].CBOT
flabel metal4 1066 2958 1092 2990 0 FreeSans 320 0 0 0 x1[0].CTOP
flabel pwell 1602 3874 1654 3898 0 FreeSans 160 0 0 0 SUB
port 1 nsew
<< end >>
