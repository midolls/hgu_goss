magic
tech sky130A
magscale 1 2
timestamp 1699352056
<< nwell >>
rect -270 -833 1830 -767
rect -233 -834 1830 -833
rect -233 -902 1795 -834
rect -5 -2078 29 -2072
rect 88 -2078 122 -2072
rect 177 -2078 211 -2072
rect 269 -2078 303 -2071
rect 360 -2078 394 -2072
rect 453 -2078 487 -2071
rect 545 -2078 579 -2071
rect 639 -2078 673 -2072
rect 718 -2078 752 -2072
rect 809 -2078 843 -2071
rect 901 -2078 935 -2072
rect 993 -2078 1027 -2072
rect 1085 -2078 1119 -2072
rect 1176 -2078 1210 -2072
rect 1269 -2078 1303 -2072
rect 1362 -2078 1396 -2072
rect 1454 -2078 1488 -2072
rect 1545 -2078 1579 -2072
rect 1637 -2078 1671 -2071
rect 1724 -2078 1758 -2071
rect 1780 -2078 1830 -1830
rect -178 -2143 1830 -2078
rect -178 -2420 1795 -2143
<< psubdiff >>
rect -118 -1463 -89 -1429
rect -55 -1430 85 -1429
rect -55 -1463 -5 -1430
rect -118 -1464 -5 -1463
rect 29 -1463 85 -1430
rect 119 -1463 177 -1429
rect 211 -1430 545 -1429
rect 211 -1463 267 -1430
rect 29 -1464 267 -1463
rect 301 -1464 361 -1430
rect 395 -1464 452 -1430
rect 486 -1463 545 -1430
rect 579 -1430 1453 -1429
rect 579 -1463 636 -1430
rect 486 -1464 636 -1463
rect 670 -1464 716 -1430
rect 750 -1464 809 -1430
rect 843 -1464 901 -1430
rect 935 -1464 994 -1430
rect 1028 -1464 1085 -1430
rect 1119 -1464 1177 -1430
rect 1211 -1464 1270 -1430
rect 1304 -1464 1361 -1430
rect 1395 -1463 1453 -1430
rect 1487 -1430 1790 -1429
rect 1487 -1463 1545 -1430
rect 1395 -1464 1545 -1463
rect 1579 -1464 1640 -1430
rect 1674 -1464 1728 -1430
rect 1762 -1464 1790 -1430
rect -133 -2698 -19 -2697
rect -133 -2732 -109 -2698
rect -75 -2731 -19 -2698
rect 15 -2731 73 -2697
rect 107 -2731 165 -2697
rect 199 -2731 257 -2697
rect 291 -2731 349 -2697
rect 383 -2731 441 -2697
rect 475 -2731 533 -2697
rect 567 -2731 625 -2697
rect 659 -2731 717 -2697
rect 751 -2731 809 -2697
rect 843 -2731 901 -2697
rect 935 -2731 993 -2697
rect 1027 -2731 1085 -2697
rect 1119 -2731 1177 -2697
rect 1211 -2698 1361 -2697
rect 1211 -2731 1269 -2698
rect -75 -2732 1269 -2731
rect 1303 -2731 1361 -2698
rect 1395 -2731 1453 -2697
rect 1487 -2731 1545 -2697
rect 1579 -2731 1637 -2697
rect 1671 -2731 1717 -2697
rect 1751 -2731 1775 -2697
rect 1303 -2732 1775 -2731
<< nsubdiff >>
rect -151 -805 1757 -804
rect -151 -839 -111 -805
rect -77 -839 -19 -805
rect 15 -839 73 -805
rect 107 -839 165 -805
rect 199 -839 257 -805
rect 291 -839 349 -805
rect 383 -839 441 -805
rect 475 -839 533 -805
rect 567 -839 625 -805
rect 659 -839 717 -805
rect 751 -839 809 -805
rect 843 -839 901 -805
rect 935 -839 993 -805
rect 1027 -839 1085 -805
rect 1119 -839 1177 -805
rect 1211 -839 1269 -805
rect 1303 -839 1361 -805
rect 1395 -839 1453 -805
rect 1487 -839 1545 -805
rect 1579 -839 1637 -805
rect 1671 -839 1757 -805
rect -125 -2105 -101 -2071
rect -67 -2072 269 -2071
rect -67 -2105 -5 -2072
rect -125 -2106 -5 -2105
rect 29 -2106 88 -2072
rect 122 -2106 177 -2072
rect 211 -2105 269 -2072
rect 303 -2072 453 -2071
rect 303 -2105 360 -2072
rect 211 -2106 360 -2105
rect 394 -2105 453 -2072
rect 487 -2105 545 -2071
rect 579 -2072 809 -2071
rect 579 -2105 639 -2072
rect 394 -2106 639 -2105
rect 673 -2106 718 -2072
rect 752 -2105 809 -2072
rect 843 -2072 1637 -2071
rect 843 -2105 901 -2072
rect 752 -2106 901 -2105
rect 935 -2106 993 -2072
rect 1027 -2106 1085 -2072
rect 1119 -2106 1176 -2072
rect 1210 -2106 1269 -2072
rect 1303 -2106 1362 -2072
rect 1396 -2106 1454 -2072
rect 1488 -2106 1545 -2072
rect 1579 -2105 1637 -2072
rect 1671 -2105 1724 -2071
rect 1758 -2105 1783 -2071
rect 1579 -2106 1783 -2105
<< psubdiffcont >>
rect -89 -1463 -55 -1429
rect -5 -1464 29 -1430
rect 85 -1463 119 -1429
rect 177 -1463 211 -1429
rect 267 -1464 301 -1430
rect 361 -1464 395 -1430
rect 452 -1464 486 -1430
rect 545 -1463 579 -1429
rect 636 -1464 670 -1430
rect 716 -1464 750 -1430
rect 809 -1464 843 -1430
rect 901 -1464 935 -1430
rect 994 -1464 1028 -1430
rect 1085 -1464 1119 -1430
rect 1177 -1464 1211 -1430
rect 1270 -1464 1304 -1430
rect 1361 -1464 1395 -1430
rect 1453 -1463 1487 -1429
rect 1545 -1464 1579 -1430
rect 1640 -1464 1674 -1430
rect 1728 -1464 1762 -1430
rect -109 -2732 -75 -2698
rect -19 -2731 15 -2697
rect 73 -2731 107 -2697
rect 165 -2731 199 -2697
rect 257 -2731 291 -2697
rect 349 -2731 383 -2697
rect 441 -2731 475 -2697
rect 533 -2731 567 -2697
rect 625 -2731 659 -2697
rect 717 -2731 751 -2697
rect 809 -2731 843 -2697
rect 901 -2731 935 -2697
rect 993 -2731 1027 -2697
rect 1085 -2731 1119 -2697
rect 1177 -2731 1211 -2697
rect 1269 -2732 1303 -2698
rect 1361 -2731 1395 -2697
rect 1453 -2731 1487 -2697
rect 1545 -2731 1579 -2697
rect 1637 -2731 1671 -2697
rect 1717 -2731 1751 -2697
<< nsubdiffcont >>
rect -111 -839 -77 -805
rect -19 -839 15 -805
rect 73 -839 107 -805
rect 165 -839 199 -805
rect 257 -839 291 -805
rect 349 -839 383 -805
rect 441 -839 475 -805
rect 533 -839 567 -805
rect 625 -839 659 -805
rect 717 -839 751 -805
rect 809 -839 843 -805
rect 901 -839 935 -805
rect 993 -839 1027 -805
rect 1085 -839 1119 -805
rect 1177 -839 1211 -805
rect 1269 -839 1303 -805
rect 1361 -839 1395 -805
rect 1453 -839 1487 -805
rect 1545 -839 1579 -805
rect 1637 -839 1671 -805
rect -101 -2105 -67 -2071
rect -5 -2106 29 -2072
rect 88 -2106 122 -2072
rect 177 -2106 211 -2072
rect 269 -2105 303 -2071
rect 360 -2106 394 -2072
rect 453 -2105 487 -2071
rect 545 -2105 579 -2071
rect 639 -2106 673 -2072
rect 718 -2106 752 -2072
rect 809 -2105 843 -2071
rect 901 -2106 935 -2072
rect 993 -2106 1027 -2072
rect 1085 -2106 1119 -2072
rect 1176 -2106 1210 -2072
rect 1269 -2106 1303 -2072
rect 1362 -2106 1396 -2072
rect 1454 -2106 1488 -2072
rect 1545 -2106 1579 -2072
rect 1637 -2105 1671 -2071
rect 1724 -2105 1758 -2071
<< locali >>
rect -232 -805 1792 -804
rect -232 -839 -111 -805
rect -77 -839 -19 -805
rect 15 -839 73 -805
rect 107 -839 165 -805
rect 199 -839 257 -805
rect 291 -839 349 -805
rect 383 -839 441 -805
rect 475 -839 533 -805
rect 567 -839 625 -805
rect 659 -839 717 -805
rect 751 -839 809 -805
rect 843 -839 901 -805
rect 935 -839 993 -805
rect 1027 -839 1085 -805
rect 1119 -839 1177 -805
rect 1211 -839 1269 -805
rect 1303 -839 1361 -805
rect 1395 -839 1453 -805
rect 1487 -839 1545 -805
rect 1579 -839 1637 -805
rect 1671 -839 1792 -805
rect -232 -841 1792 -839
rect -128 -1429 1792 -1400
rect -128 -1463 -89 -1429
rect -55 -1430 85 -1429
rect -55 -1463 -5 -1430
rect -128 -1464 -5 -1463
rect 29 -1463 85 -1430
rect 119 -1463 177 -1429
rect 211 -1430 545 -1429
rect 211 -1463 267 -1430
rect 29 -1464 267 -1463
rect 301 -1464 361 -1430
rect 395 -1464 452 -1430
rect 486 -1463 545 -1430
rect 579 -1430 1453 -1429
rect 579 -1463 636 -1430
rect 486 -1464 636 -1463
rect 670 -1464 716 -1430
rect 750 -1464 809 -1430
rect 843 -1464 901 -1430
rect 935 -1464 994 -1430
rect 1028 -1464 1085 -1430
rect 1119 -1464 1177 -1430
rect 1211 -1464 1270 -1430
rect 1304 -1464 1361 -1430
rect 1395 -1463 1453 -1430
rect 1487 -1430 1792 -1429
rect 1487 -1463 1545 -1430
rect 1395 -1464 1545 -1463
rect 1579 -1464 1640 -1430
rect 1674 -1464 1728 -1430
rect 1762 -1464 1792 -1430
rect -128 -1485 1792 -1464
rect -128 -2071 1792 -2056
rect -128 -2105 -101 -2071
rect -67 -2072 269 -2071
rect -67 -2105 -5 -2072
rect -128 -2106 -5 -2105
rect 29 -2106 88 -2072
rect 122 -2106 177 -2072
rect 211 -2105 269 -2072
rect 303 -2072 453 -2071
rect 303 -2105 360 -2072
rect 211 -2106 360 -2105
rect 394 -2105 453 -2072
rect 487 -2105 545 -2071
rect 579 -2072 809 -2071
rect 579 -2105 639 -2072
rect 394 -2106 639 -2105
rect 673 -2106 718 -2072
rect 752 -2105 809 -2072
rect 843 -2072 1637 -2071
rect 843 -2105 901 -2072
rect 752 -2106 901 -2105
rect 935 -2106 993 -2072
rect 1027 -2106 1085 -2072
rect 1119 -2106 1176 -2072
rect 1210 -2106 1269 -2072
rect 1303 -2106 1362 -2072
rect 1396 -2106 1454 -2072
rect 1488 -2106 1545 -2072
rect 1579 -2105 1637 -2072
rect 1671 -2105 1724 -2071
rect 1758 -2105 1792 -2071
rect 1579 -2106 1792 -2105
rect -128 -2125 1792 -2106
rect -140 -2698 -19 -2697
rect -140 -2732 -109 -2698
rect -75 -2731 -19 -2698
rect 15 -2731 73 -2697
rect 107 -2731 165 -2697
rect 199 -2731 257 -2697
rect 291 -2731 349 -2697
rect 383 -2731 441 -2697
rect 475 -2731 533 -2697
rect 567 -2731 625 -2697
rect 659 -2731 717 -2697
rect 751 -2731 809 -2697
rect 843 -2731 901 -2697
rect 935 -2731 993 -2697
rect 1027 -2731 1085 -2697
rect 1119 -2731 1177 -2697
rect 1211 -2698 1361 -2697
rect 1211 -2731 1269 -2698
rect -75 -2732 1269 -2731
rect 1303 -2731 1361 -2698
rect 1395 -2731 1453 -2697
rect 1487 -2731 1545 -2697
rect 1579 -2731 1637 -2697
rect 1671 -2731 1717 -2697
rect 1751 -2731 1792 -2697
rect 1303 -2732 1792 -2731
rect -140 -2733 1792 -2732
<< viali >>
rect -200 -1176 -166 -1142
rect 1419 -1183 1453 -1149
rect -97 -1745 -63 -1711
rect 302 -1748 336 -1714
rect 632 -1752 666 -1718
rect 872 -1754 906 -1720
rect 1160 -1757 1194 -1723
rect 1425 -1747 1459 -1713
rect 1712 -1754 1746 -1720
rect 86 -1969 120 -1935
rect 716 -2241 750 -2207
rect 1268 -2241 1302 -2207
rect 78 -2310 112 -2276
rect 353 -2307 387 -2273
rect 627 -2307 661 -2273
rect 1185 -2304 1219 -2270
rect 1733 -2306 1767 -2272
rect -110 -2467 -76 -2433
rect 166 -2467 200 -2433
rect 442 -2467 476 -2433
rect 899 -2465 933 -2431
rect 994 -2465 1028 -2431
rect 1451 -2465 1485 -2431
rect 1547 -2465 1581 -2431
<< metal1 >>
rect -19 -839 15 -805
rect 73 -839 107 -805
rect 165 -839 199 -805
rect 257 -839 291 -805
rect 349 -839 383 -805
rect 441 -839 475 -805
rect 533 -839 567 -805
rect 625 -839 659 -805
rect 717 -839 751 -805
rect 809 -839 843 -805
rect 901 -839 935 -805
rect 993 -829 1027 -805
rect 967 -881 974 -829
rect 1026 -881 1032 -829
rect 1085 -839 1119 -805
rect 1177 -828 1211 -805
rect 1168 -880 1175 -828
rect 1227 -880 1233 -828
rect 1269 -839 1303 -805
rect 1361 -825 1395 -805
rect 1361 -839 1375 -825
rect 1368 -877 1375 -839
rect 1427 -877 1433 -825
rect 1453 -839 1487 -805
rect 1545 -839 1579 -805
rect 1637 -826 1671 -805
rect 1368 -878 1433 -877
rect 1592 -878 1599 -826
rect 1651 -839 1671 -826
rect 1651 -878 1657 -839
rect 1592 -879 1657 -878
rect 1168 -881 1233 -880
rect 967 -882 1032 -881
rect -209 -1133 -157 -1127
rect -209 -1191 -157 -1185
rect 1410 -1140 1462 -1134
rect 1410 -1198 1462 -1192
rect -68 -1474 -61 -1422
rect -9 -1430 -3 -1422
rect -9 -1464 29 -1430
rect 85 -1463 119 -1429
rect 177 -1463 211 -1429
rect 267 -1464 301 -1430
rect 361 -1464 395 -1430
rect -9 -1474 -3 -1464
rect 425 -1471 432 -1419
rect 484 -1471 490 -1419
rect 545 -1463 579 -1429
rect 425 -1472 490 -1471
rect 611 -1472 618 -1420
rect 670 -1472 676 -1420
rect 716 -1464 750 -1430
rect 809 -1464 843 -1430
rect 901 -1464 935 -1430
rect 994 -1464 1028 -1430
rect 1085 -1464 1119 -1430
rect 1177 -1464 1211 -1430
rect 1270 -1464 1304 -1430
rect 1361 -1464 1395 -1430
rect 1453 -1463 1487 -1429
rect 1545 -1464 1579 -1430
rect 1640 -1464 1674 -1430
rect 1728 -1464 1762 -1430
rect 611 -1473 676 -1472
rect -68 -1475 -3 -1474
rect -108 -1711 -51 -1521
rect -108 -1745 -97 -1711
rect -63 -1745 -51 -1711
rect -108 -1757 -51 -1745
rect 201 -1705 253 -1699
rect 295 -1709 349 -1706
rect 253 -1714 349 -1709
rect 253 -1748 302 -1714
rect 336 -1748 349 -1714
rect 253 -1752 349 -1748
rect 295 -1755 349 -1752
rect 623 -1709 675 -1703
rect 1416 -1704 1468 -1698
rect 201 -1763 253 -1757
rect 623 -1767 675 -1761
rect 863 -1711 915 -1705
rect 863 -1769 915 -1763
rect 1151 -1714 1203 -1708
rect 1416 -1762 1468 -1756
rect 1703 -1711 1755 -1705
rect 1151 -1772 1203 -1766
rect 1703 -1769 1755 -1763
rect 79 -1935 128 -1922
rect 79 -1969 86 -1935
rect 120 -1969 128 -1935
rect 79 -2008 128 -1969
rect -5 -2106 29 -2072
rect 88 -2106 122 -2072
rect 177 -2106 211 -2072
rect 269 -2105 303 -2071
rect 360 -2106 394 -2072
rect 453 -2105 487 -2071
rect 545 -2105 579 -2071
rect 639 -2106 673 -2072
rect 718 -2106 752 -2072
rect 809 -2105 843 -2071
rect 872 -2114 879 -2062
rect 931 -2114 937 -2062
rect 993 -2106 1027 -2072
rect 1057 -2113 1064 -2061
rect 1116 -2113 1122 -2061
rect 1176 -2106 1210 -2072
rect 1057 -2114 1122 -2113
rect 1247 -2113 1254 -2061
rect 1306 -2113 1312 -2061
rect 1431 -2072 1438 -2062
rect 1362 -2106 1438 -2072
rect 1247 -2114 1312 -2113
rect 1431 -2114 1438 -2106
rect 1490 -2114 1496 -2062
rect 1545 -2106 1579 -2072
rect 872 -2115 937 -2114
rect 1431 -2115 1496 -2114
rect 1615 -2117 1622 -2065
rect 1674 -2117 1680 -2065
rect 1724 -2105 1758 -2071
rect 1615 -2118 1680 -2117
rect 708 -2207 757 -2168
rect 708 -2241 716 -2207
rect 750 -2241 757 -2207
rect 708 -2254 757 -2241
rect 1260 -2207 1309 -2168
rect 1260 -2241 1268 -2207
rect 1302 -2241 1309 -2207
rect 1260 -2254 1309 -2241
rect 69 -2267 121 -2261
rect 69 -2325 121 -2319
rect 344 -2264 396 -2258
rect 344 -2322 396 -2316
rect 618 -2264 670 -2258
rect 618 -2322 670 -2316
rect 1176 -2261 1228 -2255
rect 1176 -2319 1228 -2313
rect 1724 -2263 1776 -2257
rect 1724 -2321 1776 -2315
rect -119 -2424 -67 -2418
rect -119 -2482 -67 -2476
rect 157 -2424 209 -2418
rect 157 -2482 209 -2476
rect 433 -2424 485 -2418
rect 433 -2482 485 -2476
rect 887 -2431 944 -2419
rect 887 -2465 899 -2431
rect 933 -2465 944 -2431
rect 4 -2697 11 -2654
rect -19 -2706 11 -2697
rect 63 -2706 69 -2654
rect 887 -2655 944 -2465
rect 985 -2422 1037 -2416
rect 985 -2480 1037 -2474
rect 1439 -2431 1496 -2419
rect 1439 -2465 1451 -2431
rect 1485 -2465 1496 -2431
rect 1439 -2655 1496 -2465
rect 1538 -2422 1590 -2416
rect 1538 -2480 1590 -2474
rect 263 -2697 270 -2658
rect -19 -2707 69 -2706
rect -19 -2731 15 -2707
rect 73 -2731 107 -2697
rect 165 -2731 199 -2697
rect 257 -2710 270 -2697
rect 322 -2710 328 -2658
rect 257 -2711 328 -2710
rect 257 -2731 291 -2711
rect 349 -2731 383 -2697
rect 441 -2731 475 -2697
rect 533 -2731 567 -2697
rect 568 -2710 575 -2658
rect 627 -2710 633 -2658
rect 568 -2711 633 -2710
rect 625 -2731 659 -2711
rect 717 -2731 751 -2697
rect 809 -2731 843 -2697
rect 901 -2731 935 -2697
rect 993 -2731 1027 -2697
rect 1085 -2731 1119 -2697
rect 1177 -2731 1211 -2697
rect 1269 -2732 1303 -2698
rect 1361 -2731 1395 -2697
rect 1453 -2731 1487 -2697
rect 1545 -2731 1579 -2697
rect 1637 -2731 1671 -2697
rect 1716 -2731 1750 -2697
<< via1 >>
rect 974 -881 1026 -829
rect 1175 -880 1227 -828
rect 1375 -877 1427 -825
rect 1599 -878 1651 -826
rect -209 -1142 -157 -1133
rect -209 -1176 -200 -1142
rect -200 -1176 -166 -1142
rect -166 -1176 -157 -1142
rect -209 -1185 -157 -1176
rect 1410 -1149 1462 -1140
rect 1410 -1183 1419 -1149
rect 1419 -1183 1453 -1149
rect 1453 -1183 1462 -1149
rect 1410 -1192 1462 -1183
rect -61 -1474 -9 -1422
rect 432 -1471 484 -1419
rect 618 -1472 670 -1420
rect 201 -1757 253 -1705
rect 623 -1718 675 -1709
rect 623 -1752 632 -1718
rect 632 -1752 666 -1718
rect 666 -1752 675 -1718
rect 623 -1761 675 -1752
rect 863 -1720 915 -1711
rect 863 -1754 872 -1720
rect 872 -1754 906 -1720
rect 906 -1754 915 -1720
rect 863 -1763 915 -1754
rect 1151 -1723 1203 -1714
rect 1151 -1757 1160 -1723
rect 1160 -1757 1194 -1723
rect 1194 -1757 1203 -1723
rect 1151 -1766 1203 -1757
rect 1416 -1713 1468 -1704
rect 1416 -1747 1425 -1713
rect 1425 -1747 1459 -1713
rect 1459 -1747 1468 -1713
rect 1416 -1756 1468 -1747
rect 1703 -1720 1755 -1711
rect 1703 -1754 1712 -1720
rect 1712 -1754 1746 -1720
rect 1746 -1754 1755 -1720
rect 1703 -1763 1755 -1754
rect 879 -2114 931 -2062
rect 1064 -2113 1116 -2061
rect 1254 -2113 1306 -2061
rect 1438 -2114 1490 -2062
rect 1622 -2117 1674 -2065
rect 69 -2276 121 -2267
rect 69 -2310 78 -2276
rect 78 -2310 112 -2276
rect 112 -2310 121 -2276
rect 69 -2319 121 -2310
rect 344 -2273 396 -2264
rect 344 -2307 353 -2273
rect 353 -2307 387 -2273
rect 387 -2307 396 -2273
rect 344 -2316 396 -2307
rect 618 -2273 670 -2264
rect 618 -2307 627 -2273
rect 627 -2307 661 -2273
rect 661 -2307 670 -2273
rect 618 -2316 670 -2307
rect 1176 -2270 1228 -2261
rect 1176 -2304 1185 -2270
rect 1185 -2304 1219 -2270
rect 1219 -2304 1228 -2270
rect 1176 -2313 1228 -2304
rect 1724 -2272 1776 -2263
rect 1724 -2306 1733 -2272
rect 1733 -2306 1767 -2272
rect 1767 -2306 1776 -2272
rect 1724 -2315 1776 -2306
rect -119 -2433 -67 -2424
rect -119 -2467 -110 -2433
rect -110 -2467 -76 -2433
rect -76 -2467 -67 -2433
rect -119 -2476 -67 -2467
rect 157 -2433 209 -2424
rect 157 -2467 166 -2433
rect 166 -2467 200 -2433
rect 200 -2467 209 -2433
rect 157 -2476 209 -2467
rect 433 -2433 485 -2424
rect 433 -2467 442 -2433
rect 442 -2467 476 -2433
rect 476 -2467 485 -2433
rect 433 -2476 485 -2467
rect 11 -2706 63 -2654
rect 985 -2431 1037 -2422
rect 985 -2465 994 -2431
rect 994 -2465 1028 -2431
rect 1028 -2465 1037 -2431
rect 985 -2474 1037 -2465
rect 1538 -2431 1590 -2422
rect 1538 -2465 1547 -2431
rect 1547 -2465 1581 -2431
rect 1581 -2465 1590 -2431
rect 1538 -2474 1590 -2465
rect 270 -2710 322 -2658
rect 575 -2710 627 -2658
<< metal2 >>
rect -204 -1127 -163 -714
rect -209 -1133 -157 -1127
rect -209 -1191 -157 -1185
rect -72 -1476 -63 -1420
rect -7 -1476 2 -1420
rect 74 -2261 115 -714
rect 206 -1699 247 -714
rect 201 -1705 253 -1699
rect 201 -1763 253 -1757
rect 350 -2258 391 -714
rect 421 -1473 430 -1417
rect 486 -1473 495 -1417
rect 607 -1474 616 -1418
rect 672 -1474 681 -1418
rect 623 -1709 675 -1703
rect 869 -1705 910 -714
rect 963 -883 972 -827
rect 1028 -883 1037 -827
rect 1164 -882 1173 -826
rect 1229 -882 1238 -826
rect 1364 -879 1373 -823
rect 1429 -879 1438 -823
rect 1588 -880 1597 -824
rect 1653 -880 1662 -824
rect 1410 -1140 1462 -1134
rect 1462 -1192 1466 -1170
rect 1410 -1198 1466 -1192
rect 1416 -1698 1466 -1198
rect 1416 -1704 1468 -1698
rect 621 -1761 623 -1730
rect 621 -1767 675 -1761
rect 863 -1711 915 -1705
rect 621 -2258 671 -1767
rect 863 -1769 915 -1763
rect 1151 -1714 1203 -1708
rect 1203 -1766 1215 -1735
rect 1416 -1762 1468 -1756
rect 1703 -1711 1755 -1705
rect 1151 -1772 1215 -1766
rect 1755 -1763 1765 -1736
rect 1703 -1769 1765 -1763
rect 868 -2116 877 -2060
rect 933 -2116 942 -2060
rect 1053 -2115 1062 -2059
rect 1118 -2115 1127 -2059
rect 69 -2267 121 -2261
rect 69 -2325 121 -2319
rect 344 -2264 396 -2258
rect 344 -2322 396 -2316
rect 618 -2264 671 -2258
rect 670 -2298 671 -2264
rect 1165 -2255 1215 -1772
rect 1243 -2115 1252 -2059
rect 1308 -2115 1317 -2059
rect 1427 -2116 1436 -2060
rect 1492 -2116 1501 -2060
rect 1611 -2119 1620 -2063
rect 1676 -2119 1685 -2063
rect 1165 -2261 1228 -2255
rect 1165 -2303 1176 -2261
rect 618 -2322 670 -2316
rect 1715 -2257 1765 -1769
rect 1715 -2263 1776 -2257
rect 1715 -2304 1724 -2263
rect 1176 -2319 1228 -2313
rect 1724 -2321 1776 -2315
rect -119 -2424 -67 -2418
rect -119 -2482 -67 -2476
rect 157 -2424 209 -2418
rect 157 -2482 209 -2476
rect 433 -2424 485 -2418
rect 433 -2482 485 -2476
rect 985 -2422 1037 -2416
rect 985 -2480 1037 -2474
rect 1538 -2422 1590 -2416
rect 1538 -2480 1590 -2474
rect -106 -2798 -78 -2482
rect 0 -2708 9 -2652
rect 65 -2708 74 -2652
rect 171 -2798 199 -2482
rect 259 -2712 268 -2656
rect 324 -2712 333 -2656
rect 446 -2793 474 -2482
rect 564 -2712 573 -2656
rect 629 -2712 638 -2656
rect 991 -2788 1019 -2480
rect 1550 -2793 1578 -2480
<< via2 >>
rect -63 -1422 -7 -1420
rect -63 -1474 -61 -1422
rect -61 -1474 -9 -1422
rect -9 -1474 -7 -1422
rect -63 -1476 -7 -1474
rect 430 -1419 486 -1417
rect 430 -1471 432 -1419
rect 432 -1471 484 -1419
rect 484 -1471 486 -1419
rect 430 -1473 486 -1471
rect 616 -1420 672 -1418
rect 616 -1472 618 -1420
rect 618 -1472 670 -1420
rect 670 -1472 672 -1420
rect 616 -1474 672 -1472
rect 972 -829 1028 -827
rect 972 -881 974 -829
rect 974 -881 1026 -829
rect 1026 -881 1028 -829
rect 972 -883 1028 -881
rect 1173 -828 1229 -826
rect 1173 -880 1175 -828
rect 1175 -880 1227 -828
rect 1227 -880 1229 -828
rect 1173 -882 1229 -880
rect 1373 -825 1429 -823
rect 1373 -877 1375 -825
rect 1375 -877 1427 -825
rect 1427 -877 1429 -825
rect 1373 -879 1429 -877
rect 1597 -826 1653 -824
rect 1597 -878 1599 -826
rect 1599 -878 1651 -826
rect 1651 -878 1653 -826
rect 1597 -880 1653 -878
rect 877 -2062 933 -2060
rect 877 -2114 879 -2062
rect 879 -2114 931 -2062
rect 931 -2114 933 -2062
rect 877 -2116 933 -2114
rect 1062 -2061 1118 -2059
rect 1062 -2113 1064 -2061
rect 1064 -2113 1116 -2061
rect 1116 -2113 1118 -2061
rect 1062 -2115 1118 -2113
rect 1252 -2061 1308 -2059
rect 1252 -2113 1254 -2061
rect 1254 -2113 1306 -2061
rect 1306 -2113 1308 -2061
rect 1252 -2115 1308 -2113
rect 1436 -2062 1492 -2060
rect 1436 -2114 1438 -2062
rect 1438 -2114 1490 -2062
rect 1490 -2114 1492 -2062
rect 1436 -2116 1492 -2114
rect 1620 -2065 1676 -2063
rect 1620 -2117 1622 -2065
rect 1622 -2117 1674 -2065
rect 1674 -2117 1676 -2065
rect 1620 -2119 1676 -2117
rect 9 -2654 65 -2652
rect 9 -2706 11 -2654
rect 11 -2706 63 -2654
rect 63 -2706 65 -2654
rect 9 -2708 65 -2706
rect 268 -2658 324 -2656
rect 268 -2710 270 -2658
rect 270 -2710 322 -2658
rect 322 -2710 324 -2658
rect 268 -2712 324 -2710
rect 573 -2658 629 -2656
rect 573 -2710 575 -2658
rect 575 -2710 627 -2658
rect 627 -2710 629 -2658
rect 573 -2712 629 -2710
<< metal3 >>
rect 942 -824 1066 -818
rect 942 -888 968 -824
rect 1032 -888 1066 -824
rect 942 -896 1066 -888
rect 1143 -823 1267 -817
rect 1143 -887 1169 -823
rect 1233 -887 1267 -823
rect 1143 -895 1267 -887
rect 1343 -820 1467 -814
rect 1343 -884 1369 -820
rect 1433 -884 1467 -820
rect 1343 -892 1467 -884
rect 1567 -821 1691 -815
rect 1567 -885 1593 -821
rect 1657 -885 1691 -821
rect 1567 -893 1691 -885
rect -93 -1417 31 -1411
rect -93 -1481 -67 -1417
rect -3 -1481 31 -1417
rect -93 -1489 31 -1481
rect 400 -1414 524 -1408
rect 400 -1478 426 -1414
rect 490 -1478 524 -1414
rect 400 -1486 524 -1478
rect 586 -1415 710 -1409
rect 586 -1479 612 -1415
rect 676 -1479 710 -1415
rect 586 -1487 710 -1479
rect 847 -2057 971 -2051
rect 847 -2121 873 -2057
rect 937 -2121 971 -2057
rect 847 -2129 971 -2121
rect 1032 -2056 1156 -2050
rect 1032 -2120 1058 -2056
rect 1122 -2120 1156 -2056
rect 1032 -2128 1156 -2120
rect 1222 -2056 1346 -2050
rect 1222 -2120 1248 -2056
rect 1312 -2120 1346 -2056
rect 1222 -2128 1346 -2120
rect 1406 -2057 1530 -2051
rect 1406 -2121 1432 -2057
rect 1496 -2121 1530 -2057
rect 1406 -2129 1530 -2121
rect 1590 -2060 1714 -2054
rect 1590 -2124 1616 -2060
rect 1680 -2124 1714 -2060
rect 1590 -2132 1714 -2124
rect -21 -2649 103 -2643
rect -21 -2713 5 -2649
rect 69 -2713 103 -2649
rect -21 -2721 103 -2713
rect 238 -2653 362 -2647
rect 238 -2717 264 -2653
rect 328 -2717 362 -2653
rect 238 -2725 362 -2717
rect 543 -2653 667 -2647
rect 543 -2717 569 -2653
rect 633 -2717 667 -2653
rect 543 -2725 667 -2717
<< via3 >>
rect 968 -827 1032 -824
rect 968 -883 972 -827
rect 972 -883 1028 -827
rect 1028 -883 1032 -827
rect 968 -888 1032 -883
rect 1169 -826 1233 -823
rect 1169 -882 1173 -826
rect 1173 -882 1229 -826
rect 1229 -882 1233 -826
rect 1169 -887 1233 -882
rect 1369 -823 1433 -820
rect 1369 -879 1373 -823
rect 1373 -879 1429 -823
rect 1429 -879 1433 -823
rect 1369 -884 1433 -879
rect 1593 -824 1657 -821
rect 1593 -880 1597 -824
rect 1597 -880 1653 -824
rect 1653 -880 1657 -824
rect 1593 -885 1657 -880
rect -67 -1420 -3 -1417
rect -67 -1476 -63 -1420
rect -63 -1476 -7 -1420
rect -7 -1476 -3 -1420
rect -67 -1481 -3 -1476
rect 426 -1417 490 -1414
rect 426 -1473 430 -1417
rect 430 -1473 486 -1417
rect 486 -1473 490 -1417
rect 426 -1478 490 -1473
rect 612 -1418 676 -1415
rect 612 -1474 616 -1418
rect 616 -1474 672 -1418
rect 672 -1474 676 -1418
rect 612 -1479 676 -1474
rect 873 -2060 937 -2057
rect 873 -2116 877 -2060
rect 877 -2116 933 -2060
rect 933 -2116 937 -2060
rect 873 -2121 937 -2116
rect 1058 -2059 1122 -2056
rect 1058 -2115 1062 -2059
rect 1062 -2115 1118 -2059
rect 1118 -2115 1122 -2059
rect 1058 -2120 1122 -2115
rect 1248 -2059 1312 -2056
rect 1248 -2115 1252 -2059
rect 1252 -2115 1308 -2059
rect 1308 -2115 1312 -2059
rect 1248 -2120 1312 -2115
rect 1432 -2060 1496 -2057
rect 1432 -2116 1436 -2060
rect 1436 -2116 1492 -2060
rect 1492 -2116 1496 -2060
rect 1432 -2121 1496 -2116
rect 1616 -2063 1680 -2060
rect 1616 -2119 1620 -2063
rect 1620 -2119 1676 -2063
rect 1676 -2119 1680 -2063
rect 1616 -2124 1680 -2119
rect 5 -2652 69 -2649
rect 5 -2708 9 -2652
rect 9 -2708 65 -2652
rect 65 -2708 69 -2652
rect 5 -2713 69 -2708
rect 264 -2656 328 -2653
rect 264 -2712 268 -2656
rect 268 -2712 324 -2656
rect 324 -2712 328 -2656
rect 264 -2717 328 -2712
rect 569 -2656 633 -2653
rect 569 -2712 573 -2656
rect 573 -2712 629 -2656
rect 629 -2712 633 -2656
rect 569 -2717 633 -2712
<< metal4 >>
rect -233 -1414 746 -804
rect -233 -1417 426 -1414
rect -233 -1481 -67 -1417
rect -3 -1478 426 -1417
rect 490 -1415 746 -1414
rect 490 -1478 612 -1415
rect -3 -1479 612 -1478
rect 676 -1479 746 -1415
rect -3 -1481 746 -1479
rect -233 -2649 746 -1481
rect -233 -2713 5 -2649
rect 69 -2653 746 -2649
rect 69 -2713 264 -2653
rect -233 -2717 264 -2713
rect 328 -2717 569 -2653
rect 633 -2717 746 -2653
rect -233 -2732 746 -2717
rect 826 -820 1795 -808
rect 826 -823 1369 -820
rect 826 -824 1169 -823
rect 826 -888 968 -824
rect 1032 -887 1169 -824
rect 1233 -884 1369 -823
rect 1433 -821 1795 -820
rect 1433 -884 1593 -821
rect 1233 -885 1593 -884
rect 1657 -885 1795 -821
rect 1233 -887 1795 -885
rect 1032 -888 1795 -887
rect 826 -2056 1795 -888
rect 826 -2057 1058 -2056
rect 826 -2121 873 -2057
rect 937 -2120 1058 -2057
rect 1122 -2120 1248 -2056
rect 1312 -2057 1795 -2056
rect 1312 -2120 1432 -2057
rect 937 -2121 1432 -2120
rect 1496 -2060 1795 -2057
rect 1496 -2121 1616 -2060
rect 826 -2124 1616 -2121
rect 1680 -2124 1795 -2060
rect 826 -2736 1795 -2124
use sky130_fd_sc_hd__buf_4  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698323353
transform -1 0 1240 0 -1 -1496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  x2
timestamp 1698323353
transform -1 0 700 0 -1 -1496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698323353
transform 1 0 964 0 1 -2680
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x4
timestamp 1698323353
transform 1 0 412 0 1 -2680
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x5
timestamp 1698323353
transform 1 0 -140 0 1 -2680
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x6
timestamp 1698323353
transform 1 0 136 0 1 -2680
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x7
timestamp 1698323353
transform 1 0 -128 0 -1 -1496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x8
timestamp 1698323353
transform -1 0 1516 0 1 -2680
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x9
timestamp 1698323353
transform 1 0 1516 0 1 -2680
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  x10
timestamp 1698323353
transform -1 0 1792 0 -1 -1496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_16  x11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698323353
transform -1 0 1792 0 1 -1400
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_1  x12
timestamp 1698323353
transform -1 0 964 0 1 -2680
box -38 -48 314 592
<< labels >>
flabel metal4 1680 -2736 1795 -808 0 FreeSans 320 0 0 0 VDD
port 0 nsew
flabel metal4 -233 -2732 -67 -804 0 FreeSans 320 0 0 0 VSS
port 1 nsew
flabel metal2 1550 -2793 1578 -2474 0 FreeSans 320 0 0 0 sar_val<7>
port 2 nsew
flabel metal2 991 -2788 1019 -2474 0 FreeSans 320 0 0 0 sar_val<6>
port 3 nsew
flabel metal2 446 -2793 474 -2476 0 FreeSans 320 0 0 0 sar_val<5>
port 4 nsew
flabel metal2 171 -2798 199 -2476 0 FreeSans 320 0 0 0 sar_val<4>
port 5 nsew
flabel metal2 -106 -2798 -78 -2476 0 FreeSans 320 0 0 0 sar_val<3>
port 6 nsew
flabel metal2 -204 -1133 -163 -714 0 FreeSans 320 0 0 0 sw<6>
port 7 nsew
flabel metal2 74 -2267 115 -714 0 FreeSans 320 0 0 0 sw<2>
port 8 nsew
flabel metal2 350 -2264 391 -714 0 FreeSans 320 0 0 0 sw<3>
port 9 nsew
flabel metal2 206 -1705 247 -714 0 FreeSans 320 0 0 0 sw<4>
port 10 nsew
flabel metal2 869 -1711 910 -714 0 FreeSans 320 0 0 0 sw<5>
port 11 nsew
<< end >>
