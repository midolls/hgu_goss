magic
tech sky130A
magscale 1 2
timestamp 1698584986
<< pwell >>
rect 689 963 715 995
<< nmos >>
rect 691 1701 721 1785
<< ndiff >>
rect 633 1773 691 1785
rect 633 1713 645 1773
rect 679 1713 691 1773
rect 633 1701 691 1713
rect 721 1773 779 1785
rect 721 1713 733 1773
rect 767 1713 779 1773
rect 721 1701 779 1713
<< ndiffc >>
rect 645 1713 679 1773
rect 733 1713 767 1773
<< poly >>
rect 691 1785 721 1811
rect 691 1679 721 1701
rect 673 1663 739 1679
rect 673 1629 689 1663
rect 723 1629 739 1663
rect 673 1613 739 1629
<< polycont >>
rect 689 1629 723 1663
<< locali >>
rect 645 1773 679 1789
rect 645 1697 679 1713
rect 733 1773 767 1789
rect 733 1697 767 1713
rect 673 1629 689 1663
rect 723 1629 739 1663
<< viali >>
rect 645 1713 679 1773
rect 733 1713 767 1773
rect 689 1629 723 1663
<< metal1 >>
rect 617 1723 623 1787
rect 687 1723 694 1787
rect 727 1773 773 1854
rect 639 1713 645 1723
rect 679 1713 685 1723
rect 639 1701 685 1713
rect 727 1713 733 1773
rect 767 1713 773 1773
rect 727 1701 773 1713
rect 677 1663 736 1669
rect 677 1629 689 1663
rect 723 1629 736 1663
rect 677 540 736 1629
<< via1 >>
rect 623 1773 687 1787
rect 623 1723 645 1773
rect 645 1723 679 1773
rect 679 1723 687 1773
<< metal2 >>
rect 614 1723 623 1787
rect 687 1723 696 1787
rect 614 1722 696 1723
<< via2 >>
rect 623 1723 687 1787
<< metal3 >>
rect 614 1787 696 1794
rect 614 1775 623 1787
rect 369 1773 623 1775
rect 687 1775 696 1787
rect 687 1773 1041 1775
rect 369 1709 473 1773
rect 537 1709 553 1773
rect 617 1723 623 1773
rect 617 1709 633 1723
rect 697 1709 713 1773
rect 777 1709 793 1773
rect 857 1709 873 1773
rect 937 1709 1041 1773
rect 369 1707 1041 1709
rect 369 1553 435 1707
rect 369 1489 370 1553
rect 434 1489 435 1553
rect 369 1473 435 1489
rect 369 1409 370 1473
rect 434 1409 435 1473
rect 369 1393 435 1409
rect 369 1329 370 1393
rect 434 1329 435 1393
rect 369 1313 435 1329
rect 369 1249 370 1313
rect 434 1249 435 1313
rect 369 1233 435 1249
rect 369 1169 370 1233
rect 434 1169 435 1233
rect 369 1153 435 1169
rect 369 1089 370 1153
rect 434 1089 435 1153
rect 369 1073 435 1089
rect 369 1009 370 1073
rect 434 1009 435 1073
rect 369 993 435 1009
rect 369 929 370 993
rect 434 929 435 993
rect 369 913 435 929
rect 369 849 370 913
rect 434 849 435 913
rect 369 833 435 849
rect 369 769 370 833
rect 434 769 435 833
rect 369 679 435 769
rect 495 675 555 1707
rect 615 615 675 1645
rect 735 675 795 1707
rect 855 615 915 1645
rect 975 1553 1041 1707
rect 975 1489 976 1553
rect 1040 1489 1041 1553
rect 975 1473 1041 1489
rect 975 1409 976 1473
rect 1040 1409 1041 1473
rect 975 1393 1041 1409
rect 975 1329 976 1393
rect 1040 1329 1041 1393
rect 975 1313 1041 1329
rect 975 1249 976 1313
rect 1040 1249 1041 1313
rect 975 1233 1041 1249
rect 975 1169 976 1233
rect 1040 1169 1041 1233
rect 975 1153 1041 1169
rect 975 1089 976 1153
rect 1040 1089 1041 1153
rect 975 1073 1041 1089
rect 975 1009 976 1073
rect 1040 1009 1041 1073
rect 975 993 1041 1009
rect 975 929 976 993
rect 1040 929 1041 993
rect 975 913 1041 929
rect 975 849 976 913
rect 1040 849 1041 913
rect 975 833 1041 849
rect 975 769 976 833
rect 1040 769 1041 833
rect 975 679 1041 769
rect 369 613 1041 615
rect 369 549 473 613
rect 537 549 553 613
rect 617 549 633 613
rect 697 549 713 613
rect 777 549 793 613
rect 857 549 873 613
rect 937 549 1041 613
rect 369 547 1041 549
<< via3 >>
rect 473 1709 537 1773
rect 553 1709 617 1773
rect 633 1723 687 1773
rect 687 1723 697 1773
rect 633 1709 697 1723
rect 713 1709 777 1773
rect 793 1709 857 1773
rect 873 1709 937 1773
rect 370 1489 434 1553
rect 370 1409 434 1473
rect 370 1329 434 1393
rect 370 1249 434 1313
rect 370 1169 434 1233
rect 370 1089 434 1153
rect 370 1009 434 1073
rect 370 929 434 993
rect 370 849 434 913
rect 370 769 434 833
rect 976 1489 1040 1553
rect 976 1409 1040 1473
rect 976 1329 1040 1393
rect 976 1249 1040 1313
rect 976 1169 1040 1233
rect 976 1089 1040 1153
rect 976 1009 1040 1073
rect 976 929 1040 993
rect 976 849 1040 913
rect 976 769 1040 833
rect 473 549 537 613
rect 553 549 617 613
rect 633 549 697 613
rect 713 549 777 613
rect 793 549 857 613
rect 873 549 937 613
<< metal4 >>
rect 369 1773 1041 1775
rect 369 1709 473 1773
rect 537 1709 553 1773
rect 617 1709 633 1773
rect 697 1709 713 1773
rect 777 1709 793 1773
rect 857 1709 873 1773
rect 937 1709 1041 1773
rect 369 1707 1041 1709
rect 369 1553 435 1707
rect 369 1489 370 1553
rect 434 1489 435 1553
rect 369 1473 435 1489
rect 369 1409 370 1473
rect 434 1409 435 1473
rect 369 1393 435 1409
rect 369 1329 370 1393
rect 434 1329 435 1393
rect 369 1313 435 1329
rect 369 1249 370 1313
rect 434 1249 435 1313
rect 369 1233 435 1249
rect 369 1169 370 1233
rect 434 1169 435 1233
rect 369 1153 435 1169
rect 369 1089 370 1153
rect 434 1089 435 1153
rect 369 1073 435 1089
rect 369 1009 370 1073
rect 434 1009 435 1073
rect 369 993 435 1009
rect 369 929 370 993
rect 434 929 435 993
rect 369 913 435 929
rect 369 849 370 913
rect 434 849 435 913
rect 369 833 435 849
rect 369 769 370 833
rect 434 769 435 833
rect 369 679 435 769
rect 495 615 555 1645
rect 615 675 675 1707
rect 735 615 795 1645
rect 855 675 915 1707
rect 975 1553 1041 1707
rect 975 1489 976 1553
rect 1040 1489 1041 1553
rect 975 1473 1041 1489
rect 975 1409 976 1473
rect 1040 1409 1041 1473
rect 975 1393 1041 1409
rect 975 1329 976 1393
rect 1040 1329 1041 1393
rect 975 1313 1041 1329
rect 975 1249 976 1313
rect 1040 1249 1041 1313
rect 975 1233 1041 1249
rect 975 1169 976 1233
rect 1040 1169 1041 1233
rect 975 1153 1041 1169
rect 975 1089 976 1153
rect 1040 1089 1041 1153
rect 975 1073 1041 1089
rect 975 1009 976 1073
rect 1040 1009 1041 1073
rect 975 993 1041 1009
rect 975 929 976 993
rect 1040 929 1041 993
rect 975 913 1041 929
rect 975 849 976 913
rect 1040 849 1041 913
rect 975 833 1041 849
rect 975 769 976 833
rect 1040 769 1041 833
rect 975 679 1041 769
rect 369 613 1041 615
rect 369 549 473 613
rect 537 549 553 613
rect 617 549 633 613
rect 697 549 713 613
rect 777 549 793 613
rect 857 549 873 613
rect 937 549 1041 613
rect 369 547 1041 549
<< labels >>
flabel pwell 689 963 715 995 0 FreeSans 160 0 0 0 x2.SUB
flabel metal4 631 1297 657 1329 0 FreeSans 320 0 0 0 x2.CBOT
flabel metal4 749 707 775 739 0 FreeSans 320 0 0 0 x2.CTOP
<< end >>
