magic
tech sky130A
magscale 1 2
timestamp 1698843163
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
use sky130_fd_pr__pfet_01v8_M479BZ  XM16
timestamp 0
transform 1 0 158 0 1 808
box 0 0 1 1
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 SW
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 DELAY_SIGNAL
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 VDD
port 2 nsew
<< end >>
