magic
tech sky130A
timestamp 1698475227
<< end >>
