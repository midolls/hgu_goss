* NGSPICE file created from hgu_delay_no_code_flat.ext - technology: sky130A

.subckt hgu_delay_no_code_flat IN OUT VDD code[3] code_offset code[0] code[1] code[2]
+ VSS
X0 a_9939_2268# IN a_9851_2130# x5.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X1 a_9939_2130# x1.Y x5[7].x1.CBOT x5.VPB sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X2 x5[7].x1.CBOT x1.Y a_9939_2130# x5.VPB sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X3 a_15703_1340# OUT VDD x5.VNB sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_9939_2130# code[2] x4[3].x2.CBOT x5.VNB sky130_fd_pr__nfet_01v8 ad=0.0987 pd=0.89 as=0.122 ps=1.42 w=0.42 l=0.15
X5 a_9893_879# IN a_9805_879# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X6 a_9965_465# IN a_9893_465# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X7 a_9939_2544# IN a_9851_2682# x5.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X8 a_9965_1017# IN a_9893_1017# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 a_15703_1340# a_9939_2130# VSS x5.VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X10 a_15703_1681# a_9939_2130# OUT x5.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X11 VDD OUT a_15703_1340# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X12 a_9893_465# IN a_9805_327# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X13 VDD code_offset x5.Y x5.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X14 x2.x2.CBOT code[0] a_9939_2130# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X15 VSS IN a_9893_327# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X16 a_9939_2544# IN a_9851_2406# x5.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X17 x3[1].x2.CBOT code[1] a_9939_2130# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0987 ps=0.89 w=0.42 l=0.15
X18 a_9939_2130# x1.Y x5[7].x1.CBOT x5.VPB sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X19 x5[7].x1.CBOT x1.Y a_9939_2130# x5.VPB sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X20 a_9965_741# IN a_9893_741# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X21 a_9893_327# IN a_9805_327# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X22 x1.Y code[3] VDD x5.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X23 a_15703_1681# a_9939_2130# VDD x5.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X24 a_9939_2130# code_offset x7.x2.CBOT x5.VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X25 a_9939_2130# code[2] x4[3].x2.CBOT x5.VNB sky130_fd_pr__nfet_01v8 ad=0.0987 pd=0.89 as=0.122 ps=1.42 w=0.42 l=0.15
X26 x4[3].x2.CBOT code[2] a_9939_2130# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0987 ps=0.89 w=0.42 l=0.15
X27 a_9939_2130# IN a_9851_2130# x5.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X28 a_9939_2130# x5.Y x6.x1.CBOT x5.VPB sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X29 a_9939_2268# IN a_9851_2406# x5.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X30 VSS code_offset x5.Y x5.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X31 a_9893_1293# IN a_9805_1155# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X32 x5[7].x1.CBOT x1.Y a_9939_2130# x5.VPB sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X33 a_15703_1681# OUT VSS x5.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 a_9893_741# IN a_9805_603# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X35 x5[7].x1.CBOT x1.Y a_9939_2130# x5.VPB sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X36 a_9939_2130# x1.Y x5[7].x1.CBOT x5.VPB sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X37 a_9965_465# IN a_9893_603# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X38 VDD IN a_9851_2682# x5.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X39 a_15703_1340# a_9939_2130# OUT x5.VNB sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X40 a_9939_2130# IN a_9893_1293# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X41 x1.Y code[3] VSS x5.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X42 a_9893_1155# IN a_9805_1155# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X43 a_9939_2130# x1.Y x5[7].x1.CBOT x5.VPB sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X44 VSS OUT a_15703_1681# x5.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X45 a_9893_603# IN a_9805_603# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X46 x4[3].x2.CBOT code[2] a_9939_2130# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0987 ps=0.89 w=0.42 l=0.15
X47 a_9965_1017# IN a_9893_1155# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X48 a_9965_741# IN a_9893_879# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X49 a_9939_2130# code[1] x3[1].x2.CBOT x5.VNB sky130_fd_pr__nfet_01v8 ad=0.0987 pd=0.89 as=0.122 ps=1.42 w=0.42 l=0.15
X50 a_9893_1017# IN a_9805_879# x5.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
.ends

