magic
tech sky130A
magscale 1 2
timestamp 1699514362
<< nwell >>
rect 2532 94 2608 112
rect 1406 76 1434 78
rect 1044 -42 1110 24
rect 1434 12 1498 76
rect 1928 12 1966 34
rect 338 -1944 2010 -1508
<< psubdiff >>
rect 826 -336 1338 -324
rect 826 -370 868 -336
rect 902 -370 968 -336
rect 1002 -370 1068 -336
rect 1102 -370 1168 -336
rect 1202 -370 1268 -336
rect 1302 -370 1338 -336
rect 826 -382 1338 -370
rect 2028 -336 2540 -324
rect 2028 -370 2070 -336
rect 2104 -370 2170 -336
rect 2204 -370 2270 -336
rect 2304 -370 2370 -336
rect 2404 -370 2470 -336
rect 2504 -370 2540 -336
rect 2028 -382 2540 -370
rect 544 -836 2834 -812
rect 544 -870 568 -836
rect 602 -870 668 -836
rect 702 -870 768 -836
rect 802 -870 868 -836
rect 902 -870 968 -836
rect 1002 -870 1068 -836
rect 1102 -870 1168 -836
rect 1202 -870 1268 -836
rect 1302 -870 1368 -836
rect 1402 -870 1468 -836
rect 1502 -870 1568 -836
rect 1602 -870 1668 -836
rect 1702 -870 1768 -836
rect 1802 -870 1868 -836
rect 1902 -870 1968 -836
rect 2002 -870 2068 -836
rect 2102 -870 2168 -836
rect 2202 -870 2268 -836
rect 2302 -870 2368 -836
rect 2402 -870 2468 -836
rect 2502 -870 2568 -836
rect 2602 -870 2668 -836
rect 2702 -870 2768 -836
rect 2802 -870 2834 -836
rect 544 -952 2834 -870
rect 472 -976 2834 -952
rect 472 -1010 496 -976
rect 530 -1010 568 -976
rect 602 -1010 668 -976
rect 702 -980 2834 -976
rect 702 -1010 1568 -980
rect 472 -1014 1568 -1010
rect 1602 -1014 1668 -980
rect 1702 -1014 1768 -980
rect 1802 -1014 2834 -980
rect 472 -1034 2834 -1014
rect 764 -1038 2834 -1034
rect 764 -1062 1516 -1038
rect 764 -1096 770 -1062
rect 804 -1096 868 -1062
rect 902 -1096 968 -1062
rect 1002 -1096 1068 -1062
rect 1102 -1096 1168 -1062
rect 1202 -1096 1268 -1062
rect 1302 -1096 1368 -1062
rect 1402 -1096 1468 -1062
rect 1502 -1096 1516 -1062
rect 764 -1120 1516 -1096
rect 1860 -1062 2834 -1038
rect 1860 -1096 1868 -1062
rect 1902 -1096 1968 -1062
rect 2002 -1096 2068 -1062
rect 2102 -1096 2168 -1062
rect 2202 -1096 2268 -1062
rect 2302 -1096 2368 -1062
rect 2402 -1096 2468 -1062
rect 2502 -1096 2568 -1062
rect 2602 -1096 2668 -1062
rect 2702 -1096 2768 -1062
rect 2802 -1096 2834 -1062
rect 1860 -1120 2834 -1096
<< nsubdiff >>
rect 762 412 2624 428
rect 762 378 802 412
rect 836 378 958 412
rect 992 378 1114 412
rect 1148 378 1270 412
rect 1304 378 1426 412
rect 1460 378 1582 412
rect 1616 378 1738 412
rect 1772 378 1894 412
rect 1928 378 2050 412
rect 2084 378 2206 412
rect 2240 378 2362 412
rect 2396 378 2518 412
rect 2552 378 2624 412
rect 762 364 2624 378
rect 758 -1792 2440 -1776
rect 758 -1826 818 -1792
rect 852 -1826 958 -1792
rect 992 -1826 1114 -1792
rect 1148 -1826 1270 -1792
rect 1304 -1826 1426 -1792
rect 1460 -1826 1582 -1792
rect 1616 -1826 1738 -1792
rect 1772 -1826 1894 -1792
rect 1928 -1826 2050 -1792
rect 2084 -1826 2206 -1792
rect 2240 -1826 2362 -1792
rect 2396 -1826 2440 -1792
rect 758 -1840 2440 -1826
<< psubdiffcont >>
rect 868 -370 902 -336
rect 968 -370 1002 -336
rect 1068 -370 1102 -336
rect 1168 -370 1202 -336
rect 1268 -370 1302 -336
rect 2070 -370 2104 -336
rect 2170 -370 2204 -336
rect 2270 -370 2304 -336
rect 2370 -370 2404 -336
rect 2470 -370 2504 -336
rect 568 -870 602 -836
rect 668 -870 702 -836
rect 768 -870 802 -836
rect 868 -870 902 -836
rect 968 -870 1002 -836
rect 1068 -870 1102 -836
rect 1168 -870 1202 -836
rect 1268 -870 1302 -836
rect 1368 -870 1402 -836
rect 1468 -870 1502 -836
rect 1568 -870 1602 -836
rect 1668 -870 1702 -836
rect 1768 -870 1802 -836
rect 1868 -870 1902 -836
rect 1968 -870 2002 -836
rect 2068 -870 2102 -836
rect 2168 -870 2202 -836
rect 2268 -870 2302 -836
rect 2368 -870 2402 -836
rect 2468 -870 2502 -836
rect 2568 -870 2602 -836
rect 2668 -870 2702 -836
rect 2768 -870 2802 -836
rect 496 -1010 530 -976
rect 568 -1010 602 -976
rect 668 -1010 702 -976
rect 1568 -1014 1602 -980
rect 1668 -1014 1702 -980
rect 1768 -1014 1802 -980
rect 770 -1096 804 -1062
rect 868 -1096 902 -1062
rect 968 -1096 1002 -1062
rect 1068 -1096 1102 -1062
rect 1168 -1096 1202 -1062
rect 1268 -1096 1302 -1062
rect 1368 -1096 1402 -1062
rect 1468 -1096 1502 -1062
rect 1868 -1096 1902 -1062
rect 1968 -1096 2002 -1062
rect 2068 -1096 2102 -1062
rect 2168 -1096 2202 -1062
rect 2268 -1096 2302 -1062
rect 2368 -1096 2402 -1062
rect 2468 -1096 2502 -1062
rect 2568 -1096 2602 -1062
rect 2668 -1096 2702 -1062
rect 2768 -1096 2802 -1062
<< nsubdiffcont >>
rect 802 378 836 412
rect 958 378 992 412
rect 1114 378 1148 412
rect 1270 378 1304 412
rect 1426 378 1460 412
rect 1582 378 1616 412
rect 1738 378 1772 412
rect 1894 378 1928 412
rect 2050 378 2084 412
rect 2206 378 2240 412
rect 2362 378 2396 412
rect 2518 378 2552 412
rect 818 -1826 852 -1792
rect 958 -1826 992 -1792
rect 1114 -1826 1148 -1792
rect 1270 -1826 1304 -1792
rect 1426 -1826 1460 -1792
rect 1582 -1826 1616 -1792
rect 1738 -1826 1772 -1792
rect 1894 -1826 1928 -1792
rect 2050 -1826 2084 -1792
rect 2206 -1826 2240 -1792
rect 2362 -1826 2396 -1792
<< poly >>
rect 1044 24 1074 96
rect 1044 8 1110 24
rect 1044 -26 1060 8
rect 1094 -26 1110 8
rect 1044 -42 1110 -26
rect 1248 -22 1278 114
rect 1432 64 1566 94
rect 1432 62 1498 64
rect 1432 28 1448 62
rect 1482 28 1498 62
rect 1432 12 1498 28
rect 1624 -8 1654 78
rect 1248 -38 1328 -22
rect 1536 -38 1654 -8
rect 1044 -132 1074 -42
rect 1248 -72 1278 -38
rect 1312 -72 1328 -38
rect 1248 -88 1328 -72
rect 1488 -50 1566 -38
rect 1488 -84 1504 -50
rect 1538 -84 1566 -50
rect 1248 -152 1278 -88
rect 1488 -96 1566 -84
rect 1536 -154 1566 -96
rect 1712 -86 1742 78
rect 1800 64 1934 94
rect 1868 62 1934 64
rect 1868 28 1884 62
rect 1918 28 1934 62
rect 1868 12 1934 28
rect 2088 -86 2118 114
rect 2292 24 2322 96
rect 2256 8 2322 24
rect 2256 -26 2272 8
rect 2306 -26 2322 8
rect 2256 -42 2322 -26
rect 1712 -94 1832 -86
rect 1712 -106 1880 -94
rect 1712 -116 1830 -106
rect 1800 -140 1830 -116
rect 1864 -140 1880 -106
rect 1800 -150 1880 -140
rect 2036 -102 2118 -86
rect 2036 -136 2052 -102
rect 2086 -136 2118 -102
rect 2292 -132 2322 -42
rect 1800 -152 1878 -150
rect 2036 -152 2118 -136
rect 1800 -160 1830 -152
rect 1650 -398 1716 -384
rect 1650 -432 1666 -398
rect 1700 -432 1716 -398
rect 1650 -446 1716 -432
rect 534 -1526 564 -1292
rect 622 -1456 652 -1292
rect 768 -1306 852 -1290
rect 768 -1340 784 -1306
rect 818 -1340 852 -1306
rect 768 -1356 852 -1340
rect 622 -1472 704 -1456
rect 622 -1506 654 -1472
rect 688 -1506 704 -1472
rect 622 -1522 704 -1506
rect 822 -1522 852 -1356
rect 1216 -1394 1248 -1312
rect 1422 -1394 1452 -1292
rect 1592 -1300 1658 -1286
rect 1592 -1334 1608 -1300
rect 1642 -1334 1658 -1300
rect 1592 -1348 1658 -1334
rect 1716 -1300 1782 -1286
rect 1716 -1334 1732 -1300
rect 1766 -1334 1782 -1300
rect 1716 -1348 1782 -1334
rect 1216 -1408 1314 -1394
rect 1216 -1442 1264 -1408
rect 1298 -1442 1314 -1408
rect 1216 -1456 1314 -1442
rect 1422 -1408 1506 -1394
rect 1422 -1442 1456 -1408
rect 1490 -1442 1506 -1408
rect 1422 -1456 1506 -1442
rect 1716 -1404 1782 -1390
rect 1920 -1394 1950 -1292
rect 2124 -1394 2156 -1312
rect 1716 -1438 1732 -1404
rect 1766 -1438 1782 -1404
rect 1716 -1452 1782 -1438
rect 1872 -1408 1950 -1394
rect 1872 -1442 1888 -1408
rect 1922 -1442 1950 -1408
rect 1216 -1508 1248 -1456
rect 1422 -1522 1452 -1456
rect 1592 -1472 1658 -1458
rect 1592 -1506 1608 -1472
rect 1642 -1506 1658 -1472
rect 1592 -1520 1658 -1506
rect 622 -1526 652 -1522
rect 1628 -1532 1658 -1520
rect 1716 -1526 1746 -1452
rect 1872 -1456 1950 -1442
rect 2060 -1408 2156 -1394
rect 2060 -1442 2076 -1408
rect 2110 -1442 2156 -1408
rect 2060 -1456 2156 -1442
rect 1920 -1526 1950 -1456
rect 2124 -1508 2156 -1456
rect 534 -1752 564 -1748
rect 482 -1768 564 -1752
rect 482 -1802 498 -1768
rect 532 -1802 564 -1768
rect 482 -1818 564 -1802
<< polycont >>
rect 1060 -26 1094 8
rect 1448 28 1482 62
rect 1278 -72 1312 -38
rect 1504 -84 1538 -50
rect 1884 28 1918 62
rect 2272 -26 2306 8
rect 1830 -140 1864 -106
rect 2052 -136 2086 -102
rect 1666 -432 1700 -398
rect 784 -1340 818 -1306
rect 654 -1506 688 -1472
rect 1608 -1334 1642 -1300
rect 1732 -1334 1766 -1300
rect 1264 -1442 1298 -1408
rect 1456 -1442 1490 -1408
rect 1732 -1438 1766 -1404
rect 1888 -1442 1922 -1408
rect 1608 -1506 1642 -1472
rect 2076 -1442 2110 -1408
rect 498 -1802 532 -1768
<< locali >>
rect 762 412 2624 428
rect 762 378 802 412
rect 836 378 958 412
rect 992 378 1114 412
rect 1148 378 1270 412
rect 1304 378 1426 412
rect 1460 378 1582 412
rect 1616 378 1738 412
rect 1772 378 1894 412
rect 1928 378 2050 412
rect 2084 378 2206 412
rect 2240 378 2362 412
rect 2396 378 2518 412
rect 2552 378 2624 412
rect 762 364 2624 378
rect 1432 28 1448 62
rect 1482 28 1498 62
rect 1868 28 1884 62
rect 1918 28 1934 62
rect 1044 -26 1060 8
rect 1094 -26 1110 8
rect 2256 -26 2272 8
rect 2306 -26 2322 8
rect 1262 -72 1278 -38
rect 1312 -72 1328 -38
rect 1488 -84 1504 -50
rect 1538 -84 1554 -50
rect 1812 -140 1830 -106
rect 1864 -140 1880 -106
rect 2036 -136 2052 -102
rect 2086 -136 2102 -102
rect 826 -336 1338 -324
rect 826 -370 868 -336
rect 902 -370 968 -336
rect 1002 -370 1068 -336
rect 1102 -370 1168 -336
rect 1202 -370 1268 -336
rect 1302 -370 1338 -336
rect 826 -382 1338 -370
rect 2028 -336 2540 -324
rect 2028 -370 2070 -336
rect 2104 -370 2170 -336
rect 2204 -370 2270 -336
rect 2304 -370 2370 -336
rect 2404 -370 2470 -336
rect 2504 -370 2540 -336
rect 2028 -382 2540 -370
rect 1650 -432 1666 -398
rect 1700 -432 1716 -398
rect 1570 -812 1604 -690
rect 1762 -812 1796 -690
rect 544 -836 2834 -812
rect 544 -870 568 -836
rect 602 -870 668 -836
rect 702 -870 768 -836
rect 802 -870 868 -836
rect 902 -870 968 -836
rect 1002 -870 1068 -836
rect 1102 -870 1168 -836
rect 1202 -870 1268 -836
rect 1302 -870 1368 -836
rect 1402 -870 1468 -836
rect 1502 -870 1568 -836
rect 1602 -870 1668 -836
rect 1702 -870 1768 -836
rect 1802 -870 1868 -836
rect 1902 -870 1968 -836
rect 2002 -870 2068 -836
rect 2102 -870 2168 -836
rect 2202 -870 2268 -836
rect 2302 -870 2368 -836
rect 2402 -870 2468 -836
rect 2502 -870 2568 -836
rect 2602 -870 2668 -836
rect 2702 -870 2768 -836
rect 2802 -870 2834 -836
rect 544 -952 2834 -870
rect 472 -976 2834 -952
rect 472 -1010 496 -976
rect 530 -1010 568 -976
rect 602 -1010 668 -976
rect 702 -980 2834 -976
rect 702 -1010 1568 -980
rect 472 -1014 1568 -1010
rect 1602 -1014 1668 -980
rect 1702 -1014 1768 -980
rect 1802 -1014 2834 -980
rect 472 -1034 2834 -1014
rect 488 -1108 522 -1034
rect 764 -1038 2834 -1034
rect 764 -1062 1516 -1038
rect 764 -1096 770 -1062
rect 804 -1096 868 -1062
rect 902 -1096 968 -1062
rect 1002 -1096 1068 -1062
rect 1102 -1096 1168 -1062
rect 1202 -1096 1268 -1062
rect 1302 -1096 1368 -1062
rect 1402 -1096 1468 -1062
rect 1502 -1096 1516 -1062
rect 764 -1120 1516 -1096
rect 1860 -1062 2834 -1038
rect 1860 -1096 1868 -1062
rect 1902 -1096 1968 -1062
rect 2002 -1096 2068 -1062
rect 2102 -1096 2168 -1062
rect 2202 -1096 2268 -1062
rect 2302 -1096 2368 -1062
rect 2402 -1096 2468 -1062
rect 2502 -1096 2568 -1062
rect 2602 -1096 2668 -1062
rect 2702 -1096 2768 -1062
rect 2802 -1096 2834 -1062
rect 1860 -1120 2834 -1096
rect 1874 -1122 1908 -1120
rect 768 -1340 784 -1306
rect 818 -1340 834 -1306
rect 1592 -1334 1608 -1300
rect 1642 -1334 1658 -1300
rect 1716 -1334 1732 -1300
rect 1766 -1334 1782 -1300
rect 1248 -1442 1264 -1408
rect 1298 -1442 1314 -1408
rect 1440 -1442 1456 -1408
rect 1490 -1442 1506 -1408
rect 1716 -1438 1732 -1404
rect 1766 -1438 1782 -1404
rect 1872 -1442 1888 -1408
rect 1922 -1442 1938 -1408
rect 2060 -1442 2076 -1408
rect 2110 -1442 2126 -1408
rect 488 -1506 654 -1472
rect 688 -1506 704 -1472
rect 1592 -1506 1608 -1472
rect 1642 -1506 1658 -1472
rect 488 -1550 522 -1506
rect 664 -1768 698 -1709
rect 482 -1802 498 -1768
rect 532 -1802 698 -1768
rect 758 -1792 2440 -1776
rect 758 -1826 818 -1792
rect 852 -1826 958 -1792
rect 992 -1826 1114 -1792
rect 1148 -1826 1270 -1792
rect 1304 -1826 1426 -1792
rect 1460 -1826 1582 -1792
rect 1616 -1826 1738 -1792
rect 1772 -1826 1894 -1792
rect 1928 -1826 2050 -1792
rect 2084 -1826 2206 -1792
rect 2240 -1826 2362 -1792
rect 2396 -1826 2440 -1792
rect 758 -1840 2440 -1826
<< viali >>
rect 802 378 836 412
rect 958 378 992 412
rect 1114 378 1148 412
rect 1270 378 1304 412
rect 1426 378 1460 412
rect 1582 378 1616 412
rect 1738 378 1772 412
rect 1894 378 1928 412
rect 2050 378 2084 412
rect 2206 378 2240 412
rect 2362 378 2396 412
rect 2518 378 2552 412
rect 1448 28 1482 62
rect 1884 28 1918 62
rect 1060 -26 1094 8
rect 2272 -26 2306 8
rect 1278 -72 1312 -38
rect 1504 -84 1538 -50
rect 1830 -140 1864 -106
rect 2052 -136 2086 -102
rect 868 -370 902 -336
rect 968 -370 1002 -336
rect 1068 -370 1102 -336
rect 1168 -370 1202 -336
rect 1268 -370 1302 -336
rect 2070 -370 2104 -336
rect 2170 -370 2204 -336
rect 2270 -370 2304 -336
rect 2370 -370 2404 -336
rect 2470 -370 2504 -336
rect 1666 -432 1700 -398
rect 568 -870 602 -836
rect 668 -870 702 -836
rect 768 -870 802 -836
rect 868 -870 902 -836
rect 968 -870 1002 -836
rect 1068 -870 1102 -836
rect 1168 -870 1202 -836
rect 1268 -870 1302 -836
rect 1368 -870 1402 -836
rect 1468 -870 1502 -836
rect 1568 -870 1602 -836
rect 1668 -870 1702 -836
rect 1768 -870 1802 -836
rect 1868 -870 1902 -836
rect 1968 -870 2002 -836
rect 2068 -870 2102 -836
rect 2168 -870 2202 -836
rect 2268 -870 2302 -836
rect 2368 -870 2402 -836
rect 2468 -870 2502 -836
rect 2568 -870 2602 -836
rect 2668 -870 2702 -836
rect 2768 -870 2802 -836
rect 496 -1010 530 -976
rect 568 -1010 602 -976
rect 668 -1010 702 -976
rect 1568 -1014 1602 -980
rect 1668 -1014 1702 -980
rect 1768 -1014 1802 -980
rect 770 -1096 804 -1062
rect 868 -1096 902 -1062
rect 968 -1096 1002 -1062
rect 1068 -1096 1102 -1062
rect 1168 -1096 1202 -1062
rect 1268 -1096 1302 -1062
rect 1368 -1096 1402 -1062
rect 1468 -1096 1502 -1062
rect 1868 -1096 1902 -1062
rect 1968 -1096 2002 -1062
rect 2068 -1096 2102 -1062
rect 2168 -1096 2202 -1062
rect 2268 -1096 2302 -1062
rect 2368 -1096 2402 -1062
rect 2468 -1096 2502 -1062
rect 2568 -1096 2602 -1062
rect 2668 -1096 2702 -1062
rect 2768 -1096 2802 -1062
rect 784 -1340 818 -1306
rect 1608 -1334 1642 -1300
rect 1732 -1334 1766 -1300
rect 1264 -1442 1298 -1408
rect 1456 -1442 1490 -1408
rect 1732 -1438 1766 -1404
rect 1888 -1442 1922 -1408
rect 2076 -1442 2110 -1408
rect 654 -1506 688 -1472
rect 1608 -1506 1642 -1472
rect 498 -1802 532 -1768
rect 818 -1826 852 -1792
rect 958 -1826 992 -1792
rect 1114 -1826 1148 -1792
rect 1270 -1826 1304 -1792
rect 1426 -1826 1460 -1792
rect 1582 -1826 1616 -1792
rect 1738 -1826 1772 -1792
rect 1894 -1826 1928 -1792
rect 2050 -1826 2084 -1792
rect 2206 -1826 2240 -1792
rect 2362 -1826 2396 -1792
<< metal1 >>
rect 762 424 2624 428
rect 762 422 1104 424
rect 762 370 794 422
rect 846 370 952 422
rect 1004 372 1104 422
rect 1156 372 1264 424
rect 1316 372 1418 424
rect 1470 422 2200 424
rect 1470 372 1574 422
rect 1004 370 1574 372
rect 1626 370 1728 422
rect 1780 370 1886 422
rect 1938 370 2040 422
rect 2092 372 2200 422
rect 2252 422 2624 424
rect 2252 372 2354 422
rect 2092 370 2354 372
rect 2406 370 2510 422
rect 2562 370 2624 422
rect 762 364 2624 370
rect 898 297 932 364
rect 1090 297 1124 364
rect 1290 297 1324 364
rect 1490 304 1524 364
rect 1666 290 1700 364
rect 1842 297 1876 364
rect 2042 297 2076 364
rect 2242 297 2276 364
rect 2434 297 2468 364
rect 802 100 836 150
rect 994 100 1028 142
rect 802 66 1028 100
rect 802 -60 836 66
rect 1044 16 1108 22
rect 1044 -36 1050 16
rect 1102 8 1108 16
rect 1202 8 1236 154
rect 1102 -26 1236 8
rect 1102 -36 1108 -26
rect 1044 -42 1108 -36
rect 802 -72 878 -60
rect 802 -124 814 -72
rect 866 -102 878 -72
rect 866 -124 1028 -102
rect 802 -136 1028 -124
rect 802 -188 836 -136
rect 994 -178 1028 -136
rect 1202 -218 1236 -26
rect 1264 -28 1328 -22
rect 1264 -80 1270 -28
rect 1322 -80 1328 -28
rect 1264 -86 1328 -80
rect 898 -324 932 -218
rect 1090 -324 1124 -228
rect 1290 -324 1324 -240
rect 826 -330 1338 -324
rect 566 -390 642 -372
rect 826 -382 860 -330
rect 912 -336 1338 -330
rect 912 -370 968 -336
rect 1002 -370 1068 -336
rect 1102 -370 1168 -336
rect 1202 -370 1268 -336
rect 1302 -370 1338 -336
rect 912 -382 1338 -370
rect 566 -442 578 -390
rect 630 -442 642 -390
rect 1374 -418 1402 138
rect 1434 70 1498 76
rect 1434 68 1440 70
rect 1432 22 1440 68
rect 1434 18 1440 22
rect 1492 18 1498 70
rect 1434 12 1498 18
rect 1486 -40 1550 -34
rect 1486 -92 1492 -40
rect 1544 -92 1550 -40
rect 1486 -98 1550 -92
rect 1578 -86 1612 112
rect 1650 74 1714 80
rect 1650 22 1656 74
rect 1708 22 1714 74
rect 1650 16 1714 22
rect 1578 -92 1642 -86
rect 1578 -144 1584 -92
rect 1636 -144 1642 -92
rect 1578 -150 1642 -144
rect 1578 -184 1612 -150
rect 1670 -214 1698 16
rect 1754 -18 1788 110
rect 1868 70 1932 76
rect 1868 18 1874 70
rect 1926 18 1932 70
rect 1868 12 1932 18
rect 1726 -24 1790 -18
rect 1726 -76 1732 -24
rect 1784 -76 1790 -24
rect 1726 -82 1790 -76
rect 1754 -180 1788 -82
rect 1818 -92 1882 -86
rect 1818 -144 1824 -92
rect 1876 -144 1882 -92
rect 1818 -150 1882 -144
rect 1650 -220 1714 -214
rect 1650 -272 1656 -220
rect 1708 -272 1714 -220
rect 1650 -278 1714 -272
rect 1490 -418 1524 -376
rect 1670 -382 1698 -278
rect 566 -448 642 -442
rect 690 -446 1524 -418
rect 1650 -388 1714 -382
rect 1650 -440 1656 -388
rect 1708 -440 1714 -388
rect 1650 -446 1714 -440
rect 1842 -418 1876 -364
rect 1960 -418 1988 138
rect 2130 8 2164 142
rect 2338 100 2372 142
rect 2530 112 2564 142
rect 2530 100 2608 112
rect 2338 66 2544 100
rect 2530 48 2544 66
rect 2596 48 2608 100
rect 2530 36 2608 48
rect 2256 16 2320 22
rect 2256 8 2262 16
rect 2130 -26 2262 8
rect 2036 -92 2100 -86
rect 2036 -144 2042 -92
rect 2094 -144 2100 -92
rect 2036 -150 2100 -144
rect 2130 -178 2164 -26
rect 2256 -36 2262 -26
rect 2314 -36 2320 16
rect 2256 -42 2320 -36
rect 2530 -102 2564 36
rect 2338 -136 2564 -102
rect 2338 -178 2372 -136
rect 2530 -178 2564 -136
rect 2042 -324 2076 -178
rect 2242 -324 2276 -258
rect 2434 -324 2468 -258
rect 2028 -330 2540 -324
rect 2028 -336 2460 -330
rect 2028 -370 2070 -336
rect 2104 -370 2170 -336
rect 2204 -370 2270 -336
rect 2304 -370 2370 -336
rect 2404 -370 2460 -336
rect 2028 -382 2460 -370
rect 2512 -382 2540 -330
rect 2454 -388 2518 -382
rect 2724 -390 2788 -384
rect 1842 -446 2676 -418
rect 690 -502 724 -446
rect 882 -506 916 -446
rect 1074 -506 1108 -446
rect 1266 -504 1300 -446
rect 2066 -506 2100 -446
rect 2258 -504 2292 -446
rect 2450 -508 2484 -446
rect 2642 -508 2676 -446
rect 2724 -442 2730 -390
rect 2782 -442 2788 -390
rect 2724 -448 2788 -442
rect 594 -756 628 -694
rect 786 -756 820 -694
rect 978 -756 1012 -696
rect 1170 -756 1204 -694
rect 1362 -756 1396 -698
rect 1474 -756 1508 -694
rect 1666 -756 1700 -690
rect 1858 -756 1892 -696
rect 1970 -756 2004 -694
rect 2162 -756 2196 -698
rect 2354 -756 2388 -694
rect 2546 -756 2580 -692
rect 2738 -756 2772 -692
rect 594 -784 2772 -756
rect 544 -818 2834 -812
rect 544 -836 860 -818
rect 912 -836 2460 -818
rect 2512 -836 2834 -818
rect 544 -870 568 -836
rect 602 -870 668 -836
rect 702 -870 768 -836
rect 802 -870 860 -836
rect 912 -870 968 -836
rect 1002 -870 1068 -836
rect 1102 -870 1168 -836
rect 1202 -870 1268 -836
rect 1302 -870 1368 -836
rect 1402 -870 1468 -836
rect 1502 -870 1568 -836
rect 1602 -870 1668 -836
rect 1702 -870 1768 -836
rect 1802 -870 1868 -836
rect 1902 -870 1968 -836
rect 2002 -870 2068 -836
rect 2102 -870 2168 -836
rect 2202 -870 2268 -836
rect 2302 -870 2368 -836
rect 2402 -870 2460 -836
rect 2512 -870 2568 -836
rect 2602 -870 2668 -836
rect 2702 -870 2768 -836
rect 2802 -870 2834 -836
rect 544 -900 2834 -870
rect 544 -952 2676 -900
rect 472 -976 2676 -952
rect 472 -1010 496 -976
rect 530 -1010 568 -976
rect 602 -1010 668 -976
rect 702 -980 2676 -976
rect 702 -1010 1568 -980
rect 472 -1014 1568 -1010
rect 1602 -1014 1668 -980
rect 1702 -1014 1768 -980
rect 1802 -1010 2676 -980
rect 2786 -1010 2834 -900
rect 1802 -1014 2834 -1010
rect 472 -1034 2834 -1014
rect 764 -1038 2834 -1034
rect 764 -1062 1516 -1038
rect 764 -1096 770 -1062
rect 804 -1096 868 -1062
rect 902 -1096 968 -1062
rect 1002 -1096 1068 -1062
rect 1102 -1096 1168 -1062
rect 1202 -1096 1268 -1062
rect 1302 -1096 1368 -1062
rect 1402 -1096 1468 -1062
rect 1502 -1096 1516 -1062
rect 764 -1120 1516 -1096
rect 1670 -1104 1704 -1038
rect 1860 -1062 2834 -1038
rect 1860 -1096 1868 -1062
rect 1902 -1096 1968 -1062
rect 2002 -1096 2068 -1062
rect 2102 -1096 2168 -1062
rect 2202 -1096 2268 -1062
rect 2302 -1096 2368 -1062
rect 2402 -1096 2468 -1062
rect 2502 -1096 2568 -1062
rect 2602 -1096 2668 -1062
rect 2702 -1096 2768 -1062
rect 2802 -1096 2834 -1062
rect 1860 -1120 2834 -1096
rect 776 -1196 810 -1120
rect 1072 -1186 1106 -1120
rect 1264 -1186 1298 -1120
rect 1464 -1194 1498 -1120
rect 1874 -1194 1908 -1120
rect 2074 -1186 2108 -1120
rect 2266 -1186 2300 -1120
rect 1576 -1232 1582 -1226
rect 1752 -1232 1758 -1226
rect 1792 -1232 1798 -1226
rect 664 -1306 698 -1252
rect 768 -1306 830 -1300
rect 576 -1340 784 -1306
rect 818 -1340 830 -1306
rect 576 -1600 610 -1340
rect 768 -1346 830 -1340
rect 864 -1452 898 -1254
rect 976 -1294 1010 -1255
rect 1168 -1294 1202 -1255
rect 976 -1322 1202 -1294
rect 976 -1356 1010 -1322
rect 976 -1362 1040 -1356
rect 976 -1414 982 -1362
rect 1034 -1414 1040 -1362
rect 976 -1420 1040 -1414
rect 1252 -1408 1310 -1402
rect 1376 -1408 1410 -1254
rect 1532 -1260 1616 -1232
rect 1752 -1260 1840 -1232
rect 640 -1458 704 -1456
rect 638 -1462 704 -1458
rect 638 -1512 646 -1462
rect 640 -1514 646 -1512
rect 698 -1514 704 -1462
rect 640 -1520 704 -1514
rect 864 -1458 930 -1452
rect 864 -1510 872 -1458
rect 924 -1510 930 -1458
rect 864 -1516 930 -1510
rect 976 -1496 1010 -1420
rect 1252 -1442 1264 -1408
rect 1298 -1442 1410 -1408
rect 1252 -1448 1310 -1442
rect 864 -1560 898 -1516
rect 976 -1524 1202 -1496
rect 976 -1566 1010 -1524
rect 1168 -1564 1202 -1524
rect 1376 -1597 1410 -1442
rect 1444 -1408 1502 -1402
rect 1532 -1404 1566 -1260
rect 1596 -1294 1660 -1288
rect 1596 -1346 1602 -1294
rect 1654 -1346 1660 -1294
rect 1596 -1352 1660 -1346
rect 1714 -1294 1778 -1288
rect 1714 -1346 1720 -1294
rect 1772 -1346 1778 -1294
rect 1714 -1352 1778 -1346
rect 1720 -1404 1778 -1398
rect 1532 -1408 1732 -1404
rect 1444 -1442 1456 -1408
rect 1490 -1438 1732 -1408
rect 1766 -1438 1778 -1404
rect 1490 -1442 1566 -1438
rect 1444 -1448 1502 -1442
rect 1532 -1552 1566 -1442
rect 1720 -1444 1778 -1438
rect 1806 -1408 1840 -1260
rect 1876 -1408 1934 -1402
rect 1806 -1442 1888 -1408
rect 1922 -1442 1934 -1408
rect 1596 -1472 1654 -1466
rect 1806 -1472 1840 -1442
rect 1876 -1448 1934 -1442
rect 1962 -1408 1996 -1254
rect 2170 -1294 2204 -1266
rect 2362 -1294 2396 -1254
rect 2170 -1328 2396 -1294
rect 2064 -1408 2122 -1402
rect 1962 -1442 2076 -1408
rect 2110 -1442 2122 -1408
rect 1596 -1506 1608 -1472
rect 1642 -1506 1840 -1472
rect 1596 -1512 1654 -1506
rect 1806 -1552 1840 -1506
rect 1532 -1586 1616 -1552
rect 1752 -1586 1840 -1552
rect 1962 -1597 1996 -1442
rect 2064 -1448 2122 -1442
rect 2362 -1490 2396 -1328
rect 2170 -1524 2396 -1490
rect 2170 -1558 2204 -1524
rect 2362 -1609 2396 -1524
rect 482 -1758 546 -1752
rect 482 -1810 488 -1758
rect 540 -1810 546 -1758
rect 776 -1776 810 -1705
rect 1072 -1776 1106 -1642
rect 1264 -1776 1298 -1642
rect 1464 -1776 1498 -1705
rect 1670 -1776 1704 -1660
rect 1874 -1776 1908 -1709
rect 2074 -1776 2108 -1709
rect 2266 -1776 2300 -1709
rect 482 -1816 546 -1810
rect 758 -1780 2440 -1776
rect 758 -1782 948 -1780
rect 758 -1834 808 -1782
rect 860 -1832 948 -1782
rect 1000 -1832 1104 -1780
rect 1156 -1832 1260 -1780
rect 1312 -1832 1420 -1780
rect 1472 -1832 1572 -1780
rect 1624 -1832 1726 -1780
rect 1778 -1832 1884 -1780
rect 1936 -1782 2194 -1780
rect 1936 -1832 2036 -1782
rect 860 -1834 2036 -1832
rect 2088 -1832 2194 -1782
rect 2246 -1832 2348 -1780
rect 2400 -1832 2440 -1780
rect 2088 -1834 2440 -1832
rect 758 -1840 2440 -1834
<< via1 >>
rect 794 412 846 422
rect 794 378 802 412
rect 802 378 836 412
rect 836 378 846 412
rect 794 370 846 378
rect 952 412 1004 422
rect 952 378 958 412
rect 958 378 992 412
rect 992 378 1004 412
rect 952 370 1004 378
rect 1104 412 1156 424
rect 1104 378 1114 412
rect 1114 378 1148 412
rect 1148 378 1156 412
rect 1104 372 1156 378
rect 1264 412 1316 424
rect 1264 378 1270 412
rect 1270 378 1304 412
rect 1304 378 1316 412
rect 1264 372 1316 378
rect 1418 412 1470 424
rect 1418 378 1426 412
rect 1426 378 1460 412
rect 1460 378 1470 412
rect 1418 372 1470 378
rect 1574 412 1626 422
rect 1574 378 1582 412
rect 1582 378 1616 412
rect 1616 378 1626 412
rect 1574 370 1626 378
rect 1728 412 1780 422
rect 1728 378 1738 412
rect 1738 378 1772 412
rect 1772 378 1780 412
rect 1728 370 1780 378
rect 1886 412 1938 422
rect 1886 378 1894 412
rect 1894 378 1928 412
rect 1928 378 1938 412
rect 1886 370 1938 378
rect 2040 412 2092 422
rect 2040 378 2050 412
rect 2050 378 2084 412
rect 2084 378 2092 412
rect 2040 370 2092 378
rect 2200 412 2252 424
rect 2200 378 2206 412
rect 2206 378 2240 412
rect 2240 378 2252 412
rect 2200 372 2252 378
rect 2354 412 2406 422
rect 2354 378 2362 412
rect 2362 378 2396 412
rect 2396 378 2406 412
rect 2354 370 2406 378
rect 2510 412 2562 422
rect 2510 378 2518 412
rect 2518 378 2552 412
rect 2552 378 2562 412
rect 2510 370 2562 378
rect 1050 8 1102 16
rect 1050 -26 1060 8
rect 1060 -26 1094 8
rect 1094 -26 1102 8
rect 1050 -36 1102 -26
rect 814 -124 866 -72
rect 1270 -38 1322 -28
rect 1270 -72 1278 -38
rect 1278 -72 1312 -38
rect 1312 -72 1322 -38
rect 1270 -80 1322 -72
rect 860 -336 912 -330
rect 860 -370 868 -336
rect 868 -370 902 -336
rect 902 -370 912 -336
rect 860 -382 912 -370
rect 578 -442 630 -390
rect 1440 62 1492 70
rect 1440 28 1448 62
rect 1448 28 1482 62
rect 1482 28 1492 62
rect 1440 18 1492 28
rect 1492 -50 1544 -40
rect 1492 -84 1504 -50
rect 1504 -84 1538 -50
rect 1538 -84 1544 -50
rect 1492 -92 1544 -84
rect 1656 22 1708 74
rect 1584 -144 1636 -92
rect 1874 62 1926 70
rect 1874 28 1884 62
rect 1884 28 1918 62
rect 1918 28 1926 62
rect 1874 18 1926 28
rect 1732 -76 1784 -24
rect 1824 -106 1876 -92
rect 1824 -140 1830 -106
rect 1830 -140 1864 -106
rect 1864 -140 1876 -106
rect 1824 -144 1876 -140
rect 1656 -272 1708 -220
rect 1656 -398 1708 -388
rect 1656 -432 1666 -398
rect 1666 -432 1700 -398
rect 1700 -432 1708 -398
rect 1656 -440 1708 -432
rect 2544 48 2596 100
rect 2262 8 2314 16
rect 2262 -26 2272 8
rect 2272 -26 2306 8
rect 2306 -26 2314 8
rect 2042 -102 2094 -92
rect 2042 -136 2052 -102
rect 2052 -136 2086 -102
rect 2086 -136 2094 -102
rect 2042 -144 2094 -136
rect 2262 -36 2314 -26
rect 2460 -336 2512 -330
rect 2460 -370 2470 -336
rect 2470 -370 2504 -336
rect 2504 -370 2512 -336
rect 2460 -382 2512 -370
rect 2730 -442 2782 -390
rect 860 -836 912 -818
rect 2460 -836 2512 -818
rect 860 -870 868 -836
rect 868 -870 902 -836
rect 902 -870 912 -836
rect 2460 -870 2468 -836
rect 2468 -870 2502 -836
rect 2502 -870 2512 -836
rect 2676 -1010 2786 -900
rect 982 -1414 1034 -1362
rect 646 -1472 698 -1462
rect 646 -1506 654 -1472
rect 654 -1506 688 -1472
rect 688 -1506 698 -1472
rect 646 -1514 698 -1506
rect 872 -1510 924 -1458
rect 1602 -1300 1654 -1294
rect 1602 -1334 1608 -1300
rect 1608 -1334 1642 -1300
rect 1642 -1334 1654 -1300
rect 1602 -1346 1654 -1334
rect 1720 -1300 1772 -1294
rect 1720 -1334 1732 -1300
rect 1732 -1334 1766 -1300
rect 1766 -1334 1772 -1300
rect 1720 -1346 1772 -1334
rect 488 -1768 540 -1758
rect 488 -1802 498 -1768
rect 498 -1802 532 -1768
rect 532 -1802 540 -1768
rect 488 -1810 540 -1802
rect 808 -1792 860 -1782
rect 808 -1826 818 -1792
rect 818 -1826 852 -1792
rect 852 -1826 860 -1792
rect 808 -1834 860 -1826
rect 948 -1792 1000 -1780
rect 948 -1826 958 -1792
rect 958 -1826 992 -1792
rect 992 -1826 1000 -1792
rect 948 -1832 1000 -1826
rect 1104 -1792 1156 -1780
rect 1104 -1826 1114 -1792
rect 1114 -1826 1148 -1792
rect 1148 -1826 1156 -1792
rect 1104 -1832 1156 -1826
rect 1260 -1792 1312 -1780
rect 1260 -1826 1270 -1792
rect 1270 -1826 1304 -1792
rect 1304 -1826 1312 -1792
rect 1260 -1832 1312 -1826
rect 1420 -1792 1472 -1780
rect 1420 -1826 1426 -1792
rect 1426 -1826 1460 -1792
rect 1460 -1826 1472 -1792
rect 1420 -1832 1472 -1826
rect 1572 -1792 1624 -1780
rect 1572 -1826 1582 -1792
rect 1582 -1826 1616 -1792
rect 1616 -1826 1624 -1792
rect 1572 -1832 1624 -1826
rect 1726 -1792 1778 -1780
rect 1726 -1826 1738 -1792
rect 1738 -1826 1772 -1792
rect 1772 -1826 1778 -1792
rect 1726 -1832 1778 -1826
rect 1884 -1792 1936 -1780
rect 1884 -1826 1894 -1792
rect 1894 -1826 1928 -1792
rect 1928 -1826 1936 -1792
rect 1884 -1832 1936 -1826
rect 2036 -1792 2088 -1782
rect 2036 -1826 2050 -1792
rect 2050 -1826 2084 -1792
rect 2084 -1826 2088 -1792
rect 2036 -1834 2088 -1826
rect 2194 -1792 2246 -1780
rect 2194 -1826 2206 -1792
rect 2206 -1826 2240 -1792
rect 2240 -1826 2246 -1792
rect 2194 -1832 2246 -1826
rect 2348 -1792 2400 -1780
rect 2348 -1826 2362 -1792
rect 2362 -1826 2396 -1792
rect 2396 -1826 2400 -1792
rect 2348 -1832 2400 -1826
<< metal2 >>
rect 762 428 2624 482
rect 762 426 1104 428
rect 762 370 794 426
rect 850 370 952 426
rect 1008 372 1104 426
rect 1160 372 1264 428
rect 1320 372 1418 428
rect 1474 426 2200 428
rect 1474 372 1574 426
rect 1008 370 1574 372
rect 1630 370 1728 426
rect 1784 370 1886 426
rect 1942 370 2040 426
rect 2096 372 2200 426
rect 2256 426 2624 428
rect 2256 372 2354 426
rect 2096 370 2354 372
rect 2410 370 2510 426
rect 2566 370 2624 426
rect 762 364 2624 370
rect 488 100 564 110
rect 488 44 498 100
rect 554 44 564 100
rect 488 34 564 44
rect 488 -1752 516 34
rect 670 -60 698 112
rect 2532 102 2608 112
rect 1434 70 1498 76
rect 1044 16 1108 22
rect 1044 -36 1050 16
rect 1102 -36 1108 16
rect 1434 18 1440 70
rect 1492 62 1498 70
rect 1650 74 1714 80
rect 1650 62 1656 74
rect 1492 28 1656 62
rect 1492 18 1498 28
rect 1434 12 1498 18
rect 1650 22 1656 28
rect 1708 62 1714 74
rect 1868 70 1932 76
rect 1868 62 1874 70
rect 1708 28 1874 62
rect 1708 22 1714 28
rect 1650 16 1714 22
rect 1868 18 1874 28
rect 1926 18 1932 70
rect 2532 46 2542 102
rect 2598 46 2608 102
rect 2532 36 2608 46
rect 1868 12 1932 18
rect 2256 16 2320 22
rect 1044 -42 1108 -36
rect 1264 -24 1486 -22
rect 1726 -24 1790 -18
rect 1264 -28 1732 -24
rect 658 -70 734 -60
rect 658 -126 668 -70
rect 724 -126 734 -70
rect 658 -136 734 -126
rect 802 -70 878 -60
rect 802 -126 812 -70
rect 868 -126 878 -70
rect 802 -136 878 -126
rect 566 -382 642 -372
rect 566 -438 576 -382
rect 632 -438 642 -382
rect 566 -442 578 -438
rect 630 -442 642 -438
rect 566 -448 642 -442
rect 572 -764 600 -448
rect 670 -1456 698 -136
rect 854 -330 918 -324
rect 854 -382 860 -330
rect 912 -382 918 -330
rect 854 -388 918 -382
rect 854 -812 882 -388
rect 854 -818 918 -812
rect 854 -870 860 -818
rect 912 -870 918 -818
rect 854 -876 918 -870
rect 1066 -982 1094 -42
rect 1264 -80 1270 -28
rect 1322 -40 1732 -28
rect 1322 -56 1492 -40
rect 1322 -80 1328 -56
rect 1264 -86 1328 -80
rect 1486 -92 1492 -56
rect 1544 -58 1732 -40
rect 1544 -70 1554 -58
rect 1544 -92 1550 -70
rect 1726 -76 1732 -58
rect 1784 -76 1790 -24
rect 2256 -36 2262 16
rect 2314 -36 2320 16
rect 2256 -42 2320 -36
rect 1726 -82 1790 -76
rect 1486 -98 1550 -92
rect 1578 -92 1642 -86
rect 1578 -144 1584 -92
rect 1636 -116 1642 -92
rect 1818 -92 1882 -86
rect 1818 -116 1824 -92
rect 1636 -144 1824 -116
rect 1876 -116 1882 -92
rect 2036 -92 2100 -86
rect 2036 -116 2042 -92
rect 1876 -144 2042 -116
rect 2094 -144 2100 -92
rect 1578 -150 2100 -144
rect 1646 -216 1722 -206
rect 1646 -272 1656 -216
rect 1712 -272 1722 -216
rect 1646 -282 1722 -272
rect 1650 -388 1714 -382
rect 1650 -440 1656 -388
rect 1708 -440 1714 -388
rect 1650 -446 1714 -440
rect 2272 -982 2300 -42
rect 2744 -206 2772 618
rect 2706 -216 2782 -206
rect 2706 -272 2716 -216
rect 2772 -272 2782 -216
rect 2706 -282 2782 -272
rect 2454 -330 2518 -324
rect 2454 -382 2460 -330
rect 2512 -382 2518 -330
rect 2454 -388 2518 -382
rect 2490 -812 2518 -388
rect 2724 -390 2788 -384
rect 2724 -442 2730 -390
rect 2782 -442 2788 -390
rect 2724 -448 2788 -442
rect 2734 -688 2762 -448
rect 2696 -698 2772 -688
rect 2696 -754 2706 -698
rect 2762 -754 2772 -698
rect 2696 -764 2772 -754
rect 2454 -818 2518 -812
rect 2454 -870 2460 -818
rect 2512 -870 2518 -818
rect 2454 -876 2518 -870
rect 1066 -1012 1622 -982
rect 1594 -1286 1622 -1012
rect 1744 -1012 2300 -982
rect 2660 -894 2802 -884
rect 1594 -1288 1630 -1286
rect 1744 -1288 1772 -1012
rect 2660 -1016 2670 -894
rect 2792 -1016 2802 -894
rect 2660 -1026 2802 -1016
rect 1590 -1294 1660 -1288
rect 1590 -1346 1602 -1294
rect 1654 -1346 1660 -1294
rect 1590 -1352 1660 -1346
rect 1714 -1294 1784 -1288
rect 1714 -1346 1720 -1294
rect 1772 -1346 1784 -1294
rect 1714 -1352 1784 -1346
rect 976 -1362 1040 -1356
rect 976 -1414 982 -1362
rect 1034 -1386 1040 -1362
rect 1034 -1414 3788 -1386
rect 976 -1420 1040 -1414
rect 640 -1462 704 -1456
rect 640 -1514 646 -1462
rect 698 -1514 704 -1462
rect 640 -1520 704 -1514
rect 866 -1458 930 -1452
rect 866 -1510 872 -1458
rect 924 -1486 3788 -1458
rect 924 -1510 930 -1486
rect 866 -1516 930 -1510
rect 482 -1758 546 -1752
rect 482 -1810 488 -1758
rect 540 -1810 546 -1758
rect 482 -1816 546 -1810
rect 670 -1816 698 -1520
rect 758 -1780 2440 -1776
rect 758 -1782 948 -1780
rect 758 -1784 808 -1782
rect 860 -1784 948 -1782
rect 1000 -1784 1104 -1780
rect 1156 -1784 1260 -1780
rect 1312 -1784 1420 -1780
rect 1472 -1784 1572 -1780
rect 1624 -1784 1726 -1780
rect 1778 -1784 1884 -1780
rect 1936 -1782 2194 -1780
rect 1936 -1784 2036 -1782
rect 2088 -1784 2194 -1782
rect 2246 -1784 2348 -1780
rect 2400 -1784 2440 -1780
rect 758 -1840 806 -1784
rect 862 -1840 948 -1784
rect 1004 -1840 1104 -1784
rect 1160 -1840 1260 -1784
rect 1316 -1840 1420 -1784
rect 1476 -1840 1572 -1784
rect 1628 -1840 1726 -1784
rect 1782 -1840 1884 -1784
rect 1940 -1840 2036 -1784
rect 2092 -1840 2194 -1784
rect 2250 -1840 2348 -1784
rect 2404 -1840 2440 -1784
rect 758 -1892 2440 -1840
<< via2 >>
rect 794 422 850 426
rect 794 370 846 422
rect 846 370 850 422
rect 952 422 1008 426
rect 952 370 1004 422
rect 1004 370 1008 422
rect 1104 424 1160 428
rect 1104 372 1156 424
rect 1156 372 1160 424
rect 1264 424 1320 428
rect 1264 372 1316 424
rect 1316 372 1320 424
rect 1418 424 1474 428
rect 1418 372 1470 424
rect 1470 372 1474 424
rect 1574 422 1630 426
rect 1574 370 1626 422
rect 1626 370 1630 422
rect 1728 422 1784 426
rect 1728 370 1780 422
rect 1780 370 1784 422
rect 1886 422 1942 426
rect 1886 370 1938 422
rect 1938 370 1942 422
rect 2040 422 2096 426
rect 2040 370 2092 422
rect 2092 370 2096 422
rect 2200 424 2256 428
rect 2200 372 2252 424
rect 2252 372 2256 424
rect 2354 422 2410 426
rect 2354 370 2406 422
rect 2406 370 2410 422
rect 2510 422 2566 426
rect 2510 370 2562 422
rect 2562 370 2566 422
rect 498 44 554 100
rect 2542 100 2598 102
rect 2542 48 2544 100
rect 2544 48 2596 100
rect 2596 48 2598 100
rect 2542 46 2598 48
rect 668 -126 724 -70
rect 812 -72 868 -70
rect 812 -124 814 -72
rect 814 -124 866 -72
rect 866 -124 868 -72
rect 812 -126 868 -124
rect 576 -390 632 -382
rect 576 -438 578 -390
rect 578 -438 630 -390
rect 630 -438 632 -390
rect 1656 -220 1712 -216
rect 1656 -272 1708 -220
rect 1708 -272 1712 -220
rect 2716 -272 2772 -216
rect 2706 -754 2762 -698
rect 2670 -900 2792 -894
rect 2670 -1010 2676 -900
rect 2676 -1010 2786 -900
rect 2786 -1010 2792 -900
rect 2670 -1016 2792 -1010
rect 806 -1834 808 -1784
rect 808 -1834 860 -1784
rect 860 -1834 862 -1784
rect 806 -1840 862 -1834
rect 948 -1832 1000 -1784
rect 1000 -1832 1004 -1784
rect 948 -1840 1004 -1832
rect 1104 -1832 1156 -1784
rect 1156 -1832 1160 -1784
rect 1104 -1840 1160 -1832
rect 1260 -1832 1312 -1784
rect 1312 -1832 1316 -1784
rect 1260 -1840 1316 -1832
rect 1420 -1832 1472 -1784
rect 1472 -1832 1476 -1784
rect 1420 -1840 1476 -1832
rect 1572 -1832 1624 -1784
rect 1624 -1832 1628 -1784
rect 1572 -1840 1628 -1832
rect 1726 -1832 1778 -1784
rect 1778 -1832 1782 -1784
rect 1726 -1840 1782 -1832
rect 1884 -1832 1936 -1784
rect 1936 -1832 1940 -1784
rect 1884 -1840 1940 -1832
rect 2036 -1834 2088 -1784
rect 2088 -1834 2092 -1784
rect 2036 -1840 2092 -1834
rect 2194 -1832 2246 -1784
rect 2246 -1832 2250 -1784
rect 2194 -1840 2250 -1832
rect 2348 -1832 2400 -1784
rect 2400 -1832 2404 -1784
rect 2348 -1840 2404 -1832
<< metal3 >>
rect 762 478 3612 482
rect 762 428 3336 478
rect 762 426 1104 428
rect 762 370 794 426
rect 850 370 952 426
rect 1008 372 1104 426
rect 1160 372 1264 428
rect 1320 372 1418 428
rect 1474 426 2200 428
rect 1474 372 1574 426
rect 1008 370 1574 372
rect 1630 370 1728 426
rect 1784 370 1886 426
rect 1942 370 2040 426
rect 2096 372 2200 426
rect 2256 426 3336 428
rect 2256 372 2354 426
rect 2096 370 2354 372
rect 2410 370 2510 426
rect 2566 370 3336 426
rect 762 368 3336 370
rect 3602 368 3612 478
rect 762 364 3612 368
rect 488 104 564 110
rect 2532 104 2608 112
rect 488 102 2608 104
rect 488 100 2542 102
rect 488 44 498 100
rect 554 46 2542 100
rect 2598 46 2608 102
rect 554 44 2608 46
rect 488 34 564 44
rect 2532 36 2608 44
rect 658 -66 734 -60
rect 802 -66 878 -60
rect 488 -70 2608 -66
rect 488 -126 668 -70
rect 724 -126 812 -70
rect 868 -126 2608 -70
rect 658 -136 734 -126
rect 802 -136 878 -126
rect 1646 -214 1722 -206
rect 2706 -214 2782 -206
rect 1646 -216 2782 -214
rect 1646 -272 1656 -216
rect 1712 -272 2716 -216
rect 2772 -272 2782 -216
rect 1646 -274 2782 -272
rect 1646 -282 1722 -274
rect 2706 -282 2782 -274
rect 566 -380 642 -372
rect 338 -382 2790 -380
rect 338 -438 576 -382
rect 632 -438 2790 -382
rect 338 -440 2790 -438
rect 566 -448 642 -440
rect 2696 -698 2772 -688
rect 338 -754 2706 -698
rect 2762 -754 2772 -698
rect 338 -758 2772 -754
rect 2696 -764 2772 -758
rect 2654 -884 2808 -878
rect 2654 -1026 2660 -884
rect 2802 -1026 2808 -884
rect 2654 -1032 2808 -1026
rect 742 -1778 3612 -1776
rect 742 -1784 3336 -1778
rect 742 -1840 806 -1784
rect 862 -1840 948 -1784
rect 1004 -1840 1104 -1784
rect 1160 -1840 1260 -1784
rect 1316 -1840 1420 -1784
rect 1476 -1840 1572 -1784
rect 1628 -1840 1726 -1784
rect 1782 -1840 1884 -1784
rect 1940 -1840 2036 -1784
rect 2092 -1840 2194 -1784
rect 2250 -1840 2348 -1784
rect 2404 -1840 3336 -1784
rect 742 -1888 3336 -1840
rect 3602 -1888 3612 -1778
rect 742 -1892 3612 -1888
<< via3 >>
rect 3336 368 3602 478
rect 2660 -894 2802 -884
rect 2660 -1016 2670 -894
rect 2670 -1016 2792 -894
rect 2792 -1016 2802 -894
rect 2660 -1026 2802 -1016
rect 3336 -1888 3602 -1778
<< metal4 >>
rect 3326 478 3612 534
rect 2654 -884 2808 -878
rect 2940 -884 3226 444
rect 2654 -1026 2660 -884
rect 2802 -1026 3226 -884
rect 2654 -1032 2808 -1026
rect 2940 -1928 3226 -1026
rect 3326 368 3336 478
rect 3602 368 3612 478
rect 3326 -1778 3612 368
rect 3326 -1888 3336 -1778
rect 3602 -1888 3612 -1778
rect 3326 -1928 3612 -1888
use sky130_fd_pr__nfet_01v8_HNLS5R  XM1
timestamp 1697527592
transform 1 0 1683 0 1 -602
box -221 -126 221 156
use sky130_fd_pr__nfet_01v8_4HESND  XM2
timestamp 1698714739
transform -1 0 995 0 1 -600
box -413 -128 417 188
use sky130_fd_pr__nfet_01v8_4HESND  XM3
timestamp 1698714739
transform 1 0 2371 0 1 -602
box -413 -128 417 188
use sky130_fd_pr__nfet_01v8_648S5X  XM4
timestamp 1697700693
transform 1 0 1551 0 1 -278
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_648S5X  XM5
timestamp 1697700693
transform 1 0 1815 0 1 -278
box -73 -126 73 126
use sky130_fd_pr__pfet_01v8_XGS3BL  XM6
timestamp 1697700693
transform 1 0 1639 0 1 209
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM7
timestamp 1697700693
transform 1 0 1727 0 1 209
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM8
timestamp 1697700693
transform 1 0 1551 0 1 209
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM9
timestamp 1697700693
transform 1 0 1463 0 1 209
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM10
timestamp 1697700693
transform 1 0 1815 0 1 209
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM11
timestamp 1697700693
transform 1 0 1903 0 1 209
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_MQX2PY  XM12
timestamp 1698734556
transform 1 0 2103 0 1 255
box -152 -152 153 232
use sky130_fd_pr__nfet_01v8_EDB9KC  XM13
timestamp 1698718954
transform 1 0 2103 0 1 -220
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_MQP8BZ  XM14
timestamp 1698237672
transform 1 0 2403 0 1 225
box -311 -303 311 303
use sky130_fd_pr__nfet_01v8_PK34ES  XM15
timestamp 1697705701
transform 1 0 2403 0 1 -224
box -173 -72 173 92
use sky130_fd_pr__pfet_01v8_MQX2PY  XM16
timestamp 1698734556
transform -1 0 1731 0 -1 -1667
box -152 -152 153 232
use sky130_fd_pr__pfet_01v8_MQX2PY  XM17
timestamp 1698734556
transform -1 0 1643 0 -1 -1667
box -152 -152 153 232
use sky130_fd_pr__pfet_01v8_MQX2PY  XM18
timestamp 1698734556
transform 1 0 1263 0 1 255
box -152 -152 153 232
use sky130_fd_pr__nfet_01v8_9NW3WL  XM19
timestamp 1697452276
transform -1 0 1643 0 -1 -1176
box -73 -110 73 110
use sky130_fd_pr__nfet_01v8_EDB9KC  XM20
timestamp 1698718954
transform 1 0 1263 0 1 -220
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_MQP8BZ  XM21
timestamp 1698237672
transform -1 0 963 0 1 225
box -311 -303 311 303
use sky130_fd_pr__nfet_01v8_PK34ES  XM22
timestamp 1697705701
transform 1 0 963 0 1 -224
box -173 -72 173 92
use sky130_fd_pr__nfet_01v8_9NW3WL  XM23
timestamp 1697452276
transform -1 0 1731 0 -1 -1176
box -73 -110 73 110
use sky130_fd_pr__pfet_01v8_MQX2PY  XM24
timestamp 1698734556
transform 1 0 637 0 -1 -1667
box -152 -152 153 232
use sky130_fd_pr__pfet_01v8_MQX2PY  XM25
timestamp 1698734556
transform 1 0 549 0 -1 -1667
box -152 -152 153 232
use sky130_fd_pr__nfet_01v8_9NW3WL  XM26
timestamp 1697452276
transform 1 0 637 0 -1 -1182
box -73 -110 73 110
use sky130_fd_pr__nfet_01v8_9NW3WL  XM27
timestamp 1697452276
transform 1 0 549 0 -1 -1182
box -73 -110 73 110
use sky130_fd_pr__pfet_01v8_MQX2PY  XM28
timestamp 1698734556
transform 1 0 837 0 -1 -1663
box -152 -152 153 232
use sky130_fd_pr__nfet_01v8_EDB9KC  XM29
timestamp 1698718954
transform 1 0 837 0 -1 -1222
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_MQX2PY  XM30
timestamp 1698734556
transform -1 0 1437 0 -1 -1663
box -152 -152 153 232
use sky130_fd_pr__nfet_01v8_EDB9KC  XM31
timestamp 1698718954
transform 1 0 1935 0 -1 -1224
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_MQP8BZ  XM32
timestamp 1698237672
transform -1 0 1137 0 -1 -1637
box -311 -303 311 303
use sky130_fd_pr__nfet_01v8_PK34ES  XM33
timestamp 1697705701
transform -1 0 1137 0 -1 -1220
box -173 -72 173 92
use sky130_fd_pr__pfet_01v8_MQX2PY  XM34
timestamp 1698734556
transform 1 0 1935 0 -1 -1667
box -152 -152 153 232
use sky130_fd_pr__nfet_01v8_EDB9KC  XM35
timestamp 1698718954
transform 1 0 1437 0 -1 -1224
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_MQP8BZ  XM36
timestamp 1698237672
transform 1 0 2235 0 -1 -1637
box -311 -303 311 303
use sky130_fd_pr__nfet_01v8_PK34ES  XM37
timestamp 1697705701
transform 1 0 2235 0 -1 -1220
box -173 -72 173 92
<< labels >>
flabel space 1202 -220 1236 153 0 FreeSans 240 0 0 0 Y_inv
flabel space 802 -72 836 153 0 FreeSans 240 0 0 0 Y_drive
flabel metal1 1806 -1586 1840 -1232 0 FreeSans 240 0 0 0 RS_n
flabel metal1 1532 -1586 1566 -1232 0 FreeSans 240 0 0 0 RS_p
flabel space 1578 -92 1612 121 0 FreeSans 288 0 0 0 X
flabel space 1754 -24 1788 121 0 FreeSans 288 0 0 0 Y
flabel space 2530 -190 2564 48 0 FreeSans 288 0 0 0 X_drive
flabel metal4 2940 -1928 3226 444 0 FreeSans 800 0 0 0 VSS
port 15 nsew
flabel metal4 3326 -1928 3612 534 0 FreeSans 800 0 0 0 VDD
port 16 nsew
flabel metal3 338 -758 408 -698 0 FreeSans 240 0 0 0 cdac_vn
port 20 nsew
flabel metal1 2362 -1609 2396 -1254 0 FreeSans 240 0 0 0 comp_outn
port 21 nsew
flabel metal2 3662 -1486 3788 -1458 0 FreeSans 160 0 0 0 ready
port 22 nsew
flabel metal2 3662 -1414 3788 -1386 0 FreeSans 160 0 0 0 comp_outp
port 25 nsew
flabel metal2 2744 536 2772 618 0 FreeSans 160 0 0 0 clk
port 26 nsew
flabel metal1 690 -446 1524 -418 0 FreeSans 160 0 0 0 P
flabel metal3 338 -440 408 -380 0 FreeSans 240 0 0 0 cdac_vp
port 19 nsew
flabel metal1 1842 -446 2676 -418 0 FreeSans 160 0 0 0 Q
<< end >>
