magic
tech sky130A
magscale 1 2
timestamp 1697348449
<< error_p >>
rect -29 379 29 385
rect -29 345 -17 379
rect -29 339 29 345
rect -29 -345 29 -339
rect -29 -379 -17 -345
rect -29 -385 29 -379
<< nwell >>
rect -211 -517 211 517
<< pmos >>
rect -15 -298 15 298
<< pdiff >>
rect -73 286 -15 298
rect -73 -286 -61 286
rect -27 -286 -15 286
rect -73 -298 -15 -286
rect 15 286 73 298
rect 15 -286 27 286
rect 61 -286 73 286
rect 15 -298 73 -286
<< pdiffc >>
rect -61 -286 -27 286
rect 27 -286 61 286
<< nsubdiff >>
rect -175 447 -79 481
rect 79 447 175 481
rect -175 385 -141 447
rect 141 385 175 447
rect -175 -447 -141 -385
rect 141 -447 175 -385
rect -175 -481 -79 -447
rect 79 -481 175 -447
<< nsubdiffcont >>
rect -79 447 79 481
rect -175 -385 -141 385
rect 141 -385 175 385
rect -79 -481 79 -447
<< poly >>
rect -33 379 33 395
rect -33 345 -17 379
rect 17 345 33 379
rect -33 329 33 345
rect -15 298 15 329
rect -15 -329 15 -298
rect -33 -345 33 -329
rect -33 -379 -17 -345
rect 17 -379 33 -345
rect -33 -395 33 -379
<< polycont >>
rect -17 345 17 379
rect -17 -379 17 -345
<< locali >>
rect -175 447 -79 481
rect 79 447 175 481
rect -175 385 -141 447
rect 141 385 175 447
rect -33 345 -17 379
rect 17 345 33 379
rect -61 286 -27 302
rect -61 -302 -27 -286
rect 27 286 61 302
rect 27 -302 61 -286
rect -33 -379 -17 -345
rect 17 -379 33 -345
rect -175 -447 -141 -385
rect 141 -447 175 -385
rect -175 -481 -79 -447
rect 79 -481 175 -447
<< viali >>
rect -17 345 17 379
rect -61 -286 -27 286
rect 27 -286 61 286
rect -17 -379 17 -345
<< metal1 >>
rect -29 379 29 385
rect -29 345 -17 379
rect 17 345 29 379
rect -29 339 29 345
rect -67 286 -21 298
rect -67 -286 -61 286
rect -27 -286 -21 286
rect -67 -298 -21 -286
rect 21 286 67 298
rect 21 -286 27 286
rect 61 -286 67 286
rect 21 -298 67 -286
rect -29 -345 29 -339
rect -29 -379 -17 -345
rect 17 -379 29 -345
rect -29 -385 29 -379
<< properties >>
string FIXED_BBOX -158 -464 158 464
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.98 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
