magic
tech sky130A
timestamp 1698026957
use hgu_cdac_unit  x1
timestamp 1698026957
transform 1 0 376 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x2[0]
timestamp 1698026957
transform 1 0 1478 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x2[1]
timestamp 1698026957
transform 1 0 739 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x3[0]
timestamp 1698026957
transform 1 0 4434 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x3[1]
timestamp 1698026957
transform 1 0 3695 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x3[2]
timestamp 1698026957
transform 1 0 2956 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x3[3]
timestamp 1698026957
transform 1 0 2217 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x4[0]
timestamp 1698026957
transform 1 0 10346 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x4[1]
timestamp 1698026957
transform 1 0 9607 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x4[2]
timestamp 1698026957
transform 1 0 8868 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x4[3]
timestamp 1698026957
transform 1 0 8129 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x4[4]
timestamp 1698026957
transform 1 0 7390 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x4[5]
timestamp 1698026957
transform 1 0 6651 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x4[6]
timestamp 1698026957
transform 1 0 5912 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x4[7]
timestamp 1698026957
transform 1 0 5173 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x5[0]
timestamp 1698026957
transform 1 0 22170 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x5[1]
timestamp 1698026957
transform 1 0 21431 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x5[2]
timestamp 1698026957
transform 1 0 20692 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x5[3]
timestamp 1698026957
transform 1 0 19953 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x5[4]
timestamp 1698026957
transform 1 0 19214 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x5[5]
timestamp 1698026957
transform 1 0 18475 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x5[6]
timestamp 1698026957
transform 1 0 17736 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x5[7]
timestamp 1698026957
transform 1 0 16997 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x5[8]
timestamp 1698026957
transform 1 0 16258 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x5[9]
timestamp 1698026957
transform 1 0 15519 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x5[10]
timestamp 1698026957
transform 1 0 14780 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x5[11]
timestamp 1698026957
transform 1 0 14041 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x5[12]
timestamp 1698026957
transform 1 0 13302 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x5[13]
timestamp 1698026957
transform 1 0 12563 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x5[14]
timestamp 1698026957
transform 1 0 11824 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x5[15]
timestamp 1698026957
transform 1 0 11085 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[0]
timestamp 1698026957
transform 1 0 45818 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[1]
timestamp 1698026957
transform 1 0 45079 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[2]
timestamp 1698026957
transform 1 0 44340 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[3]
timestamp 1698026957
transform 1 0 43601 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[4]
timestamp 1698026957
transform 1 0 42862 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[5]
timestamp 1698026957
transform 1 0 42123 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[6]
timestamp 1698026957
transform 1 0 41384 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[7]
timestamp 1698026957
transform 1 0 40645 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[8]
timestamp 1698026957
transform 1 0 39906 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[9]
timestamp 1698026957
transform 1 0 39167 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[10]
timestamp 1698026957
transform 1 0 38428 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[11]
timestamp 1698026957
transform 1 0 37689 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[12]
timestamp 1698026957
transform 1 0 36950 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[13]
timestamp 1698026957
transform 1 0 36211 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[14]
timestamp 1698026957
transform 1 0 35472 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[15]
timestamp 1698026957
transform 1 0 34733 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[16]
timestamp 1698026957
transform 1 0 33994 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[17]
timestamp 1698026957
transform 1 0 33255 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[18]
timestamp 1698026957
transform 1 0 32516 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[19]
timestamp 1698026957
transform 1 0 31777 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[20]
timestamp 1698026957
transform 1 0 31038 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[21]
timestamp 1698026957
transform 1 0 30299 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[22]
timestamp 1698026957
transform 1 0 29560 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[23]
timestamp 1698026957
transform 1 0 28821 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[24]
timestamp 1698026957
transform 1 0 28082 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[25]
timestamp 1698026957
transform 1 0 27343 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[26]
timestamp 1698026957
transform 1 0 26604 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[27]
timestamp 1698026957
transform 1 0 25865 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[28]
timestamp 1698026957
transform 1 0 25126 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[29]
timestamp 1698026957
transform 1 0 24387 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[30]
timestamp 1698026957
transform 1 0 23648 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x6[31]
timestamp 1698026957
transform 1 0 22909 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[0]
timestamp 1698026957
transform 1 0 93114 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[1]
timestamp 1698026957
transform 1 0 92375 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[2]
timestamp 1698026957
transform 1 0 91636 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[3]
timestamp 1698026957
transform 1 0 90897 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[4]
timestamp 1698026957
transform 1 0 90158 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[5]
timestamp 1698026957
transform 1 0 89419 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[6]
timestamp 1698026957
transform 1 0 88680 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[7]
timestamp 1698026957
transform 1 0 87941 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[8]
timestamp 1698026957
transform 1 0 87202 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[9]
timestamp 1698026957
transform 1 0 86463 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[10]
timestamp 1698026957
transform 1 0 85724 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[11]
timestamp 1698026957
transform 1 0 84985 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[12]
timestamp 1698026957
transform 1 0 84246 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[13]
timestamp 1698026957
transform 1 0 83507 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[14]
timestamp 1698026957
transform 1 0 82768 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[15]
timestamp 1698026957
transform 1 0 82029 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[16]
timestamp 1698026957
transform 1 0 81290 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[17]
timestamp 1698026957
transform 1 0 80551 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[18]
timestamp 1698026957
transform 1 0 79812 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[19]
timestamp 1698026957
transform 1 0 79073 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[20]
timestamp 1698026957
transform 1 0 78334 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[21]
timestamp 1698026957
transform 1 0 77595 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[22]
timestamp 1698026957
transform 1 0 76856 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[23]
timestamp 1698026957
transform 1 0 76117 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[24]
timestamp 1698026957
transform 1 0 75378 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[25]
timestamp 1698026957
transform 1 0 74639 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[26]
timestamp 1698026957
transform 1 0 73900 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[27]
timestamp 1698026957
transform 1 0 73161 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[28]
timestamp 1698026957
transform 1 0 72422 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[29]
timestamp 1698026957
transform 1 0 71683 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[30]
timestamp 1698026957
transform 1 0 70944 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[31]
timestamp 1698026957
transform 1 0 70205 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[32]
timestamp 1698026957
transform 1 0 69466 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[33]
timestamp 1698026957
transform 1 0 68727 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[34]
timestamp 1698026957
transform 1 0 67988 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[35]
timestamp 1698026957
transform 1 0 67249 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[36]
timestamp 1698026957
transform 1 0 66510 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[37]
timestamp 1698026957
transform 1 0 65771 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[38]
timestamp 1698026957
transform 1 0 65032 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[39]
timestamp 1698026957
transform 1 0 64293 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[40]
timestamp 1698026957
transform 1 0 63554 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[41]
timestamp 1698026957
transform 1 0 62815 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[42]
timestamp 1698026957
transform 1 0 62076 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[43]
timestamp 1698026957
transform 1 0 61337 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[44]
timestamp 1698026957
transform 1 0 60598 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[45]
timestamp 1698026957
transform 1 0 59859 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[46]
timestamp 1698026957
transform 1 0 59120 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[47]
timestamp 1698026957
transform 1 0 58381 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[48]
timestamp 1698026957
transform 1 0 57642 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[49]
timestamp 1698026957
transform 1 0 56903 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[50]
timestamp 1698026957
transform 1 0 56164 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[51]
timestamp 1698026957
transform 1 0 55425 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[52]
timestamp 1698026957
transform 1 0 54686 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[53]
timestamp 1698026957
transform 1 0 53947 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[54]
timestamp 1698026957
transform 1 0 53208 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[55]
timestamp 1698026957
transform 1 0 52469 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[56]
timestamp 1698026957
transform 1 0 51730 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[57]
timestamp 1698026957
transform 1 0 50991 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[58]
timestamp 1698026957
transform 1 0 50252 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[59]
timestamp 1698026957
transform 1 0 49513 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[60]
timestamp 1698026957
transform 1 0 48774 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[61]
timestamp 1698026957
transform 1 0 48035 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[62]
timestamp 1698026957
transform 1 0 47296 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x7[63]
timestamp 1698026957
transform 1 0 46557 0 1 1100
box 343 298 739 758
<< end >>
