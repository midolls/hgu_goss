magic
tech sky130A
magscale 1 2
timestamp 1698622076
<< pwell >>
rect 19408 -940 19434 -908
rect 20014 -940 20040 -908
rect 20620 -940 20646 -908
rect 21226 -940 21252 -908
rect 21832 -940 21858 -908
rect 22438 -940 22464 -908
rect 23044 -940 23070 -908
rect 23650 -940 23676 -908
rect 24256 -940 24282 -908
rect 24862 -940 24888 -908
rect 25468 -940 25494 -908
rect 26074 -940 26100 -908
rect 26680 -940 26706 -908
rect 27286 -940 27312 -908
rect 27892 -940 27918 -908
rect 28498 -940 28524 -908
rect 23654 -1110 23676 -1070
rect 19408 -2100 19434 -2068
rect 20014 -2100 20040 -2068
rect 20620 -2100 20646 -2068
rect 21226 -2100 21252 -2068
rect 21832 -2100 21858 -2068
rect 22438 -2100 22464 -2068
rect 23044 -2100 23070 -2068
rect 23650 -2100 23676 -2068
rect 24256 -2100 24282 -2068
rect 24862 -2100 24888 -2068
rect 25468 -2100 25494 -2068
rect 26074 -2100 26100 -2068
rect 26680 -2100 26706 -2068
rect 27286 -2100 27312 -2068
rect 27892 -2100 27918 -2068
rect 28498 -2100 28524 -2068
<< metal3 >>
rect 19088 -130 28850 -128
rect 19088 -194 19192 -130
rect 19256 -194 19272 -130
rect 19336 -194 19352 -130
rect 19416 -194 19432 -130
rect 19496 -194 19512 -130
rect 19576 -194 19592 -130
rect 19656 -194 19798 -130
rect 19862 -194 19878 -130
rect 19942 -194 19958 -130
rect 20022 -194 20038 -130
rect 20102 -194 20118 -130
rect 20182 -194 20198 -130
rect 20262 -194 20404 -130
rect 20468 -194 20484 -130
rect 20548 -194 20564 -130
rect 20628 -194 20644 -130
rect 20708 -194 20724 -130
rect 20788 -194 20804 -130
rect 20868 -194 21010 -130
rect 21074 -194 21090 -130
rect 21154 -194 21170 -130
rect 21234 -194 21250 -130
rect 21314 -194 21330 -130
rect 21394 -194 21410 -130
rect 21474 -194 21616 -130
rect 21680 -194 21696 -130
rect 21760 -194 21776 -130
rect 21840 -194 21856 -130
rect 21920 -194 21936 -130
rect 22000 -194 22016 -130
rect 22080 -194 22222 -130
rect 22286 -194 22302 -130
rect 22366 -194 22382 -130
rect 22446 -194 22462 -130
rect 22526 -194 22542 -130
rect 22606 -194 22622 -130
rect 22686 -194 22828 -130
rect 22892 -194 22908 -130
rect 22972 -194 22988 -130
rect 23052 -194 23068 -130
rect 23132 -194 23148 -130
rect 23212 -194 23228 -130
rect 23292 -194 23434 -130
rect 23498 -194 23514 -130
rect 23578 -194 23594 -130
rect 23658 -194 23674 -130
rect 23738 -194 23754 -130
rect 23818 -194 23834 -130
rect 23898 -194 24040 -130
rect 24104 -194 24120 -130
rect 24184 -194 24200 -130
rect 24264 -194 24280 -130
rect 24344 -194 24360 -130
rect 24424 -194 24440 -130
rect 24504 -194 24646 -130
rect 24710 -194 24726 -130
rect 24790 -194 24806 -130
rect 24870 -194 24886 -130
rect 24950 -194 24966 -130
rect 25030 -194 25046 -130
rect 25110 -194 25252 -130
rect 25316 -194 25332 -130
rect 25396 -194 25412 -130
rect 25476 -194 25492 -130
rect 25556 -194 25572 -130
rect 25636 -194 25652 -130
rect 25716 -194 25858 -130
rect 25922 -194 25938 -130
rect 26002 -194 26018 -130
rect 26082 -194 26098 -130
rect 26162 -194 26178 -130
rect 26242 -194 26258 -130
rect 26322 -194 26464 -130
rect 26528 -194 26544 -130
rect 26608 -194 26624 -130
rect 26688 -194 26704 -130
rect 26768 -194 26784 -130
rect 26848 -194 26864 -130
rect 26928 -194 27070 -130
rect 27134 -194 27150 -130
rect 27214 -194 27230 -130
rect 27294 -194 27310 -130
rect 27374 -194 27390 -130
rect 27454 -194 27470 -130
rect 27534 -194 27676 -130
rect 27740 -194 27756 -130
rect 27820 -194 27836 -130
rect 27900 -194 27916 -130
rect 27980 -194 27996 -130
rect 28060 -194 28076 -130
rect 28140 -194 28282 -130
rect 28346 -194 28362 -130
rect 28426 -194 28442 -130
rect 28506 -194 28522 -130
rect 28586 -194 28602 -130
rect 28666 -194 28682 -130
rect 28746 -194 28850 -130
rect 19088 -196 28850 -194
rect 19088 -350 19154 -196
rect 19088 -414 19089 -350
rect 19153 -414 19154 -350
rect 19088 -430 19154 -414
rect 19088 -494 19089 -430
rect 19153 -494 19154 -430
rect 19088 -510 19154 -494
rect 19088 -574 19089 -510
rect 19153 -574 19154 -510
rect 19088 -590 19154 -574
rect 19088 -654 19089 -590
rect 19153 -654 19154 -590
rect 19088 -670 19154 -654
rect 19088 -734 19089 -670
rect 19153 -734 19154 -670
rect 19088 -750 19154 -734
rect 19088 -814 19089 -750
rect 19153 -814 19154 -750
rect 19088 -830 19154 -814
rect 19088 -894 19089 -830
rect 19153 -894 19154 -830
rect 19088 -910 19154 -894
rect 19088 -974 19089 -910
rect 19153 -974 19154 -910
rect 19088 -990 19154 -974
rect 19088 -1054 19089 -990
rect 19153 -1054 19154 -990
rect 19088 -1070 19154 -1054
rect 19088 -1134 19089 -1070
rect 19153 -1134 19154 -1070
rect 19088 -1224 19154 -1134
rect 19214 -1228 19274 -196
rect 19334 -1288 19394 -258
rect 19454 -1228 19514 -196
rect 19574 -1288 19634 -258
rect 19694 -350 19760 -196
rect 19694 -414 19695 -350
rect 19759 -414 19760 -350
rect 19694 -430 19760 -414
rect 19694 -494 19695 -430
rect 19759 -494 19760 -430
rect 19694 -510 19760 -494
rect 19694 -574 19695 -510
rect 19759 -574 19760 -510
rect 19694 -590 19760 -574
rect 19694 -654 19695 -590
rect 19759 -654 19760 -590
rect 19694 -670 19760 -654
rect 19694 -734 19695 -670
rect 19759 -734 19760 -670
rect 19694 -750 19760 -734
rect 19694 -814 19695 -750
rect 19759 -814 19760 -750
rect 19694 -830 19760 -814
rect 19694 -894 19695 -830
rect 19759 -894 19760 -830
rect 19694 -910 19760 -894
rect 19694 -974 19695 -910
rect 19759 -974 19760 -910
rect 19694 -990 19760 -974
rect 19694 -1054 19695 -990
rect 19759 -1054 19760 -990
rect 19694 -1070 19760 -1054
rect 19694 -1134 19695 -1070
rect 19759 -1134 19760 -1070
rect 19694 -1224 19760 -1134
rect 19820 -1228 19880 -196
rect 19940 -1288 20000 -258
rect 20060 -1228 20120 -196
rect 20180 -1288 20240 -258
rect 20300 -350 20366 -196
rect 20300 -414 20301 -350
rect 20365 -414 20366 -350
rect 20300 -430 20366 -414
rect 20300 -494 20301 -430
rect 20365 -494 20366 -430
rect 20300 -510 20366 -494
rect 20300 -574 20301 -510
rect 20365 -574 20366 -510
rect 20300 -590 20366 -574
rect 20300 -654 20301 -590
rect 20365 -654 20366 -590
rect 20300 -670 20366 -654
rect 20300 -734 20301 -670
rect 20365 -734 20366 -670
rect 20300 -750 20366 -734
rect 20300 -814 20301 -750
rect 20365 -814 20366 -750
rect 20300 -830 20366 -814
rect 20300 -894 20301 -830
rect 20365 -894 20366 -830
rect 20300 -910 20366 -894
rect 20300 -974 20301 -910
rect 20365 -974 20366 -910
rect 20300 -990 20366 -974
rect 20300 -1054 20301 -990
rect 20365 -1054 20366 -990
rect 20300 -1070 20366 -1054
rect 20300 -1134 20301 -1070
rect 20365 -1134 20366 -1070
rect 20300 -1224 20366 -1134
rect 20426 -1228 20486 -196
rect 20546 -1288 20606 -258
rect 20666 -1228 20726 -196
rect 20786 -1288 20846 -258
rect 20906 -350 20972 -196
rect 20906 -414 20907 -350
rect 20971 -414 20972 -350
rect 20906 -430 20972 -414
rect 20906 -494 20907 -430
rect 20971 -494 20972 -430
rect 20906 -510 20972 -494
rect 20906 -574 20907 -510
rect 20971 -574 20972 -510
rect 20906 -590 20972 -574
rect 20906 -654 20907 -590
rect 20971 -654 20972 -590
rect 20906 -670 20972 -654
rect 20906 -734 20907 -670
rect 20971 -734 20972 -670
rect 20906 -750 20972 -734
rect 20906 -814 20907 -750
rect 20971 -814 20972 -750
rect 20906 -830 20972 -814
rect 20906 -894 20907 -830
rect 20971 -894 20972 -830
rect 20906 -910 20972 -894
rect 20906 -974 20907 -910
rect 20971 -974 20972 -910
rect 20906 -990 20972 -974
rect 20906 -1054 20907 -990
rect 20971 -1054 20972 -990
rect 20906 -1070 20972 -1054
rect 20906 -1134 20907 -1070
rect 20971 -1134 20972 -1070
rect 20906 -1224 20972 -1134
rect 21032 -1228 21092 -196
rect 21152 -1288 21212 -258
rect 21272 -1228 21332 -196
rect 21392 -1288 21452 -258
rect 21512 -350 21578 -196
rect 21512 -414 21513 -350
rect 21577 -414 21578 -350
rect 21512 -430 21578 -414
rect 21512 -494 21513 -430
rect 21577 -494 21578 -430
rect 21512 -510 21578 -494
rect 21512 -574 21513 -510
rect 21577 -574 21578 -510
rect 21512 -590 21578 -574
rect 21512 -654 21513 -590
rect 21577 -654 21578 -590
rect 21512 -670 21578 -654
rect 21512 -734 21513 -670
rect 21577 -734 21578 -670
rect 21512 -750 21578 -734
rect 21512 -814 21513 -750
rect 21577 -814 21578 -750
rect 21512 -830 21578 -814
rect 21512 -894 21513 -830
rect 21577 -894 21578 -830
rect 21512 -910 21578 -894
rect 21512 -974 21513 -910
rect 21577 -974 21578 -910
rect 21512 -990 21578 -974
rect 21512 -1054 21513 -990
rect 21577 -1054 21578 -990
rect 21512 -1070 21578 -1054
rect 21512 -1134 21513 -1070
rect 21577 -1134 21578 -1070
rect 21512 -1224 21578 -1134
rect 21638 -1228 21698 -196
rect 21758 -1288 21818 -258
rect 21878 -1228 21938 -196
rect 21998 -1288 22058 -258
rect 22118 -350 22184 -196
rect 22118 -414 22119 -350
rect 22183 -414 22184 -350
rect 22118 -430 22184 -414
rect 22118 -494 22119 -430
rect 22183 -494 22184 -430
rect 22118 -510 22184 -494
rect 22118 -574 22119 -510
rect 22183 -574 22184 -510
rect 22118 -590 22184 -574
rect 22118 -654 22119 -590
rect 22183 -654 22184 -590
rect 22118 -670 22184 -654
rect 22118 -734 22119 -670
rect 22183 -734 22184 -670
rect 22118 -750 22184 -734
rect 22118 -814 22119 -750
rect 22183 -814 22184 -750
rect 22118 -830 22184 -814
rect 22118 -894 22119 -830
rect 22183 -894 22184 -830
rect 22118 -910 22184 -894
rect 22118 -974 22119 -910
rect 22183 -974 22184 -910
rect 22118 -990 22184 -974
rect 22118 -1054 22119 -990
rect 22183 -1054 22184 -990
rect 22118 -1070 22184 -1054
rect 22118 -1134 22119 -1070
rect 22183 -1134 22184 -1070
rect 22118 -1224 22184 -1134
rect 22244 -1228 22304 -196
rect 22364 -1288 22424 -258
rect 22484 -1228 22544 -196
rect 22604 -1288 22664 -258
rect 22724 -350 22790 -196
rect 22724 -414 22725 -350
rect 22789 -414 22790 -350
rect 22724 -430 22790 -414
rect 22724 -494 22725 -430
rect 22789 -494 22790 -430
rect 22724 -510 22790 -494
rect 22724 -574 22725 -510
rect 22789 -574 22790 -510
rect 22724 -590 22790 -574
rect 22724 -654 22725 -590
rect 22789 -654 22790 -590
rect 22724 -670 22790 -654
rect 22724 -734 22725 -670
rect 22789 -734 22790 -670
rect 22724 -750 22790 -734
rect 22724 -814 22725 -750
rect 22789 -814 22790 -750
rect 22724 -830 22790 -814
rect 22724 -894 22725 -830
rect 22789 -894 22790 -830
rect 22724 -910 22790 -894
rect 22724 -974 22725 -910
rect 22789 -974 22790 -910
rect 22724 -990 22790 -974
rect 22724 -1054 22725 -990
rect 22789 -1054 22790 -990
rect 22724 -1070 22790 -1054
rect 22724 -1134 22725 -1070
rect 22789 -1134 22790 -1070
rect 22724 -1224 22790 -1134
rect 22850 -1228 22910 -196
rect 22970 -1288 23030 -258
rect 23090 -1228 23150 -196
rect 23210 -1288 23270 -258
rect 23330 -350 23396 -196
rect 23330 -414 23331 -350
rect 23395 -414 23396 -350
rect 23330 -430 23396 -414
rect 23330 -494 23331 -430
rect 23395 -494 23396 -430
rect 23330 -510 23396 -494
rect 23330 -574 23331 -510
rect 23395 -574 23396 -510
rect 23330 -590 23396 -574
rect 23330 -654 23331 -590
rect 23395 -654 23396 -590
rect 23330 -670 23396 -654
rect 23330 -734 23331 -670
rect 23395 -734 23396 -670
rect 23330 -750 23396 -734
rect 23330 -814 23331 -750
rect 23395 -814 23396 -750
rect 23330 -830 23396 -814
rect 23330 -894 23331 -830
rect 23395 -894 23396 -830
rect 23330 -910 23396 -894
rect 23330 -974 23331 -910
rect 23395 -974 23396 -910
rect 23330 -990 23396 -974
rect 23330 -1054 23331 -990
rect 23395 -1054 23396 -990
rect 23330 -1070 23396 -1054
rect 23330 -1134 23331 -1070
rect 23395 -1134 23396 -1070
rect 23330 -1224 23396 -1134
rect 23456 -1228 23516 -196
rect 23576 -1288 23636 -258
rect 23696 -1228 23756 -196
rect 23816 -1288 23876 -258
rect 23936 -350 24002 -196
rect 23936 -414 23937 -350
rect 24001 -414 24002 -350
rect 23936 -430 24002 -414
rect 23936 -494 23937 -430
rect 24001 -494 24002 -430
rect 23936 -510 24002 -494
rect 23936 -574 23937 -510
rect 24001 -574 24002 -510
rect 23936 -590 24002 -574
rect 23936 -654 23937 -590
rect 24001 -654 24002 -590
rect 23936 -670 24002 -654
rect 23936 -734 23937 -670
rect 24001 -734 24002 -670
rect 23936 -750 24002 -734
rect 23936 -814 23937 -750
rect 24001 -814 24002 -750
rect 23936 -830 24002 -814
rect 23936 -894 23937 -830
rect 24001 -894 24002 -830
rect 23936 -910 24002 -894
rect 23936 -974 23937 -910
rect 24001 -974 24002 -910
rect 23936 -990 24002 -974
rect 23936 -1054 23937 -990
rect 24001 -1054 24002 -990
rect 23936 -1070 24002 -1054
rect 23936 -1134 23937 -1070
rect 24001 -1134 24002 -1070
rect 23936 -1224 24002 -1134
rect 24062 -1228 24122 -196
rect 24182 -1288 24242 -258
rect 24302 -1228 24362 -196
rect 24422 -1288 24482 -258
rect 24542 -350 24608 -196
rect 24542 -414 24543 -350
rect 24607 -414 24608 -350
rect 24542 -430 24608 -414
rect 24542 -494 24543 -430
rect 24607 -494 24608 -430
rect 24542 -510 24608 -494
rect 24542 -574 24543 -510
rect 24607 -574 24608 -510
rect 24542 -590 24608 -574
rect 24542 -654 24543 -590
rect 24607 -654 24608 -590
rect 24542 -670 24608 -654
rect 24542 -734 24543 -670
rect 24607 -734 24608 -670
rect 24542 -750 24608 -734
rect 24542 -814 24543 -750
rect 24607 -814 24608 -750
rect 24542 -830 24608 -814
rect 24542 -894 24543 -830
rect 24607 -894 24608 -830
rect 24542 -910 24608 -894
rect 24542 -974 24543 -910
rect 24607 -974 24608 -910
rect 24542 -990 24608 -974
rect 24542 -1054 24543 -990
rect 24607 -1054 24608 -990
rect 24542 -1070 24608 -1054
rect 24542 -1134 24543 -1070
rect 24607 -1134 24608 -1070
rect 24542 -1224 24608 -1134
rect 24668 -1228 24728 -196
rect 24788 -1288 24848 -258
rect 24908 -1228 24968 -196
rect 25028 -1288 25088 -258
rect 25148 -350 25214 -196
rect 25148 -414 25149 -350
rect 25213 -414 25214 -350
rect 25148 -430 25214 -414
rect 25148 -494 25149 -430
rect 25213 -494 25214 -430
rect 25148 -510 25214 -494
rect 25148 -574 25149 -510
rect 25213 -574 25214 -510
rect 25148 -590 25214 -574
rect 25148 -654 25149 -590
rect 25213 -654 25214 -590
rect 25148 -670 25214 -654
rect 25148 -734 25149 -670
rect 25213 -734 25214 -670
rect 25148 -750 25214 -734
rect 25148 -814 25149 -750
rect 25213 -814 25214 -750
rect 25148 -830 25214 -814
rect 25148 -894 25149 -830
rect 25213 -894 25214 -830
rect 25148 -910 25214 -894
rect 25148 -974 25149 -910
rect 25213 -974 25214 -910
rect 25148 -990 25214 -974
rect 25148 -1054 25149 -990
rect 25213 -1054 25214 -990
rect 25148 -1070 25214 -1054
rect 25148 -1134 25149 -1070
rect 25213 -1134 25214 -1070
rect 25148 -1224 25214 -1134
rect 25274 -1228 25334 -196
rect 25394 -1288 25454 -258
rect 25514 -1228 25574 -196
rect 25634 -1288 25694 -258
rect 25754 -350 25820 -196
rect 25754 -414 25755 -350
rect 25819 -414 25820 -350
rect 25754 -430 25820 -414
rect 25754 -494 25755 -430
rect 25819 -494 25820 -430
rect 25754 -510 25820 -494
rect 25754 -574 25755 -510
rect 25819 -574 25820 -510
rect 25754 -590 25820 -574
rect 25754 -654 25755 -590
rect 25819 -654 25820 -590
rect 25754 -670 25820 -654
rect 25754 -734 25755 -670
rect 25819 -734 25820 -670
rect 25754 -750 25820 -734
rect 25754 -814 25755 -750
rect 25819 -814 25820 -750
rect 25754 -830 25820 -814
rect 25754 -894 25755 -830
rect 25819 -894 25820 -830
rect 25754 -910 25820 -894
rect 25754 -974 25755 -910
rect 25819 -974 25820 -910
rect 25754 -990 25820 -974
rect 25754 -1054 25755 -990
rect 25819 -1054 25820 -990
rect 25754 -1070 25820 -1054
rect 25754 -1134 25755 -1070
rect 25819 -1134 25820 -1070
rect 25754 -1224 25820 -1134
rect 25880 -1228 25940 -196
rect 26000 -1288 26060 -258
rect 26120 -1228 26180 -196
rect 26240 -1288 26300 -258
rect 26360 -350 26426 -196
rect 26360 -414 26361 -350
rect 26425 -414 26426 -350
rect 26360 -430 26426 -414
rect 26360 -494 26361 -430
rect 26425 -494 26426 -430
rect 26360 -510 26426 -494
rect 26360 -574 26361 -510
rect 26425 -574 26426 -510
rect 26360 -590 26426 -574
rect 26360 -654 26361 -590
rect 26425 -654 26426 -590
rect 26360 -670 26426 -654
rect 26360 -734 26361 -670
rect 26425 -734 26426 -670
rect 26360 -750 26426 -734
rect 26360 -814 26361 -750
rect 26425 -814 26426 -750
rect 26360 -830 26426 -814
rect 26360 -894 26361 -830
rect 26425 -894 26426 -830
rect 26360 -910 26426 -894
rect 26360 -974 26361 -910
rect 26425 -974 26426 -910
rect 26360 -990 26426 -974
rect 26360 -1054 26361 -990
rect 26425 -1054 26426 -990
rect 26360 -1070 26426 -1054
rect 26360 -1134 26361 -1070
rect 26425 -1134 26426 -1070
rect 26360 -1224 26426 -1134
rect 26486 -1228 26546 -196
rect 26606 -1288 26666 -258
rect 26726 -1228 26786 -196
rect 26846 -1288 26906 -258
rect 26966 -350 27032 -196
rect 26966 -414 26967 -350
rect 27031 -414 27032 -350
rect 26966 -430 27032 -414
rect 26966 -494 26967 -430
rect 27031 -494 27032 -430
rect 26966 -510 27032 -494
rect 26966 -574 26967 -510
rect 27031 -574 27032 -510
rect 26966 -590 27032 -574
rect 26966 -654 26967 -590
rect 27031 -654 27032 -590
rect 26966 -670 27032 -654
rect 26966 -734 26967 -670
rect 27031 -734 27032 -670
rect 26966 -750 27032 -734
rect 26966 -814 26967 -750
rect 27031 -814 27032 -750
rect 26966 -830 27032 -814
rect 26966 -894 26967 -830
rect 27031 -894 27032 -830
rect 26966 -910 27032 -894
rect 26966 -974 26967 -910
rect 27031 -974 27032 -910
rect 26966 -990 27032 -974
rect 26966 -1054 26967 -990
rect 27031 -1054 27032 -990
rect 26966 -1070 27032 -1054
rect 26966 -1134 26967 -1070
rect 27031 -1134 27032 -1070
rect 26966 -1224 27032 -1134
rect 27092 -1228 27152 -196
rect 27212 -1288 27272 -258
rect 27332 -1228 27392 -196
rect 27452 -1288 27512 -258
rect 27572 -350 27638 -196
rect 27572 -414 27573 -350
rect 27637 -414 27638 -350
rect 27572 -430 27638 -414
rect 27572 -494 27573 -430
rect 27637 -494 27638 -430
rect 27572 -510 27638 -494
rect 27572 -574 27573 -510
rect 27637 -574 27638 -510
rect 27572 -590 27638 -574
rect 27572 -654 27573 -590
rect 27637 -654 27638 -590
rect 27572 -670 27638 -654
rect 27572 -734 27573 -670
rect 27637 -734 27638 -670
rect 27572 -750 27638 -734
rect 27572 -814 27573 -750
rect 27637 -814 27638 -750
rect 27572 -830 27638 -814
rect 27572 -894 27573 -830
rect 27637 -894 27638 -830
rect 27572 -910 27638 -894
rect 27572 -974 27573 -910
rect 27637 -974 27638 -910
rect 27572 -990 27638 -974
rect 27572 -1054 27573 -990
rect 27637 -1054 27638 -990
rect 27572 -1070 27638 -1054
rect 27572 -1134 27573 -1070
rect 27637 -1134 27638 -1070
rect 27572 -1224 27638 -1134
rect 27698 -1228 27758 -196
rect 27818 -1288 27878 -258
rect 27938 -1228 27998 -196
rect 28058 -1288 28118 -258
rect 28178 -350 28244 -196
rect 28178 -414 28179 -350
rect 28243 -414 28244 -350
rect 28178 -430 28244 -414
rect 28178 -494 28179 -430
rect 28243 -494 28244 -430
rect 28178 -510 28244 -494
rect 28178 -574 28179 -510
rect 28243 -574 28244 -510
rect 28178 -590 28244 -574
rect 28178 -654 28179 -590
rect 28243 -654 28244 -590
rect 28178 -670 28244 -654
rect 28178 -734 28179 -670
rect 28243 -734 28244 -670
rect 28178 -750 28244 -734
rect 28178 -814 28179 -750
rect 28243 -814 28244 -750
rect 28178 -830 28244 -814
rect 28178 -894 28179 -830
rect 28243 -894 28244 -830
rect 28178 -910 28244 -894
rect 28178 -974 28179 -910
rect 28243 -974 28244 -910
rect 28178 -990 28244 -974
rect 28178 -1054 28179 -990
rect 28243 -1054 28244 -990
rect 28178 -1070 28244 -1054
rect 28178 -1134 28179 -1070
rect 28243 -1134 28244 -1070
rect 28178 -1224 28244 -1134
rect 28304 -1228 28364 -196
rect 28424 -1288 28484 -258
rect 28544 -1228 28604 -196
rect 28664 -1288 28724 -258
rect 28784 -350 28850 -196
rect 28784 -414 28785 -350
rect 28849 -414 28850 -350
rect 28784 -430 28850 -414
rect 28784 -494 28785 -430
rect 28849 -494 28850 -430
rect 28784 -510 28850 -494
rect 28784 -574 28785 -510
rect 28849 -574 28850 -510
rect 28784 -590 28850 -574
rect 28784 -654 28785 -590
rect 28849 -654 28850 -590
rect 28784 -670 28850 -654
rect 28784 -734 28785 -670
rect 28849 -734 28850 -670
rect 28784 -750 28850 -734
rect 28784 -814 28785 -750
rect 28849 -814 28850 -750
rect 28784 -830 28850 -814
rect 28784 -894 28785 -830
rect 28849 -894 28850 -830
rect 28784 -910 28850 -894
rect 28784 -974 28785 -910
rect 28849 -974 28850 -910
rect 28784 -990 28850 -974
rect 28784 -1054 28785 -990
rect 28849 -1054 28850 -990
rect 28784 -1070 28850 -1054
rect 28784 -1134 28785 -1070
rect 28849 -1134 28850 -1070
rect 28784 -1224 28850 -1134
rect 19088 -1290 28850 -1288
rect 19088 -1354 19192 -1290
rect 19256 -1354 19272 -1290
rect 19336 -1354 19352 -1290
rect 19416 -1354 19432 -1290
rect 19496 -1354 19512 -1290
rect 19576 -1354 19592 -1290
rect 19656 -1354 19798 -1290
rect 19862 -1354 19878 -1290
rect 19942 -1354 19958 -1290
rect 20022 -1354 20038 -1290
rect 20102 -1354 20118 -1290
rect 20182 -1354 20198 -1290
rect 20262 -1354 20404 -1290
rect 20468 -1354 20484 -1290
rect 20548 -1354 20564 -1290
rect 20628 -1354 20644 -1290
rect 20708 -1354 20724 -1290
rect 20788 -1354 20804 -1290
rect 20868 -1354 21010 -1290
rect 21074 -1354 21090 -1290
rect 21154 -1354 21170 -1290
rect 21234 -1354 21250 -1290
rect 21314 -1354 21330 -1290
rect 21394 -1354 21410 -1290
rect 21474 -1354 21616 -1290
rect 21680 -1354 21696 -1290
rect 21760 -1354 21776 -1290
rect 21840 -1354 21856 -1290
rect 21920 -1354 21936 -1290
rect 22000 -1354 22016 -1290
rect 22080 -1354 22222 -1290
rect 22286 -1354 22302 -1290
rect 22366 -1354 22382 -1290
rect 22446 -1354 22462 -1290
rect 22526 -1354 22542 -1290
rect 22606 -1354 22622 -1290
rect 22686 -1354 22828 -1290
rect 22892 -1354 22908 -1290
rect 22972 -1354 22988 -1290
rect 23052 -1354 23068 -1290
rect 23132 -1354 23148 -1290
rect 23212 -1354 23228 -1290
rect 23292 -1354 23434 -1290
rect 23498 -1354 23514 -1290
rect 23578 -1354 23594 -1290
rect 23658 -1354 23674 -1290
rect 23738 -1354 23754 -1290
rect 23818 -1354 23834 -1290
rect 23898 -1354 24040 -1290
rect 24104 -1354 24120 -1290
rect 24184 -1354 24200 -1290
rect 24264 -1354 24280 -1290
rect 24344 -1354 24360 -1290
rect 24424 -1354 24440 -1290
rect 24504 -1354 24646 -1290
rect 24710 -1354 24726 -1290
rect 24790 -1354 24806 -1290
rect 24870 -1354 24886 -1290
rect 24950 -1354 24966 -1290
rect 25030 -1354 25046 -1290
rect 25110 -1354 25252 -1290
rect 25316 -1354 25332 -1290
rect 25396 -1354 25412 -1290
rect 25476 -1354 25492 -1290
rect 25556 -1354 25572 -1290
rect 25636 -1354 25652 -1290
rect 25716 -1354 25858 -1290
rect 25922 -1354 25938 -1290
rect 26002 -1354 26018 -1290
rect 26082 -1354 26098 -1290
rect 26162 -1354 26178 -1290
rect 26242 -1354 26258 -1290
rect 26322 -1354 26464 -1290
rect 26528 -1354 26544 -1290
rect 26608 -1354 26624 -1290
rect 26688 -1354 26704 -1290
rect 26768 -1354 26784 -1290
rect 26848 -1354 26864 -1290
rect 26928 -1354 27070 -1290
rect 27134 -1354 27150 -1290
rect 27214 -1354 27230 -1290
rect 27294 -1354 27310 -1290
rect 27374 -1354 27390 -1290
rect 27454 -1354 27470 -1290
rect 27534 -1354 27676 -1290
rect 27740 -1354 27756 -1290
rect 27820 -1354 27836 -1290
rect 27900 -1354 27916 -1290
rect 27980 -1354 27996 -1290
rect 28060 -1354 28076 -1290
rect 28140 -1354 28282 -1290
rect 28346 -1354 28362 -1290
rect 28426 -1354 28442 -1290
rect 28506 -1354 28522 -1290
rect 28586 -1354 28602 -1290
rect 28666 -1354 28682 -1290
rect 28746 -1354 28850 -1290
rect 19088 -1356 28850 -1354
rect 19088 -1510 19154 -1356
rect 19088 -1574 19089 -1510
rect 19153 -1574 19154 -1510
rect 19088 -1590 19154 -1574
rect 19088 -1654 19089 -1590
rect 19153 -1654 19154 -1590
rect 19088 -1670 19154 -1654
rect 19088 -1734 19089 -1670
rect 19153 -1734 19154 -1670
rect 19088 -1750 19154 -1734
rect 19088 -1814 19089 -1750
rect 19153 -1814 19154 -1750
rect 19088 -1830 19154 -1814
rect 19088 -1894 19089 -1830
rect 19153 -1894 19154 -1830
rect 19088 -1910 19154 -1894
rect 19088 -1974 19089 -1910
rect 19153 -1974 19154 -1910
rect 19088 -1990 19154 -1974
rect 19088 -2054 19089 -1990
rect 19153 -2054 19154 -1990
rect 19088 -2070 19154 -2054
rect 19088 -2134 19089 -2070
rect 19153 -2134 19154 -2070
rect 19088 -2150 19154 -2134
rect 19088 -2214 19089 -2150
rect 19153 -2214 19154 -2150
rect 19088 -2230 19154 -2214
rect 19088 -2294 19089 -2230
rect 19153 -2294 19154 -2230
rect 19088 -2384 19154 -2294
rect 19214 -2388 19274 -1356
rect 19334 -2448 19394 -1418
rect 19454 -2388 19514 -1356
rect 19574 -2448 19634 -1418
rect 19694 -1510 19760 -1356
rect 19694 -1574 19695 -1510
rect 19759 -1574 19760 -1510
rect 19694 -1590 19760 -1574
rect 19694 -1654 19695 -1590
rect 19759 -1654 19760 -1590
rect 19694 -1670 19760 -1654
rect 19694 -1734 19695 -1670
rect 19759 -1734 19760 -1670
rect 19694 -1750 19760 -1734
rect 19694 -1814 19695 -1750
rect 19759 -1814 19760 -1750
rect 19694 -1830 19760 -1814
rect 19694 -1894 19695 -1830
rect 19759 -1894 19760 -1830
rect 19694 -1910 19760 -1894
rect 19694 -1974 19695 -1910
rect 19759 -1974 19760 -1910
rect 19694 -1990 19760 -1974
rect 19694 -2054 19695 -1990
rect 19759 -2054 19760 -1990
rect 19694 -2070 19760 -2054
rect 19694 -2134 19695 -2070
rect 19759 -2134 19760 -2070
rect 19694 -2150 19760 -2134
rect 19694 -2214 19695 -2150
rect 19759 -2214 19760 -2150
rect 19694 -2230 19760 -2214
rect 19694 -2294 19695 -2230
rect 19759 -2294 19760 -2230
rect 19694 -2384 19760 -2294
rect 19820 -2388 19880 -1356
rect 19940 -2448 20000 -1418
rect 20060 -2388 20120 -1356
rect 20180 -2448 20240 -1418
rect 20300 -1510 20366 -1356
rect 20300 -1574 20301 -1510
rect 20365 -1574 20366 -1510
rect 20300 -1590 20366 -1574
rect 20300 -1654 20301 -1590
rect 20365 -1654 20366 -1590
rect 20300 -1670 20366 -1654
rect 20300 -1734 20301 -1670
rect 20365 -1734 20366 -1670
rect 20300 -1750 20366 -1734
rect 20300 -1814 20301 -1750
rect 20365 -1814 20366 -1750
rect 20300 -1830 20366 -1814
rect 20300 -1894 20301 -1830
rect 20365 -1894 20366 -1830
rect 20300 -1910 20366 -1894
rect 20300 -1974 20301 -1910
rect 20365 -1974 20366 -1910
rect 20300 -1990 20366 -1974
rect 20300 -2054 20301 -1990
rect 20365 -2054 20366 -1990
rect 20300 -2070 20366 -2054
rect 20300 -2134 20301 -2070
rect 20365 -2134 20366 -2070
rect 20300 -2150 20366 -2134
rect 20300 -2214 20301 -2150
rect 20365 -2214 20366 -2150
rect 20300 -2230 20366 -2214
rect 20300 -2294 20301 -2230
rect 20365 -2294 20366 -2230
rect 20300 -2384 20366 -2294
rect 20426 -2388 20486 -1356
rect 20546 -2448 20606 -1418
rect 20666 -2388 20726 -1356
rect 20786 -2448 20846 -1418
rect 20906 -1510 20972 -1356
rect 20906 -1574 20907 -1510
rect 20971 -1574 20972 -1510
rect 20906 -1590 20972 -1574
rect 20906 -1654 20907 -1590
rect 20971 -1654 20972 -1590
rect 20906 -1670 20972 -1654
rect 20906 -1734 20907 -1670
rect 20971 -1734 20972 -1670
rect 20906 -1750 20972 -1734
rect 20906 -1814 20907 -1750
rect 20971 -1814 20972 -1750
rect 20906 -1830 20972 -1814
rect 20906 -1894 20907 -1830
rect 20971 -1894 20972 -1830
rect 20906 -1910 20972 -1894
rect 20906 -1974 20907 -1910
rect 20971 -1974 20972 -1910
rect 20906 -1990 20972 -1974
rect 20906 -2054 20907 -1990
rect 20971 -2054 20972 -1990
rect 20906 -2070 20972 -2054
rect 20906 -2134 20907 -2070
rect 20971 -2134 20972 -2070
rect 20906 -2150 20972 -2134
rect 20906 -2214 20907 -2150
rect 20971 -2214 20972 -2150
rect 20906 -2230 20972 -2214
rect 20906 -2294 20907 -2230
rect 20971 -2294 20972 -2230
rect 20906 -2384 20972 -2294
rect 21032 -2388 21092 -1356
rect 21152 -2448 21212 -1418
rect 21272 -2388 21332 -1356
rect 21392 -2448 21452 -1418
rect 21512 -1510 21578 -1356
rect 21512 -1574 21513 -1510
rect 21577 -1574 21578 -1510
rect 21512 -1590 21578 -1574
rect 21512 -1654 21513 -1590
rect 21577 -1654 21578 -1590
rect 21512 -1670 21578 -1654
rect 21512 -1734 21513 -1670
rect 21577 -1734 21578 -1670
rect 21512 -1750 21578 -1734
rect 21512 -1814 21513 -1750
rect 21577 -1814 21578 -1750
rect 21512 -1830 21578 -1814
rect 21512 -1894 21513 -1830
rect 21577 -1894 21578 -1830
rect 21512 -1910 21578 -1894
rect 21512 -1974 21513 -1910
rect 21577 -1974 21578 -1910
rect 21512 -1990 21578 -1974
rect 21512 -2054 21513 -1990
rect 21577 -2054 21578 -1990
rect 21512 -2070 21578 -2054
rect 21512 -2134 21513 -2070
rect 21577 -2134 21578 -2070
rect 21512 -2150 21578 -2134
rect 21512 -2214 21513 -2150
rect 21577 -2214 21578 -2150
rect 21512 -2230 21578 -2214
rect 21512 -2294 21513 -2230
rect 21577 -2294 21578 -2230
rect 21512 -2384 21578 -2294
rect 21638 -2388 21698 -1356
rect 21758 -2448 21818 -1418
rect 21878 -2388 21938 -1356
rect 21998 -2448 22058 -1418
rect 22118 -1510 22184 -1356
rect 22118 -1574 22119 -1510
rect 22183 -1574 22184 -1510
rect 22118 -1590 22184 -1574
rect 22118 -1654 22119 -1590
rect 22183 -1654 22184 -1590
rect 22118 -1670 22184 -1654
rect 22118 -1734 22119 -1670
rect 22183 -1734 22184 -1670
rect 22118 -1750 22184 -1734
rect 22118 -1814 22119 -1750
rect 22183 -1814 22184 -1750
rect 22118 -1830 22184 -1814
rect 22118 -1894 22119 -1830
rect 22183 -1894 22184 -1830
rect 22118 -1910 22184 -1894
rect 22118 -1974 22119 -1910
rect 22183 -1974 22184 -1910
rect 22118 -1990 22184 -1974
rect 22118 -2054 22119 -1990
rect 22183 -2054 22184 -1990
rect 22118 -2070 22184 -2054
rect 22118 -2134 22119 -2070
rect 22183 -2134 22184 -2070
rect 22118 -2150 22184 -2134
rect 22118 -2214 22119 -2150
rect 22183 -2214 22184 -2150
rect 22118 -2230 22184 -2214
rect 22118 -2294 22119 -2230
rect 22183 -2294 22184 -2230
rect 22118 -2384 22184 -2294
rect 22244 -2388 22304 -1356
rect 22364 -2448 22424 -1418
rect 22484 -2388 22544 -1356
rect 22604 -2448 22664 -1418
rect 22724 -1510 22790 -1356
rect 22724 -1574 22725 -1510
rect 22789 -1574 22790 -1510
rect 22724 -1590 22790 -1574
rect 22724 -1654 22725 -1590
rect 22789 -1654 22790 -1590
rect 22724 -1670 22790 -1654
rect 22724 -1734 22725 -1670
rect 22789 -1734 22790 -1670
rect 22724 -1750 22790 -1734
rect 22724 -1814 22725 -1750
rect 22789 -1814 22790 -1750
rect 22724 -1830 22790 -1814
rect 22724 -1894 22725 -1830
rect 22789 -1894 22790 -1830
rect 22724 -1910 22790 -1894
rect 22724 -1974 22725 -1910
rect 22789 -1974 22790 -1910
rect 22724 -1990 22790 -1974
rect 22724 -2054 22725 -1990
rect 22789 -2054 22790 -1990
rect 22724 -2070 22790 -2054
rect 22724 -2134 22725 -2070
rect 22789 -2134 22790 -2070
rect 22724 -2150 22790 -2134
rect 22724 -2214 22725 -2150
rect 22789 -2214 22790 -2150
rect 22724 -2230 22790 -2214
rect 22724 -2294 22725 -2230
rect 22789 -2294 22790 -2230
rect 22724 -2384 22790 -2294
rect 22850 -2388 22910 -1356
rect 22970 -2448 23030 -1418
rect 23090 -2388 23150 -1356
rect 23210 -2448 23270 -1418
rect 23330 -1510 23396 -1356
rect 23330 -1574 23331 -1510
rect 23395 -1574 23396 -1510
rect 23330 -1590 23396 -1574
rect 23330 -1654 23331 -1590
rect 23395 -1654 23396 -1590
rect 23330 -1670 23396 -1654
rect 23330 -1734 23331 -1670
rect 23395 -1734 23396 -1670
rect 23330 -1750 23396 -1734
rect 23330 -1814 23331 -1750
rect 23395 -1814 23396 -1750
rect 23330 -1830 23396 -1814
rect 23330 -1894 23331 -1830
rect 23395 -1894 23396 -1830
rect 23330 -1910 23396 -1894
rect 23330 -1974 23331 -1910
rect 23395 -1974 23396 -1910
rect 23330 -1990 23396 -1974
rect 23330 -2054 23331 -1990
rect 23395 -2054 23396 -1990
rect 23330 -2070 23396 -2054
rect 23330 -2134 23331 -2070
rect 23395 -2134 23396 -2070
rect 23330 -2150 23396 -2134
rect 23330 -2214 23331 -2150
rect 23395 -2214 23396 -2150
rect 23330 -2230 23396 -2214
rect 23330 -2294 23331 -2230
rect 23395 -2294 23396 -2230
rect 23330 -2384 23396 -2294
rect 23456 -2388 23516 -1356
rect 23576 -2448 23636 -1418
rect 23696 -2388 23756 -1356
rect 23816 -2448 23876 -1418
rect 23936 -1510 24002 -1356
rect 23936 -1574 23937 -1510
rect 24001 -1574 24002 -1510
rect 23936 -1590 24002 -1574
rect 23936 -1654 23937 -1590
rect 24001 -1654 24002 -1590
rect 23936 -1670 24002 -1654
rect 23936 -1734 23937 -1670
rect 24001 -1734 24002 -1670
rect 23936 -1750 24002 -1734
rect 23936 -1814 23937 -1750
rect 24001 -1814 24002 -1750
rect 23936 -1830 24002 -1814
rect 23936 -1894 23937 -1830
rect 24001 -1894 24002 -1830
rect 23936 -1910 24002 -1894
rect 23936 -1974 23937 -1910
rect 24001 -1974 24002 -1910
rect 23936 -1990 24002 -1974
rect 23936 -2054 23937 -1990
rect 24001 -2054 24002 -1990
rect 23936 -2070 24002 -2054
rect 23936 -2134 23937 -2070
rect 24001 -2134 24002 -2070
rect 23936 -2150 24002 -2134
rect 23936 -2214 23937 -2150
rect 24001 -2214 24002 -2150
rect 23936 -2230 24002 -2214
rect 23936 -2294 23937 -2230
rect 24001 -2294 24002 -2230
rect 23936 -2384 24002 -2294
rect 24062 -2388 24122 -1356
rect 24182 -2448 24242 -1418
rect 24302 -2388 24362 -1356
rect 24422 -2448 24482 -1418
rect 24542 -1510 24608 -1356
rect 24542 -1574 24543 -1510
rect 24607 -1574 24608 -1510
rect 24542 -1590 24608 -1574
rect 24542 -1654 24543 -1590
rect 24607 -1654 24608 -1590
rect 24542 -1670 24608 -1654
rect 24542 -1734 24543 -1670
rect 24607 -1734 24608 -1670
rect 24542 -1750 24608 -1734
rect 24542 -1814 24543 -1750
rect 24607 -1814 24608 -1750
rect 24542 -1830 24608 -1814
rect 24542 -1894 24543 -1830
rect 24607 -1894 24608 -1830
rect 24542 -1910 24608 -1894
rect 24542 -1974 24543 -1910
rect 24607 -1974 24608 -1910
rect 24542 -1990 24608 -1974
rect 24542 -2054 24543 -1990
rect 24607 -2054 24608 -1990
rect 24542 -2070 24608 -2054
rect 24542 -2134 24543 -2070
rect 24607 -2134 24608 -2070
rect 24542 -2150 24608 -2134
rect 24542 -2214 24543 -2150
rect 24607 -2214 24608 -2150
rect 24542 -2230 24608 -2214
rect 24542 -2294 24543 -2230
rect 24607 -2294 24608 -2230
rect 24542 -2384 24608 -2294
rect 24668 -2388 24728 -1356
rect 24788 -2448 24848 -1418
rect 24908 -2388 24968 -1356
rect 25028 -2448 25088 -1418
rect 25148 -1510 25214 -1356
rect 25148 -1574 25149 -1510
rect 25213 -1574 25214 -1510
rect 25148 -1590 25214 -1574
rect 25148 -1654 25149 -1590
rect 25213 -1654 25214 -1590
rect 25148 -1670 25214 -1654
rect 25148 -1734 25149 -1670
rect 25213 -1734 25214 -1670
rect 25148 -1750 25214 -1734
rect 25148 -1814 25149 -1750
rect 25213 -1814 25214 -1750
rect 25148 -1830 25214 -1814
rect 25148 -1894 25149 -1830
rect 25213 -1894 25214 -1830
rect 25148 -1910 25214 -1894
rect 25148 -1974 25149 -1910
rect 25213 -1974 25214 -1910
rect 25148 -1990 25214 -1974
rect 25148 -2054 25149 -1990
rect 25213 -2054 25214 -1990
rect 25148 -2070 25214 -2054
rect 25148 -2134 25149 -2070
rect 25213 -2134 25214 -2070
rect 25148 -2150 25214 -2134
rect 25148 -2214 25149 -2150
rect 25213 -2214 25214 -2150
rect 25148 -2230 25214 -2214
rect 25148 -2294 25149 -2230
rect 25213 -2294 25214 -2230
rect 25148 -2384 25214 -2294
rect 25274 -2388 25334 -1356
rect 25394 -2448 25454 -1418
rect 25514 -2388 25574 -1356
rect 25634 -2448 25694 -1418
rect 25754 -1510 25820 -1356
rect 25754 -1574 25755 -1510
rect 25819 -1574 25820 -1510
rect 25754 -1590 25820 -1574
rect 25754 -1654 25755 -1590
rect 25819 -1654 25820 -1590
rect 25754 -1670 25820 -1654
rect 25754 -1734 25755 -1670
rect 25819 -1734 25820 -1670
rect 25754 -1750 25820 -1734
rect 25754 -1814 25755 -1750
rect 25819 -1814 25820 -1750
rect 25754 -1830 25820 -1814
rect 25754 -1894 25755 -1830
rect 25819 -1894 25820 -1830
rect 25754 -1910 25820 -1894
rect 25754 -1974 25755 -1910
rect 25819 -1974 25820 -1910
rect 25754 -1990 25820 -1974
rect 25754 -2054 25755 -1990
rect 25819 -2054 25820 -1990
rect 25754 -2070 25820 -2054
rect 25754 -2134 25755 -2070
rect 25819 -2134 25820 -2070
rect 25754 -2150 25820 -2134
rect 25754 -2214 25755 -2150
rect 25819 -2214 25820 -2150
rect 25754 -2230 25820 -2214
rect 25754 -2294 25755 -2230
rect 25819 -2294 25820 -2230
rect 25754 -2384 25820 -2294
rect 25880 -2388 25940 -1356
rect 26000 -2448 26060 -1418
rect 26120 -2388 26180 -1356
rect 26240 -2448 26300 -1418
rect 26360 -1510 26426 -1356
rect 26360 -1574 26361 -1510
rect 26425 -1574 26426 -1510
rect 26360 -1590 26426 -1574
rect 26360 -1654 26361 -1590
rect 26425 -1654 26426 -1590
rect 26360 -1670 26426 -1654
rect 26360 -1734 26361 -1670
rect 26425 -1734 26426 -1670
rect 26360 -1750 26426 -1734
rect 26360 -1814 26361 -1750
rect 26425 -1814 26426 -1750
rect 26360 -1830 26426 -1814
rect 26360 -1894 26361 -1830
rect 26425 -1894 26426 -1830
rect 26360 -1910 26426 -1894
rect 26360 -1974 26361 -1910
rect 26425 -1974 26426 -1910
rect 26360 -1990 26426 -1974
rect 26360 -2054 26361 -1990
rect 26425 -2054 26426 -1990
rect 26360 -2070 26426 -2054
rect 26360 -2134 26361 -2070
rect 26425 -2134 26426 -2070
rect 26360 -2150 26426 -2134
rect 26360 -2214 26361 -2150
rect 26425 -2214 26426 -2150
rect 26360 -2230 26426 -2214
rect 26360 -2294 26361 -2230
rect 26425 -2294 26426 -2230
rect 26360 -2384 26426 -2294
rect 26486 -2388 26546 -1356
rect 26606 -2448 26666 -1418
rect 26726 -2388 26786 -1356
rect 26846 -2448 26906 -1418
rect 26966 -1510 27032 -1356
rect 26966 -1574 26967 -1510
rect 27031 -1574 27032 -1510
rect 26966 -1590 27032 -1574
rect 26966 -1654 26967 -1590
rect 27031 -1654 27032 -1590
rect 26966 -1670 27032 -1654
rect 26966 -1734 26967 -1670
rect 27031 -1734 27032 -1670
rect 26966 -1750 27032 -1734
rect 26966 -1814 26967 -1750
rect 27031 -1814 27032 -1750
rect 26966 -1830 27032 -1814
rect 26966 -1894 26967 -1830
rect 27031 -1894 27032 -1830
rect 26966 -1910 27032 -1894
rect 26966 -1974 26967 -1910
rect 27031 -1974 27032 -1910
rect 26966 -1990 27032 -1974
rect 26966 -2054 26967 -1990
rect 27031 -2054 27032 -1990
rect 26966 -2070 27032 -2054
rect 26966 -2134 26967 -2070
rect 27031 -2134 27032 -2070
rect 26966 -2150 27032 -2134
rect 26966 -2214 26967 -2150
rect 27031 -2214 27032 -2150
rect 26966 -2230 27032 -2214
rect 26966 -2294 26967 -2230
rect 27031 -2294 27032 -2230
rect 26966 -2384 27032 -2294
rect 27092 -2388 27152 -1356
rect 27212 -2448 27272 -1418
rect 27332 -2388 27392 -1356
rect 27452 -2448 27512 -1418
rect 27572 -1510 27638 -1356
rect 27572 -1574 27573 -1510
rect 27637 -1574 27638 -1510
rect 27572 -1590 27638 -1574
rect 27572 -1654 27573 -1590
rect 27637 -1654 27638 -1590
rect 27572 -1670 27638 -1654
rect 27572 -1734 27573 -1670
rect 27637 -1734 27638 -1670
rect 27572 -1750 27638 -1734
rect 27572 -1814 27573 -1750
rect 27637 -1814 27638 -1750
rect 27572 -1830 27638 -1814
rect 27572 -1894 27573 -1830
rect 27637 -1894 27638 -1830
rect 27572 -1910 27638 -1894
rect 27572 -1974 27573 -1910
rect 27637 -1974 27638 -1910
rect 27572 -1990 27638 -1974
rect 27572 -2054 27573 -1990
rect 27637 -2054 27638 -1990
rect 27572 -2070 27638 -2054
rect 27572 -2134 27573 -2070
rect 27637 -2134 27638 -2070
rect 27572 -2150 27638 -2134
rect 27572 -2214 27573 -2150
rect 27637 -2214 27638 -2150
rect 27572 -2230 27638 -2214
rect 27572 -2294 27573 -2230
rect 27637 -2294 27638 -2230
rect 27572 -2384 27638 -2294
rect 27698 -2388 27758 -1356
rect 27818 -2448 27878 -1418
rect 27938 -2388 27998 -1356
rect 28058 -2448 28118 -1418
rect 28178 -1510 28244 -1356
rect 28178 -1574 28179 -1510
rect 28243 -1574 28244 -1510
rect 28178 -1590 28244 -1574
rect 28178 -1654 28179 -1590
rect 28243 -1654 28244 -1590
rect 28178 -1670 28244 -1654
rect 28178 -1734 28179 -1670
rect 28243 -1734 28244 -1670
rect 28178 -1750 28244 -1734
rect 28178 -1814 28179 -1750
rect 28243 -1814 28244 -1750
rect 28178 -1830 28244 -1814
rect 28178 -1894 28179 -1830
rect 28243 -1894 28244 -1830
rect 28178 -1910 28244 -1894
rect 28178 -1974 28179 -1910
rect 28243 -1974 28244 -1910
rect 28178 -1990 28244 -1974
rect 28178 -2054 28179 -1990
rect 28243 -2054 28244 -1990
rect 28178 -2070 28244 -2054
rect 28178 -2134 28179 -2070
rect 28243 -2134 28244 -2070
rect 28178 -2150 28244 -2134
rect 28178 -2214 28179 -2150
rect 28243 -2214 28244 -2150
rect 28178 -2230 28244 -2214
rect 28178 -2294 28179 -2230
rect 28243 -2294 28244 -2230
rect 28178 -2384 28244 -2294
rect 28304 -2388 28364 -1356
rect 28424 -2448 28484 -1418
rect 28544 -2388 28604 -1356
rect 28664 -2448 28724 -1418
rect 28784 -1510 28850 -1356
rect 28784 -1574 28785 -1510
rect 28849 -1574 28850 -1510
rect 28784 -1590 28850 -1574
rect 28784 -1654 28785 -1590
rect 28849 -1654 28850 -1590
rect 28784 -1670 28850 -1654
rect 28784 -1734 28785 -1670
rect 28849 -1734 28850 -1670
rect 28784 -1750 28850 -1734
rect 28784 -1814 28785 -1750
rect 28849 -1814 28850 -1750
rect 28784 -1830 28850 -1814
rect 28784 -1894 28785 -1830
rect 28849 -1894 28850 -1830
rect 28784 -1910 28850 -1894
rect 28784 -1974 28785 -1910
rect 28849 -1974 28850 -1910
rect 28784 -1990 28850 -1974
rect 28784 -2054 28785 -1990
rect 28849 -2054 28850 -1990
rect 28784 -2070 28850 -2054
rect 28784 -2134 28785 -2070
rect 28849 -2134 28850 -2070
rect 28784 -2150 28850 -2134
rect 28784 -2214 28785 -2150
rect 28849 -2214 28850 -2150
rect 28784 -2230 28850 -2214
rect 28784 -2294 28785 -2230
rect 28849 -2294 28850 -2230
rect 28784 -2384 28850 -2294
rect 19088 -2450 28850 -2448
rect 19088 -2514 19192 -2450
rect 19256 -2514 19272 -2450
rect 19336 -2514 19352 -2450
rect 19416 -2514 19432 -2450
rect 19496 -2514 19512 -2450
rect 19576 -2514 19592 -2450
rect 19656 -2514 19798 -2450
rect 19862 -2514 19878 -2450
rect 19942 -2514 19958 -2450
rect 20022 -2514 20038 -2450
rect 20102 -2514 20118 -2450
rect 20182 -2514 20198 -2450
rect 20262 -2514 20404 -2450
rect 20468 -2514 20484 -2450
rect 20548 -2514 20564 -2450
rect 20628 -2514 20644 -2450
rect 20708 -2514 20724 -2450
rect 20788 -2514 20804 -2450
rect 20868 -2514 21010 -2450
rect 21074 -2514 21090 -2450
rect 21154 -2514 21170 -2450
rect 21234 -2514 21250 -2450
rect 21314 -2514 21330 -2450
rect 21394 -2514 21410 -2450
rect 21474 -2514 21616 -2450
rect 21680 -2514 21696 -2450
rect 21760 -2514 21776 -2450
rect 21840 -2514 21856 -2450
rect 21920 -2514 21936 -2450
rect 22000 -2514 22016 -2450
rect 22080 -2514 22222 -2450
rect 22286 -2514 22302 -2450
rect 22366 -2514 22382 -2450
rect 22446 -2514 22462 -2450
rect 22526 -2514 22542 -2450
rect 22606 -2514 22622 -2450
rect 22686 -2514 22828 -2450
rect 22892 -2514 22908 -2450
rect 22972 -2514 22988 -2450
rect 23052 -2514 23068 -2450
rect 23132 -2514 23148 -2450
rect 23212 -2514 23228 -2450
rect 23292 -2514 23434 -2450
rect 23498 -2514 23514 -2450
rect 23578 -2514 23594 -2450
rect 23658 -2514 23674 -2450
rect 23738 -2514 23754 -2450
rect 23818 -2514 23834 -2450
rect 23898 -2514 24040 -2450
rect 24104 -2514 24120 -2450
rect 24184 -2514 24200 -2450
rect 24264 -2514 24280 -2450
rect 24344 -2514 24360 -2450
rect 24424 -2514 24440 -2450
rect 24504 -2514 24646 -2450
rect 24710 -2514 24726 -2450
rect 24790 -2514 24806 -2450
rect 24870 -2514 24886 -2450
rect 24950 -2514 24966 -2450
rect 25030 -2514 25046 -2450
rect 25110 -2514 25252 -2450
rect 25316 -2514 25332 -2450
rect 25396 -2514 25412 -2450
rect 25476 -2514 25492 -2450
rect 25556 -2514 25572 -2450
rect 25636 -2514 25652 -2450
rect 25716 -2514 25858 -2450
rect 25922 -2514 25938 -2450
rect 26002 -2514 26018 -2450
rect 26082 -2514 26098 -2450
rect 26162 -2514 26178 -2450
rect 26242 -2514 26258 -2450
rect 26322 -2514 26464 -2450
rect 26528 -2514 26544 -2450
rect 26608 -2514 26624 -2450
rect 26688 -2514 26704 -2450
rect 26768 -2514 26784 -2450
rect 26848 -2514 26864 -2450
rect 26928 -2514 27070 -2450
rect 27134 -2514 27150 -2450
rect 27214 -2514 27230 -2450
rect 27294 -2514 27310 -2450
rect 27374 -2514 27390 -2450
rect 27454 -2514 27470 -2450
rect 27534 -2514 27676 -2450
rect 27740 -2514 27756 -2450
rect 27820 -2514 27836 -2450
rect 27900 -2514 27916 -2450
rect 27980 -2514 27996 -2450
rect 28060 -2514 28076 -2450
rect 28140 -2514 28282 -2450
rect 28346 -2514 28362 -2450
rect 28426 -2514 28442 -2450
rect 28506 -2514 28522 -2450
rect 28586 -2514 28602 -2450
rect 28666 -2514 28682 -2450
rect 28746 -2514 28850 -2450
rect 19088 -2516 28850 -2514
<< via3 >>
rect 19192 -194 19256 -130
rect 19272 -194 19336 -130
rect 19352 -194 19416 -130
rect 19432 -194 19496 -130
rect 19512 -194 19576 -130
rect 19592 -194 19656 -130
rect 19798 -194 19862 -130
rect 19878 -194 19942 -130
rect 19958 -194 20022 -130
rect 20038 -194 20102 -130
rect 20118 -194 20182 -130
rect 20198 -194 20262 -130
rect 20404 -194 20468 -130
rect 20484 -194 20548 -130
rect 20564 -194 20628 -130
rect 20644 -194 20708 -130
rect 20724 -194 20788 -130
rect 20804 -194 20868 -130
rect 21010 -194 21074 -130
rect 21090 -194 21154 -130
rect 21170 -194 21234 -130
rect 21250 -194 21314 -130
rect 21330 -194 21394 -130
rect 21410 -194 21474 -130
rect 21616 -194 21680 -130
rect 21696 -194 21760 -130
rect 21776 -194 21840 -130
rect 21856 -194 21920 -130
rect 21936 -194 22000 -130
rect 22016 -194 22080 -130
rect 22222 -194 22286 -130
rect 22302 -194 22366 -130
rect 22382 -194 22446 -130
rect 22462 -194 22526 -130
rect 22542 -194 22606 -130
rect 22622 -194 22686 -130
rect 22828 -194 22892 -130
rect 22908 -194 22972 -130
rect 22988 -194 23052 -130
rect 23068 -194 23132 -130
rect 23148 -194 23212 -130
rect 23228 -194 23292 -130
rect 23434 -194 23498 -130
rect 23514 -194 23578 -130
rect 23594 -194 23658 -130
rect 23674 -194 23738 -130
rect 23754 -194 23818 -130
rect 23834 -194 23898 -130
rect 24040 -194 24104 -130
rect 24120 -194 24184 -130
rect 24200 -194 24264 -130
rect 24280 -194 24344 -130
rect 24360 -194 24424 -130
rect 24440 -194 24504 -130
rect 24646 -194 24710 -130
rect 24726 -194 24790 -130
rect 24806 -194 24870 -130
rect 24886 -194 24950 -130
rect 24966 -194 25030 -130
rect 25046 -194 25110 -130
rect 25252 -194 25316 -130
rect 25332 -194 25396 -130
rect 25412 -194 25476 -130
rect 25492 -194 25556 -130
rect 25572 -194 25636 -130
rect 25652 -194 25716 -130
rect 25858 -194 25922 -130
rect 25938 -194 26002 -130
rect 26018 -194 26082 -130
rect 26098 -194 26162 -130
rect 26178 -194 26242 -130
rect 26258 -194 26322 -130
rect 26464 -194 26528 -130
rect 26544 -194 26608 -130
rect 26624 -194 26688 -130
rect 26704 -194 26768 -130
rect 26784 -194 26848 -130
rect 26864 -194 26928 -130
rect 27070 -194 27134 -130
rect 27150 -194 27214 -130
rect 27230 -194 27294 -130
rect 27310 -194 27374 -130
rect 27390 -194 27454 -130
rect 27470 -194 27534 -130
rect 27676 -194 27740 -130
rect 27756 -194 27820 -130
rect 27836 -194 27900 -130
rect 27916 -194 27980 -130
rect 27996 -194 28060 -130
rect 28076 -194 28140 -130
rect 28282 -194 28346 -130
rect 28362 -194 28426 -130
rect 28442 -194 28506 -130
rect 28522 -194 28586 -130
rect 28602 -194 28666 -130
rect 28682 -194 28746 -130
rect 19089 -414 19153 -350
rect 19089 -494 19153 -430
rect 19089 -574 19153 -510
rect 19089 -654 19153 -590
rect 19089 -734 19153 -670
rect 19089 -814 19153 -750
rect 19089 -894 19153 -830
rect 19089 -974 19153 -910
rect 19089 -1054 19153 -990
rect 19089 -1134 19153 -1070
rect 19695 -414 19759 -350
rect 19695 -494 19759 -430
rect 19695 -574 19759 -510
rect 19695 -654 19759 -590
rect 19695 -734 19759 -670
rect 19695 -814 19759 -750
rect 19695 -894 19759 -830
rect 19695 -974 19759 -910
rect 19695 -1054 19759 -990
rect 19695 -1134 19759 -1070
rect 20301 -414 20365 -350
rect 20301 -494 20365 -430
rect 20301 -574 20365 -510
rect 20301 -654 20365 -590
rect 20301 -734 20365 -670
rect 20301 -814 20365 -750
rect 20301 -894 20365 -830
rect 20301 -974 20365 -910
rect 20301 -1054 20365 -990
rect 20301 -1134 20365 -1070
rect 20907 -414 20971 -350
rect 20907 -494 20971 -430
rect 20907 -574 20971 -510
rect 20907 -654 20971 -590
rect 20907 -734 20971 -670
rect 20907 -814 20971 -750
rect 20907 -894 20971 -830
rect 20907 -974 20971 -910
rect 20907 -1054 20971 -990
rect 20907 -1134 20971 -1070
rect 21513 -414 21577 -350
rect 21513 -494 21577 -430
rect 21513 -574 21577 -510
rect 21513 -654 21577 -590
rect 21513 -734 21577 -670
rect 21513 -814 21577 -750
rect 21513 -894 21577 -830
rect 21513 -974 21577 -910
rect 21513 -1054 21577 -990
rect 21513 -1134 21577 -1070
rect 22119 -414 22183 -350
rect 22119 -494 22183 -430
rect 22119 -574 22183 -510
rect 22119 -654 22183 -590
rect 22119 -734 22183 -670
rect 22119 -814 22183 -750
rect 22119 -894 22183 -830
rect 22119 -974 22183 -910
rect 22119 -1054 22183 -990
rect 22119 -1134 22183 -1070
rect 22725 -414 22789 -350
rect 22725 -494 22789 -430
rect 22725 -574 22789 -510
rect 22725 -654 22789 -590
rect 22725 -734 22789 -670
rect 22725 -814 22789 -750
rect 22725 -894 22789 -830
rect 22725 -974 22789 -910
rect 22725 -1054 22789 -990
rect 22725 -1134 22789 -1070
rect 23331 -414 23395 -350
rect 23331 -494 23395 -430
rect 23331 -574 23395 -510
rect 23331 -654 23395 -590
rect 23331 -734 23395 -670
rect 23331 -814 23395 -750
rect 23331 -894 23395 -830
rect 23331 -974 23395 -910
rect 23331 -1054 23395 -990
rect 23331 -1134 23395 -1070
rect 23937 -414 24001 -350
rect 23937 -494 24001 -430
rect 23937 -574 24001 -510
rect 23937 -654 24001 -590
rect 23937 -734 24001 -670
rect 23937 -814 24001 -750
rect 23937 -894 24001 -830
rect 23937 -974 24001 -910
rect 23937 -1054 24001 -990
rect 23937 -1134 24001 -1070
rect 24543 -414 24607 -350
rect 24543 -494 24607 -430
rect 24543 -574 24607 -510
rect 24543 -654 24607 -590
rect 24543 -734 24607 -670
rect 24543 -814 24607 -750
rect 24543 -894 24607 -830
rect 24543 -974 24607 -910
rect 24543 -1054 24607 -990
rect 24543 -1134 24607 -1070
rect 25149 -414 25213 -350
rect 25149 -494 25213 -430
rect 25149 -574 25213 -510
rect 25149 -654 25213 -590
rect 25149 -734 25213 -670
rect 25149 -814 25213 -750
rect 25149 -894 25213 -830
rect 25149 -974 25213 -910
rect 25149 -1054 25213 -990
rect 25149 -1134 25213 -1070
rect 25755 -414 25819 -350
rect 25755 -494 25819 -430
rect 25755 -574 25819 -510
rect 25755 -654 25819 -590
rect 25755 -734 25819 -670
rect 25755 -814 25819 -750
rect 25755 -894 25819 -830
rect 25755 -974 25819 -910
rect 25755 -1054 25819 -990
rect 25755 -1134 25819 -1070
rect 26361 -414 26425 -350
rect 26361 -494 26425 -430
rect 26361 -574 26425 -510
rect 26361 -654 26425 -590
rect 26361 -734 26425 -670
rect 26361 -814 26425 -750
rect 26361 -894 26425 -830
rect 26361 -974 26425 -910
rect 26361 -1054 26425 -990
rect 26361 -1134 26425 -1070
rect 26967 -414 27031 -350
rect 26967 -494 27031 -430
rect 26967 -574 27031 -510
rect 26967 -654 27031 -590
rect 26967 -734 27031 -670
rect 26967 -814 27031 -750
rect 26967 -894 27031 -830
rect 26967 -974 27031 -910
rect 26967 -1054 27031 -990
rect 26967 -1134 27031 -1070
rect 27573 -414 27637 -350
rect 27573 -494 27637 -430
rect 27573 -574 27637 -510
rect 27573 -654 27637 -590
rect 27573 -734 27637 -670
rect 27573 -814 27637 -750
rect 27573 -894 27637 -830
rect 27573 -974 27637 -910
rect 27573 -1054 27637 -990
rect 27573 -1134 27637 -1070
rect 28179 -414 28243 -350
rect 28179 -494 28243 -430
rect 28179 -574 28243 -510
rect 28179 -654 28243 -590
rect 28179 -734 28243 -670
rect 28179 -814 28243 -750
rect 28179 -894 28243 -830
rect 28179 -974 28243 -910
rect 28179 -1054 28243 -990
rect 28179 -1134 28243 -1070
rect 28785 -414 28849 -350
rect 28785 -494 28849 -430
rect 28785 -574 28849 -510
rect 28785 -654 28849 -590
rect 28785 -734 28849 -670
rect 28785 -814 28849 -750
rect 28785 -894 28849 -830
rect 28785 -974 28849 -910
rect 28785 -1054 28849 -990
rect 28785 -1134 28849 -1070
rect 19192 -1354 19256 -1290
rect 19272 -1354 19336 -1290
rect 19352 -1354 19416 -1290
rect 19432 -1354 19496 -1290
rect 19512 -1354 19576 -1290
rect 19592 -1354 19656 -1290
rect 19798 -1354 19862 -1290
rect 19878 -1354 19942 -1290
rect 19958 -1354 20022 -1290
rect 20038 -1354 20102 -1290
rect 20118 -1354 20182 -1290
rect 20198 -1354 20262 -1290
rect 20404 -1354 20468 -1290
rect 20484 -1354 20548 -1290
rect 20564 -1354 20628 -1290
rect 20644 -1354 20708 -1290
rect 20724 -1354 20788 -1290
rect 20804 -1354 20868 -1290
rect 21010 -1354 21074 -1290
rect 21090 -1354 21154 -1290
rect 21170 -1354 21234 -1290
rect 21250 -1354 21314 -1290
rect 21330 -1354 21394 -1290
rect 21410 -1354 21474 -1290
rect 21616 -1354 21680 -1290
rect 21696 -1354 21760 -1290
rect 21776 -1354 21840 -1290
rect 21856 -1354 21920 -1290
rect 21936 -1354 22000 -1290
rect 22016 -1354 22080 -1290
rect 22222 -1354 22286 -1290
rect 22302 -1354 22366 -1290
rect 22382 -1354 22446 -1290
rect 22462 -1354 22526 -1290
rect 22542 -1354 22606 -1290
rect 22622 -1354 22686 -1290
rect 22828 -1354 22892 -1290
rect 22908 -1354 22972 -1290
rect 22988 -1354 23052 -1290
rect 23068 -1354 23132 -1290
rect 23148 -1354 23212 -1290
rect 23228 -1354 23292 -1290
rect 23434 -1354 23498 -1290
rect 23514 -1354 23578 -1290
rect 23594 -1354 23658 -1290
rect 23674 -1354 23738 -1290
rect 23754 -1354 23818 -1290
rect 23834 -1354 23898 -1290
rect 24040 -1354 24104 -1290
rect 24120 -1354 24184 -1290
rect 24200 -1354 24264 -1290
rect 24280 -1354 24344 -1290
rect 24360 -1354 24424 -1290
rect 24440 -1354 24504 -1290
rect 24646 -1354 24710 -1290
rect 24726 -1354 24790 -1290
rect 24806 -1354 24870 -1290
rect 24886 -1354 24950 -1290
rect 24966 -1354 25030 -1290
rect 25046 -1354 25110 -1290
rect 25252 -1354 25316 -1290
rect 25332 -1354 25396 -1290
rect 25412 -1354 25476 -1290
rect 25492 -1354 25556 -1290
rect 25572 -1354 25636 -1290
rect 25652 -1354 25716 -1290
rect 25858 -1354 25922 -1290
rect 25938 -1354 26002 -1290
rect 26018 -1354 26082 -1290
rect 26098 -1354 26162 -1290
rect 26178 -1354 26242 -1290
rect 26258 -1354 26322 -1290
rect 26464 -1354 26528 -1290
rect 26544 -1354 26608 -1290
rect 26624 -1354 26688 -1290
rect 26704 -1354 26768 -1290
rect 26784 -1354 26848 -1290
rect 26864 -1354 26928 -1290
rect 27070 -1354 27134 -1290
rect 27150 -1354 27214 -1290
rect 27230 -1354 27294 -1290
rect 27310 -1354 27374 -1290
rect 27390 -1354 27454 -1290
rect 27470 -1354 27534 -1290
rect 27676 -1354 27740 -1290
rect 27756 -1354 27820 -1290
rect 27836 -1354 27900 -1290
rect 27916 -1354 27980 -1290
rect 27996 -1354 28060 -1290
rect 28076 -1354 28140 -1290
rect 28282 -1354 28346 -1290
rect 28362 -1354 28426 -1290
rect 28442 -1354 28506 -1290
rect 28522 -1354 28586 -1290
rect 28602 -1354 28666 -1290
rect 28682 -1354 28746 -1290
rect 19089 -1574 19153 -1510
rect 19089 -1654 19153 -1590
rect 19089 -1734 19153 -1670
rect 19089 -1814 19153 -1750
rect 19089 -1894 19153 -1830
rect 19089 -1974 19153 -1910
rect 19089 -2054 19153 -1990
rect 19089 -2134 19153 -2070
rect 19089 -2214 19153 -2150
rect 19089 -2294 19153 -2230
rect 19695 -1574 19759 -1510
rect 19695 -1654 19759 -1590
rect 19695 -1734 19759 -1670
rect 19695 -1814 19759 -1750
rect 19695 -1894 19759 -1830
rect 19695 -1974 19759 -1910
rect 19695 -2054 19759 -1990
rect 19695 -2134 19759 -2070
rect 19695 -2214 19759 -2150
rect 19695 -2294 19759 -2230
rect 20301 -1574 20365 -1510
rect 20301 -1654 20365 -1590
rect 20301 -1734 20365 -1670
rect 20301 -1814 20365 -1750
rect 20301 -1894 20365 -1830
rect 20301 -1974 20365 -1910
rect 20301 -2054 20365 -1990
rect 20301 -2134 20365 -2070
rect 20301 -2214 20365 -2150
rect 20301 -2294 20365 -2230
rect 20907 -1574 20971 -1510
rect 20907 -1654 20971 -1590
rect 20907 -1734 20971 -1670
rect 20907 -1814 20971 -1750
rect 20907 -1894 20971 -1830
rect 20907 -1974 20971 -1910
rect 20907 -2054 20971 -1990
rect 20907 -2134 20971 -2070
rect 20907 -2214 20971 -2150
rect 20907 -2294 20971 -2230
rect 21513 -1574 21577 -1510
rect 21513 -1654 21577 -1590
rect 21513 -1734 21577 -1670
rect 21513 -1814 21577 -1750
rect 21513 -1894 21577 -1830
rect 21513 -1974 21577 -1910
rect 21513 -2054 21577 -1990
rect 21513 -2134 21577 -2070
rect 21513 -2214 21577 -2150
rect 21513 -2294 21577 -2230
rect 22119 -1574 22183 -1510
rect 22119 -1654 22183 -1590
rect 22119 -1734 22183 -1670
rect 22119 -1814 22183 -1750
rect 22119 -1894 22183 -1830
rect 22119 -1974 22183 -1910
rect 22119 -2054 22183 -1990
rect 22119 -2134 22183 -2070
rect 22119 -2214 22183 -2150
rect 22119 -2294 22183 -2230
rect 22725 -1574 22789 -1510
rect 22725 -1654 22789 -1590
rect 22725 -1734 22789 -1670
rect 22725 -1814 22789 -1750
rect 22725 -1894 22789 -1830
rect 22725 -1974 22789 -1910
rect 22725 -2054 22789 -1990
rect 22725 -2134 22789 -2070
rect 22725 -2214 22789 -2150
rect 22725 -2294 22789 -2230
rect 23331 -1574 23395 -1510
rect 23331 -1654 23395 -1590
rect 23331 -1734 23395 -1670
rect 23331 -1814 23395 -1750
rect 23331 -1894 23395 -1830
rect 23331 -1974 23395 -1910
rect 23331 -2054 23395 -1990
rect 23331 -2134 23395 -2070
rect 23331 -2214 23395 -2150
rect 23331 -2294 23395 -2230
rect 23937 -1574 24001 -1510
rect 23937 -1654 24001 -1590
rect 23937 -1734 24001 -1670
rect 23937 -1814 24001 -1750
rect 23937 -1894 24001 -1830
rect 23937 -1974 24001 -1910
rect 23937 -2054 24001 -1990
rect 23937 -2134 24001 -2070
rect 23937 -2214 24001 -2150
rect 23937 -2294 24001 -2230
rect 24543 -1574 24607 -1510
rect 24543 -1654 24607 -1590
rect 24543 -1734 24607 -1670
rect 24543 -1814 24607 -1750
rect 24543 -1894 24607 -1830
rect 24543 -1974 24607 -1910
rect 24543 -2054 24607 -1990
rect 24543 -2134 24607 -2070
rect 24543 -2214 24607 -2150
rect 24543 -2294 24607 -2230
rect 25149 -1574 25213 -1510
rect 25149 -1654 25213 -1590
rect 25149 -1734 25213 -1670
rect 25149 -1814 25213 -1750
rect 25149 -1894 25213 -1830
rect 25149 -1974 25213 -1910
rect 25149 -2054 25213 -1990
rect 25149 -2134 25213 -2070
rect 25149 -2214 25213 -2150
rect 25149 -2294 25213 -2230
rect 25755 -1574 25819 -1510
rect 25755 -1654 25819 -1590
rect 25755 -1734 25819 -1670
rect 25755 -1814 25819 -1750
rect 25755 -1894 25819 -1830
rect 25755 -1974 25819 -1910
rect 25755 -2054 25819 -1990
rect 25755 -2134 25819 -2070
rect 25755 -2214 25819 -2150
rect 25755 -2294 25819 -2230
rect 26361 -1574 26425 -1510
rect 26361 -1654 26425 -1590
rect 26361 -1734 26425 -1670
rect 26361 -1814 26425 -1750
rect 26361 -1894 26425 -1830
rect 26361 -1974 26425 -1910
rect 26361 -2054 26425 -1990
rect 26361 -2134 26425 -2070
rect 26361 -2214 26425 -2150
rect 26361 -2294 26425 -2230
rect 26967 -1574 27031 -1510
rect 26967 -1654 27031 -1590
rect 26967 -1734 27031 -1670
rect 26967 -1814 27031 -1750
rect 26967 -1894 27031 -1830
rect 26967 -1974 27031 -1910
rect 26967 -2054 27031 -1990
rect 26967 -2134 27031 -2070
rect 26967 -2214 27031 -2150
rect 26967 -2294 27031 -2230
rect 27573 -1574 27637 -1510
rect 27573 -1654 27637 -1590
rect 27573 -1734 27637 -1670
rect 27573 -1814 27637 -1750
rect 27573 -1894 27637 -1830
rect 27573 -1974 27637 -1910
rect 27573 -2054 27637 -1990
rect 27573 -2134 27637 -2070
rect 27573 -2214 27637 -2150
rect 27573 -2294 27637 -2230
rect 28179 -1574 28243 -1510
rect 28179 -1654 28243 -1590
rect 28179 -1734 28243 -1670
rect 28179 -1814 28243 -1750
rect 28179 -1894 28243 -1830
rect 28179 -1974 28243 -1910
rect 28179 -2054 28243 -1990
rect 28179 -2134 28243 -2070
rect 28179 -2214 28243 -2150
rect 28179 -2294 28243 -2230
rect 28785 -1574 28849 -1510
rect 28785 -1654 28849 -1590
rect 28785 -1734 28849 -1670
rect 28785 -1814 28849 -1750
rect 28785 -1894 28849 -1830
rect 28785 -1974 28849 -1910
rect 28785 -2054 28849 -1990
rect 28785 -2134 28849 -2070
rect 28785 -2214 28849 -2150
rect 28785 -2294 28849 -2230
rect 19192 -2514 19256 -2450
rect 19272 -2514 19336 -2450
rect 19352 -2514 19416 -2450
rect 19432 -2514 19496 -2450
rect 19512 -2514 19576 -2450
rect 19592 -2514 19656 -2450
rect 19798 -2514 19862 -2450
rect 19878 -2514 19942 -2450
rect 19958 -2514 20022 -2450
rect 20038 -2514 20102 -2450
rect 20118 -2514 20182 -2450
rect 20198 -2514 20262 -2450
rect 20404 -2514 20468 -2450
rect 20484 -2514 20548 -2450
rect 20564 -2514 20628 -2450
rect 20644 -2514 20708 -2450
rect 20724 -2514 20788 -2450
rect 20804 -2514 20868 -2450
rect 21010 -2514 21074 -2450
rect 21090 -2514 21154 -2450
rect 21170 -2514 21234 -2450
rect 21250 -2514 21314 -2450
rect 21330 -2514 21394 -2450
rect 21410 -2514 21474 -2450
rect 21616 -2514 21680 -2450
rect 21696 -2514 21760 -2450
rect 21776 -2514 21840 -2450
rect 21856 -2514 21920 -2450
rect 21936 -2514 22000 -2450
rect 22016 -2514 22080 -2450
rect 22222 -2514 22286 -2450
rect 22302 -2514 22366 -2450
rect 22382 -2514 22446 -2450
rect 22462 -2514 22526 -2450
rect 22542 -2514 22606 -2450
rect 22622 -2514 22686 -2450
rect 22828 -2514 22892 -2450
rect 22908 -2514 22972 -2450
rect 22988 -2514 23052 -2450
rect 23068 -2514 23132 -2450
rect 23148 -2514 23212 -2450
rect 23228 -2514 23292 -2450
rect 23434 -2514 23498 -2450
rect 23514 -2514 23578 -2450
rect 23594 -2514 23658 -2450
rect 23674 -2514 23738 -2450
rect 23754 -2514 23818 -2450
rect 23834 -2514 23898 -2450
rect 24040 -2514 24104 -2450
rect 24120 -2514 24184 -2450
rect 24200 -2514 24264 -2450
rect 24280 -2514 24344 -2450
rect 24360 -2514 24424 -2450
rect 24440 -2514 24504 -2450
rect 24646 -2514 24710 -2450
rect 24726 -2514 24790 -2450
rect 24806 -2514 24870 -2450
rect 24886 -2514 24950 -2450
rect 24966 -2514 25030 -2450
rect 25046 -2514 25110 -2450
rect 25252 -2514 25316 -2450
rect 25332 -2514 25396 -2450
rect 25412 -2514 25476 -2450
rect 25492 -2514 25556 -2450
rect 25572 -2514 25636 -2450
rect 25652 -2514 25716 -2450
rect 25858 -2514 25922 -2450
rect 25938 -2514 26002 -2450
rect 26018 -2514 26082 -2450
rect 26098 -2514 26162 -2450
rect 26178 -2514 26242 -2450
rect 26258 -2514 26322 -2450
rect 26464 -2514 26528 -2450
rect 26544 -2514 26608 -2450
rect 26624 -2514 26688 -2450
rect 26704 -2514 26768 -2450
rect 26784 -2514 26848 -2450
rect 26864 -2514 26928 -2450
rect 27070 -2514 27134 -2450
rect 27150 -2514 27214 -2450
rect 27230 -2514 27294 -2450
rect 27310 -2514 27374 -2450
rect 27390 -2514 27454 -2450
rect 27470 -2514 27534 -2450
rect 27676 -2514 27740 -2450
rect 27756 -2514 27820 -2450
rect 27836 -2514 27900 -2450
rect 27916 -2514 27980 -2450
rect 27996 -2514 28060 -2450
rect 28076 -2514 28140 -2450
rect 28282 -2514 28346 -2450
rect 28362 -2514 28426 -2450
rect 28442 -2514 28506 -2450
rect 28522 -2514 28586 -2450
rect 28602 -2514 28666 -2450
rect 28682 -2514 28746 -2450
<< metal4 >>
rect 19088 -130 28850 -128
rect 19088 -194 19192 -130
rect 19256 -194 19272 -130
rect 19336 -194 19352 -130
rect 19416 -194 19432 -130
rect 19496 -194 19512 -130
rect 19576 -194 19592 -130
rect 19656 -194 19798 -130
rect 19862 -194 19878 -130
rect 19942 -194 19958 -130
rect 20022 -194 20038 -130
rect 20102 -194 20118 -130
rect 20182 -194 20198 -130
rect 20262 -194 20404 -130
rect 20468 -194 20484 -130
rect 20548 -194 20564 -130
rect 20628 -194 20644 -130
rect 20708 -194 20724 -130
rect 20788 -194 20804 -130
rect 20868 -194 21010 -130
rect 21074 -194 21090 -130
rect 21154 -194 21170 -130
rect 21234 -194 21250 -130
rect 21314 -194 21330 -130
rect 21394 -194 21410 -130
rect 21474 -194 21616 -130
rect 21680 -194 21696 -130
rect 21760 -194 21776 -130
rect 21840 -194 21856 -130
rect 21920 -194 21936 -130
rect 22000 -194 22016 -130
rect 22080 -194 22222 -130
rect 22286 -194 22302 -130
rect 22366 -194 22382 -130
rect 22446 -194 22462 -130
rect 22526 -194 22542 -130
rect 22606 -194 22622 -130
rect 22686 -194 22828 -130
rect 22892 -194 22908 -130
rect 22972 -194 22988 -130
rect 23052 -194 23068 -130
rect 23132 -194 23148 -130
rect 23212 -194 23228 -130
rect 23292 -194 23434 -130
rect 23498 -194 23514 -130
rect 23578 -194 23594 -130
rect 23658 -194 23674 -130
rect 23738 -194 23754 -130
rect 23818 -194 23834 -130
rect 23898 -194 24040 -130
rect 24104 -194 24120 -130
rect 24184 -194 24200 -130
rect 24264 -194 24280 -130
rect 24344 -194 24360 -130
rect 24424 -194 24440 -130
rect 24504 -194 24646 -130
rect 24710 -194 24726 -130
rect 24790 -194 24806 -130
rect 24870 -194 24886 -130
rect 24950 -194 24966 -130
rect 25030 -194 25046 -130
rect 25110 -194 25252 -130
rect 25316 -194 25332 -130
rect 25396 -194 25412 -130
rect 25476 -194 25492 -130
rect 25556 -194 25572 -130
rect 25636 -194 25652 -130
rect 25716 -194 25858 -130
rect 25922 -194 25938 -130
rect 26002 -194 26018 -130
rect 26082 -194 26098 -130
rect 26162 -194 26178 -130
rect 26242 -194 26258 -130
rect 26322 -194 26464 -130
rect 26528 -194 26544 -130
rect 26608 -194 26624 -130
rect 26688 -194 26704 -130
rect 26768 -194 26784 -130
rect 26848 -194 26864 -130
rect 26928 -194 27070 -130
rect 27134 -194 27150 -130
rect 27214 -194 27230 -130
rect 27294 -194 27310 -130
rect 27374 -194 27390 -130
rect 27454 -194 27470 -130
rect 27534 -194 27676 -130
rect 27740 -194 27756 -130
rect 27820 -194 27836 -130
rect 27900 -194 27916 -130
rect 27980 -194 27996 -130
rect 28060 -194 28076 -130
rect 28140 -194 28282 -130
rect 28346 -194 28362 -130
rect 28426 -194 28442 -130
rect 28506 -194 28522 -130
rect 28586 -194 28602 -130
rect 28666 -194 28682 -130
rect 28746 -194 28850 -130
rect 19088 -196 28850 -194
rect 19088 -350 19154 -196
rect 19088 -414 19089 -350
rect 19153 -414 19154 -350
rect 19088 -430 19154 -414
rect 19088 -494 19089 -430
rect 19153 -494 19154 -430
rect 19088 -510 19154 -494
rect 19088 -574 19089 -510
rect 19153 -574 19154 -510
rect 19088 -590 19154 -574
rect 19088 -654 19089 -590
rect 19153 -654 19154 -590
rect 19088 -670 19154 -654
rect 19088 -734 19089 -670
rect 19153 -734 19154 -670
rect 19088 -750 19154 -734
rect 19088 -814 19089 -750
rect 19153 -814 19154 -750
rect 19088 -830 19154 -814
rect 19088 -894 19089 -830
rect 19153 -894 19154 -830
rect 19088 -910 19154 -894
rect 19088 -974 19089 -910
rect 19153 -974 19154 -910
rect 19088 -990 19154 -974
rect 19088 -1054 19089 -990
rect 19153 -1054 19154 -990
rect 19088 -1070 19154 -1054
rect 19088 -1134 19089 -1070
rect 19153 -1134 19154 -1070
rect 19088 -1224 19154 -1134
rect 19214 -1288 19274 -258
rect 19334 -1228 19394 -196
rect 19454 -1288 19514 -258
rect 19574 -1228 19634 -196
rect 19694 -350 19760 -196
rect 19694 -414 19695 -350
rect 19759 -414 19760 -350
rect 19694 -430 19760 -414
rect 19694 -494 19695 -430
rect 19759 -494 19760 -430
rect 19694 -510 19760 -494
rect 19694 -574 19695 -510
rect 19759 -574 19760 -510
rect 19694 -590 19760 -574
rect 19694 -654 19695 -590
rect 19759 -654 19760 -590
rect 19694 -670 19760 -654
rect 19694 -734 19695 -670
rect 19759 -734 19760 -670
rect 19694 -750 19760 -734
rect 19694 -814 19695 -750
rect 19759 -814 19760 -750
rect 19694 -830 19760 -814
rect 19694 -894 19695 -830
rect 19759 -894 19760 -830
rect 19694 -910 19760 -894
rect 19694 -974 19695 -910
rect 19759 -974 19760 -910
rect 19694 -990 19760 -974
rect 19694 -1054 19695 -990
rect 19759 -1054 19760 -990
rect 19694 -1070 19760 -1054
rect 19694 -1134 19695 -1070
rect 19759 -1134 19760 -1070
rect 19694 -1224 19760 -1134
rect 19820 -1288 19880 -258
rect 19940 -1228 20000 -196
rect 20060 -1288 20120 -258
rect 20180 -1228 20240 -196
rect 20300 -350 20366 -196
rect 20300 -414 20301 -350
rect 20365 -414 20366 -350
rect 20300 -430 20366 -414
rect 20300 -494 20301 -430
rect 20365 -494 20366 -430
rect 20300 -510 20366 -494
rect 20300 -574 20301 -510
rect 20365 -574 20366 -510
rect 20300 -590 20366 -574
rect 20300 -654 20301 -590
rect 20365 -654 20366 -590
rect 20300 -670 20366 -654
rect 20300 -734 20301 -670
rect 20365 -734 20366 -670
rect 20300 -750 20366 -734
rect 20300 -814 20301 -750
rect 20365 -814 20366 -750
rect 20300 -830 20366 -814
rect 20300 -894 20301 -830
rect 20365 -894 20366 -830
rect 20300 -910 20366 -894
rect 20300 -974 20301 -910
rect 20365 -974 20366 -910
rect 20300 -990 20366 -974
rect 20300 -1054 20301 -990
rect 20365 -1054 20366 -990
rect 20300 -1070 20366 -1054
rect 20300 -1134 20301 -1070
rect 20365 -1134 20366 -1070
rect 20300 -1224 20366 -1134
rect 20426 -1288 20486 -258
rect 20546 -1228 20606 -196
rect 20666 -1288 20726 -258
rect 20786 -1228 20846 -196
rect 20906 -350 20972 -196
rect 20906 -414 20907 -350
rect 20971 -414 20972 -350
rect 20906 -430 20972 -414
rect 20906 -494 20907 -430
rect 20971 -494 20972 -430
rect 20906 -510 20972 -494
rect 20906 -574 20907 -510
rect 20971 -574 20972 -510
rect 20906 -590 20972 -574
rect 20906 -654 20907 -590
rect 20971 -654 20972 -590
rect 20906 -670 20972 -654
rect 20906 -734 20907 -670
rect 20971 -734 20972 -670
rect 20906 -750 20972 -734
rect 20906 -814 20907 -750
rect 20971 -814 20972 -750
rect 20906 -830 20972 -814
rect 20906 -894 20907 -830
rect 20971 -894 20972 -830
rect 20906 -910 20972 -894
rect 20906 -974 20907 -910
rect 20971 -974 20972 -910
rect 20906 -990 20972 -974
rect 20906 -1054 20907 -990
rect 20971 -1054 20972 -990
rect 20906 -1070 20972 -1054
rect 20906 -1134 20907 -1070
rect 20971 -1134 20972 -1070
rect 20906 -1224 20972 -1134
rect 21032 -1288 21092 -258
rect 21152 -1228 21212 -196
rect 21272 -1288 21332 -258
rect 21392 -1228 21452 -196
rect 21512 -350 21578 -196
rect 21512 -414 21513 -350
rect 21577 -414 21578 -350
rect 21512 -430 21578 -414
rect 21512 -494 21513 -430
rect 21577 -494 21578 -430
rect 21512 -510 21578 -494
rect 21512 -574 21513 -510
rect 21577 -574 21578 -510
rect 21512 -590 21578 -574
rect 21512 -654 21513 -590
rect 21577 -654 21578 -590
rect 21512 -670 21578 -654
rect 21512 -734 21513 -670
rect 21577 -734 21578 -670
rect 21512 -750 21578 -734
rect 21512 -814 21513 -750
rect 21577 -814 21578 -750
rect 21512 -830 21578 -814
rect 21512 -894 21513 -830
rect 21577 -894 21578 -830
rect 21512 -910 21578 -894
rect 21512 -974 21513 -910
rect 21577 -974 21578 -910
rect 21512 -990 21578 -974
rect 21512 -1054 21513 -990
rect 21577 -1054 21578 -990
rect 21512 -1070 21578 -1054
rect 21512 -1134 21513 -1070
rect 21577 -1134 21578 -1070
rect 21512 -1224 21578 -1134
rect 21638 -1288 21698 -258
rect 21758 -1228 21818 -196
rect 21878 -1288 21938 -258
rect 21998 -1228 22058 -196
rect 22118 -350 22184 -196
rect 22118 -414 22119 -350
rect 22183 -414 22184 -350
rect 22118 -430 22184 -414
rect 22118 -494 22119 -430
rect 22183 -494 22184 -430
rect 22118 -510 22184 -494
rect 22118 -574 22119 -510
rect 22183 -574 22184 -510
rect 22118 -590 22184 -574
rect 22118 -654 22119 -590
rect 22183 -654 22184 -590
rect 22118 -670 22184 -654
rect 22118 -734 22119 -670
rect 22183 -734 22184 -670
rect 22118 -750 22184 -734
rect 22118 -814 22119 -750
rect 22183 -814 22184 -750
rect 22118 -830 22184 -814
rect 22118 -894 22119 -830
rect 22183 -894 22184 -830
rect 22118 -910 22184 -894
rect 22118 -974 22119 -910
rect 22183 -974 22184 -910
rect 22118 -990 22184 -974
rect 22118 -1054 22119 -990
rect 22183 -1054 22184 -990
rect 22118 -1070 22184 -1054
rect 22118 -1134 22119 -1070
rect 22183 -1134 22184 -1070
rect 22118 -1224 22184 -1134
rect 22244 -1288 22304 -258
rect 22364 -1228 22424 -196
rect 22484 -1288 22544 -258
rect 22604 -1228 22664 -196
rect 22724 -350 22790 -196
rect 22724 -414 22725 -350
rect 22789 -414 22790 -350
rect 22724 -430 22790 -414
rect 22724 -494 22725 -430
rect 22789 -494 22790 -430
rect 22724 -510 22790 -494
rect 22724 -574 22725 -510
rect 22789 -574 22790 -510
rect 22724 -590 22790 -574
rect 22724 -654 22725 -590
rect 22789 -654 22790 -590
rect 22724 -670 22790 -654
rect 22724 -734 22725 -670
rect 22789 -734 22790 -670
rect 22724 -750 22790 -734
rect 22724 -814 22725 -750
rect 22789 -814 22790 -750
rect 22724 -830 22790 -814
rect 22724 -894 22725 -830
rect 22789 -894 22790 -830
rect 22724 -910 22790 -894
rect 22724 -974 22725 -910
rect 22789 -974 22790 -910
rect 22724 -990 22790 -974
rect 22724 -1054 22725 -990
rect 22789 -1054 22790 -990
rect 22724 -1070 22790 -1054
rect 22724 -1134 22725 -1070
rect 22789 -1134 22790 -1070
rect 22724 -1224 22790 -1134
rect 22850 -1288 22910 -258
rect 22970 -1228 23030 -196
rect 23090 -1288 23150 -258
rect 23210 -1228 23270 -196
rect 23330 -350 23396 -196
rect 23330 -414 23331 -350
rect 23395 -414 23396 -350
rect 23330 -430 23396 -414
rect 23330 -494 23331 -430
rect 23395 -494 23396 -430
rect 23330 -510 23396 -494
rect 23330 -574 23331 -510
rect 23395 -574 23396 -510
rect 23330 -590 23396 -574
rect 23330 -654 23331 -590
rect 23395 -654 23396 -590
rect 23330 -670 23396 -654
rect 23330 -734 23331 -670
rect 23395 -734 23396 -670
rect 23330 -750 23396 -734
rect 23330 -814 23331 -750
rect 23395 -814 23396 -750
rect 23330 -830 23396 -814
rect 23330 -894 23331 -830
rect 23395 -894 23396 -830
rect 23330 -910 23396 -894
rect 23330 -974 23331 -910
rect 23395 -974 23396 -910
rect 23330 -990 23396 -974
rect 23330 -1054 23331 -990
rect 23395 -1054 23396 -990
rect 23330 -1070 23396 -1054
rect 23330 -1134 23331 -1070
rect 23395 -1134 23396 -1070
rect 23330 -1224 23396 -1134
rect 23456 -1288 23516 -258
rect 23576 -1228 23636 -196
rect 23696 -1288 23756 -258
rect 23816 -1228 23876 -196
rect 23936 -350 24002 -196
rect 23936 -414 23937 -350
rect 24001 -414 24002 -350
rect 23936 -430 24002 -414
rect 23936 -494 23937 -430
rect 24001 -494 24002 -430
rect 23936 -510 24002 -494
rect 23936 -574 23937 -510
rect 24001 -574 24002 -510
rect 23936 -590 24002 -574
rect 23936 -654 23937 -590
rect 24001 -654 24002 -590
rect 23936 -670 24002 -654
rect 23936 -734 23937 -670
rect 24001 -734 24002 -670
rect 23936 -750 24002 -734
rect 23936 -814 23937 -750
rect 24001 -814 24002 -750
rect 23936 -830 24002 -814
rect 23936 -894 23937 -830
rect 24001 -894 24002 -830
rect 23936 -910 24002 -894
rect 23936 -974 23937 -910
rect 24001 -974 24002 -910
rect 23936 -990 24002 -974
rect 23936 -1054 23937 -990
rect 24001 -1054 24002 -990
rect 23936 -1070 24002 -1054
rect 23936 -1134 23937 -1070
rect 24001 -1134 24002 -1070
rect 23936 -1224 24002 -1134
rect 24062 -1288 24122 -258
rect 24182 -1228 24242 -196
rect 24302 -1288 24362 -258
rect 24422 -1228 24482 -196
rect 24542 -350 24608 -196
rect 24542 -414 24543 -350
rect 24607 -414 24608 -350
rect 24542 -430 24608 -414
rect 24542 -494 24543 -430
rect 24607 -494 24608 -430
rect 24542 -510 24608 -494
rect 24542 -574 24543 -510
rect 24607 -574 24608 -510
rect 24542 -590 24608 -574
rect 24542 -654 24543 -590
rect 24607 -654 24608 -590
rect 24542 -670 24608 -654
rect 24542 -734 24543 -670
rect 24607 -734 24608 -670
rect 24542 -750 24608 -734
rect 24542 -814 24543 -750
rect 24607 -814 24608 -750
rect 24542 -830 24608 -814
rect 24542 -894 24543 -830
rect 24607 -894 24608 -830
rect 24542 -910 24608 -894
rect 24542 -974 24543 -910
rect 24607 -974 24608 -910
rect 24542 -990 24608 -974
rect 24542 -1054 24543 -990
rect 24607 -1054 24608 -990
rect 24542 -1070 24608 -1054
rect 24542 -1134 24543 -1070
rect 24607 -1134 24608 -1070
rect 24542 -1224 24608 -1134
rect 24668 -1288 24728 -258
rect 24788 -1228 24848 -196
rect 24908 -1288 24968 -258
rect 25028 -1228 25088 -196
rect 25148 -350 25214 -196
rect 25148 -414 25149 -350
rect 25213 -414 25214 -350
rect 25148 -430 25214 -414
rect 25148 -494 25149 -430
rect 25213 -494 25214 -430
rect 25148 -510 25214 -494
rect 25148 -574 25149 -510
rect 25213 -574 25214 -510
rect 25148 -590 25214 -574
rect 25148 -654 25149 -590
rect 25213 -654 25214 -590
rect 25148 -670 25214 -654
rect 25148 -734 25149 -670
rect 25213 -734 25214 -670
rect 25148 -750 25214 -734
rect 25148 -814 25149 -750
rect 25213 -814 25214 -750
rect 25148 -830 25214 -814
rect 25148 -894 25149 -830
rect 25213 -894 25214 -830
rect 25148 -910 25214 -894
rect 25148 -974 25149 -910
rect 25213 -974 25214 -910
rect 25148 -990 25214 -974
rect 25148 -1054 25149 -990
rect 25213 -1054 25214 -990
rect 25148 -1070 25214 -1054
rect 25148 -1134 25149 -1070
rect 25213 -1134 25214 -1070
rect 25148 -1224 25214 -1134
rect 25274 -1288 25334 -258
rect 25394 -1228 25454 -196
rect 25514 -1288 25574 -258
rect 25634 -1228 25694 -196
rect 25754 -350 25820 -196
rect 25754 -414 25755 -350
rect 25819 -414 25820 -350
rect 25754 -430 25820 -414
rect 25754 -494 25755 -430
rect 25819 -494 25820 -430
rect 25754 -510 25820 -494
rect 25754 -574 25755 -510
rect 25819 -574 25820 -510
rect 25754 -590 25820 -574
rect 25754 -654 25755 -590
rect 25819 -654 25820 -590
rect 25754 -670 25820 -654
rect 25754 -734 25755 -670
rect 25819 -734 25820 -670
rect 25754 -750 25820 -734
rect 25754 -814 25755 -750
rect 25819 -814 25820 -750
rect 25754 -830 25820 -814
rect 25754 -894 25755 -830
rect 25819 -894 25820 -830
rect 25754 -910 25820 -894
rect 25754 -974 25755 -910
rect 25819 -974 25820 -910
rect 25754 -990 25820 -974
rect 25754 -1054 25755 -990
rect 25819 -1054 25820 -990
rect 25754 -1070 25820 -1054
rect 25754 -1134 25755 -1070
rect 25819 -1134 25820 -1070
rect 25754 -1224 25820 -1134
rect 25880 -1288 25940 -258
rect 26000 -1228 26060 -196
rect 26120 -1288 26180 -258
rect 26240 -1228 26300 -196
rect 26360 -350 26426 -196
rect 26360 -414 26361 -350
rect 26425 -414 26426 -350
rect 26360 -430 26426 -414
rect 26360 -494 26361 -430
rect 26425 -494 26426 -430
rect 26360 -510 26426 -494
rect 26360 -574 26361 -510
rect 26425 -574 26426 -510
rect 26360 -590 26426 -574
rect 26360 -654 26361 -590
rect 26425 -654 26426 -590
rect 26360 -670 26426 -654
rect 26360 -734 26361 -670
rect 26425 -734 26426 -670
rect 26360 -750 26426 -734
rect 26360 -814 26361 -750
rect 26425 -814 26426 -750
rect 26360 -830 26426 -814
rect 26360 -894 26361 -830
rect 26425 -894 26426 -830
rect 26360 -910 26426 -894
rect 26360 -974 26361 -910
rect 26425 -974 26426 -910
rect 26360 -990 26426 -974
rect 26360 -1054 26361 -990
rect 26425 -1054 26426 -990
rect 26360 -1070 26426 -1054
rect 26360 -1134 26361 -1070
rect 26425 -1134 26426 -1070
rect 26360 -1224 26426 -1134
rect 26486 -1288 26546 -258
rect 26606 -1228 26666 -196
rect 26726 -1288 26786 -258
rect 26846 -1228 26906 -196
rect 26966 -350 27032 -196
rect 26966 -414 26967 -350
rect 27031 -414 27032 -350
rect 26966 -430 27032 -414
rect 26966 -494 26967 -430
rect 27031 -494 27032 -430
rect 26966 -510 27032 -494
rect 26966 -574 26967 -510
rect 27031 -574 27032 -510
rect 26966 -590 27032 -574
rect 26966 -654 26967 -590
rect 27031 -654 27032 -590
rect 26966 -670 27032 -654
rect 26966 -734 26967 -670
rect 27031 -734 27032 -670
rect 26966 -750 27032 -734
rect 26966 -814 26967 -750
rect 27031 -814 27032 -750
rect 26966 -830 27032 -814
rect 26966 -894 26967 -830
rect 27031 -894 27032 -830
rect 26966 -910 27032 -894
rect 26966 -974 26967 -910
rect 27031 -974 27032 -910
rect 26966 -990 27032 -974
rect 26966 -1054 26967 -990
rect 27031 -1054 27032 -990
rect 26966 -1070 27032 -1054
rect 26966 -1134 26967 -1070
rect 27031 -1134 27032 -1070
rect 26966 -1224 27032 -1134
rect 27092 -1288 27152 -258
rect 27212 -1228 27272 -196
rect 27332 -1288 27392 -258
rect 27452 -1228 27512 -196
rect 27572 -350 27638 -196
rect 27572 -414 27573 -350
rect 27637 -414 27638 -350
rect 27572 -430 27638 -414
rect 27572 -494 27573 -430
rect 27637 -494 27638 -430
rect 27572 -510 27638 -494
rect 27572 -574 27573 -510
rect 27637 -574 27638 -510
rect 27572 -590 27638 -574
rect 27572 -654 27573 -590
rect 27637 -654 27638 -590
rect 27572 -670 27638 -654
rect 27572 -734 27573 -670
rect 27637 -734 27638 -670
rect 27572 -750 27638 -734
rect 27572 -814 27573 -750
rect 27637 -814 27638 -750
rect 27572 -830 27638 -814
rect 27572 -894 27573 -830
rect 27637 -894 27638 -830
rect 27572 -910 27638 -894
rect 27572 -974 27573 -910
rect 27637 -974 27638 -910
rect 27572 -990 27638 -974
rect 27572 -1054 27573 -990
rect 27637 -1054 27638 -990
rect 27572 -1070 27638 -1054
rect 27572 -1134 27573 -1070
rect 27637 -1134 27638 -1070
rect 27572 -1224 27638 -1134
rect 27698 -1288 27758 -258
rect 27818 -1228 27878 -196
rect 27938 -1288 27998 -258
rect 28058 -1228 28118 -196
rect 28178 -350 28244 -196
rect 28178 -414 28179 -350
rect 28243 -414 28244 -350
rect 28178 -430 28244 -414
rect 28178 -494 28179 -430
rect 28243 -494 28244 -430
rect 28178 -510 28244 -494
rect 28178 -574 28179 -510
rect 28243 -574 28244 -510
rect 28178 -590 28244 -574
rect 28178 -654 28179 -590
rect 28243 -654 28244 -590
rect 28178 -670 28244 -654
rect 28178 -734 28179 -670
rect 28243 -734 28244 -670
rect 28178 -750 28244 -734
rect 28178 -814 28179 -750
rect 28243 -814 28244 -750
rect 28178 -830 28244 -814
rect 28178 -894 28179 -830
rect 28243 -894 28244 -830
rect 28178 -910 28244 -894
rect 28178 -974 28179 -910
rect 28243 -974 28244 -910
rect 28178 -990 28244 -974
rect 28178 -1054 28179 -990
rect 28243 -1054 28244 -990
rect 28178 -1070 28244 -1054
rect 28178 -1134 28179 -1070
rect 28243 -1134 28244 -1070
rect 28178 -1224 28244 -1134
rect 28304 -1288 28364 -258
rect 28424 -1228 28484 -196
rect 28544 -1288 28604 -258
rect 28664 -1228 28724 -196
rect 28784 -350 28850 -196
rect 28784 -414 28785 -350
rect 28849 -414 28850 -350
rect 28784 -430 28850 -414
rect 28784 -494 28785 -430
rect 28849 -494 28850 -430
rect 28784 -510 28850 -494
rect 28784 -574 28785 -510
rect 28849 -574 28850 -510
rect 28784 -590 28850 -574
rect 28784 -654 28785 -590
rect 28849 -654 28850 -590
rect 28784 -670 28850 -654
rect 28784 -734 28785 -670
rect 28849 -734 28850 -670
rect 28784 -750 28850 -734
rect 28784 -814 28785 -750
rect 28849 -814 28850 -750
rect 28784 -830 28850 -814
rect 28784 -894 28785 -830
rect 28849 -894 28850 -830
rect 28784 -910 28850 -894
rect 28784 -974 28785 -910
rect 28849 -974 28850 -910
rect 28784 -990 28850 -974
rect 28784 -1054 28785 -990
rect 28849 -1054 28850 -990
rect 28784 -1070 28850 -1054
rect 28784 -1134 28785 -1070
rect 28849 -1134 28850 -1070
rect 28784 -1224 28850 -1134
rect 19088 -1290 28850 -1288
rect 19088 -1354 19192 -1290
rect 19256 -1354 19272 -1290
rect 19336 -1354 19352 -1290
rect 19416 -1354 19432 -1290
rect 19496 -1354 19512 -1290
rect 19576 -1354 19592 -1290
rect 19656 -1354 19798 -1290
rect 19862 -1354 19878 -1290
rect 19942 -1354 19958 -1290
rect 20022 -1354 20038 -1290
rect 20102 -1354 20118 -1290
rect 20182 -1354 20198 -1290
rect 20262 -1354 20404 -1290
rect 20468 -1354 20484 -1290
rect 20548 -1354 20564 -1290
rect 20628 -1354 20644 -1290
rect 20708 -1354 20724 -1290
rect 20788 -1354 20804 -1290
rect 20868 -1354 21010 -1290
rect 21074 -1354 21090 -1290
rect 21154 -1354 21170 -1290
rect 21234 -1354 21250 -1290
rect 21314 -1354 21330 -1290
rect 21394 -1354 21410 -1290
rect 21474 -1354 21616 -1290
rect 21680 -1354 21696 -1290
rect 21760 -1354 21776 -1290
rect 21840 -1354 21856 -1290
rect 21920 -1354 21936 -1290
rect 22000 -1354 22016 -1290
rect 22080 -1354 22222 -1290
rect 22286 -1354 22302 -1290
rect 22366 -1354 22382 -1290
rect 22446 -1354 22462 -1290
rect 22526 -1354 22542 -1290
rect 22606 -1354 22622 -1290
rect 22686 -1354 22828 -1290
rect 22892 -1354 22908 -1290
rect 22972 -1354 22988 -1290
rect 23052 -1354 23068 -1290
rect 23132 -1354 23148 -1290
rect 23212 -1354 23228 -1290
rect 23292 -1354 23434 -1290
rect 23498 -1354 23514 -1290
rect 23578 -1354 23594 -1290
rect 23658 -1354 23674 -1290
rect 23738 -1354 23754 -1290
rect 23818 -1354 23834 -1290
rect 23898 -1354 24040 -1290
rect 24104 -1354 24120 -1290
rect 24184 -1354 24200 -1290
rect 24264 -1354 24280 -1290
rect 24344 -1354 24360 -1290
rect 24424 -1354 24440 -1290
rect 24504 -1354 24646 -1290
rect 24710 -1354 24726 -1290
rect 24790 -1354 24806 -1290
rect 24870 -1354 24886 -1290
rect 24950 -1354 24966 -1290
rect 25030 -1354 25046 -1290
rect 25110 -1354 25252 -1290
rect 25316 -1354 25332 -1290
rect 25396 -1354 25412 -1290
rect 25476 -1354 25492 -1290
rect 25556 -1354 25572 -1290
rect 25636 -1354 25652 -1290
rect 25716 -1354 25858 -1290
rect 25922 -1354 25938 -1290
rect 26002 -1354 26018 -1290
rect 26082 -1354 26098 -1290
rect 26162 -1354 26178 -1290
rect 26242 -1354 26258 -1290
rect 26322 -1354 26464 -1290
rect 26528 -1354 26544 -1290
rect 26608 -1354 26624 -1290
rect 26688 -1354 26704 -1290
rect 26768 -1354 26784 -1290
rect 26848 -1354 26864 -1290
rect 26928 -1354 27070 -1290
rect 27134 -1354 27150 -1290
rect 27214 -1354 27230 -1290
rect 27294 -1354 27310 -1290
rect 27374 -1354 27390 -1290
rect 27454 -1354 27470 -1290
rect 27534 -1354 27676 -1290
rect 27740 -1354 27756 -1290
rect 27820 -1354 27836 -1290
rect 27900 -1354 27916 -1290
rect 27980 -1354 27996 -1290
rect 28060 -1354 28076 -1290
rect 28140 -1354 28282 -1290
rect 28346 -1354 28362 -1290
rect 28426 -1354 28442 -1290
rect 28506 -1354 28522 -1290
rect 28586 -1354 28602 -1290
rect 28666 -1354 28682 -1290
rect 28746 -1354 28850 -1290
rect 19088 -1356 28850 -1354
rect 19088 -1510 19154 -1356
rect 19088 -1574 19089 -1510
rect 19153 -1574 19154 -1510
rect 19088 -1590 19154 -1574
rect 19088 -1654 19089 -1590
rect 19153 -1654 19154 -1590
rect 19088 -1670 19154 -1654
rect 19088 -1734 19089 -1670
rect 19153 -1734 19154 -1670
rect 19088 -1750 19154 -1734
rect 19088 -1814 19089 -1750
rect 19153 -1814 19154 -1750
rect 19088 -1830 19154 -1814
rect 19088 -1894 19089 -1830
rect 19153 -1894 19154 -1830
rect 19088 -1910 19154 -1894
rect 19088 -1974 19089 -1910
rect 19153 -1974 19154 -1910
rect 19088 -1990 19154 -1974
rect 19088 -2054 19089 -1990
rect 19153 -2054 19154 -1990
rect 19088 -2070 19154 -2054
rect 19088 -2134 19089 -2070
rect 19153 -2134 19154 -2070
rect 19088 -2150 19154 -2134
rect 19088 -2214 19089 -2150
rect 19153 -2214 19154 -2150
rect 19088 -2230 19154 -2214
rect 19088 -2294 19089 -2230
rect 19153 -2294 19154 -2230
rect 19088 -2384 19154 -2294
rect 19214 -2448 19274 -1418
rect 19334 -2388 19394 -1356
rect 19454 -2448 19514 -1418
rect 19574 -2388 19634 -1356
rect 19694 -1510 19760 -1356
rect 19694 -1574 19695 -1510
rect 19759 -1574 19760 -1510
rect 19694 -1590 19760 -1574
rect 19694 -1654 19695 -1590
rect 19759 -1654 19760 -1590
rect 19694 -1670 19760 -1654
rect 19694 -1734 19695 -1670
rect 19759 -1734 19760 -1670
rect 19694 -1750 19760 -1734
rect 19694 -1814 19695 -1750
rect 19759 -1814 19760 -1750
rect 19694 -1830 19760 -1814
rect 19694 -1894 19695 -1830
rect 19759 -1894 19760 -1830
rect 19694 -1910 19760 -1894
rect 19694 -1974 19695 -1910
rect 19759 -1974 19760 -1910
rect 19694 -1990 19760 -1974
rect 19694 -2054 19695 -1990
rect 19759 -2054 19760 -1990
rect 19694 -2070 19760 -2054
rect 19694 -2134 19695 -2070
rect 19759 -2134 19760 -2070
rect 19694 -2150 19760 -2134
rect 19694 -2214 19695 -2150
rect 19759 -2214 19760 -2150
rect 19694 -2230 19760 -2214
rect 19694 -2294 19695 -2230
rect 19759 -2294 19760 -2230
rect 19694 -2384 19760 -2294
rect 19820 -2448 19880 -1418
rect 19940 -2388 20000 -1356
rect 20060 -2448 20120 -1418
rect 20180 -2388 20240 -1356
rect 20300 -1510 20366 -1356
rect 20300 -1574 20301 -1510
rect 20365 -1574 20366 -1510
rect 20300 -1590 20366 -1574
rect 20300 -1654 20301 -1590
rect 20365 -1654 20366 -1590
rect 20300 -1670 20366 -1654
rect 20300 -1734 20301 -1670
rect 20365 -1734 20366 -1670
rect 20300 -1750 20366 -1734
rect 20300 -1814 20301 -1750
rect 20365 -1814 20366 -1750
rect 20300 -1830 20366 -1814
rect 20300 -1894 20301 -1830
rect 20365 -1894 20366 -1830
rect 20300 -1910 20366 -1894
rect 20300 -1974 20301 -1910
rect 20365 -1974 20366 -1910
rect 20300 -1990 20366 -1974
rect 20300 -2054 20301 -1990
rect 20365 -2054 20366 -1990
rect 20300 -2070 20366 -2054
rect 20300 -2134 20301 -2070
rect 20365 -2134 20366 -2070
rect 20300 -2150 20366 -2134
rect 20300 -2214 20301 -2150
rect 20365 -2214 20366 -2150
rect 20300 -2230 20366 -2214
rect 20300 -2294 20301 -2230
rect 20365 -2294 20366 -2230
rect 20300 -2384 20366 -2294
rect 20426 -2448 20486 -1418
rect 20546 -2388 20606 -1356
rect 20666 -2448 20726 -1418
rect 20786 -2388 20846 -1356
rect 20906 -1510 20972 -1356
rect 20906 -1574 20907 -1510
rect 20971 -1574 20972 -1510
rect 20906 -1590 20972 -1574
rect 20906 -1654 20907 -1590
rect 20971 -1654 20972 -1590
rect 20906 -1670 20972 -1654
rect 20906 -1734 20907 -1670
rect 20971 -1734 20972 -1670
rect 20906 -1750 20972 -1734
rect 20906 -1814 20907 -1750
rect 20971 -1814 20972 -1750
rect 20906 -1830 20972 -1814
rect 20906 -1894 20907 -1830
rect 20971 -1894 20972 -1830
rect 20906 -1910 20972 -1894
rect 20906 -1974 20907 -1910
rect 20971 -1974 20972 -1910
rect 20906 -1990 20972 -1974
rect 20906 -2054 20907 -1990
rect 20971 -2054 20972 -1990
rect 20906 -2070 20972 -2054
rect 20906 -2134 20907 -2070
rect 20971 -2134 20972 -2070
rect 20906 -2150 20972 -2134
rect 20906 -2214 20907 -2150
rect 20971 -2214 20972 -2150
rect 20906 -2230 20972 -2214
rect 20906 -2294 20907 -2230
rect 20971 -2294 20972 -2230
rect 20906 -2384 20972 -2294
rect 21032 -2448 21092 -1418
rect 21152 -2388 21212 -1356
rect 21272 -2448 21332 -1418
rect 21392 -2388 21452 -1356
rect 21512 -1510 21578 -1356
rect 21512 -1574 21513 -1510
rect 21577 -1574 21578 -1510
rect 21512 -1590 21578 -1574
rect 21512 -1654 21513 -1590
rect 21577 -1654 21578 -1590
rect 21512 -1670 21578 -1654
rect 21512 -1734 21513 -1670
rect 21577 -1734 21578 -1670
rect 21512 -1750 21578 -1734
rect 21512 -1814 21513 -1750
rect 21577 -1814 21578 -1750
rect 21512 -1830 21578 -1814
rect 21512 -1894 21513 -1830
rect 21577 -1894 21578 -1830
rect 21512 -1910 21578 -1894
rect 21512 -1974 21513 -1910
rect 21577 -1974 21578 -1910
rect 21512 -1990 21578 -1974
rect 21512 -2054 21513 -1990
rect 21577 -2054 21578 -1990
rect 21512 -2070 21578 -2054
rect 21512 -2134 21513 -2070
rect 21577 -2134 21578 -2070
rect 21512 -2150 21578 -2134
rect 21512 -2214 21513 -2150
rect 21577 -2214 21578 -2150
rect 21512 -2230 21578 -2214
rect 21512 -2294 21513 -2230
rect 21577 -2294 21578 -2230
rect 21512 -2384 21578 -2294
rect 21638 -2448 21698 -1418
rect 21758 -2388 21818 -1356
rect 21878 -2448 21938 -1418
rect 21998 -2388 22058 -1356
rect 22118 -1510 22184 -1356
rect 22118 -1574 22119 -1510
rect 22183 -1574 22184 -1510
rect 22118 -1590 22184 -1574
rect 22118 -1654 22119 -1590
rect 22183 -1654 22184 -1590
rect 22118 -1670 22184 -1654
rect 22118 -1734 22119 -1670
rect 22183 -1734 22184 -1670
rect 22118 -1750 22184 -1734
rect 22118 -1814 22119 -1750
rect 22183 -1814 22184 -1750
rect 22118 -1830 22184 -1814
rect 22118 -1894 22119 -1830
rect 22183 -1894 22184 -1830
rect 22118 -1910 22184 -1894
rect 22118 -1974 22119 -1910
rect 22183 -1974 22184 -1910
rect 22118 -1990 22184 -1974
rect 22118 -2054 22119 -1990
rect 22183 -2054 22184 -1990
rect 22118 -2070 22184 -2054
rect 22118 -2134 22119 -2070
rect 22183 -2134 22184 -2070
rect 22118 -2150 22184 -2134
rect 22118 -2214 22119 -2150
rect 22183 -2214 22184 -2150
rect 22118 -2230 22184 -2214
rect 22118 -2294 22119 -2230
rect 22183 -2294 22184 -2230
rect 22118 -2384 22184 -2294
rect 22244 -2448 22304 -1418
rect 22364 -2388 22424 -1356
rect 22484 -2448 22544 -1418
rect 22604 -2388 22664 -1356
rect 22724 -1510 22790 -1356
rect 22724 -1574 22725 -1510
rect 22789 -1574 22790 -1510
rect 22724 -1590 22790 -1574
rect 22724 -1654 22725 -1590
rect 22789 -1654 22790 -1590
rect 22724 -1670 22790 -1654
rect 22724 -1734 22725 -1670
rect 22789 -1734 22790 -1670
rect 22724 -1750 22790 -1734
rect 22724 -1814 22725 -1750
rect 22789 -1814 22790 -1750
rect 22724 -1830 22790 -1814
rect 22724 -1894 22725 -1830
rect 22789 -1894 22790 -1830
rect 22724 -1910 22790 -1894
rect 22724 -1974 22725 -1910
rect 22789 -1974 22790 -1910
rect 22724 -1990 22790 -1974
rect 22724 -2054 22725 -1990
rect 22789 -2054 22790 -1990
rect 22724 -2070 22790 -2054
rect 22724 -2134 22725 -2070
rect 22789 -2134 22790 -2070
rect 22724 -2150 22790 -2134
rect 22724 -2214 22725 -2150
rect 22789 -2214 22790 -2150
rect 22724 -2230 22790 -2214
rect 22724 -2294 22725 -2230
rect 22789 -2294 22790 -2230
rect 22724 -2384 22790 -2294
rect 22850 -2448 22910 -1418
rect 22970 -2388 23030 -1356
rect 23090 -2448 23150 -1418
rect 23210 -2388 23270 -1356
rect 23330 -1510 23396 -1356
rect 23330 -1574 23331 -1510
rect 23395 -1574 23396 -1510
rect 23330 -1590 23396 -1574
rect 23330 -1654 23331 -1590
rect 23395 -1654 23396 -1590
rect 23330 -1670 23396 -1654
rect 23330 -1734 23331 -1670
rect 23395 -1734 23396 -1670
rect 23330 -1750 23396 -1734
rect 23330 -1814 23331 -1750
rect 23395 -1814 23396 -1750
rect 23330 -1830 23396 -1814
rect 23330 -1894 23331 -1830
rect 23395 -1894 23396 -1830
rect 23330 -1910 23396 -1894
rect 23330 -1974 23331 -1910
rect 23395 -1974 23396 -1910
rect 23330 -1990 23396 -1974
rect 23330 -2054 23331 -1990
rect 23395 -2054 23396 -1990
rect 23330 -2070 23396 -2054
rect 23330 -2134 23331 -2070
rect 23395 -2134 23396 -2070
rect 23330 -2150 23396 -2134
rect 23330 -2214 23331 -2150
rect 23395 -2214 23396 -2150
rect 23330 -2230 23396 -2214
rect 23330 -2294 23331 -2230
rect 23395 -2294 23396 -2230
rect 23330 -2384 23396 -2294
rect 23456 -2448 23516 -1418
rect 23576 -2388 23636 -1356
rect 23696 -2448 23756 -1418
rect 23816 -2388 23876 -1356
rect 23936 -1510 24002 -1356
rect 23936 -1574 23937 -1510
rect 24001 -1574 24002 -1510
rect 23936 -1590 24002 -1574
rect 23936 -1654 23937 -1590
rect 24001 -1654 24002 -1590
rect 23936 -1670 24002 -1654
rect 23936 -1734 23937 -1670
rect 24001 -1734 24002 -1670
rect 23936 -1750 24002 -1734
rect 23936 -1814 23937 -1750
rect 24001 -1814 24002 -1750
rect 23936 -1830 24002 -1814
rect 23936 -1894 23937 -1830
rect 24001 -1894 24002 -1830
rect 23936 -1910 24002 -1894
rect 23936 -1974 23937 -1910
rect 24001 -1974 24002 -1910
rect 23936 -1990 24002 -1974
rect 23936 -2054 23937 -1990
rect 24001 -2054 24002 -1990
rect 23936 -2070 24002 -2054
rect 23936 -2134 23937 -2070
rect 24001 -2134 24002 -2070
rect 23936 -2150 24002 -2134
rect 23936 -2214 23937 -2150
rect 24001 -2214 24002 -2150
rect 23936 -2230 24002 -2214
rect 23936 -2294 23937 -2230
rect 24001 -2294 24002 -2230
rect 23936 -2384 24002 -2294
rect 24062 -2448 24122 -1418
rect 24182 -2388 24242 -1356
rect 24302 -2448 24362 -1418
rect 24422 -2388 24482 -1356
rect 24542 -1510 24608 -1356
rect 24542 -1574 24543 -1510
rect 24607 -1574 24608 -1510
rect 24542 -1590 24608 -1574
rect 24542 -1654 24543 -1590
rect 24607 -1654 24608 -1590
rect 24542 -1670 24608 -1654
rect 24542 -1734 24543 -1670
rect 24607 -1734 24608 -1670
rect 24542 -1750 24608 -1734
rect 24542 -1814 24543 -1750
rect 24607 -1814 24608 -1750
rect 24542 -1830 24608 -1814
rect 24542 -1894 24543 -1830
rect 24607 -1894 24608 -1830
rect 24542 -1910 24608 -1894
rect 24542 -1974 24543 -1910
rect 24607 -1974 24608 -1910
rect 24542 -1990 24608 -1974
rect 24542 -2054 24543 -1990
rect 24607 -2054 24608 -1990
rect 24542 -2070 24608 -2054
rect 24542 -2134 24543 -2070
rect 24607 -2134 24608 -2070
rect 24542 -2150 24608 -2134
rect 24542 -2214 24543 -2150
rect 24607 -2214 24608 -2150
rect 24542 -2230 24608 -2214
rect 24542 -2294 24543 -2230
rect 24607 -2294 24608 -2230
rect 24542 -2384 24608 -2294
rect 24668 -2448 24728 -1418
rect 24788 -2388 24848 -1356
rect 24908 -2448 24968 -1418
rect 25028 -2388 25088 -1356
rect 25148 -1510 25214 -1356
rect 25148 -1574 25149 -1510
rect 25213 -1574 25214 -1510
rect 25148 -1590 25214 -1574
rect 25148 -1654 25149 -1590
rect 25213 -1654 25214 -1590
rect 25148 -1670 25214 -1654
rect 25148 -1734 25149 -1670
rect 25213 -1734 25214 -1670
rect 25148 -1750 25214 -1734
rect 25148 -1814 25149 -1750
rect 25213 -1814 25214 -1750
rect 25148 -1830 25214 -1814
rect 25148 -1894 25149 -1830
rect 25213 -1894 25214 -1830
rect 25148 -1910 25214 -1894
rect 25148 -1974 25149 -1910
rect 25213 -1974 25214 -1910
rect 25148 -1990 25214 -1974
rect 25148 -2054 25149 -1990
rect 25213 -2054 25214 -1990
rect 25148 -2070 25214 -2054
rect 25148 -2134 25149 -2070
rect 25213 -2134 25214 -2070
rect 25148 -2150 25214 -2134
rect 25148 -2214 25149 -2150
rect 25213 -2214 25214 -2150
rect 25148 -2230 25214 -2214
rect 25148 -2294 25149 -2230
rect 25213 -2294 25214 -2230
rect 25148 -2384 25214 -2294
rect 25274 -2448 25334 -1418
rect 25394 -2388 25454 -1356
rect 25514 -2448 25574 -1418
rect 25634 -2388 25694 -1356
rect 25754 -1510 25820 -1356
rect 25754 -1574 25755 -1510
rect 25819 -1574 25820 -1510
rect 25754 -1590 25820 -1574
rect 25754 -1654 25755 -1590
rect 25819 -1654 25820 -1590
rect 25754 -1670 25820 -1654
rect 25754 -1734 25755 -1670
rect 25819 -1734 25820 -1670
rect 25754 -1750 25820 -1734
rect 25754 -1814 25755 -1750
rect 25819 -1814 25820 -1750
rect 25754 -1830 25820 -1814
rect 25754 -1894 25755 -1830
rect 25819 -1894 25820 -1830
rect 25754 -1910 25820 -1894
rect 25754 -1974 25755 -1910
rect 25819 -1974 25820 -1910
rect 25754 -1990 25820 -1974
rect 25754 -2054 25755 -1990
rect 25819 -2054 25820 -1990
rect 25754 -2070 25820 -2054
rect 25754 -2134 25755 -2070
rect 25819 -2134 25820 -2070
rect 25754 -2150 25820 -2134
rect 25754 -2214 25755 -2150
rect 25819 -2214 25820 -2150
rect 25754 -2230 25820 -2214
rect 25754 -2294 25755 -2230
rect 25819 -2294 25820 -2230
rect 25754 -2384 25820 -2294
rect 25880 -2448 25940 -1418
rect 26000 -2388 26060 -1356
rect 26120 -2448 26180 -1418
rect 26240 -2388 26300 -1356
rect 26360 -1510 26426 -1356
rect 26360 -1574 26361 -1510
rect 26425 -1574 26426 -1510
rect 26360 -1590 26426 -1574
rect 26360 -1654 26361 -1590
rect 26425 -1654 26426 -1590
rect 26360 -1670 26426 -1654
rect 26360 -1734 26361 -1670
rect 26425 -1734 26426 -1670
rect 26360 -1750 26426 -1734
rect 26360 -1814 26361 -1750
rect 26425 -1814 26426 -1750
rect 26360 -1830 26426 -1814
rect 26360 -1894 26361 -1830
rect 26425 -1894 26426 -1830
rect 26360 -1910 26426 -1894
rect 26360 -1974 26361 -1910
rect 26425 -1974 26426 -1910
rect 26360 -1990 26426 -1974
rect 26360 -2054 26361 -1990
rect 26425 -2054 26426 -1990
rect 26360 -2070 26426 -2054
rect 26360 -2134 26361 -2070
rect 26425 -2134 26426 -2070
rect 26360 -2150 26426 -2134
rect 26360 -2214 26361 -2150
rect 26425 -2214 26426 -2150
rect 26360 -2230 26426 -2214
rect 26360 -2294 26361 -2230
rect 26425 -2294 26426 -2230
rect 26360 -2384 26426 -2294
rect 26486 -2448 26546 -1418
rect 26606 -2388 26666 -1356
rect 26726 -2448 26786 -1418
rect 26846 -2388 26906 -1356
rect 26966 -1510 27032 -1356
rect 26966 -1574 26967 -1510
rect 27031 -1574 27032 -1510
rect 26966 -1590 27032 -1574
rect 26966 -1654 26967 -1590
rect 27031 -1654 27032 -1590
rect 26966 -1670 27032 -1654
rect 26966 -1734 26967 -1670
rect 27031 -1734 27032 -1670
rect 26966 -1750 27032 -1734
rect 26966 -1814 26967 -1750
rect 27031 -1814 27032 -1750
rect 26966 -1830 27032 -1814
rect 26966 -1894 26967 -1830
rect 27031 -1894 27032 -1830
rect 26966 -1910 27032 -1894
rect 26966 -1974 26967 -1910
rect 27031 -1974 27032 -1910
rect 26966 -1990 27032 -1974
rect 26966 -2054 26967 -1990
rect 27031 -2054 27032 -1990
rect 26966 -2070 27032 -2054
rect 26966 -2134 26967 -2070
rect 27031 -2134 27032 -2070
rect 26966 -2150 27032 -2134
rect 26966 -2214 26967 -2150
rect 27031 -2214 27032 -2150
rect 26966 -2230 27032 -2214
rect 26966 -2294 26967 -2230
rect 27031 -2294 27032 -2230
rect 26966 -2384 27032 -2294
rect 27092 -2448 27152 -1418
rect 27212 -2388 27272 -1356
rect 27332 -2448 27392 -1418
rect 27452 -2388 27512 -1356
rect 27572 -1510 27638 -1356
rect 27572 -1574 27573 -1510
rect 27637 -1574 27638 -1510
rect 27572 -1590 27638 -1574
rect 27572 -1654 27573 -1590
rect 27637 -1654 27638 -1590
rect 27572 -1670 27638 -1654
rect 27572 -1734 27573 -1670
rect 27637 -1734 27638 -1670
rect 27572 -1750 27638 -1734
rect 27572 -1814 27573 -1750
rect 27637 -1814 27638 -1750
rect 27572 -1830 27638 -1814
rect 27572 -1894 27573 -1830
rect 27637 -1894 27638 -1830
rect 27572 -1910 27638 -1894
rect 27572 -1974 27573 -1910
rect 27637 -1974 27638 -1910
rect 27572 -1990 27638 -1974
rect 27572 -2054 27573 -1990
rect 27637 -2054 27638 -1990
rect 27572 -2070 27638 -2054
rect 27572 -2134 27573 -2070
rect 27637 -2134 27638 -2070
rect 27572 -2150 27638 -2134
rect 27572 -2214 27573 -2150
rect 27637 -2214 27638 -2150
rect 27572 -2230 27638 -2214
rect 27572 -2294 27573 -2230
rect 27637 -2294 27638 -2230
rect 27572 -2384 27638 -2294
rect 27698 -2448 27758 -1418
rect 27818 -2388 27878 -1356
rect 27938 -2448 27998 -1418
rect 28058 -2388 28118 -1356
rect 28178 -1510 28244 -1356
rect 28178 -1574 28179 -1510
rect 28243 -1574 28244 -1510
rect 28178 -1590 28244 -1574
rect 28178 -1654 28179 -1590
rect 28243 -1654 28244 -1590
rect 28178 -1670 28244 -1654
rect 28178 -1734 28179 -1670
rect 28243 -1734 28244 -1670
rect 28178 -1750 28244 -1734
rect 28178 -1814 28179 -1750
rect 28243 -1814 28244 -1750
rect 28178 -1830 28244 -1814
rect 28178 -1894 28179 -1830
rect 28243 -1894 28244 -1830
rect 28178 -1910 28244 -1894
rect 28178 -1974 28179 -1910
rect 28243 -1974 28244 -1910
rect 28178 -1990 28244 -1974
rect 28178 -2054 28179 -1990
rect 28243 -2054 28244 -1990
rect 28178 -2070 28244 -2054
rect 28178 -2134 28179 -2070
rect 28243 -2134 28244 -2070
rect 28178 -2150 28244 -2134
rect 28178 -2214 28179 -2150
rect 28243 -2214 28244 -2150
rect 28178 -2230 28244 -2214
rect 28178 -2294 28179 -2230
rect 28243 -2294 28244 -2230
rect 28178 -2384 28244 -2294
rect 28304 -2448 28364 -1418
rect 28424 -2388 28484 -1356
rect 28544 -2448 28604 -1418
rect 28664 -2388 28724 -1356
rect 28784 -1510 28850 -1356
rect 28784 -1574 28785 -1510
rect 28849 -1574 28850 -1510
rect 28784 -1590 28850 -1574
rect 28784 -1654 28785 -1590
rect 28849 -1654 28850 -1590
rect 28784 -1670 28850 -1654
rect 28784 -1734 28785 -1670
rect 28849 -1734 28850 -1670
rect 28784 -1750 28850 -1734
rect 28784 -1814 28785 -1750
rect 28849 -1814 28850 -1750
rect 28784 -1830 28850 -1814
rect 28784 -1894 28785 -1830
rect 28849 -1894 28850 -1830
rect 28784 -1910 28850 -1894
rect 28784 -1974 28785 -1910
rect 28849 -1974 28850 -1910
rect 28784 -1990 28850 -1974
rect 28784 -2054 28785 -1990
rect 28849 -2054 28850 -1990
rect 28784 -2070 28850 -2054
rect 28784 -2134 28785 -2070
rect 28849 -2134 28850 -2070
rect 28784 -2150 28850 -2134
rect 28784 -2214 28785 -2150
rect 28849 -2214 28850 -2150
rect 28784 -2230 28850 -2214
rect 28784 -2294 28785 -2230
rect 28849 -2294 28850 -2230
rect 28784 -2384 28850 -2294
rect 19088 -2450 28850 -2448
rect 19088 -2514 19192 -2450
rect 19256 -2514 19272 -2450
rect 19336 -2514 19352 -2450
rect 19416 -2514 19432 -2450
rect 19496 -2514 19512 -2450
rect 19576 -2514 19592 -2450
rect 19656 -2514 19798 -2450
rect 19862 -2514 19878 -2450
rect 19942 -2514 19958 -2450
rect 20022 -2514 20038 -2450
rect 20102 -2514 20118 -2450
rect 20182 -2514 20198 -2450
rect 20262 -2514 20404 -2450
rect 20468 -2514 20484 -2450
rect 20548 -2514 20564 -2450
rect 20628 -2514 20644 -2450
rect 20708 -2514 20724 -2450
rect 20788 -2514 20804 -2450
rect 20868 -2514 21010 -2450
rect 21074 -2514 21090 -2450
rect 21154 -2514 21170 -2450
rect 21234 -2514 21250 -2450
rect 21314 -2514 21330 -2450
rect 21394 -2514 21410 -2450
rect 21474 -2514 21616 -2450
rect 21680 -2514 21696 -2450
rect 21760 -2514 21776 -2450
rect 21840 -2514 21856 -2450
rect 21920 -2514 21936 -2450
rect 22000 -2514 22016 -2450
rect 22080 -2514 22222 -2450
rect 22286 -2514 22302 -2450
rect 22366 -2514 22382 -2450
rect 22446 -2514 22462 -2450
rect 22526 -2514 22542 -2450
rect 22606 -2514 22622 -2450
rect 22686 -2514 22828 -2450
rect 22892 -2514 22908 -2450
rect 22972 -2514 22988 -2450
rect 23052 -2514 23068 -2450
rect 23132 -2514 23148 -2450
rect 23212 -2514 23228 -2450
rect 23292 -2514 23434 -2450
rect 23498 -2514 23514 -2450
rect 23578 -2514 23594 -2450
rect 23658 -2514 23674 -2450
rect 23738 -2514 23754 -2450
rect 23818 -2514 23834 -2450
rect 23898 -2514 24040 -2450
rect 24104 -2514 24120 -2450
rect 24184 -2514 24200 -2450
rect 24264 -2514 24280 -2450
rect 24344 -2514 24360 -2450
rect 24424 -2514 24440 -2450
rect 24504 -2514 24646 -2450
rect 24710 -2514 24726 -2450
rect 24790 -2514 24806 -2450
rect 24870 -2514 24886 -2450
rect 24950 -2514 24966 -2450
rect 25030 -2514 25046 -2450
rect 25110 -2514 25252 -2450
rect 25316 -2514 25332 -2450
rect 25396 -2514 25412 -2450
rect 25476 -2514 25492 -2450
rect 25556 -2514 25572 -2450
rect 25636 -2514 25652 -2450
rect 25716 -2514 25858 -2450
rect 25922 -2514 25938 -2450
rect 26002 -2514 26018 -2450
rect 26082 -2514 26098 -2450
rect 26162 -2514 26178 -2450
rect 26242 -2514 26258 -2450
rect 26322 -2514 26464 -2450
rect 26528 -2514 26544 -2450
rect 26608 -2514 26624 -2450
rect 26688 -2514 26704 -2450
rect 26768 -2514 26784 -2450
rect 26848 -2514 26864 -2450
rect 26928 -2514 27070 -2450
rect 27134 -2514 27150 -2450
rect 27214 -2514 27230 -2450
rect 27294 -2514 27310 -2450
rect 27374 -2514 27390 -2450
rect 27454 -2514 27470 -2450
rect 27534 -2514 27676 -2450
rect 27740 -2514 27756 -2450
rect 27820 -2514 27836 -2450
rect 27900 -2514 27916 -2450
rect 27980 -2514 27996 -2450
rect 28060 -2514 28076 -2450
rect 28140 -2514 28282 -2450
rect 28346 -2514 28362 -2450
rect 28426 -2514 28442 -2450
rect 28506 -2514 28522 -2450
rect 28586 -2514 28602 -2450
rect 28666 -2514 28682 -2450
rect 28746 -2514 28850 -2450
rect 19088 -2516 28850 -2514
<< labels >>
flabel pwell 19408 -2100 19434 -2068 0 FreeSans 160 0 0 0 x1[0].SUB
flabel metal4 19350 -1766 19376 -1734 0 FreeSans 320 0 0 0 x1[0].CBOT
flabel metal4 19468 -2356 19494 -2324 0 FreeSans 320 0 0 0 x1[0].CTOP
flabel pwell 21832 -2100 21858 -2068 0 FreeSans 160 0 0 0 x1[8].SUB
flabel metal4 21774 -1766 21800 -1734 0 FreeSans 320 0 0 0 x1[8].CBOT
flabel metal4 21892 -2356 21918 -2324 0 FreeSans 320 0 0 0 x1[8].CTOP
flabel pwell 21226 -2100 21252 -2068 0 FreeSans 160 0 0 0 x1[6].SUB
flabel metal4 21168 -1766 21194 -1734 0 FreeSans 320 0 0 0 x1[6].CBOT
flabel metal4 21286 -2356 21312 -2324 0 FreeSans 320 0 0 0 x1[6].CTOP
flabel pwell 20620 -2100 20646 -2068 0 FreeSans 160 0 0 0 x1[4].SUB
flabel metal4 20562 -1766 20588 -1734 0 FreeSans 320 0 0 0 x1[4].CBOT
flabel metal4 20680 -2356 20706 -2324 0 FreeSans 320 0 0 0 x1[4].CTOP
flabel pwell 20014 -2100 20040 -2068 0 FreeSans 160 0 0 0 x1[2].SUB
flabel metal4 19956 -1766 19982 -1734 0 FreeSans 320 0 0 0 x1[2].CBOT
flabel metal4 20074 -2356 20100 -2324 0 FreeSans 320 0 0 0 x1[2].CTOP
flabel pwell 19408 -940 19434 -908 0 FreeSans 160 0 0 0 x1[1].SUB
flabel metal4 19350 -606 19376 -574 0 FreeSans 320 0 0 0 x1[1].CBOT
flabel metal4 19468 -1196 19494 -1164 0 FreeSans 320 0 0 0 x1[1].CTOP
flabel pwell 21832 -940 21858 -908 0 FreeSans 160 0 0 0 x1[9].SUB
flabel metal4 21774 -606 21800 -574 0 FreeSans 320 0 0 0 x1[9].CBOT
flabel metal4 21892 -1196 21918 -1164 0 FreeSans 320 0 0 0 x1[9].CTOP
flabel pwell 21226 -940 21252 -908 0 FreeSans 160 0 0 0 x1[7].SUB
flabel metal4 21168 -606 21194 -574 0 FreeSans 320 0 0 0 x1[7].CBOT
flabel metal4 21286 -1196 21312 -1164 0 FreeSans 320 0 0 0 x1[7].CTOP
flabel pwell 20620 -940 20646 -908 0 FreeSans 160 0 0 0 x1[5].SUB
flabel metal4 20562 -606 20588 -574 0 FreeSans 320 0 0 0 x1[5].CBOT
flabel metal4 20680 -1196 20706 -1164 0 FreeSans 320 0 0 0 x1[5].CTOP
flabel pwell 20014 -940 20040 -908 0 FreeSans 160 0 0 0 x1[3].SUB
flabel metal4 19956 -606 19982 -574 0 FreeSans 320 0 0 0 x1[3].CBOT
flabel metal4 20074 -1196 20100 -1164 0 FreeSans 320 0 0 0 x1[3].CTOP
flabel pwell 24256 -2100 24282 -2068 0 FreeSans 160 0 0 0 x1[16].SUB
flabel metal4 24198 -1766 24224 -1734 0 FreeSans 320 0 0 0 x1[16].CBOT
flabel metal4 24316 -2356 24342 -2324 0 FreeSans 320 0 0 0 x1[16].CTOP
flabel pwell 23650 -2100 23676 -2068 0 FreeSans 160 0 0 0 x1[14].SUB
flabel metal4 23592 -1766 23618 -1734 0 FreeSans 320 0 0 0 x1[14].CBOT
flabel metal4 23710 -2356 23736 -2324 0 FreeSans 320 0 0 0 x1[14].CTOP
flabel pwell 23044 -2100 23070 -2068 0 FreeSans 160 0 0 0 x1[12].SUB
flabel metal4 22986 -1766 23012 -1734 0 FreeSans 320 0 0 0 x1[12].CBOT
flabel metal4 23104 -2356 23130 -2324 0 FreeSans 320 0 0 0 x1[12].CTOP
flabel pwell 22438 -2100 22464 -2068 0 FreeSans 160 0 0 0 x1[10].SUB
flabel metal4 22380 -1766 22406 -1734 0 FreeSans 320 0 0 0 x1[10].CBOT
flabel metal4 22498 -2356 22524 -2324 0 FreeSans 320 0 0 0 x1[10].CTOP
flabel pwell 26074 -2100 26100 -2068 0 FreeSans 160 0 0 0 x1[22].SUB
flabel metal4 26016 -1766 26042 -1734 0 FreeSans 320 0 0 0 x1[22].CBOT
flabel metal4 26134 -2356 26160 -2324 0 FreeSans 320 0 0 0 x1[22].CTOP
flabel pwell 25468 -2100 25494 -2068 0 FreeSans 160 0 0 0 x1[20].SUB
flabel metal4 25410 -1766 25436 -1734 0 FreeSans 320 0 0 0 x1[20].CBOT
flabel metal4 25528 -2356 25554 -2324 0 FreeSans 320 0 0 0 x1[20].CTOP
flabel pwell 24862 -2100 24888 -2068 0 FreeSans 160 0 0 0 x1[18].SUB
flabel metal4 24804 -1766 24830 -1734 0 FreeSans 320 0 0 0 x1[18].CBOT
flabel metal4 24922 -2356 24948 -2324 0 FreeSans 320 0 0 0 x1[18].CTOP
flabel pwell 28498 -2100 28524 -2068 0 FreeSans 160 0 0 0 x1[30].SUB
flabel metal4 28440 -1766 28466 -1734 0 FreeSans 320 0 0 0 x1[30].CBOT
flabel metal4 28558 -2356 28584 -2324 0 FreeSans 320 0 0 0 x1[30].CTOP
flabel pwell 27892 -2100 27918 -2068 0 FreeSans 160 0 0 0 x1[28].SUB
flabel metal4 27834 -1766 27860 -1734 0 FreeSans 320 0 0 0 x1[28].CBOT
flabel metal4 27952 -2356 27978 -2324 0 FreeSans 320 0 0 0 x1[28].CTOP
flabel pwell 27286 -2100 27312 -2068 0 FreeSans 160 0 0 0 x1[26].SUB
flabel metal4 27228 -1766 27254 -1734 0 FreeSans 320 0 0 0 x1[26].CBOT
flabel metal4 27346 -2356 27372 -2324 0 FreeSans 320 0 0 0 x1[26].CTOP
flabel pwell 26680 -2100 26706 -2068 0 FreeSans 160 0 0 0 x1[24].SUB
flabel metal4 26622 -1766 26648 -1734 0 FreeSans 320 0 0 0 x1[24].CBOT
flabel metal4 26740 -2356 26766 -2324 0 FreeSans 320 0 0 0 x1[24].CTOP
flabel pwell 24256 -940 24282 -908 0 FreeSans 160 0 0 0 x1[17].SUB
flabel metal4 24198 -606 24224 -574 0 FreeSans 320 0 0 0 x1[17].CBOT
flabel metal4 24316 -1196 24342 -1164 0 FreeSans 320 0 0 0 x1[17].CTOP
flabel pwell 23650 -940 23676 -908 0 FreeSans 160 0 0 0 x1[15].SUB
flabel metal4 23592 -606 23618 -574 0 FreeSans 320 0 0 0 x1[15].CBOT
flabel metal4 23710 -1196 23736 -1164 0 FreeSans 320 0 0 0 x1[15].CTOP
flabel pwell 23044 -940 23070 -908 0 FreeSans 160 0 0 0 x1[13].SUB
flabel metal4 22986 -606 23012 -574 0 FreeSans 320 0 0 0 x1[13].CBOT
flabel metal4 23104 -1196 23130 -1164 0 FreeSans 320 0 0 0 x1[13].CTOP
flabel pwell 22438 -940 22464 -908 0 FreeSans 160 0 0 0 x1[11].SUB
flabel metal4 22380 -606 22406 -574 0 FreeSans 320 0 0 0 x1[11].CBOT
flabel metal4 22498 -1196 22524 -1164 0 FreeSans 320 0 0 0 x1[11].CTOP
flabel pwell 26074 -940 26100 -908 0 FreeSans 160 0 0 0 x1[23].SUB
flabel metal4 26016 -606 26042 -574 0 FreeSans 320 0 0 0 x1[23].CBOT
flabel metal4 26134 -1196 26160 -1164 0 FreeSans 320 0 0 0 x1[23].CTOP
flabel pwell 25468 -940 25494 -908 0 FreeSans 160 0 0 0 x1[21].SUB
flabel metal4 25410 -606 25436 -574 0 FreeSans 320 0 0 0 x1[21].CBOT
flabel metal4 25528 -1196 25554 -1164 0 FreeSans 320 0 0 0 x1[21].CTOP
flabel pwell 24862 -940 24888 -908 0 FreeSans 160 0 0 0 x1[19].SUB
flabel metal4 24804 -606 24830 -574 0 FreeSans 320 0 0 0 x1[19].CBOT
flabel metal4 24922 -1196 24948 -1164 0 FreeSans 320 0 0 0 x1[19].CTOP
flabel pwell 28498 -940 28524 -908 0 FreeSans 160 0 0 0 x1[31].SUB
flabel metal4 28440 -606 28466 -574 0 FreeSans 320 0 0 0 x1[31].CBOT
flabel metal4 28558 -1196 28584 -1164 0 FreeSans 320 0 0 0 x1[31].CTOP
flabel pwell 27892 -940 27918 -908 0 FreeSans 160 0 0 0 x1[29].SUB
flabel metal4 27834 -606 27860 -574 0 FreeSans 320 0 0 0 x1[29].CBOT
flabel metal4 27952 -1196 27978 -1164 0 FreeSans 320 0 0 0 x1[29].CTOP
flabel pwell 27286 -940 27312 -908 0 FreeSans 160 0 0 0 x1[27].SUB
flabel metal4 27228 -606 27254 -574 0 FreeSans 320 0 0 0 x1[27].CBOT
flabel metal4 27346 -1196 27372 -1164 0 FreeSans 320 0 0 0 x1[27].CTOP
flabel pwell 26680 -940 26706 -908 0 FreeSans 160 0 0 0 x1[25].SUB
flabel metal4 26622 -606 26648 -574 0 FreeSans 320 0 0 0 x1[25].CBOT
flabel metal4 26740 -1196 26766 -1164 0 FreeSans 320 0 0 0 x1[25].CTOP
flabel pwell 23654 -1110 23676 -1070 0 FreeSans 160 0 0 0 SUB
port 3 nsew
<< end >>
