magic
tech sky130A
magscale 1 2
timestamp 1697710383
<< nwell >>
rect -311 -303 311 303
<< pmos >>
rect -111 -84 -81 84
rect -15 -84 15 84
rect 81 -84 111 84
<< pdiff >>
rect -173 72 -111 84
rect -173 -72 -161 72
rect -127 -72 -111 72
rect -173 -84 -111 -72
rect -81 72 -15 84
rect -81 -72 -65 72
rect -31 -72 -15 72
rect -81 -84 -15 -72
rect 15 72 81 84
rect 15 -72 31 72
rect 65 -72 81 72
rect 15 -84 81 -72
rect 111 72 173 84
rect 111 -72 127 72
rect 161 -72 173 72
rect 111 -84 173 -72
<< pdiffc >>
rect -161 -72 -127 72
rect -65 -72 -31 72
rect 31 -72 65 72
rect 127 -72 161 72
<< poly >>
rect -111 84 -81 110
rect -15 84 15 115
rect 81 84 111 110
rect -111 -99 -81 -84
rect -15 -99 15 -84
rect 81 -99 111 -84
rect -111 -129 111 -99
<< locali >>
rect -161 72 -127 88
rect -161 -88 -127 -72
rect -65 72 -31 88
rect -65 -88 -31 -72
rect 31 72 65 88
rect 31 -88 65 -72
rect 127 72 161 88
rect 127 -88 161 -72
<< viali >>
rect -161 -72 -127 72
rect -65 -72 -31 72
rect 31 -72 65 72
rect 127 -72 161 72
<< metal1 >>
rect -167 72 -121 84
rect -167 -72 -161 72
rect -127 -72 -121 72
rect -167 -84 -121 -72
rect -71 72 -25 84
rect -71 -72 -65 72
rect -31 -72 -25 72
rect -71 -84 -25 -72
rect 25 72 71 84
rect 25 -72 31 72
rect 65 -72 71 72
rect 25 -84 71 -72
rect 121 72 167 84
rect 121 -72 127 72
rect 161 -72 167 72
rect 121 -84 167 -72
<< properties >>
string FIXED_BBOX -258 -250 258 250
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.84 l 0.15 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
