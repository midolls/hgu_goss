magic
tech sky130A
magscale 1 2
timestamp 1696942209
<< error_s >>
rect 4760 -700 4818 -694
rect 4760 -734 4772 -700
rect 4760 -740 4818 -734
rect 718 -800 896 -766
rect 656 -904 714 -898
rect 656 -938 668 -904
rect 656 -944 714 -938
rect 656 -1432 714 -1426
rect 656 -1466 668 -1432
rect 656 -1472 714 -1466
rect 972 -1604 1150 -800
rect 1446 -916 1648 -784
rect 2480 -904 2538 -898
rect 1446 -922 1686 -916
rect 1154 -938 1212 -932
rect 1154 -972 1166 -938
rect 1446 -956 1648 -922
rect 2480 -938 2492 -904
rect 2480 -944 2538 -938
rect 1446 -962 1686 -956
rect 1154 -978 1212 -972
rect 1446 -1444 1648 -962
rect 2480 -1432 2538 -1426
rect 1446 -1450 1686 -1444
rect 1154 -1466 1212 -1460
rect 1154 -1500 1166 -1466
rect 1446 -1484 1648 -1450
rect 2480 -1466 2492 -1432
rect 2480 -1472 2538 -1466
rect 1446 -1490 1686 -1484
rect 1154 -1506 1212 -1500
rect 1446 -1622 1648 -1490
rect 2874 -1588 2974 -750
rect 3228 -776 3296 -750
rect 3056 -888 3114 -882
rect 3056 -922 3068 -888
rect 3056 -928 3114 -922
rect 3056 -1416 3114 -1410
rect 3056 -1450 3068 -1416
rect 3056 -1456 3114 -1450
rect 3482 -1588 3550 -776
rect 3664 -914 3722 -908
rect 3664 -948 3676 -914
rect 3664 -954 3722 -948
rect 4760 -996 4818 -990
rect 4760 -1030 4772 -996
rect 4760 -1036 4818 -1030
rect 5250 -1066 5254 -494
rect 6542 -534 6646 -516
rect 5532 -632 5590 -626
rect 5532 -666 5544 -632
rect 6406 -654 6464 -648
rect 5532 -672 5590 -666
rect 6406 -688 6418 -654
rect 6406 -694 6464 -688
rect 5436 -894 5494 -888
rect 5628 -894 5686 -888
rect 5436 -928 5448 -894
rect 5628 -928 5640 -894
rect 5436 -934 5494 -928
rect 5628 -934 5686 -928
rect 6406 -950 6464 -944
rect 6406 -984 6418 -950
rect 6406 -990 6464 -984
rect 5296 -1066 5718 -1058
rect 6796 -1122 6900 -534
rect 6978 -672 7036 -666
rect 6978 -706 6990 -672
rect 6978 -712 7036 -706
rect 6978 -968 7036 -962
rect 6978 -1002 6990 -968
rect 6978 -1008 7036 -1002
rect 5478 -1196 5536 -1190
rect 5478 -1230 5490 -1196
rect 5478 -1236 5536 -1230
rect 9906 -1246 9964 -1240
rect 9906 -1280 9918 -1246
rect 9906 -1286 9964 -1280
rect 4742 -1318 4800 -1312
rect 4742 -1352 4754 -1318
rect 4742 -1358 4800 -1352
rect 6430 -1422 6488 -1416
rect 3664 -1442 3722 -1436
rect 3664 -1476 3676 -1442
rect 6430 -1456 6442 -1422
rect 6430 -1462 6488 -1456
rect 7024 -1470 7082 -1464
rect 3664 -1482 3722 -1476
rect 5478 -1506 5536 -1500
rect 7024 -1504 7036 -1470
rect 4742 -1512 4800 -1506
rect 4742 -1546 4754 -1512
rect 5478 -1540 5490 -1506
rect 7024 -1510 7082 -1504
rect 5478 -1546 5536 -1540
rect 9906 -1542 9964 -1536
rect 4742 -1552 4800 -1546
rect 9906 -1576 9918 -1542
rect 9906 -1582 9964 -1576
rect 10318 -1644 10400 -1072
rect 10600 -1210 10658 -1204
rect 10600 -1244 10612 -1210
rect 10600 -1250 10658 -1244
rect 10504 -1472 10562 -1466
rect 10696 -1472 10754 -1466
rect 10504 -1506 10516 -1472
rect 10696 -1506 10708 -1472
rect 10504 -1512 10562 -1506
rect 10696 -1512 10754 -1506
rect 6430 -1700 6488 -1694
rect 6430 -1734 6442 -1700
rect 6430 -1740 6488 -1734
rect 7024 -1748 7082 -1742
rect 7024 -1782 7036 -1748
rect 7024 -1788 7082 -1782
rect 10536 -1802 10594 -1796
rect 10536 -1836 10548 -1802
rect 10536 -1842 10594 -1836
rect 9930 -1884 9988 -1878
rect 9930 -1918 9942 -1884
rect 9930 -1924 9988 -1918
rect 4704 -2148 4762 -2142
rect 4704 -2182 4716 -2148
rect 4704 -2188 4762 -2182
rect 2912 -2370 2970 -2364
rect 2912 -2404 2924 -2370
rect 2912 -2410 2970 -2404
rect 1512 -2430 1570 -2424
rect 2194 -2430 2252 -2424
rect 1512 -2464 1524 -2430
rect 2194 -2464 2206 -2430
rect 4704 -2444 4762 -2438
rect 1512 -2470 1570 -2464
rect 2194 -2470 2252 -2464
rect 4704 -2478 4716 -2444
rect 4704 -2484 4762 -2478
rect 5192 -2566 5198 -1994
rect 7614 -2064 7672 -2058
rect 6812 -2082 6870 -2076
rect 6812 -2116 6824 -2082
rect 7614 -2098 7626 -2064
rect 9930 -2078 9988 -2072
rect 7614 -2104 7672 -2098
rect 9930 -2112 9942 -2078
rect 10536 -2112 10594 -2106
rect 6812 -2122 6870 -2116
rect 9930 -2118 9988 -2112
rect 5474 -2132 5532 -2126
rect 5474 -2166 5486 -2132
rect 10536 -2146 10548 -2112
rect 10536 -2152 10594 -2146
rect 5474 -2172 5532 -2166
rect 8484 -2180 8542 -2174
rect 8484 -2214 8496 -2180
rect 8484 -2220 8542 -2214
rect 7614 -2360 7672 -2354
rect 6812 -2378 6870 -2372
rect 5378 -2394 5436 -2388
rect 5570 -2394 5628 -2388
rect 5378 -2428 5390 -2394
rect 5570 -2428 5582 -2394
rect 6812 -2412 6824 -2378
rect 7614 -2394 7626 -2360
rect 7614 -2400 7672 -2394
rect 6812 -2418 6870 -2412
rect 5378 -2434 5436 -2428
rect 5570 -2434 5628 -2428
rect 8484 -2476 8542 -2470
rect 8484 -2510 8496 -2476
rect 8484 -2516 8542 -2510
rect 3588 -2588 3646 -2582
rect 3780 -2588 3838 -2582
rect 3588 -2622 3600 -2588
rect 3780 -2622 3792 -2588
rect 3588 -2628 3646 -2622
rect 3780 -2628 3838 -2622
rect 792 -2654 850 -2648
rect 984 -2654 1042 -2648
rect 792 -2688 804 -2654
rect 984 -2688 996 -2654
rect 792 -2694 850 -2688
rect 984 -2694 1042 -2688
rect 7262 -2812 7320 -2806
rect 10030 -2808 10216 -2752
rect 5474 -2822 5532 -2816
rect 4704 -2854 4762 -2848
rect 4704 -2888 4716 -2854
rect 5474 -2856 5486 -2822
rect 7262 -2846 7274 -2812
rect 7262 -2852 7320 -2846
rect 5474 -2862 5532 -2856
rect 4704 -2894 4762 -2888
rect 9976 -2890 10034 -2884
rect 8484 -2928 8542 -2922
rect 9976 -2924 9988 -2890
rect 8484 -2962 8496 -2928
rect 9976 -2930 10034 -2924
rect 8484 -2968 8542 -2962
rect 4704 -3048 4762 -3042
rect 4704 -3082 4716 -3048
rect 4704 -3088 4762 -3082
rect 7262 -3090 7320 -3084
rect 3492 -3098 3550 -3092
rect 3684 -3098 3742 -3092
rect 3492 -3132 3504 -3098
rect 3684 -3132 3696 -3098
rect 7262 -3124 7274 -3090
rect 8484 -3122 8542 -3116
rect 5474 -3132 5532 -3126
rect 7262 -3130 7320 -3124
rect 3492 -3138 3550 -3132
rect 3684 -3138 3742 -3132
rect 696 -3164 754 -3158
rect 888 -3164 946 -3158
rect 696 -3198 708 -3164
rect 888 -3198 900 -3164
rect 5474 -3166 5486 -3132
rect 8484 -3156 8496 -3122
rect 8484 -3162 8542 -3156
rect 5474 -3172 5532 -3166
rect 9976 -3186 10034 -3180
rect 696 -3204 754 -3198
rect 888 -3204 946 -3198
rect 9976 -3220 9988 -3186
rect 10284 -3202 10470 -2808
rect 10566 -2946 10624 -2940
rect 10566 -2980 10578 -2946
rect 10566 -2986 10624 -2980
rect 10284 -3208 10528 -3202
rect 10662 -3208 10720 -3202
rect 9976 -3226 10034 -3220
rect 10284 -3242 10482 -3208
rect 10662 -3242 10674 -3208
rect 10284 -3248 10528 -3242
rect 10662 -3248 10720 -3242
rect 2912 -3280 2970 -3274
rect 2912 -3314 2924 -3280
rect 2912 -3320 2970 -3314
rect 1512 -3340 1570 -3334
rect 2194 -3340 2252 -3334
rect 1512 -3374 1524 -3340
rect 2194 -3374 2206 -3340
rect 10284 -3358 10470 -3248
rect 1512 -3380 1570 -3374
rect 2194 -3380 2252 -3374
rect 7258 -3482 7316 -3476
rect 7258 -3516 7270 -3482
rect 7258 -3522 7316 -3516
rect 10010 -3528 10068 -3522
rect 10010 -3562 10022 -3528
rect 10570 -3540 10628 -3534
rect 10010 -3568 10068 -3562
rect 10570 -3574 10582 -3540
rect 10570 -3580 10628 -3574
rect 10010 -3722 10068 -3716
rect 7258 -3760 7316 -3754
rect 10010 -3756 10022 -3722
rect 7258 -3794 7270 -3760
rect 10010 -3762 10068 -3756
rect 7258 -3800 7316 -3794
rect 10570 -3850 10628 -3844
rect 10570 -3884 10582 -3850
rect 10570 -3890 10628 -3884
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
use sky130_fd_pr__nfet_01v8_PWNS5P  XM1
timestamp 1696942209
transform 1 0 2223 0 1 -2902
box -211 -610 211 610
use sky130_fd_pr__nfet_01v8_lvt_F5PS5H  XM2
timestamp 1696942209
transform 1 0 3665 0 1 -2860
box -359 -410 359 410
use sky130_fd_pr__nfet_01v8_lvt_F5PS5H  XM3
timestamp 1696942209
transform 1 0 869 0 1 -2926
box -359 -410 359 410
use sky130_fd_pr__nfet_01v8_PWNS5P  XM4
timestamp 1696942209
transform 1 0 1541 0 1 -2902
box -211 -610 211 610
use sky130_fd_pr__nfet_01v8_PWNS5P  XM5
timestamp 1696942209
transform 1 0 2941 0 1 -2842
box -211 -610 211 610
use sky130_fd_pr__pfet_01v8_XGAKDL  XM6
timestamp 1696942209
transform 1 0 1657 0 1 -1203
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XGAKDL  XM7
timestamp 1696942209
transform 1 0 2509 0 1 -1185
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XGAKDL  XM8
timestamp 1696942209
transform 1 0 1183 0 1 -1219
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XGAKDL  XM9
timestamp 1696942209
transform 1 0 685 0 1 -1185
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XGAKDL  XM10
timestamp 1696942209
transform 1 0 3085 0 1 -1169
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XGAKDL  XM11
timestamp 1696942209
transform 1 0 3693 0 1 -1195
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_MQX2PY  XM12
timestamp 1696942209
transform 1 0 4789 0 1 -865
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_L7T3GD  XM13
timestamp 1696942209
transform 1 0 4771 0 1 -1432
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_HFBCFR  XM14
timestamp 1696942209
transform 1 0 5561 0 1 -780
box -311 -286 311 286
use sky130_fd_pr__nfet_01v8_648S5X  XM15
timestamp 1696942209
transform 1 0 5507 0 1 -1368
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_MQX2PY  XM16
timestamp 1696942209
transform 1 0 6435 0 1 -819
box -211 -303 211 303
use sky130_fd_pr__pfet_01v8_MQX2PY  XM17
timestamp 1696942209
transform 1 0 7007 0 1 -837
box -211 -303 211 303
use sky130_fd_pr__pfet_01v8_MQX2PY  XM18
timestamp 1696942209
transform 1 0 4733 0 1 -2313
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_9NW3WL  XM19
timestamp 1696942209
transform 1 0 7053 0 1 -1626
box -211 -294 211 294
use sky130_fd_pr__nfet_01v8_L7T3GD  XM20
timestamp 1696942209
transform 1 0 4733 0 1 -2968
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_HFBCFR  XM21
timestamp 1696942209
transform 1 0 5503 0 1 -2280
box -311 -286 311 286
use sky130_fd_pr__nfet_01v8_648S5X  XM22
timestamp 1696942209
transform 1 0 5503 0 1 -2994
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_9NW3WL  XM23
timestamp 1696942209
transform 1 0 6459 0 1 -1578
box -211 -294 211 294
use sky130_fd_pr__pfet_01v8_MQX2PY  XM24
timestamp 1696942209
transform 1 0 6841 0 1 -2247
box -211 -303 211 303
use sky130_fd_pr__pfet_01v8_MQX2PY  XM25
timestamp 1696942209
transform 1 0 7643 0 1 -2229
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_9NW3WL  XM26
timestamp 1696942209
transform 1 0 7291 0 1 -2968
box -211 -294 211 294
use sky130_fd_pr__nfet_01v8_9NW3WL  XM27
timestamp 1696942209
transform 1 0 7287 0 1 -3638
box -211 -294 211 294
use sky130_fd_pr__pfet_01v8_MQX2PY  XM28
timestamp 1696942209
transform 1 0 8513 0 1 -2345
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_L7T3GD  XM29
timestamp 1696942209
transform 1 0 8513 0 1 -3042
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_MQX2PY  XM30
timestamp 1696942209
transform 1 0 9935 0 1 -1411
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_L7T3GD  XM31
timestamp 1696942209
transform 1 0 9959 0 1 -1998
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_HFBCFR  XM32
timestamp 1696942209
transform 1 0 10629 0 1 -1358
box -311 -286 311 286
use sky130_fd_pr__nfet_01v8_648S5X  XM33
timestamp 1696942209
transform 1 0 10565 0 1 -1974
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_MQX2PY  XM34
timestamp 1696942209
transform 1 0 10005 0 1 -3055
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_L7T3GD  XM35
timestamp 1696942209
transform 1 0 10039 0 1 -3642
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_HFBCFR  XM36
timestamp 1696942209
transform 1 0 10595 0 1 -3094
box -311 -286 311 286
use sky130_fd_pr__nfet_01v8_648S5X  XM37
timestamp 1696942209
transform 1 0 10599 0 1 -3712
box -211 -310 211 310
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 cdac_vn
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 cdac_vp
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 VDD
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 clk
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 X
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 Y
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 P
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 Q
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 ready
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 X_drive
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 Y_drive
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 comp_outp
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 comp_outn
port 13 nsew
<< end >>
