* NGSPICE file created from hgu_comp_flat.ext - technology: sky130A

.subckt hgu_comp ready cdac_vn comp_outp comp_outn cdac_vp clk VDD VSS P Q a_1566_n378# a_1248_n288#
X0 ready.t0 a_564_n1721# VDD.t38 VDD.t37 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X1 a_564_n1721# a_476_n1721# a_564_n1266# VSS.t62 sky130_fd_pr__nfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X2 comp_outn.t2 a_1950_n1721# VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X3 Q cdac_vn.t0 a_582_n700# VSS.t65 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X4 a_1950_n1721# RS_n VDD.t10 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X5 a_482_n1818# a_1716_n1348# VSS.t37 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X6 P cdac_vp.t0 a_582_n700# VSS.t52 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X7 a_564_n1721# a_482_n1818# a_476_n1721# VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
X8 VDD.t36 a_1026_n1747# comp_outp.t2 VDD.t35 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X9 VSS.t56 RS_p a_1026_n1747# VSS.t55 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X10 VDD.t50 clk.t0 a_1248_n288# VDD.t49 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X11 a_582_n700# cdac_vp.t1 P VSS.t61 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X12 a_582_n700# cdac_vn.t1 Q VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X13 VDD.t24 a_852_n296# a_476_n1721# VDD.t23 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X14 ready.t1 a_564_n1721# VSS.t47 VSS.t46 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X15 comp_outp.t1 a_1026_n1747# VDD.t34 VDD.t33 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X16 a_476_n1721# a_852_n296# VDD.t22 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X17 comp_outn.t5 a_1950_n1721# VSS.t17 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X18 VDD.t48 RS_p a_1026_n1747# VDD.t47 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X19 VDD.t20 a_852_n296# a_476_n1721# VDD.t19 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X20 a_582_n700# cdac_vp.t2 P VSS.t59 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X21 a_582_n700# cdac_vn.t2 Q VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X22 a_564_n1266# a_482_n1818# VSS.t6 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
X23 VSS.t44 a_1026_n1747# comp_outp.t5 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X24 a_1950_n1721# RS_n VSS.t11 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X25 a_1566_n378# clk.t1 VDD.t12 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X26 VSS.t27 a_852_n296# a_476_n1721# VSS.t26 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X27 Q cdac_vn.t3 a_582_n700# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X28 VDD.t6 a_1248_n288# a_852_n296# VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X29 a_482_n1818# a_1716_n1348# VSS.t35 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X30 a_582_n700# clk.t2 VSS.t64 VSS.t63 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X31 comp_outp.t4 a_1026_n1747# VSS.t42 VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X32 VSS.t9 a_1248_n288# a_852_n296# VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X33 P cdac_vp.t3 a_582_n700# VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X34 a_1248_n288# a_1566_n378# VDD.t44 VDD.t43 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X35 Q clk.t3 VDD.t2 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X36 VDD.t32 a_1026_n1747# comp_outp.t0 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X37 RS_n a_1716_n1348# VSS.t33 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X38 comp_outn.t1 a_1950_n1721# VDD.t16 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X39 a_582_n700# cdac_vp.t4 P VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X40 a_582_n700# cdac_vn.t4 Q VSS.t57 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X41 a_1716_n1348# a_1566_n378# VSS.t51 VSS.t50 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X42 VSS.t31 a_1716_n1348# a_482_n1818# VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X43 VSS.t3 clk.t4 a_582_n700# VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X44 VSS.t25 a_852_n296# a_476_n1721# VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X45 Q a_1566_n378# a_1248_n288# VSS.t49 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X46 P cdac_vp.t5 a_582_n700# VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X47 RS_n RS_p VDD.t46 VDD.t45 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X48 VDD.t14 a_1950_n1721# comp_outn.t0 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X49 a_1716_n1348# a_1566_n378# VDD.t42 VDD.t41 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X50 a_582_n700# clk.t5 VSS.t19 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X51 a_582_n700# cdac_vn.t5 Q VSS.t58 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X52 VDD.t40 clk.t6 P VDD.t39 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X53 VSS.t40 a_1026_n1747# comp_outp.t3 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X54 Q cdac_vn.t6 a_582_n700# VSS.t60 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X55 comp_outn.t4 a_1950_n1721# VSS.t15 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
X56 a_482_n1818# a_1716_n1348# VDD.t30 VDD.t29 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X57 a_482_n1818# a_1716_n1348# VDD.t28 VDD.t27 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
X58 P cdac_vp.t6 a_582_n700# VSS.t54 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X59 VSS.t23 a_852_n296# RS_p VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
X60 VDD.t26 a_1716_n1348# a_482_n1818# VDD.t25 sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X61 a_482_n1818# a_476_n1721# a_564_n1721# VDD.t51 sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.122 ps=1.13 w=0.84 l=0.15
X62 a_582_n700# cdac_vp.t7 P VSS.t53 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X63 VSS.t13 a_1950_n1721# comp_outn.t3 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X64 a_476_n1721# a_852_n296# VSS.t21 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X65 VDD.t4 a_1248_n288# a_1566_n378# VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X66 a_1566_n378# a_1248_n288# P VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X67 VSS.t48 clk.t7 a_582_n700# VSS.t32 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X68 Q cdac_vn.t7 a_582_n700# VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X69 VDD.t8 RS_n RS_p VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.13 as=0.244 ps=2.26 w=0.84 l=0.15
R0 VDD.n242 VDD.t51 425.812
R1 VDD.t51 VDD.t0 183.923
R2 VDD.n171 VDD.t29 112.871
R3 VDD.n17 VDD.t19 112.871
R4 VDD.n334 VDD.t15 112.871
R5 VDD.n230 VDD.t35 103.466
R6 VDD.n281 VDD.t7 97.2098
R7 VDD.n99 VDD.t49 89.3422
R8 VDD.n201 VDD.t31 84.654
R9 VDD.n33 VDD.t23 84.1029
R10 VDD.n363 VDD.t17 84.1029
R11 VDD.n85 VDD.t11 71.4739
R12 VDD.n187 VDD.t27 65.291
R13 VDD.n85 VDD.t3 59.5616
R14 VDD.n135 VDD.t41 53.6055
R15 VDD.n298 VDD.t45 53.5216
R16 VDD.n99 VDD.t43 41.6933
R17 VDD.n23 VDD.t20 39.1333
R18 VDD.n152 VDD.t30 39.1333
R19 VDD.n332 VDD.t16 39.1333
R20 VDD.n206 VDD.t32 39.1333
R21 VDD.n315 VDD.t9 39.1171
R22 VDD.n14 VDD.t22 38.6969
R23 VDD.n14 VDD.t24 38.6969
R24 VDD.n184 VDD.t28 38.6969
R25 VDD.n184 VDD.t26 38.6969
R26 VDD.n366 VDD.t18 38.6969
R27 VDD.n366 VDD.t14 38.6969
R28 VDD.n227 VDD.t34 38.6969
R29 VDD.n227 VDD.t36 38.6969
R30 VDD.n171 VDD.t25 37.6243
R31 VDD.n51 VDD.t5 35.7372
R32 VDD.n246 VDD.t38 34.4966
R33 VDD.n264 VDD.t48 34.4575
R34 VDD.n50 VDD.t6 34.4428
R35 VDD.n140 VDD.t42 34.4428
R36 VDD.n320 VDD.t10 34.4428
R37 VDD.n302 VDD.t46 34.0065
R38 VDD.n302 VDD.t8 34.0065
R39 VDD.n67 VDD.t39 29.7811
R40 VDD.n82 VDD.t12 28.5655
R41 VDD.n82 VDD.t40 28.5655
R42 VDD.n103 VDD.t44 28.5655
R43 VDD.n103 VDD.t4 28.5655
R44 VDD.n118 VDD.t2 28.5655
R45 VDD.n118 VDD.t50 28.5655
R46 VDD.n26 VDD.t21 18.8124
R47 VDD.n350 VDD.t13 18.8124
R48 VDD.n121 VDD.t1 11.9127
R49 VDD.n268 VDD.n267 10.6304
R50 VDD.n243 VDD.n242 9.92059
R51 VDD.n215 VDD.t33 9.40644
R52 VDD.n28 VDD.n27 8.85536
R53 VDD.n27 VDD.n26 8.85536
R54 VDD.n19 VDD.n18 8.85536
R55 VDD.n18 VDD.n17 8.85536
R56 VDD.n53 VDD.n52 8.85536
R57 VDD.n52 VDD.n51 8.85536
R58 VDD.n69 VDD.n68 8.85536
R59 VDD.n68 VDD.n67 8.85536
R60 VDD.n87 VDD.n86 8.85536
R61 VDD.n86 VDD.n85 8.85536
R62 VDD.n101 VDD.n100 8.85536
R63 VDD.n100 VDD.n99 8.85536
R64 VDD.n123 VDD.n122 8.85536
R65 VDD.n122 VDD.n121 8.85536
R66 VDD.n137 VDD.n136 8.85536
R67 VDD.n136 VDD.n135 8.85536
R68 VDD.n188 VDD.n187 8.85536
R69 VDD.n173 VDD.n172 8.85536
R70 VDD.n172 VDD.n171 8.85536
R71 VDD.n157 VDD.n156 8.85536
R72 VDD.n156 VDD.n155 8.85536
R73 VDD.n34 VDD.n33 8.85536
R74 VDD.n336 VDD.n335 8.85536
R75 VDD.n335 VDD.n334 8.85536
R76 VDD.n217 VDD.n216 8.85536
R77 VDD.n216 VDD.n215 8.85536
R78 VDD.n203 VDD.n202 8.85536
R79 VDD.n202 VDD.n201 8.85536
R80 VDD.n269 VDD.n268 8.85536
R81 VDD.n283 VDD.n282 8.85536
R82 VDD.n282 VDD.n281 8.85536
R83 VDD.n300 VDD.n299 8.85536
R84 VDD.n299 VDD.n298 8.85536
R85 VDD.n317 VDD.n316 8.85536
R86 VDD.n316 VDD.n315 8.85536
R87 VDD.n232 VDD.n231 8.85536
R88 VDD.n231 VDD.n230 8.85536
R89 VDD.n244 VDD.n243 8.85536
R90 VDD.n364 VDD.n363 8.85536
R91 VDD.n352 VDD.n351 8.85536
R92 VDD.n351 VDD.n350 8.85536
R93 VDD.n267 VDD.t47 5.50293
R94 VDD.n35 VDD.n34 3.03483
R95 VDD.n29 VDD.n28 3.03311
R96 VDD.n88 VDD.n87 3.03311
R97 VDD.n102 VDD.n101 3.03311
R98 VDD.n124 VDD.n123 3.03311
R99 VDD.n138 VDD.n137 3.03311
R100 VDD.n174 VDD.n173 3.03311
R101 VDD.n189 VDD.n188 3.03311
R102 VDD.n20 VDD.n19 3.03311
R103 VDD.n54 VDD.n53 3.03311
R104 VDD.n70 VDD.n69 3.03311
R105 VDD.n158 VDD.n157 3.03311
R106 VDD.n218 VDD.n217 3.03311
R107 VDD.n365 VDD.n364 3.03311
R108 VDD.n245 VDD.n244 3.03311
R109 VDD.n204 VDD.n203 3.03311
R110 VDD.n270 VDD.n269 3.03311
R111 VDD.n284 VDD.n283 3.03311
R112 VDD.n301 VDD.n300 3.03311
R113 VDD.n318 VDD.n317 3.03311
R114 VDD.n337 VDD.n336 3.03311
R115 VDD.n233 VDD.n232 3.03311
R116 VDD.n353 VDD.n352 3.03311
R117 VDD.n242 VDD.t37 1.83498
R118 VDD.n58 VDD.n57 1.7055
R119 VDD.n74 VDD.n73 1.7055
R120 VDD.n162 VDD.n161 1.7055
R121 VDD.n193 VDD.n192 1.7055
R122 VDD.n178 VDD.n177 1.7055
R123 VDD.n145 VDD.n144 1.7055
R124 VDD.n128 VDD.n127 1.7055
R125 VDD.n110 VDD.n109 1.7055
R126 VDD.n92 VDD.n91 1.7055
R127 VDD.n358 VDD.n357 1.7055
R128 VDD.n342 VDD.n341 1.7055
R129 VDD.n325 VDD.n324 1.7055
R130 VDD.n308 VDD.n307 1.7055
R131 VDD.n290 VDD.n289 1.7055
R132 VDD.n274 VDD.n273 1.7055
R133 VDD.n372 VDD.n371 1.7055
R134 VDD.n56 VDD.n55 1.35607
R135 VDD.n72 VDD.n71 1.35607
R136 VDD.n160 VDD.n159 1.35607
R137 VDD.n191 VDD.n190 1.35607
R138 VDD.n176 VDD.n175 1.35607
R139 VDD.n142 VDD.n141 1.35607
R140 VDD.n126 VDD.n125 1.35607
R141 VDD.n107 VDD.n106 1.35607
R142 VDD.n90 VDD.n89 1.35607
R143 VDD.n37 VDD.n36 1.14764
R144 VDD.n248 VDD.n247 1.04225
R145 VDD.n370 VDD.n369 1.04225
R146 VDD.n236 VDD.n235 1.04225
R147 VDD.n221 VDD.n220 1.04225
R148 VDD.n208 VDD.n207 1.04225
R149 VDD.n272 VDD.n271 1.04225
R150 VDD.n287 VDD.n286 1.04225
R151 VDD.n306 VDD.n305 1.04225
R152 VDD.n322 VDD.n321 1.04225
R153 VDD.n340 VDD.n339 1.04225
R154 VDD.n356 VDD.n355 1.04225
R155 VDD.n250 VDD.n249 0.861312
R156 VDD.n36 VDD.n35 0.850734
R157 VDD.n374 VDD.n194 0.731708
R158 VDD.n83 VDD.n82 0.479026
R159 VDD.n104 VDD.n103 0.479026
R160 VDD.n119 VDD.n118 0.479026
R161 VDD.n31 VDD.n14 0.436881
R162 VDD.n185 VDD.n184 0.436881
R163 VDD.n367 VDD.n366 0.436881
R164 VDD.n303 VDD.n302 0.436881
R165 VDD.n228 VDD.n227 0.436881
R166 VDD.n374 VDD.n373 0.43282
R167 VDD.n16 VDD.n15 0.225109
R168 VDD.n24 VDD.n23 0.213391
R169 VDD.n229 VDD.n228 0.182141
R170 VDD.n32 VDD.n31 0.145031
R171 VDD.n368 VDD.n367 0.141125
R172 VDD.n84 VDD.n83 0.139172
R173 VDD.n186 VDD.n185 0.123547
R174 VDD.n196 VDD.n195 0.117957
R175 VDD.n210 VDD.n209 0.115802
R176 VDD.n223 VDD.n222 0.115802
R177 VDD.n12 VDD.n11 0.113847
R178 VDD.n6 VDD.n5 0.10961
R179 VDD.n238 VDD.n237 0.0996379
R180 VDD.n105 VDD.n104 0.0981562
R181 VDD.n304 VDD.n303 0.0883906
R182 VDD.n31 VDD.n30 0.078625
R183 VDD.n120 VDD.n119 0.0610469
R184 VDD.n260 VDD.n259 0.0539828
R185 VDD.n344 VDD.n343 0.0531724
R186 VDD.n310 VDD.n309 0.0531724
R187 VDD.n147 VDD.n146 0.0530763
R188 VDD.n44 VDD.n43 0.0530763
R189 VDD.n257 VDD.n256 0.0523621
R190 VDD.n254 VDD.n253 0.0523621
R191 VDD.n112 VDD.n111 0.0522797
R192 VDD.n38 VDD.n37 0.0522797
R193 VDD.n360 VDD.n359 0.0515517
R194 VDD.n292 VDD.n291 0.0515517
R195 VDD.n180 VDD.n179 0.0514831
R196 VDD.n76 VDD.n75 0.0514831
R197 VDD.n327 VDD.n326 0.0507414
R198 VDD.n276 VDD.n275 0.0507414
R199 VDD.n164 VDD.n163 0.0506864
R200 VDD.n130 VDD.n129 0.0506864
R201 VDD.n94 VDD.n93 0.0506864
R202 VDD.n60 VDD.n59 0.0506864
R203 VDD.n41 VDD.n40 0.0498898
R204 VDD.n251 VDD.n250 0.0462845
R205 VDD.n35 VDD.n32 0.0427461
R206 VDD.n189 VDD.n186 0.0415156
R207 VDD.n175 VDD.n169 0.0415156
R208 VDD.n174 VDD.n170 0.0415156
R209 VDD.n138 VDD.n134 0.0415156
R210 VDD.n125 VDD.n117 0.0415156
R211 VDD.n124 VDD.n120 0.0415156
R212 VDD.n102 VDD.n98 0.0415156
R213 VDD.n106 VDD.n105 0.0415156
R214 VDD.n89 VDD.n81 0.0415156
R215 VDD.n88 VDD.n84 0.0415156
R216 VDD.n71 VDD.n65 0.0415156
R217 VDD.n70 VDD.n66 0.0415156
R218 VDD.n20 VDD.n16 0.0415156
R219 VDD.n22 VDD.n21 0.0415156
R220 VDD.n318 VDD.n314 0.0415156
R221 VDD.n284 VDD.n280 0.0415156
R222 VDD.n286 VDD.n285 0.0415156
R223 VDD.n204 VDD.n200 0.0415156
R224 VDD.n218 VDD.n214 0.0415156
R225 VDD.n220 VDD.n219 0.0415156
R226 VDD.n233 VDD.n229 0.0415156
R227 VDD.n235 VDD.n234 0.0415156
R228 VDD.n245 VDD.n241 0.0415156
R229 VDD.n247 VDD.n246 0.0415156
R230 VDD.n159 VDD.n153 0.0395625
R231 VDD.n158 VDD.n154 0.0395625
R232 VDD.n25 VDD.n24 0.0395625
R233 VDD.n30 VDD.n29 0.0395625
R234 VDD.n353 VDD.n349 0.0395625
R235 VDD.n355 VDD.n354 0.0395625
R236 VDD.n301 VDD.n297 0.0395625
R237 VDD.n305 VDD.n304 0.0395625
R238 VDD.n271 VDD.n265 0.0395625
R239 VDD.n270 VDD.n266 0.0395625
R240 VDD.n369 VDD.n368 0.0376094
R241 VDD.n337 VDD.n333 0.0376094
R242 VDD.n339 VDD.n338 0.0376094
R243 VDD.n321 VDD.n320 0.0376094
R244 VDD.n55 VDD.n50 0.0337031
R245 VDD.n206 VDD.n205 0.03175
R246 VDD.n265 VDD.n264 0.0297969
R247 VDD.n140 VDD.n139 0.0278438
R248 VDD.n153 VDD.n152 0.0258906
R249 VDD.n322 VDD.n313 0.0231293
R250 VDD.n287 VDD.n279 0.0231293
R251 VDD.n209 VDD.n208 0.0231293
R252 VDD.n222 VDD.n221 0.0231293
R253 VDD.n237 VDD.n236 0.0231293
R254 VDD.n240 VDD.n239 0.0231293
R255 VDD.n183 VDD.n182 0.0227458
R256 VDD.n168 VDD.n167 0.0227458
R257 VDD.n142 VDD.n133 0.0227458
R258 VDD.n116 VDD.n115 0.0227458
R259 VDD.n107 VDD.n97 0.0227458
R260 VDD.n80 VDD.n79 0.0227458
R261 VDD.n64 VDD.n63 0.0227458
R262 VDD.n5 VDD.n4 0.0227458
R263 VDD.n347 VDD.n346 0.0220517
R264 VDD.n356 VDD.n348 0.0220517
R265 VDD.n324 VDD.n312 0.0220517
R266 VDD.n295 VDD.n294 0.0220517
R267 VDD.n306 VDD.n296 0.0220517
R268 VDD.n289 VDD.n278 0.0220517
R269 VDD.n198 VDD.n197 0.0220517
R270 VDD.n212 VDD.n211 0.0220517
R271 VDD.n225 VDD.n224 0.0220517
R272 VDD.n36 VDD.n13 0.0218329
R273 VDD.n151 VDD.n150 0.0216864
R274 VDD.n144 VDD.n132 0.0216864
R275 VDD.n109 VDD.n96 0.0216864
R276 VDD.n48 VDD.n47 0.0216864
R277 VDD.n2 VDD.n1 0.0216864
R278 VDD.n11 VDD.n10 0.0216864
R279 VDD.n370 VDD.n362 0.0209741
R280 VDD.n330 VDD.n329 0.0209741
R281 VDD.n340 VDD.n331 0.0209741
R282 VDD.n192 VDD.n181 0.0206271
R283 VDD.n177 VDD.n166 0.0206271
R284 VDD.n127 VDD.n114 0.0206271
R285 VDD.n91 VDD.n78 0.0206271
R286 VDD.n73 VDD.n62 0.0206271
R287 VDD.n273 VDD.n262 0.0198966
R288 VDD.n161 VDD.n149 0.0195678
R289 VDD.n57 VDD.n46 0.0195678
R290 VDD.n8 VDD.n7 0.0195678
R291 VDD VDD.n374 0.0161119
R292 VDD.n371 VDD.n361 0.0144047
R293 VDD.n141 VDD.n140 0.0141719
R294 VDD.n373 VDD.n372 0.0110345
R295 VDD.n359 VDD.n358 0.0110345
R296 VDD.n343 VDD.n342 0.0110345
R297 VDD.n326 VDD.n325 0.0110345
R298 VDD.n309 VDD.n308 0.0110345
R299 VDD.n291 VDD.n290 0.0110345
R300 VDD.n275 VDD.n274 0.0110345
R301 VDD.n259 VDD.n258 0.0110345
R302 VDD.n256 VDD.n255 0.0110345
R303 VDD.n253 VDD.n252 0.0110345
R304 VDD.n194 VDD.n193 0.0108559
R305 VDD.n179 VDD.n178 0.0108559
R306 VDD.n163 VDD.n162 0.0108559
R307 VDD.n146 VDD.n145 0.0108559
R308 VDD.n129 VDD.n128 0.0108559
R309 VDD.n111 VDD.n110 0.0108559
R310 VDD.n93 VDD.n92 0.0108559
R311 VDD.n75 VDD.n74 0.0108559
R312 VDD.n59 VDD.n58 0.0108559
R313 VDD.n43 VDD.n42 0.0108559
R314 VDD.n40 VDD.n39 0.0108559
R315 VDD.n369 VDD.n365 0.0102656
R316 VDD.n333 VDD.n332 0.0102656
R317 VDD.n339 VDD.n337 0.0102656
R318 VDD.n207 VDD.n206 0.0102656
R319 VDD.n262 VDD.n261 0.00912069
R320 VDD.n149 VDD.n148 0.00897458
R321 VDD.n46 VDD.n45 0.00897458
R322 VDD.n7 VDD.n6 0.00897458
R323 VDD.n166 VDD.n165 0.00791525
R324 VDD.n114 VDD.n113 0.00791525
R325 VDD.n78 VDD.n77 0.00791525
R326 VDD.n62 VDD.n61 0.00791525
R327 VDD.n13 VDD.n12 0.00791525
R328 VDD.n312 VDD.n311 0.00696552
R329 VDD.n278 VDD.n277 0.00696552
R330 VDD.n197 VDD.n196 0.00696552
R331 VDD.n211 VDD.n210 0.00696552
R332 VDD.n224 VDD.n223 0.00696552
R333 VDD.n132 VDD.n131 0.00685593
R334 VDD.n96 VDD.n95 0.00685593
R335 VDD.n1 VDD.n0 0.00685593
R336 VDD.n249 VDD.n248 0.00660795
R337 VDD.n159 VDD.n158 0.00635938
R338 VDD.n50 VDD.n49 0.00635938
R339 VDD.n55 VDD.n54 0.00635938
R340 VDD.n29 VDD.n25 0.00635938
R341 VDD.n355 VDD.n353 0.00635938
R342 VDD.n305 VDD.n301 0.00635938
R343 VDD.n271 VDD.n270 0.00635938
R344 VDD.n346 VDD.n345 0.00588793
R345 VDD.n294 VDD.n293 0.00588793
R346 VDD.n239 VDD.n238 0.00588793
R347 VDD.n329 VDD.n328 0.00481034
R348 VDD.n23 VDD.n22 0.00440625
R349 VDD.n320 VDD.n319 0.00440625
R350 VDD.n341 VDD.n330 0.00373276
R351 VDD.n272 VDD.n263 0.00373276
R352 VDD.n160 VDD.n151 0.00367797
R353 VDD.n56 VDD.n48 0.00367797
R354 VDD.n10 VDD.n9 0.00367797
R355 VDD.n371 VDD.n370 0.00265517
R356 VDD.n357 VDD.n356 0.00265517
R357 VDD.n341 VDD.n340 0.00265517
R358 VDD.n307 VDD.n306 0.00265517
R359 VDD.n273 VDD.n272 0.00265517
R360 VDD.n192 VDD.n191 0.00261864
R361 VDD.n177 VDD.n176 0.00261864
R362 VDD.n161 VDD.n160 0.00261864
R363 VDD.n127 VDD.n126 0.00261864
R364 VDD.n91 VDD.n90 0.00261864
R365 VDD.n73 VDD.n72 0.00261864
R366 VDD.n57 VDD.n56 0.00261864
R367 VDD.n9 VDD.n8 0.00261864
R368 VDD.n190 VDD.n189 0.00245312
R369 VDD.n175 VDD.n174 0.00245312
R370 VDD.n141 VDD.n138 0.00245312
R371 VDD.n125 VDD.n124 0.00245312
R372 VDD.n106 VDD.n102 0.00245312
R373 VDD.n89 VDD.n88 0.00245312
R374 VDD.n71 VDD.n70 0.00245312
R375 VDD.n21 VDD.n20 0.00245312
R376 VDD.n321 VDD.n318 0.00245312
R377 VDD.n286 VDD.n284 0.00245312
R378 VDD.n207 VDD.n204 0.00245312
R379 VDD.n220 VDD.n218 0.00245312
R380 VDD.n235 VDD.n233 0.00245312
R381 VDD.n247 VDD.n245 0.00245312
R382 VDD.n357 VDD.n347 0.00157759
R383 VDD.n324 VDD.n323 0.00157759
R384 VDD.n323 VDD.n322 0.00157759
R385 VDD.n307 VDD.n295 0.00157759
R386 VDD.n289 VDD.n288 0.00157759
R387 VDD.n288 VDD.n287 0.00157759
R388 VDD.n199 VDD.n198 0.00157759
R389 VDD.n208 VDD.n199 0.00157759
R390 VDD.n213 VDD.n212 0.00157759
R391 VDD.n221 VDD.n213 0.00157759
R392 VDD.n226 VDD.n225 0.00157759
R393 VDD.n236 VDD.n226 0.00157759
R394 VDD.n248 VDD.n240 0.00157759
R395 VDD.n191 VDD.n183 0.00155932
R396 VDD.n176 VDD.n168 0.00155932
R397 VDD.n144 VDD.n143 0.00155932
R398 VDD.n143 VDD.n142 0.00155932
R399 VDD.n126 VDD.n116 0.00155932
R400 VDD.n109 VDD.n108 0.00155932
R401 VDD.n108 VDD.n107 0.00155932
R402 VDD.n90 VDD.n80 0.00155932
R403 VDD.n72 VDD.n64 0.00155932
R404 VDD.n3 VDD.n2 0.00155932
R405 VDD.n4 VDD.n3 0.00155932
R406 VDD.n372 VDD.n360 0.00131035
R407 VDD.n358 VDD.n344 0.00131035
R408 VDD.n342 VDD.n327 0.00131035
R409 VDD.n325 VDD.n310 0.00131035
R410 VDD.n308 VDD.n292 0.00131035
R411 VDD.n290 VDD.n276 0.00131035
R412 VDD.n274 VDD.n260 0.00131035
R413 VDD.n258 VDD.n257 0.00131035
R414 VDD.n255 VDD.n254 0.00131035
R415 VDD.n252 VDD.n251 0.00131035
R416 VDD.n193 VDD.n180 0.00129661
R417 VDD.n178 VDD.n164 0.00129661
R418 VDD.n162 VDD.n147 0.00129661
R419 VDD.n145 VDD.n130 0.00129661
R420 VDD.n128 VDD.n112 0.00129661
R421 VDD.n110 VDD.n94 0.00129661
R422 VDD.n92 VDD.n76 0.00129661
R423 VDD.n74 VDD.n60 0.00129661
R424 VDD.n58 VDD.n44 0.00129661
R425 VDD.n42 VDD.n41 0.00129661
R426 VDD.n39 VDD.n38 0.00129661
R427 ready.n0 ready.t1 42.3194
R428 ready.n0 ready.t0 34.4226
R429 ready ready.n0 14.5094
R430 VSS.n109 VSS.t60 179.739
R431 VSS.n104 VSS.t10 179.739
R432 VSS.n121 VSS.t12 175.16
R433 VSS.n81 VSS.t55 172.549
R434 VSS.n67 VSS.t39 172.549
R435 VSS.n72 VSS.t61 165.359
R436 VSS.n67 VSS.t53 165.359
R437 VSS.n91 VSS.t32 165.359
R438 VSS.n115 VSS.t14 161.147
R439 VSS.n91 VSS.t22 150.981
R440 VSS.n114 VSS.t65 140.127
R441 VSS.n34 VSS.t5 129.412
R442 VSS.n87 VSS.t7 122.222
R443 VSS.n98 VSS.t49 107.844
R444 VSS.n42 VSS.t59 107.844
R445 VSS.t8 VSS.t29 100.654
R446 VSS.n62 VSS.t24 93.4646
R447 VSS.n38 VSS.t45 93.4646
R448 VSS.n162 VSS.t1 91.0833
R449 VSS.n33 VSS.t6 83.725
R450 VSS.n72 VSS.t8 79.0855
R451 VSS.n58 VSS.t20 79.0855
R452 VSS.t45 VSS.t62 79.0855
R453 VSS.t50 VSS.t38 79.0708
R454 VSS.n97 VSS.n96 79.0622
R455 VSS.n86 VSS.n85 79.0622
R456 VSS.n166 VSS.t58 77.0706
R457 VSS.n120 VSS.t36 70.0642
R458 VSS.n53 VSS.t26 64.7064
R459 VSS.n108 VSS.t50 57.5168
R460 VSS.t24 VSS.t52 57.5168
R461 VSS.t20 VSS.t4 57.5168
R462 VSS.t26 VSS.t54 57.5168
R463 VSS.t34 VSS.t28 56.0515
R464 VSS.t30 VSS.t0 56.0515
R465 VSS.n125 VSS.t30 56.0515
R466 VSS.t36 VSS.t57 56.0515
R467 VSS.t54 VSS.t46 50.3273
R468 VSS.n19 VSS.t25 43.3862
R469 VSS.n147 VSS.t37 43.3862
R470 VSS.n71 VSS.t40 43.3862
R471 VSS.n113 VSS.t15 43.3862
R472 VSS.t49 VSS.t18 43.1378
R473 VSS.t7 VSS.t2 43.1378
R474 VSS.n12 VSS.t21 43.044
R475 VSS.n12 VSS.t27 43.044
R476 VSS.n138 VSS.t35 43.044
R477 VSS.n138 VSS.t31 43.044
R478 VSS.n8 VSS.t42 43.044
R479 VSS.n8 VSS.t44 43.044
R480 VSS.n3 VSS.t17 43.044
R481 VSS.n3 VSS.t13 43.044
R482 VSS.n131 VSS.t34 42.0387
R483 VSS.n143 VSS.t51 41.8559
R484 VSS.n15 VSS.t9 41.843
R485 VSS.n80 VSS.t56 41.7956
R486 VSS.n103 VSS.t11 41.7956
R487 VSS.n51 VSS.t47 41.7882
R488 VSS.t22 VSS.t63 28.7587
R489 VSS.n47 VSS.n46 28.7587
R490 VSS.t57 VSS.t16 28.026
R491 VSS.n7 VSS.t33 20.7148
R492 VSS.n7 VSS.t23 20.7148
R493 VSS.n96 VSS.t19 19.8005
R494 VSS.n96 VSS.t48 19.8005
R495 VSS.n85 VSS.t64 19.8005
R496 VSS.n85 VSS.t3 19.8005
R497 VSS.n140 VSS.n139 9.15497
R498 VSS.n145 VSS.n144 9.15497
R499 VSS.n137 VSS.n136 9.15497
R500 VSS.n150 VSS.n149 9.15497
R501 VSS.n14 VSS.n13 9.15497
R502 VSS.n17 VSS.n16 9.15497
R503 VSS.n21 VSS.n20 9.15497
R504 VSS.n24 VSS.n23 9.15497
R505 VSS.n10 VSS.n9 9.15497
R506 VSS.n142 VSS.n141 9.15497
R507 VSS.n33 VSS.n32 9.15497
R508 VSS.n49 VSS.n48 9.15497
R509 VSS.n48 VSS.n47 9.15497
R510 VSS.n44 VSS.n43 9.15497
R511 VSS.n43 VSS.n42 9.15497
R512 VSS.n109 VSS.n108 7.19004
R513 VSS.t53 VSS.t41 7.19004
R514 VSS.t52 VSS.t43 7.19004
R515 VSS.n132 VSS.n131 7.00687
R516 VSS.n126 VSS.n125 7.00687
R517 VSS.n121 VSS.n120 7.00687
R518 VSS.n115 VSS.n114 7.00687
R519 VSS.n25 VSS.n24 4.6505
R520 VSS.n15 VSS.n14 4.6505
R521 VSS.n148 VSS.n140 4.6505
R522 VSS.n146 VSS.n145 4.6505
R523 VSS.n151 VSS.n150 4.6505
R524 VSS.n18 VSS.n17 4.6505
R525 VSS.n22 VSS.n21 4.6505
R526 VSS.n143 VSS.n142 4.6505
R527 VSS.n50 VSS.n49 4.6505
R528 VSS.n45 VSS.n44 4.6505
R529 VSS.n6 VSS.n5 4.57773
R530 VSS.n5 VSS.n4 4.57773
R531 VSS.n36 VSS.n35 4.57773
R532 VSS.n35 VSS.n34 4.57773
R533 VSS.n40 VSS.n39 4.57773
R534 VSS.n39 VSS.n38 4.57773
R535 VSS.n83 VSS.n82 4.57773
R536 VSS.n82 VSS.n81 4.57773
R537 VSS.n78 VSS.n77 4.57773
R538 VSS.n77 VSS.n76 4.57773
R539 VSS.n74 VSS.n73 4.57773
R540 VSS.n73 VSS.n72 4.57773
R541 VSS.n69 VSS.n68 4.57773
R542 VSS.n68 VSS.n67 4.57773
R543 VSS.n64 VSS.n63 4.57773
R544 VSS.n63 VSS.n62 4.57773
R545 VSS.n60 VSS.n59 4.57773
R546 VSS.n59 VSS.n58 4.57773
R547 VSS.n55 VSS.n54 4.57773
R548 VSS.n54 VSS.n53 4.57773
R549 VSS.n100 VSS.n99 4.57773
R550 VSS.n99 VSS.n98 4.57773
R551 VSS.n93 VSS.n92 4.57773
R552 VSS.n92 VSS.n91 4.57773
R553 VSS.n89 VSS.n88 4.57773
R554 VSS.n88 VSS.n87 4.57773
R555 VSS.n2 VSS.n1 4.57773
R556 VSS.n1 VSS.n0 4.57773
R557 VSS.n168 VSS.n167 4.57773
R558 VSS.n167 VSS.n166 4.57773
R559 VSS.n164 VSS.n163 4.57773
R560 VSS.n163 VSS.n162 4.57773
R561 VSS.n134 VSS.n133 4.57773
R562 VSS.n133 VSS.n132 4.57773
R563 VSS.n128 VSS.n127 4.57773
R564 VSS.n127 VSS.n126 4.57773
R565 VSS.n123 VSS.n122 4.57773
R566 VSS.n122 VSS.n121 4.57773
R567 VSS.n117 VSS.n116 4.57773
R568 VSS.n116 VSS.n115 4.57773
R569 VSS.n111 VSS.n110 4.57773
R570 VSS.n110 VSS.n109 4.57773
R571 VSS.n106 VSS.n105 4.57773
R572 VSS.n105 VSS.n104 4.57773
R573 VSS.n155 VSS.n137 3.03433
R574 VSS.n11 VSS.n10 3.03311
R575 VSS.n170 VSS.n2 2.34742
R576 VSS.n41 VSS.n40 2.3255
R577 VSS.n84 VSS.n83 2.3255
R578 VSS.n79 VSS.n78 2.3255
R579 VSS.n75 VSS.n74 2.3255
R580 VSS.n70 VSS.n69 2.3255
R581 VSS.n65 VSS.n64 2.3255
R582 VSS.n61 VSS.n60 2.3255
R583 VSS.n101 VSS.n100 2.3255
R584 VSS.n94 VSS.n93 2.3255
R585 VSS.n90 VSS.n89 2.3255
R586 VSS.n102 VSS.n6 2.3255
R587 VSS.n169 VSS.n168 2.3255
R588 VSS.n165 VSS.n164 2.3255
R589 VSS.n129 VSS.n128 2.3255
R590 VSS.n124 VSS.n123 2.3255
R591 VSS.n118 VSS.n117 2.3255
R592 VSS.n112 VSS.n111 2.3255
R593 VSS.n107 VSS.n106 2.3255
R594 VSS.n160 VSS.n159 2.2505
R595 VSS.n30 VSS.n28 2.24128
R596 VSS.n31 VSS.n30 1.93674
R597 VSS.n158 VSS.n157 1.93674
R598 VSS.n56 VSS.n55 1.83603
R599 VSS.n135 VSS.n134 1.83603
R600 VSS.n156 VSS.n155 1.51031
R601 VSS.n41 VSS.n37 1.22368
R602 VSS.n37 VSS.n33 1.18692
R603 VSS.n57 VSS.n31 1.16137
R604 VSS.n37 VSS.n36 0.585126
R605 VSS.n95 VSS.n7 0.433079
R606 VSS.n26 VSS.n12 0.342742
R607 VSS.n152 VSS.n138 0.342742
R608 VSS.n66 VSS.n8 0.342742
R609 VSS.n119 VSS.n3 0.342742
R610 VSS.n100 VSS.n97 0.340323
R611 VSS VSS.n170 0.231462
R612 VSS.n18 VSS.n15 0.216017
R613 VSS.n25 VSS.n22 0.216017
R614 VSS.n151 VSS.n148 0.216017
R615 VSS.n146 VSS.n143 0.216017
R616 VSS.n19 VSS.n18 0.168603
R617 VSS.n147 VSS.n146 0.155672
R618 VSS.n26 VSS.n25 0.151362
R619 VSS.n152 VSS.n151 0.138431
R620 VSS.n89 VSS.n86 0.113774
R621 VSS.n148 VSS.n147 0.0608448
R622 VSS.n94 VSS.n90 0.0558097
R623 VSS.n101 VSS.n95 0.0547035
R624 VSS.n45 VSS.n41 0.0535047
R625 VSS.n102 VSS.n101 0.0521284
R626 VSS.n90 VSS.n84 0.0512449
R627 VSS.n22 VSS.n19 0.0479138
R628 VSS.n154 VSS.n153 0.0457586
R629 VSS.n79 VSS.n75 0.0410844
R630 VSS.n65 VSS.n61 0.0410844
R631 VSS.n169 VSS.n165 0.0410844
R632 VSS.n129 VSS.n124 0.0410844
R633 VSS.n112 VSS.n107 0.0410844
R634 VSS.n27 VSS.n26 0.0406606
R635 VSS.n61 VSS.n57 0.0405313
R636 VSS.n119 VSS.n118 0.0402727
R637 VSS.n80 VSS.n79 0.039461
R638 VSS.n71 VSS.n70 0.039461
R639 VSS.n70 VSS.n66 0.039461
R640 VSS.n118 VSS.n113 0.0386493
R641 VSS.n107 VSS.n103 0.0386493
R642 VSS.n130 VSS.n129 0.0373384
R643 VSS.n159 VSS.n158 0.0356562
R644 VSS.n165 VSS.n161 0.0321558
R645 VSS.n153 VSS.n152 0.0306724
R646 VSS.n52 VSS.n51 0.0293149
R647 VSS.n30 VSS.n29 0.0263062
R648 VSS.n157 VSS.n156 0.0263062
R649 VSS.n28 VSS.n27 0.0236139
R650 VSS.n170 VSS.n169 0.0191688
R651 VSS.n56 VSS.n52 0.00902273
R652 VSS.n161 VSS.n160 0.00902273
R653 VSS.n135 VSS.n130 0.00523804
R654 VSS.n57 VSS.n56 0.00403904
R655 VSS.n51 VSS.n50 0.00293507
R656 VSS.n113 VSS.n112 0.00293507
R657 VSS.n103 VSS.n102 0.00293507
R658 VSS.n28 VSS.n11 0.00265517
R659 VSS.n155 VSS.n154 0.00243786
R660 VSS.n84 VSS.n80 0.00212338
R661 VSS.n75 VSS.n71 0.00212338
R662 VSS.n66 VSS.n65 0.00212338
R663 VSS.n95 VSS.n94 0.00160619
R664 VSS.n50 VSS.n45 0.00131169
R665 VSS.n124 VSS.n119 0.00131169
R666 VSS.n160 VSS.n135 0.000905844
R667 comp_outn.n0 comp_outn.t5 43.1877
R668 comp_outn.n1 comp_outn.t3 43.044
R669 comp_outn.n1 comp_outn.t4 43.044
R670 comp_outn comp_outn.t2 38.7789
R671 comp_outn.n4 comp_outn.t0 38.6969
R672 comp_outn.n4 comp_outn.t1 38.6969
R673 comp_outn.n2 comp_outn 1.15859
R674 comp_outn comp_outn.n4 0.984675
R675 comp_outn.n0 comp_outn 0.932565
R676 comp_outn.n5 comp_outn.n3 0.596088
R677 comp_outn.n5 comp_outn 0.438
R678 comp_outn.n2 comp_outn.n1 0.247153
R679 comp_outn comp_outn.n6 0.206382
R680 comp_outn.n3 comp_outn 0.15592
R681 comp_outn.n6 comp_outn 0.152674
R682 comp_outn.n6 comp_outn.n5 0.107118
R683 comp_outn.n2 comp_outn.n0 0.103441
R684 comp_outn.n5 comp_outn 0.063
R685 comp_outn.n3 comp_outn.n2 0.0193053
R686 cdac_vn.n0 cdac_vn.t6 350.253
R687 cdac_vn.n0 cdac_vn.t2 196.013
R688 cdac_vn.n1 cdac_vn.t0 196.013
R689 cdac_vn.n2 cdac_vn.t4 196.013
R690 cdac_vn.n3 cdac_vn.t3 196.013
R691 cdac_vn.n4 cdac_vn.t1 196.013
R692 cdac_vn.n5 cdac_vn.t7 196.013
R693 cdac_vn.n6 cdac_vn.t5 196.013
R694 cdac_vn.n6 cdac_vn.n5 154.24
R695 cdac_vn.n5 cdac_vn.n4 154.24
R696 cdac_vn.n4 cdac_vn.n3 154.24
R697 cdac_vn.n3 cdac_vn.n2 154.24
R698 cdac_vn.n2 cdac_vn.n1 154.24
R699 cdac_vn.n1 cdac_vn.n0 154.24
R700 cdac_vn cdac_vn.n6 65.4199
R701 cdac_vp.n0 cdac_vp.t1 350.253
R702 cdac_vp.n6 cdac_vp.t3 196.013
R703 cdac_vp.n5 cdac_vp.t2 196.013
R704 cdac_vp.n4 cdac_vp.t6 196.013
R705 cdac_vp.n3 cdac_vp.t4 196.013
R706 cdac_vp.n2 cdac_vp.t0 196.013
R707 cdac_vp.n1 cdac_vp.t7 196.013
R708 cdac_vp.n0 cdac_vp.t5 196.013
R709 cdac_vp.n1 cdac_vp.n0 154.24
R710 cdac_vp.n2 cdac_vp.n1 154.24
R711 cdac_vp.n3 cdac_vp.n2 154.24
R712 cdac_vp.n4 cdac_vp.n3 154.24
R713 cdac_vp.n5 cdac_vp.n4 154.24
R714 cdac_vp.n6 cdac_vp.n5 154.24
R715 cdac_vp cdac_vp.n6 61.3876
R716 comp_outp.n1 comp_outp.t5 43.3421
R717 comp_outp.n0 comp_outp.t3 43.044
R718 comp_outp.n0 comp_outp.t4 43.044
R719 comp_outp.n3 comp_outp.t2 39.1234
R720 comp_outp.n2 comp_outp.t0 38.6969
R721 comp_outp.n2 comp_outp.t1 38.6969
R722 comp_outp comp_outp.n4 14.0184
R723 comp_outp.n3 comp_outp.n2 1.09812
R724 comp_outp.n1 comp_outp.n0 1.00398
R725 comp_outp.n4 comp_outp.n3 0.449029
R726 comp_outp.n4 comp_outp.n1 0.294618
R727 clk.n4 clk.t4 356.68
R728 clk.n3 clk.t5 356.68
R729 clk.n1 clk.t1 269.921
R730 clk.n0 clk.t0 269.921
R731 clk.n4 clk.t2 202.44
R732 clk.n3 clk.t7 202.44
R733 clk.n1 clk.t6 195.721
R734 clk.n0 clk.t3 195.721
R735 clk.n5 clk.n4 41.3896
R736 clk.n5 clk.n3 41.3896
R737 clk.n2 clk.n0 38.0628
R738 clk.n2 clk.n1 38.0536
R739 clk.n6 clk.n5 12.3898
R740 clk clk.n6 8.69013
R741 clk.n6 clk.n2 3.40229
C0 a_1566_n378# a_582_n700# 0.00889f
C1 a_1566_n378# a_476_n1721# 0.117f
C2 a_564_n1721# a_564_n1266# 0.161f
C3 a_1566_n378# a_852_n296# 0.011f
C4 a_582_n700# VDD 0.0192f
C5 VDD a_476_n1721# 0.799f
C6 P a_1716_n1348# 9.22e-19
C7 cdac_vp a_564_n1266# 8.1e-19
C8 a_852_n296# VDD 0.78f
C9 a_1026_n1747# RS_n 7.1e-19
C10 P RS_p 8.56e-20
C11 a_1716_n1348# a_1026_n1747# 2.23e-21
C12 P Q 0.00291f
C13 a_1026_n1747# RS_p 0.144f
C14 a_1950_n1721# a_1026_n1747# 1.46e-19
C15 a_482_n1818# comp_outp 0.00346f
C16 P ready 1.69e-19
C17 a_582_n700# cdac_vn 0.426f
C18 cdac_vn a_476_n1721# 0.037f
C19 a_852_n296# cdac_vn 0.0563f
C20 cdac_vp a_1248_n288# 0.0187f
C21 a_1566_n378# comp_outp 6.13e-21
C22 ready a_1026_n1747# 0.0565f
C23 VDD comp_outp 0.671f
C24 clk a_582_n700# 0.0956f
C25 clk a_476_n1721# 0.459f
C26 a_564_n1721# cdac_vp 0.00295f
C27 clk a_852_n296# 0.0265f
C28 a_1566_n378# a_482_n1818# 0.0257f
C29 a_582_n700# RS_n 1.88e-19
C30 a_476_n1721# RS_n 0.00191f
C31 a_852_n296# RS_n 0.0212f
C32 VDD a_482_n1818# 1.48f
C33 a_582_n700# a_1716_n1348# 0.0758f
C34 a_1716_n1348# a_476_n1721# 0.0571f
C35 a_852_n296# a_1716_n1348# 0.215f
C36 a_582_n700# RS_p 2.41e-19
C37 a_476_n1721# RS_p 0.00222f
C38 cdac_vn comp_outp 0.0118f
C39 a_582_n700# Q 1.45f
C40 a_476_n1721# Q 0.00932f
C41 a_1566_n378# VDD 0.8f
C42 a_582_n700# a_1950_n1721# 5.87e-19
C43 a_852_n296# RS_p 0.158f
C44 a_1950_n1721# a_476_n1721# 5.72e-19
C45 a_852_n296# Q 9.24e-19
C46 a_1026_n1747# a_564_n1266# 1.23e-20
C47 clk comp_outp 0.00305f
C48 a_582_n700# ready 1.98e-19
C49 ready a_476_n1721# 0.0403f
C50 cdac_vn a_482_n1818# 0.0389f
C51 a_852_n296# ready 5.98e-19
C52 a_476_n1721# comp_outn 1.55e-19
C53 comp_outp RS_n 0.0437f
C54 a_1566_n378# cdac_vn 0.00873f
C55 a_1716_n1348# comp_outp 0.0993f
C56 P a_1248_n288# 0.133f
C57 clk a_482_n1818# 0.171f
C58 cdac_vn VDD 0.19f
C59 comp_outp RS_p 0.0759f
C60 comp_outp Q 7.56e-19
C61 a_1950_n1721# comp_outp 0.0559f
C62 a_482_n1818# RS_n 3.41e-20
C63 a_1566_n378# clk 0.525f
C64 cdac_vp P 0.224f
C65 a_1716_n1348# a_482_n1818# 0.197f
C66 clk VDD 0.772f
C67 a_564_n1721# a_1026_n1747# 0.0214f
C68 cdac_vp a_1026_n1747# 0.00718f
C69 a_1566_n378# RS_n 1.34e-19
C70 a_482_n1818# RS_p 4.35e-20
C71 ready comp_outp 1.69f
C72 a_482_n1818# Q 0.0247f
C73 a_476_n1721# a_564_n1266# 0.0214f
C74 a_1950_n1721# a_482_n1818# 1.15e-20
C75 a_1566_n378# a_1716_n1348# 0.135f
C76 VDD RS_n 0.581f
C77 a_852_n296# a_564_n1266# 1.58e-21
C78 comp_outp comp_outn 0.053f
C79 a_1716_n1348# VDD 0.786f
C80 a_1566_n378# RS_p 4.77e-20
C81 a_1566_n378# Q 0.155f
C82 VDD RS_p 0.536f
C83 VDD Q 0.368f
C84 ready a_482_n1818# 2.42e-20
C85 a_1950_n1721# VDD 0.767f
C86 clk cdac_vn 0.0494f
C87 a_1566_n378# ready 6.39e-21
C88 a_582_n700# a_1248_n288# 0.00749f
C89 cdac_vn RS_n 0.00684f
C90 a_476_n1721# a_1248_n288# 0.11f
C91 a_852_n296# a_1248_n288# 0.134f
C92 ready VDD 0.614f
C93 cdac_vn a_1716_n1348# 0.0947f
C94 VDD comp_outn 0.608f
C95 a_564_n1721# a_582_n700# 3.54e-19
C96 a_564_n1721# a_476_n1721# 0.386f
C97 cdac_vn RS_p 0.00693f
C98 a_564_n1721# a_852_n296# 0.00167f
C99 cdac_vn Q 0.216f
C100 cdac_vn a_1950_n1721# 0.0166f
C101 clk RS_n 0.00117f
C102 cdac_vp a_582_n700# 0.265f
C103 cdac_vp a_476_n1721# 0.484f
C104 cdac_vp a_852_n296# 0.087f
C105 clk a_1716_n1348# 0.113f
C106 a_482_n1818# a_564_n1266# 0.0164f
C107 clk RS_p 0.00116f
C108 clk Q 0.114f
C109 a_1716_n1348# RS_n 0.133f
C110 cdac_vn ready 0.00514f
C111 P a_1026_n1747# 3.42e-19
C112 cdac_vn comp_outn 0.00606f
C113 RS_n RS_p 0.314f
C114 comp_outp a_1248_n288# 4.23e-21
C115 RS_n Q 6.73e-20
C116 a_1950_n1721# RS_n 0.147f
C117 a_1716_n1348# RS_p 0.0744f
C118 VDD a_564_n1266# 5.28e-20
C119 a_1716_n1348# Q 0.141f
C120 a_1950_n1721# a_1716_n1348# 0.011f
C121 clk ready 2.93e-20
C122 a_564_n1721# comp_outp 0.00536f
C123 a_1950_n1721# RS_p 1.26e-19
C124 a_1950_n1721# Q 3.44e-19
C125 cdac_vp comp_outp 0.00146f
C126 ready RS_n 0.0795f
C127 a_482_n1818# a_1248_n288# 0.0534f
C128 RS_n comp_outn 1.64e-19
C129 a_1716_n1348# comp_outn 0.00481f
C130 a_564_n1721# a_482_n1818# 0.201f
C131 a_1566_n378# a_1248_n288# 0.406f
C132 ready RS_p 0.0658f
C133 cdac_vn a_564_n1266# 0.00183f
C134 ready a_1950_n1721# 0.0553f
C135 cdac_vp a_482_n1818# 0.207f
C136 RS_p comp_outn 8.63e-21
C137 VDD a_1248_n288# 0.851f
C138 a_1950_n1721# comp_outn 0.116f
C139 a_582_n700# P 1.45f
C140 P a_476_n1721# 0.0817f
C141 P a_852_n296# 0.142f
C142 a_1566_n378# cdac_vp 0.016f
C143 a_564_n1721# VDD 0.156f
C144 cdac_vp VDD 0.0194f
C145 a_582_n700# a_1026_n1747# 5.9e-19
C146 a_476_n1721# a_1026_n1747# 0.00774f
C147 ready comp_outn 0.0692f
C148 a_852_n296# a_1026_n1747# 0.0111f
C149 cdac_vn a_1248_n288# 9.58e-19
C150 a_564_n1266# RS_p 1.21e-21
C151 a_564_n1721# cdac_vn 0.00596f
C152 clk a_1248_n288# 0.602f
C153 cdac_vp cdac_vn 0.63f
C154 P comp_outp 1.61e-19
C155 comp_outp a_1026_n1747# 0.17f
C156 a_1716_n1348# a_1248_n288# 0.00907f
C157 cdac_vp clk 0.517f
C158 a_564_n1721# RS_n 3.53e-20
C159 a_582_n700# a_476_n1721# 0.0604f
C160 P a_482_n1818# 0.0143f
C161 a_1248_n288# RS_p 2.46e-19
C162 Q a_1248_n288# 0.195f
C163 a_582_n700# a_852_n296# 0.0763f
C164 a_852_n296# a_476_n1721# 0.309f
C165 a_564_n1721# a_1716_n1348# 1.33e-20
C166 cdac_vp RS_n 4.37e-20
C167 cdac_vp a_1716_n1348# 0.0393f
C168 a_482_n1818# a_1026_n1747# 2.77e-19
C169 a_564_n1721# RS_p 0.00175f
C170 a_1566_n378# P 0.194f
C171 a_564_n1721# a_1950_n1721# 3.46e-21
C172 P VDD 0.369f
C173 cdac_vp RS_p 4.07e-20
C174 cdac_vp Q 0.0612f
C175 ready a_1248_n288# 3.55e-21
C176 VDD a_1026_n1747# 0.762f
C177 a_564_n1721# ready 0.0708f
C178 cdac_vp ready 9.23e-19
C179 a_564_n1721# comp_outn 8.24e-22
C180 a_582_n700# comp_outp 0.00262f
C181 a_476_n1721# comp_outp 0.0165f
C182 a_852_n296# comp_outp 0.105f
C183 P cdac_vn 0.0279f
C184 cdac_vn a_1026_n1747# 0.0095f
C185 a_582_n700# a_482_n1818# 0.0121f
C186 a_482_n1818# a_476_n1721# 1.63f
C187 clk P 0.0966f
C188 a_852_n296# a_482_n1818# 0.042f
.ends

