* NGSPICE file created from hgu_sarlogic_sw_ctrl_flat.ext - technology: sky130A

.subckt hgu_sarlogic_sw_ctrl_flat VSS_SW[1] VSS_SW[2] VSS_SW[3] VSS_SW[4] VSS_SW[5]
+ VSS_SW[6] VSS_SW[7] VDD_SW[2] VDD_SW[3] VDD_SW[4] VDD_SW[5] VDD_SW[6] VDD_SW[7]
+ D[4] D[6] D[7] check[0] check[1] check[2] check[3] check[4] check[6] VDD_SW_b[1]
+ VDD_SW_b[2] VDD_SW_b[3] VDD_SW_b[4] VDD_SW_b[5] VDD_SW_b[6] VDD_SW_b[7] VSS_SW_b[1]
+ VSS_SW_b[2] VSS_SW_b[3] VSS_SW_b[4] VSS_SW_b[5] VSS_SW_b[6] VSS_SW_b[7] D[1] VDD_SW[1]
+ ready reset D[2] check[5] D[3] D[5] VSS VDD
X0 a_3420_212# x9.X VSS.t11 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VSS.t617 VDD.t753 a_10509_601# VSS.t616 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_11539_1642# VSS.t718 a_11325_1642# VDD.t475 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X3 VSS.t619 VDD.t754 a_7769_n62# VSS.t618 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X4 VDD.t57 a_15293_601# a_16024_909# VDD.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X5 VSS.t200 a_5812_212# a_5813_n88# VSS.t199 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6 a_5927_n62# a_5812_212# a_5504_106# VSS.t198 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X7 a_5323_2457# x30.A VSS.t670 VSS.t669 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VDD.t616 x3.X a_939_2457# VDD.t615 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_5271_n62# x2.X.t32 VSS.t504 VSS.t503 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X10 a_13300_993# a_11987_627# a_13216_993# VDD.t583 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VDD.t554 VDD.t552 a_10509_601# VDD.t553 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X12 VDD.t670 x16.X a_11987_627# VDD.t669 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X13 a_14887_1642# x9.A1.t32 a_14428_1467# VDD.t350 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X14 a_7896_106# a_8205_n88# a_8140_n62# VSS.t190 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X15 VSS.t285 a_9742_n88# VSS_SW_b[3].t0 VSS.t284 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X16 VSS.t333 a_14857_1289# a_14791_1315# VSS.t332 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 VDD.t649 a_1415_895# a_2136_627# VDD.t648 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X18 VDD.t622 a_8591_895# a_8516_993# VDD.t621 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X19 x7.X a_1757_1642# VSS.t416 VSS.t415 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X20 a_1501_122# a_1029_n88# a_1745_304# VDD.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X21 a_8933_1642# x9.A1.t33 a_8861_1642# VDD.t351 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X22 a_8933_1315# a_8679_1642# VSS.t308 VSS.t307 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X23 a_9154_1315# x9.A1.t34 a_8933_1642# VSS.t263 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X24 VSS.t68 D[6].t0 a_4338_n62# VSS.t67 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X25 VDD.t660 check[1].t0 a_13461_1642# VDD.t659 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X26 a_10983_895# a_10824_993# a_11123_627# VSS.t694 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X27 VSS.t615 check[1].t1 a_13461_1642# VSS.t614 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X28 VDD.t283 D[2].t0 a_13906_n62# VDD.t282 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X29 a_16298_n62# a_15381_n88# a_15853_122# VSS.t436 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X30 a_15518_304# a_15381_n88# a_15072_106# VDD.t438 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X31 VDD_SW_b[6].t1 a_3807_895# VDD.t572 VDD.t571 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X32 a_8731_627# a_8117_601# a_8591_895# VSS.t641 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X33 a_10041_993# a_9595_627# a_9949_627# VDD.t326 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X34 a_5462_220# a_5271_n62# VDD.t637 VDD.t636 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X35 VSS.t637 x16.X a_11987_627# VSS.t636 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X36 x9.A1.t15 a_5323_2457# VSS.t240 VSS.t239 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X37 a_15608_993# a_14545_627# a_15464_909# VDD.t741 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X38 a_9949_627# D[3].t0 VDD.t343 VDD.t342 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X39 VDD.t44 a_76_1467# x6.X VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X40 VDD.t55 a_15293_601# a_15243_909# VDD.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X41 a_8545_n62# a_8677_122# a_8409_n88# VSS.t301 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X42 a_11325_1642# x9.A1.t35 a_11253_1642# VDD.t272 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X43 VDD.t589 a_12134_n88# VSS_SW_b[2].t1 VDD.t588 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X44 a_15585_n88# a_15853_122# a_15799_220# VDD.t681 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X45 a_11325_1315# a_11071_1642# VSS.t292 VSS.t291 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X46 VDD.t444 a_13193_n88# a_13126_304# VDD.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X47 VDD.t701 x30.A a_5323_2457# VDD.t700 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X48 a_10532_n62# a_9742_n88# VSS.t283 VSS.t282 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X49 a_1028_212# x7.X VSS.t88 VSS.t87 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X50 a_5319_1642# x9.A1.t36 a_4860_1467# VDD.t273 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X51 a_10801_n88# a_10055_n62# a_10937_n62# VSS.t95 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X52 a_8921_304# a_8409_n88# VDD.t726 VDD.t725 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X53 VSS.t9 a_3420_212# a_3421_n88# VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X54 VSS.t535 a_5289_1289# a_5223_1315# VSS.t534 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X55 a_3807_895# x2.X.t33 VDD.t491 VDD.t490 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X56 a_15380_212# x20.X VSS.t631 VSS.t630 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X57 VSS.t318 a_7823_601# a_7757_627# VSS.t317 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X58 a_2773_627# D[6].t1 VSS.t70 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X59 a_12433_993# a_12153_627# a_12341_627# VSS.t696 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X60 VDD.t678 check[4].t0 a_6753_1642# VDD.t677 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X61 VSS.t621 VDD.t755 a_8545_n62# VSS.t620 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X62 a_12134_n88# a_12680_106# a_12638_220# VDD.t424 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X63 VSS.t643 check[4].t1 a_6760_1315# VSS.t642 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X64 VSS.t345 a_305_2457# x3.X VSS.t344 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X65 VDD.t254 a_12607_601# a_12517_993# VDD.t253 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X66 a_6753_1642# VSS.t719 a_6539_1642# VDD.t474 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X67 a_7757_627# a_7203_627# a_7649_993# VSS.t136 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X68 VDD_SW[4].t0 a_9312_627# VSS.t355 VSS.t354 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X69 VSS.t623 VDD.t756 a_8117_601# VSS.t622 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X70 VSS.t571 x3.X a_939_2457# VSS.t570 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X71 a_2927_1642# x9.A1.t37 a_2468_1467# VDD.t269 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X72 a_4862_90# a_4958_n88# VDD.t85 VDD.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X73 VDD.t262 a_13375_895# a_14096_627# VDD.t261 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X74 VSS.t275 D[7].t0 a_1946_n62# VSS.t274 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X75 a_487_n62# x2.X.t34 VSS.t359 VSS.t358 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X76 x30.A a_4689_2457# VDD.t750 VDD.t749 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X77 VDD.t247 a_5323_2457# x9.A1.t31 VDD.t246 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X78 x9.A1.t14 a_5323_2457# VSS.t238 VSS.t237 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X79 VSS.t151 a_2897_1289# a_2831_1315# VSS.t150 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X80 VDD.t385 check[3].t0 a_8679_1642# VDD.t384 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X81 VDD.t551 VDD.t549 a_1233_n88# VDD.t550 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X82 VDD.t87 a_7681_1289# a_7711_1642# VDD.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X83 VSS.t371 check[3].t1 a_8679_1642# VSS.t370 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X84 VDD.t685 check[0].t0 a_16323_1642# VDD.t684 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X85 VSS.t625 VDD.t757 a_941_601# VSS.t624 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X86 VSS.t654 check[0].t1 a_16330_1315# VSS.t653 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X87 a_6730_n62# a_5813_n88# a_6285_122# VSS.t140 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X88 a_10596_212# x15.X VDD.t93 VDD.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X89 a_5950_304# a_5813_n88# a_5504_106# VDD.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X90 a_15143_627# a_15293_601# a_14999_601# VSS.t50 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X91 a_3732_993# a_2419_627# a_3648_993# VDD.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X92 a_13126_304# a_12989_n88# a_12680_106# VDD.t209 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X93 VSS.t403 a_939_2457# x2.X.t15 VSS.t402 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X94 a_16323_1642# VSS.t720 a_16109_1642# VDD.t473 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X95 VDD.t548 VDD.t546 a_941_601# VDD.t547 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X96 a_3070_220# a_2879_n62# VDD.t22 VDD.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X97 VDD.t79 reset.t0 a_29_2457# VDD.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X98 a_13216_993# a_12153_627# a_13072_909# VDD.t729 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X99 a_7557_627# D[4].t0 VDD.t564 VDD.t563 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X100 VSS.t579 a_14428_1467# x18.X VSS.t578 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X101 a_14945_n62# a_15072_106# a_14526_n88# VSS.t302 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X102 x9.A1.t13 a_5323_2457# VSS.t236 VSS.t235 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X103 VSS.t577 a_8591_895# a_8539_627# VSS.t576 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X104 VDD.t643 a_6199_895# a_6124_993# VDD.t642 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X105 VSS.t702 a_7350_n88# VSS_SW_b[4].t0 VSS.t701 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X106 VDD_SW_b[1].t1 a_15767_895# VDD.t168 VDD.t167 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X107 VSS.t693 a_8409_n88# a_8319_n62# VSS.t692 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X108 a_13193_n88# a_13461_122# a_13407_220# VDD.t709 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X109 VDD.t699 x30.A a_5323_2457# VDD.t698 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X110 VSS.t401 a_939_2457# x2.X.t14 VSS.t400 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X111 a_678_220# a_487_n62# VDD.t320 VDD.t319 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X112 a_1415_895# x2.X.t35 VDD.t381 VDD.t380 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X113 VDD.t545 VDD.t543 a_8117_601# VDD.t544 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X114 a_9644_1467# VSS.t721 a_9786_1642# VDD.t472 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X115 a_12937_304# a_12134_n88# VDD.t587 VDD.t586 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X116 a_4862_90# a_4958_n88# VSS.t76 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X117 a_12988_212# x17.X VSS.t165 VSS.t164 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X118 VSS.t298 a_10983_895# a_11704_627# VSS.t297 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X119 VSS.t457 a_5431_601# a_5365_627# VSS.t456 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X120 a_15495_n62# a_15380_212# a_15072_106# VSS.t26 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X121 VSS.t25 a_15380_212# a_15381_n88# VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X122 VDD.t345 D[3].t1 a_11514_n62# VDD.t344 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X123 a_10041_993# a_9761_627# a_9949_627# VSS.t177 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X124 VSS.t627 VDD.t758 a_6153_n62# VSS.t626 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X125 VDD.t287 a_9644_1467# x14.X VDD.t286 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X126 a_9786_1642# check[2].t0 VDD.t383 VDD.t382 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X127 VDD.t355 a_14857_1289# a_14887_1642# VDD.t354 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X128 x2.X.t31 a_939_2457# VDD.t417 VDD.t416 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X129 a_9786_1315# check[2].t1 VSS.t363 VSS.t362 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X130 x17.X a_13715_1642# VDD.t188 VDD.t187 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X131 VDD.t708 a_10215_601# a_10125_993# VDD.t707 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X132 a_7769_n62# a_7896_106# a_7350_n88# VSS.t487 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X133 a_939_2457# x3.X VDD.t614 VDD.t613 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X134 VDD.t722 a_5725_601# a_5675_909# VDD.t721 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X135 a_5365_627# a_4811_627# a_5257_993# VSS.t103 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X136 VDD_SW[5].t0 a_6920_627# VSS.t717 VSS.t716 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X137 a_8140_n62# a_7350_n88# VSS.t700 VSS.t699 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X138 a_14733_627# D[1].t0 VSS.t551 VSS.t550 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X139 VDD.t245 a_5323_2457# x9.A1.t30 VDD.t244 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X140 a_6153_n62# a_6285_122# a_6017_n88# VSS.t523 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X141 VSS.t60 x3.A a_305_2457# VSS.t59 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X142 a_2470_90# a_2566_n88# VDD.t716 VDD.t715 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X143 a_8409_n88# a_7663_n62# a_8545_n62# VSS.t434 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X144 VSS.t273 D[2].t1 a_13906_n62# VSS.t272 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X145 a_11069_122# a_10597_n88# a_11313_304# VDD.t683 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X146 a_76_1467# x9.A1.t38 a_218_1315# VSS.t259 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X147 a_15799_220# a_14839_n62# VDD.t316 VDD.t315 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X148 x9.A1.t12 a_5323_2457# VSS.t234 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X149 VDD.t330 a_3333_601# a_4064_909# VDD.t329 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X150 a_10931_627# a_9761_627# a_10824_993# VSS.t176 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X151 a_6529_304# a_6017_n88# VDD.t42 VDD.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X152 VSS.t54 a_1028_212# a_1029_n88# VSS.t53 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X153 a_7615_1315# VSS.t485 a_7252_1467# VSS.t486 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X154 a_1340_993# a_27_627# a_1256_993# VDD.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X155 VDD.t243 a_5323_2457# x9.A1.t29 VDD.t242 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X156 a_1978_1315# x9.A1.t39 a_1757_1642# VSS.t260 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X157 a_12036_1467# VSS.t722 a_12178_1642# VDD.t471 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X158 a_5165_627# D[5].t0 VDD.t264 VDD.t263 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X159 x2.X.t30 a_939_2457# VDD.t415 VDD.t414 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X160 VSS.t399 a_939_2457# x2.X.t13 VSS.t398 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X161 VDD_SW[6].t1 a_4528_627# VDD.t656 VDD.t655 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X162 VSS.t598 a_6199_895# a_6147_627# VSS.t597 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X163 a_9742_n88# a_10288_106# a_10246_220# VDD.t445 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X164 a_15030_220# a_14839_n62# VDD.t314 VDD.t313 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X165 VSS.t74 a_4958_n88# VSS_SW_b[5].t0 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X166 VSS.t244 reset.t1 a_29_2457# VSS.t243 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X167 VDD.t542 VDD.t540 a_14526_n88# VDD.t541 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X168 VSS.t39 a_6017_n88# a_5927_n62# VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X169 a_8335_627# a_7823_601# VSS.t316 VSS.t315 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X170 a_8921_n62# a_8409_n88# VSS.t691 VSS.t690 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X171 x9.A1.t11 a_5323_2457# VSS.t232 VSS.t231 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X172 a_13715_1642# x9.A1.t40 a_13643_1642# VDD.t627 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X173 VSS.t290 a_2468_1467# x8.X VSS.t289 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X174 a_13715_1315# a_13461_1642# VSS.t92 VSS.t91 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X175 a_8848_909# a_8432_993# a_8591_895# VDD.t123 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X176 a_10545_304# a_9742_n88# VDD.t295 VDD.t294 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X177 a_2470_90# a_2566_n88# VSS.t685 VSS.t684 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X178 VDD.t697 x30.A a_5323_2457# VDD.t696 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X179 VSS.t397 a_939_2457# x2.X.t12 VSS.t396 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X180 VDD.t668 a_941_601# a_891_909# VDD.t667 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X181 a_581_627# a_27_627# a_473_993# VSS.t99 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X182 a_4338_n62# a_3421_n88# a_3893_122# VSS.t288 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X183 x9.A1.t10 a_5323_2457# VSS.t230 VSS.t229 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X184 a_5575_627# a_5725_601# a_5431_601# VSS.t689 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X185 a_13103_n62# a_12988_212# a_12680_106# VSS.t271 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X186 a_3558_304# a_3421_n88# a_3112_106# VDD.t298 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X187 VDD.t138 a_10596_212# a_10597_n88# VDD.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X188 a_15072_106# a_15381_n88# a_15316_n62# VSS.t435 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X189 x3.X a_305_2457# VDD.t369 VDD.t368 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X190 a_3648_993# a_2585_627# a_3504_909# VDD.t423 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X191 a_8677_122# a_8204_212# a_8921_n62# VSS.t608 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X192 a_5504_106# a_5812_212# a_5761_304# VDD.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X193 VSS.t325 a_12036_1467# x16.X VSS.t324 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X194 a_5377_n62# a_5504_106# a_4958_n88# VSS.t323 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X195 a_12341_627# D[2].t2 VSS.t124 VSS.t123 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X196 a_939_2457# x3.X VDD.t612 VDD.t611 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X197 VDD.t328 a_3333_601# a_3283_909# VDD.t327 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X198 a_7350_n88# a_7663_n62# a_7769_n62# VSS.t433 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X199 a_5675_909# a_5257_993# a_5431_601# VDD.t742 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X200 a_7967_627# x2.X.t36 VSS.t361 VSS.t360 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X201 VDD.t241 a_5323_2457# x9.A1.t28 VDD.t240 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X202 VDD.t160 a_2897_1289# a_2927_1642# VDD.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X203 a_10801_n88# a_11069_122# a_11015_220# VDD.t189 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X204 VDD.t239 a_5323_2457# x9.A1.t27 VDD.t238 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X205 a_9761_627# a_9595_627# VDD.t325 VDD.t324 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X206 a_13407_220# a_12447_n62# VDD.t361 VDD.t360 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X207 a_381_627# D[7].t1 VDD.t285 VDD.t284 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X208 VSS.t48 a_647_601# a_581_627# VSS.t47 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X209 VSS.t575 a_8591_895# a_9312_627# VSS.t574 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X210 VDD.t489 check[2].t2 a_11539_1642# VDD.t488 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X211 a_14430_90# a_14526_n88# VDD.t122 VDD.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X212 a_8204_212# x13.X VDD.t421 VDD.t420 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X213 VDD.t566 D[4].t1 a_9122_n62# VDD.t565 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X214 VSS.t498 check[2].t3 a_11546_1315# VSS.t497 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X215 VSS.t629 VDD.t759 a_14945_n62# VSS.t628 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X216 VSS.t175 a_174_n88# VSS_SW_b[7].t0 VSS.t174 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X217 VSS.t186 a_3039_601# a_2973_627# VSS.t185 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X218 x13.X a_8933_1642# VSS.t22 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X219 VSS.t270 a_12988_212# a_12989_n88# VSS.t269 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X220 VDD.t237 a_5323_2457# x9.A1.t26 VDD.t236 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X221 VSS.t343 a_305_2457# x3.X VSS.t342 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X222 VDD_SW[7].t1 a_2136_627# VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X223 VDD_SW_b[5].t0 a_6199_895# VSS.t596 VSS.t595 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X224 VDD.t539 VDD.t537 a_4958_n88# VDD.t538 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X225 a_8677_122# a_8205_n88# a_8921_304# VDD.t199 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X226 VSS.t395 a_939_2457# x2.X.t11 VSS.t394 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X227 a_16037_1642# a_15855_1642# VDD.t453 VDD.t452 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X228 a_14857_1289# check[0].t2 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X229 VDD_SW[1].t1 a_16488_627# VDD.t604 VDD.t603 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X230 x30.A a_4689_2457# VDD.t748 VDD.t747 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X231 a_791_627# a_941_601# a_647_601# VSS.t635 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X232 x2.X.t29 a_939_2457# VDD.t413 VDD.t412 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X233 a_14857_1289# check[0].t3 VSS.t13 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X234 a_4149_1642# VSS.t483 a_4149_1315# VSS.t484 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X235 x20.X a_16109_1642# VDD.t213 VDD.t212 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X236 a_7823_601# x2.X.t37 VDD.t89 VDD.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X237 a_9761_627# a_9595_627# VSS.t312 VSS.t311 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X238 a_6456_909# a_6040_993# a_6199_895# VDD.t296 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X239 VSS.t28 D[3].t2 a_11514_n62# VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X240 x9.A1.t9 a_5323_2457# VSS.t228 VSS.t227 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X241 a_8731_627# x2.X.t38 VSS.t80 VSS.t79 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X242 a_891_909# a_473_993# a_647_601# VDD.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X243 a_3183_627# a_3333_601# a_3039_601# VSS.t314 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X244 a_10824_993# a_9595_627# a_10727_627# VSS.t310 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X245 VSS.t393 a_939_2457# x2.X.t10 VSS.t392 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X246 a_1166_304# a_1029_n88# a_720_106# VDD.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X247 a_10983_895# x2.X.t39 VDD.t91 VDD.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X248 a_5431_601# a_5257_993# a_5575_627# VSS.t707 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X249 a_14430_90# a_14526_n88# VSS.t115 VSS.t114 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X250 VDD.t5 a_9646_90# VSS_SW[3].t1 VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X251 a_1256_993# a_193_627# a_1112_909# VDD.t428 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X252 a_6285_122# a_5812_212# a_6529_n62# VSS.t197 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X253 VSS.t182 a_4862_90# VSS_SW[5].t0 VSS.t181 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X254 a_3112_106# a_3420_212# a_3369_304# VDD.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X255 VSS.t1 x27.A a_4689_2457# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X256 a_12465_1289# check[1].t2 VDD.t375 VDD.t374 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X257 a_2985_n62# a_3112_106# a_2566_n88# VSS.t93 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X258 VDD.t170 check[6].t0 a_1971_1642# VDD.t169 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X259 a_7252_1467# x9.A1.t41 a_7394_1315# VSS.t582 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X260 a_12465_1289# check[1].t3 VSS.t351 VSS.t350 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X261 a_5896_909# a_5431_601# VDD.t459 VDD.t458 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X262 a_15907_627# a_15293_601# a_15767_895# VSS.t49 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X263 a_1757_1642# VSS.t481 a_1757_1315# VSS.t482 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X264 VSS.t161 check[6].t1 a_1978_1315# VSS.t160 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X265 a_3283_909# a_2865_993# a_3039_601# VDD.t654 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X266 a_5575_627# x2.X.t40 VSS.t32 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X267 a_1233_n88# a_1501_122# a_1447_220# VDD.t481 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X268 a_939_2457# x3.X VDD.t610 VDD.t609 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X269 a_6529_n62# a_6017_n88# VSS.t37 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X270 a_8153_304# a_7350_n88# VDD.t735 VDD.t734 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X271 VSS.t391 a_939_2457# x2.X.t9 VSS.t390 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X272 a_8539_627# a_7369_627# a_8432_993# VSS.t86 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X273 a_12038_90# a_12134_n88# VDD.t585 VDD.t584 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X274 a_7733_993# a_7369_627# a_7649_993# VDD.t97 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X275 a_5812_212# x11.X VDD.t289 VDD.t288 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X276 VSS.t537 VDD.t760 a_5377_n62# VSS.t536 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X277 VDD.t739 a_12901_601# a_13632_909# VDD.t738 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X278 VDD.t653 a_8204_212# a_8205_n88# VDD.t652 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X279 a_593_n62# a_720_106# a_174_n88# VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X280 a_2831_1315# VSS.t479 a_2468_1467# VSS.t480 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X281 VDD.t46 ready.t0 a_4413_2457# VDD.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X282 a_3535_n62# a_3420_212# a_3112_106# VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X283 x2.X.t28 a_939_2457# VDD.t411 VDD.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X284 a_16097_304# a_15585_n88# VDD.t154 VDD.t153 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X285 VSS.t349 a_14999_601# a_14933_627# VSS.t348 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X286 a_5504_106# a_5813_n88# a_5748_n62# VSS.t139 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X287 VDD_SW_b[6].t0 a_3807_895# VSS.t518 VSS.t517 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X288 a_16330_1315# x9.A1.t42 a_16109_1642# VSS.t583 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X289 a_7663_n62# x2.X.t41 VDD.t30 VDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X290 VSS.t159 a_15767_895# a_15715_627# VSS.t158 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X291 VDD.t235 a_5323_2457# x9.A1.t25 VDD.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X292 a_5323_2457# x30.A VSS.t668 VSS.t667 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X293 VDD.t536 VDD.t534 a_8409_n88# VDD.t535 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X294 VSS.t145 a_15585_n88# a_15495_n62# VSS.t144 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X295 VSS.t41 a_76_1467# x6.X VSS.t40 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X296 a_4958_n88# a_5271_n62# a_5377_n62# VSS.t592 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X297 VDD_SW[2].t1 a_14096_627# VDD.t310 VDD.t309 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X298 a_5431_601# x2.X.t42 VDD.t32 VDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X299 a_4064_909# a_3648_993# a_3807_895# VDD.t704 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X300 a_3839_220# a_2879_n62# VDD.t20 VDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X301 x2.X.t27 a_939_2457# VDD.t409 VDD.t408 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X302 a_4077_1642# a_3895_1642# VDD.t672 VDD.t671 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X303 a_7369_627# a_7203_627# VDD.t143 VDD.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X304 a_14428_1467# x9.A1.t43 a_14570_1315# VSS.t554 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X305 a_2897_1289# check[5].t0 VDD.t357 VDD.t356 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X306 VDD.t664 x14.X a_9595_627# VDD.t663 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X307 VDD.t533 VDD.t531 a_174_n88# VDD.t532 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X308 VDD.t233 a_5323_2457# x9.A1.t24 VDD.t232 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X309 x9.A1.t8 a_5323_2457# VSS.t226 VSS.t225 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X310 a_2897_1289# check[5].t1 VSS.t335 VSS.t334 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X311 a_791_627# x2.X.t43 VSS.t105 VSS.t104 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X312 a_13906_n62# a_12989_n88# a_13461_122# VSS.t202 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X313 x9.X a_4149_1642# VDD.t101 VDD.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X314 a_10908_993# a_9595_627# a_10824_993# VDD.t323 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X315 a_12038_90# a_12134_n88# VSS.t533 VSS.t532 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X316 VDD.t626 a_7254_90# VSS_SW[4].t1 VDD.t625 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X317 a_2879_n62# x2.X.t44 VSS.t107 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X318 a_720_106# a_1028_212# a_977_304# VDD.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X319 VSS.t449 a_2470_90# VSS_SW[6].t0 VSS.t448 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X320 VDD_SW_b[7].t1 a_1415_895# VDD.t647 VDD.t646 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X321 a_6339_627# a_5725_601# a_6199_895# VSS.t688 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X322 a_3504_909# a_3039_601# VDD.t195 VDD.t194 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X323 VDD.t530 VDD.t528 a_2566_n88# VDD.t529 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X324 a_3183_627# x2.X.t45 VSS.t109 VSS.t108 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X325 a_15072_106# a_15380_212# a_15329_304# VDD.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X326 VSS.t500 D[4].t2 a_9122_n62# VSS.t499 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X327 VSS.t389 a_939_2457# x2.X.t8 VSS.t388 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X328 a_12495_1642# x9.A1.t44 a_12036_1467# VDD.t598 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X329 a_1685_1642# a_1503_1642# VDD.t432 VDD.t431 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X330 VSS.t453 a_12465_1289# a_12399_1315# VSS.t452 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X331 a_6147_627# a_4977_627# a_6040_993# VSS.t672 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X332 a_15243_909# a_14825_993# a_14999_601# VDD.t215 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X333 a_218_1642# check[6].t2 VDD.t485 VDD.t484 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X334 a_647_601# a_473_993# a_791_627# VSS.t62 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X335 a_5341_993# a_4977_627# a_5257_993# VDD.t703 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X336 a_7369_627# a_7203_627# VSS.t135 VSS.t134 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X337 a_8432_993# a_7203_627# a_8335_627# VSS.t133 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X338 VDD.t576 a_10509_601# a_11240_909# VDD.t575 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X339 a_218_1315# check[6].t3 VSS.t494 VSS.t493 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X340 VSS.t633 x14.X a_9595_627# VSS.t632 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X341 a_13929_1642# VSS.t723 a_13715_1642# VDD.t470 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X342 a_1143_n62# a_1028_212# a_720_106# VSS.t52 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X343 a_174_n88# a_487_n62# a_593_n62# VSS.t306 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X344 a_6339_627# x2.X.t46 VSS.t489 VSS.t488 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X345 a_3112_106# a_3421_n88# a_3356_n62# VSS.t287 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X346 a_647_601# x2.X.t47 VDD.t478 VDD.t477 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X347 a_3039_601# a_2865_993# a_3183_627# VSS.t609 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X348 VDD.t293 a_9742_n88# VSS_SW_b[3].t1 VDD.t292 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X349 VSS.t353 ready.t1 a_4413_2457# VSS.t352 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X350 a_16298_n62# a_15380_212# a_15853_122# VDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X351 a_5271_n62# x2.X.t48 VDD.t480 VDD.t479 sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X352 VSS.t442 a_13193_n88# a_13103_n62# VSS.t441 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X353 VDD.t527 VDD.t525 a_6017_n88# VDD.t526 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X354 VDD.t256 check[0].t4 a_15855_1642# VDD.t255 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X355 a_4860_1467# x9.A1.t45 a_5002_1315# VSS.t555 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X356 VSS.t250 check[0].t5 a_15855_1642# VSS.t249 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X357 a_15511_627# a_14999_601# VSS.t347 VSS.t346 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X358 a_5323_2457# x30.A VSS.t666 VSS.t665 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X359 a_15316_n62# a_14526_n88# VSS.t113 VSS.t112 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X360 a_2566_n88# a_2879_n62# a_2985_n62# VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X361 VSS.t539 VDD.t761 a_593_n62# VSS.t538 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X362 VDD_SW_b[1].t0 a_15767_895# VSS.t157 VSS.t156 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X363 VDD.t308 a_10983_895# a_11704_627# VDD.t307 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X364 a_4370_1315# x9.A1.t46 a_4149_1642# VSS.t586 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X365 a_8591_895# a_8432_993# a_8731_627# VSS.t116 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X366 a_3039_601# x2.X.t49 VDD.t203 VDD.t202 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X367 x3.X a_305_2457# VSS.t341 VSS.t340 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X368 VDD.t562 a_10801_n88# a_10734_304# VDD.t561 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X369 a_1447_220# a_487_n62# VDD.t318 VDD.t317 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X370 a_16024_909# a_15608_993# a_15767_895# VDD.t710 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X371 a_6539_1642# VSS.t477 a_6539_1315# VSS.t478 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X372 VDD.t201 x12.X a_7203_627# VDD.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X373 VSS.t541 VDD.t762 a_2985_n62# VSS.t540 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X374 x2.X.t26 a_939_2457# VDD.t407 VDD.t406 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X375 VDD.t746 a_4689_2457# x30.A VDD.t745 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X376 VSS.t569 x3.X a_939_2457# VSS.t568 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X377 a_11514_n62# a_10597_n88# a_11069_122# VSS.t648 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X378 a_7649_993# a_7203_627# a_7557_627# VDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X379 a_2468_1467# x9.A1.t47 a_2610_1315# VSS.t587 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X380 a_10824_993# a_9761_627# a_10680_909# VDD.t186 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X381 VSS.t277 a_9644_1467# x14.X VSS.t276 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X382 a_1112_909# a_647_601# VDD.t53 VDD.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X383 a_14839_n62# x2.X.t50 VSS.t194 VSS.t193 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X384 VSS.t256 a_13375_895# a_13323_627# VSS.t255 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X385 VDD_SW_b[2].t1 a_13375_895# VDD.t260 VDD.t259 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X386 x2.X.t7 a_939_2457# VSS.t387 VSS.t386 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X387 x17.X a_13715_1642# VSS.t179 VSS.t178 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X388 a_16109_1642# VSS.t475 a_16109_1315# VSS.t476 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X389 a_12680_106# a_12988_212# a_12937_304# VDD.t281 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X390 VSS.t188 a_14430_90# VSS_SW[1].t0 VSS.t187 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X391 a_15853_122# a_15380_212# a_16097_n62# VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X392 VSS.t543 VDD.t763 a_5725_601# VSS.t542 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X393 a_15464_909# a_14999_601# VDD.t373 VDD.t372 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X394 a_15143_627# x2.X.t51 VSS.t196 VSS.t195 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X395 a_6040_993# a_4811_627# a_5943_627# VSS.t102 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X396 a_16097_n62# a_15585_n88# VSS.t143 VSS.t142 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X397 VSS.t192 x12.X a_7203_627# VSS.t191 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X398 a_8516_993# a_7203_627# a_8432_993# VDD.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X399 VDD.t524 VDD.t522 a_5725_601# VDD.t523 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X400 a_10596_212# x15.X VSS.t82 VSS.t81 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X401 a_11546_1315# x9.A1.t48 a_11325_1642# VSS.t588 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X402 VDD.t591 a_5289_1289# a_5319_1642# VDD.t590 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X403 a_5323_2457# x30.A VDD.t695 VDD.t694 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X404 VSS.t545 VDD.t764 a_3761_n62# VSS.t544 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X405 VSS.t715 a_4689_2457# x30.A VSS.t714 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X406 a_193_627# a_27_627# VDD.t111 VDD.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X407 a_2973_627# a_2419_627# a_2865_993# VSS.t149 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X408 VDD_SW[6].t0 a_4528_627# VSS.t611 VSS.t610 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X409 a_12553_n62# a_12680_106# a_12134_n88# VSS.t410 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X410 a_557_993# a_193_627# a_473_993# VDD.t427 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X411 a_3947_627# a_3333_601# a_3807_895# VSS.t313 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X412 a_14999_601# a_14825_993# a_15143_627# VSS.t208 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X413 a_14526_n88# a_14839_n62# a_14945_n62# VSS.t304 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X414 a_3761_n62# a_3893_122# a_3625_n88# VSS.t61 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X415 a_6199_895# a_6040_993# a_6339_627# VSS.t286 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X416 VDD.t172 check[5].t2 a_3895_1642# VDD.t171 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X417 a_14791_1315# VSS.t473 a_14428_1467# VSS.t474 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X418 a_4149_1642# x9.A1.t49 a_4077_1642# VDD.t249 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X419 VSS.t163 check[5].t3 a_3895_1642# VSS.t162 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X420 a_6467_1642# a_6285_1642# VDD.t556 VDD.t555 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X421 VDD.t666 a_941_601# a_1672_909# VDD.t665 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X422 a_7649_993# a_7369_627# a_7557_627# VSS.t85 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X423 a_6017_n88# a_5271_n62# a_6153_n62# VSS.t591 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X424 a_4149_1315# a_3895_1642# VSS.t639 VSS.t638 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X425 a_14999_601# x2.X.t52 VDD.t600 VDD.t599 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X426 a_5257_993# a_4811_627# a_5165_627# VDD.t116 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X427 VSS.t167 a_78_90# VSS_SW[7].t0 VSS.t166 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X428 a_487_n62# x2.X.t53 VDD.t602 VDD.t601 sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X429 VDD.t334 a_7823_601# a_7733_993# VDD.t333 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X430 x11.X a_6539_1642# VDD.t658 VDD.t657 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X431 a_7252_1467# VSS.t724 a_7394_1642# VDD.t469 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X432 a_2773_627# D[6].t2 VDD.t67 VDD.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X433 a_4137_304# a_3625_n88# VDD.t65 VDD.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X434 a_193_627# a_27_627# VSS.t98 VSS.t97 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X435 VDD.t620 a_8591_895# a_9312_627# VDD.t619 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X436 a_6730_n62# a_5812_212# a_6285_122# VDD.t206 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X437 a_720_106# a_1029_n88# a_964_n62# VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X438 VSS.t516 a_3807_895# a_3755_627# VSS.t515 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X439 a_12447_n62# x2.X.t54 VSS.t557 VSS.t556 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X440 VDD.t733 a_7350_n88# VSS_SW_b[4].t1 VDD.t732 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X441 VSS.t683 a_2566_n88# VSS_SW_b[6].t0 VSS.t682 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X442 x9.A1.t23 a_5323_2457# VDD.t231 VDD.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X443 VDD.t521 VDD.t519 a_12134_n88# VDD.t520 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X444 VSS.t58 a_3625_n88# a_3535_n62# VSS.t57 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X445 a_15853_122# a_15381_n88# a_16097_304# VDD.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X446 VDD.t724 a_8409_n88# a_8342_304# VDD.t723 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X447 VDD.t449 a_7252_1467# x12.X VDD.t448 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X448 a_7394_1642# check[3].t2 VDD.t633 VDD.t632 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X449 VDD.t455 a_12465_1289# a_12495_1642# VDD.t454 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X450 a_5943_627# a_5431_601# VSS.t455 VSS.t454 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X451 a_13119_627# a_12607_601# VSS.t248 VSS.t247 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X452 a_1757_1642# x9.A1.t50 a_1685_1642# VDD.t250 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X453 a_7394_1315# check[3].t3 VSS.t590 VSS.t589 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X454 a_5748_n62# a_4958_n88# VSS.t72 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X455 x2.X.t6 a_939_2457# VSS.t385 VSS.t384 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X456 VSS.t547 VDD.t765 a_3333_601# VSS.t546 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X457 VDD.t166 a_15767_895# a_15692_993# VDD.t165 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X458 a_13072_909# a_12607_601# VDD.t252 VDD.t251 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X459 a_1757_1315# a_1503_1642# VSS.t418 VSS.t417 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X460 a_15715_627# a_14545_627# a_15608_993# VSS.t706 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X461 a_9122_n62# a_8205_n88# a_8677_122# VSS.t189 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X462 a_6124_993# a_4811_627# a_6040_993# VDD.t115 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X463 VSS.t567 x3.X a_939_2457# VSS.t566 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X464 VDD.t518 VDD.t516 a_3333_601# VDD.t517 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X465 a_10711_n62# a_10596_212# a_10288_106# VSS.t131 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X466 a_7350_n88# a_7896_106# a_7854_220# VDD.t476 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X467 a_1946_n62# a_1029_n88# a_1501_122# VSS.t43 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0675 ps=0.735 w=0.36 l=0.15
X468 a_15907_627# x2.X.t55 VSS.t365 VSS.t364 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X469 VDD.t447 a_4860_1467# x10.X VDD.t446 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X470 a_5002_1642# check[4].t2 VDD.t353 VDD.t352 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X471 a_5002_1315# check[4].t3 VSS.t331 VSS.t330 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X472 a_5223_1315# VSS.t471 a_4860_1467# VSS.t472 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X473 a_9147_1642# VSS.t725 a_8933_1642# VDD.t468 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X474 VDD_SW[7].t0 a_2136_627# VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X475 VSS.t549 VDD.t766 a_15721_n62# VSS.t548 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X476 a_10161_n62# a_10288_106# a_9742_n88# VSS.t443 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0864 ps=0.91 w=0.64 l=0.15
X477 VDD_SW_b[3].t1 a_10983_895# VDD.t306 VDD.t305 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X478 a_12638_220# a_12447_n62# VDD.t359 VDD.t358 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X479 VSS.t262 a_12038_90# VSS_SW[2].t0 VSS.t261 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X480 VDD.t367 a_305_2457# x3.X VDD.t366 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X481 a_473_993# a_27_627# a_381_627# VDD.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X482 a_3807_895# a_3648_993# a_3947_627# VSS.t673 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X483 a_14933_627# a_14379_627# a_14825_993# VSS.t122 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X484 VDD.t608 x3.X a_939_2457# VDD.t607 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X485 a_6760_1315# x9.A1.t51 a_6539_1642# VSS.t242 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X486 VSS.t594 a_6199_895# a_6920_627# VSS.t593 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X487 a_15329_304# a_14526_n88# VDD.t120 VDD.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X488 a_11015_220# a_10055_n62# VDD.t108 VDD.t107 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X489 VDD_SW[1].t0 a_16488_627# VSS.t559 VSS.t558 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X490 a_15721_n62# a_15853_122# a_15585_n88# VSS.t646 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X491 a_5257_993# a_4977_627# a_5165_627# VSS.t671 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X492 VDD.t266 D[5].t1 a_6730_n62# VDD.t265 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X493 x9.A1.t22 a_5323_2457# VDD.t229 VDD.t228 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X494 x20.X a_16109_1642# VSS.t206 VSS.t205 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X495 VSS.t420 VDD.t767 a_12553_n62# VSS.t419 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X496 a_14909_993# a_14545_627# a_14825_993# VDD.t740 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X497 a_535_1642# x9.A1.t52 a_76_1467# VDD.t460 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X498 VDD.t457 a_5431_601# a_5341_993# VDD.t456 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X499 a_964_n62# a_174_n88# VSS.t173 VSS.t172 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X500 VSS.t169 a_505_1289# a_439_1315# VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X501 VSS.t130 a_10596_212# a_10597_n88# VSS.t129 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X502 a_12680_106# a_12989_n88# a_12924_n62# VSS.t201 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X503 a_4338_n62# a_3420_212# a_3893_122# VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X504 VDD.t405 a_939_2457# x2.X.t25 VDD.t404 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X505 a_10055_n62# x2.X.t56 VSS.t367 VSS.t366 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X506 VDD.t83 a_4958_n88# VSS_SW_b[5].t1 VDD.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X507 VDD.t515 VDD.t513 a_9742_n88# VDD.t514 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X508 a_8409_n88# a_8677_122# a_8623_220# VDD.t311 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X509 VDD.t40 a_6017_n88# a_5950_304# VDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X510 VSS.t322 a_1233_n88# a_1143_n62# VSS.t321 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X511 a_3551_627# a_3039_601# VSS.t184 VSS.t183 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X512 a_14733_627# D[1].t1 VDD.t593 VDD.t592 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X513 x9.A1.t21 a_5323_2457# VDD.t227 VDD.t226 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X514 VSS.t664 x30.A a_5323_2457# VSS.t663 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X515 a_3356_n62# a_2566_n88# VSS.t681 VSS.t680 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X516 VSS.t111 a_14526_n88# VSS_SW_b[1].t0 VSS.t110 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X517 VDD.t258 a_13375_895# a_13300_993# VDD.t257 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X518 a_13323_627# a_12153_627# a_13216_993# VSS.t695 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X519 VDD.t75 check[6].t4 a_1503_1642# VDD.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X520 a_12399_1315# VSS.t469 a_12036_1467# VSS.t470 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X521 VSS.t64 check[6].t5 a_1503_1642# VSS.t63 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X522 a_8204_212# x13.X VSS.t407 VSS.t406 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X523 VSS.t422 VDD.t768 a_15293_601# VSS.t421 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X524 VDD.t403 a_939_2457# x2.X.t24 VDD.t402 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X525 a_13515_627# x2.X.t57 VSS.t369 VSS.t368 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X526 a_13936_1315# x9.A1.t53 a_13715_1642# VSS.t458 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X527 VDD.t512 VDD.t510 a_15293_601# VDD.t511 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X528 a_9949_627# D[3].t3 VSS.t30 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X529 VSS.t424 VDD.t769 a_13329_n62# VSS.t423 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X530 a_7681_1289# check[3].t4 VDD.t268 VDD.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X531 VSS.t604 a_1415_895# a_1363_627# VSS.t603 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X532 a_10246_220# a_10055_n62# VDD.t106 VDD.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X533 a_3893_122# a_3420_212# a_4137_n62# VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X534 a_13515_627# a_12901_601# a_13375_895# VSS.t704 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X535 a_7681_1289# check[3].t5 VSS.t258 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X536 a_6285_122# a_5813_n88# a_6529_304# VDD.t148 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X537 a_15767_895# a_15608_993# a_15907_627# VSS.t679 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X538 x30.A a_4689_2457# VSS.t713 VSS.t712 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X539 VSS.t224 a_5323_2457# x9.A1.t7 VSS.t223 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X540 a_5761_304# a_4958_n88# VDD.t81 VDD.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X541 VDD_SW[2].t0 a_14096_627# VSS.t300 VSS.t299 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X542 a_12541_627# a_11987_627# a_12433_993# VSS.t527 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X543 VSS.t514 a_3807_895# a_4528_627# VSS.t513 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X544 VDD.t737 a_12901_601# a_12851_909# VDD.t736 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X545 VDD.t71 x3.A a_305_2457# VDD.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X546 a_76_1467# VSS.t726 a_218_1642# VDD.t467 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X547 a_13329_n62# a_13461_122# a_13193_n88# VSS.t678 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X548 a_15585_n88# a_14839_n62# a_15721_n62# VSS.t303 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X549 a_4137_n62# a_3625_n88# VSS.t56 VSS.t55 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X550 a_3420_212# x9.X VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X551 VDD.t184 a_174_n88# VSS_SW_b[7].t1 VDD.t183 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X552 a_12517_993# a_12153_627# a_12433_993# VDD.t728 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X553 a_6539_1642# x9.A1.t54 a_6467_1642# VDD.t461 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X554 a_8591_895# x2.X.t58 VDD.t145 VDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X555 a_6539_1315# a_6285_1642# VSS.t506 VSS.t505 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X556 VDD.t205 a_5812_212# a_5813_n88# VDD.t204 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X557 a_14825_993# a_14379_627# a_14733_627# VDD.t129 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X558 x9.A1.t20 a_5323_2457# VDD.t225 VDD.t224 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X559 a_13705_304# a_13193_n88# VDD.t442 VDD.t441 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X560 VDD_SW_b[4].t1 a_8591_895# VDD.t618 VDD.t617 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X561 x9.X a_4149_1642# VSS.t90 VSS.t89 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X562 a_10288_106# a_10597_n88# a_10532_n62# VSS.t647 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.066 ps=0.745 w=0.36 l=0.15
X563 a_6017_n88# a_6285_122# a_6231_220# VDD.t579 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X564 a_8623_220# a_7663_n62# VDD.t436 VDD.t435 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X565 VSS.t246 a_12607_601# a_12541_627# VSS.t245 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X566 a_12341_627# D[2].t3 VDD.t131 VDD.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X567 VDD.t401 a_939_2457# x2.X.t23 VDD.t400 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X568 a_11253_1642# a_11071_1642# VDD.t302 VDD.t301 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X569 a_16109_1642# x9.A1.t55 a_16037_1642# VDD.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X570 a_473_993# a_193_627# a_381_627# VSS.t414 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X571 VDD_SW_b[7].t0 a_1415_895# VSS.t602 VSS.t601 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X572 a_9646_90# a_9742_n88# VDD.t291 VDD.t290 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X573 VDD_SW[3].t1 a_11704_627# VDD.t718 VDD.t717 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X574 VSS.t531 a_12134_n88# VSS_SW_b[2].t0 VSS.t530 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X575 a_10073_1289# check[2].t4 VDD.t77 VDD.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X576 a_16109_1315# a_15855_1642# VSS.t451 VSS.t450 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X577 x9.A1.t19 a_5323_2457# VDD.t223 VDD.t222 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X578 VSS.t662 x30.A a_5323_2457# VSS.t661 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X579 a_10073_1289# check[2].t5 VSS.t66 VSS.t65 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X580 x15.X a_11325_1642# VDD.t277 VDD.t276 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X581 VDD.t51 a_647_601# a_557_993# VDD.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X582 a_1672_909# a_1256_993# a_1415_895# VDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X583 a_4977_627# a_4811_627# VDD.t114 VDD.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X584 a_5812_212# x11.X VSS.t279 VSS.t278 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X585 VSS.t607 a_8204_212# a_8205_n88# VSS.t606 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X586 a_8319_n62# a_8204_212# a_7896_106# VSS.t605 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.0486 ps=0.63 w=0.36 l=0.15
X587 a_11123_627# x2.X.t59 VSS.t138 VSS.t137 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X588 VDD.t399 a_939_2457# x2.X.t22 VDD.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X589 x2.X.t5 a_939_2457# VSS.t383 VSS.t382 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X590 VDD.t193 a_3039_601# a_2949_993# VDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X591 VDD.t191 a_4862_90# VSS_SW[5].t1 VDD.t190 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X592 a_7557_627# D[4].t3 VSS.t502 VSS.t501 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X593 x9.A1.t18 a_5323_2457# VDD.t221 VDD.t220 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X594 a_12751_627# a_12901_601# a_12607_601# VSS.t703 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X595 a_939_2457# x3.X VSS.t565 VSS.t564 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X596 VSS.t222 a_5323_2457# x9.A1.t6 VSS.t221 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X597 a_10734_304# a_10597_n88# a_10288_106# VDD.t682 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X598 a_11123_627# a_10509_601# a_10983_895# VSS.t520 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X599 VSS.t650 D[5].t2 a_6730_n62# VSS.t649 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X600 a_3893_122# a_3421_n88# a_4137_304# VDD.t297 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X601 a_13375_895# a_13216_993# a_13515_627# VSS.t241 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X602 a_1159_627# a_647_601# VSS.t46 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X603 VDD.t570 a_3807_895# a_3732_993# VDD.t569 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X604 VDD.t574 a_10509_601# a_10459_909# VDD.t573 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X605 a_10937_n62# a_11069_122# a_10801_n88# VSS.t180 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X606 a_3755_627# a_2585_627# a_3648_993# VSS.t409 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X607 a_12851_909# a_12433_993# a_12607_601# VDD.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X608 a_13193_n88# a_12447_n62# a_13329_n62# VSS.t337 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X609 a_4977_627# a_4811_627# VSS.t101 VSS.t100 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X610 a_6199_895# x2.X.t60 VDD.t147 VDD.t146 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X611 a_10125_993# a_9761_627# a_10041_993# VDD.t185 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X612 a_1028_212# x7.X VDD.t99 VDD.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X613 VDD.t7 a_3420_212# a_3421_n88# VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X614 VSS.t220 a_5323_2457# x9.A1.t5 VSS.t219 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X615 a_9646_90# a_9742_n88# VSS.t281 VSS.t280 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X616 VSS.t155 a_15767_895# a_16488_627# VSS.t154 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X617 VDD.t689 D[1].t2 a_16298_n62# VDD.t688 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X618 a_3947_627# x2.X.t61 VSS.t16 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X619 a_15380_212# x20.X VDD.t662 VDD.t661 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X620 a_11313_304# a_10801_n88# VDD.t560 VDD.t559 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X621 x2.X.t4 a_939_2457# VSS.t381 VSS.t380 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X622 a_12036_1467# x9.A1.t56 a_12178_1315# VSS.t35 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X623 a_2879_n62# x2.X.t62 VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X624 a_977_304# a_174_n88# VDD.t182 VDD.t181 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X625 x7.X a_1757_1642# VDD.t430 VDD.t429 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X626 VDD.t379 check[1].t4 a_13929_1642# VDD.t378 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X627 VSS.t677 a_10215_601# a_10149_627# VSS.t676 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X628 VSS.t426 VDD.t770 a_10937_n62# VSS.t425 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X629 VDD.t365 a_305_2457# x3.X VDD.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X630 VSS.t357 check[1].t5 a_13936_1315# VSS.t356 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X631 a_7254_90# a_7350_n88# VDD.t731 VDD.t730 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X632 a_12924_n62# a_12134_n88# VSS.t529 VSS.t528 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0703 ps=0.755 w=0.42 l=0.15
X633 VDD_SW_b[2].t0 a_13375_895# VSS.t254 VSS.t253 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X634 VDD.t676 a_8117_601# a_8848_909# VDD.t675 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X635 VDD.t509 VDD.t507 a_3625_n88# VDD.t508 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X636 VDD.t397 a_939_2457# x2.X.t21 VDD.t396 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X637 a_3369_304# a_2566_n88# VDD.t714 VDD.t713 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0956 ps=0.875 w=0.42 l=0.15
X638 a_10149_627# a_9595_627# a_10041_993# VSS.t309 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X639 a_10103_1642# x9.A1.t57 a_9644_1467# VDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X640 a_2585_627# a_2419_627# VDD.t157 VDD.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X641 VSS.t600 a_1415_895# a_2136_627# VSS.t599 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X642 VSS.t660 x30.A a_5323_2457# VSS.t659 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X643 VSS.t438 a_10073_1289# a_10007_1315# VSS.t437 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X644 VDD.t275 x10.X a_4811_627# VDD.t274 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X645 a_2949_993# a_2585_627# a_2865_993# VDD.t422 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X646 a_14825_993# a_14545_627# a_14733_627# VSS.t705 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X647 a_505_1289# check[6].t6 VDD.t483 VDD.t482 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X648 a_505_1289# check[6].t7 VSS.t492 VSS.t491 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X649 a_13632_909# a_13216_993# a_13375_895# VDD.t248 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X650 x9.A1.t17 a_5323_2457# VDD.t219 VDD.t218 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X651 x3.X a_305_2457# VSS.t339 VSS.t338 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X652 VDD.t451 a_2470_90# VSS_SW[6].t1 VDD.t450 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X653 a_5165_627# D[5].t3 VSS.t652 VSS.t651 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X654 VDD.t371 a_14999_601# a_14909_993# VDD.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X655 a_14526_n88# a_15072_106# a_15030_220# VDD.t312 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X656 x3.A a_29_2457# VDD.t558 VDD.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X657 VDD.t395 a_939_2457# x2.X.t20 VDD.t394 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X658 a_939_2457# x3.X VSS.t563 VSS.t562 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X659 a_13906_n62# a_12988_212# a_13461_122# VDD.t280 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X660 VDD.t1 x27.A a_4689_2457# VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X661 VSS.t218 a_5323_2457# x9.A1.t4 VSS.t217 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X662 a_10288_106# a_10596_212# a_10545_304# VDD.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X663 VSS.t296 a_10983_895# a_10931_627# VSS.t295 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X664 a_13461_122# a_12988_212# a_13705_n62# VSS.t268 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X665 VSS.t216 a_5323_2457# x9.A1.t3 VSS.t215 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X666 VDD.t645 a_1415_895# a_1340_993# VDD.t644 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X667 a_1363_627# a_193_627# a_1256_993# VSS.t413 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X668 a_2585_627# a_2419_627# VSS.t148 VSS.t147 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X669 a_12751_627# x2.X.t63 VSS.t18 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X670 a_3648_993# a_2419_627# a_3551_627# VSS.t146 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X671 a_13705_n62# a_13193_n88# VSS.t440 VSS.t439 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X672 VDD.t393 a_939_2457# x2.X.t19 VDD.t392 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X673 VSS.t265 x10.X a_4811_627# VSS.t264 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X674 a_7254_90# a_7350_n88# VSS.t698 VSS.t697 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X675 VSS.t214 a_5323_2457# x9.A1.t2 VSS.t213 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X676 a_1555_627# x2.X.t64 VSS.t34 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X677 a_12988_212# x17.X VDD.t174 VDD.t173 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X678 a_8342_304# a_8205_n88# a_7896_106# VDD.t198 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X679 a_8432_993# a_7369_627# a_8288_909# VDD.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X680 VDD.t26 a_15380_212# a_15381_n88# VDD.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X681 x11.X a_6539_1642# VSS.t613 VSS.t612 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X682 a_8933_1642# VSS.t467 a_8933_1315# VSS.t468 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X683 a_439_1315# VSS.t465 a_76_1467# VSS.t466 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X684 VDD.t674 a_8117_601# a_8067_909# VDD.t673 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X685 VDD.t133 check[3].t6 a_9147_1642# VDD.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X686 VDD_SW[4].t1 a_9312_627# VDD.t377 VDD.t376 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X687 VSS.t428 VDD.t771 a_1369_n62# VSS.t427 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0974 ps=0.97 w=0.42 l=0.15
X688 a_10359_627# a_10509_601# a_10215_601# VSS.t519 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X689 x30.A a_4689_2457# VSS.t711 VSS.t710 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X690 VSS.t126 check[3].t7 a_9154_1315# VSS.t125 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X691 a_1555_627# a_941_601# a_1415_895# VSS.t634 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X692 a_12607_601# a_12433_993# a_12751_627# VSS.t132 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X693 a_5323_2457# x30.A VDD.t693 VDD.t692 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X694 x2.X.t3 a_939_2457# VSS.t379 VSS.t378 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X695 a_13643_1642# a_13461_1642# VDD.t103 VDD.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X696 a_14839_n62# x2.X.t65 VDD.t34 VDD.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X697 VSS.t447 a_7252_1467# x12.X VSS.t446 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X698 VDD.t506 VDD.t504 a_15585_n88# VDD.t505 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X699 a_381_627# D[7].t2 VSS.t329 VSS.t328 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X700 a_1369_n62# a_1501_122# a_1233_n88# VSS.t490 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X701 a_12134_n88# a_12447_n62# a_12553_n62# VSS.t336 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X702 a_10007_1315# VSS.t463 a_9644_1467# VSS.t464 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X703 VDD.t578 x8.X a_2419_627# VDD.t577 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X704 a_10459_909# a_10041_993# a_10215_601# VDD.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X705 a_3625_n88# a_2879_n62# a_3761_n62# VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X706 a_14428_1467# VSS.t727 a_14570_1642# VDD.t466 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X707 a_12607_601# x2.X.t66 VDD.t36 VDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X708 a_2865_993# a_2419_627# a_2773_627# VDD.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X709 VDD.t60 a_1028_212# a_1029_n88# VDD.t59 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X710 VSS.t252 a_13375_895# a_14096_627# VSS.t251 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X711 a_14545_627# a_14379_627# VDD.t128 VDD.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X712 a_11240_909# a_10824_993# a_10983_895# VDD.t727 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X713 VDD.t624 a_14428_1467# x18.X VDD.t623 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X714 a_14570_1642# check[0].t6 VDD.t347 VDD.t346 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X715 a_1745_304# a_1233_n88# VDD.t338 VDD.t337 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X716 x9.A1.t16 a_5323_2457# VDD.t217 VDD.t216 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X717 a_14570_1315# check[0].t7 VSS.t327 VSS.t326 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X718 VDD.t641 a_6199_895# a_6920_627# VDD.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X719 a_11514_n62# a_10596_212# a_11069_122# VDD.t135 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X720 VSS.t445 a_4860_1467# x10.X VSS.t444 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X721 VDD.t197 a_14430_90# VSS_SW[1].t1 VDD.t196 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X722 a_939_2457# x3.X VSS.t561 VSS.t560 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X723 a_13461_122# a_12989_n88# a_13705_304# VDD.t208 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X724 x3.A a_29_2457# VSS.t508 VSS.t507 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X725 a_11325_1642# VSS.t461 a_11325_1315# VSS.t462 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X726 a_10727_627# a_10215_601# VSS.t675 VSS.t674 sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X727 a_10680_909# a_10215_601# VDD.t706 VDD.t705 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X728 VDD_SW_b[3].t0 a_10983_895# VSS.t294 VSS.t293 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X729 VDD.t391 a_939_2457# x2.X.t18 VDD.t390 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X730 VDD.t720 a_5725_601# a_6456_909# VDD.t719 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X731 VSS.t658 D[1].t3 a_16298_n62# VSS.t657 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X732 a_11313_n62# a_10801_n88# VSS.t512 VSS.t511 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X733 VSS.t522 x8.X a_2419_627# VSS.t521 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X734 x2.X.t2 a_939_2457# VSS.t377 VSS.t376 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X735 a_15608_993# a_14379_627# a_15511_627# VSS.t121 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X736 a_14545_627# a_14379_627# VSS.t120 VSS.t119 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X737 a_6040_993# a_4977_627# a_5896_909# VDD.t702 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X738 VSS.t212 a_5323_2457# x9.A1.t1 VSS.t211 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X739 a_4958_n88# a_5504_106# a_5462_220# VDD.t339 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X740 VDD_SW[5].t1 a_6920_627# VDD.t752 VDD.t751 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X741 a_10215_601# a_10041_993# a_10359_627# VSS.t141 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X742 a_4860_1467# VSS.t728 a_5002_1642# VDD.t465 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X743 a_1415_895# a_1256_993# a_1555_627# VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
X744 a_11069_122# a_10596_212# a_11313_n62# VSS.t128 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X745 a_8861_1642# a_8679_1642# VDD.t322 VDD.t321 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X746 VDD.t162 check[2].t6 a_11071_1642# VDD.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X747 a_5323_2457# x30.A VDD.t691 VDD.t690 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X748 x2.X.t1 a_939_2457# VSS.t375 VSS.t374 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X749 a_9742_n88# a_10055_n62# a_10161_n62# VSS.t94 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X750 VDD.t440 a_10073_1289# a_10103_1642# VDD.t439 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X751 VSS.t153 check[2].t7 a_11071_1642# VSS.t152 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X752 a_1233_n88# a_487_n62# a_1369_n62# VSS.t305 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X753 a_10359_627# x2.X.t67 VSS.t585 VSS.t584 sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X754 x3.X a_305_2457# VDD.t363 VDD.t362 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X755 a_1256_993# a_27_627# a_1159_627# VSS.t96 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X756 a_10215_601# x2.X.t68 VDD.t629 VDD.t628 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X757 VSS.t210 a_5323_2457# x9.A1.t0 VSS.t209 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X758 VDD.t176 a_78_90# VSS_SW[7].t1 VDD.t175 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X759 x27.A a_4413_2457# VDD.t95 VDD.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X760 a_15767_895# x2.X.t69 VDD.t631 VDD.t630 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X761 a_12153_627# a_11987_627# VDD.t582 VDD.t581 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X762 a_7967_627# a_8117_601# a_7823_601# VSS.t640 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X763 VDD.t69 D[6].t3 a_4338_n62# VDD.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X764 VDD.t419 x18.X a_14379_627# VDD.t418 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X765 VDD.t606 x3.X a_939_2457# VDD.t605 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X766 VSS.t430 VDD.t772 a_10161_n62# VSS.t429 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.109 ps=1.03 w=0.42 l=0.15
X767 a_78_90# a_174_n88# VDD.t180 VDD.t179 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X768 a_2468_1467# VSS.t729 a_2610_1642# VDD.t464 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X769 VDD.t279 a_12988_212# a_12989_n88# VDD.t278 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X770 VSS.t5 a_9646_90# VSS_SW[3].t0 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X771 a_7896_106# a_8204_212# a_8153_304# VDD.t651 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0787 ps=0.795 w=0.42 l=0.15
X772 VDD.t568 a_3807_895# a_4528_627# VDD.t567 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X773 VDD.t712 a_2566_n88# VSS_SW_b[6].t1 VDD.t711 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X774 VDD.t63 a_3625_n88# a_3558_304# VDD.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X775 VDD.t300 a_2468_1467# x8.X VDD.t299 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X776 a_2610_1642# check[5].t4 VDD.t687 VDD.t686 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X777 a_8067_909# a_7649_993# a_7823_601# VDD.t214 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X778 x2.X.t17 a_939_2457# VDD.t389 VDD.t388 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X779 a_2610_1315# check[5].t5 VSS.t656 VSS.t655 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X780 VDD.t304 a_10983_895# a_10908_993# VDD.t303 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X781 a_12447_n62# x2.X.t70 VDD.t595 VDD.t594 sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X782 VDD.t503 VDD.t501 a_13193_n88# VDD.t502 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X783 a_174_n88# a_720_106# a_678_220# VDD.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X784 VSS.t432 VDD.t773 a_12901_601# VSS.t431 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X785 a_2865_993# a_2585_627# a_2773_627# VSS.t408 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X786 a_12153_627# a_11987_627# VSS.t526 VSS.t525 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X787 a_7663_n62# x2.X.t71 VSS.t553 VSS.t552 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X788 a_9122_n62# a_8204_212# a_8677_122# VDD.t650 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X789 a_15692_993# a_14379_627# a_15608_993# VDD.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X790 VSS.t405 x18.X a_14379_627# VSS.t404 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X791 VDD.t487 check[5].t6 a_4363_1642# VDD.t486 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X792 VDD.t500 VDD.t498 a_12901_601# VDD.t499 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X793 VDD.t341 a_12036_1467# x16.X VDD.t340 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X794 a_12178_1642# check[1].t6 VDD.t125 VDD.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X795 a_9644_1467# x9.A1.t58 a_9786_1315# VSS.t127 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X796 VSS.t496 check[5].t7 a_4370_1315# VSS.t495 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X797 a_12178_1315# check[1].t7 VSS.t118 VSS.t117 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X798 a_2566_n88# a_3112_106# a_3070_220# VDD.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0882 ps=1.05 w=0.84 l=0.15
X799 VDD_SW_b[4].t0 a_8591_895# VSS.t573 VSS.t572 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X800 VDD.t744 a_4689_2457# x30.A VDD.t743 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X801 VDD.t497 VDD.t495 a_7350_n88# VDD.t496 sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.132 ps=1.22 w=0.42 l=0.15
X802 a_1946_n62# a_1028_212# a_1501_122# VDD.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X803 a_4363_1642# VSS.t730 a_4149_1642# VDD.t463 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X804 VDD.t271 a_12038_90# VSS_SW[2].t1 VDD.t270 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X805 a_1501_122# a_1028_212# a_1745_n62# VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.0671 ps=0.75 w=0.36 l=0.15
X806 a_78_90# a_174_n88# VSS.t171 VSS.t170 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X807 VDD.t211 x6.X a_27_627# VDD.t210 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X808 VDD_SW[3].t0 a_11704_627# VSS.t687 VSS.t686 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X809 x2.X.t0 a_939_2457# VSS.t373 VSS.t372 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X810 a_7711_1642# x9.A1.t59 a_7252_1467# VDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X811 a_1745_n62# a_1233_n88# VSS.t320 VSS.t319 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0882 ps=0.84 w=0.42 l=0.15
X812 VSS.t709 a_4689_2457# x30.A VSS.t708 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X813 x15.X a_11325_1642# VSS.t267 VSS.t266 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X814 VSS.t78 a_7681_1289# a_7615_1315# VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X815 a_13375_895# x2.X.t72 VDD.t597 VDD.t596 sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X816 VDD.t349 D[7].t3 a_1946_n62# VDD.t348 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X817 VDD.t178 a_505_1289# a_535_1642# VDD.t177 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X818 x13.X a_8933_1642# VDD.t24 VDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X819 a_13216_993# a_11987_627# a_13119_627# VSS.t524 sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X820 a_7823_601# a_7649_993# a_7967_627# VSS.t207 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X821 x27.A a_4413_2457# VSS.t84 VSS.t83 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X822 a_1971_1642# VSS.t731 a_1757_1642# VDD.t462 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X823 VDD_SW_b[5].t1 a_6199_895# VDD.t639 VDD.t638 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X824 VSS.t581 a_7254_90# VSS_SW[4].t0 VSS.t580 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X825 a_12433_993# a_11987_627# a_12341_627# VDD.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X826 a_7854_220# a_7663_n62# VDD.t434 VDD.t433 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X827 VDD.t426 check[4].t4 a_6285_1642# VDD.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X828 a_3625_n88# a_3893_122# a_3839_220# VDD.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X829 VSS.t412 check[4].t5 a_6285_1642# VSS.t411 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X830 VDD.t336 a_1233_n88# a_1166_304# VDD.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X831 a_8288_909# a_7823_601# VDD.t332 VDD.t331 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X832 a_13715_1642# VSS.t459 a_13715_1315# VSS.t460 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X833 VDD.t118 a_14526_n88# VSS_SW_b[1].t1 VDD.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X834 VDD.t164 a_15767_895# a_16488_627# VDD.t163 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X835 a_10055_n62# x2.X.t73 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.154 ps=1.34 w=0.64 l=0.15
X836 VSS.t204 x6.X a_27_627# VSS.t203 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X837 VSS.t510 a_10801_n88# a_10711_n62# VSS.t509 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.116 ps=1.09 w=0.64 l=0.15
X838 VDD.t152 a_15585_n88# a_15518_304# VDD.t151 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X839 VDD.t494 VDD.t492 a_10801_n88# VDD.t493 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X840 a_6231_220# a_5271_n62# VDD.t635 VDD.t634 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X841 a_5289_1289# check[4].t6 VDD.t680 VDD.t679 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X842 x2.X.t16 a_939_2457# VDD.t387 VDD.t386 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X843 a_5289_1289# check[4].t7 VSS.t645 VSS.t644 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
R0 VSS.n3198 VSS.n3196 51421.5
R1 VSS.n2902 VSS.n6 47892.9
R2 VSS.n2200 VSS.n2199 6286.08
R3 VSS VSS.n2893 5198.5
R4 VSS.n3196 VSS.n6 4543.55
R5 VSS.n3198 VSS.n3197 3810.55
R6 VSS VSS.n3198 2123.94
R7 VSS.n18 VSS.n14 1597.54
R8 VSS.n2893 VSS.n2892 1126.83
R9 VSS VSS.n717 1056
R10 VSS VSS.n557 1056
R11 VSS.n1514 VSS 1006.1
R12 VSS.n1628 VSS 1006.1
R13 VSS.n1742 VSS 1006.1
R14 VSS.n1856 VSS 1006.1
R15 VSS.n1970 VSS 1006.1
R16 VSS.n2084 VSS 1006.1
R17 VSS.n464 VSS 1001.85
R18 VSS.n357 VSS 1001.85
R19 VSS.n2199 VSS 898.782
R20 VSS.n2794 VSS 817.779
R21 VSS.n2695 VSS 817.779
R22 VSS.n2596 VSS 817.779
R23 VSS.n2497 VSS 817.779
R24 VSS.n2398 VSS 817.779
R25 VSS.n2299 VSS 817.779
R26 VSS.t578 VSS.n70 744.615
R27 VSS.t324 VSS.n137 744.615
R28 VSS.n549 VSS.t612 649.846
R29 VSS VSS.t404 643.903
R30 VSS VSS.t636 643.903
R31 VSS VSS.t632 643.903
R32 VSS VSS.t191 643.903
R33 VSS VSS.t264 643.903
R34 VSS VSS.t521 643.903
R35 VSS VSS.t203 643.903
R36 VSS.n1489 VSS.t705 603.659
R37 VSS.n1603 VSS.t696 603.659
R38 VSS.n1717 VSS.t177 603.659
R39 VSS.n1831 VSS.t85 603.659
R40 VSS.n1945 VSS.t671 603.659
R41 VSS.n2059 VSS.t408 603.659
R42 VSS.n2173 VSS.t414 603.659
R43 VSS.t444 VSS.n480 595.692
R44 VSS.n441 VSS.t484 595.692
R45 VSS.t289 VSS.n373 595.692
R46 VSS.n334 VSS.t482 595.692
R47 VSS.t40 VSS.n266 595.692
R48 VSS.n1404 VSS.t558 590.245
R49 VSS.n1497 VSS.t550 590.245
R50 VSS.t404 VSS.n1512 590.245
R51 VSS.n1518 VSS.t299 590.245
R52 VSS.n1611 VSS.t123 590.245
R53 VSS.t636 VSS.n1626 590.245
R54 VSS.n1632 VSS.t686 590.245
R55 VSS.n1725 VSS.t29 590.245
R56 VSS.t632 VSS.n1740 590.245
R57 VSS.n1746 VSS.t354 590.245
R58 VSS.n1839 VSS.t501 590.245
R59 VSS.t191 VSS.n1854 590.245
R60 VSS.n1860 VSS.t716 590.245
R61 VSS.n1953 VSS.t651 590.245
R62 VSS.t264 VSS.n1968 590.245
R63 VSS.n1974 VSS.t610 590.245
R64 VSS.n2067 VSS.t69 590.245
R65 VSS.t521 VSS.n2082 590.245
R66 VSS.n2088 VSS.t2 590.245
R67 VSS.n2181 VSS.t328 590.245
R68 VSS.n2190 VSS.t203 590.245
R69 VSS.n1277 VSS.t653 582.154
R70 VSS.n1067 VSS.t356 568.615
R71 VSS.n739 VSS.t464 568.615
R72 VSS.n579 VSS.t486 568.615
R73 VSS.n1410 VSS.t154 550
R74 VSS.n1524 VSS.t251 550
R75 VSS.n1638 VSS.t297 550
R76 VSS.n1752 VSS.t574 550
R77 VSS.n1866 VSS.t593 550
R78 VSS.n1980 VSS.t513 550
R79 VSS.n2094 VSS.t599 550
R80 VSS.n433 VSS.t638 541.538
R81 VSS.n326 VSS.t417 541.538
R82 VSS.n1512 VSS.t119 536.586
R83 VSS.n1626 VSS.t525 536.586
R84 VSS.n1740 VSS.t311 536.586
R85 VSS.n1854 VSS.t134 536.586
R86 VSS.n1968 VSS.t100 536.586
R87 VSS.n2082 VSS.t147 536.586
R88 VSS.n2190 VSS.t97 536.586
R89 VSS.n3041 VSS.n3038 533.059
R90 VSS.n3061 VSS.n3058 533.059
R91 VSS.n1263 VSS.t583 528
R92 VSS.n1100 VSS.t326 514.462
R93 VSS.n1053 VSS.t458 514.462
R94 VSS.n889 VSS.t117 514.462
R95 VSS.n745 VSS.t65 514.462
R96 VSS.n747 VSS.t437 514.462
R97 VSS.n585 VSS.t257 514.462
R98 VSS.n587 VSS.t77 514.462
R99 VSS.n481 VSS 514.462
R100 VSS.n374 VSS 514.462
R101 VSS.n267 VSS 514.462
R102 VSS.n1436 VSS.t679 509.757
R103 VSS.n1550 VSS.t241 509.757
R104 VSS.n1664 VSS.t694 509.757
R105 VSS.n1778 VSS.t116 509.757
R106 VSS.n1892 VSS.t286 509.757
R107 VSS.n2006 VSS.t673 509.757
R108 VSS.n2120 VSS.t14 509.757
R109 VSS.n1418 VSS.t156 496.341
R110 VSS.n1532 VSS.t253 496.341
R111 VSS.n1646 VSS.t293 496.341
R112 VSS.n1760 VSS.t572 496.341
R113 VSS.n1874 VSS.t595 496.341
R114 VSS.n1988 VSS.t517 496.341
R115 VSS.n2102 VSS.t601 496.341
R116 VSS.n23 VSS 487.385
R117 VSS.n436 VSS.t162 487.385
R118 VSS.n329 VSS.t63 487.385
R119 VSS.n89 VSS 473.846
R120 VSS.n2903 VSS.n2902 473.24
R121 VSS.n3196 VSS.n3195 473.24
R122 VSS.n911 VSS.t722 471.289
R123 VSS.n1122 VSS.t727 471.289
R124 VSS.n1240 VSS.t720 471.289
R125 VSS.n1030 VSS.t723 471.289
R126 VSS.n823 VSS.t718 471.289
R127 VSS.n731 VSS.t721 471.289
R128 VSS.n663 VSS.t725 471.289
R129 VSS.n571 VSS.t724 471.289
R130 VSS.n530 VSS.t719 471.289
R131 VSS.n494 VSS.t728 471.289
R132 VSS.n449 VSS.t730 471.289
R133 VSS.n387 VSS.t729 471.289
R134 VSS.n342 VSS.t731 471.289
R135 VSS.n280 VSS.t726 471.289
R136 VSS.n1114 VSS.t554 460.308
R137 VSS.n903 VSS.t35 460.308
R138 VSS.n1424 VSS.t421 456.099
R139 VSS.n1538 VSS.t431 456.099
R140 VSS.n1652 VSS.t616 456.099
R141 VSS.n1766 VSS.t622 456.099
R142 VSS.n1880 VSS.t542 456.099
R143 VSS.n1994 VSS.t546 456.099
R144 VSS.n2108 VSS.t624 456.099
R145 VSS.n1485 VSS.t122 429.269
R146 VSS.n1599 VSS.t527 429.269
R147 VSS.n1713 VSS.t309 429.269
R148 VSS.n1827 VSS.t136 429.269
R149 VSS.n1941 VSS.t103 429.269
R150 VSS.n2055 VSS.t149 429.269
R151 VSS.n2169 VSS.t99 429.269
R152 VSS.n3011 VSS 428.17
R153 VSS.n3040 VSS 428.17
R154 VSS VSS.n3087 428.17
R155 VSS VSS.n3059 428.17
R156 VSS.t266 VSS.n153 406.154
R157 VSS.t21 VSS.n195 406.154
R158 VSS.n1432 VSS.t49 402.44
R159 VSS.n1546 VSS.t704 402.44
R160 VSS.n1660 VSS.t520 402.44
R161 VSS.n1774 VSS.t641 402.44
R162 VSS.n1888 VSS.t688 402.44
R163 VSS.n2002 VSS.t313 402.44
R164 VSS.n2116 VSS.t634 402.44
R165 VSS.n2873 VSS.t436 400
R166 VSS.n2774 VSS.t202 400
R167 VSS.n2675 VSS.t648 400
R168 VSS.n2576 VSS.t189 400
R169 VSS.n2477 VSS.t140 400
R170 VSS.n2378 VSS.t288 400
R171 VSS.n2279 VSS.t43 400
R172 VSS.t630 VSS.n2895 391.111
R173 VSS.n1288 VSS.t657 391.111
R174 VSS.n1297 VSS.t187 391.111
R175 VSS.t164 VSS.n2792 391.111
R176 VSS.n1304 VSS.t272 391.111
R177 VSS.n1313 VSS.t261 391.111
R178 VSS.t81 VSS.n2693 391.111
R179 VSS.n1320 VSS.t27 391.111
R180 VSS.n1329 VSS.t4 391.111
R181 VSS.t406 VSS.n2594 391.111
R182 VSS.n1336 VSS.t499 391.111
R183 VSS.n1345 VSS.t580 391.111
R184 VSS.t278 VSS.n2495 391.111
R185 VSS.n1352 VSS.t649 391.111
R186 VSS.n1361 VSS.t181 391.111
R187 VSS.t10 VSS.n2396 391.111
R188 VSS.n1368 VSS.t67 391.111
R189 VSS.n1377 VSS.t448 391.111
R190 VSS.t87 VSS.n2297 391.111
R191 VSS.n1384 VSS.t274 391.111
R192 VSS.n1393 VSS.t166 391.111
R193 VSS VSS.n6 388.733
R194 VSS.n859 VSS.t497 379.077
R195 VSS.n699 VSS.t125 379.077
R196 VSS.n1481 VSS.t348 375.611
R197 VSS.n1595 VSS.t245 375.611
R198 VSS.n1709 VSS.t676 375.611
R199 VSS.n1823 VSS.t317 375.611
R200 VSS.n1937 VSS.t456 375.611
R201 VSS.n2051 VSS.t185 375.611
R202 VSS.n2165 VSS.t47 375.611
R203 VSS.n541 VSS.t642 365.538
R204 VSS.n486 VSS.t330 365.538
R205 VSS.n379 VSS.t655 365.538
R206 VSS.n272 VSS.t493 365.538
R207 VSS.n2799 VSS.t114 364.445
R208 VSS.n2700 VSS.t532 364.445
R209 VSS.n2601 VSS.t280 364.445
R210 VSS.n2502 VSS.t697 364.445
R211 VSS.n2403 VSS.t75 364.445
R212 VSS.n2304 VSS.t684 364.445
R213 VSS.n2205 VSS.t170 364.445
R214 VSS.n2895 VSS.t24 355.557
R215 VSS.n2792 VSS.t269 355.557
R216 VSS.n2693 VSS.t129 355.557
R217 VSS.n2594 VSS.t606 355.557
R218 VSS.n2495 VSS.t199 355.557
R219 VSS.n2396 VSS.t8 355.557
R220 VSS.n2297 VSS.t53 355.557
R221 VSS.n2820 VSS.t302 337.779
R222 VSS.n2721 VSS.t410 337.779
R223 VSS.n2622 VSS.t443 337.779
R224 VSS.n2523 VSS.t487 337.779
R225 VSS.n2424 VSS.t323 337.779
R226 VSS.n2325 VSS.t93 337.779
R227 VSS.n2226 VSS.t42 337.779
R228 VSS.n1292 VSS.t110 328.889
R229 VSS.n1308 VSS.t530 328.889
R230 VSS.n1324 VSS.t284 328.889
R231 VSS.n1340 VSS.t701 328.889
R232 VSS.n1356 VSS.t73 328.889
R233 VSS.n1372 VSS.t682 328.889
R234 VSS.n1388 VSS.t174 328.889
R235 VSS VSS.t205 324.923
R236 VSS VSS.t178 324.923
R237 VSS VSS.t266 324.923
R238 VSS.n846 VSS.t588 324.923
R239 VSS VSS.t21 324.923
R240 VSS.n686 VSS.t263 324.923
R241 VSS.t612 VSS 324.923
R242 VSS.n537 VSS.t242 311.385
R243 VSS.n490 VSS.t555 311.385
R244 VSS.n383 VSS.t587 311.385
R245 VSS.n276 VSS.t259 311.385
R246 VSS.n2808 VSS.t193 302.223
R247 VSS.n2709 VSS.t556 302.223
R248 VSS.n2610 VSS.t366 302.223
R249 VSS.n2511 VSS.t552 302.223
R250 VSS.n2412 VSS.t503 302.223
R251 VSS.n2313 VSS.t106 302.223
R252 VSS.n2214 VSS.t358 302.223
R253 VSS.n1442 VSS.t364 295.123
R254 VSS.n1454 VSS.t121 295.123
R255 VSS.n1556 VSS.t368 295.123
R256 VSS.n1568 VSS.t524 295.123
R257 VSS.n1670 VSS.t137 295.123
R258 VSS.n1682 VSS.t310 295.123
R259 VSS.n1784 VSS.t79 295.123
R260 VSS.n1796 VSS.t133 295.123
R261 VSS.n1898 VSS.t488 295.123
R262 VSS.n1910 VSS.t102 295.123
R263 VSS.n2012 VSS.t15 295.123
R264 VSS.n2024 VSS.t146 295.123
R265 VSS.n2126 VSS.t33 295.123
R266 VSS.n2138 VSS.t96 295.123
R267 VSS.n750 VSS.n746 294.007
R268 VSS.n590 VSS.n586 294.007
R269 VSS.n438 VSS.n437 294.007
R270 VSS.n331 VSS.n330 294.007
R271 VSS.n302 VSS.n301 292.5
R272 VSS.n301 VSS.n300 292.5
R273 VSS.n305 VSS.n304 292.5
R274 VSS.n304 VSS.n303 292.5
R275 VSS.n308 VSS.n307 292.5
R276 VSS.n307 VSS.n306 292.5
R277 VSS.n311 VSS.n310 292.5
R278 VSS.n310 VSS.n309 292.5
R279 VSS.n314 VSS.n313 292.5
R280 VSS.n313 VSS.n312 292.5
R281 VSS.n317 VSS.n316 292.5
R282 VSS.n316 VSS.n315 292.5
R283 VSS.n320 VSS.n319 292.5
R284 VSS.n319 VSS.n318 292.5
R285 VSS.n256 VSS.n255 292.5
R286 VSS.n255 VSS.n254 292.5
R287 VSS.n330 VSS.n329 292.5
R288 VSS.n328 VSS.n327 292.5
R289 VSS.n327 VSS.n326 292.5
R290 VSS.n336 VSS.n335 292.5
R291 VSS.n335 VSS.n334 292.5
R292 VSS.n341 VSS.n340 292.5
R293 VSS.n340 VSS.n339 292.5
R294 VSS.n349 VSS.n348 292.5
R295 VSS.n348 VSS.n347 292.5
R296 VSS.n359 VSS.n358 292.5
R297 VSS.n358 VSS.n357 292.5
R298 VSS.n355 VSS.n253 292.5
R299 VSS.n356 VSS.n355 292.5
R300 VSS.n367 VSS.n366 292.5
R301 VSS.n366 VSS.n365 292.5
R302 VSS.n370 VSS.n369 292.5
R303 VSS.n369 VSS.n368 292.5
R304 VSS.n409 VSS.n408 292.5
R305 VSS.n408 VSS.n407 292.5
R306 VSS.n412 VSS.n411 292.5
R307 VSS.n411 VSS.n410 292.5
R308 VSS.n415 VSS.n414 292.5
R309 VSS.n414 VSS.n413 292.5
R310 VSS.n418 VSS.n417 292.5
R311 VSS.n417 VSS.n416 292.5
R312 VSS.n421 VSS.n420 292.5
R313 VSS.n420 VSS.n419 292.5
R314 VSS.n424 VSS.n423 292.5
R315 VSS.n423 VSS.n422 292.5
R316 VSS.n427 VSS.n426 292.5
R317 VSS.n426 VSS.n425 292.5
R318 VSS.n245 VSS.n244 292.5
R319 VSS.n244 VSS.n243 292.5
R320 VSS.n437 VSS.n436 292.5
R321 VSS.n435 VSS.n434 292.5
R322 VSS.n434 VSS.n433 292.5
R323 VSS.n443 VSS.n442 292.5
R324 VSS.n442 VSS.n441 292.5
R325 VSS.n448 VSS.n447 292.5
R326 VSS.n447 VSS.n446 292.5
R327 VSS.n456 VSS.n455 292.5
R328 VSS.n455 VSS.n454 292.5
R329 VSS.n466 VSS.n465 292.5
R330 VSS.n465 VSS.n464 292.5
R331 VSS.n462 VSS.n242 292.5
R332 VSS.n463 VSS.n462 292.5
R333 VSS.n474 VSS.n473 292.5
R334 VSS.n473 VSS.n472 292.5
R335 VSS.n477 VSS.n476 292.5
R336 VSS.n476 VSS.n475 292.5
R337 VSS.n516 VSS.n515 292.5
R338 VSS.n515 VSS.n514 292.5
R339 VSS.n554 VSS.n553 292.5
R340 VSS.n553 VSS.n552 292.5
R341 VSS.n556 VSS.n555 292.5
R342 VSS.n557 VSS.n556 292.5
R343 VSS.n560 VSS.n559 292.5
R344 VSS.n559 VSS.n558 292.5
R345 VSS.n225 VSS.n224 292.5
R346 VSS.n224 VSS.n223 292.5
R347 VSS.n568 VSS.n567 292.5
R348 VSS.n567 VSS.n566 292.5
R349 VSS.n576 VSS.n575 292.5
R350 VSS.n575 VSS.n574 292.5
R351 VSS.n581 VSS.n580 292.5
R352 VSS.n580 VSS.n579 292.5
R353 VSS.n589 VSS.n588 292.5
R354 VSS.n588 VSS.n587 292.5
R355 VSS.n586 VSS.n585 292.5
R356 VSS.n220 VSS.n219 292.5
R357 VSS.n219 VSS.n218 292.5
R358 VSS.n599 VSS.n598 292.5
R359 VSS.n598 VSS.n597 292.5
R360 VSS.n602 VSS.n601 292.5
R361 VSS.n601 VSS.n600 292.5
R362 VSS.n605 VSS.n604 292.5
R363 VSS.n604 VSS.n603 292.5
R364 VSS.n608 VSS.n607 292.5
R365 VSS.n607 VSS.n606 292.5
R366 VSS.n611 VSS.n610 292.5
R367 VSS.n610 VSS.n609 292.5
R368 VSS.n614 VSS.n613 292.5
R369 VSS.n613 VSS.n612 292.5
R370 VSS.n617 VSS.n616 292.5
R371 VSS.n616 VSS.n615 292.5
R372 VSS.n714 VSS.n713 292.5
R373 VSS.n713 VSS.n712 292.5
R374 VSS.n716 VSS.n715 292.5
R375 VSS.n717 VSS.n716 292.5
R376 VSS.n720 VSS.n719 292.5
R377 VSS.n719 VSS.n718 292.5
R378 VSS.n183 VSS.n182 292.5
R379 VSS.n182 VSS.n181 292.5
R380 VSS.n728 VSS.n727 292.5
R381 VSS.n727 VSS.n726 292.5
R382 VSS.n736 VSS.n735 292.5
R383 VSS.n735 VSS.n734 292.5
R384 VSS.n741 VSS.n740 292.5
R385 VSS.n740 VSS.n739 292.5
R386 VSS.n749 VSS.n748 292.5
R387 VSS.n748 VSS.n747 292.5
R388 VSS.n746 VSS.n745 292.5
R389 VSS.n178 VSS.n177 292.5
R390 VSS.n177 VSS.n176 292.5
R391 VSS.n759 VSS.n758 292.5
R392 VSS.n758 VSS.n757 292.5
R393 VSS.n762 VSS.n761 292.5
R394 VSS.n761 VSS.n760 292.5
R395 VSS.n765 VSS.n764 292.5
R396 VSS.n764 VSS.n763 292.5
R397 VSS.n768 VSS.n767 292.5
R398 VSS.n767 VSS.n766 292.5
R399 VSS.n771 VSS.n770 292.5
R400 VSS.n770 VSS.n769 292.5
R401 VSS.n774 VSS.n773 292.5
R402 VSS.n773 VSS.n772 292.5
R403 VSS.n777 VSS.n776 292.5
R404 VSS.n776 VSS.n775 292.5
R405 VSS.n874 VSS.n873 292.5
R406 VSS.n873 VSS.n872 292.5
R407 VSS.n970 VSS.n969 292.5
R408 VSS.n969 VSS.n968 292.5
R409 VSS.n973 VSS.n972 292.5
R410 VSS.n972 VSS.n971 292.5
R411 VSS.n976 VSS.n975 292.5
R412 VSS.n975 VSS.n974 292.5
R413 VSS.n979 VSS.n978 292.5
R414 VSS.n978 VSS.n977 292.5
R415 VSS.n982 VSS.n981 292.5
R416 VSS.n981 VSS.n980 292.5
R417 VSS.n985 VSS.n984 292.5
R418 VSS.n984 VSS.n983 292.5
R419 VSS.n1082 VSS.n1081 292.5
R420 VSS.n1081 VSS.n1080 292.5
R421 VSS.n1085 VSS.n1084 292.5
R422 VSS.n1084 VSS.n1083 292.5
R423 VSS.n1181 VSS.n1180 292.5
R424 VSS.n1180 VSS.n1179 292.5
R425 VSS.n1184 VSS.n1183 292.5
R426 VSS.n1183 VSS.n1182 292.5
R427 VSS.n1187 VSS.n1186 292.5
R428 VSS.n1186 VSS.n1185 292.5
R429 VSS.n1190 VSS.n1189 292.5
R430 VSS.n1189 VSS.n1188 292.5
R431 VSS.n1193 VSS.n1192 292.5
R432 VSS.n1192 VSS.n1191 292.5
R433 VSS.n1196 VSS.n1195 292.5
R434 VSS.n1195 VSS.n1194 292.5
R435 VSS.n2869 VSS.t23 284.445
R436 VSS.n2770 VSS.t268 284.445
R437 VSS.n2671 VSS.t128 284.445
R438 VSS.n2572 VSS.t608 284.445
R439 VSS.n2473 VSS.t197 284.445
R440 VSS.n2374 VSS.t6 284.445
R441 VSS.n2275 VSS.t51 284.445
R442 VSS.n156 VSS 284.308
R443 VSS.n198 VSS 284.308
R444 VSS VSS.t630 275.557
R445 VSS VSS.t164 275.557
R446 VSS VSS.t81 275.557
R447 VSS VSS.t406 275.557
R448 VSS VSS.t278 275.557
R449 VSS VSS.t10 275.557
R450 VSS VSS.t87 275.557
R451 VSS VSS.n548 270.769
R452 VSS.n3040 VSS.t83 270.423
R453 VSS.n3060 VSS.t59 270.423
R454 VSS.n2816 VSS.t304 266.668
R455 VSS.n2717 VSS.t336 266.668
R456 VSS.n2618 VSS.t94 266.668
R457 VSS.n2519 VSS.t433 266.668
R458 VSS.n2420 VSS.t592 266.668
R459 VSS.n2321 VSS.t20 266.668
R460 VSS.n2222 VSS.t306 266.668
R461 VSS.n2865 VSS.t142 248.889
R462 VSS.n2766 VSS.t439 248.889
R463 VSS.n2667 VSS.t511 248.889
R464 VSS.n2568 VSS.t690 248.889
R465 VSS.n2469 VSS.t36 248.889
R466 VSS.n2370 VSS.t55 248.889
R467 VSS.n2271 VSS.t319 248.889
R468 VSS.n2954 VSS.t227 247.887
R469 VSS.n3003 VSS.t665 247.887
R470 VSS.n3030 VSS.t0 247.887
R471 VSS.n3044 VSS.t352 247.887
R472 VSS.n3143 VSS.t386 247.887
R473 VSS.n3092 VSS.t564 247.887
R474 VSS.n1 VSS.t507 247.887
R475 VSS.n1 VSS.t243 247.887
R476 VSS.n1217 VSS.t249 243.692
R477 VSS VSS.n463 243.692
R478 VSS VSS.n356 243.692
R479 VSS.n1006 VSS.t614 230.155
R480 VSS.n726 VSS.t127 230.155
R481 VSS.n566 VSS.t582 230.155
R482 VSS.n1446 VSS.t158 228.049
R483 VSS.n1560 VSS.t255 228.049
R484 VSS.n1674 VSS.t295 228.049
R485 VSS.n1788 VSS.t576 228.049
R486 VSS.n1902 VSS.t597 228.049
R487 VSS.n2016 VSS.t515 228.049
R488 VSS.n2130 VSS.t603 228.049
R489 VSS.n2954 VSS.t221 225.352
R490 VSS.n3003 VSS.t659 225.352
R491 VSS.n3030 VSS.t712 225.352
R492 VSS.n3143 VSS.t402 225.352
R493 VSS.n3092 VSS.t566 225.352
R494 VSS.n3064 VSS.t338 225.352
R495 VSS.n19 VSS.n18 216.615
R496 VSS.n23 VSS.n22 216.615
R497 VSS.n1277 VSS.n1276 216.615
R498 VSS.n1263 VSS.n1262 216.615
R499 VSS.n1248 VSS.n1247 216.615
R500 VSS.n1232 VSS.n1231 216.615
R501 VSS.n34 VSS.n33 216.615
R502 VSS.n1217 VSS.n1216 216.615
R503 VSS.n1203 VSS.n1202 216.615
R504 VSS.t178 VSS.n86 216.615
R505 VSS.n153 VSS.n152 216.615
R506 VSS.n155 VSS.n154 216.615
R507 VSS.n858 VSS.n857 216.615
R508 VSS.n845 VSS.n844 216.615
R509 VSS.n169 VSS.n168 216.615
R510 VSS.n797 VSS.n796 216.615
R511 VSS.n783 VSS.n782 216.615
R512 VSS.n195 VSS.n194 216.615
R513 VSS.n197 VSS.n196 216.615
R514 VSS.n698 VSS.n697 216.615
R515 VSS.n685 VSS.n684 216.615
R516 VSS.n211 VSS.n210 216.615
R517 VSS.n637 VSS.n636 216.615
R518 VSS.n623 VSS.n622 216.615
R519 VSS.t205 VSS.n20 203.077
R520 VSS.n85 VSS.n84 203.077
R521 VSS.n89 VSS.n88 203.077
R522 VSS.n1067 VSS.n1066 203.077
R523 VSS.n1053 VSS.n1052 203.077
R524 VSS.n1038 VSS.n1037 203.077
R525 VSS.n1022 VSS.n1021 203.077
R526 VSS.n101 VSS.n100 203.077
R527 VSS.n1006 VSS.n1005 203.077
R528 VSS.n992 VSS.n991 203.077
R529 VSS.n454 VSS.t586 203.077
R530 VSS.n347 VSS.t260 203.077
R531 VSS.n2948 VSS.t211 202.817
R532 VSS.n3147 VSS.t388 202.817
R533 VSS.n2838 VSS.t26 195.556
R534 VSS.n2826 VSS.t628 195.556
R535 VSS.n2739 VSS.t271 195.556
R536 VSS.n2727 VSS.t419 195.556
R537 VSS.n2640 VSS.t131 195.556
R538 VSS.n2628 VSS.t429 195.556
R539 VSS.n2541 VSS.t605 195.556
R540 VSS.n2529 VSS.t618 195.556
R541 VSS.n2442 VSS.t198 195.556
R542 VSS.n2430 VSS.t536 195.556
R543 VSS.n2343 VSS.t7 195.556
R544 VSS.n2331 VSS.t540 195.556
R545 VSS.n2244 VSS.t52 195.556
R546 VSS.n2232 VSS.t538 195.556
R547 VSS.n3187 VSS.t391 190.065
R548 VSS.n2907 VSS.t210 190.065
R549 VSS.n526 VSS.t505 189.538
R550 VSS.n501 VSS.t534 189.538
R551 VSS.n394 VSS.t150 189.538
R552 VSS.n287 VSS.t168 189.538
R553 VSS.n2846 VSS.t145 189.362
R554 VSS.n2747 VSS.t442 189.362
R555 VSS.n2648 VSS.t510 189.362
R556 VSS.n2549 VSS.t693 189.362
R557 VSS.n2450 VSS.t39 189.362
R558 VSS.n2351 VSS.t58 189.362
R559 VSS.n2252 VSS.t322 189.362
R560 VSS.n1462 VSS.t347 189.362
R561 VSS.n1576 VSS.t248 189.362
R562 VSS.n1690 VSS.t675 189.362
R563 VSS.n1804 VSS.t316 189.362
R564 VSS.n1918 VSS.t455 189.362
R565 VSS.n2032 VSS.t184 189.362
R566 VSS.n2146 VSS.t46 189.362
R567 VSS.n1450 VSS.t706 187.805
R568 VSS.n1564 VSS.t695 187.805
R569 VSS.n1678 VSS.t176 187.805
R570 VSS.n1792 VSS.t86 187.805
R571 VSS.n1906 VSS.t672 187.805
R572 VSS.n2020 VSS.t409 187.805
R573 VSS.n2134 VSS.t413 187.805
R574 VSS.n2958 VSS.t225 180.282
R575 VSS.n2999 VSS.t667 180.282
R576 VSS.n3026 VSS.t708 180.282
R577 VSS.n3137 VSS.t384 180.282
R578 VSS.n3098 VSS.t560 180.282
R579 VSS.n3070 VSS.t344 180.282
R580 VSS.n1160 VSS.t12 176
R581 VSS.n949 VSS.t350 176
R582 VSS.n181 VSS.t362 176
R583 VSS.n223 VSS.t589 176
R584 VSS.n814 VSS.t291 162.463
R585 VSS.n654 VSS.t307 162.463
R586 VSS.n2908 VSS.t209 157.746
R587 VSS.n2942 VSS.t231 157.746
R588 VSS.n3188 VSS.t390 157.746
R589 VSS.n3151 VSS.t372 157.746
R590 VSS.n519 VSS.n516 155.916
R591 VSS.n2830 VSS.t112 151.112
R592 VSS.n2731 VSS.t528 151.112
R593 VSS.n2632 VSS.t282 151.112
R594 VSS.n2533 VSS.t699 151.112
R595 VSS.n2434 VSS.t71 151.112
R596 VSS.n2335 VSS.t680 151.112
R597 VSS.n2236 VSS.t172 151.112
R598 VSS.n1174 VSS.n1173 148.923
R599 VSS.n1160 VSS.n1159 148.923
R600 VSS.n49 VSS.n48 148.923
R601 VSS.n1130 VSS.n1129 148.923
R602 VSS.n1114 VSS.n1113 148.923
R603 VSS.n1100 VSS.n1099 148.923
R604 VSS.n70 VSS.n64 148.923
R605 VSS.n73 VSS.n72 148.923
R606 VSS.n963 VSS.n962 148.923
R607 VSS.n949 VSS.n948 148.923
R608 VSS.n116 VSS.n115 148.923
R609 VSS.n919 VSS.n918 148.923
R610 VSS.n903 VSS.n902 148.923
R611 VSS.n889 VSS.n888 148.923
R612 VSS.n137 VSS.n131 148.923
R613 VSS.n140 VSS.n139 148.923
R614 VSS.n464 VSS.t495 148.923
R615 VSS.n357 VSS.t160 148.923
R616 VSS.n911 VSS.t469 148.35
R617 VSS.n1122 VSS.t473 148.35
R618 VSS.n1240 VSS.t475 148.35
R619 VSS.n1030 VSS.t459 148.35
R620 VSS.n823 VSS.t461 148.35
R621 VSS.n731 VSS.t463 148.35
R622 VSS.n663 VSS.t467 148.35
R623 VSS.n571 VSS.t485 148.35
R624 VSS.n530 VSS.t477 148.35
R625 VSS.n494 VSS.t471 148.35
R626 VSS.n449 VSS.t483 148.35
R627 VSS.n387 VSS.t479 148.35
R628 VSS.n342 VSS.t481 148.35
R629 VSS.n280 VSS.t465 148.35
R630 VSS.n1291 VSS.t658 145.006
R631 VSS.n1307 VSS.t273 145.006
R632 VSS.n1323 VSS.t28 145.006
R633 VSS.n1339 VSS.t500 145.006
R634 VSS.n1355 VSS.t650 145.006
R635 VSS.n1371 VSS.t68 145.006
R636 VSS.n1387 VSS.t275 145.006
R637 VSS.n1500 VSS.t551 145.006
R638 VSS.n1614 VSS.t124 145.006
R639 VSS.n1728 VSS.t30 145.006
R640 VSS.n1842 VSS.t502 145.006
R641 VSS.n1956 VSS.t652 145.006
R642 VSS.n2070 VSS.t70 145.006
R643 VSS.n2184 VSS.t329 145.006
R644 VSS VSS.t578 135.386
R645 VSS.n71 VSS 135.386
R646 VSS VSS.t324 135.386
R647 VSS.n138 VSS 135.386
R648 VSS.t276 VSS 135.386
R649 VSS.t446 VSS 135.386
R650 VSS.n533 VSS.t478 135.386
R651 VSS.n497 VSS.t472 135.386
R652 VSS VSS.t444 135.386
R653 VSS.n390 VSS.t480 135.386
R654 VSS VSS.t289 135.386
R655 VSS.n283 VSS.t466 135.386
R656 VSS VSS.t40 135.386
R657 VSS.n2964 VSS.t215 135.212
R658 VSS.n2993 VSS.t661 135.212
R659 VSS.n3020 VSS.t710 135.212
R660 VSS.n3133 VSS.t398 135.212
R661 VSS.n3102 VSS.t568 135.212
R662 VSS.n3074 VSS.t340 135.212
R663 VSS.n1467 VSS.t50 134.147
R664 VSS.n1581 VSS.t703 134.147
R665 VSS.n1695 VSS.t519 134.147
R666 VSS.n1809 VSS.t640 134.147
R667 VSS.n1923 VSS.t689 134.147
R668 VSS.n2037 VSS.t314 134.147
R669 VSS.n2151 VSS.t635 134.147
R670 VSS.n2834 VSS.t435 124.445
R671 VSS.n2735 VSS.t201 124.445
R672 VSS.n2636 VSS.t647 124.445
R673 VSS.n2537 VSS.t190 124.445
R674 VSS.n2438 VSS.t139 124.445
R675 VSS.n2339 VSS.t287 124.445
R676 VSS.n2240 VSS.t44 124.445
R677 VSS.n3178 VSS.n3177 116.219
R678 VSS.n3168 VSS.n3167 116.219
R679 VSS.n3164 VSS.n3163 116.219
R680 VSS.n3154 VSS.n3153 116.219
R681 VSS.n3142 VSS.n3141 116.219
R682 VSS.n3132 VSS.n3131 116.219
R683 VSS.n3122 VSS.n3121 116.219
R684 VSS.n3117 VSS.n3116 116.219
R685 VSS.n3107 VSS.n3106 116.219
R686 VSS.n3097 VSS.n3096 116.219
R687 VSS.n2917 VSS.n2916 116.219
R688 VSS.n2925 VSS.n2924 116.219
R689 VSS.n2935 VSS.n2934 116.219
R690 VSS.n2945 VSS.n2944 116.219
R691 VSS.n2953 VSS.n2952 116.219
R692 VSS.n2963 VSS.n2962 116.219
R693 VSS.n2973 VSS.n2972 116.219
R694 VSS.n2979 VSS.n2978 116.219
R695 VSS.n2988 VSS.n2987 116.219
R696 VSS.n2998 VSS.n2997 116.219
R697 VSS.n3054 VSS.t565 114.775
R698 VSS.n7 VSS.t666 114.775
R699 VSS.n2864 VSS.n2863 113.207
R700 VSS.n2765 VSS.n2764 113.207
R701 VSS.n2666 VSS.n2665 113.207
R702 VSS.n2567 VSS.n2566 113.207
R703 VSS.n2468 VSS.n2467 113.207
R704 VSS.n2369 VSS.n2368 113.207
R705 VSS.n2270 VSS.n2269 113.207
R706 VSS.n1480 VSS.n1479 113.207
R707 VSS.n1594 VSS.n1593 113.207
R708 VSS.n1708 VSS.n1707 113.207
R709 VSS.n1822 VSS.n1821 113.207
R710 VSS.n1936 VSS.n1935 113.207
R711 VSS.n2050 VSS.n2049 113.207
R712 VSS.n2164 VSS.n2163 113.207
R713 VSS.n2912 VSS.t229 112.677
R714 VSS.n2938 VSS.t213 112.677
R715 VSS.n3183 VSS.t380 112.677
R716 VSS.n3157 VSS.t392 112.677
R717 VSS.n3067 VSS.n3066 109.3
R718 VSS.n3033 VSS.n3032 109.3
R719 VSS.n1301 VSS.n1300 109.231
R720 VSS.n1317 VSS.n1316 109.231
R721 VSS.n1333 VSS.n1332 109.231
R722 VSS.n1349 VSS.n1348 109.231
R723 VSS.n1365 VSS.n1364 109.231
R724 VSS.n1381 VSS.n1380 109.231
R725 VSS.n1397 VSS.n1396 109.231
R726 VSS.n1522 VSS.n1521 109.231
R727 VSS.n1636 VSS.n1635 109.231
R728 VSS.n1750 VSS.n1749 109.231
R729 VSS.n1864 VSS.n1863 109.231
R730 VSS.n1978 VSS.n1977 109.231
R731 VSS.n2092 VSS.n2091 109.231
R732 VSS.n1408 VSS.n1407 109.231
R733 VSS.n2825 VSS.n2824 109.043
R734 VSS.n2726 VSS.n2725 109.043
R735 VSS.n2627 VSS.n2626 109.043
R736 VSS.n2528 VSS.n2527 109.043
R737 VSS.n2429 VSS.n2428 109.043
R738 VSS.n2330 VSS.n2329 109.043
R739 VSS.n2231 VSS.n2230 109.043
R740 VSS.n1441 VSS.n1440 109.043
R741 VSS.n1555 VSS.n1554 109.043
R742 VSS.n1669 VSS.n1668 109.043
R743 VSS.n1783 VSS.n1782 109.043
R744 VSS.n1897 VSS.n1896 109.043
R745 VSS.n2011 VSS.n2010 109.043
R746 VSS.n2125 VSS.n2124 109.043
R747 VSS.n1296 VSS.n1295 108.689
R748 VSS.n1312 VSS.n1311 108.689
R749 VSS.n1328 VSS.n1327 108.689
R750 VSS.n1344 VSS.n1343 108.689
R751 VSS.n1360 VSS.n1359 108.689
R752 VSS.n1376 VSS.n1375 108.689
R753 VSS.n1392 VSS.n1391 108.689
R754 VSS.n1422 VSS.n1421 108.689
R755 VSS.n1536 VSS.n1535 108.689
R756 VSS.n1650 VSS.n1649 108.689
R757 VSS.n1764 VSS.n1763 108.689
R758 VSS.n1878 VSS.n1877 108.689
R759 VSS.n1992 VSS.n1991 108.689
R760 VSS.n2106 VSS.n2105 108.689
R761 VSS.t332 VSS.n1143 108.308
R762 VSS.t452 VSS.n932 108.308
R763 VSS.n831 VSS.t462 108.308
R764 VSS.t462 VSS.n830 108.308
R765 VSS.n671 VSS.t468 108.308
R766 VSS.t468 VSS.n670 108.308
R767 VSS.n3078 VSS.n3077 108.254
R768 VSS.n3024 VSS.n3023 108.254
R769 VSS.n4 VSS.n0 107.478
R770 VSS.n2789 VSS.n2788 107.478
R771 VSS.n2690 VSS.n2689 107.478
R772 VSS.n2591 VSS.n2590 107.478
R773 VSS.n2492 VSS.n2491 107.478
R774 VSS.n2393 VSS.n2392 107.478
R775 VSS.n2294 VSS.n2293 107.478
R776 VSS.n2888 VSS.n2887 107.478
R777 VSS.n1509 VSS.n1508 107.478
R778 VSS.n1623 VSS.n1622 107.478
R779 VSS.n1737 VSS.n1736 107.478
R780 VSS.n1851 VSS.n1850 107.478
R781 VSS.n1965 VSS.n1964 107.478
R782 VSS.n2079 VSS.n2078 107.478
R783 VSS.n2194 VSS.n2193 107.478
R784 VSS.n229 VSS.n228 107.478
R785 VSS.n241 VSS.n240 107.478
R786 VSS.n252 VSS.n251 107.478
R787 VSS.n263 VSS.n262 107.478
R788 VSS.n3048 VSS.n3047 107.478
R789 VSS.n722 VSS.n180 107.24
R790 VSS.n562 VSS.n222 107.24
R791 VSS.n468 VSS.n461 107.24
R792 VSS.n361 VSS.n354 107.24
R793 VSS.n57 VSS.n56 106.731
R794 VSS.n96 VSS.n78 106.731
R795 VSS.n124 VSS.n123 106.731
R796 VSS.n163 VSS.n145 106.731
R797 VSS.n205 VSS.n187 106.731
R798 VSS.n28 VSS.n9 106.731
R799 VSS.n3055 VSS.t343 105.835
R800 VSS.n3016 VSS.t715 105.835
R801 VSS.n29 VSS.t451 93.2783
R802 VSS.n97 VSS.t92 93.2783
R803 VSS.n164 VSS.t292 93.2783
R804 VSS.n206 VSS.t308 93.2783
R805 VSS.n233 VSS.t506 93.2783
R806 VSS.n432 VSS.t639 93.2783
R807 VSS.n325 VSS.t418 93.2783
R808 VSS.n46 VSS.t333 93.2779
R809 VSS.n113 VSS.t453 93.2779
R810 VSS.n744 VSS.t438 93.2779
R811 VSS.n584 VSS.t78 93.2779
R812 VSS.n238 VSS.t535 93.2779
R813 VSS.n249 VSS.t151 93.2779
R814 VSS.n260 VSS.t169 93.2779
R815 VSS.n149 VSS.n148 92.7064
R816 VSS.n159 VSS.n158 92.7064
R817 VSS.n856 VSS.n855 92.7064
R818 VSS.n843 VSS.n842 92.7064
R819 VSS.n829 VSS.n828 92.7064
R820 VSS.n812 VSS.n811 92.7064
R821 VSS.n795 VSS.n794 92.7064
R822 VSS.n781 VSS.n780 92.7064
R823 VSS.n191 VSS.n190 92.7064
R824 VSS.n201 VSS.n200 92.7064
R825 VSS.n696 VSS.n695 92.7064
R826 VSS.n683 VSS.n682 92.7064
R827 VSS.n669 VSS.n668 92.7064
R828 VSS.n652 VSS.n651 92.7064
R829 VSS.n635 VSS.n634 92.7064
R830 VSS.n621 VSS.n620 92.7064
R831 VSS.n17 VSS.n16 92.7064
R832 VSS.n24 VSS.n13 92.7064
R833 VSS.n1278 VSS.n1274 92.7064
R834 VSS.n1264 VSS.n1260 92.7064
R835 VSS.n1249 VSS.n1245 92.7064
R836 VSS.n1233 VSS.n1229 92.7064
R837 VSS.n1218 VSS.n1214 92.7064
R838 VSS.n1204 VSS.n1200 92.7064
R839 VSS.n2968 VSS.t237 90.1413
R840 VSS.n2989 VSS.t669 90.1413
R841 VSS VSS.n3010 90.1413
R842 VSS.n3013 VSS.t714 90.1413
R843 VSS VSS.n3039 90.1413
R844 VSS.n3127 VSS.t376 90.1413
R845 VSS.n3108 VSS.t562 90.1413
R846 VSS.n3088 VSS 90.1413
R847 VSS.n3080 VSS.t342 90.1413
R848 VSS.n3060 VSS 90.1413
R849 VSS.n2851 VSS.t303 88.8894
R850 VSS.n2752 VSS.t337 88.8894
R851 VSS.n2653 VSS.t95 88.8894
R852 VSS.n2554 VSS.t434 88.8894
R853 VSS.n2455 VSS.t591 88.8894
R854 VSS.n2356 VSS.t19 88.8894
R855 VSS.n2257 VSS.t305 88.8894
R856 VSS.n83 VSS.n82 86.9123
R857 VSS.n1068 VSS.n1064 86.9123
R858 VSS.n1054 VSS.n1050 86.9123
R859 VSS.n1039 VSS.n1035 86.9123
R860 VSS.n1023 VSS.n1019 86.9123
R861 VSS.n1007 VSS.n1003 86.9123
R862 VSS.n993 VSS.n989 86.9123
R863 VSS.n3050 VSS 84.5075
R864 VSS.n3199 VSS 84.5075
R865 VSS.n2863 VSS.t143 81.4291
R866 VSS.n2764 VSS.t440 81.4291
R867 VSS.n2665 VSS.t512 81.4291
R868 VSS.n2566 VSS.t691 81.4291
R869 VSS.n2467 VSS.t37 81.4291
R870 VSS.n2368 VSS.t56 81.4291
R871 VSS.n2269 VSS.t320 81.4291
R872 VSS.n1479 VSS.t349 81.4291
R873 VSS.n1593 VSS.t246 81.4291
R874 VSS.n1707 VSS.t677 81.4291
R875 VSS.n1821 VSS.t318 81.4291
R876 VSS.n1935 VSS.t457 81.4291
R877 VSS.n2049 VSS.t186 81.4291
R878 VSS.n2163 VSS.t48 81.4291
R879 VSS.n1248 VSS.t476 81.2313
R880 VSS.n1173 VSS.n1172 81.2313
R881 VSS.n1159 VSS.n1158 81.2313
R882 VSS.n48 VSS.n47 81.2313
R883 VSS.n1143 VSS.n1142 81.2313
R884 VSS.n1129 VSS.n1128 81.2313
R885 VSS.n1113 VSS.n1112 81.2313
R886 VSS.n1099 VSS.n1098 81.2313
R887 VSS.n64 VSS.n63 81.2313
R888 VSS.n72 VSS.n71 81.2313
R889 VSS.n962 VSS.n961 81.2313
R890 VSS.n948 VSS.n947 81.2313
R891 VSS.n115 VSS.n114 81.2313
R892 VSS.n932 VSS.n931 81.2313
R893 VSS.n918 VSS.n917 81.2313
R894 VSS.n902 VSS.n901 81.2313
R895 VSS.n888 VSS.n887 81.2313
R896 VSS.n131 VSS.n130 81.2313
R897 VSS.n139 VSS.n138 81.2313
R898 VSS.n463 VSS.t89 81.2313
R899 VSS.n356 VSS.t415 81.2313
R900 VSS.n1458 VSS.t346 80.4883
R901 VSS.n1475 VSS.t195 80.4883
R902 VSS.n1572 VSS.t247 80.4883
R903 VSS.n1589 VSS.t17 80.4883
R904 VSS.n1686 VSS.t674 80.4883
R905 VSS.n1703 VSS.t584 80.4883
R906 VSS.n1800 VSS.t315 80.4883
R907 VSS.n1817 VSS.t360 80.4883
R908 VSS.n1914 VSS.t454 80.4883
R909 VSS.n1931 VSS.t31 80.4883
R910 VSS.n2028 VSS.t183 80.4883
R911 VSS.n2045 VSS.t108 80.4883
R912 VSS.n2142 VSS.t45 80.4883
R913 VSS.n2159 VSS.t104 80.4883
R914 VSS.n912 VSS.n911 76.0005
R915 VSS.n1123 VSS.n1122 76.0005
R916 VSS.n1241 VSS.n1240 76.0005
R917 VSS.n1031 VSS.n1030 76.0005
R918 VSS.n824 VSS.n823 76.0005
R919 VSS.n732 VSS.n731 76.0005
R920 VSS.n664 VSS.n663 76.0005
R921 VSS.n572 VSS.n571 76.0005
R922 VSS.n531 VSS.n530 76.0005
R923 VSS.n495 VSS.n494 76.0005
R924 VSS.n450 VSS.n449 76.0005
R925 VSS.n388 VSS.n387 76.0005
R926 VSS.n343 VSS.n342 76.0005
R927 VSS.n281 VSS.n280 76.0005
R928 VSS.n9 VSS.t654 74.2862
R929 VSS.n56 VSS.t327 74.2862
R930 VSS.n78 VSS.t357 74.2862
R931 VSS.n123 VSS.t118 74.2862
R932 VSS.n145 VSS.t498 74.2862
R933 VSS.n180 VSS.t363 74.2862
R934 VSS.n187 VSS.t126 74.2862
R935 VSS.n222 VSS.t590 74.2862
R936 VSS.n228 VSS.t643 74.2862
R937 VSS.n240 VSS.t331 74.2862
R938 VSS.n461 VSS.t496 74.2862
R939 VSS.n251 VSS.t656 74.2862
R940 VSS.n354 VSS.t161 74.2862
R941 VSS.n262 VSS.t494 74.2862
R942 VSS.n46 VSS.t13 70.4212
R943 VSS.n113 VSS.t351 70.4212
R944 VSS.n744 VSS.t66 70.4212
R945 VSS.n584 VSS.t258 70.4212
R946 VSS.n238 VSS.t645 70.4212
R947 VSS.n249 VSS.t335 70.4212
R948 VSS.n260 VSS.t492 70.4212
R949 VSS.n29 VSS.t250 70.4207
R950 VSS.n97 VSS.t615 70.4207
R951 VSS.n164 VSS.t153 70.4207
R952 VSS.n206 VSS.t371 70.4207
R953 VSS.n233 VSS.t412 70.4207
R954 VSS.n432 VSS.t163 70.4207
R955 VSS.n325 VSS.t64 70.4207
R956 VSS.n38 VSS.n37 68.8369
R957 VSS.n1038 VSS.t460 67.6928
R958 VSS.n2918 VSS.t223 67.6061
R959 VSS.n2932 VSS.t235 67.6061
R960 VSS.n3179 VSS.t400 67.6061
R961 VSS.n3161 VSS.t374 67.6061
R962 VSS.n93 VSS.n92 65.5421
R963 VSS.n105 VSS.n104 65.4925
R964 VSS.n1175 VSS.n1171 63.7358
R965 VSS.n1161 VSS.n1157 63.7358
R966 VSS.n1145 VSS.n1141 63.7358
R967 VSS.n1131 VSS.n1127 63.7358
R968 VSS.n1115 VSS.n1111 63.7358
R969 VSS.n1101 VSS.n1097 63.7358
R970 VSS.n69 VSS.n67 63.7358
R971 VSS.n74 VSS.n62 63.7358
R972 VSS.n964 VSS.n960 63.7358
R973 VSS.n950 VSS.n946 63.7358
R974 VSS.n934 VSS.n930 63.7358
R975 VSS.n920 VSS.n916 63.7358
R976 VSS.n904 VSS.n900 63.7358
R977 VSS.n890 VSS.n886 63.7358
R978 VSS.n136 VSS.n134 63.7358
R979 VSS.n141 VSS.n129 63.7358
R980 VSS.n2824 VSS.t113 57.1434
R981 VSS.n2725 VSS.t529 57.1434
R982 VSS.n2626 VSS.t283 57.1434
R983 VSS.n2527 VSS.t700 57.1434
R984 VSS.n2428 VSS.t72 57.1434
R985 VSS.n2329 VSS.t681 57.1434
R986 VSS.n2230 VSS.t173 57.1434
R987 VSS.n1440 VSS.t159 57.1434
R988 VSS.n1554 VSS.t256 57.1434
R989 VSS.n1668 VSS.t296 57.1434
R990 VSS.n1782 VSS.t577 57.1434
R991 VSS.n1896 VSS.t598 57.1434
R992 VSS.n2010 VSS.t516 57.1434
R993 VSS.n2124 VSS.t604 57.1434
R994 VSS.n166 VSS.n165 55.8038
R995 VSS.n208 VSS.n207 55.8038
R996 VSS.n1295 VSS.t194 54.2862
R997 VSS.n1300 VSS.t115 54.2862
R998 VSS.n1311 VSS.t557 54.2862
R999 VSS.n1316 VSS.t533 54.2862
R1000 VSS.n1327 VSS.t367 54.2862
R1001 VSS.n1332 VSS.t281 54.2862
R1002 VSS.n1343 VSS.t553 54.2862
R1003 VSS.n1348 VSS.t698 54.2862
R1004 VSS.n1359 VSS.t504 54.2862
R1005 VSS.n1364 VSS.t76 54.2862
R1006 VSS.n1375 VSS.t107 54.2862
R1007 VSS.n1380 VSS.t685 54.2862
R1008 VSS.n1391 VSS.t359 54.2862
R1009 VSS.n1396 VSS.t171 54.2862
R1010 VSS.n1407 VSS.t155 54.2862
R1011 VSS.n1421 VSS.t422 54.2862
R1012 VSS.n1521 VSS.t252 54.2862
R1013 VSS.n1535 VSS.t432 54.2862
R1014 VSS.n1635 VSS.t298 54.2862
R1015 VSS.n1649 VSS.t617 54.2862
R1016 VSS.n1749 VSS.t575 54.2862
R1017 VSS.n1763 VSS.t623 54.2862
R1018 VSS.n1863 VSS.t594 54.2862
R1019 VSS.n1877 VSS.t543 54.2862
R1020 VSS.n1977 VSS.t514 54.2862
R1021 VSS.n1991 VSS.t547 54.2862
R1022 VSS.n2091 VSS.t600 54.2862
R1023 VSS.n2105 VSS.t625 54.2862
R1024 VSS.t291 VSS.n813 54.1543
R1025 VSS.n718 VSS.t276 54.1543
R1026 VSS.t307 VSS.n653 54.1543
R1027 VSS.n558 VSS.t446 54.1543
R1028 VSS.n2859 VSS.t548 53.3338
R1029 VSS.n2842 VSS.t144 53.3338
R1030 VSS.n2760 VSS.t423 53.3338
R1031 VSS.n2743 VSS.t441 53.3338
R1032 VSS.n2661 VSS.t425 53.3338
R1033 VSS.n2644 VSS.t509 53.3338
R1034 VSS.n2562 VSS.t620 53.3338
R1035 VSS.n2545 VSS.t692 53.3338
R1036 VSS.n2463 VSS.t626 53.3338
R1037 VSS.n2446 VSS.t38 53.3338
R1038 VSS.n2364 VSS.t544 53.3338
R1039 VSS.n2347 VSS.t57 53.3338
R1040 VSS.n2265 VSS.t427 53.3338
R1041 VSS.n2248 VSS.t321 53.3338
R1042 VSS.n53 VSS.n52 51.0594
R1043 VSS.n120 VSS.n119 51.0594
R1044 VSS.n2974 VSS.t217 45.0709
R1045 VSS.n2983 VSS.t663 45.0709
R1046 VSS.n3123 VSS.t394 45.0709
R1047 VSS.n3112 VSS.t570 45.0709
R1048 VSS.n234 VSS.n233 41.945
R1049 VSS.n239 VSS.n238 41.945
R1050 VSS.n250 VSS.n249 41.945
R1051 VSS.n261 VSS.n260 41.945
R1052 VSS.n751 VSS.n744 41.7468
R1053 VSS.n591 VSS.n584 41.7468
R1054 VSS.n439 VSS.n432 41.7468
R1055 VSS.n332 VSS.n325 41.7468
R1056 VSS.n921 VSS.n912 41.6587
R1057 VSS.n1132 VSS.n1123 41.6587
R1058 VSS.n1251 VSS.n1241 41.6587
R1059 VSS.n1041 VSS.n1031 41.6587
R1060 VSS.n826 VSS.n824 41.6587
R1061 VSS.n733 VSS.n732 41.6587
R1062 VSS.n666 VSS.n664 41.6587
R1063 VSS.n573 VSS.n572 41.6587
R1064 VSS.n532 VSS.n531 41.6587
R1065 VSS.n496 VSS.n495 41.6587
R1066 VSS.n451 VSS.n450 41.6587
R1067 VSS.n389 VSS.n388 41.6587
R1068 VSS.n344 VSS.n343 41.6587
R1069 VSS.n282 VSS.n281 41.6587
R1070 VSS.n40 VSS.n29 41.4233
R1071 VSS.n55 VSS.n46 41.4233
R1072 VSS.n107 VSS.n97 41.4233
R1073 VSS.n122 VSS.n113 41.4233
R1074 VSS.n173 VSS.n164 41.4233
R1075 VSS.n215 VSS.n206 41.4233
R1076 VSS.n1144 VSS.t332 40.6159
R1077 VSS.n933 VSS.t452 40.6159
R1078 VSS.n798 VSS.t152 40.6159
R1079 VSS.n638 VSS.t370 40.6159
R1080 VSS.n2887 VSS.t631 38.5719
R1081 VSS.n2887 VSS.t25 38.5719
R1082 VSS.n2863 VSS.t549 38.5719
R1083 VSS.n2824 VSS.t629 38.5719
R1084 VSS.n2788 VSS.t165 38.5719
R1085 VSS.n2788 VSS.t270 38.5719
R1086 VSS.n2764 VSS.t424 38.5719
R1087 VSS.n2725 VSS.t420 38.5719
R1088 VSS.n2689 VSS.t82 38.5719
R1089 VSS.n2689 VSS.t130 38.5719
R1090 VSS.n2665 VSS.t426 38.5719
R1091 VSS.n2626 VSS.t430 38.5719
R1092 VSS.n2590 VSS.t407 38.5719
R1093 VSS.n2590 VSS.t607 38.5719
R1094 VSS.n2566 VSS.t621 38.5719
R1095 VSS.n2527 VSS.t619 38.5719
R1096 VSS.n2491 VSS.t279 38.5719
R1097 VSS.n2491 VSS.t200 38.5719
R1098 VSS.n2467 VSS.t627 38.5719
R1099 VSS.n2428 VSS.t537 38.5719
R1100 VSS.n2392 VSS.t11 38.5719
R1101 VSS.n2392 VSS.t9 38.5719
R1102 VSS.n2368 VSS.t545 38.5719
R1103 VSS.n2329 VSS.t541 38.5719
R1104 VSS.n2293 VSS.t88 38.5719
R1105 VSS.n2293 VSS.t54 38.5719
R1106 VSS.n2269 VSS.t428 38.5719
R1107 VSS.n2230 VSS.t539 38.5719
R1108 VSS.n1440 VSS.t365 38.5719
R1109 VSS.n1479 VSS.t196 38.5719
R1110 VSS.n1508 VSS.t120 38.5719
R1111 VSS.n1508 VSS.t405 38.5719
R1112 VSS.n1554 VSS.t369 38.5719
R1113 VSS.n1593 VSS.t18 38.5719
R1114 VSS.n1622 VSS.t526 38.5719
R1115 VSS.n1622 VSS.t637 38.5719
R1116 VSS.n1668 VSS.t138 38.5719
R1117 VSS.n1707 VSS.t585 38.5719
R1118 VSS.n1736 VSS.t312 38.5719
R1119 VSS.n1736 VSS.t633 38.5719
R1120 VSS.n1782 VSS.t80 38.5719
R1121 VSS.n1821 VSS.t361 38.5719
R1122 VSS.n1850 VSS.t135 38.5719
R1123 VSS.n1850 VSS.t192 38.5719
R1124 VSS.n1896 VSS.t489 38.5719
R1125 VSS.n1935 VSS.t32 38.5719
R1126 VSS.n1964 VSS.t101 38.5719
R1127 VSS.n1964 VSS.t265 38.5719
R1128 VSS.n2010 VSS.t16 38.5719
R1129 VSS.n2049 VSS.t109 38.5719
R1130 VSS.n2078 VSS.t148 38.5719
R1131 VSS.n2078 VSS.t522 38.5719
R1132 VSS.n2124 VSS.t34 38.5719
R1133 VSS.n2163 VSS.t105 38.5719
R1134 VSS.n2193 VSS.t98 38.5719
R1135 VSS.n2193 VSS.t204 38.5719
R1136 VSS.n1171 VSS.n1170 34.7652
R1137 VSS.n1157 VSS.n1156 34.7652
R1138 VSS.n52 VSS.n51 34.7652
R1139 VSS.n1141 VSS.n1140 34.7652
R1140 VSS.n1127 VSS.n1126 34.7652
R1141 VSS.n1111 VSS.n1110 34.7652
R1142 VSS.n1097 VSS.n1096 34.7652
R1143 VSS.n62 VSS.n61 34.7652
R1144 VSS.n960 VSS.n959 34.7652
R1145 VSS.n946 VSS.n945 34.7652
R1146 VSS.n119 VSS.n118 34.7652
R1147 VSS.n930 VSS.n929 34.7652
R1148 VSS.n916 VSS.n915 34.7652
R1149 VSS.n900 VSS.n899 34.7652
R1150 VSS.n886 VSS.n885 34.7652
R1151 VSS.n129 VSS.n128 34.7652
R1152 VSS.n0 VSS.t508 33.462
R1153 VSS.n0 VSS.t244 33.462
R1154 VSS.n3047 VSS.t84 33.462
R1155 VSS.n3047 VSS.t353 33.462
R1156 VSS.n875 VSS.n874 31.2934
R1157 VSS.n167 VSS.n166 28.061
R1158 VSS.n209 VSS.n208 28.061
R1159 VSS.n1232 VSS.t450 27.0774
R1160 VSS.n86 VSS.n85 27.0774
R1161 VSS.n88 VSS.n87 27.0774
R1162 VSS.n1066 VSS.n1065 27.0774
R1163 VSS.n1052 VSS.n1051 27.0774
R1164 VSS.n1037 VSS.n1036 27.0774
R1165 VSS.n1021 VSS.n1020 27.0774
R1166 VSS.n100 VSS.n99 27.0774
R1167 VSS.n1005 VSS.n1004 27.0774
R1168 VSS.n991 VSS.n990 27.0774
R1169 VSS.n521 VSS.t411 27.0774
R1170 VSS.n506 VSS.t644 27.0774
R1171 VSS.n399 VSS.t334 27.0774
R1172 VSS.n292 VSS.t491 27.0774
R1173 VSS.n1471 VSS.t208 26.8298
R1174 VSS.n1585 VSS.t132 26.8298
R1175 VSS.n1699 VSS.t141 26.8298
R1176 VSS.n1813 VSS.t207 26.8298
R1177 VSS.n1927 VSS.t707 26.8298
R1178 VSS.n2041 VSS.t609 26.8298
R1179 VSS.n2155 VSS.t62 26.8298
R1180 VSS.n1295 VSS.t111 25.9346
R1181 VSS.n1300 VSS.t188 25.9346
R1182 VSS.n1311 VSS.t531 25.9346
R1183 VSS.n1316 VSS.t262 25.9346
R1184 VSS.n1327 VSS.t285 25.9346
R1185 VSS.n1332 VSS.t5 25.9346
R1186 VSS.n1343 VSS.t702 25.9346
R1187 VSS.n1348 VSS.t581 25.9346
R1188 VSS.n1359 VSS.t74 25.9346
R1189 VSS.n1364 VSS.t182 25.9346
R1190 VSS.n1375 VSS.t683 25.9346
R1191 VSS.n1380 VSS.t449 25.9346
R1192 VSS.n1391 VSS.t175 25.9346
R1193 VSS.n1396 VSS.t167 25.9346
R1194 VSS.n1407 VSS.t559 25.9346
R1195 VSS.n1421 VSS.t157 25.9346
R1196 VSS.n1521 VSS.t300 25.9346
R1197 VSS.n1535 VSS.t254 25.9346
R1198 VSS.n1635 VSS.t687 25.9346
R1199 VSS.n1649 VSS.t294 25.9346
R1200 VSS.n1749 VSS.t355 25.9346
R1201 VSS.n1763 VSS.t573 25.9346
R1202 VSS.n1863 VSS.t717 25.9346
R1203 VSS.n1877 VSS.t596 25.9346
R1204 VSS.n1977 VSS.t611 25.9346
R1205 VSS.n1991 VSS.t518 25.9346
R1206 VSS.n2091 VSS.t3 25.9346
R1207 VSS.n2105 VSS.t602 25.9346
R1208 VSS.n9 VSS.t206 25.4291
R1209 VSS.n56 VSS.t579 25.4291
R1210 VSS.n78 VSS.t179 25.4291
R1211 VSS.n123 VSS.t325 25.4291
R1212 VSS.n145 VSS.t267 25.4291
R1213 VSS.n180 VSS.t277 25.4291
R1214 VSS.n187 VSS.t22 25.4291
R1215 VSS.n222 VSS.t447 25.4291
R1216 VSS.n228 VSS.t613 25.4291
R1217 VSS.n240 VSS.t445 25.4291
R1218 VSS.n461 VSS.t90 25.4291
R1219 VSS.n251 VSS.t290 25.4291
R1220 VSS.n354 VSS.t416 25.4291
R1221 VSS.n262 VSS.t41 25.4291
R1222 VSS.n3066 VSS.t339 24.9236
R1223 VSS.n3066 VSS.t60 24.9236
R1224 VSS.n3077 VSS.t341 24.9236
R1225 VSS.n3077 VSS.t345 24.9236
R1226 VSS.n3177 VSS.t381 24.9236
R1227 VSS.n3177 VSS.t401 24.9236
R1228 VSS.n3167 VSS.t379 24.9236
R1229 VSS.n3167 VSS.t397 24.9236
R1230 VSS.n3163 VSS.t375 24.9236
R1231 VSS.n3163 VSS.t393 24.9236
R1232 VSS.n3153 VSS.t373 24.9236
R1233 VSS.n3153 VSS.t389 24.9236
R1234 VSS.n3141 VSS.t387 24.9236
R1235 VSS.n3141 VSS.t403 24.9236
R1236 VSS.n3131 VSS.t385 24.9236
R1237 VSS.n3131 VSS.t399 24.9236
R1238 VSS.n3121 VSS.t377 24.9236
R1239 VSS.n3121 VSS.t395 24.9236
R1240 VSS.n3116 VSS.t383 24.9236
R1241 VSS.n3116 VSS.t571 24.9236
R1242 VSS.n3106 VSS.t563 24.9236
R1243 VSS.n3106 VSS.t569 24.9236
R1244 VSS.n3096 VSS.t561 24.9236
R1245 VSS.n3096 VSS.t567 24.9236
R1246 VSS.n2916 VSS.t230 24.9236
R1247 VSS.n2916 VSS.t224 24.9236
R1248 VSS.n2924 VSS.t240 24.9236
R1249 VSS.n2924 VSS.t220 24.9236
R1250 VSS.n2934 VSS.t236 24.9236
R1251 VSS.n2934 VSS.t214 24.9236
R1252 VSS.n2944 VSS.t232 24.9236
R1253 VSS.n2944 VSS.t212 24.9236
R1254 VSS.n2952 VSS.t228 24.9236
R1255 VSS.n2952 VSS.t222 24.9236
R1256 VSS.n2962 VSS.t226 24.9236
R1257 VSS.n2962 VSS.t216 24.9236
R1258 VSS.n2972 VSS.t238 24.9236
R1259 VSS.n2972 VSS.t218 24.9236
R1260 VSS.n2978 VSS.t234 24.9236
R1261 VSS.n2978 VSS.t664 24.9236
R1262 VSS.n2987 VSS.t670 24.9236
R1263 VSS.n2987 VSS.t662 24.9236
R1264 VSS.n2997 VSS.t668 24.9236
R1265 VSS.n2997 VSS.t660 24.9236
R1266 VSS.n3023 VSS.t711 24.9236
R1267 VSS.n3023 VSS.t709 24.9236
R1268 VSS.n3032 VSS.t713 24.9236
R1269 VSS.n3032 VSS.t1 24.9236
R1270 VSS.n1196 VSS.n1193 24.0332
R1271 VSS.n1193 VSS.n1190 24.0332
R1272 VSS.n1190 VSS.n1187 24.0332
R1273 VSS.n1187 VSS.n1184 24.0332
R1274 VSS.n1184 VSS.n1181 24.0332
R1275 VSS.n1085 VSS.n1082 24.0332
R1276 VSS.n985 VSS.n982 24.0332
R1277 VSS.n982 VSS.n979 24.0332
R1278 VSS.n979 VSS.n976 24.0332
R1279 VSS.n976 VSS.n973 24.0332
R1280 VSS.n973 VSS.n970 24.0332
R1281 VSS.n777 VSS.n774 24.0332
R1282 VSS.n774 VSS.n771 24.0332
R1283 VSS.n771 VSS.n768 24.0332
R1284 VSS.n768 VSS.n765 24.0332
R1285 VSS.n765 VSS.n762 24.0332
R1286 VSS.n762 VSS.n759 24.0332
R1287 VSS.n617 VSS.n614 24.0332
R1288 VSS.n614 VSS.n611 24.0332
R1289 VSS.n611 VSS.n608 24.0332
R1290 VSS.n608 VSS.n605 24.0332
R1291 VSS.n605 VSS.n602 24.0332
R1292 VSS.n602 VSS.n599 24.0332
R1293 VSS.n427 VSS.n424 24.0332
R1294 VSS.n424 VSS.n421 24.0332
R1295 VSS.n421 VSS.n418 24.0332
R1296 VSS.n418 VSS.n415 24.0332
R1297 VSS.n415 VSS.n412 24.0332
R1298 VSS.n412 VSS.n409 24.0332
R1299 VSS.n320 VSS.n317 24.0332
R1300 VSS.n317 VSS.n314 24.0332
R1301 VSS.n314 VSS.n311 24.0332
R1302 VSS.n311 VSS.n308 24.0332
R1303 VSS.n308 VSS.n305 24.0332
R1304 VSS.n305 VSS.n302 24.0332
R1305 VSS.n715 VSS.n714 23.7899
R1306 VSS.n555 VSS.n554 23.7899
R1307 VSS.n477 VSS.n474 23.7089
R1308 VSS.n370 VSS.n367 23.7089
R1309 VSS.n1197 VSS.n1196 23.245
R1310 VSS.n986 VSS.n985 22.9432
R1311 VSS.n2922 VSS.t239 22.5357
R1312 VSS.n2928 VSS.t219 22.5357
R1313 VSS.n3173 VSS.t378 22.5357
R1314 VSS.n3169 VSS.t396 22.5357
R1315 VSS.n66 VSS.n65 22.2316
R1316 VSS.n133 VSS.n132 22.2316
R1317 VSS.n554 VSS.n551 22.1686
R1318 VSS.n516 VSS.n513 22.1686
R1319 VSS.n483 VSS.n477 22.1686
R1320 VSS.n409 VSS.n406 22.1686
R1321 VSS.n376 VSS.n370 22.1686
R1322 VSS.n302 VSS.n299 22.1686
R1323 VSS.n1181 VSS.n1178 21.7362
R1324 VSS.n970 VSS.n967 21.7362
R1325 VSS.n3090 VSS.n3085 20.3039
R1326 VSS.n2796 VSS.n1302 20.3039
R1327 VSS.n2697 VSS.n1318 20.3039
R1328 VSS.n2598 VSS.n1334 20.3039
R1329 VSS.n2499 VSS.n1350 20.3039
R1330 VSS.n2400 VSS.n1366 20.3039
R1331 VSS.n2301 VSS.n1382 20.3039
R1332 VSS.n1516 VSS.n1403 20.3039
R1333 VSS.n1630 VSS.n1402 20.3039
R1334 VSS.n1744 VSS.n1401 20.3039
R1335 VSS.n1858 VSS.n1400 20.3039
R1336 VSS.n1972 VSS.n1399 20.3039
R1337 VSS.n2086 VSS.n1398 20.3039
R1338 VSS.n3017 VSS.n3008 20.3039
R1339 VSS.n778 VSS.n777 18.7186
R1340 VSS.n618 VSS.n617 18.7186
R1341 VSS.n874 VSS.n871 18.1151
R1342 VSS.n714 VSS.n711 18.1151
R1343 VSS.n2855 VSS.t646 17.7783
R1344 VSS.n2756 VSS.t678 17.7783
R1345 VSS.n2657 VSS.t180 17.7783
R1346 VSS.n2558 VSS.t301 17.7783
R1347 VSS.n2459 VSS.t523 17.7783
R1348 VSS.n2360 VSS.t61 17.7783
R1349 VSS.n2261 VSS.t490 17.7783
R1350 VSS.n3057 VSS 16.7729
R1351 VSS.n3042 VSS 16.7729
R1352 VSS.n1086 VSS.n1085 15.0975
R1353 VSS.n1082 VSS.n1079 13.8904
R1354 VSS.n20 VSS.n19 13.539
R1355 VSS.n22 VSS.n21 13.539
R1356 VSS.n1276 VSS.n1275 13.539
R1357 VSS.n1262 VSS.n1261 13.539
R1358 VSS.n1247 VSS.n1246 13.539
R1359 VSS.n1231 VSS.n1230 13.539
R1360 VSS.n33 VSS.n32 13.539
R1361 VSS.n1216 VSS.n1215 13.539
R1362 VSS.n1202 VSS.n1201 13.539
R1363 VSS.n1130 VSS.t474 13.539
R1364 VSS.n1022 VSS.t91 13.539
R1365 VSS.n919 VSS.t470 13.539
R1366 VSS.n152 VSS.n151 13.539
R1367 VSS.n156 VSS.n155 13.539
R1368 VSS.n859 VSS.n858 13.539
R1369 VSS.n846 VSS.n845 13.539
R1370 VSS.n832 VSS.n831 13.539
R1371 VSS.n815 VSS.n814 13.539
R1372 VSS.n170 VSS.n169 13.539
R1373 VSS.n798 VSS.n797 13.539
R1374 VSS.n784 VSS.n783 13.539
R1375 VSS.n194 VSS.n193 13.539
R1376 VSS.n198 VSS.n197 13.539
R1377 VSS.n699 VSS.n698 13.539
R1378 VSS.n686 VSS.n685 13.539
R1379 VSS.n672 VSS.n671 13.539
R1380 VSS.n655 VSS.n654 13.539
R1381 VSS.n212 VSS.n211 13.539
R1382 VSS.n638 VSS.n637 13.539
R1383 VSS.n624 VSS.n623 13.539
R1384 VSS.n2906 VSS.n2901 13.0559
R1385 VSS.n44 VSS.n43 12.8005
R1386 VSS.n111 VSS.n110 12.8005
R1387 VSS.n2790 VSS.n1302 12.5798
R1388 VSS.n2691 VSS.n1318 12.5798
R1389 VSS.n2592 VSS.n1334 12.5798
R1390 VSS.n2493 VSS.n1350 12.5798
R1391 VSS.n2394 VSS.n1366 12.5798
R1392 VSS.n2295 VSS.n1382 12.5798
R1393 VSS.n2897 VSS.n2889 12.5798
R1394 VSS.n551 VSS.n227 12.5798
R1395 VSS.n428 VSS.n427 12.242
R1396 VSS.n321 VSS.n320 12.242
R1397 VSS.n471 VSS.n242 11.9177
R1398 VSS.n364 VSS.n253 11.9177
R1399 VSS.n759 VSS.n756 11.7196
R1400 VSS.n599 VSS.n596 11.7196
R1401 VSS.n82 VSS.n81 11.5887
R1402 VSS.n92 VSS.n91 11.5887
R1403 VSS.n1064 VSS.n1063 11.5887
R1404 VSS.n1050 VSS.n1049 11.5887
R1405 VSS.n1035 VSS.n1034 11.5887
R1406 VSS.n1019 VSS.n1018 11.5887
R1407 VSS.n104 VSS.n103 11.5887
R1408 VSS.n1003 VSS.n1002 11.5887
R1409 VSS.n989 VSS.n988 11.5887
R1410 VSS.n67 VSS.n66 11.214
R1411 VSS.n134 VSS.n133 11.214
R1412 VSS.n3171 VSS.n3168 10.1522
R1413 VSS.n2926 VSS.n2925 10.1522
R1414 VSS.n162 VSS.n161 9.93153
R1415 VSS.n204 VSS.n203 9.93153
R1416 VSS.n2867 VSS.n2864 9.71084
R1417 VSS.n2768 VSS.n2765 9.71084
R1418 VSS.n2669 VSS.n2666 9.71084
R1419 VSS.n2570 VSS.n2567 9.71084
R1420 VSS.n2471 VSS.n2468 9.71084
R1421 VSS.n2372 VSS.n2369 9.71084
R1422 VSS.n2273 VSS.n2270 9.71084
R1423 VSS.n1483 VSS.n1480 9.71084
R1424 VSS.n1597 VSS.n1594 9.71084
R1425 VSS.n1711 VSS.n1708 9.71084
R1426 VSS.n1825 VSS.n1822 9.71084
R1427 VSS.n1939 VSS.n1936 9.71084
R1428 VSS.n2053 VSS.n2050 9.71084
R1429 VSS.n2167 VSS.n2164 9.71084
R1430 VSS.n27 VSS.n24 9.3005
R1431 VSS.n24 VSS.n23 9.3005
R1432 VSS.n1265 VSS.n1264 9.3005
R1433 VSS.n1264 VSS.n1263 9.3005
R1434 VSS.n1234 VSS.n1233 9.3005
R1435 VSS.n1233 VSS.n1232 9.3005
R1436 VSS.n1219 VSS.n1218 9.3005
R1437 VSS.n1218 VSS.n1217 9.3005
R1438 VSS.n1176 VSS.n1175 9.3005
R1439 VSS.n1175 VSS.n1174 9.3005
R1440 VSS.n1162 VSS.n1161 9.3005
R1441 VSS.n1161 VSS.n1160 9.3005
R1442 VSS.n50 VSS.n49 9.3005
R1443 VSS.n1146 VSS.n1145 9.3005
R1444 VSS.n1145 VSS.n1144 9.3005
R1445 VSS.n1132 VSS.n1131 9.3005
R1446 VSS.n1131 VSS.n1130 9.3005
R1447 VSS.n1116 VSS.n1115 9.3005
R1448 VSS.n1115 VSS.n1114 9.3005
R1449 VSS.n1102 VSS.n1101 9.3005
R1450 VSS.n1101 VSS.n1100 9.3005
R1451 VSS.n69 VSS.n68 9.3005
R1452 VSS.n70 VSS.n69 9.3005
R1453 VSS.n75 VSS.n74 9.3005
R1454 VSS.n74 VSS.n73 9.3005
R1455 VSS.n90 VSS.n89 9.3005
R1456 VSS.n1055 VSS.n1054 9.3005
R1457 VSS.n1054 VSS.n1053 9.3005
R1458 VSS.n1024 VSS.n1023 9.3005
R1459 VSS.n1023 VSS.n1022 9.3005
R1460 VSS.n1008 VSS.n1007 9.3005
R1461 VSS.n1007 VSS.n1006 9.3005
R1462 VSS.n965 VSS.n964 9.3005
R1463 VSS.n964 VSS.n963 9.3005
R1464 VSS.n951 VSS.n950 9.3005
R1465 VSS.n950 VSS.n949 9.3005
R1466 VSS.n117 VSS.n116 9.3005
R1467 VSS.n935 VSS.n934 9.3005
R1468 VSS.n934 VSS.n933 9.3005
R1469 VSS.n921 VSS.n920 9.3005
R1470 VSS.n920 VSS.n919 9.3005
R1471 VSS.n905 VSS.n904 9.3005
R1472 VSS.n904 VSS.n903 9.3005
R1473 VSS.n891 VSS.n890 9.3005
R1474 VSS.n890 VSS.n889 9.3005
R1475 VSS.n136 VSS.n135 9.3005
R1476 VSS.n137 VSS.n136 9.3005
R1477 VSS.n142 VSS.n141 9.3005
R1478 VSS.n141 VSS.n140 9.3005
R1479 VSS.n150 VSS.n143 9.3005
R1480 VSS.n151 VSS.n150 9.3005
R1481 VSS.n157 VSS.n156 9.3005
R1482 VSS.n861 VSS.n860 9.3005
R1483 VSS.n860 VSS.n859 9.3005
R1484 VSS.n848 VSS.n847 9.3005
R1485 VSS.n847 VSS.n846 9.3005
R1486 VSS.n834 VSS.n833 9.3005
R1487 VSS.n833 VSS.n832 9.3005
R1488 VSS.n817 VSS.n816 9.3005
R1489 VSS.n816 VSS.n815 9.3005
R1490 VSS.n172 VSS.n171 9.3005
R1491 VSS.n171 VSS.n170 9.3005
R1492 VSS.n800 VSS.n799 9.3005
R1493 VSS.n799 VSS.n798 9.3005
R1494 VSS.n786 VSS.n785 9.3005
R1495 VSS.n785 VSS.n784 9.3005
R1496 VSS.n192 VSS.n185 9.3005
R1497 VSS.n193 VSS.n192 9.3005
R1498 VSS.n199 VSS.n198 9.3005
R1499 VSS.n701 VSS.n700 9.3005
R1500 VSS.n700 VSS.n699 9.3005
R1501 VSS.n688 VSS.n687 9.3005
R1502 VSS.n687 VSS.n686 9.3005
R1503 VSS.n674 VSS.n673 9.3005
R1504 VSS.n673 VSS.n672 9.3005
R1505 VSS.n657 VSS.n656 9.3005
R1506 VSS.n656 VSS.n655 9.3005
R1507 VSS.n214 VSS.n213 9.3005
R1508 VSS.n213 VSS.n212 9.3005
R1509 VSS.n640 VSS.n639 9.3005
R1510 VSS.n639 VSS.n638 9.3005
R1511 VSS.n626 VSS.n625 9.3005
R1512 VSS.n625 VSS.n624 9.3005
R1513 VSS.n994 VSS.n993 9.3005
R1514 VSS.n993 VSS.n992 9.3005
R1515 VSS.n102 VSS.n101 9.3005
R1516 VSS.n1040 VSS.n1039 9.3005
R1517 VSS.n1039 VSS.n1038 9.3005
R1518 VSS.n1069 VSS.n1068 9.3005
R1519 VSS.n1068 VSS.n1067 9.3005
R1520 VSS.n83 VSS.n76 9.3005
R1521 VSS.n84 VSS.n83 9.3005
R1522 VSS.n1205 VSS.n1204 9.3005
R1523 VSS.n1204 VSS.n1203 9.3005
R1524 VSS.n35 VSS.n34 9.3005
R1525 VSS.n1250 VSS.n1249 9.3005
R1526 VSS.n1249 VSS.n1248 9.3005
R1527 VSS.n1279 VSS.n1278 9.3005
R1528 VSS.n1278 VSS.n1277 9.3005
R1529 VSS.n17 VSS.n8 9.3005
R1530 VSS.n18 VSS.n17 9.3005
R1531 VSS.n3119 VSS.n3117 9.26947
R1532 VSS.n2981 VSS.n2979 9.26947
R1533 VSS.n3022 VSS.n3021 9.01832
R1534 VSS.n3076 VSS.n3075 9.01832
R1535 VSS.n3 VSS.n2 9.01734
R1536 VSS.n1299 VSS.n1298 9.01662
R1537 VSS.n1315 VSS.n1314 9.01662
R1538 VSS.n1331 VSS.n1330 9.01662
R1539 VSS.n1347 VSS.n1346 9.01662
R1540 VSS.n1363 VSS.n1362 9.01662
R1541 VSS.n1379 VSS.n1378 9.01662
R1542 VSS.n1395 VSS.n1394 9.01662
R1543 VSS.n1520 VSS.n1519 9.01662
R1544 VSS.n1634 VSS.n1633 9.01662
R1545 VSS.n1748 VSS.n1747 9.01662
R1546 VSS.n1862 VSS.n1861 9.01662
R1547 VSS.n1976 VSS.n1975 9.01662
R1548 VSS.n2090 VSS.n2089 9.01662
R1549 VSS.n1406 VSS.n1405 9.01662
R1550 VSS.n1294 VSS.n1293 9.01654
R1551 VSS.n1310 VSS.n1309 9.01654
R1552 VSS.n1326 VSS.n1325 9.01654
R1553 VSS.n1342 VSS.n1341 9.01654
R1554 VSS.n1358 VSS.n1357 9.01654
R1555 VSS.n1374 VSS.n1373 9.01654
R1556 VSS.n1390 VSS.n1389 9.01654
R1557 VSS.n1420 VSS.n1419 9.01654
R1558 VSS.n1534 VSS.n1533 9.01654
R1559 VSS.n1648 VSS.n1647 9.01654
R1560 VSS.n1762 VSS.n1761 9.01654
R1561 VSS.n1876 VSS.n1875 9.01654
R1562 VSS.n1990 VSS.n1989 9.01654
R1563 VSS.n2104 VSS.n2103 9.01654
R1564 VSS.n2791 VSS.n2790 9.01634
R1565 VSS.n2692 VSS.n2691 9.01634
R1566 VSS.n2593 VSS.n2592 9.01634
R1567 VSS.n2494 VSS.n2493 9.01634
R1568 VSS.n2395 VSS.n2394 9.01634
R1569 VSS.n2296 VSS.n2295 9.01634
R1570 VSS.n2894 VSS.n2889 9.01634
R1571 VSS.n1511 VSS.n1510 9.01634
R1572 VSS.n1625 VSS.n1624 9.01634
R1573 VSS.n1739 VSS.n1738 9.01634
R1574 VSS.n1853 VSS.n1852 9.01634
R1575 VSS.n1967 VSS.n1966 9.01634
R1576 VSS.n2081 VSS.n2080 9.01634
R1577 VSS.n2192 VSS.n2191 9.01634
R1578 VSS.n547 VSS.n227 9.01634
R1579 VSS.n479 VSS.n478 9.01634
R1580 VSS.n372 VSS.n371 9.01634
R1581 VSS.n265 VSS.n264 9.01634
R1582 VSS.n3046 VSS.n3045 9.01634
R1583 VSS.n1290 VSS.n1289 9.01617
R1584 VSS.n1306 VSS.n1305 9.01617
R1585 VSS.n1322 VSS.n1321 9.01617
R1586 VSS.n1338 VSS.n1337 9.01617
R1587 VSS.n1354 VSS.n1353 9.01617
R1588 VSS.n1370 VSS.n1369 9.01617
R1589 VSS.n1386 VSS.n1385 9.01617
R1590 VSS.n1499 VSS.n1498 9.01617
R1591 VSS.n1613 VSS.n1612 9.01617
R1592 VSS.n1727 VSS.n1726 9.01617
R1593 VSS.n1841 VSS.n1840 9.01617
R1594 VSS.n1955 VSS.n1954 9.01617
R1595 VSS.n2069 VSS.n2068 9.01617
R1596 VSS.n2183 VSS.n2182 9.01617
R1597 VSS.n232 VSS.n231 9.01549
R1598 VSS.n237 VSS.n236 9.01549
R1599 VSS.n248 VSS.n247 9.01549
R1600 VSS.n259 VSS.n258 9.01549
R1601 VSS.n2891 VSS.n2890 9.01392
R1602 VSS.n2892 VSS.n2891 9.01392
R1603 VSS.n1412 VSS.n1411 9.01392
R1604 VSS.n1416 VSS.n1415 9.01392
R1605 VSS.n1426 VSS.n1425 9.01392
R1606 VSS.n1430 VSS.n1429 9.01392
R1607 VSS.n1434 VSS.n1433 9.01392
R1608 VSS.n1438 VSS.n1437 9.01392
R1609 VSS.n1444 VSS.n1443 9.01392
R1610 VSS.n1448 VSS.n1447 9.01392
R1611 VSS.n1452 VSS.n1451 9.01392
R1612 VSS.n1456 VSS.n1455 9.01392
R1613 VSS.n1460 VSS.n1459 9.01392
R1614 VSS.n1465 VSS.n1464 9.01392
R1615 VSS.n1469 VSS.n1468 9.01392
R1616 VSS.n1473 VSS.n1472 9.01392
R1617 VSS.n1477 VSS.n1476 9.01392
R1618 VSS.n1483 VSS.n1482 9.01392
R1619 VSS.n1487 VSS.n1486 9.01392
R1620 VSS.n1491 VSS.n1490 9.01392
R1621 VSS.n1495 VSS.n1494 9.01392
R1622 VSS.n1504 VSS.n1503 9.01392
R1623 VSS.n1513 VSS.n1403 9.01392
R1624 VSS VSS.n1513 9.01392
R1625 VSS.n1516 VSS.n1515 9.01392
R1626 VSS.n1526 VSS.n1525 9.01392
R1627 VSS.n1530 VSS.n1529 9.01392
R1628 VSS.n1540 VSS.n1539 9.01392
R1629 VSS.n1544 VSS.n1543 9.01392
R1630 VSS.n1548 VSS.n1547 9.01392
R1631 VSS.n1552 VSS.n1551 9.01392
R1632 VSS.n1558 VSS.n1557 9.01392
R1633 VSS.n1562 VSS.n1561 9.01392
R1634 VSS.n1566 VSS.n1565 9.01392
R1635 VSS.n1570 VSS.n1569 9.01392
R1636 VSS.n1574 VSS.n1573 9.01392
R1637 VSS.n1579 VSS.n1578 9.01392
R1638 VSS.n1583 VSS.n1582 9.01392
R1639 VSS.n1587 VSS.n1586 9.01392
R1640 VSS.n1591 VSS.n1590 9.01392
R1641 VSS.n1597 VSS.n1596 9.01392
R1642 VSS.n1601 VSS.n1600 9.01392
R1643 VSS.n1605 VSS.n1604 9.01392
R1644 VSS.n1609 VSS.n1608 9.01392
R1645 VSS.n1618 VSS.n1617 9.01392
R1646 VSS.n1627 VSS.n1402 9.01392
R1647 VSS VSS.n1627 9.01392
R1648 VSS.n1630 VSS.n1629 9.01392
R1649 VSS.n1640 VSS.n1639 9.01392
R1650 VSS.n1644 VSS.n1643 9.01392
R1651 VSS.n1654 VSS.n1653 9.01392
R1652 VSS.n1658 VSS.n1657 9.01392
R1653 VSS.n1662 VSS.n1661 9.01392
R1654 VSS.n1666 VSS.n1665 9.01392
R1655 VSS.n1672 VSS.n1671 9.01392
R1656 VSS.n1676 VSS.n1675 9.01392
R1657 VSS.n1680 VSS.n1679 9.01392
R1658 VSS.n1684 VSS.n1683 9.01392
R1659 VSS.n1688 VSS.n1687 9.01392
R1660 VSS.n1693 VSS.n1692 9.01392
R1661 VSS.n1697 VSS.n1696 9.01392
R1662 VSS.n1701 VSS.n1700 9.01392
R1663 VSS.n1705 VSS.n1704 9.01392
R1664 VSS.n1711 VSS.n1710 9.01392
R1665 VSS.n1715 VSS.n1714 9.01392
R1666 VSS.n1719 VSS.n1718 9.01392
R1667 VSS.n1723 VSS.n1722 9.01392
R1668 VSS.n1732 VSS.n1731 9.01392
R1669 VSS.n1741 VSS.n1401 9.01392
R1670 VSS VSS.n1741 9.01392
R1671 VSS.n1744 VSS.n1743 9.01392
R1672 VSS.n1754 VSS.n1753 9.01392
R1673 VSS.n1758 VSS.n1757 9.01392
R1674 VSS.n1768 VSS.n1767 9.01392
R1675 VSS.n1772 VSS.n1771 9.01392
R1676 VSS.n1776 VSS.n1775 9.01392
R1677 VSS.n1780 VSS.n1779 9.01392
R1678 VSS.n1786 VSS.n1785 9.01392
R1679 VSS.n1790 VSS.n1789 9.01392
R1680 VSS.n1794 VSS.n1793 9.01392
R1681 VSS.n1798 VSS.n1797 9.01392
R1682 VSS.n1802 VSS.n1801 9.01392
R1683 VSS.n1807 VSS.n1806 9.01392
R1684 VSS.n1811 VSS.n1810 9.01392
R1685 VSS.n1815 VSS.n1814 9.01392
R1686 VSS.n1819 VSS.n1818 9.01392
R1687 VSS.n1825 VSS.n1824 9.01392
R1688 VSS.n1829 VSS.n1828 9.01392
R1689 VSS.n1833 VSS.n1832 9.01392
R1690 VSS.n1837 VSS.n1836 9.01392
R1691 VSS.n1846 VSS.n1845 9.01392
R1692 VSS.n1855 VSS.n1400 9.01392
R1693 VSS VSS.n1855 9.01392
R1694 VSS.n1858 VSS.n1857 9.01392
R1695 VSS.n1868 VSS.n1867 9.01392
R1696 VSS.n1872 VSS.n1871 9.01392
R1697 VSS.n1882 VSS.n1881 9.01392
R1698 VSS.n1886 VSS.n1885 9.01392
R1699 VSS.n1890 VSS.n1889 9.01392
R1700 VSS.n1894 VSS.n1893 9.01392
R1701 VSS.n1900 VSS.n1899 9.01392
R1702 VSS.n1904 VSS.n1903 9.01392
R1703 VSS.n1908 VSS.n1907 9.01392
R1704 VSS.n1912 VSS.n1911 9.01392
R1705 VSS.n1916 VSS.n1915 9.01392
R1706 VSS.n1921 VSS.n1920 9.01392
R1707 VSS.n1925 VSS.n1924 9.01392
R1708 VSS.n1929 VSS.n1928 9.01392
R1709 VSS.n1933 VSS.n1932 9.01392
R1710 VSS.n1939 VSS.n1938 9.01392
R1711 VSS.n1943 VSS.n1942 9.01392
R1712 VSS.n1947 VSS.n1946 9.01392
R1713 VSS.n1951 VSS.n1950 9.01392
R1714 VSS.n1960 VSS.n1959 9.01392
R1715 VSS.n1969 VSS.n1399 9.01392
R1716 VSS VSS.n1969 9.01392
R1717 VSS.n1972 VSS.n1971 9.01392
R1718 VSS.n1982 VSS.n1981 9.01392
R1719 VSS.n1986 VSS.n1985 9.01392
R1720 VSS.n1996 VSS.n1995 9.01392
R1721 VSS.n2000 VSS.n1999 9.01392
R1722 VSS.n2004 VSS.n2003 9.01392
R1723 VSS.n2008 VSS.n2007 9.01392
R1724 VSS.n2014 VSS.n2013 9.01392
R1725 VSS.n2018 VSS.n2017 9.01392
R1726 VSS.n2022 VSS.n2021 9.01392
R1727 VSS.n2026 VSS.n2025 9.01392
R1728 VSS.n2030 VSS.n2029 9.01392
R1729 VSS.n2035 VSS.n2034 9.01392
R1730 VSS.n2039 VSS.n2038 9.01392
R1731 VSS.n2043 VSS.n2042 9.01392
R1732 VSS.n2047 VSS.n2046 9.01392
R1733 VSS.n2053 VSS.n2052 9.01392
R1734 VSS.n2057 VSS.n2056 9.01392
R1735 VSS.n2061 VSS.n2060 9.01392
R1736 VSS.n2065 VSS.n2064 9.01392
R1737 VSS.n2074 VSS.n2073 9.01392
R1738 VSS.n2083 VSS.n1398 9.01392
R1739 VSS VSS.n2083 9.01392
R1740 VSS.n2086 VSS.n2085 9.01392
R1741 VSS.n2096 VSS.n2095 9.01392
R1742 VSS.n2100 VSS.n2099 9.01392
R1743 VSS.n2110 VSS.n2109 9.01392
R1744 VSS.n2114 VSS.n2113 9.01392
R1745 VSS.n2118 VSS.n2117 9.01392
R1746 VSS.n2122 VSS.n2121 9.01392
R1747 VSS.n2128 VSS.n2127 9.01392
R1748 VSS.n2132 VSS.n2131 9.01392
R1749 VSS.n2136 VSS.n2135 9.01392
R1750 VSS.n2140 VSS.n2139 9.01392
R1751 VSS.n2144 VSS.n2143 9.01392
R1752 VSS.n2149 VSS.n2148 9.01392
R1753 VSS.n2153 VSS.n2152 9.01392
R1754 VSS.n2157 VSS.n2156 9.01392
R1755 VSS.n2161 VSS.n2160 9.01392
R1756 VSS.n2167 VSS.n2166 9.01392
R1757 VSS.n2171 VSS.n2170 9.01392
R1758 VSS.n2175 VSS.n2174 9.01392
R1759 VSS.n2179 VSS.n2178 9.01392
R1760 VSS.n2188 VSS.n2187 9.01392
R1761 VSS.n289 VSS.n288 9.01392
R1762 VSS.n285 VSS.n284 9.01392
R1763 VSS.n278 VSS.n277 9.01392
R1764 VSS.n274 VSS.n273 9.01392
R1765 VSS.n294 VSS.n293 9.01392
R1766 VSS.n396 VSS.n395 9.01392
R1767 VSS.n392 VSS.n391 9.01392
R1768 VSS.n385 VSS.n384 9.01392
R1769 VSS.n381 VSS.n380 9.01392
R1770 VSS.n376 VSS.n375 9.01392
R1771 VSS.n401 VSS.n400 9.01392
R1772 VSS.n508 VSS.n507 9.01392
R1773 VSS.n503 VSS.n502 9.01392
R1774 VSS.n499 VSS.n498 9.01392
R1775 VSS.n492 VSS.n491 9.01392
R1776 VSS.n488 VSS.n487 9.01392
R1777 VSS.n483 VSS.n482 9.01392
R1778 VSS.n513 VSS.n512 9.01392
R1779 VSS.n543 VSS.n542 9.01392
R1780 VSS.n539 VSS.n538 9.01392
R1781 VSS.n535 VSS.n534 9.01392
R1782 VSS.n528 VSS.n527 9.01392
R1783 VSS.n523 VSS.n522 9.01392
R1784 VSS.n519 VSS.n518 9.01392
R1785 VSS.n551 VSS.n550 9.01392
R1786 VSS.n3052 VSS.n3051 9.01392
R1787 VSS.n3051 VSS.n3050 9.01392
R1788 VSS.n2897 VSS.n2896 9.01392
R1789 VSS.n2896 VSS 9.01392
R1790 VSS.n2884 VSS.n2883 9.01392
R1791 VSS.n2879 VSS.n2878 9.01392
R1792 VSS.n2875 VSS.n2874 9.01392
R1793 VSS.n2871 VSS.n2870 9.01392
R1794 VSS.n2867 VSS.n2866 9.01392
R1795 VSS.n2861 VSS.n2860 9.01392
R1796 VSS.n2857 VSS.n2856 9.01392
R1797 VSS.n2853 VSS.n2852 9.01392
R1798 VSS.n2849 VSS.n2848 9.01392
R1799 VSS.n2844 VSS.n2843 9.01392
R1800 VSS.n2840 VSS.n2839 9.01392
R1801 VSS.n2836 VSS.n2835 9.01392
R1802 VSS.n2832 VSS.n2831 9.01392
R1803 VSS.n2828 VSS.n2827 9.01392
R1804 VSS.n2822 VSS.n2821 9.01392
R1805 VSS.n2818 VSS.n2817 9.01392
R1806 VSS.n2814 VSS.n2813 9.01392
R1807 VSS.n2810 VSS.n2809 9.01392
R1808 VSS.n2805 VSS.n2804 9.01392
R1809 VSS.n2801 VSS.n2800 9.01392
R1810 VSS.n2796 VSS.n2795 9.01392
R1811 VSS.n2793 VSS.n1302 9.01392
R1812 VSS VSS.n2793 9.01392
R1813 VSS.n2785 VSS.n2784 9.01392
R1814 VSS.n2780 VSS.n2779 9.01392
R1815 VSS.n2776 VSS.n2775 9.01392
R1816 VSS.n2772 VSS.n2771 9.01392
R1817 VSS.n2768 VSS.n2767 9.01392
R1818 VSS.n2762 VSS.n2761 9.01392
R1819 VSS.n2758 VSS.n2757 9.01392
R1820 VSS.n2754 VSS.n2753 9.01392
R1821 VSS.n2750 VSS.n2749 9.01392
R1822 VSS.n2745 VSS.n2744 9.01392
R1823 VSS.n2741 VSS.n2740 9.01392
R1824 VSS.n2737 VSS.n2736 9.01392
R1825 VSS.n2733 VSS.n2732 9.01392
R1826 VSS.n2729 VSS.n2728 9.01392
R1827 VSS.n2723 VSS.n2722 9.01392
R1828 VSS.n2719 VSS.n2718 9.01392
R1829 VSS.n2715 VSS.n2714 9.01392
R1830 VSS.n2711 VSS.n2710 9.01392
R1831 VSS.n2706 VSS.n2705 9.01392
R1832 VSS.n2702 VSS.n2701 9.01392
R1833 VSS.n2697 VSS.n2696 9.01392
R1834 VSS.n2694 VSS.n1318 9.01392
R1835 VSS VSS.n2694 9.01392
R1836 VSS.n2686 VSS.n2685 9.01392
R1837 VSS.n2681 VSS.n2680 9.01392
R1838 VSS.n2677 VSS.n2676 9.01392
R1839 VSS.n2673 VSS.n2672 9.01392
R1840 VSS.n2669 VSS.n2668 9.01392
R1841 VSS.n2663 VSS.n2662 9.01392
R1842 VSS.n2659 VSS.n2658 9.01392
R1843 VSS.n2655 VSS.n2654 9.01392
R1844 VSS.n2651 VSS.n2650 9.01392
R1845 VSS.n2646 VSS.n2645 9.01392
R1846 VSS.n2642 VSS.n2641 9.01392
R1847 VSS.n2638 VSS.n2637 9.01392
R1848 VSS.n2634 VSS.n2633 9.01392
R1849 VSS.n2630 VSS.n2629 9.01392
R1850 VSS.n2624 VSS.n2623 9.01392
R1851 VSS.n2620 VSS.n2619 9.01392
R1852 VSS.n2616 VSS.n2615 9.01392
R1853 VSS.n2612 VSS.n2611 9.01392
R1854 VSS.n2607 VSS.n2606 9.01392
R1855 VSS.n2603 VSS.n2602 9.01392
R1856 VSS.n2598 VSS.n2597 9.01392
R1857 VSS.n2595 VSS.n1334 9.01392
R1858 VSS VSS.n2595 9.01392
R1859 VSS.n2587 VSS.n2586 9.01392
R1860 VSS.n2582 VSS.n2581 9.01392
R1861 VSS.n2578 VSS.n2577 9.01392
R1862 VSS.n2574 VSS.n2573 9.01392
R1863 VSS.n2570 VSS.n2569 9.01392
R1864 VSS.n2564 VSS.n2563 9.01392
R1865 VSS.n2560 VSS.n2559 9.01392
R1866 VSS.n2556 VSS.n2555 9.01392
R1867 VSS.n2552 VSS.n2551 9.01392
R1868 VSS.n2547 VSS.n2546 9.01392
R1869 VSS.n2543 VSS.n2542 9.01392
R1870 VSS.n2539 VSS.n2538 9.01392
R1871 VSS.n2535 VSS.n2534 9.01392
R1872 VSS.n2531 VSS.n2530 9.01392
R1873 VSS.n2525 VSS.n2524 9.01392
R1874 VSS.n2521 VSS.n2520 9.01392
R1875 VSS.n2517 VSS.n2516 9.01392
R1876 VSS.n2513 VSS.n2512 9.01392
R1877 VSS.n2508 VSS.n2507 9.01392
R1878 VSS.n2504 VSS.n2503 9.01392
R1879 VSS.n2499 VSS.n2498 9.01392
R1880 VSS.n2496 VSS.n1350 9.01392
R1881 VSS VSS.n2496 9.01392
R1882 VSS.n2488 VSS.n2487 9.01392
R1883 VSS.n2483 VSS.n2482 9.01392
R1884 VSS.n2479 VSS.n2478 9.01392
R1885 VSS.n2475 VSS.n2474 9.01392
R1886 VSS.n2471 VSS.n2470 9.01392
R1887 VSS.n2465 VSS.n2464 9.01392
R1888 VSS.n2461 VSS.n2460 9.01392
R1889 VSS.n2457 VSS.n2456 9.01392
R1890 VSS.n2453 VSS.n2452 9.01392
R1891 VSS.n2448 VSS.n2447 9.01392
R1892 VSS.n2444 VSS.n2443 9.01392
R1893 VSS.n2440 VSS.n2439 9.01392
R1894 VSS.n2436 VSS.n2435 9.01392
R1895 VSS.n2432 VSS.n2431 9.01392
R1896 VSS.n2426 VSS.n2425 9.01392
R1897 VSS.n2422 VSS.n2421 9.01392
R1898 VSS.n2418 VSS.n2417 9.01392
R1899 VSS.n2414 VSS.n2413 9.01392
R1900 VSS.n2409 VSS.n2408 9.01392
R1901 VSS.n2405 VSS.n2404 9.01392
R1902 VSS.n2400 VSS.n2399 9.01392
R1903 VSS.n2397 VSS.n1366 9.01392
R1904 VSS VSS.n2397 9.01392
R1905 VSS.n2389 VSS.n2388 9.01392
R1906 VSS.n2384 VSS.n2383 9.01392
R1907 VSS.n2380 VSS.n2379 9.01392
R1908 VSS.n2376 VSS.n2375 9.01392
R1909 VSS.n2372 VSS.n2371 9.01392
R1910 VSS.n2366 VSS.n2365 9.01392
R1911 VSS.n2362 VSS.n2361 9.01392
R1912 VSS.n2358 VSS.n2357 9.01392
R1913 VSS.n2354 VSS.n2353 9.01392
R1914 VSS.n2349 VSS.n2348 9.01392
R1915 VSS.n2345 VSS.n2344 9.01392
R1916 VSS.n2341 VSS.n2340 9.01392
R1917 VSS.n2337 VSS.n2336 9.01392
R1918 VSS.n2333 VSS.n2332 9.01392
R1919 VSS.n2327 VSS.n2326 9.01392
R1920 VSS.n2323 VSS.n2322 9.01392
R1921 VSS.n2319 VSS.n2318 9.01392
R1922 VSS.n2315 VSS.n2314 9.01392
R1923 VSS.n2310 VSS.n2309 9.01392
R1924 VSS.n2306 VSS.n2305 9.01392
R1925 VSS.n2301 VSS.n2300 9.01392
R1926 VSS.n2298 VSS.n1382 9.01392
R1927 VSS VSS.n2298 9.01392
R1928 VSS.n2290 VSS.n2289 9.01392
R1929 VSS.n2285 VSS.n2284 9.01392
R1930 VSS.n2281 VSS.n2280 9.01392
R1931 VSS.n2277 VSS.n2276 9.01392
R1932 VSS.n2273 VSS.n2272 9.01392
R1933 VSS.n2267 VSS.n2266 9.01392
R1934 VSS.n2263 VSS.n2262 9.01392
R1935 VSS.n2259 VSS.n2258 9.01392
R1936 VSS.n2255 VSS.n2254 9.01392
R1937 VSS.n2250 VSS.n2249 9.01392
R1938 VSS.n2246 VSS.n2245 9.01392
R1939 VSS.n2242 VSS.n2241 9.01392
R1940 VSS.n2238 VSS.n2237 9.01392
R1941 VSS.n2234 VSS.n2233 9.01392
R1942 VSS.n2228 VSS.n2227 9.01392
R1943 VSS.n2224 VSS.n2223 9.01392
R1944 VSS.n2220 VSS.n2219 9.01392
R1945 VSS.n2216 VSS.n2215 9.01392
R1946 VSS.n2211 VSS.n2210 9.01392
R1947 VSS.n2207 VSS.n2206 9.01392
R1948 VSS.n3201 VSS.n3200 9.01392
R1949 VSS.n3200 VSS.n3199 9.01392
R1950 VSS.n3194 VSS.n3193 9.01392
R1951 VSS.n3118 VSS.t382 9.01392
R1952 VSS.n2 VSS.n1 9.01392
R1953 VSS.n1405 VSS.n1404 9.01392
R1954 VSS.n1411 VSS.n1410 9.01392
R1955 VSS.n1415 VSS.n1414 9.01392
R1956 VSS.n1419 VSS.n1418 9.01392
R1957 VSS.n1425 VSS.n1424 9.01392
R1958 VSS.n1429 VSS.n1428 9.01392
R1959 VSS.n1433 VSS.n1432 9.01392
R1960 VSS.n1437 VSS.n1436 9.01392
R1961 VSS.n1443 VSS.n1442 9.01392
R1962 VSS.n1447 VSS.n1446 9.01392
R1963 VSS.n1451 VSS.n1450 9.01392
R1964 VSS.n1455 VSS.n1454 9.01392
R1965 VSS.n1459 VSS.n1458 9.01392
R1966 VSS.n1464 VSS.n1463 9.01392
R1967 VSS.n1468 VSS.n1467 9.01392
R1968 VSS.n1472 VSS.n1471 9.01392
R1969 VSS.n1476 VSS.n1475 9.01392
R1970 VSS.n1482 VSS.n1481 9.01392
R1971 VSS.n1486 VSS.n1485 9.01392
R1972 VSS.n1490 VSS.n1489 9.01392
R1973 VSS.n1494 VSS.n1493 9.01392
R1974 VSS.n1498 VSS.n1497 9.01392
R1975 VSS.n1503 VSS.n1502 9.01392
R1976 VSS.n1512 VSS.n1511 9.01392
R1977 VSS.n1515 VSS.n1514 9.01392
R1978 VSS.n1519 VSS.n1518 9.01392
R1979 VSS.n1525 VSS.n1524 9.01392
R1980 VSS.n1529 VSS.n1528 9.01392
R1981 VSS.n1533 VSS.n1532 9.01392
R1982 VSS.n1539 VSS.n1538 9.01392
R1983 VSS.n1543 VSS.n1542 9.01392
R1984 VSS.n1547 VSS.n1546 9.01392
R1985 VSS.n1551 VSS.n1550 9.01392
R1986 VSS.n1557 VSS.n1556 9.01392
R1987 VSS.n1561 VSS.n1560 9.01392
R1988 VSS.n1565 VSS.n1564 9.01392
R1989 VSS.n1569 VSS.n1568 9.01392
R1990 VSS.n1573 VSS.n1572 9.01392
R1991 VSS.n1578 VSS.n1577 9.01392
R1992 VSS.n1582 VSS.n1581 9.01392
R1993 VSS.n1586 VSS.n1585 9.01392
R1994 VSS.n1590 VSS.n1589 9.01392
R1995 VSS.n1596 VSS.n1595 9.01392
R1996 VSS.n1600 VSS.n1599 9.01392
R1997 VSS.n1604 VSS.n1603 9.01392
R1998 VSS.n1608 VSS.n1607 9.01392
R1999 VSS.n1612 VSS.n1611 9.01392
R2000 VSS.n1617 VSS.n1616 9.01392
R2001 VSS.n1626 VSS.n1625 9.01392
R2002 VSS.n1629 VSS.n1628 9.01392
R2003 VSS.n1633 VSS.n1632 9.01392
R2004 VSS.n1639 VSS.n1638 9.01392
R2005 VSS.n1643 VSS.n1642 9.01392
R2006 VSS.n1647 VSS.n1646 9.01392
R2007 VSS.n1653 VSS.n1652 9.01392
R2008 VSS.n1657 VSS.n1656 9.01392
R2009 VSS.n1661 VSS.n1660 9.01392
R2010 VSS.n1665 VSS.n1664 9.01392
R2011 VSS.n1671 VSS.n1670 9.01392
R2012 VSS.n1675 VSS.n1674 9.01392
R2013 VSS.n1679 VSS.n1678 9.01392
R2014 VSS.n1683 VSS.n1682 9.01392
R2015 VSS.n1687 VSS.n1686 9.01392
R2016 VSS.n1692 VSS.n1691 9.01392
R2017 VSS.n1696 VSS.n1695 9.01392
R2018 VSS.n1700 VSS.n1699 9.01392
R2019 VSS.n1704 VSS.n1703 9.01392
R2020 VSS.n1710 VSS.n1709 9.01392
R2021 VSS.n1714 VSS.n1713 9.01392
R2022 VSS.n1718 VSS.n1717 9.01392
R2023 VSS.n1722 VSS.n1721 9.01392
R2024 VSS.n1726 VSS.n1725 9.01392
R2025 VSS.n1731 VSS.n1730 9.01392
R2026 VSS.n1740 VSS.n1739 9.01392
R2027 VSS.n1743 VSS.n1742 9.01392
R2028 VSS.n1747 VSS.n1746 9.01392
R2029 VSS.n1753 VSS.n1752 9.01392
R2030 VSS.n1757 VSS.n1756 9.01392
R2031 VSS.n1761 VSS.n1760 9.01392
R2032 VSS.n1767 VSS.n1766 9.01392
R2033 VSS.n1771 VSS.n1770 9.01392
R2034 VSS.n1775 VSS.n1774 9.01392
R2035 VSS.n1779 VSS.n1778 9.01392
R2036 VSS.n1785 VSS.n1784 9.01392
R2037 VSS.n1789 VSS.n1788 9.01392
R2038 VSS.n1793 VSS.n1792 9.01392
R2039 VSS.n1797 VSS.n1796 9.01392
R2040 VSS.n1801 VSS.n1800 9.01392
R2041 VSS.n1806 VSS.n1805 9.01392
R2042 VSS.n1810 VSS.n1809 9.01392
R2043 VSS.n1814 VSS.n1813 9.01392
R2044 VSS.n1818 VSS.n1817 9.01392
R2045 VSS.n1824 VSS.n1823 9.01392
R2046 VSS.n1828 VSS.n1827 9.01392
R2047 VSS.n1832 VSS.n1831 9.01392
R2048 VSS.n1836 VSS.n1835 9.01392
R2049 VSS.n1840 VSS.n1839 9.01392
R2050 VSS.n1845 VSS.n1844 9.01392
R2051 VSS.n1854 VSS.n1853 9.01392
R2052 VSS.n1857 VSS.n1856 9.01392
R2053 VSS.n1861 VSS.n1860 9.01392
R2054 VSS.n1867 VSS.n1866 9.01392
R2055 VSS.n1871 VSS.n1870 9.01392
R2056 VSS.n1875 VSS.n1874 9.01392
R2057 VSS.n1881 VSS.n1880 9.01392
R2058 VSS.n1885 VSS.n1884 9.01392
R2059 VSS.n1889 VSS.n1888 9.01392
R2060 VSS.n1893 VSS.n1892 9.01392
R2061 VSS.n1899 VSS.n1898 9.01392
R2062 VSS.n1903 VSS.n1902 9.01392
R2063 VSS.n1907 VSS.n1906 9.01392
R2064 VSS.n1911 VSS.n1910 9.01392
R2065 VSS.n1915 VSS.n1914 9.01392
R2066 VSS.n1920 VSS.n1919 9.01392
R2067 VSS.n1924 VSS.n1923 9.01392
R2068 VSS.n1928 VSS.n1927 9.01392
R2069 VSS.n1932 VSS.n1931 9.01392
R2070 VSS.n1938 VSS.n1937 9.01392
R2071 VSS.n1942 VSS.n1941 9.01392
R2072 VSS.n1946 VSS.n1945 9.01392
R2073 VSS.n1950 VSS.n1949 9.01392
R2074 VSS.n1954 VSS.n1953 9.01392
R2075 VSS.n1959 VSS.n1958 9.01392
R2076 VSS.n1968 VSS.n1967 9.01392
R2077 VSS.n1971 VSS.n1970 9.01392
R2078 VSS.n1975 VSS.n1974 9.01392
R2079 VSS.n1981 VSS.n1980 9.01392
R2080 VSS.n1985 VSS.n1984 9.01392
R2081 VSS.n1989 VSS.n1988 9.01392
R2082 VSS.n1995 VSS.n1994 9.01392
R2083 VSS.n1999 VSS.n1998 9.01392
R2084 VSS.n2003 VSS.n2002 9.01392
R2085 VSS.n2007 VSS.n2006 9.01392
R2086 VSS.n2013 VSS.n2012 9.01392
R2087 VSS.n2017 VSS.n2016 9.01392
R2088 VSS.n2021 VSS.n2020 9.01392
R2089 VSS.n2025 VSS.n2024 9.01392
R2090 VSS.n2029 VSS.n2028 9.01392
R2091 VSS.n2034 VSS.n2033 9.01392
R2092 VSS.n2038 VSS.n2037 9.01392
R2093 VSS.n2042 VSS.n2041 9.01392
R2094 VSS.n2046 VSS.n2045 9.01392
R2095 VSS.n2052 VSS.n2051 9.01392
R2096 VSS.n2056 VSS.n2055 9.01392
R2097 VSS.n2060 VSS.n2059 9.01392
R2098 VSS.n2064 VSS.n2063 9.01392
R2099 VSS.n2068 VSS.n2067 9.01392
R2100 VSS.n2073 VSS.n2072 9.01392
R2101 VSS.n2082 VSS.n2081 9.01392
R2102 VSS.n2085 VSS.n2084 9.01392
R2103 VSS.n2089 VSS.n2088 9.01392
R2104 VSS.n2095 VSS.n2094 9.01392
R2105 VSS.n2099 VSS.n2098 9.01392
R2106 VSS.n2103 VSS.n2102 9.01392
R2107 VSS.n2109 VSS.n2108 9.01392
R2108 VSS.n2113 VSS.n2112 9.01392
R2109 VSS.n2117 VSS.n2116 9.01392
R2110 VSS.n2121 VSS.n2120 9.01392
R2111 VSS.n2127 VSS.n2126 9.01392
R2112 VSS.n2131 VSS.n2130 9.01392
R2113 VSS.n2135 VSS.n2134 9.01392
R2114 VSS.n2139 VSS.n2138 9.01392
R2115 VSS.n2143 VSS.n2142 9.01392
R2116 VSS.n2148 VSS.n2147 9.01392
R2117 VSS.n2152 VSS.n2151 9.01392
R2118 VSS.n2156 VSS.n2155 9.01392
R2119 VSS.n2160 VSS.n2159 9.01392
R2120 VSS.n2166 VSS.n2165 9.01392
R2121 VSS.n2170 VSS.n2169 9.01392
R2122 VSS.n2174 VSS.n2173 9.01392
R2123 VSS.n2178 VSS.n2177 9.01392
R2124 VSS.n2182 VSS.n2181 9.01392
R2125 VSS.n2187 VSS.n2186 9.01392
R2126 VSS.n2191 VSS.n2190 9.01392
R2127 VSS.n2198 VSS.n2197 9.01392
R2128 VSS VSS.n2198 9.01392
R2129 VSS.n550 VSS.n549 9.01392
R2130 VSS.n548 VSS.n547 9.01392
R2131 VSS.n542 VSS.n541 9.01392
R2132 VSS.n538 VSS.n537 9.01392
R2133 VSS.n534 VSS.n533 9.01392
R2134 VSS.n527 VSS.n526 9.01392
R2135 VSS.n231 VSS.n230 9.01392
R2136 VSS.n522 VSS.n521 9.01392
R2137 VSS.n518 VSS.n517 9.01392
R2138 VSS.n512 VSS.n511 9.01392
R2139 VSS.n507 VSS.n506 9.01392
R2140 VSS.n236 VSS.n235 9.01392
R2141 VSS.n502 VSS.n501 9.01392
R2142 VSS.n498 VSS.n497 9.01392
R2143 VSS.n491 VSS.n490 9.01392
R2144 VSS.n487 VSS.n486 9.01392
R2145 VSS.n480 VSS.n479 9.01392
R2146 VSS.n482 VSS.n481 9.01392
R2147 VSS.n400 VSS.n399 9.01392
R2148 VSS.n247 VSS.n246 9.01392
R2149 VSS.n395 VSS.n394 9.01392
R2150 VSS.n391 VSS.n390 9.01392
R2151 VSS.n384 VSS.n383 9.01392
R2152 VSS.n380 VSS.n379 9.01392
R2153 VSS.n373 VSS.n372 9.01392
R2154 VSS.n375 VSS.n374 9.01392
R2155 VSS.n293 VSS.n292 9.01392
R2156 VSS.n258 VSS.n257 9.01392
R2157 VSS.n288 VSS.n287 9.01392
R2158 VSS.n284 VSS.n283 9.01392
R2159 VSS.n277 VSS.n276 9.01392
R2160 VSS.n273 VSS.n272 9.01392
R2161 VSS.n266 VSS.n265 9.01392
R2162 VSS.n269 VSS.n268 9.01392
R2163 VSS.n268 VSS.n267 9.01392
R2164 VSS.n299 VSS.n298 9.01392
R2165 VSS.n298 VSS.n297 9.01392
R2166 VSS.n406 VSS.n405 9.01392
R2167 VSS.n405 VSS.n404 9.01392
R2168 VSS.n2895 VSS.n2894 9.01392
R2169 VSS.n2883 VSS.n2882 9.01392
R2170 VSS.n1289 VSS.n1288 9.01392
R2171 VSS.n2878 VSS.n2877 9.01392
R2172 VSS.n2874 VSS.n2873 9.01392
R2173 VSS.n2870 VSS.n2869 9.01392
R2174 VSS.n2866 VSS.n2865 9.01392
R2175 VSS.n2860 VSS.n2859 9.01392
R2176 VSS.n2856 VSS.n2855 9.01392
R2177 VSS.n2852 VSS.n2851 9.01392
R2178 VSS.n2848 VSS.n2847 9.01392
R2179 VSS.n2843 VSS.n2842 9.01392
R2180 VSS.n2839 VSS.n2838 9.01392
R2181 VSS.n2835 VSS.n2834 9.01392
R2182 VSS.n2831 VSS.n2830 9.01392
R2183 VSS.n2827 VSS.n2826 9.01392
R2184 VSS.n2821 VSS.n2820 9.01392
R2185 VSS.n2817 VSS.n2816 9.01392
R2186 VSS.n2813 VSS.n2812 9.01392
R2187 VSS.n2809 VSS.n2808 9.01392
R2188 VSS.n1293 VSS.n1292 9.01392
R2189 VSS.n2804 VSS.n2803 9.01392
R2190 VSS.n2800 VSS.n2799 9.01392
R2191 VSS.n1298 VSS.n1297 9.01392
R2192 VSS.n2795 VSS.n2794 9.01392
R2193 VSS.n2792 VSS.n2791 9.01392
R2194 VSS.n2784 VSS.n2783 9.01392
R2195 VSS.n1305 VSS.n1304 9.01392
R2196 VSS.n2779 VSS.n2778 9.01392
R2197 VSS.n2775 VSS.n2774 9.01392
R2198 VSS.n2771 VSS.n2770 9.01392
R2199 VSS.n2767 VSS.n2766 9.01392
R2200 VSS.n2761 VSS.n2760 9.01392
R2201 VSS.n2757 VSS.n2756 9.01392
R2202 VSS.n2753 VSS.n2752 9.01392
R2203 VSS.n2749 VSS.n2748 9.01392
R2204 VSS.n2744 VSS.n2743 9.01392
R2205 VSS.n2740 VSS.n2739 9.01392
R2206 VSS.n2736 VSS.n2735 9.01392
R2207 VSS.n2732 VSS.n2731 9.01392
R2208 VSS.n2728 VSS.n2727 9.01392
R2209 VSS.n2722 VSS.n2721 9.01392
R2210 VSS.n2718 VSS.n2717 9.01392
R2211 VSS.n2714 VSS.n2713 9.01392
R2212 VSS.n2710 VSS.n2709 9.01392
R2213 VSS.n1309 VSS.n1308 9.01392
R2214 VSS.n2705 VSS.n2704 9.01392
R2215 VSS.n2701 VSS.n2700 9.01392
R2216 VSS.n1314 VSS.n1313 9.01392
R2217 VSS.n2696 VSS.n2695 9.01392
R2218 VSS.n2693 VSS.n2692 9.01392
R2219 VSS.n2685 VSS.n2684 9.01392
R2220 VSS.n1321 VSS.n1320 9.01392
R2221 VSS.n2680 VSS.n2679 9.01392
R2222 VSS.n2676 VSS.n2675 9.01392
R2223 VSS.n2672 VSS.n2671 9.01392
R2224 VSS.n2668 VSS.n2667 9.01392
R2225 VSS.n2662 VSS.n2661 9.01392
R2226 VSS.n2658 VSS.n2657 9.01392
R2227 VSS.n2654 VSS.n2653 9.01392
R2228 VSS.n2650 VSS.n2649 9.01392
R2229 VSS.n2645 VSS.n2644 9.01392
R2230 VSS.n2641 VSS.n2640 9.01392
R2231 VSS.n2637 VSS.n2636 9.01392
R2232 VSS.n2633 VSS.n2632 9.01392
R2233 VSS.n2629 VSS.n2628 9.01392
R2234 VSS.n2623 VSS.n2622 9.01392
R2235 VSS.n2619 VSS.n2618 9.01392
R2236 VSS.n2615 VSS.n2614 9.01392
R2237 VSS.n2611 VSS.n2610 9.01392
R2238 VSS.n1325 VSS.n1324 9.01392
R2239 VSS.n2606 VSS.n2605 9.01392
R2240 VSS.n2602 VSS.n2601 9.01392
R2241 VSS.n1330 VSS.n1329 9.01392
R2242 VSS.n2597 VSS.n2596 9.01392
R2243 VSS.n2594 VSS.n2593 9.01392
R2244 VSS.n2586 VSS.n2585 9.01392
R2245 VSS.n1337 VSS.n1336 9.01392
R2246 VSS.n2581 VSS.n2580 9.01392
R2247 VSS.n2577 VSS.n2576 9.01392
R2248 VSS.n2573 VSS.n2572 9.01392
R2249 VSS.n2569 VSS.n2568 9.01392
R2250 VSS.n2563 VSS.n2562 9.01392
R2251 VSS.n2559 VSS.n2558 9.01392
R2252 VSS.n2555 VSS.n2554 9.01392
R2253 VSS.n2551 VSS.n2550 9.01392
R2254 VSS.n2546 VSS.n2545 9.01392
R2255 VSS.n2542 VSS.n2541 9.01392
R2256 VSS.n2538 VSS.n2537 9.01392
R2257 VSS.n2534 VSS.n2533 9.01392
R2258 VSS.n2530 VSS.n2529 9.01392
R2259 VSS.n2524 VSS.n2523 9.01392
R2260 VSS.n2520 VSS.n2519 9.01392
R2261 VSS.n2516 VSS.n2515 9.01392
R2262 VSS.n2512 VSS.n2511 9.01392
R2263 VSS.n1341 VSS.n1340 9.01392
R2264 VSS.n2507 VSS.n2506 9.01392
R2265 VSS.n2503 VSS.n2502 9.01392
R2266 VSS.n1346 VSS.n1345 9.01392
R2267 VSS.n2498 VSS.n2497 9.01392
R2268 VSS.n2495 VSS.n2494 9.01392
R2269 VSS.n2487 VSS.n2486 9.01392
R2270 VSS.n1353 VSS.n1352 9.01392
R2271 VSS.n2482 VSS.n2481 9.01392
R2272 VSS.n2478 VSS.n2477 9.01392
R2273 VSS.n2474 VSS.n2473 9.01392
R2274 VSS.n2470 VSS.n2469 9.01392
R2275 VSS.n2464 VSS.n2463 9.01392
R2276 VSS.n2460 VSS.n2459 9.01392
R2277 VSS.n2456 VSS.n2455 9.01392
R2278 VSS.n2452 VSS.n2451 9.01392
R2279 VSS.n2447 VSS.n2446 9.01392
R2280 VSS.n2443 VSS.n2442 9.01392
R2281 VSS.n2439 VSS.n2438 9.01392
R2282 VSS.n2435 VSS.n2434 9.01392
R2283 VSS.n2431 VSS.n2430 9.01392
R2284 VSS.n2425 VSS.n2424 9.01392
R2285 VSS.n2421 VSS.n2420 9.01392
R2286 VSS.n2417 VSS.n2416 9.01392
R2287 VSS.n2413 VSS.n2412 9.01392
R2288 VSS.n1357 VSS.n1356 9.01392
R2289 VSS.n2408 VSS.n2407 9.01392
R2290 VSS.n2404 VSS.n2403 9.01392
R2291 VSS.n1362 VSS.n1361 9.01392
R2292 VSS.n2399 VSS.n2398 9.01392
R2293 VSS.n2396 VSS.n2395 9.01392
R2294 VSS.n2388 VSS.n2387 9.01392
R2295 VSS.n1369 VSS.n1368 9.01392
R2296 VSS.n2383 VSS.n2382 9.01392
R2297 VSS.n2379 VSS.n2378 9.01392
R2298 VSS.n2375 VSS.n2374 9.01392
R2299 VSS.n2371 VSS.n2370 9.01392
R2300 VSS.n2365 VSS.n2364 9.01392
R2301 VSS.n2361 VSS.n2360 9.01392
R2302 VSS.n2357 VSS.n2356 9.01392
R2303 VSS.n2353 VSS.n2352 9.01392
R2304 VSS.n2348 VSS.n2347 9.01392
R2305 VSS.n2344 VSS.n2343 9.01392
R2306 VSS.n2340 VSS.n2339 9.01392
R2307 VSS.n2336 VSS.n2335 9.01392
R2308 VSS.n2332 VSS.n2331 9.01392
R2309 VSS.n2326 VSS.n2325 9.01392
R2310 VSS.n2322 VSS.n2321 9.01392
R2311 VSS.n2318 VSS.n2317 9.01392
R2312 VSS.n2314 VSS.n2313 9.01392
R2313 VSS.n1373 VSS.n1372 9.01392
R2314 VSS.n2309 VSS.n2308 9.01392
R2315 VSS.n2305 VSS.n2304 9.01392
R2316 VSS.n1378 VSS.n1377 9.01392
R2317 VSS.n2300 VSS.n2299 9.01392
R2318 VSS.n2297 VSS.n2296 9.01392
R2319 VSS.n2289 VSS.n2288 9.01392
R2320 VSS.n1385 VSS.n1384 9.01392
R2321 VSS.n2284 VSS.n2283 9.01392
R2322 VSS.n2280 VSS.n2279 9.01392
R2323 VSS.n2276 VSS.n2275 9.01392
R2324 VSS.n2272 VSS.n2271 9.01392
R2325 VSS.n2266 VSS.n2265 9.01392
R2326 VSS.n2262 VSS.n2261 9.01392
R2327 VSS.n2258 VSS.n2257 9.01392
R2328 VSS.n2254 VSS.n2253 9.01392
R2329 VSS.n2249 VSS.n2248 9.01392
R2330 VSS.n2245 VSS.n2244 9.01392
R2331 VSS.n2241 VSS.n2240 9.01392
R2332 VSS.n2237 VSS.n2236 9.01392
R2333 VSS.n2233 VSS.n2232 9.01392
R2334 VSS.n2227 VSS.n2226 9.01392
R2335 VSS.n2223 VSS.n2222 9.01392
R2336 VSS.n2219 VSS.n2218 9.01392
R2337 VSS.n2215 VSS.n2214 9.01392
R2338 VSS.n1389 VSS.n1388 9.01392
R2339 VSS.n2210 VSS.n2209 9.01392
R2340 VSS.n2206 VSS.n2205 9.01392
R2341 VSS.n1394 VSS.n1393 9.01392
R2342 VSS.n2202 VSS.n2201 9.01392
R2343 VSS.n2201 VSS.n2200 9.01392
R2344 VSS.n3058 VSS.n3057 9.01392
R2345 VSS.n3059 VSS.n3058 9.01392
R2346 VSS.n3062 VSS.n3061 9.01392
R2347 VSS.n3061 VSS.n3060 9.01392
R2348 VSS.n3068 VSS.n3065 9.01392
R2349 VSS.n3065 VSS.n3064 9.01392
R2350 VSS.n3072 VSS.n3071 9.01392
R2351 VSS.n3071 VSS.n3070 9.01392
R2352 VSS.n3075 VSS.n3074 9.01392
R2353 VSS.n3082 VSS.n3081 9.01392
R2354 VSS.n3081 VSS.n3080 9.01392
R2355 VSS.n3086 VSS.n3085 9.01392
R2356 VSS.n3087 VSS.n3086 9.01392
R2357 VSS.n3090 VSS.n3089 9.01392
R2358 VSS.n3089 VSS.n3088 9.01392
R2359 VSS.n3094 VSS.n3093 9.01392
R2360 VSS.n3093 VSS.n3092 9.01392
R2361 VSS.n3100 VSS.n3099 9.01392
R2362 VSS.n3099 VSS.n3098 9.01392
R2363 VSS.n3104 VSS.n3103 9.01392
R2364 VSS.n3103 VSS.n3102 9.01392
R2365 VSS.n3110 VSS.n3109 9.01392
R2366 VSS.n3109 VSS.n3108 9.01392
R2367 VSS.n3114 VSS.n3113 9.01392
R2368 VSS.n3113 VSS.n3112 9.01392
R2369 VSS.n3119 VSS.n3118 9.01392
R2370 VSS.n3125 VSS.n3124 9.01392
R2371 VSS.n3124 VSS.n3123 9.01392
R2372 VSS.n3129 VSS.n3128 9.01392
R2373 VSS.n3128 VSS.n3127 9.01392
R2374 VSS.n3135 VSS.n3134 9.01392
R2375 VSS.n3134 VSS.n3133 9.01392
R2376 VSS.n3139 VSS.n3138 9.01392
R2377 VSS.n3138 VSS.n3137 9.01392
R2378 VSS.n3145 VSS.n3144 9.01392
R2379 VSS.n3144 VSS.n3143 9.01392
R2380 VSS.n3149 VSS.n3148 9.01392
R2381 VSS.n3148 VSS.n3147 9.01392
R2382 VSS.n3155 VSS.n3152 9.01392
R2383 VSS.n3152 VSS.n3151 9.01392
R2384 VSS.n3159 VSS.n3158 9.01392
R2385 VSS.n3158 VSS.n3157 9.01392
R2386 VSS.n3165 VSS.n3162 9.01392
R2387 VSS.n3162 VSS.n3161 9.01392
R2388 VSS.n3171 VSS.n3170 9.01392
R2389 VSS.n3170 VSS.n3169 9.01392
R2390 VSS.n3175 VSS.n3174 9.01392
R2391 VSS.n3174 VSS.n3173 9.01392
R2392 VSS.n3181 VSS.n3180 9.01392
R2393 VSS.n3180 VSS.n3179 9.01392
R2394 VSS.n3185 VSS.n3184 9.01392
R2395 VSS.n3184 VSS.n3183 9.01392
R2396 VSS.n3190 VSS.n3189 9.01392
R2397 VSS.n3189 VSS.n3188 9.01392
R2398 VSS.n3045 VSS.n3044 9.01392
R2399 VSS.n3042 VSS.n3041 9.01392
R2400 VSS.n3041 VSS.n3040 9.01392
R2401 VSS.n3038 VSS.n3037 9.01392
R2402 VSS.n3039 VSS.n3038 9.01392
R2403 VSS.n3034 VSS.n3031 9.01392
R2404 VSS.n3031 VSS.n3030 9.01392
R2405 VSS.n3028 VSS.n3027 9.01392
R2406 VSS.n3027 VSS.n3026 9.01392
R2407 VSS.n3021 VSS.n3020 9.01392
R2408 VSS.n3015 VSS.n3014 9.01392
R2409 VSS.n3014 VSS.n3013 9.01392
R2410 VSS.n3017 VSS.n3012 9.01392
R2411 VSS.n3012 VSS.n3011 9.01392
R2412 VSS.n3009 VSS.n3008 9.01392
R2413 VSS.n3010 VSS.n3009 9.01392
R2414 VSS.n3005 VSS.n3004 9.01392
R2415 VSS.n3004 VSS.n3003 9.01392
R2416 VSS.n3001 VSS.n3000 9.01392
R2417 VSS.n3000 VSS.n2999 9.01392
R2418 VSS.n2995 VSS.n2994 9.01392
R2419 VSS.n2994 VSS.n2993 9.01392
R2420 VSS.n2991 VSS.n2990 9.01392
R2421 VSS.n2990 VSS.n2989 9.01392
R2422 VSS.n2985 VSS.n2984 9.01392
R2423 VSS.n2984 VSS.n2983 9.01392
R2424 VSS.n2981 VSS.n2980 9.01392
R2425 VSS.n2980 VSS.t233 9.01392
R2426 VSS.n2976 VSS.n2975 9.01392
R2427 VSS.n2975 VSS.n2974 9.01392
R2428 VSS.n2970 VSS.n2969 9.01392
R2429 VSS.n2969 VSS.n2968 9.01392
R2430 VSS.n2966 VSS.n2965 9.01392
R2431 VSS.n2965 VSS.n2964 9.01392
R2432 VSS.n2960 VSS.n2959 9.01392
R2433 VSS.n2959 VSS.n2958 9.01392
R2434 VSS.n2956 VSS.n2955 9.01392
R2435 VSS.n2955 VSS.n2954 9.01392
R2436 VSS.n2950 VSS.n2949 9.01392
R2437 VSS.n2949 VSS.n2948 9.01392
R2438 VSS.n2946 VSS.n2943 9.01392
R2439 VSS.n2943 VSS.n2942 9.01392
R2440 VSS.n2940 VSS.n2939 9.01392
R2441 VSS.n2939 VSS.n2938 9.01392
R2442 VSS.n2936 VSS.n2933 9.01392
R2443 VSS.n2933 VSS.n2932 9.01392
R2444 VSS.n2930 VSS.n2929 9.01392
R2445 VSS.n2929 VSS.n2928 9.01392
R2446 VSS.n2926 VSS.n2923 9.01392
R2447 VSS.n2923 VSS.n2922 9.01392
R2448 VSS.n2920 VSS.n2919 9.01392
R2449 VSS.n2919 VSS.n2918 9.01392
R2450 VSS.n2914 VSS.n2913 9.01392
R2451 VSS.n2913 VSS.n2912 9.01392
R2452 VSS.n2910 VSS.n2909 9.01392
R2453 VSS.n2909 VSS.n2908 9.01392
R2454 VSS.n2905 VSS.n2904 9.01392
R2455 VSS.n2904 VSS.n2903 9.01392
R2456 VSS.n3195 VSS.n3194 9.01392
R2457 VSS.n204 VSS.n202 8.84842
R2458 VSS.n162 VSS.n160 8.84842
R2459 VSS.n756 VSS.n178 8.82809
R2460 VSS.n742 VSS.n741 8.82809
R2461 VSS.n737 VSS.n736 8.82809
R2462 VSS.n729 VSS.n728 8.82809
R2463 VSS.n715 VSS.n184 8.82809
R2464 VSS.n596 VSS.n220 8.82809
R2465 VSS.n582 VSS.n581 8.82809
R2466 VSS.n577 VSS.n576 8.82809
R2467 VSS.n569 VSS.n568 8.82809
R2468 VSS.n555 VSS.n226 8.82809
R2469 VSS.n162 VSS.n147 8.6074
R2470 VSS.n204 VSS.n189 8.6074
R2471 VSS.n474 VSS.n471 8.38671
R2472 VSS.n457 VSS.n456 8.38671
R2473 VSS.n452 VSS.n448 8.38671
R2474 VSS.n444 VSS.n443 8.38671
R2475 VSS.n428 VSS.n245 8.38671
R2476 VSS.n367 VSS.n364 8.38671
R2477 VSS.n350 VSS.n349 8.38671
R2478 VSS.n345 VSS.n341 8.38671
R2479 VSS.n337 VSS.n336 8.38671
R2480 VSS.n321 VSS.n256 8.38671
R2481 VSS.n3125 VSS.n3122 7.50395
R2482 VSS.n2976 VSS.n2973 7.50395
R2483 VSS.n54 VSS.n53 7.45124
R2484 VSS.n121 VSS.n120 7.45124
R2485 VSS.n95 VSS.n93 7.01423
R2486 VSS.n106 VSS.n105 7.00892
R2487 VSS.n39 VSS.n38 6.90643
R2488 VSS.n3181 VSS.n3178 6.62119
R2489 VSS.n3165 VSS.n3164 6.62119
R2490 VSS.n2920 VSS.n2917 6.62119
R2491 VSS.n2936 VSS.n2935 6.62119
R2492 VSS.n912 VSS 5.81868
R2493 VSS.n1123 VSS 5.81868
R2494 VSS.n1241 VSS 5.81868
R2495 VSS.n1031 VSS 5.81868
R2496 VSS.n824 VSS 5.81868
R2497 VSS.n732 VSS 5.81868
R2498 VSS.n664 VSS 5.81868
R2499 VSS.n572 VSS 5.81868
R2500 VSS.n531 VSS 5.81868
R2501 VSS.n495 VSS 5.81868
R2502 VSS.n450 VSS 5.81868
R2503 VSS.n388 VSS 5.81868
R2504 VSS.n343 VSS 5.81868
R2505 VSS.n281 VSS 5.81868
R2506 VSS.n150 VSS.n149 5.79462
R2507 VSS.n860 VSS.n856 5.79462
R2508 VSS.n847 VSS.n843 5.79462
R2509 VSS.n833 VSS.n829 5.79462
R2510 VSS.n816 VSS.n812 5.79462
R2511 VSS.n171 VSS.n167 5.79462
R2512 VSS.n799 VSS.n795 5.79462
R2513 VSS.n785 VSS.n781 5.79462
R2514 VSS.n192 VSS.n191 5.79462
R2515 VSS.n700 VSS.n696 5.79462
R2516 VSS.n687 VSS.n683 5.79462
R2517 VSS.n673 VSS.n669 5.79462
R2518 VSS.n656 VSS.n652 5.79462
R2519 VSS.n213 VSS.n209 5.79462
R2520 VSS.n639 VSS.n635 5.79462
R2521 VSS.n625 VSS.n621 5.79462
R2522 VSS.n16 VSS.n15 5.79462
R2523 VSS.n13 VSS.n12 5.79462
R2524 VSS.n1274 VSS.n1273 5.79462
R2525 VSS.n1260 VSS.n1259 5.79462
R2526 VSS.n1245 VSS.n1244 5.79462
R2527 VSS.n1229 VSS.n1228 5.79462
R2528 VSS.n37 VSS.n36 5.79462
R2529 VSS.n1214 VSS.n1213 5.79462
R2530 VSS.n1200 VSS.n1199 5.79462
R2531 VSS.n3110 VSS.n3107 5.73843
R2532 VSS.n2991 VSS.n2988 5.73843
R2533 VSS.n95 VSS.n80 5.51774
R2534 VSS.n3016 VSS.n3015 5.51774
R2535 VSS.n160 VSS.n159 5.51315
R2536 VSS.n202 VSS.n201 5.51315
R2537 VSS.n27 VSS.n26 5.29705
R2538 VSS.n106 VSS.n98 5.07636
R2539 VSS.n467 VSS.n466 5.07636
R2540 VSS.n360 VSS.n359 5.07636
R2541 VSS.n39 VSS.n31 4.85567
R2542 VSS.n1281 VSS.n1280 4.6505
R2543 VSS.n1253 VSS.n1252 4.6505
R2544 VSS.n1207 VSS.n1206 4.6505
R2545 VSS.n1169 VSS.n1168 4.6505
R2546 VSS.n1165 VSS.n1164 4.6505
R2547 VSS.n1149 VSS.n1148 4.6505
R2548 VSS.n1135 VSS.n1134 4.6505
R2549 VSS.n1119 VSS.n1118 4.6505
R2550 VSS.n1105 VSS.n1104 4.6505
R2551 VSS.n1088 VSS.n1087 4.6505
R2552 VSS.n1078 VSS.n1077 4.6505
R2553 VSS.n1071 VSS.n1070 4.6505
R2554 VSS.n1043 VSS.n1042 4.6505
R2555 VSS.n996 VSS.n995 4.6505
R2556 VSS.n958 VSS.n957 4.6505
R2557 VSS.n954 VSS.n953 4.6505
R2558 VSS.n938 VSS.n937 4.6505
R2559 VSS.n924 VSS.n923 4.6505
R2560 VSS.n908 VSS.n907 4.6505
R2561 VSS.n894 VSS.n893 4.6505
R2562 VSS.n877 VSS.n876 4.6505
R2563 VSS.n870 VSS.n869 4.6505
R2564 VSS.n863 VSS.n862 4.6505
R2565 VSS.n850 VSS.n849 4.6505
R2566 VSS.n836 VSS.n835 4.6505
R2567 VSS.n819 VSS.n818 4.6505
R2568 VSS.n802 VSS.n801 4.6505
R2569 VSS.n788 VSS.n787 4.6505
R2570 VSS.n752 VSS.n751 4.6505
R2571 VSS.n738 VSS.n737 4.6505
R2572 VSS.n725 VSS.n724 4.6505
R2573 VSS.n184 VSS.n179 4.6505
R2574 VSS.n710 VSS.n709 4.6505
R2575 VSS.n703 VSS.n702 4.6505
R2576 VSS.n690 VSS.n689 4.6505
R2577 VSS.n676 VSS.n675 4.6505
R2578 VSS.n659 VSS.n658 4.6505
R2579 VSS.n642 VSS.n641 4.6505
R2580 VSS.n628 VSS.n627 4.6505
R2581 VSS.n592 VSS.n591 4.6505
R2582 VSS.n578 VSS.n577 4.6505
R2583 VSS.n565 VSS.n564 4.6505
R2584 VSS.n226 VSS.n221 4.6505
R2585 VSS.n471 VSS.n470 4.6505
R2586 VSS.n460 VSS.n459 4.6505
R2587 VSS.n453 VSS.n452 4.6505
R2588 VSS.n440 VSS.n439 4.6505
R2589 VSS.n429 VSS.n428 4.6505
R2590 VSS.n364 VSS.n363 4.6505
R2591 VSS.n353 VSS.n352 4.6505
R2592 VSS.n346 VSS.n345 4.6505
R2593 VSS.n333 VSS.n332 4.6505
R2594 VSS.n322 VSS.n321 4.6505
R2595 VSS.n324 VSS.n323 4.6505
R2596 VSS.n338 VSS.n337 4.6505
R2597 VSS.n351 VSS.n350 4.6505
R2598 VSS.n362 VSS.n361 4.6505
R2599 VSS.n431 VSS.n430 4.6505
R2600 VSS.n445 VSS.n444 4.6505
R2601 VSS.n458 VSS.n457 4.6505
R2602 VSS.n469 VSS.n468 4.6505
R2603 VSS.n563 VSS.n562 4.6505
R2604 VSS.n570 VSS.n569 4.6505
R2605 VSS.n583 VSS.n582 4.6505
R2606 VSS.n594 VSS.n593 4.6505
R2607 VSS.n596 VSS.n595 4.6505
R2608 VSS.n723 VSS.n722 4.6505
R2609 VSS.n730 VSS.n729 4.6505
R2610 VSS.n743 VSS.n742 4.6505
R2611 VSS.n754 VSS.n753 4.6505
R2612 VSS.n756 VSS.n755 4.6505
R2613 VSS.n1010 VSS.n1009 4.6505
R2614 VSS.n1026 VSS.n1025 4.6505
R2615 VSS.n1057 VSS.n1056 4.6505
R2616 VSS.n1221 VSS.n1220 4.6505
R2617 VSS.n1236 VSS.n1235 4.6505
R2618 VSS.n1267 VSS.n1266 4.6505
R2619 VSS.n721 VSS.n183 4.63498
R2620 VSS.n561 VSS.n225 4.63498
R2621 VSS.n645 VSS.n215 4.49926
R2622 VSS.n805 VSS.n173 4.49926
R2623 VSS.n941 VSS.n122 4.49926
R2624 VSS.n1013 VSS.n107 4.49926
R2625 VSS.n1152 VSS.n55 4.49926
R2626 VSS.n1224 VSS.n40 4.49926
R2627 VSS.n706 VSS.n205 4.42059
R2628 VSS.n866 VSS.n163 4.42059
R2629 VSS.n880 VSS.n124 4.42059
R2630 VSS.n1074 VSS.n96 4.42059
R2631 VSS.n1091 VSS.n57 4.42059
R2632 VSS.n1284 VSS.n28 4.42059
R2633 VSS.n3135 VSS.n3132 3.97291
R2634 VSS.n2966 VSS.n2963 3.97291
R2635 VSS.n1286 VSS.n8 3.87498
R2636 VSS.n3062 VSS 3.53153
R2637 VSS.n1280 VSS.n1279 3.53153
R2638 VSS.n1279 VSS.n1272 3.53153
R2639 VSS.n1266 VSS.n1265 3.53153
R2640 VSS.n1265 VSS.n1258 3.53153
R2641 VSS.n1250 VSS.n1243 3.53153
R2642 VSS.n1235 VSS.n1234 3.53153
R2643 VSS.n1220 VSS.n1219 3.53153
R2644 VSS.n1219 VSS.n1212 3.53153
R2645 VSS.n1206 VSS.n1205 3.53153
R2646 VSS.n1205 VSS.n1198 3.53153
R2647 VSS.n871 VSS.n870 3.53153
R2648 VSS.n147 VSS.n146 3.53153
R2649 VSS.n854 VSS.n853 3.53153
R2650 VSS.n849 VSS.n839 3.53153
R2651 VSS.n841 VSS.n840 3.53153
R2652 VSS.n835 VSS.n822 3.53153
R2653 VSS.n818 VSS.n808 3.53153
R2654 VSS.n810 VSS.n809 3.53153
R2655 VSS.n801 VSS.n791 3.53153
R2656 VSS.n793 VSS.n792 3.53153
R2657 VSS.n787 VSS.n175 3.53153
R2658 VSS.n779 VSS.n778 3.53153
R2659 VSS.n711 VSS.n710 3.53153
R2660 VSS.n189 VSS.n188 3.53153
R2661 VSS.n694 VSS.n693 3.53153
R2662 VSS.n689 VSS.n679 3.53153
R2663 VSS.n681 VSS.n680 3.53153
R2664 VSS.n675 VSS.n662 3.53153
R2665 VSS.n658 VSS.n648 3.53153
R2666 VSS.n650 VSS.n649 3.53153
R2667 VSS.n641 VSS.n631 3.53153
R2668 VSS.n633 VSS.n632 3.53153
R2669 VSS.n627 VSS.n217 3.53153
R2670 VSS.n619 VSS.n618 3.53153
R2671 VSS.n25 VSS.n8 3.53153
R2672 VSS.n3037 VSS 3.53153
R2673 VSS.n1078 VSS.n76 3.31084
R2674 VSS.n79 VSS.n76 3.31084
R2675 VSS.n1070 VSS.n1069 3.31084
R2676 VSS.n1069 VSS.n1062 3.31084
R2677 VSS.n1056 VSS.n1055 3.31084
R2678 VSS.n1055 VSS.n1048 3.31084
R2679 VSS.n1040 VSS.n1033 3.31084
R2680 VSS.n1025 VSS.n1024 3.31084
R2681 VSS.n1024 VSS.n1017 3.31084
R2682 VSS.n1009 VSS.n1008 3.31084
R2683 VSS.n1008 VSS.n1001 3.31084
R2684 VSS.n995 VSS.n994 3.31084
R2685 VSS.n994 VSS.n987 3.31084
R2686 VSS.n3052 VSS 3.31084
R2687 VSS.n3201 VSS 3.31084
R2688 VSS.n2203 VSS.n2202 3.1005
R2689 VSS.n2898 VSS.n2897 3.1005
R2690 VSS.n2197 VSS.n2196 3.1005
R2691 VSS.n2890 VSS.n1287 3.1005
R2692 VSS.n1413 VSS.n1412 3.1005
R2693 VSS.n1417 VSS.n1416 3.1005
R2694 VSS.n1427 VSS.n1426 3.1005
R2695 VSS.n1431 VSS.n1430 3.1005
R2696 VSS.n1435 VSS.n1434 3.1005
R2697 VSS.n1439 VSS.n1438 3.1005
R2698 VSS.n1445 VSS.n1444 3.1005
R2699 VSS.n1449 VSS.n1448 3.1005
R2700 VSS.n1453 VSS.n1452 3.1005
R2701 VSS.n1457 VSS.n1456 3.1005
R2702 VSS.n1461 VSS.n1460 3.1005
R2703 VSS.n1466 VSS.n1465 3.1005
R2704 VSS.n1470 VSS.n1469 3.1005
R2705 VSS.n1474 VSS.n1473 3.1005
R2706 VSS.n1478 VSS.n1477 3.1005
R2707 VSS.n1484 VSS.n1483 3.1005
R2708 VSS.n1488 VSS.n1487 3.1005
R2709 VSS.n1492 VSS.n1491 3.1005
R2710 VSS.n1496 VSS.n1495 3.1005
R2711 VSS.n1505 VSS.n1504 3.1005
R2712 VSS.n1506 VSS.n1403 3.1005
R2713 VSS.n1517 VSS.n1516 3.1005
R2714 VSS.n1527 VSS.n1526 3.1005
R2715 VSS.n1531 VSS.n1530 3.1005
R2716 VSS.n1541 VSS.n1540 3.1005
R2717 VSS.n1545 VSS.n1544 3.1005
R2718 VSS.n1549 VSS.n1548 3.1005
R2719 VSS.n1553 VSS.n1552 3.1005
R2720 VSS.n1559 VSS.n1558 3.1005
R2721 VSS.n1563 VSS.n1562 3.1005
R2722 VSS.n1567 VSS.n1566 3.1005
R2723 VSS.n1571 VSS.n1570 3.1005
R2724 VSS.n1575 VSS.n1574 3.1005
R2725 VSS.n1580 VSS.n1579 3.1005
R2726 VSS.n1584 VSS.n1583 3.1005
R2727 VSS.n1588 VSS.n1587 3.1005
R2728 VSS.n1592 VSS.n1591 3.1005
R2729 VSS.n1598 VSS.n1597 3.1005
R2730 VSS.n1602 VSS.n1601 3.1005
R2731 VSS.n1606 VSS.n1605 3.1005
R2732 VSS.n1610 VSS.n1609 3.1005
R2733 VSS.n1619 VSS.n1618 3.1005
R2734 VSS.n1620 VSS.n1402 3.1005
R2735 VSS.n1631 VSS.n1630 3.1005
R2736 VSS.n1641 VSS.n1640 3.1005
R2737 VSS.n1645 VSS.n1644 3.1005
R2738 VSS.n1655 VSS.n1654 3.1005
R2739 VSS.n1659 VSS.n1658 3.1005
R2740 VSS.n1663 VSS.n1662 3.1005
R2741 VSS.n1667 VSS.n1666 3.1005
R2742 VSS.n1673 VSS.n1672 3.1005
R2743 VSS.n1677 VSS.n1676 3.1005
R2744 VSS.n1681 VSS.n1680 3.1005
R2745 VSS.n1685 VSS.n1684 3.1005
R2746 VSS.n1689 VSS.n1688 3.1005
R2747 VSS.n1694 VSS.n1693 3.1005
R2748 VSS.n1698 VSS.n1697 3.1005
R2749 VSS.n1702 VSS.n1701 3.1005
R2750 VSS.n1706 VSS.n1705 3.1005
R2751 VSS.n1712 VSS.n1711 3.1005
R2752 VSS.n1716 VSS.n1715 3.1005
R2753 VSS.n1720 VSS.n1719 3.1005
R2754 VSS.n1724 VSS.n1723 3.1005
R2755 VSS.n1733 VSS.n1732 3.1005
R2756 VSS.n1734 VSS.n1401 3.1005
R2757 VSS.n1745 VSS.n1744 3.1005
R2758 VSS.n1755 VSS.n1754 3.1005
R2759 VSS.n1759 VSS.n1758 3.1005
R2760 VSS.n1769 VSS.n1768 3.1005
R2761 VSS.n1773 VSS.n1772 3.1005
R2762 VSS.n1777 VSS.n1776 3.1005
R2763 VSS.n1781 VSS.n1780 3.1005
R2764 VSS.n1787 VSS.n1786 3.1005
R2765 VSS.n1791 VSS.n1790 3.1005
R2766 VSS.n1795 VSS.n1794 3.1005
R2767 VSS.n1799 VSS.n1798 3.1005
R2768 VSS.n1803 VSS.n1802 3.1005
R2769 VSS.n1808 VSS.n1807 3.1005
R2770 VSS.n1812 VSS.n1811 3.1005
R2771 VSS.n1816 VSS.n1815 3.1005
R2772 VSS.n1820 VSS.n1819 3.1005
R2773 VSS.n1826 VSS.n1825 3.1005
R2774 VSS.n1830 VSS.n1829 3.1005
R2775 VSS.n1834 VSS.n1833 3.1005
R2776 VSS.n1838 VSS.n1837 3.1005
R2777 VSS.n1847 VSS.n1846 3.1005
R2778 VSS.n1848 VSS.n1400 3.1005
R2779 VSS.n1859 VSS.n1858 3.1005
R2780 VSS.n1869 VSS.n1868 3.1005
R2781 VSS.n1873 VSS.n1872 3.1005
R2782 VSS.n1883 VSS.n1882 3.1005
R2783 VSS.n1887 VSS.n1886 3.1005
R2784 VSS.n1891 VSS.n1890 3.1005
R2785 VSS.n1895 VSS.n1894 3.1005
R2786 VSS.n1901 VSS.n1900 3.1005
R2787 VSS.n1905 VSS.n1904 3.1005
R2788 VSS.n1909 VSS.n1908 3.1005
R2789 VSS.n1913 VSS.n1912 3.1005
R2790 VSS.n1917 VSS.n1916 3.1005
R2791 VSS.n1922 VSS.n1921 3.1005
R2792 VSS.n1926 VSS.n1925 3.1005
R2793 VSS.n1930 VSS.n1929 3.1005
R2794 VSS.n1934 VSS.n1933 3.1005
R2795 VSS.n1940 VSS.n1939 3.1005
R2796 VSS.n1944 VSS.n1943 3.1005
R2797 VSS.n1948 VSS.n1947 3.1005
R2798 VSS.n1952 VSS.n1951 3.1005
R2799 VSS.n1961 VSS.n1960 3.1005
R2800 VSS.n1962 VSS.n1399 3.1005
R2801 VSS.n1973 VSS.n1972 3.1005
R2802 VSS.n1983 VSS.n1982 3.1005
R2803 VSS.n1987 VSS.n1986 3.1005
R2804 VSS.n1997 VSS.n1996 3.1005
R2805 VSS.n2001 VSS.n2000 3.1005
R2806 VSS.n2005 VSS.n2004 3.1005
R2807 VSS.n2009 VSS.n2008 3.1005
R2808 VSS.n2015 VSS.n2014 3.1005
R2809 VSS.n2019 VSS.n2018 3.1005
R2810 VSS.n2023 VSS.n2022 3.1005
R2811 VSS.n2027 VSS.n2026 3.1005
R2812 VSS.n2031 VSS.n2030 3.1005
R2813 VSS.n2036 VSS.n2035 3.1005
R2814 VSS.n2040 VSS.n2039 3.1005
R2815 VSS.n2044 VSS.n2043 3.1005
R2816 VSS.n2048 VSS.n2047 3.1005
R2817 VSS.n2054 VSS.n2053 3.1005
R2818 VSS.n2058 VSS.n2057 3.1005
R2819 VSS.n2062 VSS.n2061 3.1005
R2820 VSS.n2066 VSS.n2065 3.1005
R2821 VSS.n2075 VSS.n2074 3.1005
R2822 VSS.n2076 VSS.n1398 3.1005
R2823 VSS.n2087 VSS.n2086 3.1005
R2824 VSS.n2097 VSS.n2096 3.1005
R2825 VSS.n2101 VSS.n2100 3.1005
R2826 VSS.n2111 VSS.n2110 3.1005
R2827 VSS.n2115 VSS.n2114 3.1005
R2828 VSS.n2119 VSS.n2118 3.1005
R2829 VSS.n2123 VSS.n2122 3.1005
R2830 VSS.n2129 VSS.n2128 3.1005
R2831 VSS.n2133 VSS.n2132 3.1005
R2832 VSS.n2137 VSS.n2136 3.1005
R2833 VSS.n2141 VSS.n2140 3.1005
R2834 VSS.n2145 VSS.n2144 3.1005
R2835 VSS.n2150 VSS.n2149 3.1005
R2836 VSS.n2154 VSS.n2153 3.1005
R2837 VSS.n2158 VSS.n2157 3.1005
R2838 VSS.n2162 VSS.n2161 3.1005
R2839 VSS.n2168 VSS.n2167 3.1005
R2840 VSS.n2172 VSS.n2171 3.1005
R2841 VSS.n2176 VSS.n2175 3.1005
R2842 VSS.n2180 VSS.n2179 3.1005
R2843 VSS.n2189 VSS.n2188 3.1005
R2844 VSS.n270 VSS.n269 3.1005
R2845 VSS.n551 VSS.n546 3.1005
R2846 VSS.n544 VSS.n543 3.1005
R2847 VSS.n540 VSS.n539 3.1005
R2848 VSS.n536 VSS.n535 3.1005
R2849 VSS.n529 VSS.n528 3.1005
R2850 VSS.n524 VSS.n523 3.1005
R2851 VSS.n520 VSS.n519 3.1005
R2852 VSS.n513 VSS.n510 3.1005
R2853 VSS.n509 VSS.n508 3.1005
R2854 VSS.n504 VSS.n503 3.1005
R2855 VSS.n500 VSS.n499 3.1005
R2856 VSS.n493 VSS.n492 3.1005
R2857 VSS.n489 VSS.n488 3.1005
R2858 VSS.n484 VSS.n483 3.1005
R2859 VSS.n402 VSS.n401 3.1005
R2860 VSS.n397 VSS.n396 3.1005
R2861 VSS.n393 VSS.n392 3.1005
R2862 VSS.n386 VSS.n385 3.1005
R2863 VSS.n382 VSS.n381 3.1005
R2864 VSS.n377 VSS.n376 3.1005
R2865 VSS.n295 VSS.n294 3.1005
R2866 VSS.n290 VSS.n289 3.1005
R2867 VSS.n286 VSS.n285 3.1005
R2868 VSS.n279 VSS.n278 3.1005
R2869 VSS.n275 VSS.n274 3.1005
R2870 VSS.n299 VSS.n296 3.1005
R2871 VSS.n406 VSS.n403 3.1005
R2872 VSS.n2885 VSS.n2884 3.1005
R2873 VSS.n2880 VSS.n2879 3.1005
R2874 VSS.n2876 VSS.n2875 3.1005
R2875 VSS.n2872 VSS.n2871 3.1005
R2876 VSS.n2868 VSS.n2867 3.1005
R2877 VSS.n2862 VSS.n2861 3.1005
R2878 VSS.n2858 VSS.n2857 3.1005
R2879 VSS.n2854 VSS.n2853 3.1005
R2880 VSS.n2850 VSS.n2849 3.1005
R2881 VSS.n2845 VSS.n2844 3.1005
R2882 VSS.n2841 VSS.n2840 3.1005
R2883 VSS.n2837 VSS.n2836 3.1005
R2884 VSS.n2833 VSS.n2832 3.1005
R2885 VSS.n2829 VSS.n2828 3.1005
R2886 VSS.n2823 VSS.n2822 3.1005
R2887 VSS.n2819 VSS.n2818 3.1005
R2888 VSS.n2815 VSS.n2814 3.1005
R2889 VSS.n2811 VSS.n2810 3.1005
R2890 VSS.n2806 VSS.n2805 3.1005
R2891 VSS.n2802 VSS.n2801 3.1005
R2892 VSS.n2797 VSS.n2796 3.1005
R2893 VSS.n1303 VSS.n1302 3.1005
R2894 VSS.n2786 VSS.n2785 3.1005
R2895 VSS.n2781 VSS.n2780 3.1005
R2896 VSS.n2777 VSS.n2776 3.1005
R2897 VSS.n2773 VSS.n2772 3.1005
R2898 VSS.n2769 VSS.n2768 3.1005
R2899 VSS.n2763 VSS.n2762 3.1005
R2900 VSS.n2759 VSS.n2758 3.1005
R2901 VSS.n2755 VSS.n2754 3.1005
R2902 VSS.n2751 VSS.n2750 3.1005
R2903 VSS.n2746 VSS.n2745 3.1005
R2904 VSS.n2742 VSS.n2741 3.1005
R2905 VSS.n2738 VSS.n2737 3.1005
R2906 VSS.n2734 VSS.n2733 3.1005
R2907 VSS.n2730 VSS.n2729 3.1005
R2908 VSS.n2724 VSS.n2723 3.1005
R2909 VSS.n2720 VSS.n2719 3.1005
R2910 VSS.n2716 VSS.n2715 3.1005
R2911 VSS.n2712 VSS.n2711 3.1005
R2912 VSS.n2707 VSS.n2706 3.1005
R2913 VSS.n2703 VSS.n2702 3.1005
R2914 VSS.n2698 VSS.n2697 3.1005
R2915 VSS.n1319 VSS.n1318 3.1005
R2916 VSS.n2687 VSS.n2686 3.1005
R2917 VSS.n2682 VSS.n2681 3.1005
R2918 VSS.n2678 VSS.n2677 3.1005
R2919 VSS.n2674 VSS.n2673 3.1005
R2920 VSS.n2670 VSS.n2669 3.1005
R2921 VSS.n2664 VSS.n2663 3.1005
R2922 VSS.n2660 VSS.n2659 3.1005
R2923 VSS.n2656 VSS.n2655 3.1005
R2924 VSS.n2652 VSS.n2651 3.1005
R2925 VSS.n2647 VSS.n2646 3.1005
R2926 VSS.n2643 VSS.n2642 3.1005
R2927 VSS.n2639 VSS.n2638 3.1005
R2928 VSS.n2635 VSS.n2634 3.1005
R2929 VSS.n2631 VSS.n2630 3.1005
R2930 VSS.n2625 VSS.n2624 3.1005
R2931 VSS.n2621 VSS.n2620 3.1005
R2932 VSS.n2617 VSS.n2616 3.1005
R2933 VSS.n2613 VSS.n2612 3.1005
R2934 VSS.n2608 VSS.n2607 3.1005
R2935 VSS.n2604 VSS.n2603 3.1005
R2936 VSS.n2599 VSS.n2598 3.1005
R2937 VSS.n1335 VSS.n1334 3.1005
R2938 VSS.n2588 VSS.n2587 3.1005
R2939 VSS.n2583 VSS.n2582 3.1005
R2940 VSS.n2579 VSS.n2578 3.1005
R2941 VSS.n2575 VSS.n2574 3.1005
R2942 VSS.n2571 VSS.n2570 3.1005
R2943 VSS.n2565 VSS.n2564 3.1005
R2944 VSS.n2561 VSS.n2560 3.1005
R2945 VSS.n2557 VSS.n2556 3.1005
R2946 VSS.n2553 VSS.n2552 3.1005
R2947 VSS.n2548 VSS.n2547 3.1005
R2948 VSS.n2544 VSS.n2543 3.1005
R2949 VSS.n2540 VSS.n2539 3.1005
R2950 VSS.n2536 VSS.n2535 3.1005
R2951 VSS.n2532 VSS.n2531 3.1005
R2952 VSS.n2526 VSS.n2525 3.1005
R2953 VSS.n2522 VSS.n2521 3.1005
R2954 VSS.n2518 VSS.n2517 3.1005
R2955 VSS.n2514 VSS.n2513 3.1005
R2956 VSS.n2509 VSS.n2508 3.1005
R2957 VSS.n2505 VSS.n2504 3.1005
R2958 VSS.n2500 VSS.n2499 3.1005
R2959 VSS.n1351 VSS.n1350 3.1005
R2960 VSS.n2489 VSS.n2488 3.1005
R2961 VSS.n2484 VSS.n2483 3.1005
R2962 VSS.n2480 VSS.n2479 3.1005
R2963 VSS.n2476 VSS.n2475 3.1005
R2964 VSS.n2472 VSS.n2471 3.1005
R2965 VSS.n2466 VSS.n2465 3.1005
R2966 VSS.n2462 VSS.n2461 3.1005
R2967 VSS.n2458 VSS.n2457 3.1005
R2968 VSS.n2454 VSS.n2453 3.1005
R2969 VSS.n2449 VSS.n2448 3.1005
R2970 VSS.n2445 VSS.n2444 3.1005
R2971 VSS.n2441 VSS.n2440 3.1005
R2972 VSS.n2437 VSS.n2436 3.1005
R2973 VSS.n2433 VSS.n2432 3.1005
R2974 VSS.n2427 VSS.n2426 3.1005
R2975 VSS.n2423 VSS.n2422 3.1005
R2976 VSS.n2419 VSS.n2418 3.1005
R2977 VSS.n2415 VSS.n2414 3.1005
R2978 VSS.n2410 VSS.n2409 3.1005
R2979 VSS.n2406 VSS.n2405 3.1005
R2980 VSS.n2401 VSS.n2400 3.1005
R2981 VSS.n1367 VSS.n1366 3.1005
R2982 VSS.n2390 VSS.n2389 3.1005
R2983 VSS.n2385 VSS.n2384 3.1005
R2984 VSS.n2381 VSS.n2380 3.1005
R2985 VSS.n2377 VSS.n2376 3.1005
R2986 VSS.n2373 VSS.n2372 3.1005
R2987 VSS.n2367 VSS.n2366 3.1005
R2988 VSS.n2363 VSS.n2362 3.1005
R2989 VSS.n2359 VSS.n2358 3.1005
R2990 VSS.n2355 VSS.n2354 3.1005
R2991 VSS.n2350 VSS.n2349 3.1005
R2992 VSS.n2346 VSS.n2345 3.1005
R2993 VSS.n2342 VSS.n2341 3.1005
R2994 VSS.n2338 VSS.n2337 3.1005
R2995 VSS.n2334 VSS.n2333 3.1005
R2996 VSS.n2328 VSS.n2327 3.1005
R2997 VSS.n2324 VSS.n2323 3.1005
R2998 VSS.n2320 VSS.n2319 3.1005
R2999 VSS.n2316 VSS.n2315 3.1005
R3000 VSS.n2311 VSS.n2310 3.1005
R3001 VSS.n2307 VSS.n2306 3.1005
R3002 VSS.n2302 VSS.n2301 3.1005
R3003 VSS.n1383 VSS.n1382 3.1005
R3004 VSS.n2291 VSS.n2290 3.1005
R3005 VSS.n2286 VSS.n2285 3.1005
R3006 VSS.n2282 VSS.n2281 3.1005
R3007 VSS.n2278 VSS.n2277 3.1005
R3008 VSS.n2274 VSS.n2273 3.1005
R3009 VSS.n2268 VSS.n2267 3.1005
R3010 VSS.n2264 VSS.n2263 3.1005
R3011 VSS.n2260 VSS.n2259 3.1005
R3012 VSS.n2256 VSS.n2255 3.1005
R3013 VSS.n2251 VSS.n2250 3.1005
R3014 VSS.n2247 VSS.n2246 3.1005
R3015 VSS.n2243 VSS.n2242 3.1005
R3016 VSS.n2239 VSS.n2238 3.1005
R3017 VSS.n2235 VSS.n2234 3.1005
R3018 VSS.n2229 VSS.n2228 3.1005
R3019 VSS.n2225 VSS.n2224 3.1005
R3020 VSS.n2221 VSS.n2220 3.1005
R3021 VSS.n2217 VSS.n2216 3.1005
R3022 VSS.n2212 VSS.n2211 3.1005
R3023 VSS.n2208 VSS.n2207 3.1005
R3024 VSS.n3193 VSS.n3192 3.1005
R3025 VSS.n3191 VSS.n3190 3.1005
R3026 VSS.n3186 VSS.n3185 3.1005
R3027 VSS.n3182 VSS.n3181 3.1005
R3028 VSS.n3176 VSS.n3175 3.1005
R3029 VSS.n3172 VSS.n3171 3.1005
R3030 VSS.n3166 VSS.n3165 3.1005
R3031 VSS.n3160 VSS.n3159 3.1005
R3032 VSS.n3156 VSS.n3155 3.1005
R3033 VSS.n3150 VSS.n3149 3.1005
R3034 VSS.n3146 VSS.n3145 3.1005
R3035 VSS.n3140 VSS.n3139 3.1005
R3036 VSS.n3136 VSS.n3135 3.1005
R3037 VSS.n3130 VSS.n3129 3.1005
R3038 VSS.n3126 VSS.n3125 3.1005
R3039 VSS.n3120 VSS.n3119 3.1005
R3040 VSS.n3115 VSS.n3114 3.1005
R3041 VSS.n3111 VSS.n3110 3.1005
R3042 VSS.n3105 VSS.n3104 3.1005
R3043 VSS.n3101 VSS.n3100 3.1005
R3044 VSS.n3095 VSS.n3094 3.1005
R3045 VSS.n3091 VSS.n3090 3.1005
R3046 VSS.n3085 VSS.n3084 3.1005
R3047 VSS.n3083 VSS.n3082 3.1005
R3048 VSS.n3073 VSS.n3072 3.1005
R3049 VSS.n3069 VSS.n3068 3.1005
R3050 VSS.n3063 VSS.n3062 3.1005
R3051 VSS.n3057 VSS.n3056 3.1005
R3052 VSS.n3202 VSS.n3201 3.1005
R3053 VSS.n3053 VSS.n3052 3.1005
R3054 VSS.n3043 VSS.n3042 3.1005
R3055 VSS.n3037 VSS.n3036 3.1005
R3056 VSS.n3035 VSS.n3034 3.1005
R3057 VSS.n3029 VSS.n3028 3.1005
R3058 VSS.n3018 VSS.n3017 3.1005
R3059 VSS.n3008 VSS.n3007 3.1005
R3060 VSS.n3006 VSS.n3005 3.1005
R3061 VSS.n3002 VSS.n3001 3.1005
R3062 VSS.n2996 VSS.n2995 3.1005
R3063 VSS.n2992 VSS.n2991 3.1005
R3064 VSS.n2986 VSS.n2985 3.1005
R3065 VSS.n2982 VSS.n2981 3.1005
R3066 VSS.n2977 VSS.n2976 3.1005
R3067 VSS.n2971 VSS.n2970 3.1005
R3068 VSS.n2967 VSS.n2966 3.1005
R3069 VSS.n2961 VSS.n2960 3.1005
R3070 VSS.n2957 VSS.n2956 3.1005
R3071 VSS.n2951 VSS.n2950 3.1005
R3072 VSS.n2947 VSS.n2946 3.1005
R3073 VSS.n2941 VSS.n2940 3.1005
R3074 VSS.n2937 VSS.n2936 3.1005
R3075 VSS.n2931 VSS.n2930 3.1005
R3076 VSS.n2927 VSS.n2926 3.1005
R3077 VSS.n2921 VSS.n2920 3.1005
R3078 VSS.n2915 VSS.n2914 3.1005
R3079 VSS.n2911 VSS.n2910 3.1005
R3080 VSS.n2906 VSS.n2905 3.1005
R3081 VSS.n3190 VSS.n3187 3.09016
R3082 VSS.n3155 VSS.n3154 3.09016
R3083 VSS.n2910 VSS.n2907 3.09016
R3084 VSS.n2946 VSS.n2945 3.09016
R3085 VSS.n68 VSS.n57 2.7891
R3086 VSS.n96 VSS.n95 2.7891
R3087 VSS.n135 VSS.n124 2.7891
R3088 VSS.n163 VSS.n162 2.7891
R3089 VSS.n205 VSS.n204 2.7891
R3090 VSS.n28 VSS.n27 2.7891
R3091 VSS.n291 VSS.n261 2.68147
R3092 VSS.n398 VSS.n250 2.68147
R3093 VSS.n505 VSS.n239 2.68147
R3094 VSS.n525 VSS.n234 2.68147
R3095 VSS.n1252 VSS.n1251 2.64878
R3096 VSS.n1042 VSS.n1041 2.64878
R3097 VSS.n535 VSS.n532 2.64878
R3098 VSS.n452 VSS.n451 2.64878
R3099 VSS.n345 VSS.n344 2.64878
R3100 VSS.n2287 VSS.n1387 2.52719
R3101 VSS.n2386 VSS.n1371 2.52719
R3102 VSS.n2485 VSS.n1355 2.52719
R3103 VSS.n2584 VSS.n1339 2.52719
R3104 VSS.n2683 VSS.n1323 2.52719
R3105 VSS.n2782 VSS.n1307 2.52719
R3106 VSS.n2881 VSS.n1291 2.52719
R3107 VSS.n2185 VSS.n2184 2.52719
R3108 VSS.n2071 VSS.n2070 2.52719
R3109 VSS.n1957 VSS.n1956 2.52719
R3110 VSS.n1843 VSS.n1842 2.52719
R3111 VSS.n1729 VSS.n1728 2.52719
R3112 VSS.n1615 VSS.n1614 2.52719
R3113 VSS.n1501 VSS.n1500 2.52719
R3114 VSS.n2294 VSS.n2292 2.49102
R3115 VSS.n2393 VSS.n2391 2.49102
R3116 VSS.n2492 VSS.n2490 2.49102
R3117 VSS.n2591 VSS.n2589 2.49102
R3118 VSS.n2690 VSS.n2688 2.49102
R3119 VSS.n2789 VSS.n2787 2.49102
R3120 VSS.n2888 VSS.n2886 2.49102
R3121 VSS.n2195 VSS.n2194 2.49102
R3122 VSS.n2079 VSS.n2077 2.49102
R3123 VSS.n1965 VSS.n1963 2.49102
R3124 VSS.n1851 VSS.n1849 2.49102
R3125 VSS.n1737 VSS.n1735 2.49102
R3126 VSS.n1623 VSS.n1621 2.49102
R3127 VSS.n1509 VSS.n1507 2.49102
R3128 VSS.n271 VSS.n263 2.49102
R3129 VSS.n378 VSS.n252 2.49102
R3130 VSS.n485 VSS.n241 2.49102
R3131 VSS.n545 VSS.n229 2.49102
R3132 VSS.n3079 VSS.n3078 2.49102
R3133 VSS.n3049 VSS.n3048 2.49102
R3134 VSS.n3025 VSS.n3024 2.49102
R3135 VSS.n5 VSS.n4 2.49101
R3136 VSS.n2213 VSS.n1392 2.45
R3137 VSS.n2312 VSS.n1376 2.45
R3138 VSS.n2411 VSS.n1360 2.45
R3139 VSS.n2510 VSS.n1344 2.45
R3140 VSS.n2609 VSS.n1328 2.45
R3141 VSS.n2708 VSS.n1312 2.45
R3142 VSS.n2807 VSS.n1296 2.45
R3143 VSS.n2107 VSS.n2106 2.45
R3144 VSS.n1993 VSS.n1992 2.45
R3145 VSS.n1879 VSS.n1878 2.45
R3146 VSS.n1765 VSS.n1764 2.45
R3147 VSS.n1651 VSS.n1650 2.45
R3148 VSS.n1537 VSS.n1536 2.45
R3149 VSS.n1423 VSS.n1422 2.45
R3150 VSS.n2204 VSS.n1397 2.43201
R3151 VSS.n2303 VSS.n1381 2.43201
R3152 VSS.n2402 VSS.n1365 2.43201
R3153 VSS.n2501 VSS.n1349 2.43201
R3154 VSS.n2600 VSS.n1333 2.43201
R3155 VSS.n2699 VSS.n1317 2.43201
R3156 VSS.n2798 VSS.n1301 2.43201
R3157 VSS.n2093 VSS.n2092 2.43201
R3158 VSS.n1979 VSS.n1978 2.43201
R3159 VSS.n1865 VSS.n1864 2.43201
R3160 VSS.n1751 VSS.n1750 2.43201
R3161 VSS.n1637 VSS.n1636 2.43201
R3162 VSS.n1523 VSS.n1522 2.43201
R3163 VSS.n1409 VSS.n1408 2.43201
R3164 VSS.n1177 VSS.n1176 2.42809
R3165 VSS.n1176 VSS.n1169 2.42809
R3166 VSS.n1162 VSS.n1155 2.42809
R3167 VSS.n1164 VSS.n1162 2.42809
R3168 VSS.n1146 VSS.n1139 2.42809
R3169 VSS.n1148 VSS.n1146 2.42809
R3170 VSS.n1132 VSS.n1125 2.42809
R3171 VSS.n1134 VSS.n1132 2.42809
R3172 VSS.n1116 VSS.n1109 2.42809
R3173 VSS.n1118 VSS.n1116 2.42809
R3174 VSS.n1102 VSS.n1095 2.42809
R3175 VSS.n1104 VSS.n1102 2.42809
R3176 VSS.n75 VSS.n60 2.42809
R3177 VSS.n1087 VSS.n75 2.42809
R3178 VSS.n966 VSS.n965 2.42809
R3179 VSS.n965 VSS.n958 2.42809
R3180 VSS.n951 VSS.n944 2.42809
R3181 VSS.n953 VSS.n951 2.42809
R3182 VSS.n935 VSS.n928 2.42809
R3183 VSS.n937 VSS.n935 2.42809
R3184 VSS.n921 VSS.n914 2.42809
R3185 VSS.n923 VSS.n921 2.42809
R3186 VSS.n905 VSS.n898 2.42809
R3187 VSS.n907 VSS.n905 2.42809
R3188 VSS.n891 VSS.n884 2.42809
R3189 VSS.n893 VSS.n891 2.42809
R3190 VSS.n142 VSS.n127 2.42809
R3191 VSS.n876 VSS.n142 2.42809
R3192 VSS.n737 VSS.n733 2.42809
R3193 VSS.n577 VSS.n573 2.42809
R3194 VSS.n499 VSS.n496 2.42809
R3195 VSS.n392 VSS.n389 2.42809
R3196 VSS.n285 VSS.n282 2.42809
R3197 VSS.n722 VSS.n721 2.32777
R3198 VSS.n562 VSS.n561 2.32777
R3199 VSS.n468 VSS.n467 2.32777
R3200 VSS.n361 VSS.n360 2.32777
R3201 VSS.n3100 VSS.n3097 2.2074
R3202 VSS.n827 VSS.n826 2.2074
R3203 VSS.n667 VSS.n666 2.2074
R3204 VSS.n3001 VSS.n2998 2.2074
R3205 VSS.n38 VSS.n35 2.17726
R3206 VSS.n105 VSS.n102 2.07152
R3207 VSS.n93 VSS.n90 2.06672
R3208 VSS.n3192 VSS 2.05519
R3209 VSS.n3068 VSS.n3067 1.98671
R3210 VSS.n3034 VSS.n3033 1.98671
R3211 VSS.n40 VSS.n39 1.81037
R3212 VSS.n55 VSS.n54 1.81037
R3213 VSS.n107 VSS.n106 1.81037
R3214 VSS.n122 VSS.n121 1.81037
R3215 VSS.n173 VSS.n172 1.81037
R3216 VSS.n215 VSS.n214 1.81037
R3217 VSS.n1408 VSS.n1406 1.72554
R3218 VSS.n1522 VSS.n1520 1.72554
R3219 VSS.n1636 VSS.n1634 1.72554
R3220 VSS.n1750 VSS.n1748 1.72554
R3221 VSS.n1864 VSS.n1862 1.72554
R3222 VSS.n1978 VSS.n1976 1.72554
R3223 VSS.n2092 VSS.n2090 1.72554
R3224 VSS.n1301 VSS.n1299 1.72554
R3225 VSS.n1317 VSS.n1315 1.72554
R3226 VSS.n1333 VSS.n1331 1.72554
R3227 VSS.n1349 VSS.n1347 1.72554
R3228 VSS.n1365 VSS.n1363 1.72554
R3229 VSS.n1381 VSS.n1379 1.72554
R3230 VSS.n1397 VSS.n1395 1.72554
R3231 VSS.n1422 VSS.n1420 1.67882
R3232 VSS.n1536 VSS.n1534 1.67882
R3233 VSS.n1650 VSS.n1648 1.67882
R3234 VSS.n1764 VSS.n1762 1.67882
R3235 VSS.n1878 VSS.n1876 1.67882
R3236 VSS.n1992 VSS.n1990 1.67882
R3237 VSS.n2106 VSS.n2104 1.67882
R3238 VSS.n1296 VSS.n1294 1.67882
R3239 VSS.n1312 VSS.n1310 1.67882
R3240 VSS.n1328 VSS.n1326 1.67882
R3241 VSS.n1344 VSS.n1342 1.67882
R3242 VSS.n1360 VSS.n1358 1.67882
R3243 VSS.n1376 VSS.n1374 1.67882
R3244 VSS.n1392 VSS.n1390 1.67882
R3245 VSS.n53 VSS.n50 1.61522
R3246 VSS.n120 VSS.n117 1.61522
R3247 VSS.n2889 VSS.n2888 1.57241
R3248 VSS.n1510 VSS.n1509 1.57241
R3249 VSS.n1624 VSS.n1623 1.57241
R3250 VSS.n1738 VSS.n1737 1.57241
R3251 VSS.n1852 VSS.n1851 1.57241
R3252 VSS.n1966 VSS.n1965 1.57241
R3253 VSS.n2080 VSS.n2079 1.57241
R3254 VSS.n2194 VSS.n2192 1.57241
R3255 VSS.n229 VSS.n227 1.57241
R3256 VSS.n478 VSS.n241 1.57241
R3257 VSS.n371 VSS.n252 1.57241
R3258 VSS.n264 VSS.n263 1.57241
R3259 VSS.n2790 VSS.n2789 1.57241
R3260 VSS.n2691 VSS.n2690 1.57241
R3261 VSS.n2592 VSS.n2591 1.57241
R3262 VSS.n2493 VSS.n2492 1.57241
R3263 VSS.n2394 VSS.n2393 1.57241
R3264 VSS.n2295 VSS.n2294 1.57241
R3265 VSS.n3078 VSS.n3076 1.57241
R3266 VSS.n3048 VSS.n3046 1.57241
R3267 VSS.n3024 VSS.n3022 1.57241
R3268 VSS.n4 VSS.n3 1.57193
R3269 VSS.n2849 VSS.n2846 1.54533
R3270 VSS.n2750 VSS.n2747 1.54533
R3271 VSS.n2651 VSS.n2648 1.54533
R3272 VSS.n2552 VSS.n2549 1.54533
R3273 VSS.n2453 VSS.n2450 1.54533
R3274 VSS.n2354 VSS.n2351 1.54533
R3275 VSS.n2255 VSS.n2252 1.54533
R3276 VSS.n1465 VSS.n1462 1.54533
R3277 VSS.n1579 VSS.n1576 1.54533
R3278 VSS.n1693 VSS.n1690 1.54533
R3279 VSS.n1807 VSS.n1804 1.54533
R3280 VSS.n1921 VSS.n1918 1.54533
R3281 VSS.n2035 VSS.n2032 1.54533
R3282 VSS.n2149 VSS.n2146 1.54533
R3283 VSS.n751 VSS.n750 1.50638
R3284 VSS.n591 VSS.n590 1.50638
R3285 VSS.n439 VSS.n438 1.50638
R3286 VSS.n332 VSS.n331 1.50638
R3287 VSS.n1500 VSS.n1499 1.47868
R3288 VSS.n1614 VSS.n1613 1.47868
R3289 VSS.n1728 VSS.n1727 1.47868
R3290 VSS.n1842 VSS.n1841 1.47868
R3291 VSS.n1956 VSS.n1955 1.47868
R3292 VSS.n2070 VSS.n2069 1.47868
R3293 VSS.n2184 VSS.n2183 1.47868
R3294 VSS.n1291 VSS.n1290 1.47868
R3295 VSS.n1307 VSS.n1306 1.47868
R3296 VSS.n1323 VSS.n1322 1.47868
R3297 VSS.n1339 VSS.n1338 1.47868
R3298 VSS.n1355 VSS.n1354 1.47868
R3299 VSS.n1371 VSS.n1370 1.47868
R3300 VSS.n1387 VSS.n1386 1.47868
R3301 VSS.n3090 VSS.n3054 1.32464
R3302 VSS.n1178 VSS.n1177 1.32464
R3303 VSS.n1169 VSS.n44 1.32464
R3304 VSS.n1164 VSS.n1163 1.32464
R3305 VSS.n1139 VSS.n1138 1.32464
R3306 VSS.n1148 VSS.n1147 1.32464
R3307 VSS.n1125 VSS.n1124 1.32464
R3308 VSS.n1134 VSS.n1133 1.32464
R3309 VSS.n1109 VSS.n1108 1.32464
R3310 VSS.n1118 VSS.n1117 1.32464
R3311 VSS.n1095 VSS.n1094 1.32464
R3312 VSS.n1104 VSS.n1103 1.32464
R3313 VSS.n60 VSS.n59 1.32464
R3314 VSS.n1087 VSS.n1086 1.32464
R3315 VSS.n967 VSS.n966 1.32464
R3316 VSS.n958 VSS.n111 1.32464
R3317 VSS.n953 VSS.n952 1.32464
R3318 VSS.n928 VSS.n927 1.32464
R3319 VSS.n937 VSS.n936 1.32464
R3320 VSS.n914 VSS.n913 1.32464
R3321 VSS.n923 VSS.n922 1.32464
R3322 VSS.n898 VSS.n897 1.32464
R3323 VSS.n907 VSS.n906 1.32464
R3324 VSS.n884 VSS.n883 1.32464
R3325 VSS.n893 VSS.n892 1.32464
R3326 VSS.n127 VSS.n126 1.32464
R3327 VSS.n876 VSS.n875 1.32464
R3328 VSS.n826 VSS.n825 1.32464
R3329 VSS.n666 VSS.n665 1.32464
R3330 VSS.n3008 VSS.n7 1.32464
R3331 VSS.n721 VSS.n720 1.10395
R3332 VSS.n561 VSS.n560 1.10395
R3333 VSS.n234 VSS.n232 1.0798
R3334 VSS.n239 VSS.n237 1.0798
R3335 VSS.n250 VSS.n248 1.0798
R3336 VSS.n261 VSS.n259 1.0798
R3337 VSS.n1251 VSS.n1250 0.883259
R3338 VSS.n755 VSS 0.849458
R3339 VSS.n595 VSS 0.849458
R3340 VSS.n403 VSS 0.849458
R3341 VSS.n296 VSS 0.849458
R3342 VSS.n510 VSS 0.846854
R3343 VSS.n45 VSS 0.835135
R3344 VSS.n112 VSS 0.832531
R3345 VSS.n2828 VSS.n2825 0.662569
R3346 VSS.n2729 VSS.n2726 0.662569
R3347 VSS.n2630 VSS.n2627 0.662569
R3348 VSS.n2531 VSS.n2528 0.662569
R3349 VSS.n2432 VSS.n2429 0.662569
R3350 VSS.n2333 VSS.n2330 0.662569
R3351 VSS.n2234 VSS.n2231 0.662569
R3352 VSS.n1444 VSS.n1441 0.662569
R3353 VSS.n1558 VSS.n1555 0.662569
R3354 VSS.n1672 VSS.n1669 0.662569
R3355 VSS.n1786 VSS.n1783 0.662569
R3356 VSS.n1900 VSS.n1897 0.662569
R3357 VSS.n2014 VSS.n2011 0.662569
R3358 VSS.n2128 VSS.n2125 0.662569
R3359 VSS.n1041 VSS.n1040 0.662569
R3360 VSS.n750 VSS.n749 0.662569
R3361 VSS.n590 VSS.n589 0.662569
R3362 VSS.n467 VSS.n242 0.662569
R3363 VSS.n360 VSS.n253 0.662569
R3364 VSS.n2901 VSS.n1286 0.596589
R3365 VSS.n3145 VSS.n3142 0.441879
R3366 VSS.n1079 VSS.n1078 0.441879
R3367 VSS.n80 VSS.n79 0.441879
R3368 VSS.n1070 VSS.n1060 0.441879
R3369 VSS.n1062 VSS.n1061 0.441879
R3370 VSS.n1056 VSS.n1046 0.441879
R3371 VSS.n1048 VSS.n1047 0.441879
R3372 VSS.n1042 VSS.n1029 0.441879
R3373 VSS.n1033 VSS.n1032 0.441879
R3374 VSS.n1025 VSS.n1016 0.441879
R3375 VSS.n1009 VSS.n999 0.441879
R3376 VSS.n1001 VSS.n1000 0.441879
R3377 VSS.n995 VSS.n109 0.441879
R3378 VSS.n987 VSS.n986 0.441879
R3379 VSS.n2956 VSS.n2953 0.441879
R3380 VSS.n2899 VSS.n2898 0.417681
R3381 VSS.n2900 VSS.n1287 0.417681
R3382 VSS.n546 VSS 0.232271
R3383 VSS.n77 VSS 0.229667
R3384 VSS.n470 VSS 0.229667
R3385 VSS.n363 VSS 0.229667
R3386 VSS.n3085 VSS.n3055 0.22119
R3387 VSS.n27 VSS.n11 0.22119
R3388 VSS.n11 VSS.n10 0.22119
R3389 VSS.n1280 VSS.n1270 0.22119
R3390 VSS.n1272 VSS.n1271 0.22119
R3391 VSS.n1266 VSS.n1256 0.22119
R3392 VSS.n1258 VSS.n1257 0.22119
R3393 VSS.n1252 VSS.n1239 0.22119
R3394 VSS.n1243 VSS.n1242 0.22119
R3395 VSS.n1235 VSS.n1227 0.22119
R3396 VSS.n31 VSS.n30 0.22119
R3397 VSS.n1220 VSS.n1210 0.22119
R3398 VSS.n1212 VSS.n1211 0.22119
R3399 VSS.n1206 VSS.n42 0.22119
R3400 VSS.n1198 VSS.n1197 0.22119
R3401 VSS.n95 VSS.n94 0.22119
R3402 VSS.n870 VSS.n143 0.22119
R3403 VSS.n146 VSS.n143 0.22119
R3404 VSS.n862 VSS.n861 0.22119
R3405 VSS.n861 VSS.n854 0.22119
R3406 VSS.n849 VSS.n848 0.22119
R3407 VSS.n848 VSS.n841 0.22119
R3408 VSS.n835 VSS.n834 0.22119
R3409 VSS.n834 VSS.n827 0.22119
R3410 VSS.n818 VSS.n817 0.22119
R3411 VSS.n817 VSS.n810 0.22119
R3412 VSS.n801 VSS.n800 0.22119
R3413 VSS.n800 VSS.n793 0.22119
R3414 VSS.n787 VSS.n786 0.22119
R3415 VSS.n786 VSS.n779 0.22119
R3416 VSS.n710 VSS.n185 0.22119
R3417 VSS.n188 VSS.n185 0.22119
R3418 VSS.n702 VSS.n701 0.22119
R3419 VSS.n701 VSS.n694 0.22119
R3420 VSS.n689 VSS.n688 0.22119
R3421 VSS.n688 VSS.n681 0.22119
R3422 VSS.n675 VSS.n674 0.22119
R3423 VSS.n674 VSS.n667 0.22119
R3424 VSS.n658 VSS.n657 0.22119
R3425 VSS.n657 VSS.n650 0.22119
R3426 VSS.n641 VSS.n640 0.22119
R3427 VSS.n640 VSS.n633 0.22119
R3428 VSS.n627 VSS.n626 0.22119
R3429 VSS.n626 VSS.n619 0.22119
R3430 VSS.n438 VSS.n435 0.22119
R3431 VSS.n331 VSS.n328 0.22119
R3432 VSS.n26 VSS.n25 0.22119
R3433 VSS.n3017 VSS.n3016 0.22119
R3434 VSS.n144 VSS 0.208833
R3435 VSS.n186 VSS 0.208833
R3436 VSS.n160 VSS.n157 0.174731
R3437 VSS.n202 VSS.n199 0.174731
R3438 VSS.n2900 VSS.n2899 0.159507
R3439 VSS.n2901 VSS.n2900 0.158129
R3440 VSS.n2886 VSS.n2885 0.120292
R3441 VSS.n2885 VSS.n2881 0.120292
R3442 VSS.n2881 VSS.n2880 0.120292
R3443 VSS.n2880 VSS.n2876 0.120292
R3444 VSS.n2876 VSS.n2872 0.120292
R3445 VSS.n2872 VSS.n2868 0.120292
R3446 VSS.n2868 VSS.n2862 0.120292
R3447 VSS.n2862 VSS.n2858 0.120292
R3448 VSS.n2858 VSS.n2854 0.120292
R3449 VSS.n2854 VSS.n2850 0.120292
R3450 VSS.n2850 VSS.n2845 0.120292
R3451 VSS.n2845 VSS.n2841 0.120292
R3452 VSS.n2841 VSS.n2837 0.120292
R3453 VSS.n2837 VSS.n2833 0.120292
R3454 VSS.n2833 VSS.n2829 0.120292
R3455 VSS.n2829 VSS.n2823 0.120292
R3456 VSS.n2823 VSS.n2819 0.120292
R3457 VSS.n2819 VSS.n2815 0.120292
R3458 VSS.n2815 VSS.n2811 0.120292
R3459 VSS.n2811 VSS.n2807 0.120292
R3460 VSS.n2807 VSS.n2806 0.120292
R3461 VSS.n2806 VSS.n2802 0.120292
R3462 VSS.n2802 VSS.n2798 0.120292
R3463 VSS.n2798 VSS.n2797 0.120292
R3464 VSS.n2787 VSS.n2786 0.120292
R3465 VSS.n2786 VSS.n2782 0.120292
R3466 VSS.n2782 VSS.n2781 0.120292
R3467 VSS.n2781 VSS.n2777 0.120292
R3468 VSS.n2777 VSS.n2773 0.120292
R3469 VSS.n2773 VSS.n2769 0.120292
R3470 VSS.n2769 VSS.n2763 0.120292
R3471 VSS.n2763 VSS.n2759 0.120292
R3472 VSS.n2759 VSS.n2755 0.120292
R3473 VSS.n2755 VSS.n2751 0.120292
R3474 VSS.n2751 VSS.n2746 0.120292
R3475 VSS.n2746 VSS.n2742 0.120292
R3476 VSS.n2742 VSS.n2738 0.120292
R3477 VSS.n2738 VSS.n2734 0.120292
R3478 VSS.n2734 VSS.n2730 0.120292
R3479 VSS.n2730 VSS.n2724 0.120292
R3480 VSS.n2724 VSS.n2720 0.120292
R3481 VSS.n2720 VSS.n2716 0.120292
R3482 VSS.n2716 VSS.n2712 0.120292
R3483 VSS.n2712 VSS.n2708 0.120292
R3484 VSS.n2708 VSS.n2707 0.120292
R3485 VSS.n2707 VSS.n2703 0.120292
R3486 VSS.n2703 VSS.n2699 0.120292
R3487 VSS.n2699 VSS.n2698 0.120292
R3488 VSS.n2688 VSS.n2687 0.120292
R3489 VSS.n2687 VSS.n2683 0.120292
R3490 VSS.n2683 VSS.n2682 0.120292
R3491 VSS.n2682 VSS.n2678 0.120292
R3492 VSS.n2678 VSS.n2674 0.120292
R3493 VSS.n2674 VSS.n2670 0.120292
R3494 VSS.n2670 VSS.n2664 0.120292
R3495 VSS.n2664 VSS.n2660 0.120292
R3496 VSS.n2660 VSS.n2656 0.120292
R3497 VSS.n2656 VSS.n2652 0.120292
R3498 VSS.n2652 VSS.n2647 0.120292
R3499 VSS.n2647 VSS.n2643 0.120292
R3500 VSS.n2643 VSS.n2639 0.120292
R3501 VSS.n2639 VSS.n2635 0.120292
R3502 VSS.n2635 VSS.n2631 0.120292
R3503 VSS.n2631 VSS.n2625 0.120292
R3504 VSS.n2625 VSS.n2621 0.120292
R3505 VSS.n2621 VSS.n2617 0.120292
R3506 VSS.n2617 VSS.n2613 0.120292
R3507 VSS.n2613 VSS.n2609 0.120292
R3508 VSS.n2609 VSS.n2608 0.120292
R3509 VSS.n2608 VSS.n2604 0.120292
R3510 VSS.n2604 VSS.n2600 0.120292
R3511 VSS.n2600 VSS.n2599 0.120292
R3512 VSS.n2589 VSS.n2588 0.120292
R3513 VSS.n2588 VSS.n2584 0.120292
R3514 VSS.n2584 VSS.n2583 0.120292
R3515 VSS.n2583 VSS.n2579 0.120292
R3516 VSS.n2579 VSS.n2575 0.120292
R3517 VSS.n2575 VSS.n2571 0.120292
R3518 VSS.n2571 VSS.n2565 0.120292
R3519 VSS.n2565 VSS.n2561 0.120292
R3520 VSS.n2561 VSS.n2557 0.120292
R3521 VSS.n2557 VSS.n2553 0.120292
R3522 VSS.n2553 VSS.n2548 0.120292
R3523 VSS.n2548 VSS.n2544 0.120292
R3524 VSS.n2544 VSS.n2540 0.120292
R3525 VSS.n2540 VSS.n2536 0.120292
R3526 VSS.n2536 VSS.n2532 0.120292
R3527 VSS.n2532 VSS.n2526 0.120292
R3528 VSS.n2526 VSS.n2522 0.120292
R3529 VSS.n2522 VSS.n2518 0.120292
R3530 VSS.n2518 VSS.n2514 0.120292
R3531 VSS.n2514 VSS.n2510 0.120292
R3532 VSS.n2510 VSS.n2509 0.120292
R3533 VSS.n2509 VSS.n2505 0.120292
R3534 VSS.n2505 VSS.n2501 0.120292
R3535 VSS.n2501 VSS.n2500 0.120292
R3536 VSS.n2490 VSS.n2489 0.120292
R3537 VSS.n2489 VSS.n2485 0.120292
R3538 VSS.n2485 VSS.n2484 0.120292
R3539 VSS.n2484 VSS.n2480 0.120292
R3540 VSS.n2480 VSS.n2476 0.120292
R3541 VSS.n2476 VSS.n2472 0.120292
R3542 VSS.n2472 VSS.n2466 0.120292
R3543 VSS.n2466 VSS.n2462 0.120292
R3544 VSS.n2462 VSS.n2458 0.120292
R3545 VSS.n2458 VSS.n2454 0.120292
R3546 VSS.n2454 VSS.n2449 0.120292
R3547 VSS.n2449 VSS.n2445 0.120292
R3548 VSS.n2445 VSS.n2441 0.120292
R3549 VSS.n2441 VSS.n2437 0.120292
R3550 VSS.n2437 VSS.n2433 0.120292
R3551 VSS.n2433 VSS.n2427 0.120292
R3552 VSS.n2427 VSS.n2423 0.120292
R3553 VSS.n2423 VSS.n2419 0.120292
R3554 VSS.n2419 VSS.n2415 0.120292
R3555 VSS.n2415 VSS.n2411 0.120292
R3556 VSS.n2411 VSS.n2410 0.120292
R3557 VSS.n2410 VSS.n2406 0.120292
R3558 VSS.n2406 VSS.n2402 0.120292
R3559 VSS.n2402 VSS.n2401 0.120292
R3560 VSS.n2391 VSS.n2390 0.120292
R3561 VSS.n2390 VSS.n2386 0.120292
R3562 VSS.n2386 VSS.n2385 0.120292
R3563 VSS.n2385 VSS.n2381 0.120292
R3564 VSS.n2381 VSS.n2377 0.120292
R3565 VSS.n2377 VSS.n2373 0.120292
R3566 VSS.n2373 VSS.n2367 0.120292
R3567 VSS.n2367 VSS.n2363 0.120292
R3568 VSS.n2363 VSS.n2359 0.120292
R3569 VSS.n2359 VSS.n2355 0.120292
R3570 VSS.n2355 VSS.n2350 0.120292
R3571 VSS.n2350 VSS.n2346 0.120292
R3572 VSS.n2346 VSS.n2342 0.120292
R3573 VSS.n2342 VSS.n2338 0.120292
R3574 VSS.n2338 VSS.n2334 0.120292
R3575 VSS.n2334 VSS.n2328 0.120292
R3576 VSS.n2328 VSS.n2324 0.120292
R3577 VSS.n2324 VSS.n2320 0.120292
R3578 VSS.n2320 VSS.n2316 0.120292
R3579 VSS.n2316 VSS.n2312 0.120292
R3580 VSS.n2312 VSS.n2311 0.120292
R3581 VSS.n2311 VSS.n2307 0.120292
R3582 VSS.n2307 VSS.n2303 0.120292
R3583 VSS.n2303 VSS.n2302 0.120292
R3584 VSS.n2292 VSS.n2291 0.120292
R3585 VSS.n2291 VSS.n2287 0.120292
R3586 VSS.n2287 VSS.n2286 0.120292
R3587 VSS.n2286 VSS.n2282 0.120292
R3588 VSS.n2282 VSS.n2278 0.120292
R3589 VSS.n2278 VSS.n2274 0.120292
R3590 VSS.n2274 VSS.n2268 0.120292
R3591 VSS.n2268 VSS.n2264 0.120292
R3592 VSS.n2264 VSS.n2260 0.120292
R3593 VSS.n2260 VSS.n2256 0.120292
R3594 VSS.n2256 VSS.n2251 0.120292
R3595 VSS.n2251 VSS.n2247 0.120292
R3596 VSS.n2247 VSS.n2243 0.120292
R3597 VSS.n2243 VSS.n2239 0.120292
R3598 VSS.n2239 VSS.n2235 0.120292
R3599 VSS.n2235 VSS.n2229 0.120292
R3600 VSS.n2229 VSS.n2225 0.120292
R3601 VSS.n2225 VSS.n2221 0.120292
R3602 VSS.n2221 VSS.n2217 0.120292
R3603 VSS.n2217 VSS.n2213 0.120292
R3604 VSS.n2213 VSS.n2212 0.120292
R3605 VSS.n2212 VSS.n2208 0.120292
R3606 VSS.n2208 VSS.n2204 0.120292
R3607 VSS.n2204 VSS.n2203 0.120292
R3608 VSS.n1409 VSS.n1287 0.120292
R3609 VSS.n1413 VSS.n1409 0.120292
R3610 VSS.n1417 VSS.n1413 0.120292
R3611 VSS.n1423 VSS.n1417 0.120292
R3612 VSS.n1427 VSS.n1423 0.120292
R3613 VSS.n1431 VSS.n1427 0.120292
R3614 VSS.n1435 VSS.n1431 0.120292
R3615 VSS.n1439 VSS.n1435 0.120292
R3616 VSS.n1445 VSS.n1439 0.120292
R3617 VSS.n1449 VSS.n1445 0.120292
R3618 VSS.n1453 VSS.n1449 0.120292
R3619 VSS.n1457 VSS.n1453 0.120292
R3620 VSS.n1461 VSS.n1457 0.120292
R3621 VSS.n1466 VSS.n1461 0.120292
R3622 VSS.n1470 VSS.n1466 0.120292
R3623 VSS.n1474 VSS.n1470 0.120292
R3624 VSS.n1478 VSS.n1474 0.120292
R3625 VSS.n1484 VSS.n1478 0.120292
R3626 VSS.n1488 VSS.n1484 0.120292
R3627 VSS.n1492 VSS.n1488 0.120292
R3628 VSS.n1496 VSS.n1492 0.120292
R3629 VSS.n1501 VSS.n1496 0.120292
R3630 VSS.n1505 VSS.n1501 0.120292
R3631 VSS.n1507 VSS.n1505 0.120292
R3632 VSS.n1507 VSS.n1506 0.120292
R3633 VSS.n1523 VSS.n1517 0.120292
R3634 VSS.n1527 VSS.n1523 0.120292
R3635 VSS.n1531 VSS.n1527 0.120292
R3636 VSS.n1537 VSS.n1531 0.120292
R3637 VSS.n1541 VSS.n1537 0.120292
R3638 VSS.n1545 VSS.n1541 0.120292
R3639 VSS.n1549 VSS.n1545 0.120292
R3640 VSS.n1553 VSS.n1549 0.120292
R3641 VSS.n1559 VSS.n1553 0.120292
R3642 VSS.n1563 VSS.n1559 0.120292
R3643 VSS.n1567 VSS.n1563 0.120292
R3644 VSS.n1571 VSS.n1567 0.120292
R3645 VSS.n1575 VSS.n1571 0.120292
R3646 VSS.n1580 VSS.n1575 0.120292
R3647 VSS.n1584 VSS.n1580 0.120292
R3648 VSS.n1588 VSS.n1584 0.120292
R3649 VSS.n1592 VSS.n1588 0.120292
R3650 VSS.n1598 VSS.n1592 0.120292
R3651 VSS.n1602 VSS.n1598 0.120292
R3652 VSS.n1606 VSS.n1602 0.120292
R3653 VSS.n1610 VSS.n1606 0.120292
R3654 VSS.n1615 VSS.n1610 0.120292
R3655 VSS.n1619 VSS.n1615 0.120292
R3656 VSS.n1621 VSS.n1619 0.120292
R3657 VSS.n1621 VSS.n1620 0.120292
R3658 VSS.n1637 VSS.n1631 0.120292
R3659 VSS.n1641 VSS.n1637 0.120292
R3660 VSS.n1645 VSS.n1641 0.120292
R3661 VSS.n1651 VSS.n1645 0.120292
R3662 VSS.n1655 VSS.n1651 0.120292
R3663 VSS.n1659 VSS.n1655 0.120292
R3664 VSS.n1663 VSS.n1659 0.120292
R3665 VSS.n1667 VSS.n1663 0.120292
R3666 VSS.n1673 VSS.n1667 0.120292
R3667 VSS.n1677 VSS.n1673 0.120292
R3668 VSS.n1681 VSS.n1677 0.120292
R3669 VSS.n1685 VSS.n1681 0.120292
R3670 VSS.n1689 VSS.n1685 0.120292
R3671 VSS.n1694 VSS.n1689 0.120292
R3672 VSS.n1698 VSS.n1694 0.120292
R3673 VSS.n1702 VSS.n1698 0.120292
R3674 VSS.n1706 VSS.n1702 0.120292
R3675 VSS.n1712 VSS.n1706 0.120292
R3676 VSS.n1716 VSS.n1712 0.120292
R3677 VSS.n1720 VSS.n1716 0.120292
R3678 VSS.n1724 VSS.n1720 0.120292
R3679 VSS.n1729 VSS.n1724 0.120292
R3680 VSS.n1733 VSS.n1729 0.120292
R3681 VSS.n1735 VSS.n1733 0.120292
R3682 VSS.n1735 VSS.n1734 0.120292
R3683 VSS.n1751 VSS.n1745 0.120292
R3684 VSS.n1755 VSS.n1751 0.120292
R3685 VSS.n1759 VSS.n1755 0.120292
R3686 VSS.n1765 VSS.n1759 0.120292
R3687 VSS.n1769 VSS.n1765 0.120292
R3688 VSS.n1773 VSS.n1769 0.120292
R3689 VSS.n1777 VSS.n1773 0.120292
R3690 VSS.n1781 VSS.n1777 0.120292
R3691 VSS.n1787 VSS.n1781 0.120292
R3692 VSS.n1791 VSS.n1787 0.120292
R3693 VSS.n1795 VSS.n1791 0.120292
R3694 VSS.n1799 VSS.n1795 0.120292
R3695 VSS.n1803 VSS.n1799 0.120292
R3696 VSS.n1808 VSS.n1803 0.120292
R3697 VSS.n1812 VSS.n1808 0.120292
R3698 VSS.n1816 VSS.n1812 0.120292
R3699 VSS.n1820 VSS.n1816 0.120292
R3700 VSS.n1826 VSS.n1820 0.120292
R3701 VSS.n1830 VSS.n1826 0.120292
R3702 VSS.n1834 VSS.n1830 0.120292
R3703 VSS.n1838 VSS.n1834 0.120292
R3704 VSS.n1843 VSS.n1838 0.120292
R3705 VSS.n1847 VSS.n1843 0.120292
R3706 VSS.n1849 VSS.n1847 0.120292
R3707 VSS.n1849 VSS.n1848 0.120292
R3708 VSS.n1865 VSS.n1859 0.120292
R3709 VSS.n1869 VSS.n1865 0.120292
R3710 VSS.n1873 VSS.n1869 0.120292
R3711 VSS.n1879 VSS.n1873 0.120292
R3712 VSS.n1883 VSS.n1879 0.120292
R3713 VSS.n1887 VSS.n1883 0.120292
R3714 VSS.n1891 VSS.n1887 0.120292
R3715 VSS.n1895 VSS.n1891 0.120292
R3716 VSS.n1901 VSS.n1895 0.120292
R3717 VSS.n1905 VSS.n1901 0.120292
R3718 VSS.n1909 VSS.n1905 0.120292
R3719 VSS.n1913 VSS.n1909 0.120292
R3720 VSS.n1917 VSS.n1913 0.120292
R3721 VSS.n1922 VSS.n1917 0.120292
R3722 VSS.n1926 VSS.n1922 0.120292
R3723 VSS.n1930 VSS.n1926 0.120292
R3724 VSS.n1934 VSS.n1930 0.120292
R3725 VSS.n1940 VSS.n1934 0.120292
R3726 VSS.n1944 VSS.n1940 0.120292
R3727 VSS.n1948 VSS.n1944 0.120292
R3728 VSS.n1952 VSS.n1948 0.120292
R3729 VSS.n1957 VSS.n1952 0.120292
R3730 VSS.n1961 VSS.n1957 0.120292
R3731 VSS.n1963 VSS.n1961 0.120292
R3732 VSS.n1963 VSS.n1962 0.120292
R3733 VSS.n1979 VSS.n1973 0.120292
R3734 VSS.n1983 VSS.n1979 0.120292
R3735 VSS.n1987 VSS.n1983 0.120292
R3736 VSS.n1993 VSS.n1987 0.120292
R3737 VSS.n1997 VSS.n1993 0.120292
R3738 VSS.n2001 VSS.n1997 0.120292
R3739 VSS.n2005 VSS.n2001 0.120292
R3740 VSS.n2009 VSS.n2005 0.120292
R3741 VSS.n2015 VSS.n2009 0.120292
R3742 VSS.n2019 VSS.n2015 0.120292
R3743 VSS.n2023 VSS.n2019 0.120292
R3744 VSS.n2027 VSS.n2023 0.120292
R3745 VSS.n2031 VSS.n2027 0.120292
R3746 VSS.n2036 VSS.n2031 0.120292
R3747 VSS.n2040 VSS.n2036 0.120292
R3748 VSS.n2044 VSS.n2040 0.120292
R3749 VSS.n2048 VSS.n2044 0.120292
R3750 VSS.n2054 VSS.n2048 0.120292
R3751 VSS.n2058 VSS.n2054 0.120292
R3752 VSS.n2062 VSS.n2058 0.120292
R3753 VSS.n2066 VSS.n2062 0.120292
R3754 VSS.n2071 VSS.n2066 0.120292
R3755 VSS.n2075 VSS.n2071 0.120292
R3756 VSS.n2077 VSS.n2075 0.120292
R3757 VSS.n2077 VSS.n2076 0.120292
R3758 VSS.n2093 VSS.n2087 0.120292
R3759 VSS.n2097 VSS.n2093 0.120292
R3760 VSS.n2101 VSS.n2097 0.120292
R3761 VSS.n2107 VSS.n2101 0.120292
R3762 VSS.n2111 VSS.n2107 0.120292
R3763 VSS.n2115 VSS.n2111 0.120292
R3764 VSS.n2119 VSS.n2115 0.120292
R3765 VSS.n2123 VSS.n2119 0.120292
R3766 VSS.n2129 VSS.n2123 0.120292
R3767 VSS.n2133 VSS.n2129 0.120292
R3768 VSS.n2137 VSS.n2133 0.120292
R3769 VSS.n2141 VSS.n2137 0.120292
R3770 VSS.n2145 VSS.n2141 0.120292
R3771 VSS.n2150 VSS.n2145 0.120292
R3772 VSS.n2154 VSS.n2150 0.120292
R3773 VSS.n2158 VSS.n2154 0.120292
R3774 VSS.n2162 VSS.n2158 0.120292
R3775 VSS.n2168 VSS.n2162 0.120292
R3776 VSS.n2172 VSS.n2168 0.120292
R3777 VSS.n2176 VSS.n2172 0.120292
R3778 VSS.n2180 VSS.n2176 0.120292
R3779 VSS.n2185 VSS.n2180 0.120292
R3780 VSS.n2189 VSS.n2185 0.120292
R3781 VSS.n2195 VSS.n2189 0.120292
R3782 VSS.n2196 VSS.n2195 0.120292
R3783 VSS.n755 VSS.n754 0.120292
R3784 VSS.n754 VSS.n752 0.120292
R3785 VSS.n752 VSS.n743 0.120292
R3786 VSS.n743 VSS.n738 0.120292
R3787 VSS.n738 VSS.n730 0.120292
R3788 VSS.n730 VSS.n725 0.120292
R3789 VSS.n725 VSS.n723 0.120292
R3790 VSS.n723 VSS.n179 0.120292
R3791 VSS.n595 VSS.n594 0.120292
R3792 VSS.n594 VSS.n592 0.120292
R3793 VSS.n592 VSS.n583 0.120292
R3794 VSS.n583 VSS.n578 0.120292
R3795 VSS.n578 VSS.n570 0.120292
R3796 VSS.n570 VSS.n565 0.120292
R3797 VSS.n565 VSS.n563 0.120292
R3798 VSS.n563 VSS.n221 0.120292
R3799 VSS.n545 VSS.n544 0.120292
R3800 VSS.n544 VSS.n540 0.120292
R3801 VSS.n540 VSS.n536 0.120292
R3802 VSS.n536 VSS.n529 0.120292
R3803 VSS.n529 VSS.n525 0.120292
R3804 VSS.n525 VSS.n524 0.120292
R3805 VSS.n524 VSS.n520 0.120292
R3806 VSS.n510 VSS.n509 0.120292
R3807 VSS.n509 VSS.n505 0.120292
R3808 VSS.n505 VSS.n504 0.120292
R3809 VSS.n504 VSS.n500 0.120292
R3810 VSS.n500 VSS.n493 0.120292
R3811 VSS.n493 VSS.n489 0.120292
R3812 VSS.n489 VSS.n485 0.120292
R3813 VSS.n485 VSS.n484 0.120292
R3814 VSS.n469 VSS.n460 0.120292
R3815 VSS.n460 VSS.n458 0.120292
R3816 VSS.n458 VSS.n453 0.120292
R3817 VSS.n453 VSS.n445 0.120292
R3818 VSS.n445 VSS.n440 0.120292
R3819 VSS.n440 VSS.n431 0.120292
R3820 VSS.n431 VSS.n429 0.120292
R3821 VSS.n403 VSS.n402 0.120292
R3822 VSS.n402 VSS.n398 0.120292
R3823 VSS.n398 VSS.n397 0.120292
R3824 VSS.n397 VSS.n393 0.120292
R3825 VSS.n393 VSS.n386 0.120292
R3826 VSS.n386 VSS.n382 0.120292
R3827 VSS.n382 VSS.n378 0.120292
R3828 VSS.n378 VSS.n377 0.120292
R3829 VSS.n362 VSS.n353 0.120292
R3830 VSS.n353 VSS.n351 0.120292
R3831 VSS.n351 VSS.n346 0.120292
R3832 VSS.n346 VSS.n338 0.120292
R3833 VSS.n338 VSS.n333 0.120292
R3834 VSS.n333 VSS.n324 0.120292
R3835 VSS.n324 VSS.n322 0.120292
R3836 VSS.n296 VSS.n295 0.120292
R3837 VSS.n295 VSS.n291 0.120292
R3838 VSS.n291 VSS.n290 0.120292
R3839 VSS.n290 VSS.n286 0.120292
R3840 VSS.n286 VSS.n279 0.120292
R3841 VSS.n279 VSS.n275 0.120292
R3842 VSS.n275 VSS.n271 0.120292
R3843 VSS.n271 VSS.n270 0.120292
R3844 VSS.n2911 VSS.n2906 0.120292
R3845 VSS.n2915 VSS.n2911 0.120292
R3846 VSS.n2921 VSS.n2915 0.120292
R3847 VSS.n2927 VSS.n2921 0.120292
R3848 VSS.n2931 VSS.n2927 0.120292
R3849 VSS.n2937 VSS.n2931 0.120292
R3850 VSS.n2941 VSS.n2937 0.120292
R3851 VSS.n2947 VSS.n2941 0.120292
R3852 VSS.n2951 VSS.n2947 0.120292
R3853 VSS.n2957 VSS.n2951 0.120292
R3854 VSS.n2961 VSS.n2957 0.120292
R3855 VSS.n2967 VSS.n2961 0.120292
R3856 VSS.n2971 VSS.n2967 0.120292
R3857 VSS.n2977 VSS.n2971 0.120292
R3858 VSS.n2982 VSS.n2977 0.120292
R3859 VSS.n2986 VSS.n2982 0.120292
R3860 VSS.n2992 VSS.n2986 0.120292
R3861 VSS.n2996 VSS.n2992 0.120292
R3862 VSS.n3002 VSS.n2996 0.120292
R3863 VSS.n3006 VSS.n3002 0.120292
R3864 VSS.n3007 VSS.n3006 0.120292
R3865 VSS.n3019 VSS.n3018 0.120292
R3866 VSS.n3025 VSS.n3019 0.120292
R3867 VSS.n3029 VSS.n3025 0.120292
R3868 VSS.n3035 VSS.n3029 0.120292
R3869 VSS.n3036 VSS.n3035 0.120292
R3870 VSS.n3049 VSS.n3043 0.120292
R3871 VSS.n3053 VSS.n3049 0.120292
R3872 VSS.n3192 VSS.n3191 0.120292
R3873 VSS.n3191 VSS.n3186 0.120292
R3874 VSS.n3186 VSS.n3182 0.120292
R3875 VSS.n3182 VSS.n3176 0.120292
R3876 VSS.n3176 VSS.n3172 0.120292
R3877 VSS.n3172 VSS.n3166 0.120292
R3878 VSS.n3166 VSS.n3160 0.120292
R3879 VSS.n3160 VSS.n3156 0.120292
R3880 VSS.n3156 VSS.n3150 0.120292
R3881 VSS.n3150 VSS.n3146 0.120292
R3882 VSS.n3146 VSS.n3140 0.120292
R3883 VSS.n3140 VSS.n3136 0.120292
R3884 VSS.n3136 VSS.n3130 0.120292
R3885 VSS.n3130 VSS.n3126 0.120292
R3886 VSS.n3126 VSS.n3120 0.120292
R3887 VSS.n3120 VSS.n3115 0.120292
R3888 VSS.n3115 VSS.n3111 0.120292
R3889 VSS.n3111 VSS.n3105 0.120292
R3890 VSS.n3105 VSS.n3101 0.120292
R3891 VSS.n3101 VSS.n3095 0.120292
R3892 VSS.n3095 VSS.n3091 0.120292
R3893 VSS.n3084 VSS.n3083 0.120292
R3894 VSS.n3083 VSS.n3079 0.120292
R3895 VSS.n3079 VSS.n3073 0.120292
R3896 VSS.n3073 VSS.n3069 0.120292
R3897 VSS.n3069 VSS.n3063 0.120292
R3898 VSS.n3056 VSS.n5 0.120292
R3899 VSS.n3202 VSS.n5 0.120292
R3900 VSS.n2886 VSS 0.0981562
R3901 VSS.n2787 VSS 0.0981562
R3902 VSS.n2688 VSS 0.0981562
R3903 VSS.n2589 VSS 0.0981562
R3904 VSS.n2490 VSS 0.0981562
R3905 VSS.n2391 VSS 0.0981562
R3906 VSS.n2292 VSS 0.0981562
R3907 VSS.n1283 VSS.n1282 0.0981562
R3908 VSS.n1269 VSS.n1268 0.0981562
R3909 VSS.n1255 VSS.n1254 0.0981562
R3910 VSS.n1238 VSS.n1237 0.0981562
R3911 VSS.n1226 VSS.n1225 0.0981562
R3912 VSS.n1223 VSS.n1222 0.0981562
R3913 VSS.n1209 VSS.n1208 0.0981562
R3914 VSS.n1167 VSS.n1166 0.0981562
R3915 VSS.n1154 VSS.n1153 0.0981562
R3916 VSS.n1151 VSS.n1150 0.0981562
R3917 VSS.n1137 VSS.n1136 0.0981562
R3918 VSS.n1121 VSS.n1120 0.0981562
R3919 VSS.n1107 VSS.n1106 0.0981562
R3920 VSS.n1093 VSS.n1092 0.0981562
R3921 VSS.n1090 VSS.n1089 0.0981562
R3922 VSS.n1073 VSS.n1072 0.0981562
R3923 VSS.n1059 VSS.n1058 0.0981562
R3924 VSS.n1045 VSS.n1044 0.0981562
R3925 VSS.n1028 VSS.n1027 0.0981562
R3926 VSS.n1015 VSS.n1014 0.0981562
R3927 VSS.n1012 VSS.n1011 0.0981562
R3928 VSS.n998 VSS.n997 0.0981562
R3929 VSS.n956 VSS.n955 0.0981562
R3930 VSS.n943 VSS.n942 0.0981562
R3931 VSS.n940 VSS.n939 0.0981562
R3932 VSS.n926 VSS.n925 0.0981562
R3933 VSS.n910 VSS.n909 0.0981562
R3934 VSS.n896 VSS.n895 0.0981562
R3935 VSS.n882 VSS.n881 0.0981562
R3936 VSS.n879 VSS.n878 0.0981562
R3937 VSS.n865 VSS.n864 0.0981562
R3938 VSS.n852 VSS.n851 0.0981562
R3939 VSS.n838 VSS.n837 0.0981562
R3940 VSS.n821 VSS.n820 0.0981562
R3941 VSS.n807 VSS.n806 0.0981562
R3942 VSS.n804 VSS.n803 0.0981562
R3943 VSS.n790 VSS.n789 0.0981562
R3944 VSS.n705 VSS.n704 0.0981562
R3945 VSS.n692 VSS.n691 0.0981562
R3946 VSS.n678 VSS.n677 0.0981562
R3947 VSS.n661 VSS.n660 0.0981562
R3948 VSS.n647 VSS.n646 0.0981562
R3949 VSS.n644 VSS.n643 0.0981562
R3950 VSS.n630 VSS.n629 0.0981562
R3951 VSS VSS.n545 0.0968542
R3952 VSS VSS.n469 0.0968542
R3953 VSS VSS.n362 0.0968542
R3954 VSS VSS.n1285 0.0955521
R3955 VSS VSS.n1075 0.09425
R3956 VSS VSS.n867 0.0760208
R3957 VSS VSS.n707 0.0760208
R3958 VSS.n2797 VSS 0.0603958
R3959 VSS.n1303 VSS 0.0603958
R3960 VSS.n2698 VSS 0.0603958
R3961 VSS.n1319 VSS 0.0603958
R3962 VSS.n2599 VSS 0.0603958
R3963 VSS.n1335 VSS 0.0603958
R3964 VSS.n2500 VSS 0.0603958
R3965 VSS.n1351 VSS 0.0603958
R3966 VSS.n2401 VSS 0.0603958
R3967 VSS.n1367 VSS 0.0603958
R3968 VSS.n2302 VSS 0.0603958
R3969 VSS.n1383 VSS 0.0603958
R3970 VSS.n2203 VSS 0.0603958
R3971 VSS.n1517 VSS 0.0603958
R3972 VSS.n1631 VSS 0.0603958
R3973 VSS.n1745 VSS 0.0603958
R3974 VSS.n1859 VSS 0.0603958
R3975 VSS.n1973 VSS 0.0603958
R3976 VSS.n2087 VSS 0.0603958
R3977 VSS.n520 VSS 0.0603958
R3978 VSS.n429 VSS 0.0603958
R3979 VSS.n322 VSS 0.0603958
R3980 VSS.n3018 VSS 0.0603958
R3981 VSS.n3036 VSS 0.0603958
R3982 VSS.n3043 VSS 0.0603958
R3983 VSS VSS.n3053 0.0603958
R3984 VSS.n3084 VSS 0.0603958
R3985 VSS.n3063 VSS 0.0603958
R3986 VSS.n3056 VSS 0.0603958
R3987 VSS VSS.n3202 0.0603958
R3988 VSS VSS.n174 0.0590938
R3989 VSS VSS.n216 0.0590938
R3990 VSS VSS.n108 0.0408646
R3991 VSS VSS.n41 0.0395625
R3992 VSS.n546 VSS 0.0239375
R3993 VSS.n470 VSS 0.0239375
R3994 VSS.n363 VSS 0.0239375
R3995 VSS.n2898 VSS 0.0226354
R3996 VSS VSS.n1303 0.0226354
R3997 VSS VSS.n1319 0.0226354
R3998 VSS VSS.n1335 0.0226354
R3999 VSS VSS.n1351 0.0226354
R4000 VSS VSS.n1367 0.0226354
R4001 VSS VSS.n1383 0.0226354
R4002 VSS.n1506 VSS 0.0226354
R4003 VSS.n1620 VSS 0.0226354
R4004 VSS.n1734 VSS 0.0226354
R4005 VSS.n1848 VSS 0.0226354
R4006 VSS.n1962 VSS 0.0226354
R4007 VSS.n2076 VSS 0.0226354
R4008 VSS.n2196 VSS 0.0226354
R4009 VSS.n868 VSS 0.0226354
R4010 VSS.n708 VSS 0.0226354
R4011 VSS.n1284 VSS.n1283 0.0213333
R4012 VSS.n1281 VSS.n1269 0.0213333
R4013 VSS.n1267 VSS.n1255 0.0213333
R4014 VSS.n1236 VSS.n1226 0.0213333
R4015 VSS.n1224 VSS.n1223 0.0213333
R4016 VSS.n1221 VSS.n1209 0.0213333
R4017 VSS.n1207 VSS.n41 0.0213333
R4018 VSS.n869 VSS.n144 0.0213333
R4019 VSS.n867 VSS.n866 0.0213333
R4020 VSS.n864 VSS.n863 0.0213333
R4021 VSS.n851 VSS.n850 0.0213333
R4022 VSS.n837 VSS.n836 0.0213333
R4023 VSS.n820 VSS.n819 0.0213333
R4024 VSS.n806 VSS.n805 0.0213333
R4025 VSS.n803 VSS.n802 0.0213333
R4026 VSS.n789 VSS.n788 0.0213333
R4027 VSS VSS.n179 0.0213333
R4028 VSS.n709 VSS.n186 0.0213333
R4029 VSS.n707 VSS.n706 0.0213333
R4030 VSS.n704 VSS.n703 0.0213333
R4031 VSS.n691 VSS.n690 0.0213333
R4032 VSS.n677 VSS.n676 0.0213333
R4033 VSS.n660 VSS.n659 0.0213333
R4034 VSS.n646 VSS.n645 0.0213333
R4035 VSS.n643 VSS.n642 0.0213333
R4036 VSS.n629 VSS.n628 0.0213333
R4037 VSS VSS.n221 0.0213333
R4038 VSS.n484 VSS 0.0213333
R4039 VSS.n377 VSS 0.0213333
R4040 VSS.n270 VSS 0.0213333
R4041 VSS.n3007 VSS 0.0213333
R4042 VSS.n3091 VSS 0.0213333
R4043 VSS.n1253 VSS.n1238 0.0213333
R4044 VSS.n1077 VSS.n1076 0.0200312
R4045 VSS.n1074 VSS.n1073 0.0200312
R4046 VSS.n1071 VSS.n1059 0.0200312
R4047 VSS.n1057 VSS.n1045 0.0200312
R4048 VSS.n1043 VSS.n1028 0.0200312
R4049 VSS.n1026 VSS.n1015 0.0200312
R4050 VSS.n1013 VSS.n1012 0.0200312
R4051 VSS.n1010 VSS.n998 0.0200312
R4052 VSS.n996 VSS.n108 0.0200312
R4053 VSS.n2899 VSS 0.0195717
R4054 VSS.n1286 VSS 0.0162706
R4055 VSS.n1168 VSS.n45 0.0148229
R4056 VSS.n1166 VSS.n1165 0.0148229
R4057 VSS.n1153 VSS.n1152 0.0148229
R4058 VSS.n1150 VSS.n1149 0.0148229
R4059 VSS.n1136 VSS.n1135 0.0148229
R4060 VSS.n1120 VSS.n1119 0.0148229
R4061 VSS.n1106 VSS.n1105 0.0148229
R4062 VSS.n1092 VSS.n1091 0.0148229
R4063 VSS.n1089 VSS.n1088 0.0148229
R4064 VSS.n957 VSS.n112 0.0148229
R4065 VSS.n955 VSS.n954 0.0148229
R4066 VSS.n942 VSS.n941 0.0148229
R4067 VSS.n939 VSS.n938 0.0148229
R4068 VSS.n925 VSS.n924 0.0148229
R4069 VSS.n909 VSS.n908 0.0148229
R4070 VSS.n895 VSS.n894 0.0148229
R4071 VSS.n881 VSS.n880 0.0148229
R4072 VSS.n878 VSS.n877 0.0148229
R4073 VSS VSS.n58 0.0135208
R4074 VSS VSS.n125 0.0135208
R4075 VSS.n1168 VSS.n1167 0.0083125
R4076 VSS.n1165 VSS.n1154 0.0083125
R4077 VSS.n1152 VSS.n1151 0.0083125
R4078 VSS.n1149 VSS.n1137 0.0083125
R4079 VSS.n1135 VSS.n1121 0.0083125
R4080 VSS.n1119 VSS.n1107 0.0083125
R4081 VSS.n1105 VSS.n1093 0.0083125
R4082 VSS.n1091 VSS.n1090 0.0083125
R4083 VSS.n1088 VSS.n58 0.0083125
R4084 VSS.n957 VSS.n956 0.0083125
R4085 VSS.n954 VSS.n943 0.0083125
R4086 VSS.n941 VSS.n940 0.0083125
R4087 VSS.n938 VSS.n926 0.0083125
R4088 VSS.n924 VSS.n910 0.0083125
R4089 VSS.n908 VSS.n896 0.0083125
R4090 VSS.n894 VSS.n882 0.0083125
R4091 VSS.n880 VSS.n879 0.0083125
R4092 VSS.n877 VSS.n125 0.0083125
R4093 VSS.n1076 VSS 0.00440625
R4094 VSS.n1077 VSS.n77 0.00310417
R4095 VSS.n1075 VSS.n1074 0.00310417
R4096 VSS.n1072 VSS.n1071 0.00310417
R4097 VSS.n1058 VSS.n1057 0.00310417
R4098 VSS.n1044 VSS.n1043 0.00310417
R4099 VSS.n1027 VSS.n1026 0.00310417
R4100 VSS.n1014 VSS.n1013 0.00310417
R4101 VSS.n1011 VSS.n1010 0.00310417
R4102 VSS.n997 VSS.n996 0.00310417
R4103 VSS.n1285 VSS.n1284 0.00180208
R4104 VSS.n1282 VSS.n1281 0.00180208
R4105 VSS.n1268 VSS.n1267 0.00180208
R4106 VSS.n1254 VSS.n1253 0.00180208
R4107 VSS.n1237 VSS.n1236 0.00180208
R4108 VSS.n1225 VSS.n1224 0.00180208
R4109 VSS.n1222 VSS.n1221 0.00180208
R4110 VSS.n1208 VSS.n1207 0.00180208
R4111 VSS.n869 VSS.n868 0.00180208
R4112 VSS.n866 VSS.n865 0.00180208
R4113 VSS.n863 VSS.n852 0.00180208
R4114 VSS.n850 VSS.n838 0.00180208
R4115 VSS.n836 VSS.n821 0.00180208
R4116 VSS.n819 VSS.n807 0.00180208
R4117 VSS.n805 VSS.n804 0.00180208
R4118 VSS.n802 VSS.n790 0.00180208
R4119 VSS.n788 VSS.n174 0.00180208
R4120 VSS.n709 VSS.n708 0.00180208
R4121 VSS.n706 VSS.n705 0.00180208
R4122 VSS.n703 VSS.n692 0.00180208
R4123 VSS.n690 VSS.n678 0.00180208
R4124 VSS.n676 VSS.n661 0.00180208
R4125 VSS.n659 VSS.n647 0.00180208
R4126 VSS.n645 VSS.n644 0.00180208
R4127 VSS.n642 VSS.n630 0.00180208
R4128 VSS.n628 VSS.n216 0.00180208
R4129 VDD.n2924 VDD.n1924 2372.71
R4130 VDD.n2926 VDD.n2925 1576.37
R4131 VDD.n2622 VDD.n2074 533.883
R4132 VDD.n940 VDD.t320 507.748
R4133 VDD.n1025 VDD.t666 500.865
R4134 VDD.n1068 VDD.t330 500.865
R4135 VDD.n1110 VDD.t720 500.865
R4136 VDD.n1152 VDD.t676 500.865
R4137 VDD.n1194 VDD.t576 500.865
R4138 VDD.n1236 VDD.t739 500.865
R4139 VDD.n1278 VDD.t57 500.865
R4140 VDD.n251 VDD.t359 500.865
R4141 VDD.n111 VDD.t314 500.865
R4142 VDD.n386 VDD.t106 500.865
R4143 VDD.n529 VDD.t434 500.865
R4144 VDD.n662 VDD.t637 500.865
R4145 VDD.n797 VDD.t22 500.865
R4146 VDD.n1761 VDD.n1760 440.25
R4147 VDD.n1680 VDD.n1679 440.25
R4148 VDD.n1603 VDD.n1602 440.25
R4149 VDD.n1526 VDD.n1525 440.25
R4150 VDD.n1449 VDD.n1448 440.25
R4151 VDD.n1372 VDD.n1371 440.25
R4152 VDD.n1295 VDD.n1294 440.25
R4153 VDD.n270 VDD.n269 440.25
R4154 VDD.n131 VDD.n130 440.25
R4155 VDD.n406 VDD.n405 440.25
R4156 VDD.n540 VDD.n539 440.25
R4157 VDD.n674 VDD.n673 440.25
R4158 VDD.n817 VDD.n816 440.25
R4159 VDD.n963 VDD.n962 440.25
R4160 VDD.t501 VDD.n200 396.851
R4161 VDD.t504 VDD.n60 396.851
R4162 VDD.t492 VDD.n335 396.851
R4163 VDD.t534 VDD.n478 396.851
R4164 VDD.t525 VDD.n611 396.851
R4165 VDD.t507 VDD.n746 396.851
R4166 VDD.t549 VDD.n889 396.851
R4167 VDD.n192 VDD.t519 391.606
R4168 VDD.n52 VDD.t540 391.606
R4169 VDD.n327 VDD.t513 391.606
R4170 VDD.n470 VDD.t495 391.606
R4171 VDD.n603 VDD.t537 391.606
R4172 VDD.n738 VDD.t528 391.606
R4173 VDD.n881 VDD.t531 391.606
R4174 VDD.n1814 VDD.t285 374.084
R4175 VDD.n1041 VDD.t67 374.084
R4176 VDD.n1081 VDD.t264 374.084
R4177 VDD.n1123 VDD.t564 374.084
R4178 VDD.n1165 VDD.t343 374.084
R4179 VDD.n1207 VDD.t131 374.084
R4180 VDD.n1249 VDD.t593 374.084
R4181 VDD.n861 VDD.t349 374.084
R4182 VDD.n718 VDD.t69 374.084
R4183 VDD.n583 VDD.t266 374.084
R4184 VDD.n450 VDD.t566 374.084
R4185 VDD.n307 VDD.t345 374.084
R4186 VDD.n32 VDD.t689 374.084
R4187 VDD.n172 VDD.t283 374.084
R4188 VDD.n2621 VDD.n2073 373.214
R4189 VDD.n2322 VDD.n2228 337.3
R4190 VDD.n2210 VDD.n2209 337.3
R4191 VDD.n2511 VDD.n2137 337.3
R4192 VDD.n2561 VDD.n2560 337.3
R4193 VDD.n2696 VDD.n2042 337.3
R4194 VDD.n2735 VDD.n2734 337.3
R4195 VDD.n2832 VDD.n1975 337.3
R4196 VDD.n2871 VDD.n2870 337.3
R4197 VDD.n1931 VDD.n1930 337.3
R4198 VDD.n1921 VDD.n1920 337.3
R4199 VDD.n1891 VDD.n1890 337.3
R4200 VDD.n1878 VDD.n1877 337.3
R4201 VDD.n1849 VDD.n1848 337.3
R4202 VDD.n1836 VDD.n1835 337.3
R4203 VDD.n1305 VDD.t511 327.223
R4204 VDD.n1382 VDD.t499 327.223
R4205 VDD.n1459 VDD.t553 327.223
R4206 VDD.n1536 VDD.t544 327.223
R4207 VDD.n1613 VDD.t523 327.223
R4208 VDD.n1690 VDD.t517 327.223
R4209 VDD.n1771 VDD.t547 327.223
R4210 VDD.n3217 VDD.n3211 324.707
R4211 VDD.n3217 VDD.n3203 324.707
R4212 VDD.n3223 VDD.n3203 324.707
R4213 VDD.n3223 VDD.n3202 324.707
R4214 VDD.n3228 VDD.n3202 324.707
R4215 VDD.n3228 VDD.n3194 324.707
R4216 VDD.n3236 VDD.n3194 324.707
R4217 VDD.n3236 VDD.n3193 324.707
R4218 VDD.n3241 VDD.n3193 324.707
R4219 VDD.n3241 VDD.n3186 324.707
R4220 VDD.n3248 VDD.n3186 324.707
R4221 VDD.n3248 VDD.n3185 324.707
R4222 VDD.n3252 VDD.n3185 324.707
R4223 VDD.n3252 VDD.n3178 324.707
R4224 VDD.n3259 VDD.n3178 324.707
R4225 VDD.n3259 VDD.n3177 324.707
R4226 VDD.n3264 VDD.n3177 324.707
R4227 VDD.n3264 VDD.n3170 324.707
R4228 VDD.n3271 VDD.n3170 324.707
R4229 VDD.n3271 VDD.n3169 324.707
R4230 VDD.n3276 VDD.n3169 324.707
R4231 VDD.n3276 VDD.n3163 324.707
R4232 VDD.n3284 VDD.n3163 324.707
R4233 VDD.n3284 VDD.n3162 324.707
R4234 VDD.n3289 VDD.n3162 324.707
R4235 VDD.n3289 VDD.n3158 324.707
R4236 VDD.n3295 VDD.n3158 324.707
R4237 VDD.n3295 VDD.n3157 324.707
R4238 VDD.n3299 VDD.n3157 324.707
R4239 VDD.n3307 VDD.n3151 324.707
R4240 VDD.n3307 VDD.n3143 324.707
R4241 VDD.n3313 VDD.n3143 324.707
R4242 VDD.n3313 VDD.n3142 324.707
R4243 VDD.n3318 VDD.n3142 324.707
R4244 VDD.n3318 VDD.n3134 324.707
R4245 VDD.n3326 VDD.n3134 324.707
R4246 VDD.n3326 VDD.n3133 324.707
R4247 VDD.n3331 VDD.n3133 324.707
R4248 VDD.n3331 VDD.n3126 324.707
R4249 VDD.n3338 VDD.n3126 324.707
R4250 VDD.n3338 VDD.n3125 324.707
R4251 VDD.n3342 VDD.n3125 324.707
R4252 VDD.n3342 VDD.n3118 324.707
R4253 VDD.n3349 VDD.n3118 324.707
R4254 VDD.n3349 VDD.n3117 324.707
R4255 VDD.n3354 VDD.n3117 324.707
R4256 VDD.n3354 VDD.n3110 324.707
R4257 VDD.n3361 VDD.n3110 324.707
R4258 VDD.n3361 VDD.n3109 324.707
R4259 VDD.n3366 VDD.n3109 324.707
R4260 VDD.n3366 VDD.n3103 324.707
R4261 VDD.n3374 VDD.n3103 324.707
R4262 VDD.n3374 VDD.n3102 324.707
R4263 VDD.n3379 VDD.n3102 324.707
R4264 VDD.n3379 VDD.n3098 324.707
R4265 VDD.n3385 VDD.n3098 324.707
R4266 VDD.n3385 VDD.n3097 324.707
R4267 VDD.n3389 VDD.n3097 324.707
R4268 VDD.n2990 VDD.n1885 324.707
R4269 VDD.n2990 VDD.n1883 324.707
R4270 VDD.n2994 VDD.n1883 324.707
R4271 VDD.n2994 VDD.n1881 324.707
R4272 VDD.n2999 VDD.n1881 324.707
R4273 VDD.n2999 VDD.n1876 324.707
R4274 VDD.n3005 VDD.n1876 324.707
R4275 VDD.n3005 VDD.n1875 324.707
R4276 VDD.n3010 VDD.n1875 324.707
R4277 VDD.n3010 VDD.n1870 324.707
R4278 VDD.n3016 VDD.n1870 324.707
R4279 VDD.n3016 VDD.n1869 324.707
R4280 VDD.n3023 VDD.n1869 324.707
R4281 VDD.n3023 VDD.n3022 324.707
R4282 VDD.n3022 VDD.n1860 324.707
R4283 VDD.n3031 VDD.n1860 324.707
R4284 VDD.n3031 VDD.n1859 324.707
R4285 VDD.n3035 VDD.n1859 324.707
R4286 VDD.n3035 VDD.n1853 324.707
R4287 VDD.n3044 VDD.n1853 324.707
R4288 VDD.n3044 VDD.n1850 324.707
R4289 VDD.n3049 VDD.n1850 324.707
R4290 VDD.n3049 VDD.n1851 324.707
R4291 VDD.n1851 VDD.n1845 324.707
R4292 VDD.n3057 VDD.n1845 324.707
R4293 VDD.n3057 VDD.n1843 324.707
R4294 VDD.n3061 VDD.n1843 324.707
R4295 VDD.n3061 VDD.n1841 324.707
R4296 VDD.n3065 VDD.n1841 324.707
R4297 VDD.n3065 VDD.n1839 324.707
R4298 VDD.n3070 VDD.n1839 324.707
R4299 VDD.n3070 VDD.n1834 324.707
R4300 VDD.n3076 VDD.n1834 324.707
R4301 VDD.n3076 VDD.n1833 324.707
R4302 VDD.n3081 VDD.n1833 324.707
R4303 VDD.n3081 VDD.n1828 324.707
R4304 VDD.n3087 VDD.n1828 324.707
R4305 VDD.n3087 VDD.n1827 324.707
R4306 VDD.n3090 VDD.n1827 324.707
R4307 VDD.n2929 VDD.n1924 324.707
R4308 VDD.n2929 VDD.n1919 324.707
R4309 VDD.n2935 VDD.n1919 324.707
R4310 VDD.n2935 VDD.n1918 324.707
R4311 VDD.n2940 VDD.n1918 324.707
R4312 VDD.n2940 VDD.n1913 324.707
R4313 VDD.n2946 VDD.n1913 324.707
R4314 VDD.n2946 VDD.n1911 324.707
R4315 VDD.n2952 VDD.n1911 324.707
R4316 VDD.n2952 VDD.n1912 324.707
R4317 VDD.n1912 VDD.n1902 324.707
R4318 VDD.n2960 VDD.n1902 324.707
R4319 VDD.n2960 VDD.n1901 324.707
R4320 VDD.n2964 VDD.n1901 324.707
R4321 VDD.n2964 VDD.n1895 324.707
R4322 VDD.n2973 VDD.n1895 324.707
R4323 VDD.n2973 VDD.n1892 324.707
R4324 VDD.n2978 VDD.n1892 324.707
R4325 VDD.n2978 VDD.n1893 324.707
R4326 VDD.n1893 VDD.n1887 324.707
R4327 VDD.n2718 VDD.n2030 324.707
R4328 VDD.n2718 VDD.n2028 324.707
R4329 VDD.n2722 VDD.n2028 324.707
R4330 VDD.n2722 VDD.n2026 324.707
R4331 VDD.n2727 VDD.n2026 324.707
R4332 VDD.n2727 VDD.n2024 324.707
R4333 VDD.n2732 VDD.n2024 324.707
R4334 VDD.n2732 VDD.n2019 324.707
R4335 VDD.n2743 VDD.n2019 324.707
R4336 VDD.n2743 VDD.n2018 324.707
R4337 VDD.n2748 VDD.n2018 324.707
R4338 VDD.n2748 VDD.n2011 324.707
R4339 VDD.n2758 VDD.n2011 324.707
R4340 VDD.n2758 VDD.n2010 324.707
R4341 VDD.n2762 VDD.n2010 324.707
R4342 VDD.n2762 VDD.n2007 324.707
R4343 VDD.n2854 VDD.n1963 324.707
R4344 VDD.n2854 VDD.n1961 324.707
R4345 VDD.n2858 VDD.n1961 324.707
R4346 VDD.n2858 VDD.n1959 324.707
R4347 VDD.n2863 VDD.n1959 324.707
R4348 VDD.n2863 VDD.n1957 324.707
R4349 VDD.n2868 VDD.n1957 324.707
R4350 VDD.n2868 VDD.n1952 324.707
R4351 VDD.n2879 VDD.n1952 324.707
R4352 VDD.n2879 VDD.n1951 324.707
R4353 VDD.n2884 VDD.n1951 324.707
R4354 VDD.n2884 VDD.n1947 324.707
R4355 VDD.n2894 VDD.n1947 324.707
R4356 VDD.n2894 VDD.n1946 324.707
R4357 VDD.n2898 VDD.n1946 324.707
R4358 VDD.n2898 VDD.n1940 324.707
R4359 VDD.n2904 VDD.n1940 324.707
R4360 VDD.n2904 VDD.n1938 324.707
R4361 VDD.n2908 VDD.n1938 324.707
R4362 VDD.n2908 VDD.n1934 324.707
R4363 VDD.n2914 VDD.n1934 324.707
R4364 VDD.n2914 VDD.n1932 324.707
R4365 VDD.n2918 VDD.n1932 324.707
R4366 VDD.n2918 VDD.n1926 324.707
R4367 VDD.n2924 VDD.n1926 324.707
R4368 VDD.n2349 VDD.n2335 324.707
R4369 VDD.n2349 VDD.n2337 324.707
R4370 VDD.n2345 VDD.n2337 324.707
R4371 VDD.n2345 VDD.n2339 324.707
R4372 VDD.n2341 VDD.n2339 324.707
R4373 VDD.n2442 VDD.n2169 324.707
R4374 VDD.n2533 VDD.n2125 324.707
R4375 VDD.n2533 VDD.n2123 324.707
R4376 VDD.n2537 VDD.n2123 324.707
R4377 VDD.n2537 VDD.n2121 324.707
R4378 VDD.n2541 VDD.n2121 324.707
R4379 VDD.n1288 VDD.n1286 324.707
R4380 VDD.n1288 VDD.n1280 324.707
R4381 VDD.n1303 VDD.n1280 324.707
R4382 VDD.n1309 VDD.n1308 324.707
R4383 VDD.n1308 VDD.n1272 324.707
R4384 VDD.n1317 VDD.n1272 324.707
R4385 VDD.n1317 VDD.n1271 324.707
R4386 VDD.n1322 VDD.n1271 324.707
R4387 VDD.n1322 VDD.n1266 324.707
R4388 VDD.n1328 VDD.n1266 324.707
R4389 VDD.n1328 VDD.n1265 324.707
R4390 VDD.n1332 VDD.n1265 324.707
R4391 VDD.n1332 VDD.n1260 324.707
R4392 VDD.n1338 VDD.n1260 324.707
R4393 VDD.n1338 VDD.n1258 324.707
R4394 VDD.n1343 VDD.n1258 324.707
R4395 VDD.n1343 VDD.n1252 324.707
R4396 VDD.n1349 VDD.n1252 324.707
R4397 VDD.n1349 VDD.n1251 324.707
R4398 VDD.n1354 VDD.n1251 324.707
R4399 VDD.n1354 VDD.n1245 324.707
R4400 VDD.n1362 VDD.n1245 324.707
R4401 VDD.n1362 VDD.n1244 324.707
R4402 VDD.n1365 VDD.n1244 324.707
R4403 VDD.n1365 VDD.n1238 324.707
R4404 VDD.n1380 VDD.n1238 324.707
R4405 VDD.n1386 VDD.n1385 324.707
R4406 VDD.n1385 VDD.n1230 324.707
R4407 VDD.n1394 VDD.n1230 324.707
R4408 VDD.n1394 VDD.n1229 324.707
R4409 VDD.n1399 VDD.n1229 324.707
R4410 VDD.n1399 VDD.n1224 324.707
R4411 VDD.n1405 VDD.n1224 324.707
R4412 VDD.n1405 VDD.n1223 324.707
R4413 VDD.n1409 VDD.n1223 324.707
R4414 VDD.n1409 VDD.n1218 324.707
R4415 VDD.n1415 VDD.n1218 324.707
R4416 VDD.n1415 VDD.n1216 324.707
R4417 VDD.n1420 VDD.n1216 324.707
R4418 VDD.n1420 VDD.n1210 324.707
R4419 VDD.n1426 VDD.n1210 324.707
R4420 VDD.n1426 VDD.n1209 324.707
R4421 VDD.n1431 VDD.n1209 324.707
R4422 VDD.n1431 VDD.n1203 324.707
R4423 VDD.n1439 VDD.n1203 324.707
R4424 VDD.n1439 VDD.n1202 324.707
R4425 VDD.n1442 VDD.n1202 324.707
R4426 VDD.n1442 VDD.n1196 324.707
R4427 VDD.n1457 VDD.n1196 324.707
R4428 VDD.n1463 VDD.n1462 324.707
R4429 VDD.n1462 VDD.n1188 324.707
R4430 VDD.n1471 VDD.n1188 324.707
R4431 VDD.n1471 VDD.n1187 324.707
R4432 VDD.n1476 VDD.n1187 324.707
R4433 VDD.n1476 VDD.n1182 324.707
R4434 VDD.n1482 VDD.n1182 324.707
R4435 VDD.n1482 VDD.n1181 324.707
R4436 VDD.n1486 VDD.n1181 324.707
R4437 VDD.n1486 VDD.n1176 324.707
R4438 VDD.n1492 VDD.n1176 324.707
R4439 VDD.n1492 VDD.n1174 324.707
R4440 VDD.n1497 VDD.n1174 324.707
R4441 VDD.n1497 VDD.n1168 324.707
R4442 VDD.n1503 VDD.n1168 324.707
R4443 VDD.n1503 VDD.n1167 324.707
R4444 VDD.n1508 VDD.n1167 324.707
R4445 VDD.n1508 VDD.n1161 324.707
R4446 VDD.n1516 VDD.n1161 324.707
R4447 VDD.n1516 VDD.n1160 324.707
R4448 VDD.n1519 VDD.n1160 324.707
R4449 VDD.n1519 VDD.n1154 324.707
R4450 VDD.n1534 VDD.n1154 324.707
R4451 VDD.n1540 VDD.n1539 324.707
R4452 VDD.n1539 VDD.n1146 324.707
R4453 VDD.n1548 VDD.n1146 324.707
R4454 VDD.n1548 VDD.n1145 324.707
R4455 VDD.n1553 VDD.n1145 324.707
R4456 VDD.n1553 VDD.n1140 324.707
R4457 VDD.n1559 VDD.n1140 324.707
R4458 VDD.n1559 VDD.n1139 324.707
R4459 VDD.n1563 VDD.n1139 324.707
R4460 VDD.n1563 VDD.n1134 324.707
R4461 VDD.n1569 VDD.n1134 324.707
R4462 VDD.n1569 VDD.n1132 324.707
R4463 VDD.n1574 VDD.n1132 324.707
R4464 VDD.n1574 VDD.n1126 324.707
R4465 VDD.n1580 VDD.n1126 324.707
R4466 VDD.n1580 VDD.n1125 324.707
R4467 VDD.n1585 VDD.n1125 324.707
R4468 VDD.n1585 VDD.n1119 324.707
R4469 VDD.n1593 VDD.n1119 324.707
R4470 VDD.n1593 VDD.n1118 324.707
R4471 VDD.n1596 VDD.n1118 324.707
R4472 VDD.n1596 VDD.n1112 324.707
R4473 VDD.n1611 VDD.n1112 324.707
R4474 VDD.n1617 VDD.n1616 324.707
R4475 VDD.n1616 VDD.n1104 324.707
R4476 VDD.n1625 VDD.n1104 324.707
R4477 VDD.n1625 VDD.n1103 324.707
R4478 VDD.n1630 VDD.n1103 324.707
R4479 VDD.n1630 VDD.n1098 324.707
R4480 VDD.n1636 VDD.n1098 324.707
R4481 VDD.n1636 VDD.n1097 324.707
R4482 VDD.n1640 VDD.n1097 324.707
R4483 VDD.n1640 VDD.n1092 324.707
R4484 VDD.n1646 VDD.n1092 324.707
R4485 VDD.n1646 VDD.n1090 324.707
R4486 VDD.n1651 VDD.n1090 324.707
R4487 VDD.n1651 VDD.n1084 324.707
R4488 VDD.n1657 VDD.n1084 324.707
R4489 VDD.n1657 VDD.n1083 324.707
R4490 VDD.n1662 VDD.n1083 324.707
R4491 VDD.n1662 VDD.n1077 324.707
R4492 VDD.n1670 VDD.n1077 324.707
R4493 VDD.n1670 VDD.n1076 324.707
R4494 VDD.n1673 VDD.n1076 324.707
R4495 VDD.n1673 VDD.n1070 324.707
R4496 VDD.n1688 VDD.n1070 324.707
R4497 VDD.n1694 VDD.n1693 324.707
R4498 VDD.n1693 VDD.n1062 324.707
R4499 VDD.n1702 VDD.n1062 324.707
R4500 VDD.n1702 VDD.n1061 324.707
R4501 VDD.n1707 VDD.n1061 324.707
R4502 VDD.n1707 VDD.n1056 324.707
R4503 VDD.n1713 VDD.n1056 324.707
R4504 VDD.n1713 VDD.n1055 324.707
R4505 VDD.n1717 VDD.n1055 324.707
R4506 VDD.n1717 VDD.n1050 324.707
R4507 VDD.n1723 VDD.n1050 324.707
R4508 VDD.n1723 VDD.n1047 324.707
R4509 VDD.n1729 VDD.n1047 324.707
R4510 VDD.n1729 VDD.n1048 324.707
R4511 VDD.n1048 VDD.n1040 324.707
R4512 VDD.n1737 VDD.n1040 324.707
R4513 VDD.n1737 VDD.n1039 324.707
R4514 VDD.n1741 VDD.n1039 324.707
R4515 VDD.n1741 VDD.n1032 324.707
R4516 VDD.n1748 VDD.n1032 324.707
R4517 VDD.n1748 VDD.n1031 324.707
R4518 VDD.n1754 VDD.n1031 324.707
R4519 VDD.n1754 VDD.n1753 324.707
R4520 VDD.n1770 VDD.n1023 324.707
R4521 VDD.n1775 VDD.n1023 324.707
R4522 VDD.n1775 VDD.n1021 324.707
R4523 VDD.n1021 VDD.n1017 324.707
R4524 VDD.n1784 VDD.n1017 324.707
R4525 VDD.n1784 VDD.n1015 324.707
R4526 VDD.n1788 VDD.n1015 324.707
R4527 VDD.n1788 VDD.n1010 324.707
R4528 VDD.n1794 VDD.n1010 324.707
R4529 VDD.n1794 VDD.n1008 324.707
R4530 VDD.n1799 VDD.n1008 324.707
R4531 VDD.n1799 VDD.n1004 324.707
R4532 VDD.n1807 VDD.n1004 324.707
R4533 VDD.n1807 VDD.n1003 324.707
R4534 VDD.n1811 VDD.n1003 324.707
R4535 VDD.n1811 VDD.n999 324.707
R4536 VDD.n1818 VDD.n999 324.707
R4537 VDD.n1818 VDD.n997 324.707
R4538 VDD.n1821 VDD.n997 324.707
R4539 VDD.n2634 VDD.n2074 321.176
R4540 VDD.n2770 VDD.n2007 321.176
R4541 VDD.n2353 VDD.n2335 321.176
R4542 VDD.n2529 VDD.n2125 317.647
R4543 VDD.n1358 VDD.n1357 312.132
R4544 VDD.n1435 VDD.n1434 312.132
R4545 VDD.n1512 VDD.n1511 312.132
R4546 VDD.n1589 VDD.n1588 312.132
R4547 VDD.n1666 VDD.n1665 312.132
R4548 VDD.n1743 VDD.n1037 312.132
R4549 VDD.n995 VDD.n994 312.132
R4550 VDD.n163 VDD.n14 312.132
R4551 VDD.n852 VDD.n0 312.132
R4552 VDD.n709 VDD.n3 312.132
R4553 VDD.n574 VDD.n6 312.132
R4554 VDD.n441 VDD.n9 312.132
R4555 VDD.n298 VDD.n12 312.132
R4556 VDD.n23 VDD.n17 312.132
R4557 VDD.n1803 VDD.n1802 307.212
R4558 VDD.n1045 VDD.n1044 307.212
R4559 VDD.n1088 VDD.n1087 307.212
R4560 VDD.n1130 VDD.n1129 307.212
R4561 VDD.n1172 VDD.n1171 307.212
R4562 VDD.n1214 VDD.n1213 307.212
R4563 VDD.n1256 VDD.n1255 307.212
R4564 VDD.n877 VDD.n876 306.985
R4565 VDD.n734 VDD.n733 306.985
R4566 VDD.n599 VDD.n598 306.985
R4567 VDD.n466 VDD.n465 306.985
R4568 VDD.n323 VDD.n322 306.985
R4569 VDD.n48 VDD.n47 306.985
R4570 VDD.n188 VDD.n187 306.985
R4571 VDD.n1778 VDD.n1020 305.529
R4572 VDD.n1064 VDD.n1063 305.529
R4573 VDD.n1106 VDD.n1105 305.529
R4574 VDD.n1148 VDD.n1147 305.529
R4575 VDD.n1190 VDD.n1189 305.529
R4576 VDD.n1232 VDD.n1231 305.529
R4577 VDD.n1274 VDD.n1273 305.529
R4578 VDD.n101 VDD.n97 305.529
R4579 VDD.n930 VDD.n926 305.529
R4580 VDD.n787 VDD.n783 305.529
R4581 VDD.n652 VDD.n648 305.529
R4582 VDD.n519 VDD.n515 305.529
R4583 VDD.n376 VDD.n372 305.529
R4584 VDD.n241 VDD.n237 305.529
R4585 VDD.n2341 VDD.n2217 303.529
R4586 VDD.n2541 VDD.n2119 303.529
R4587 VDD.n2986 VDD.n1885 300.937
R4588 VDD.n2986 VDD.n1887 291.212
R4589 VDD.n1450 VDD.t552 287.159
R4590 VDD.n1527 VDD.t543 287.159
R4591 VDD.n1762 VDD.t546 287.159
R4592 VDD.n1296 VDD.t510 286.277
R4593 VDD.n1373 VDD.t498 286.277
R4594 VDD.n1604 VDD.t522 286.277
R4595 VDD.n1681 VDD.t516 286.277
R4596 VDD.n2442 VDD.n2172 285.882
R4597 VDD.n67 VDD.t505 278.947
R4598 VDD.n207 VDD.t502 278.947
R4599 VDD.n342 VDD.t493 278.947
R4600 VDD.n485 VDD.t535 278.947
R4601 VDD.n618 VDD.t526 278.947
R4602 VDD.n753 VDD.t508 278.947
R4603 VDD.n896 VDD.t550 278.947
R4604 VDD.n2450 VDD.n2169 271.765
R4605 VDD.n2714 VDD.n2030 268.236
R4606 VDD.n2850 VDD.n1963 268.236
R4607 VDD.n2638 VDD.n2067 264.707
R4608 VDD.n2653 VDD.n2065 264.707
R4609 VDD.n2660 VDD.n2058 264.707
R4610 VDD.n2672 VDD.n2054 264.707
R4611 VDD.n2676 VDD.n2048 264.707
R4612 VDD.n2690 VDD.n2046 264.707
R4613 VDD.n2698 VDD.n2038 264.707
R4614 VDD.n2710 VDD.n2034 264.707
R4615 VDD.n2774 VDD.n2000 264.707
R4616 VDD.n2789 VDD.n1998 264.707
R4617 VDD.n2796 VDD.n1991 264.707
R4618 VDD.n2808 VDD.n1987 264.707
R4619 VDD.n2812 VDD.n1981 264.707
R4620 VDD.n2826 VDD.n1979 264.707
R4621 VDD.n2834 VDD.n1971 264.707
R4622 VDD.n2846 VDD.n1967 264.707
R4623 VDD.n2265 VDD.n2253 264.707
R4624 VDD.n2278 VDD.n2249 264.707
R4625 VDD.n2282 VDD.n2244 264.707
R4626 VDD.n2296 VDD.n2242 264.707
R4627 VDD.n2303 VDD.n2235 264.707
R4628 VDD.n2316 VDD.n2231 264.707
R4629 VDD.n2320 VDD.n2225 264.707
R4630 VDD.n2357 VDD.n2222 264.707
R4631 VDD.n2367 VDD.n2215 264.707
R4632 VDD.n2374 VDD.n2205 264.707
R4633 VDD.n2387 VDD.n2201 264.707
R4634 VDD.n2391 VDD.n2195 264.707
R4635 VDD.n2403 VDD.n2193 264.707
R4636 VDD.n2410 VDD.n2185 264.707
R4637 VDD.n2423 VDD.n2181 264.707
R4638 VDD.n2427 VDD.n2173 264.707
R4639 VDD.n2454 VDD.n2162 264.707
R4640 VDD.n2468 VDD.n2160 264.707
R4641 VDD.n2475 VDD.n2153 264.707
R4642 VDD.n2487 VDD.n2149 264.707
R4643 VDD.n2491 VDD.n2143 264.707
R4644 VDD.n2505 VDD.n2141 264.707
R4645 VDD.n2513 VDD.n2133 264.707
R4646 VDD.n2525 VDD.n2129 264.707
R4647 VDD.n2553 VDD.n2116 264.707
R4648 VDD.n2557 VDD.n2109 264.707
R4649 VDD.n2572 VDD.n2107 264.707
R4650 VDD.n2579 VDD.n2100 264.707
R4651 VDD.n2591 VDD.n2096 264.707
R4652 VDD.n2595 VDD.n2089 264.707
R4653 VDD.n2609 VDD.n2086 264.707
R4654 VDD.n2619 VDD.n2080 264.707
R4655 VDD.t511 VDD.t167 255.972
R4656 VDD.t499 VDD.t259 255.972
R4657 VDD.t553 VDD.t305 255.972
R4658 VDD.t544 VDD.t617 255.972
R4659 VDD.t523 VDD.t638 255.972
R4660 VDD.t517 VDD.t571 255.972
R4661 VDD.t646 VDD.t547 255.972
R4662 VDD.n1304 VDD.n1279 242.779
R4663 VDD.n1321 VDD.n1319 242.779
R4664 VDD.n1331 VDD.n1330 242.779
R4665 VDD.n1339 VDD.n1259 242.779
R4666 VDD.n1353 VDD.n1351 242.779
R4667 VDD.n1381 VDD.n1237 242.779
R4668 VDD.n1398 VDD.n1396 242.779
R4669 VDD.n1408 VDD.n1407 242.779
R4670 VDD.n1416 VDD.n1217 242.779
R4671 VDD.n1430 VDD.n1428 242.779
R4672 VDD.n1458 VDD.n1195 242.779
R4673 VDD.n1475 VDD.n1473 242.779
R4674 VDD.n1485 VDD.n1484 242.779
R4675 VDD.n1493 VDD.n1175 242.779
R4676 VDD.n1507 VDD.n1505 242.779
R4677 VDD.n1535 VDD.n1153 242.779
R4678 VDD.n1552 VDD.n1550 242.779
R4679 VDD.n1562 VDD.n1561 242.779
R4680 VDD.n1570 VDD.n1133 242.779
R4681 VDD.n1584 VDD.n1582 242.779
R4682 VDD.n1612 VDD.n1111 242.779
R4683 VDD.n1629 VDD.n1627 242.779
R4684 VDD.n1639 VDD.n1638 242.779
R4685 VDD.n1647 VDD.n1091 242.779
R4686 VDD.n1661 VDD.n1659 242.779
R4687 VDD.n1689 VDD.n1069 242.779
R4688 VDD.n1706 VDD.n1704 242.779
R4689 VDD.n1716 VDD.n1715 242.779
R4690 VDD.n1724 VDD.n1049 242.779
R4691 VDD.n1739 VDD.n1738 242.779
R4692 VDD.n1752 VDD.n1751 242.779
R4693 VDD.n1785 VDD.n1016 242.779
R4694 VDD.n1795 VDD.n1009 242.779
R4695 VDD.n1798 VDD.n1796 242.779
R4696 VDD.n1819 VDD.n998 242.779
R4697 VDD VDD.n158 242.106
R4698 VDD VDD.n293 242.106
R4699 VDD VDD.n436 242.106
R4700 VDD VDD.n569 242.106
R4701 VDD VDD.n704 242.106
R4702 VDD VDD.n847 242.106
R4703 VDD.n1329 VDD.t741 240.139
R4704 VDD.n1406 VDD.t729 240.139
R4705 VDD.n1483 VDD.t186 240.139
R4706 VDD.n1560 VDD.t96 240.139
R4707 VDD.n1637 VDD.t702 240.139
R4708 VDD.n1714 VDD.t423 240.139
R4709 VDD.n1787 VDD.t428 240.139
R4710 VDD.n2348 VDD.n2334 240.111
R4711 VDD.n2348 VDD.n2347 240.111
R4712 VDD.n2347 VDD.n2346 240.111
R4713 VDD.n2346 VDD.n2338 240.111
R4714 VDD.n2340 VDD.n2338 240.111
R4715 VDD.n2441 VDD.n2168 240.111
R4716 VDD.n2534 VDD.n2124 240.111
R4717 VDD.n2535 VDD.n2534 240.111
R4718 VDD.n2536 VDD.n2535 240.111
R4719 VDD.n2536 VDD.n2120 240.111
R4720 VDD.n2542 VDD.n2120 240.111
R4721 VDD.n2719 VDD.n2029 240.111
R4722 VDD.n2720 VDD.n2719 240.111
R4723 VDD.n2721 VDD.n2720 240.111
R4724 VDD.n2721 VDD.n2025 240.111
R4725 VDD.n2728 VDD.n2025 240.111
R4726 VDD.n2729 VDD.n2728 240.111
R4727 VDD.n2731 VDD.n2729 240.111
R4728 VDD.n2747 VDD.n2745 240.111
R4729 VDD.n2760 VDD.n2759 240.111
R4730 VDD.n2761 VDD.n2006 240.111
R4731 VDD.n2855 VDD.n1962 240.111
R4732 VDD.n2856 VDD.n2855 240.111
R4733 VDD.n2857 VDD.n2856 240.111
R4734 VDD.n2857 VDD.n1958 240.111
R4735 VDD.n2864 VDD.n1958 240.111
R4736 VDD.n2865 VDD.n2864 240.111
R4737 VDD.n2867 VDD.n2865 240.111
R4738 VDD.n2883 VDD.n2881 240.111
R4739 VDD.n2896 VDD.n2895 240.111
R4740 VDD.n2897 VDD.n1939 240.111
R4741 VDD.n2905 VDD.n1939 240.111
R4742 VDD.n2915 VDD.n1933 240.111
R4743 VDD.n2916 VDD.n2915 240.111
R4744 VDD.n2925 VDD.n1925 240.111
R4745 VDD.n2928 VDD.n2926 240.111
R4746 VDD.n2928 VDD.n2927 240.111
R4747 VDD.n2939 VDD.n2937 240.111
R4748 VDD.n2939 VDD.n2938 240.111
R4749 VDD.n2951 VDD.n2950 240.111
R4750 VDD.n2950 VDD.n2949 240.111
R4751 VDD.n2974 VDD.n1894 240.111
R4752 VDD.n2976 VDD.n1886 240.111
R4753 VDD.n2987 VDD.n1886 240.111
R4754 VDD.n2988 VDD.n2987 240.111
R4755 VDD.n2989 VDD.n2988 240.111
R4756 VDD.n2989 VDD.n1882 240.111
R4757 VDD.n2995 VDD.n1882 240.111
R4758 VDD.n2996 VDD.n2995 240.111
R4759 VDD.n2998 VDD.n2996 240.111
R4760 VDD.n2998 VDD.n2997 240.111
R4761 VDD.n3009 VDD.n3007 240.111
R4762 VDD.n3009 VDD.n3008 240.111
R4763 VDD.n3021 VDD.n3019 240.111
R4764 VDD.n3021 VDD.n3020 240.111
R4765 VDD.n3045 VDD.n1852 240.111
R4766 VDD.n3047 VDD.n1844 240.111
R4767 VDD.n3058 VDD.n1844 240.111
R4768 VDD.n3059 VDD.n3058 240.111
R4769 VDD.n3060 VDD.n3059 240.111
R4770 VDD.n3060 VDD.n1840 240.111
R4771 VDD.n3066 VDD.n1840 240.111
R4772 VDD.n3067 VDD.n3066 240.111
R4773 VDD.n3069 VDD.n3067 240.111
R4774 VDD.n3069 VDD.n3068 240.111
R4775 VDD.n3080 VDD.n3078 240.111
R4776 VDD.n3080 VDD.n3079 240.111
R4777 VDD.n2354 VDD.n2334 237.5
R4778 VDD.n2635 VDD.n2073 237.5
R4779 VDD.n2771 VDD.n2006 237.5
R4780 VDD.n2528 VDD.n2124 234.891
R4781 VDD.n2917 VDD.t425 234.891
R4782 VDD.n2936 VDD.t679 234.891
R4783 VDD.n3006 VDD.t356 234.891
R4784 VDD.n3077 VDD.t482 234.891
R4785 VDD.t165 VDD.n1318 232.222
R4786 VDD.t257 VDD.n1395 232.222
R4787 VDD.t303 VDD.n1472 232.222
R4788 VDD.t621 VDD.n1549 232.222
R4789 VDD.t642 VDD.n1626 232.222
R4790 VDD.t569 VDD.n1703 232.222
R4791 VDD.n1773 VDD.t644 232.222
R4792 VDD.n2340 VDD.n2216 224.452
R4793 VDD.n2543 VDD.n2542 224.452
R4794 VDD.n2949 VDD.t100 224.452
R4795 VDD.n3020 VDD.t429 224.452
R4796 VDD.t242 VDD.t230 221.667
R4797 VDD.t240 VDD.t224 221.667
R4798 VDD.t224 VDD.t700 221.667
R4799 VDD.t398 VDD.t412 221.667
R4800 VDD.t396 VDD.t416 221.667
R4801 VDD.t416 VDD.t607 221.667
R4802 VDD.t54 VDD.t215 221.667
R4803 VDD.t736 VDD.t139 221.667
R4804 VDD.t573 VDD.t150 221.667
R4805 VDD.t673 VDD.t214 221.667
R4806 VDD.t721 VDD.t742 221.667
R4807 VDD.t327 VDD.t654 221.667
R4808 VDD.t73 VDD.t667 221.667
R4809 VDD.n2962 VDD 219.232
R4810 VDD.n3033 VDD 219.232
R4811 VDD.t126 VDD.n1320 219.029
R4812 VDD.t583 VDD.n1397 219.029
R4813 VDD.t323 VDD.n1474 219.029
R4814 VDD.t140 VDD.n1551 219.029
R4815 VDD.t115 VDD.n1628 219.029
R4816 VDD.t158 VDD.n1705 219.029
R4817 VDD.n1786 VDD.t112 219.029
R4818 VDD.n2441 VDD.n2440 211.401
R4819 VDD.n2963 VDD.t486 211.401
R4820 VDD.n3034 VDD.t169 211.401
R4821 VDD.n3224 VDD.t246 211.112
R4822 VDD.t226 VDD.n3225 211.112
R4823 VDD.n3314 VDD.t402 211.112
R4824 VDD.t408 VDD.n3315 211.112
R4825 VDD.n2746 VDD.t382 206.181
R4826 VDD.n2882 VDD.t632 206.181
R4827 VDD.n1340 VDD.t599 205.833
R4828 VDD.n1417 VDD.t35 205.833
R4829 VDD.n1494 VDD.t628 205.833
R4830 VDD.n1571 VDD.t88 205.833
R4831 VDD.n1648 VDD.t31 205.833
R4832 VDD.n1725 VDD.t202 205.833
R4833 VDD.t477 VDD.n1797 205.833
R4834 VDD.n1027 VDD.t757 202.559
R4835 VDD.n1678 VDD.t765 202.559
R4836 VDD.n1601 VDD.t763 202.559
R4837 VDD.n1524 VDD.t756 202.559
R4838 VDD.n1447 VDD.t753 202.559
R4839 VDD.n1370 VDD.t773 202.559
R4840 VDD.n1293 VDD.t768 202.559
R4841 VDD.n3212 VDD.t233 201.19
R4842 VDD.n3152 VDD.t393 201.19
R4843 VDD.n2451 VDD.n2168 200.963
R4844 VDD.n3251 VDD.t228 200.556
R4845 VDD.t694 VDD.n3260 200.556
R4846 VDD.n3275 VDD 200.556
R4847 VDD.n3275 VDD.t743 200.556
R4848 VDD.n3296 VDD 200.556
R4849 VDD.n3341 VDD.t410 200.556
R4850 VDD.t611 VDD.n3350 200.556
R4851 VDD.n3365 VDD 200.556
R4852 VDD.n3365 VDD.t364 200.556
R4853 VDD.n3386 VDD 200.556
R4854 VDD.n2713 VDD.n2029 198.352
R4855 VDD.n2849 VDD.n1962 198.352
R4856 VDD.n2907 VDD.t474 198.352
R4857 VDD.n2947 VDD.t465 198.352
R4858 VDD.n3017 VDD.t464 198.352
R4859 VDD.n3088 VDD.t467 198.352
R4860 VDD.n1363 VDD 197.917
R4861 VDD.n1440 VDD 197.917
R4862 VDD.n1517 VDD 197.917
R4863 VDD.n1594 VDD 197.917
R4864 VDD.n1671 VDD 197.917
R4865 VDD.n1749 VDD 197.917
R4866 VDD.n2295 VDD.n2294 195.743
R4867 VDD.n2356 VDD.n2333 195.743
R4868 VDD.n2366 VDD.n2365 195.743
R4869 VDD.n2390 VDD.n2194 195.743
R4870 VDD.n2402 VDD.n2401 195.743
R4871 VDD.n2488 VDD.n2148 195.743
R4872 VDD.n2526 VDD.n2128 195.743
R4873 VDD.n2554 VDD.n2115 195.743
R4874 VDD.n2581 VDD.n2580 195.743
R4875 VDD.n2592 VDD.n2095 195.743
R4876 VDD.n2673 VDD.n2053 195.743
R4877 VDD.n2675 VDD.n2047 195.743
R4878 VDD.n2711 VDD.n2033 195.743
R4879 VDD.n2809 VDD.n1986 195.743
R4880 VDD.n2811 VDD.n1980 195.743
R4881 VDD.n2847 VDD.n1966 195.743
R4882 VDD.n2490 VDD.t627 193.132
R4883 VDD.t37 VDD.n2304 190.523
R4884 VDD.t220 VDD.n3215 190
R4885 VDD.n3227 VDD.t236 190
R4886 VDD.t414 VDD.n3305 190
R4887 VDD.n3317 VDD.t394 190
R4888 VDD.t161 VDD.n2699 187.912
R4889 VDD.t384 VDD.n2835 187.912
R4890 VDD.t555 VDD.t461 187.912
R4891 VDD.t273 VDD.t590 187.912
R4892 VDD.t269 VDD.t159 187.912
R4893 VDD.t460 VDD.t177 187.912
R4894 VDD.n2265 VDD.n2264 185
R4895 VDD.n2266 VDD.n2265 185
R4896 VDD.n2283 VDD.n2282 185
R4897 VDD.n2282 VDD.n2281 185
R4898 VDD.n2290 VDD.n2242 185
R4899 VDD.n2294 VDD.n2242 185
R4900 VDD.n2303 VDD.n2302 185
R4901 VDD.n2304 VDD.n2303 185
R4902 VDD.n2310 VDD.n2231 185
R4903 VDD.n2306 VDD.n2231 185
R4904 VDD.n2321 VDD.n2320 185
R4905 VDD.n2320 VDD.n2319 185
R4906 VDD.n2329 VDD.n2222 185
R4907 VDD.n2333 VDD.n2222 185
R4908 VDD.n2353 VDD.n2352 185
R4909 VDD.n2354 VDD.n2353 185
R4910 VDD.n2272 VDD.n2249 185
R4911 VDD.n2268 VDD.n2249 185
R4912 VDD.n2218 VDD.n2217 185
R4913 VDD.n2217 VDD.n2216 185
R4914 VDD.n2368 VDD.n2367 185
R4915 VDD.n2367 VDD.n2366 185
R4916 VDD.n2205 VDD.n2204 185
R4917 VDD.n2376 VDD.n2205 185
R4918 VDD.n2387 VDD.n2386 185
R4919 VDD.n2388 VDD.n2387 185
R4920 VDD.n2196 VDD.n2195 185
R4921 VDD.n2195 VDD.n2194 185
R4922 VDD.n2404 VDD.n2403 185
R4923 VDD.n2403 VDD.n2402 185
R4924 VDD.n2185 VDD.n2184 185
R4925 VDD.n2412 VDD.n2185 185
R4926 VDD.n2423 VDD.n2422 185
R4927 VDD.n2424 VDD.n2423 185
R4928 VDD.n2174 VDD.n2173 185
R4929 VDD.n2173 VDD 185
R4930 VDD.n2455 VDD.n2454 185
R4931 VDD.n2454 VDD.n2453 185
R4932 VDD.n2462 VDD.n2160 185
R4933 VDD.n2466 VDD.n2160 185
R4934 VDD.n2475 VDD.n2474 185
R4935 VDD.n2476 VDD.n2475 185
R4936 VDD.n2481 VDD.n2149 185
R4937 VDD.n2149 VDD.n2148 185
R4938 VDD.n2492 VDD.n2491 185
R4939 VDD.n2491 VDD.n2490 185
R4940 VDD.n2499 VDD.n2141 185
R4941 VDD.n2503 VDD.n2141 185
R4942 VDD.n2513 VDD.n2512 185
R4943 VDD.n2514 VDD.n2513 185
R4944 VDD.n2519 VDD.n2129 185
R4945 VDD.n2129 VDD.n2128 185
R4946 VDD.n2530 VDD.n2529 185
R4947 VDD.n2529 VDD.n2528 185
R4948 VDD.n2119 VDD.n2118 185
R4949 VDD.n2543 VDD.n2119 185
R4950 VDD.n2553 VDD.n2552 185
R4951 VDD.n2554 VDD.n2553 185
R4952 VDD.n2110 VDD.n2109 185
R4953 VDD.n2109 VDD.n2108 185
R4954 VDD.n2573 VDD.n2572 185
R4955 VDD.n2572 VDD.n2571 185
R4956 VDD.n2100 VDD.n2099 185
R4957 VDD.n2581 VDD.n2100 185
R4958 VDD.n2591 VDD.n2590 185
R4959 VDD.n2592 VDD.n2591 185
R4960 VDD.n2090 VDD.n2089 185
R4961 VDD.n2089 VDD.n2088 185
R4962 VDD.n2610 VDD.n2609 185
R4963 VDD.n2609 VDD.n2608 185
R4964 VDD.n2619 VDD.n2618 185
R4965 VDD VDD.n2619 185
R4966 VDD.n2639 VDD.n2638 185
R4967 VDD.n2638 VDD.n2637 185
R4968 VDD.n2647 VDD.n2065 185
R4969 VDD.n2651 VDD.n2065 185
R4970 VDD.n2660 VDD.n2659 185
R4971 VDD.n2661 VDD.n2660 185
R4972 VDD.n2666 VDD.n2054 185
R4973 VDD.n2054 VDD.n2053 185
R4974 VDD.n2677 VDD.n2676 185
R4975 VDD.n2676 VDD.n2675 185
R4976 VDD.n2684 VDD.n2046 185
R4977 VDD.n2688 VDD.n2046 185
R4978 VDD.n2698 VDD.n2697 185
R4979 VDD.n2699 VDD.n2698 185
R4980 VDD.n2704 VDD.n2034 185
R4981 VDD.n2034 VDD.n2033 185
R4982 VDD.n2715 VDD.n2714 185
R4983 VDD.n2714 VDD.n2713 185
R4984 VDD.n2775 VDD.n2774 185
R4985 VDD.n2774 VDD.n2773 185
R4986 VDD.n2783 VDD.n1998 185
R4987 VDD.n2787 VDD.n1998 185
R4988 VDD.n2796 VDD.n2795 185
R4989 VDD.n2797 VDD.n2796 185
R4990 VDD.n2802 VDD.n1987 185
R4991 VDD.n1987 VDD.n1986 185
R4992 VDD.n2813 VDD.n2812 185
R4993 VDD.n2812 VDD.n2811 185
R4994 VDD.n2820 VDD.n1979 185
R4995 VDD.n2824 VDD.n1979 185
R4996 VDD.n2834 VDD.n2833 185
R4997 VDD.n2835 VDD.n2834 185
R4998 VDD.n2840 VDD.n1967 185
R4999 VDD.n1967 VDD.n1966 185
R5000 VDD.n2851 VDD.n2850 185
R5001 VDD.n2850 VDD.n2849 185
R5002 VDD.t463 VDD.n1894 182.692
R5003 VDD.t462 VDD.n1852 182.692
R5004 VDD.n3250 VDD.t238 179.445
R5005 VDD.t698 VDD.n3261 179.445
R5006 VDD.n3274 VDD.t747 179.445
R5007 VDD.n3340 VDD.t400 179.445
R5008 VDD.t605 VDD.n3351 179.445
R5009 VDD.n3364 VDD.t362 179.445
R5010 VDD.t301 VDD.n2688 177.474
R5011 VDD.n2747 VDD.t472 177.474
R5012 VDD.n2761 VDD 177.474
R5013 VDD.t321 VDD.n2824 177.474
R5014 VDD.n2883 VDD.t469 177.474
R5015 VDD.n2897 VDD 177.474
R5016 VDD.n3172 VDD.n3171 174.595
R5017 VDD.n3176 VDD.n3175 174.595
R5018 VDD.n3180 VDD.n3179 174.595
R5019 VDD.n3184 VDD.n3183 174.595
R5020 VDD.n3188 VDD.n3187 174.595
R5021 VDD.n3192 VDD.n3191 174.595
R5022 VDD.n3197 VDD.n3196 174.595
R5023 VDD.n3201 VDD.n3200 174.595
R5024 VDD.n3206 VDD.n3205 174.595
R5025 VDD.n3210 VDD.n3209 174.595
R5026 VDD.n3112 VDD.n3111 174.595
R5027 VDD.n3116 VDD.n3115 174.595
R5028 VDD.n3120 VDD.n3119 174.595
R5029 VDD.n3124 VDD.n3123 174.595
R5030 VDD.n3128 VDD.n3127 174.595
R5031 VDD.n3132 VDD.n3131 174.595
R5032 VDD.n3137 VDD.n3136 174.595
R5033 VDD.n3141 VDD.n3140 174.595
R5034 VDD.n3146 VDD.n3145 174.595
R5035 VDD.n3150 VDD.n3149 174.595
R5036 VDD.t546 VDD.n1027 173.638
R5037 VDD.t516 VDD.n1678 173.638
R5038 VDD.t522 VDD.n1601 173.638
R5039 VDD.t543 VDD.n1524 173.638
R5040 VDD.t552 VDD.n1447 173.638
R5041 VDD.t498 VDD.n1370 173.638
R5042 VDD.t510 VDD.n1293 173.638
R5043 VDD.t56 VDD.n1305 171.529
R5044 VDD.t738 VDD.n1382 171.529
R5045 VDD.t575 VDD.n1459 171.529
R5046 VDD.t675 VDD.n1536 171.529
R5047 VDD.t719 VDD.n1613 171.529
R5048 VDD.t329 VDD.n1690 171.529
R5049 VDD.t665 VDD.n1771 171.529
R5050 VDD.t677 VDD.n2906 169.643
R5051 VDD.n2948 VDD.t352 169.643
R5052 VDD.n3018 VDD.t686 169.643
R5053 VDD.n3089 VDD.t484 169.643
R5054 VDD.n3216 VDD.t232 168.889
R5055 VDD.n3226 VDD.t222 168.889
R5056 VDD.n3306 VDD.t392 168.889
R5057 VDD.n3316 VDD.t406 168.889
R5058 VDD.n1342 VDD.t370 168.889
R5059 VDD.n1419 VDD.t253 168.889
R5060 VDD.n1496 VDD.t707 168.889
R5061 VDD.n1573 VDD.t333 168.889
R5062 VDD.n1650 VDD.t456 168.889
R5063 VDD.n1728 VDD.t192 168.889
R5064 VDD.n1808 VDD.t50 168.889
R5065 VDD.n42 VDD.t153 168.422
R5066 VDD.n182 VDD.t441 168.422
R5067 VDD.n317 VDD.t559 168.422
R5068 VDD.n460 VDD.t725 168.422
R5069 VDD.n593 VDD.t41 168.422
R5070 VDD.n728 VDD.t64 168.422
R5071 VDD.n871 VDD.t337 168.422
R5072 VDD.n1012 VDD.n1011 166.542
R5073 VDD.n1054 VDD.n1053 166.542
R5074 VDD.n1096 VDD.n1095 166.542
R5075 VDD.n1138 VDD.n1137 166.542
R5076 VDD.n1180 VDD.n1179 166.542
R5077 VDD.n1222 VDD.n1221 166.542
R5078 VDD.n1264 VDD.n1263 166.542
R5079 VDD.n212 VDD.n211 166.542
R5080 VDD.n72 VDD.n71 166.542
R5081 VDD.n901 VDD.n900 166.542
R5082 VDD.n758 VDD.n757 166.542
R5083 VDD.n623 VDD.n622 166.542
R5084 VDD.n490 VDD.n489 166.542
R5085 VDD.n347 VDD.n346 166.542
R5086 VDD.n3161 VDD.n3160 166.381
R5087 VDD.n3101 VDD.n3100 166.381
R5088 VDD.n3155 VDD.n3154 166.006
R5089 VDD.n3095 VDD.n3094 166.006
R5090 VDD.n1285 VDD.n1284 165.578
R5091 VDD.n1243 VDD.n1242 165.578
R5092 VDD.n1201 VDD.n1200 165.578
R5093 VDD.n1159 VDD.n1158 165.578
R5094 VDD.n1117 VDD.n1116 165.578
R5095 VDD.n1075 VDD.n1074 165.578
R5096 VDD.n1035 VDD.n1034 165.578
R5097 VDD.n150 VDD.n149 165.578
R5098 VDD.n985 VDD.n984 165.578
R5099 VDD.n839 VDD.n838 165.578
R5100 VDD.n696 VDD.n695 165.578
R5101 VDD.n561 VDD.n560 165.578
R5102 VDD.n428 VDD.n427 165.578
R5103 VDD.n284 VDD.n283 165.578
R5104 VDD.n3166 VDD.n3165 164.453
R5105 VDD.n3106 VDD.n3105 164.453
R5106 VDD.n2376 VDD.t14 161.814
R5107 VDD.t374 VDD.n2108 161.814
R5108 VDD.n3173 VDD.t691 159.46
R5109 VDD.n3113 VDD.t614 159.46
R5110 VDD.n3249 VDD.t216 158.333
R5111 VDD.n3263 VDD.t692 158.333
R5112 VDD.t745 VDD.n3285 158.333
R5113 VDD.n3339 VDD.t386 158.333
R5114 VDD.n3353 VDD.t609 158.333
R5115 VDD.t366 VDD.n3375 158.333
R5116 VDD.n2977 VDD.t671 156.594
R5117 VDD.n3048 VDD.t431 156.594
R5118 VDD.n2923 VDD.n1923 155.916
R5119 VDD.n1306 VDD.t630 155.695
R5120 VDD.n1383 VDD.t596 155.695
R5121 VDD.n1460 VDD.t90 155.695
R5122 VDD.n1537 VDD.t144 155.695
R5123 VDD.n1614 VDD.t146 155.695
R5124 VDD.n1691 VDD.t490 155.695
R5125 VDD.n1774 VDD.t380 155.695
R5126 VDD.n2388 VDD.t354 151.375
R5127 VDD.t659 VDD.n2514 151.375
R5128 VDD.n2571 VDD.t454 151.375
R5129 VDD.t475 VDD.n2661 151.375
R5130 VDD.n2730 VDD.t439 151.375
R5131 VDD.t468 VDD.n2797 151.375
R5132 VDD.n2866 VDD.t86 151.375
R5133 VDD.n2319 VDD.t255 148.764
R5134 VDD.n3168 VDD.t744 148.195
R5135 VDD.n3108 VDD.t365 148.195
R5136 VDD.n3214 VDD.n3213 148.043
R5137 VDD.n3304 VDD.n3303 148.043
R5138 VDD.t234 VDD.n3237 147.779
R5139 VDD.t390 VDD.n3327 147.779
R5140 VDD.n1342 VDD.t740 147.779
R5141 VDD.n1419 VDD.t728 147.779
R5142 VDD.n1496 VDD.t185 147.779
R5143 VDD.n1573 VDD.t97 147.779
R5144 VDD.n1650 VDD.t703 147.779
R5145 VDD.n1728 VDD.t422 147.779
R5146 VDD.t427 VDD.n1808 147.779
R5147 VDD.n201 VDD.t501 146.553
R5148 VDD.n336 VDD.t492 146.553
R5149 VDD.n479 VDD.t534 146.553
R5150 VDD.n612 VDD.t525 146.553
R5151 VDD.n747 VDD.t507 146.553
R5152 VDD.n890 VDD.t549 146.553
R5153 VDD.t171 VDD.n2976 146.155
R5154 VDD.t74 VDD.n3047 146.155
R5155 VDD.t167 VDD.n1304 145.139
R5156 VDD.t259 VDD.n1381 145.139
R5157 VDD.t305 VDD.n1458 145.139
R5158 VDD.t617 VDD.n1535 145.139
R5159 VDD.t638 VDD.n1612 145.139
R5160 VDD.t571 VDD.n1689 145.139
R5161 VDD.n1752 VDD.t646 145.139
R5162 VDD.n2426 VDD.t623 143.544
R5163 VDD.n2606 VDD.t340 143.544
R5164 VDD.n61 VDD.t504 142.458
R5165 VDD.t102 VDD.n2503 140.935
R5166 VDD.n2731 VDD.t76 140.935
R5167 VDD.n2745 VDD.t38 140.935
R5168 VDD.n2867 VDD.t267 140.935
R5169 VDD.n2881 VDD.t134 140.935
R5170 VDD.t372 VDD.n1329 139.862
R5171 VDD.t251 VDD.n1406 139.862
R5172 VDD.t705 VDD.n1483 139.862
R5173 VDD.t331 VDD.n1560 139.862
R5174 VDD.t458 VDD.n1637 139.862
R5175 VDD.t194 VDD.n1714 139.862
R5176 VDD.n1787 VDD.t52 139.862
R5177 VDD.n2306 VDD.t452 138.325
R5178 VDD.n192 VDD.t767 137.93
R5179 VDD.n52 VDD.t759 137.93
R5180 VDD.n327 VDD.t772 137.93
R5181 VDD.n470 VDD.t754 137.93
R5182 VDD.n603 VDD.t760 137.93
R5183 VDD.n738 VDD.t762 137.93
R5184 VDD.n881 VDD.t761 137.93
R5185 VDD.n2456 VDD.n2165 137.606
R5186 VDD.n2263 VDD.n2257 137.606
R5187 VDD.n2430 VDD.n2177 137.606
R5188 VDD.n2616 VDD.n2081 137.606
R5189 VDD.n2641 VDD.n2070 137.606
R5190 VDD.n2015 VDD.n2013 137.606
R5191 VDD.n2777 VDD.n2003 137.606
R5192 VDD.n2891 VDD.n2890 137.606
R5193 VDD.n1943 VDD.n1942 137.606
R5194 VDD.n1908 VDD.n1907 137.606
R5195 VDD.n2958 VDD.n1904 137.606
R5196 VDD.n1866 VDD.n1865 137.606
R5197 VDD.n3029 VDD.n1862 137.606
R5198 VDD.n1826 VDD.n1825 137.606
R5199 VDD.t244 VDD.n3239 137.222
R5200 VDD.n3262 VDD.t696 137.222
R5201 VDD.t749 VDD.n3286 137.222
R5202 VDD.t404 VDD.n3329 137.222
R5203 VDD.n3352 VDD.t615 137.222
R5204 VDD.t368 VDD.n3376 137.222
R5205 VDD.n1353 VDD.t127 137.222
R5206 VDD.n1430 VDD.t581 137.222
R5207 VDD.n1507 VDD.t324 137.222
R5208 VDD.n1584 VDD.t142 137.222
R5209 VDD.n1661 VDD.t113 137.222
R5210 VDD.t156 VDD.n1739 137.222
R5211 VDD.t110 VDD.n1819 137.222
R5212 VDD.t249 VDD.n2974 135.714
R5213 VDD.t250 VDD.n3045 135.714
R5214 VDD.t603 VDD.n1286 135.118
R5215 VDD.n1287 VDD.t163 134.583
R5216 VDD.n1364 VDD.t261 134.583
R5217 VDD.n1441 VDD.t307 134.583
R5218 VDD.n1518 VDD.t619 134.583
R5219 VDD.n1595 VDD.t640 134.583
R5220 VDD.n1672 VDD.t567 134.583
R5221 VDD.t648 VDD.n1750 134.583
R5222 VDD.n200 VDD.t769 134.047
R5223 VDD.n60 VDD.t766 134.047
R5224 VDD.n335 VDD.t770 134.047
R5225 VDD.n478 VDD.t755 134.047
R5226 VDD.n611 VDD.t758 134.047
R5227 VDD.n746 VDD.t764 134.047
R5228 VDD.n889 VDD.t771 134.047
R5229 VDD.t218 VDD.n3238 126.668
R5230 VDD.n3273 VDD.t690 126.668
R5231 VDD.t0 VDD.n3287 126.668
R5232 VDD.t94 VDD.n3296 126.668
R5233 VDD.n3298 VDD.t45 126.668
R5234 VDD.t388 VDD.n3328 126.668
R5235 VDD.n3363 VDD.t613 126.668
R5236 VDD.t70 VDD.n3377 126.668
R5237 VDD.t557 VDD.n3386 126.668
R5238 VDD.n3388 VDD.t78 126.668
R5239 VDD.n1341 VDD.t129 126.668
R5240 VDD.t592 VDD.n1350 126.668
R5241 VDD VDD.t418 126.668
R5242 VDD.t309 VDD.n1363 126.668
R5243 VDD.n1418 VDD.t580 126.668
R5244 VDD.t130 VDD.n1427 126.668
R5245 VDD VDD.t669 126.668
R5246 VDD.t717 VDD.n1440 126.668
R5247 VDD.n1495 VDD.t326 126.668
R5248 VDD.t342 VDD.n1504 126.668
R5249 VDD VDD.t663 126.668
R5250 VDD.t376 VDD.n1517 126.668
R5251 VDD.n1572 VDD.t141 126.668
R5252 VDD.t563 VDD.n1581 126.668
R5253 VDD VDD.t200 126.668
R5254 VDD.t751 VDD.n1594 126.668
R5255 VDD.n1649 VDD.t116 126.668
R5256 VDD.t263 VDD.n1658 126.668
R5257 VDD VDD.t274 126.668
R5258 VDD.t655 VDD.n1671 126.668
R5259 VDD.n1727 VDD.t155 126.668
R5260 VDD.n1726 VDD.t66 126.668
R5261 VDD.t577 VDD 126.668
R5262 VDD.t2 VDD.n1749 126.668
R5263 VDD.t109 VDD.n1809 126.668
R5264 VDD.n1810 VDD.t284 126.668
R5265 VDD VDD.t210 126.668
R5266 VDD.n2412 VDD.t466 125.275
R5267 VDD.t471 VDD.n2088 125.275
R5268 VDD.t657 VDD.n2905 125.275
R5269 VDD.t710 VDD.n1306 124.028
R5270 VDD.t248 VDD.n1383 124.028
R5271 VDD.t727 VDD.n1460 124.028
R5272 VDD.t123 VDD.n1537 124.028
R5273 VDD.t296 VDD.n1614 124.028
R5274 VDD.t704 VDD.n1691 124.028
R5275 VDD.n1774 VDD.t16 124.028
R5276 VDD.n2165 VDD.t379 123.496
R5277 VDD.n2257 VDD.t685 123.496
R5278 VDD.n2177 VDD.t347 123.496
R5279 VDD.n2081 VDD.t125 123.496
R5280 VDD.n2070 VDD.t489 123.496
R5281 VDD.n2013 VDD.t383 123.496
R5282 VDD.n2003 VDD.t133 123.496
R5283 VDD.n2890 VDD.t633 123.496
R5284 VDD.n1942 VDD.t678 123.496
R5285 VDD.n1907 VDD.t353 123.496
R5286 VDD.n1904 VDD.t487 123.496
R5287 VDD.n1865 VDD.t687 123.496
R5288 VDD.n1862 VDD.t170 123.496
R5289 VDD.n1825 VDD.t485 123.496
R5290 VDD.t488 VDD.n2651 122.665
R5291 VDD.t132 VDD.n2787 122.665
R5292 VDD.n1020 VDD.t645 121.953
R5293 VDD.n1063 VDD.t570 121.953
R5294 VDD.n1105 VDD.t643 121.953
R5295 VDD.n1147 VDD.t622 121.953
R5296 VDD.n1189 VDD.t304 121.953
R5297 VDD.n1231 VDD.t258 121.953
R5298 VDD.n1273 VDD.t166 121.953
R5299 VDD.n237 VDD.t587 121.953
R5300 VDD.n97 VDD.t120 121.953
R5301 VDD.n926 VDD.t182 121.953
R5302 VDD.n783 VDD.t714 121.953
R5303 VDD.n648 VDD.t81 121.953
R5304 VDD.n515 VDD.t735 121.953
R5305 VDD.n372 VDD.t295 121.953
R5306 VDD.n2267 VDD 120.055
R5307 VDD.n1307 VDD.t710 118.751
R5308 VDD.n1384 VDD.t248 118.751
R5309 VDD.n1461 VDD.t727 118.751
R5310 VDD.n1538 VDD.t123 118.751
R5311 VDD.n1615 VDD.t296 118.751
R5312 VDD.n1692 VDD.t704 118.751
R5313 VDD.t16 VDD.n1772 118.751
R5314 VDD.n107 VDD.t312 118.421
R5315 VDD.n247 VDD.t424 118.421
R5316 VDD.n382 VDD.t445 118.421
R5317 VDD.n525 VDD.t476 118.421
R5318 VDD.n658 VDD.t339 118.421
R5319 VDD.n793 VDD.t104 118.421
R5320 VDD.n936 VDD.t47 118.421
R5321 VDD VDD.n2161 117.445
R5322 VDD.n3240 VDD.t218 116.112
R5323 VDD.t690 VDD.n3272 116.112
R5324 VDD.n3288 VDD.t0 116.112
R5325 VDD.n3297 VDD.t94 116.112
R5326 VDD.t45 VDD.n3297 116.112
R5327 VDD.n3330 VDD.t388 116.112
R5328 VDD.t613 VDD.n3362 116.112
R5329 VDD.n3378 VDD.t70 116.112
R5330 VDD.n3387 VDD.t557 116.112
R5331 VDD.t78 VDD.n3387 116.112
R5332 VDD.n1287 VDD.t603 116.112
R5333 VDD.n1350 VDD.t129 116.112
R5334 VDD.n1351 VDD.t592 116.112
R5335 VDD.n1352 VDD.t418 116.112
R5336 VDD.n1364 VDD.t309 116.112
R5337 VDD.n1427 VDD.t580 116.112
R5338 VDD.n1428 VDD.t130 116.112
R5339 VDD.n1429 VDD.t669 116.112
R5340 VDD.n1441 VDD.t717 116.112
R5341 VDD.n1504 VDD.t326 116.112
R5342 VDD.n1505 VDD.t342 116.112
R5343 VDD.n1506 VDD.t663 116.112
R5344 VDD.n1518 VDD.t376 116.112
R5345 VDD.n1581 VDD.t141 116.112
R5346 VDD.n1582 VDD.t563 116.112
R5347 VDD.n1583 VDD.t200 116.112
R5348 VDD.n1595 VDD.t751 116.112
R5349 VDD.n1658 VDD.t116 116.112
R5350 VDD.n1659 VDD.t263 116.112
R5351 VDD.n1660 VDD.t274 116.112
R5352 VDD.n1672 VDD.t655 116.112
R5353 VDD.t155 VDD.n1726 116.112
R5354 VDD.n1738 VDD.t66 116.112
R5355 VDD.n1740 VDD.t577 116.112
R5356 VDD.n1750 VDD.t2 116.112
R5357 VDD.n1810 VDD.t109 116.112
R5358 VDD.t284 VDD.n998 116.112
R5359 VDD.t210 VDD.n1820 116.112
R5360 VDD.n20 VDD.t661 115.79
R5361 VDD.n29 VDD.t688 115.79
R5362 VDD.n34 VDD.t27 115.79
R5363 VDD.n151 VDD.t196 115.79
R5364 VDD.t173 VDD.n159 115.79
R5365 VDD.n169 VDD.t282 115.79
R5366 VDD.n174 VDD.t280 115.79
R5367 VDD.n285 VDD.t270 115.79
R5368 VDD.n295 VDD.t92 115.79
R5369 VDD.n304 VDD.t344 115.79
R5370 VDD.n309 VDD.t135 115.79
R5371 VDD.n429 VDD.t4 115.79
R5372 VDD.t420 VDD.n437 115.79
R5373 VDD.n447 VDD.t565 115.79
R5374 VDD.n452 VDD.t650 115.79
R5375 VDD.n562 VDD.t625 115.79
R5376 VDD.t288 VDD.n570 115.79
R5377 VDD.n580 VDD.t265 115.79
R5378 VDD.n585 VDD.t206 115.79
R5379 VDD.n697 VDD.t190 115.79
R5380 VDD.t10 VDD.n705 115.79
R5381 VDD.n715 VDD.t68 115.79
R5382 VDD.n720 VDD.t8 115.79
R5383 VDD.n840 VDD.t450 115.79
R5384 VDD.t98 VDD.n848 115.79
R5385 VDD.n858 VDD.t348 115.79
R5386 VDD.n863 VDD.t58 115.79
R5387 VDD.n986 VDD.t175 115.79
R5388 VDD.t470 VDD.n2476 114.835
R5389 VDD.t446 VDD.n2948 114.835
R5390 VDD.t299 VDD.n3018 114.835
R5391 VDD.t43 VDD.n3089 114.835
R5392 VDD.n2279 VDD.t684 112.225
R5393 VDD.n2281 VDD.t473 112.225
R5394 VDD.n2467 VDD.t378 109.615
R5395 VDD.t163 VDD.n1279 108.195
R5396 VDD.t261 VDD.n1237 108.195
R5397 VDD.t307 VDD.n1195 108.195
R5398 VDD.t619 VDD.n1153 108.195
R5399 VDD.t640 VDD.n1111 108.195
R5400 VDD.t567 VDD.n1069 108.195
R5401 VDD.n1751 VDD.t648 108.195
R5402 VDD.n145 VDD.t121 107.895
R5403 VDD.n279 VDD.t584 107.895
R5404 VDD.n423 VDD.t290 107.895
R5405 VDD.n556 VDD.t730 107.895
R5406 VDD.n691 VDD.t84 107.895
R5407 VDD.n834 VDD.t715 107.895
R5408 VDD.n980 VDD.t179 107.895
R5409 VDD.n3240 VDD.t244 105.556
R5410 VDD.n3272 VDD.t696 105.556
R5411 VDD.n3288 VDD.t749 105.556
R5412 VDD.n3330 VDD.t404 105.556
R5413 VDD.n3362 VDD.t615 105.556
R5414 VDD.n3378 VDD.t368 105.556
R5415 VDD.t127 VDD.n1352 105.556
R5416 VDD.t581 VDD.n1429 105.556
R5417 VDD.t324 VDD.n1506 105.556
R5418 VDD.t142 VDD.n1583 105.556
R5419 VDD.t113 VDD.n1660 105.556
R5420 VDD.n1740 VDD.t156 105.556
R5421 VDD.n1820 VDD.t110 105.556
R5422 VDD.n20 VDD.t25 105.263
R5423 VDD.n159 VDD.t278 105.263
R5424 VDD.n295 VDD.t137 105.263
R5425 VDD.n437 VDD.t652 105.263
R5426 VDD.n570 VDD.t204 105.263
R5427 VDD.n705 VDD.t6 105.263
R5428 VDD.n848 VDD.t59 105.263
R5429 VDD.n2975 VDD.t249 104.397
R5430 VDD.n3046 VDD.t250 104.397
R5431 VDD.n1330 VDD.t372 102.918
R5432 VDD.n1407 VDD.t251 102.918
R5433 VDD.n1484 VDD.t705 102.918
R5434 VDD.n1561 VDD.t331 102.918
R5435 VDD.n1638 VDD.t458 102.918
R5436 VDD.n1715 VDD.t194 102.918
R5437 VDD.t52 VDD.n1009 102.918
R5438 VDD.n77 VDD.t151 102.632
R5439 VDD.n217 VDD.t443 102.632
R5440 VDD.n352 VDD.t561 102.632
R5441 VDD.n495 VDD.t723 102.632
R5442 VDD.n628 VDD.t39 102.632
R5443 VDD.n763 VDD.t62 102.632
R5444 VDD.n906 VDD.t335 102.632
R5445 VDD.n823 VDD.t711 100.001
R5446 VDD.n2413 VDD.t346 99.1763
R5447 VDD.t124 VDD.n2605 99.1763
R5448 VDD.t76 VDD.n2730 99.1763
R5449 VDD.t38 VDD.n2744 99.1763
R5450 VDD.t267 VDD.n2866 99.1763
R5451 VDD.t134 VDD.n2880 99.1763
R5452 VDD.n271 VDD.t588 97.3689
R5453 VDD.n547 VDD.t732 97.3689
R5454 VDD.n2424 VDD.t346 96.5664
R5455 VDD.n2608 VDD.t124 96.5664
R5456 VDD.n3238 VDD.t234 95.0005
R5457 VDD.n3328 VDD.t390 95.0005
R5458 VDD.t740 VDD.n1341 95.0005
R5459 VDD.t728 VDD.n1418 95.0005
R5460 VDD.t185 VDD.n1495 95.0005
R5461 VDD.t97 VDD.n1572 95.0005
R5462 VDD.t703 VDD.n1649 95.0005
R5463 VDD.t422 VDD.n1727 95.0005
R5464 VDD.n1809 VDD.t427 95.0005
R5465 VDD.n38 VDD.t437 94.7373
R5466 VDD.n178 VDD.t208 94.7373
R5467 VDD.n313 VDD.t683 94.7373
R5468 VDD.n456 VDD.t199 94.7373
R5469 VDD.n589 VDD.t148 94.7373
R5470 VDD.n724 VDD.t297 94.7373
R5471 VDD.n867 VDD.t49 94.7373
R5472 VDD.n2977 VDD.t171 93.9565
R5473 VDD.n3048 VDD.t74 93.9565
R5474 VDD.n2270 VDD.n2269 92.5005
R5475 VDD.n2280 VDD.n2248 92.5005
R5476 VDD.n2293 VDD.n2292 92.5005
R5477 VDD.n2237 VDD.n2236 92.5005
R5478 VDD.n2308 VDD.n2307 92.5005
R5479 VDD.n2318 VDD.n2230 92.5005
R5480 VDD.n2332 VDD.n2331 92.5005
R5481 VDD.n2355 VDD.n2223 92.5005
R5482 VDD.n2248 VDD.n2247 92.5005
R5483 VDD.n2292 VDD.n2291 92.5005
R5484 VDD.n2238 VDD.n2237 92.5005
R5485 VDD.n2309 VDD.n2308 92.5005
R5486 VDD.n2230 VDD.n2229 92.5005
R5487 VDD.n2331 VDD.n2330 92.5005
R5488 VDD.n2223 VDD.n2221 92.5005
R5489 VDD.n2271 VDD.n2270 92.5005
R5490 VDD.n2256 VDD.n2255 92.5005
R5491 VDD.n2351 VDD.n2335 92.5005
R5492 VDD.n2335 VDD.n2334 92.5005
R5493 VDD.n2350 VDD.n2349 92.5005
R5494 VDD.n2349 VDD.n2348 92.5005
R5495 VDD.n2337 VDD.n2336 92.5005
R5496 VDD.n2347 VDD.n2337 92.5005
R5497 VDD.n2345 VDD.n2344 92.5005
R5498 VDD.n2346 VDD.n2345 92.5005
R5499 VDD.n2343 VDD.n2339 92.5005
R5500 VDD.n2339 VDD.n2338 92.5005
R5501 VDD.n2342 VDD.n2341 92.5005
R5502 VDD.n2341 VDD.n2340 92.5005
R5503 VDD.n2364 VDD.n2363 92.5005
R5504 VDD.n2207 VDD.n2206 92.5005
R5505 VDD.n2379 VDD.n2378 92.5005
R5506 VDD.n2389 VDD.n2200 92.5005
R5507 VDD.n2400 VDD.n2399 92.5005
R5508 VDD.n2187 VDD.n2186 92.5005
R5509 VDD.n2415 VDD.n2414 92.5005
R5510 VDD.n2425 VDD.n2180 92.5005
R5511 VDD.n2439 VDD.n2438 92.5005
R5512 VDD.n2363 VDD.n2362 92.5005
R5513 VDD.n2208 VDD.n2207 92.5005
R5514 VDD.n2380 VDD.n2379 92.5005
R5515 VDD.n2200 VDD.n2198 92.5005
R5516 VDD.n2399 VDD.n2398 92.5005
R5517 VDD.n2188 VDD.n2187 92.5005
R5518 VDD.n2416 VDD.n2415 92.5005
R5519 VDD.n2180 VDD.n2178 92.5005
R5520 VDD.n2438 VDD.n2437 92.5005
R5521 VDD.n2443 VDD.n2442 92.5005
R5522 VDD.n2442 VDD.n2441 92.5005
R5523 VDD.n2444 VDD.n2169 92.5005
R5524 VDD.n2169 VDD.n2168 92.5005
R5525 VDD.n2452 VDD.n2167 92.5005
R5526 VDD.n2465 VDD.n2464 92.5005
R5527 VDD.n2155 VDD.n2154 92.5005
R5528 VDD.n2479 VDD.n2478 92.5005
R5529 VDD.n2489 VDD.n2147 92.5005
R5530 VDD.n2502 VDD.n2501 92.5005
R5531 VDD.n2135 VDD.n2134 92.5005
R5532 VDD.n2517 VDD.n2516 92.5005
R5533 VDD.n2527 VDD.n2127 92.5005
R5534 VDD.n2167 VDD.n2166 92.5005
R5535 VDD.n2464 VDD.n2463 92.5005
R5536 VDD.n2156 VDD.n2155 92.5005
R5537 VDD.n2480 VDD.n2479 92.5005
R5538 VDD.n2147 VDD.n2146 92.5005
R5539 VDD.n2501 VDD.n2500 92.5005
R5540 VDD.n2136 VDD.n2135 92.5005
R5541 VDD.n2518 VDD.n2517 92.5005
R5542 VDD.n2127 VDD.n2126 92.5005
R5543 VDD.n2531 VDD.n2125 92.5005
R5544 VDD.n2125 VDD.n2124 92.5005
R5545 VDD.n2533 VDD.n2532 92.5005
R5546 VDD.n2534 VDD.n2533 92.5005
R5547 VDD.n2123 VDD.n2122 92.5005
R5548 VDD.n2535 VDD.n2123 92.5005
R5549 VDD.n2538 VDD.n2537 92.5005
R5550 VDD.n2537 VDD.n2536 92.5005
R5551 VDD.n2539 VDD.n2121 92.5005
R5552 VDD.n2121 VDD.n2120 92.5005
R5553 VDD.n2541 VDD.n2540 92.5005
R5554 VDD.n2542 VDD.n2541 92.5005
R5555 VDD.n2545 VDD.n2544 92.5005
R5556 VDD.n2555 VDD.n2114 92.5005
R5557 VDD.n2568 VDD.n2567 92.5005
R5558 VDD.n2570 VDD.n2101 92.5005
R5559 VDD.n2583 VDD.n2582 92.5005
R5560 VDD.n2593 VDD.n2094 92.5005
R5561 VDD.n2604 VDD.n2603 92.5005
R5562 VDD.n2607 VDD.n2087 92.5005
R5563 VDD.n2620 VDD.n2079 92.5005
R5564 VDD.n2546 VDD.n2545 92.5005
R5565 VDD.n2114 VDD.n2112 92.5005
R5566 VDD.n2567 VDD.n2566 92.5005
R5567 VDD.n2102 VDD.n2101 92.5005
R5568 VDD.n2584 VDD.n2583 92.5005
R5569 VDD.n2094 VDD.n2092 92.5005
R5570 VDD.n2603 VDD.n2602 92.5005
R5571 VDD.n2087 VDD.n2085 92.5005
R5572 VDD.n2079 VDD.n2078 92.5005
R5573 VDD.n2628 VDD.n2074 92.5005
R5574 VDD.n2074 VDD.n2073 92.5005
R5575 VDD.n2636 VDD.n2072 92.5005
R5576 VDD.n2650 VDD.n2649 92.5005
R5577 VDD.n2060 VDD.n2059 92.5005
R5578 VDD.n2664 VDD.n2663 92.5005
R5579 VDD.n2674 VDD.n2052 92.5005
R5580 VDD.n2687 VDD.n2686 92.5005
R5581 VDD.n2040 VDD.n2039 92.5005
R5582 VDD.n2702 VDD.n2701 92.5005
R5583 VDD.n2712 VDD.n2032 92.5005
R5584 VDD.n2072 VDD.n2071 92.5005
R5585 VDD.n2649 VDD.n2648 92.5005
R5586 VDD.n2061 VDD.n2060 92.5005
R5587 VDD.n2665 VDD.n2664 92.5005
R5588 VDD.n2052 VDD.n2051 92.5005
R5589 VDD.n2686 VDD.n2685 92.5005
R5590 VDD.n2041 VDD.n2040 92.5005
R5591 VDD.n2703 VDD.n2702 92.5005
R5592 VDD.n2032 VDD.n2031 92.5005
R5593 VDD.n2716 VDD.n2030 92.5005
R5594 VDD.n2030 VDD.n2029 92.5005
R5595 VDD.n2718 VDD.n2717 92.5005
R5596 VDD.n2719 VDD.n2718 92.5005
R5597 VDD.n2028 VDD.n2027 92.5005
R5598 VDD.n2720 VDD.n2028 92.5005
R5599 VDD.n2723 VDD.n2722 92.5005
R5600 VDD.n2722 VDD.n2721 92.5005
R5601 VDD.n2724 VDD.n2026 92.5005
R5602 VDD.n2026 VDD.n2025 92.5005
R5603 VDD.n2727 VDD.n2726 92.5005
R5604 VDD.n2728 VDD.n2727 92.5005
R5605 VDD.n2725 VDD.n2024 92.5005
R5606 VDD.n2729 VDD.n2024 92.5005
R5607 VDD.n2763 VDD.n2762 92.5005
R5608 VDD.n2762 VDD.n2761 92.5005
R5609 VDD.n2014 VDD.n2010 92.5005
R5610 VDD.n2760 VDD.n2010 92.5005
R5611 VDD.n2758 VDD.n2757 92.5005
R5612 VDD.n2759 VDD.n2758 92.5005
R5613 VDD.n2750 VDD.n2011 92.5005
R5614 VDD.n2746 VDD.n2011 92.5005
R5615 VDD.n2749 VDD.n2748 92.5005
R5616 VDD.n2748 VDD.n2747 92.5005
R5617 VDD.n2021 VDD.n2018 92.5005
R5618 VDD.n2745 VDD.n2018 92.5005
R5619 VDD.n2743 VDD.n2742 92.5005
R5620 VDD.n2744 VDD.n2743 92.5005
R5621 VDD.n2736 VDD.n2019 92.5005
R5622 VDD.n2730 VDD.n2019 92.5005
R5623 VDD.n2733 VDD.n2732 92.5005
R5624 VDD.n2732 VDD.n2731 92.5005
R5625 VDD.n2764 VDD.n2007 92.5005
R5626 VDD.n2007 VDD.n2006 92.5005
R5627 VDD.n2772 VDD.n2005 92.5005
R5628 VDD.n2786 VDD.n2785 92.5005
R5629 VDD.n1993 VDD.n1992 92.5005
R5630 VDD.n2800 VDD.n2799 92.5005
R5631 VDD.n2810 VDD.n1985 92.5005
R5632 VDD.n2823 VDD.n2822 92.5005
R5633 VDD.n1973 VDD.n1972 92.5005
R5634 VDD.n2838 VDD.n2837 92.5005
R5635 VDD.n2848 VDD.n1965 92.5005
R5636 VDD.n2005 VDD.n2004 92.5005
R5637 VDD.n2785 VDD.n2784 92.5005
R5638 VDD.n1994 VDD.n1993 92.5005
R5639 VDD.n2801 VDD.n2800 92.5005
R5640 VDD.n1985 VDD.n1984 92.5005
R5641 VDD.n2822 VDD.n2821 92.5005
R5642 VDD.n1974 VDD.n1973 92.5005
R5643 VDD.n2839 VDD.n2838 92.5005
R5644 VDD.n1965 VDD.n1964 92.5005
R5645 VDD.n2852 VDD.n1963 92.5005
R5646 VDD.n1963 VDD.n1962 92.5005
R5647 VDD.n2854 VDD.n2853 92.5005
R5648 VDD.n2855 VDD.n2854 92.5005
R5649 VDD.n1961 VDD.n1960 92.5005
R5650 VDD.n2856 VDD.n1961 92.5005
R5651 VDD.n2859 VDD.n2858 92.5005
R5652 VDD.n2858 VDD.n2857 92.5005
R5653 VDD.n2860 VDD.n1959 92.5005
R5654 VDD.n1959 VDD.n1958 92.5005
R5655 VDD.n2863 VDD.n2862 92.5005
R5656 VDD.n2864 VDD.n2863 92.5005
R5657 VDD.n2861 VDD.n1957 92.5005
R5658 VDD.n2865 VDD.n1957 92.5005
R5659 VDD.n2899 VDD.n2898 92.5005
R5660 VDD.n2898 VDD.n2897 92.5005
R5661 VDD.n1946 VDD.n1945 92.5005
R5662 VDD.n2896 VDD.n1946 92.5005
R5663 VDD.n2894 VDD.n2893 92.5005
R5664 VDD.n2895 VDD.n2894 92.5005
R5665 VDD.n1948 VDD.n1947 92.5005
R5666 VDD.n2882 VDD.n1947 92.5005
R5667 VDD.n2885 VDD.n2884 92.5005
R5668 VDD.n2884 VDD.n2883 92.5005
R5669 VDD.n1954 VDD.n1951 92.5005
R5670 VDD.n2881 VDD.n1951 92.5005
R5671 VDD.n2879 VDD.n2878 92.5005
R5672 VDD.n2880 VDD.n2879 92.5005
R5673 VDD.n2872 VDD.n1952 92.5005
R5674 VDD.n2866 VDD.n1952 92.5005
R5675 VDD.n2869 VDD.n2868 92.5005
R5676 VDD.n2868 VDD.n2867 92.5005
R5677 VDD.n1941 VDD.n1940 92.5005
R5678 VDD.n1940 VDD.n1939 92.5005
R5679 VDD.n1924 VDD.n1923 92.5005
R5680 VDD.n2926 VDD.n1924 92.5005
R5681 VDD.n1912 VDD.n1910 92.5005
R5682 VDD.n2950 VDD.n1912 92.5005
R5683 VDD.n1893 VDD.n1888 92.5005
R5684 VDD.n2976 VDD.n1893 92.5005
R5685 VDD.n2979 VDD.n2978 92.5005
R5686 VDD.n2978 VDD.n2977 92.5005
R5687 VDD.n1898 VDD.n1892 92.5005
R5688 VDD.n2975 VDD.n1892 92.5005
R5689 VDD.n2973 VDD.n2972 92.5005
R5690 VDD.n2974 VDD.n2973 92.5005
R5691 VDD.n2966 VDD.n1895 92.5005
R5692 VDD.n1895 VDD.n1894 92.5005
R5693 VDD.n2965 VDD.n2964 92.5005
R5694 VDD.n2964 VDD.n2963 92.5005
R5695 VDD.n1905 VDD.n1901 92.5005
R5696 VDD.n2962 VDD.n1901 92.5005
R5697 VDD.n1909 VDD.n1902 92.5005
R5698 VDD.n2949 VDD.n1902 92.5005
R5699 VDD.n2960 VDD.n2959 92.5005
R5700 VDD.n2961 VDD.n2960 92.5005
R5701 VDD.n1881 VDD.n1880 92.5005
R5702 VDD.n2996 VDD.n1881 92.5005
R5703 VDD.n2994 VDD.n2993 92.5005
R5704 VDD.n2995 VDD.n2994 92.5005
R5705 VDD.n2992 VDD.n1883 92.5005
R5706 VDD.n1883 VDD.n1882 92.5005
R5707 VDD.n2991 VDD.n2990 92.5005
R5708 VDD.n2990 VDD.n2989 92.5005
R5709 VDD.n2986 VDD.n2985 92.5005
R5710 VDD.n2987 VDD.n2986 92.5005
R5711 VDD.n1885 VDD.n1884 92.5005
R5712 VDD.n2988 VDD.n1885 92.5005
R5713 VDD.n2984 VDD.n1887 92.5005
R5714 VDD.n1887 VDD.n1886 92.5005
R5715 VDD.n3022 VDD.n1868 92.5005
R5716 VDD.n3022 VDD.n3021 92.5005
R5717 VDD.n1851 VDD.n1846 92.5005
R5718 VDD.n3047 VDD.n1851 92.5005
R5719 VDD.n3050 VDD.n3049 92.5005
R5720 VDD.n3049 VDD.n3048 92.5005
R5721 VDD.n1856 VDD.n1850 92.5005
R5722 VDD.n3046 VDD.n1850 92.5005
R5723 VDD.n3044 VDD.n3043 92.5005
R5724 VDD.n3045 VDD.n3044 92.5005
R5725 VDD.n3037 VDD.n1853 92.5005
R5726 VDD.n1853 VDD.n1852 92.5005
R5727 VDD.n3036 VDD.n3035 92.5005
R5728 VDD.n3035 VDD.n3034 92.5005
R5729 VDD.n1863 VDD.n1859 92.5005
R5730 VDD.n3033 VDD.n1859 92.5005
R5731 VDD.n1867 VDD.n1860 92.5005
R5732 VDD.n3020 VDD.n1860 92.5005
R5733 VDD.n3031 VDD.n3030 92.5005
R5734 VDD.n3032 VDD.n3031 92.5005
R5735 VDD.n1839 VDD.n1838 92.5005
R5736 VDD.n3067 VDD.n1839 92.5005
R5737 VDD.n3065 VDD.n3064 92.5005
R5738 VDD.n3066 VDD.n3065 92.5005
R5739 VDD.n3063 VDD.n1841 92.5005
R5740 VDD.n1841 VDD.n1840 92.5005
R5741 VDD.n3062 VDD.n3061 92.5005
R5742 VDD.n3061 VDD.n3060 92.5005
R5743 VDD.n1843 VDD.n1842 92.5005
R5744 VDD.n3059 VDD.n1843 92.5005
R5745 VDD.n3057 VDD.n3056 92.5005
R5746 VDD.n3058 VDD.n3057 92.5005
R5747 VDD.n3055 VDD.n1845 92.5005
R5748 VDD.n1845 VDD.n1844 92.5005
R5749 VDD.n953 VDD.t601 92.1058
R5750 VDD.n1802 VDD.t478 91.4648
R5751 VDD.n1020 VDD.t381 91.4648
R5752 VDD.n1044 VDD.t203 91.4648
R5753 VDD.n1063 VDD.t491 91.4648
R5754 VDD.n1087 VDD.t32 91.4648
R5755 VDD.n1105 VDD.t147 91.4648
R5756 VDD.n1129 VDD.t89 91.4648
R5757 VDD.n1147 VDD.t145 91.4648
R5758 VDD.n1171 VDD.t629 91.4648
R5759 VDD.n1189 VDD.t91 91.4648
R5760 VDD.n1213 VDD.t36 91.4648
R5761 VDD.n1231 VDD.t597 91.4648
R5762 VDD.n1255 VDD.t600 91.4648
R5763 VDD.n1273 VDD.t631 91.4648
R5764 VDD.n237 VDD.t521 91.4648
R5765 VDD.n97 VDD.t542 91.4648
R5766 VDD.n926 VDD.t533 91.4648
R5767 VDD.n876 VDD.t551 91.4648
R5768 VDD.n783 VDD.t530 91.4648
R5769 VDD.n733 VDD.t509 91.4648
R5770 VDD.n648 VDD.t539 91.4648
R5771 VDD.n598 VDD.t527 91.4648
R5772 VDD.n515 VDD.t497 91.4648
R5773 VDD.n465 VDD.t536 91.4648
R5774 VDD.n372 VDD.t515 91.4648
R5775 VDD.n322 VDD.t494 91.4648
R5776 VDD.n47 VDD.t506 91.4648
R5777 VDD.n187 VDD.t503 91.4648
R5778 VDD.n2744 VDD.t439 88.7368
R5779 VDD.n2880 VDD.t86 88.7368
R5780 VDD.n1318 VDD.t630 87.0838
R5781 VDD.n1395 VDD.t596 87.0838
R5782 VDD.n1472 VDD.t90 87.0838
R5783 VDD.n1549 VDD.t144 87.0838
R5784 VDD.n1626 VDD.t146 87.0838
R5785 VDD.n1703 VDD.t490 87.0838
R5786 VDD.t380 VDD.n1773 87.0838
R5787 VDD.n98 VDD.t541 86.8426
R5788 VDD.n238 VDD.t520 86.8426
R5789 VDD.n373 VDD.t514 86.8426
R5790 VDD.n516 VDD.t496 86.8426
R5791 VDD.n649 VDD.t538 86.8426
R5792 VDD.n784 VDD.t529 86.8426
R5793 VDD.n927 VDD.t532 86.8426
R5794 VDD.n2228 VDD.t453 86.7743
R5795 VDD.n2209 VDD.t355 86.7743
R5796 VDD.n2137 VDD.t103 86.7743
R5797 VDD.n2560 VDD.t455 86.7743
R5798 VDD.n2042 VDD.t302 86.7743
R5799 VDD.n2734 VDD.t440 86.7743
R5800 VDD.n1975 VDD.t322 86.7743
R5801 VDD.n2870 VDD.t87 86.7743
R5802 VDD.n1930 VDD.t556 86.7743
R5803 VDD.n1920 VDD.t591 86.7743
R5804 VDD.n1890 VDD.t672 86.7743
R5805 VDD.n1877 VDD.t160 86.7743
R5806 VDD.n1848 VDD.t432 86.7743
R5807 VDD.n1835 VDD.t178 86.7743
R5808 VDD.n1802 VDD.t51 86.7743
R5809 VDD.n1011 VDD.t53 86.7743
R5810 VDD.n1044 VDD.t193 86.7743
R5811 VDD.n1053 VDD.t195 86.7743
R5812 VDD.n1087 VDD.t457 86.7743
R5813 VDD.n1095 VDD.t459 86.7743
R5814 VDD.n1129 VDD.t334 86.7743
R5815 VDD.n1137 VDD.t332 86.7743
R5816 VDD.n1171 VDD.t708 86.7743
R5817 VDD.n1179 VDD.t706 86.7743
R5818 VDD.n1213 VDD.t254 86.7743
R5819 VDD.n1221 VDD.t252 86.7743
R5820 VDD.n1255 VDD.t371 86.7743
R5821 VDD.n1263 VDD.t373 86.7743
R5822 VDD.n211 VDD.t444 86.7743
R5823 VDD.n71 VDD.t152 86.7743
R5824 VDD.n900 VDD.t336 86.7743
R5825 VDD.n876 VDD.t338 86.7743
R5826 VDD.n757 VDD.t63 86.7743
R5827 VDD.n733 VDD.t65 86.7743
R5828 VDD.n622 VDD.t40 86.7743
R5829 VDD.n598 VDD.t42 86.7743
R5830 VDD.n489 VDD.t724 86.7743
R5831 VDD.n465 VDD.t726 86.7743
R5832 VDD.n346 VDD.t562 86.7743
R5833 VDD.n322 VDD.t560 86.7743
R5834 VDD.n47 VDD.t154 86.7743
R5835 VDD.n187 VDD.t442 86.7743
R5836 VDD.t378 VDD.n2466 86.1269
R5837 VDD.n3239 VDD.t216 84.4449
R5838 VDD.t692 VDD.n3262 84.4449
R5839 VDD.n3286 VDD.t745 84.4449
R5840 VDD.n3329 VDD.t386 84.4449
R5841 VDD.t609 VDD.n3352 84.4449
R5842 VDD.n3376 VDD.t366 84.4449
R5843 VDD.n123 VDD.t33 84.211
R5844 VDD.n398 VDD.t12 84.211
R5845 VDD.n534 VDD.t29 84.211
R5846 VDD.n667 VDD.t479 84.211
R5847 VDD.n809 VDD.t17 84.211
R5848 VDD.n2268 VDD.t684 83.517
R5849 VDD.t473 VDD.n2243 83.517
R5850 VDD.t671 VDD.n2975 83.517
R5851 VDD.t431 VDD.n3046 83.517
R5852 VDD.t661 VDD 81.5794
R5853 VDD VDD.t173 81.5794
R5854 VDD.t92 VDD 81.5794
R5855 VDD VDD.t420 81.5794
R5856 VDD VDD.t288 81.5794
R5857 VDD VDD.t10 81.5794
R5858 VDD VDD.t98 81.5794
R5859 VDD.n3090 VDD 81.5278
R5860 VDD.n2477 VDD.t470 80.9071
R5861 VDD VDD.n2066 80.9071
R5862 VDD VDD.n1999 80.9071
R5863 VDD.n2637 VDD.t276 78.2972
R5864 VDD.n2773 VDD.t23 78.2972
R5865 VDD.n2906 VDD 78.2972
R5866 VDD.n1027 VDD 78.1104
R5867 VDD.n1678 VDD 78.1104
R5868 VDD.n1601 VDD 78.1104
R5869 VDD.n1524 VDD 78.1104
R5870 VDD.n1447 VDD 78.1104
R5871 VDD.n1370 VDD 78.1104
R5872 VDD.n1293 VDD 78.1104
R5873 VDD.t232 VDD.n3214 77.5227
R5874 VDD.t392 VDD.n3304 77.5227
R5875 VDD.n3237 VDD.t222 73.8894
R5876 VDD.n3327 VDD.t406 73.8894
R5877 VDD.t370 VDD.n1340 73.8894
R5878 VDD.t253 VDD.n1417 73.8894
R5879 VDD.t707 VDD.n1494 73.8894
R5880 VDD.t333 VDD.n1571 73.8894
R5881 VDD.t456 VDD.n1648 73.8894
R5882 VDD.t192 VDD.n1725 73.8894
R5883 VDD.n1797 VDD.t50 73.8894
R5884 VDD.n2652 VDD.t488 73.0774
R5885 VDD.n2788 VDD.t132 73.0774
R5886 VDD.n2951 VDD 73.0774
R5887 VDD.n3019 VDD 73.0774
R5888 VDD.n1307 VDD.t56 71.2505
R5889 VDD.n1384 VDD.t738 71.2505
R5890 VDD.n1461 VDD.t575 71.2505
R5891 VDD.n1538 VDD.t675 71.2505
R5892 VDD.n1615 VDD.t719 71.2505
R5893 VDD.n1692 VDD.t329 71.2505
R5894 VDD.n1772 VDD.t665 71.2505
R5895 VDD.n107 VDD.t313 71.0531
R5896 VDD.n247 VDD.t358 71.0531
R5897 VDD.n382 VDD.t105 71.0531
R5898 VDD.n525 VDD.t433 71.0531
R5899 VDD.n658 VDD.t636 71.0531
R5900 VDD.n793 VDD.t21 71.0531
R5901 VDD.n936 VDD.t319 71.0531
R5902 VDD.t466 VDD.n2411 70.4675
R5903 VDD.n2594 VDD.t471 70.4675
R5904 VDD.n2907 VDD.t677 70.4675
R5905 VDD.t352 VDD.n2947 70.4675
R5906 VDD.t686 VDD.n3017 70.4675
R5907 VDD.t484 VDD.n3088 70.4675
R5908 VDD.n2228 VDD.t256 68.0124
R5909 VDD.n2209 VDD.t15 68.0124
R5910 VDD.n2137 VDD.t660 68.0124
R5911 VDD.n2560 VDD.t375 68.0124
R5912 VDD.n2042 VDD.t162 68.0124
R5913 VDD.n2734 VDD.t77 68.0124
R5914 VDD.n1975 VDD.t385 68.0124
R5915 VDD.n2870 VDD.t268 68.0124
R5916 VDD.n1930 VDD.t426 68.0124
R5917 VDD.n1920 VDD.t680 68.0124
R5918 VDD.n1890 VDD.t172 68.0124
R5919 VDD.n1877 VDD.t357 68.0124
R5920 VDD.n1848 VDD.t75 68.0124
R5921 VDD.n1835 VDD.t483 68.0124
R5922 VDD.t238 VDD.n3249 63.3338
R5923 VDD.n3263 VDD.t698 63.3338
R5924 VDD.n3285 VDD.t747 63.3338
R5925 VDD.t400 VDD.n3339 63.3338
R5926 VDD.n3353 VDD.t605 63.3338
R5927 VDD.n3375 VDD.t362 63.3338
R5928 VDD.n1760 VDD.t548 63.1021
R5929 VDD.n1679 VDD.t518 63.1021
R5930 VDD.n1602 VDD.t524 63.1021
R5931 VDD.n1525 VDD.t545 63.1021
R5932 VDD.n1448 VDD.t554 63.1021
R5933 VDD.n1371 VDD.t500 63.1021
R5934 VDD.n1294 VDD.t512 63.1021
R5935 VDD.n269 VDD.t595 63.1021
R5936 VDD.n130 VDD.t34 63.1021
R5937 VDD.n405 VDD.t13 63.1021
R5938 VDD.n539 VDD.t30 63.1021
R5939 VDD.n673 VDD.t480 63.1021
R5940 VDD.n816 VDD.t18 63.1021
R5941 VDD.n962 VDD.t602 63.1021
R5942 VDD.t472 VDD.n2746 62.6379
R5943 VDD.t469 VDD.n2882 62.6379
R5944 VDD.n136 VDD.n133 60.0005
R5945 VDD.n263 VDD.n260 60.0005
R5946 VDD.n1284 VDD.t164 58.4849
R5947 VDD.n1242 VDD.t262 58.4849
R5948 VDD.n1200 VDD.t308 58.4849
R5949 VDD.n1158 VDD.t620 58.4849
R5950 VDD.n1116 VDD.t641 58.4849
R5951 VDD.n1074 VDD.t568 58.4849
R5952 VDD.n1034 VDD.t649 58.4849
R5953 VDD.n149 VDD.t122 58.4849
R5954 VDD.n984 VDD.t180 58.4849
R5955 VDD.n838 VDD.t716 58.4849
R5956 VDD.n695 VDD.t85 58.4849
R5957 VDD.n560 VDD.t731 58.4849
R5958 VDD.n427 VDD.t291 58.4849
R5959 VDD.n283 VDD.t585 58.4849
R5960 VDD.n2317 VDD.t452 57.4181
R5961 VDD.n2963 VDD.t463 57.4181
R5962 VDD.n3034 VDD.t462 57.4181
R5963 VDD.n2638 VDD.n2072 56.4711
R5964 VDD.n2649 VDD.n2065 56.4711
R5965 VDD.n2660 VDD.n2060 56.4711
R5966 VDD.n2664 VDD.n2054 56.4711
R5967 VDD.n2676 VDD.n2052 56.4711
R5968 VDD.n2686 VDD.n2046 56.4711
R5969 VDD.n2698 VDD.n2040 56.4711
R5970 VDD.n2702 VDD.n2034 56.4711
R5971 VDD.n2714 VDD.n2032 56.4711
R5972 VDD.n2774 VDD.n2005 56.4711
R5973 VDD.n2785 VDD.n1998 56.4711
R5974 VDD.n2796 VDD.n1993 56.4711
R5975 VDD.n2800 VDD.n1987 56.4711
R5976 VDD.n2812 VDD.n1985 56.4711
R5977 VDD.n2822 VDD.n1979 56.4711
R5978 VDD.n2834 VDD.n1973 56.4711
R5979 VDD.n2838 VDD.n1967 56.4711
R5980 VDD.n2850 VDD.n1965 56.4711
R5981 VDD.n2270 VDD.n2253 56.4711
R5982 VDD.n2278 VDD.n2248 56.4711
R5983 VDD.n2292 VDD.n2244 56.4711
R5984 VDD.n2296 VDD.n2237 56.4711
R5985 VDD.n2308 VDD.n2235 56.4711
R5986 VDD.n2316 VDD.n2230 56.4711
R5987 VDD.n2331 VDD.n2225 56.4711
R5988 VDD.n2357 VDD.n2223 56.4711
R5989 VDD.n806 VDD.n805 56.4711
R5990 VDD.n820 VDD.n819 56.4711
R5991 VDD.n678 VDD.n677 56.4711
R5992 VDD.n544 VDD.n543 56.4711
R5993 VDD.n395 VDD.n394 56.4711
R5994 VDD.n410 VDD.n409 56.4711
R5995 VDD.n120 VDD.n119 56.4711
R5996 VDD.n967 VDD.n966 54.8576
R5997 VDD.n2504 VDD.t102 54.8082
R5998 VDD.n2450 VDD.n2167 52.9417
R5999 VDD.n2464 VDD.n2162 52.9417
R6000 VDD.n2468 VDD.n2155 52.9417
R6001 VDD.n2479 VDD.n2153 52.9417
R6002 VDD.n2487 VDD.n2147 52.9417
R6003 VDD.n2501 VDD.n2143 52.9417
R6004 VDD.n2505 VDD.n2135 52.9417
R6005 VDD.n2517 VDD.n2133 52.9417
R6006 VDD.n2525 VDD.n2127 52.9417
R6007 VDD.n3216 VDD.t220 52.7783
R6008 VDD.t236 VDD.n3226 52.7783
R6009 VDD.n3306 VDD.t414 52.7783
R6010 VDD.t394 VDD.n3316 52.7783
R6011 VDD.t623 VDD 52.1983
R6012 VDD VDD.t340 52.1983
R6013 VDD VDD.t286 52.1983
R6014 VDD VDD.t448 52.1983
R6015 VDD VDD.t446 52.1983
R6016 VDD VDD.t299 52.1983
R6017 VDD VDD.t43 52.1983
R6018 VDD.n134 VDD.t117 50.0005
R6019 VDD.n411 VDD.t292 50.0005
R6020 VDD.n679 VDD.t82 50.0005
R6021 VDD.n968 VDD.t183 47.3689
R6022 VDD.t255 VDD.n2224 46.9785
R6023 VDD.n3298 VDD 44.8616
R6024 VDD.n3388 VDD 44.8616
R6025 VDD.n135 VDD.n134 44.7373
R6026 VDD.n262 VDD.n261 44.7373
R6027 VDD.n950 VDD.n949 44.5719
R6028 VDD.n2377 VDD.t354 44.3686
R6029 VDD.n2515 VDD.t659 44.3686
R6030 VDD.t454 VDD.n2569 44.3686
R6031 VDD.n2662 VDD.t475 44.3686
R6032 VDD.n2798 VDD.t468 44.3686
R6033 VDD.t228 VDD.n3250 42.2227
R6034 VDD.n3261 VDD.t694 42.2227
R6035 VDD VDD.n3273 42.2227
R6036 VDD.t743 VDD.n3274 42.2227
R6037 VDD.n3287 VDD 42.2227
R6038 VDD.t410 VDD.n3340 42.2227
R6039 VDD.n3351 VDD.t611 42.2227
R6040 VDD VDD.n3363 42.2227
R6041 VDD.t364 VDD.n3364 42.2227
R6042 VDD.n3377 VDD 42.2227
R6043 VDD.n122 VDD.n121 42.1058
R6044 VDD.n397 VDD.n396 42.1058
R6045 VDD.n412 VDD.n411 42.1058
R6046 VDD.n546 VDD.n545 42.1058
R6047 VDD.n680 VDD.n679 42.1058
R6048 VDD.n808 VDD.n807 42.1058
R6049 VDD.n822 VDD.n821 42.1058
R6050 VDD.n969 VDD.n968 42.1058
R6051 VDD.n2269 VDD.n2267 41.7587
R6052 VDD.n2280 VDD.n2279 41.7587
R6053 VDD.n2293 VDD.n2243 41.7587
R6054 VDD.n2295 VDD.n2236 41.7587
R6055 VDD.n2307 VDD.n2305 41.7587
R6056 VDD.n2318 VDD.n2317 41.7587
R6057 VDD.n2332 VDD.n2224 41.7587
R6058 VDD.n2356 VDD.n2355 41.7587
R6059 VDD.n2453 VDD.t187 41.7587
R6060 VDD.n2637 VDD.n2636 41.7587
R6061 VDD.n2651 VDD.n2650 41.7587
R6062 VDD.n2661 VDD.n2059 41.7587
R6063 VDD.n2663 VDD.n2053 41.7587
R6064 VDD.n2675 VDD.n2674 41.7587
R6065 VDD.n2699 VDD.n2039 41.7587
R6066 VDD.n2701 VDD.n2033 41.7587
R6067 VDD.n2713 VDD.n2712 41.7587
R6068 VDD.n2773 VDD.n2772 41.7587
R6069 VDD.n2787 VDD.n2786 41.7587
R6070 VDD.n2797 VDD.n1992 41.7587
R6071 VDD.n2799 VDD.n1986 41.7587
R6072 VDD.n2811 VDD.n2810 41.7587
R6073 VDD.n2835 VDD.n1972 41.7587
R6074 VDD.n2837 VDD.n1966 41.7587
R6075 VDD.n2849 VDD.n2848 41.7587
R6076 VDD.t474 VDD.n1933 41.7587
R6077 VDD.n2938 VDD.t465 41.7587
R6078 VDD.n3008 VDD.t464 41.7587
R6079 VDD.n3079 VDD.t467 41.7587
R6080 VDD.n994 VDD.t111 41.5552
R6081 VDD.n994 VDD.t211 41.5552
R6082 VDD.n1037 VDD.t157 41.5552
R6083 VDD.n1037 VDD.t578 41.5552
R6084 VDD.n1665 VDD.t114 41.5552
R6085 VDD.n1665 VDD.t275 41.5552
R6086 VDD.n1588 VDD.t143 41.5552
R6087 VDD.n1588 VDD.t201 41.5552
R6088 VDD.n1511 VDD.t325 41.5552
R6089 VDD.n1511 VDD.t664 41.5552
R6090 VDD.n1434 VDD.t582 41.5552
R6091 VDD.n1434 VDD.t670 41.5552
R6092 VDD.n1357 VDD.t128 41.5552
R6093 VDD.n1357 VDD.t419 41.5552
R6094 VDD.n14 VDD.t174 41.5552
R6095 VDD.n14 VDD.t279 41.5552
R6096 VDD.n0 VDD.t99 41.5552
R6097 VDD.n0 VDD.t60 41.5552
R6098 VDD.n3 VDD.t11 41.5552
R6099 VDD.n3 VDD.t7 41.5552
R6100 VDD.n6 VDD.t289 41.5552
R6101 VDD.n6 VDD.t205 41.5552
R6102 VDD.n9 VDD.t421 41.5552
R6103 VDD.n9 VDD.t653 41.5552
R6104 VDD.n12 VDD.t93 41.5552
R6105 VDD.n12 VDD.t138 41.5552
R6106 VDD.n17 VDD.t662 41.5552
R6107 VDD.n17 VDD.t26 41.5552
R6108 VDD.t212 VDD.n2266 39.1488
R6109 VDD.n2452 VDD.n2451 39.1488
R6110 VDD.n2465 VDD.n2161 39.1488
R6111 VDD.n2467 VDD.n2154 39.1488
R6112 VDD.n2478 VDD.n2477 39.1488
R6113 VDD.n2489 VDD.n2488 39.1488
R6114 VDD.n2502 VDD.n2142 39.1488
R6115 VDD.n2504 VDD.n2134 39.1488
R6116 VDD.n2516 VDD.n2515 39.1488
R6117 VDD.n2527 VDD.n2526 39.1488
R6118 VDD.n2363 VDD.n2215 38.824
R6119 VDD.n2374 VDD.n2207 38.824
R6120 VDD.n2379 VDD.n2201 38.824
R6121 VDD.n2391 VDD.n2200 38.824
R6122 VDD.n2399 VDD.n2193 38.824
R6123 VDD.n2410 VDD.n2187 38.824
R6124 VDD.n2415 VDD.n2181 38.824
R6125 VDD.n2427 VDD.n2180 38.824
R6126 VDD.n2438 VDD.n2172 38.824
R6127 VDD.n2545 VDD.n2116 38.824
R6128 VDD.n2557 VDD.n2114 38.824
R6129 VDD.n2567 VDD.n2107 38.824
R6130 VDD.n2579 VDD.n2101 38.824
R6131 VDD.n2583 VDD.n2096 38.824
R6132 VDD.n2595 VDD.n2094 38.824
R6133 VDD.n2603 VDD.n2086 38.824
R6134 VDD.n2087 VDD.n2080 38.824
R6135 VDD.n2622 VDD.n2079 38.824
R6136 VDD.n1011 VDD.t668 38.6969
R6137 VDD.n1053 VDD.t328 38.6969
R6138 VDD.n1095 VDD.t722 38.6969
R6139 VDD.n1137 VDD.t674 38.6969
R6140 VDD.n1179 VDD.t574 38.6969
R6141 VDD.n1221 VDD.t737 38.6969
R6142 VDD.n1263 VDD.t55 38.6969
R6143 VDD.n211 VDD.t361 38.6969
R6144 VDD.n71 VDD.t316 38.6969
R6145 VDD.n900 VDD.t318 38.6969
R6146 VDD.n757 VDD.t20 38.6969
R6147 VDD.n622 VDD.t635 38.6969
R6148 VDD.n489 VDD.t436 38.6969
R6149 VDD.n346 VDD.t108 38.6969
R6150 VDD.t599 VDD.n1339 36.9449
R6151 VDD.t35 VDD.n1416 36.9449
R6152 VDD.t628 VDD.n1493 36.9449
R6153 VDD.t88 VDD.n1570 36.9449
R6154 VDD.t31 VDD.n1647 36.9449
R6155 VDD.t202 VDD.n1724 36.9449
R6156 VDD.n1798 VDD.t477 36.9449
R6157 VDD.n261 VDD.t594 36.8426
R6158 VDD VDD.t212 36.539
R6159 VDD.t187 VDD 36.539
R6160 VDD.t276 VDD 36.539
R6161 VDD.t23 VDD 36.539
R6162 VDD VDD.t657 36.539
R6163 VDD.t461 VDD.n2916 36.539
R6164 VDD.n2937 VDD.t273 36.539
R6165 VDD.n3007 VDD.t269 36.539
R6166 VDD.n3078 VDD.t460 36.539
R6167 VDD.n3154 VDD.t95 36.1587
R6168 VDD.n3154 VDD.t46 36.1587
R6169 VDD.n3094 VDD.t558 36.1587
R6170 VDD.n3094 VDD.t79 36.1587
R6171 VDD.n952 VDD.n951 34.211
R6172 VDD.t14 VDD.n2375 33.9291
R6173 VDD.n2556 VDD.t374 33.9291
R6174 VDD.n2759 VDD.t382 33.9291
R6175 VDD.n2895 VDD.t632 33.9291
R6176 VDD.n1284 VDD.t604 31.831
R6177 VDD.n1242 VDD.t310 31.831
R6178 VDD.n1200 VDD.t718 31.831
R6179 VDD.n1158 VDD.t377 31.831
R6180 VDD.n1116 VDD.t752 31.831
R6181 VDD.n1074 VDD.t656 31.831
R6182 VDD.n1034 VDD.t3 31.831
R6183 VDD.n149 VDD.t197 31.831
R6184 VDD.n984 VDD.t176 31.831
R6185 VDD.n838 VDD.t451 31.831
R6186 VDD.n695 VDD.t191 31.831
R6187 VDD.n560 VDD.t626 31.831
R6188 VDD.n427 VDD.t5 31.831
R6189 VDD.n283 VDD.t271 31.831
R6190 VDD.n3215 VDD.t246 31.6672
R6191 VDD.n3227 VDD.t226 31.6672
R6192 VDD.n3305 VDD.t402 31.6672
R6193 VDD.n3317 VDD.t408 31.6672
R6194 VDD.t272 VDD.n2687 31.3192
R6195 VDD.t351 VDD.n2823 31.3192
R6196 VDD.n2628 VDD.n2627 31.2934
R6197 VDD.n2165 VDD.t188 28.7575
R6198 VDD.n2257 VDD.t213 28.7575
R6199 VDD.n2177 VDD.t624 28.7575
R6200 VDD.n2081 VDD.t341 28.7575
R6201 VDD.n2070 VDD.t277 28.7575
R6202 VDD.n2013 VDD.t287 28.7575
R6203 VDD.n2003 VDD.t24 28.7575
R6204 VDD.n2890 VDD.t449 28.7575
R6205 VDD.n1942 VDD.t658 28.7575
R6206 VDD.n1907 VDD.t447 28.7575
R6207 VDD.n1904 VDD.t101 28.7575
R6208 VDD.n1865 VDD.t300 28.7575
R6209 VDD.n1862 VDD.t430 28.7575
R6210 VDD.n1825 VDD.t44 28.7575
R6211 VDD.n2365 VDD.n2364 28.7093
R6212 VDD.n2375 VDD.n2206 28.7093
R6213 VDD.n2378 VDD.n2377 28.7093
R6214 VDD.n2401 VDD.n2400 28.7093
R6215 VDD.n2411 VDD.n2186 28.7093
R6216 VDD.n2414 VDD.n2413 28.7093
R6217 VDD.n2426 VDD.n2425 28.7093
R6218 VDD.n2440 VDD.n2439 28.7093
R6219 VDD.n2544 VDD.n2115 28.7093
R6220 VDD.n2556 VDD.n2555 28.7093
R6221 VDD.n2569 VDD.n2568 28.7093
R6222 VDD.n2582 VDD.n2095 28.7093
R6223 VDD.n2594 VDD.n2593 28.7093
R6224 VDD.n2605 VDD.n2604 28.7093
R6225 VDD.n2607 VDD.n2606 28.7093
R6226 VDD.n2621 VDD.n2620 28.7093
R6227 VDD.t486 VDD.n2962 28.7093
R6228 VDD.t169 VDD.n3033 28.7093
R6229 VDD.n1760 VDD.t647 28.0332
R6230 VDD.n1679 VDD.t572 28.0332
R6231 VDD.n1602 VDD.t639 28.0332
R6232 VDD.n1525 VDD.t618 28.0332
R6233 VDD.n1448 VDD.t306 28.0332
R6234 VDD.n1371 VDD.t260 28.0332
R6235 VDD.n1294 VDD.t168 28.0332
R6236 VDD.n269 VDD.t589 28.0332
R6237 VDD.n130 VDD.t118 28.0332
R6238 VDD.n405 VDD.t293 28.0332
R6239 VDD.n539 VDD.t733 28.0332
R6240 VDD.n673 VDD.t83 28.0332
R6241 VDD.n816 VDD.t712 28.0332
R6242 VDD.n962 VDD.t184 28.0332
R6243 VDD.n3171 VDD.t693 26.5955
R6244 VDD.n3171 VDD.t697 26.5955
R6245 VDD.n3175 VDD.t695 26.5955
R6246 VDD.n3175 VDD.t699 26.5955
R6247 VDD.n3179 VDD.t225 26.5955
R6248 VDD.n3179 VDD.t701 26.5955
R6249 VDD.n3183 VDD.t229 26.5955
R6250 VDD.n3183 VDD.t241 26.5955
R6251 VDD.n3187 VDD.t217 26.5955
R6252 VDD.n3187 VDD.t239 26.5955
R6253 VDD.n3191 VDD.t219 26.5955
R6254 VDD.n3191 VDD.t245 26.5955
R6255 VDD.n3196 VDD.t223 26.5955
R6256 VDD.n3196 VDD.t235 26.5955
R6257 VDD.n3200 VDD.t227 26.5955
R6258 VDD.n3200 VDD.t237 26.5955
R6259 VDD.n3205 VDD.t231 26.5955
R6260 VDD.n3205 VDD.t243 26.5955
R6261 VDD.n3209 VDD.t221 26.5955
R6262 VDD.n3209 VDD.t247 26.5955
R6263 VDD.n3165 VDD.t748 26.5955
R6264 VDD.n3165 VDD.t746 26.5955
R6265 VDD.n3160 VDD.t750 26.5955
R6266 VDD.n3160 VDD.t1 26.5955
R6267 VDD.n3111 VDD.t610 26.5955
R6268 VDD.n3111 VDD.t616 26.5955
R6269 VDD.n3115 VDD.t612 26.5955
R6270 VDD.n3115 VDD.t606 26.5955
R6271 VDD.n3119 VDD.t417 26.5955
R6272 VDD.n3119 VDD.t608 26.5955
R6273 VDD.n3123 VDD.t411 26.5955
R6274 VDD.n3123 VDD.t397 26.5955
R6275 VDD.n3127 VDD.t387 26.5955
R6276 VDD.n3127 VDD.t401 26.5955
R6277 VDD.n3131 VDD.t389 26.5955
R6278 VDD.n3131 VDD.t405 26.5955
R6279 VDD.n3136 VDD.t407 26.5955
R6280 VDD.n3136 VDD.t391 26.5955
R6281 VDD.n3140 VDD.t409 26.5955
R6282 VDD.n3140 VDD.t395 26.5955
R6283 VDD.n3145 VDD.t413 26.5955
R6284 VDD.n3145 VDD.t399 26.5955
R6285 VDD.n3149 VDD.t415 26.5955
R6286 VDD.n3149 VDD.t403 26.5955
R6287 VDD.n3105 VDD.t363 26.5955
R6288 VDD.n3105 VDD.t367 26.5955
R6289 VDD.n3100 VDD.t369 26.5955
R6290 VDD.n3100 VDD.t71 26.5955
R6291 VDD.n2266 VDD.n2254 26.2219
R6292 VDD.n2255 VDD.n2254 26.1149
R6293 VDD.n2351 VDD.n2350 24.0332
R6294 VDD.n2350 VDD.n2336 24.0332
R6295 VDD.n2344 VDD.n2336 24.0332
R6296 VDD.n2344 VDD.n2343 24.0332
R6297 VDD.n2343 VDD.n2342 24.0332
R6298 VDD.n2444 VDD.n2443 24.0332
R6299 VDD.n2532 VDD.n2531 24.0332
R6300 VDD.n2532 VDD.n2122 24.0332
R6301 VDD.n2538 VDD.n2122 24.0332
R6302 VDD.n2539 VDD.n2538 24.0332
R6303 VDD.n2540 VDD.n2539 24.0332
R6304 VDD.n2717 VDD.n2716 24.0332
R6305 VDD.n2717 VDD.n2027 24.0332
R6306 VDD.n2723 VDD.n2027 24.0332
R6307 VDD.n2724 VDD.n2723 24.0332
R6308 VDD.n2726 VDD.n2724 24.0332
R6309 VDD.n2726 VDD.n2725 24.0332
R6310 VDD.n2853 VDD.n2852 24.0332
R6311 VDD.n2853 VDD.n1960 24.0332
R6312 VDD.n2859 VDD.n1960 24.0332
R6313 VDD.n2860 VDD.n2859 24.0332
R6314 VDD.n2862 VDD.n2860 24.0332
R6315 VDD.n2862 VDD.n2861 24.0332
R6316 VDD.n2985 VDD.n2984 24.0332
R6317 VDD.n2985 VDD.n1884 24.0332
R6318 VDD.n2991 VDD.n1884 24.0332
R6319 VDD.n2992 VDD.n2991 24.0332
R6320 VDD.n2993 VDD.n2992 24.0332
R6321 VDD.n2993 VDD.n1880 24.0332
R6322 VDD.n3056 VDD.n3055 24.0332
R6323 VDD.n3056 VDD.n1842 24.0332
R6324 VDD.n3062 VDD.n1842 24.0332
R6325 VDD.n3063 VDD.n3062 24.0332
R6326 VDD.n3064 VDD.n3063 24.0332
R6327 VDD.n3064 VDD.n1838 24.0332
R6328 VDD.n2764 VDD.n2763 23.7899
R6329 VDD.n2899 VDD.n1941 23.7899
R6330 VDD.n1321 VDD.t126 23.7505
R6331 VDD.n1398 VDD.t583 23.7505
R6332 VDD.n1475 VDD.t323 23.7505
R6333 VDD.n1552 VDD.t140 23.7505
R6334 VDD.n1629 VDD.t115 23.7505
R6335 VDD.n1706 VDD.t158 23.7505
R6336 VDD.t112 VDD.n1785 23.7505
R6337 VDD.n2259 VDD.n2254 23.7154
R6338 VDD.n1910 VDD.n1909 23.7089
R6339 VDD.n1868 VDD.n1867 23.7089
R6340 VDD.n89 VDD.t28 23.6847
R6341 VDD.n229 VDD.t281 23.6847
R6342 VDD.n364 VDD.t136 23.6847
R6343 VDD.n507 VDD.t651 23.6847
R6344 VDD.n640 VDD.t207 23.6847
R6345 VDD.n775 VDD.t9 23.6847
R6346 VDD.n918 VDD.t61 23.6847
R6347 VDD.n2352 VDD.n2351 23.245
R6348 VDD.n2531 VDD.n2530 22.9432
R6349 VDD.n2903 VDD.n1941 22.1686
R6350 VDD.n2930 VDD.n1923 22.1686
R6351 VDD.n2953 VDD.n1910 22.1686
R6352 VDD.n3000 VDD.n1880 22.1686
R6353 VDD.n3024 VDD.n1868 22.1686
R6354 VDD.n3071 VDD.n1838 22.1686
R6355 VDD.n2342 VDD.n2218 21.7362
R6356 VDD.n2540 VDD.n2118 21.7362
R6357 VDD.n2363 VDD.n2217 21.177
R6358 VDD.n2367 VDD.n2207 21.177
R6359 VDD.n2379 VDD.n2205 21.177
R6360 VDD.n2387 VDD.n2200 21.177
R6361 VDD.n2399 VDD.n2195 21.177
R6362 VDD.n2403 VDD.n2187 21.177
R6363 VDD.n2415 VDD.n2185 21.177
R6364 VDD.n2423 VDD.n2180 21.177
R6365 VDD.n2438 VDD.n2173 21.177
R6366 VDD.n2545 VDD.n2119 21.177
R6367 VDD.n2553 VDD.n2114 21.177
R6368 VDD.n2567 VDD.n2109 21.177
R6369 VDD.n2572 VDD.n2101 21.177
R6370 VDD.n2583 VDD.n2100 21.177
R6371 VDD.n2591 VDD.n2094 21.177
R6372 VDD.n2603 VDD.n2089 21.177
R6373 VDD.n2609 VDD.n2087 21.177
R6374 VDD.n2619 VDD.n2079 21.177
R6375 VDD.n3251 VDD.t240 21.1116
R6376 VDD.n3260 VDD.t700 21.1116
R6377 VDD.n3341 VDD.t396 21.1116
R6378 VDD.n3350 VDD.t607 21.1116
R6379 VDD.t350 VDD.n2389 20.8796
R6380 VDD.n2570 VDD.t598 20.8796
R6381 VDD VDD.n2961 20.8796
R6382 VDD VDD.n3032 20.8796
R6383 VDD.n3218 VDD.n3208 20.3039
R6384 VDD.n3222 VDD.n3204 20.3039
R6385 VDD.n3229 VDD.n3199 20.3039
R6386 VDD.n3235 VDD.n3195 20.3039
R6387 VDD.n3243 VDD.n3242 20.3039
R6388 VDD.n3247 VDD.n3189 20.3039
R6389 VDD.n3254 VDD.n3253 20.3039
R6390 VDD.n3258 VDD.n3181 20.3039
R6391 VDD.n3266 VDD.n3265 20.3039
R6392 VDD.n3277 VDD.n3167 20.3039
R6393 VDD.n3291 VDD.n3290 20.3039
R6394 VDD.n3308 VDD.n3148 20.3039
R6395 VDD.n3312 VDD.n3144 20.3039
R6396 VDD.n3319 VDD.n3139 20.3039
R6397 VDD.n3325 VDD.n3135 20.3039
R6398 VDD.n3333 VDD.n3332 20.3039
R6399 VDD.n3337 VDD.n3129 20.3039
R6400 VDD.n3344 VDD.n3343 20.3039
R6401 VDD.n3348 VDD.n3121 20.3039
R6402 VDD.n3356 VDD.n3355 20.3039
R6403 VDD.n3367 VDD.n3107 20.3039
R6404 VDD.n3381 VDD.n3380 20.3039
R6405 VDD.n2909 VDD.n1937 20.3039
R6406 VDD.n2909 VDD.n1935 20.3039
R6407 VDD.n2913 VDD.n1935 20.3039
R6408 VDD.n2913 VDD.n1929 20.3039
R6409 VDD.n2919 VDD.n1929 20.3039
R6410 VDD.n2923 VDD.n1927 20.3039
R6411 VDD.n2931 VDD.n2930 20.3039
R6412 VDD.n2934 VDD.n1917 20.3039
R6413 VDD.n2941 VDD.n1917 20.3039
R6414 VDD.n2941 VDD.n1914 20.3039
R6415 VDD.n2945 VDD.n1914 20.3039
R6416 VDD.n2945 VDD.n1915 20.3039
R6417 VDD.n3001 VDD.n3000 20.3039
R6418 VDD.n3004 VDD.n1874 20.3039
R6419 VDD.n3011 VDD.n1874 20.3039
R6420 VDD.n3011 VDD.n1871 20.3039
R6421 VDD.n3015 VDD.n1871 20.3039
R6422 VDD.n3015 VDD.n1872 20.3039
R6423 VDD.n3072 VDD.n3071 20.3039
R6424 VDD.n3075 VDD.n1832 20.3039
R6425 VDD.n3082 VDD.n1832 20.3039
R6426 VDD.n3082 VDD.n1829 20.3039
R6427 VDD.n3086 VDD.n1829 20.3039
R6428 VDD.n3086 VDD.n1830 20.3039
R6429 VDD.n1806 VDD.n1002 20.3039
R6430 VDD.n1812 VDD.n1002 20.3039
R6431 VDD.n1793 VDD.n1007 20.3039
R6432 VDD.n1800 VDD.n1007 20.3039
R6433 VDD.n1783 VDD.n1018 20.3039
R6434 VDD.n1783 VDD.n1014 20.3039
R6435 VDD.n1789 VDD.n1014 20.3039
R6436 VDD.n1790 VDD.n1789 20.3039
R6437 VDD.n1730 VDD.n1042 20.3039
R6438 VDD.n1735 VDD.n1042 20.3039
R6439 VDD.n1718 VDD.n1051 20.3039
R6440 VDD.n1722 VDD.n1051 20.3039
R6441 VDD.n1708 VDD.n1060 20.3039
R6442 VDD.n1708 VDD.n1057 20.3039
R6443 VDD.n1712 VDD.n1057 20.3039
R6444 VDD.n1712 VDD.n1058 20.3039
R6445 VDD.n1652 VDD.n1085 20.3039
R6446 VDD.n1656 VDD.n1085 20.3039
R6447 VDD.n1641 VDD.n1093 20.3039
R6448 VDD.n1645 VDD.n1093 20.3039
R6449 VDD.n1631 VDD.n1102 20.3039
R6450 VDD.n1631 VDD.n1099 20.3039
R6451 VDD.n1635 VDD.n1099 20.3039
R6452 VDD.n1635 VDD.n1100 20.3039
R6453 VDD.n1575 VDD.n1127 20.3039
R6454 VDD.n1579 VDD.n1127 20.3039
R6455 VDD.n1564 VDD.n1135 20.3039
R6456 VDD.n1568 VDD.n1135 20.3039
R6457 VDD.n1554 VDD.n1144 20.3039
R6458 VDD.n1554 VDD.n1141 20.3039
R6459 VDD.n1558 VDD.n1141 20.3039
R6460 VDD.n1558 VDD.n1142 20.3039
R6461 VDD.n1498 VDD.n1169 20.3039
R6462 VDD.n1502 VDD.n1169 20.3039
R6463 VDD.n1487 VDD.n1177 20.3039
R6464 VDD.n1491 VDD.n1177 20.3039
R6465 VDD.n1477 VDD.n1186 20.3039
R6466 VDD.n1477 VDD.n1183 20.3039
R6467 VDD.n1481 VDD.n1183 20.3039
R6468 VDD.n1481 VDD.n1184 20.3039
R6469 VDD.n1421 VDD.n1211 20.3039
R6470 VDD.n1425 VDD.n1211 20.3039
R6471 VDD.n1410 VDD.n1219 20.3039
R6472 VDD.n1414 VDD.n1219 20.3039
R6473 VDD.n1400 VDD.n1228 20.3039
R6474 VDD.n1400 VDD.n1225 20.3039
R6475 VDD.n1404 VDD.n1225 20.3039
R6476 VDD.n1404 VDD.n1226 20.3039
R6477 VDD.n1344 VDD.n1253 20.3039
R6478 VDD.n1348 VDD.n1253 20.3039
R6479 VDD.n1333 VDD.n1261 20.3039
R6480 VDD.n1337 VDD.n1261 20.3039
R6481 VDD.n1323 VDD.n1270 20.3039
R6482 VDD.n1323 VDD.n1267 20.3039
R6483 VDD.n1327 VDD.n1267 20.3039
R6484 VDD.n1327 VDD.n1268 20.3039
R6485 VDD.n1289 VDD.n1281 20.3039
R6486 VDD.n1302 VDD.n1281 20.3039
R6487 VDD.n1315 VDD.n1275 20.3039
R6488 VDD.n1361 VDD.n1247 20.3039
R6489 VDD.n1366 VDD.n1239 20.3039
R6490 VDD.n1379 VDD.n1239 20.3039
R6491 VDD.n1392 VDD.n1233 20.3039
R6492 VDD.n1438 VDD.n1205 20.3039
R6493 VDD.n1443 VDD.n1197 20.3039
R6494 VDD.n1456 VDD.n1197 20.3039
R6495 VDD.n1469 VDD.n1191 20.3039
R6496 VDD.n1515 VDD.n1163 20.3039
R6497 VDD.n1520 VDD.n1155 20.3039
R6498 VDD.n1533 VDD.n1155 20.3039
R6499 VDD.n1546 VDD.n1149 20.3039
R6500 VDD.n1592 VDD.n1121 20.3039
R6501 VDD.n1597 VDD.n1113 20.3039
R6502 VDD.n1610 VDD.n1113 20.3039
R6503 VDD.n1623 VDD.n1107 20.3039
R6504 VDD.n1669 VDD.n1079 20.3039
R6505 VDD.n1674 VDD.n1071 20.3039
R6506 VDD.n1687 VDD.n1071 20.3039
R6507 VDD.n1700 VDD.n1065 20.3039
R6508 VDD.n1747 VDD.n1033 20.3039
R6509 VDD.n1755 VDD.n1030 20.3039
R6510 VDD.n1755 VDD.n1028 20.3039
R6511 VDD.n1776 VDD.n1022 20.3039
R6512 VDD.n161 VDD.n16 20.3039
R6513 VDD.n850 VDD.n2 20.3039
R6514 VDD.n707 VDD.n5 20.3039
R6515 VDD.n572 VDD.n8 20.3039
R6516 VDD.n439 VDD.n11 20.3039
R6517 VDD.n291 VDD.n13 20.3039
R6518 VDD.n3232 VDD.n3192 19.8626
R6519 VDD.n3322 VDD.n3132 19.8626
R6520 VDD.n2903 VDD.n1943 19.8626
R6521 VDD.n2953 VDD.n1908 19.8626
R6522 VDD.n3024 VDD.n1866 19.8626
R6523 VDD.n3091 VDD.n1826 19.8626
R6524 VDD.n3282 VDD.n3161 19.2005
R6525 VDD.n3372 VDD.n3101 19.2005
R6526 VDD.n3270 VDD.n3173 18.9798
R6527 VDD.n3360 VDD.n3113 18.9798
R6528 VDD.n1285 VDD.n1283 18.9798
R6529 VDD.n1247 VDD.n1243 18.9798
R6530 VDD.n1205 VDD.n1201 18.9798
R6531 VDD.n1163 VDD.n1159 18.9798
R6532 VDD.n1121 VDD.n1117 18.9798
R6533 VDD.n1079 VDD.n1075 18.9798
R6534 VDD.n1747 VDD.n1035 18.9798
R6535 VDD.n2716 VDD.n2715 18.7186
R6536 VDD.n2852 VDD.n2851 18.7186
R6537 VDD.n1806 VDD.n1005 18.3177
R6538 VDD.n1730 VDD.n1046 18.3177
R6539 VDD.n1652 VDD.n1089 18.3177
R6540 VDD.n1575 VDD.n1131 18.3177
R6541 VDD.n1498 VDD.n1173 18.3177
R6542 VDD.n1421 VDD.n1215 18.3177
R6543 VDD.n1344 VDD.n1257 18.3177
R6544 VDD.n2689 VDD.t301 18.2697
R6545 VDD.n2825 VDD.t321 18.2697
R6546 VDD.n2629 VDD.n2628 18.1151
R6547 VDD.n2765 VDD.n2764 18.1151
R6548 VDD.n3270 VDD.n3172 18.097
R6549 VDD.n3360 VDD.n3112 18.097
R6550 VDD.n3213 VDD.n3212 17.2143
R6551 VDD.n3232 VDD.n3197 17.2143
R6552 VDD.n3303 VDD.n3152 17.2143
R6553 VDD.n3322 VDD.n3137 17.2143
R6554 VDD.n3283 VDD.n3164 16.9936
R6555 VDD.n3373 VDD.n3104 16.9936
R6556 VDD.n1302 VDD.n1282 16.7993
R6557 VDD.n1379 VDD.n1240 16.7993
R6558 VDD.n1456 VDD.n1198 16.7993
R6559 VDD.n1533 VDD.n1156 16.7993
R6560 VDD.n1610 VDD.n1114 16.7993
R6561 VDD.n1687 VDD.n1072 16.7993
R6562 VDD.n1759 VDD.n1028 16.7993
R6563 VDD.n3294 VDD 16.7729
R6564 VDD.n3384 VDD 16.7729
R6565 VDD.n3243 VDD.n3188 16.3315
R6566 VDD.n3333 VDD.n3128 16.3315
R6567 VDD.n1331 VDD.t54 15.8338
R6568 VDD.n1408 VDD.t736 15.8338
R6569 VDD.n1485 VDD.t573 15.8338
R6570 VDD.n1562 VDD.t673 15.8338
R6571 VDD.n1639 VDD.t721 15.8338
R6572 VDD.n1716 VDD.t327 15.8338
R6573 VDD.t667 VDD.n1795 15.8338
R6574 VDD.n73 VDD.t315 15.79
R6575 VDD.n213 VDD.t360 15.79
R6576 VDD.n348 VDD.t107 15.79
R6577 VDD.n491 VDD.t435 15.79
R6578 VDD.n624 VDD.t634 15.79
R6579 VDD.n759 VDD.t19 15.79
R6580 VDD.n902 VDD.t317 15.79
R6581 VDD.n2364 VDD.n2216 15.6598
R6582 VDD.n2366 VDD.n2206 15.6598
R6583 VDD.n2378 VDD.n2376 15.6598
R6584 VDD.n2389 VDD.n2388 15.6598
R6585 VDD.n2400 VDD.n2194 15.6598
R6586 VDD.n2402 VDD.n2186 15.6598
R6587 VDD.n2414 VDD.n2412 15.6598
R6588 VDD.n2425 VDD.n2424 15.6598
R6589 VDD.n2439 VDD 15.6598
R6590 VDD.n2544 VDD.n2543 15.6598
R6591 VDD.n2555 VDD.n2554 15.6598
R6592 VDD.n2568 VDD.n2108 15.6598
R6593 VDD.n2571 VDD.n2570 15.6598
R6594 VDD.n2582 VDD.n2581 15.6598
R6595 VDD.n2593 VDD.n2592 15.6598
R6596 VDD.n2604 VDD.n2088 15.6598
R6597 VDD.n2608 VDD.n2607 15.6598
R6598 VDD.n2620 VDD 15.6598
R6599 VDD.n2917 VDD.t555 15.6598
R6600 VDD.t590 VDD.n2936 15.6598
R6601 VDD.n2961 VDD.t100 15.6598
R6602 VDD.t159 VDD.n3006 15.6598
R6603 VDD.n3032 VDD.t429 15.6598
R6604 VDD.t177 VDD.n3077 15.6598
R6605 VDD.n1316 VDD.n1315 15.4488
R6606 VDD.n1393 VDD.n1392 15.4488
R6607 VDD.n1470 VDD.n1469 15.4488
R6608 VDD.n1547 VDD.n1546 15.4488
R6609 VDD.n1624 VDD.n1623 15.4488
R6610 VDD.n1701 VDD.n1700 15.4488
R6611 VDD.n1777 VDD.n1776 15.4488
R6612 VDD.n2443 VDD.n2171 15.0975
R6613 VDD.n3265 VDD.n3176 14.566
R6614 VDD.n3355 VDD.n3116 14.566
R6615 VDD.n2445 VDD.n2444 13.8904
R6616 VDD.n954 VDD.n950 13.7148
R6617 VDD.n3218 VDD.n3210 13.6833
R6618 VDD.n3201 VDD.n3195 13.6833
R6619 VDD.n3308 VDD.n3150 13.6833
R6620 VDD.n3141 VDD.n3135 13.6833
R6621 VDD.n198 VDD 13.6005
R6622 VDD.n58 VDD 13.6005
R6623 VDD.n333 VDD 13.6005
R6624 VDD.n476 VDD 13.6005
R6625 VDD.n609 VDD 13.6005
R6626 VDD.n744 VDD 13.6005
R6627 VDD.n887 VDD 13.6005
R6628 VDD.n1817 VDD.n996 13.4626
R6629 VDD.n1742 VDD.n1038 13.4626
R6630 VDD.n1663 VDD.n1078 13.4626
R6631 VDD.n1586 VDD.n1120 13.4626
R6632 VDD.n1509 VDD.n1162 13.4626
R6633 VDD.n1432 VDD.n1204 13.4626
R6634 VDD.n1355 VDD.n1246 13.4626
R6635 VDD.n3294 VDD.n3156 13.0212
R6636 VDD.n3300 VDD.n3156 13.0212
R6637 VDD.n3384 VDD.n3096 13.0212
R6638 VDD.n3390 VDD.n3096 13.0212
R6639 VDD.n3189 VDD.n3184 12.8005
R6640 VDD.n3129 VDD.n3124 12.8005
R6641 VDD.n2273 VDD.n2272 12.8005
R6642 VDD.n2284 VDD.n2283 12.8005
R6643 VDD.n2290 VDD.n2289 12.8005
R6644 VDD.n2302 VDD.n2301 12.8005
R6645 VDD.n2311 VDD.n2310 12.8005
R6646 VDD.n2329 VDD.n2328 12.8005
R6647 VDD.n2369 VDD.n2368 12.8005
R6648 VDD.n2386 VDD.n2385 12.8005
R6649 VDD.n2394 VDD.n2196 12.8005
R6650 VDD.n2405 VDD.n2404 12.8005
R6651 VDD.n2189 VDD.n2184 12.8005
R6652 VDD.n2422 VDD.n2421 12.8005
R6653 VDD.n2431 VDD.n2174 12.8005
R6654 VDD.n2456 VDD.n2455 12.8005
R6655 VDD.n2462 VDD.n2461 12.8005
R6656 VDD.n2474 VDD.n2473 12.8005
R6657 VDD.n2482 VDD.n2481 12.8005
R6658 VDD.n2493 VDD.n2492 12.8005
R6659 VDD.n2499 VDD.n2498 12.8005
R6660 VDD.n2520 VDD.n2519 12.8005
R6661 VDD.n2552 VDD.n2551 12.8005
R6662 VDD.n2574 VDD.n2573 12.8005
R6663 VDD.n2103 VDD.n2099 12.8005
R6664 VDD.n2590 VDD.n2589 12.8005
R6665 VDD.n2598 VDD.n2090 12.8005
R6666 VDD.n2611 VDD.n2610 12.8005
R6667 VDD.n2618 VDD.n2617 12.8005
R6668 VDD.n2640 VDD.n2639 12.8005
R6669 VDD.n2647 VDD.n2646 12.8005
R6670 VDD.n2659 VDD.n2658 12.8005
R6671 VDD.n2667 VDD.n2666 12.8005
R6672 VDD.n2678 VDD.n2677 12.8005
R6673 VDD.n2684 VDD.n2683 12.8005
R6674 VDD.n2705 VDD.n2704 12.8005
R6675 VDD.n2776 VDD.n2775 12.8005
R6676 VDD.n2783 VDD.n2782 12.8005
R6677 VDD.n2795 VDD.n2794 12.8005
R6678 VDD.n2803 VDD.n2802 12.8005
R6679 VDD.n2814 VDD.n2813 12.8005
R6680 VDD.n2820 VDD.n2819 12.8005
R6681 VDD.n2841 VDD.n2840 12.8005
R6682 VDD.n2264 VDD.n2263 12.5798
R6683 VDD.n1812 VDD.n1000 12.5798
R6684 VDD.n1736 VDD.n1735 12.5798
R6685 VDD.n1656 VDD.n1082 12.5798
R6686 VDD.n1579 VDD.n1124 12.5798
R6687 VDD.n1502 VDD.n1166 12.5798
R6688 VDD.n1425 VDD.n1208 12.5798
R6689 VDD.n1348 VDD.n1250 12.5798
R6690 VDD.n1361 VDD.n1246 12.5798
R6691 VDD.n1438 VDD.n1204 12.5798
R6692 VDD.n1515 VDD.n1162 12.5798
R6693 VDD.n1592 VDD.n1120 12.5798
R6694 VDD.n1669 VDD.n1078 12.5798
R6695 VDD.n1742 VDD.n1033 12.5798
R6696 VDD.n1822 VDD.n996 12.5798
R6697 VDD.n162 VDD.n161 12.5798
R6698 VDD.n22 VDD.n18 12.5798
R6699 VDD.n851 VDD.n850 12.5798
R6700 VDD.n708 VDD.n707 12.5798
R6701 VDD.n573 VDD.n572 12.5798
R6702 VDD.n440 VDD.n439 12.5798
R6703 VDD.n297 VDD.n13 12.5798
R6704 VDD.n1817 VDD.n1000 12.3591
R6705 VDD.n1736 VDD.n1038 12.3591
R6706 VDD.n1663 VDD.n1082 12.3591
R6707 VDD.n1586 VDD.n1124 12.3591
R6708 VDD.n1509 VDD.n1166 12.3591
R6709 VDD.n1432 VDD.n1208 12.3591
R6710 VDD.n1355 VDD.n1250 12.3591
R6711 VDD.n2984 VDD.n2983 12.242
R6712 VDD.n3055 VDD.n3054 12.242
R6713 VDD.n2959 VDD.n1903 11.9177
R6714 VDD.n2957 VDD.n1905 11.9177
R6715 VDD.n2965 VDD.n1900 11.9177
R6716 VDD.n2967 VDD.n2966 11.9177
R6717 VDD.n2972 VDD.n1896 11.9177
R6718 VDD.n2971 VDD.n1898 11.9177
R6719 VDD.n2980 VDD.n1888 11.9177
R6720 VDD.n3030 VDD.n1861 11.9177
R6721 VDD.n3028 VDD.n1863 11.9177
R6722 VDD.n3036 VDD.n1858 11.9177
R6723 VDD.n3038 VDD.n3037 11.9177
R6724 VDD.n3043 VDD.n1854 11.9177
R6725 VDD.n3042 VDD.n1856 11.9177
R6726 VDD.n3051 VDD.n1846 11.9177
R6727 VDD.n2725 VDD.n2023 11.7196
R6728 VDD.n2861 VDD.n1956 11.7196
R6729 VDD.n2737 VDD.n2733 11.4764
R6730 VDD.n2742 VDD.n2741 11.4764
R6731 VDD.n2021 VDD.n2017 11.4764
R6732 VDD.n2751 VDD.n2749 11.4764
R6733 VDD.n2750 VDD.n2012 11.4764
R6734 VDD.n2757 VDD.n2756 11.4764
R6735 VDD.n2014 VDD.n2009 11.4764
R6736 VDD.n2873 VDD.n2869 11.4764
R6737 VDD.n2878 VDD.n2877 11.4764
R6738 VDD.n1954 VDD.n1950 11.4764
R6739 VDD.n2886 VDD.n2885 11.4764
R6740 VDD.n2889 VDD.n1948 11.4764
R6741 VDD.n2893 VDD.n2892 11.4764
R6742 VDD.n2900 VDD.n1945 11.4764
R6743 VDD.n3258 VDD.n3180 11.035
R6744 VDD.n3348 VDD.n3120 11.035
R6745 VDD.t230 VDD.n3224 10.5561
R6746 VDD.n3225 VDD.t242 10.5561
R6747 VDD.t412 VDD.n3314 10.5561
R6748 VDD.n3315 VDD.t398 10.5561
R6749 VDD.n1319 VDD.t165 10.5561
R6750 VDD.n1396 VDD.t257 10.5561
R6751 VDD.n1473 VDD.t303 10.5561
R6752 VDD.n1550 VDD.t621 10.5561
R6753 VDD.n1627 VDD.t642 10.5561
R6754 VDD.n1704 VDD.t569 10.5561
R6755 VDD.t644 VDD.n1016 10.5561
R6756 VDD.n93 VDD.t119 10.5268
R6757 VDD.n233 VDD.t586 10.5268
R6758 VDD.n368 VDD.t294 10.5268
R6759 VDD.n511 VDD.t734 10.5268
R6760 VDD.n644 VDD.t80 10.5268
R6761 VDD.n779 VDD.t713 10.5268
R6762 VDD.n922 VDD.t181 10.5268
R6763 VDD.n953 VDD.n952 10.5268
R6764 VDD.n2688 VDD.t272 10.4401
R6765 VDD.t286 VDD.n2760 10.4401
R6766 VDD.n2824 VDD.t351 10.4401
R6767 VDD.t448 VDD.n2896 10.4401
R6768 VDD.n3222 VDD.n3206 10.1522
R6769 VDD.n3206 VDD.n3199 10.1522
R6770 VDD.n3312 VDD.n3146 10.1522
R6771 VDD.n3146 VDD.n3139 10.1522
R6772 VDD.n2735 VDD.n2020 10.1522
R6773 VDD.n2871 VDD.n1953 10.1522
R6774 VDD.n2919 VDD.n1931 10.1522
R6775 VDD.n1931 VDD.n1927 10.1522
R6776 VDD.n2931 VDD.n1921 10.1522
R6777 VDD.n2934 VDD.n1921 10.1522
R6778 VDD.n1897 VDD.n1891 10.1522
R6779 VDD.n3001 VDD.n1878 10.1522
R6780 VDD.n3004 VDD.n1878 10.1522
R6781 VDD.n1855 VDD.n1849 10.1522
R6782 VDD.n3072 VDD.n1836 10.1522
R6783 VDD.n3075 VDD.n1836 10.1522
R6784 VDD.n2323 VDD.n2322 9.93153
R6785 VDD.n1278 VDD.n1275 9.84589
R6786 VDD.n1236 VDD.n1233 9.84589
R6787 VDD.n1194 VDD.n1191 9.84589
R6788 VDD.n1152 VDD.n1149 9.84589
R6789 VDD.n1110 VDD.n1107 9.84589
R6790 VDD.n1068 VDD.n1065 9.84589
R6791 VDD.n1025 VDD.n1022 9.84589
R6792 VDD.n2511 VDD.n2510 9.71084
R6793 VDD.n2274 VDD.n2273 9.3005
R6794 VDD.n2277 VDD.n2276 9.3005
R6795 VDD.n2278 VDD.n2277 9.3005
R6796 VDD.n2279 VDD.n2278 9.3005
R6797 VDD.n2284 VDD.n2246 9.3005
R6798 VDD.n2287 VDD.n2245 9.3005
R6799 VDD.n2245 VDD.n2244 9.3005
R6800 VDD.n2244 VDD.n2243 9.3005
R6801 VDD.n2289 VDD.n2288 9.3005
R6802 VDD.n2298 VDD.n2297 9.3005
R6803 VDD.n2297 VDD.n2296 9.3005
R6804 VDD.n2296 VDD.n2295 9.3005
R6805 VDD.n2301 VDD.n2300 9.3005
R6806 VDD.n2234 VDD.n2233 9.3005
R6807 VDD.n2235 VDD.n2234 9.3005
R6808 VDD.n2305 VDD.n2235 9.3005
R6809 VDD.n2312 VDD.n2311 9.3005
R6810 VDD.n2315 VDD.n2314 9.3005
R6811 VDD.n2316 VDD.n2315 9.3005
R6812 VDD.n2317 VDD.n2316 9.3005
R6813 VDD.n2323 VDD.n2227 9.3005
R6814 VDD.n2326 VDD.n2226 9.3005
R6815 VDD.n2226 VDD.n2225 9.3005
R6816 VDD.n2225 VDD.n2224 9.3005
R6817 VDD.n2328 VDD.n2327 9.3005
R6818 VDD.n2359 VDD.n2358 9.3005
R6819 VDD.n2358 VDD.n2357 9.3005
R6820 VDD.n2357 VDD.n2356 9.3005
R6821 VDD.n2361 VDD.n2360 9.3005
R6822 VDD.n2361 VDD.n2215 9.3005
R6823 VDD.n2365 VDD.n2215 9.3005
R6824 VDD.n2370 VDD.n2369 9.3005
R6825 VDD.n2373 VDD.n2372 9.3005
R6826 VDD.n2374 VDD.n2373 9.3005
R6827 VDD.n2375 VDD.n2374 9.3005
R6828 VDD.n2211 VDD.n2203 9.3005
R6829 VDD.n2382 VDD.n2381 9.3005
R6830 VDD.n2381 VDD.n2201 9.3005
R6831 VDD.n2377 VDD.n2201 9.3005
R6832 VDD.n2385 VDD.n2384 9.3005
R6833 VDD.n2392 VDD.n2199 9.3005
R6834 VDD.n2392 VDD.n2391 9.3005
R6835 VDD.n2391 VDD.n2390 9.3005
R6836 VDD.n2395 VDD.n2394 9.3005
R6837 VDD.n2397 VDD.n2396 9.3005
R6838 VDD.n2397 VDD.n2193 9.3005
R6839 VDD.n2401 VDD.n2193 9.3005
R6840 VDD.n2406 VDD.n2405 9.3005
R6841 VDD.n2409 VDD.n2408 9.3005
R6842 VDD.n2410 VDD.n2409 9.3005
R6843 VDD.n2411 VDD.n2410 9.3005
R6844 VDD.n2189 VDD.n2183 9.3005
R6845 VDD.n2418 VDD.n2417 9.3005
R6846 VDD.n2417 VDD.n2181 9.3005
R6847 VDD.n2413 VDD.n2181 9.3005
R6848 VDD.n2421 VDD.n2420 9.3005
R6849 VDD.n2428 VDD.n2179 9.3005
R6850 VDD.n2428 VDD.n2427 9.3005
R6851 VDD.n2427 VDD.n2426 9.3005
R6852 VDD.n2432 VDD.n2431 9.3005
R6853 VDD.n2436 VDD.n2435 9.3005
R6854 VDD.n2436 VDD.n2172 9.3005
R6855 VDD.n2440 VDD.n2172 9.3005
R6856 VDD.n2433 VDD.n2171 9.3005
R6857 VDD.n2446 VDD.n2445 9.3005
R6858 VDD.n2449 VDD.n2448 9.3005
R6859 VDD.n2450 VDD.n2449 9.3005
R6860 VDD.n2451 VDD.n2450 9.3005
R6861 VDD.n2456 VDD.n2164 9.3005
R6862 VDD.n2459 VDD.n2163 9.3005
R6863 VDD.n2163 VDD.n2162 9.3005
R6864 VDD.n2162 VDD.n2161 9.3005
R6865 VDD.n2461 VDD.n2460 9.3005
R6866 VDD.n2470 VDD.n2469 9.3005
R6867 VDD.n2469 VDD.n2468 9.3005
R6868 VDD.n2468 VDD.n2467 9.3005
R6869 VDD.n2473 VDD.n2472 9.3005
R6870 VDD.n2152 VDD.n2151 9.3005
R6871 VDD.n2153 VDD.n2152 9.3005
R6872 VDD.n2477 VDD.n2153 9.3005
R6873 VDD.n2483 VDD.n2482 9.3005
R6874 VDD.n2486 VDD.n2485 9.3005
R6875 VDD.n2487 VDD.n2486 9.3005
R6876 VDD.n2488 VDD.n2487 9.3005
R6877 VDD.n2493 VDD.n2145 9.3005
R6878 VDD.n2496 VDD.n2144 9.3005
R6879 VDD.n2144 VDD.n2143 9.3005
R6880 VDD.n2143 VDD.n2142 9.3005
R6881 VDD.n2498 VDD.n2497 9.3005
R6882 VDD.n2507 VDD.n2506 9.3005
R6883 VDD.n2506 VDD.n2505 9.3005
R6884 VDD.n2505 VDD.n2504 9.3005
R6885 VDD.n2510 VDD.n2509 9.3005
R6886 VDD.n2132 VDD.n2131 9.3005
R6887 VDD.n2133 VDD.n2132 9.3005
R6888 VDD.n2515 VDD.n2133 9.3005
R6889 VDD.n2521 VDD.n2520 9.3005
R6890 VDD.n2524 VDD.n2523 9.3005
R6891 VDD.n2525 VDD.n2524 9.3005
R6892 VDD.n2526 VDD.n2525 9.3005
R6893 VDD.n2548 VDD.n2547 9.3005
R6894 VDD.n2547 VDD.n2116 9.3005
R6895 VDD.n2116 VDD.n2115 9.3005
R6896 VDD.n2551 VDD.n2550 9.3005
R6897 VDD.n2558 VDD.n2113 9.3005
R6898 VDD.n2558 VDD.n2557 9.3005
R6899 VDD.n2557 VDD.n2556 9.3005
R6900 VDD.n2563 VDD.n2562 9.3005
R6901 VDD.n2565 VDD.n2564 9.3005
R6902 VDD.n2565 VDD.n2107 9.3005
R6903 VDD.n2569 VDD.n2107 9.3005
R6904 VDD.n2575 VDD.n2574 9.3005
R6905 VDD.n2578 VDD.n2577 9.3005
R6906 VDD.n2579 VDD.n2578 9.3005
R6907 VDD.n2580 VDD.n2579 9.3005
R6908 VDD.n2103 VDD.n2098 9.3005
R6909 VDD.n2586 VDD.n2585 9.3005
R6910 VDD.n2585 VDD.n2096 9.3005
R6911 VDD.n2096 VDD.n2095 9.3005
R6912 VDD.n2589 VDD.n2588 9.3005
R6913 VDD.n2596 VDD.n2093 9.3005
R6914 VDD.n2596 VDD.n2595 9.3005
R6915 VDD.n2595 VDD.n2594 9.3005
R6916 VDD.n2599 VDD.n2598 9.3005
R6917 VDD.n2601 VDD.n2600 9.3005
R6918 VDD.n2601 VDD.n2086 9.3005
R6919 VDD.n2605 VDD.n2086 9.3005
R6920 VDD.n2612 VDD.n2611 9.3005
R6921 VDD.n2613 VDD.n2082 9.3005
R6922 VDD.n2082 VDD.n2080 9.3005
R6923 VDD.n2606 VDD.n2080 9.3005
R6924 VDD.n2617 VDD.n2077 9.3005
R6925 VDD.n2624 VDD.n2623 9.3005
R6926 VDD.n2623 VDD.n2622 9.3005
R6927 VDD.n2622 VDD.n2621 9.3005
R6928 VDD.n2627 VDD.n2626 9.3005
R6929 VDD.n2630 VDD.n2629 9.3005
R6930 VDD.n2633 VDD.n2632 9.3005
R6931 VDD.n2634 VDD.n2633 9.3005
R6932 VDD.n2635 VDD.n2634 9.3005
R6933 VDD.n2640 VDD.n2069 9.3005
R6934 VDD.n2644 VDD.n2068 9.3005
R6935 VDD.n2068 VDD.n2067 9.3005
R6936 VDD.n2067 VDD.n2066 9.3005
R6937 VDD.n2646 VDD.n2645 9.3005
R6938 VDD.n2655 VDD.n2654 9.3005
R6939 VDD.n2654 VDD.n2653 9.3005
R6940 VDD.n2653 VDD.n2652 9.3005
R6941 VDD.n2658 VDD.n2657 9.3005
R6942 VDD.n2057 VDD.n2056 9.3005
R6943 VDD.n2058 VDD.n2057 9.3005
R6944 VDD.n2662 VDD.n2058 9.3005
R6945 VDD.n2668 VDD.n2667 9.3005
R6946 VDD.n2671 VDD.n2670 9.3005
R6947 VDD.n2672 VDD.n2671 9.3005
R6948 VDD.n2673 VDD.n2672 9.3005
R6949 VDD.n2678 VDD.n2050 9.3005
R6950 VDD.n2681 VDD.n2049 9.3005
R6951 VDD.n2049 VDD.n2048 9.3005
R6952 VDD.n2048 VDD.n2047 9.3005
R6953 VDD.n2683 VDD.n2682 9.3005
R6954 VDD.n2692 VDD.n2691 9.3005
R6955 VDD.n2691 VDD.n2690 9.3005
R6956 VDD.n2690 VDD.n2689 9.3005
R6957 VDD.n2695 VDD.n2694 9.3005
R6958 VDD.n2037 VDD.n2036 9.3005
R6959 VDD.n2038 VDD.n2037 9.3005
R6960 VDD.n2700 VDD.n2038 9.3005
R6961 VDD.n2706 VDD.n2705 9.3005
R6962 VDD.n2709 VDD.n2708 9.3005
R6963 VDD.n2710 VDD.n2709 9.3005
R6964 VDD.n2711 VDD.n2710 9.3005
R6965 VDD.n2769 VDD.n2768 9.3005
R6966 VDD.n2770 VDD.n2769 9.3005
R6967 VDD.n2771 VDD.n2770 9.3005
R6968 VDD.n2776 VDD.n2002 9.3005
R6969 VDD.n2780 VDD.n2001 9.3005
R6970 VDD.n2001 VDD.n2000 9.3005
R6971 VDD.n2000 VDD.n1999 9.3005
R6972 VDD.n2782 VDD.n2781 9.3005
R6973 VDD.n2791 VDD.n2790 9.3005
R6974 VDD.n2790 VDD.n2789 9.3005
R6975 VDD.n2789 VDD.n2788 9.3005
R6976 VDD.n2794 VDD.n2793 9.3005
R6977 VDD.n1990 VDD.n1989 9.3005
R6978 VDD.n1991 VDD.n1990 9.3005
R6979 VDD.n2798 VDD.n1991 9.3005
R6980 VDD.n2804 VDD.n2803 9.3005
R6981 VDD.n2807 VDD.n2806 9.3005
R6982 VDD.n2808 VDD.n2807 9.3005
R6983 VDD.n2809 VDD.n2808 9.3005
R6984 VDD.n2814 VDD.n1983 9.3005
R6985 VDD.n2817 VDD.n1982 9.3005
R6986 VDD.n1982 VDD.n1981 9.3005
R6987 VDD.n1981 VDD.n1980 9.3005
R6988 VDD.n2819 VDD.n2818 9.3005
R6989 VDD.n2828 VDD.n2827 9.3005
R6990 VDD.n2827 VDD.n2826 9.3005
R6991 VDD.n2826 VDD.n2825 9.3005
R6992 VDD.n2831 VDD.n2830 9.3005
R6993 VDD.n1970 VDD.n1969 9.3005
R6994 VDD.n1971 VDD.n1970 9.3005
R6995 VDD.n2836 VDD.n1971 9.3005
R6996 VDD.n2842 VDD.n2841 9.3005
R6997 VDD.n2845 VDD.n2844 9.3005
R6998 VDD.n2846 VDD.n2845 9.3005
R6999 VDD.n2847 VDD.n2846 9.3005
R7000 VDD.n2766 VDD.n2765 9.3005
R7001 VDD.n2262 VDD.n2261 9.3005
R7002 VDD.n2252 VDD.n2251 9.3005
R7003 VDD.n2253 VDD.n2252 9.3005
R7004 VDD.n2267 VDD.n2253 9.3005
R7005 VDD.n1766 VDD.n1024 9.3005
R7006 VDD.n1763 VDD.n1026 9.3005
R7007 VDD.n1067 VDD.n1066 9.3005
R7008 VDD.n1684 VDD.n1683 9.3005
R7009 VDD.n1109 VDD.n1108 9.3005
R7010 VDD.n1607 VDD.n1606 9.3005
R7011 VDD.n1151 VDD.n1150 9.3005
R7012 VDD.n1530 VDD.n1529 9.3005
R7013 VDD.n1193 VDD.n1192 9.3005
R7014 VDD.n1453 VDD.n1452 9.3005
R7015 VDD.n1235 VDD.n1234 9.3005
R7016 VDD.n1376 VDD.n1375 9.3005
R7017 VDD.n1277 VDD.n1276 9.3005
R7018 VDD.n1299 VDD.n1298 9.3005
R7019 VDD.n196 VDD.n195 9.3005
R7020 VDD.n195 VDD.n193 9.3005
R7021 VDD.n56 VDD.n55 9.3005
R7022 VDD.n55 VDD.n53 9.3005
R7023 VDD.n331 VDD.n330 9.3005
R7024 VDD.n330 VDD.n328 9.3005
R7025 VDD.n474 VDD.n473 9.3005
R7026 VDD.n473 VDD.n471 9.3005
R7027 VDD.n607 VDD.n606 9.3005
R7028 VDD.n606 VDD.n604 9.3005
R7029 VDD.n742 VDD.n741 9.3005
R7030 VDD.n741 VDD.n739 9.3005
R7031 VDD.n885 VDD.n884 9.3005
R7032 VDD.n884 VDD.n882 9.3005
R7033 VDD.n125 VDD.n124 9.3005
R7034 VDD.n124 VDD.n123 9.3005
R7035 VDD.n972 VDD.n971 9.3005
R7036 VDD.n971 VDD.n970 9.3005
R7037 VDD.n955 VDD.n954 9.3005
R7038 VDD.n954 VDD.n953 9.3005
R7039 VDD.n811 VDD.n810 9.3005
R7040 VDD.n810 VDD.n809 9.3005
R7041 VDD.n825 VDD.n824 9.3005
R7042 VDD.n824 VDD.n823 9.3005
R7043 VDD.n683 VDD.n682 9.3005
R7044 VDD.n682 VDD.n681 9.3005
R7045 VDD.n549 VDD.n548 9.3005
R7046 VDD.n548 VDD.n547 9.3005
R7047 VDD.n415 VDD.n414 9.3005
R7048 VDD.n414 VDD.n413 9.3005
R7049 VDD.n400 VDD.n399 9.3005
R7050 VDD.n399 VDD.n398 9.3005
R7051 VDD.n3254 VDD.n3180 9.26947
R7052 VDD.n3344 VDD.n3120 9.26947
R7053 VDD.n3283 VDD.n3282 9.04877
R7054 VDD.n3373 VDD.n3372 9.04877
R7055 VDD.n200 VDD.n199 8.94661
R7056 VDD.n60 VDD.n59 8.94661
R7057 VDD.n335 VDD.n334 8.94661
R7058 VDD.n478 VDD.n477 8.94661
R7059 VDD.n611 VDD.n610 8.94661
R7060 VDD.n746 VDD.n745 8.94661
R7061 VDD.n889 VDD.n888 8.94661
R7062 VDD.n2211 VDD.n2210 8.82809
R7063 VDD.n2562 VDD.n2561 8.82809
R7064 VDD.n2733 VDD.n2023 8.82809
R7065 VDD.n2737 VDD.n2736 8.82809
R7066 VDD.n2742 VDD.n2020 8.82809
R7067 VDD.n2741 VDD.n2021 8.82809
R7068 VDD.n2749 VDD.n2017 8.82809
R7069 VDD.n2751 VDD.n2750 8.82809
R7070 VDD.n2757 VDD.n2012 8.82809
R7071 VDD.n2763 VDD.n2009 8.82809
R7072 VDD.n2869 VDD.n1956 8.82809
R7073 VDD.n2873 VDD.n2872 8.82809
R7074 VDD.n2878 VDD.n1953 8.82809
R7075 VDD.n2877 VDD.n1954 8.82809
R7076 VDD.n2885 VDD.n1950 8.82809
R7077 VDD.n2886 VDD.n1948 8.82809
R7078 VDD.n2893 VDD.n2889 8.82809
R7079 VDD.n2900 VDD.n2899 8.82809
R7080 VDD.n1310 VDD.n1277 8.69304
R7081 VDD.n1387 VDD.n1235 8.69304
R7082 VDD.n1464 VDD.n1193 8.69304
R7083 VDD.n1541 VDD.n1151 8.69304
R7084 VDD.n1618 VDD.n1109 8.69304
R7085 VDD.n1695 VDD.n1067 8.69304
R7086 VDD.n1769 VDD.n1024 8.69304
R7087 VDD.n3157 VDD.n3156 8.47281
R7088 VDD.n3097 VDD.n3096 8.47281
R7089 VDD.n1246 VDD.n1245 8.47281
R7090 VDD.n1204 VDD.n1203 8.47281
R7091 VDD.n1162 VDD.n1161 8.47281
R7092 VDD.n1120 VDD.n1119 8.47281
R7093 VDD.n1078 VDD.n1077 8.47281
R7094 VDD.n1742 VDD.n1741 8.47281
R7095 VDD.n997 VDD.n996 8.47281
R7096 VDD.n3374 VDD.n3373 8.47276
R7097 VDD.n3284 VDD.n3283 8.47276
R7098 VDD.n162 VDD.n15 8.47276
R7099 VDD.n297 VDD.n296 8.47276
R7100 VDD.n22 VDD.n21 8.47181
R7101 VDD.n440 VDD.n10 8.47181
R7102 VDD.n573 VDD.n7 8.47181
R7103 VDD.n708 VDD.n4 8.47181
R7104 VDD.n851 VDD.n1 8.47181
R7105 VDD.n31 VDD.n30 8.47137
R7106 VDD.n171 VDD.n170 8.47137
R7107 VDD.n1251 VDD.n1250 8.47133
R7108 VDD.n1209 VDD.n1208 8.47133
R7109 VDD.n1167 VDD.n1166 8.47133
R7110 VDD.n1125 VDD.n1124 8.47133
R7111 VDD.n1083 VDD.n1082 8.47133
R7112 VDD.n1737 VDD.n1736 8.47133
R7113 VDD.n1000 VDD.n999 8.47133
R7114 VDD.n306 VDD.n305 8.47133
R7115 VDD.n860 VDD.n859 8.47037
R7116 VDD.n717 VDD.n716 8.47037
R7117 VDD.n582 VDD.n581 8.47037
R7118 VDD.n449 VDD.n448 8.47037
R7119 VDD.n240 VDD.n239 8.47011
R7120 VDD.n1258 VDD.n1257 8.47007
R7121 VDD.n1216 VDD.n1215 8.47007
R7122 VDD.n1174 VDD.n1173 8.47007
R7123 VDD.n1132 VDD.n1131 8.47007
R7124 VDD.n1090 VDD.n1089 8.47007
R7125 VDD.n1047 VDD.n1046 8.47007
R7126 VDD.n1005 VDD.n1004 8.47007
R7127 VDD.n1777 VDD.n1021 8.47007
R7128 VDD.n1702 VDD.n1701 8.47007
R7129 VDD.n1625 VDD.n1624 8.47007
R7130 VDD.n1548 VDD.n1547 8.47007
R7131 VDD.n1471 VDD.n1470 8.47007
R7132 VDD.n1394 VDD.n1393 8.47007
R7133 VDD.n1317 VDD.n1316 8.47007
R7134 VDD.n100 VDD.n99 8.47007
R7135 VDD.n929 VDD.n928 8.46911
R7136 VDD.n786 VDD.n785 8.46911
R7137 VDD.n651 VDD.n650 8.46911
R7138 VDD.n518 VDD.n517 8.46911
R7139 VDD.n375 VDD.n374 8.46911
R7140 VDD.n943 VDD.n942 8.46584
R7141 VDD.n3295 VDD.n3294 8.45089
R7142 VDD.n3296 VDD.n3295 8.45089
R7143 VDD.n3287 VDD.n3158 8.45089
R7144 VDD.n3289 VDD.n3288 8.45089
R7145 VDD.n3286 VDD.n3162 8.45089
R7146 VDD.n3285 VDD.n3284 8.45089
R7147 VDD.n3274 VDD.n3163 8.45089
R7148 VDD.n3276 VDD.n3275 8.45089
R7149 VDD.n3273 VDD.n3169 8.45089
R7150 VDD.n3272 VDD.n3271 8.45089
R7151 VDD.n3262 VDD.n3170 8.45089
R7152 VDD.n3264 VDD.n3263 8.45089
R7153 VDD.n3261 VDD.n3177 8.45089
R7154 VDD.n3260 VDD.n3259 8.45089
R7155 VDD.t224 VDD.n3178 8.45089
R7156 VDD.n3252 VDD.n3251 8.45089
R7157 VDD.n3250 VDD.n3185 8.45089
R7158 VDD.n3249 VDD.n3248 8.45089
R7159 VDD.n3239 VDD.n3186 8.45089
R7160 VDD.n3241 VDD.n3240 8.45089
R7161 VDD.n3238 VDD.n3193 8.45089
R7162 VDD.n3237 VDD.n3236 8.45089
R7163 VDD.n3226 VDD.n3194 8.45089
R7164 VDD.n3228 VDD.n3227 8.45089
R7165 VDD.n3225 VDD.n3202 8.45089
R7166 VDD.n3224 VDD.n3223 8.45089
R7167 VDD.n3215 VDD.n3203 8.45089
R7168 VDD.n3217 VDD.n3216 8.45089
R7169 VDD.n3297 VDD.n3157 8.45089
R7170 VDD.n3299 VDD.n3298 8.45089
R7171 VDD.n3385 VDD.n3384 8.45089
R7172 VDD.n3386 VDD.n3385 8.45089
R7173 VDD.n3377 VDD.n3098 8.45089
R7174 VDD.n3379 VDD.n3378 8.45089
R7175 VDD.n3376 VDD.n3102 8.45089
R7176 VDD.n3375 VDD.n3374 8.45089
R7177 VDD.n3364 VDD.n3103 8.45089
R7178 VDD.n3366 VDD.n3365 8.45089
R7179 VDD.n3363 VDD.n3109 8.45089
R7180 VDD.n3362 VDD.n3361 8.45089
R7181 VDD.n3352 VDD.n3110 8.45089
R7182 VDD.n3354 VDD.n3353 8.45089
R7183 VDD.n3351 VDD.n3117 8.45089
R7184 VDD.n3350 VDD.n3349 8.45089
R7185 VDD.t416 VDD.n3118 8.45089
R7186 VDD.n3342 VDD.n3341 8.45089
R7187 VDD.n3340 VDD.n3125 8.45089
R7188 VDD.n3339 VDD.n3338 8.45089
R7189 VDD.n3329 VDD.n3126 8.45089
R7190 VDD.n3331 VDD.n3330 8.45089
R7191 VDD.n3328 VDD.n3133 8.45089
R7192 VDD.n3327 VDD.n3326 8.45089
R7193 VDD.n3316 VDD.n3134 8.45089
R7194 VDD.n3318 VDD.n3317 8.45089
R7195 VDD.n3315 VDD.n3142 8.45089
R7196 VDD.n3314 VDD.n3313 8.45089
R7197 VDD.n3305 VDD.n3143 8.45089
R7198 VDD.n3307 VDD.n3306 8.45089
R7199 VDD.n3387 VDD.n3097 8.45089
R7200 VDD.n3390 VDD.n3389 8.45089
R7201 VDD.n3389 VDD.n3388 8.45089
R7202 VDD.n2906 VDD.n1938 8.45089
R7203 VDD.n1934 VDD.n1933 8.45089
R7204 VDD.n2916 VDD.n1932 8.45089
R7205 VDD.n1926 VDD.n1925 8.45089
R7206 VDD.n2925 VDD.n2924 8.45089
R7207 VDD.n2918 VDD.n2917 8.45089
R7208 VDD.n2915 VDD.n2914 8.45089
R7209 VDD.n2908 VDD.n2907 8.45089
R7210 VDD.n2905 VDD.n2904 8.45089
R7211 VDD.n2927 VDD.n1919 8.45089
R7212 VDD.n2936 VDD.n2935 8.45089
R7213 VDD.n2940 VDD.n2939 8.45089
R7214 VDD.n2947 VDD.n2946 8.45089
R7215 VDD.n2952 VDD.n2951 8.45089
R7216 VDD.n2948 VDD.n1911 8.45089
R7217 VDD.n2938 VDD.n1913 8.45089
R7218 VDD.n2937 VDD.n1918 8.45089
R7219 VDD.n2929 VDD.n2928 8.45089
R7220 VDD.n2997 VDD.n1876 8.45089
R7221 VDD.n3007 VDD.n1875 8.45089
R7222 VDD.n3008 VDD.n1870 8.45089
R7223 VDD.n3018 VDD.n1869 8.45089
R7224 VDD.n3023 VDD.n3019 8.45089
R7225 VDD.n3017 VDD.n3016 8.45089
R7226 VDD.n3010 VDD.n3009 8.45089
R7227 VDD.n3006 VDD.n3005 8.45089
R7228 VDD.n2999 VDD.n2998 8.45089
R7229 VDD.n3070 VDD.n3069 8.45089
R7230 VDD.n3077 VDD.n3076 8.45089
R7231 VDD.n3081 VDD.n3080 8.45089
R7232 VDD.n3088 VDD.n3087 8.45089
R7233 VDD.n3091 VDD.n3090 8.45089
R7234 VDD.n3089 VDD.n1827 8.45089
R7235 VDD.n3079 VDD.n1828 8.45089
R7236 VDD.n3078 VDD.n1833 8.45089
R7237 VDD.n3068 VDD.n1834 8.45089
R7238 VDD.n1289 VDD.n1288 8.45089
R7239 VDD.n1288 VDD.n1287 8.45089
R7240 VDD.n1304 VDD.n1303 8.45089
R7241 VDD.n1280 VDD.n1279 8.45089
R7242 VDD.n1308 VDD.n1275 8.45089
R7243 VDD.n1308 VDD.n1307 8.45089
R7244 VDD.n1318 VDD.n1317 8.45089
R7245 VDD.n1322 VDD.n1321 8.45089
R7246 VDD.n1329 VDD.n1328 8.45089
R7247 VDD.n1332 VDD.n1331 8.45089
R7248 VDD.n1339 VDD.n1338 8.45089
R7249 VDD.n1343 VDD.n1342 8.45089
R7250 VDD.n1350 VDD.n1349 8.45089
R7251 VDD.n1351 VDD.n1251 8.45089
R7252 VDD.n1354 VDD.n1353 8.45089
R7253 VDD.n1341 VDD.n1252 8.45089
R7254 VDD.n1340 VDD.n1258 8.45089
R7255 VDD.n1260 VDD.n1259 8.45089
R7256 VDD.n1330 VDD.n1265 8.45089
R7257 VDD.n1320 VDD.n1266 8.45089
R7258 VDD.n1319 VDD.n1271 8.45089
R7259 VDD.n1306 VDD.n1272 8.45089
R7260 VDD.n1309 VDD.n1305 8.45089
R7261 VDD.n1352 VDD.n1245 8.45089
R7262 VDD.n1363 VDD.n1244 8.45089
R7263 VDD.n1365 VDD.n1364 8.45089
R7264 VDD.n1381 VDD.n1380 8.45089
R7265 VDD.n1238 VDD.n1237 8.45089
R7266 VDD.n1385 VDD.n1233 8.45089
R7267 VDD.n1385 VDD.n1384 8.45089
R7268 VDD.n1395 VDD.n1394 8.45089
R7269 VDD.n1399 VDD.n1398 8.45089
R7270 VDD.n1406 VDD.n1405 8.45089
R7271 VDD.n1409 VDD.n1408 8.45089
R7272 VDD.n1416 VDD.n1415 8.45089
R7273 VDD.n1420 VDD.n1419 8.45089
R7274 VDD.n1427 VDD.n1426 8.45089
R7275 VDD.n1428 VDD.n1209 8.45089
R7276 VDD.n1431 VDD.n1430 8.45089
R7277 VDD.n1418 VDD.n1210 8.45089
R7278 VDD.n1417 VDD.n1216 8.45089
R7279 VDD.n1218 VDD.n1217 8.45089
R7280 VDD.n1407 VDD.n1223 8.45089
R7281 VDD.n1397 VDD.n1224 8.45089
R7282 VDD.n1396 VDD.n1229 8.45089
R7283 VDD.n1383 VDD.n1230 8.45089
R7284 VDD.n1386 VDD.n1382 8.45089
R7285 VDD.n1429 VDD.n1203 8.45089
R7286 VDD.n1440 VDD.n1202 8.45089
R7287 VDD.n1442 VDD.n1441 8.45089
R7288 VDD.n1458 VDD.n1457 8.45089
R7289 VDD.n1196 VDD.n1195 8.45089
R7290 VDD.n1462 VDD.n1191 8.45089
R7291 VDD.n1462 VDD.n1461 8.45089
R7292 VDD.n1472 VDD.n1471 8.45089
R7293 VDD.n1476 VDD.n1475 8.45089
R7294 VDD.n1483 VDD.n1482 8.45089
R7295 VDD.n1486 VDD.n1485 8.45089
R7296 VDD.n1493 VDD.n1492 8.45089
R7297 VDD.n1497 VDD.n1496 8.45089
R7298 VDD.n1504 VDD.n1503 8.45089
R7299 VDD.n1505 VDD.n1167 8.45089
R7300 VDD.n1508 VDD.n1507 8.45089
R7301 VDD.n1495 VDD.n1168 8.45089
R7302 VDD.n1494 VDD.n1174 8.45089
R7303 VDD.n1176 VDD.n1175 8.45089
R7304 VDD.n1484 VDD.n1181 8.45089
R7305 VDD.n1474 VDD.n1182 8.45089
R7306 VDD.n1473 VDD.n1187 8.45089
R7307 VDD.n1460 VDD.n1188 8.45089
R7308 VDD.n1463 VDD.n1459 8.45089
R7309 VDD.n1506 VDD.n1161 8.45089
R7310 VDD.n1517 VDD.n1160 8.45089
R7311 VDD.n1519 VDD.n1518 8.45089
R7312 VDD.n1535 VDD.n1534 8.45089
R7313 VDD.n1154 VDD.n1153 8.45089
R7314 VDD.n1539 VDD.n1149 8.45089
R7315 VDD.n1539 VDD.n1538 8.45089
R7316 VDD.n1549 VDD.n1548 8.45089
R7317 VDD.n1553 VDD.n1552 8.45089
R7318 VDD.n1560 VDD.n1559 8.45089
R7319 VDD.n1563 VDD.n1562 8.45089
R7320 VDD.n1570 VDD.n1569 8.45089
R7321 VDD.n1574 VDD.n1573 8.45089
R7322 VDD.n1581 VDD.n1580 8.45089
R7323 VDD.n1582 VDD.n1125 8.45089
R7324 VDD.n1585 VDD.n1584 8.45089
R7325 VDD.n1572 VDD.n1126 8.45089
R7326 VDD.n1571 VDD.n1132 8.45089
R7327 VDD.n1134 VDD.n1133 8.45089
R7328 VDD.n1561 VDD.n1139 8.45089
R7329 VDD.n1551 VDD.n1140 8.45089
R7330 VDD.n1550 VDD.n1145 8.45089
R7331 VDD.n1537 VDD.n1146 8.45089
R7332 VDD.n1540 VDD.n1536 8.45089
R7333 VDD.n1583 VDD.n1119 8.45089
R7334 VDD.n1594 VDD.n1118 8.45089
R7335 VDD.n1596 VDD.n1595 8.45089
R7336 VDD.n1612 VDD.n1611 8.45089
R7337 VDD.n1112 VDD.n1111 8.45089
R7338 VDD.n1616 VDD.n1107 8.45089
R7339 VDD.n1616 VDD.n1615 8.45089
R7340 VDD.n1626 VDD.n1625 8.45089
R7341 VDD.n1630 VDD.n1629 8.45089
R7342 VDD.n1637 VDD.n1636 8.45089
R7343 VDD.n1640 VDD.n1639 8.45089
R7344 VDD.n1647 VDD.n1646 8.45089
R7345 VDD.n1651 VDD.n1650 8.45089
R7346 VDD.n1658 VDD.n1657 8.45089
R7347 VDD.n1659 VDD.n1083 8.45089
R7348 VDD.n1662 VDD.n1661 8.45089
R7349 VDD.n1649 VDD.n1084 8.45089
R7350 VDD.n1648 VDD.n1090 8.45089
R7351 VDD.n1092 VDD.n1091 8.45089
R7352 VDD.n1638 VDD.n1097 8.45089
R7353 VDD.n1628 VDD.n1098 8.45089
R7354 VDD.n1627 VDD.n1103 8.45089
R7355 VDD.n1614 VDD.n1104 8.45089
R7356 VDD.n1617 VDD.n1613 8.45089
R7357 VDD.n1660 VDD.n1077 8.45089
R7358 VDD.n1671 VDD.n1076 8.45089
R7359 VDD.n1673 VDD.n1672 8.45089
R7360 VDD.n1689 VDD.n1688 8.45089
R7361 VDD.n1070 VDD.n1069 8.45089
R7362 VDD.n1693 VDD.n1065 8.45089
R7363 VDD.n1693 VDD.n1692 8.45089
R7364 VDD.n1703 VDD.n1702 8.45089
R7365 VDD.n1707 VDD.n1706 8.45089
R7366 VDD.n1714 VDD.n1713 8.45089
R7367 VDD.n1717 VDD.n1716 8.45089
R7368 VDD.n1724 VDD.n1723 8.45089
R7369 VDD.n1729 VDD.n1728 8.45089
R7370 VDD.n1726 VDD.n1040 8.45089
R7371 VDD.n1738 VDD.n1737 8.45089
R7372 VDD.n1739 VDD.n1039 8.45089
R7373 VDD.n1727 VDD.n1048 8.45089
R7374 VDD.n1725 VDD.n1047 8.45089
R7375 VDD.n1050 VDD.n1049 8.45089
R7376 VDD.n1715 VDD.n1055 8.45089
R7377 VDD.n1705 VDD.n1056 8.45089
R7378 VDD.n1704 VDD.n1061 8.45089
R7379 VDD.n1691 VDD.n1062 8.45089
R7380 VDD.n1694 VDD.n1690 8.45089
R7381 VDD.n1741 VDD.n1740 8.45089
R7382 VDD.n1749 VDD.n1748 8.45089
R7383 VDD.n1750 VDD.n1031 8.45089
R7384 VDD.n1753 VDD.n1752 8.45089
R7385 VDD.n1754 VDD.n1751 8.45089
R7386 VDD.n1023 VDD.n1022 8.45089
R7387 VDD.n1772 VDD.n1023 8.45089
R7388 VDD.n1773 VDD.n1021 8.45089
R7389 VDD.n1785 VDD.n1784 8.45089
R7390 VDD.n1788 VDD.n1787 8.45089
R7391 VDD.n1795 VDD.n1794 8.45089
R7392 VDD.n1799 VDD.n1798 8.45089
R7393 VDD.n1808 VDD.n1807 8.45089
R7394 VDD.n1811 VDD.n1810 8.45089
R7395 VDD.n999 VDD.n998 8.45089
R7396 VDD.n1819 VDD.n1818 8.45089
R7397 VDD.n1809 VDD.n1003 8.45089
R7398 VDD.n1797 VDD.n1004 8.45089
R7399 VDD.n1796 VDD.n1008 8.45089
R7400 VDD.n1010 VDD.n1009 8.45089
R7401 VDD.n1786 VDD.n1015 8.45089
R7402 VDD.n1017 VDD.n1016 8.45089
R7403 VDD.n1775 VDD.n1774 8.45089
R7404 VDD.n1771 VDD.n1770 8.45089
R7405 VDD.n1820 VDD.n997 8.45089
R7406 VDD.n1822 VDD.n1821 8.45089
R7407 VDD.n344 VDD.n343 8.45089
R7408 VDD.n343 VDD.n342 8.45089
R7409 VDD.n349 VDD.n348 8.45089
R7410 VDD.n357 VDD.n356 8.45089
R7411 VDD.n365 VDD.n364 8.45089
R7412 VDD.n374 VDD.n373 8.45089
R7413 VDD.n383 VDD.n382 8.45089
R7414 VDD.n388 VDD.n387 8.45089
R7415 VDD.n424 VDD.n423 8.45089
R7416 VDD.n430 VDD.n429 8.45089
R7417 VDD.n437 VDD.n10 8.45089
R7418 VDD.n448 VDD.n447 8.45089
R7419 VDD.n457 VDD.n456 8.45089
R7420 VDD.n487 VDD.n486 8.45089
R7421 VDD.n486 VDD.n485 8.45089
R7422 VDD.n492 VDD.n491 8.45089
R7423 VDD.n500 VDD.n499 8.45089
R7424 VDD.n508 VDD.n507 8.45089
R7425 VDD.n517 VDD.n516 8.45089
R7426 VDD.n526 VDD.n525 8.45089
R7427 VDD.n531 VDD.n530 8.45089
R7428 VDD.n557 VDD.n556 8.45089
R7429 VDD.n563 VDD.n562 8.45089
R7430 VDD.n570 VDD.n7 8.45089
R7431 VDD.n581 VDD.n580 8.45089
R7432 VDD.n590 VDD.n589 8.45089
R7433 VDD.n620 VDD.n619 8.45089
R7434 VDD.n619 VDD.n618 8.45089
R7435 VDD.n625 VDD.n624 8.45089
R7436 VDD.n633 VDD.n632 8.45089
R7437 VDD.n641 VDD.n640 8.45089
R7438 VDD.n650 VDD.n649 8.45089
R7439 VDD.n659 VDD.n658 8.45089
R7440 VDD.n664 VDD.n663 8.45089
R7441 VDD.n692 VDD.n691 8.45089
R7442 VDD.n698 VDD.n697 8.45089
R7443 VDD.n705 VDD.n4 8.45089
R7444 VDD.n716 VDD.n715 8.45089
R7445 VDD.n725 VDD.n724 8.45089
R7446 VDD.n755 VDD.n754 8.45089
R7447 VDD.n754 VDD.n753 8.45089
R7448 VDD.n760 VDD.n759 8.45089
R7449 VDD.n768 VDD.n767 8.45089
R7450 VDD.n776 VDD.n775 8.45089
R7451 VDD.n785 VDD.n784 8.45089
R7452 VDD.n794 VDD.n793 8.45089
R7453 VDD.n799 VDD.n798 8.45089
R7454 VDD.n835 VDD.n834 8.45089
R7455 VDD.n841 VDD.n840 8.45089
R7456 VDD.n848 VDD.n1 8.45089
R7457 VDD.n859 VDD.n858 8.45089
R7458 VDD.n868 VDD.n867 8.45089
R7459 VDD.n898 VDD.n897 8.45089
R7460 VDD.n897 VDD.n896 8.45089
R7461 VDD.n903 VDD.n902 8.45089
R7462 VDD.n911 VDD.n910 8.45089
R7463 VDD.n919 VDD.n918 8.45089
R7464 VDD.n928 VDD.n927 8.45089
R7465 VDD.n937 VDD.n936 8.45089
R7466 VDD.n942 VDD.n941 8.45089
R7467 VDD.n981 VDD.n980 8.45089
R7468 VDD.n987 VDD.n986 8.45089
R7469 VDD.n977 VDD.n976 8.45089
R7470 VDD.n933 VDD.n932 8.45089
R7471 VDD.n923 VDD.n922 8.45089
R7472 VDD.n915 VDD.n914 8.45089
R7473 VDD.n907 VDD.n906 8.45089
R7474 VDD.n872 VDD.n871 8.45089
R7475 VDD.n864 VDD.n863 8.45089
R7476 VDD.n855 VDD.n854 8.45089
R7477 VDD.n847 VDD.n846 8.45089
R7478 VDD.n831 VDD.n830 8.45089
R7479 VDD.n790 VDD.n789 8.45089
R7480 VDD.n780 VDD.n779 8.45089
R7481 VDD.n772 VDD.n771 8.45089
R7482 VDD.n764 VDD.n763 8.45089
R7483 VDD.n729 VDD.n728 8.45089
R7484 VDD.n721 VDD.n720 8.45089
R7485 VDD.n712 VDD.n711 8.45089
R7486 VDD.n704 VDD.n703 8.45089
R7487 VDD.n668 VDD.n667 8.45089
R7488 VDD.n688 VDD.n687 8.45089
R7489 VDD.n655 VDD.n654 8.45089
R7490 VDD.n645 VDD.n644 8.45089
R7491 VDD.n637 VDD.n636 8.45089
R7492 VDD.n629 VDD.n628 8.45089
R7493 VDD.n594 VDD.n593 8.45089
R7494 VDD.n586 VDD.n585 8.45089
R7495 VDD.n577 VDD.n576 8.45089
R7496 VDD.n569 VDD.n568 8.45089
R7497 VDD.n553 VDD.n552 8.45089
R7498 VDD.n535 VDD.n534 8.45089
R7499 VDD.n522 VDD.n521 8.45089
R7500 VDD.n512 VDD.n511 8.45089
R7501 VDD.n504 VDD.n503 8.45089
R7502 VDD.n496 VDD.n495 8.45089
R7503 VDD.n461 VDD.n460 8.45089
R7504 VDD.n453 VDD.n452 8.45089
R7505 VDD.n444 VDD.n443 8.45089
R7506 VDD.n436 VDD.n435 8.45089
R7507 VDD.n420 VDD.n419 8.45089
R7508 VDD.n379 VDD.n378 8.45089
R7509 VDD.n369 VDD.n368 8.45089
R7510 VDD.n361 VDD.n360 8.45089
R7511 VDD.n353 VDD.n352 8.45089
R7512 VDD.n21 VDD.n20 8.45089
R7513 VDD.n27 VDD.n26 8.45089
R7514 VDD.n26 VDD.n25 8.45089
R7515 VDD.n19 VDD.n18 8.45089
R7516 VDD.n30 VDD.n29 8.45089
R7517 VDD.n39 VDD.n38 8.45089
R7518 VDD.n43 VDD.n42 8.45089
R7519 VDD.n35 VDD.n34 8.45089
R7520 VDD.n69 VDD.n68 8.45089
R7521 VDD.n68 VDD.n67 8.45089
R7522 VDD.n74 VDD.n73 8.45089
R7523 VDD.n82 VDD.n81 8.45089
R7524 VDD.n90 VDD.n89 8.45089
R7525 VDD.n99 VDD.n98 8.45089
R7526 VDD.n108 VDD.n107 8.45089
R7527 VDD.n113 VDD.n112 8.45089
R7528 VDD.n146 VDD.n145 8.45089
R7529 VDD.n152 VDD.n151 8.45089
R7530 VDD.n159 VDD.n15 8.45089
R7531 VDD.n166 VDD.n165 8.45089
R7532 VDD.n158 VDD.n157 8.45089
R7533 VDD.n136 VDD.n135 8.45089
R7534 VDD.n142 VDD.n141 8.45089
R7535 VDD.n104 VDD.n103 8.45089
R7536 VDD.n94 VDD.n93 8.45089
R7537 VDD.n86 VDD.n85 8.45089
R7538 VDD.n78 VDD.n77 8.45089
R7539 VDD.n170 VDD.n169 8.45089
R7540 VDD.n179 VDD.n178 8.45089
R7541 VDD.n183 VDD.n182 8.45089
R7542 VDD.n175 VDD.n174 8.45089
R7543 VDD.n209 VDD.n208 8.45089
R7544 VDD.n208 VDD.n207 8.45089
R7545 VDD.n214 VDD.n213 8.45089
R7546 VDD.n222 VDD.n221 8.45089
R7547 VDD.n230 VDD.n229 8.45089
R7548 VDD.n276 VDD.n275 8.45089
R7549 VDD.n280 VDD.n279 8.45089
R7550 VDD.n286 VDD.n285 8.45089
R7551 VDD.n296 VDD.n295 8.45089
R7552 VDD.n305 VDD.n304 8.45089
R7553 VDD.n314 VDD.n313 8.45089
R7554 VDD.n318 VDD.n317 8.45089
R7555 VDD.n310 VDD.n309 8.45089
R7556 VDD.n301 VDD.n300 8.45089
R7557 VDD.n293 VDD.n292 8.45089
R7558 VDD.n234 VDD.n233 8.45089
R7559 VDD.n226 VDD.n225 8.45089
R7560 VDD.n218 VDD.n217 8.45089
R7561 VDD.n239 VDD.n238 8.45089
R7562 VDD.n248 VDD.n247 8.45089
R7563 VDD.n244 VDD.n243 8.45089
R7564 VDD.n254 VDD.n253 8.45089
R7565 VDD.n253 VDD.n252 8.45089
R7566 VDD.n272 VDD.n271 8.45089
R7567 VDD.n263 VDD.n262 8.45089
R7568 VDD.n3381 VDD.n3098 8.45089
R7569 VDD.n3380 VDD.n3379 8.45089
R7570 VDD.n3372 VDD.n3102 8.45089
R7571 VDD.n3104 VDD.n3103 8.45089
R7572 VDD.n3367 VDD.n3366 8.45089
R7573 VDD.n3109 VDD.n3107 8.45089
R7574 VDD.n3361 VDD.n3360 8.45089
R7575 VDD.n3356 VDD.n3110 8.45089
R7576 VDD.n3355 VDD.n3354 8.45089
R7577 VDD.n3121 VDD.n3117 8.45089
R7578 VDD.n3349 VDD.n3348 8.45089
R7579 VDD.n3344 VDD.n3118 8.45089
R7580 VDD.n3343 VDD.n3342 8.45089
R7581 VDD.n3129 VDD.n3125 8.45089
R7582 VDD.n3338 VDD.n3337 8.45089
R7583 VDD.n3333 VDD.n3126 8.45089
R7584 VDD.n3332 VDD.n3331 8.45089
R7585 VDD.n3322 VDD.n3133 8.45089
R7586 VDD.n3326 VDD.n3325 8.45089
R7587 VDD.n3135 VDD.n3134 8.45089
R7588 VDD.n3319 VDD.n3318 8.45089
R7589 VDD.n3142 VDD.n3139 8.45089
R7590 VDD.n3313 VDD.n3312 8.45089
R7591 VDD.n3144 VDD.n3143 8.45089
R7592 VDD.n3308 VDD.n3307 8.45089
R7593 VDD.n3151 VDD.n3148 8.45089
R7594 VDD.n3300 VDD.n3299 8.45089
R7595 VDD.n3291 VDD.n3158 8.45089
R7596 VDD.n3290 VDD.n3289 8.45089
R7597 VDD.n3282 VDD.n3162 8.45089
R7598 VDD.n3164 VDD.n3163 8.45089
R7599 VDD.n3277 VDD.n3276 8.45089
R7600 VDD.n3169 VDD.n3167 8.45089
R7601 VDD.n3271 VDD.n3270 8.45089
R7602 VDD.n3266 VDD.n3170 8.45089
R7603 VDD.n3265 VDD.n3264 8.45089
R7604 VDD.n3181 VDD.n3177 8.45089
R7605 VDD.n3259 VDD.n3258 8.45089
R7606 VDD.n3254 VDD.n3178 8.45089
R7607 VDD.n3253 VDD.n3252 8.45089
R7608 VDD.n3189 VDD.n3185 8.45089
R7609 VDD.n3248 VDD.n3247 8.45089
R7610 VDD.n3243 VDD.n3186 8.45089
R7611 VDD.n3242 VDD.n3241 8.45089
R7612 VDD.n3232 VDD.n3193 8.45089
R7613 VDD.n3236 VDD.n3235 8.45089
R7614 VDD.n3195 VDD.n3194 8.45089
R7615 VDD.n3229 VDD.n3228 8.45089
R7616 VDD.n3202 VDD.n3199 8.45089
R7617 VDD.n3223 VDD.n3222 8.45089
R7618 VDD.n3204 VDD.n3203 8.45089
R7619 VDD.n3218 VDD.n3217 8.45089
R7620 VDD.n3211 VDD.n3208 8.45089
R7621 VDD.n2904 VDD.n2903 8.45089
R7622 VDD.n2909 VDD.n2908 8.45089
R7623 VDD.n2914 VDD.n2913 8.45089
R7624 VDD.n2919 VDD.n2918 8.45089
R7625 VDD.n2924 VDD.n2923 8.45089
R7626 VDD.n2930 VDD.n2929 8.45089
R7627 VDD.n2931 VDD.n1919 8.45089
R7628 VDD.n1918 VDD.n1917 8.45089
R7629 VDD.n1914 VDD.n1913 8.45089
R7630 VDD.n1915 VDD.n1911 8.45089
R7631 VDD.n3000 VDD.n2999 8.45089
R7632 VDD.n3005 VDD.n3004 8.45089
R7633 VDD.n3011 VDD.n3010 8.45089
R7634 VDD.n3016 VDD.n3015 8.45089
R7635 VDD.n3024 VDD.n3023 8.45089
R7636 VDD.n3072 VDD.n1834 8.45089
R7637 VDD.n1833 VDD.n1832 8.45089
R7638 VDD.n1829 VDD.n1828 8.45089
R7639 VDD.n1830 VDD.n1827 8.45089
R7640 VDD.n3087 VDD.n3086 8.45089
R7641 VDD.n3082 VDD.n3081 8.45089
R7642 VDD.n3076 VDD.n3075 8.45089
R7643 VDD.n3071 VDD.n3070 8.45089
R7644 VDD.n1872 VDD.n1869 8.45089
R7645 VDD.n1871 VDD.n1870 8.45089
R7646 VDD.n1875 VDD.n1874 8.45089
R7647 VDD.n3001 VDD.n1876 8.45089
R7648 VDD.n2953 VDD.n2952 8.45089
R7649 VDD.n2946 VDD.n2945 8.45089
R7650 VDD.n2941 VDD.n2940 8.45089
R7651 VDD.n2935 VDD.n2934 8.45089
R7652 VDD.n1927 VDD.n1926 8.45089
R7653 VDD.n1932 VDD.n1929 8.45089
R7654 VDD.n1935 VDD.n1934 8.45089
R7655 VDD.n1938 VDD.n1937 8.45089
R7656 VDD.n1286 VDD.n1283 8.45089
R7657 VDD.n1281 VDD.n1280 8.45089
R7658 VDD.n1310 VDD.n1309 8.45089
R7659 VDD.n1315 VDD.n1272 8.45089
R7660 VDD.n1271 VDD.n1270 8.45089
R7661 VDD.n1267 VDD.n1266 8.45089
R7662 VDD.n1268 VDD.n1265 8.45089
R7663 VDD.n1261 VDD.n1260 8.45089
R7664 VDD.n1253 VDD.n1252 8.45089
R7665 VDD.n1355 VDD.n1354 8.45089
R7666 VDD.n1362 VDD.n1361 8.45089
R7667 VDD VDD.n1362 8.45089
R7668 VDD.n1366 VDD.n1365 8.45089
R7669 VDD.n1239 VDD.n1238 8.45089
R7670 VDD.n1387 VDD.n1386 8.45089
R7671 VDD.n1392 VDD.n1230 8.45089
R7672 VDD.n1229 VDD.n1228 8.45089
R7673 VDD.n1225 VDD.n1224 8.45089
R7674 VDD.n1226 VDD.n1223 8.45089
R7675 VDD.n1219 VDD.n1218 8.45089
R7676 VDD.n1211 VDD.n1210 8.45089
R7677 VDD.n1432 VDD.n1431 8.45089
R7678 VDD.n1439 VDD.n1438 8.45089
R7679 VDD VDD.n1439 8.45089
R7680 VDD.n1443 VDD.n1442 8.45089
R7681 VDD.n1197 VDD.n1196 8.45089
R7682 VDD.n1464 VDD.n1463 8.45089
R7683 VDD.n1469 VDD.n1188 8.45089
R7684 VDD.n1187 VDD.n1186 8.45089
R7685 VDD.n1183 VDD.n1182 8.45089
R7686 VDD.n1184 VDD.n1181 8.45089
R7687 VDD.n1177 VDD.n1176 8.45089
R7688 VDD.n1169 VDD.n1168 8.45089
R7689 VDD.n1509 VDD.n1508 8.45089
R7690 VDD.n1516 VDD.n1515 8.45089
R7691 VDD VDD.n1516 8.45089
R7692 VDD.n1520 VDD.n1519 8.45089
R7693 VDD.n1155 VDD.n1154 8.45089
R7694 VDD.n1541 VDD.n1540 8.45089
R7695 VDD.n1546 VDD.n1146 8.45089
R7696 VDD.n1145 VDD.n1144 8.45089
R7697 VDD.n1141 VDD.n1140 8.45089
R7698 VDD.n1142 VDD.n1139 8.45089
R7699 VDD.n1135 VDD.n1134 8.45089
R7700 VDD.n1127 VDD.n1126 8.45089
R7701 VDD.n1586 VDD.n1585 8.45089
R7702 VDD.n1593 VDD.n1592 8.45089
R7703 VDD VDD.n1593 8.45089
R7704 VDD.n1597 VDD.n1596 8.45089
R7705 VDD.n1113 VDD.n1112 8.45089
R7706 VDD.n1618 VDD.n1617 8.45089
R7707 VDD.n1623 VDD.n1104 8.45089
R7708 VDD.n1103 VDD.n1102 8.45089
R7709 VDD.n1099 VDD.n1098 8.45089
R7710 VDD.n1100 VDD.n1097 8.45089
R7711 VDD.n1093 VDD.n1092 8.45089
R7712 VDD.n1085 VDD.n1084 8.45089
R7713 VDD.n1663 VDD.n1662 8.45089
R7714 VDD.n1670 VDD.n1669 8.45089
R7715 VDD VDD.n1670 8.45089
R7716 VDD.n1674 VDD.n1673 8.45089
R7717 VDD.n1071 VDD.n1070 8.45089
R7718 VDD.n1695 VDD.n1694 8.45089
R7719 VDD.n1700 VDD.n1062 8.45089
R7720 VDD.n1061 VDD.n1060 8.45089
R7721 VDD.n1057 VDD.n1056 8.45089
R7722 VDD.n1058 VDD.n1055 8.45089
R7723 VDD.n1051 VDD.n1050 8.45089
R7724 VDD.n1048 VDD.n1042 8.45089
R7725 VDD.n1039 VDD.n1038 8.45089
R7726 VDD.n1033 VDD.n1032 8.45089
R7727 VDD VDD.n1032 8.45089
R7728 VDD.n1031 VDD.n1030 8.45089
R7729 VDD.n1755 VDD.n1754 8.45089
R7730 VDD.n1770 VDD.n1769 8.45089
R7731 VDD.n1776 VDD.n1775 8.45089
R7732 VDD.n1018 VDD.n1017 8.45089
R7733 VDD.n1015 VDD.n1014 8.45089
R7734 VDD.n1790 VDD.n1010 8.45089
R7735 VDD.n1008 VDD.n1007 8.45089
R7736 VDD.n1003 VDD.n1002 8.45089
R7737 VDD.n1818 VDD.n1817 8.45089
R7738 VDD.n1821 VDD 8.45089
R7739 VDD.n1812 VDD.n1811 8.45089
R7740 VDD.n1807 VDD.n1806 8.45089
R7741 VDD.n1800 VDD.n1799 8.45089
R7742 VDD.n1794 VDD.n1793 8.45089
R7743 VDD.n1789 VDD.n1788 8.45089
R7744 VDD.n1784 VDD.n1783 8.45089
R7745 VDD.n1753 VDD.n1028 8.45089
R7746 VDD.n1748 VDD.n1747 8.45089
R7747 VDD.n1735 VDD.n1040 8.45089
R7748 VDD.n1730 VDD.n1729 8.45089
R7749 VDD.n1723 VDD.n1722 8.45089
R7750 VDD.n1718 VDD.n1717 8.45089
R7751 VDD.n1713 VDD.n1712 8.45089
R7752 VDD.n1708 VDD.n1707 8.45089
R7753 VDD.n1688 VDD.n1687 8.45089
R7754 VDD.n1079 VDD.n1076 8.45089
R7755 VDD.n1657 VDD.n1656 8.45089
R7756 VDD.n1652 VDD.n1651 8.45089
R7757 VDD.n1646 VDD.n1645 8.45089
R7758 VDD.n1641 VDD.n1640 8.45089
R7759 VDD.n1636 VDD.n1635 8.45089
R7760 VDD.n1631 VDD.n1630 8.45089
R7761 VDD.n1611 VDD.n1610 8.45089
R7762 VDD.n1121 VDD.n1118 8.45089
R7763 VDD.n1580 VDD.n1579 8.45089
R7764 VDD.n1575 VDD.n1574 8.45089
R7765 VDD.n1569 VDD.n1568 8.45089
R7766 VDD.n1564 VDD.n1563 8.45089
R7767 VDD.n1559 VDD.n1558 8.45089
R7768 VDD.n1554 VDD.n1553 8.45089
R7769 VDD.n1534 VDD.n1533 8.45089
R7770 VDD.n1163 VDD.n1160 8.45089
R7771 VDD.n1503 VDD.n1502 8.45089
R7772 VDD.n1498 VDD.n1497 8.45089
R7773 VDD.n1492 VDD.n1491 8.45089
R7774 VDD.n1487 VDD.n1486 8.45089
R7775 VDD.n1482 VDD.n1481 8.45089
R7776 VDD.n1477 VDD.n1476 8.45089
R7777 VDD.n1457 VDD.n1456 8.45089
R7778 VDD.n1205 VDD.n1202 8.45089
R7779 VDD.n1426 VDD.n1425 8.45089
R7780 VDD.n1421 VDD.n1420 8.45089
R7781 VDD.n1415 VDD.n1414 8.45089
R7782 VDD.n1410 VDD.n1409 8.45089
R7783 VDD.n1405 VDD.n1404 8.45089
R7784 VDD.n1400 VDD.n1399 8.45089
R7785 VDD.n1380 VDD.n1379 8.45089
R7786 VDD.n1247 VDD.n1244 8.45089
R7787 VDD.n1349 VDD.n1348 8.45089
R7788 VDD.n1344 VDD.n1343 8.45089
R7789 VDD.n1338 VDD.n1337 8.45089
R7790 VDD.n1333 VDD.n1332 8.45089
R7791 VDD.n1328 VDD.n1327 8.45089
R7792 VDD.n1323 VDD.n1322 8.45089
R7793 VDD.n1303 VDD.n1302 8.45089
R7794 VDD VDD.n19 8.45089
R7795 VDD.n36 VDD.n35 8.45089
R7796 VDD.n44 VDD.n43 8.45089
R7797 VDD.n79 VDD.n78 8.45089
R7798 VDD.n87 VDD.n86 8.45089
R7799 VDD.n95 VDD.n94 8.45089
R7800 VDD.n105 VDD.n104 8.45089
R7801 VDD.n114 VDD.n113 8.45089
R7802 VDD.n143 VDD.n142 8.45089
R7803 VDD.n147 VDD.n146 8.45089
R7804 VDD.n157 VDD.n16 8.45089
R7805 VDD.n167 VDD.n166 8.45089
R7806 VDD.n176 VDD.n175 8.45089
R7807 VDD.n184 VDD.n183 8.45089
R7808 VDD.n219 VDD.n218 8.45089
R7809 VDD.n227 VDD.n226 8.45089
R7810 VDD.n235 VDD.n234 8.45089
R7811 VDD.n245 VDD.n244 8.45089
R7812 VDD.n249 VDD.n248 8.45089
R7813 VDD.n231 VDD.n230 8.45089
R7814 VDD.n223 VDD.n222 8.45089
R7815 VDD.n215 VDD.n214 8.45089
R7816 VDD.n180 VDD.n179 8.45089
R7817 VDD.n161 VDD.n160 8.45089
R7818 VDD.n160 VDD 8.45089
R7819 VDD.n153 VDD.n152 8.45089
R7820 VDD.n137 VDD.n136 8.45089
R7821 VDD.n109 VDD.n108 8.45089
R7822 VDD.n91 VDD.n90 8.45089
R7823 VDD.n83 VDD.n82 8.45089
R7824 VDD.n75 VDD.n74 8.45089
R7825 VDD.n40 VDD.n39 8.45089
R7826 VDD.n264 VDD.n263 8.45089
R7827 VDD.n277 VDD.n276 8.45089
R7828 VDD.n287 VDD.n286 8.45089
R7829 VDD.n292 VDD.n291 8.45089
R7830 VDD.n302 VDD.n301 8.45089
R7831 VDD.n311 VDD.n310 8.45089
R7832 VDD.n319 VDD.n318 8.45089
R7833 VDD.n354 VDD.n353 8.45089
R7834 VDD.n362 VDD.n361 8.45089
R7835 VDD.n370 VDD.n369 8.45089
R7836 VDD.n380 VDD.n379 8.45089
R7837 VDD.n389 VDD.n388 8.45089
R7838 VDD.n421 VDD.n420 8.45089
R7839 VDD.n425 VDD.n424 8.45089
R7840 VDD.n435 VDD.n11 8.45089
R7841 VDD.n445 VDD.n444 8.45089
R7842 VDD.n454 VDD.n453 8.45089
R7843 VDD.n462 VDD.n461 8.45089
R7844 VDD.n497 VDD.n496 8.45089
R7845 VDD.n505 VDD.n504 8.45089
R7846 VDD.n513 VDD.n512 8.45089
R7847 VDD.n523 VDD.n522 8.45089
R7848 VDD.n532 VDD.n531 8.45089
R7849 VDD.n554 VDD.n553 8.45089
R7850 VDD.n564 VDD.n563 8.45089
R7851 VDD.n568 VDD.n8 8.45089
R7852 VDD.n578 VDD.n577 8.45089
R7853 VDD.n587 VDD.n586 8.45089
R7854 VDD.n595 VDD.n594 8.45089
R7855 VDD.n630 VDD.n629 8.45089
R7856 VDD.n638 VDD.n637 8.45089
R7857 VDD.n646 VDD.n645 8.45089
R7858 VDD.n656 VDD.n655 8.45089
R7859 VDD.n665 VDD.n664 8.45089
R7860 VDD.n689 VDD.n688 8.45089
R7861 VDD.n693 VDD.n692 8.45089
R7862 VDD.n703 VDD.n5 8.45089
R7863 VDD.n713 VDD.n712 8.45089
R7864 VDD.n722 VDD.n721 8.45089
R7865 VDD.n730 VDD.n729 8.45089
R7866 VDD.n765 VDD.n764 8.45089
R7867 VDD.n773 VDD.n772 8.45089
R7868 VDD.n781 VDD.n780 8.45089
R7869 VDD.n791 VDD.n790 8.45089
R7870 VDD.n800 VDD.n799 8.45089
R7871 VDD.n832 VDD.n831 8.45089
R7872 VDD.n842 VDD.n841 8.45089
R7873 VDD.n846 VDD.n2 8.45089
R7874 VDD.n856 VDD.n855 8.45089
R7875 VDD.n865 VDD.n864 8.45089
R7876 VDD.n873 VDD.n872 8.45089
R7877 VDD.n908 VDD.n907 8.45089
R7878 VDD.n916 VDD.n915 8.45089
R7879 VDD.n924 VDD.n923 8.45089
R7880 VDD.n934 VDD.n933 8.45089
R7881 VDD.n978 VDD.n977 8.45089
R7882 VDD.n982 VDD.n981 8.45089
R7883 VDD.n991 VDD.n990 8.45089
R7884 VDD.n988 VDD.n987 8.45089
R7885 VDD.n938 VDD.n937 8.45089
R7886 VDD.n920 VDD.n919 8.45089
R7887 VDD.n912 VDD.n911 8.45089
R7888 VDD.n904 VDD.n903 8.45089
R7889 VDD.n869 VDD.n868 8.45089
R7890 VDD.n850 VDD.n849 8.45089
R7891 VDD.n849 VDD 8.45089
R7892 VDD.n836 VDD.n835 8.45089
R7893 VDD.n795 VDD.n794 8.45089
R7894 VDD.n777 VDD.n776 8.45089
R7895 VDD.n769 VDD.n768 8.45089
R7896 VDD.n761 VDD.n760 8.45089
R7897 VDD.n726 VDD.n725 8.45089
R7898 VDD.n707 VDD.n706 8.45089
R7899 VDD.n706 VDD 8.45089
R7900 VDD.n699 VDD.n698 8.45089
R7901 VDD.n669 VDD.n668 8.45089
R7902 VDD.n660 VDD.n659 8.45089
R7903 VDD.n642 VDD.n641 8.45089
R7904 VDD.n634 VDD.n633 8.45089
R7905 VDD.n626 VDD.n625 8.45089
R7906 VDD.n591 VDD.n590 8.45089
R7907 VDD.n572 VDD.n571 8.45089
R7908 VDD.n571 VDD 8.45089
R7909 VDD.n558 VDD.n557 8.45089
R7910 VDD.n536 VDD.n535 8.45089
R7911 VDD.n527 VDD.n526 8.45089
R7912 VDD.n509 VDD.n508 8.45089
R7913 VDD.n501 VDD.n500 8.45089
R7914 VDD.n493 VDD.n492 8.45089
R7915 VDD.n458 VDD.n457 8.45089
R7916 VDD.n439 VDD.n438 8.45089
R7917 VDD.n438 VDD 8.45089
R7918 VDD.n431 VDD.n430 8.45089
R7919 VDD.n384 VDD.n383 8.45089
R7920 VDD.n366 VDD.n365 8.45089
R7921 VDD.n358 VDD.n357 8.45089
R7922 VDD.n350 VDD.n349 8.45089
R7923 VDD.n315 VDD.n314 8.45089
R7924 VDD.n294 VDD.n13 8.45089
R7925 VDD VDD.n294 8.45089
R7926 VDD.n281 VDD.n280 8.45089
R7927 VDD.n273 VDD.n272 8.45089
R7928 VDD.n2015 VDD.n2014 8.38671
R7929 VDD.n2891 VDD.n1945 8.38671
R7930 VDD.n1909 VDD.n1903 8.38671
R7931 VDD.n1905 VDD.n1900 8.38671
R7932 VDD.n2967 VDD.n2965 8.38671
R7933 VDD.n2966 VDD.n1896 8.38671
R7934 VDD.n2972 VDD.n2971 8.38671
R7935 VDD.n1898 VDD.n1897 8.38671
R7936 VDD.n2980 VDD.n2979 8.38671
R7937 VDD.n2983 VDD.n1888 8.38671
R7938 VDD.n1867 VDD.n1861 8.38671
R7939 VDD.n1863 VDD.n1858 8.38671
R7940 VDD.n3038 VDD.n3036 8.38671
R7941 VDD.n3037 VDD.n1854 8.38671
R7942 VDD.n3043 VDD.n3042 8.38671
R7943 VDD.n1856 VDD.n1855 8.38671
R7944 VDD.n3051 VDD.n3050 8.38671
R7945 VDD.n3054 VDD.n1846 8.38671
R7946 VDD.n1777 VDD.n1018 8.38671
R7947 VDD.n1701 VDD.n1060 8.38671
R7948 VDD.n1624 VDD.n1102 8.38671
R7949 VDD.n1547 VDD.n1144 8.38671
R7950 VDD.n1470 VDD.n1186 8.38671
R7951 VDD.n1393 VDD.n1228 8.38671
R7952 VDD.n1316 VDD.n1270 8.38671
R7953 VDD.n2959 VDD.n2958 7.94533
R7954 VDD.n3030 VDD.n3029 7.94533
R7955 VDD.n2390 VDD.t350 7.83017
R7956 VDD.n2580 VDD.t598 7.83017
R7957 VDD.n2700 VDD.t161 7.83017
R7958 VDD.n2836 VDD.t384 7.83017
R7959 VDD.n3253 VDD.n3184 7.50395
R7960 VDD.n3343 VDD.n3124 7.50395
R7961 VDD.n2454 VDD.n2167 7.05932
R7962 VDD.n2464 VDD.n2160 7.05932
R7963 VDD.n2475 VDD.n2155 7.05932
R7964 VDD.n2479 VDD.n2149 7.05932
R7965 VDD.n2491 VDD.n2147 7.05932
R7966 VDD.n2501 VDD.n2141 7.05932
R7967 VDD.n2513 VDD.n2135 7.05932
R7968 VDD.n2517 VDD.n2129 7.05932
R7969 VDD.n2529 VDD.n2127 7.05932
R7970 VDD.n195 VDD.n192 6.80365
R7971 VDD.n55 VDD.n52 6.80365
R7972 VDD.n330 VDD.n327 6.80365
R7973 VDD.n473 VDD.n470 6.80365
R7974 VDD.n606 VDD.n603 6.80365
R7975 VDD.n741 VDD.n738 6.80365
R7976 VDD.n884 VDD.n881 6.80365
R7977 VDD.n3210 VDD.n3204 6.62119
R7978 VDD.n3229 VDD.n3201 6.62119
R7979 VDD.n3150 VDD.n3144 6.62119
R7980 VDD.n3319 VDD.n3141 6.62119
R7981 VDD.n2696 VDD.n2695 6.62119
R7982 VDD.n2832 VDD.n2831 6.62119
R7983 VDD.n1450 VDD.n1449 6.5222
R7984 VDD.n1527 VDD.n1526 6.5222
R7985 VDD.n1762 VDD.n1761 6.5222
R7986 VDD.n1296 VDD.n1295 6.5213
R7987 VDD.n1373 VDD.n1372 6.5213
R7988 VDD.n1604 VDD.n1603 6.5213
R7989 VDD.n1681 VDD.n1680 6.5213
R7990 VDD.n2697 VDD.n2696 6.17981
R7991 VDD.n2833 VDD.n2832 6.17981
R7992 VDD.n3181 VDD.n3176 5.73843
R7993 VDD.n3121 VDD.n3116 5.73843
R7994 VDD.n3168 VDD.n3164 5.51774
R7995 VDD.n3108 VDD.n3104 5.51774
R7996 VDD.n1800 VDD.n1005 5.51774
R7997 VDD.n1722 VDD.n1046 5.51774
R7998 VDD.n1645 VDD.n1089 5.51774
R7999 VDD.n1568 VDD.n1131 5.51774
R8000 VDD.n1491 VDD.n1173 5.51774
R8001 VDD.n1414 VDD.n1215 5.51774
R8002 VDD.n1337 VDD.n1257 5.51774
R8003 VDD.t215 VDD.n1259 5.27828
R8004 VDD.t139 VDD.n1217 5.27828
R8005 VDD.t150 VDD.n1175 5.27828
R8006 VDD.t214 VDD.n1133 5.27828
R8007 VDD.t742 VDD.n1091 5.27828
R8008 VDD.t654 VDD.n1049 5.27828
R8009 VDD.n1796 VDD.t73 5.27828
R8010 VDD.n67 VDD.t681 5.26366
R8011 VDD.n207 VDD.t709 5.26366
R8012 VDD.n342 VDD.t189 5.26366
R8013 VDD.n485 VDD.t311 5.26366
R8014 VDD.n618 VDD.t579 5.26366
R8015 VDD.n753 VDD.t72 5.26366
R8016 VDD.n896 VDD.t481 5.26366
R8017 VDD.n2305 VDD.t37 5.22028
R8018 VDD.n2453 VDD.n2452 5.22028
R8019 VDD.n2466 VDD.n2465 5.22028
R8020 VDD.n2476 VDD.n2154 5.22028
R8021 VDD.n2478 VDD.n2148 5.22028
R8022 VDD.n2490 VDD.n2489 5.22028
R8023 VDD.n2503 VDD.n2502 5.22028
R8024 VDD.n2514 VDD.n2134 5.22028
R8025 VDD.n2516 VDD.n2128 5.22028
R8026 VDD.n2528 VDD.n2527 5.22028
R8027 VDD.t425 VDD.n1925 5.22028
R8028 VDD.n2927 VDD.t679 5.22028
R8029 VDD.n2997 VDD.t356 5.22028
R8030 VDD.n3068 VDD.t482 5.22028
R8031 VDD.n3214 VDD.n3211 4.69636
R8032 VDD.n3304 VDD.n3151 4.69636
R8033 VDD.n3054 VDD.n3053 4.6505
R8034 VDD.n3052 VDD.n3051 4.6505
R8035 VDD.n1855 VDD.n1847 4.6505
R8036 VDD.n3042 VDD.n3041 4.6505
R8037 VDD.n3040 VDD.n1854 4.6505
R8038 VDD.n3039 VDD.n3038 4.6505
R8039 VDD.n1858 VDD.n1857 4.6505
R8040 VDD.n3028 VDD.n3027 4.6505
R8041 VDD.n3026 VDD.n1861 4.6505
R8042 VDD.n2983 VDD.n2982 4.6505
R8043 VDD.n2981 VDD.n2980 4.6505
R8044 VDD.n1897 VDD.n1889 4.6505
R8045 VDD.n2971 VDD.n2970 4.6505
R8046 VDD.n2969 VDD.n1896 4.6505
R8047 VDD.n2968 VDD.n2967 4.6505
R8048 VDD.n1900 VDD.n1899 4.6505
R8049 VDD.n2957 VDD.n2956 4.6505
R8050 VDD.n2955 VDD.n1903 4.6505
R8051 VDD.n2901 VDD.n2900 4.6505
R8052 VDD.n2892 VDD.n1944 4.6505
R8053 VDD.n2889 VDD.n2888 4.6505
R8054 VDD.n2887 VDD.n2886 4.6505
R8055 VDD.n1950 VDD.n1949 4.6505
R8056 VDD.n2877 VDD.n2876 4.6505
R8057 VDD.n2875 VDD.n1953 4.6505
R8058 VDD.n2874 VDD.n2873 4.6505
R8059 VDD.n1956 VDD.n1955 4.6505
R8060 VDD.n2843 VDD.n1968 4.6505
R8061 VDD.n2829 VDD.n1976 4.6505
R8062 VDD.n1978 VDD.n1977 4.6505
R8063 VDD.n2816 VDD.n2815 4.6505
R8064 VDD.n2805 VDD.n1988 4.6505
R8065 VDD.n2792 VDD.n1995 4.6505
R8066 VDD.n1997 VDD.n1996 4.6505
R8067 VDD.n2779 VDD.n2778 4.6505
R8068 VDD.n2767 VDD.n2008 4.6505
R8069 VDD.n2754 VDD.n2009 4.6505
R8070 VDD.n2756 VDD.n2755 4.6505
R8071 VDD.n2753 VDD.n2012 4.6505
R8072 VDD.n2752 VDD.n2751 4.6505
R8073 VDD.n2017 VDD.n2016 4.6505
R8074 VDD.n2741 VDD.n2740 4.6505
R8075 VDD.n2739 VDD.n2020 4.6505
R8076 VDD.n2738 VDD.n2737 4.6505
R8077 VDD.n2023 VDD.n2022 4.6505
R8078 VDD.n2707 VDD.n2035 4.6505
R8079 VDD.n2693 VDD.n2043 4.6505
R8080 VDD.n2045 VDD.n2044 4.6505
R8081 VDD.n2680 VDD.n2679 4.6505
R8082 VDD.n2669 VDD.n2055 4.6505
R8083 VDD.n2656 VDD.n2062 4.6505
R8084 VDD.n2064 VDD.n2063 4.6505
R8085 VDD.n2643 VDD.n2642 4.6505
R8086 VDD.n2631 VDD.n2075 4.6505
R8087 VDD.n2625 VDD.n2076 4.6505
R8088 VDD.n2615 VDD.n2614 4.6505
R8089 VDD.n2084 VDD.n2083 4.6505
R8090 VDD.n2597 VDD.n2091 4.6505
R8091 VDD.n2587 VDD.n2097 4.6505
R8092 VDD.n2576 VDD.n2104 4.6505
R8093 VDD.n2106 VDD.n2105 4.6505
R8094 VDD.n2559 VDD.n2111 4.6505
R8095 VDD.n2549 VDD.n2117 4.6505
R8096 VDD.n2522 VDD.n2130 4.6505
R8097 VDD.n2508 VDD.n2138 4.6505
R8098 VDD.n2140 VDD.n2139 4.6505
R8099 VDD.n2495 VDD.n2494 4.6505
R8100 VDD.n2484 VDD.n2150 4.6505
R8101 VDD.n2471 VDD.n2157 4.6505
R8102 VDD.n2159 VDD.n2158 4.6505
R8103 VDD.n2458 VDD.n2457 4.6505
R8104 VDD.n2447 VDD.n2170 4.6505
R8105 VDD.n2434 VDD.n2175 4.6505
R8106 VDD.n2429 VDD.n2176 4.6505
R8107 VDD.n2419 VDD.n2182 4.6505
R8108 VDD.n2407 VDD.n2190 4.6505
R8109 VDD.n2192 VDD.n2191 4.6505
R8110 VDD.n2393 VDD.n2197 4.6505
R8111 VDD.n2383 VDD.n2202 4.6505
R8112 VDD.n2371 VDD.n2212 4.6505
R8113 VDD.n2214 VDD.n2213 4.6505
R8114 VDD.n2220 VDD.n2219 4.6505
R8115 VDD.n2325 VDD.n2324 4.6505
R8116 VDD.n2313 VDD.n2232 4.6505
R8117 VDD.n2299 VDD.n2239 4.6505
R8118 VDD.n2241 VDD.n2240 4.6505
R8119 VDD.n2286 VDD.n2285 4.6505
R8120 VDD.n2275 VDD.n2250 4.6505
R8121 VDD.n2260 VDD.n2258 4.6505
R8122 VDD.n1300 VDD.n1282 4.6505
R8123 VDD.n1297 VDD.n1292 4.6505
R8124 VDD.n1377 VDD.n1240 4.6505
R8125 VDD.n1374 VDD.n1369 4.6505
R8126 VDD.n1454 VDD.n1198 4.6505
R8127 VDD.n1451 VDD.n1446 4.6505
R8128 VDD.n1531 VDD.n1156 4.6505
R8129 VDD.n1528 VDD.n1523 4.6505
R8130 VDD.n1608 VDD.n1114 4.6505
R8131 VDD.n1605 VDD.n1600 4.6505
R8132 VDD.n1685 VDD.n1072 4.6505
R8133 VDD.n1682 VDD.n1677 4.6505
R8134 VDD.n1759 VDD.n1758 4.6505
R8135 VDD.n1765 VDD.n1764 4.6505
R8136 VDD.n139 VDD.n138 4.6505
R8137 VDD.n205 VDD.n204 4.6505
R8138 VDD.n189 VDD.n188 4.6505
R8139 VDD.n65 VDD.n64 4.6505
R8140 VDD.n49 VDD.n48 4.6505
R8141 VDD.n266 VDD.n265 4.6505
R8142 VDD.n417 VDD.n416 4.6505
R8143 VDD.n685 VDD.n684 4.6505
R8144 VDD.n828 VDD.n827 4.6505
R8145 VDD.n958 VDD.n957 4.6505
R8146 VDD.n974 VDD.n973 4.6505
R8147 VDD.n894 VDD.n893 4.6505
R8148 VDD.n878 VDD.n877 4.6505
R8149 VDD.n751 VDD.n750 4.6505
R8150 VDD.n735 VDD.n734 4.6505
R8151 VDD.n616 VDD.n615 4.6505
R8152 VDD.n600 VDD.n599 4.6505
R8153 VDD.n483 VDD.n482 4.6505
R8154 VDD.n467 VDD.n466 4.6505
R8155 VDD.n340 VDD.n339 4.6505
R8156 VDD.n324 VDD.n323 4.6505
R8157 VDD.n194 VDD.n191 4.53646
R8158 VDD.n54 VDD.n51 4.53646
R8159 VDD.n329 VDD.n326 4.53646
R8160 VDD.n472 VDD.n469 4.53646
R8161 VDD.n605 VDD.n602 4.53646
R8162 VDD.n740 VDD.n737 4.53646
R8163 VDD.n883 VDD.n880 4.53646
R8164 VDD.n3247 VDD.n3188 3.97291
R8165 VDD.n3337 VDD.n3128 3.97291
R8166 VDD.n2210 VDD.n2204 3.97291
R8167 VDD.n2561 VDD.n2110 3.97291
R8168 VDD VDD.n2259 3.89041
R8169 VDD.n944 VDD.n940 3.78744
R8170 VDD.n3300 VDD 3.75222
R8171 VDD.n3390 VDD 3.75222
R8172 VDD.n1790 VDD.n1012 3.75222
R8173 VDD.n1058 VDD.n1054 3.75222
R8174 VDD.n1100 VDD.n1096 3.75222
R8175 VDD.n1142 VDD.n1138 3.75222
R8176 VDD.n1184 VDD.n1180 3.75222
R8177 VDD.n1226 VDD.n1222 3.75222
R8178 VDD.n1268 VDD.n1264 3.75222
R8179 VDD.n3291 VDD 3.53153
R8180 VDD.n3381 VDD 3.53153
R8181 VDD.n2259 VDD.n2256 3.53153
R8182 VDD.n2258 VDD.n2252 3.53153
R8183 VDD.n2271 VDD.n2252 3.53153
R8184 VDD.n2277 VDD.n2250 3.53153
R8185 VDD.n2277 VDD.n2247 3.53153
R8186 VDD.n2285 VDD.n2245 3.53153
R8187 VDD.n2291 VDD.n2245 3.53153
R8188 VDD.n2297 VDD.n2241 3.53153
R8189 VDD.n2297 VDD.n2238 3.53153
R8190 VDD.n2239 VDD.n2234 3.53153
R8191 VDD.n2309 VDD.n2234 3.53153
R8192 VDD.n2315 VDD.n2232 3.53153
R8193 VDD.n2315 VDD.n2229 3.53153
R8194 VDD.n2324 VDD.n2226 3.53153
R8195 VDD.n2330 VDD.n2226 3.53153
R8196 VDD.n2358 VDD.n2220 3.53153
R8197 VDD.n2358 VDD.n2221 3.53153
R8198 VDD.n2629 VDD.n2075 3.53153
R8199 VDD.n2639 VDD.n2071 3.53153
R8200 VDD.n2648 VDD.n2647 3.53153
R8201 VDD.n2646 VDD.n2064 3.53153
R8202 VDD.n2659 VDD.n2061 3.53153
R8203 VDD.n2658 VDD.n2062 3.53153
R8204 VDD.n2666 VDD.n2665 3.53153
R8205 VDD.n2667 VDD.n2055 3.53153
R8206 VDD.n2677 VDD.n2051 3.53153
R8207 VDD.n2679 VDD.n2678 3.53153
R8208 VDD.n2685 VDD.n2684 3.53153
R8209 VDD.n2683 VDD.n2045 3.53153
R8210 VDD.n2697 VDD.n2041 3.53153
R8211 VDD.n2695 VDD.n2043 3.53153
R8212 VDD.n2704 VDD.n2703 3.53153
R8213 VDD.n2705 VDD.n2035 3.53153
R8214 VDD.n2715 VDD.n2031 3.53153
R8215 VDD.n2765 VDD.n2008 3.53153
R8216 VDD.n2775 VDD.n2004 3.53153
R8217 VDD.n2784 VDD.n2783 3.53153
R8218 VDD.n2782 VDD.n1997 3.53153
R8219 VDD.n2795 VDD.n1994 3.53153
R8220 VDD.n2794 VDD.n1995 3.53153
R8221 VDD.n2802 VDD.n2801 3.53153
R8222 VDD.n2803 VDD.n1988 3.53153
R8223 VDD.n2813 VDD.n1984 3.53153
R8224 VDD.n2815 VDD.n2814 3.53153
R8225 VDD.n2821 VDD.n2820 3.53153
R8226 VDD.n2819 VDD.n1978 3.53153
R8227 VDD.n2833 VDD.n1974 3.53153
R8228 VDD.n2831 VDD.n1976 3.53153
R8229 VDD.n2840 VDD.n2839 3.53153
R8230 VDD.n2841 VDD.n1968 3.53153
R8231 VDD.n2851 VDD.n1964 3.53153
R8232 VDD.n2634 VDD.n2072 3.52991
R8233 VDD.n2649 VDD.n2067 3.52991
R8234 VDD.n2653 VDD.n2060 3.52991
R8235 VDD.n2664 VDD.n2058 3.52991
R8236 VDD.n2672 VDD.n2052 3.52991
R8237 VDD.n2686 VDD.n2048 3.52991
R8238 VDD.n2690 VDD.n2040 3.52991
R8239 VDD.n2702 VDD.n2038 3.52991
R8240 VDD.n2710 VDD.n2032 3.52991
R8241 VDD.n2770 VDD.n2005 3.52991
R8242 VDD.n2785 VDD.n2000 3.52991
R8243 VDD.n2789 VDD.n1993 3.52991
R8244 VDD.n2800 VDD.n1991 3.52991
R8245 VDD.n2808 VDD.n1985 3.52991
R8246 VDD.n2822 VDD.n1981 3.52991
R8247 VDD.n2826 VDD.n1973 3.52991
R8248 VDD.n2838 VDD.n1971 3.52991
R8249 VDD.n2846 VDD.n1965 3.52991
R8250 VDD.n2265 VDD.n2255 3.52991
R8251 VDD.n2270 VDD.n2249 3.52991
R8252 VDD.n2282 VDD.n2248 3.52991
R8253 VDD.n2292 VDD.n2242 3.52991
R8254 VDD.n2303 VDD.n2237 3.52991
R8255 VDD.n2308 VDD.n2231 3.52991
R8256 VDD.n2320 VDD.n2230 3.52991
R8257 VDD.n2331 VDD.n2222 3.52991
R8258 VDD.n2353 VDD.n2223 3.52991
R8259 VDD.n810 VDD.n806 3.52991
R8260 VDD.n824 VDD.n820 3.52991
R8261 VDD.n682 VDD.n678 3.52991
R8262 VDD.n548 VDD.n544 3.52991
R8263 VDD.n399 VDD.n395 3.52991
R8264 VDD.n414 VDD.n410 3.52991
R8265 VDD.n124 VDD.n120 3.52991
R8266 VDD.n971 VDD.n967 3.42907
R8267 VDD.n2449 VDD.n2170 3.31084
R8268 VDD.n2449 VDD.n2166 3.31084
R8269 VDD.n2457 VDD.n2163 3.31084
R8270 VDD.n2463 VDD.n2163 3.31084
R8271 VDD.n2469 VDD.n2159 3.31084
R8272 VDD.n2469 VDD.n2156 3.31084
R8273 VDD.n2157 VDD.n2152 3.31084
R8274 VDD.n2480 VDD.n2152 3.31084
R8275 VDD.n2486 VDD.n2150 3.31084
R8276 VDD.n2486 VDD.n2146 3.31084
R8277 VDD.n2494 VDD.n2144 3.31084
R8278 VDD.n2500 VDD.n2144 3.31084
R8279 VDD.n2506 VDD.n2140 3.31084
R8280 VDD.n2506 VDD.n2136 3.31084
R8281 VDD.n2138 VDD.n2132 3.31084
R8282 VDD.n2518 VDD.n2132 3.31084
R8283 VDD.n2524 VDD.n2130 3.31084
R8284 VDD.n2524 VDD.n2126 3.31084
R8285 VDD.n3213 VDD.n3207 3.22029
R8286 VDD.n1290 VDD.n1283 3.22029
R8287 VDD.n18 VDD 3.12264
R8288 VDD.n198 VDD 3.10353
R8289 VDD.n58 VDD 3.10353
R8290 VDD.n333 VDD 3.10353
R8291 VDD.n476 VDD 3.10353
R8292 VDD.n609 VDD 3.10353
R8293 VDD.n744 VDD 3.10353
R8294 VDD.n887 VDD 3.10353
R8295 VDD.n3391 VDD.n3390 3.1005
R8296 VDD.n3384 VDD.n3383 3.1005
R8297 VDD.n3301 VDD.n3300 3.1005
R8298 VDD.n3294 VDD.n3293 3.1005
R8299 VDD.n3208 VDD.n3207 3.1005
R8300 VDD.n3219 VDD.n3218 3.1005
R8301 VDD.n3220 VDD.n3204 3.1005
R8302 VDD.n3222 VDD.n3221 3.1005
R8303 VDD.n3199 VDD.n3198 3.1005
R8304 VDD.n3230 VDD.n3229 3.1005
R8305 VDD.n3231 VDD.n3195 3.1005
R8306 VDD.n3235 VDD.n3234 3.1005
R8307 VDD.n3233 VDD.n3232 3.1005
R8308 VDD.n3242 VDD.n3190 3.1005
R8309 VDD.n3244 VDD.n3243 3.1005
R8310 VDD.n3247 VDD.n3246 3.1005
R8311 VDD.n3245 VDD.n3189 3.1005
R8312 VDD.n3253 VDD.n3182 3.1005
R8313 VDD.n3255 VDD.n3254 3.1005
R8314 VDD.n3258 VDD.n3257 3.1005
R8315 VDD.n3256 VDD.n3181 3.1005
R8316 VDD.n3265 VDD.n3174 3.1005
R8317 VDD.n3267 VDD.n3266 3.1005
R8318 VDD.n3270 VDD.n3269 3.1005
R8319 VDD.n3268 VDD.n3167 3.1005
R8320 VDD.n3278 VDD.n3277 3.1005
R8321 VDD.n3279 VDD.n3164 3.1005
R8322 VDD.n3282 VDD.n3281 3.1005
R8323 VDD.n3290 VDD.n3159 3.1005
R8324 VDD.n3292 VDD.n3291 3.1005
R8325 VDD.n3303 VDD.n3302 3.1005
R8326 VDD.n3148 VDD.n3147 3.1005
R8327 VDD.n3309 VDD.n3308 3.1005
R8328 VDD.n3310 VDD.n3144 3.1005
R8329 VDD.n3312 VDD.n3311 3.1005
R8330 VDD.n3139 VDD.n3138 3.1005
R8331 VDD.n3320 VDD.n3319 3.1005
R8332 VDD.n3321 VDD.n3135 3.1005
R8333 VDD.n3325 VDD.n3324 3.1005
R8334 VDD.n3323 VDD.n3322 3.1005
R8335 VDD.n3332 VDD.n3130 3.1005
R8336 VDD.n3334 VDD.n3333 3.1005
R8337 VDD.n3337 VDD.n3336 3.1005
R8338 VDD.n3335 VDD.n3129 3.1005
R8339 VDD.n3343 VDD.n3122 3.1005
R8340 VDD.n3345 VDD.n3344 3.1005
R8341 VDD.n3348 VDD.n3347 3.1005
R8342 VDD.n3346 VDD.n3121 3.1005
R8343 VDD.n3355 VDD.n3114 3.1005
R8344 VDD.n3357 VDD.n3356 3.1005
R8345 VDD.n3360 VDD.n3359 3.1005
R8346 VDD.n3358 VDD.n3107 3.1005
R8347 VDD.n3368 VDD.n3367 3.1005
R8348 VDD.n3369 VDD.n3104 3.1005
R8349 VDD.n3372 VDD.n3371 3.1005
R8350 VDD.n3380 VDD.n3099 3.1005
R8351 VDD.n3382 VDD.n3381 3.1005
R8352 VDD.n3092 VDD.n3091 3.1005
R8353 VDD.n2903 VDD.n2902 3.1005
R8354 VDD.n2910 VDD.n2909 3.1005
R8355 VDD.n2913 VDD.n2912 3.1005
R8356 VDD.n2920 VDD.n2919 3.1005
R8357 VDD.n2923 VDD.n2922 3.1005
R8358 VDD.n2932 VDD.n2931 3.1005
R8359 VDD.n1917 VDD.n1916 3.1005
R8360 VDD.n2943 VDD.n1914 3.1005
R8361 VDD.n1915 VDD.n1906 3.1005
R8362 VDD.n3000 VDD.n1879 3.1005
R8363 VDD.n3004 VDD.n3003 3.1005
R8364 VDD.n3012 VDD.n3011 3.1005
R8365 VDD.n3015 VDD.n3014 3.1005
R8366 VDD.n3025 VDD.n3024 3.1005
R8367 VDD.n3073 VDD.n3072 3.1005
R8368 VDD.n1832 VDD.n1831 3.1005
R8369 VDD.n3084 VDD.n1829 3.1005
R8370 VDD.n1830 VDD.n1824 3.1005
R8371 VDD.n3086 VDD.n3085 3.1005
R8372 VDD.n3083 VDD.n3082 3.1005
R8373 VDD.n3075 VDD.n3074 3.1005
R8374 VDD.n3071 VDD.n1837 3.1005
R8375 VDD.n1872 VDD.n1864 3.1005
R8376 VDD.n3013 VDD.n1871 3.1005
R8377 VDD.n1874 VDD.n1873 3.1005
R8378 VDD.n3002 VDD.n3001 3.1005
R8379 VDD.n2954 VDD.n2953 3.1005
R8380 VDD.n2945 VDD.n2944 3.1005
R8381 VDD.n2942 VDD.n2941 3.1005
R8382 VDD.n2934 VDD.n2933 3.1005
R8383 VDD.n2930 VDD.n1922 3.1005
R8384 VDD.n2921 VDD.n1927 3.1005
R8385 VDD.n1929 VDD.n1928 3.1005
R8386 VDD.n2911 VDD.n1935 3.1005
R8387 VDD.n1937 VDD.n1936 3.1005
R8388 VDD.n1823 VDD.n1822 3.1005
R8389 VDD.n1767 VDD.n1022 3.1005
R8390 VDD.n1697 VDD.n1065 3.1005
R8391 VDD.n1620 VDD.n1107 3.1005
R8392 VDD.n1543 VDD.n1149 3.1005
R8393 VDD.n1466 VDD.n1191 3.1005
R8394 VDD.n1389 VDD.n1233 3.1005
R8395 VDD.n1312 VDD.n1275 3.1005
R8396 VDD.n1291 VDD.n1281 3.1005
R8397 VDD.n1311 VDD.n1310 3.1005
R8398 VDD.n1315 VDD.n1314 3.1005
R8399 VDD.n1270 VDD.n1269 3.1005
R8400 VDD.n1325 VDD.n1267 3.1005
R8401 VDD.n1268 VDD.n1262 3.1005
R8402 VDD.n1335 VDD.n1261 3.1005
R8403 VDD.n1346 VDD.n1253 3.1005
R8404 VDD.n1356 VDD.n1355 3.1005
R8405 VDD.n1361 VDD.n1360 3.1005
R8406 VDD.n1367 VDD.n1366 3.1005
R8407 VDD.n1368 VDD.n1239 3.1005
R8408 VDD.n1388 VDD.n1387 3.1005
R8409 VDD.n1392 VDD.n1391 3.1005
R8410 VDD.n1228 VDD.n1227 3.1005
R8411 VDD.n1402 VDD.n1225 3.1005
R8412 VDD.n1226 VDD.n1220 3.1005
R8413 VDD.n1412 VDD.n1219 3.1005
R8414 VDD.n1423 VDD.n1211 3.1005
R8415 VDD.n1433 VDD.n1432 3.1005
R8416 VDD.n1438 VDD.n1437 3.1005
R8417 VDD.n1444 VDD.n1443 3.1005
R8418 VDD.n1445 VDD.n1197 3.1005
R8419 VDD.n1465 VDD.n1464 3.1005
R8420 VDD.n1469 VDD.n1468 3.1005
R8421 VDD.n1186 VDD.n1185 3.1005
R8422 VDD.n1479 VDD.n1183 3.1005
R8423 VDD.n1184 VDD.n1178 3.1005
R8424 VDD.n1489 VDD.n1177 3.1005
R8425 VDD.n1500 VDD.n1169 3.1005
R8426 VDD.n1510 VDD.n1509 3.1005
R8427 VDD.n1515 VDD.n1514 3.1005
R8428 VDD.n1521 VDD.n1520 3.1005
R8429 VDD.n1522 VDD.n1155 3.1005
R8430 VDD.n1542 VDD.n1541 3.1005
R8431 VDD.n1546 VDD.n1545 3.1005
R8432 VDD.n1144 VDD.n1143 3.1005
R8433 VDD.n1556 VDD.n1141 3.1005
R8434 VDD.n1142 VDD.n1136 3.1005
R8435 VDD.n1566 VDD.n1135 3.1005
R8436 VDD.n1577 VDD.n1127 3.1005
R8437 VDD.n1587 VDD.n1586 3.1005
R8438 VDD.n1592 VDD.n1591 3.1005
R8439 VDD.n1598 VDD.n1597 3.1005
R8440 VDD.n1599 VDD.n1113 3.1005
R8441 VDD.n1619 VDD.n1618 3.1005
R8442 VDD.n1623 VDD.n1622 3.1005
R8443 VDD.n1102 VDD.n1101 3.1005
R8444 VDD.n1633 VDD.n1099 3.1005
R8445 VDD.n1100 VDD.n1094 3.1005
R8446 VDD.n1643 VDD.n1093 3.1005
R8447 VDD.n1654 VDD.n1085 3.1005
R8448 VDD.n1664 VDD.n1663 3.1005
R8449 VDD.n1669 VDD.n1668 3.1005
R8450 VDD.n1675 VDD.n1674 3.1005
R8451 VDD.n1676 VDD.n1071 3.1005
R8452 VDD.n1696 VDD.n1695 3.1005
R8453 VDD.n1700 VDD.n1699 3.1005
R8454 VDD.n1060 VDD.n1059 3.1005
R8455 VDD.n1710 VDD.n1057 3.1005
R8456 VDD.n1058 VDD.n1052 3.1005
R8457 VDD.n1720 VDD.n1051 3.1005
R8458 VDD.n1732 VDD.n1042 3.1005
R8459 VDD.n1038 VDD.n1036 3.1005
R8460 VDD.n1745 VDD.n1033 3.1005
R8461 VDD.n1030 VDD.n1029 3.1005
R8462 VDD.n1756 VDD.n1755 3.1005
R8463 VDD.n1769 VDD.n1768 3.1005
R8464 VDD.n1776 VDD.n1019 3.1005
R8465 VDD.n1780 VDD.n1018 3.1005
R8466 VDD.n1781 VDD.n1014 3.1005
R8467 VDD.n1791 VDD.n1790 3.1005
R8468 VDD.n1007 VDD.n1006 3.1005
R8469 VDD.n1002 VDD.n1001 3.1005
R8470 VDD.n1817 VDD.n1816 3.1005
R8471 VDD.n1813 VDD.n1812 3.1005
R8472 VDD.n1806 VDD.n1805 3.1005
R8473 VDD.n1801 VDD.n1800 3.1005
R8474 VDD.n1793 VDD.n1792 3.1005
R8475 VDD.n1789 VDD.n1013 3.1005
R8476 VDD.n1783 VDD.n1782 3.1005
R8477 VDD.n1757 VDD.n1028 3.1005
R8478 VDD.n1747 VDD.n1746 3.1005
R8479 VDD.n1735 VDD.n1734 3.1005
R8480 VDD.n1731 VDD.n1730 3.1005
R8481 VDD.n1722 VDD.n1721 3.1005
R8482 VDD.n1719 VDD.n1718 3.1005
R8483 VDD.n1712 VDD.n1711 3.1005
R8484 VDD.n1709 VDD.n1708 3.1005
R8485 VDD.n1687 VDD.n1686 3.1005
R8486 VDD.n1079 VDD.n1073 3.1005
R8487 VDD.n1656 VDD.n1655 3.1005
R8488 VDD.n1653 VDD.n1652 3.1005
R8489 VDD.n1645 VDD.n1644 3.1005
R8490 VDD.n1642 VDD.n1641 3.1005
R8491 VDD.n1635 VDD.n1634 3.1005
R8492 VDD.n1632 VDD.n1631 3.1005
R8493 VDD.n1610 VDD.n1609 3.1005
R8494 VDD.n1121 VDD.n1115 3.1005
R8495 VDD.n1579 VDD.n1578 3.1005
R8496 VDD.n1576 VDD.n1575 3.1005
R8497 VDD.n1568 VDD.n1567 3.1005
R8498 VDD.n1565 VDD.n1564 3.1005
R8499 VDD.n1558 VDD.n1557 3.1005
R8500 VDD.n1555 VDD.n1554 3.1005
R8501 VDD.n1533 VDD.n1532 3.1005
R8502 VDD.n1163 VDD.n1157 3.1005
R8503 VDD.n1502 VDD.n1501 3.1005
R8504 VDD.n1499 VDD.n1498 3.1005
R8505 VDD.n1491 VDD.n1490 3.1005
R8506 VDD.n1488 VDD.n1487 3.1005
R8507 VDD.n1481 VDD.n1480 3.1005
R8508 VDD.n1478 VDD.n1477 3.1005
R8509 VDD.n1456 VDD.n1455 3.1005
R8510 VDD.n1205 VDD.n1199 3.1005
R8511 VDD.n1425 VDD.n1424 3.1005
R8512 VDD.n1422 VDD.n1421 3.1005
R8513 VDD.n1414 VDD.n1413 3.1005
R8514 VDD.n1411 VDD.n1410 3.1005
R8515 VDD.n1404 VDD.n1403 3.1005
R8516 VDD.n1401 VDD.n1400 3.1005
R8517 VDD.n1379 VDD.n1378 3.1005
R8518 VDD.n1247 VDD.n1241 3.1005
R8519 VDD.n1348 VDD.n1347 3.1005
R8520 VDD.n1345 VDD.n1344 3.1005
R8521 VDD.n1337 VDD.n1336 3.1005
R8522 VDD.n1334 VDD.n1333 3.1005
R8523 VDD.n1327 VDD.n1326 3.1005
R8524 VDD.n1324 VDD.n1323 3.1005
R8525 VDD.n1302 VDD.n1301 3.1005
R8526 VDD.n1290 VDD.n1289 3.1005
R8527 VDD.n255 VDD.n254 3.1005
R8528 VDD.n210 VDD.n209 3.1005
R8529 VDD.n70 VDD.n69 3.1005
R8530 VDD.n28 VDD.n27 3.1005
R8531 VDD.n37 VDD.n36 3.1005
R8532 VDD.n45 VDD.n44 3.1005
R8533 VDD.n80 VDD.n79 3.1005
R8534 VDD.n88 VDD.n87 3.1005
R8535 VDD.n96 VDD.n95 3.1005
R8536 VDD.n106 VDD.n105 3.1005
R8537 VDD.n115 VDD.n114 3.1005
R8538 VDD.n148 VDD.n147 3.1005
R8539 VDD.n155 VDD.n16 3.1005
R8540 VDD.n168 VDD.n167 3.1005
R8541 VDD.n177 VDD.n176 3.1005
R8542 VDD.n185 VDD.n184 3.1005
R8543 VDD.n220 VDD.n219 3.1005
R8544 VDD.n228 VDD.n227 3.1005
R8545 VDD.n236 VDD.n235 3.1005
R8546 VDD.n246 VDD.n245 3.1005
R8547 VDD.n250 VDD.n249 3.1005
R8548 VDD.n232 VDD.n231 3.1005
R8549 VDD.n224 VDD.n223 3.1005
R8550 VDD.n216 VDD.n215 3.1005
R8551 VDD.n181 VDD.n180 3.1005
R8552 VDD.n161 VDD.n156 3.1005
R8553 VDD.n154 VDD.n153 3.1005
R8554 VDD.n126 VDD.n125 3.1005
R8555 VDD.n144 VDD.n143 3.1005
R8556 VDD.n110 VDD.n109 3.1005
R8557 VDD.n92 VDD.n91 3.1005
R8558 VDD.n84 VDD.n83 3.1005
R8559 VDD.n76 VDD.n75 3.1005
R8560 VDD.n41 VDD.n40 3.1005
R8561 VDD.n345 VDD.n344 3.1005
R8562 VDD.n278 VDD.n277 3.1005
R8563 VDD.n288 VDD.n287 3.1005
R8564 VDD.n291 VDD.n290 3.1005
R8565 VDD.n303 VDD.n302 3.1005
R8566 VDD.n312 VDD.n311 3.1005
R8567 VDD.n320 VDD.n319 3.1005
R8568 VDD.n355 VDD.n354 3.1005
R8569 VDD.n363 VDD.n362 3.1005
R8570 VDD.n371 VDD.n370 3.1005
R8571 VDD.n381 VDD.n380 3.1005
R8572 VDD.n390 VDD.n389 3.1005
R8573 VDD.n426 VDD.n425 3.1005
R8574 VDD.n433 VDD.n11 3.1005
R8575 VDD.n446 VDD.n445 3.1005
R8576 VDD.n455 VDD.n454 3.1005
R8577 VDD.n463 VDD.n462 3.1005
R8578 VDD.n498 VDD.n497 3.1005
R8579 VDD.n506 VDD.n505 3.1005
R8580 VDD.n514 VDD.n513 3.1005
R8581 VDD.n524 VDD.n523 3.1005
R8582 VDD.n533 VDD.n532 3.1005
R8583 VDD.n555 VDD.n554 3.1005
R8584 VDD.n565 VDD.n564 3.1005
R8585 VDD.n566 VDD.n8 3.1005
R8586 VDD.n579 VDD.n578 3.1005
R8587 VDD.n588 VDD.n587 3.1005
R8588 VDD.n596 VDD.n595 3.1005
R8589 VDD.n631 VDD.n630 3.1005
R8590 VDD.n639 VDD.n638 3.1005
R8591 VDD.n647 VDD.n646 3.1005
R8592 VDD.n657 VDD.n656 3.1005
R8593 VDD.n666 VDD.n665 3.1005
R8594 VDD.n694 VDD.n693 3.1005
R8595 VDD.n701 VDD.n5 3.1005
R8596 VDD.n714 VDD.n713 3.1005
R8597 VDD.n723 VDD.n722 3.1005
R8598 VDD.n731 VDD.n730 3.1005
R8599 VDD.n766 VDD.n765 3.1005
R8600 VDD.n774 VDD.n773 3.1005
R8601 VDD.n782 VDD.n781 3.1005
R8602 VDD.n792 VDD.n791 3.1005
R8603 VDD.n801 VDD.n800 3.1005
R8604 VDD.n833 VDD.n832 3.1005
R8605 VDD.n843 VDD.n842 3.1005
R8606 VDD.n844 VDD.n2 3.1005
R8607 VDD.n857 VDD.n856 3.1005
R8608 VDD.n866 VDD.n865 3.1005
R8609 VDD.n874 VDD.n873 3.1005
R8610 VDD.n909 VDD.n908 3.1005
R8611 VDD.n917 VDD.n916 3.1005
R8612 VDD.n925 VDD.n924 3.1005
R8613 VDD.n935 VDD.n934 3.1005
R8614 VDD.n983 VDD.n982 3.1005
R8615 VDD.n992 VDD.n991 3.1005
R8616 VDD.n989 VDD.n988 3.1005
R8617 VDD.n979 VDD.n978 3.1005
R8618 VDD.n939 VDD.n938 3.1005
R8619 VDD.n921 VDD.n920 3.1005
R8620 VDD.n913 VDD.n912 3.1005
R8621 VDD.n905 VDD.n904 3.1005
R8622 VDD.n899 VDD.n898 3.1005
R8623 VDD.n870 VDD.n869 3.1005
R8624 VDD.n850 VDD.n845 3.1005
R8625 VDD.n837 VDD.n836 3.1005
R8626 VDD.n812 VDD.n811 3.1005
R8627 VDD.n796 VDD.n795 3.1005
R8628 VDD.n778 VDD.n777 3.1005
R8629 VDD.n770 VDD.n769 3.1005
R8630 VDD.n762 VDD.n761 3.1005
R8631 VDD.n756 VDD.n755 3.1005
R8632 VDD.n727 VDD.n726 3.1005
R8633 VDD.n707 VDD.n702 3.1005
R8634 VDD.n700 VDD.n699 3.1005
R8635 VDD.n670 VDD.n669 3.1005
R8636 VDD.n690 VDD.n689 3.1005
R8637 VDD.n661 VDD.n660 3.1005
R8638 VDD.n643 VDD.n642 3.1005
R8639 VDD.n635 VDD.n634 3.1005
R8640 VDD.n627 VDD.n626 3.1005
R8641 VDD.n621 VDD.n620 3.1005
R8642 VDD.n592 VDD.n591 3.1005
R8643 VDD.n572 VDD.n567 3.1005
R8644 VDD.n559 VDD.n558 3.1005
R8645 VDD.n537 VDD.n536 3.1005
R8646 VDD.n550 VDD.n549 3.1005
R8647 VDD.n528 VDD.n527 3.1005
R8648 VDD.n510 VDD.n509 3.1005
R8649 VDD.n502 VDD.n501 3.1005
R8650 VDD.n494 VDD.n493 3.1005
R8651 VDD.n488 VDD.n487 3.1005
R8652 VDD.n459 VDD.n458 3.1005
R8653 VDD.n439 VDD.n434 3.1005
R8654 VDD.n432 VDD.n431 3.1005
R8655 VDD.n401 VDD.n400 3.1005
R8656 VDD.n422 VDD.n421 3.1005
R8657 VDD.n385 VDD.n384 3.1005
R8658 VDD.n367 VDD.n366 3.1005
R8659 VDD.n359 VDD.n358 3.1005
R8660 VDD.n351 VDD.n350 3.1005
R8661 VDD.n316 VDD.n315 3.1005
R8662 VDD.n289 VDD.n13 3.1005
R8663 VDD.n282 VDD.n281 3.1005
R8664 VDD.n274 VDD.n273 3.1005
R8665 VDD.n3212 VDD.n3208 3.09016
R8666 VDD.n3235 VDD.n3197 3.09016
R8667 VDD.n3152 VDD.n3148 3.09016
R8668 VDD.n3325 VDD.n3137 3.09016
R8669 VDD.n2512 VDD.n2511 3.09016
R8670 VDD.n2641 VDD.n2640 3.09016
R8671 VDD.n2777 VDD.n2776 3.09016
R8672 VDD VDD.n197 3.08979
R8673 VDD VDD.n57 3.08979
R8674 VDD VDD.n332 3.08979
R8675 VDD VDD.n475 3.08979
R8676 VDD VDD.n608 3.08979
R8677 VDD VDD.n743 3.08979
R8678 VDD VDD.n886 3.08979
R8679 VDD.n2322 VDD.n2321 2.86947
R8680 VDD.n945 VDD.n944 2.64594
R8681 VDD.n1320 VDD.t741 2.63939
R8682 VDD.n1397 VDD.t729 2.63939
R8683 VDD.n1474 VDD.t186 2.63939
R8684 VDD.n1551 VDD.t96 2.63939
R8685 VDD.n1628 VDD.t702 2.63939
R8686 VDD.n1705 VDD.t423 2.63939
R8687 VDD.t428 VDD.n1786 2.63939
R8688 VDD.n85 VDD.t438 2.63208
R8689 VDD.n123 VDD.n122 2.63208
R8690 VDD.n225 VDD.t209 2.63208
R8691 VDD.n360 VDD.t682 2.63208
R8692 VDD.n398 VDD.n397 2.63208
R8693 VDD.n413 VDD.n412 2.63208
R8694 VDD.n503 VDD.t198 2.63208
R8695 VDD.n547 VDD.n546 2.63208
R8696 VDD.n636 VDD.t149 2.63208
R8697 VDD.n681 VDD.n680 2.63208
R8698 VDD.n771 VDD.t298 2.63208
R8699 VDD.n809 VDD.n808 2.63208
R8700 VDD.n823 VDD.n822 2.63208
R8701 VDD.n914 VDD.t48 2.63208
R8702 VDD.n970 VDD.n969 2.63208
R8703 VDD.n2269 VDD.n2268 2.61039
R8704 VDD.n2281 VDD.n2280 2.61039
R8705 VDD.n2294 VDD.n2293 2.61039
R8706 VDD.n2304 VDD.n2236 2.61039
R8707 VDD.n2307 VDD.n2306 2.61039
R8708 VDD.n2319 VDD.n2318 2.61039
R8709 VDD.n2333 VDD.n2332 2.61039
R8710 VDD.n2355 VDD.n2354 2.61039
R8711 VDD.t627 VDD.n2142 2.61039
R8712 VDD.n2636 VDD.n2635 2.61039
R8713 VDD.n2650 VDD.n2066 2.61039
R8714 VDD.n2652 VDD.n2059 2.61039
R8715 VDD.n2663 VDD.n2662 2.61039
R8716 VDD.n2674 VDD.n2673 2.61039
R8717 VDD.n2687 VDD.n2047 2.61039
R8718 VDD.n2689 VDD.n2039 2.61039
R8719 VDD.n2701 VDD.n2700 2.61039
R8720 VDD.n2712 VDD.n2711 2.61039
R8721 VDD.n2772 VDD.n2771 2.61039
R8722 VDD.n2786 VDD.n1999 2.61039
R8723 VDD.n2788 VDD.n1992 2.61039
R8724 VDD.n2799 VDD.n2798 2.61039
R8725 VDD.n2810 VDD.n2809 2.61039
R8726 VDD.n2823 VDD.n1980 2.61039
R8727 VDD.n2825 VDD.n1972 2.61039
R8728 VDD.n2837 VDD.n2836 2.61039
R8729 VDD.n2848 VDD.n2847 2.61039
R8730 VDD.n1256 VDD.n1254 2.55931
R8731 VDD.n1214 VDD.n1212 2.55931
R8732 VDD.n1172 VDD.n1170 2.55931
R8733 VDD.n1130 VDD.n1128 2.55931
R8734 VDD.n1088 VDD.n1086 2.55931
R8735 VDD.n1045 VDD.n1043 2.55931
R8736 VDD.n1804 VDD.n1803 2.55931
R8737 VDD.n1779 VDD.n1778 2.55931
R8738 VDD.n1698 VDD.n1064 2.55931
R8739 VDD.n1621 VDD.n1106 2.55931
R8740 VDD.n1544 VDD.n1148 2.55931
R8741 VDD.n1467 VDD.n1190 2.55931
R8742 VDD.n1390 VDD.n1232 2.55931
R8743 VDD.n1313 VDD.n1274 2.55931
R8744 VDD.n242 VDD.n241 2.55931
R8745 VDD.n102 VDD.n101 2.55931
R8746 VDD.n931 VDD.n930 2.55931
R8747 VDD.n788 VDD.n787 2.55931
R8748 VDD.n653 VDD.n652 2.55931
R8749 VDD.n520 VDD.n519 2.55931
R8750 VDD.n377 VDD.n376 2.55931
R8751 VDD.n1249 VDD.n1248 2.52719
R8752 VDD.n1207 VDD.n1206 2.52719
R8753 VDD.n1165 VDD.n1164 2.52719
R8754 VDD.n1123 VDD.n1122 2.52719
R8755 VDD.n1081 VDD.n1080 2.52719
R8756 VDD.n1733 VDD.n1041 2.52719
R8757 VDD.n1815 VDD.n1814 2.52719
R8758 VDD.n173 VDD.n172 2.52719
R8759 VDD.n33 VDD.n32 2.52719
R8760 VDD.n862 VDD.n861 2.52719
R8761 VDD.n719 VDD.n718 2.52719
R8762 VDD.n584 VDD.n583 2.52719
R8763 VDD.n451 VDD.n450 2.52719
R8764 VDD.n308 VDD.n307 2.52719
R8765 VDD.n3280 VDD.n3166 2.49102
R8766 VDD.n3155 VDD.n3153 2.49102
R8767 VDD.n3370 VDD.n3106 2.49102
R8768 VDD.n3095 VDD.n3093 2.49102
R8769 VDD.n995 VDD.n993 2.49102
R8770 VDD.n1744 VDD.n1743 2.49102
R8771 VDD.n1667 VDD.n1666 2.49102
R8772 VDD.n1590 VDD.n1589 2.49102
R8773 VDD.n1513 VDD.n1512 2.49102
R8774 VDD.n1436 VDD.n1435 2.49102
R8775 VDD.n1359 VDD.n1358 2.49102
R8776 VDD.n164 VDD.n163 2.49102
R8777 VDD.n24 VDD.n23 2.49102
R8778 VDD.n299 VDD.n298 2.49102
R8779 VDD.n442 VDD.n441 2.49102
R8780 VDD.n575 VDD.n574 2.49102
R8781 VDD.n710 VDD.n709 2.49102
R8782 VDD.n853 VDD.n852 2.49102
R8783 VDD.n194 VDD 2.46127
R8784 VDD.n54 VDD 2.46127
R8785 VDD.n329 VDD 2.46127
R8786 VDD.n472 VDD 2.46127
R8787 VDD.n605 VDD 2.46127
R8788 VDD.n740 VDD 2.46127
R8789 VDD.n883 VDD 2.46127
R8790 VDD.n2362 VDD.n2361 2.42809
R8791 VDD.n2361 VDD.n2214 2.42809
R8792 VDD.n2373 VDD.n2208 2.42809
R8793 VDD.n2373 VDD.n2212 2.42809
R8794 VDD.n2381 VDD.n2380 2.42809
R8795 VDD.n2381 VDD.n2202 2.42809
R8796 VDD.n2392 VDD.n2198 2.42809
R8797 VDD.n2393 VDD.n2392 2.42809
R8798 VDD.n2398 VDD.n2397 2.42809
R8799 VDD.n2397 VDD.n2192 2.42809
R8800 VDD.n2409 VDD.n2188 2.42809
R8801 VDD.n2409 VDD.n2190 2.42809
R8802 VDD.n2417 VDD.n2416 2.42809
R8803 VDD.n2417 VDD.n2182 2.42809
R8804 VDD.n2428 VDD.n2178 2.42809
R8805 VDD.n2429 VDD.n2428 2.42809
R8806 VDD.n2437 VDD.n2436 2.42809
R8807 VDD.n2436 VDD.n2175 2.42809
R8808 VDD.n2547 VDD.n2546 2.42809
R8809 VDD.n2547 VDD.n2117 2.42809
R8810 VDD.n2558 VDD.n2112 2.42809
R8811 VDD.n2559 VDD.n2558 2.42809
R8812 VDD.n2566 VDD.n2565 2.42809
R8813 VDD.n2565 VDD.n2106 2.42809
R8814 VDD.n2578 VDD.n2102 2.42809
R8815 VDD.n2578 VDD.n2104 2.42809
R8816 VDD.n2585 VDD.n2584 2.42809
R8817 VDD.n2585 VDD.n2097 2.42809
R8818 VDD.n2596 VDD.n2092 2.42809
R8819 VDD.n2597 VDD.n2596 2.42809
R8820 VDD.n2602 VDD.n2601 2.42809
R8821 VDD.n2601 VDD.n2084 2.42809
R8822 VDD.n2085 VDD.n2082 2.42809
R8823 VDD.n2615 VDD.n2082 2.42809
R8824 VDD.n2623 VDD.n2078 2.42809
R8825 VDD.n2623 VDD.n2076 2.42809
R8826 VDD.n3266 VDD.n3172 2.2074
R8827 VDD.n3356 VDD.n3112 2.2074
R8828 VDD.n893 VDD.n892 2.2074
R8829 VDD.n750 VDD.n749 2.2074
R8830 VDD.n615 VDD.n614 2.2074
R8831 VDD.n482 VDD.n481 2.2074
R8832 VDD.n339 VDD.n338 2.2074
R8833 VDD.n64 VDD.n63 2.2074
R8834 VDD.n204 VDD.n203 2.2074
R8835 VDD.n1310 VDD.n1278 2.19751
R8836 VDD.n1387 VDD.n1236 2.19751
R8837 VDD.n1464 VDD.n1194 2.19751
R8838 VDD.n1541 VDD.n1152 2.19751
R8839 VDD.n1618 VDD.n1110 2.19751
R8840 VDD.n1695 VDD.n1068 2.19751
R8841 VDD.n1769 VDD.n1025 2.19751
R8842 VDD.n114 VDD.n111 2.19751
R8843 VDD.n800 VDD.n797 2.19751
R8844 VDD.n665 VDD.n662 2.19751
R8845 VDD.n532 VDD.n529 2.19751
R8846 VDD.n389 VDD.n386 2.19751
R8847 VDD.n254 VDD.n251 2.19751
R8848 VDD.n3302 VDD 2.05519
R8849 VDD.n877 VDD.n875 2.02155
R8850 VDD.n734 VDD.n732 2.02155
R8851 VDD.n599 VDD.n597 2.02155
R8852 VDD.n466 VDD.n464 2.02155
R8853 VDD.n323 VDD.n321 2.02155
R8854 VDD.n48 VDD.n46 2.02155
R8855 VDD.n188 VDD.n186 2.02155
R8856 VDD.n1793 VDD.n1012 1.98671
R8857 VDD.n1718 VDD.n1054 1.98671
R8858 VDD.n1641 VDD.n1096 1.98671
R8859 VDD.n1564 VDD.n1138 1.98671
R8860 VDD.n1487 VDD.n1180 1.98671
R8861 VDD.n1410 VDD.n1222 1.98671
R8862 VDD.n1333 VDD.n1264 1.98671
R8863 VDD.n904 VDD.n901 1.98671
R8864 VDD.n761 VDD.n758 1.98671
R8865 VDD.n626 VDD.n623 1.98671
R8866 VDD.n493 VDD.n490 1.98671
R8867 VDD.n350 VDD.n347 1.98671
R8868 VDD.n75 VDD.n72 1.98671
R8869 VDD.n215 VDD.n212 1.98671
R8870 VDD.n199 VDD 1.91393
R8871 VDD.n59 VDD 1.91393
R8872 VDD.n334 VDD 1.91393
R8873 VDD.n477 VDD 1.91393
R8874 VDD.n610 VDD 1.91393
R8875 VDD.n745 VDD 1.91393
R8876 VDD.n888 VDD 1.91393
R8877 VDD.n2979 VDD.n1891 1.76602
R8878 VDD.n3050 VDD.n1849 1.76602
R8879 VDD.n195 VDD.n194 1.75668
R8880 VDD.n55 VDD.n54 1.75668
R8881 VDD.n330 VDD.n329 1.75668
R8882 VDD.n473 VDD.n472 1.75668
R8883 VDD.n606 VDD.n605 1.75668
R8884 VDD.n741 VDD.n740 1.75668
R8885 VDD.n884 VDD.n883 1.75668
R8886 VDD.n125 VDD.n118 1.62438
R8887 VDD.n137 VDD.n132 1.62438
R8888 VDD.n811 VDD.n804 1.62438
R8889 VDD.n549 VDD.n542 1.62438
R8890 VDD.n400 VDD.n393 1.62438
R8891 VDD.n264 VDD.n259 1.62438
R8892 VDD.n3283 VDD.n3166 1.57241
R8893 VDD.n3156 VDD.n3155 1.57241
R8894 VDD.n3373 VDD.n3106 1.57241
R8895 VDD.n3096 VDD.n3095 1.57241
R8896 VDD.n996 VDD.n995 1.57241
R8897 VDD.n1743 VDD.n1742 1.57241
R8898 VDD.n1666 VDD.n1078 1.57241
R8899 VDD.n1589 VDD.n1120 1.57241
R8900 VDD.n1512 VDD.n1162 1.57241
R8901 VDD.n1435 VDD.n1204 1.57241
R8902 VDD.n1358 VDD.n1246 1.57241
R8903 VDD.n163 VDD.n162 1.57241
R8904 VDD.n23 VDD.n22 1.57241
R8905 VDD.n852 VDD.n851 1.57241
R8906 VDD.n709 VDD.n708 1.57241
R8907 VDD.n574 VDD.n573 1.57241
R8908 VDD.n441 VDD.n440 1.57241
R8909 VDD.n298 VDD.n297 1.57241
R8910 VDD.n893 VDD.n891 1.54533
R8911 VDD.n750 VDD.n748 1.54533
R8912 VDD.n615 VDD.n613 1.54533
R8913 VDD.n482 VDD.n480 1.54533
R8914 VDD.n339 VDD.n337 1.54533
R8915 VDD.n64 VDD.n62 1.54533
R8916 VDD.n204 VDD.n202 1.54533
R8917 VDD.n1298 VDD.n1297 1.52886
R8918 VDD.n1375 VDD.n1374 1.52886
R8919 VDD.n1452 VDD.n1451 1.52886
R8920 VDD.n1529 VDD.n1528 1.52886
R8921 VDD.n1606 VDD.n1605 1.52886
R8922 VDD.n1683 VDD.n1682 1.52886
R8923 VDD.n1764 VDD.n1763 1.52886
R8924 VDD.n117 VDD.n116 1.52886
R8925 VDD.n803 VDD.n802 1.52886
R8926 VDD.n827 VDD.n826 1.52886
R8927 VDD.n676 VDD.n675 1.52886
R8928 VDD.n392 VDD.n391 1.52886
R8929 VDD.n408 VDD.n407 1.52886
R8930 VDD.n265 VDD.n258 1.52886
R8931 VDD.n965 VDD.n964 1.51754
R8932 VDD.n1814 VDD.n1000 1.47868
R8933 VDD.n1736 VDD.n1041 1.47868
R8934 VDD.n1082 VDD.n1081 1.47868
R8935 VDD.n1124 VDD.n1123 1.47868
R8936 VDD.n1166 VDD.n1165 1.47868
R8937 VDD.n1208 VDD.n1207 1.47868
R8938 VDD.n1250 VDD.n1249 1.47868
R8939 VDD.n172 VDD.n171 1.47868
R8940 VDD.n32 VDD.n31 1.47868
R8941 VDD.n861 VDD.n860 1.47868
R8942 VDD.n718 VDD.n717 1.47868
R8943 VDD.n583 VDD.n582 1.47868
R8944 VDD.n450 VDD.n449 1.47868
R8945 VDD.n307 VDD.n306 1.47868
R8946 VDD.n1803 VDD.n1005 1.39551
R8947 VDD.n1778 VDD.n1777 1.39551
R8948 VDD.n1046 VDD.n1045 1.39551
R8949 VDD.n1701 VDD.n1064 1.39551
R8950 VDD.n1089 VDD.n1088 1.39551
R8951 VDD.n1624 VDD.n1106 1.39551
R8952 VDD.n1131 VDD.n1130 1.39551
R8953 VDD.n1547 VDD.n1148 1.39551
R8954 VDD.n1173 VDD.n1172 1.39551
R8955 VDD.n1470 VDD.n1190 1.39551
R8956 VDD.n1215 VDD.n1214 1.39551
R8957 VDD.n1393 VDD.n1232 1.39551
R8958 VDD.n1257 VDD.n1256 1.39551
R8959 VDD.n1316 VDD.n1274 1.39551
R8960 VDD.n241 VDD.n240 1.39551
R8961 VDD.n101 VDD.n100 1.39551
R8962 VDD.n930 VDD.n929 1.39551
R8963 VDD.n787 VDD.n786 1.39551
R8964 VDD.n652 VDD.n651 1.39551
R8965 VDD.n519 VDD.n518 1.39551
R8966 VDD.n376 VDD.n375 1.39551
R8967 VDD.n957 VDD.n956 1.32791
R8968 VDD.n3173 VDD.n3167 1.32464
R8969 VDD.n3113 VDD.n3107 1.32464
R8970 VDD.n2362 VDD.n2218 1.32464
R8971 VDD.n2369 VDD.n2214 1.32464
R8972 VDD.n2368 VDD.n2208 1.32464
R8973 VDD.n2212 VDD.n2211 1.32464
R8974 VDD.n2380 VDD.n2204 1.32464
R8975 VDD.n2385 VDD.n2202 1.32464
R8976 VDD.n2386 VDD.n2198 1.32464
R8977 VDD.n2394 VDD.n2393 1.32464
R8978 VDD.n2398 VDD.n2196 1.32464
R8979 VDD.n2405 VDD.n2192 1.32464
R8980 VDD.n2404 VDD.n2188 1.32464
R8981 VDD.n2190 VDD.n2189 1.32464
R8982 VDD.n2416 VDD.n2184 1.32464
R8983 VDD.n2421 VDD.n2182 1.32464
R8984 VDD.n2422 VDD.n2178 1.32464
R8985 VDD.n2437 VDD.n2174 1.32464
R8986 VDD.n2175 VDD.n2171 1.32464
R8987 VDD.n2546 VDD.n2118 1.32464
R8988 VDD.n2551 VDD.n2117 1.32464
R8989 VDD.n2552 VDD.n2112 1.32464
R8990 VDD.n2562 VDD.n2559 1.32464
R8991 VDD.n2566 VDD.n2110 1.32464
R8992 VDD.n2574 VDD.n2106 1.32464
R8993 VDD.n2573 VDD.n2102 1.32464
R8994 VDD.n2104 VDD.n2103 1.32464
R8995 VDD.n2584 VDD.n2099 1.32464
R8996 VDD.n2589 VDD.n2097 1.32464
R8997 VDD.n2590 VDD.n2092 1.32464
R8998 VDD.n2598 VDD.n2597 1.32464
R8999 VDD.n2602 VDD.n2090 1.32464
R9000 VDD.n2611 VDD.n2084 1.32464
R9001 VDD.n2610 VDD.n2085 1.32464
R9002 VDD.n2618 VDD.n2078 1.32464
R9003 VDD.n2627 VDD.n2076 1.32464
R9004 VDD.n2736 VDD.n2735 1.32464
R9005 VDD.n2872 VDD.n2871 1.32464
R9006 VDD.n1289 VDD.n1285 1.32464
R9007 VDD.n1366 VDD.n1243 1.32464
R9008 VDD.n1443 VDD.n1201 1.32464
R9009 VDD.n1520 VDD.n1159 1.32464
R9010 VDD.n1597 VDD.n1117 1.32464
R9011 VDD.n1674 VDD.n1075 1.32464
R9012 VDD.n1035 VDD.n1030 1.32464
R9013 VDD.n153 VDD.n150 1.32464
R9014 VDD.n842 VDD.n839 1.32464
R9015 VDD.n699 VDD.n696 1.32464
R9016 VDD.n564 VDD.n561 1.32464
R9017 VDD.n431 VDD.n428 1.32464
R9018 VDD.n287 VDD.n284 1.32464
R9019 VDD.n988 VDD.n985 1.30219
R9020 VDD.n817 VDD.n815 1.24229
R9021 VDD.n948 VDD.n947 1.23309
R9022 VDD.n944 VDD.n943 1.17153
R9023 VDD.n540 VDD.n538 1.14677
R9024 VDD.n3290 VDD.n3161 1.10395
R9025 VDD.n3380 VDD.n3101 1.10395
R9026 VDD.n131 VDD.n129 1.05125
R9027 VDD.n674 VDD.n672 1.05125
R9028 VDD.n406 VDD.n404 1.05125
R9029 VDD.n963 VDD.n961 0.948648
R9030 VDD.n2431 VDD.n2430 0.883259
R9031 VDD.n2617 VDD.n2616 0.883259
R9032 VDD VDD.n2022 0.849458
R9033 VDD VDD.n1955 0.849458
R9034 VDD VDD.n1879 0.849458
R9035 VDD VDD.n1837 0.849458
R9036 VDD VDD.n1922 0.846854
R9037 VDD.n3392 VDD 0.838032
R9038 VDD.n2360 VDD 0.835135
R9039 VDD.n2548 VDD 0.832531
R9040 VDD.n199 VDD.n198 0.750619
R9041 VDD.n59 VDD.n58 0.750619
R9042 VDD.n334 VDD.n333 0.750619
R9043 VDD.n477 VDD.n476 0.750619
R9044 VDD.n610 VDD.n609 0.750619
R9045 VDD.n745 VDD.n744 0.750619
R9046 VDD.n888 VDD.n887 0.750619
R9047 VDD.n257 VDD 0.678885
R9048 VDD.n268 VDD 0.546892
R9049 VDD.n1295 VDD.n1282 0.478112
R9050 VDD.n1372 VDD.n1240 0.478112
R9051 VDD.n1449 VDD.n1198 0.478112
R9052 VDD.n1526 VDD.n1156 0.478112
R9053 VDD.n1603 VDD.n1114 0.478112
R9054 VDD.n1680 VDD.n1072 0.478112
R9055 VDD.n1761 VDD.n1759 0.478112
R9056 VDD.n138 VDD.n131 0.478112
R9057 VDD.n684 VDD.n674 0.478112
R9058 VDD.n416 VDD.n406 0.478112
R9059 VDD.n273 VDD.n270 0.478112
R9060 VDD.n973 VDD.n963 0.474574
R9061 VDD.n3242 VDD.n3192 0.441879
R9062 VDD.n3332 VDD.n3132 0.441879
R9063 VDD.n2430 VDD.n2429 0.441879
R9064 VDD.n2445 VDD.n2170 0.441879
R9065 VDD.n2455 VDD.n2166 0.441879
R9066 VDD.n2457 VDD.n2456 0.441879
R9067 VDD.n2463 VDD.n2462 0.441879
R9068 VDD.n2461 VDD.n2159 0.441879
R9069 VDD.n2474 VDD.n2156 0.441879
R9070 VDD.n2473 VDD.n2157 0.441879
R9071 VDD.n2481 VDD.n2480 0.441879
R9072 VDD.n2482 VDD.n2150 0.441879
R9073 VDD.n2492 VDD.n2146 0.441879
R9074 VDD.n2494 VDD.n2493 0.441879
R9075 VDD.n2500 VDD.n2499 0.441879
R9076 VDD.n2498 VDD.n2140 0.441879
R9077 VDD.n2512 VDD.n2136 0.441879
R9078 VDD.n2510 VDD.n2138 0.441879
R9079 VDD.n2519 VDD.n2518 0.441879
R9080 VDD.n2520 VDD.n2130 0.441879
R9081 VDD.n2530 VDD.n2126 0.441879
R9082 VDD.n2616 VDD.n2615 0.441879
R9083 VDD.n2642 VDD.n2641 0.441879
R9084 VDD.n2756 VDD.n2015 0.441879
R9085 VDD.n2778 VDD.n2777 0.441879
R9086 VDD.n2892 VDD.n2891 0.441879
R9087 VDD.n1943 VDD.n1937 0.441879
R9088 VDD.n1915 VDD.n1908 0.441879
R9089 VDD.n2958 VDD.n2957 0.441879
R9090 VDD.n1872 VDD.n1866 0.441879
R9091 VDD.n3029 VDD.n3028 0.441879
R9092 VDD.n1830 VDD.n1826 0.441879
R9093 VDD.n541 VDD.n540 0.38259
R9094 VDD.n955 VDD.n948 0.379759
R9095 VDD.n3392 VDD 0.344795
R9096 VDD.n3393 VDD 0.344795
R9097 VDD VDD.n3394 0.344795
R9098 VDD.n62 VDD.n61 0.332294
R9099 VDD.n891 VDD.n890 0.331593
R9100 VDD.n748 VDD.n747 0.331593
R9101 VDD.n613 VDD.n612 0.331593
R9102 VDD.n480 VDD.n479 0.331593
R9103 VDD.n337 VDD.n336 0.331593
R9104 VDD.n202 VDD.n201 0.331593
R9105 VDD.n818 VDD.n817 0.287067
R9106 VDD.n957 VDD.n955 0.284944
R9107 VDD.n197 VDD 0.259429
R9108 VDD.n57 VDD 0.259429
R9109 VDD.n332 VDD 0.259429
R9110 VDD.n475 VDD 0.259429
R9111 VDD.n608 VDD 0.259429
R9112 VDD.n743 VDD 0.259429
R9113 VDD.n886 VDD 0.259429
R9114 VDD.n2902 VDD 0.232271
R9115 VDD.n2446 VDD 0.229667
R9116 VDD.n2955 VDD 0.229667
R9117 VDD.n3026 VDD 0.229667
R9118 VDD.n1683 VDD.n1681 0.226033
R9119 VDD.n1606 VDD.n1604 0.226033
R9120 VDD.n1375 VDD.n1373 0.226033
R9121 VDD.n1298 VDD.n1296 0.226033
R9122 VDD.n1763 VDD.n1762 0.225256
R9123 VDD.n1529 VDD.n1527 0.225256
R9124 VDD.n1452 VDD.n1450 0.225256
R9125 VDD.n3277 VDD.n3168 0.22119
R9126 VDD.n3367 VDD.n3108 0.22119
R9127 VDD.n2264 VDD.n2256 0.22119
R9128 VDD.n2263 VDD.n2262 0.22119
R9129 VDD.n2262 VDD.n2258 0.22119
R9130 VDD.n2272 VDD.n2271 0.22119
R9131 VDD.n2273 VDD.n2250 0.22119
R9132 VDD.n2283 VDD.n2247 0.22119
R9133 VDD.n2285 VDD.n2284 0.22119
R9134 VDD.n2291 VDD.n2290 0.22119
R9135 VDD.n2289 VDD.n2241 0.22119
R9136 VDD.n2302 VDD.n2238 0.22119
R9137 VDD.n2301 VDD.n2239 0.22119
R9138 VDD.n2310 VDD.n2309 0.22119
R9139 VDD.n2311 VDD.n2232 0.22119
R9140 VDD.n2321 VDD.n2229 0.22119
R9141 VDD.n2324 VDD.n2323 0.22119
R9142 VDD.n2330 VDD.n2329 0.22119
R9143 VDD.n2328 VDD.n2220 0.22119
R9144 VDD.n2352 VDD.n2221 0.22119
R9145 VDD.n2633 VDD.n2075 0.22119
R9146 VDD.n2633 VDD.n2071 0.22119
R9147 VDD.n2642 VDD.n2068 0.22119
R9148 VDD.n2648 VDD.n2068 0.22119
R9149 VDD.n2654 VDD.n2064 0.22119
R9150 VDD.n2654 VDD.n2061 0.22119
R9151 VDD.n2062 VDD.n2057 0.22119
R9152 VDD.n2665 VDD.n2057 0.22119
R9153 VDD.n2671 VDD.n2055 0.22119
R9154 VDD.n2671 VDD.n2051 0.22119
R9155 VDD.n2679 VDD.n2049 0.22119
R9156 VDD.n2685 VDD.n2049 0.22119
R9157 VDD.n2691 VDD.n2045 0.22119
R9158 VDD.n2691 VDD.n2041 0.22119
R9159 VDD.n2043 VDD.n2037 0.22119
R9160 VDD.n2703 VDD.n2037 0.22119
R9161 VDD.n2709 VDD.n2035 0.22119
R9162 VDD.n2709 VDD.n2031 0.22119
R9163 VDD.n2769 VDD.n2008 0.22119
R9164 VDD.n2769 VDD.n2004 0.22119
R9165 VDD.n2778 VDD.n2001 0.22119
R9166 VDD.n2784 VDD.n2001 0.22119
R9167 VDD.n2790 VDD.n1997 0.22119
R9168 VDD.n2790 VDD.n1994 0.22119
R9169 VDD.n1995 VDD.n1990 0.22119
R9170 VDD.n2801 VDD.n1990 0.22119
R9171 VDD.n2807 VDD.n1988 0.22119
R9172 VDD.n2807 VDD.n1984 0.22119
R9173 VDD.n2815 VDD.n1982 0.22119
R9174 VDD.n2821 VDD.n1982 0.22119
R9175 VDD.n2827 VDD.n1978 0.22119
R9176 VDD.n2827 VDD.n1974 0.22119
R9177 VDD.n1976 VDD.n1970 0.22119
R9178 VDD.n2839 VDD.n1970 0.22119
R9179 VDD.n2845 VDD.n1968 0.22119
R9180 VDD.n2845 VDD.n1964 0.22119
R9181 VDD.n3393 VDD.n3392 0.215674
R9182 VDD.n3394 VDD.n3393 0.21443
R9183 VDD.n2630 VDD 0.208833
R9184 VDD.n2766 VDD 0.208833
R9185 VDD.n973 VDD.n972 0.19013
R9186 VDD.n3394 VDD 0.151308
R9187 VDD.n3219 VDD.n3207 0.120292
R9188 VDD.n3220 VDD.n3219 0.120292
R9189 VDD.n3221 VDD.n3220 0.120292
R9190 VDD.n3221 VDD.n3198 0.120292
R9191 VDD.n3230 VDD.n3198 0.120292
R9192 VDD.n3231 VDD.n3230 0.120292
R9193 VDD.n3234 VDD.n3231 0.120292
R9194 VDD.n3234 VDD.n3233 0.120292
R9195 VDD.n3233 VDD.n3190 0.120292
R9196 VDD.n3244 VDD.n3190 0.120292
R9197 VDD.n3246 VDD.n3244 0.120292
R9198 VDD.n3246 VDD.n3245 0.120292
R9199 VDD.n3245 VDD.n3182 0.120292
R9200 VDD.n3255 VDD.n3182 0.120292
R9201 VDD.n3257 VDD.n3255 0.120292
R9202 VDD.n3257 VDD.n3256 0.120292
R9203 VDD.n3256 VDD.n3174 0.120292
R9204 VDD.n3267 VDD.n3174 0.120292
R9205 VDD.n3269 VDD.n3267 0.120292
R9206 VDD.n3269 VDD.n3268 0.120292
R9207 VDD.n3279 VDD.n3278 0.120292
R9208 VDD.n3280 VDD.n3279 0.120292
R9209 VDD.n3281 VDD.n3280 0.120292
R9210 VDD.n3281 VDD.n3159 0.120292
R9211 VDD.n3292 VDD.n3159 0.120292
R9212 VDD.n3293 VDD.n3153 0.120292
R9213 VDD.n3301 VDD.n3153 0.120292
R9214 VDD.n3302 VDD.n3147 0.120292
R9215 VDD.n3309 VDD.n3147 0.120292
R9216 VDD.n3310 VDD.n3309 0.120292
R9217 VDD.n3311 VDD.n3310 0.120292
R9218 VDD.n3311 VDD.n3138 0.120292
R9219 VDD.n3320 VDD.n3138 0.120292
R9220 VDD.n3321 VDD.n3320 0.120292
R9221 VDD.n3324 VDD.n3321 0.120292
R9222 VDD.n3324 VDD.n3323 0.120292
R9223 VDD.n3323 VDD.n3130 0.120292
R9224 VDD.n3334 VDD.n3130 0.120292
R9225 VDD.n3336 VDD.n3334 0.120292
R9226 VDD.n3336 VDD.n3335 0.120292
R9227 VDD.n3335 VDD.n3122 0.120292
R9228 VDD.n3345 VDD.n3122 0.120292
R9229 VDD.n3347 VDD.n3345 0.120292
R9230 VDD.n3347 VDD.n3346 0.120292
R9231 VDD.n3346 VDD.n3114 0.120292
R9232 VDD.n3357 VDD.n3114 0.120292
R9233 VDD.n3359 VDD.n3357 0.120292
R9234 VDD.n3359 VDD.n3358 0.120292
R9235 VDD.n3369 VDD.n3368 0.120292
R9236 VDD.n3370 VDD.n3369 0.120292
R9237 VDD.n3371 VDD.n3370 0.120292
R9238 VDD.n3371 VDD.n3099 0.120292
R9239 VDD.n3382 VDD.n3099 0.120292
R9240 VDD.n3383 VDD.n3093 0.120292
R9241 VDD.n3391 VDD.n3093 0.120292
R9242 VDD.n2738 VDD.n2022 0.120292
R9243 VDD.n2739 VDD.n2738 0.120292
R9244 VDD.n2740 VDD.n2739 0.120292
R9245 VDD.n2740 VDD.n2016 0.120292
R9246 VDD.n2752 VDD.n2016 0.120292
R9247 VDD.n2753 VDD.n2752 0.120292
R9248 VDD.n2755 VDD.n2753 0.120292
R9249 VDD.n2755 VDD.n2754 0.120292
R9250 VDD.n2874 VDD.n1955 0.120292
R9251 VDD.n2875 VDD.n2874 0.120292
R9252 VDD.n2876 VDD.n2875 0.120292
R9253 VDD.n2876 VDD.n1949 0.120292
R9254 VDD.n2887 VDD.n1949 0.120292
R9255 VDD.n2888 VDD.n2887 0.120292
R9256 VDD.n2888 VDD.n1944 0.120292
R9257 VDD.n2901 VDD.n1944 0.120292
R9258 VDD.n2910 VDD.n1936 0.120292
R9259 VDD.n2911 VDD.n2910 0.120292
R9260 VDD.n2912 VDD.n2911 0.120292
R9261 VDD.n2912 VDD.n1928 0.120292
R9262 VDD.n2920 VDD.n1928 0.120292
R9263 VDD.n2921 VDD.n2920 0.120292
R9264 VDD.n2922 VDD.n2921 0.120292
R9265 VDD.n2932 VDD.n1922 0.120292
R9266 VDD.n2933 VDD.n2932 0.120292
R9267 VDD.n2933 VDD.n1916 0.120292
R9268 VDD.n2942 VDD.n1916 0.120292
R9269 VDD.n2943 VDD.n2942 0.120292
R9270 VDD.n2944 VDD.n2943 0.120292
R9271 VDD.n2944 VDD.n1906 0.120292
R9272 VDD.n2954 VDD.n1906 0.120292
R9273 VDD.n2956 VDD.n1899 0.120292
R9274 VDD.n2968 VDD.n1899 0.120292
R9275 VDD.n2969 VDD.n2968 0.120292
R9276 VDD.n2970 VDD.n2969 0.120292
R9277 VDD.n2970 VDD.n1889 0.120292
R9278 VDD.n2981 VDD.n1889 0.120292
R9279 VDD.n2982 VDD.n2981 0.120292
R9280 VDD.n3002 VDD.n1879 0.120292
R9281 VDD.n3003 VDD.n3002 0.120292
R9282 VDD.n3003 VDD.n1873 0.120292
R9283 VDD.n3012 VDD.n1873 0.120292
R9284 VDD.n3013 VDD.n3012 0.120292
R9285 VDD.n3014 VDD.n3013 0.120292
R9286 VDD.n3014 VDD.n1864 0.120292
R9287 VDD.n3025 VDD.n1864 0.120292
R9288 VDD.n3027 VDD.n1857 0.120292
R9289 VDD.n3039 VDD.n1857 0.120292
R9290 VDD.n3040 VDD.n3039 0.120292
R9291 VDD.n3041 VDD.n3040 0.120292
R9292 VDD.n3041 VDD.n1847 0.120292
R9293 VDD.n3052 VDD.n1847 0.120292
R9294 VDD.n3053 VDD.n3052 0.120292
R9295 VDD.n3073 VDD.n1837 0.120292
R9296 VDD.n3074 VDD.n3073 0.120292
R9297 VDD.n3074 VDD.n1831 0.120292
R9298 VDD.n3083 VDD.n1831 0.120292
R9299 VDD.n3084 VDD.n3083 0.120292
R9300 VDD.n3085 VDD.n3084 0.120292
R9301 VDD.n3085 VDD.n1824 0.120292
R9302 VDD.n3092 VDD.n1824 0.120292
R9303 VDD.n1291 VDD.n1290 0.120292
R9304 VDD.n1301 VDD.n1291 0.120292
R9305 VDD.n1301 VDD.n1300 0.120292
R9306 VDD.n1312 VDD.n1311 0.120292
R9307 VDD.n1314 VDD.n1312 0.120292
R9308 VDD.n1314 VDD.n1313 0.120292
R9309 VDD.n1313 VDD.n1269 0.120292
R9310 VDD.n1324 VDD.n1269 0.120292
R9311 VDD.n1325 VDD.n1324 0.120292
R9312 VDD.n1326 VDD.n1325 0.120292
R9313 VDD.n1326 VDD.n1262 0.120292
R9314 VDD.n1334 VDD.n1262 0.120292
R9315 VDD.n1335 VDD.n1334 0.120292
R9316 VDD.n1336 VDD.n1335 0.120292
R9317 VDD.n1336 VDD.n1254 0.120292
R9318 VDD.n1345 VDD.n1254 0.120292
R9319 VDD.n1346 VDD.n1345 0.120292
R9320 VDD.n1347 VDD.n1346 0.120292
R9321 VDD.n1347 VDD.n1248 0.120292
R9322 VDD.n1356 VDD.n1248 0.120292
R9323 VDD.n1359 VDD.n1356 0.120292
R9324 VDD.n1360 VDD.n1359 0.120292
R9325 VDD.n1367 VDD.n1241 0.120292
R9326 VDD.n1368 VDD.n1367 0.120292
R9327 VDD.n1378 VDD.n1368 0.120292
R9328 VDD.n1378 VDD.n1377 0.120292
R9329 VDD.n1389 VDD.n1388 0.120292
R9330 VDD.n1391 VDD.n1389 0.120292
R9331 VDD.n1391 VDD.n1390 0.120292
R9332 VDD.n1390 VDD.n1227 0.120292
R9333 VDD.n1401 VDD.n1227 0.120292
R9334 VDD.n1402 VDD.n1401 0.120292
R9335 VDD.n1403 VDD.n1402 0.120292
R9336 VDD.n1403 VDD.n1220 0.120292
R9337 VDD.n1411 VDD.n1220 0.120292
R9338 VDD.n1412 VDD.n1411 0.120292
R9339 VDD.n1413 VDD.n1412 0.120292
R9340 VDD.n1413 VDD.n1212 0.120292
R9341 VDD.n1422 VDD.n1212 0.120292
R9342 VDD.n1423 VDD.n1422 0.120292
R9343 VDD.n1424 VDD.n1423 0.120292
R9344 VDD.n1424 VDD.n1206 0.120292
R9345 VDD.n1433 VDD.n1206 0.120292
R9346 VDD.n1436 VDD.n1433 0.120292
R9347 VDD.n1437 VDD.n1436 0.120292
R9348 VDD.n1444 VDD.n1199 0.120292
R9349 VDD.n1445 VDD.n1444 0.120292
R9350 VDD.n1455 VDD.n1445 0.120292
R9351 VDD.n1455 VDD.n1454 0.120292
R9352 VDD.n1466 VDD.n1465 0.120292
R9353 VDD.n1468 VDD.n1466 0.120292
R9354 VDD.n1468 VDD.n1467 0.120292
R9355 VDD.n1467 VDD.n1185 0.120292
R9356 VDD.n1478 VDD.n1185 0.120292
R9357 VDD.n1479 VDD.n1478 0.120292
R9358 VDD.n1480 VDD.n1479 0.120292
R9359 VDD.n1480 VDD.n1178 0.120292
R9360 VDD.n1488 VDD.n1178 0.120292
R9361 VDD.n1489 VDD.n1488 0.120292
R9362 VDD.n1490 VDD.n1489 0.120292
R9363 VDD.n1490 VDD.n1170 0.120292
R9364 VDD.n1499 VDD.n1170 0.120292
R9365 VDD.n1500 VDD.n1499 0.120292
R9366 VDD.n1501 VDD.n1500 0.120292
R9367 VDD.n1501 VDD.n1164 0.120292
R9368 VDD.n1510 VDD.n1164 0.120292
R9369 VDD.n1513 VDD.n1510 0.120292
R9370 VDD.n1514 VDD.n1513 0.120292
R9371 VDD.n1521 VDD.n1157 0.120292
R9372 VDD.n1522 VDD.n1521 0.120292
R9373 VDD.n1532 VDD.n1522 0.120292
R9374 VDD.n1532 VDD.n1531 0.120292
R9375 VDD.n1543 VDD.n1542 0.120292
R9376 VDD.n1545 VDD.n1543 0.120292
R9377 VDD.n1545 VDD.n1544 0.120292
R9378 VDD.n1544 VDD.n1143 0.120292
R9379 VDD.n1555 VDD.n1143 0.120292
R9380 VDD.n1556 VDD.n1555 0.120292
R9381 VDD.n1557 VDD.n1556 0.120292
R9382 VDD.n1557 VDD.n1136 0.120292
R9383 VDD.n1565 VDD.n1136 0.120292
R9384 VDD.n1566 VDD.n1565 0.120292
R9385 VDD.n1567 VDD.n1566 0.120292
R9386 VDD.n1567 VDD.n1128 0.120292
R9387 VDD.n1576 VDD.n1128 0.120292
R9388 VDD.n1577 VDD.n1576 0.120292
R9389 VDD.n1578 VDD.n1577 0.120292
R9390 VDD.n1578 VDD.n1122 0.120292
R9391 VDD.n1587 VDD.n1122 0.120292
R9392 VDD.n1590 VDD.n1587 0.120292
R9393 VDD.n1591 VDD.n1590 0.120292
R9394 VDD.n1598 VDD.n1115 0.120292
R9395 VDD.n1599 VDD.n1598 0.120292
R9396 VDD.n1609 VDD.n1599 0.120292
R9397 VDD.n1609 VDD.n1608 0.120292
R9398 VDD.n1620 VDD.n1619 0.120292
R9399 VDD.n1622 VDD.n1620 0.120292
R9400 VDD.n1622 VDD.n1621 0.120292
R9401 VDD.n1621 VDD.n1101 0.120292
R9402 VDD.n1632 VDD.n1101 0.120292
R9403 VDD.n1633 VDD.n1632 0.120292
R9404 VDD.n1634 VDD.n1633 0.120292
R9405 VDD.n1634 VDD.n1094 0.120292
R9406 VDD.n1642 VDD.n1094 0.120292
R9407 VDD.n1643 VDD.n1642 0.120292
R9408 VDD.n1644 VDD.n1643 0.120292
R9409 VDD.n1644 VDD.n1086 0.120292
R9410 VDD.n1653 VDD.n1086 0.120292
R9411 VDD.n1654 VDD.n1653 0.120292
R9412 VDD.n1655 VDD.n1654 0.120292
R9413 VDD.n1655 VDD.n1080 0.120292
R9414 VDD.n1664 VDD.n1080 0.120292
R9415 VDD.n1667 VDD.n1664 0.120292
R9416 VDD.n1668 VDD.n1667 0.120292
R9417 VDD.n1675 VDD.n1073 0.120292
R9418 VDD.n1676 VDD.n1675 0.120292
R9419 VDD.n1686 VDD.n1676 0.120292
R9420 VDD.n1686 VDD.n1685 0.120292
R9421 VDD.n1697 VDD.n1696 0.120292
R9422 VDD.n1699 VDD.n1697 0.120292
R9423 VDD.n1699 VDD.n1698 0.120292
R9424 VDD.n1698 VDD.n1059 0.120292
R9425 VDD.n1709 VDD.n1059 0.120292
R9426 VDD.n1710 VDD.n1709 0.120292
R9427 VDD.n1711 VDD.n1710 0.120292
R9428 VDD.n1711 VDD.n1052 0.120292
R9429 VDD.n1719 VDD.n1052 0.120292
R9430 VDD.n1720 VDD.n1719 0.120292
R9431 VDD.n1721 VDD.n1720 0.120292
R9432 VDD.n1721 VDD.n1043 0.120292
R9433 VDD.n1731 VDD.n1043 0.120292
R9434 VDD.n1732 VDD.n1731 0.120292
R9435 VDD.n1734 VDD.n1732 0.120292
R9436 VDD.n1734 VDD.n1733 0.120292
R9437 VDD.n1733 VDD.n1036 0.120292
R9438 VDD.n1744 VDD.n1036 0.120292
R9439 VDD.n1745 VDD.n1744 0.120292
R9440 VDD.n1746 VDD.n1029 0.120292
R9441 VDD.n1756 VDD.n1029 0.120292
R9442 VDD.n1757 VDD.n1756 0.120292
R9443 VDD.n1758 VDD.n1757 0.120292
R9444 VDD.n1768 VDD.n1767 0.120292
R9445 VDD.n1767 VDD.n1019 0.120292
R9446 VDD.n1779 VDD.n1019 0.120292
R9447 VDD.n1780 VDD.n1779 0.120292
R9448 VDD.n1782 VDD.n1780 0.120292
R9449 VDD.n1782 VDD.n1781 0.120292
R9450 VDD.n1781 VDD.n1013 0.120292
R9451 VDD.n1791 VDD.n1013 0.120292
R9452 VDD.n1792 VDD.n1791 0.120292
R9453 VDD.n1792 VDD.n1006 0.120292
R9454 VDD.n1801 VDD.n1006 0.120292
R9455 VDD.n1804 VDD.n1801 0.120292
R9456 VDD.n1805 VDD.n1804 0.120292
R9457 VDD.n1805 VDD.n1001 0.120292
R9458 VDD.n1813 VDD.n1001 0.120292
R9459 VDD.n1815 VDD.n1813 0.120292
R9460 VDD.n1816 VDD.n1815 0.120292
R9461 VDD.n1816 VDD.n993 0.120292
R9462 VDD.n1823 VDD.n993 0.120292
R9463 VDD.n28 VDD.n24 0.120292
R9464 VDD.n33 VDD.n28 0.120292
R9465 VDD.n37 VDD.n33 0.120292
R9466 VDD.n41 VDD.n37 0.120292
R9467 VDD.n45 VDD.n41 0.120292
R9468 VDD.n49 VDD.n45 0.120292
R9469 VDD.n76 VDD.n70 0.120292
R9470 VDD.n80 VDD.n76 0.120292
R9471 VDD.n84 VDD.n80 0.120292
R9472 VDD.n88 VDD.n84 0.120292
R9473 VDD.n92 VDD.n88 0.120292
R9474 VDD.n96 VDD.n92 0.120292
R9475 VDD.n102 VDD.n96 0.120292
R9476 VDD.n106 VDD.n102 0.120292
R9477 VDD.n110 VDD.n106 0.120292
R9478 VDD.n115 VDD.n110 0.120292
R9479 VDD.n126 VDD.n115 0.120292
R9480 VDD.n148 VDD.n144 0.120292
R9481 VDD.n154 VDD.n148 0.120292
R9482 VDD.n155 VDD.n154 0.120292
R9483 VDD.n168 VDD.n164 0.120292
R9484 VDD.n173 VDD.n168 0.120292
R9485 VDD.n177 VDD.n173 0.120292
R9486 VDD.n181 VDD.n177 0.120292
R9487 VDD.n185 VDD.n181 0.120292
R9488 VDD.n189 VDD.n185 0.120292
R9489 VDD.n216 VDD.n210 0.120292
R9490 VDD.n220 VDD.n216 0.120292
R9491 VDD.n224 VDD.n220 0.120292
R9492 VDD.n228 VDD.n224 0.120292
R9493 VDD.n232 VDD.n228 0.120292
R9494 VDD.n236 VDD.n232 0.120292
R9495 VDD.n242 VDD.n236 0.120292
R9496 VDD.n246 VDD.n242 0.120292
R9497 VDD.n250 VDD.n246 0.120292
R9498 VDD.n255 VDD.n250 0.120292
R9499 VDD.n278 VDD.n274 0.120292
R9500 VDD.n282 VDD.n278 0.120292
R9501 VDD.n288 VDD.n282 0.120292
R9502 VDD.n290 VDD.n288 0.120292
R9503 VDD.n303 VDD.n299 0.120292
R9504 VDD.n308 VDD.n303 0.120292
R9505 VDD.n312 VDD.n308 0.120292
R9506 VDD.n316 VDD.n312 0.120292
R9507 VDD.n320 VDD.n316 0.120292
R9508 VDD.n324 VDD.n320 0.120292
R9509 VDD.n351 VDD.n345 0.120292
R9510 VDD.n355 VDD.n351 0.120292
R9511 VDD.n359 VDD.n355 0.120292
R9512 VDD.n363 VDD.n359 0.120292
R9513 VDD.n367 VDD.n363 0.120292
R9514 VDD.n371 VDD.n367 0.120292
R9515 VDD.n377 VDD.n371 0.120292
R9516 VDD.n381 VDD.n377 0.120292
R9517 VDD.n385 VDD.n381 0.120292
R9518 VDD.n390 VDD.n385 0.120292
R9519 VDD.n401 VDD.n390 0.120292
R9520 VDD.n426 VDD.n422 0.120292
R9521 VDD.n432 VDD.n426 0.120292
R9522 VDD.n433 VDD.n432 0.120292
R9523 VDD.n446 VDD.n442 0.120292
R9524 VDD.n451 VDD.n446 0.120292
R9525 VDD.n455 VDD.n451 0.120292
R9526 VDD.n459 VDD.n455 0.120292
R9527 VDD.n463 VDD.n459 0.120292
R9528 VDD.n467 VDD.n463 0.120292
R9529 VDD.n494 VDD.n488 0.120292
R9530 VDD.n498 VDD.n494 0.120292
R9531 VDD.n502 VDD.n498 0.120292
R9532 VDD.n506 VDD.n502 0.120292
R9533 VDD.n510 VDD.n506 0.120292
R9534 VDD.n514 VDD.n510 0.120292
R9535 VDD.n520 VDD.n514 0.120292
R9536 VDD.n524 VDD.n520 0.120292
R9537 VDD.n528 VDD.n524 0.120292
R9538 VDD.n533 VDD.n528 0.120292
R9539 VDD.n537 VDD.n533 0.120292
R9540 VDD.n550 VDD.n537 0.120292
R9541 VDD.n559 VDD.n555 0.120292
R9542 VDD.n565 VDD.n559 0.120292
R9543 VDD.n566 VDD.n565 0.120292
R9544 VDD.n579 VDD.n575 0.120292
R9545 VDD.n584 VDD.n579 0.120292
R9546 VDD.n588 VDD.n584 0.120292
R9547 VDD.n592 VDD.n588 0.120292
R9548 VDD.n596 VDD.n592 0.120292
R9549 VDD.n600 VDD.n596 0.120292
R9550 VDD.n627 VDD.n621 0.120292
R9551 VDD.n631 VDD.n627 0.120292
R9552 VDD.n635 VDD.n631 0.120292
R9553 VDD.n639 VDD.n635 0.120292
R9554 VDD.n643 VDD.n639 0.120292
R9555 VDD.n647 VDD.n643 0.120292
R9556 VDD.n653 VDD.n647 0.120292
R9557 VDD.n657 VDD.n653 0.120292
R9558 VDD.n661 VDD.n657 0.120292
R9559 VDD.n666 VDD.n661 0.120292
R9560 VDD.n670 VDD.n666 0.120292
R9561 VDD.n694 VDD.n690 0.120292
R9562 VDD.n700 VDD.n694 0.120292
R9563 VDD.n701 VDD.n700 0.120292
R9564 VDD.n714 VDD.n710 0.120292
R9565 VDD.n719 VDD.n714 0.120292
R9566 VDD.n723 VDD.n719 0.120292
R9567 VDD.n727 VDD.n723 0.120292
R9568 VDD.n731 VDD.n727 0.120292
R9569 VDD.n735 VDD.n731 0.120292
R9570 VDD.n762 VDD.n756 0.120292
R9571 VDD.n766 VDD.n762 0.120292
R9572 VDD.n770 VDD.n766 0.120292
R9573 VDD.n774 VDD.n770 0.120292
R9574 VDD.n778 VDD.n774 0.120292
R9575 VDD.n782 VDD.n778 0.120292
R9576 VDD.n788 VDD.n782 0.120292
R9577 VDD.n792 VDD.n788 0.120292
R9578 VDD.n796 VDD.n792 0.120292
R9579 VDD.n801 VDD.n796 0.120292
R9580 VDD.n812 VDD.n801 0.120292
R9581 VDD.n837 VDD.n833 0.120292
R9582 VDD.n843 VDD.n837 0.120292
R9583 VDD.n844 VDD.n843 0.120292
R9584 VDD.n857 VDD.n853 0.120292
R9585 VDD.n862 VDD.n857 0.120292
R9586 VDD.n866 VDD.n862 0.120292
R9587 VDD.n870 VDD.n866 0.120292
R9588 VDD.n874 VDD.n870 0.120292
R9589 VDD.n878 VDD.n874 0.120292
R9590 VDD.n905 VDD.n899 0.120292
R9591 VDD.n909 VDD.n905 0.120292
R9592 VDD.n913 VDD.n909 0.120292
R9593 VDD.n917 VDD.n913 0.120292
R9594 VDD.n921 VDD.n917 0.120292
R9595 VDD.n925 VDD.n921 0.120292
R9596 VDD.n931 VDD.n925 0.120292
R9597 VDD.n935 VDD.n931 0.120292
R9598 VDD.n939 VDD.n935 0.120292
R9599 VDD.n945 VDD.n939 0.120292
R9600 VDD.n983 VDD.n979 0.120292
R9601 VDD.n989 VDD.n983 0.120292
R9602 VDD.n992 VDD.n989 0.120292
R9603 VDD.n1311 VDD.n1276 0.11899
R9604 VDD.n1388 VDD.n1234 0.11899
R9605 VDD.n1465 VDD.n1192 0.11899
R9606 VDD.n1542 VDD.n1150 0.11899
R9607 VDD.n1619 VDD.n1108 0.11899
R9608 VDD.n1696 VDD.n1066 0.11899
R9609 VDD.n1768 VDD.n1766 0.11899
R9610 VDD.n144 VDD.n140 0.11899
R9611 VDD.n422 VDD.n418 0.11899
R9612 VDD.n690 VDD.n686 0.11899
R9613 VDD.n979 VDD.n975 0.117688
R9614 VDD.n946 VDD.n945 0.116385
R9615 VDD.n50 VDD.n49 0.111177
R9616 VDD.n190 VDD.n189 0.111177
R9617 VDD.n325 VDD.n324 0.111177
R9618 VDD.n468 VDD.n467 0.111177
R9619 VDD.n601 VDD.n600 0.111177
R9620 VDD.n736 VDD.n735 0.111177
R9621 VDD.n879 VDD.n878 0.111177
R9622 VDD.n70 VDD.n66 0.107271
R9623 VDD.n210 VDD.n206 0.107271
R9624 VDD.n345 VDD.n341 0.107271
R9625 VDD.n488 VDD.n484 0.107271
R9626 VDD.n621 VDD.n617 0.107271
R9627 VDD.n756 VDD.n752 0.107271
R9628 VDD.n899 VDD.n895 0.107271
R9629 VDD.n268 VDD.n267 0.104881
R9630 VDD.n1300 VDD.n1299 0.0994583
R9631 VDD.n1377 VDD.n1376 0.0994583
R9632 VDD.n1454 VDD.n1453 0.0994583
R9633 VDD.n1531 VDD.n1530 0.0994583
R9634 VDD.n1608 VDD.n1607 0.0994583
R9635 VDD.n1685 VDD.n1684 0.0994583
R9636 VDD.n1758 VDD.n1026 0.0994583
R9637 VDD.n256 VDD.n255 0.0994583
R9638 VDD.n671 VDD.n670 0.0994583
R9639 VDD.n833 VDD.n829 0.0994583
R9640 VDD.n2274 VDD.n2251 0.0981562
R9641 VDD.n2276 VDD.n2246 0.0981562
R9642 VDD.n2288 VDD.n2287 0.0981562
R9643 VDD.n2300 VDD.n2298 0.0981562
R9644 VDD.n2312 VDD.n2233 0.0981562
R9645 VDD.n2314 VDD.n2227 0.0981562
R9646 VDD.n2327 VDD.n2326 0.0981562
R9647 VDD.n2372 VDD.n2370 0.0981562
R9648 VDD.n2382 VDD.n2203 0.0981562
R9649 VDD.n2384 VDD.n2199 0.0981562
R9650 VDD.n2396 VDD.n2395 0.0981562
R9651 VDD.n2408 VDD.n2406 0.0981562
R9652 VDD.n2418 VDD.n2183 0.0981562
R9653 VDD.n2420 VDD.n2179 0.0981562
R9654 VDD.n2435 VDD.n2432 0.0981562
R9655 VDD.n2460 VDD.n2459 0.0981562
R9656 VDD.n2472 VDD.n2470 0.0981562
R9657 VDD.n2483 VDD.n2151 0.0981562
R9658 VDD.n2485 VDD.n2145 0.0981562
R9659 VDD.n2497 VDD.n2496 0.0981562
R9660 VDD.n2509 VDD.n2507 0.0981562
R9661 VDD.n2521 VDD.n2131 0.0981562
R9662 VDD.n2550 VDD.n2113 0.0981562
R9663 VDD.n2564 VDD.n2563 0.0981562
R9664 VDD.n2577 VDD.n2575 0.0981562
R9665 VDD.n2586 VDD.n2098 0.0981562
R9666 VDD.n2588 VDD.n2093 0.0981562
R9667 VDD.n2600 VDD.n2599 0.0981562
R9668 VDD.n2613 VDD.n2612 0.0981562
R9669 VDD.n2624 VDD.n2077 0.0981562
R9670 VDD.n2645 VDD.n2644 0.0981562
R9671 VDD.n2657 VDD.n2655 0.0981562
R9672 VDD.n2668 VDD.n2056 0.0981562
R9673 VDD.n2670 VDD.n2050 0.0981562
R9674 VDD.n2682 VDD.n2681 0.0981562
R9675 VDD.n2694 VDD.n2692 0.0981562
R9676 VDD.n2706 VDD.n2036 0.0981562
R9677 VDD.n2781 VDD.n2780 0.0981562
R9678 VDD.n2793 VDD.n2791 0.0981562
R9679 VDD.n2804 VDD.n1989 0.0981562
R9680 VDD.n2806 VDD.n1983 0.0981562
R9681 VDD.n2818 VDD.n2817 0.0981562
R9682 VDD.n2830 VDD.n2828 0.0981562
R9683 VDD.n2842 VDD.n1969 0.0981562
R9684 VDD.n24 VDD 0.0981562
R9685 VDD.n164 VDD 0.0981562
R9686 VDD.n299 VDD 0.0981562
R9687 VDD.n442 VDD 0.0981562
R9688 VDD.n555 VDD.n551 0.0981562
R9689 VDD.n575 VDD 0.0981562
R9690 VDD.n710 VDD 0.0981562
R9691 VDD.n853 VDD 0.0981562
R9692 VDD VDD.n1936 0.0968542
R9693 VDD.n2956 VDD 0.0968542
R9694 VDD.n3027 VDD 0.0968542
R9695 VDD.n814 VDD.n813 0.0968542
R9696 VDD.n1297 VDD.n1277 0.0960224
R9697 VDD.n1374 VDD.n1235 0.0960224
R9698 VDD.n1451 VDD.n1193 0.0960224
R9699 VDD.n1528 VDD.n1151 0.0960224
R9700 VDD.n1605 VDD.n1109 0.0960224
R9701 VDD.n1682 VDD.n1067 0.0960224
R9702 VDD.n1764 VDD.n1024 0.0960224
R9703 VDD.n125 VDD.n117 0.0960224
R9704 VDD.n138 VDD.n137 0.0960224
R9705 VDD.n811 VDD.n803 0.0960224
R9706 VDD.n825 VDD.n818 0.0960224
R9707 VDD.n827 VDD.n825 0.0960224
R9708 VDD.n684 VDD.n683 0.0960224
R9709 VDD.n683 VDD.n676 0.0960224
R9710 VDD.n549 VDD.n541 0.0960224
R9711 VDD.n400 VDD.n392 0.0960224
R9712 VDD.n416 VDD.n415 0.0960224
R9713 VDD.n415 VDD.n408 0.0960224
R9714 VDD.n265 VDD.n264 0.0960224
R9715 VDD.n2261 VDD 0.0955521
R9716 VDD.n972 VDD.n965 0.0953148
R9717 VDD VDD.n2164 0.09425
R9718 VDD.n960 VDD.n959 0.0825312
R9719 VDD.n128 VDD.n127 0.0773229
R9720 VDD.n403 VDD.n402 0.0773229
R9721 VDD VDD.n2069 0.0760208
R9722 VDD VDD.n2002 0.0760208
R9723 VDD.n197 VDD.n196 0.0738696
R9724 VDD.n57 VDD.n56 0.0738696
R9725 VDD.n332 VDD.n331 0.0738696
R9726 VDD.n475 VDD.n474 0.0738696
R9727 VDD.n608 VDD.n607 0.0738696
R9728 VDD.n743 VDD.n742 0.0738696
R9729 VDD.n886 VDD.n885 0.0738696
R9730 VDD.n3278 VDD 0.0603958
R9731 VDD VDD.n3292 0.0603958
R9732 VDD.n3293 VDD 0.0603958
R9733 VDD VDD.n3301 0.0603958
R9734 VDD.n3368 VDD 0.0603958
R9735 VDD VDD.n3382 0.0603958
R9736 VDD.n3383 VDD 0.0603958
R9737 VDD VDD.n3391 0.0603958
R9738 VDD.n2922 VDD 0.0603958
R9739 VDD.n2982 VDD 0.0603958
R9740 VDD.n3053 VDD 0.0603958
R9741 VDD VDD.n1241 0.0603958
R9742 VDD VDD.n1199 0.0603958
R9743 VDD VDD.n1157 0.0603958
R9744 VDD VDD.n1115 0.0603958
R9745 VDD VDD.n1073 0.0603958
R9746 VDD.n1746 VDD 0.0603958
R9747 VDD VDD.n155 0.0603958
R9748 VDD.n156 VDD 0.0603958
R9749 VDD.n290 VDD 0.0603958
R9750 VDD VDD.n289 0.0603958
R9751 VDD VDD.n433 0.0603958
R9752 VDD.n434 VDD 0.0603958
R9753 VDD VDD.n566 0.0603958
R9754 VDD.n567 VDD 0.0603958
R9755 VDD VDD.n701 0.0603958
R9756 VDD.n702 VDD 0.0603958
R9757 VDD VDD.n844 0.0603958
R9758 VDD.n845 VDD 0.0603958
R9759 VDD VDD.n992 0.0603958
R9760 VDD.n2708 VDD 0.0590938
R9761 VDD.n2844 VDD 0.0590938
R9762 VDD.n193 VDD.n191 0.0412609
R9763 VDD.n53 VDD.n51 0.0412609
R9764 VDD.n328 VDD.n326 0.0412609
R9765 VDD.n471 VDD.n469 0.0412609
R9766 VDD.n604 VDD.n602 0.0412609
R9767 VDD.n739 VDD.n737 0.0412609
R9768 VDD.n882 VDD.n880 0.0412609
R9769 VDD.n2523 VDD 0.0408646
R9770 VDD VDD.n2359 0.0395625
R9771 VDD.n193 VDD 0.0385435
R9772 VDD.n53 VDD 0.0385435
R9773 VDD.n328 VDD 0.0385435
R9774 VDD.n471 VDD 0.0385435
R9775 VDD.n604 VDD 0.0385435
R9776 VDD.n739 VDD 0.0385435
R9777 VDD.n882 VDD 0.0385435
R9778 VDD.n2902 VDD 0.0239375
R9779 VDD VDD.n2955 0.0239375
R9780 VDD VDD.n3026 0.0239375
R9781 VDD.n2632 VDD 0.0226354
R9782 VDD.n2768 VDD 0.0226354
R9783 VDD.n1360 VDD 0.0226354
R9784 VDD.n1437 VDD 0.0226354
R9785 VDD.n1514 VDD 0.0226354
R9786 VDD.n1591 VDD 0.0226354
R9787 VDD.n1668 VDD 0.0226354
R9788 VDD VDD.n1745 0.0226354
R9789 VDD VDD.n1823 0.0226354
R9790 VDD.n127 VDD.n126 0.0226354
R9791 VDD.n156 VDD 0.0226354
R9792 VDD.n289 VDD 0.0226354
R9793 VDD.n402 VDD.n401 0.0226354
R9794 VDD.n434 VDD 0.0226354
R9795 VDD.n551 VDD.n550 0.0226354
R9796 VDD.n567 VDD 0.0226354
R9797 VDD.n702 VDD 0.0226354
R9798 VDD.n813 VDD.n812 0.0226354
R9799 VDD.n845 VDD 0.0226354
R9800 VDD.n3268 VDD 0.0213333
R9801 VDD.n3358 VDD 0.0213333
R9802 VDD.n2260 VDD.n2251 0.0213333
R9803 VDD.n2276 VDD.n2275 0.0213333
R9804 VDD.n2287 VDD.n2286 0.0213333
R9805 VDD.n2298 VDD.n2240 0.0213333
R9806 VDD.n2299 VDD.n2233 0.0213333
R9807 VDD.n2314 VDD.n2313 0.0213333
R9808 VDD.n2326 VDD.n2325 0.0213333
R9809 VDD.n2359 VDD.n2219 0.0213333
R9810 VDD.n2631 VDD.n2630 0.0213333
R9811 VDD.n2643 VDD.n2069 0.0213333
R9812 VDD.n2645 VDD.n2063 0.0213333
R9813 VDD.n2657 VDD.n2656 0.0213333
R9814 VDD.n2669 VDD.n2668 0.0213333
R9815 VDD.n2680 VDD.n2050 0.0213333
R9816 VDD.n2682 VDD.n2044 0.0213333
R9817 VDD.n2694 VDD.n2693 0.0213333
R9818 VDD.n2707 VDD.n2706 0.0213333
R9819 VDD.n2754 VDD 0.0213333
R9820 VDD.n2767 VDD.n2766 0.0213333
R9821 VDD.n2779 VDD.n2002 0.0213333
R9822 VDD.n2781 VDD.n1996 0.0213333
R9823 VDD.n2793 VDD.n2792 0.0213333
R9824 VDD.n2805 VDD.n2804 0.0213333
R9825 VDD.n2816 VDD.n1983 0.0213333
R9826 VDD.n2818 VDD.n1977 0.0213333
R9827 VDD.n2830 VDD.n2829 0.0213333
R9828 VDD.n2843 VDD.n2842 0.0213333
R9829 VDD VDD.n2901 0.0213333
R9830 VDD VDD.n2954 0.0213333
R9831 VDD VDD.n3025 0.0213333
R9832 VDD VDD.n3092 0.0213333
R9833 VDD.n1299 VDD.n1292 0.0213333
R9834 VDD.n1376 VDD.n1369 0.0213333
R9835 VDD.n1453 VDD.n1446 0.0213333
R9836 VDD.n1530 VDD.n1523 0.0213333
R9837 VDD.n1607 VDD.n1600 0.0213333
R9838 VDD.n1684 VDD.n1677 0.0213333
R9839 VDD.n1765 VDD.n1026 0.0213333
R9840 VDD.n139 VDD.n128 0.0213333
R9841 VDD.n417 VDD.n403 0.0213333
R9842 VDD.n685 VDD.n671 0.0213333
R9843 VDD.n829 VDD.n828 0.0213333
R9844 VDD.n2448 VDD.n2447 0.0200312
R9845 VDD.n2459 VDD.n2458 0.0200312
R9846 VDD.n2470 VDD.n2158 0.0200312
R9847 VDD.n2471 VDD.n2151 0.0200312
R9848 VDD.n2485 VDD.n2484 0.0200312
R9849 VDD.n2496 VDD.n2495 0.0200312
R9850 VDD.n2507 VDD.n2139 0.0200312
R9851 VDD.n2508 VDD.n2131 0.0200312
R9852 VDD.n2523 VDD.n2522 0.0200312
R9853 VDD.n974 VDD.n960 0.0200312
R9854 VDD.n266 VDD.n257 0.0198299
R9855 VDD.n959 VDD.n958 0.0187292
R9856 VDD.n2360 VDD.n2213 0.0148229
R9857 VDD.n2372 VDD.n2371 0.0148229
R9858 VDD.n2383 VDD.n2382 0.0148229
R9859 VDD.n2199 VDD.n2197 0.0148229
R9860 VDD.n2396 VDD.n2191 0.0148229
R9861 VDD.n2408 VDD.n2407 0.0148229
R9862 VDD.n2419 VDD.n2418 0.0148229
R9863 VDD.n2179 VDD.n2176 0.0148229
R9864 VDD.n2435 VDD.n2434 0.0148229
R9865 VDD.n2549 VDD.n2548 0.0148229
R9866 VDD.n2113 VDD.n2111 0.0148229
R9867 VDD.n2564 VDD.n2105 0.0148229
R9868 VDD.n2577 VDD.n2576 0.0148229
R9869 VDD.n2587 VDD.n2586 0.0148229
R9870 VDD.n2093 VDD.n2091 0.0148229
R9871 VDD.n2600 VDD.n2083 0.0148229
R9872 VDD.n2614 VDD.n2613 0.0148229
R9873 VDD.n2625 VDD.n2624 0.0148229
R9874 VDD.n2433 VDD 0.0135208
R9875 VDD.n2626 VDD 0.0135208
R9876 VDD.n66 VDD.n65 0.0135208
R9877 VDD.n206 VDD.n205 0.0135208
R9878 VDD.n274 VDD.n268 0.0135208
R9879 VDD.n341 VDD.n340 0.0135208
R9880 VDD.n484 VDD.n483 0.0135208
R9881 VDD.n617 VDD.n616 0.0135208
R9882 VDD.n752 VDD.n751 0.0135208
R9883 VDD.n895 VDD.n894 0.0135208
R9884 VDD.n65 VDD.n50 0.00961458
R9885 VDD.n205 VDD.n190 0.00961458
R9886 VDD.n340 VDD.n325 0.00961458
R9887 VDD.n483 VDD.n468 0.00961458
R9888 VDD.n616 VDD.n601 0.00961458
R9889 VDD.n751 VDD.n736 0.00961458
R9890 VDD.n894 VDD.n879 0.00961458
R9891 VDD.n2370 VDD.n2213 0.0083125
R9892 VDD.n2371 VDD.n2203 0.0083125
R9893 VDD.n2384 VDD.n2383 0.0083125
R9894 VDD.n2395 VDD.n2197 0.0083125
R9895 VDD.n2406 VDD.n2191 0.0083125
R9896 VDD.n2407 VDD.n2183 0.0083125
R9897 VDD.n2420 VDD.n2419 0.0083125
R9898 VDD.n2432 VDD.n2176 0.0083125
R9899 VDD.n2434 VDD.n2433 0.0083125
R9900 VDD.n2550 VDD.n2549 0.0083125
R9901 VDD.n2563 VDD.n2111 0.0083125
R9902 VDD.n2575 VDD.n2105 0.0083125
R9903 VDD.n2576 VDD.n2098 0.0083125
R9904 VDD.n2588 VDD.n2587 0.0083125
R9905 VDD.n2599 VDD.n2091 0.0083125
R9906 VDD.n2612 VDD.n2083 0.0083125
R9907 VDD.n2614 VDD.n2077 0.0083125
R9908 VDD.n2626 VDD.n2625 0.0083125
R9909 VDD.n196 VDD.n191 0.00593478
R9910 VDD.n56 VDD.n51 0.00593478
R9911 VDD.n331 VDD.n326 0.00593478
R9912 VDD.n474 VDD.n469 0.00593478
R9913 VDD.n607 VDD.n602 0.00593478
R9914 VDD.n742 VDD.n737 0.00593478
R9915 VDD.n885 VDD.n880 0.00593478
R9916 VDD.n2448 VDD 0.00440625
R9917 VDD.n958 VDD.n946 0.00440625
R9918 VDD.n2447 VDD.n2446 0.00310417
R9919 VDD.n2458 VDD.n2164 0.00310417
R9920 VDD.n2460 VDD.n2158 0.00310417
R9921 VDD.n2472 VDD.n2471 0.00310417
R9922 VDD.n2484 VDD.n2483 0.00310417
R9923 VDD.n2495 VDD.n2145 0.00310417
R9924 VDD.n2497 VDD.n2139 0.00310417
R9925 VDD.n2509 VDD.n2508 0.00310417
R9926 VDD.n2522 VDD.n2521 0.00310417
R9927 VDD.n975 VDD.n974 0.00310417
R9928 VDD.n2261 VDD.n2260 0.00180208
R9929 VDD.n2275 VDD.n2274 0.00180208
R9930 VDD.n2286 VDD.n2246 0.00180208
R9931 VDD.n2288 VDD.n2240 0.00180208
R9932 VDD.n2300 VDD.n2299 0.00180208
R9933 VDD.n2313 VDD.n2312 0.00180208
R9934 VDD.n2325 VDD.n2227 0.00180208
R9935 VDD.n2327 VDD.n2219 0.00180208
R9936 VDD.n2632 VDD.n2631 0.00180208
R9937 VDD.n2644 VDD.n2643 0.00180208
R9938 VDD.n2655 VDD.n2063 0.00180208
R9939 VDD.n2656 VDD.n2056 0.00180208
R9940 VDD.n2670 VDD.n2669 0.00180208
R9941 VDD.n2681 VDD.n2680 0.00180208
R9942 VDD.n2692 VDD.n2044 0.00180208
R9943 VDD.n2693 VDD.n2036 0.00180208
R9944 VDD.n2708 VDD.n2707 0.00180208
R9945 VDD.n2768 VDD.n2767 0.00180208
R9946 VDD.n2780 VDD.n2779 0.00180208
R9947 VDD.n2791 VDD.n1996 0.00180208
R9948 VDD.n2792 VDD.n1989 0.00180208
R9949 VDD.n2806 VDD.n2805 0.00180208
R9950 VDD.n2817 VDD.n2816 0.00180208
R9951 VDD.n2828 VDD.n1977 0.00180208
R9952 VDD.n2829 VDD.n1969 0.00180208
R9953 VDD.n2844 VDD.n2843 0.00180208
R9954 VDD.n1292 VDD.n1276 0.00180208
R9955 VDD.n1369 VDD.n1234 0.00180208
R9956 VDD.n1446 VDD.n1192 0.00180208
R9957 VDD.n1523 VDD.n1150 0.00180208
R9958 VDD.n1600 VDD.n1108 0.00180208
R9959 VDD.n1677 VDD.n1066 0.00180208
R9960 VDD.n1766 VDD.n1765 0.00180208
R9961 VDD.n140 VDD.n139 0.00180208
R9962 VDD.n257 VDD.n256 0.00180208
R9963 VDD.n418 VDD.n417 0.00180208
R9964 VDD.n686 VDD.n685 0.00180208
R9965 VDD.n828 VDD.n814 0.00180208
R9966 VDD.n267 VDD.n266 0.00178866
R9967 x2.X.n138 x2.X.t47 396.834
R9968 x2.X.n117 x2.X.t49 396.834
R9969 x2.X.n96 x2.X.t42 396.834
R9970 x2.X.n75 x2.X.t37 396.834
R9971 x2.X.n54 x2.X.t68 396.834
R9972 x2.X.n33 x2.X.t66 396.834
R9973 x2.X.n13 x2.X.t52 396.834
R9974 x2.X.n133 x2.X.t35 381.228
R9975 x2.X.n112 x2.X.t33 381.228
R9976 x2.X.n91 x2.X.t60 381.228
R9977 x2.X.n70 x2.X.t58 381.228
R9978 x2.X.n49 x2.X.t39 381.228
R9979 x2.X.n28 x2.X.t72 381.228
R9980 x2.X.n8 x2.X.t69 381.228
R9981 x2.X.n127 x2.X.t44 198.335
R9982 x2.X.n106 x2.X.t32 198.335
R9983 x2.X.n85 x2.X.t71 198.335
R9984 x2.X.n64 x2.X.t56 198.335
R9985 x2.X.n43 x2.X.t54 198.335
R9986 x2.X.n23 x2.X.t50 198.335
R9987 x2.X.n148 x2.X.t34 198.025
R9988 x2.X.n149 x2.X.t53 172.463
R9989 x2.X.n128 x2.X.t62 171.875
R9990 x2.X.n107 x2.X.t48 171.875
R9991 x2.X.n86 x2.X.t41 171.875
R9992 x2.X.n65 x2.X.t73 171.875
R9993 x2.X.n44 x2.X.t70 171.875
R9994 x2.X.n24 x2.X.t65 171.875
R9995 x2.X.n135 x2.X.n134 152
R9996 x2.X.n114 x2.X.n113 152
R9997 x2.X.n93 x2.X.n92 152
R9998 x2.X.n72 x2.X.n71 152
R9999 x2.X.n51 x2.X.n50 152
R10000 x2.X.n30 x2.X.n29 152
R10001 x2.X.n10 x2.X.n9 152
R10002 x2.X.n161 x2.X.n160 146.812
R10003 x2.X.n135 x2.X.t64 136.745
R10004 x2.X.n114 x2.X.t61 136.745
R10005 x2.X.n93 x2.X.t46 136.745
R10006 x2.X.n72 x2.X.t38 136.745
R10007 x2.X.n51 x2.X.t59 136.745
R10008 x2.X.n30 x2.X.t57 136.745
R10009 x2.X.n10 x2.X.t55 136.745
R10010 x2.X.n138 x2.X.t43 134.065
R10011 x2.X.n117 x2.X.t45 134.065
R10012 x2.X.n96 x2.X.t40 134.065
R10013 x2.X.n75 x2.X.t36 134.065
R10014 x2.X.n54 x2.X.t67 134.065
R10015 x2.X.n33 x2.X.t63 134.065
R10016 x2.X.n13 x2.X.t51 134.065
R10017 x2.X.n167 x2.X.n153 108.412
R10018 x2.X.n166 x2.X.n154 108.412
R10019 x2.X.n165 x2.X.n155 108.412
R10020 x2.X.n164 x2.X.n156 108.412
R10021 x2.X.n163 x2.X.n157 108.412
R10022 x2.X.n162 x2.X.n158 108.412
R10023 x2.X.n161 x2.X.n159 108.412
R10024 x2.X.n171 x2.X.n169 90.8321
R10025 x2.X.n133 x2.X.n132 75.1188
R10026 x2.X.n112 x2.X.n111 75.1188
R10027 x2.X.n91 x2.X.n90 75.1188
R10028 x2.X.n70 x2.X.n69 75.1188
R10029 x2.X.n49 x2.X.n48 75.1188
R10030 x2.X.n28 x2.X.n27 75.1188
R10031 x2.X.n8 x2.X.n7 75.1188
R10032 x2.X.n171 x2.X.n170 52.4321
R10033 x2.X.n173 x2.X.n172 52.4321
R10034 x2.X.n175 x2.X.n174 52.4321
R10035 x2.X.n177 x2.X.n176 52.4321
R10036 x2.X.n179 x2.X.n178 52.4321
R10037 x2.X.n181 x2.X.n180 52.4321
R10038 x2.X.n183 x2.X.n182 52.4321
R10039 x2.X x2.X.n183 40.4711
R10040 x2.X.n173 x2.X.n171 38.4005
R10041 x2.X.n175 x2.X.n173 38.4005
R10042 x2.X.n177 x2.X.n175 38.4005
R10043 x2.X.n179 x2.X.n177 38.4005
R10044 x2.X.n181 x2.X.n179 38.4005
R10045 x2.X.n183 x2.X.n181 38.4005
R10046 x2.X.n167 x2.X.n166 38.4005
R10047 x2.X.n166 x2.X.n165 38.4005
R10048 x2.X.n165 x2.X.n164 38.4005
R10049 x2.X.n164 x2.X.n163 38.4005
R10050 x2.X.n163 x2.X.n162 38.4005
R10051 x2.X.n162 x2.X.n161 38.4005
R10052 x2.X x2.X.n167 33.7342
R10053 x2.X.n168 x2.X.n152 26.8074
R10054 x2.X.n153 x2.X.t19 26.5955
R10055 x2.X.n153 x2.X.t30 26.5955
R10056 x2.X.n154 x2.X.t24 26.5955
R10057 x2.X.n154 x2.X.t29 26.5955
R10058 x2.X.n155 x2.X.t22 26.5955
R10059 x2.X.n155 x2.X.t27 26.5955
R10060 x2.X.n156 x2.X.t20 26.5955
R10061 x2.X.n156 x2.X.t26 26.5955
R10062 x2.X.n157 x2.X.t18 26.5955
R10063 x2.X.n157 x2.X.t17 26.5955
R10064 x2.X.n158 x2.X.t25 26.5955
R10065 x2.X.n158 x2.X.t16 26.5955
R10066 x2.X.n159 x2.X.t23 26.5955
R10067 x2.X.n159 x2.X.t28 26.5955
R10068 x2.X.n160 x2.X.t21 26.5955
R10069 x2.X.n160 x2.X.t31 26.5955
R10070 x2.X.n169 x2.X.t11 24.9236
R10071 x2.X.n169 x2.X.t5 24.9236
R10072 x2.X.n170 x2.X.t13 24.9236
R10073 x2.X.n170 x2.X.t2 24.9236
R10074 x2.X.n172 x2.X.t15 24.9236
R10075 x2.X.n172 x2.X.t6 24.9236
R10076 x2.X.n174 x2.X.t8 24.9236
R10077 x2.X.n174 x2.X.t7 24.9236
R10078 x2.X.n176 x2.X.t10 24.9236
R10079 x2.X.n176 x2.X.t0 24.9236
R10080 x2.X.n178 x2.X.t12 24.9236
R10081 x2.X.n178 x2.X.t1 24.9236
R10082 x2.X.n180 x2.X.t14 24.9236
R10083 x2.X.n180 x2.X.t3 24.9236
R10084 x2.X.n182 x2.X.t9 24.9236
R10085 x2.X.n182 x2.X.t4 24.9236
R10086 x2.X.n140 x2.X 13.6005
R10087 x2.X.n119 x2.X 13.6005
R10088 x2.X.n98 x2.X 13.6005
R10089 x2.X.n77 x2.X 13.6005
R10090 x2.X.n56 x2.X 13.6005
R10091 x2.X.n35 x2.X 13.6005
R10092 x2.X.n15 x2.X 13.6005
R10093 x2.X.n135 x2.X.n133 13.3692
R10094 x2.X.n114 x2.X.n112 13.3692
R10095 x2.X.n93 x2.X.n91 13.3692
R10096 x2.X.n72 x2.X.n70 13.3692
R10097 x2.X.n51 x2.X.n49 13.3692
R10098 x2.X.n30 x2.X.n28 13.3692
R10099 x2.X.n10 x2.X.n8 13.3692
R10100 x2.X.n47 x2.X.n26 13.2412
R10101 x2.X.n152 x2.X.n151 11.2004
R10102 x2.X.n134 x2.X 11.055
R10103 x2.X.n113 x2.X 11.055
R10104 x2.X.n92 x2.X 11.055
R10105 x2.X.n71 x2.X 11.055
R10106 x2.X.n50 x2.X 11.055
R10107 x2.X.n29 x2.X 11.055
R10108 x2.X.n9 x2.X 11.055
R10109 x2.X.n136 x2.X.n135 9.3005
R10110 x2.X.n150 x2.X.n149 9.3005
R10111 x2.X.n115 x2.X.n114 9.3005
R10112 x2.X.n129 x2.X.n128 9.3005
R10113 x2.X.n94 x2.X.n93 9.3005
R10114 x2.X.n108 x2.X.n107 9.3005
R10115 x2.X.n73 x2.X.n72 9.3005
R10116 x2.X.n87 x2.X.n86 9.3005
R10117 x2.X.n52 x2.X.n51 9.3005
R10118 x2.X.n66 x2.X.n65 9.3005
R10119 x2.X.n31 x2.X.n30 9.3005
R10120 x2.X.n45 x2.X.n44 9.3005
R10121 x2.X.n11 x2.X.n10 9.3005
R10122 x2.X.n25 x2.X.n24 9.3005
R10123 x2.X.n151 x2.X.n150 9.23046
R10124 x2.X.n46 x2.X.n45 9.10496
R10125 x2.X.n26 x2.X.n25 9.10496
R10126 x2.X.n109 x2.X.n108 9.10363
R10127 x2.X.n88 x2.X.n87 9.10363
R10128 x2.X.n67 x2.X.n66 9.1023
R10129 x2.X.n130 x2.X.n129 8.98032
R10130 x2.X.n168 x2.X 8.75839
R10131 x2.X.n89 x2.X.n68 8.70611
R10132 x2.X.n68 x2.X.n47 8.70243
R10133 x2.X.n131 x2.X.n110 8.70243
R10134 x2.X.n110 x2.X.n89 8.69014
R10135 x2.X.n139 x2.X.n138 6.98562
R10136 x2.X.n118 x2.X.n117 6.98562
R10137 x2.X.n97 x2.X.n96 6.98562
R10138 x2.X.n76 x2.X.n75 6.98562
R10139 x2.X.n55 x2.X.n54 6.98562
R10140 x2.X.n34 x2.X.n33 6.98562
R10141 x2.X.n14 x2.X.n13 6.98562
R10142 x2.X.n128 x2.X.n127 5.7706
R10143 x2.X.n107 x2.X.n106 5.7706
R10144 x2.X.n86 x2.X.n85 5.7706
R10145 x2.X.n65 x2.X.n64 5.7706
R10146 x2.X.n44 x2.X.n43 5.7706
R10147 x2.X.n24 x2.X.n23 5.7706
R10148 x2.X.n149 x2.X.n148 5.46089
R10149 x2.X.n131 x2.X.n130 4.53188
R10150 x2.X.n110 x2.X.n109 4.53188
R10151 x2.X.n89 x2.X.n88 4.53188
R10152 x2.X.n68 x2.X.n67 4.53188
R10153 x2.X.n47 x2.X.n46 4.53188
R10154 x2.X.n0 x2.X.n141 4.46483
R10155 x2.X.n1 x2.X.n120 4.46483
R10156 x2.X.n2 x2.X.n99 4.46483
R10157 x2.X.n3 x2.X.n78 4.46483
R10158 x2.X.n4 x2.X.n57 4.46483
R10159 x2.X.n5 x2.X.n36 4.46483
R10160 x2.X.n6 x2.X.n16 4.46483
R10161 x2.X.n126 x2.X.n125 4.17441
R10162 x2.X.n105 x2.X.n104 4.17441
R10163 x2.X.n63 x2.X.n62 4.17441
R10164 x2.X.n22 x2.X.n21 4.17441
R10165 x2.X.n147 x2.X.n146 3.89615
R10166 x2.X.n84 x2.X.n83 3.89615
R10167 x2.X.n42 x2.X.n41 3.89615
R10168 x2.X.n134 x2.X.n132 2.90959
R10169 x2.X.n113 x2.X.n111 2.90959
R10170 x2.X.n92 x2.X.n90 2.90959
R10171 x2.X.n71 x2.X.n69 2.90959
R10172 x2.X.n50 x2.X.n48 2.90959
R10173 x2.X.n29 x2.X.n27 2.90959
R10174 x2.X.n9 x2.X.n7 2.90959
R10175 x2.X.n141 x2.X 2.89456
R10176 x2.X.n120 x2.X 2.89456
R10177 x2.X.n99 x2.X 2.89456
R10178 x2.X.n78 x2.X 2.89456
R10179 x2.X.n57 x2.X 2.89456
R10180 x2.X.n36 x2.X 2.89456
R10181 x2.X.n16 x2.X 2.89456
R10182 x2.X x2.X.n136 2.75432
R10183 x2.X x2.X.n115 2.75432
R10184 x2.X x2.X.n94 2.75432
R10185 x2.X x2.X.n73 2.75432
R10186 x2.X x2.X.n52 2.75432
R10187 x2.X x2.X.n31 2.75432
R10188 x2.X x2.X.n11 2.75432
R10189 x2.X x2.X.n168 2.69524
R10190 x2.X.n140 x2.X.n139 2.52171
R10191 x2.X.n119 x2.X.n118 2.52171
R10192 x2.X.n98 x2.X.n97 2.52171
R10193 x2.X.n77 x2.X.n76 2.52171
R10194 x2.X.n56 x2.X.n55 2.52171
R10195 x2.X.n35 x2.X.n34 2.52171
R10196 x2.X.n15 x2.X.n14 2.52171
R10197 x2.X.n146 x2.X 2.50485
R10198 x2.X.n83 x2.X 2.50485
R10199 x2.X.n41 x2.X 2.50485
R10200 x2.X.n151 x2.X.n145 2.2505
R10201 x2.X.n130 x2.X.n124 2.2505
R10202 x2.X.n109 x2.X.n103 2.2505
R10203 x2.X.n88 x2.X.n82 2.2505
R10204 x2.X.n67 x2.X.n61 2.2505
R10205 x2.X.n46 x2.X.n40 2.2505
R10206 x2.X.n26 x2.X.n20 2.2505
R10207 x2.X.n125 x2.X 2.22659
R10208 x2.X.n104 x2.X 2.22659
R10209 x2.X.n62 x2.X 2.22659
R10210 x2.X.n21 x2.X 2.22659
R10211 x2.X.n152 x2.X.n131 1.94561
R10212 x2.X.n137 x2.X 1.89782
R10213 x2.X.n53 x2.X 1.89782
R10214 x2.X.n32 x2.X 1.89782
R10215 x2.X.n12 x2.X 1.89782
R10216 x2.X.n116 x2.X 1.89336
R10217 x2.X.n95 x2.X 1.89336
R10218 x2.X.n74 x2.X 1.89336
R10219 x2.X.n116 x2.X 1.45586
R10220 x2.X.n95 x2.X 1.45586
R10221 x2.X.n74 x2.X 1.45586
R10222 x2.X.n137 x2.X 1.45139
R10223 x2.X.n53 x2.X 1.45139
R10224 x2.X.n32 x2.X 1.45139
R10225 x2.X.n12 x2.X 1.45139
R10226 x2.X.n123 x2.X.n122 0.955857
R10227 x2.X.n102 x2.X.n101 0.955857
R10228 x2.X.n81 x2.X.n80 0.955857
R10229 x2.X.n144 x2.X.n143 0.951393
R10230 x2.X.n60 x2.X.n59 0.951393
R10231 x2.X.n39 x2.X.n38 0.951393
R10232 x2.X.n19 x2.X.n18 0.951393
R10233 x2.X.n150 x2.X.n147 0.835283
R10234 x2.X.n87 x2.X.n84 0.835283
R10235 x2.X.n45 x2.X.n42 0.835283
R10236 x2.X.n129 x2.X.n126 0.557022
R10237 x2.X.n108 x2.X.n105 0.557022
R10238 x2.X.n66 x2.X.n63 0.557022
R10239 x2.X.n25 x2.X.n22 0.557022
R10240 x2.X.n123 x2.X 0.53175
R10241 x2.X.n102 x2.X 0.53175
R10242 x2.X.n81 x2.X 0.53175
R10243 x2.X.n144 x2.X 0.529797
R10244 x2.X.n39 x2.X 0.529797
R10245 x2.X.n19 x2.X 0.529797
R10246 x2.X.n60 x2.X 0.513758
R10247 x2.X.n136 x2.X.n132 0.388379
R10248 x2.X.n115 x2.X.n111 0.388379
R10249 x2.X.n94 x2.X.n90 0.388379
R10250 x2.X.n73 x2.X.n69 0.388379
R10251 x2.X.n52 x2.X.n48 0.388379
R10252 x2.X.n31 x2.X.n27 0.388379
R10253 x2.X.n11 x2.X.n7 0.388379
R10254 x2.X.n141 x2.X.n140 0.373349
R10255 x2.X.n120 x2.X.n119 0.373349
R10256 x2.X.n99 x2.X.n98 0.373349
R10257 x2.X.n78 x2.X.n77 0.373349
R10258 x2.X.n57 x2.X.n56 0.373349
R10259 x2.X.n36 x2.X.n35 0.373349
R10260 x2.X.n16 x2.X.n15 0.373349
R10261 x2.X.n143 x2.X 0.259429
R10262 x2.X.n122 x2.X 0.259429
R10263 x2.X.n101 x2.X 0.259429
R10264 x2.X.n80 x2.X 0.259429
R10265 x2.X.n59 x2.X 0.259429
R10266 x2.X.n38 x2.X 0.259429
R10267 x2.X.n18 x2.X 0.259429
R10268 x2.X.n143 x2.X.n0 0.076587
R10269 x2.X.n122 x2.X.n1 0.076587
R10270 x2.X.n101 x2.X.n2 0.076587
R10271 x2.X.n80 x2.X.n3 0.076587
R10272 x2.X.n59 x2.X.n4 0.076587
R10273 x2.X.n38 x2.X.n5 0.076587
R10274 x2.X.n18 x2.X.n6 0.076587
R10275 x2.X.n145 x2.X.n137 0.0532344
R10276 x2.X.n145 x2.X.n144 0.0532344
R10277 x2.X.n124 x2.X.n116 0.0532344
R10278 x2.X.n124 x2.X.n123 0.0532344
R10279 x2.X.n103 x2.X.n95 0.0532344
R10280 x2.X.n103 x2.X.n102 0.0532344
R10281 x2.X.n82 x2.X.n74 0.0532344
R10282 x2.X.n82 x2.X.n81 0.0532344
R10283 x2.X.n40 x2.X.n32 0.0532344
R10284 x2.X.n40 x2.X.n39 0.0532344
R10285 x2.X.n20 x2.X.n12 0.0532344
R10286 x2.X.n20 x2.X.n19 0.0532344
R10287 x2.X.n61 x2.X.n53 0.0516364
R10288 x2.X.n61 x2.X.n60 0.0516364
R10289 x2.X.n6 x2.X.n17 0.0466957
R10290 x2.X.n5 x2.X.n37 0.0466957
R10291 x2.X.n4 x2.X.n58 0.0466957
R10292 x2.X.n3 x2.X.n79 0.0466957
R10293 x2.X.n2 x2.X.n100 0.0466957
R10294 x2.X.n1 x2.X.n121 0.0466957
R10295 x2.X.n0 x2.X.n142 0.0466957
R10296 x2.X.n142 x2.X 0.0358261
R10297 x2.X.n121 x2.X 0.0358261
R10298 x2.X.n100 x2.X 0.0358261
R10299 x2.X.n79 x2.X 0.0358261
R10300 x2.X.n58 x2.X 0.0358261
R10301 x2.X.n37 x2.X 0.0358261
R10302 x2.X.n17 x2.X 0.0358261
R10303 x9.A1.n88 x9.A1.t41 327.974
R10304 x9.A1.n105 x9.A1.t45 327.961
R10305 x9.A1.n121 x9.A1.t47 327.961
R10306 x9.A1.n137 x9.A1.t38 327.599
R10307 x9.A1.n70 x9.A1.t58 327.584
R10308 x9.A1.n34 x9.A1.t43 327.584
R10309 x9.A1.n52 x9.A1.t56 327.57
R10310 x9.A1.n76 x9.A1.t34 327.361
R10311 x9.A1.n40 x9.A1.t53 327.361
R10312 x9.A1.n110 x9.A1.t46 327.337
R10313 x9.A1.n126 x9.A1.t39 327.337
R10314 x9.A1.n94 x9.A1.t51 326.986
R10315 x9.A1.n58 x9.A1.t48 326.986
R10316 x9.A1.n23 x9.A1.t42 326.986
R10317 x9.A1.n50 x9.A1.t44 151.681
R10318 x9.A1.n103 x9.A1.t36 150.825
R10319 x9.A1.n119 x9.A1.t37 150.825
R10320 x9.A1.n86 x9.A1.t59 150.81
R10321 x9.A1.n68 x9.A1.t57 150.794
R10322 x9.A1.n32 x9.A1.t32 150.794
R10323 x9.A1.n111 x9.A1.t49 150.78
R10324 x9.A1.n127 x9.A1.t50 150.78
R10325 x9.A1.n135 x9.A1.t52 150.78
R10326 x9.A1.n77 x9.A1.t33 149.893
R10327 x9.A1.n41 x9.A1.t40 149.893
R10328 x9.A1.n95 x9.A1.t54 149.862
R10329 x9.A1.n59 x9.A1.t35 149.862
R10330 x9.A1.n24 x9.A1.t55 149.862
R10331 x9.A1.n10 x9.A1.n8 146.811
R10332 x9.A1.n20 x9.A1.n19 108.412
R10333 x9.A1.n21 x9.A1.n7 108.412
R10334 x9.A1.n10 x9.A1.n9 108.412
R10335 x9.A1.n12 x9.A1.n11 108.412
R10336 x9.A1.n14 x9.A1.n13 108.412
R10337 x9.A1.n16 x9.A1.n15 108.412
R10338 x9.A1.n18 x9.A1.n17 108.412
R10339 x9.A1.n150 x9.A1.n148 90.8321
R10340 x9.A1.n150 x9.A1.n149 52.4321
R10341 x9.A1.n152 x9.A1.n151 52.4321
R10342 x9.A1.n154 x9.A1.n153 52.4321
R10343 x9.A1.n156 x9.A1.n155 52.4321
R10344 x9.A1.n158 x9.A1.n157 52.4321
R10345 x9.A1.n160 x9.A1.n159 52.4321
R10346 x9.A1.n162 x9.A1.n161 52.4321
R10347 x9.A1 x9.A1.n162 40.4711
R10348 x9.A1.n152 x9.A1.n150 38.4005
R10349 x9.A1.n154 x9.A1.n152 38.4005
R10350 x9.A1.n156 x9.A1.n154 38.4005
R10351 x9.A1.n158 x9.A1.n156 38.4005
R10352 x9.A1.n160 x9.A1.n158 38.4005
R10353 x9.A1.n162 x9.A1.n160 38.4005
R10354 x9.A1.n12 x9.A1.n10 38.4005
R10355 x9.A1.n14 x9.A1.n12 38.4005
R10356 x9.A1.n16 x9.A1.n14 38.4005
R10357 x9.A1.n18 x9.A1.n16 38.4005
R10358 x9.A1.n20 x9.A1.n18 38.4005
R10359 x9.A1.n21 x9.A1.n20 38.4005
R10360 x9.A1 x9.A1.n21 33.7342
R10361 x9.A1.n95 x9.A1 29.1167
R10362 x9.A1.n59 x9.A1 29.1167
R10363 x9.A1.n24 x9.A1 29.1167
R10364 x9.A1.n77 x9.A1 28.9113
R10365 x9.A1.n41 x9.A1 28.9113
R10366 x9.A1.n111 x9.A1 28.5657
R10367 x9.A1.n127 x9.A1 28.5657
R10368 x9.A1.n135 x9.A1 28.5657
R10369 x9.A1.n86 x9.A1 28.3628
R10370 x9.A1.n68 x9.A1 28.246
R10371 x9.A1.n32 x9.A1 28.246
R10372 x9.A1.n103 x9.A1 28.0462
R10373 x9.A1.n119 x9.A1 28.0462
R10374 x9.A1.n50 x9.A1 27.901
R10375 x9.A1.n7 x9.A1.t24 26.5955
R10376 x9.A1.n7 x9.A1.t18 26.5955
R10377 x9.A1.n8 x9.A1.t28 26.5955
R10378 x9.A1.n8 x9.A1.t20 26.5955
R10379 x9.A1.n9 x9.A1.t27 26.5955
R10380 x9.A1.n9 x9.A1.t22 26.5955
R10381 x9.A1.n11 x9.A1.t30 26.5955
R10382 x9.A1.n11 x9.A1.t16 26.5955
R10383 x9.A1.n13 x9.A1.t25 26.5955
R10384 x9.A1.n13 x9.A1.t17 26.5955
R10385 x9.A1.n15 x9.A1.t26 26.5955
R10386 x9.A1.n15 x9.A1.t19 26.5955
R10387 x9.A1.n17 x9.A1.t29 26.5955
R10388 x9.A1.n17 x9.A1.t21 26.5955
R10389 x9.A1.n19 x9.A1.t31 26.5955
R10390 x9.A1.n19 x9.A1.t23 26.5955
R10391 x9.A1.n148 x9.A1.t4 24.9236
R10392 x9.A1.n148 x9.A1.t12 24.9236
R10393 x9.A1.n149 x9.A1.t3 24.9236
R10394 x9.A1.n149 x9.A1.t14 24.9236
R10395 x9.A1.n151 x9.A1.t6 24.9236
R10396 x9.A1.n151 x9.A1.t8 24.9236
R10397 x9.A1.n153 x9.A1.t1 24.9236
R10398 x9.A1.n153 x9.A1.t9 24.9236
R10399 x9.A1.n155 x9.A1.t2 24.9236
R10400 x9.A1.n155 x9.A1.t11 24.9236
R10401 x9.A1.n157 x9.A1.t5 24.9236
R10402 x9.A1.n157 x9.A1.t13 24.9236
R10403 x9.A1.n159 x9.A1.t7 24.9236
R10404 x9.A1.n159 x9.A1.t15 24.9236
R10405 x9.A1.n161 x9.A1.t0 24.9236
R10406 x9.A1.n161 x9.A1.t10 24.9236
R10407 x9.A1.n147 x9.A1.n146 11.2712
R10408 x9.A1.n147 x9.A1 8.42155
R10409 x9.A1.n38 x9.A1.n30 8.31458
R10410 x9.A1.n141 x9.A1.n140 8.3109
R10411 x9.A1.n74 x9.A1.n66 4.55989
R10412 x9.A1.n143 x9.A1.n142 4.55254
R10413 x9.A1.n92 x9.A1.n84 4.55254
R10414 x9.A1.n145 x9.A1.n144 4.54886
R10415 x9.A1.n56 x9.A1.n48 4.54886
R10416 x9.A1.n48 x9.A1.n38 4.07827
R10417 x9.A1.n142 x9.A1.n141 4.07459
R10418 x9.A1.n144 x9.A1.n143 4.07459
R10419 x9.A1.n84 x9.A1.n74 4.07092
R10420 x9.A1.n66 x9.A1.n56 4.06724
R10421 x9.A1.n145 x9.A1.n101 3.75519
R10422 x9.A1.n144 x9.A1.n108 3.75519
R10423 x9.A1.n143 x9.A1.n117 3.75519
R10424 x9.A1.n142 x9.A1.n124 3.75519
R10425 x9.A1.n141 x9.A1.n133 3.75519
R10426 x9.A1.n92 x9.A1.n91 3.75519
R10427 x9.A1.n84 x9.A1.n83 3.75519
R10428 x9.A1.n74 x9.A1.n73 3.75519
R10429 x9.A1.n66 x9.A1.n65 3.75519
R10430 x9.A1.n56 x9.A1.n55 3.75519
R10431 x9.A1.n48 x9.A1.n47 3.75519
R10432 x9.A1.n38 x9.A1.n37 3.75519
R10433 x9.A1.n138 x9.A1.n137 3.44665
R10434 x9.A1.n89 x9.A1.n88 3.44665
R10435 x9.A1.n106 x9.A1.n105 3.38163
R10436 x9.A1.n122 x9.A1.n121 3.38163
R10437 x9.A1.n71 x9.A1.n70 3.38163
R10438 x9.A1.n35 x9.A1.n34 3.38163
R10439 x9.A1.n53 x9.A1.n52 3.31902
R10440 x9.A1.n146 x9.A1.n145 3.25601
R10441 x9.A1.n98 x9.A1.n97 3.03311
R10442 x9.A1.n0 x9.A1.n106 3.03311
R10443 x9.A1.n114 x9.A1.n113 3.03311
R10444 x9.A1.n1 x9.A1.n122 3.03311
R10445 x9.A1.n130 x9.A1.n129 3.03311
R10446 x9.A1.n2 x9.A1.n138 3.03311
R10447 x9.A1.n3 x9.A1.n89 3.03311
R10448 x9.A1.n80 x9.A1.n79 3.03311
R10449 x9.A1.n4 x9.A1.n71 3.03311
R10450 x9.A1.n62 x9.A1.n61 3.03311
R10451 x9.A1.n5 x9.A1.n53 3.03311
R10452 x9.A1.n44 x9.A1.n43 3.03311
R10453 x9.A1.n6 x9.A1.n35 3.03311
R10454 x9.A1.n27 x9.A1.n26 3.03311
R10455 x9.A1 x9.A1.n147 3.03208
R10456 x9.A1.n97 x9.A1.n94 3.01226
R10457 x9.A1.n79 x9.A1.n76 3.01226
R10458 x9.A1.n61 x9.A1.n58 3.01226
R10459 x9.A1.n43 x9.A1.n40 3.01226
R10460 x9.A1.n26 x9.A1.n23 3.01226
R10461 x9.A1.n113 x9.A1.n110 2.95435
R10462 x9.A1.n129 x9.A1.n126 2.95435
R10463 x9.A1.n107 x9.A1.n0 1.50871
R10464 x9.A1.n123 x9.A1.n1 1.50871
R10465 x9.A1.n139 x9.A1.n2 1.50871
R10466 x9.A1.n90 x9.A1.n3 1.50871
R10467 x9.A1.n72 x9.A1.n4 1.50871
R10468 x9.A1.n54 x9.A1.n5 1.50871
R10469 x9.A1.n36 x9.A1.n6 1.50871
R10470 x9.A1.n100 x9.A1.n99 1.50153
R10471 x9.A1.n116 x9.A1.n115 1.50153
R10472 x9.A1.n132 x9.A1.n131 1.50153
R10473 x9.A1.n82 x9.A1.n81 1.50153
R10474 x9.A1.n64 x9.A1.n63 1.50153
R10475 x9.A1.n46 x9.A1.n45 1.50153
R10476 x9.A1.n29 x9.A1.n28 1.50153
R10477 x9.A1.n97 x9.A1.n96 1.2554
R10478 x9.A1.n79 x9.A1.n78 1.2554
R10479 x9.A1.n61 x9.A1.n60 1.2554
R10480 x9.A1.n43 x9.A1.n42 1.2554
R10481 x9.A1.n26 x9.A1.n25 1.2554
R10482 x9.A1.n113 x9.A1.n112 1.23127
R10483 x9.A1.n129 x9.A1.n128 1.23127
R10484 x9.A1.n146 x9.A1.n92 0.741309
R10485 x9.A1.n138 x9.A1.n136 0.738962
R10486 x9.A1.n89 x9.A1.n87 0.738962
R10487 x9.A1.n106 x9.A1.n104 0.725028
R10488 x9.A1.n122 x9.A1.n120 0.725028
R10489 x9.A1.n71 x9.A1.n69 0.725028
R10490 x9.A1.n35 x9.A1.n33 0.725028
R10491 x9.A1.n53 x9.A1.n51 0.711611
R10492 x9.A1.n96 x9.A1.n95 0.213762
R10493 x9.A1.n60 x9.A1.n59 0.213762
R10494 x9.A1.n25 x9.A1.n24 0.213762
R10495 x9.A1.n78 x9.A1.n77 0.178608
R10496 x9.A1.n42 x9.A1.n41 0.178608
R10497 x9.A1.n112 x9.A1.n111 0.178047
R10498 x9.A1.n128 x9.A1.n127 0.178047
R10499 x9.A1.n136 x9.A1.n135 0.178047
R10500 x9.A1.n69 x9.A1.n68 0.161787
R10501 x9.A1.n33 x9.A1.n32 0.161787
R10502 x9.A1.n51 x9.A1.n50 0.161251
R10503 x9.A1.n87 x9.A1.n86 0.143169
R10504 x9.A1.n104 x9.A1.n103 0.127479
R10505 x9.A1.n120 x9.A1.n119 0.127479
R10506 x9.A1.n6 x9.A1.n31 0.0373802
R10507 x9.A1.n5 x9.A1.n49 0.0373802
R10508 x9.A1.n4 x9.A1.n67 0.0373802
R10509 x9.A1.n3 x9.A1.n85 0.0373802
R10510 x9.A1.n2 x9.A1.n134 0.0373802
R10511 x9.A1.n1 x9.A1.n118 0.0373802
R10512 x9.A1.n0 x9.A1.n102 0.0373802
R10513 x9.A1.n101 x9.A1.n100 0.0226928
R10514 x9.A1.n108 x9.A1.n107 0.0226928
R10515 x9.A1.n117 x9.A1.n116 0.0226928
R10516 x9.A1.n124 x9.A1.n123 0.0226928
R10517 x9.A1.n133 x9.A1.n132 0.0226928
R10518 x9.A1.n140 x9.A1.n139 0.0226928
R10519 x9.A1.n91 x9.A1.n90 0.0226928
R10520 x9.A1.n83 x9.A1.n82 0.0226928
R10521 x9.A1.n73 x9.A1.n72 0.0226928
R10522 x9.A1.n65 x9.A1.n64 0.0226928
R10523 x9.A1.n55 x9.A1.n54 0.0226928
R10524 x9.A1.n47 x9.A1.n46 0.0226928
R10525 x9.A1.n37 x9.A1.n36 0.0226928
R10526 x9.A1.n30 x9.A1.n29 0.0226928
R10527 x9.A1.n98 x9.A1.n93 0.0125192
R10528 x9.A1.n114 x9.A1.n109 0.0125192
R10529 x9.A1.n130 x9.A1.n125 0.0125192
R10530 x9.A1.n80 x9.A1.n75 0.0125192
R10531 x9.A1.n62 x9.A1.n57 0.0125192
R10532 x9.A1.n44 x9.A1.n39 0.0125192
R10533 x9.A1.n27 x9.A1.n22 0.0125192
R10534 x9.A1.n99 x9.A1.n98 0.0109043
R10535 x9.A1.n115 x9.A1.n114 0.0109043
R10536 x9.A1.n131 x9.A1.n130 0.0109043
R10537 x9.A1.n81 x9.A1.n80 0.0109043
R10538 x9.A1.n63 x9.A1.n62 0.0109043
R10539 x9.A1.n45 x9.A1.n44 0.0109043
R10540 x9.A1.n28 x9.A1.n27 0.0109043
R10541 VSS_SW_b[3].n4 VSS_SW_b[3].n3 641.827
R10542 VSS_SW_b[3] VSS_SW_b[3].t1 422.656
R10543 VSS_SW_b[3].t1 VSS_SW_b[3].n5 121.231
R10544 VSS_SW_b[3].n2 VSS_SW_b[3].t0 117.424
R10545 VSS_SW_b[3].n3 VSS_SW_b[3].n2 77.418
R10546 VSS_SW_b[3].n6 VSS_SW_b[3] 11.3827
R10547 VSS_SW_b[3].n5 VSS_SW_b[3].n0 9.15497
R10548 VSS_SW_b[3].n5 VSS_SW_b[3].n4 7.57742
R10549 VSS_SW_b[3].n2 VSS_SW_b[3] 5.61454
R10550 VSS_SW_b[3].n8 VSS_SW_b[3].n6 2.47092
R10551 VSS_SW_b[3].n3 VSS_SW_b[3] 2.02155
R10552 VSS_SW_b[3].n12 VSS_SW_b[3] 1.6999
R10553 VSS_SW_b[3].n6 VSS_SW_b[3].n0 1.50964
R10554 VSS_SW_b[3].n10 VSS_SW_b[3].n9 1.5083
R10555 VSS_SW_b[3] VSS_SW_b[3].n12 1.3731
R10556 VSS_SW_b[3] VSS_SW_b[3].n1 1.34787
R10557 VSS_SW_b[3].n1 VSS_SW_b[3].n0 0.449623
R10558 VSS_SW_b[3].n12 VSS_SW_b[3].n11 0.0501381
R10559 VSS_SW_b[3].n11 VSS_SW_b[3].n10 0.0260996
R10560 VSS_SW_b[3].n8 VSS_SW_b[3].n7 0.0219844
R10561 VSS_SW_b[3].n9 VSS_SW_b[3].n8 0.00489987
R10562 D[6].n0 D[6].t2 331.51
R10563 D[6].n5 D[6].t3 331.51
R10564 D[6].n0 D[6].t1 209.403
R10565 D[6].n5 D[6].t0 209.403
R10566 D[6].n1 D[6].n0 76.0005
R10567 D[6].n6 D[6].n5 76.0005
R10568 D[6].n3 D[6].n2 14.0187
R10569 D[6].n2 D[6].n1 8.11757
R10570 D[6].n4 D[6] 7.49318
R10571 D[6].n4 D[6].n3 6.97656
R10572 D[6].n1 D[6] 2.02977
R10573 D[6] D[6].n6 2.02977
R10574 D[6].n6 D[6].n4 1.09318
R10575 D[6].n2 D[6] 0.468793
R10576 D[6].n3 D[6] 0.0519212
R10577 check[1] check[1].n3 363.457
R10578 check[1] check[1].n1 352.005
R10579 check[1].n0 check[1].t3 329.762
R10580 check[1].n7 check[1].t1 328.118
R10581 check[1].n3 check[1].t4 272.062
R10582 check[1].n1 check[1].t6 272.062
R10583 check[1].n3 check[1].t5 206.19
R10584 check[1].n1 check[1].t7 206.19
R10585 check[1].n0 check[1].t2 147.188
R10586 check[1].n6 check[1].t0 141.374
R10587 check[1].n16 check[1] 28.0657
R10588 check[1].n4 check[1] 15.1584
R10589 check[1].n8 check[1].n7 9.3005
R10590 check[1].n7 check[1].n6 8.19823
R10591 check[1] check[1].n0 7.17927
R10592 check[1].n5 check[1].n4 5.05313
R10593 check[1].n10 check[1].n9 5.05313
R10594 check[1].n16 check[1].n15 4.77557
R10595 check[1].n9 check[1] 4.37945
R10596 check[1].n13 check[1].n10 3.03311
R10597 check[1] check[1].n16 1.31653
R10598 check[1].n8 check[1].n5 0.674184
R10599 check[1].n10 check[1].n8 0.674184
R10600 check[1].n13 check[1].n12 0.166613
R10601 check[1].n12 check[1] 0.0531797
R10602 check[1].n14 check[1].n13 0.0352222
R10603 check[1].n15 check[1].n14 0.0167037
R10604 check[1].n12 check[1].n11 0.00485575
R10605 check[1].n13 check[1].n2 0.00331272
R10606 D[2].n0 D[2].t3 331.51
R10607 D[2].n5 D[2].t0 331.51
R10608 D[2].n0 D[2].t2 209.403
R10609 D[2].n5 D[2].t1 209.403
R10610 D[2].n1 D[2].n0 76.0005
R10611 D[2].n6 D[2].n5 76.0005
R10612 D[2].n3 D[2].n2 14.0187
R10613 D[2].n2 D[2].n1 8.27367
R10614 D[2].n4 D[2] 7.49318
R10615 D[2].n4 D[2].n3 6.97953
R10616 D[2].n1 D[2] 2.02977
R10617 D[2] D[2].n6 2.02977
R10618 D[2].n6 D[2].n4 1.09318
R10619 D[2].n2 D[2] 0.312695
R10620 D[2].n3 D[2] 0.051922
R10621 VDD_SW_b[6].n3 VDD_SW_b[6].t0 117.424
R10622 VDD_SW_b[6].n0 VDD_SW_b[6].t1 100.715
R10623 VDD_SW_b[6].n4 VDD_SW_b[6].n3 76.5198
R10624 VDD_SW_b[6].n0 VDD_SW_b[6] 10.2646
R10625 VDD_SW_b[6].n6 VDD_SW_b[6].n4 9.3005
R10626 VDD_SW_b[6].n3 VDD_SW_b[6] 5.61454
R10627 VDD_SW_b[6].n6 VDD_SW_b[6].n2 4.5005
R10628 VDD_SW_b[6].n1 VDD_SW_b[6].n0 3.75113
R10629 VDD_SW_b[6].n10 VDD_SW_b[6] 3.66121
R10630 VDD_SW_b[6] VDD_SW_b[6].n10 2.95723
R10631 VDD_SW_b[6].n4 VDD_SW_b[6] 2.9198
R10632 VDD_SW_b[6].n8 VDD_SW_b[6].n7 1.50505
R10633 VDD_SW_b[6].n2 VDD_SW_b[6].n1 0.449623
R10634 VDD_SW_b[6] VDD_SW_b[6].n2 0.449623
R10635 VDD_SW_b[6].n10 VDD_SW_b[6].n9 0.0501381
R10636 VDD_SW_b[6].n9 VDD_SW_b[6].n8 0.0260996
R10637 VDD_SW_b[6].n6 VDD_SW_b[6].n5 0.0122188
R10638 VDD_SW_b[6].n7 VDD_SW_b[6].n6 0.00814977
R10639 D[3].n0 D[3].t0 331.51
R10640 D[3].n5 D[3].t1 331.51
R10641 D[3].n0 D[3].t3 209.403
R10642 D[3].n5 D[3].t2 209.403
R10643 D[3].n1 D[3].n0 76.0005
R10644 D[3].n6 D[3].n5 76.0005
R10645 D[3].n3 D[3].n2 14.0217
R10646 D[3].n2 D[3].n1 8.11757
R10647 D[3].n4 D[3] 7.49318
R10648 D[3].n4 D[3].n3 6.97953
R10649 D[3].n1 D[3] 2.02977
R10650 D[3] D[3].n6 2.02977
R10651 D[3].n6 D[3].n4 1.09318
R10652 D[3].n2 D[3] 0.468793
R10653 D[3].n3 D[3] 0.051922
R10654 VSS_SW_b[2].n4 VSS_SW_b[2].n3 638.038
R10655 VSS_SW_b[2] VSS_SW_b[2].t1 422.656
R10656 VSS_SW_b[2].t1 VSS_SW_b[2].n5 117.442
R10657 VSS_SW_b[2].n2 VSS_SW_b[2].t0 117.424
R10658 VSS_SW_b[2].n3 VSS_SW_b[2].n2 77.6426
R10659 VSS_SW_b[2].n5 VSS_SW_b[2].n4 11.3659
R10660 VSS_SW_b[2].n6 VSS_SW_b[2] 11.1582
R10661 VSS_SW_b[2].n5 VSS_SW_b[2].n0 9.15497
R10662 VSS_SW_b[2].n2 VSS_SW_b[2] 5.61454
R10663 VSS_SW_b[2].n8 VSS_SW_b[2].n6 2.47092
R10664 VSS_SW_b[2].n3 VSS_SW_b[2] 1.79699
R10665 VSS_SW_b[2].n12 VSS_SW_b[2] 1.70288
R10666 VSS_SW_b[2].n6 VSS_SW_b[2].n0 1.50964
R10667 VSS_SW_b[2].n10 VSS_SW_b[2].n9 1.5083
R10668 VSS_SW_b[2] VSS_SW_b[2].n12 1.3755
R10669 VSS_SW_b[2] VSS_SW_b[2].n1 1.34787
R10670 VSS_SW_b[2].n1 VSS_SW_b[2].n0 0.674184
R10671 VSS_SW_b[2].n12 VSS_SW_b[2].n11 0.0501381
R10672 VSS_SW_b[2].n11 VSS_SW_b[2].n10 0.0260996
R10673 VSS_SW_b[2].n8 VSS_SW_b[2].n7 0.0219844
R10674 VSS_SW_b[2].n9 VSS_SW_b[2].n8 0.00489987
R10675 check[4] check[4].n3 363.457
R10676 check[4] check[4].n1 352.005
R10677 check[4].n0 check[4].t7 328.911
R10678 check[4].n7 check[4].t5 328.118
R10679 check[4].n3 check[4].t0 272.062
R10680 check[4].n1 check[4].t2 272.062
R10681 check[4].n3 check[4].t1 206.19
R10682 check[4].n1 check[4].t3 206.19
R10683 check[4].n0 check[4].t6 148.035
R10684 check[4].n6 check[4].t4 141.374
R10685 check[4].n16 check[4] 28.0656
R10686 check[4].n4 check[4] 15.1584
R10687 check[4].n8 check[4].n7 9.3005
R10688 check[4].n7 check[4].n6 8.19823
R10689 check[4] check[4].n0 7.14463
R10690 check[4].n10 check[4].n9 5.38997
R10691 check[4].n16 check[4].n15 5.06786
R10692 check[4].n5 check[4].n4 5.05313
R10693 check[4].n9 check[4] 4.37945
R10694 check[4].n13 check[4].n10 3.03311
R10695 check[4] check[4].n16 1.31656
R10696 check[4].n8 check[4].n5 0.674184
R10697 check[4].n10 check[4].n8 0.337342
R10698 check[4].n13 check[4].n12 0.166613
R10699 check[4].n12 check[4] 0.0531797
R10700 check[4].n14 check[4].n13 0.037537
R10701 check[4].n15 check[4].n14 0.0143889
R10702 check[4].n12 check[4].n11 0.00485575
R10703 check[4].n13 check[4].n2 0.00215636
R10704 VDD_SW[4].n8 VDD_SW[4].t0 117.424
R10705 VDD_SW[4].n6 VDD_SW[4].t1 75.7697
R10706 VDD_SW[4].n7 VDD_SW[4].n6 73.0808
R10707 VDD_SW[4] VDD_SW[4].n8 67.6928
R10708 VDD_SW[4].n10 VDD_SW[4].n9 13.0467
R10709 VDD_SW[4].n8 VDD_SW[4] 6.64665
R10710 VDD_SW[4].n5 VDD_SW[4].n4 2.82795
R10711 VDD_SW[4] VDD_SW[4].n7 2.2023
R10712 VDD_SW[4] VDD_SW[4].n10 1.96973
R10713 VDD_SW[4].n9 VDD_SW[4] 1.72358
R10714 VDD_SW[4].n3 VDD_SW[4].n1 1.49691
R10715 VDD_SW[4].n1 VDD_SW[4] 0.0595299
R10716 VDD_SW[4].n1 VDD_SW[4].n0 0.0177811
R10717 VDD_SW[4].n7 VDD_SW[4].n5 0.0146776
R10718 VDD_SW[4].n3 VDD_SW[4].n2 0.0102656
R10719 VDD_SW[4].n4 VDD_SW[4].n3 0.00635152
R10720 D[7].n0 D[7].t1 331.51
R10721 D[7].n5 D[7].t3 331.51
R10722 D[7].n0 D[7].t2 209.403
R10723 D[7].n5 D[7].t0 209.403
R10724 D[7].n1 D[7].n0 76.0005
R10725 D[7].n6 D[7].n5 76.0005
R10726 D[7].n3 D[7].n2 14.0187
R10727 D[7].n2 D[7].n1 8.11757
R10728 D[7].n4 D[7] 7.49318
R10729 D[7].n4 D[7].n3 6.97656
R10730 D[7].n1 D[7] 2.02977
R10731 D[7] D[7].n6 2.02977
R10732 D[7].n6 D[7].n4 1.09318
R10733 D[7].n2 D[7] 0.468793
R10734 D[7].n3 D[7] 0.0519212
R10735 check[3] check[3].n3 363.457
R10736 check[3] check[3].n1 352.005
R10737 check[3].n7 check[3].t1 329.01
R10738 check[3].n0 check[3].t5 328.911
R10739 check[3].n3 check[3].t6 272.062
R10740 check[3].n1 check[3].t2 272.062
R10741 check[3].n3 check[3].t7 206.19
R10742 check[3].n1 check[3].t3 206.19
R10743 check[3].n0 check[3].t4 148.035
R10744 check[3].n6 check[3].t0 140.888
R10745 check[3].n16 check[3] 28.1395
R10746 check[3].n4 check[3] 15.1584
R10747 check[3].n8 check[3].n7 9.3005
R10748 check[3].n7 check[3].n6 7.71392
R10749 check[3] check[3].n0 7.14463
R10750 check[3].n10 check[3].n9 5.38997
R10751 check[3].n5 check[3].n4 5.05313
R10752 check[3].n16 check[3].n15 4.87033
R10753 check[3].n9 check[3] 4.37945
R10754 check[3].n13 check[3].n10 3.03311
R10755 check[3] check[3].n16 1.15253
R10756 check[3].n8 check[3].n5 0.674184
R10757 check[3].n10 check[3].n8 0.337342
R10758 check[3].n13 check[3].n12 0.166613
R10759 check[3].n12 check[3] 0.0531806
R10760 check[3].n14 check[3].n13 0.037537
R10761 check[3].n15 check[3].n14 0.0143889
R10762 check[3].n12 check[3].n11 0.00485575
R10763 check[3].n13 check[3].n2 0.00215636
R10764 check[0] check[0].n3 363.457
R10765 check[0] check[0].n1 352.005
R10766 check[0].n0 check[0].t3 329.762
R10767 check[0].n7 check[0].t5 329.01
R10768 check[0].n3 check[0].t0 272.062
R10769 check[0].n1 check[0].t6 272.062
R10770 check[0].n3 check[0].t1 206.19
R10771 check[0].n1 check[0].t7 206.19
R10772 check[0].n0 check[0].t2 147.188
R10773 check[0].n6 check[0].t4 140.888
R10774 check[0].n16 check[0] 28.1411
R10775 check[0].n4 check[0] 15.1584
R10776 check[0].n8 check[0].n7 9.3005
R10777 check[0].n7 check[0].n6 7.71392
R10778 check[0] check[0].n0 7.17927
R10779 check[0].n10 check[0].n9 5.38997
R10780 check[0].n5 check[0].n4 5.05313
R10781 check[0].n16 check[0].n15 4.81189
R10782 check[0].n9 check[0] 4.37945
R10783 check[0].n13 check[0].n10 3.03311
R10784 check[0] check[0].n16 1.15191
R10785 check[0].n8 check[0].n5 0.674184
R10786 check[0].n10 check[0].n8 0.337342
R10787 check[0].n13 check[0].n12 0.166613
R10788 check[0].n12 check[0] 0.0531806
R10789 check[0].n14 check[0].n13 0.037537
R10790 check[0].n15 check[0].n14 0.0143889
R10791 check[0].n12 check[0].n11 0.00485575
R10792 check[0].n13 check[0].n2 0.00215636
R10793 reset.n2 reset.t0 255.25
R10794 reset.n0 reset.t1 169.462
R10795 reset.n3 reset.n2 9.3005
R10796 reset.n1 reset.n0 5.70839
R10797 reset.n3 reset 5.61776
R10798 reset.n2 reset.n1 5.07418
R10799 reset.n5 reset.n4 1.69462
R10800 reset.n4 reset.n3 1.50638
R10801 reset reset.n5 0.376971
R10802 D[4].n0 D[4].t0 331.51
R10803 D[4].n5 D[4].t1 331.51
R10804 D[4].n0 D[4].t3 209.403
R10805 D[4].n5 D[4].t2 209.403
R10806 D[4].n1 D[4].n0 76.0005
R10807 D[4].n6 D[4].n5 76.0005
R10808 D[4].n3 D[4].n2 14.0157
R10809 D[4].n2 D[4].n1 8.27367
R10810 D[4].n4 D[4] 7.49318
R10811 D[4].n4 D[4].n3 6.97656
R10812 D[4].n1 D[4] 2.02977
R10813 D[4] D[4].n6 2.02977
R10814 D[4].n6 D[4].n4 1.09318
R10815 D[4].n2 D[4] 0.312695
R10816 D[4].n3 D[4] 0.0519212
R10817 VSS_SW_b[4].n4 VSS_SW_b[4].n3 641.827
R10818 VSS_SW_b[4] VSS_SW_b[4].t1 422.656
R10819 VSS_SW_b[4].t1 VSS_SW_b[4].n5 121.231
R10820 VSS_SW_b[4].n2 VSS_SW_b[4].t0 117.424
R10821 VSS_SW_b[4].n3 VSS_SW_b[4].n2 77.418
R10822 VSS_SW_b[4].n6 VSS_SW_b[4] 11.3827
R10823 VSS_SW_b[4].n5 VSS_SW_b[4].n0 9.15497
R10824 VSS_SW_b[4].n5 VSS_SW_b[4].n4 7.57742
R10825 VSS_SW_b[4].n2 VSS_SW_b[4] 5.61454
R10826 VSS_SW_b[4].n8 VSS_SW_b[4].n6 2.47092
R10827 VSS_SW_b[4].n3 VSS_SW_b[4] 2.02155
R10828 VSS_SW_b[4].n12 VSS_SW_b[4] 1.6999
R10829 VSS_SW_b[4].n6 VSS_SW_b[4].n0 1.50964
R10830 VSS_SW_b[4].n10 VSS_SW_b[4].n9 1.5083
R10831 VSS_SW_b[4] VSS_SW_b[4].n12 1.3731
R10832 VSS_SW_b[4] VSS_SW_b[4].n1 1.34787
R10833 VSS_SW_b[4].n1 VSS_SW_b[4].n0 0.449623
R10834 VSS_SW_b[4].n12 VSS_SW_b[4].n11 0.0501381
R10835 VSS_SW_b[4].n11 VSS_SW_b[4].n10 0.0260996
R10836 VSS_SW_b[4].n8 VSS_SW_b[4].n7 0.0219844
R10837 VSS_SW_b[4].n9 VSS_SW_b[4].n8 0.00489987
R10838 VDD_SW_b[1].n3 VDD_SW_b[1].t0 117.424
R10839 VDD_SW_b[1].n0 VDD_SW_b[1].t1 100.715
R10840 VDD_SW_b[1].n4 VDD_SW_b[1].n3 76.5198
R10841 VDD_SW_b[1].n0 VDD_SW_b[1] 10.2646
R10842 VDD_SW_b[1].n6 VDD_SW_b[1].n4 9.3005
R10843 VDD_SW_b[1].n3 VDD_SW_b[1] 5.61454
R10844 VDD_SW_b[1].n6 VDD_SW_b[1].n2 4.5005
R10845 VDD_SW_b[1].n1 VDD_SW_b[1].n0 3.75113
R10846 VDD_SW_b[1].n10 VDD_SW_b[1] 3.66419
R10847 VDD_SW_b[1] VDD_SW_b[1].n10 2.95963
R10848 VDD_SW_b[1].n4 VDD_SW_b[1] 2.9198
R10849 VDD_SW_b[1].n8 VDD_SW_b[1].n7 1.50505
R10850 VDD_SW_b[1] VDD_SW_b[1].n2 0.674184
R10851 VDD_SW_b[1].n2 VDD_SW_b[1].n1 0.225061
R10852 VDD_SW_b[1].n10 VDD_SW_b[1].n9 0.0501381
R10853 VDD_SW_b[1].n9 VDD_SW_b[1].n8 0.0260996
R10854 VDD_SW_b[1].n6 VDD_SW_b[1].n5 0.0122188
R10855 VDD_SW_b[1].n7 VDD_SW_b[1].n6 0.00814977
R10856 check[2] check[2].n3 363.457
R10857 check[2] check[2].n1 352.005
R10858 check[2].n0 check[2].t5 329.762
R10859 check[2].n7 check[2].t7 328.118
R10860 check[2].n3 check[2].t2 272.062
R10861 check[2].n1 check[2].t0 272.062
R10862 check[2].n3 check[2].t3 206.19
R10863 check[2].n1 check[2].t1 206.19
R10864 check[2].n0 check[2].t4 147.188
R10865 check[2].n6 check[2].t6 141.374
R10866 check[2].n16 check[2] 28.0653
R10867 check[2].n4 check[2] 15.1584
R10868 check[2].n8 check[2].n7 9.3005
R10869 check[2].n7 check[2].n6 8.19823
R10870 check[2] check[2].n0 7.17927
R10871 check[2].n10 check[2].n9 5.38997
R10872 check[2].n5 check[2].n4 5.05313
R10873 check[2].n16 check[2].n15 4.97041
R10874 check[2].n9 check[2] 4.37945
R10875 check[2].n13 check[2].n10 3.03311
R10876 check[2] check[2].n16 1.31669
R10877 check[2].n8 check[2].n5 0.674184
R10878 check[2].n10 check[2].n8 0.337342
R10879 check[2].n13 check[2].n12 0.166613
R10880 check[2].n12 check[2] 0.0531797
R10881 check[2].n14 check[2].n13 0.037537
R10882 check[2].n15 check[2].n14 0.0143889
R10883 check[2].n12 check[2].n11 0.00485575
R10884 check[2].n13 check[2].n2 0.00215636
R10885 VDD_SW[5].n8 VDD_SW[5].t0 117.424
R10886 VDD_SW[5].n6 VDD_SW[5].t1 75.7697
R10887 VDD_SW[5].n7 VDD_SW[5].n6 73.0808
R10888 VDD_SW[5] VDD_SW[5].n8 67.6928
R10889 VDD_SW[5].n10 VDD_SW[5].n9 13.0467
R10890 VDD_SW[5].n8 VDD_SW[5] 6.64665
R10891 VDD_SW[5].n5 VDD_SW[5].n4 2.82795
R10892 VDD_SW[5] VDD_SW[5].n7 2.2023
R10893 VDD_SW[5] VDD_SW[5].n10 1.96973
R10894 VDD_SW[5].n9 VDD_SW[5] 1.72358
R10895 VDD_SW[5].n3 VDD_SW[5].n1 1.49691
R10896 VDD_SW[5].n1 VDD_SW[5] 0.0595299
R10897 VDD_SW[5].n1 VDD_SW[5].n0 0.0177811
R10898 VDD_SW[5].n7 VDD_SW[5].n5 0.0146776
R10899 VDD_SW[5].n3 VDD_SW[5].n2 0.0102656
R10900 VDD_SW[5].n4 VDD_SW[5].n3 0.00635152
R10901 D[1].n0 D[1].t1 331.51
R10902 D[1].n5 D[1].t2 331.51
R10903 D[1].n0 D[1].t0 209.403
R10904 D[1].n5 D[1].t3 209.403
R10905 D[1].n1 D[1].n0 76.0005
R10906 D[1].n6 D[1].n5 76.0005
R10907 D[1].n3 D[1].n2 14.0217
R10908 D[1].n2 D[1].n1 8.11757
R10909 D[1].n4 D[1] 7.49318
R10910 D[1].n4 D[1].n3 6.97953
R10911 D[1].n1 D[1] 2.02977
R10912 D[1] D[1].n6 2.02977
R10913 D[1].n6 D[1].n4 1.09318
R10914 D[1].n2 D[1] 0.468793
R10915 D[1].n3 D[1] 0.051922
R10916 D[5].n0 D[5].t0 331.51
R10917 D[5].n5 D[5].t1 331.51
R10918 D[5].n0 D[5].t3 209.403
R10919 D[5].n5 D[5].t2 209.403
R10920 D[5].n1 D[5].n0 76.0005
R10921 D[5].n6 D[5].n5 76.0005
R10922 D[5].n3 D[5].n2 14.0187
R10923 D[5].n2 D[5].n1 8.27367
R10924 D[5].n4 D[5] 7.33709
R10925 D[5].n4 D[5].n3 6.97656
R10926 D[5].n1 D[5] 2.02977
R10927 D[5] D[5].n6 2.02977
R10928 D[5].n6 D[5].n4 1.24928
R10929 D[5].n2 D[5] 0.312695
R10930 D[5].n3 D[5] 0.051922
R10931 VDD_SW[6].n8 VDD_SW[6].t0 117.424
R10932 VDD_SW[6].n6 VDD_SW[6].t1 75.7697
R10933 VDD_SW[6].n7 VDD_SW[6].n6 73.0808
R10934 VDD_SW[6] VDD_SW[6].n8 67.6928
R10935 VDD_SW[6].n10 VDD_SW[6].n9 13.0467
R10936 VDD_SW[6].n8 VDD_SW[6] 6.64665
R10937 VDD_SW[6].n5 VDD_SW[6].n4 2.82795
R10938 VDD_SW[6] VDD_SW[6].n7 2.2023
R10939 VDD_SW[6] VDD_SW[6].n10 1.96973
R10940 VDD_SW[6].n9 VDD_SW[6] 1.72358
R10941 VDD_SW[6].n3 VDD_SW[6].n1 1.49691
R10942 VDD_SW[6].n1 VDD_SW[6] 0.0595299
R10943 VDD_SW[6].n1 VDD_SW[6].n0 0.0177811
R10944 VDD_SW[6].n7 VDD_SW[6].n5 0.0146776
R10945 VDD_SW[6].n3 VDD_SW[6].n2 0.0102656
R10946 VDD_SW[6].n4 VDD_SW[6].n3 0.00635152
R10947 VSS_SW_b[5].n4 VSS_SW_b[5].n3 641.827
R10948 VSS_SW_b[5] VSS_SW_b[5].t1 422.656
R10949 VSS_SW_b[5].t1 VSS_SW_b[5].n5 121.231
R10950 VSS_SW_b[5].n2 VSS_SW_b[5].t0 117.424
R10951 VSS_SW_b[5].n3 VSS_SW_b[5].n2 77.418
R10952 VSS_SW_b[5].n6 VSS_SW_b[5] 11.3827
R10953 VSS_SW_b[5].n5 VSS_SW_b[5].n0 9.15497
R10954 VSS_SW_b[5].n5 VSS_SW_b[5].n4 7.57742
R10955 VSS_SW_b[5].n2 VSS_SW_b[5] 5.61454
R10956 VSS_SW_b[5].n8 VSS_SW_b[5].n6 2.47092
R10957 VSS_SW_b[5].n3 VSS_SW_b[5] 2.02155
R10958 VSS_SW_b[5].n12 VSS_SW_b[5] 1.6999
R10959 VSS_SW_b[5].n6 VSS_SW_b[5].n0 1.50964
R10960 VSS_SW_b[5].n10 VSS_SW_b[5].n9 1.5083
R10961 VSS_SW_b[5] VSS_SW_b[5].n12 1.3731
R10962 VSS_SW_b[5] VSS_SW_b[5].n1 1.34787
R10963 VSS_SW_b[5].n1 VSS_SW_b[5].n0 0.449623
R10964 VSS_SW_b[5].n12 VSS_SW_b[5].n11 0.0501381
R10965 VSS_SW_b[5].n11 VSS_SW_b[5].n10 0.0260996
R10966 VSS_SW_b[5].n8 VSS_SW_b[5].n7 0.0219844
R10967 VSS_SW_b[5].n9 VSS_SW_b[5].n8 0.00489987
R10968 VSS_SW_b[7].n4 VSS_SW_b[7].n3 641.827
R10969 VSS_SW_b[7] VSS_SW_b[7].t1 422.656
R10970 VSS_SW_b[7].t1 VSS_SW_b[7].n5 121.231
R10971 VSS_SW_b[7].n2 VSS_SW_b[7].t0 117.424
R10972 VSS_SW_b[7].n3 VSS_SW_b[7].n2 77.418
R10973 VSS_SW_b[7].n6 VSS_SW_b[7] 11.3827
R10974 VSS_SW_b[7].n5 VSS_SW_b[7].n0 9.15497
R10975 VSS_SW_b[7].n5 VSS_SW_b[7].n4 7.57742
R10976 VSS_SW_b[7].n2 VSS_SW_b[7] 5.61454
R10977 VSS_SW_b[7].n8 VSS_SW_b[7].n6 2.47092
R10978 VSS_SW_b[7].n3 VSS_SW_b[7] 2.02155
R10979 VSS_SW_b[7].n12 VSS_SW_b[7] 1.6999
R10980 VSS_SW_b[7].n6 VSS_SW_b[7].n0 1.50964
R10981 VSS_SW_b[7].n10 VSS_SW_b[7].n9 1.5083
R10982 VSS_SW_b[7] VSS_SW_b[7].n12 1.3731
R10983 VSS_SW_b[7] VSS_SW_b[7].n1 1.34787
R10984 VSS_SW_b[7].n1 VSS_SW_b[7].n0 0.449623
R10985 VSS_SW_b[7].n12 VSS_SW_b[7].n11 0.0501381
R10986 VSS_SW_b[7].n11 VSS_SW_b[7].n10 0.0260996
R10987 VSS_SW_b[7].n8 VSS_SW_b[7].n7 0.0219844
R10988 VSS_SW_b[7].n9 VSS_SW_b[7].n8 0.00489987
R10989 VDD_SW[7].n8 VDD_SW[7].t0 117.424
R10990 VDD_SW[7].n6 VDD_SW[7].t1 75.7697
R10991 VDD_SW[7].n7 VDD_SW[7].n6 73.0808
R10992 VDD_SW[7] VDD_SW[7].n8 67.6928
R10993 VDD_SW[7].n10 VDD_SW[7].n9 13.0467
R10994 VDD_SW[7].n8 VDD_SW[7] 6.64665
R10995 VDD_SW[7].n5 VDD_SW[7].n4 2.82795
R10996 VDD_SW[7] VDD_SW[7].n7 2.2023
R10997 VDD_SW[7] VDD_SW[7].n10 1.96973
R10998 VDD_SW[7].n9 VDD_SW[7] 1.72358
R10999 VDD_SW[7].n3 VDD_SW[7].n1 1.49691
R11000 VDD_SW[7].n1 VDD_SW[7] 0.0595299
R11001 VDD_SW[7].n1 VDD_SW[7].n0 0.0177811
R11002 VDD_SW[7].n7 VDD_SW[7].n5 0.0146776
R11003 VDD_SW[7].n3 VDD_SW[7].n2 0.0102656
R11004 VDD_SW[7].n4 VDD_SW[7].n3 0.00635152
R11005 VDD_SW_b[5].n3 VDD_SW_b[5].t0 117.424
R11006 VDD_SW_b[5].n0 VDD_SW_b[5].t1 100.715
R11007 VDD_SW_b[5].n4 VDD_SW_b[5].n3 76.5198
R11008 VDD_SW_b[5].n0 VDD_SW_b[5] 10.2646
R11009 VDD_SW_b[5].n6 VDD_SW_b[5].n4 9.3005
R11010 VDD_SW_b[5].n3 VDD_SW_b[5] 5.61454
R11011 VDD_SW_b[5].n6 VDD_SW_b[5].n2 4.5005
R11012 VDD_SW_b[5].n1 VDD_SW_b[5].n0 3.75113
R11013 VDD_SW_b[5].n10 VDD_SW_b[5] 3.66121
R11014 VDD_SW_b[5] VDD_SW_b[5].n10 2.95723
R11015 VDD_SW_b[5].n4 VDD_SW_b[5] 2.9198
R11016 VDD_SW_b[5].n8 VDD_SW_b[5].n7 1.5044
R11017 VDD_SW_b[5].n2 VDD_SW_b[5].n1 0.449623
R11018 VDD_SW_b[5] VDD_SW_b[5].n2 0.449623
R11019 VDD_SW_b[5].n10 VDD_SW_b[5].n9 0.0501381
R11020 VDD_SW_b[5].n9 VDD_SW_b[5].n8 0.0260996
R11021 VDD_SW_b[5].n6 VDD_SW_b[5].n5 0.0102656
R11022 VDD_SW_b[5].n7 VDD_SW_b[5].n6 0.00879975
R11023 VDD_SW[1].n8 VDD_SW[1].t0 117.424
R11024 VDD_SW[1].n6 VDD_SW[1].t1 75.7697
R11025 VDD_SW[1].n7 VDD_SW[1].n6 73.0808
R11026 VDD_SW[1] VDD_SW[1].n8 67.6928
R11027 VDD_SW[1].n10 VDD_SW[1].n9 13.0467
R11028 VDD_SW[1].n8 VDD_SW[1] 6.64665
R11029 VDD_SW[1].n5 VDD_SW[1].n4 2.82795
R11030 VDD_SW[1] VDD_SW[1].n7 2.2023
R11031 VDD_SW[1] VDD_SW[1].n10 1.96973
R11032 VDD_SW[1].n9 VDD_SW[1] 1.72358
R11033 VDD_SW[1].n3 VDD_SW[1].n1 1.49691
R11034 VDD_SW[1].n1 VDD_SW[1] 0.0595299
R11035 VDD_SW[1].n1 VDD_SW[1].n0 0.0177811
R11036 VDD_SW[1].n7 VDD_SW[1].n5 0.0146776
R11037 VDD_SW[1].n3 VDD_SW[1].n2 0.0102656
R11038 VDD_SW[1].n4 VDD_SW[1].n3 0.00635152
R11039 VSS_SW[3].n3 VSS_SW[3].n2 585
R11040 VSS_SW[3].n1 VSS_SW[3].t1 417.519
R11041 VSS_SW[3].n0 VSS_SW[3].t0 117.424
R11042 VSS_SW[3].n4 VSS_SW[3].n3 73.4178
R11043 VSS_SW[3].n3 VSS_SW[3].t1 68.1928
R11044 VSS_SW[3] VSS_SW[3].n0 67.6928
R11045 VSS_SW[3].n2 VSS_SW[3].n1 12.5543
R11046 VSS_SW[3].n0 VSS_SW[3] 6.64665
R11047 VSS_SW[3] VSS_SW[3].n4 3.039
R11048 VSS_SW[3].n2 VSS_SW[3] 2.46204
R11049 VSS_SW[3].n4 VSS_SW[3] 1.72358
R11050 VSS_SW[3].n1 VSS_SW[3] 1.72358
R11051 VSS_SW[5].n3 VSS_SW[5].n0 585
R11052 VSS_SW[5].n2 VSS_SW[5].t1 417.519
R11053 VSS_SW[5].n1 VSS_SW[5].t0 117.424
R11054 VSS_SW[5].n4 VSS_SW[5].n0 73.2739
R11055 VSS_SW[5].t1 VSS_SW[5].n0 71.9813
R11056 VSS_SW[5] VSS_SW[5].n1 67.6928
R11057 VSS_SW[5].n3 VSS_SW[5].n2 12.8005
R11058 VSS_SW[5].n1 VSS_SW[5] 6.64665
R11059 VSS_SW[5] VSS_SW[5].n4 3.04482
R11060 VSS_SW[5] VSS_SW[5].n3 2.21588
R11061 VSS_SW[5].n4 VSS_SW[5] 1.9648
R11062 VSS_SW[5].n2 VSS_SW[5] 1.72358
R11063 check[6] check[6].n3 363.457
R11064 check[6] check[6].n1 352.005
R11065 check[6].n7 check[6].t5 329.01
R11066 check[6].n0 check[6].t7 328.911
R11067 check[6].n3 check[6].t0 272.062
R11068 check[6].n1 check[6].t2 272.062
R11069 check[6].n3 check[6].t1 206.19
R11070 check[6].n1 check[6].t3 206.19
R11071 check[6].n0 check[6].t6 148.035
R11072 check[6].n6 check[6].t4 140.888
R11073 check[6].n16 check[6] 28.1391
R11074 check[6].n4 check[6] 15.1584
R11075 check[6].n8 check[6].n7 9.3005
R11076 check[6].n7 check[6].n6 7.71392
R11077 check[6] check[6].n0 7.14463
R11078 check[6].n10 check[6].n9 5.38997
R11079 check[6].n5 check[6].n4 5.05313
R11080 check[6].n16 check[6].n15 4.76728
R11081 check[6].n9 check[6] 4.37945
R11082 check[6].n13 check[6].n10 3.03311
R11083 check[6] check[6].n16 1.15267
R11084 check[6].n8 check[6].n5 0.674184
R11085 check[6].n10 check[6].n8 0.337342
R11086 check[6].n13 check[6].n12 0.166672
R11087 check[6].n12 check[6] 0.0532291
R11088 check[6].n14 check[6].n13 0.037537
R11089 check[6].n15 check[6].n14 0.0143889
R11090 check[6].n12 check[6].n11 0.00481511
R11091 check[6].n13 check[6].n2 0.00215119
R11092 ready.n0 ready.t0 259.723
R11093 ready.n0 ready.t1 175.108
R11094 ready.n1 ready 19.9175
R11095 ready.n1 ready.n0 8.27037
R11096 ready ready.n1 1.16637
R11097 VDD_SW[2].n8 VDD_SW[2].t0 117.424
R11098 VDD_SW[2].n6 VDD_SW[2].t1 75.7697
R11099 VDD_SW[2].n7 VDD_SW[2].n6 73.0808
R11100 VDD_SW[2] VDD_SW[2].n8 67.6928
R11101 VDD_SW[2].n10 VDD_SW[2].n9 13.0467
R11102 VDD_SW[2].n8 VDD_SW[2] 6.64665
R11103 VDD_SW[2].n5 VDD_SW[2].n4 2.82795
R11104 VDD_SW[2] VDD_SW[2].n7 2.2023
R11105 VDD_SW[2] VDD_SW[2].n10 1.96973
R11106 VDD_SW[2].n9 VDD_SW[2] 1.72358
R11107 VDD_SW[2].n3 VDD_SW[2].n1 1.49691
R11108 VDD_SW[2].n1 VDD_SW[2] 0.0595299
R11109 VDD_SW[2].n1 VDD_SW[2].n0 0.0177811
R11110 VDD_SW[2].n7 VDD_SW[2].n5 0.0146776
R11111 VDD_SW[2].n3 VDD_SW[2].n2 0.0102656
R11112 VDD_SW[2].n4 VDD_SW[2].n3 0.00635152
R11113 check[5] check[5].n3 363.457
R11114 check[5] check[5].n1 352.005
R11115 check[5].n0 check[5].t1 328.911
R11116 check[5].n7 check[5].t3 328.118
R11117 check[5].n3 check[5].t6 272.062
R11118 check[5].n1 check[5].t4 272.062
R11119 check[5].n3 check[5].t7 206.19
R11120 check[5].n1 check[5].t5 206.19
R11121 check[5].n0 check[5].t0 148.035
R11122 check[5].n6 check[5].t2 141.374
R11123 check[5].n16 check[5] 28.1388
R11124 check[5].n4 check[5] 15.1584
R11125 check[5].n8 check[5].n7 9.3005
R11126 check[5].n7 check[5].n6 8.19823
R11127 check[5] check[5].n0 7.14463
R11128 check[5].n10 check[5].n9 5.38997
R11129 check[5].n5 check[5].n4 5.05313
R11130 check[5].n16 check[5].n15 4.76129
R11131 check[5].n9 check[5] 4.37945
R11132 check[5].n13 check[5].n10 3.03311
R11133 check[5] check[5].n16 1.15277
R11134 check[5].n8 check[5].n5 0.674184
R11135 check[5].n10 check[5].n8 0.337342
R11136 check[5].n13 check[5].n12 0.166672
R11137 check[5].n12 check[5] 0.0532282
R11138 check[5].n14 check[5].n13 0.037537
R11139 check[5].n15 check[5].n14 0.0143889
R11140 check[5].n12 check[5].n11 0.00481511
R11141 check[5].n13 check[5].n2 0.00215119
R11142 VSS_SW[4].n3 VSS_SW[4].n0 585
R11143 VSS_SW[4].n2 VSS_SW[4].t1 417.519
R11144 VSS_SW[4].n1 VSS_SW[4].t0 117.424
R11145 VSS_SW[4].n4 VSS_SW[4].n0 73.2739
R11146 VSS_SW[4].t1 VSS_SW[4].n0 71.9813
R11147 VSS_SW[4] VSS_SW[4].n1 67.6928
R11148 VSS_SW[4].n3 VSS_SW[4].n2 12.8005
R11149 VSS_SW[4].n1 VSS_SW[4] 6.64665
R11150 VSS_SW[4] VSS_SW[4].n4 3.04482
R11151 VSS_SW[4] VSS_SW[4].n3 2.21588
R11152 VSS_SW[4].n4 VSS_SW[4] 1.9648
R11153 VSS_SW[4].n2 VSS_SW[4] 1.72358
R11154 VSS_SW[6].n3 VSS_SW[6].n0 585
R11155 VSS_SW[6].n2 VSS_SW[6].t1 417.519
R11156 VSS_SW[6].n1 VSS_SW[6].t0 117.424
R11157 VSS_SW[6].n4 VSS_SW[6].n0 73.2739
R11158 VSS_SW[6].t1 VSS_SW[6].n0 71.9813
R11159 VSS_SW[6] VSS_SW[6].n1 67.6928
R11160 VSS_SW[6].n3 VSS_SW[6].n2 12.8005
R11161 VSS_SW[6].n1 VSS_SW[6] 6.64665
R11162 VSS_SW[6] VSS_SW[6].n4 3.04482
R11163 VSS_SW[6] VSS_SW[6].n3 2.21588
R11164 VSS_SW[6].n4 VSS_SW[6] 1.9648
R11165 VSS_SW[6].n2 VSS_SW[6] 1.72358
R11166 VDD_SW_b[7].n3 VDD_SW_b[7].t0 117.424
R11167 VDD_SW_b[7].n0 VDD_SW_b[7].t1 102.686
R11168 VDD_SW_b[7].n4 VDD_SW_b[7].n3 76.2952
R11169 VDD_SW_b[7].n0 VDD_SW_b[7] 10.3552
R11170 VDD_SW_b[7].n6 VDD_SW_b[7].n4 9.3005
R11171 VDD_SW_b[7].n3 VDD_SW_b[7] 5.61454
R11172 VDD_SW_b[7].n6 VDD_SW_b[7].n2 4.5005
R11173 VDD_SW_b[7].n1 VDD_SW_b[7].n0 3.87653
R11174 VDD_SW_b[7].n10 VDD_SW_b[7] 3.65824
R11175 VDD_SW_b[7].n4 VDD_SW_b[7] 3.14436
R11176 VDD_SW_b[7] VDD_SW_b[7].n10 2.95483
R11177 VDD_SW_b[7].n8 VDD_SW_b[7].n7 1.50505
R11178 VDD_SW_b[7].n2 VDD_SW_b[7].n1 0.449623
R11179 VDD_SW_b[7] VDD_SW_b[7].n2 0.225061
R11180 VDD_SW_b[7].n10 VDD_SW_b[7].n9 0.0501381
R11181 VDD_SW_b[7].n9 VDD_SW_b[7].n8 0.0260996
R11182 VDD_SW_b[7].n6 VDD_SW_b[7].n5 0.0122188
R11183 VDD_SW_b[7].n7 VDD_SW_b[7].n6 0.00814977
R11184 VDD_SW_b[2].n3 VDD_SW_b[2].t0 117.424
R11185 VDD_SW_b[2].n0 VDD_SW_b[2].t1 102.686
R11186 VDD_SW_b[2].n4 VDD_SW_b[2].n3 76.2952
R11187 VDD_SW_b[2].n0 VDD_SW_b[2] 10.3552
R11188 VDD_SW_b[2].n6 VDD_SW_b[2].n4 9.3005
R11189 VDD_SW_b[2].n3 VDD_SW_b[2] 5.61454
R11190 VDD_SW_b[2].n6 VDD_SW_b[2].n2 4.5005
R11191 VDD_SW_b[2].n1 VDD_SW_b[2].n0 3.87653
R11192 VDD_SW_b[2].n10 VDD_SW_b[2] 3.65824
R11193 VDD_SW_b[2].n4 VDD_SW_b[2] 3.14436
R11194 VDD_SW_b[2] VDD_SW_b[2].n10 2.95483
R11195 VDD_SW_b[2].n8 VDD_SW_b[2].n7 1.50505
R11196 VDD_SW_b[2].n2 VDD_SW_b[2].n1 0.449623
R11197 VDD_SW_b[2] VDD_SW_b[2].n2 0.225061
R11198 VDD_SW_b[2].n10 VDD_SW_b[2].n9 0.0501381
R11199 VDD_SW_b[2].n9 VDD_SW_b[2].n8 0.0260996
R11200 VDD_SW_b[2].n6 VDD_SW_b[2].n5 0.0122188
R11201 VDD_SW_b[2].n7 VDD_SW_b[2].n6 0.00814977
R11202 VSS_SW[1].n3 VSS_SW[1].n0 585
R11203 VSS_SW[1].n2 VSS_SW[1].t1 417.519
R11204 VSS_SW[1].n1 VSS_SW[1].t0 117.424
R11205 VSS_SW[1].n4 VSS_SW[1].n0 73.2739
R11206 VSS_SW[1].t1 VSS_SW[1].n0 71.9813
R11207 VSS_SW[1] VSS_SW[1].n1 67.6928
R11208 VSS_SW[1].n3 VSS_SW[1].n2 12.8005
R11209 VSS_SW[1].n1 VSS_SW[1] 6.64665
R11210 VSS_SW[1] VSS_SW[1].n4 3.11587
R11211 VSS_SW[1] VSS_SW[1].n3 2.21588
R11212 VSS_SW[1].n4 VSS_SW[1] 1.9648
R11213 VSS_SW[1].n2 VSS_SW[1] 1.72358
R11214 VSS_SW[7].n3 VSS_SW[7].n0 585
R11215 VSS_SW[7].n2 VSS_SW[7].t1 417.519
R11216 VSS_SW[7].n1 VSS_SW[7].t0 117.424
R11217 VSS_SW[7].n4 VSS_SW[7].n0 73.2739
R11218 VSS_SW[7].t1 VSS_SW[7].n0 71.9813
R11219 VSS_SW[7] VSS_SW[7].n1 67.6928
R11220 VSS_SW[7].n3 VSS_SW[7].n2 12.8005
R11221 VSS_SW[7].n1 VSS_SW[7] 6.64665
R11222 VSS_SW[7] VSS_SW[7].n4 3.04482
R11223 VSS_SW[7] VSS_SW[7].n3 2.21588
R11224 VSS_SW[7].n4 VSS_SW[7] 1.9648
R11225 VSS_SW[7].n2 VSS_SW[7] 1.72358
R11226 VSS_SW_b[6].n4 VSS_SW_b[6].n3 641.827
R11227 VSS_SW_b[6] VSS_SW_b[6].t1 422.656
R11228 VSS_SW_b[6].t1 VSS_SW_b[6].n5 121.231
R11229 VSS_SW_b[6].n2 VSS_SW_b[6].t0 117.424
R11230 VSS_SW_b[6].n3 VSS_SW_b[6].n2 77.418
R11231 VSS_SW_b[6].n6 VSS_SW_b[6] 11.3827
R11232 VSS_SW_b[6].n5 VSS_SW_b[6].n0 9.15497
R11233 VSS_SW_b[6].n5 VSS_SW_b[6].n4 7.57742
R11234 VSS_SW_b[6].n2 VSS_SW_b[6] 5.61454
R11235 VSS_SW_b[6].n8 VSS_SW_b[6].n6 2.47092
R11236 VSS_SW_b[6].n3 VSS_SW_b[6] 2.02155
R11237 VSS_SW_b[6].n12 VSS_SW_b[6] 1.6999
R11238 VSS_SW_b[6].n6 VSS_SW_b[6].n0 1.50964
R11239 VSS_SW_b[6].n10 VSS_SW_b[6].n9 1.5083
R11240 VSS_SW_b[6] VSS_SW_b[6].n12 1.3731
R11241 VSS_SW_b[6] VSS_SW_b[6].n1 1.34787
R11242 VSS_SW_b[6].n1 VSS_SW_b[6].n0 0.449623
R11243 VSS_SW_b[6].n12 VSS_SW_b[6].n11 0.0501381
R11244 VSS_SW_b[6].n11 VSS_SW_b[6].n10 0.0260996
R11245 VSS_SW_b[6].n8 VSS_SW_b[6].n7 0.0219844
R11246 VSS_SW_b[6].n9 VSS_SW_b[6].n8 0.00489987
R11247 VDD_SW_b[3].n3 VDD_SW_b[3].t0 117.424
R11248 VDD_SW_b[3].n0 VDD_SW_b[3].t1 100.715
R11249 VDD_SW_b[3].n4 VDD_SW_b[3].n3 76.5198
R11250 VDD_SW_b[3].n0 VDD_SW_b[3] 10.2646
R11251 VDD_SW_b[3].n6 VDD_SW_b[3].n4 9.3005
R11252 VDD_SW_b[3].n3 VDD_SW_b[3] 5.61454
R11253 VDD_SW_b[3].n6 VDD_SW_b[3].n2 4.5005
R11254 VDD_SW_b[3].n1 VDD_SW_b[3].n0 3.75113
R11255 VDD_SW_b[3].n10 VDD_SW_b[3] 3.66121
R11256 VDD_SW_b[3] VDD_SW_b[3].n10 2.95723
R11257 VDD_SW_b[3].n4 VDD_SW_b[3] 2.9198
R11258 VDD_SW_b[3].n8 VDD_SW_b[3].n7 1.5044
R11259 VDD_SW_b[3].n2 VDD_SW_b[3].n1 0.449623
R11260 VDD_SW_b[3] VDD_SW_b[3].n2 0.449623
R11261 VDD_SW_b[3].n10 VDD_SW_b[3].n9 0.0501381
R11262 VDD_SW_b[3].n9 VDD_SW_b[3].n8 0.0260996
R11263 VDD_SW_b[3].n6 VDD_SW_b[3].n5 0.0102656
R11264 VDD_SW_b[3].n7 VDD_SW_b[3].n6 0.00879975
R11265 VSS_SW[2].n3 VSS_SW[2].n0 585
R11266 VSS_SW[2].n2 VSS_SW[2].t1 417.519
R11267 VSS_SW[2].n1 VSS_SW[2].t0 117.424
R11268 VSS_SW[2].n4 VSS_SW[2].n0 73.2739
R11269 VSS_SW[2].t1 VSS_SW[2].n0 71.9813
R11270 VSS_SW[2] VSS_SW[2].n1 67.6928
R11271 VSS_SW[2].n3 VSS_SW[2].n2 12.8005
R11272 VSS_SW[2].n1 VSS_SW[2] 6.64665
R11273 VSS_SW[2] VSS_SW[2].n4 3.11587
R11274 VSS_SW[2] VSS_SW[2].n3 2.21588
R11275 VSS_SW[2].n4 VSS_SW[2] 1.9648
R11276 VSS_SW[2].n2 VSS_SW[2] 1.72358
R11277 VSS_SW_b[1].n4 VSS_SW_b[1].n3 641.827
R11278 VSS_SW_b[1] VSS_SW_b[1].t1 422.656
R11279 VSS_SW_b[1].t1 VSS_SW_b[1].n5 121.231
R11280 VSS_SW_b[1].n2 VSS_SW_b[1].t0 117.424
R11281 VSS_SW_b[1].n3 VSS_SW_b[1].n2 77.418
R11282 VSS_SW_b[1].n6 VSS_SW_b[1] 11.3827
R11283 VSS_SW_b[1].n5 VSS_SW_b[1].n0 9.15497
R11284 VSS_SW_b[1].n5 VSS_SW_b[1].n4 7.57742
R11285 VSS_SW_b[1].n2 VSS_SW_b[1] 5.61454
R11286 VSS_SW_b[1].n8 VSS_SW_b[1].n6 2.47092
R11287 VSS_SW_b[1].n3 VSS_SW_b[1] 2.02155
R11288 VSS_SW_b[1].n12 VSS_SW_b[1] 1.6999
R11289 VSS_SW_b[1].n6 VSS_SW_b[1].n0 1.50964
R11290 VSS_SW_b[1].n10 VSS_SW_b[1].n9 1.5083
R11291 VSS_SW_b[1] VSS_SW_b[1].n12 1.3731
R11292 VSS_SW_b[1] VSS_SW_b[1].n1 1.34787
R11293 VSS_SW_b[1].n1 VSS_SW_b[1].n0 0.449623
R11294 VSS_SW_b[1].n12 VSS_SW_b[1].n11 0.0501381
R11295 VSS_SW_b[1].n11 VSS_SW_b[1].n10 0.0260996
R11296 VSS_SW_b[1].n8 VSS_SW_b[1].n7 0.0219844
R11297 VSS_SW_b[1].n9 VSS_SW_b[1].n8 0.00489987
R11298 VDD_SW_b[4].n3 VDD_SW_b[4].t0 117.424
R11299 VDD_SW_b[4].n0 VDD_SW_b[4].t1 100.715
R11300 VDD_SW_b[4].n4 VDD_SW_b[4].n3 76.5198
R11301 VDD_SW_b[4].n0 VDD_SW_b[4] 10.2646
R11302 VDD_SW_b[4].n6 VDD_SW_b[4].n4 9.3005
R11303 VDD_SW_b[4].n3 VDD_SW_b[4] 5.61454
R11304 VDD_SW_b[4].n6 VDD_SW_b[4].n2 4.5005
R11305 VDD_SW_b[4].n1 VDD_SW_b[4].n0 3.75113
R11306 VDD_SW_b[4].n10 VDD_SW_b[4] 3.66419
R11307 VDD_SW_b[4] VDD_SW_b[4].n10 2.95963
R11308 VDD_SW_b[4].n4 VDD_SW_b[4] 2.9198
R11309 VDD_SW_b[4].n8 VDD_SW_b[4].n7 1.50505
R11310 VDD_SW_b[4] VDD_SW_b[4].n2 0.674184
R11311 VDD_SW_b[4].n2 VDD_SW_b[4].n1 0.225061
R11312 VDD_SW_b[4].n10 VDD_SW_b[4].n9 0.0501381
R11313 VDD_SW_b[4].n9 VDD_SW_b[4].n8 0.0260996
R11314 VDD_SW_b[4].n6 VDD_SW_b[4].n5 0.0122188
R11315 VDD_SW_b[4].n7 VDD_SW_b[4].n6 0.00814977
R11316 VDD_SW[3].n8 VDD_SW[3].t0 117.424
R11317 VDD_SW[3].n6 VDD_SW[3].t1 75.7697
R11318 VDD_SW[3].n7 VDD_SW[3].n6 73.0808
R11319 VDD_SW[3] VDD_SW[3].n8 67.6928
R11320 VDD_SW[3].n10 VDD_SW[3].n9 13.0467
R11321 VDD_SW[3].n8 VDD_SW[3] 6.64665
R11322 VDD_SW[3].n5 VDD_SW[3].n4 2.82795
R11323 VDD_SW[3] VDD_SW[3].n7 2.2023
R11324 VDD_SW[3] VDD_SW[3].n10 1.96973
R11325 VDD_SW[3].n9 VDD_SW[3] 1.72358
R11326 VDD_SW[3].n3 VDD_SW[3].n1 1.49691
R11327 VDD_SW[3].n1 VDD_SW[3] 0.0595299
R11328 VDD_SW[3].n1 VDD_SW[3].n0 0.0177811
R11329 VDD_SW[3].n7 VDD_SW[3].n5 0.0146776
R11330 VDD_SW[3].n3 VDD_SW[3].n2 0.0102656
R11331 VDD_SW[3].n4 VDD_SW[3].n3 0.00635152
C0 a_2419_627# a_5165_627# 4.46e-21
C1 VDD a_2610_1642# 0.00177f
C2 a_3420_212# a_5504_106# 5.86e-20
C3 a_11546_1315# D[3] 0.0012f
C4 a_3421_n88# a_5271_n62# 4.56e-21
C5 VDD a_15721_n62# 0.0301f
C6 VSS_SW[2] a_12447_n62# 3.44e-19
C7 x2.X a_977_304# 0.00167f
C8 a_3039_601# a_2566_n88# 4.37e-19
C9 a_2585_627# a_2879_n62# 2.38e-19
C10 VDD a_9154_1315# 3.89e-19
C11 D[1] a_15293_601# 0.0189f
C12 a_14379_627# a_15767_895# 0.0321f
C13 VSS_SW_b[3] a_10937_n62# 5.35e-19
C14 a_11069_122# VSS_SW[2] 6.75e-20
C15 a_1672_909# VDD_SW[7] 2.12e-20
C16 check[1] x17.X 0.00967f
C17 a_10824_993# a_10596_212# 8.94e-21
C18 a_10509_601# a_10801_n88# 0.00251f
C19 a_10983_895# a_10597_n88# 6.35e-19
C20 x13.X D[4] 0.0996f
C21 D[3] a_10597_n88# 0.159f
C22 x12.X a_7557_627# 6.12e-19
C23 a_14430_90# a_14839_n62# 4.24e-20
C24 ready check[6] 0.0393f
C25 x9.A1 a_5725_601# 0.00103f
C26 check[3] a_8409_n88# 2.51e-19
C27 VSS_SW[3] a_9742_n88# 0.00683f
C28 a_3535_n62# a_3761_n62# 3.34e-19
C29 check[1] a_12134_n88# 5.26e-19
C30 x7.X a_1029_n88# 0.019f
C31 reset a_76_1467# 8.22e-19
C32 a_7252_1467# check[3] 0.318f
C33 check[6] a_1501_122# 6.43e-20
C34 VDD_SW[3] a_12433_993# 7.03e-20
C35 check[2] a_11123_627# 4.06e-19
C36 a_15243_909# VDD_SW_b[1] 3.6e-21
C37 check[4] VSS_SW_b[5] 3.18e-20
C38 check[3] x14.X 5.82e-19
C39 x15.X a_10288_106# 1.89e-20
C40 x9.A1 VDD_SW[4] 0.0329f
C41 VDD a_1757_1642# 0.115f
C42 x2.X a_10215_601# 0.2f
C43 a_15608_993# a_14839_n62# 3.59e-19
C44 a_14857_1289# a_14839_n62# 3.44e-19
C45 a_15293_601# a_15380_212# 6.03e-19
C46 check[5] VSS_SW[5] 1.43e-19
C47 a_14733_627# a_14526_n88# 3.32e-19
C48 x3.X a_647_601# 3.71e-19
C49 a_1028_212# a_3421_n88# 5.48e-21
C50 a_1029_n88# a_3420_212# 8.02e-22
C51 VDD a_2773_627# 0.109f
C52 a_305_2457# a_473_993# 4.56e-21
C53 a_29_2457# VSS_SW[7] 0.0221f
C54 D[7] a_2585_627# 7.7e-21
C55 a_5431_601# a_5341_993# 6.69e-20
C56 a_4977_627# a_5675_909# 0.00276f
C57 a_5725_601# a_6040_993# 0.13f
C58 a_5257_993# a_5165_627# 0.0369f
C59 x2.X a_16298_n62# 1.24e-19
C60 x18.X a_12153_627# 6.35e-20
C61 a_381_627# VSS_SW[7] 0.00595f
C62 VDD a_487_n62# 0.327f
C63 x30.A D[5] 1.01e-19
C64 a_4689_2457# a_5323_2457# 8.37e-20
C65 check[4] VDD_SW[5] 0.0039f
C66 x3.X x9.A1 9e-19
C67 a_2468_1467# VDD_SW[7] 0.00487f
C68 D[6] a_5812_212# 2.89e-20
C69 VSS_SW[2] a_13126_304# 1.97e-20
C70 a_12989_n88# a_13461_122# 0.15f
C71 a_12988_212# VSS_SW_b[2] 0.00119f
C72 VDD_SW[5] a_8432_993# 1.08e-20
C73 a_7203_627# a_8205_n88# 1.06e-19
C74 D[4] a_8204_212# 0.158f
C75 VSS_SW[4] a_8204_212# 5.9e-22
C76 VDD_SW_b[3] a_11514_n62# 0.0145f
C77 a_2419_627# a_2585_627# 0.786f
C78 a_4149_1315# D[6] 0.00195f
C79 a_9761_627# a_10359_627# 6.04e-20
C80 a_6199_895# VDD_SW_b[5] 0.129f
C81 D[5] a_7203_627# 9.94e-20
C82 a_4811_627# D[4] 1.19e-20
C83 ready D[7] 0.038f
C84 a_9595_627# a_10459_909# 2.46e-19
C85 x2.X VSS_SW_b[4] 0.0279f
C86 a_4811_627# VSS_SW[4] 4.66e-21
C87 a_5289_1289# x11.X 1.7e-20
C88 VDD a_10734_304# 0.0164f
C89 a_9595_627# VSS_SW[3] 0.0577f
C90 x3.X a_505_1289# 2.51e-20
C91 check[3] a_8591_895# 0.00271f
C92 a_27_627# VSS_SW_b[7] 1.08e-19
C93 a_8117_601# a_10509_601# 1.08e-20
C94 a_12036_1467# VDD_SW[3] 0.00487f
C95 D[7] a_1501_122# 0.00928f
C96 x9.A1 a_5271_n62# 1.54e-20
C97 a_4528_627# a_4811_627# 0.0011f
C98 VSS_SW_b[6] a_4137_n62# 6.94e-20
C99 a_4862_90# a_4958_n88# 0.0967f
C100 a_11987_627# a_12751_627# 0.00134f
C101 D[2] a_13300_993# 2.53e-19
C102 x9.A1 a_10073_1289# 0.104f
C103 x20.X a_16109_1315# 1.98e-19
C104 a_16024_909# VDD_SW[1] 2.12e-20
C105 x12.X a_4977_627# 6.35e-20
C106 x11.X a_4958_n88# 1.53e-21
C107 D[6] a_3732_993# 2.53e-19
C108 a_2419_627# a_3183_627# 0.00134f
C109 ready a_2419_627# 1.4e-20
C110 VDD a_5462_220# 0.0041f
C111 a_1757_1642# a_941_601# 7.12e-21
C112 VDD_SW[7] a_3039_601# 7.64e-20
C113 a_14999_601# a_14945_n62# 1.07e-20
C114 VDD a_12851_909# 0.00984f
C115 a_14933_627# VSS_SW[1] 3.79e-19
C116 a_1415_895# a_3648_993# 1.86e-21
C117 a_941_601# a_2773_627# 2.34e-20
C118 a_13936_1315# D[2] 0.0012f
C119 VDD_SW_b[2] a_14379_627# 5.97e-19
C120 a_13515_627# a_13323_627# 4.19e-20
C121 a_14096_627# VDD_SW[2] 0.0729f
C122 x9.X a_3112_106# 2.38e-20
C123 check[3] VDD_SW_b[4] 0.00218f
C124 a_10596_212# a_10734_304# 1.09e-19
C125 a_5165_627# a_4958_n88# 3.32e-19
C126 a_5725_601# a_5812_212# 6.03e-19
C127 a_6040_993# a_5271_n62# 3.59e-19
C128 VSS_SW[5] a_6285_122# 2.79e-21
C129 a_941_601# a_487_n62# 3.74e-20
C130 a_647_601# a_1028_212# 4.51e-19
C131 a_193_627# a_1029_n88# 1.27e-19
C132 a_473_993# a_720_106# 4.96e-20
C133 x7.X a_2470_90# 0.0273f
C134 a_13461_122# a_13906_n62# 0.0369f
C135 x9.A1 a_12988_212# 1.36e-20
C136 VDD_SW[6] a_3420_212# 4.31e-19
C137 a_3947_627# a_3625_n88# 7.32e-20
C138 a_12901_601# a_12988_212# 6.03e-19
C139 VDD D[4] 0.771f
C140 a_12341_627# a_12134_n88# 3.32e-19
C141 a_13216_993# a_12447_n62# 3.59e-19
C142 a_11704_627# D[2] 4.42e-19
C143 VDD VSS_SW[4] 0.526f
C144 a_11123_627# a_11987_627# 1.09e-19
C145 D[4] a_7649_993# 0.00874f
C146 a_7203_627# a_8117_601# 0.14f
C147 a_7649_993# VSS_SW[4] 0.00299f
C148 a_7350_n88# a_7663_n62# 0.245f
C149 a_6730_n62# a_6529_n62# 3.81e-19
C150 check[2] VSS_SW_b[3] 3.18e-20
C151 x14.X a_10215_601# 2.39e-20
C152 x9.A1 a_1028_212# 1.41e-20
C153 a_2468_1467# a_2610_1642# 0.00557f
C154 a_10073_1289# a_9742_n88# 5.67e-21
C155 a_1946_n62# a_3421_n88# 3.67e-21
C156 a_1166_304# VSS_SW_b[6] 9.89e-21
C157 VDD a_4528_627# 0.194f
C158 a_2470_90# a_3420_212# 2.02e-20
C159 x2.X a_7557_627# 0.0014f
C160 VDD_SW_b[5] a_5504_106# 5.26e-19
C161 a_14379_627# a_15072_106# 3.88e-21
C162 D[1] a_14839_n62# 0.00257f
C163 check[5] a_3648_993# 3.41e-19
C164 VDD_SW[4] a_9595_627# 0.0865f
C165 VDD_SW_b[7] a_174_n88# 3.21e-19
C166 a_9644_1467# a_10103_1642# 6.64e-19
C167 VDD a_1447_220# 0.00984f
C168 a_7681_1289# a_7896_106# 5.3e-21
C169 x30.A a_4860_1467# 6.58e-20
C170 x16.X a_12433_993# 1.03e-19
C171 ready a_4149_1642# 6.63e-21
C172 VDD_SW_b[6] a_3535_n62# 5.2e-19
C173 D[4] a_10596_212# 2.89e-20
C174 x27.A x9.A1 1.25e-19
C175 x2.X a_13375_895# 0.148f
C176 a_6760_1315# D[5] 0.0012f
C177 x2.X check[2] 0.148f
C178 D[4] a_8335_627# 6.12e-19
C179 x2.X a_5223_1315# 3.19e-19
C180 D[4] a_8921_304# 8.38e-19
C181 a_8409_n88# VSS_SW_b[4] 9.21e-19
C182 VDD_SW_b[1] a_15853_122# 0.00443f
C183 x20.X a_15853_122# 2.61e-19
C184 a_76_1467# a_78_90# 1e-19
C185 a_12038_90# VSS_SW[2] 0.082f
C186 a_7252_1467# VSS_SW_b[4] 2.13e-19
C187 a_5575_627# a_6147_627# 2.46e-21
C188 x2.X a_8140_n62# 3.68e-20
C189 check[0] VDD_SW[2] 4.27e-19
C190 x18.X a_14379_627# 0.236f
C191 a_10215_601# a_10680_909# 9.46e-19
C192 x17.X a_14096_627# 0.0338f
C193 x18.X VDD_SW_b[2] 7.23e-19
C194 a_13461_1642# x18.X 9.44e-21
C195 D[3] a_11313_304# 8.39e-19
C196 x9.X D[6] 0.0992f
C197 x2.X a_14887_1642# 2.63e-19
C198 x2.X a_15243_909# 0.00138f
C199 a_14526_n88# a_15381_n88# 0.0477f
C200 check[4] a_6753_1642# 0.00688f
C201 a_14839_n62# a_15380_212# 0.138f
C202 a_10041_993# VSS_SW[3] 0.00296f
C203 a_1757_1642# a_2468_1467# 0.00963f
C204 VDD_SW_b[6] a_5896_909# 2.96e-21
C205 a_5271_n62# a_5812_212# 0.138f
C206 a_4958_n88# a_5813_n88# 0.0477f
C207 a_8432_993# a_9761_627# 3.24e-21
C208 x9.A1 a_13705_304# 4.37e-21
C209 a_78_90# a_174_n88# 0.0967f
C210 a_8204_212# a_10597_n88# 5.48e-21
C211 a_12153_627# a_12433_993# 0.15f
C212 a_12541_627# VSS_SW[2] 3.8e-19
C213 x7.X a_1757_1315# 2.09e-19
C214 x2.X a_3070_220# 0.0028f
C215 check[5] a_2897_1289# 0.251f
C216 x9.A1 a_7394_1642# 9.48e-19
C217 x3.A x2.X 2.91e-19
C218 a_4689_2457# D[6] 0.00292f
C219 x3.X a_939_2457# 0.619f
C220 x2.X a_1363_627# 0.00111f
C221 a_8679_1642# check[2] 8.62e-21
C222 a_305_2457# ready 0.0596f
C223 a_7369_627# a_7350_n88# 4.91e-19
C224 x2.X a_557_993# 5.31e-19
C225 a_10073_1289# a_9595_627# 0.00104f
C226 D[1] a_15518_304# 9.65e-19
C227 a_12036_1467# x16.X 0.0876f
C228 x9.A1 a_15293_601# 0.00103f
C229 a_13375_895# a_14825_993# 8e-21
C230 a_12153_627# a_14733_627# 3.67e-21
C231 a_12901_601# a_15293_601# 9.37e-21
C232 x2.X a_14428_1467# 2.88e-19
C233 VDD_SW_b[4] a_8921_n62# 5.22e-19
C234 VDD_SW_b[4] a_10215_601# 2.46e-20
C235 a_7681_1289# a_7823_601# 8.76e-20
C236 x2.X a_4977_627# 0.0537f
C237 x2.X VSS_SW[5] 0.0861f
C238 a_12680_106# a_12924_n62# 0.00707f
C239 a_4413_2457# VSS_SW[5] 3.26e-20
C240 a_12447_n62# a_13103_n62# 3.73e-19
C241 VDD check[6] 1.68f
C242 a_8432_993# a_8677_122# 1.51e-20
C243 a_7967_627# a_7350_n88# 1.08e-19
C244 VDD a_11546_1315# 3.89e-19
C245 a_11987_627# a_12680_106# 3.88e-21
C246 D[2] a_12447_n62# 0.00257f
C247 VDD_SW_b[1] a_15316_n62# 8.09e-20
C248 a_3039_601# a_2773_627# 8.07e-20
C249 x9.A1 a_1946_n62# 1.9e-20
C250 a_2585_627# a_2949_993# 0.0018f
C251 a_3333_601# a_3807_895# 0.265f
C252 x9.X a_5725_601# 4.04e-21
C253 a_3420_212# a_3421_n88# 0.785f
C254 a_2879_n62# a_3893_122# 0.0633f
C255 a_3112_106# a_3625_n88# 0.00189f
C256 a_2566_n88# VSS_SW_b[6] 0.135f
C257 a_15855_1642# a_15767_895# 5.45e-19
C258 a_14999_601# a_15464_909# 9.46e-19
C259 a_10215_601# VDD_SW[3] 2.07e-20
C260 a_10509_601# a_11123_627# 0.0526f
C261 a_10983_895# a_11704_627# 0.0967f
C262 x17.X check[0] 5.47e-19
C263 x2.X a_9312_627# 3.88e-19
C264 D[3] a_11704_627# 0.00234f
C265 x2.X a_16109_1315# 2.32e-19
C266 x2.X a_15715_627# 0.00111f
C267 a_15380_212# a_15518_304# 1.09e-19
C268 VDD_SW[4] a_10041_993# 7.03e-20
C269 VDD a_2879_n62# 0.326f
C270 x9.A1 a_8933_1642# 0.195f
C271 x2.X a_5575_627# 0.0388f
C272 VDD_SW[6] a_6199_895# 1.27e-20
C273 VDD_SW_b[6] VSS_SW_b[5] 0.0382f
C274 VDD a_10597_n88# 0.66f
C275 reset x6.X 2.16e-19
C276 a_13461_1642# a_13461_122# 1.57e-21
C277 VDD_SW_b[2] a_13461_122# 0.00445f
C278 x2.X a_12924_n62# 3.67e-20
C279 a_11539_1642# VDD_SW[3] 5.44e-19
C280 x14.X check[2] 0.00901f
C281 a_7896_106# VSS_SW[3] 9.06e-21
C282 x2.X a_11987_627# 0.354f
C283 a_8204_212# a_8545_n62# 0.00134f
C284 a_8205_n88# a_8319_n62# 2.14e-20
C285 a_3333_601# VDD_SW_b[6] 0.00635f
C286 a_2419_627# a_4811_627# 1.63e-20
C287 a_2773_627# a_2973_627# 3.81e-19
C288 a_3807_895# a_4064_909# 0.00869f
C289 a_3648_993# a_3551_627# 0.00386f
C290 x2.X VDD_SW_b[3] 7.39e-19
C291 x12.X a_7615_1315# 2.41e-19
C292 a_5323_2457# x11.X 3.12e-19
C293 a_10288_106# a_12134_n88# 1.86e-21
C294 a_14096_627# a_14545_627# 5.39e-19
C295 x9.A1 a_7350_n88# 7.41e-19
C296 reset a_27_627# 7.49e-21
C297 a_2897_1289# a_2865_993# 4.54e-19
C298 a_5812_212# a_5950_304# 1.09e-19
C299 a_10055_n62# a_11069_122# 0.0633f
C300 a_10288_106# a_10801_n88# 0.00189f
C301 a_10596_212# a_10597_n88# 0.784f
C302 a_487_n62# VSS_SW_b[7] 0.0142f
C303 a_1028_212# a_1233_n88# 0.15f
C304 VSS_SW[7] a_977_304# 8.35e-20
C305 check[3] VDD_SW[5] 4.37e-19
C306 x12.X a_7203_627# 0.236f
C307 VDD D[7] 0.791f
C308 a_12447_n62# VSS_SW_b[1] 1.09e-20
C309 a_12989_n88# a_15381_n88# 1.33e-19
C310 VDD a_8067_909# 0.00984f
C311 a_4064_909# VDD_SW_b[6] 3.4e-20
C312 a_8205_n88# a_10288_106# 1.67e-21
C313 D[2] a_13126_304# 9.67e-19
C314 check[6] a_941_601# 2.14e-19
C315 a_7823_601# a_8288_909# 9.46e-19
C316 a_14999_601# VDD_SW[1] 2.07e-20
C317 a_15293_601# a_15907_627# 0.0526f
C318 a_15767_895# a_16488_627# 0.0967f
C319 x9.A1 a_6467_1642# 5.26e-19
C320 x10.X a_5431_601# 2.7e-20
C321 a_10073_1289# a_10041_993# 4.54e-19
C322 D[6] a_3625_n88# 0.00546f
C323 check[3] a_7711_1642# 0.00526f
C324 x9.X a_5271_n62# 4.43e-20
C325 x9.A1 a_439_1315# 0.00504f
C326 VDD a_12638_220# 0.00411f
C327 x9.A1 x7.X 6.79e-19
C328 a_6017_n88# VSS_SW[4] 8.81e-20
C329 a_6285_122# a_6153_n62# 0.025f
C330 VSS_SW_b[5] a_5927_n62# 5.23e-19
C331 VDD a_2419_627# 0.393f
C332 x9.A1 a_12465_1289# 0.104f
C333 D[5] a_5431_601# 0.00583f
C334 a_4811_627# a_5257_993# 0.159f
C335 x2.X a_15853_122# 0.00427f
C336 a_12433_993# VDD_SW_b[2] 3.93e-21
C337 a_12901_601# a_13632_909# 0.0016f
C338 x2.X a_76_1467# 2.67e-19
C339 VDD a_8545_n62# 0.0301f
C340 VDD a_4077_1642# 8.63e-19
C341 VDD a_535_1642# 9.76e-19
C342 x2.X a_3648_993# 0.187f
C343 x9.A1 a_3420_212# 1.41e-20
C344 a_3421_n88# a_4137_304# 0.0018f
C345 a_3625_n88# a_3839_220# 0.0104f
C346 a_2879_n62# a_2985_n62# 0.0526f
C347 a_3420_212# a_4338_n62# 0.0453f
C348 VSS_SW[2] a_12988_212# 1.18e-21
C349 a_505_1289# x7.X 1.75e-20
C350 a_14379_627# a_14733_627# 0.0455f
C351 x14.X a_9312_627# 0.0285f
C352 check[0] a_14545_627# 5.41e-19
C353 a_14857_1289# D[1] 0.0662f
C354 x2.X a_174_n88# 0.178f
C355 D[1] a_15608_993# 0.00606f
C356 a_3895_1642# a_3947_627# 1.92e-20
C357 D[3] a_12447_n62# 3.12e-21
C358 VDD_SW_b[7] a_2566_n88# 5.91e-19
C359 VDD a_3558_304# 0.0164f
C360 VDD_SW_b[2] a_14733_627# 9.33e-21
C361 check[2] a_9646_90# 2.5e-20
C362 x15.X a_11546_1315# 0.00143f
C363 a_10824_993# a_10801_n88# 1.86e-19
C364 a_10983_895# a_11069_122# 4.53e-22
C365 a_4811_627# a_5943_627# 0.00272f
C366 D[3] a_11069_122# 0.00933f
C367 x8.X D[6] 0.00886f
C368 a_13126_304# VSS_SW_b[1] 9.89e-21
C369 a_13906_n62# a_15381_n88# 3.67e-21
C370 VDD a_1112_909# 0.0166f
C371 a_14430_90# a_15380_212# 2.02e-20
C372 check[5] a_2566_n88# 5.27e-19
C373 a_12988_212# a_14945_n62# 1.09e-19
C374 x9.A1 a_14839_n62# 1.54e-20
C375 D[7] a_941_601# 0.019f
C376 a_27_627# a_1415_895# 0.0321f
C377 VDD_SW_b[4] a_8140_n62# 8.1e-20
C378 a_8623_220# VSS_SW[3] 1.57e-20
C379 a_9644_1467# check[3] 1.56e-19
C380 a_3504_909# VDD_SW[6] 2.82e-20
C381 check[1] a_12680_106# 8.64e-22
C382 a_6539_1642# x11.X 0.0845f
C383 VDD_SW[3] a_13375_895# 1.27e-20
C384 check[2] VDD_SW[3] 0.00394f
C385 x16.X a_10215_601# 1.98e-20
C386 x15.X a_10597_n88# 0.0189f
C387 x2.X a_10509_601# 0.119f
C388 a_5289_1289# a_4811_627# 0.00104f
C389 x12.X a_6760_1315# 4.97e-20
C390 VDD a_4149_1642# 0.115f
C391 VDD a_5257_993# 0.18f
C392 a_5725_601# a_7823_601# 1.55e-20
C393 a_6199_895# a_7369_627# 2.8e-19
C394 x27.A x9.X 9.96e-20
C395 a_15767_895# a_15381_n88# 6.35e-19
C396 a_15293_601# a_15585_n88# 0.00251f
C397 a_15608_993# a_15380_212# 8.94e-21
C398 a_2468_1467# check[6] 1.54e-19
C399 x2.X a_2897_1289# 0.0112f
C400 a_5812_212# a_7350_n88# 6.19e-19
C401 a_941_601# a_2419_627# 3.79e-19
C402 VSS_SW_b[7] a_1447_220# 1.12e-20
C403 a_5323_2457# a_6920_627# 3.86e-19
C404 a_1233_n88# a_1946_n62# 8.07e-20
C405 x2.X a_15316_n62# 3.67e-20
C406 a_720_106# a_964_n62# 0.00707f
C407 a_487_n62# a_1143_n62# 3.73e-19
C408 a_1501_122# a_1745_304# 0.00972f
C409 a_1029_n88# a_2470_90# 5.39e-19
C410 D[7] a_1672_909# 8.06e-19
C411 a_27_627# VDD_SW_b[7] 1.09e-19
C412 a_12851_909# VDD_SW[2] 1.01e-20
C413 x18.X a_12433_993# 1.55e-20
C414 x2.X check[1] 0.15f
C415 a_4811_627# a_4958_n88# 0.00176f
C416 a_193_627# a_647_601# 0.117f
C417 x2.X a_7615_1315# 3.2e-19
C418 a_8117_601# a_8731_627# 0.0526f
C419 a_8591_895# a_9312_627# 0.0967f
C420 a_7823_601# VDD_SW[4] 2.07e-20
C421 x30.A x2.X 0.002f
C422 x27.A a_4689_2457# 0.3f
C423 ready a_5323_2457# 4.34e-19
C424 a_4413_2457# x30.A 6.66e-19
C425 a_13193_n88# VSS_SW_b[2] 9.26e-19
C426 x6.X a_78_90# 0.00259f
C427 VDD a_5943_627# 6.2e-19
C428 D[6] a_4862_90# 8.78e-19
C429 VDD_SW_b[5] a_7369_627# 0.00336f
C430 a_14379_627# a_16488_627# 1.75e-19
C431 a_10680_909# VDD_SW_b[3] 7.05e-21
C432 a_10359_627# a_10727_627# 3.34e-19
C433 x18.X a_15855_1642# 1.97e-20
C434 x9.A1 a_193_627# 3.22e-19
C435 x18.X a_14733_627# 6.12e-19
C436 a_7254_90# VSS_SW[4] 0.082f
C437 a_9761_627# a_10727_627# 2.14e-20
C438 a_9595_627# a_10908_993# 2.13e-19
C439 a_1256_993# a_1363_627# 0.00707f
C440 a_1415_895# VDD_SW[7] 0.00356f
C441 VDD a_305_2457# 0.359f
C442 a_14428_1467# a_14526_n88# 6.87e-20
C443 x2.X a_7203_627# 0.354f
C444 VDD a_11313_304# 0.00421f
C445 a_647_601# a_791_627# 0.0697f
C446 a_941_601# a_1112_909# 0.00652f
C447 VDD a_5289_1289# 0.191f
C448 VDD_SW_b[4] a_9312_627# 0.186f
C449 x9.A1 a_9786_1642# 8.64e-19
C450 a_11987_627# a_13119_627# 0.00272f
C451 x9.A1 a_4137_304# 6.9e-21
C452 a_27_627# a_78_90# 6.13e-19
C453 check[2] a_11071_1642# 0.257f
C454 a_3421_n88# a_5504_106# 1.67e-21
C455 a_3893_122# a_4958_n88# 8e-21
C456 a_3420_212# a_5812_212# 9.5e-22
C457 a_4137_304# a_4338_n62# 8.99e-19
C458 a_505_1289# a_193_627# 0.00323f
C459 a_9786_1315# VSS_SW[3] 7.95e-19
C460 a_2468_1467# D[7] 2.91e-19
C461 x2.X a_1166_304# 0.00334f
C462 VDD a_13300_993# 0.00281f
C463 a_3039_601# a_2879_n62# 0.0026f
C464 a_2865_993# a_2566_n88# 8.71e-20
C465 VDD a_4958_n88# 0.69f
C466 a_15767_895# a_16298_n62# 4.06e-19
C467 VDD_SW_b[7] VDD_SW[7] 3.64e-19
C468 a_891_909# VDD_SW_b[7] 2.4e-21
C469 a_10597_n88# a_11015_220# 0.00276f
C470 a_10801_n88# a_10734_304# 9.46e-19
C471 a_10596_212# a_11313_304# 4.45e-20
C472 VSS_SW_b[3] a_10246_220# 5.34e-20
C473 a_10055_n62# a_12038_90# 3.67e-21
C474 a_9742_n88# a_10161_n62# 0.0383f
C475 a_939_2457# x7.X 2.98e-19
C476 check[5] VDD_SW[7] 4.38e-19
C477 x9.A1 a_6199_895# 2.54e-19
C478 check[3] a_8677_122# 6.43e-20
C479 VSS_SW[3] a_10055_n62# 3.44e-19
C480 x7.X a_1233_n88# 1.81e-19
C481 VDD a_16024_909# 0.00438f
C482 VDD a_13936_1315# 3.62e-19
C483 x9.A1 a_13193_n88# 3.88e-20
C484 check[6] VSS_SW_b[7] 3.18e-20
C485 a_2468_1467# a_2419_627# 5.32e-19
C486 a_12901_601# a_13193_n88# 0.00251f
C487 a_13375_895# a_12989_n88# 6.35e-19
C488 a_13216_993# a_12988_212# 8.94e-21
C489 x11.X a_5725_601# 1.29e-19
C490 VDD_SW[3] a_11987_627# 0.0865f
C491 check[0] VDD_SW_b[1] 0.00215f
C492 VDD_SW_b[3] VDD_SW[3] 3.63e-19
C493 a_2773_627# VSS_SW_b[6] 5.82e-19
C494 check[0] x20.X 0.00965f
C495 x18.X a_14570_1315# 8.21e-19
C496 x2.X a_10246_220# 0.00279f
C497 x14.X a_10509_601# 4.89e-20
C498 a_6539_1642# a_6920_627# 5.84e-19
C499 x3.X a_473_993# 4.27e-21
C500 VDD a_2949_993# 0.0042f
C501 a_487_n62# VSS_SW_b[6] 1.09e-20
C502 a_1029_n88# a_3421_n88# 1.33e-19
C503 VDD a_11704_627# 0.194f
C504 D[1] a_15380_212# 0.157f
C505 x3.A VSS_SW[7] 0.0165f
C506 a_14379_627# a_15381_n88# 1.06e-19
C507 x9.A1 VDD_SW_b[5] 1.13e-19
C508 a_5431_601# a_5675_909# 0.0104f
C509 a_5725_601# a_5165_627# 1.15e-20
C510 a_4977_627# a_5896_909# 0.00907f
C511 a_6199_895# a_6040_993# 0.207f
C512 a_5257_993# a_5341_993# 0.00972f
C513 VDD_SW_b[2] a_15381_n88# 2.44e-21
C514 D[5] a_5462_220# 1.98e-20
C515 a_11325_1642# a_11253_1642# 6.64e-19
C516 VDD a_720_106# 0.356f
C517 check[2] x16.X 6.04e-19
C518 x2.X a_12341_627# 0.00141f
C519 D[6] a_5813_n88# 4.83e-22
C520 VDD_SW[5] a_7557_627# 6.11e-20
C521 a_7203_627# a_8409_n88# 0.00204f
C522 D[4] a_8205_n88# 0.158f
C523 a_2419_627# a_3039_601# 0.149f
C524 VSS_SW[4] a_8205_n88# 9.29e-21
C525 D[6] a_2585_627# 0.168f
C526 x10.X a_4528_627# 0.0285f
C527 a_7252_1467# a_7203_627# 5.32e-19
C528 a_10509_601# a_10680_909# 0.00652f
C529 a_10215_601# a_10359_627# 0.0697f
C530 a_11704_627# a_10596_212# 6.63e-19
C531 a_6040_993# VDD_SW_b[5] 5e-20
C532 D[5] D[4] 0.00183f
C533 D[3] a_10459_909# 6.77e-19
C534 D[3] a_12038_90# 8.76e-19
C535 a_9761_627# a_10215_601# 0.117f
C536 x2.X a_15692_993# 4.67e-19
C537 D[5] VSS_SW[4] 4.85e-19
C538 check[4] check[3] 0.00525f
C539 a_15072_106# a_15381_n88# 0.0327f
C540 x14.X a_7203_627# 0.00113f
C541 a_14526_n88# a_15853_122# 4.59e-22
C542 a_14839_n62# a_15585_n88# 0.199f
C543 a_3895_1642# D[6] 0.0681f
C544 check[3] a_8432_993# 3.41e-19
C545 D[3] VSS_SW[3] 0.134f
C546 D[7] VSS_SW_b[7] 5.32e-19
C547 a_8591_895# a_10509_601# 1.54e-20
C548 a_3947_627# a_4811_627# 1.09e-19
C549 a_4528_627# D[5] 4.42e-19
C550 a_13375_895# a_13906_n62# 4.06e-19
C551 x9.A1 a_12607_601# 2.81e-20
C552 a_4862_90# a_5271_n62# 4.24e-20
C553 a_12607_601# a_12901_601# 0.199f
C554 a_12153_627# a_13375_895# 0.0494f
C555 a_12465_1289# VSS_SW[2] 0.00187f
C556 check[5] a_2610_1642# 0.00688f
C557 x9.A1 a_8861_1642# 5.26e-19
C558 x12.X a_5431_601# 1.98e-20
C559 x11.X a_5271_n62# 0.002f
C560 x2.X a_2566_n88# 0.178f
C561 a_2419_627# a_2973_627# 0.00206f
C562 ready D[6] 0.0519f
C563 a_7681_1289# x13.X 1.75e-20
C564 a_1757_1642# a_1415_895# 0.00232f
C565 VDD a_5761_304# 0.00266f
C566 VDD_SW[7] a_2865_993# 7.03e-20
C567 a_1415_895# a_2773_627# 8.26e-21
C568 D[1] a_16097_304# 8.37e-19
C569 a_939_2457# a_193_627# 2.84e-21
C570 x9.X a_3420_212# 0.244f
C571 x9.A1 a_14857_1289# 0.105f
C572 x9.A1 a_15608_993# 4.84e-21
C573 VDD_SW_b[4] a_10509_601# 2.26e-20
C574 x2.X x6.X 2.59e-20
C575 a_5725_601# a_5813_n88# 3.89e-19
C576 a_4977_627# VSS_SW_b[5] 5.23e-20
C577 a_6199_895# a_5812_212# 0.00165f
C578 x2.X a_14096_627# 3.85e-19
C579 a_647_601# a_1029_n88# 0.00322f
C580 a_941_601# a_720_106# 3.46e-19
C581 a_193_627# a_1233_n88# 8.75e-19
C582 VSS_SW[5] VSS_SW_b[5] 0.00723f
C583 a_1415_895# a_487_n62# 0.00219f
C584 a_5323_2457# a_4811_627# 4.8e-19
C585 a_8677_122# a_8921_n62# 0.00807f
C586 a_3333_601# a_4977_627# 6.25e-20
C587 a_12680_106# a_13329_n62# 0.00316f
C588 a_12988_212# a_13103_n62# 0.00272f
C589 a_12447_n62# VSS_SW[1] 1.64e-20
C590 a_3947_627# a_3893_122# 2.54e-20
C591 a_3333_601# VSS_SW[5] 2.89e-20
C592 a_3807_895# a_3761_n62# 1.65e-20
C593 a_1757_1642# VDD_SW_b[7] 2.58e-19
C594 D[2] a_12988_212# 0.158f
C595 a_7203_627# a_8591_895# 0.0321f
C596 D[4] a_8117_601# 0.0191f
C597 a_11987_627# a_12989_n88# 1.06e-19
C598 VDD_SW_b[1] a_15721_n62# 0.00178f
C599 VDD_SW_b[3] a_12989_n88# 2.44e-21
C600 a_8117_601# VSS_SW[4] 2.17e-19
C601 a_14999_601# a_15143_627# 0.0697f
C602 x9.A1 a_1029_n88# 8.52e-21
C603 a_15293_601# a_15464_909# 0.00652f
C604 a_7350_n88# a_7896_106# 0.207f
C605 a_10824_993# a_11123_627# 0.0256f
C606 a_10509_601# VDD_SW[3] 1.79e-19
C607 VDD_SW_b[7] a_2773_627# 9.33e-21
C608 VDD a_3947_627# 6.99e-19
C609 a_10073_1289# a_10055_n62# 3.44e-19
C610 D[3] a_10931_627# 2e-19
C611 a_1447_220# VSS_SW_b[6] 3.96e-21
C612 a_1757_1642# check[5] 1.67e-19
C613 a_2470_90# a_3421_n88# 9.87e-21
C614 x2.X a_27_627# 0.352f
C615 a_5725_601# a_6920_627# 5.73e-19
C616 a_4977_627# VDD_SW[5] 1.96e-20
C617 x2.X a_7733_993# 5.31e-19
C618 a_15380_212# a_16097_304# 4.45e-20
C619 a_15585_n88# a_15518_304# 9.46e-19
C620 VSS_SW_b[1] a_15030_220# 5.34e-20
C621 a_14839_n62# a_14945_n62# 0.0526f
C622 a_15381_n88# a_15799_220# 0.00276f
C623 VDD a_12447_n62# 0.326f
C624 VDD_SW_b[5] a_5812_212# 0.0417f
C625 VDD_SW[4] a_10983_895# 1.27e-20
C626 VDD_SW_b[7] a_487_n62# 5.22e-19
C627 VDD_SW[4] D[3] 4.43e-19
C628 x9.A1 a_11325_1642# 0.195f
C629 VDD a_1745_304# 0.0042f
C630 VDD a_11069_122# 0.313f
C631 a_9644_1467# check[2] 0.318f
C632 VDD_SW_b[6] a_3761_n62# 0.00179f
C633 check[1] VDD_SW[3] 4.32e-19
C634 x16.X a_11987_627# 0.236f
C635 x16.X VDD_SW_b[3] 7.25e-19
C636 x15.X a_11704_627# 0.0338f
C637 D[4] a_8848_909# 8.06e-19
C638 a_7203_627# VDD_SW_b[4] 1.15e-19
C639 a_1503_1642# a_1028_212# 1.39e-21
C640 D[4] a_9122_n62# 0.158f
C641 a_8677_122# VSS_SW_b[4] 7.15e-19
C642 a_76_1467# VSS_SW[7] 0.0274f
C643 a_10532_n62# a_10937_n62# 2.46e-21
C644 a_16109_1642# a_15293_601# 7.12e-21
C645 VDD a_5323_2457# 1.38f
C646 a_10041_993# a_10161_n62# 6.88e-22
C647 a_10597_n88# a_12134_n88# 1.98e-19
C648 a_10596_212# a_12447_n62# 2.62e-19
C649 x2.X check[0] 0.149f
C650 a_10288_106# VSS_SW_b[3] 0.00322f
C651 VSS_SW[3] a_10545_304# 8.35e-20
C652 a_10597_n88# a_10801_n88# 0.117f
C653 a_10596_212# a_11069_122# 0.159f
C654 x2.X a_10007_1315# 3.2e-19
C655 a_5271_n62# a_5813_n88# 0.125f
C656 a_5504_106# a_5812_212# 0.14f
C657 a_12988_212# VSS_SW_b[1] 0.00377f
C658 a_13126_304# VSS_SW[1] 2.77e-20
C659 VSS_SW[7] a_174_n88# 0.00677f
C660 a_78_90# a_487_n62# 4.24e-20
C661 a_12607_601# a_12553_n62# 1.07e-20
C662 a_8205_n88# a_10597_n88# 1.33e-19
C663 D[2] a_13705_304# 8.38e-19
C664 a_11987_627# a_12153_627# 0.786f
C665 x2.X a_3369_304# 0.00168f
C666 VDD_SW_b[3] a_12153_627# 0.00336f
C667 a_15293_601# VDD_SW[1] 1.83e-19
C668 a_15608_993# a_15907_627# 0.0256f
C669 x2.X VDD_SW[7] 0.0768f
C670 x3.X ready 0.127f
C671 a_7823_601# a_7350_n88# 4.37e-19
C672 a_7369_627# a_7663_n62# 2.38e-19
C673 a_11071_1642# a_10509_601# 0.00263f
C674 a_10073_1289# D[3] 0.0662f
C675 x2.X a_891_909# 0.00138f
C676 check[2] a_9761_627# 5.35e-19
C677 check[3] a_9147_1642# 0.00688f
C678 x2.X a_10288_106# 0.0385f
C679 VDD a_13126_304# 0.0164f
C680 x13.X VSS_SW[3] 0.149f
C681 a_5431_601# a_5377_n62# 1.07e-20
C682 a_14999_601# VSS_SW[1] 6.23e-19
C683 VDD a_7681_1289# 0.191f
C684 x9.A1 D[1] 0.268f
C685 D[2] a_15293_601# 2.67e-21
C686 a_13375_895# a_14379_627# 6.9e-19
C687 a_12901_601# D[1] 8.7e-19
C688 a_7681_1289# a_7649_993# 4.54e-19
C689 x9.A1 a_12178_1642# 8.64e-19
C690 a_13461_1642# a_13375_895# 5.55e-19
C691 a_13375_895# VDD_SW_b[2] 0.128f
C692 a_11071_1642# check[1] 6.17e-21
C693 reset check[6] 1.32e-20
C694 x9.A1 VDD_SW[6] 0.0329f
C695 x2.X a_5431_601# 0.2f
C696 VDD a_218_1315# 6.87e-19
C697 a_12134_n88# a_12638_220# 0.00869f
C698 VDD a_14999_601# 0.313f
C699 a_3039_601# a_2949_993# 6.69e-20
C700 a_7663_n62# a_8342_304# 0.00652f
C701 a_2585_627# a_3283_909# 0.00276f
C702 a_3333_601# a_3648_993# 0.13f
C703 a_2865_993# a_2773_627# 0.0369f
C704 a_7896_106# a_8153_304# 0.00857f
C705 VSS_SW[2] a_13193_n88# 9.93e-21
C706 a_3420_212# a_3625_n88# 0.15f
C707 VSS_SW[6] a_3070_220# 4.25e-19
C708 a_2879_n62# VSS_SW_b[6] 0.0142f
C709 D[1] a_14909_993# 8.12e-19
C710 check[0] a_14825_993# 7.14e-20
C711 a_14379_627# a_15243_909# 2.46e-19
C712 x2.X a_8731_627# 0.0151f
C713 a_11069_122# a_11313_n62# 0.00807f
C714 D[3] a_12988_212# 5.78e-20
C715 VDD_SW_b[2] a_15243_909# 2.1e-21
C716 x10.X a_2419_627# 0.00117f
C717 VDD a_3112_106# 0.356f
C718 VDD_SW[6] a_6040_993# 1.08e-20
C719 x2.X a_5365_627# 3.94e-19
C720 x9.A1 a_15380_212# 1.41e-20
C721 check[1] a_12989_n88# 2.51e-20
C722 x15.X a_12447_n62# 4.73e-20
C723 VDD_SW[3] a_12341_627# 6.11e-20
C724 VSS_SW_b[4] a_7769_n62# 0.00335f
C725 a_2419_627# D[5] 1.19e-20
C726 D[6] a_4811_627# 9.98e-20
C727 a_3807_895# VDD_SW_b[6] 0.129f
C728 a_8205_n88# a_8545_n62# 6.04e-20
C729 a_8409_n88# a_8319_n62# 9.75e-19
C730 a_8204_212# VSS_SW[3] 0.0872f
C731 x16.X a_10509_601# 0.00124f
C732 x7.X x8.X 0.11f
C733 x15.X a_11069_122# 2.61e-19
C734 x2.X a_10824_993# 0.187f
C735 VDD a_6539_1642# 0.115f
C736 x13.X VDD_SW[4] 0.177f
C737 a_15608_993# a_15585_n88# 1.86e-19
C738 a_15767_895# a_15853_122# 4.53e-22
C739 a_14428_1467# a_14379_627# 5.32e-19
C740 a_13715_1642# D[1] 1.62e-19
C741 D[7] VSS_SW_b[6] 2.02e-19
C742 a_8679_1642# a_8731_627# 1.92e-20
C743 a_12036_1467# a_12495_1642# 6.64e-19
C744 x9.A1 a_7663_n62# 1.53e-20
C745 a_12751_627# a_13323_627# 2.46e-21
C746 x18.X a_13375_895# 0.00863f
C747 a_9312_627# a_9761_627# 5.39e-19
C748 a_5812_212# a_6231_220# 2.46e-19
C749 a_5813_n88# a_5950_304# 0.00907f
C750 a_5271_n62# a_6730_n62# 3.79e-20
C751 x16.X check[1] 0.00902f
C752 a_720_106# VSS_SW_b[7] 0.00322f
C753 a_1029_n88# a_1233_n88# 0.117f
C754 VSS_SW[7] a_1166_304# 1.97e-20
C755 a_1028_212# a_1501_122# 0.159f
C756 x14.X a_10007_1315# 2.35e-19
C757 x12.X D[4] 0.00875f
C758 a_9122_n62# a_10597_n88# 3.67e-21
C759 x12.X VSS_SW[4] 0.253f
C760 x11.X a_7350_n88# 0.00864f
C761 VDD a_8288_909# 0.0164f
C762 VDD a_7854_220# 0.0041f
C763 a_8117_601# a_8067_909# 1.21e-20
C764 a_7369_627# a_7967_627# 6.04e-20
C765 check[6] a_1415_895# 0.00271f
C766 ready x27.A 0.00414f
C767 a_12607_601# VSS_SW[2] 6.25e-19
C768 a_4149_1642# x10.X 7.97e-19
C769 x10.X a_5257_993# 1.03e-19
C770 D[1] a_15907_627# 0.0043f
C771 a_14791_1315# D[1] 0.00202f
C772 D[6] a_3893_122# 0.00928f
C773 a_10509_601# a_12153_627# 6.25e-20
C774 a_2419_627# VSS_SW_b[6] 1.08e-19
C775 a_9761_627# a_11987_627# 1.36e-20
C776 x9.A1 a_1757_1315# 0.00499f
C777 a_9761_627# VDD_SW_b[3] 0.00226f
C778 a_9595_627# a_10149_627# 0.00206f
C779 a_6285_122# VSS_SW[4] 6.66e-20
C780 VSS_SW_b[5] a_6153_n62# 5.34e-19
C781 VDD D[6] 0.784f
C782 x9.A1 a_16097_304# 8.15e-21
C783 VDD a_10459_909# 0.00984f
C784 VDD a_12038_90# 0.189f
C785 a_4811_627# a_5725_601# 0.14f
C786 D[5] a_5257_993# 0.00874f
C787 a_4149_1642# D[5] 1.74e-19
C788 VDD_SW_b[2] a_12924_n62# 8.1e-20
C789 VDD a_5002_1642# 0.00177f
C790 a_11987_627# a_14379_627# 1.74e-20
C791 x2.X a_1757_1642# 5.76e-19
C792 D[2] a_13632_909# 8.06e-19
C793 check[1] a_12153_627# 5.41e-19
C794 VDD VSS_SW[3] 0.523f
C795 a_11987_627# VDD_SW_b[2] 1.09e-19
C796 a_12465_1289# D[2] 0.0662f
C797 x9.A1 a_11253_1642# 5.26e-19
C798 check[6] VDD_SW_b[7] 0.00217f
C799 a_8731_627# a_8409_n88# 7.32e-20
C800 VDD_SW[4] a_8204_212# 4.35e-19
C801 check[2] a_10103_1642# 0.00526f
C802 x9.A1 a_3421_n88# 8.52e-21
C803 x2.X a_2773_627# 0.0014f
C804 VDD a_1685_1642# 8.63e-19
C805 a_7663_n62# a_9742_n88# 5.13e-21
C806 a_3625_n88# a_4137_304# 6.69e-20
C807 a_3420_212# a_4862_90# 0.00101f
C808 VSS_SW_b[6] a_3558_304# 3.58e-20
C809 a_3112_106# a_2985_n62# 0.0256f
C810 a_2879_n62# a_3356_n62# 1.96e-20
C811 a_3421_n88# a_4338_n62# 0.189f
C812 VDD_SW[5] a_7203_627# 0.0865f
C813 a_1503_1642# x7.X 1.35e-19
C814 check[6] check[5] 0.00521f
C815 a_15907_627# a_15380_212# 7.07e-21
C816 a_14428_1467# x18.X 0.0878f
C817 x2.X a_487_n62# 0.374f
C818 VDD a_3839_220# 0.00984f
C819 x9.A1 a_7369_627# 3.48e-19
C820 a_10801_n88# a_11313_304# 6.69e-20
C821 a_10596_212# a_12038_90# 0.00101f
C822 VSS_SW_b[3] a_10734_304# 3.58e-20
C823 a_10597_n88# a_11514_n62# 0.189f
C824 D[5] a_5943_627# 6.13e-19
C825 a_27_627# a_2136_627# 1.75e-19
C826 check[5] a_2879_n62# 1.43e-20
C827 VDD a_1340_993# 0.00281f
C828 a_174_n88# a_678_220# 0.00869f
C829 x10.X a_5289_1289# 1.54e-19
C830 VSS_SW[3] a_10596_212# 5.9e-22
C831 a_1971_1642# VDD_SW[7] 5.38e-19
C832 VDD_SW_b[4] a_8319_n62# 5.2e-19
C833 a_27_627# a_1256_993# 0.14f
C834 D[7] a_1415_895# 0.0294f
C835 D[2] a_14839_n62# 3.12e-21
C836 a_3183_627# a_3755_627# 2.46e-21
C837 a_8921_304# VSS_SW[3] 6.59e-21
C838 a_7769_n62# a_8140_n62# 4.19e-20
C839 x9.A1 VSS_SW_b[2] 2.85e-19
C840 a_13216_993# a_13193_n88# 1.86e-19
C841 a_13375_895# a_13461_122# 4.53e-22
C842 x8.X a_193_627# 6.39e-20
C843 a_8933_1642# D[3] 1.65e-19
C844 check[6] a_78_90# 2.5e-20
C845 x17.X a_13936_1315# 0.00145f
C846 x2.X a_10734_304# 0.00334f
C847 check[4] a_4977_627# 5.33e-19
C848 a_5289_1289# D[5] 0.0662f
C849 VDD a_5725_601# 0.46f
C850 a_4149_1642# a_4363_1642# 0.00557f
C851 check[4] VSS_SW[5] 0.0495f
C852 a_6040_993# a_7369_627# 3.63e-21
C853 a_5725_601# a_7649_993# 1.11e-20
C854 a_5812_212# a_7663_n62# 2.63e-19
C855 a_5813_n88# a_7350_n88# 1.98e-19
C856 D[1] a_15585_n88# 0.00544f
C857 check[0] a_14526_n88# 5.26e-19
C858 a_941_601# D[6] 9.16e-19
C859 a_1415_895# a_2419_627# 6.86e-19
C860 a_174_n88# VSS_SW[6] 4.28e-21
C861 a_487_n62# a_1369_n62# 0.00926f
C862 a_1501_122# a_1946_n62# 0.0369f
C863 a_720_106# a_1143_n62# 0.00386f
C864 D[7] VDD_SW_b[7] 0.453f
C865 x18.X a_11987_627# 0.00113f
C866 D[5] a_4958_n88# 0.00506f
C867 x2.X a_5462_220# 0.00279f
C868 a_4811_627# a_5271_n62# 7.27e-19
C869 VDD VDD_SW[4] 0.374f
C870 x16.X a_12341_627# 6.07e-19
C871 a_193_627# a_473_993# 0.15f
C872 a_8117_601# a_8539_627# 1.96e-20
C873 a_7649_993# VDD_SW[4] 4.17e-21
C874 x2.X a_12851_909# 0.00138f
C875 D[4] VSS_SW_b[3] 1.99e-19
C876 a_8591_895# a_8731_627# 0.0383f
C877 x14.X a_9154_1315# 3.14e-20
C878 check[5] D[7] 6.16e-20
C879 VDD a_6456_909# 0.00438f
C880 x6.X VSS_SW[7] 0.253f
C881 VDD_SW_b[5] a_7823_601# 2.22e-20
C882 a_29_2457# x3.A 0.129f
C883 VDD_SW_b[3] a_10532_n62# 8.12e-20
C884 reset a_305_2457# 0.0023f
C885 x9.A1 a_647_601# 2.81e-20
C886 a_5748_n62# a_6153_n62# 2.46e-21
C887 a_10509_601# a_10359_627# 0.00926f
C888 a_2136_627# VDD_SW[7] 0.0729f
C889 VDD_SW_b[7] a_2419_627# 5.96e-19
C890 a_1555_627# a_1363_627# 4.19e-20
C891 a_10215_601# a_10727_627# 9.75e-19
C892 a_10824_993# a_10680_909# 0.00412f
C893 a_10041_993# a_10149_627# 0.00807f
C894 D[3] a_10908_993# 2.53e-19
C895 a_1256_993# VDD_SW[7] 3.28e-20
C896 x2.X a_12399_1315# 3.21e-19
C897 VDD x3.X 0.703f
C898 x2.X a_14933_627# 3.94e-19
C899 a_9761_627# a_10509_601# 0.126f
C900 x2.X D[4] 0.199f
C901 a_9949_627# VSS_SW[3] 0.00595f
C902 a_15380_212# a_15585_n88# 0.15f
C903 a_14839_n62# VSS_SW_b[1] 0.0142f
C904 VSS_SW[1] a_15030_220# 4.25e-19
C905 a_4149_1642# a_4860_1467# 0.00963f
C906 x2.X VSS_SW[4] 0.0687f
C907 a_2927_1642# D[6] 5.72e-19
C908 a_941_601# a_1340_993# 9.41e-19
C909 a_473_993# a_791_627# 0.025f
C910 a_193_627# a_1159_627# 2.14e-20
C911 a_381_627# a_557_993# 8.99e-19
C912 check[5] a_2419_627# 0.00121f
C913 a_2897_1289# VSS_SW[6] 0.00189f
C914 x7.X a_2585_627# 1.68e-19
C915 a_8591_895# a_10824_993# 1.86e-21
C916 a_13515_627# a_12988_212# 7.07e-21
C917 a_27_627# VSS_SW[7] 0.0576f
C918 x9.A1 a_12901_601# 0.00103f
C919 a_12178_1642# VSS_SW[2] 0.00105f
C920 a_12607_601# a_13216_993# 0.00189f
C921 x9.A1 a_4338_n62# 1.9e-20
C922 x2.X a_4528_627# 3.85e-19
C923 a_12153_627# a_12341_627# 0.189f
C924 a_4413_2457# a_4528_627# 1.19e-21
C925 a_3421_n88# a_5812_212# 4.01e-22
C926 a_3420_212# a_5813_n88# 5.48e-21
C927 check[5] a_4077_1642# 0.00577f
C928 a_505_1289# a_647_601# 8.76e-20
C929 x15.X a_12038_90# 0.0273f
C930 a_12465_1289# D[3] 5.1e-21
C931 VDD a_15030_220# 0.0041f
C932 a_3333_601# a_2566_n88# 0.00259f
C933 a_2865_993# a_2879_n62# 2.63e-19
C934 a_2585_627# a_3420_212# 1.02e-19
C935 a_3039_601# a_3112_106# 1.01e-19
C936 x2.X a_1447_220# 9.51e-19
C937 x9.X VDD_SW[6] 0.179f
C938 VDD a_5271_n62# 0.326f
C939 VDD a_10073_1289# 0.191f
C940 x9.A1 a_14570_1642# 8.64e-19
C941 a_1112_909# VDD_SW_b[7] 4.69e-21
C942 a_10055_n62# a_10161_n62# 0.0526f
C943 a_791_627# a_1159_627# 3.34e-19
C944 a_13375_895# a_14733_627# 8.26e-21
C945 x9.A1 a_505_1289# 0.104f
C946 ready x7.X 5.93e-21
C947 a_3895_1642# a_3420_212# 1.39e-21
C948 check[1] VDD_SW_b[2] 0.0021f
C949 check[1] a_13461_1642# 0.257f
C950 x9.A1 a_6040_993# 4.84e-21
C951 x2.X a_13323_627# 0.00111f
C952 check[3] VSS_SW_b[4] 3.18e-20
C953 a_8679_1642# D[4] 0.0682f
C954 a_7203_627# a_9761_627# 1.08e-20
C955 a_7369_627# a_9595_627# 1.14e-20
C956 a_4689_2457# VDD_SW[6] 0.0305f
C957 x7.X a_1501_122# 2.79e-19
C958 a_12989_n88# a_13329_n62# 6.04e-20
C959 a_13193_n88# a_13103_n62# 9.75e-19
C960 VSS_SW_b[2] a_12553_n62# 0.00334f
C961 a_12988_212# VSS_SW[1] 0.0872f
C962 a_2468_1467# D[6] 0.0183f
C963 x11.X a_6199_895# 0.00663f
C964 a_218_1642# VSS_SW[7] 0.00105f
C965 D[2] a_13193_n88# 0.00546f
C966 a_15608_993# a_15464_909# 0.00412f
C967 a_15293_601# a_15143_627# 0.00926f
C968 a_14999_601# a_15511_627# 9.75e-19
C969 a_14825_993# a_14933_627# 0.00807f
C970 a_14545_627# a_16024_909# 7.17e-20
C971 a_10824_993# VDD_SW[3] 3.28e-20
C972 a_9154_1315# VDD_SW_b[4] 2.65e-20
C973 x9.A1 a_9742_n88# 7.41e-19
C974 a_6285_122# a_6529_n62# 0.00807f
C975 a_6730_n62# a_7350_n88# 8.26e-21
C976 a_4149_1642# check[5] 0.318f
C977 a_1757_1642# a_1971_1642# 0.00557f
C978 a_15381_n88# a_16298_n62# 0.189f
C979 a_15585_n88# a_16097_304# 6.69e-20
C980 a_14839_n62# a_15495_n62# 3.73e-19
C981 a_1166_304# VSS_SW[6] 2.77e-20
C982 VDD a_3283_909# 0.00984f
C983 x3.X a_941_601# 6.38e-19
C984 VSS_SW_b[1] a_15518_304# 3.58e-20
C985 a_15072_106# a_15316_n62# 0.00707f
C986 VDD a_12988_212# 0.687f
C987 VDD_SW[4] a_9949_627# 6.11e-20
C988 a_5431_601# a_5896_909# 9.46e-19
C989 x9.A1 a_13715_1642# 0.195f
C990 a_13715_1642# a_12901_601# 7.56e-21
C991 a_4860_1467# a_4958_n88# 6.87e-20
C992 a_12036_1467# check[2] 1.58e-19
C993 a_12153_627# a_14096_627# 2.2e-20
C994 x17.X a_12447_n62# 0.00192f
C995 a_8933_1642# x13.X 0.0843f
C996 VDD a_1028_212# 0.687f
C997 x11.X VDD_SW_b[5] 0.24f
C998 VDD_SW[5] a_7733_993# 6.61e-21
C999 D[4] a_8409_n88# 0.00546f
C1000 a_12134_n88# a_12447_n62# 0.245f
C1001 VSS_SW[4] a_8409_n88# 9.92e-21
C1002 D[6] a_3039_601# 0.00583f
C1003 a_2419_627# a_2865_993# 0.159f
C1004 a_7252_1467# D[4] 0.0183f
C1005 a_10596_212# a_12988_212# 1.9e-21
C1006 a_11069_122# a_12134_n88# 8e-21
C1007 a_11313_304# a_11514_n62# 8.99e-19
C1008 a_10597_n88# a_12680_106# 1.67e-21
C1009 x9.A1 a_15907_627# 5.3e-20
C1010 x9.A1 a_14791_1315# 0.00504f
C1011 VDD_SW[2] a_14999_601# 7.64e-20
C1012 a_7252_1467# VSS_SW[4] 0.0274f
C1013 VDD x27.A 0.166f
C1014 check[1] x18.X 5.77e-19
C1015 a_193_627# a_2585_627# 3.26e-19
C1016 a_10597_n88# VSS_SW_b[3] 7.59e-19
C1017 VSS_SW[3] a_11015_220# 6.42e-21
C1018 x14.X D[4] 0.00106f
C1019 a_10801_n88# a_11069_122# 0.206f
C1020 x2.X check[6] 0.193f
C1021 x13.X a_7350_n88# 1.64e-21
C1022 a_5289_1289# a_6285_1642# 0.0146f
C1023 a_13705_304# VSS_SW[1] 6.59e-21
C1024 a_13193_n88# VSS_SW_b[1] 4.54e-20
C1025 x9.A1 a_5812_212# 1.36e-20
C1026 a_4338_n62# a_5812_212# 2.79e-22
C1027 check[5] a_5289_1289# 4.15e-21
C1028 D[2] a_14430_90# 8.78e-19
C1029 a_29_2457# a_76_1467# 1.6e-20
C1030 a_11987_627# a_12433_993# 0.159f
C1031 D[2] a_12607_601# 0.00583f
C1032 x12.X a_5257_993# 1.55e-20
C1033 a_1757_1642# a_2136_627# 5.9e-19
C1034 VDD_SW_b[3] a_12433_993# 8.18e-21
C1035 x11.X a_5504_106# 1.89e-20
C1036 a_15608_993# VDD_SW[1] 3.28e-20
C1037 x2.X a_2879_n62# 0.371f
C1038 a_2419_627# a_3551_627# 0.00272f
C1039 x9.A1 a_4149_1315# 0.00499f
C1040 a_11071_1642# a_10824_993# 0.00176f
C1041 check[3] check[2] 0.00521f
C1042 VDD a_5950_304# 0.0164f
C1043 a_9761_627# a_12341_627# 3.67e-21
C1044 x9.A1 a_9595_627# 8.16e-19
C1045 VDD_SW[7] a_3333_601# 2.55e-20
C1046 x2.X a_10597_n88# 0.0213f
C1047 x30.A check[4] 0.00702f
C1048 VDD a_13705_304# 0.0042f
C1049 a_8933_1642# a_8204_212# 1.17e-22
C1050 ready a_193_627# 6.76e-21
C1051 a_939_2457# a_647_601# 2.7e-21
C1052 a_15293_601# VSS_SW[1] 2.13e-19
C1053 x9.X a_3421_n88# 0.0186f
C1054 VDD a_7394_1642# 0.00177f
C1055 a_6199_895# a_5813_n88# 6.35e-19
C1056 a_5725_601# a_6017_n88# 0.00251f
C1057 a_11987_627# a_14733_627# 4.74e-21
C1058 a_14857_1289# D[2] 5.1e-21
C1059 a_6040_993# a_5812_212# 8.94e-21
C1060 x9.A1 a_13643_1642# 5.26e-19
C1061 a_381_627# a_174_n88# 3.32e-19
C1062 a_1256_993# a_487_n62# 3.59e-19
C1063 a_941_601# a_1028_212# 6.03e-19
C1064 VSS_SW_b[4] a_8921_n62# 6.94e-20
C1065 check[6] a_1369_n62# 9.72e-20
C1066 a_5323_2457# D[5] 0.038f
C1067 a_10073_1289# x15.X 1.7e-20
C1068 a_3807_895# a_4977_627# 2.8e-19
C1069 a_3333_601# a_5431_601# 1.55e-20
C1070 a_939_2457# x9.A1 0.00366f
C1071 a_3807_895# VSS_SW[5] 7.52e-21
C1072 check[4] a_6153_n62# 1.02e-19
C1073 VDD a_15293_601# 0.46f
C1074 a_7203_627# a_8432_993# 0.14f
C1075 D[4] a_8591_895# 0.0294f
C1076 VSS_SW[2] VSS_SW_b[2] 0.00722f
C1077 a_14428_1467# a_14570_1315# 0.00783f
C1078 a_7350_n88# a_8204_212# 0.0319f
C1079 a_7663_n62# a_7896_106# 0.124f
C1080 x9.A1 a_1233_n88# 3.89e-20
C1081 a_14379_627# a_15692_993# 2.13e-19
C1082 check[0] a_15767_895# 0.00271f
C1083 D[1] a_15464_909# 8.49e-19
C1084 a_16037_1642# D[1] 5.74e-19
C1085 a_1028_212# a_2985_n62# 1.09e-19
C1086 VSS_SW[6] a_2566_n88# 0.00677f
C1087 x2.X D[7] 0.252f
C1088 a_5725_601# a_6339_627# 0.0526f
C1089 a_6199_895# a_6920_627# 0.0967f
C1090 x2.X a_8067_909# 0.00138f
C1091 a_5431_601# VDD_SW[5] 2.07e-20
C1092 VDD_SW_b[5] a_5813_n88# 0.0406f
C1093 VDD_SW_b[7] a_720_106# 5.23e-19
C1094 a_14430_90# VSS_SW_b[1] 0.19f
C1095 x9.A1 a_15585_n88# 3.88e-20
C1096 VDD a_1946_n62# 0.109f
C1097 a_9595_627# a_9742_n88# 0.00176f
C1098 a_11325_1642# D[2] 1.73e-19
C1099 a_12036_1467# a_11987_627# 5.32e-19
C1100 VDD_SW_b[6] a_4977_627# 0.00337f
C1101 x8.X a_2610_1315# 8.34e-19
C1102 VDD_SW_b[6] VSS_SW[5] 0.00248f
C1103 check[1] a_13461_122# 6.52e-20
C1104 VDD_SW[3] a_12851_909# 2.16e-20
C1105 x15.X a_12988_212# 1.68e-21
C1106 x2.X a_12638_220# 0.0028f
C1107 D[4] VDD_SW_b[4] 0.454f
C1108 a_7681_1289# D[5] 1.02e-20
C1109 a_16024_909# VDD_SW_b[1] 3.65e-20
C1110 D[4] a_9646_90# 8.78e-19
C1111 x16.X a_10824_993# 2.81e-19
C1112 x2.X a_2419_627# 0.355f
C1113 VDD a_8933_1642# 0.115f
C1114 VDD_SW_b[5] a_6920_627# 0.185f
C1115 a_15855_1642# a_15853_122# 1.57e-21
C1116 a_16109_1642# D[1] 0.061f
C1117 a_13715_1642# a_13643_1642# 6.64e-19
C1118 a_14096_627# a_14379_627# 0.00111f
C1119 VDD_SW_b[2] a_14096_627# 0.185f
C1120 x2.X a_535_1642# 2.63e-19
C1121 a_27_627# VSS_SW[6] 4.66e-21
C1122 x9.A1 a_6529_304# 5.63e-21
C1123 a_5271_n62# a_6017_n88# 0.199f
C1124 a_5504_106# a_5813_n88# 0.0327f
C1125 a_4958_n88# a_6285_122# 4.59e-22
C1126 x8.X a_2470_90# 0.00259f
C1127 VSS_SW[7] a_487_n62# 3.44e-19
C1128 x2.X a_3558_304# 0.00338f
C1129 x9.A1 VSS_SW[2] 0.113f
C1130 a_12901_601# VSS_SW[2] 2.17e-19
C1131 VDD a_7350_n88# 0.69f
C1132 check[2] a_10937_n62# 9.81e-20
C1133 D[1] VDD_SW[1] 0.246f
C1134 a_16330_1315# D[1] 0.0012f
C1135 a_7823_601# a_7663_n62# 0.0026f
C1136 x9.A1 a_10041_993# 1.42e-19
C1137 a_4370_1315# VDD_SW_b[6] 2.65e-20
C1138 a_7649_993# a_7350_n88# 8.71e-20
C1139 a_10509_601# a_12433_993# 1.11e-20
C1140 a_10824_993# a_12153_627# 3.63e-21
C1141 x2.X a_1112_909# 0.00309f
C1142 check[2] a_10215_601# 0.00262f
C1143 x9.A1 x9.X 6.77e-19
C1144 x9.X a_4338_n62# 0.00158f
C1145 a_16109_1642# a_15380_212# 1.17e-22
C1146 a_5257_993# a_5377_n62# 6.88e-22
C1147 a_6199_895# a_6730_n62# 4.06e-19
C1148 VDD a_10908_993# 0.00281f
C1149 a_647_601# a_593_n62# 1.07e-20
C1150 a_6539_1642# D[5] 0.0605f
C1151 VDD_SW_b[2] a_13329_n62# 0.00179f
C1152 D[2] D[1] 0.00183f
C1153 VDD a_6467_1642# 8.63e-19
C1154 x2.X a_5257_993# 0.15f
C1155 x2.X a_4149_1642# 5.23e-19
C1156 check[1] a_12433_993# 7.12e-20
C1157 x9.A1 a_7394_1315# 4.35e-20
C1158 VDD a_439_1315# 9.49e-20
C1159 a_4413_2457# a_4149_1642# 9.92e-19
C1160 a_4689_2457# x9.A1 5.5e-19
C1161 check[2] a_11539_1642# 0.00688f
C1162 VDD x7.X 0.458f
C1163 a_7557_627# VSS_SW_b[4] 5.82e-19
C1164 a_7663_n62# a_8623_220# 1.21e-20
C1165 a_8204_212# a_8153_304# 2.13e-19
C1166 a_7896_106# a_8342_304# 0.00412f
C1167 a_8205_n88# a_7854_220# 4.48e-20
C1168 a_3039_601# a_3283_909# 0.0104f
C1169 a_3807_895# a_3648_993# 0.207f
C1170 a_3333_601# a_2773_627# 1.24e-20
C1171 a_2865_993# a_2949_993# 0.00972f
C1172 a_2585_627# a_3504_909# 0.00907f
C1173 a_3421_n88# a_3625_n88# 0.117f
C1174 a_3112_106# VSS_SW_b[6] 0.00322f
C1175 a_3420_212# a_3893_122# 0.159f
C1176 VSS_SW[6] a_3369_304# 8.28e-20
C1177 a_15767_895# a_15721_n62# 1.65e-20
C1178 VDD_SW[1] a_15380_212# 4.35e-19
C1179 VDD a_13632_909# 0.00438f
C1180 VDD a_12465_1289# 0.191f
C1181 a_15907_627# a_15585_n88# 7.32e-20
C1182 check[6] a_1971_1642# 0.00688f
C1183 a_12038_90# a_12134_n88# 0.0967f
C1184 x2.X a_8539_627# 0.00111f
C1185 VDD_SW[7] VSS_SW[6] 0.429f
C1186 VDD_SW_b[5] a_6730_n62# 0.0145f
C1187 check[0] a_14379_627# 0.00121f
C1188 a_14545_627# a_14999_601# 0.117f
C1189 check[5] a_3947_627# 4.06e-19
C1190 x18.X a_14096_627# 0.0285f
C1191 a_13461_1642# check[0] 2.07e-21
C1192 a_11069_122# a_11514_n62# 0.0369f
C1193 a_9742_n88# VSS_SW[2] 4.18e-21
C1194 x10.X D[6] 9.68e-19
C1195 VDD a_3420_212# 0.687f
C1196 a_10041_993# a_9742_n88# 8.71e-20
C1197 VSS_SW[1] a_14839_n62# 3.44e-19
C1198 x2.X a_5943_627# 0.00702f
C1199 VDD_SW[6] a_5165_627# 6.11e-20
C1200 VSS_SW[3] a_10801_n88# 9.92e-21
C1201 a_8204_212# a_10161_n62# 1.09e-19
C1202 D[2] a_15380_212# 5.78e-20
C1203 VSS_SW_b[4] a_8140_n62# 1.68e-19
C1204 a_11325_1642# a_10983_895# 0.00232f
C1205 x8.X a_1757_1315# 1.78e-20
C1206 a_8409_n88# a_8545_n62# 0.0697f
C1207 a_8205_n88# VSS_SW[3] 9.23e-19
C1208 a_3648_993# VDD_SW_b[6] 4.99e-20
C1209 D[6] D[5] 0.00189f
C1210 a_11325_1642# D[3] 0.0604f
C1211 a_305_2457# x2.X 0.00106f
C1212 a_7369_627# a_7823_601# 0.117f
C1213 x2.X a_11313_304# 3.34e-19
C1214 VDD a_14839_n62# 0.326f
C1215 x2.X a_5289_1289# 0.0112f
C1216 a_5323_2457# a_6285_1642# 0.00184f
C1217 D[1] VSS_SW_b[1] 4.85e-19
C1218 check[0] a_15072_106# 8.65e-22
C1219 a_12036_1467# check[1] 0.318f
C1220 a_5812_212# a_6529_304# 4.45e-20
C1221 a_5271_n62# a_7254_90# 3.67e-21
C1222 a_4958_n88# a_5377_n62# 0.0383f
C1223 a_6017_n88# a_5950_304# 9.46e-19
C1224 a_5813_n88# a_6231_220# 0.00276f
C1225 VSS_SW_b[5] a_5462_220# 5.33e-20
C1226 a_1028_212# VSS_SW_b[7] 0.00119f
C1227 VSS_SW[7] a_1447_220# 6.42e-21
C1228 a_1029_n88# a_1501_122# 0.15f
C1229 VDD_SW_b[4] a_10597_n88# 2.44e-21
C1230 a_9646_90# a_10597_n88# 9.87e-21
C1231 x11.X a_7663_n62# 4.73e-20
C1232 x2.X a_13300_993# 4.66e-19
C1233 x2.X a_4958_n88# 0.178f
C1234 VDD a_8516_993# 0.00281f
C1235 x7.X a_941_601# 1.26e-19
C1236 VDD a_8153_304# 0.00266f
C1237 a_8117_601# a_8288_909# 0.00652f
C1238 a_7823_601# a_7967_627# 0.0697f
C1239 check[6] a_1256_993# 3.41e-19
C1240 a_1971_1642# D[7] 0.00163f
C1241 x10.X a_5725_601# 5e-20
C1242 VDD_SW_b[3] a_10937_n62# 0.00179f
C1243 D[6] VSS_SW_b[6] 5.32e-19
C1244 x9.X a_5812_212# 8.4e-22
C1245 x18.X check[0] 0.009f
C1246 a_10509_601# a_10727_627# 3.73e-19
C1247 a_11123_627# a_11069_122# 2.54e-20
C1248 a_10215_601# VDD_SW_b[3] 1.75e-20
C1249 a_10824_993# a_10359_627# 0.00316f
C1250 x16.X a_12399_1315# 2.4e-19
C1251 a_9595_627# VSS_SW[2] 4.66e-21
C1252 x2.X a_16024_909# 4.02e-19
C1253 a_9761_627# a_10824_993# 0.0334f
C1254 VSS_SW[1] a_15518_304# 1.97e-20
C1255 a_15380_212# VSS_SW_b[1] 0.00119f
C1256 a_15381_n88# a_15853_122# 0.15f
C1257 a_9595_627# a_10041_993# 0.159f
C1258 a_4363_1642# D[6] 0.00163f
C1259 VDD a_10161_n62# 0.0133f
C1260 x9.X a_4149_1315# 2.08e-19
C1261 a_4811_627# a_6199_895# 0.0321f
C1262 D[5] a_5725_601# 0.0192f
C1263 a_2610_1642# VSS_SW[6] 0.00105f
C1264 VDD_SW_b[6] a_4137_n62# 5.22e-19
C1265 a_29_2457# x6.X 2.77e-19
C1266 VDD_SW[2] a_12988_212# 4.35e-19
C1267 a_13515_627# a_13193_n88# 7.32e-20
C1268 a_8067_909# VDD_SW_b[4] 3.61e-21
C1269 x9.A1 a_13216_993# 4.84e-21
C1270 VDD a_193_627# 0.664f
C1271 a_12607_601# a_12517_993# 6.69e-20
C1272 a_12433_993# a_12341_627# 0.0369f
C1273 a_12153_627# a_12851_909# 0.00276f
C1274 a_12901_601# a_13216_993# 0.13f
C1275 a_8731_627# a_8677_122# 2.54e-20
C1276 a_8591_895# a_8545_n62# 1.65e-20
C1277 a_8117_601# VSS_SW[3] 2.9e-20
C1278 a_7896_106# a_9742_n88# 1.86e-21
C1279 x9.A1 a_6539_1315# 0.00496f
C1280 a_3333_601# a_4528_627# 5.73e-19
C1281 x6.X a_381_627# 6.12e-19
C1282 x2.X a_2949_993# 5.29e-19
C1283 x9.A1 a_3625_n88# 3.89e-20
C1284 a_2585_627# VDD_SW[6] 1.96e-20
C1285 x2.X a_11704_627# 3.88e-19
C1286 a_3421_n88# a_4862_90# 5.39e-19
C1287 a_3893_122# a_4137_304# 0.00972f
C1288 a_3112_106# a_3356_n62# 0.00707f
C1289 a_3625_n88# a_4338_n62# 8.07e-20
C1290 a_2879_n62# a_3535_n62# 3.73e-19
C1291 VSS_SW_b[6] a_3839_220# 1.12e-20
C1292 VDD a_15518_304# 0.0164f
C1293 VDD_SW[5] D[4] 4.55e-19
C1294 VDD_SW[5] VSS_SW[4] 0.429f
C1295 VDD_SW_b[5] a_8204_212# 2.29e-22
C1296 x2.X a_720_106# 0.0385f
C1297 VDD a_9786_1642# 0.00177f
C1298 VDD a_4137_304# 0.0042f
C1299 x9.A1 a_7823_601# 2.81e-20
C1300 a_10288_106# a_10532_n62# 0.00707f
C1301 a_10055_n62# a_10711_n62# 3.73e-19
C1302 x9.A1 a_16037_1642# 5.26e-19
C1303 D[5] a_6456_909# 8.07e-19
C1304 a_4811_627# VDD_SW_b[5] 1.12e-19
C1305 a_29_2457# a_27_627# 1.01e-19
C1306 check[1] a_12495_1642# 0.00526f
C1307 D[7] a_2136_627# 0.00238f
C1308 check[5] a_3112_106# 8.68e-22
C1309 a_487_n62# a_678_220# 3.24e-19
C1310 VDD a_791_627# 4.58e-19
C1311 a_7711_1642# D[4] 5.72e-19
C1312 a_27_627# a_381_627# 0.0455f
C1313 D[7] a_1256_993# 0.00608f
C1314 x11.X a_7369_627# 1.68e-19
C1315 check[3] a_7203_627# 0.0012f
C1316 VDD_SW_b[4] a_8545_n62# 0.00179f
C1317 a_9122_n62# VSS_SW[3] 6.09e-20
C1318 a_13461_122# a_13329_n62# 0.025f
C1319 a_13193_n88# VSS_SW[1] 8.41e-20
C1320 VSS_SW_b[2] a_13103_n62# 5.23e-19
C1321 ready VDD_SW[6] 0.00397f
C1322 x8.X a_647_601# 1.98e-20
C1323 a_4860_1467# D[6] 2.91e-19
C1324 D[2] VSS_SW_b[2] 5.22e-19
C1325 check[6] VSS_SW[7] 0.0495f
C1326 a_4860_1467# a_5002_1642# 0.00557f
C1327 a_15293_601# a_15511_627# 3.73e-19
C1328 check[4] a_5431_601# 0.00262f
C1329 a_15608_993# a_15143_627# 0.00316f
C1330 a_14999_601# VDD_SW_b[1] 2.14e-20
C1331 VDD a_6199_895# 0.671f
C1332 a_2773_627# VSS_SW[6] 0.00595f
C1333 a_5725_601# a_8117_601# 9.37e-21
C1334 a_4977_627# a_7557_627# 3.67e-21
C1335 a_6199_895# a_7649_993# 8e-21
C1336 a_2136_627# a_2419_627# 0.0011f
C1337 x12.X a_7681_1289# 1.51e-19
C1338 a_15853_122# a_16298_n62# 0.0369f
C1339 a_15072_106# a_15721_n62# 0.00316f
C1340 a_2468_1467# x7.X 4.97e-19
C1341 a_15380_212# a_15495_n62# 0.00272f
C1342 x9.A1 x8.X 9.17e-19
C1343 VDD a_13193_n88# 0.48f
C1344 a_5813_n88# a_7663_n62# 4.56e-21
C1345 a_5812_212# a_7896_106# 5.96e-20
C1346 a_1256_993# a_2419_627# 7.46e-20
C1347 a_1415_895# D[6] 2.13e-19
C1348 x9.A1 a_16109_1642# 0.195f
C1349 a_487_n62# VSS_SW[6] 1.64e-20
C1350 a_1028_212# a_1143_n62# 0.00272f
C1351 a_720_106# a_1369_n62# 0.00316f
C1352 x2.X a_5761_304# 0.00166f
C1353 a_4811_627# a_5504_106# 3.88e-21
C1354 x17.X a_12988_212# 0.245f
C1355 D[5] a_5271_n62# 0.00258f
C1356 a_193_627# a_941_601# 0.126f
C1357 a_647_601# a_473_993# 0.206f
C1358 a_8432_993# a_8731_627# 0.0256f
C1359 a_8117_601# VDD_SW[4] 1.83e-19
C1360 VDD VDD_SW_b[5] 0.157f
C1361 a_12447_n62# a_12680_106# 0.124f
C1362 a_12134_n88# a_12988_212# 0.0319f
C1363 VDD_SW_b[5] a_7649_993# 8.18e-21
C1364 reset x3.X 0.00166f
C1365 x9.A1 a_473_993# 1.42e-19
C1366 a_14428_1467# a_14887_1642# 6.64e-19
C1367 a_9644_1467# D[4] 2.78e-19
C1368 a_5927_n62# a_6153_n62# 3.34e-19
C1369 x9.A1 VDD_SW[1] 0.0323f
C1370 a_10055_n62# VSS_SW_b[2] 9.32e-21
C1371 VDD_SW_b[7] D[6] 1.53e-19
C1372 a_10597_n88# a_12989_n88# 1.33e-19
C1373 VDD_SW[2] a_15293_601# 2.55e-20
C1374 a_10215_601# a_10509_601# 0.199f
C1375 x16.X a_11546_1315# 5.02e-20
C1376 a_11069_122# VSS_SW_b[3] 7.15e-19
C1377 a_941_601# a_791_627# 0.00926f
C1378 a_193_627# a_1672_909# 7.17e-20
C1379 a_647_601# a_1159_627# 9.75e-19
C1380 a_1256_993# a_1112_909# 0.00412f
C1381 a_473_993# a_581_627# 0.00807f
C1382 check[5] D[6] 0.465f
C1383 a_8848_909# VDD_SW[4] 2.12e-20
C1384 a_14430_90# VSS_SW[1] 0.0819f
C1385 D[7] VSS_SW[7] 0.134f
C1386 x2.X a_3947_627# 0.0151f
C1387 x9.A1 D[2] 0.267f
C1388 D[2] a_12901_601# 0.0191f
C1389 a_2879_n62# VSS_SW_b[5] 1.09e-20
C1390 a_6539_1642# x12.X 7.67e-19
C1391 a_11987_627# a_13375_895# 0.0321f
C1392 a_3421_n88# a_5813_n88# 1.33e-19
C1393 a_505_1289# a_473_993# 4.54e-19
C1394 x2.X a_12447_n62# 0.371f
C1395 x9.A1 x11.X 7.59e-19
C1396 check[2] VDD_SW_b[3] 0.0022f
C1397 a_3039_601# a_3420_212# 4.51e-19
C1398 a_2865_993# a_3112_106# 4.96e-20
C1399 x2.X a_1745_304# 3.34e-19
C1400 a_11253_1642# D[3] 5.74e-19
C1401 a_3333_601# a_2879_n62# 3.74e-20
C1402 a_2585_627# a_3421_n88# 1.27e-19
C1403 x2.X a_11069_122# 0.0043f
C1404 VDD a_5504_106# 0.356f
C1405 VDD a_14430_90# 0.189f
C1406 VDD a_12607_601# 0.313f
C1407 a_14857_1289# VSS_SW[1] 0.00186f
C1408 VDD a_8861_1642# 8.63e-19
C1409 x9.A1 a_1503_1642# 0.101f
C1410 a_12851_909# VDD_SW_b[2] 2.4e-21
C1411 x9.A1 a_5165_627# 4.11e-19
C1412 a_4977_627# VSS_SW[5] 0.0232f
C1413 D[4] a_9761_627# 5.14e-21
C1414 a_5323_2457# x2.X 0.00627f
C1415 a_4413_2457# a_5323_2457# 2.64e-19
C1416 VDD a_14857_1289# 0.191f
C1417 a_12680_106# a_13126_304# 0.00412f
C1418 a_12447_n62# a_13407_220# 1.21e-20
C1419 a_12989_n88# a_12638_220# 4.71e-20
C1420 a_12988_212# a_12937_304# 2.13e-19
C1421 VDD a_15608_993# 0.189f
C1422 VDD_SW_b[6] a_2566_n88# 3.21e-19
C1423 a_6285_1642# a_5725_601# 0.00263f
C1424 a_6920_627# a_7369_627# 5.39e-19
C1425 a_505_1289# a_1503_1642# 0.0146f
C1426 a_14379_627# a_14933_627# 0.00206f
C1427 check[0] a_15855_1642# 0.257f
C1428 x9.A1 a_10055_n62# 1.54e-20
C1429 D[3] VSS_SW_b[2] 2.05e-19
C1430 VSS_SW_b[5] a_6529_n62# 6.93e-20
C1431 a_7254_90# a_7350_n88# 0.0967f
C1432 x17.X a_15293_601# 4.31e-21
C1433 VDD a_3504_909# 0.0164f
C1434 a_1447_220# VSS_SW[6] 1.57e-20
C1435 a_1028_212# VSS_SW_b[6] 0.00377f
C1436 VDD_SW[4] a_10125_993# 6.61e-21
C1437 D[7] a_3333_601# 2.67e-21
C1438 a_5725_601# a_5675_909# 1.21e-20
C1439 a_4977_627# a_5575_627# 6.04e-20
C1440 D[5] a_5950_304# 9.69e-19
C1441 a_5575_627# VSS_SW[5] 0.0012f
C1442 x9.A1 VSS_SW_b[1] 2.86e-19
C1443 a_13715_1642# D[2] 0.0607f
C1444 VDD a_1029_n88# 0.66f
C1445 x2.X a_13126_304# 0.00338f
C1446 VDD_SW[5] a_8067_909# 2.16e-20
C1447 x2.X a_7681_1289# 0.0113f
C1448 VDD a_11325_1642# 0.115f
C1449 D[4] a_8677_122# 0.00928f
C1450 a_7203_627# VSS_SW_b[4] 1.08e-19
C1451 VSS_SW[4] a_8677_122# 2.79e-21
C1452 a_2419_627# a_3333_601# 0.14f
C1453 D[6] a_2865_993# 0.00884f
C1454 a_13632_909# VDD_SW[2] 2.12e-20
C1455 a_939_2457# x8.X 8.68e-19
C1456 x2.X a_14999_601# 0.2f
C1457 x13.X a_7663_n62# 0.00192f
C1458 a_9742_n88# a_10055_n62# 0.245f
C1459 VDD_SW[6] a_4811_627# 0.0865f
C1460 x9.A1 a_5813_n88# 8.59e-21
C1461 a_3558_304# VSS_SW_b[5] 9.9e-21
C1462 a_4338_n62# a_5813_n88# 3.67e-21
C1463 a_4862_90# a_5812_212# 1.66e-20
C1464 x3.A a_76_1467# 2.66e-20
C1465 x9.A1 a_2585_627# 3.23e-19
C1466 x12.X a_5725_601# 0.00124f
C1467 a_11325_1642# a_10596_212# 1.17e-22
C1468 x11.X a_5812_212# 0.245f
C1469 VDD_SW_b[3] a_11987_627# 5.95e-19
C1470 a_11704_627# VDD_SW[3] 0.0729f
C1471 a_11123_627# a_10931_627# 4.19e-20
C1472 x2.X a_3112_106# 0.0385f
C1473 D[6] a_3551_627# 6.12e-19
C1474 x9.A1 a_10983_895# 2.64e-19
C1475 a_10983_895# a_12901_601# 1.38e-20
C1476 VDD a_6231_220# 0.00984f
C1477 x9.A1 D[3] 0.269f
C1478 check[2] a_10509_601# 2.09e-19
C1479 VDD_SW[7] a_3807_895# 1.27e-20
C1480 D[3] a_12901_601# 2.67e-21
C1481 a_7681_1289# a_8679_1642# 0.0146f
C1482 a_9595_627# D[2] 1.19e-20
C1483 x9.A1 a_3895_1642# 0.101f
C1484 ready a_647_601# 3.47e-22
C1485 x9.X a_3625_n88# 1.8e-19
C1486 x9.A1 a_6920_627# 2.14e-20
C1487 a_305_2457# VSS_SW[7] 0.0177f
C1488 D[1] VSS_SW[1] 0.133f
C1489 a_5725_601# a_6285_122# 2.7e-19
C1490 a_6199_895# a_6017_n88# 4.26e-19
C1491 VDD a_2610_1315# 4.95e-19
C1492 a_941_601# a_1029_n88# 3.89e-19
C1493 x2.X a_6539_1642# 5.27e-19
C1494 a_1415_895# a_1028_212# 0.00165f
C1495 a_193_627# VSS_SW_b[7] 5.23e-20
C1496 x9.A1 a_8933_1315# 0.00499f
C1497 a_13643_1642# D[2] 5.74e-19
C1498 check[1] a_13375_895# 0.00266f
C1499 check[2] check[1] 0.0052f
C1500 check[6] VSS_SW[6] 1.39e-19
C1501 a_4149_1642# a_3333_601# 7.12e-21
C1502 a_3648_993# a_4977_627# 3.63e-21
C1503 a_3333_601# a_5257_993# 1.11e-20
C1504 ready x9.A1 3.55e-19
C1505 check[4] D[4] 3.66e-20
C1506 check[4] VSS_SW[4] 1.4e-19
C1507 D[4] a_8432_993# 0.00608f
C1508 a_7203_627# a_7557_627# 0.0455f
C1509 VDD D[1] 0.767f
C1510 VDD a_12178_1642# 0.00177f
C1511 a_7350_n88# a_8205_n88# 0.0477f
C1512 a_7663_n62# a_8204_212# 0.138f
C1513 VDD_SW_b[7] a_3283_909# 2.1e-21
C1514 x9.A1 a_1501_122# 4.39e-20
C1515 a_11514_n62# a_12988_212# 5.58e-22
C1516 VDD VDD_SW[6] 0.39f
C1517 a_1946_n62# VSS_SW_b[6] 2.63e-19
C1518 VSS_SW[6] a_2879_n62# 3.44e-19
C1519 a_14999_601# a_14825_993# 0.206f
C1520 a_14545_627# a_15293_601# 0.126f
C1521 x2.X a_8288_909# 0.00309f
C1522 a_6199_895# a_6339_627# 0.0383f
C1523 a_5257_993# VDD_SW[5] 4.17e-21
C1524 a_5725_601# a_6147_627# 1.96e-20
C1525 a_12465_1289# x17.X 1.79e-20
C1526 D[5] a_7350_n88# 4.26e-19
C1527 x2.X a_7854_220# 0.00279f
C1528 VDD_SW_b[5] a_6017_n88# 0.00133f
C1529 a_9761_627# a_10597_n88# 1.27e-19
C1530 VDD_SW_b[7] a_1028_212# 0.0416f
C1531 x13.X a_7369_627# 1.02e-20
C1532 VSS_SW[1] a_15380_212# 1.18e-21
C1533 VDD a_2470_90# 0.189f
C1534 a_939_2457# a_1503_1642# 0.00188f
C1535 ready a_505_1289# 2.39e-20
C1536 VSS_SW[3] VSS_SW_b[3] 0.0075f
C1537 a_9595_627# a_10055_n62# 7.27e-19
C1538 D[3] a_9742_n88# 0.00507f
C1539 D[7] a_678_220# 1.98e-20
C1540 VDD_SW_b[6] a_5431_601# 2.23e-20
C1541 a_12465_1289# a_12134_n88# 5.67e-21
C1542 a_1503_1642# a_1233_n88# 4.63e-19
C1543 x2.X D[6] 0.199f
C1544 a_6467_1642# D[5] 5.74e-19
C1545 x2.X a_10459_909# 0.00138f
C1546 x2.X a_12038_90# 0.00366f
C1547 a_4413_2457# D[6] 0.0191f
C1548 VDD a_15380_212# 0.686f
C1549 a_8933_1642# a_8117_601# 7.12e-21
C1550 x2.X VSS_SW[3] 0.086f
C1551 check[0] a_15381_n88# 2.51e-20
C1552 a_14428_1467# check[1] 1.57e-19
C1553 x17.X a_14839_n62# 4.41e-20
C1554 check[3] a_8731_627# 4.05e-19
C1555 a_11325_1642# x15.X 0.0847f
C1556 a_9312_627# a_10509_601# 1.84e-20
C1557 D[7] VSS_SW[6] 4.85e-19
C1558 x9.A1 a_6730_n62# 1.56e-20
C1559 a_5812_212# a_5813_n88# 0.784f
C1560 a_5271_n62# a_6285_122# 0.0633f
C1561 a_5504_106# a_6017_n88# 0.00189f
C1562 a_4958_n88# VSS_SW_b[5] 0.134f
C1563 x2.X a_12541_627# 3.94e-19
C1564 x30.A a_4977_627# 1.19e-21
C1565 VSS_SW[7] a_720_106# 4.63e-19
C1566 a_78_90# a_1028_212# 1.66e-20
C1567 x30.A VSS_SW[5] 0.0445f
C1568 a_12447_n62# a_14526_n88# 5.13e-21
C1569 x2.X a_3839_220# 9.61e-19
C1570 VDD a_7663_n62# 0.326f
C1571 D[2] VSS_SW[2] 0.134f
C1572 a_7369_627# a_8204_212# 1.02e-19
C1573 a_8117_601# a_7350_n88# 0.00259f
C1574 a_7649_993# a_7663_n62# 2.63e-19
C1575 a_7823_601# a_7896_106# 1.01e-19
C1576 x2.X a_1340_993# 4.67e-19
C1577 a_10509_601# a_11987_627# 3.81e-19
C1578 a_9949_627# a_10149_627# 3.81e-19
C1579 a_10509_601# VDD_SW_b[3] 0.00636f
C1580 a_10983_895# a_11240_909# 0.00869f
C1581 a_10824_993# a_10727_627# 0.00386f
C1582 a_2419_627# VSS_SW[6] 0.0576f
C1583 x9.X a_4862_90# 0.0273f
C1584 D[3] a_11240_909# 8.07e-19
C1585 a_4811_627# a_7369_627# 1.09e-20
C1586 a_4977_627# a_7203_627# 1.36e-20
C1587 a_15585_n88# VSS_SW_b[1] 9.21e-19
C1588 a_6920_627# a_5812_212# 6.63e-19
C1589 a_6539_1642# a_7252_1467# 0.00957f
C1590 a_9595_627# a_10983_895# 0.0321f
C1591 VDD a_10711_n62# 0.00521f
C1592 a_1415_895# a_1946_n62# 4.06e-19
C1593 a_9595_627# D[3] 0.138f
C1594 a_473_993# a_593_n62# 6.88e-22
C1595 x7.X VSS_SW_b[6] 0.0172f
C1596 x2.X a_5725_601# 0.119f
C1597 a_12607_601# a_13072_909# 9.46e-19
C1598 check[1] a_11987_627# 0.00121f
C1599 x9.A1 x13.X 6.78e-19
C1600 x16.X a_11704_627# 0.0286f
C1601 a_7203_627# a_9312_627# 1.75e-19
C1602 x2.X a_10931_627# 0.00111f
C1603 a_8204_212# a_8342_304# 1.09e-19
C1604 VDD a_16097_304# 0.0042f
C1605 a_3039_601# a_3504_909# 9.46e-19
C1606 a_939_2457# a_2585_627# 4.92e-21
C1607 VSS_SW[6] a_3558_304# 1.97e-20
C1608 a_3421_n88# a_3893_122# 0.15f
C1609 a_3420_212# VSS_SW_b[6] 0.00119f
C1610 a_76_1467# a_174_n88# 6.87e-20
C1611 x2.X VDD_SW[4] 0.0327f
C1612 VDD a_11253_1642# 8.63e-19
C1613 VDD_SW_b[5] a_7254_90# 0.00346f
C1614 a_10596_212# a_10711_n62# 0.00272f
C1615 a_10055_n62# VSS_SW[2] 1.46e-20
C1616 VDD_SW_b[7] a_1946_n62# 0.0144f
C1617 a_10288_106# a_10937_n62# 0.00316f
C1618 VDD a_3421_n88# 0.66f
C1619 check[1] a_13929_1642# 0.00688f
C1620 a_10215_601# a_10288_106# 1.01e-19
C1621 x2.X a_6456_909# 4.03e-19
C1622 a_10041_993# a_10055_n62# 2.63e-19
C1623 a_9147_1642# D[4] 0.00163f
C1624 VDD_SW[6] a_5341_993# 6.61e-21
C1625 a_12988_212# a_13705_n62# 0.00206f
C1626 VSS_SW_b[4] a_8319_n62# 5.24e-19
C1627 a_8677_122# a_8545_n62# 0.025f
C1628 a_8409_n88# VSS_SW[3] 8.81e-20
C1629 VDD a_7369_627# 0.659f
C1630 x3.X x2.X 0.00477f
C1631 a_11704_627# a_12153_627# 5.39e-19
C1632 a_2468_1467# a_2610_1315# 0.00783f
C1633 a_7369_627# a_7649_993# 0.15f
C1634 a_939_2457# ready 0.262f
C1635 a_14733_627# a_14933_627# 3.81e-19
C1636 a_15767_895# a_16024_909# 0.00869f
C1637 x20.X a_15293_601# 1.31e-19
C1638 a_15293_601# VDD_SW_b[1] 0.00622f
C1639 a_15608_993# a_15511_627# 0.00386f
C1640 a_11071_1642# a_11069_122# 1.57e-21
C1641 a_15585_n88# a_15495_n62# 9.75e-19
C1642 a_15380_212# a_16097_n62# 0.00206f
C1643 a_15381_n88# a_15721_n62# 6.04e-20
C1644 VSS_SW_b[1] a_14945_n62# 0.00335f
C1645 x14.X VSS_SW[3] 0.251f
C1646 x13.X a_9742_n88# 0.00862f
C1647 VDD VSS_SW_b[2] 0.0969f
C1648 a_14545_627# a_14839_n62# 2.38e-19
C1649 x9.A1 a_8204_212# 1.41e-20
C1650 a_14999_601# a_14526_n88# 4.37e-19
C1651 a_5813_n88# a_6529_304# 0.0018f
C1652 a_6017_n88# a_6231_220# 0.0104f
C1653 a_5812_212# a_6730_n62# 0.0453f
C1654 a_5271_n62# a_5377_n62# 0.0526f
C1655 x9.A1 a_13515_627# 5.03e-20
C1656 a_1029_n88# VSS_SW_b[7] 7.59e-19
C1657 x2.X a_15030_220# 0.0028f
C1658 a_1233_n88# a_1501_122# 0.206f
C1659 x17.X a_13193_n88# 1.81e-19
C1660 a_12607_601# VDD_SW[2] 2.07e-20
C1661 a_12901_601# a_13515_627# 0.0526f
C1662 a_13375_895# a_14096_627# 0.0967f
C1663 a_29_2457# check[6] 7.65e-19
C1664 x9.A1 a_4811_627# 8.11e-19
C1665 VDD a_7967_627# 1.8e-19
C1666 check[6] a_1555_627# 4.05e-19
C1667 x2.X a_5271_n62# 0.373f
C1668 VDD a_8342_304# 0.0164f
C1669 x7.X a_1415_895# 0.00659f
C1670 x2.X a_10073_1289# 0.0112f
C1671 a_7369_627# a_8335_627# 2.14e-20
C1672 a_8117_601# a_8516_993# 9.41e-19
C1673 a_7649_993# a_7967_627# 0.025f
C1674 a_7557_627# a_7733_993# 8.99e-19
C1675 a_2468_1467# a_2470_90# 1e-19
C1676 a_12447_n62# a_12989_n88# 0.125f
C1677 a_12680_106# a_12988_212# 0.14f
C1678 a_2566_n88# a_3070_220# 0.00869f
C1679 a_16109_1642# a_16037_1642# 6.64e-19
C1680 a_10983_895# VSS_SW[2] 7.52e-21
C1681 a_10596_212# VSS_SW_b[2] 0.0038f
C1682 VDD_SW[2] a_15608_993# 1.08e-20
C1683 D[3] VSS_SW[2] 4.86e-19
C1684 x9.X a_2585_627# 1.07e-20
C1685 a_10215_601# a_10824_993# 0.00189f
C1686 D[3] a_10041_993# 0.00884f
C1687 D[5] a_6199_895# 0.0294f
C1688 a_4811_627# a_6040_993# 0.14f
C1689 x7.X VDD_SW_b[7] 0.242f
C1690 x9.A1 VSS_SW[1] 0.113f
C1691 a_13375_895# a_13329_n62# 1.65e-20
C1692 VDD a_647_601# 0.314f
C1693 a_12901_601# VSS_SW[1] 2.72e-20
C1694 a_8288_909# VDD_SW_b[4] 9.38e-21
C1695 a_7967_627# a_8335_627# 3.34e-19
C1696 a_3895_1642# x9.X 1.34e-19
C1697 a_8591_895# VSS_SW[3] 7.03e-21
C1698 D[2] a_13216_993# 0.00608f
C1699 a_11987_627# a_12341_627# 0.0455f
C1700 x9.A1 a_3893_122# 4.39e-20
C1701 a_3807_895# a_4528_627# 0.0967f
C1702 x2.X a_3283_909# 0.00137f
C1703 a_3039_601# VDD_SW[6] 2.07e-20
C1704 a_8204_212# a_9742_n88# 6.15e-19
C1705 a_3333_601# a_3947_627# 0.0526f
C1706 VDD_SW_b[3] a_12341_627# 9.3e-21
C1707 x2.X a_12988_212# 0.0126f
C1708 a_15464_909# VDD_SW[1] 2.82e-20
C1709 x7.X check[5] 5.61e-19
C1710 a_2566_n88# VSS_SW[5] 4.18e-21
C1711 a_3112_106# a_3535_n62# 0.00386f
C1712 a_2879_n62# a_3761_n62# 0.00926f
C1713 a_3893_122# a_4338_n62# 0.0369f
C1714 x11.X a_6539_1315# 1.97e-19
C1715 VDD_SW_b[5] a_8205_n88# 2.44e-21
C1716 x13.X a_9595_627# 0.00295f
C1717 x14.X VDD_SW[4] 0.308f
C1718 x2.X a_1028_212# 0.0128f
C1719 VDD x9.A1 4.51f
C1720 VDD a_12901_601# 0.46f
C1721 VDD_SW_b[7] a_3420_212# 4.59e-22
C1722 VDD a_4338_n62# 0.109f
C1723 x9.A1 a_7649_993# 1.48e-19
C1724 a_14570_1642# VSS_SW[1] 0.00105f
C1725 D[5] VDD_SW_b[5] 0.453f
C1726 VDD a_5002_1315# 4.95e-19
C1727 VDD_SW_b[4] a_10459_909# 3.15e-21
C1728 x9.A1 a_11325_1315# 0.00496f
C1729 D[7] a_1555_627# 0.00431f
C1730 x17.X a_14430_90# 0.0273f
C1731 check[5] a_3420_212# 3.24e-20
C1732 VDD a_581_627# 1.28e-19
C1733 a_27_627# a_557_993# 4.45e-20
C1734 D[7] a_381_627# 0.161f
C1735 check[3] D[4] 0.462f
C1736 VDD_SW_b[4] VSS_SW[3] 0.00248f
C1737 a_7369_627# a_9949_627# 3.67e-21
C1738 check[3] VSS_SW[4] 0.0367f
C1739 VDD_SW_b[6] a_4528_627# 0.186f
C1740 a_9646_90# VSS_SW[3] 0.082f
C1741 a_218_1315# VSS_SW[7] 7.95e-19
C1742 x8.X a_473_993# 1.55e-20
C1743 x27.A x2.X 2.91e-19
C1744 a_12988_212# a_13407_220# 2.46e-19
C1745 a_12447_n62# a_13906_n62# 3.79e-20
C1746 VDD a_14570_1642# 0.00177f
C1747 VDD a_14909_993# 0.0042f
C1748 a_12989_n88# a_13126_304# 0.00907f
C1749 VDD a_505_1289# 0.192f
C1750 ready a_4689_2457# 0.00228f
C1751 a_4413_2457# x27.A 0.129f
C1752 a_12153_627# a_12447_n62# 2.38e-19
C1753 a_12607_601# a_12134_n88# 4.37e-19
C1754 a_16109_1642# VDD_SW[1] 0.00494f
C1755 a_16109_1642# a_16330_1315# 0.00783f
C1756 check[4] a_5257_993# 6.52e-20
C1757 a_4149_1642# check[4] 1.58e-19
C1758 VDD a_6040_993# 0.189f
C1759 x9.A1 a_10596_212# 1.41e-20
C1760 a_10459_909# VDD_SW[3] 1.01e-20
C1761 check[0] a_14887_1642# 0.00526f
C1762 a_1757_1642# a_1978_1315# 0.00783f
C1763 D[1] a_15511_627# 6.11e-19
C1764 a_6199_895# a_8117_601# 1.38e-20
C1765 a_1555_627# a_2419_627# 1.09e-19
C1766 a_2136_627# D[6] 4.35e-19
C1767 check[2] a_10288_106# 8.14e-22
C1768 x9.A1 a_8921_304# 6.89e-21
C1769 a_9761_627# a_11704_627# 2e-20
C1770 a_5813_n88# a_7896_106# 1.67e-21
C1771 a_5812_212# a_8204_212# 9.5e-22
C1772 a_6285_122# a_7350_n88# 8e-21
C1773 a_6529_304# a_6730_n62# 8.99e-19
C1774 VDD_SW[4] a_10680_909# 2.77e-20
C1775 a_1028_212# a_1369_n62# 0.00134f
C1776 a_720_106# VSS_SW[6] 9.06e-21
C1777 a_5323_2457# VDD_SW[5] 0.0154f
C1778 a_1029_n88# a_1143_n62# 2.14e-20
C1779 x2.X a_5950_304# 0.00334f
C1780 a_4811_627# a_5812_212# 6.99e-20
C1781 D[5] a_5504_106# 8.77e-19
C1782 a_193_627# a_1415_895# 0.0494f
C1783 a_647_601# a_941_601# 0.199f
C1784 VDD a_9742_n88# 0.69f
C1785 a_11987_627# a_14096_627# 1.75e-19
C1786 a_8432_993# a_8539_627# 0.00707f
C1787 a_8591_895# VDD_SW[4] 0.00356f
C1788 x15.X VSS_SW_b[2] 0.0171f
C1789 x2.X a_13705_304# 3.38e-19
C1790 x14.X a_10073_1289# 1.5e-19
C1791 VDD a_13715_1642# 0.115f
C1792 VDD_SW_b[5] a_8117_601# 5.19e-20
C1793 a_1503_1642# x8.X 1.14e-20
C1794 x9.A1 a_941_601# 0.00103f
C1795 VDD_SW_b[1] a_14839_n62# 5.21e-19
C1796 x20.X a_14839_n62# 0.002f
C1797 a_14428_1467# check[0] 0.318f
C1798 VDD_SW[2] D[1] 4.41e-19
C1799 x2.X a_15293_601# 0.119f
C1800 a_1256_993# a_1340_993# 0.00857f
C1801 a_193_627# VDD_SW_b[7] 0.0022f
C1802 VDD_SW_b[4] VDD_SW[4] 3.64e-19
C1803 check[4] a_5289_1289# 0.247f
C1804 a_9742_n88# a_10596_212# 0.0319f
C1805 a_12924_n62# a_13329_n62# 2.46e-21
C1806 x2.X a_3755_627# 0.00111f
C1807 VDD a_15907_627# 6.88e-19
C1808 x9.A1 a_11313_n62# 5.47e-21
C1809 x9.A1 a_9949_627# 4.11e-19
C1810 a_10509_601# a_12341_627# 2.42e-20
C1811 a_10983_895# a_13216_993# 1.86e-21
C1812 x18.X a_13936_1315# 3.11e-20
C1813 a_3039_601# a_3421_n88# 0.00322f
C1814 a_3333_601# a_3112_106# 3.46e-19
C1815 x2.X a_1946_n62# 1.87e-19
C1816 a_3807_895# a_2879_n62# 0.00219f
C1817 a_2585_627# a_3625_n88# 8.75e-19
C1818 check[2] a_10824_993# 3.41e-19
C1819 check[4] a_4958_n88# 5.26e-19
C1820 VDD a_5812_212# 0.687f
C1821 VDD a_12553_n62# 0.0133f
C1822 x9.A1 a_2927_1642# 5.26e-19
C1823 x9.A1 a_16097_n62# 5.47e-21
C1824 a_76_1467# x6.X 0.0876f
C1825 VDD a_11240_909# 0.00438f
C1826 a_3895_1642# a_3625_n88# 4.63e-19
C1827 a_4977_627# a_5431_601# 0.117f
C1828 a_12178_1315# VSS_SW[2] 7.96e-19
C1829 x2.X a_8933_1642# 5.21e-19
C1830 a_5431_601# VSS_SW[5] 6.28e-19
C1831 VDD a_9595_627# 0.393f
C1832 x9.A1 x15.X 6.84e-19
C1833 x15.X a_12901_601# 4.02e-21
C1834 VDD_SW_b[6] a_2879_n62# 5.22e-19
C1835 a_6285_1642# a_6199_895# 5.55e-19
C1836 VDD a_13643_1642# 8.63e-19
C1837 a_29_2457# a_305_2457# 0.00202f
C1838 a_11015_220# VSS_SW_b[2] 4.16e-21
C1839 a_10596_212# a_12553_n62# 1.09e-19
C1840 a_12038_90# a_12989_n88# 9.87e-21
C1841 a_76_1467# a_27_627# 5.32e-19
C1842 a_14857_1289# a_14545_627# 0.00323f
C1843 a_14545_627# a_15608_993# 0.0334f
C1844 a_7254_90# a_7663_n62# 4.24e-20
C1845 a_14825_993# a_15293_601# 0.0633f
C1846 a_6539_1642# VDD_SW[5] 0.00492f
C1847 x17.X D[1] 2.04e-19
C1848 VDD a_3732_993# 0.00281f
C1849 x3.X a_1256_993# 9.79e-21
C1850 a_593_n62# a_964_n62# 4.19e-20
C1851 VDD_SW_b[3] a_10288_106# 5.24e-19
C1852 a_1745_304# VSS_SW[6] 6.59e-21
C1853 a_1029_n88# VSS_SW_b[6] 0.00485f
C1854 VDD a_939_2457# 1.37f
C1855 a_5431_601# a_5575_627# 0.0697f
C1856 a_5725_601# a_5896_909# 0.00652f
C1857 a_14526_n88# a_15030_220# 0.00869f
C1858 a_9949_627# a_9742_n88# 3.32e-19
C1859 D[5] a_6231_220# 7.13e-19
C1860 x2.X a_7350_n88# 0.178f
C1861 a_5365_627# VSS_SW[5] 3.8e-19
C1862 VSS_SW[1] a_15585_n88# 9.92e-21
C1863 a_9595_627# a_10596_212# 6.99e-20
C1864 a_2897_1289# a_2566_n88# 5.67e-21
C1865 x8.X a_2585_627# 0.00315f
C1866 x9.A1 a_2468_1467# 0.197f
C1867 D[2] VSS_SW_b[1] 2.02e-19
C1868 VDD a_1233_n88# 0.48f
C1869 a_27_627# a_174_n88# 0.00176f
C1870 a_12465_1289# a_12680_106# 5.3e-21
C1871 VDD_SW_b[2] a_12447_n62# 5.22e-19
C1872 a_7252_1467# a_7394_1642# 0.00557f
C1873 D[6] VSS_SW_b[5] 2.03e-19
C1874 x16.X a_12038_90# 0.00259f
C1875 x8.X a_3895_1642# 1.98e-20
C1876 VDD_SW[5] a_8288_909# 2.77e-20
C1877 x2.X a_10908_993# 4.67e-19
C1878 D[4] VSS_SW_b[4] 5.32e-19
C1879 VDD a_15585_n88# 0.48f
C1880 x15.X a_9742_n88# 1.53e-21
C1881 a_2419_627# a_3807_895# 0.0321f
C1882 D[6] a_3333_601# 0.019f
C1883 VSS_SW[4] VSS_SW_b[4] 0.0072f
C1884 x9.X a_4811_627# 0.00299f
C1885 x10.X VDD_SW[6] 0.305f
C1886 check[0] a_15853_122# 6.43e-20
C1887 x2.X a_439_1315# 3.2e-19
C1888 a_5675_909# VDD_SW_b[5] 3.01e-21
C1889 x17.X a_15380_212# 1.68e-21
C1890 a_76_1467# a_218_1642# 0.00557f
C1891 x2.X x7.X 0.0046f
C1892 ready x8.X 2.31e-20
C1893 x13.X a_7896_106# 2.38e-20
C1894 VDD_SW[6] D[5] 4.59e-19
C1895 x9.A1 a_6017_n88# 3.88e-20
C1896 x2.X a_12465_1289# 0.0112f
C1897 x2.X a_13632_909# 4.01e-19
C1898 a_3420_212# a_5377_n62# 1.09e-19
C1899 a_3839_220# VSS_SW_b[5] 3.96e-21
C1900 a_4862_90# a_5813_n88# 9.87e-21
C1901 a_4689_2457# a_4811_627# 3.76e-19
C1902 a_12988_212# a_14526_n88# 6.15e-19
C1903 x12.X a_6199_895# 0.00864f
C1904 x9.A1 a_3039_601# 2.81e-20
C1905 x11.X a_5813_n88# 0.0189f
C1906 x2.X a_3420_212# 0.0127f
C1907 a_2419_627# VDD_SW_b[6] 1.12e-19
C1908 D[6] a_4064_909# 8.06e-19
C1909 VDD a_6529_304# 0.0042f
C1910 VDD_SW[7] a_3648_993# 1.08e-20
C1911 a_10824_993# a_11987_627# 7.46e-20
C1912 a_10983_895# D[2] 2.17e-19
C1913 a_10824_993# VDD_SW_b[3] 5e-20
C1914 D[3] D[2] 0.00189f
C1915 a_939_2457# a_941_601# 2.13e-20
C1916 ready a_473_993# 7.59e-22
C1917 x9.X a_3893_122# 2.77e-19
C1918 x3.X VSS_SW[7] 0.0128f
C1919 a_9595_627# a_9949_627# 0.0455f
C1920 x9.A1 a_6339_627# 5.12e-20
C1921 VDD VSS_SW[2] 0.523f
C1922 a_2136_627# a_1028_212# 6.63e-19
C1923 check[3] a_8545_n62# 9.72e-20
C1924 a_6040_993# a_6017_n88# 1.86e-19
C1925 a_6199_895# a_6285_122# 4.53e-22
C1926 VDD a_10041_993# 0.18f
C1927 check[1] a_13329_n62# 1.04e-19
C1928 a_1256_993# a_1028_212# 8.94e-21
C1929 a_1415_895# a_1029_n88# 6.35e-19
C1930 a_941_601# a_1233_n88# 0.00251f
C1931 a_8933_1642# x14.X 8.08e-19
C1932 x2.X a_14839_n62# 0.371f
C1933 a_12901_601# a_13072_909# 0.00652f
C1934 a_12607_601# a_12751_627# 0.0697f
C1935 VDD x9.X 0.458f
C1936 x11.X a_6920_627# 0.0338f
C1937 x12.X VDD_SW_b[5] 7.21e-19
C1938 a_3807_895# a_5257_993# 8e-21
C1939 a_4149_1642# a_3807_895# 0.00232f
C1940 a_2585_627# a_5165_627# 3.67e-21
C1941 a_3333_601# a_5725_601# 9.37e-21
C1942 a_10073_1289# a_11071_1642# 0.0146f
C1943 a_9786_1315# D[3] 7.54e-19
C1944 a_7203_627# a_7733_993# 4.45e-20
C1945 D[4] a_7557_627# 0.161f
C1946 VDD a_14945_n62# 0.0133f
C1947 a_7557_627# VSS_SW[4] 0.00595f
C1948 x15.X a_9595_627# 2.67e-20
C1949 a_7663_n62# a_8205_n88# 0.125f
C1950 a_7896_106# a_8204_212# 0.14f
C1951 x9.A1 VSS_SW_b[7] 2.86e-19
C1952 VDD_SW_b[7] a_3504_909# 1.97e-21
C1953 VSS_SW[6] a_3112_106# 4.63e-19
C1954 a_2470_90# VSS_SW_b[6] 0.19f
C1955 a_4363_1642# VDD_SW[6] 5.38e-19
C1956 VDD a_7394_1315# 4.95e-19
C1957 a_7252_1467# a_7350_n88# 6.87e-20
C1958 a_6040_993# a_6339_627# 0.0256f
C1959 x2.X a_8516_993# 4.67e-19
C1960 D[1] a_14545_627# 0.168f
C1961 a_5725_601# VDD_SW[5] 1.79e-19
C1962 a_14379_627# a_14999_601# 0.149f
C1963 VDD a_4689_2457# 0.359f
C1964 x9.A1 a_13715_1315# 0.00499f
C1965 x2.X a_8153_304# 0.00166f
C1966 a_10597_n88# a_10937_n62# 6.04e-20
C1967 a_10801_n88# a_10711_n62# 9.75e-19
C1968 check[1] check[0] 0.00509f
C1969 VDD_SW_b[5] a_6285_122# 0.00447f
C1970 VSS_SW_b[3] a_10161_n62# 0.00335f
C1971 VDD_SW_b[2] a_14999_601# 1.99e-20
C1972 a_10596_212# VSS_SW[2] 0.0872f
C1973 a_10983_895# a_10055_n62# 0.00219f
C1974 a_10509_601# a_10288_106# 3.46e-19
C1975 VDD_SW_b[7] a_1029_n88# 0.0406f
C1976 a_10215_601# a_10597_n88# 0.00322f
C1977 check[2] D[4] 6.03e-20
C1978 VDD a_593_n62# 0.0138f
C1979 D[3] a_10055_n62# 0.00258f
C1980 ready a_1503_1642# 9.79e-21
C1981 a_4149_1642# VDD_SW_b[6] 2.59e-19
C1982 VDD_SW_b[6] a_5257_993# 8.2e-21
C1983 a_1503_1642# a_1501_122# 1.57e-21
C1984 a_6539_1642# a_6753_1642# 0.00557f
C1985 x2.X a_10161_n62# 5.57e-20
C1986 a_15608_993# VDD_SW_b[1] 5.61e-20
C1987 a_9644_1467# VSS_SW[3] 0.0274f
C1988 a_14857_1289# x20.X 1.7e-20
C1989 a_6456_909# VDD_SW[5] 2.12e-20
C1990 a_8933_1642# a_8591_895# 0.00232f
C1991 a_5323_2457# check[4] 0.0505f
C1992 x2.X a_193_627# 0.0537f
C1993 a_15853_122# a_15721_n62# 0.025f
C1994 VSS_SW_b[1] a_15495_n62# 5.24e-19
C1995 a_15293_601# a_14526_n88# 0.00259f
C1996 a_14999_601# a_15072_106# 1.01e-19
C1997 a_14825_993# a_14839_n62# 2.63e-19
C1998 a_14545_627# a_15380_212# 1.02e-19
C1999 x2.X a_15518_304# 0.00338f
C2000 x9.A1 VDD_SW[2] 0.0329f
C2001 a_13216_993# a_13515_627# 0.0256f
C2002 a_4860_1467# VDD_SW[6] 0.00487f
C2003 a_12901_601# VDD_SW[2] 1.75e-19
C2004 a_5271_n62# VSS_SW_b[5] 0.0142f
C2005 a_5812_212# a_6017_n88# 0.15f
C2006 VSS_SW[5] a_5462_220# 4.26e-19
C2007 VSS_SW[7] a_1028_212# 5.9e-22
C2008 a_78_90# a_1029_n88# 9.87e-21
C2009 a_1978_1315# D[7] 0.0012f
C2010 x30.A a_5431_601# 7.99e-20
C2011 a_939_2457# a_2468_1467# 0.0011f
C2012 x11.X a_6730_n62# 0.00162f
C2013 x2.X a_4137_304# 3.38e-19
C2014 VDD a_7896_106# 0.356f
C2015 a_8117_601# a_7663_n62# 3.74e-20
C2016 a_8933_1642# VDD_SW_b[4] 2.6e-19
C2017 a_7369_627# a_8205_n88# 1.27e-19
C2018 a_12447_n62# a_13461_122# 0.0633f
C2019 a_7823_601# a_8204_212# 4.51e-19
C2020 a_12680_106# a_13193_n88# 0.00189f
C2021 a_12988_212# a_12989_n88# 0.785f
C2022 a_7649_993# a_7896_106# 4.96e-20
C2023 a_12134_n88# VSS_SW_b[2] 0.135f
C2024 x2.X a_791_627# 0.0388f
C2025 D[6] VSS_SW[6] 0.134f
C2026 x18.X a_14999_601# 2.4e-20
C2027 VDD_SW[2] a_14909_993# 6.61e-21
C2028 a_10801_n88# VSS_SW_b[2] 5.04e-20
C2029 D[5] a_7369_627# 6.4e-21
C2030 a_10041_993# a_9949_627# 0.0369f
C2031 a_10509_601# a_10824_993# 0.13f
C2032 a_9761_627# a_10459_909# 0.00276f
C2033 a_6339_627# a_5812_212# 7.07e-21
C2034 a_4977_627# VSS_SW[4] 5.07e-21
C2035 check[4] a_7681_1289# 4.13e-21
C2036 a_10359_627# VSS_SW[3] 0.0012f
C2037 D[3] a_10983_895# 0.0294f
C2038 a_9761_627# VSS_SW[3] 0.023f
C2039 x2.X a_6199_895# 0.148f
C2040 a_4528_627# a_4977_627# 5.39e-19
C2041 VDD_SW_b[6] a_4958_n88# 5.91e-19
C2042 a_4528_627# VSS_SW[5] 0.00162f
C2043 D[2] a_12517_993# 8.11e-19
C2044 a_11987_627# a_12851_909# 2.46e-19
C2045 D[4] a_9312_627# 0.00232f
C2046 VDD_SW_b[3] a_12851_909# 2.62e-21
C2047 x15.X VSS_SW[2] 0.148f
C2048 VDD_SW_b[4] a_7350_n88# 3.21e-19
C2049 x2.X a_13193_n88# 0.00372f
C2050 a_9644_1467# VDD_SW[4] 0.00484f
C2051 a_3333_601# a_3283_909# 1.21e-20
C2052 a_8205_n88# a_8342_304# 0.00907f
C2053 a_7663_n62# a_9122_n62# 3.79e-20
C2054 a_8204_212# a_8623_220# 2.46e-19
C2055 a_2585_627# a_3183_627# 6.04e-20
C2056 a_3625_n88# a_3893_122# 0.206f
C2057 ready a_2585_627# 9.49e-21
C2058 a_3421_n88# VSS_SW_b[6] 7.59e-19
C2059 VSS_SW[6] a_3839_220# 6.42e-21
C2060 a_15316_n62# a_15721_n62# 2.46e-21
C2061 VDD_SW_b[5] a_5377_n62# 4.78e-19
C2062 VDD a_13216_993# 0.189f
C2063 check[5] VDD_SW[6] 0.00393f
C2064 VDD_SW_b[7] a_2470_90# 0.00345f
C2065 a_13715_1642# VDD_SW[2] 0.00502f
C2066 VDD a_3625_n88# 0.48f
C2067 a_12178_1315# D[2] 7.54e-19
C2068 ready a_3895_1642# 4.05e-20
C2069 x9.A1 x17.X 6.87e-19
C2070 x2.X VDD_SW_b[5] 7.37e-19
C2071 VDD_SW[6] a_5675_909# 2.16e-20
C2072 x17.X a_12901_601# 1.26e-19
C2073 check[5] a_2470_90# 2.5e-20
C2074 a_174_n88# a_487_n62# 0.245f
C2075 VDD a_7823_601# 0.313f
C2076 a_8677_122# VSS_SW[3] 6.66e-20
C2077 VSS_SW_b[4] a_8545_n62# 5.35e-19
C2078 a_12988_212# a_13906_n62# 0.0453f
C2079 VDD a_16037_1642# 8.63e-19
C2080 VDD a_15464_909# 0.0164f
C2081 x9.A1 a_12134_n88# 7.4e-19
C2082 a_12989_n88# a_13705_304# 0.0018f
C2083 a_13193_n88# a_13407_220# 0.0104f
C2084 a_12433_993# a_12447_n62# 2.63e-19
C2085 a_12607_601# a_12680_106# 1.01e-19
C2086 a_12153_627# a_12988_212# 1.02e-19
C2087 a_12901_601# a_12134_n88# 0.00259f
C2088 a_7369_627# a_8117_601# 0.126f
C2089 a_7823_601# a_7649_993# 0.206f
C2090 x6.X a_27_627# 0.236f
C2091 a_6539_1642# check[4] 0.318f
C2092 a_10359_627# a_10931_627# 2.46e-21
C2093 x20.X D[1] 0.101f
C2094 x9.A1 a_10801_n88# 3.88e-20
C2095 check[0] a_16323_1642# 0.00688f
C2096 D[1] VDD_SW_b[1] 0.454f
C2097 x9.A1 x10.X 9.2e-19
C2098 check[2] a_10597_n88# 2.47e-20
C2099 x13.X a_10055_n62# 4.41e-20
C2100 x10.X a_5002_1315# 8.34e-19
C2101 x9.A1 a_8205_n88# 8.52e-21
C2102 a_5504_106# a_5377_n62# 0.0256f
C2103 a_5271_n62# a_5748_n62# 1.96e-20
C2104 a_6017_n88# a_6529_304# 6.69e-20
C2105 a_5812_212# a_7254_90# 0.00102f
C2106 VSS_SW_b[5] a_5950_304# 3.57e-20
C2107 a_5813_n88# a_6730_n62# 0.189f
C2108 VDD_SW[4] a_9761_627# 9.25e-19
C2109 a_1233_n88# VSS_SW_b[7] 9.21e-19
C2110 x3.A check[6] 9.84e-19
C2111 x7.X a_2136_627# 0.0338f
C2112 x9.A1 D[5] 0.324f
C2113 D[2] a_13515_627# 0.00431f
C2114 x11.X a_8204_212# 8.4e-22
C2115 x2.X a_5504_106# 0.0385f
C2116 a_4811_627# a_4862_90# 6.13e-19
C2117 x2.X a_14430_90# 0.00368f
C2118 VDD a_8623_220# 0.00984f
C2119 a_7369_627# a_8848_909# 7.17e-20
C2120 a_8432_993# a_8288_909# 0.00412f
C2121 a_8117_601# a_7967_627# 0.00926f
C2122 a_5002_1315# D[5] 7.54e-19
C2123 a_7823_601# a_8335_627# 9.75e-19
C2124 x2.X a_12607_601# 0.2f
C2125 a_7649_993# a_7757_627# 0.00807f
C2126 VDD x8.X 0.338f
C2127 x11.X a_4811_627# 2.67e-20
C2128 VDD a_16109_1642# 0.111f
C2129 a_2879_n62# a_3070_220# 3.3e-19
C2130 x20.X a_15380_212# 0.245f
C2131 VDD_SW_b[1] a_15380_212# 0.0417f
C2132 a_11015_220# VSS_SW[2] 1.76e-20
C2133 a_13715_1642# x17.X 0.0841f
C2134 check[4] D[6] 5.94e-20
C2135 x2.X a_14857_1289# 0.0112f
C2136 x2.X a_15608_993# 0.187f
C2137 D[5] a_6040_993# 0.00609f
C2138 a_4811_627# a_5165_627# 0.0455f
C2139 check[4] a_5002_1642# 0.00688f
C2140 a_14526_n88# a_14839_n62# 0.245f
C2141 VDD a_473_993# 0.181f
C2142 D[2] VSS_SW[1] 4.85e-19
C2143 a_13705_304# a_13906_n62# 8.99e-19
C2144 VDD a_16330_1315# 3.48e-19
C2145 VDD VDD_SW[1] 0.358f
C2146 a_8204_212# a_10055_n62# 2.62e-19
C2147 a_8205_n88# a_9742_n88# 1.98e-19
C2148 x2.X a_3504_909# 0.0031f
C2149 a_3333_601# a_3755_627# 1.96e-20
C2150 a_3807_895# a_3947_627# 0.0383f
C2151 a_2865_993# VDD_SW[6] 4.17e-21
C2152 x9.A1 VSS_SW_b[6] 2.86e-19
C2153 a_2879_n62# VSS_SW[5] 1.64e-20
C2154 a_3112_106# a_3761_n62# 0.00316f
C2155 reset x9.A1 3.51e-20
C2156 a_3420_212# a_3535_n62# 0.00272f
C2157 a_10073_1289# a_9761_627# 0.00323f
C2158 VDD a_13103_n62# 0.00521f
C2159 x13.X D[3] 2.06e-19
C2160 x2.X a_1029_n88# 0.0213f
C2161 VDD_SW_b[7] a_3421_n88# 2.44e-21
C2162 VDD a_4862_90# 0.189f
C2163 x9.A1 a_8117_601# 0.00103f
C2164 VDD D[2] 0.77f
C2165 x3.A D[7] 1.17e-20
C2166 x9.A1 a_14545_627# 3.23e-19
C2167 a_27_627# VDD_SW[7] 3.29e-20
C2168 D[7] a_1363_627# 2e-19
C2169 a_12901_601# a_14545_627# 5.92e-20
C2170 check[5] a_3421_n88# 2.51e-20
C2171 VDD x11.X 0.458f
C2172 VDD a_1159_627# 7.51e-19
C2173 a_487_n62# a_1166_304# 0.00652f
C2174 a_720_106# a_977_304# 0.00857f
C2175 x2.X a_11325_1642# 5.18e-19
C2176 a_27_627# a_891_909# 2.46e-19
C2177 D[7] a_557_993# 8.11e-19
C2178 a_11546_1315# VDD_SW_b[3] 3.97e-20
C2179 D[4] a_10509_601# 3.09e-21
C2180 a_8140_n62# a_8545_n62# 2.46e-21
C2181 x13.X a_8933_1315# 2.09e-19
C2182 x8.X a_941_601# 0.00123f
C2183 a_12134_n88# a_12553_n62# 0.0383f
C2184 VDD a_1503_1642# 0.191f
C2185 VDD a_9786_1315# 4.95e-19
C2186 check[4] a_5725_601# 2.03e-19
C2187 a_11514_n62# VSS_SW_b[2] 2.8e-19
C2188 VDD a_5165_627# 0.109f
C2189 a_14857_1289# a_14825_993# 4.54e-19
C2190 a_15293_601# a_15767_895# 0.265f
C2191 a_14545_627# a_14909_993# 0.0018f
C2192 a_14999_601# a_14733_627# 8.07e-20
C2193 x9.A1 a_9122_n62# 1.9e-20
C2194 VDD_SW_b[3] a_10597_n88# 0.0406f
C2195 a_5812_212# a_8205_n88# 5.48e-21
C2196 a_5813_n88# a_8204_212# 4.92e-22
C2197 a_7615_1315# D[4] 0.00202f
C2198 a_1029_n88# a_1369_n62# 6.04e-20
C2199 a_1028_212# VSS_SW[6] 0.0872f
C2200 VSS_SW_b[7] a_593_n62# 0.00335f
C2201 a_1233_n88# a_1143_n62# 9.75e-19
C2202 a_193_627# a_2136_627# 2.2e-20
C2203 a_9595_627# a_10801_n88# 0.00204f
C2204 VSS_SW[1] VSS_SW_b[1] 0.00717f
C2205 x10.X a_4149_1315# 1.78e-20
C2206 x2.X a_6231_220# 9.51e-19
C2207 D[5] a_5812_212# 0.157f
C2208 a_4811_627# a_5813_n88# 1.06e-19
C2209 x9.A1 a_4860_1467# 0.197f
C2210 a_193_627# a_1256_993# 0.0334f
C2211 a_473_993# a_941_601# 0.0633f
C2212 VDD a_10055_n62# 0.326f
C2213 a_8432_993# VDD_SW[4] 3.28e-20
C2214 VDD_SW_b[2] a_12988_212# 0.0416f
C2215 a_13461_1642# a_12988_212# 1.39e-21
C2216 a_4860_1467# a_5002_1315# 0.00783f
C2217 a_2585_627# a_4811_627# 1.36e-20
C2218 a_2419_627# a_4977_627# 1.09e-20
C2219 a_2419_627# VSS_SW[5] 4.66e-21
C2220 x2.X a_10149_627# 3.99e-19
C2221 VDD VSS_SW_b[1] 0.0968f
C2222 a_7203_627# D[4] 0.138f
C2223 a_7203_627# VSS_SW[4] 0.0576f
C2224 x9.A1 a_1415_895# 2.64e-19
C2225 a_891_909# VDD_SW[7] 1.01e-20
C2226 a_76_1467# check[6] 0.318f
C2227 a_4811_627# a_6920_627# 1.75e-19
C2228 a_1256_993# a_791_627# 0.00316f
C2229 a_941_601# a_1159_627# 3.73e-19
C2230 a_647_601# VDD_SW_b[7] 1.36e-20
C2231 x16.X a_12465_1289# 1.54e-19
C2232 x7.X a_3333_601# 4.31e-21
C2233 x2.X D[1] 0.197f
C2234 a_10055_n62# a_10596_212# 0.138f
C2235 x12.X a_7369_627# 0.00315f
C2236 a_9122_n62# a_9742_n88# 8.26e-21
C2237 a_12989_n88# a_14839_n62# 4.56e-21
C2238 a_12988_212# a_15072_106# 5.86e-20
C2239 x2.X VDD_SW[6] 0.0327f
C2240 a_3420_212# VSS_SW_b[5] 0.00377f
C2241 a_4413_2457# VDD_SW[6] 0.0115f
C2242 a_3558_304# VSS_SW[5] 2.76e-20
C2243 a_1503_1642# a_941_601# 0.00263f
C2244 check[6] a_174_n88# 5.27e-19
C2245 x9.A1 a_11514_n62# 1.9e-20
C2246 x9.A1 VDD_SW_b[7] 2.34e-20
C2247 a_3648_993# a_2879_n62# 3.59e-19
C2248 a_2773_627# a_2566_n88# 3.32e-19
C2249 x2.X a_2470_90# 0.00368f
C2250 a_3333_601# a_3420_212# 6.03e-19
C2251 x9.A1 a_6285_1642# 0.101f
C2252 check[4] a_5271_n62# 1.31e-20
C2253 VDD a_5813_n88# 0.66f
C2254 check[3] a_7681_1289# 0.249f
C2255 a_2468_1467# x8.X 0.0876f
C2256 x9.A1 check[5] 0.412f
C2257 a_8933_1642# a_9644_1467# 0.00963f
C2258 VDD a_2585_627# 0.659f
C2259 a_487_n62# a_2566_n88# 5.13e-21
C2260 a_3895_1642# a_3893_122# 1.57e-21
C2261 VDD a_10983_895# 0.671f
C2262 a_4977_627# a_5257_993# 0.15f
C2263 a_5257_993# VSS_SW[5] 0.003f
C2264 VDD D[3] 0.771f
C2265 x2.X a_15380_212# 0.0122f
C2266 a_12607_601# a_13119_627# 9.75e-19
C2267 a_12465_1289# a_12153_627# 0.00323f
C2268 a_12433_993# a_12541_627# 0.00807f
C2269 a_12153_627# a_13632_909# 7.17e-20
C2270 a_12901_601# a_12751_627# 0.00926f
C2271 a_13216_993# a_13072_909# 0.00412f
C2272 a_193_627# VSS_SW[7] 0.023f
C2273 a_8117_601# a_9595_627# 3.84e-19
C2274 x15.X D[2] 2.14e-19
C2275 a_7663_n62# VSS_SW_b[3] 1.03e-20
C2276 VDD a_3895_1642# 0.191f
C2277 a_11325_1315# D[3] 0.00195f
C2278 VDD a_15495_n62# 0.00521f
C2279 VDD a_6920_627# 0.194f
C2280 VDD_SW_b[6] a_3112_106# 5.23e-19
C2281 a_6285_1642# a_6040_993# 0.00181f
C2282 check[6] a_2897_1289# 3.63e-21
C2283 VSS_SW[2] a_12134_n88# 0.00676f
C2284 x3.A a_305_2457# 0.3f
C2285 a_29_2457# x3.X 6.66e-19
C2286 reset a_939_2457# 4.31e-19
C2287 check[0] a_15721_n62# 9.72e-20
C2288 a_76_1467# D[7] 0.0183f
C2289 a_6730_n62# a_8204_212# 2.79e-22
C2290 a_14379_627# a_15293_601# 0.14f
C2291 D[1] a_14825_993# 0.00887f
C2292 x9.A1 x20.X 5.49e-19
C2293 a_11069_122# a_10937_n62# 0.025f
C2294 a_1946_n62# VSS_SW[6] 6.09e-20
C2295 VSS_SW_b[3] a_10711_n62# 5.24e-19
C2296 a_10801_n88# VSS_SW[2] 8.39e-20
C2297 x9.A1 VDD_SW_b[1] 2.35e-20
C2298 a_1233_n88# VSS_SW_b[6] 4.54e-20
C2299 VDD a_3183_627# 1.8e-19
C2300 VDD_SW_b[2] a_15293_601# 8.35e-20
C2301 VDD ready 0.64f
C2302 a_27_627# a_2773_627# 4.46e-21
C2303 a_5165_627# a_5341_993# 8.99e-19
C2304 a_4977_627# a_5943_627# 2.14e-20
C2305 a_5257_993# a_5575_627# 0.025f
C2306 a_5725_601# a_6124_993# 9.41e-19
C2307 a_10509_601# a_10597_n88# 3.89e-19
C2308 a_10983_895# a_10596_212# 0.00165f
C2309 x2.X a_7663_n62# 0.373f
C2310 D[5] a_6529_304# 8.39e-19
C2311 D[3] a_10596_212# 0.158f
C2312 x8.X a_3039_601# 2.4e-20
C2313 a_2897_1289# a_2879_n62# 3.44e-19
C2314 a_791_627# VSS_SW[7] 0.0012f
C2315 VSS_SW_b[2] a_13705_n62# 6.93e-20
C2316 a_14430_90# a_14526_n88# 0.0967f
C2317 x9.X x10.X 0.111f
C2318 VDD a_1501_122# 0.313f
C2319 D[7] a_174_n88# 0.00506f
C2320 a_27_627# a_487_n62# 7.27e-19
C2321 a_12036_1467# a_12038_90# 1e-19
C2322 a_6539_1642# check[3] 1.64e-19
C2323 x9.A1 a_11123_627# 5.3e-20
C2324 VDD_SW[3] a_12607_601# 7.64e-20
C2325 a_4149_1642# a_4370_1315# 0.00783f
C2326 x9.A1 x12.X 0.00118f
C2327 a_5289_1289# a_4977_627# 0.00323f
C2328 x15.X a_10055_n62# 0.002f
C2329 a_2419_627# a_3648_993# 0.14f
C2330 D[6] a_3807_895# 0.0294f
C2331 a_5289_1289# VSS_SW[5] 0.00187f
C2332 x9.X D[5] 2.11e-19
C2333 VSS_SW_b[1] a_16097_n62# 6.94e-20
C2334 a_4689_2457# x10.X 9.8e-19
C2335 a_5896_909# VDD_SW_b[5] 7.05e-21
C2336 x2.X a_1757_1315# 2.32e-19
C2337 a_5575_627# a_5943_627# 3.34e-19
C2338 a_9147_1642# VDD_SW[4] 5.38e-19
C2339 a_76_1467# a_535_1642# 6.64e-19
C2340 a_14999_601# a_15381_n88# 0.00322f
C2341 a_15767_895# a_14839_n62# 0.00219f
C2342 a_14857_1289# a_14526_n88# 5.67e-21
C2343 a_14545_627# a_15585_n88# 8.75e-19
C2344 a_15293_601# a_15072_106# 3.46e-19
C2345 a_941_601# a_2585_627# 6.03e-20
C2346 x2.X a_16097_304# 3.38e-19
C2347 x13.X a_8204_212# 0.245f
C2348 a_13216_993# VDD_SW[2] 3.28e-20
C2349 a_4977_627# a_4958_n88# 4.91e-19
C2350 x9.A1 a_6285_122# 4.73e-20
C2351 VSS_SW[5] a_4958_n88# 0.00686f
C2352 a_2897_1289# D[7] 5.1e-21
C2353 x12.X a_6040_993# 2.81e-19
C2354 a_1757_1642# VDD_SW[7] 0.00511f
C2355 x9.A1 a_2865_993# 1.48e-19
C2356 x11.X a_6017_n88# 1.87e-19
C2357 a_12680_106# VSS_SW_b[2] 0.00322f
C2358 a_12989_n88# a_13193_n88# 0.117f
C2359 D[6] VDD_SW_b[6] 0.453f
C2360 x2.X a_3421_n88# 0.0207f
C2361 VSS_SW[2] a_12937_304# 8.24e-20
C2362 a_12988_212# a_13461_122# 0.159f
C2363 VDD a_6730_n62# 0.109f
C2364 a_6285_1642# a_5812_212# 1.39e-21
C2365 VDD_SW[7] a_2773_627# 6.11e-20
C2366 x18.X a_15293_601# 4.9e-20
C2367 VDD_SW[2] a_15464_909# 2.77e-20
C2368 a_2831_1315# D[6] 0.00202f
C2369 a_1028_212# a_1745_n62# 0.00206f
C2370 a_939_2457# a_1415_895# 0.00134f
C2371 a_9595_627# a_10125_993# 4.45e-20
C2372 D[3] a_9949_627# 0.161f
C2373 x2.X a_7369_627# 0.0537f
C2374 a_1555_627# a_1028_212# 7.07e-21
C2375 check[3] VSS_SW[3] 1.4e-19
C2376 a_5575_627# a_4958_n88# 1.08e-19
C2377 a_6040_993# a_6285_122# 1.51e-20
C2378 x9.A1 a_13705_n62# 5.7e-21
C2379 VDD a_10545_304# 0.00266f
C2380 a_2897_1289# a_2419_627# 0.00104f
C2381 a_941_601# a_1501_122# 2.7e-19
C2382 a_1415_895# a_1233_n88# 4.26e-19
C2383 x7.X VSS_SW[6] 0.148f
C2384 a_8342_304# VSS_SW_b[3] 8.9e-21
C2385 a_11325_1642# VDD_SW[3] 0.00506f
C2386 a_8117_601# a_10041_993# 1.29e-20
C2387 D[2] a_13072_909# 8.51e-19
C2388 a_3807_895# a_5725_601# 1.38e-20
C2389 a_11987_627# a_13300_993# 2.13e-19
C2390 x2.X VSS_SW_b[2] 0.0278f
C2391 a_7203_627# a_8067_909# 2.46e-19
C2392 D[4] a_7733_993# 8.11e-19
C2393 x15.X a_10983_895# 0.0066f
C2394 x15.X D[3] 0.1f
C2395 a_7663_n62# a_8409_n88# 0.199f
C2396 a_7896_106# a_8205_n88# 0.0327f
C2397 a_7350_n88# a_8677_122# 4.59e-22
C2398 a_939_2457# VDD_SW_b[7] 1.96e-20
C2399 VSS_SW[6] a_3420_212# 1.18e-21
C2400 VDD a_12517_993# 0.0042f
C2401 a_6040_993# a_6147_627# 0.00707f
C2402 a_15143_627# VSS_SW[1] 0.0012f
C2403 x2.X a_7967_627# 0.0388f
C2404 a_6199_895# VDD_SW[5] 0.00356f
C2405 VDD x13.X 0.458f
C2406 x2.X a_8342_304# 0.00334f
C2407 a_13715_1315# D[2] 0.00195f
C2408 a_10055_n62# a_11015_220# 1.21e-20
C2409 a_10288_106# a_10734_304# 0.00412f
C2410 a_10596_212# a_10545_304# 2.13e-19
C2411 VDD_SW_b[7] a_1233_n88# 0.00132f
C2412 a_10597_n88# a_10246_220# 4.48e-20
C2413 a_12465_1289# a_13461_1642# 0.0146f
C2414 a_939_2457# check[5] 0.00134f
C2415 a_13632_909# VDD_SW_b[2] 3.14e-20
C2416 VDD a_964_n62# 8.23e-19
C2417 D[7] a_1166_304# 9.67e-19
C2418 VDD_SW_b[6] a_5725_601# 5.2e-20
C2419 a_12989_n88# a_14430_90# 5.39e-19
C2420 a_305_2457# a_76_1467# 1.82e-20
C2421 a_13461_122# a_13705_304# 0.00972f
C2422 VSS_SW_b[2] a_13407_220# 1.2e-20
C2423 a_13193_n88# a_13906_n62# 8.07e-20
C2424 VDD a_12178_1315# 4.95e-19
C2425 VDD a_15143_627# 1.8e-19
C2426 a_12607_601# a_12989_n88# 0.00322f
C2427 a_12901_601# a_12680_106# 3.46e-19
C2428 a_12153_627# a_13193_n88# 8.75e-19
C2429 a_13375_895# a_12447_n62# 0.00219f
C2430 a_11704_627# a_11987_627# 0.0011f
C2431 VDD_SW_b[3] a_11704_627# 0.185f
C2432 a_4860_1467# x9.X 4.97e-19
C2433 x9.A1 VSS_SW_b[3] 2.86e-19
C2434 VDD_SW_b[5] VDD_SW[5] 3.63e-19
C2435 check[2] a_11069_122# 6.44e-20
C2436 x2.X a_647_601# 0.2f
C2437 x13.X a_10596_212# 8.4e-22
C2438 check[3] VDD_SW[4] 0.00393f
C2439 D[1] a_14526_n88# 0.00508f
C2440 a_14379_627# a_14839_n62# 7.27e-19
C2441 a_5813_n88# a_6017_n88# 0.117f
C2442 VSS_SW[5] a_5761_304# 8.37e-20
C2443 a_5812_212# a_6285_122# 0.159f
C2444 a_5504_106# VSS_SW_b[5] 0.00321f
C2445 a_9644_1467# a_9786_1642# 0.00557f
C2446 D[2] VDD_SW[2] 0.246f
C2447 VSS_SW[7] a_1029_n88# 9.29e-21
C2448 x30.A a_5257_993# 5.04e-19
C2449 a_4689_2457# a_4860_1467# 0.00106f
C2450 x16.X a_12607_601# 2.69e-20
C2451 x2.X x9.A1 0.659f
C2452 a_6539_1315# D[5] 0.00195f
C2453 x2.X a_12901_601# 0.119f
C2454 D[4] a_10288_106# 1.39e-21
C2455 x11.X a_7254_90# 0.0273f
C2456 a_4413_2457# x9.A1 1.84e-19
C2457 x2.X a_4338_n62# 1.9e-19
C2458 VDD a_8204_212# 0.687f
C2459 a_7823_601# a_8205_n88# 0.00322f
C2460 a_8117_601# a_7896_106# 3.46e-19
C2461 a_7369_627# a_8409_n88# 8.75e-19
C2462 a_8591_895# a_7663_n62# 0.00219f
C2463 VDD a_13515_627# 6.99e-19
C2464 x2.X a_581_627# 3.94e-19
C2465 a_2585_627# a_3039_601# 0.117f
C2466 x20.X a_15585_n88# 1.87e-19
C2467 VDD_SW_b[1] a_15585_n88# 0.00131f
C2468 a_2566_n88# a_2879_n62# 0.245f
C2469 VDD a_4811_627# 0.393f
C2470 a_11514_n62# VSS_SW[2] 6.06e-20
C2471 a_1946_n62# a_1745_n62# 3.81e-19
C2472 x6.X check[6] 0.00903f
C2473 a_10041_993# a_10125_993# 0.00972f
C2474 a_10215_601# a_10459_909# 0.0104f
C2475 D[3] a_11015_220# 7.13e-19
C2476 x2.X a_14909_993# 5.31e-19
C2477 x14.X a_7369_627# 6.29e-20
C2478 a_193_627# VSS_SW[6] 5.36e-21
C2479 a_14526_n88# a_15380_212# 0.0319f
C2480 a_14839_n62# a_15072_106# 0.124f
C2481 x2.X a_505_1289# 0.0112f
C2482 check[4] a_6467_1642# 0.00577f
C2483 a_9742_n88# VSS_SW_b[3] 0.135f
C2484 a_10215_601# VSS_SW[3] 6.23e-19
C2485 x2.X a_6040_993# 0.187f
C2486 check[5] x9.X 0.00967f
C2487 D[4] a_8731_627# 0.00431f
C2488 a_8204_212# a_10596_212# 9.5e-22
C2489 a_12751_627# VSS_SW[2] 0.0012f
C2490 a_12153_627# a_12607_601# 0.117f
C2491 VDD_SW_b[4] a_7663_n62# 5.22e-19
C2492 a_8409_n88# a_8342_304# 9.46e-19
C2493 VSS_SW_b[4] a_7854_220# 5.34e-20
C2494 x9.A1 a_8679_1642# 0.101f
C2495 a_7663_n62# a_9646_90# 6.12e-21
C2496 a_7350_n88# a_7769_n62# 0.0383f
C2497 a_8205_n88# a_8623_220# 0.00276f
C2498 a_8204_212# a_8921_304# 4.45e-20
C2499 check[6] a_27_627# 0.00121f
C2500 a_3039_601# a_3183_627# 0.0697f
C2501 a_3333_601# a_3504_909# 0.00652f
C2502 check[3] a_10073_1289# 3.63e-21
C2503 ready a_3039_601# 7.34e-21
C2504 a_3625_n88# VSS_SW_b[6] 9.21e-19
C2505 VDD VSS_SW[1] 0.522f
C2506 x30.A a_5289_1289# 0.00187f
C2507 VDD_SW_b[5] a_5748_n62# 8.12e-20
C2508 x2.X a_9742_n88# 0.178f
C2509 VDD_SW_b[7] a_593_n62# 4.77e-19
C2510 VDD a_3893_122# 0.313f
C2511 D[7] a_2566_n88# 4.33e-19
C2512 a_11325_1642# x16.X 7.78e-19
C2513 x9.A1 a_14825_993# 1.42e-19
C2514 a_12901_601# a_14825_993# 1.11e-20
C2515 VDD_SW[6] a_5896_909# 2.77e-20
C2516 a_13216_993# a_14545_627# 4.03e-21
C2517 x2.X a_13715_1642# 5.28e-19
C2518 x17.X D[2] 0.1f
C2519 a_174_n88# a_720_106# 0.207f
C2520 a_5323_2457# a_4977_627# 7.32e-19
C2521 a_5323_2457# VSS_SW[5] 0.0134f
C2522 a_12447_n62# a_12924_n62# 1.96e-20
C2523 a_12680_106# a_12553_n62# 0.0256f
C2524 a_3283_909# VDD_SW_b[6] 3.01e-21
C2525 VDD a_7649_993# 0.18f
C2526 a_7823_601# a_8117_601# 0.199f
C2527 a_7369_627# a_8591_895# 0.0494f
C2528 x6.X D[7] 0.00886f
C2529 D[2] a_12134_n88# 0.00506f
C2530 x27.A a_3807_895# 7.61e-21
C2531 a_11987_627# a_12447_n62# 7.27e-19
C2532 VDD_SW_b[1] a_14945_n62# 4.77e-19
C2533 check[6] a_218_1642# 0.00688f
C2534 a_14545_627# a_15464_909# 0.00907f
C2535 a_15855_1642# a_15293_601# 0.00263f
C2536 a_14999_601# a_15243_909# 0.0104f
C2537 a_15767_895# a_15608_993# 0.207f
C2538 a_15293_601# a_14733_627# 1.24e-20
C2539 a_14825_993# a_14909_993# 0.00972f
C2540 a_2419_627# a_2566_n88# 0.00176f
C2541 a_10509_601# a_11704_627# 5.73e-19
C2542 x10.X a_4862_90# 0.00259f
C2543 VDD_SW_b[3] a_11069_122# 0.00446f
C2544 x2.X a_15907_627# 0.0151f
C2545 x2.X a_14791_1315# 3.2e-19
C2546 a_9154_1315# D[4] 0.0012f
C2547 a_15380_212# a_15329_304# 2.13e-19
C2548 a_14839_n62# a_15799_220# 1.21e-20
C2549 a_15381_n88# a_15030_220# 4.71e-20
C2550 a_15072_106# a_15518_304# 0.00412f
C2551 x9.A1 a_8409_n88# 3.88e-20
C2552 a_5271_n62# a_5927_n62# 3.73e-19
C2553 a_6285_122# a_6529_304# 0.00972f
C2554 VSS_SW_b[5] a_6231_220# 1.12e-20
C2555 a_5813_n88# a_7254_90# 5.39e-19
C2556 a_6017_n88# a_6730_n62# 8.07e-20
C2557 a_5504_106# a_5748_n62# 0.00707f
C2558 a_9595_627# VSS_SW_b[3] 1.08e-19
C2559 VDD_SW[4] a_10215_601# 7.64e-20
C2560 x9.A1 a_7252_1467# 0.197f
C2561 a_1501_122# VSS_SW_b[7] 7.15e-19
C2562 VDD a_10596_212# 0.687f
C2563 VDD_SW_b[2] a_13193_n88# 0.00132f
C2564 a_13461_1642# a_13193_n88# 4.63e-19
C2565 VDD a_8335_627# 6.2e-19
C2566 x2.X a_5812_212# 0.0129f
C2567 check[6] VDD_SW[7] 0.00393f
C2568 a_27_627# D[7] 0.138f
C2569 a_8933_1642# a_9147_1642# 0.00557f
C2570 x2.X a_12553_n62# 5.25e-20
C2571 VDD a_8921_304# 0.0042f
C2572 a_8432_993# a_8516_993# 0.00857f
C2573 a_7369_627# VDD_SW_b[4] 0.00231f
C2574 x9.A1 x14.X 9.22e-19
C2575 x11.X D[5] 0.1f
C2576 x2.X a_11240_909# 4.02e-19
C2577 x12.X a_7394_1315# 8.34e-19
C2578 x10.X a_5165_627# 6.12e-19
C2579 x2.X a_4149_1315# 2.33e-19
C2580 x2.X a_9595_627# 0.355f
C2581 a_10161_n62# a_10532_n62# 4.19e-20
C2582 x17.X VSS_SW_b[1] 0.0172f
C2583 a_10055_n62# a_12134_n88# 3.08e-21
C2584 a_27_627# a_2419_627# 1.63e-20
C2585 a_4811_627# a_5341_993# 4.45e-20
C2586 D[5] a_5165_627# 0.161f
C2587 a_10288_106# a_10597_n88# 0.0327f
C2588 a_10055_n62# a_10801_n88# 0.199f
C2589 VDD a_941_601# 0.461f
C2590 a_12988_212# a_15381_n88# 5.48e-21
C2591 a_12989_n88# a_15380_212# 8.02e-22
C2592 a_8205_n88# a_10055_n62# 4.56e-21
C2593 x2.X a_3732_993# 4.68e-19
C2594 a_3648_993# a_3947_627# 0.0256f
C2595 a_3333_601# VDD_SW[6] 1.79e-19
C2596 a_939_2457# x2.X 1.72f
C2597 a_3421_n88# a_3535_n62# 2.14e-20
C2598 a_3420_212# a_3761_n62# 0.00134f
C2599 a_3112_106# VSS_SW[5] 9.05e-21
C2600 a_14545_627# VDD_SW[1] 1.85e-20
C2601 a_15293_601# a_16488_627# 5.84e-19
C2602 x9.A1 a_5319_1642# 5.26e-19
C2603 a_10073_1289# a_10215_601# 8.76e-20
C2604 x2.X a_1233_n88# 0.00369f
C2605 check[3] a_7394_1642# 0.00688f
C2606 VDD a_2985_n62# 0.0133f
C2607 check[2] VSS_SW[3] 0.0493f
C2608 x9.A1 a_8591_895# 2.64e-19
C2609 D[7] VDD_SW[7] 0.246f
C2610 check[5] a_3625_n88# 2.51e-19
C2611 a_14379_627# a_14430_90# 6.13e-19
C2612 VDD a_1672_909# 0.00438f
C2613 VDD a_9949_627# 0.109f
C2614 a_487_n62# a_1447_220# 1.21e-20
C2615 a_1029_n88# a_678_220# 4.48e-20
C2616 a_1028_212# a_977_304# 2.13e-19
C2617 a_720_106# a_1166_304# 0.00412f
C2618 VDD_SW_b[2] a_14430_90# 0.00345f
C2619 D[2] a_14545_627# 7.7e-21
C2620 x11.X a_8117_601# 4.02e-21
C2621 x2.X a_15585_n88# 0.00368f
C2622 a_27_627# a_1112_909# 1.09e-19
C2623 D[7] a_891_909# 6.77e-19
C2624 a_12607_601# VDD_SW_b[2] 1.36e-20
C2625 a_12901_601# a_13119_627# 3.73e-19
C2626 a_12465_1289# a_12433_993# 4.54e-19
C2627 a_13216_993# a_12751_627# 0.00316f
C2628 a_8319_n62# a_8545_n62# 3.34e-19
C2629 a_4064_909# VDD_SW[6] 2.12e-20
C2630 VDD a_2927_1642# 8.63e-19
C2631 x8.X a_1415_895# 0.00864f
C2632 check[4] a_6199_895# 0.00267f
C2633 VDD a_5341_993# 0.0042f
C2634 D[6] a_3070_220# 2.03e-20
C2635 VSS_SW[2] a_12680_106# 4.62e-19
C2636 VDD x15.X 0.458f
C2637 x9.A1 VDD_SW_b[4] 2.35e-20
C2638 a_6199_895# a_8432_993# 1.86e-21
C2639 a_5725_601# a_7557_627# 2.42e-20
C2640 a_10596_212# a_11313_n62# 0.00206f
C2641 VDD_SW[7] a_2419_627# 0.0865f
C2642 a_14379_627# a_15608_993# 0.14f
C2643 D[1] a_15767_895# 0.0295f
C2644 a_14857_1289# a_14379_627# 0.00104f
C2645 D[3] a_12134_n88# 4.32e-19
C2646 a_5813_n88# a_8205_n88# 1.33e-19
C2647 a_5271_n62# VSS_SW_b[4] 8.69e-21
C2648 x10.X a_2585_627# 6.35e-20
C2649 a_10509_601# a_11069_122# 2.7e-19
C2650 a_1233_n88# a_1369_n62# 0.0697f
C2651 a_10983_895# a_10801_n88# 4.26e-19
C2652 VSS_SW_b[7] a_964_n62# 1.68e-19
C2653 a_1029_n88# VSS_SW[6] 9.23e-19
C2654 x15.X a_11325_1315# 1.98e-19
C2655 D[3] a_10801_n88# 0.00547f
C2656 a_4811_627# a_6017_n88# 0.00204f
C2657 a_13906_n62# a_15380_212# 5.58e-22
C2658 D[5] a_5813_n88# 0.159f
C2659 x2.X a_6529_304# 3.34e-19
C2660 x9.A1 a_14526_n88# 7.4e-19
C2661 a_193_627# a_381_627# 0.189f
C2662 a_647_601# a_1256_993# 0.00189f
C2663 x8.X VDD_SW_b[7] 7.23e-19
C2664 a_4860_1467# a_4862_90# 1e-19
C2665 a_3895_1642# x10.X 1.14e-20
C2666 check[1] a_12447_n62# 1.39e-20
C2667 a_8933_1642# check[3] 0.318f
C2668 x9.A1 VDD_SW[3] 0.0329f
C2669 D[6] a_4977_627# 6.42e-21
C2670 VDD_SW[3] a_12901_601# 2.46e-20
C2671 check[4] VDD_SW_b[5] 0.00213f
C2672 x8.X check[5] 0.00903f
C2673 D[6] VSS_SW[5] 4.85e-19
C2674 a_15464_909# VDD_SW_b[1] 9.36e-21
C2675 a_15143_627# a_15511_627# 3.34e-19
C2676 x9.A1 a_2136_627# 2e-20
C2677 x2.X VSS_SW[2] 0.0861f
C2678 x15.X a_10596_212# 0.245f
C2679 VDD a_2468_1467# 0.114f
C2680 x2.X a_10041_993# 0.15f
C2681 x9.A1 a_1256_993# 4.84e-21
C2682 a_5002_1642# VSS_SW[5] 0.00105f
C2683 D[4] VSS_SW[4] 0.133f
C2684 x12.X a_6539_1315# 2.36e-20
C2685 a_76_1467# a_218_1315# 0.00783f
C2686 x14.X a_9595_627# 0.236f
C2687 check[2] VDD_SW[4] 4.35e-19
C2688 x2.X x9.X 0.00459f
C2689 a_4413_2457# x9.X 4.53e-20
C2690 a_15293_601# a_15381_n88# 3.89e-19
C2691 a_15767_895# a_15380_212# 0.00165f
C2692 a_14857_1289# a_15072_106# 5.3e-21
C2693 a_14545_627# VSS_SW_b[1] 5.23e-20
C2694 a_1112_909# VDD_SW[7] 2.82e-20
C2695 a_1757_1642# check[6] 0.318f
C2696 a_305_2457# a_27_627# 1.18e-19
C2697 D[5] a_6920_627# 0.00234f
C2698 x18.X a_14430_90# 0.00259f
C2699 a_941_601# a_1672_909# 0.0016f
C2700 a_473_993# VDD_SW_b[7] 3.93e-21
C2701 x2.X a_14945_n62# 5.25e-20
C2702 x18.X a_12607_601# 1.98e-20
C2703 x12.X a_7823_601# 2.7e-20
C2704 a_9312_627# VSS_SW[3] 0.00166f
C2705 VDD_SW_b[4] a_9742_n88# 5.91e-19
C2706 check[3] a_7350_n88# 5.26e-19
C2707 a_9646_90# a_9742_n88# 0.0967f
C2708 a_3421_n88# VSS_SW_b[5] 0.00486f
C2709 a_3839_220# VSS_SW[5] 1.57e-20
C2710 x30.A a_5323_2457# 0.619f
C2711 a_1503_1642# a_1415_895# 5.45e-19
C2712 a_4689_2457# x2.X 0.00106f
C2713 a_4413_2457# a_4689_2457# 0.00202f
C2714 a_13193_n88# a_13461_122# 0.206f
C2715 a_12989_n88# VSS_SW_b[2] 7.6e-19
C2716 check[6] a_487_n62# 1.41e-20
C2717 VSS_SW[2] a_13407_220# 6.42e-21
C2718 a_16109_1642# x20.X 0.0846f
C2719 a_2585_627# VSS_SW_b[6] 5.23e-20
C2720 a_11987_627# a_12038_90# 6.13e-19
C2721 a_3807_895# a_3420_212# 0.00165f
C2722 a_3333_601# a_3421_n88# 3.89e-19
C2723 a_16109_1642# VDD_SW_b[1] 2.6e-19
C2724 x2.X a_593_n62# 5.57e-20
C2725 check[4] a_5504_106# 7.9e-22
C2726 a_10459_909# VDD_SW_b[3] 3.01e-21
C2727 VDD a_6017_n88# 0.48f
C2728 VDD_SW_b[3] a_12038_90# 0.00346f
C2729 x18.X a_14857_1289# 1.51e-19
C2730 a_4370_1315# D[6] 0.0012f
C2731 a_2610_1315# VSS_SW[6] 7.95e-19
C2732 a_9595_627# a_10680_909# 1.09e-19
C2733 a_6285_1642# x11.X 1.3e-19
C2734 VDD a_3039_601# 0.313f
C2735 a_720_106# a_2566_n88# 1.86e-21
C2736 a_4977_627# a_5725_601# 0.126f
C2737 VDD a_11015_220# 0.00984f
C2738 a_5431_601# a_5257_993# 0.206f
C2739 a_5725_601# VSS_SW[5] 2.18e-19
C2740 a_8591_895# a_9595_627# 6.9e-19
C2741 a_8117_601# D[3] 8.74e-19
C2742 a_647_601# VSS_SW[7] 6.23e-19
C2743 x9.A1 a_11071_1642# 0.101f
C2744 a_11987_627# a_12541_627# 0.00206f
C2745 x20.X VDD_SW[1] 0.177f
C2746 check[2] a_10073_1289# 0.248f
C2747 a_16330_1315# VDD_SW_b[1] 1.33e-20
C2748 VDD_SW_b[1] VDD_SW[1] 3.65e-19
C2749 x20.X a_16330_1315# 0.00143f
C2750 VDD a_6339_627# 6.99e-19
C2751 VDD_SW_b[6] a_3420_212# 0.0418f
C2752 a_1503_1642# check[5] 1.16e-20
C2753 a_6920_627# a_8117_601# 1.71e-20
C2754 VDD_SW[5] a_7369_627# 9.25e-19
C2755 x3.A x3.X 4.66e-19
C2756 reset ready 0.0713f
C2757 a_1757_1642# D[7] 0.0607f
C2758 VDD a_13072_909# 0.0164f
C2759 a_5950_304# VSS_SW_b[4] 9.89e-21
C2760 a_14825_993# a_14945_n62# 6.88e-22
C2761 a_7254_90# a_8204_212# 1.66e-20
C2762 a_6730_n62# a_8205_n88# 3.67e-21
C2763 x9.A1 VSS_SW[7] 0.108f
C2764 a_2470_90# VSS_SW[6] 0.082f
C2765 a_1501_122# VSS_SW_b[6] 1.09e-20
C2766 a_14379_627# D[1] 0.138f
C2767 a_5431_601# a_5943_627# 9.75e-19
C2768 a_5725_601# a_5575_627# 0.00926f
C2769 a_4977_627# a_6456_909# 7.17e-20
C2770 a_6040_993# a_5896_909# 0.00412f
C2771 a_5257_993# a_5365_627# 0.00807f
C2772 VDD_SW_b[2] D[1] 1.5e-19
C2773 a_10055_n62# a_11514_n62# 3.79e-20
C2774 a_10597_n88# a_10734_304# 0.00907f
C2775 a_10596_212# a_11015_220# 2.46e-19
C2776 D[5] a_6730_n62# 0.158f
C2777 x2.X a_7896_106# 0.0385f
C2778 x8.X a_2865_993# 9.17e-20
C2779 a_2897_1289# a_3112_106# 5.3e-21
C2780 VDD_SW_b[4] a_9595_627# 5.97e-19
C2781 a_8731_627# a_8539_627# 4.19e-20
C2782 a_9312_627# VDD_SW[4] 0.0729f
C2783 a_581_627# VSS_SW[7] 3.79e-19
C2784 VDD VSS_SW_b[7] 0.106f
C2785 a_9595_627# a_9646_90# 6.13e-19
C2786 a_7681_1289# a_7203_627# 0.00104f
C2787 D[7] a_487_n62# 0.00257f
C2788 a_27_627# a_720_106# 3.88e-21
C2789 VDD a_15511_627# 6.2e-19
C2790 x9.A1 a_12989_n88# 8.59e-21
C2791 a_12901_601# a_12989_n88# 3.89e-19
C2792 a_12153_627# VSS_SW_b[2] 5.25e-20
C2793 a_13375_895# a_12988_212# 0.00165f
C2794 a_505_1289# VSS_SW[7] 0.00189f
C2795 a_11240_909# VDD_SW[3] 2.12e-20
C2796 a_5289_1289# a_5431_601# 8.76e-20
C2797 a_2419_627# a_2773_627# 0.0455f
C2798 D[6] a_3648_993# 0.00608f
C2799 a_2468_1467# a_2927_1642# 6.64e-19
C2800 x14.X a_10041_993# 9.14e-20
C2801 a_9595_627# VDD_SW[3] 3.29e-20
C2802 x11.X x12.X 0.11f
C2803 a_1415_895# a_2585_627# 2.96e-19
C2804 a_941_601# a_3039_601# 1.52e-20
C2805 D[1] a_15072_106# 8.75e-19
C2806 a_14379_627# a_15380_212# 6.99e-20
C2807 VDD_SW_b[2] a_15380_212# 4.59e-22
C2808 VDD_SW[2] VSS_SW[1] 0.429f
C2809 x13.X a_8205_n88# 0.019f
C2810 a_7252_1467# a_7394_1315# 0.00783f
C2811 a_4977_627# a_5271_n62# 2.38e-19
C2812 x9.A1 VSS_SW_b[5] 2.85e-19
C2813 x9.A1 x16.X 9.19e-19
C2814 a_5431_601# a_4958_n88# 4.37e-19
C2815 a_4338_n62# VSS_SW_b[5] 2.64e-19
C2816 VSS_SW[5] a_5271_n62# 3.44e-19
C2817 x16.X a_12901_601# 4.99e-20
C2818 x2.X a_13216_993# 0.187f
C2819 D[4] a_10597_n88# 4.83e-22
C2820 x9.A1 a_3333_601# 0.00103f
C2821 x2.X a_6539_1315# 2.34e-19
C2822 x11.X a_6285_122# 2.61e-19
C2823 x2.X a_3625_n88# 0.00371f
C2824 a_3039_601# a_2985_n62# 1.07e-20
C2825 VDD a_7254_90# 0.189f
C2826 VDD VDD_SW[2] 0.373f
C2827 VDD_SW[7] a_2949_993# 6.61e-21
C2828 a_939_2457# a_2136_627# 6.01e-19
C2829 VDD_SW_b[7] a_2585_627# 0.00329f
C2830 x18.X D[1] 0.00892f
C2831 ready a_1415_895# 3.23e-21
C2832 a_939_2457# a_1256_993# 4.83e-21
C2833 a_10983_895# a_11514_n62# 4.06e-19
C2834 a_10509_601# a_10459_909# 1.21e-20
C2835 D[3] a_10125_993# 8.11e-19
C2836 x9.A1 VDD_SW[5] 0.0926f
C2837 x2.X a_7823_601# 0.2f
C2838 D[3] a_11514_n62# 0.158f
C2839 x2.X a_15464_909# 0.00309f
C2840 a_15072_106# a_15380_212# 0.14f
C2841 a_14839_n62# a_15381_n88# 0.125f
C2842 check[5] a_2585_627# 5.42e-19
C2843 a_10509_601# VSS_SW[3] 2.13e-19
C2844 a_2897_1289# D[6] 0.0661f
C2845 a_1256_993# a_1233_n88# 1.86e-19
C2846 a_1415_895# a_1501_122# 4.53e-22
C2847 a_8623_220# VSS_SW_b[3] 3.75e-21
C2848 a_8591_895# a_10041_993# 8e-21
C2849 x9.A1 a_13906_n62# 1.56e-20
C2850 x9.A1 a_12153_627# 3.23e-19
C2851 a_12607_601# a_12433_993# 0.206f
C2852 a_12153_627# a_12901_601# 0.126f
C2853 x7.X a_1978_1315# 0.00146f
C2854 check[1] a_12038_90# 2.5e-20
C2855 x9.A1 a_7711_1642# 5.26e-19
C2856 check[5] a_3895_1642# 0.257f
C2857 D[4] a_8067_909# 6.77e-19
C2858 a_7203_627# a_8288_909# 1.09e-19
C2859 a_7896_106# a_8409_n88# 0.00189f
C2860 a_7663_n62# a_8677_122# 0.0633f
C2861 a_7350_n88# VSS_SW_b[4] 0.135f
C2862 a_8204_212# a_8205_n88# 0.784f
C2863 check[4] VDD_SW[6] 4.33e-19
C2864 x10.X a_4811_627# 0.236f
C2865 ready VDD_SW_b[7] 1.14e-20
C2866 VSS_SW[6] a_3421_n88# 9.29e-21
C2867 x2.X a_7757_627# 3.94e-19
C2868 a_6040_993# VDD_SW[5] 3.28e-20
C2869 D[1] a_15799_220# 7.1e-19
C2870 D[5] a_8204_212# 7.45e-22
C2871 x2.X a_8623_220# 9.51e-19
C2872 x2.X x8.X 5.54e-19
C2873 x9.A1 a_15767_895# 2.64e-19
C2874 x17.X VSS_SW[1] 0.148f
C2875 x13.X a_8117_601# 1.31e-19
C2876 VDD_SW_b[7] a_1501_122# 0.00445f
C2877 ready check[5] 0.0417f
C2878 VDD a_1143_n62# 0.00535f
C2879 a_13375_895# a_15293_601# 1.42e-20
C2880 VDD_SW_b[4] a_10041_993# 8.2e-21
C2881 x2.X a_16109_1642# 5.24e-19
C2882 D[7] a_1447_220# 7.11e-19
C2883 a_4811_627# D[5] 0.137f
C2884 a_7369_627# a_9761_627# 2.62e-19
C2885 x27.A VSS_SW[5] 6.7e-19
C2886 a_12447_n62# a_13329_n62# 0.00926f
C2887 a_12680_106# a_13103_n62# 0.00386f
C2888 a_12134_n88# VSS_SW[1] 4.28e-21
C2889 a_7203_627# VSS_SW[3] 4.95e-21
C2890 a_2419_627# a_4528_627# 1.75e-19
C2891 VDD x17.X 0.458f
C2892 a_11987_627# a_12988_212# 6.99e-20
C2893 D[2] a_12680_106# 8.76e-19
C2894 VDD_SW_b[1] a_15495_n62# 5.19e-19
C2895 VDD_SW[3] VSS_SW[2] 0.427f
C2896 VDD_SW_b[3] a_12988_212# 4.59e-22
C2897 a_14857_1289# a_15855_1642# 0.0146f
C2898 a_15293_601# a_15243_909# 1.21e-20
C2899 a_15855_1642# a_15608_993# 0.00176f
C2900 a_14545_627# a_15143_627# 6.04e-20
C2901 a_10983_895# a_11123_627# 0.0383f
C2902 a_10509_601# a_10931_627# 1.96e-20
C2903 a_10041_993# VDD_SW[3] 4.17e-21
C2904 x2.X a_473_993# 0.15f
C2905 D[3] a_11123_627# 0.00433f
C2906 x2.X VDD_SW[1] 0.0322f
C2907 a_15381_n88# a_15518_304# 0.00907f
C2908 a_14839_n62# a_16298_n62# 3.79e-20
C2909 a_15380_212# a_15799_220# 2.46e-19
C2910 a_939_2457# VSS_SW[7] 0.00403f
C2911 a_14526_n88# a_14945_n62# 0.0383f
C2912 x13.X a_9122_n62# 0.0016f
C2913 VDD a_12134_n88# 0.69f
C2914 VDD_SW[4] a_10509_601# 2.55e-20
C2915 x9.A1 a_9644_1467# 0.197f
C2916 VSS_SW[5] a_5950_304# 1.97e-20
C2917 a_5813_n88# a_6285_122# 0.15f
C2918 a_5812_212# VSS_SW_b[5] 0.00119f
C2919 VDD a_10801_n88# 0.48f
C2920 a_8933_1642# check[2] 1.62e-19
C2921 VDD x10.X 0.338f
C2922 VSS_SW[7] a_1233_n88# 9.92e-21
C2923 x30.A a_5725_601# 2.1e-19
C2924 x12.X a_6920_627# 0.0285f
C2925 a_6539_1642# a_6760_1315# 0.00783f
C2926 x2.X a_4862_90# 0.00369f
C2927 x2.X D[2] 0.199f
C2928 VDD a_8205_n88# 0.66f
C2929 x6.X a_218_1315# 8.34e-19
C2930 x16.X a_9595_627# 0.00117f
C2931 a_8432_993# a_7663_n62# 3.59e-19
C2932 a_7557_627# a_7350_n88# 3.32e-19
C2933 a_8117_601# a_8204_212# 6.03e-19
C2934 x2.X x11.X 0.00457f
C2935 a_2585_627# a_2865_993# 0.15f
C2936 x2.X a_1159_627# 0.00702f
C2937 VDD D[5] 0.797f
C2938 a_2566_n88# a_3112_106# 0.207f
C2939 a_5725_601# a_7203_627# 3.81e-19
C2940 a_10596_212# a_12134_n88# 6.15e-19
C2941 a_10215_601# a_10161_n62# 1.07e-20
C2942 a_6339_627# a_6017_n88# 7.32e-20
C2943 VDD_SW[5] a_5812_212# 4.35e-19
C2944 x14.X a_7823_601# 1.98e-20
C2945 x2.X a_1503_1642# 0.00652f
C2946 a_10055_n62# VSS_SW_b[3] 0.0142f
C2947 VSS_SW[3] a_10246_220# 4.25e-19
C2948 a_10596_212# a_10801_n88# 0.15f
C2949 x2.X a_5165_627# 0.0014f
C2950 a_4149_1642# a_4528_627# 5.9e-19
C2951 D[4] a_8539_627# 2e-19
C2952 a_7203_627# VDD_SW[4] 3.29e-20
C2953 a_8205_n88# a_10596_212# 4.01e-22
C2954 D[2] a_13407_220# 7.11e-19
C2955 VDD_SW_b[4] a_7896_106# 5.23e-19
C2956 a_2773_627# a_2949_993# 8.99e-19
C2957 check[6] D[7] 0.463f
C2958 a_2585_627# a_3551_627# 2.14e-20
C2959 a_3333_601# a_3732_993# 9.41e-19
C2960 a_8409_n88# a_8623_220# 0.0104f
C2961 a_2865_993# a_3183_627# 0.025f
C2962 a_7663_n62# a_7769_n62# 0.0526f
C2963 x9.A1 VSS_SW[6] 0.113f
C2964 a_8205_n88# a_8921_304# 0.0018f
C2965 a_8204_212# a_9122_n62# 0.0453f
C2966 a_9644_1467# a_9742_n88# 6.87e-20
C2967 a_15767_895# a_15907_627# 0.0383f
C2968 ready a_2865_993# 5.7e-21
C2969 a_15293_601# a_15715_627# 1.96e-20
C2970 a_14825_993# VDD_SW[1] 4.17e-21
C2971 a_3893_122# VSS_SW_b[6] 7.15e-19
C2972 x9.A1 a_9761_627# 3.23e-19
C2973 check[3] a_8861_1642# 0.00577f
C2974 a_9595_627# a_12153_627# 1.09e-20
C2975 x2.X a_10055_n62# 0.373f
C2976 VDD_SW_b[5] a_5927_n62# 5.21e-19
C2977 VDD a_12937_304# 0.00266f
C2978 a_11325_1642# a_12036_1467# 0.00963f
C2979 VDD_SW_b[7] a_964_n62# 8.1e-20
C2980 VDD VSS_SW_b[6] 0.0968f
C2981 a_14545_627# VSS_SW[1] 0.023f
C2982 VDD reset 0.16f
C2983 D[7] a_2879_n62# 3.12e-21
C2984 x9.A1 a_14379_627# 8.16e-19
C2985 a_4860_1467# a_4811_627# 5.32e-19
C2986 a_12901_601# a_14379_627# 3.77e-19
C2987 x2.X VSS_SW_b[1] 0.0278f
C2988 x9.A1 a_13461_1642# 0.101f
C2989 x9.A1 VDD_SW_b[2] 2.34e-20
C2990 a_4958_n88# a_5462_220# 0.00869f
C2991 a_13461_1642# a_12901_601# 0.00263f
C2992 a_12901_601# VDD_SW_b[2] 0.00647f
C2993 a_12341_627# a_12541_627# 3.81e-19
C2994 a_13216_993# a_13119_627# 0.00386f
C2995 a_13375_895# a_13632_909# 0.00869f
C2996 a_174_n88# a_1028_212# 0.0319f
C2997 a_487_n62# a_720_106# 0.124f
C2998 check[2] a_12465_1289# 4.15e-21
C2999 a_5323_2457# a_5431_601# 4.92e-19
C3000 VDD a_4363_1642# 0.00177f
C3001 a_3504_909# VDD_SW_b[6] 7.04e-21
C3002 VDD a_8117_601# 0.46f
C3003 a_3183_627# a_3551_627# 3.34e-19
C3004 a_7649_993# a_8117_601# 0.0633f
C3005 a_7369_627# a_8432_993# 0.0334f
C3006 VDD a_14545_627# 0.659f
C3007 a_8933_1642# a_9312_627# 5.9e-19
C3008 VSS_SW[2] a_12989_n88# 9.3e-21
C3009 check[6] a_535_1642# 0.00526f
C3010 D[6] a_2566_n88# 0.00507f
C3011 check[0] a_14999_601# 0.00262f
C3012 a_2419_627# a_2879_n62# 7.27e-19
C3013 a_15855_1642# D[1] 0.0681f
C3014 a_14379_627# a_14909_993# 4.45e-20
C3015 D[1] a_14733_627# 0.161f
C3016 D[3] a_12680_106# 2.77e-21
C3017 x9.A1 a_8677_122# 4.36e-20
C3018 a_10824_993# a_11069_122# 1.51e-20
C3019 a_10359_627# a_9742_n88# 1.08e-19
C3020 a_4958_n88# VSS_SW[4] 4.28e-21
C3021 a_5271_n62# a_6153_n62# 0.00926f
C3022 a_6285_122# a_6730_n62# 0.0369f
C3023 a_5504_106# a_5927_n62# 0.00386f
C3024 D[3] VSS_SW_b[3] 5.32e-19
C3025 a_9761_627# a_9742_n88# 4.91e-19
C3026 a_13407_220# VSS_SW_b[1] 3.96e-21
C3027 a_14430_90# a_15381_n88# 9.87e-21
C3028 VDD a_8848_909# 0.00438f
C3029 x2.X a_5813_n88# 0.0213f
C3030 VDD a_9122_n62# 0.109f
C3031 check[1] a_12988_212# 3.22e-20
C3032 a_8432_993# a_7967_627# 0.00316f
C3033 a_7823_601# VDD_SW_b[4] 2.14e-20
C3034 a_8117_601# a_8335_627# 3.73e-19
C3035 x16.X VSS_SW[2] 0.249f
C3036 a_7252_1467# x11.X 4.9e-19
C3037 VDD_SW[3] a_13216_993# 1.08e-20
C3038 x15.X a_12134_n88# 0.00865f
C3039 a_9644_1467# a_9595_627# 5.32e-19
C3040 x16.X a_10041_993# 1.56e-20
C3041 x2.X a_2585_627# 0.0537f
C3042 x15.X a_10801_n88# 1.87e-19
C3043 x9.X VSS_SW_b[5] 0.0173f
C3044 a_3112_106# a_3369_304# 0.00857f
C3045 x2.X a_10983_895# 0.148f
C3046 a_2879_n62# a_3558_304# 0.00652f
C3047 VDD a_4860_1467# 0.114f
C3048 x2.X D[3] 0.199f
C3049 a_15767_895# a_15585_n88# 4.26e-19
C3050 a_15855_1642# a_15380_212# 1.39e-21
C3051 a_15293_601# a_15853_122# 2.7e-19
C3052 x9.X a_3333_601# 1.27e-19
C3053 x2.X a_3895_1642# 0.00651f
C3054 a_13715_1642# VDD_SW_b[2] 2.58e-19
C3055 a_12036_1467# a_12178_1642# 0.00557f
C3056 x9.A1 x18.X 9.23e-19
C3057 a_27_627# D[6] 1.19e-20
C3058 D[7] a_2419_627# 9.98e-20
C3059 a_4811_627# a_5675_909# 2.46e-19
C3060 x18.X a_12901_601# 0.00129f
C3061 D[5] a_5341_993# 8.11e-19
C3062 x2.X a_6920_627# 3.85e-19
C3063 a_13072_909# VDD_SW[2] 2.82e-20
C3064 x14.X a_9786_1315# 8.2e-19
C3065 VDD a_1415_895# 0.671f
C3066 a_9122_n62# a_10596_212# 2.79e-22
C3067 x2.X a_8933_1315# 2.32e-19
C3068 a_3648_993# a_3755_627# 0.00707f
C3069 a_8921_304# a_9122_n62# 8.99e-19
C3070 x2.X a_3183_627# 0.0388f
C3071 a_8677_122# a_9742_n88# 8e-21
C3072 a_3807_895# VDD_SW[6] 0.00356f
C3073 a_535_1642# D[7] 5.72e-19
C3074 ready x2.X 0.437f
C3075 x27.A x30.A 4.66e-19
C3076 VSS_SW_b[6] a_2985_n62# 0.00335f
C3077 a_13461_122# VSS_SW_b[2] 7.16e-19
C3078 a_3420_212# VSS_SW[5] 0.0872f
C3079 a_3625_n88# a_3535_n62# 9.75e-19
C3080 a_3421_n88# a_3761_n62# 6.04e-20
C3081 ready a_4413_2457# 0.202f
C3082 a_12153_627# VSS_SW[2] 0.0232f
C3083 a_14570_1315# D[1] 7.54e-19
C3084 VDD_SW_b[5] VSS_SW_b[4] 0.0383f
C3085 D[1] a_16488_627# 0.00233f
C3086 x9.A1 check[4] 0.473f
C3087 x2.X a_1501_122# 0.0043f
C3088 a_9761_627# a_11240_909# 7.17e-20
C3089 VDD a_3356_n62# 7.87e-19
C3090 x9.A1 a_8432_993# 4.84e-21
C3091 a_9595_627# a_10359_627# 0.00134f
C3092 a_9595_627# a_9761_627# 0.786f
C3093 VDD a_11514_n62# 0.109f
C3094 check[5] a_3893_122# 6.44e-20
C3095 VDD a_10125_993# 0.0042f
C3096 VDD VDD_SW_b[7] 0.156f
C3097 a_1028_212# a_1166_304# 1.09e-19
C3098 a_8117_601# a_9949_627# 2.42e-20
C3099 a_27_627# a_1340_993# 2.13e-19
C3100 D[7] a_1112_909# 8.51e-19
C3101 VDD_SW_b[2] a_12553_n62# 4.77e-19
C3102 x8.X a_2136_627# 0.0285f
C3103 a_305_2457# check[6] 0.00376f
C3104 VDD a_6285_1642# 0.191f
C3105 a_12465_1289# a_11987_627# 0.00104f
C3106 VDD_SW_b[6] VDD_SW[6] 3.64e-19
C3107 D[2] a_13119_627# 6.12e-19
C3108 x9.A1 a_10103_1642# 5.26e-19
C3109 x8.X a_1256_993# 2.81e-19
C3110 check[2] a_9786_1642# 0.00688f
C3111 VDD check[5] 1.65f
C3112 x12.X a_4811_627# 0.00117f
C3113 check[4] a_6040_993# 2.89e-19
C3114 VDD a_5675_909# 0.00984f
C3115 a_939_2457# VSS_SW[6] 0.0213f
C3116 a_6199_895# a_7557_627# 8.26e-21
C3117 VDD a_12751_627# 1.8e-19
C3118 a_16488_627# a_15380_212# 6.63e-19
C3119 VDD_SW[7] D[6] 4.48e-19
C3120 a_13715_1642# x18.X 7.95e-19
C3121 x10.X a_3039_601# 1.98e-20
C3122 a_10801_n88# a_11015_220# 0.0104f
C3123 a_10597_n88# a_11313_304# 0.0018f
C3124 a_1501_122# a_1369_n62# 0.025f
C3125 VSS_SW_b[7] a_1143_n62# 5.24e-19
C3126 a_10596_212# a_11514_n62# 0.0453f
C3127 a_1233_n88# VSS_SW[6] 8.81e-20
C3128 x2.X a_6730_n62# 1.83e-19
C3129 D[5] a_6017_n88# 0.00547f
C3130 a_647_601# a_381_627# 8.07e-20
C3131 a_193_627# a_557_993# 0.0018f
C3132 a_941_601# a_1415_895# 0.265f
C3133 VSS_SW[3] a_10288_106# 4.65e-19
C3134 D[2] a_14526_n88# 4.33e-19
C3135 VDD a_78_90# 0.195f
C3136 a_2468_1467# VSS_SW_b[6] 2.13e-19
C3137 VDD VDD_SW_b[1] 0.156f
C3138 VDD x20.X 0.437f
C3139 x9.A1 a_13461_122# 5.09e-20
C3140 x9.A1 a_1745_n62# 5.7e-21
C3141 a_13375_895# a_13193_n88# 4.26e-19
C3142 a_12901_601# a_13461_122# 2.7e-19
C3143 VDD_SW[3] D[2] 4.58e-19
C3144 a_29_2457# x9.A1 9.28e-20
C3145 a_2879_n62# a_4958_n88# 5.13e-21
C3146 x9.A1 a_1555_627# 5.22e-20
C3147 VDD_SW_b[5] a_7557_627# 9.3e-21
C3148 x18.X a_14791_1315# 2.35e-19
C3149 x2.X a_10545_304# 0.00167f
C3150 x17.X a_13715_1315# 2.08e-19
C3151 x9.A1 a_381_627# 4.11e-19
C3152 a_4149_1642# a_4077_1642# 6.64e-19
C3153 x14.X D[3] 0.00895f
C3154 x13.X VSS_SW_b[3] 0.0171f
C3155 a_791_627# a_1363_627# 2.46e-21
C3156 VDD a_11123_627# 6.99e-19
C3157 D[5] a_6339_627# 0.00433f
C3158 a_305_2457# D[7] 1.02e-19
C3159 D[1] a_15381_n88# 0.158f
C3160 a_14379_627# a_15585_n88# 0.00204f
C3161 x3.X a_27_627# 5.4e-19
C3162 a_941_601# VDD_SW_b[7] 0.00647f
C3163 a_1256_993# a_1159_627# 0.00386f
C3164 a_381_627# a_581_627# 3.81e-19
C3165 a_1415_895# a_1672_909# 0.00869f
C3166 VDD x12.X 0.338f
C3167 a_11325_1642# a_11539_1642# 0.00557f
C3168 x12.X a_7649_993# 1.03e-19
C3169 check[3] a_7663_n62# 1.36e-20
C3170 a_9646_90# a_10055_n62# 4.24e-20
C3171 x2.X a_12517_993# 5.32e-19
C3172 x14.X a_8933_1315# 1.48e-20
C3173 a_4137_304# VSS_SW[5] 6.58e-21
C3174 a_2985_n62# a_3356_n62# 4.19e-20
C3175 a_3625_n88# VSS_SW_b[5] 4.55e-20
C3176 a_1503_1642# a_1256_993# 0.00176f
C3177 x7.X a_174_n88# 1.64e-21
C3178 x2.X x13.X 0.00458f
C3179 check[6] a_720_106# 8.67e-22
C3180 x2.X a_964_n62# 3.68e-20
C3181 a_3648_993# a_3420_212# 8.94e-21
C3182 a_3807_895# a_3421_n88# 6.35e-19
C3183 a_3333_601# a_3625_n88# 0.00251f
C3184 check[4] a_5812_212# 3.11e-20
C3185 a_11514_n62# a_11313_n62# 3.81e-19
C3186 VDD a_6285_122# 0.313f
C3187 VDD_SW_b[3] a_10161_n62# 4.78e-19
C3188 a_10509_601# a_10908_993# 9.41e-19
C3189 a_9949_627# a_10125_993# 8.99e-19
C3190 a_10041_993# a_10359_627# 0.025f
C3191 a_9761_627# VSS_SW[2] 5.1e-21
C3192 a_11123_627# a_10596_212# 7.07e-21
C3193 x17.X VDD_SW[2] 0.177f
C3194 a_1672_909# VDD_SW_b[7] 3.14e-20
C3195 D[3] a_10680_909# 8.53e-19
C3196 x2.X a_15143_627# 0.0388f
C3197 VDD a_2865_993# 0.18f
C3198 a_1028_212# a_2566_n88# 6.15e-19
C3199 a_9761_627# a_10041_993# 0.15f
C3200 a_15072_106# a_15585_n88# 0.00189f
C3201 a_14839_n62# a_15853_122# 0.0633f
C3202 a_14526_n88# VSS_SW_b[1] 0.135f
C3203 a_15380_212# a_15381_n88# 0.785f
C3204 a_5323_2457# VSS_SW[4] 2.07e-19
C3205 a_4977_627# a_6199_895# 0.0494f
C3206 a_5431_601# a_5725_601# 0.199f
C3207 a_12036_1467# VSS_SW_b[2] 2.11e-19
C3208 a_8432_993# a_9595_627# 7.56e-20
C3209 a_473_993# VSS_SW[7] 0.00296f
C3210 a_8591_895# D[3] 2.1e-19
C3211 a_14096_627# a_12988_212# 6.63e-19
C3212 x9.A1 a_12433_993# 1.42e-19
C3213 a_12433_993# a_12901_601# 0.0633f
C3214 a_8204_212# VSS_SW_b[3] 0.00374f
C3215 a_12153_627# a_13216_993# 0.0334f
C3216 check[5] a_2927_1642# 0.00526f
C3217 x15.X a_11514_n62# 0.00162f
C3218 VDD_SW_b[6] a_3421_n88# 0.0406f
C3219 VDD_SW[5] a_7823_601# 7.64e-20
C3220 a_8679_1642# x13.X 1.35e-19
C3221 a_7203_627# a_7350_n88# 0.00176f
C3222 a_6231_220# VSS_SW_b[4] 3.96e-21
C3223 a_7254_90# a_8205_n88# 9.87e-21
C3224 a_5812_212# a_7769_n62# 1.09e-19
C3225 VDD a_3551_627# 6.2e-19
C3226 D[1] a_16298_n62# 0.158f
C3227 a_964_n62# a_1369_n62# 2.46e-21
C3228 a_6040_993# a_6124_993# 0.00857f
C3229 a_4977_627# VDD_SW_b[5] 0.00226f
C3230 x9.A1 a_15855_1642# 0.101f
C3231 x9.A1 a_14733_627# 4.11e-19
C3232 a_12901_601# a_14733_627# 2.27e-20
C3233 a_13375_895# a_15608_993# 1.86e-21
C3234 D[5] a_7254_90# 8.71e-19
C3235 x2.X a_8204_212# 0.0128f
C3236 check[1] a_12465_1289# 0.248f
C3237 x8.X a_3333_601# 4.9e-20
C3238 VDD_SW_b[4] D[3] 1.51e-19
C3239 check[3] a_7369_627# 5.38e-19
C3240 a_7681_1289# D[4] 0.0662f
C3241 x2.X a_13515_627# 0.0151f
C3242 a_27_627# a_1028_212# 6.99e-20
C3243 D[7] a_720_106# 8.74e-19
C3244 a_7681_1289# VSS_SW[4] 0.0019f
C3245 x2.X a_4811_627# 0.354f
C3246 a_12680_106# VSS_SW[1] 9.06e-21
C3247 a_12988_212# a_13329_n62# 0.00134f
C3248 a_3420_212# a_4137_n62# 0.00206f
C3249 a_12989_n88# a_13103_n62# 2.14e-20
C3250 a_1757_1642# D[6] 1.69e-19
C3251 a_11987_627# a_13193_n88# 0.00204f
C3252 D[2] a_12989_n88# 0.158f
C3253 VDD_SW_b[1] a_16097_n62# 5.21e-19
C3254 a_5289_1289# a_5257_993# 4.54e-19
C3255 a_2419_627# a_2949_993# 4.45e-20
C3256 D[6] a_2773_627# 0.161f
C3257 a_15293_601# a_15692_993# 9.41e-19
C3258 a_14545_627# a_15511_627# 2.14e-20
C3259 a_14825_993# a_15143_627# 0.025f
C3260 a_14733_627# a_14909_993# 8.99e-19
C3261 a_10824_993# a_10931_627# 0.00707f
C3262 a_10983_895# VDD_SW[3] 0.00356f
C3263 a_2136_627# a_2585_627# 5.39e-19
C3264 D[3] VDD_SW[3] 0.245f
C3265 a_10073_1289# a_10288_106# 5.3e-21
C3266 a_2468_1467# check[5] 0.318f
C3267 a_1757_1642# a_1685_1642# 6.64e-19
C3268 a_1256_993# a_2585_627# 4.03e-21
C3269 a_941_601# a_2865_993# 1.11e-20
C3270 a_15380_212# a_16298_n62# 0.0453f
C3271 a_15381_n88# a_16097_304# 0.0018f
C3272 a_15072_106# a_14945_n62# 0.0256f
C3273 a_14839_n62# a_15316_n62# 1.96e-20
C3274 a_15585_n88# a_15799_220# 0.0104f
C3275 VDD a_12680_106# 0.356f
C3276 VDD_SW[4] a_10824_993# 1.08e-20
C3277 a_14428_1467# a_14430_90# 1e-19
C3278 x13.X a_8409_n88# 1.81e-19
C3279 x9.A1 a_12036_1467# 0.197f
C3280 a_5431_601# a_5271_n62# 0.0026f
C3281 VDD VSS_SW_b[3] 0.0967f
C3282 a_5257_993# a_4958_n88# 8.71e-20
C3283 a_11325_1642# check[2] 0.318f
C3284 a_8679_1642# a_8204_212# 1.39e-21
C3285 VSS_SW[5] a_5504_106# 4.64e-19
C3286 a_4862_90# VSS_SW_b[5] 0.191f
C3287 x17.X a_12134_n88# 1.64e-21
C3288 a_193_627# a_174_n88# 4.91e-19
C3289 x2.X VSS_SW[1] 0.086f
C3290 x16.X D[2] 0.00861f
C3291 x9.A1 a_3807_895# 2.64e-19
C3292 a_2865_993# a_2985_n62# 6.88e-22
C3293 x2.X a_3893_122# 0.0043f
C3294 a_3807_895# a_4338_n62# 4.06e-19
C3295 x13.X x14.X 0.11f
C3296 VDD a_5377_n62# 0.0133f
C3297 a_6285_1642# a_6017_n88# 4.63e-19
C3298 VDD_SW[7] a_3283_909# 2.16e-20
C3299 a_29_2457# a_939_2457# 2.64e-19
C3300 a_10711_n62# a_10937_n62# 3.34e-19
C3301 a_16109_1642# a_15767_895# 0.00232f
C3302 VDD_SW_b[7] a_3039_601# 1.99e-20
C3303 a_6539_1642# D[4] 1.68e-19
C3304 x9.A1 a_16488_627# 2e-20
C3305 VDD x2.X 7.42f
C3306 a_1946_n62# a_2566_n88# 8.26e-21
C3307 a_10597_n88# a_12447_n62# 4.56e-21
C3308 a_14096_627# a_15293_601# 1.84e-20
C3309 a_10596_212# a_12680_106# 5.86e-20
C3310 VDD_SW[2] a_14545_627# 9.25e-19
C3311 VDD a_4413_2457# 0.203f
C3312 x2.X a_7649_993# 0.15f
C3313 a_1555_627# a_1233_n88# 7.32e-20
C3314 VDD_SW[7] a_1028_212# 4.35e-19
C3315 a_5165_627# VSS_SW_b[5] 6e-19
C3316 check[5] a_3039_601# 0.00264f
C3317 VSS_SW[3] a_10734_304# 1.97e-20
C3318 a_10596_212# VSS_SW_b[3] 0.00119f
C3319 a_10597_n88# a_11069_122# 0.15f
C3320 a_1256_993# a_1501_122# 1.51e-20
C3321 a_791_627# a_174_n88# 1.08e-19
C3322 x2.X a_11325_1315# 2.32e-19
C3323 x9.X check[4] 5.57e-19
C3324 a_12989_n88# VSS_SW_b[1] 0.00485f
C3325 a_13407_220# VSS_SW[1] 1.77e-20
C3326 x11.X VDD_SW[5] 0.177f
C3327 x9.A1 VDD_SW_b[6] 2.35e-20
C3328 a_3333_601# a_5165_627# 2.42e-20
C3329 a_12433_993# a_12553_n62# 6.88e-22
C3330 a_3807_895# a_6040_993# 1.86e-21
C3331 D[2] a_13906_n62# 0.158f
C3332 VDD_SW_b[6] a_4338_n62# 0.0144f
C3333 a_6285_1642# a_6339_627# 1.92e-20
C3334 a_11987_627# a_12607_601# 0.149f
C3335 D[2] a_12153_627# 0.168f
C3336 D[4] a_8288_909# 8.51e-19
C3337 a_7203_627# a_8516_993# 2.13e-19
C3338 VDD_SW_b[3] a_12607_601# 2.22e-20
C3339 x9.A1 check[3] 0.424f
C3340 D[4] a_7854_220# 1.98e-20
C3341 a_15767_895# VDD_SW[1] 0.00356f
C3342 a_15608_993# a_15715_627# 0.00707f
C3343 a_15855_1642# a_15907_627# 1.92e-20
C3344 x9.A1 a_2831_1315# 0.00507f
C3345 a_8204_212# a_8409_n88# 0.15f
C3346 a_7663_n62# VSS_SW_b[4] 0.0142f
C3347 VSS_SW[4] a_7854_220# 4.25e-19
C3348 a_11071_1642# a_10983_895# 5.45e-19
C3349 a_5289_1289# a_4958_n88# 5.67e-21
C3350 x10.X D[5] 0.00864f
C3351 a_11071_1642# D[3] 0.0682f
C3352 VSS_SW[6] a_3625_n88# 9.92e-21
C3353 x2.X a_10596_212# 0.0128f
C3354 a_16097_304# a_16298_n62# 8.99e-19
C3355 x2.X a_8335_627# 0.00702f
C3356 VDD a_13407_220# 0.00984f
C3357 a_4689_2457# check[4] 0.00137f
C3358 x2.X a_8921_304# 3.34e-19
C3359 a_14825_993# VSS_SW[1] 0.00296f
C3360 x13.X a_8591_895# 0.00658f
C3361 VDD a_8679_1642# 0.191f
C3362 VDD a_1369_n62# 0.0301f
C3363 a_13375_895# D[1] 2.1e-19
C3364 a_13216_993# a_14379_627# 7.56e-20
C3365 D[7] a_1745_304# 8.38e-19
C3366 x9.A1 a_12495_1642# 5.26e-19
C3367 a_13461_1642# a_13216_993# 0.00181f
C3368 a_13216_993# VDD_SW_b[2] 4.35e-20
C3369 D[4] VSS_SW[3] 4.86e-19
C3370 D[6] a_4528_627# 0.00235f
C3371 VDD a_14825_993# 0.18f
C3372 a_12447_n62# a_12638_220# 3.3e-19
C3373 VSS_SW[2] a_13461_122# 2.79e-21
C3374 a_14379_627# a_15464_909# 1.09e-19
C3375 a_14887_1642# D[1] 5.74e-19
C3376 D[1] a_15243_909# 6.78e-19
C3377 VSS_SW_b[3] a_11313_n62# 6.94e-20
C3378 check[0] a_15293_601# 2.14e-19
C3379 D[3] a_12989_n88# 9.65e-22
C3380 x2.X a_941_601# 0.119f
C3381 VDD_SW_b[2] a_15464_909# 1.97e-21
C3382 x17.X a_14545_627# 1.68e-19
C3383 x13.X VDD_SW_b[4] 0.242f
C3384 ready VSS_SW[7] 0.0387f
C3385 a_9949_627# VSS_SW_b[3] 5.82e-19
C3386 x13.X a_9646_90# 0.0273f
C3387 VSS_SW[5] a_6231_220# 6.42e-21
C3388 a_5813_n88# VSS_SW_b[5] 7.55e-19
C3389 a_6017_n88# a_6285_122# 0.206f
C3390 a_13906_n62# VSS_SW_b[1] 2.63e-19
C3391 x9.A1 a_15381_n88# 8.52e-21
C3392 x7.X a_2566_n88# 0.00862f
C3393 x8.X VSS_SW[6] 0.253f
C3394 VSS_SW[7] a_1501_122# 2.79e-21
C3395 a_78_90# VSS_SW_b[7] 0.19f
C3396 a_11325_1642# VDD_SW_b[3] 2.59e-19
C3397 check[1] a_13193_n88# 2.61e-19
C3398 x2.X a_2985_n62# 5.25e-20
C3399 VDD_SW[3] a_12517_993# 6.61e-21
C3400 VDD a_8409_n88# 0.48f
C3401 x16.X a_10983_895# 0.00865f
C3402 a_7369_627# VSS_SW_b[4] 5.23e-20
C3403 a_8117_601# a_8205_n88# 3.89e-19
C3404 a_8591_895# a_8204_212# 0.00165f
C3405 x6.X a_439_1315# 2.41e-19
C3406 x16.X D[3] 7.79e-19
C3407 x2.X a_9949_627# 0.00141f
C3408 a_2585_627# a_3333_601# 0.126f
C3409 VDD a_7252_1467# 0.114f
C3410 a_3039_601# a_2865_993# 0.206f
C3411 x2.X a_1672_909# 4.02e-19
C3412 a_2566_n88# a_3420_212# 0.0319f
C3413 a_2879_n62# a_3112_106# 0.124f
C3414 a_15608_993# a_15853_122# 1.51e-20
C3415 a_15143_627# a_14526_n88# 1.08e-19
C3416 a_6199_895# a_7203_627# 6.86e-19
C3417 a_5725_601# D[4] 9.63e-19
C3418 a_15855_1642# a_15585_n88# 4.63e-19
C3419 D[5] a_8117_601# 2.67e-21
C3420 a_14428_1467# D[1] 0.0177f
C3421 a_6339_627# a_6285_122# 2.54e-20
C3422 a_5725_601# VSS_SW[4] 2.9e-20
C3423 VDD x14.X 0.338f
C3424 a_6199_895# a_6153_n62# 1.65e-20
C3425 x2.X a_2927_1642# 2.62e-19
C3426 a_9644_1467# a_9786_1315# 0.00783f
C3427 x14.X a_7649_993# 1.56e-20
C3428 x18.X a_13216_993# 2.78e-19
C3429 a_3895_1642# a_3333_601# 0.00263f
C3430 VDD_SW[6] a_4977_627# 9.25e-19
C3431 a_4528_627# a_5725_601# 1.71e-20
C3432 x2.X a_5341_993# 5.3e-19
C3433 VDD_SW_b[6] a_5812_212# 2.3e-22
C3434 VDD_SW[6] VSS_SW[5] 0.427f
C3435 x2.X x15.X 0.00458f
C3436 a_218_1315# D[7] 7.54e-19
C3437 D[4] VDD_SW[4] 0.246f
C3438 VDD_SW_b[4] a_8204_212# 0.0416f
C3439 x7.X a_27_627# 2.67e-20
C3440 a_7896_106# a_7769_n62# 0.0256f
C3441 a_7663_n62# a_8140_n62# 1.96e-20
C3442 a_8204_212# a_9646_90# 0.00101f
C3443 VSS_SW_b[4] a_8342_304# 3.58e-20
C3444 a_8205_n88# a_9122_n62# 0.189f
C3445 a_8409_n88# a_8921_304# 6.69e-20
C3446 a_3648_993# a_3504_909# 0.00412f
C3447 a_12433_993# VSS_SW[2] 0.003f
C3448 a_3039_601# a_3551_627# 9.75e-19
C3449 a_2585_627# a_4064_909# 7.17e-20
C3450 a_3333_601# a_3183_627# 0.00926f
C3451 a_2865_993# a_2973_627# 0.00807f
C3452 ready a_3333_601# 5.7e-21
C3453 x9.A1 a_10215_601# 2.81e-20
C3454 a_16109_1315# D[1] 0.00195f
C3455 x9.A1 a_8921_n62# 5.7e-21
C3456 a_14379_627# VDD_SW[1] 3.29e-20
C3457 a_4860_1467# x10.X 0.0876f
C3458 D[1] a_15715_627# 2e-19
C3459 a_10509_601# a_12607_601# 1.55e-20
C3460 a_10983_895# a_12153_627# 2.8e-19
C3461 a_1757_1642# a_1028_212# 1.17e-22
C3462 a_6920_627# VDD_SW[5] 0.0729f
C3463 a_6339_627# a_6147_627# 4.19e-20
C3464 VDD_SW_b[5] a_7203_627# 5.95e-19
C3465 D[3] a_12153_627# 6.4e-21
C3466 VDD_SW_b[5] a_6153_n62# 0.00179f
C3467 VDD_SW_b[7] a_1143_n62# 5.2e-19
C3468 a_9595_627# a_10727_627# 0.00272f
C3469 D[7] a_3112_106# 2.77e-21
C3470 x9.A1 a_16298_n62# 1.9e-20
C3471 VDD a_10680_909# 0.0164f
C3472 a_5271_n62# a_5462_220# 3.24e-19
C3473 VDD_SW_b[2] a_13103_n62# 5.2e-19
C3474 a_4860_1467# D[5] 0.0184f
C3475 a_11987_627# D[1] 1.27e-20
C3476 D[2] a_14379_627# 1e-19
C3477 VDD a_5319_1642# 8.63e-19
C3478 a_174_n88# a_1029_n88# 0.0477f
C3479 a_487_n62# a_1028_212# 0.138f
C3480 check[6] D[6] 3.68e-20
C3481 a_5323_2457# a_5257_993# 8.63e-21
C3482 D[2] VDD_SW_b[2] 0.453f
C3483 a_13461_1642# D[2] 0.0681f
C3484 x2.X a_2468_1467# 3.56e-19
C3485 check[1] a_12607_601# 0.00262f
C3486 x12.X a_7254_90# 0.00259f
C3487 check[2] a_11253_1642# 0.00577f
C3488 VDD a_8591_895# 0.671f
C3489 VDD a_1971_1642# 0.00177f
C3490 a_7823_601# a_8432_993# 0.00189f
C3491 a_7369_627# a_7557_627# 0.189f
C3492 VDD a_13119_627# 6.2e-19
C3493 check[6] a_1685_1642# 0.00577f
C3494 a_2419_627# a_3112_106# 3.88e-21
C3495 D[6] a_2879_n62# 0.00257f
C3496 a_11514_n62# a_12134_n88# 8.26e-21
C3497 x9.A1 VSS_SW_b[4] 2.86e-19
C3498 check[1] a_14857_1289# 5.99e-21
C3499 a_11069_122# a_11313_304# 0.00972f
C3500 VSS_SW_b[3] a_11015_220# 1.12e-20
C3501 a_10801_n88# a_11514_n62# 8.07e-20
C3502 a_10597_n88# a_12038_90# 5.39e-19
C3503 a_5812_212# a_5927_n62# 0.00272f
C3504 a_5504_106# a_6153_n62# 0.00316f
C3505 a_5271_n62# VSS_SW[4] 1.46e-20
C3506 a_9761_627# a_10055_n62# 2.38e-19
C3507 a_10215_601# a_9742_n88# 4.37e-19
C3508 VSS_SW[1] a_14526_n88# 0.00667f
C3509 x10.X a_6285_1642# 2.02e-20
C3510 VSS_SW[3] a_10597_n88# 9.29e-21
C3511 x7.X VDD_SW[7] 0.177f
C3512 x2.X a_6017_n88# 0.00369f
C3513 VDD VDD_SW_b[4] 0.156f
C3514 D[2] a_15072_106# 2.77e-21
C3515 a_12036_1467# VSS_SW[2] 0.0274f
C3516 VDD a_9646_90# 0.189f
C3517 check[5] x10.X 5.87e-19
C3518 a_7649_993# VDD_SW_b[4] 5.9e-21
C3519 a_8117_601# a_8848_909# 0.0016f
C3520 a_12751_627# a_12134_n88# 1.08e-19
C3521 a_13216_993# a_13461_122# 1.51e-20
C3522 a_11325_1642# a_10509_601# 7.12e-21
C3523 a_7823_601# a_7769_n62# 1.07e-20
C3524 a_9644_1467# D[3] 0.0182f
C3525 x2.X a_3039_601# 0.2f
C3526 x6.X a_193_627# 0.00315f
C3527 a_3420_212# a_3369_304# 2.13e-19
C3528 a_3421_n88# a_3070_220# 4.71e-20
C3529 a_3112_106# a_3558_304# 0.00412f
C3530 a_2879_n62# a_3839_220# 1.21e-20
C3531 a_6285_1642# D[5] 0.0682f
C3532 x2.X a_11015_220# 9.52e-19
C3533 x14.X a_9949_627# 6.07e-19
C3534 VDD a_14526_n88# 0.69f
C3535 a_5323_2457# a_5289_1289# 6.83e-20
C3536 check[5] D[5] 3.88e-20
C3537 x9.X a_3807_895# 0.00641f
C3538 check[0] a_14839_n62# 1.32e-20
C3539 a_14379_627# VSS_SW_b[1] 1.08e-19
C3540 D[1] a_15853_122# 0.00923f
C3541 VDD VDD_SW[3] 0.374f
C3542 VDD_SW_b[2] VSS_SW_b[1] 0.0382f
C3543 a_11325_1642# check[1] 1.57e-19
C3544 D[7] D[6] 0.00183f
C3545 a_4811_627# a_5896_909# 1.09e-19
C3546 D[5] a_5675_909# 6.77e-19
C3547 x2.X a_6339_627# 0.0151f
C3548 VDD a_2136_627# 0.194f
C3549 a_8933_1642# a_9154_1315# 0.00783f
C3550 x18.X D[2] 0.00106f
C3551 VDD_SW_b[4] a_10596_212# 2.3e-22
C3552 a_6760_1315# VDD_SW_b[5] 1.32e-20
C3553 VDD a_1256_993# 0.189f
C3554 a_9646_90# a_10596_212# 1.66e-20
C3555 a_27_627# a_193_627# 0.786f
C3556 x2.X a_13072_909# 0.00309f
C3557 x2.X a_2973_627# 3.94e-19
C3558 a_3648_993# VDD_SW[6] 3.28e-20
C3559 a_3421_n88# VSS_SW[5] 9.22e-19
C3560 a_1685_1642# D[7] 5.72e-19
C3561 a_3625_n88# a_3761_n62# 0.0697f
C3562 VSS_SW_b[6] a_3356_n62# 1.68e-19
C3563 VDD_SW_b[3] a_10711_n62# 5.21e-19
C3564 VDD_SW_b[7] VSS_SW_b[6] 0.0382f
C3565 a_2585_627# VSS_SW[6] 0.023f
C3566 a_2419_627# D[6] 0.138f
C3567 x2.X VSS_SW_b[7] 0.0279f
C3568 check[4] a_4862_90# 2.5e-20
C3569 x9.X VDD_SW_b[6] 0.239f
C3570 VDD_SW[3] a_10596_212# 4.35e-19
C3571 a_11123_627# a_10801_n88# 7.32e-20
C3572 a_10824_993# a_10908_993# 0.00857f
C3573 VDD a_3535_n62# 0.00521f
C3574 a_4977_627# a_7369_627# 2.94e-19
C3575 x9.A1 a_7557_627# 4.44e-19
C3576 x16.X a_12178_1315# 8.32e-19
C3577 x2.X a_15511_627# 0.00702f
C3578 a_9761_627# a_10983_895# 0.0494f
C3579 x2.X a_13715_1315# 2.33e-19
C3580 a_15381_n88# a_15585_n88# 0.117f
C3581 VSS_SW[1] a_15329_304# 8.23e-20
C3582 a_15380_212# a_15853_122# 0.159f
C3583 a_15072_106# VSS_SW_b[1] 0.00322f
C3584 check[4] x11.X 0.00964f
C3585 D[3] a_9761_627# 0.168f
C3586 a_9595_627# a_10215_601# 0.149f
C3587 a_4077_1642# D[6] 5.72e-19
C3588 check[5] VSS_SW_b[6] 3.18e-20
C3589 a_1029_n88# a_1166_304# 0.00907f
C3590 a_1028_212# a_1447_220# 2.46e-19
C3591 a_487_n62# a_1946_n62# 3.79e-20
C3592 a_8591_895# a_9949_627# 8.26e-21
C3593 D[7] a_1340_993# 2.53e-19
C3594 a_27_627# a_791_627# 0.00134f
C3595 x3.X check[6] 0.0144f
C3596 x9.A1 a_13375_895# 2.41e-19
C3597 a_12607_601# a_12341_627# 8.07e-20
C3598 a_12153_627# a_12517_993# 0.0018f
C3599 a_12901_601# a_13375_895# 0.265f
C3600 x9.A1 check[2] 0.41f
C3601 a_7369_627# a_9312_627# 1.79e-20
C3602 x27.A a_4528_627# 1.61e-19
C3603 check[5] a_4363_1642# 0.00688f
C3604 x9.A1 a_5223_1315# 0.00507f
C3605 x12.X D[5] 7.76e-19
C3606 VDD a_15329_304# 0.00265f
C3607 D[6] a_3558_304# 9.67e-19
C3608 a_3183_627# VSS_SW[6] 0.0012f
C3609 VDD a_5896_909# 0.0164f
C3610 ready VSS_SW[6] 0.0361f
C3611 a_5812_212# VSS_SW_b[4] 0.00378f
C3612 VDD a_11071_1642# 0.191f
C3613 a_5950_304# VSS_SW[4] 2.77e-20
C3614 x10.X a_2865_993# 1.55e-20
C3615 VSS_SW_b[7] a_1369_n62# 5.35e-19
C3616 x9.A1 a_14887_1642# 5.26e-19
C3617 a_1501_122# VSS_SW[6] 6.66e-20
C3618 a_10055_n62# a_10532_n62# 1.96e-20
C3619 a_10288_106# a_10161_n62# 0.0256f
C3620 check[1] D[1] 3.82e-20
C3621 VDD_SW_b[4] a_9949_627# 9.33e-21
C3622 a_941_601# a_2136_627# 5.61e-19
C3623 a_193_627# VDD_SW[7] 2.07e-20
C3624 check[1] a_12178_1642# 0.00688f
C3625 a_4811_627# VSS_SW_b[5] 1.08e-19
C3626 D[5] a_6285_122# 0.00938f
C3627 x2.X a_7254_90# 0.00368f
C3628 a_941_601# a_1256_993# 0.13f
C3629 a_473_993# a_381_627# 0.0369f
C3630 a_647_601# a_557_993# 6.69e-20
C3631 a_193_627# a_891_909# 0.00276f
C3632 x2.X VDD_SW[2] 0.0327f
C3633 a_8067_909# VDD_SW[4] 1.01e-20
C3634 a_7394_1642# VSS_SW[4] 0.00105f
C3635 VDD VSS_SW[7] 0.636f
C3636 a_13193_n88# a_13329_n62# 0.0697f
C3637 VSS_SW_b[2] a_12924_n62# 1.68e-19
C3638 x30.A VDD_SW[6] 0.0077f
C3639 a_12989_n88# VSS_SW[1] 9.23e-19
C3640 a_3333_601# a_4811_627# 3.81e-19
C3641 a_4149_1642# D[6] 0.0607f
C3642 a_3112_106# a_4958_n88# 1.86e-21
C3643 D[2] a_13461_122# 0.00928f
C3644 x3.A x9.A1 1.27e-19
C3645 a_11987_627# VSS_SW_b[2] 1.08e-19
C3646 VDD_SW_b[3] VSS_SW_b[2] 0.0383f
C3647 a_14545_627# VDD_SW_b[1] 0.00231f
C3648 x20.X a_14545_627# 1.02e-20
C3649 a_15608_993# a_15692_993# 0.00857f
C3650 a_11071_1642# a_10596_212# 1.39e-21
C3651 a_4860_1467# check[5] 1.56e-19
C3652 check[2] a_9742_n88# 5.26e-19
C3653 a_15585_n88# a_16298_n62# 8.07e-20
C3654 VSS_SW_b[1] a_15799_220# 1.12e-20
C3655 a_15853_122# a_16097_304# 0.00972f
C3656 a_1757_1642# x7.X 0.0843f
C3657 a_15072_106# a_15495_n62# 0.00386f
C3658 a_14839_n62# a_15721_n62# 0.00926f
C3659 VDD a_12989_n88# 0.66f
C3660 D[5] a_6147_627# 2e-19
C3661 a_4811_627# VDD_SW[5] 3.29e-20
C3662 x3.X D[7] 1.77e-19
C3663 a_1415_895# VDD_SW_b[7] 0.128f
C3664 x9.A1 a_14428_1467# 0.197f
C3665 a_13715_1642# a_13375_895# 0.00226f
C3666 x12.X a_8117_601# 5e-20
C3667 x17.X a_12680_106# 2.38e-20
C3668 x9.A1 a_4977_627# 3.44e-19
C3669 check[3] a_7896_106# 8.41e-22
C3670 a_9644_1467# x13.X 4.97e-19
C3671 x9.A1 VSS_SW[5] 0.116f
C3672 a_1503_1642# a_1555_627# 1.92e-20
C3673 a_4338_n62# VSS_SW[5] 6.06e-20
C3674 a_3893_122# VSS_SW_b[5] 1.09e-20
C3675 x15.X VDD_SW[3] 0.177f
C3676 x7.X a_487_n62# 0.00192f
C3677 a_5002_1315# VSS_SW[5] 7.96e-19
C3678 check[6] a_1028_212# 3.24e-20
C3679 a_12134_n88# a_12680_106# 0.207f
C3680 a_3807_895# a_3625_n88# 4.26e-19
C3681 a_3333_601# a_3893_122# 2.7e-19
C3682 check[4] a_5813_n88# 2.45e-20
C3683 VDD VSS_SW_b[5] 0.0967f
C3684 VDD x16.X 0.338f
C3685 x9.A1 a_9312_627# 2e-20
C3686 a_14428_1467# a_14570_1642# 0.00557f
C3687 a_8933_1642# D[4] 0.0607f
C3688 a_10597_n88# a_12988_212# 8.02e-22
C3689 a_10596_212# a_12989_n88# 5.48e-21
C3690 x9.A1 a_16109_1315# 0.00496f
C3691 VDD_SW[2] a_14825_993# 7.03e-20
C3692 a_1029_n88# a_2566_n88# 1.98e-19
C3693 VDD a_3333_601# 0.46f
C3694 a_1028_212# a_2879_n62# 2.62e-19
C3695 a_10215_601# a_10041_993# 0.206f
C3696 x16.X a_11325_1315# 2.37e-20
C3697 a_10801_n88# VSS_SW_b[3] 9.21e-19
C3698 a_5257_993# a_5725_601# 0.0633f
C3699 a_4977_627# a_6040_993# 0.0334f
C3700 x2.X x17.X 0.00464f
C3701 a_13461_122# VSS_SW_b[1] 1.09e-20
C3702 a_13906_n62# VSS_SW[1] 6.09e-20
C3703 a_941_601# VSS_SW[7] 2.13e-19
C3704 a_12153_627# VSS_SW[1] 5.36e-21
C3705 a_8205_n88# VSS_SW_b[3] 0.00484f
C3706 a_3895_1642# check[4] 6.17e-21
C3707 x9.A1 a_11987_627# 8.17e-19
C3708 D[2] a_12433_993# 0.00874f
C3709 a_11987_627# a_12901_601# 0.14f
C3710 x9.A1 VDD_SW_b[3] 2.35e-20
C3711 VDD_SW_b[3] a_12901_601# 5.19e-20
C3712 VDD_SW_b[6] a_3625_n88# 0.00132f
C3713 VDD VDD_SW[5] 0.395f
C3714 D[6] a_4958_n88# 4.32e-19
C3715 x2.X a_12134_n88# 0.178f
C3716 VDD_SW[5] a_7649_993# 7.03e-20
C3717 D[4] a_7350_n88# 0.00506f
C3718 a_7203_627# a_7663_n62# 7.27e-19
C3719 a_10103_1642# D[3] 5.74e-19
C3720 VSS_SW[4] a_7350_n88# 0.00677f
C3721 x2.X a_10801_n88# 0.00369f
C3722 x13.X a_9761_627# 1.68e-19
C3723 check[2] a_9595_627# 0.0012f
C3724 x2.X x10.X 3.64e-19
C3725 VDD a_13906_n62# 0.109f
C3726 a_1143_n62# a_1369_n62# 3.34e-19
C3727 VDD a_4064_909# 0.00438f
C3728 VDD a_12153_627# 0.659f
C3729 a_13715_1642# a_14428_1467# 0.00957f
C3730 a_5725_601# a_5943_627# 3.73e-19
C3731 a_5431_601# VDD_SW_b[5] 1.75e-20
C3732 a_7252_1467# a_7254_90# 1e-19
C3733 a_6040_993# a_5575_627# 0.00316f
C3734 check[0] a_14430_90# 2.5e-20
C3735 x2.X a_8205_n88# 0.0213f
C3736 VDD a_7711_1642# 8.63e-19
C3737 check[3] a_7823_601# 0.00263f
C3738 a_27_627# a_1029_n88# 1.06e-19
C3739 D[7] a_1028_212# 0.158f
C3740 x2.X D[5] 0.199f
C3741 a_11071_1642# x15.X 1.31e-19
C3742 a_12680_106# a_12937_304# 0.00857f
C3743 a_12447_n62# a_13126_304# 0.00652f
C3744 VDD a_15767_895# 0.67f
C3745 a_2419_627# a_3283_909# 2.46e-19
C3746 D[6] a_2949_993# 8.11e-19
C3747 a_16109_1642# a_16488_627# 5.9e-19
C3748 D[1] a_15692_993# 2.52e-19
C3749 check[0] a_14857_1289# 0.245f
C3750 a_16323_1642# D[1] 0.00164f
C3751 check[0] a_15608_993# 3.41e-19
C3752 a_14379_627# a_15143_627# 0.00134f
C3753 a_941_601# a_3333_601# 9.37e-21
C3754 a_193_627# a_2773_627# 3.67e-21
C3755 a_1415_895# a_2865_993# 8e-21
C3756 VDD_SW_b[3] a_9742_n88# 3.21e-19
C3757 a_6285_1642# x12.X 1.51e-20
C3758 x13.X a_8677_122# 2.79e-19
C3759 x9.A1 a_15853_122# 3.99e-20
C3760 a_4977_627# a_5812_212# 1.02e-19
C3761 a_5431_601# a_5504_106# 1.01e-19
C3762 a_5257_993# a_5271_n62# 2.63e-19
C3763 a_5725_601# a_4958_n88# 0.00259f
C3764 a_12036_1467# D[2] 0.0182f
C3765 VSS_SW[5] a_5812_212# 5.9e-22
C3766 x9.A1 a_76_1467# 0.197f
C3767 x8.X a_2831_1315# 2.41e-19
C3768 a_193_627# a_487_n62# 2.38e-19
C3769 a_647_601# a_174_n88# 4.37e-19
C3770 check[1] VSS_SW_b[2] 3.19e-20
C3771 VDD_SW[3] a_13072_909# 2.77e-20
C3772 a_15907_627# a_15715_627# 4.19e-20
C3773 x2.X a_12937_304# 0.00168f
C3774 a_16488_627# VDD_SW[1] 0.0729f
C3775 x9.A1 a_3648_993# 4.84e-21
C3776 x20.X VDD_SW_b[1] 0.243f
C3777 a_4528_627# a_3420_212# 6.63e-19
C3778 x2.X VSS_SW_b[6] 0.0278f
C3779 reset x2.X 1.3e-19
C3780 VDD a_5748_n62# 7.87e-19
C3781 a_305_2457# x3.X 0.236f
C3782 a_7203_627# a_7369_627# 0.786f
C3783 a_29_2457# ready 0.0408f
C3784 a_6285_1642# a_6285_122# 1.57e-21
C3785 VDD a_9644_1467# 0.114f
C3786 VDD_SW[7] a_3504_909# 2.77e-20
C3787 VDD_SW_b[7] a_2865_993# 8.2e-21
C3788 x9.A1 a_174_n88# 7.41e-19
C3789 a_14733_627# VSS_SW_b[1] 5.82e-19
C3790 a_1501_122# a_1745_n62# 0.00807f
C3791 a_2470_90# a_2566_n88# 0.0967f
C3792 a_13715_1642# a_13929_1642# 0.00557f
C3793 a_14096_627# D[1] 4.27e-19
C3794 a_13515_627# a_14379_627# 1.09e-19
C3795 x2.X a_8117_601# 0.119f
C3796 a_1555_627# a_1501_122# 2.54e-20
C3797 a_13461_1642# a_13515_627# 1.92e-20
C3798 check[5] a_2865_993# 7.19e-20
C3799 x2.X a_14545_627# 0.0537f
C3800 a_9312_627# a_9595_627# 0.00111f
C3801 x15.X x16.X 0.11f
C3802 VDD a_678_220# 0.00415f
C3803 a_9122_n62# VSS_SW_b[3] 2.62e-19
C3804 a_12553_n62# a_12924_n62# 4.19e-20
C3805 a_3807_895# a_5165_627# 8.26e-21
C3806 VDD_SW_b[6] a_4862_90# 0.00345f
C3807 D[4] a_8516_993# 2.53e-19
C3808 a_7203_627# a_7967_627# 0.00134f
C3809 a_505_1289# a_174_n88# 5.67e-21
C3810 check[2] VSS_SW[2] 1.44e-19
C3811 VSS_SW[4] a_8153_304# 8.35e-20
C3812 a_8204_212# a_8677_122# 0.159f
C3813 a_8205_n88# a_8409_n88# 0.117f
C3814 a_7896_106# VSS_SW_b[4] 0.00322f
C3815 x9.A1 a_10509_601# 0.00103f
C3816 a_10509_601# a_12901_601# 9.37e-21
C3817 a_10983_895# a_12433_993# 8e-21
C3818 a_11240_909# VDD_SW_b[3] 3.4e-20
C3819 a_5289_1289# a_5271_n62# 3.44e-19
C3820 VSS_SW[6] a_3893_122# 2.79e-21
C3821 check[2] a_10041_993# 6.72e-20
C3822 a_9595_627# a_11987_627# 1.63e-20
C3823 x2.X a_8848_909# 4.02e-19
C3824 x11.X check[3] 5.57e-19
C3825 x9.A1 a_2897_1289# 0.104f
C3826 a_9595_627# VDD_SW_b[3] 1.12e-19
C3827 x2.X a_9122_n62# 1.88e-19
C3828 VDD a_10359_627# 1.8e-19
C3829 a_14379_627# VSS_SW[1] 0.0576f
C3830 VDD VSS_SW[6] 0.544f
C3831 a_7252_1467# D[5] 2.96e-19
C3832 VDD_SW_b[2] VSS_SW[1] 0.00248f
C3833 VDD a_6753_1642# 0.00177f
C3834 D[7] a_1946_n62# 0.158f
C3835 a_8679_1642# a_8117_601# 0.00263f
C3836 VDD a_9761_627# 0.659f
C3837 VDD_SW_b[6] a_5165_627# 9.33e-21
C3838 x9.A1 a_4137_n62# 5.7e-21
C3839 x9.A1 check[1] 0.409f
C3840 x2.X a_4860_1467# 2.87e-19
C3841 a_5323_2457# a_6539_1642# 0.00112f
C3842 a_4958_n88# a_5271_n62# 0.245f
C3843 a_12495_1642# D[2] 5.74e-19
C3844 a_4338_n62# a_4137_n62# 3.81e-19
C3845 check[1] a_12901_601# 2.11e-19
C3846 x9.A1 a_7615_1315# 0.00507f
C3847 x15.X a_12153_627# 1.68e-19
C3848 x30.A x9.A1 0.00354f
C3849 D[6] a_3947_627# 0.00431f
C3850 VDD a_14379_627# 0.393f
C3851 check[6] x7.X 0.00967f
C3852 VDD a_13461_1642# 0.191f
C3853 VDD VDD_SW_b[2] 0.156f
C3854 a_15907_627# a_15853_122# 2.54e-20
C3855 a_12038_90# a_12447_n62# 4.24e-20
C3856 x2.X a_1415_895# 0.148f
C3857 a_14545_627# a_14825_993# 0.15f
C3858 check[0] D[1] 0.461f
C3859 x9.A1 a_7203_627# 8.11e-19
C3860 a_10509_601# a_9742_n88# 0.00259f
C3861 a_9761_627# a_10596_212# 1.02e-19
C3862 VSS_SW[1] a_15072_106# 4.61e-19
C3863 a_6017_n88# VSS_SW_b[5] 9.2e-19
C3864 VSS_SW[3] a_11069_122# 2.79e-21
C3865 x7.X a_2879_n62# 4.41e-20
C3866 VSS_SW[7] VSS_SW_b[7] 0.0072f
C3867 D[2] a_15381_n88# 9.66e-22
C3868 a_12341_627# VSS_SW_b[2] 6.02e-19
C3869 x2.X a_3356_n62# 3.67e-20
C3870 x8.X a_1978_1315# 3.75e-20
C3871 VDD a_8677_122# 0.313f
C3872 a_12036_1467# D[3] 2.97e-19
C3873 a_8117_601# a_8409_n88# 0.00251f
C3874 a_8591_895# a_8205_n88# 6.35e-19
C3875 a_8432_993# a_8204_212# 8.94e-21
C3876 x2.X a_10125_993# 5.31e-19
C3877 a_5319_1642# D[5] 5.74e-19
C3878 x2.X a_11514_n62# 1.83e-19
C3879 a_3039_601# a_3333_601# 0.199f
C3880 x2.X VDD_SW_b[7] 7.38e-19
C3881 a_2585_627# a_3807_895# 0.0494f
C3882 VDD a_15072_106# 0.356f
C3883 x9.X a_4977_627# 1.69e-19
C3884 check[4] a_4811_627# 0.0012f
C3885 a_2879_n62# a_3420_212# 0.138f
C3886 x2.X a_6285_1642# 0.00651f
C3887 a_2566_n88# a_3421_n88# 0.0477f
C3888 x9.X VSS_SW[5] 0.149f
C3889 a_6199_895# D[4] 2.17e-19
C3890 a_6040_993# a_7203_627# 7.46e-20
C3891 a_6199_895# VSS_SW[4] 7.03e-21
C3892 check[0] a_15380_212# 3.24e-20
C3893 x2.X check[5] 0.167f
C3894 x18.X VSS_SW[1] 0.253f
C3895 x17.X a_14526_n88# 0.00864f
C3896 x14.X a_8117_601# 0.0013f
C3897 a_941_601# VSS_SW[6] 2.81e-20
C3898 a_4413_2457# check[5] 8.52e-19
C3899 a_13715_1642# check[1] 0.318f
C3900 a_1415_895# a_1369_n62# 1.65e-20
C3901 a_3895_1642# a_3807_895# 5.45e-19
C3902 VDD_SW[6] a_5431_601# 7.64e-20
C3903 x2.X a_5675_909# 0.00137f
C3904 VDD_SW_b[6] a_5813_n88# 2.44e-21
C3905 x2.X a_12751_627# 0.0388f
C3906 a_439_1315# D[7] 0.00202f
C3907 a_4689_2457# a_4977_627# 1.38e-20
C3908 a_4689_2457# VSS_SW[5] 0.0227f
C3909 VDD_SW_b[4] a_8205_n88# 0.0406f
C3910 x7.X D[7] 0.1f
C3911 a_7663_n62# a_8319_n62# 3.73e-19
C3912 a_7896_106# a_8140_n62# 0.00707f
C3913 a_8677_122# a_8921_304# 0.00972f
C3914 a_8205_n88# a_9646_90# 5.39e-19
C3915 a_8409_n88# a_9122_n62# 8.07e-20
C3916 VSS_SW_b[4] a_8623_220# 1.12e-20
C3917 a_3648_993# a_3732_993# 0.00857f
C3918 a_2585_627# VDD_SW_b[6] 0.00226f
C3919 VDD x18.X 0.338f
C3920 a_11987_627# VSS_SW[2] 0.0579f
C3921 ready a_3807_895# 2.44e-19
C3922 VDD_SW_b[3] VSS_SW[2] 0.00249f
C3923 VDD_SW_b[5] D[4] 1.57e-19
C3924 VDD_SW_b[5] VSS_SW[4] 0.00249f
C3925 a_10041_993# VDD_SW_b[3] 4.92e-21
C3926 a_10509_601# a_11240_909# 0.0016f
C3927 VDD_SW_b[7] a_1369_n62# 0.00179f
C3928 x2.X a_78_90# 0.00367f
C3929 D[3] a_10727_627# 6.13e-19
C3930 x2.X x20.X 1.55e-19
C3931 x2.X VDD_SW_b[1] 6.68e-19
C3932 a_9761_627# a_9949_627# 0.189f
C3933 check[3] D[3] 3.87e-20
C3934 a_15381_n88# VSS_SW_b[1] 7.59e-19
C3935 VSS_SW[1] a_15799_220# 6.42e-21
C3936 a_15585_n88# a_15853_122# 0.206f
C3937 a_9595_627# a_10509_601# 0.14f
C3938 D[7] a_3420_212# 5.78e-20
C3939 VDD a_10532_n62# 7.87e-19
C3940 x9.X a_4370_1315# 0.00145f
C3941 x7.X a_2419_627# 0.00295f
C3942 a_720_106# a_1028_212# 0.14f
C3943 VDD check[4] 1.67f
C3944 a_487_n62# a_1029_n88# 0.125f
C3945 a_13515_627# a_13461_122# 2.54e-20
C3946 a_5323_2457# a_5725_601# 4.01e-19
C3947 x9.A1 a_12341_627# 4.11e-19
C3948 a_12433_993# a_12517_993# 0.00972f
C3949 a_12901_601# a_12341_627# 1.15e-20
C3950 a_12607_601# a_12851_909# 0.0104f
C3951 a_13375_895# a_13216_993# 0.207f
C3952 a_12153_627# a_13072_909# 0.00907f
C3953 VDD a_8432_993# 0.189f
C3954 ready VDD_SW_b[6] 4.25e-20
C3955 x2.X a_11123_627# 0.0151f
C3956 a_8117_601# a_8591_895# 0.265f
C3957 a_7823_601# a_7557_627# 8.07e-20
C3958 a_7369_627# a_7733_993# 0.0018f
C3959 check[6] a_193_627# 5.41e-19
C3960 VDD a_15799_220# 0.00984f
C3961 x15.X a_9761_627# 1.08e-20
C3962 x2.X x12.X 3.64e-19
C3963 D[6] a_3112_106# 8.76e-19
C3964 a_2419_627# a_3420_212# 6.99e-20
C3965 VDD a_10103_1642# 8.63e-19
C3966 a_10288_106# a_10711_n62# 0.00386f
C3967 a_10055_n62# a_10937_n62# 0.00926f
C3968 a_5813_n88# a_5927_n62# 2.14e-20
C3969 a_5504_106# VSS_SW[4] 9.06e-21
C3970 a_5812_212# a_6153_n62# 0.00134f
C3971 check[1] a_13643_1642# 0.00577f
C3972 a_10215_601# a_10055_n62# 0.0026f
C3973 a_9742_n88# a_10246_220# 0.00869f
C3974 a_8861_1642# D[4] 5.72e-19
C3975 x11.X VSS_SW_b[4] 0.017f
C3976 x2.X a_6285_122# 0.0043f
C3977 VSS_SW_b[2] a_13329_n62# 5.34e-19
C3978 a_13461_122# VSS_SW[1] 6.77e-20
C3979 VDD a_7769_n62# 0.0133f
C3980 a_8432_993# a_8335_627# 0.00386f
C3981 a_7203_627# a_9595_627# 1.74e-20
C3982 a_8591_895# a_8848_909# 0.00869f
C3983 a_7557_627# a_7757_627# 3.81e-19
C3984 a_8117_601# VDD_SW_b[4] 0.00623f
C3985 a_7649_993# a_7769_n62# 6.88e-22
C3986 a_8591_895# a_9122_n62# 4.06e-19
C3987 a_2468_1467# VSS_SW[6] 0.0274f
C3988 x2.X a_2865_993# 0.15f
C3989 x6.X a_647_601# 2.4e-20
C3990 x9.A1 a_2566_n88# 7.4e-19
C3991 a_4860_1467# a_5319_1642# 6.64e-19
C3992 a_3420_212# a_3558_304# 1.09e-19
C3993 a_14825_993# VDD_SW_b[1] 5.89e-21
C3994 a_15293_601# a_16024_909# 0.0016f
C3995 a_11071_1642# a_10801_n88# 4.63e-19
C3996 x12.X a_8679_1642# 1.98e-20
C3997 a_15381_n88# a_15495_n62# 2.14e-20
C3998 a_15380_212# a_15721_n62# 0.00134f
C3999 VDD a_13461_122# 0.313f
C4000 VDD a_29_2457# 0.211f
C4001 a_14545_627# a_14526_n88# 4.91e-19
C4002 x2.X a_6147_627# 0.00111f
C4003 x9.A1 x6.X 6.9e-19
C4004 D[5] a_5896_909# 8.53e-19
C4005 a_4811_627# a_6124_993# 2.13e-19
C4006 VDD a_1555_627# 6.99e-19
C4007 x9.A1 a_14096_627# 2e-20
C4008 VDD a_381_627# 0.11f
C4009 x17.X a_12989_n88# 0.019f
C4010 a_12901_601# a_14096_627# 5.61e-19
C4011 a_12153_627# VDD_SW[2] 2.07e-20
C4012 a_8848_909# VDD_SW_b[4] 3.66e-20
C4013 VDD_SW_b[4] a_9122_n62# 0.0144f
C4014 a_27_627# a_647_601# 0.149f
C4015 D[7] a_193_627# 0.168f
C4016 x2.X a_3551_627# 0.00702f
C4017 a_4149_1642# a_3420_212# 1.17e-22
C4018 a_3625_n88# VSS_SW[5] 8.78e-20
C4019 a_3893_122# a_3761_n62# 0.025f
C4020 VSS_SW_b[6] a_3535_n62# 5.24e-19
C4021 a_12447_n62# a_12988_212# 0.138f
C4022 a_12134_n88# a_12989_n88# 0.0477f
C4023 a_12036_1467# a_12178_1315# 0.00783f
C4024 x6.X a_505_1289# 1.51e-19
C4025 a_3039_601# VSS_SW[6] 6.25e-19
C4026 x9.A1 a_27_627# 8.16e-19
C4027 VDD a_3761_n62# 0.0301f
C4028 a_10509_601# VSS_SW[2] 2.89e-20
C4029 a_10983_895# a_10937_n62# 1.65e-20
C4030 VDD_SW[2] a_15767_895# 1.27e-20
C4031 a_10041_993# a_10509_601# 0.0633f
C4032 a_193_627# a_2419_627# 1.58e-20
C4033 a_6539_1642# a_5725_601# 7.56e-21
C4034 D[3] a_10215_601# 0.00583f
C4035 VSS_SW_b[7] a_678_220# 5.34e-20
C4036 a_1233_n88# a_1166_304# 9.46e-19
C4037 a_1029_n88# a_1447_220# 0.00276f
C4038 a_1028_212# a_1745_304# 4.45e-20
C4039 a_174_n88# a_593_n62# 0.0383f
C4040 a_487_n62# a_2470_90# 6.12e-21
C4041 a_27_627# a_581_627# 0.00206f
C4042 a_2897_1289# x9.X 1.75e-20
C4043 a_7252_1467# x12.X 0.0876f
C4044 check[1] VSS_SW[2] 0.0496f
C4045 D[2] a_13375_895# 0.0294f
C4046 a_11987_627# a_13216_993# 0.14f
C4047 check[2] D[2] 3.87e-20
C4048 a_505_1289# a_27_627# 0.00104f
C4049 a_15243_909# VDD_SW[1] 1.01e-20
C4050 x2.X a_12680_106# 0.0385f
C4051 VDD a_6124_993# 0.00281f
C4052 D[6] a_3839_220# 7.11e-19
C4053 a_2973_627# VSS_SW[6] 3.79e-19
C4054 check[3] x13.X 0.00968f
C4055 a_11539_1642# D[3] 0.00162f
C4056 a_9595_627# a_12341_627# 4.46e-21
C4057 x2.X VSS_SW_b[3] 0.0279f
C4058 a_14945_n62# a_15316_n62# 4.19e-20
C4059 VDD a_12433_993# 0.18f
C4060 a_6231_220# VSS_SW[4] 1.57e-20
C4061 a_5813_n88# VSS_SW_b[4] 0.00486f
C4062 x10.X a_3333_601# 0.00124f
C4063 a_14733_627# VSS_SW[1] 0.00595f
C4064 x9.A1 a_218_1642# 8.64e-19
C4065 a_13715_1642# a_14096_627# 5.84e-19
C4066 VDD a_9147_1642# 0.00177f
C4067 x9.A1 check[0] 0.407f
C4068 a_647_601# VDD_SW[7] 2.07e-20
C4069 a_1415_895# a_2136_627# 0.0967f
C4070 a_941_601# a_1555_627# 0.0526f
C4071 reset VSS_SW[7] 0.0145f
C4072 x17.X a_13906_n62# 0.0016f
C4073 x9.A1 a_10007_1315# 0.00504f
C4074 x2.X a_5377_n62# 5.57e-20
C4075 a_941_601# a_381_627# 1.24e-20
C4076 a_193_627# a_1112_909# 0.00907f
C4077 a_473_993# a_557_993# 0.00972f
C4078 a_647_601# a_891_909# 0.0104f
C4079 a_13072_909# VDD_SW_b[2] 4.69e-21
C4080 D[5] VSS_SW_b[5] 5.31e-19
C4081 x17.X a_12153_627# 1.13e-20
C4082 a_1415_895# a_1256_993# 0.207f
C4083 a_12751_627# a_13119_627# 3.34e-19
C4084 a_8288_909# VDD_SW[4] 2.82e-20
C4085 a_3807_895# a_4811_627# 6.86e-19
C4086 a_3333_601# D[5] 9.63e-19
C4087 D[6] a_5725_601# 2.67e-21
C4088 a_4689_2457# x30.A 0.236f
C4089 a_4413_2457# x2.X 0.00426f
C4090 VDD a_14733_627# 0.109f
C4091 VDD a_15855_1642# 0.191f
C4092 a_12988_212# a_13126_304# 1.09e-19
C4093 a_3420_212# a_4958_n88# 6.15e-19
C4094 x9.A1 VDD_SW[7] 0.0329f
C4095 a_12153_627# a_12134_n88# 4.91e-19
C4096 VDD_SW_b[5] a_8067_909# 2.62e-21
C4097 VDD_SW_b[5] a_6529_n62# 5.22e-19
C4098 check[0] a_14570_1642# 0.00688f
C4099 a_14379_627# a_15511_627# 0.00272f
C4100 check[2] a_10055_n62# 1.35e-20
C4101 VDD_SW_b[7] a_2136_627# 0.185f
C4102 D[5] VDD_SW[5] 0.245f
C4103 VDD_SW[4] a_10459_909# 2.16e-20
C4104 a_1256_993# VDD_SW_b[7] 4.35e-20
C4105 a_14428_1467# D[2] 2.85e-19
C4106 VDD_SW[4] VSS_SW[3] 0.429f
C4107 x9.A1 a_5431_601# 3.62e-20
C4108 check[3] a_8204_212# 3.2e-20
C4109 a_3947_627# a_3755_627# 4.19e-20
C4110 a_4528_627# VDD_SW[6] 0.0729f
C4111 VDD_SW_b[6] a_4811_627# 5.96e-19
C4112 a_4862_90# VSS_SW[5] 0.082f
C4113 x2.X a_13407_220# 9.61e-19
C4114 x7.X a_720_106# 2.38e-20
C4115 check[6] a_1029_n88# 2.51e-20
C4116 x11.X a_4977_627# 1.08e-20
C4117 x2.X a_8679_1642# 0.00649f
C4118 VDD a_12036_1467# 0.114f
C4119 a_3807_895# a_3893_122# 4.53e-22
C4120 a_3648_993# a_3625_n88# 1.86e-19
C4121 check[4] a_6017_n88# 2.58e-19
C4122 x9.A1 a_8731_627# 5.21e-20
C4123 a_14570_1315# VSS_SW[1] 7.95e-19
C4124 x20.X a_14526_n88# 1.53e-21
C4125 a_13715_1642# check[0] 1.46e-19
C4126 VDD_SW_b[1] a_14526_n88# 3.21e-19
C4127 a_11325_1642# a_11546_1315# 0.00783f
C4128 a_305_2457# a_193_627# 8.93e-22
C4129 VDD_SW[2] a_14379_627# 0.0865f
C4130 VDD a_3807_895# 0.671f
C4131 a_1028_212# a_3112_106# 5.86e-20
C4132 a_1029_n88# a_2879_n62# 4.56e-21
C4133 a_1745_304# a_1946_n62# 8.99e-19
C4134 VDD_SW_b[2] VDD_SW[2] 3.64e-19
C4135 a_4977_627# a_5165_627# 0.189f
C4136 a_5431_601# a_6040_993# 0.00189f
C4137 x2.X a_14825_993# 0.15f
C4138 a_5165_627# VSS_SW[5] 0.00596f
C4139 a_9742_n88# a_10288_106# 0.207f
C4140 a_8409_n88# VSS_SW_b[3] 4.04e-20
C4141 VDD a_14570_1315# 4.95e-19
C4142 VDD a_16488_627# 0.193f
C4143 check[4] a_6339_627# 3.96e-19
C4144 a_11987_627# D[2] 0.137f
C4145 D[6] a_5271_n62# 1.56e-21
C4146 a_12341_627# VSS_SW[2] 0.00596f
C4147 VDD_SW_b[6] a_3893_122# 0.00445f
C4148 x9.A1 a_10824_993# 4.84e-21
C4149 VDD_SW_b[3] D[2] 1.57e-19
C4150 VDD_SW[5] a_8117_601# 2.46e-20
C4151 check[0] a_15907_627# 4.05e-19
C4152 x18.X a_13715_1315# 1.47e-20
C4153 a_7203_627# a_7896_106# 3.88e-21
C4154 check[2] a_10983_895# 0.00271f
C4155 D[4] a_7663_n62# 0.00257f
C4156 VSS_SW[4] a_7663_n62# 3.44e-19
C4157 a_6730_n62# VSS_SW_b[4] 2.78e-19
C4158 check[2] D[3] 0.463f
C4159 VDD VDD_SW_b[6] 0.156f
C4160 a_10073_1289# VSS_SW[3] 0.00187f
C4161 x9.A1 a_2610_1642# 8.62e-19
C4162 a_14428_1467# VSS_SW_b[1] 2.13e-19
C4163 a_5725_601# a_6456_909# 0.0016f
C4164 a_5257_993# VDD_SW_b[5] 4.92e-21
C4165 a_939_2457# a_27_627# 1.42e-20
C4166 VDD a_10727_627# 6.2e-19
C4167 x2.X a_8409_n88# 0.00369f
C4168 VDD check[3] 1.64f
C4169 a_4860_1467# VSS_SW_b[5] 2.11e-19
C4170 check[3] a_7649_993# 6.94e-20
C4171 a_12153_627# a_14545_627# 3.26e-19
C4172 x2.X a_7252_1467# 2.92e-19
C4173 check[1] a_13216_993# 2.87e-19
C4174 a_13929_1642# D[2] 0.00166f
C4175 a_27_627# a_1233_n88# 0.00204f
C4176 D[7] a_1029_n88# 0.158f
C4177 x2.X x14.X 3.61e-19
C4178 D[6] a_3283_909# 6.77e-19
C4179 a_2419_627# a_3504_909# 1.09e-19
C4180 VDD a_12495_1642# 8.63e-19
C4181 a_11514_n62# a_12989_n88# 3.67e-21
C4182 a_12038_90# a_12988_212# 2.02e-20
C4183 a_10734_304# VSS_SW_b[2] 1.09e-20
C4184 a_14999_601# a_15293_601# 0.199f
C4185 a_14545_627# a_15767_895# 0.0494f
C4186 x18.X VDD_SW[2] 0.305f
C4187 x17.X a_14379_627# 0.00295f
C4188 a_1415_895# a_3333_601# 1.42e-20
C4189 a_13461_1642# x17.X 1.37e-19
C4190 x17.X VDD_SW_b[2] 0.242f
C4191 VDD_SW_b[3] a_10055_n62# 5.23e-19
C4192 x9.X a_2566_n88# 1.49e-21
C4193 a_9761_627# a_10801_n88# 8.75e-19
C4194 VSS_SW[1] a_15381_n88# 9.29e-21
C4195 a_9595_627# a_10288_106# 3.88e-21
C4196 a_5725_601# a_5271_n62# 3.74e-20
C4197 a_5257_993# a_5504_106# 4.96e-20
C4198 a_5431_601# a_5812_212# 4.51e-19
C4199 a_4977_627# a_5813_n88# 1.27e-19
C4200 x9.A1 a_1757_1642# 0.195f
C4201 a_8679_1642# a_8409_n88# 4.63e-19
C4202 VSS_SW[5] a_5813_n88# 9.3e-21
C4203 a_647_601# a_487_n62# 0.0026f
C4204 a_473_993# a_174_n88# 8.71e-20
C4205 a_78_90# VSS_SW[7] 0.082f
C4206 a_8204_212# a_8921_n62# 0.00206f
C4207 a_12465_1289# a_12447_n62# 3.44e-19
C4208 VDD_SW_b[2] a_12134_n88# 3.21e-19
C4209 a_2585_627# a_4977_627# 2.94e-19
C4210 x9.A1 a_2773_627# 4.11e-19
C4211 a_11071_1642# a_11123_627# 1.92e-20
C4212 a_3947_627# a_3420_212# 7.07e-21
C4213 a_2585_627# VSS_SW[5] 5.1e-21
C4214 x8.X a_2897_1289# 1.51e-19
C4215 VDD a_5927_n62# 0.00521f
C4216 a_7203_627# a_7823_601# 0.149f
C4217 D[4] a_7369_627# 0.168f
C4218 x2.X a_10680_909# 0.00309f
C4219 a_6753_1642# D[5] 0.00164f
C4220 a_8679_1642# x14.X 9.51e-21
C4221 x3.A ready 0.038f
C4222 x27.A D[6] 0.00836f
C4223 VDD a_15381_n88# 0.659f
C4224 a_939_2457# VDD_SW[7] 0.0315f
C4225 a_7369_627# VSS_SW[4] 0.023f
C4226 x2.X a_5319_1642# 2.62e-19
C4227 VDD_SW_b[7] a_3333_601# 8.35e-20
C4228 x9.A1 a_487_n62# 1.53e-20
C4229 VSS_SW_b[7] a_1745_n62# 6.94e-20
C4230 a_2470_90# a_2879_n62# 4.24e-20
C4231 check[0] a_15585_n88# 2.51e-19
C4232 x2.X a_8591_895# 0.148f
C4233 a_4977_627# a_6920_627# 2e-20
C4234 a_12036_1467# x15.X 4.97e-19
C4235 VDD_SW_b[5] a_4958_n88# 3.23e-19
C4236 check[5] a_3333_601# 2.14e-19
C4237 a_381_627# VSS_SW_b[7] 5.82e-19
C4238 VDD_SW_b[4] VSS_SW_b[3] 0.0382f
C4239 a_9312_627# D[3] 4.28e-19
C4240 a_8731_627# a_9595_627# 1.09e-19
C4241 VDD a_977_304# 0.00269f
C4242 a_9646_90# VSS_SW_b[3] 0.19f
C4243 x2.X a_13119_627# 0.00702f
C4244 a_7681_1289# a_7350_n88# 5.67e-21
C4245 VDD_SW_b[6] a_2985_n62# 4.77e-19
C4246 a_12680_106# a_14526_n88# 1.86e-21
C4247 ready VSS_SW[5] 2e-19
C4248 a_7203_627# a_7757_627# 0.00206f
C4249 a_505_1289# a_487_n62# 3.44e-19
C4250 a_7967_627# VSS_SW[4] 0.0012f
C4251 D[4] a_8342_304# 9.67e-19
C4252 a_8205_n88# a_8677_122# 0.15f
C4253 a_8204_212# VSS_SW_b[4] 0.00119f
C4254 VSS_SW[4] a_8342_304# 1.97e-20
C4255 a_5289_1289# a_5504_106# 5.3e-21
C4256 VSS_SW[6] VSS_SW_b[6] 0.0072f
C4257 a_10983_895# a_11987_627# 6.86e-19
C4258 a_10509_601# D[2] 9.63e-19
C4259 x2.X VDD_SW_b[4] 7.42e-19
C4260 a_5675_909# VDD_SW[5] 1.01e-20
C4261 D[3] a_11987_627# 9.94e-20
C4262 x17.X x18.X 0.109f
C4263 a_10983_895# VDD_SW_b[3] 0.129f
C4264 x2.X a_9646_90# 0.00368f
C4265 D[3] VDD_SW_b[3] 0.453f
C4266 a_15853_122# VSS_SW_b[1] 7.15e-19
C4267 a_9595_627# a_10824_993# 0.14f
C4268 VDD a_10937_n62# 0.0301f
C4269 D[7] a_2470_90# 8.78e-19
C4270 a_8679_1642# a_8591_895# 5.45e-19
C4271 VDD a_10215_601# 0.313f
C4272 a_8117_601# a_9761_627# 6.5e-20
C4273 x2.X a_14526_n88# 0.178f
C4274 a_4958_n88# a_5504_106# 0.207f
C4275 check[1] D[2] 0.46f
C4276 VDD a_1978_1315# 3.89e-19
C4277 a_12153_627# a_12751_627# 6.04e-20
C4278 a_12901_601# a_12851_909# 1.21e-20
C4279 x2.X VDD_SW[3] 0.0327f
C4280 D[6] a_3755_627# 2e-19
C4281 a_2419_627# VDD_SW[6] 3.29e-20
C4282 x13.X check[2] 5.59e-19
C4283 VDD a_16298_n62# 0.109f
C4284 x2.X a_2136_627# 4.01e-19
C4285 x2.X a_1256_993# 0.187f
C4286 VDD a_11539_1642# 0.00177f
C4287 a_2419_627# a_2470_90# 6.13e-19
C4288 a_14379_627# a_14545_627# 0.786f
C4289 x9.A1 a_12399_1315# 0.00504f
C4290 x9.A1 D[4] 0.268f
C4291 a_10596_212# a_10937_n62# 0.00134f
C4292 a_10597_n88# a_10711_n62# 2.14e-20
C4293 a_10288_106# VSS_SW[2] 9.05e-21
C4294 VDD_SW_b[2] a_14545_627# 0.00329f
C4295 x9.A1 VSS_SW[4] 0.403f
C4296 a_10509_601# a_10055_n62# 3.74e-20
C4297 a_10041_993# a_10288_106# 4.96e-20
C4298 a_10215_601# a_10596_212# 4.51e-19
C4299 a_6285_122# VSS_SW_b[5] 7.14e-19
C4300 x10.X check[4] 0.00903f
C4301 x12.X VDD_SW[5] 0.305f
C4302 x11.X a_7203_627# 0.00295f
C4303 x9.A1 a_4528_627# 2e-20
C4304 VDD VSS_SW_b[4] 0.0968f
C4305 a_6539_1642# a_6467_1642# 6.64e-19
C4306 a_8117_601# a_8677_122# 2.7e-19
C4307 a_8591_895# a_8409_n88# 4.26e-19
C4308 x20.X a_15767_895# 0.00655f
C4309 a_7350_n88# a_7854_220# 0.00869f
C4310 a_15767_895# VDD_SW_b[1] 0.128f
C4311 a_2585_627# a_3648_993# 0.0334f
C4312 a_2865_993# a_3333_601# 0.0633f
C4313 check[4] D[5] 0.461f
C4314 a_2879_n62# a_3421_n88# 0.125f
C4315 a_3112_106# a_3420_212# 0.14f
C4316 a_4811_627# a_7557_627# 4.46e-21
C4317 VSS_SW_b[1] a_15316_n62# 1.68e-19
C4318 a_15585_n88# a_15721_n62# 0.0697f
C4319 x14.X a_8591_895# 0.00863f
C4320 a_1415_895# VSS_SW[6] 7.03e-21
C4321 a_14825_993# a_14526_n88# 8.71e-20
C4322 a_14999_601# a_14839_n62# 0.0026f
C4323 a_3895_1642# a_3648_993# 0.00176f
C4324 x2.X a_15329_304# 0.00168f
C4325 VDD_SW[6] a_5257_993# 7.03e-20
C4326 a_4149_1642# VDD_SW[6] 0.00511f
C4327 x2.X a_5896_909# 0.00309f
C4328 x17.X a_13461_122# 2.79e-19
C4329 a_12433_993# VDD_SW[2] 4.17e-21
C4330 a_13375_895# a_13515_627# 0.0383f
C4331 a_12901_601# a_13323_627# 1.96e-20
C4332 a_1757_1315# D[7] 0.00195f
C4333 a_939_2457# a_1757_1642# 0.0012f
C4334 ready a_76_1467# 3.18e-21
C4335 x2.X a_11071_1642# 0.00647f
C4336 VDD_SW_b[4] a_8409_n88# 0.00132f
C4337 D[4] a_9742_n88# 4.32e-19
C4338 a_7896_106# a_8319_n62# 0.00386f
C4339 a_7663_n62# a_8545_n62# 0.00926f
C4340 a_7350_n88# VSS_SW[3] 4.28e-21
C4341 a_3039_601# VDD_SW_b[6] 1.75e-20
C4342 a_3333_601# a_3551_627# 3.73e-19
C4343 a_3648_993# a_3183_627# 0.00316f
C4344 a_8677_122# a_9122_n62# 0.0369f
C4345 a_939_2457# a_2773_627# 1.54e-21
C4346 a_12680_106# a_12989_n88# 0.0327f
C4347 a_12447_n62# a_13193_n88# 0.199f
C4348 a_12134_n88# a_13461_122# 4.59e-22
C4349 a_16109_1642# a_16323_1642# 0.00557f
C4350 a_10597_n88# VSS_SW_b[2] 0.00487f
C4351 x18.X a_14545_627# 0.00314f
C4352 VDD_SW_b[7] VSS_SW[6] 0.00248f
C4353 VDD_SW[2] a_14733_627# 6.11e-20
C4354 x14.X VDD_SW_b[4] 7.27e-19
C4355 x13.X a_9312_627# 0.0338f
C4356 x2.X VSS_SW[7] 0.0813f
C4357 x14.X a_9646_90# 0.00259f
C4358 a_10509_601# a_10983_895# 0.265f
C4359 a_10215_601# a_9949_627# 8.07e-20
C4360 a_9761_627# a_10125_993# 0.0018f
C4361 D[3] a_10509_601# 0.0191f
C4362 D[7] a_3421_n88# 9.66e-22
C4363 a_2897_1289# a_2585_627# 0.00323f
C4364 a_5504_106# a_5761_304# 0.00857f
C4365 a_13906_n62# a_13705_n62# 3.81e-19
C4366 a_5271_n62# a_5950_304# 0.00652f
C4367 check[5] VSS_SW[6] 0.0366f
C4368 x7.X D[6] 2.1e-19
C4369 a_720_106# a_1029_n88# 0.0327f
C4370 a_174_n88# a_1501_122# 4.59e-22
C4371 a_487_n62# a_1233_n88# 0.199f
C4372 a_5323_2457# a_6199_895# 0.00152f
C4373 a_11325_1642# a_11704_627# 5.9e-19
C4374 a_13375_895# VSS_SW[1] 7.03e-21
C4375 VDD a_7557_627# 0.109f
C4376 D[2] a_12341_627# 0.161f
C4377 a_11987_627# a_12517_993# 4.45e-20
C4378 a_16323_1642# VDD_SW[1] 5.32e-19
C4379 a_7369_627# a_8067_909# 0.00276f
C4380 a_7823_601# a_7733_993# 6.69e-20
C4381 a_2897_1289# a_3895_1642# 0.0146f
C4382 x2.X a_12989_n88# 0.0207f
C4383 a_7649_993# a_7557_627# 0.0369f
C4384 a_8117_601# a_8432_993# 0.13f
C4385 check[6] a_647_601# 0.00263f
C4386 a_15143_627# a_15715_627# 2.46e-21
C4387 a_8933_1642# VDD_SW[4] 0.00511f
C4388 check[1] D[3] 6.16e-20
C4389 a_2419_627# a_3421_n88# 1.06e-19
C4390 D[6] a_3420_212# 0.158f
C4391 a_16298_n62# a_16097_n62# 3.81e-19
C4392 x11.X a_6760_1315# 0.00143f
C4393 VDD a_13375_895# 0.671f
C4394 VDD check[2] 1.64f
C4395 a_5812_212# VSS_SW[4] 0.0872f
C4396 a_6017_n88# a_5927_n62# 9.75e-19
C4397 VSS_SW_b[5] a_5377_n62# 0.00334f
C4398 VDD_SW_b[4] a_10680_909# 3.95e-21
C4399 a_5813_n88# a_6153_n62# 6.04e-20
C4400 ready a_2897_1289# 4.05e-20
C4401 x9.A1 check[6] 0.411f
C4402 a_5323_2457# VDD_SW_b[5] 1.07e-20
C4403 a_10055_n62# a_10246_220# 3.24e-19
C4404 a_4811_627# a_4977_627# 0.786f
C4405 a_4811_627# VSS_SW[5] 0.0578f
C4406 x2.X VSS_SW_b[5] 0.0278f
C4407 x2.X x16.X 3.66e-19
C4408 VDD a_8140_n62# 7.87e-19
C4409 D[4] a_9595_627# 1e-19
C4410 a_8591_895# VDD_SW_b[4] 0.129f
C4411 a_7203_627# D[3] 1.27e-20
C4412 a_9312_627# a_8204_212# 6.63e-19
C4413 x8.X a_27_627# 0.00117f
C4414 a_12988_212# a_13705_304# 4.45e-20
C4415 a_13193_n88# a_13126_304# 9.46e-19
C4416 VDD a_14887_1642# 8.63e-19
C4417 a_12989_n88# a_13407_220# 0.00276f
C4418 VSS_SW_b[2] a_12638_220# 5.56e-20
C4419 VDD a_15243_909# 0.00984f
C4420 a_12447_n62# a_14430_90# 6.12e-21
C4421 ready x30.A 0.00174f
C4422 x9.A1 a_2879_n62# 1.54e-20
C4423 x2.X a_3333_601# 0.119f
C4424 x6.X a_473_993# 9.17e-20
C4425 a_12607_601# a_12447_n62# 0.0026f
C4426 a_12433_993# a_12134_n88# 8.71e-20
C4427 a_4860_1467# check[4] 0.318f
C4428 a_3420_212# a_3839_220# 2.46e-19
C4429 a_3421_n88# a_3558_304# 0.00907f
C4430 a_2879_n62# a_4338_n62# 3.79e-20
C4431 a_10680_909# VDD_SW[3] 2.82e-20
C4432 D[1] a_16024_909# 8.04e-19
C4433 a_14379_627# VDD_SW_b[1] 1.15e-19
C4434 x9.A1 a_10597_n88# 8.52e-21
C4435 check[0] a_16037_1642# 0.00577f
C4436 x20.X a_14379_627# 2.67e-20
C4437 a_6920_627# a_7203_627# 0.0011f
C4438 reset a_29_2457# 0.201f
C4439 check[6] a_505_1289# 0.25f
C4440 check[2] a_10596_212# 3.16e-20
C4441 VDD a_3070_220# 0.0041f
C4442 VDD x3.A 0.166f
C4443 a_14428_1467# VSS_SW[1] 0.0274f
C4444 a_4811_627# a_5575_627# 0.00134f
C4445 D[5] a_6124_993# 2.53e-19
C4446 x2.X VDD_SW[5] 0.0327f
C4447 VDD a_557_993# 0.00438f
C4448 D[2] a_14096_627# 0.00238f
C4449 VDD_SW_b[4] a_9646_90# 0.00345f
C4450 a_27_627# a_473_993# 0.159f
C4451 D[7] a_647_601# 0.00584f
C4452 x2.X a_13906_n62# 1.9e-19
C4453 check[3] a_7254_90# 2.5e-20
C4454 x2.X a_4064_909# 4.04e-19
C4455 x2.X a_12153_627# 0.0537f
C4456 x14.X a_11071_1642# 1.97e-20
C4457 a_3893_122# VSS_SW[5] 6.63e-20
C4458 VSS_SW_b[6] a_3761_n62# 5.35e-19
C4459 x2.X a_7711_1642# 2.63e-19
C4460 VDD a_14428_1467# 0.114f
C4461 a_2865_993# VSS_SW[6] 0.00296f
C4462 VDD a_4977_627# 0.659f
C4463 x6.X a_1503_1642# 1.98e-20
C4464 x20.X a_15072_106# 1.89e-20
C4465 VDD_SW_b[1] a_15072_106# 5.22e-19
C4466 x9.A1 D[7] 0.268f
C4467 VDD VSS_SW[5] 0.56f
C4468 a_16109_1642# check[0] 0.318f
C4469 a_10734_304# VSS_SW[2] 2.76e-20
C4470 x9.A1 a_6529_n62# 5.7e-21
C4471 D[3] a_10246_220# 1.98e-20
C4472 a_5271_n62# a_7350_n88# 3.08e-21
C4473 a_6539_1642# a_6199_895# 0.00226f
C4474 a_1029_n88# a_1745_304# 0.0018f
C4475 a_487_n62# a_593_n62# 0.0526f
C4476 x2.X a_15767_895# 0.148f
C4477 a_1233_n88# a_1447_220# 0.0104f
C4478 a_1028_212# a_1946_n62# 0.0453f
C4479 a_27_627# a_1159_627# 0.00272f
C4480 check[4] a_6285_1642# 0.256f
C4481 x8.X VDD_SW[7] 0.305f
C4482 a_9742_n88# a_10597_n88# 0.0477f
C4483 a_13103_n62# a_13329_n62# 3.34e-19
C4484 VDD a_9312_627# 0.194f
C4485 a_12036_1467# a_12134_n88# 6.87e-20
C4486 a_11987_627# VSS_SW[1] 4.95e-21
C4487 check[5] check[4] 0.00523f
C4488 a_9644_1467# VSS_SW_b[3] 2.13e-19
C4489 a_505_1289# D[7] 0.0661f
C4490 x9.A1 a_2419_627# 8.07e-19
C4491 check[0] VDD_SW[1] 0.00392f
C4492 VDD a_5575_627# 1.8e-19
C4493 a_10983_895# a_12341_627# 8.26e-21
C4494 D[6] a_4137_304# 8.38e-19
C4495 x13.X a_10509_601# 4.31e-21
C4496 VDD a_12924_n62# 7.87e-19
C4497 a_9786_1642# VSS_SW[3] 0.00105f
C4498 x9.A1 a_4077_1642# 5.26e-19
C4499 a_6529_304# VSS_SW[4] 6.59e-21
C4500 a_5377_n62# a_5748_n62# 4.19e-20
C4501 a_6017_n88# VSS_SW_b[4] 4.54e-20
C4502 a_6539_1642# VDD_SW_b[5] 2.59e-19
C4503 x10.X a_3807_895# 0.00864f
C4504 VDD a_11987_627# 0.393f
C4505 VDD VDD_SW_b[3] 0.156f
C4506 x9.A1 a_535_1642# 5.26e-19
C4507 VDD_SW_b[2] a_13705_n62# 5.22e-19
C4508 a_1415_895# a_1555_627# 0.0383f
C4509 a_473_993# VDD_SW[7] 4.17e-21
C4510 a_941_601# a_1363_627# 1.96e-20
C4511 VDD a_4370_1315# 3.89e-19
C4512 x2.X a_5748_n62# 3.68e-20
C4513 check[0] D[2] 5.94e-20
C4514 a_647_601# a_1112_909# 9.46e-19
C4515 x2.X a_9644_1467# 2.88e-19
C4516 a_7967_627# a_8539_627# 2.46e-21
C4517 check[2] x15.X 0.00965f
C4518 a_3807_895# D[5] 2.17e-19
C4519 a_3648_993# a_4811_627# 7.46e-20
C4520 a_3420_212# a_5271_n62# 2.62e-19
C4521 a_3421_n88# a_4958_n88# 1.98e-19
C4522 VDD_SW_b[5] a_8288_909# 2.96e-21
C4523 VDD a_13929_1642# 0.00177f
C4524 a_2585_627# a_2566_n88# 4.91e-19
C4525 VDD_SW_b[7] a_1745_n62# 5.22e-19
C4526 x2.X a_678_220# 0.00279f
C4527 a_14545_627# a_14733_627# 0.189f
C4528 x10.X VDD_SW_b[6] 7.23e-19
C4529 x9.X a_4528_627# 0.0337f
C4530 a_14857_1289# a_14999_601# 8.76e-20
C4531 a_14999_601# a_15608_993# 0.00189f
C4532 a_7252_1467# VDD_SW[5] 0.00487f
C4533 VDD_SW_b[3] a_10596_212# 0.0417f
C4534 a_7394_1315# D[4] 7.54e-19
C4535 a_14839_n62# a_15030_220# 3.3e-19
C4536 check[4] x12.X 5.98e-19
C4537 a_7394_1315# VSS_SW[4] 7.95e-19
C4538 a_9761_627# VSS_SW_b[3] 5.23e-20
C4539 x13.X a_7203_627# 2.67e-20
C4540 VSS_SW[1] a_15853_122# 2.79e-21
C4541 a_9595_627# a_10597_n88# 1.06e-19
C4542 x9.A1 a_5257_993# 1.48e-19
C4543 x9.A1 a_4149_1642# 0.195f
C4544 a_939_2457# check[6] 0.0505f
C4545 check[3] a_8205_n88# 2.49e-20
C4546 VDD_SW_b[6] D[5] 1.57e-19
C4547 VDD_SW_b[2] a_12680_106# 5.23e-19
C4548 a_3356_n62# a_3761_n62# 2.46e-21
C4549 a_7252_1467# a_7711_1642# 6.64e-19
C4550 a_4689_2457# a_4528_627# 4.35e-21
C4551 x7.X a_1028_212# 0.245f
C4552 check[6] a_1233_n88# 2.51e-19
C4553 check[3] D[5] 6.36e-20
C4554 x2.X a_10359_627# 0.0391f
C4555 a_3648_993# a_3893_122# 1.51e-20
C4556 a_3183_627# a_2566_n88# 1.08e-19
C4557 x2.X VSS_SW[6] 0.184f
C4558 VDD a_15853_122# 0.313f
C4559 check[4] a_6285_122# 6.49e-20
C4560 x2.X a_9761_627# 0.0537f
C4561 VDD a_76_1467# 0.117f
C4562 a_5812_212# a_6529_n62# 0.00206f
C4563 check[0] VSS_SW_b[1] 3.18e-20
C4564 check[5] a_3761_n62# 9.81e-20
C4565 a_1029_n88# a_3112_106# 1.67e-21
C4566 a_305_2457# a_647_601# 1.12e-19
C4567 a_1501_122# a_2566_n88# 8e-21
C4568 x3.X a_193_627# 5.4e-19
C4569 a_1028_212# a_3420_212# 1.9e-21
C4570 VDD a_3648_993# 0.189f
C4571 a_27_627# a_2585_627# 1.15e-20
C4572 a_5431_601# a_5165_627# 8.07e-20
C4573 check[1] a_13515_627# 3.88e-19
C4574 a_4977_627# a_5341_993# 0.0018f
C4575 a_5725_601# a_6199_895# 0.265f
C4576 x2.X a_14379_627# 0.354f
C4577 a_10055_n62# a_10288_106# 0.124f
C4578 ready x6.X 2.32e-20
C4579 x2.X VDD_SW_b[2] 7.31e-19
C4580 x2.X a_13461_1642# 0.00643f
C4581 VDD a_174_n88# 0.693f
C4582 a_8677_122# VSS_SW_b[3] 1.02e-20
C4583 x30.A a_4811_627# 2.63e-21
C4584 a_12989_n88# a_14526_n88# 1.98e-19
C4585 a_12988_212# a_14839_n62# 2.62e-19
C4586 a_305_2457# x9.A1 0.00214f
C4587 D[6] a_5504_106# 1.39e-21
C4588 VDD_SW_b[3] a_11313_n62# 5.22e-19
C4589 VDD_SW[5] a_8591_895# 1.27e-20
C4590 x9.A1 a_11313_304# 8.15e-21
C4591 a_14545_627# a_16488_627# 1.79e-20
C4592 D[4] a_7896_106# 8.74e-19
C4593 a_7203_627# a_8204_212# 6.99e-20
C4594 VSS_SW[4] a_7896_106# 4.63e-19
C4595 x9.A1 a_5289_1289# 0.105f
C4596 a_7254_90# VSS_SW_b[4] 0.19f
C4597 a_1757_1642# x8.X 7.97e-19
C4598 a_5165_627# a_5365_627# 3.81e-19
C4599 a_6199_895# a_6456_909# 0.00869f
C4600 a_4811_627# a_7203_627# 1.63e-20
C4601 a_5725_601# VDD_SW_b[5] 0.00636f
C4602 a_6040_993# a_5943_627# 0.00386f
C4603 a_939_2457# D[7] 0.0344f
C4604 ready a_27_627# 1.42e-21
C4605 x2.X a_8677_122# 0.0043f
C4606 x8.X a_2773_627# 6.12e-19
C4607 VDD a_10509_601# 0.46f
C4608 check[1] VSS_SW[1] 1.4e-19
C4609 check[3] a_8117_601# 2.11e-19
C4610 a_305_2457# a_505_1289# 0.00165f
C4611 x2.X a_15072_106# 0.0385f
C4612 a_9644_1467# x14.X 0.0877f
C4613 D[7] a_1233_n88# 0.00546f
C4614 a_12341_627# a_12517_993# 8.99e-19
C4615 a_12901_601# a_13300_993# 9.41e-19
C4616 a_12153_627# a_13119_627# 2.14e-20
C4617 a_12433_993# a_12751_627# 0.025f
C4618 x9.A1 a_4958_n88# 7.41e-19
C4619 a_4338_n62# a_4958_n88# 8.26e-21
C4620 x16.X VDD_SW[3] 0.307f
C4621 a_3893_122# a_4137_n62# 0.00807f
C4622 x15.X a_11987_627# 0.00297f
C4623 VDD a_2897_1289# 0.191f
C4624 x15.X VDD_SW_b[3] 0.24f
C4625 a_10007_1315# D[3] 0.00202f
C4626 VDD a_15316_n62# 7.87e-19
C4627 a_2419_627# a_3732_993# 2.13e-19
C4628 D[6] a_3504_909# 8.51e-19
C4629 a_939_2457# a_2419_627# 2.48e-19
C4630 VDD check[1] 1.64f
C4631 a_2136_627# a_3333_601# 1.84e-20
C4632 VDD_SW[7] a_2585_627# 9.25e-19
C4633 a_6456_909# VDD_SW_b[5] 3.4e-20
C4634 a_14379_627# a_14825_993# 0.159f
C4635 D[1] a_14999_601# 0.00585f
C4636 VDD x30.A 0.705f
C4637 VSS_SW_b[3] a_10532_n62# 1.68e-19
C4638 VDD_SW_b[2] a_14825_993# 8.2e-21
C4639 a_10801_n88# a_10937_n62# 0.0697f
C4640 a_10597_n88# VSS_SW[2] 9.22e-19
C4641 x9.X a_2879_n62# 0.00192f
C4642 a_10509_601# a_10596_212# 6.03e-19
C4643 a_10824_993# a_10055_n62# 3.59e-19
C4644 x2.X x18.X 3.6e-19
C4645 D[3] a_10288_106# 8.76e-19
C4646 a_4977_627# a_6017_n88# 8.75e-19
C4647 a_5431_601# a_5813_n88# 0.00322f
C4648 a_6199_895# a_5271_n62# 0.00219f
C4649 a_5725_601# a_5504_106# 3.46e-19
C4650 a_8679_1642# a_8677_122# 1.57e-21
C4651 VSS_SW[5] a_6017_n88# 9.93e-21
C4652 a_941_601# a_174_n88# 0.00259f
C4653 a_473_993# a_487_n62# 2.63e-19
C4654 a_13906_n62# a_14526_n88# 8.26e-21
C4655 a_13461_122# a_13705_n62# 0.00807f
C4656 a_193_627# a_1028_212# 1.02e-19
C4657 a_647_601# a_720_106# 1.01e-19
C4658 x7.X a_1946_n62# 0.0016f
C4659 x9.A1 a_11704_627# 2e-20
C4660 VDD a_7203_627# 0.393f
C4661 VDD_SW[3] a_12153_627# 9.25e-19
C4662 a_11704_627# a_12901_601# 1.71e-20
C4663 VDD a_6153_n62# 0.0301f
C4664 a_15855_1642# x20.X 1.31e-19
C4665 a_7203_627# a_7649_993# 0.159f
C4666 D[4] a_7823_601# 0.00584f
C4667 x2.X a_10532_n62# 3.68e-20
C4668 a_7823_601# VSS_SW[4] 6.25e-19
C4669 ready VDD_SW[7] 0.0363f
C4670 x14.X a_9761_627# 0.00312f
C4671 x2.X check[4] 0.148f
C4672 VSS_SW_b[1] a_15721_n62# 5.35e-19
C4673 a_1946_n62# a_3420_212# 5.58e-22
C4674 a_15853_122# a_16097_n62# 0.00807f
C4675 x2.X a_8432_993# 0.187f
C4676 a_14999_601# a_15380_212# 4.51e-19
C4677 a_14825_993# a_15072_106# 4.96e-20
C4678 a_15293_601# a_14839_n62# 3.74e-20
C4679 a_14545_627# a_15381_n88# 1.27e-19
C4680 VDD_SW_b[5] a_5271_n62# 5.28e-19
C4681 check[5] a_3807_895# 0.00272f
C4682 x2.X a_15799_220# 9.58e-19
C4683 a_13216_993# a_13323_627# 0.00707f
C4684 a_13375_895# VDD_SW[2] 0.00356f
C4685 VDD a_1166_304# 0.0164f
C4686 a_7681_1289# a_7663_n62# 3.44e-19
C4687 a_11071_1642# x16.X 1.52e-20
C4688 VDD_SW_b[6] a_3356_n62# 8.1e-20
C4689 x2.X a_10103_1642# 2.63e-19
C4690 a_7203_627# a_8335_627# 0.00272f
C4691 a_505_1289# a_720_106# 5.3e-21
C4692 a_7757_627# VSS_SW[4] 3.79e-19
C4693 D[4] a_8623_220# 7.11e-19
C4694 a_12447_n62# VSS_SW_b[2] 0.0142f
C4695 VSS_SW[2] a_12638_220# 4.26e-19
C4696 a_12988_212# a_13193_n88# 0.15f
C4697 a_8409_n88# a_8677_122# 0.206f
C4698 VSS_SW[4] a_8623_220# 6.42e-21
C4699 a_8205_n88# VSS_SW_b[4] 7.59e-19
C4700 a_9644_1467# a_9646_90# 1e-19
C4701 a_13715_1642# a_13936_1315# 0.00783f
C4702 a_11069_122# VSS_SW_b[2] 1.16e-20
C4703 VDD_SW[2] a_15243_909# 2.16e-20
C4704 a_5896_909# VDD_SW[5] 2.82e-20
C4705 x18.X a_14825_993# 9.17e-20
C4706 x2.X a_7769_n62# 5.57e-20
C4707 D[5] VSS_SW_b[4] 2.02e-19
C4708 a_2610_1315# D[6] 7.54e-19
C4709 a_10509_601# a_9949_627# 1.24e-20
C4710 a_10983_895# a_10824_993# 0.207f
C4711 a_9761_627# a_10680_909# 0.00907f
C4712 check[5] VDD_SW_b[6] 0.00217f
C4713 D[3] a_10824_993# 0.00609f
C4714 a_10149_627# VSS_SW[3] 3.79e-19
C4715 a_6285_1642# check[3] 9.11e-21
C4716 x9.X a_2419_627# 2.64e-20
C4717 a_8679_1642# a_8432_993# 0.00176f
C4718 VDD_SW_b[6] a_5675_909# 2.62e-21
C4719 VDD a_10246_220# 0.0041f
C4720 a_5271_n62# a_5504_106# 0.124f
C4721 a_4958_n88# a_5812_212# 0.0319f
C4722 a_8591_895# a_9761_627# 2.64e-19
C4723 a_8117_601# a_10215_601# 1.75e-20
C4724 D[2] a_12851_909# 6.77e-19
C4725 a_11987_627# a_13072_909# 1.09e-19
C4726 VDD_SW_b[3] a_13072_909# 2.96e-21
C4727 VDD_SW_b[1] a_16488_627# 0.186f
C4728 x2.X a_13461_122# 0.0043f
C4729 x20.X a_16488_627# 0.0338f
C4730 D[6] VDD_SW[6] 0.246f
C4731 x15.X a_10509_601# 1.29e-19
C4732 a_29_2457# x2.X 3.13e-19
C4733 x2.X a_1555_627# 0.0151f
C4734 a_305_2457# a_939_2457# 8.52e-20
C4735 a_15495_n62# a_15721_n62# 3.34e-19
C4736 x2.X a_381_627# 0.00139f
C4737 VDD a_12341_627# 0.109f
C4738 a_14428_1467# VDD_SW[2] 0.00484f
C4739 VDD a_6760_1315# 3.75e-19
C4740 a_12399_1315# D[2] 0.00202f
C4741 a_10055_n62# a_10734_304# 0.00652f
C4742 a_10288_106# a_10545_304# 0.00857f
C4743 x17.X a_13375_895# 0.00662f
C4744 VDD_SW_b[4] a_9761_627# 0.00344f
C4745 x7.X a_3420_212# 1.68e-21
C4746 x15.X check[1] 5.58e-19
C4747 a_7681_1289# a_7369_627# 0.00323f
C4748 a_9122_n62# a_8921_n62# 3.81e-19
C4749 x11.X D[4] 2.11e-19
C4750 a_7203_627# a_9949_627# 4.74e-21
C4751 x9.A1 a_3947_627# 5.22e-20
C4752 x11.X VSS_SW[4] 0.149f
C4753 a_12988_212# a_14430_90# 0.00101f
C4754 a_13193_n88# a_13705_304# 6.69e-20
C4755 a_12989_n88# a_13906_n62# 0.189f
C4756 VSS_SW_b[2] a_13126_304# 3.87e-20
C4757 VDD a_15692_993# 0.00281f
C4758 x9.A1 a_12447_n62# 1.55e-20
C4759 VDD a_16323_1642# 0.00177f
C4760 a_12901_601# a_12447_n62# 3.74e-20
C4761 a_12433_993# a_12680_106# 4.96e-20
C4762 a_12607_601# a_12988_212# 4.51e-19
C4763 a_12153_627# a_12989_n88# 1.27e-19
C4764 a_8591_895# a_8677_122# 4.53e-22
C4765 a_8432_993# a_8409_n88# 1.86e-19
C4766 a_7663_n62# a_7854_220# 3.24e-19
C4767 a_7252_1467# check[4] 1.57e-19
C4768 a_3039_601# a_3648_993# 0.00189f
C4769 x9.A1 a_1745_304# 6.9e-21
C4770 a_2585_627# a_2773_627# 0.189f
C4771 x9.A1 a_11069_122# 3.99e-20
C4772 a_4149_1642# x9.X 0.0841f
C4773 a_2566_n88# a_3893_122# 4.59e-22
C4774 a_2879_n62# a_3625_n88# 0.199f
C4775 a_3112_106# a_3421_n88# 0.0327f
C4776 check[2] a_10801_n88# 2.51e-19
C4777 a_9761_627# VDD_SW[3] 1.96e-20
C4778 a_9595_627# a_11704_627# 1.75e-19
C4779 x12.X check[3] 0.00903f
C4780 a_2136_627# VSS_SW[6] 0.00164f
C4781 x10.X a_5223_1315# 2.41e-19
C4782 x14.X a_8432_993# 2.78e-19
C4783 a_14379_627# a_14526_n88# 0.00176f
C4784 VDD a_2566_n88# 0.69f
C4785 a_14096_627# VSS_SW[1] 0.00166f
C4786 VDD_SW_b[2] a_14526_n88# 5.91e-19
C4787 x2.X a_6124_993# 4.68e-19
C4788 VDD_SW[6] a_5725_601# 2.46e-20
C4789 D[2] a_13323_627# 2e-19
C4790 a_11987_627# VDD_SW[2] 3.29e-20
C4791 x16.X a_12153_627# 0.00313f
C4792 a_5323_2457# x9.A1 1.72f
C4793 a_5223_1315# D[5] 0.00202f
C4794 VDD_SW_b[4] a_8677_122# 0.00445f
C4795 D[4] a_10055_n62# 1.56e-21
C4796 x2.X a_12433_993# 0.15f
C4797 a_7896_106# a_8545_n62# 0.00316f
C4798 a_7663_n62# VSS_SW[3] 1.64e-20
C4799 a_8204_212# a_8319_n62# 0.00272f
C4800 a_2865_993# VDD_SW_b[6] 4.91e-21
C4801 a_3333_601# a_4064_909# 0.0016f
C4802 VDD x6.X 0.396f
C4803 a_76_1467# VSS_SW_b[7] 2.13e-19
C4804 check[6] x8.X 5.86e-19
C4805 VDD a_14096_627# 0.194f
C4806 x20.X a_15381_n88# 0.0189f
C4807 VDD_SW_b[1] a_15381_n88# 0.0406f
C4808 a_11313_304# VSS_SW[2] 6.58e-21
C4809 a_14428_1467# x17.X 4.9e-19
C4810 a_10215_601# a_10125_993# 6.69e-20
C4811 a_13929_1642# VDD_SW[2] 5.15e-19
C4812 D[3] a_10734_304# 9.69e-19
C4813 x2.X a_15855_1642# 0.00645f
C4814 x2.X a_14733_627# 0.00139f
C4815 a_5813_n88# a_5462_220# 4.48e-20
C4816 a_1978_1315# VDD_SW_b[7] 2.64e-20
C4817 a_14526_n88# a_15072_106# 0.207f
C4818 a_5504_106# a_5950_304# 0.00412f
C4819 a_5812_212# a_5761_304# 2.13e-19
C4820 a_2897_1289# a_3039_601# 8.76e-20
C4821 a_5271_n62# a_6231_220# 1.21e-20
C4822 check[4] a_5319_1642# 0.00526f
C4823 a_9742_n88# a_11069_122# 4.59e-22
C4824 a_174_n88# VSS_SW_b[7] 0.135f
C4825 a_720_106# a_1233_n88# 0.00189f
C4826 VSS_SW[7] a_678_220# 4.25e-19
C4827 a_1028_212# a_1029_n88# 0.784f
C4828 a_487_n62# a_1501_122# 0.0633f
C4829 a_5323_2457# a_6040_993# 2.04e-19
C4830 VDD a_27_627# 0.408f
C4831 VDD a_7733_993# 0.0042f
C4832 a_8204_212# a_10288_106# 5.86e-20
C4833 x7.X a_193_627# 1.13e-20
C4834 a_8117_601# a_7557_627# 1.15e-20
C4835 a_7823_601# a_8067_909# 0.0104f
C4836 a_7369_627# a_8288_909# 0.00907f
C4837 a_7649_993# a_7733_993# 0.00972f
C4838 a_8591_895# a_8432_993# 0.207f
C4839 check[6] a_473_993# 7.17e-20
C4840 x9.A1 a_7681_1289# 0.105f
C4841 x10.X a_4977_627# 0.00315f
C4842 D[6] a_3421_n88# 0.158f
C4843 a_2419_627# a_3625_n88# 0.00204f
C4844 VDD a_13329_n62# 0.0301f
C4845 x9.X a_4958_n88# 0.00863f
C4846 x10.X VSS_SW[5] 0.251f
C4847 D[1] a_15030_220# 2.03e-20
C4848 check[0] VSS_SW[1] 0.0493f
C4849 a_5813_n88# VSS_SW[4] 9.23e-19
C4850 a_6017_n88# a_6153_n62# 0.0697f
C4851 VSS_SW_b[5] a_5748_n62# 1.68e-19
C4852 x9.A1 a_14999_601# 2.81e-20
C4853 a_13375_895# a_14545_627# 2.96e-19
C4854 a_12901_601# a_14999_601# 1.52e-20
C4855 a_4811_627# a_5431_601# 0.149f
C4856 x2.X a_12036_1467# 2.86e-19
C4857 x17.X a_11987_627# 2.67e-20
C4858 D[5] a_4977_627# 0.168f
C4859 D[5] VSS_SW[5] 0.134f
C4860 VDD a_8319_n62# 0.00521f
C4861 a_8432_993# VDD_SW_b[4] 5.63e-20
C4862 D[4] D[3] 0.00183f
C4863 x13.X a_9154_1315# 0.00146f
C4864 a_7369_627# VSS_SW[3] 4.78e-21
C4865 a_8731_627# a_8204_212# 7.07e-21
C4866 a_12447_n62# a_12553_n62# 0.0526f
C4867 x8.X D[7] 9.68e-19
C4868 VDD a_218_1642# 0.00226f
C4869 x2.X a_3807_895# 0.148f
C4870 a_2585_627# a_4528_627# 2e-20
C4871 x6.X a_941_601# 4.9e-20
C4872 VDD check[0] 1.64f
C4873 a_2879_n62# a_4862_90# 6.12e-21
C4874 a_3420_212# a_4137_304# 4.45e-20
C4875 a_3625_n88# a_3558_304# 9.46e-19
C4876 VSS_SW_b[6] a_3070_220# 5.34e-20
C4877 a_3421_n88# a_3839_220# 0.00276f
C4878 a_11987_627# a_12134_n88# 0.00176f
C4879 a_2566_n88# a_2985_n62# 0.0383f
C4880 a_4413_2457# a_3807_895# 7.82e-20
C4881 VDD_SW_b[1] a_16298_n62# 0.0143f
C4882 x20.X a_16298_n62# 0.00153f
C4883 VDD_SW_b[3] a_12134_n88# 5.9e-19
C4884 a_11704_627# VSS_SW[2] 0.00163f
C4885 a_12038_90# VSS_SW_b[2] 0.191f
C4886 a_6339_627# a_7203_627# 1.09e-19
C4887 a_6920_627# D[4] 4.42e-19
C4888 reset x3.A 0.00421f
C4889 VDD_SW_b[5] a_7350_n88# 5.9e-19
C4890 check[6] a_1503_1642# 0.257f
C4891 a_14825_993# a_14733_627# 0.0369f
C4892 a_14999_601# a_14909_993# 6.69e-20
C4893 a_6920_627# VSS_SW[4] 0.00164f
C4894 a_15293_601# a_15608_993# 0.13f
C4895 a_14545_627# a_15243_909# 0.00276f
C4896 VDD_SW_b[3] a_10801_n88# 0.00132f
C4897 a_8933_1315# D[4] 0.00195f
C4898 x2.X a_16488_627# 3.63e-19
C4899 VDD a_3369_304# 0.00265f
C4900 a_15072_106# a_15329_304# 0.00857f
C4901 a_14839_n62# a_15518_304# 0.00652f
C4902 a_4811_627# a_5365_627# 0.00206f
C4903 x10.X a_4370_1315# 3.75e-20
C4904 VDD VDD_SW[7] 0.388f
C4905 x9.A1 a_6539_1642# 0.195f
C4906 x8.X a_2419_627# 0.236f
C4907 VDD a_891_909# 0.00999f
C4908 VDD a_10288_106# 0.356f
C4909 VDD_SW_b[4] a_7769_n62# 4.77e-19
C4910 a_27_627# a_941_601# 0.14f
C4911 D[7] a_473_993# 0.00884f
C4912 VDD_SW_b[2] a_12989_n88# 0.0406f
C4913 a_8933_1642# a_8861_1642# 6.64e-19
C4914 a_8342_304# VSS_SW[3] 2.77e-20
C4915 a_3283_909# VDD_SW[6] 1.01e-20
C4916 x2.X VDD_SW_b[6] 7.36e-19
C4917 a_4413_2457# VDD_SW_b[6] 7.33e-20
C4918 x2.X a_10727_627# 0.00706f
C4919 x16.X a_9761_627# 6.37e-20
C4920 x2.X check[3] 0.149f
C4921 x2.X a_2831_1315# 3.19e-19
C4922 VDD a_5431_601# 0.313f
C4923 a_3333_601# VSS_SW[6] 2.13e-19
C4924 a_5725_601# a_7369_627# 6.25e-20
C4925 a_5504_106# a_7350_n88# 1.86e-21
C4926 check[1] VDD_SW[2] 0.00389f
C4927 a_1233_n88# a_1745_304# 6.69e-20
C4928 a_1029_n88# a_1946_n62# 0.189f
C4929 VSS_SW_b[7] a_1166_304# 3.58e-20
C4930 a_487_n62# a_964_n62# 1.96e-20
C4931 a_720_106# a_593_n62# 0.0256f
C4932 a_1028_212# a_2470_90# 0.00101f
C4933 x16.X a_13461_1642# 2.02e-20
C4934 a_10055_n62# a_10597_n88# 0.125f
C4935 a_10288_106# a_10596_212# 0.14f
C4936 D[7] a_1159_627# 6.12e-19
C4937 x2.X a_12495_1642# 2.63e-19
C4938 VDD a_8731_627# 6.99e-19
C4939 a_12988_212# a_15380_212# 1.9e-21
C4940 a_12989_n88# a_15072_106# 1.67e-21
C4941 a_13461_122# a_14526_n88# 8e-21
C4942 a_7369_627# VDD_SW[4] 1.85e-20
C4943 a_6753_1642# VDD_SW[5] 5.3e-19
C4944 a_8117_601# a_9312_627# 5.84e-19
C4945 x27.A VDD_SW[6] 0.0227f
C4946 D[2] a_12638_220# 2.03e-20
C4947 a_2468_1467# a_2566_n88# 6.87e-20
C4948 a_1503_1642# D[7] 0.0682f
C4949 x9.A1 D[6] 0.268f
C4950 D[6] a_4338_n62# 0.158f
C4951 x9.A1 a_5002_1642# 8.62e-19
C4952 a_9761_627# a_12153_627# 2.94e-19
C4953 x9.A1 VSS_SW[3] 0.113f
C4954 a_7203_627# a_7254_90# 6.13e-19
C4955 check[3] a_8679_1642# 0.257f
C4956 a_6285_122# VSS_SW_b[4] 1.09e-20
C4957 a_6730_n62# VSS_SW[4] 6.09e-20
C4958 x10.X a_3648_993# 2.81e-19
C4959 x9.A1 a_1685_1642# 5.26e-19
C4960 a_1256_993# a_1555_627# 0.0256f
C4961 a_941_601# VDD_SW[7] 1.75e-19
C4962 VDD a_10824_993# 0.189f
C4963 a_941_601# a_891_909# 1.21e-20
C4964 a_193_627# a_791_627# 6.04e-20
C4965 a_4860_1467# VSS_SW[5] 0.0274f
C4966 VDD_SW_b[2] a_13906_n62# 0.0144f
C4967 a_11987_627# a_14545_627# 1.2e-20
C4968 a_12153_627# a_14379_627# 1.58e-20
C4969 x2.X a_15381_n88# 0.0206f
C4970 a_13216_993# a_13300_993# 0.00857f
C4971 a_12465_1289# a_12607_601# 8.76e-20
C4972 a_12153_627# VDD_SW_b[2] 0.0022f
C4973 a_16097_n62# VSS 0.00183f
C4974 a_15721_n62# VSS 0.176f
C4975 a_15495_n62# VSS 0.0109f
C4976 a_15316_n62# VSS 0.00193f
C4977 a_14945_n62# VSS 0.166f
C4978 a_16298_n62# VSS 0.1f
C4979 a_16097_304# VSS 1.79e-19
C4980 a_15799_220# VSS 1.48e-19
C4981 a_15518_304# VSS 6.03e-19
C4982 a_15329_304# VSS 1.17e-21
C4983 a_13705_n62# VSS 0.0017f
C4984 VSS_SW_b[1] VSS 0.32f
C4985 a_15853_122# VSS 0.263f
C4986 a_15585_n88# VSS 0.287f
C4987 a_15381_n88# VSS 0.329f
C4988 a_15380_212# VSS 0.777f
C4989 a_15072_106# VSS 0.245f
C4990 a_14839_n62# VSS 0.367f
C4991 a_14526_n88# VSS 0.454f
C4992 VSS_SW[1] VSS 0.669f
C4993 a_13329_n62# VSS 0.176f
C4994 a_13103_n62# VSS 0.0108f
C4995 a_12924_n62# VSS 0.00192f
C4996 a_12553_n62# VSS 0.166f
C4997 a_14430_90# VSS 0.224f
C4998 a_13906_n62# VSS 0.0993f
C4999 a_13126_304# VSS 3.84e-19
C5000 a_11313_n62# VSS 0.0017f
C5001 VSS_SW_b[2] VSS 0.319f
C5002 a_13461_122# VSS 0.262f
C5003 a_13193_n88# VSS 0.286f
C5004 a_12989_n88# VSS 0.321f
C5005 a_12988_212# VSS 0.713f
C5006 a_12680_106# VSS 0.245f
C5007 a_12447_n62# VSS 0.367f
C5008 a_12134_n88# VSS 0.454f
C5009 VSS_SW[2] VSS 0.669f
C5010 a_10937_n62# VSS 0.176f
C5011 a_10711_n62# VSS 0.0108f
C5012 a_10532_n62# VSS 0.00192f
C5013 a_10161_n62# VSS 0.166f
C5014 a_12038_90# VSS 0.224f
C5015 a_11514_n62# VSS 0.0993f
C5016 a_10734_304# VSS 3.84e-19
C5017 a_8921_n62# VSS 0.0017f
C5018 VSS_SW_b[3] VSS 0.319f
C5019 a_11069_122# VSS 0.262f
C5020 a_10801_n88# VSS 0.286f
C5021 a_10597_n88# VSS 0.321f
C5022 a_10596_212# VSS 0.713f
C5023 a_10288_106# VSS 0.245f
C5024 a_10055_n62# VSS 0.367f
C5025 a_9742_n88# VSS 0.454f
C5026 VSS_SW[3] VSS 0.669f
C5027 a_8545_n62# VSS 0.176f
C5028 a_8319_n62# VSS 0.0108f
C5029 a_8140_n62# VSS 0.00192f
C5030 a_7769_n62# VSS 0.166f
C5031 a_9646_90# VSS 0.224f
C5032 a_9122_n62# VSS 0.0993f
C5033 a_8342_304# VSS 3.84e-19
C5034 a_6529_n62# VSS 0.0017f
C5035 VSS_SW_b[4] VSS 0.319f
C5036 a_8677_122# VSS 0.262f
C5037 a_8409_n88# VSS 0.286f
C5038 a_8205_n88# VSS 0.321f
C5039 a_8204_212# VSS 0.713f
C5040 a_7896_106# VSS 0.245f
C5041 a_7663_n62# VSS 0.367f
C5042 a_7350_n88# VSS 0.454f
C5043 VSS_SW[4] VSS 0.585f
C5044 a_6153_n62# VSS 0.176f
C5045 a_5927_n62# VSS 0.0108f
C5046 a_5748_n62# VSS 0.00192f
C5047 a_5377_n62# VSS 0.166f
C5048 a_7254_90# VSS 0.224f
C5049 a_6730_n62# VSS 0.0993f
C5050 a_5950_304# VSS 3.84e-19
C5051 a_4137_n62# VSS 0.0017f
C5052 VSS_SW_b[5] VSS 0.319f
C5053 a_6285_122# VSS 0.262f
C5054 a_6017_n88# VSS 0.286f
C5055 a_5813_n88# VSS 0.321f
C5056 a_5812_212# VSS 0.713f
C5057 a_5504_106# VSS 0.245f
C5058 a_5271_n62# VSS 0.367f
C5059 a_4958_n88# VSS 0.454f
C5060 VSS_SW[5] VSS 0.598f
C5061 a_3761_n62# VSS 0.176f
C5062 a_3535_n62# VSS 0.0108f
C5063 a_3356_n62# VSS 0.00192f
C5064 a_2985_n62# VSS 0.166f
C5065 a_4862_90# VSS 0.224f
C5066 a_4338_n62# VSS 0.0993f
C5067 a_3558_304# VSS 3.84e-19
C5068 a_1745_n62# VSS 0.0017f
C5069 VSS_SW_b[6] VSS 0.32f
C5070 a_3893_122# VSS 0.262f
C5071 a_3625_n88# VSS 0.286f
C5072 a_3421_n88# VSS 0.321f
C5073 a_3420_212# VSS 0.713f
C5074 a_3112_106# VSS 0.245f
C5075 a_2879_n62# VSS 0.367f
C5076 a_2566_n88# VSS 0.454f
C5077 VSS_SW[6] VSS 0.593f
C5078 a_1369_n62# VSS 0.176f
C5079 a_1143_n62# VSS 0.0108f
C5080 a_964_n62# VSS 0.00192f
C5081 a_593_n62# VSS 0.166f
C5082 a_2470_90# VSS 0.224f
C5083 a_1946_n62# VSS 0.0993f
C5084 a_1166_304# VSS 3.84e-19
C5085 VSS_SW_b[7] VSS 0.378f
C5086 a_1501_122# VSS 0.262f
C5087 a_1233_n88# VSS 0.286f
C5088 a_1029_n88# VSS 0.321f
C5089 a_1028_212# VSS 0.713f
C5090 a_720_106# VSS 0.245f
C5091 a_487_n62# VSS 0.367f
C5092 a_174_n88# VSS 0.462f
C5093 VSS_SW[7] VSS 0.917f
C5094 a_78_90# VSS 0.244f
C5095 VDD_SW[1] VSS 0.903f
C5096 a_15715_627# VSS 0.00197f
C5097 a_15907_627# VSS 0.166f
C5098 a_16488_627# VSS 0.248f
C5099 VDD_SW_b[1] VSS 0.413f
C5100 a_16024_909# VSS 4.78e-20
C5101 a_15511_627# VSS 0.0109f
C5102 a_14933_627# VSS 0.0017f
C5103 a_15143_627# VSS 0.176f
C5104 a_15692_993# VSS 2.15e-20
C5105 a_15464_909# VSS 4.47e-19
C5106 a_14733_627# VSS 0.0996f
C5107 a_15608_993# VSS 0.24f
C5108 a_15767_895# VSS 0.451f
C5109 a_15293_601# VSS 0.361f
C5110 a_14825_993# VSS 0.258f
C5111 a_14999_601# VSS 0.277f
C5112 a_14545_627# VSS 0.311f
C5113 D[1] VSS 1.65f
C5114 a_14379_627# VSS 0.702f
C5115 VDD_SW[2] VSS 0.454f
C5116 a_13323_627# VSS 0.00192f
C5117 a_13515_627# VSS 0.166f
C5118 a_14096_627# VSS 0.22f
C5119 VDD_SW_b[2] VSS 0.364f
C5120 a_13119_627# VSS 0.0108f
C5121 a_12541_627# VSS 0.0017f
C5122 a_12751_627# VSS 0.176f
C5123 a_13072_909# VSS 3.84e-19
C5124 a_12341_627# VSS 0.0996f
C5125 a_13216_993# VSS 0.239f
C5126 a_13375_895# VSS 0.438f
C5127 a_12901_601# VSS 0.358f
C5128 a_12433_993# VSS 0.258f
C5129 a_12607_601# VSS 0.277f
C5130 a_12153_627# VSS 0.31f
C5131 D[2] VSS 1.64f
C5132 a_11987_627# VSS 0.7f
C5133 VDD_SW[3] VSS 0.455f
C5134 a_10931_627# VSS 0.00192f
C5135 a_11123_627# VSS 0.166f
C5136 a_11704_627# VSS 0.22f
C5137 VDD_SW_b[3] VSS 0.364f
C5138 a_10727_627# VSS 0.0108f
C5139 a_10149_627# VSS 0.0017f
C5140 a_10359_627# VSS 0.176f
C5141 a_10680_909# VSS 3.84e-19
C5142 a_9949_627# VSS 0.0996f
C5143 a_10824_993# VSS 0.239f
C5144 a_10983_895# VSS 0.438f
C5145 a_10509_601# VSS 0.358f
C5146 a_10041_993# VSS 0.258f
C5147 a_10215_601# VSS 0.277f
C5148 a_9761_627# VSS 0.31f
C5149 D[3] VSS 1.64f
C5150 a_9595_627# VSS 0.7f
C5151 VDD_SW[4] VSS 0.454f
C5152 a_8539_627# VSS 0.00192f
C5153 a_8731_627# VSS 0.166f
C5154 a_9312_627# VSS 0.22f
C5155 VDD_SW_b[4] VSS 0.364f
C5156 a_8335_627# VSS 0.0108f
C5157 a_7757_627# VSS 0.0017f
C5158 a_7967_627# VSS 0.176f
C5159 a_8288_909# VSS 3.84e-19
C5160 a_7557_627# VSS 0.0996f
C5161 a_8432_993# VSS 0.239f
C5162 a_8591_895# VSS 0.438f
C5163 a_8117_601# VSS 0.358f
C5164 a_7649_993# VSS 0.258f
C5165 a_7823_601# VSS 0.277f
C5166 a_7369_627# VSS 0.31f
C5167 D[4] VSS 1.64f
C5168 a_7203_627# VSS 0.7f
C5169 VDD_SW[5] VSS 0.417f
C5170 a_6147_627# VSS 0.00192f
C5171 a_6339_627# VSS 0.166f
C5172 a_6920_627# VSS 0.22f
C5173 VDD_SW_b[5] VSS 0.364f
C5174 a_5943_627# VSS 0.0108f
C5175 a_5365_627# VSS 0.0017f
C5176 a_5575_627# VSS 0.176f
C5177 a_5896_909# VSS 3.84e-19
C5178 a_5165_627# VSS 0.0996f
C5179 a_6040_993# VSS 0.239f
C5180 a_6199_895# VSS 0.437f
C5181 a_5725_601# VSS 0.357f
C5182 a_5257_993# VSS 0.258f
C5183 a_5431_601# VSS 0.276f
C5184 a_4977_627# VSS 0.31f
C5185 D[5] VSS 1.58f
C5186 a_4811_627# VSS 0.699f
C5187 VDD_SW[6] VSS 0.411f
C5188 a_3755_627# VSS 0.00192f
C5189 a_3947_627# VSS 0.166f
C5190 a_4528_627# VSS 0.22f
C5191 VDD_SW_b[6] VSS 0.364f
C5192 a_3551_627# VSS 0.0108f
C5193 a_2973_627# VSS 0.0017f
C5194 a_3183_627# VSS 0.176f
C5195 a_3504_909# VSS 3.84e-19
C5196 a_2773_627# VSS 0.0996f
C5197 a_3648_993# VSS 0.239f
C5198 a_3807_895# VSS 0.438f
C5199 a_3333_601# VSS 0.358f
C5200 a_2865_993# VSS 0.258f
C5201 a_3039_601# VSS 0.277f
C5202 a_2585_627# VSS 0.31f
C5203 D[6] VSS 1.61f
C5204 a_2419_627# VSS 0.7f
C5205 VDD_SW[7] VSS 0.402f
C5206 a_1363_627# VSS 0.00192f
C5207 a_1555_627# VSS 0.166f
C5208 a_2136_627# VSS 0.22f
C5209 VDD_SW_b[7] VSS 0.364f
C5210 a_1159_627# VSS 0.0108f
C5211 a_581_627# VSS 0.0017f
C5212 a_791_627# VSS 0.176f
C5213 a_1112_909# VSS 3.84e-19
C5214 a_381_627# VSS 0.0996f
C5215 a_1256_993# VSS 0.239f
C5216 a_1415_895# VSS 0.437f
C5217 a_941_601# VSS 0.357f
C5218 a_473_993# VSS 0.258f
C5219 a_647_601# VSS 0.276f
C5220 a_193_627# VSS 0.312f
C5221 D[7] VSS 1.58f
C5222 a_27_627# VSS 0.749f
C5223 a_16330_1315# VSS 0.00411f
C5224 a_16109_1315# VSS 0.008f
C5225 a_14791_1315# VSS 0.0073f
C5226 a_14570_1315# VSS 0.00337f
C5227 x20.X VSS 0.761f
C5228 a_13936_1315# VSS 0.00335f
C5229 a_13715_1315# VSS 0.00726f
C5230 a_12399_1315# VSS 0.00726f
C5231 a_12178_1315# VSS 0.00335f
C5232 a_16323_1642# VSS 6.91e-19
C5233 a_16037_1642# VSS 3.55e-19
C5234 a_14887_1642# VSS 2.7e-19
C5235 a_14570_1642# VSS 7.29e-19
C5236 a_15855_1642# VSS 0.341f
C5237 a_14857_1289# VSS 0.339f
C5238 check[0] VSS 1.02f
C5239 x18.X VSS 0.324f
C5240 x17.X VSS 0.499f
C5241 a_11546_1315# VSS 0.00335f
C5242 a_11325_1315# VSS 0.00726f
C5243 a_10007_1315# VSS 0.00726f
C5244 a_9786_1315# VSS 0.00335f
C5245 a_13929_1642# VSS 3.69e-19
C5246 a_13643_1642# VSS 2.7e-19
C5247 a_12495_1642# VSS 2.7e-19
C5248 a_12178_1642# VSS 7.29e-19
C5249 a_13461_1642# VSS 0.34f
C5250 a_12465_1289# VSS 0.339f
C5251 check[1] VSS 1f
C5252 x16.X VSS 0.325f
C5253 x15.X VSS 0.498f
C5254 a_9154_1315# VSS 0.00335f
C5255 a_8933_1315# VSS 0.00726f
C5256 a_7615_1315# VSS 0.00726f
C5257 a_7394_1315# VSS 0.00335f
C5258 a_11539_1642# VSS 4e-19
C5259 a_11253_1642# VSS 2.7e-19
C5260 a_10103_1642# VSS 2.7e-19
C5261 a_9786_1642# VSS 7.29e-19
C5262 a_11071_1642# VSS 0.34f
C5263 a_10073_1289# VSS 0.339f
C5264 check[2] VSS 1f
C5265 x14.X VSS 0.324f
C5266 x13.X VSS 0.498f
C5267 a_6760_1315# VSS 0.00335f
C5268 a_6539_1315# VSS 0.00726f
C5269 a_5223_1315# VSS 0.00726f
C5270 a_5002_1315# VSS 0.00335f
C5271 a_9147_1642# VSS 4e-19
C5272 a_8861_1642# VSS 2.7e-19
C5273 a_7711_1642# VSS 2.7e-19
C5274 a_7394_1642# VSS 7.29e-19
C5275 a_8679_1642# VSS 0.34f
C5276 a_7681_1289# VSS 0.339f
C5277 check[3] VSS 1f
C5278 x12.X VSS 0.324f
C5279 x11.X VSS 0.498f
C5280 a_4370_1315# VSS 0.00335f
C5281 a_4149_1315# VSS 0.00726f
C5282 a_2831_1315# VSS 0.00726f
C5283 a_2610_1315# VSS 0.00335f
C5284 a_6753_1642# VSS 3.84e-19
C5285 a_6467_1642# VSS 2.7e-19
C5286 a_5319_1642# VSS 2.7e-19
C5287 a_5002_1642# VSS 7.29e-19
C5288 a_6285_1642# VSS 0.338f
C5289 a_5289_1289# VSS 0.338f
C5290 check[4] VSS 0.904f
C5291 x10.X VSS 0.323f
C5292 x9.X VSS 0.498f
C5293 a_1978_1315# VSS 0.00335f
C5294 a_1757_1315# VSS 0.00726f
C5295 a_439_1315# VSS 0.00726f
C5296 a_218_1315# VSS 0.00335f
C5297 a_4363_1642# VSS 4e-19
C5298 a_4077_1642# VSS 2.7e-19
C5299 a_2927_1642# VSS 2.7e-19
C5300 a_2610_1642# VSS 7.29e-19
C5301 a_3895_1642# VSS 0.34f
C5302 a_2897_1289# VSS 0.339f
C5303 check[5] VSS 0.983f
C5304 x8.X VSS 0.323f
C5305 x7.X VSS 0.499f
C5306 a_1971_1642# VSS 4e-19
C5307 a_1685_1642# VSS 2.7e-19
C5308 a_535_1642# VSS 2.7e-19
C5309 a_218_1642# VSS 7.29e-19
C5310 a_1503_1642# VSS 0.338f
C5311 a_505_1289# VSS 0.338f
C5312 check[6] VSS 0.911f
C5313 x6.X VSS 0.538f
C5314 a_16109_1642# VSS 0.35f
C5315 a_14428_1467# VSS 0.331f
C5316 a_13715_1642# VSS 0.326f
C5317 a_12036_1467# VSS 0.331f
C5318 a_11325_1642# VSS 0.326f
C5319 a_9644_1467# VSS 0.331f
C5320 a_8933_1642# VSS 0.326f
C5321 a_7252_1467# VSS 0.331f
C5322 a_6539_1642# VSS 0.325f
C5323 a_4860_1467# VSS 0.33f
C5324 a_4149_1642# VSS 0.325f
C5325 a_2468_1467# VSS 0.33f
C5326 a_1757_1642# VSS 0.325f
C5327 a_76_1467# VSS 0.343f
C5328 x9.A1 VSS 22.9f
C5329 x2.X VSS 22.8f
C5330 a_5323_2457# VSS 2.11f
C5331 x30.A VSS 0.954f
C5332 a_4689_2457# VSS 0.532f
C5333 x27.A VSS 0.207f
C5334 a_4413_2457# VSS 0.279f
C5335 ready VSS 2.3f
C5336 a_939_2457# VSS 2.02f
C5337 x3.X VSS 0.913f
C5338 a_305_2457# VSS 0.51f
C5339 x3.A VSS 0.196f
C5340 a_29_2457# VSS 0.274f
C5341 reset VSS 0.202f
C5342 VDD VSS 0.113p
C5343 x9.A1.n0 VSS 0.00514f
C5344 x9.A1.n1 VSS 0.00514f
C5345 x9.A1.n2 VSS 0.00514f
C5346 x9.A1.n3 VSS 0.00514f
C5347 x9.A1.n4 VSS 0.00514f
C5348 x9.A1.n5 VSS 0.00514f
C5349 x9.A1.n6 VSS 0.00514f
C5350 x9.A1.t24 VSS 0.00668f
C5351 x9.A1.t18 VSS 0.00668f
C5352 x9.A1.n7 VSS 0.0165f
C5353 x9.A1.t28 VSS 0.00668f
C5354 x9.A1.t20 VSS 0.00668f
C5355 x9.A1.n8 VSS 0.0255f
C5356 x9.A1.t27 VSS 0.00668f
C5357 x9.A1.t22 VSS 0.00668f
C5358 x9.A1.n9 VSS 0.0165f
C5359 x9.A1.n10 VSS 0.0642f
C5360 x9.A1.t30 VSS 0.00668f
C5361 x9.A1.t16 VSS 0.00668f
C5362 x9.A1.n11 VSS 0.0165f
C5363 x9.A1.n12 VSS 0.0387f
C5364 x9.A1.t25 VSS 0.00668f
C5365 x9.A1.t17 VSS 0.00668f
C5366 x9.A1.n13 VSS 0.0165f
C5367 x9.A1.n14 VSS 0.0387f
C5368 x9.A1.t26 VSS 0.00668f
C5369 x9.A1.t19 VSS 0.00668f
C5370 x9.A1.n15 VSS 0.0165f
C5371 x9.A1.n16 VSS 0.0387f
C5372 x9.A1.t29 VSS 0.00668f
C5373 x9.A1.t21 VSS 0.00668f
C5374 x9.A1.n17 VSS 0.0165f
C5375 x9.A1.n18 VSS 0.0387f
C5376 x9.A1.t31 VSS 0.00668f
C5377 x9.A1.t23 VSS 0.00668f
C5378 x9.A1.n19 VSS 0.0165f
C5379 x9.A1.n20 VSS 0.0387f
C5380 x9.A1.n21 VSS 0.0369f
C5381 x9.A1.n22 VSS 0.0039f
C5382 x9.A1.t42 VSS 0.0183f
C5383 x9.A1.n23 VSS 0.0301f
C5384 x9.A1.t55 VSS 0.0052f
C5385 x9.A1.n24 VSS 0.0153f
C5386 x9.A1.n25 VSS 0.00192f
C5387 x9.A1.n26 VSS 0.00107f
C5388 x9.A1.n27 VSS 0.00111f
C5389 x9.A1.n28 VSS 0.00346f
C5390 x9.A1.n29 VSS 0.00582f
C5391 x9.A1.n30 VSS 0.0442f
C5392 x9.A1.n31 VSS 0.00334f
C5393 x9.A1.t32 VSS 0.00523f
C5394 x9.A1.n32 VSS 0.015f
C5395 x9.A1.n33 VSS 0.00195f
C5396 x9.A1.t43 VSS 0.0183f
C5397 x9.A1.n34 VSS 0.0302f
C5398 x9.A1.n35 VSS 0.00111f
C5399 x9.A1.n36 VSS 0.00582f
C5400 x9.A1.n37 VSS 0.0388f
C5401 x9.A1.n38 VSS 0.119f
C5402 x9.A1.n39 VSS 0.0039f
C5403 x9.A1.t53 VSS 0.0183f
C5404 x9.A1.n40 VSS 0.0302f
C5405 x9.A1.t40 VSS 0.0052f
C5406 x9.A1.n41 VSS 0.015f
C5407 x9.A1.n42 VSS 0.00211f
C5408 x9.A1.n43 VSS 0.00107f
C5409 x9.A1.n44 VSS 0.00111f
C5410 x9.A1.n45 VSS 0.00346f
C5411 x9.A1.n46 VSS 0.00582f
C5412 x9.A1.n47 VSS 0.0388f
C5413 x9.A1.n48 VSS 0.115f
C5414 x9.A1.n49 VSS 0.00334f
C5415 x9.A1.t44 VSS 0.00526f
C5416 x9.A1.n50 VSS 0.015f
C5417 x9.A1.n51 VSS 0.002f
C5418 x9.A1.t56 VSS 0.0183f
C5419 x9.A1.n52 VSS 0.0302f
C5420 x9.A1.n53 VSS 0.00114f
C5421 x9.A1.n54 VSS 0.00582f
C5422 x9.A1.n55 VSS 0.0388f
C5423 x9.A1.n56 VSS 0.114f
C5424 x9.A1.n57 VSS 0.0039f
C5425 x9.A1.t48 VSS 0.0183f
C5426 x9.A1.n58 VSS 0.0301f
C5427 x9.A1.t35 VSS 0.0052f
C5428 x9.A1.n59 VSS 0.0153f
C5429 x9.A1.n60 VSS 0.00192f
C5430 x9.A1.n61 VSS 0.00107f
C5431 x9.A1.n62 VSS 0.00111f
C5432 x9.A1.n63 VSS 0.00346f
C5433 x9.A1.n64 VSS 0.00582f
C5434 x9.A1.n65 VSS 0.0388f
C5435 x9.A1.n66 VSS 0.115f
C5436 x9.A1.n67 VSS 0.00334f
C5437 x9.A1.t57 VSS 0.00523f
C5438 x9.A1.n68 VSS 0.015f
C5439 x9.A1.n69 VSS 0.00195f
C5440 x9.A1.t58 VSS 0.0183f
C5441 x9.A1.n70 VSS 0.0302f
C5442 x9.A1.n71 VSS 0.00111f
C5443 x9.A1.n72 VSS 0.00582f
C5444 x9.A1.n73 VSS 0.0388f
C5445 x9.A1.n74 VSS 0.115f
C5446 x9.A1.n75 VSS 0.0039f
C5447 x9.A1.t34 VSS 0.0183f
C5448 x9.A1.n76 VSS 0.0302f
C5449 x9.A1.t33 VSS 0.0052f
C5450 x9.A1.n77 VSS 0.015f
C5451 x9.A1.n78 VSS 0.00211f
C5452 x9.A1.n79 VSS 0.00107f
C5453 x9.A1.n80 VSS 0.00111f
C5454 x9.A1.n81 VSS 0.00346f
C5455 x9.A1.n82 VSS 0.00582f
C5456 x9.A1.n83 VSS 0.0388f
C5457 x9.A1.n84 VSS 0.115f
C5458 x9.A1.n85 VSS 0.00334f
C5459 x9.A1.t59 VSS 0.00523f
C5460 x9.A1.n86 VSS 0.0146f
C5461 x9.A1.n87 VSS 0.00236f
C5462 x9.A1.t41 VSS 0.0183f
C5463 x9.A1.n88 VSS 0.0302f
C5464 x9.A1.n89 VSS 0.00109f
C5465 x9.A1.n90 VSS 0.00582f
C5466 x9.A1.n91 VSS 0.0388f
C5467 x9.A1.n92 VSS 0.0764f
C5468 x9.A1.n93 VSS 0.0039f
C5469 x9.A1.t51 VSS 0.0183f
C5470 x9.A1.n94 VSS 0.0301f
C5471 x9.A1.t54 VSS 0.0052f
C5472 x9.A1.n95 VSS 0.0153f
C5473 x9.A1.n96 VSS 0.00192f
C5474 x9.A1.n97 VSS 0.00107f
C5475 x9.A1.n98 VSS 0.00111f
C5476 x9.A1.n99 VSS 0.00346f
C5477 x9.A1.n100 VSS 0.00582f
C5478 x9.A1.n101 VSS 0.0384f
C5479 x9.A1.n102 VSS 0.00334f
C5480 x9.A1.t36 VSS 0.00524f
C5481 x9.A1.n103 VSS 0.0146f
C5482 x9.A1.n104 VSS 0.00229f
C5483 x9.A1.t45 VSS 0.0183f
C5484 x9.A1.n105 VSS 0.0303f
C5485 x9.A1.n106 VSS 0.00111f
C5486 x9.A1.n107 VSS 0.00582f
C5487 x9.A1.n108 VSS 0.0388f
C5488 x9.A1.n109 VSS 0.0039f
C5489 x9.A1.t46 VSS 0.0183f
C5490 x9.A1.n110 VSS 0.0302f
C5491 x9.A1.t49 VSS 0.00523f
C5492 x9.A1.n111 VSS 0.015f
C5493 x9.A1.n112 VSS 0.00217f
C5494 x9.A1.n113 VSS 0.00109f
C5495 x9.A1.n114 VSS 0.00111f
C5496 x9.A1.n115 VSS 0.00346f
C5497 x9.A1.n116 VSS 0.00582f
C5498 x9.A1.n117 VSS 0.0388f
C5499 x9.A1.n118 VSS 0.00334f
C5500 x9.A1.t37 VSS 0.00524f
C5501 x9.A1.n119 VSS 0.0146f
C5502 x9.A1.n120 VSS 0.00229f
C5503 x9.A1.t47 VSS 0.0183f
C5504 x9.A1.n121 VSS 0.0303f
C5505 x9.A1.n122 VSS 0.00111f
C5506 x9.A1.n123 VSS 0.00582f
C5507 x9.A1.n124 VSS 0.0388f
C5508 x9.A1.n125 VSS 0.0039f
C5509 x9.A1.t39 VSS 0.0183f
C5510 x9.A1.n126 VSS 0.0302f
C5511 x9.A1.t50 VSS 0.00523f
C5512 x9.A1.n127 VSS 0.015f
C5513 x9.A1.n128 VSS 0.00217f
C5514 x9.A1.n129 VSS 0.00109f
C5515 x9.A1.n130 VSS 0.00111f
C5516 x9.A1.n131 VSS 0.00346f
C5517 x9.A1.n132 VSS 0.00582f
C5518 x9.A1.n133 VSS 0.0388f
C5519 x9.A1.n134 VSS 0.00334f
C5520 x9.A1.t52 VSS 0.00523f
C5521 x9.A1.n135 VSS 0.015f
C5522 x9.A1.n136 VSS 0.00204f
C5523 x9.A1.t38 VSS 0.0183f
C5524 x9.A1.n137 VSS 0.0302f
C5525 x9.A1.n138 VSS 0.00109f
C5526 x9.A1.n139 VSS 0.00582f
C5527 x9.A1.n140 VSS 0.0599f
C5528 x9.A1.n141 VSS 0.132f
C5529 x9.A1.n142 VSS 0.115f
C5530 x9.A1.n143 VSS 0.115f
C5531 x9.A1.n144 VSS 0.115f
C5532 x9.A1.n145 VSS 0.105f
C5533 x9.A1.n146 VSS 0.129f
C5534 x9.A1.n147 VSS 0.0488f
C5535 x9.A1.t4 VSS 0.00434f
C5536 x9.A1.t12 VSS 0.00434f
C5537 x9.A1.n148 VSS 0.0206f
C5538 x9.A1.t3 VSS 0.00434f
C5539 x9.A1.t14 VSS 0.00434f
C5540 x9.A1.n149 VSS 0.0109f
C5541 x9.A1.n150 VSS 0.0407f
C5542 x9.A1.t6 VSS 0.00434f
C5543 x9.A1.t8 VSS 0.00434f
C5544 x9.A1.n151 VSS 0.0109f
C5545 x9.A1.n152 VSS 0.0274f
C5546 x9.A1.t1 VSS 0.00434f
C5547 x9.A1.t9 VSS 0.00434f
C5548 x9.A1.n153 VSS 0.0109f
C5549 x9.A1.n154 VSS 0.0274f
C5550 x9.A1.t2 VSS 0.00434f
C5551 x9.A1.t11 VSS 0.00434f
C5552 x9.A1.n155 VSS 0.0109f
C5553 x9.A1.n156 VSS 0.0274f
C5554 x9.A1.t5 VSS 0.00434f
C5555 x9.A1.t13 VSS 0.00434f
C5556 x9.A1.n157 VSS 0.0109f
C5557 x9.A1.n158 VSS 0.0274f
C5558 x9.A1.t7 VSS 0.00434f
C5559 x9.A1.t15 VSS 0.00434f
C5560 x9.A1.n159 VSS 0.0109f
C5561 x9.A1.n160 VSS 0.0274f
C5562 x9.A1.t0 VSS 0.00434f
C5563 x9.A1.t10 VSS 0.00434f
C5564 x9.A1.n161 VSS 0.0109f
C5565 x9.A1.n162 VSS 0.0271f
C5566 x2.X.n0 VSS 0.004f
C5567 x2.X.n1 VSS 0.004f
C5568 x2.X.n2 VSS 0.004f
C5569 x2.X.n3 VSS 0.004f
C5570 x2.X.n4 VSS 0.004f
C5571 x2.X.n5 VSS 0.004f
C5572 x2.X.n6 VSS 0.004f
C5573 x2.X.n7 VSS 0.00187f
C5574 x2.X.t69 VSS 0.0137f
C5575 x2.X.n8 VSS 0.0191f
C5576 x2.X.t55 VSS 0.00603f
C5577 x2.X.n9 VSS 0.00794f
C5578 x2.X.n10 VSS 0.00797f
C5579 x2.X.n11 VSS 0.00622f
C5580 x2.X.n12 VSS 0.038f
C5581 x2.X.t52 VSS 0.0143f
C5582 x2.X.t51 VSS 0.00602f
C5583 x2.X.n13 VSS 0.0272f
C5584 x2.X.n14 VSS 0.00786f
C5585 x2.X.n15 VSS 0.00309f
C5586 x2.X.n16 VSS 0.00163f
C5587 x2.X.n17 VSS 0.00223f
C5588 x2.X.n18 VSS 0.0148f
C5589 x2.X.n19 VSS 0.0418f
C5590 x2.X.n20 VSS 0.00577f
C5591 x2.X.n21 VSS 0.00177f
C5592 x2.X.n22 VSS 0.00131f
C5593 x2.X.t65 VSS 0.00953f
C5594 x2.X.t50 VSS 0.00804f
C5595 x2.X.n23 VSS 0.0128f
C5596 x2.X.n24 VSS 0.0141f
C5597 x2.X.n25 VSS 0.0547f
C5598 x2.X.n26 VSS 0.28f
C5599 x2.X.n27 VSS 0.00187f
C5600 x2.X.t72 VSS 0.0137f
C5601 x2.X.n28 VSS 0.0191f
C5602 x2.X.t57 VSS 0.00603f
C5603 x2.X.n29 VSS 0.00794f
C5604 x2.X.n30 VSS 0.00797f
C5605 x2.X.n31 VSS 0.00622f
C5606 x2.X.n32 VSS 0.038f
C5607 x2.X.t66 VSS 0.0143f
C5608 x2.X.t63 VSS 0.00602f
C5609 x2.X.n33 VSS 0.0272f
C5610 x2.X.n34 VSS 0.00786f
C5611 x2.X.n35 VSS 0.00309f
C5612 x2.X.n36 VSS 0.00163f
C5613 x2.X.n37 VSS 0.00223f
C5614 x2.X.n38 VSS 0.0148f
C5615 x2.X.n39 VSS 0.0418f
C5616 x2.X.n40 VSS 0.00577f
C5617 x2.X.n41 VSS 0.00177f
C5618 x2.X.n42 VSS 0.00131f
C5619 x2.X.t70 VSS 0.00953f
C5620 x2.X.t54 VSS 0.00804f
C5621 x2.X.n43 VSS 0.0128f
C5622 x2.X.n44 VSS 0.0141f
C5623 x2.X.n45 VSS 0.0546f
C5624 x2.X.n46 VSS 0.216f
C5625 x2.X.n47 VSS 0.425f
C5626 x2.X.n48 VSS 0.00187f
C5627 x2.X.t39 VSS 0.0137f
C5628 x2.X.n49 VSS 0.0191f
C5629 x2.X.t59 VSS 0.00603f
C5630 x2.X.n50 VSS 0.00794f
C5631 x2.X.n51 VSS 0.00797f
C5632 x2.X.n52 VSS 0.00622f
C5633 x2.X.n53 VSS 0.038f
C5634 x2.X.t68 VSS 0.0143f
C5635 x2.X.t67 VSS 0.00602f
C5636 x2.X.n54 VSS 0.0272f
C5637 x2.X.n55 VSS 0.00786f
C5638 x2.X.n56 VSS 0.00309f
C5639 x2.X.n57 VSS 0.00163f
C5640 x2.X.n58 VSS 0.00223f
C5641 x2.X.n59 VSS 0.0148f
C5642 x2.X.n60 VSS 0.0428f
C5643 x2.X.n61 VSS 0.00595f
C5644 x2.X.n62 VSS 0.00177f
C5645 x2.X.n63 VSS 0.00131f
C5646 x2.X.t73 VSS 0.00953f
C5647 x2.X.t56 VSS 0.00804f
C5648 x2.X.n64 VSS 0.0128f
C5649 x2.X.n65 VSS 0.0141f
C5650 x2.X.n66 VSS 0.0546f
C5651 x2.X.n67 VSS 0.216f
C5652 x2.X.n68 VSS 0.392f
C5653 x2.X.n69 VSS 0.00187f
C5654 x2.X.t58 VSS 0.0137f
C5655 x2.X.n70 VSS 0.0191f
C5656 x2.X.t38 VSS 0.00603f
C5657 x2.X.n71 VSS 0.00794f
C5658 x2.X.n72 VSS 0.00797f
C5659 x2.X.n73 VSS 0.00622f
C5660 x2.X.n74 VSS 0.038f
C5661 x2.X.t37 VSS 0.0143f
C5662 x2.X.t36 VSS 0.00602f
C5663 x2.X.n75 VSS 0.0272f
C5664 x2.X.n76 VSS 0.00786f
C5665 x2.X.n77 VSS 0.00309f
C5666 x2.X.n78 VSS 0.00163f
C5667 x2.X.n79 VSS 0.00223f
C5668 x2.X.n80 VSS 0.0149f
C5669 x2.X.n81 VSS 0.042f
C5670 x2.X.n82 VSS 0.00577f
C5671 x2.X.n83 VSS 0.00177f
C5672 x2.X.n84 VSS 0.00131f
C5673 x2.X.t41 VSS 0.00953f
C5674 x2.X.t71 VSS 0.00804f
C5675 x2.X.n85 VSS 0.0128f
C5676 x2.X.n86 VSS 0.0141f
C5677 x2.X.n87 VSS 0.0546f
C5678 x2.X.n88 VSS 0.216f
C5679 x2.X.n89 VSS 0.392f
C5680 x2.X.n90 VSS 0.00187f
C5681 x2.X.t60 VSS 0.0137f
C5682 x2.X.n91 VSS 0.0191f
C5683 x2.X.t46 VSS 0.00603f
C5684 x2.X.n92 VSS 0.00794f
C5685 x2.X.n93 VSS 0.00797f
C5686 x2.X.n94 VSS 0.00622f
C5687 x2.X.n95 VSS 0.038f
C5688 x2.X.t42 VSS 0.0143f
C5689 x2.X.t40 VSS 0.00602f
C5690 x2.X.n96 VSS 0.0272f
C5691 x2.X.n97 VSS 0.00786f
C5692 x2.X.n98 VSS 0.00309f
C5693 x2.X.n99 VSS 0.00163f
C5694 x2.X.n100 VSS 0.00223f
C5695 x2.X.n101 VSS 0.0149f
C5696 x2.X.n102 VSS 0.042f
C5697 x2.X.n103 VSS 0.00577f
C5698 x2.X.n104 VSS 0.00177f
C5699 x2.X.n105 VSS 0.00131f
C5700 x2.X.t48 VSS 0.00953f
C5701 x2.X.t32 VSS 0.00804f
C5702 x2.X.n106 VSS 0.0128f
C5703 x2.X.n107 VSS 0.0141f
C5704 x2.X.n108 VSS 0.0546f
C5705 x2.X.n109 VSS 0.216f
C5706 x2.X.n110 VSS 0.392f
C5707 x2.X.n111 VSS 0.00187f
C5708 x2.X.t33 VSS 0.0137f
C5709 x2.X.n112 VSS 0.0191f
C5710 x2.X.t61 VSS 0.00603f
C5711 x2.X.n113 VSS 0.00794f
C5712 x2.X.n114 VSS 0.00797f
C5713 x2.X.n115 VSS 0.00622f
C5714 x2.X.n116 VSS 0.038f
C5715 x2.X.t49 VSS 0.0143f
C5716 x2.X.t45 VSS 0.00602f
C5717 x2.X.n117 VSS 0.0272f
C5718 x2.X.n118 VSS 0.00786f
C5719 x2.X.n119 VSS 0.00309f
C5720 x2.X.n120 VSS 0.00163f
C5721 x2.X.n121 VSS 0.00223f
C5722 x2.X.n122 VSS 0.0149f
C5723 x2.X.n123 VSS 0.042f
C5724 x2.X.n124 VSS 0.00577f
C5725 x2.X.n125 VSS 0.00177f
C5726 x2.X.n126 VSS 0.00131f
C5727 x2.X.t62 VSS 0.00953f
C5728 x2.X.t44 VSS 0.00804f
C5729 x2.X.n127 VSS 0.0128f
C5730 x2.X.n128 VSS 0.0141f
C5731 x2.X.n129 VSS 0.0554f
C5732 x2.X.n130 VSS 0.215f
C5733 x2.X.n131 VSS 0.287f
C5734 x2.X.n132 VSS 0.00187f
C5735 x2.X.t35 VSS 0.0137f
C5736 x2.X.n133 VSS 0.0191f
C5737 x2.X.t64 VSS 0.00603f
C5738 x2.X.n134 VSS 0.00794f
C5739 x2.X.n135 VSS 0.00797f
C5740 x2.X.n136 VSS 0.00622f
C5741 x2.X.n137 VSS 0.038f
C5742 x2.X.t47 VSS 0.0143f
C5743 x2.X.t43 VSS 0.00602f
C5744 x2.X.n138 VSS 0.0272f
C5745 x2.X.n139 VSS 0.00786f
C5746 x2.X.n140 VSS 0.00309f
C5747 x2.X.n141 VSS 0.00163f
C5748 x2.X.n142 VSS 0.00223f
C5749 x2.X.n143 VSS 0.0148f
C5750 x2.X.n144 VSS 0.0418f
C5751 x2.X.n145 VSS 0.00577f
C5752 x2.X.n146 VSS 0.00177f
C5753 x2.X.n147 VSS 0.00131f
C5754 x2.X.t53 VSS 0.00957f
C5755 x2.X.t34 VSS 0.00803f
C5756 x2.X.n148 VSS 0.0125f
C5757 x2.X.n149 VSS 0.0144f
C5758 x2.X.n150 VSS 0.0541f
C5759 x2.X.n151 VSS 0.29f
C5760 x2.X.n152 VSS 0.273f
C5761 x2.X.t19 VSS 0.00902f
C5762 x2.X.t30 VSS 0.00902f
C5763 x2.X.n153 VSS 0.0223f
C5764 x2.X.t24 VSS 0.00902f
C5765 x2.X.t29 VSS 0.00902f
C5766 x2.X.n154 VSS 0.0223f
C5767 x2.X.t22 VSS 0.00902f
C5768 x2.X.t27 VSS 0.00902f
C5769 x2.X.n155 VSS 0.0223f
C5770 x2.X.t20 VSS 0.00902f
C5771 x2.X.t26 VSS 0.00902f
C5772 x2.X.n156 VSS 0.0223f
C5773 x2.X.t18 VSS 0.00902f
C5774 x2.X.t17 VSS 0.00902f
C5775 x2.X.n157 VSS 0.0223f
C5776 x2.X.t25 VSS 0.00902f
C5777 x2.X.t16 VSS 0.00902f
C5778 x2.X.n158 VSS 0.0223f
C5779 x2.X.t23 VSS 0.00902f
C5780 x2.X.t28 VSS 0.00902f
C5781 x2.X.n159 VSS 0.0223f
C5782 x2.X.t21 VSS 0.00902f
C5783 x2.X.t31 VSS 0.00902f
C5784 x2.X.n160 VSS 0.0344f
C5785 x2.X.n161 VSS 0.0867f
C5786 x2.X.n162 VSS 0.0523f
C5787 x2.X.n163 VSS 0.0523f
C5788 x2.X.n164 VSS 0.0523f
C5789 x2.X.n165 VSS 0.0523f
C5790 x2.X.n166 VSS 0.0523f
C5791 x2.X.n167 VSS 0.0498f
C5792 x2.X.n168 VSS 0.0229f
C5793 x2.X.t11 VSS 0.00586f
C5794 x2.X.t5 VSS 0.00586f
C5795 x2.X.n169 VSS 0.0278f
C5796 x2.X.t13 VSS 0.00586f
C5797 x2.X.t2 VSS 0.00586f
C5798 x2.X.n170 VSS 0.0147f
C5799 x2.X.n171 VSS 0.0549f
C5800 x2.X.t15 VSS 0.00586f
C5801 x2.X.t6 VSS 0.00586f
C5802 x2.X.n172 VSS 0.0147f
C5803 x2.X.n173 VSS 0.037f
C5804 x2.X.t8 VSS 0.00586f
C5805 x2.X.t7 VSS 0.00586f
C5806 x2.X.n174 VSS 0.0147f
C5807 x2.X.n175 VSS 0.0371f
C5808 x2.X.t10 VSS 0.00586f
C5809 x2.X.t0 VSS 0.00586f
C5810 x2.X.n176 VSS 0.0147f
C5811 x2.X.n177 VSS 0.0371f
C5812 x2.X.t12 VSS 0.00586f
C5813 x2.X.t1 VSS 0.00586f
C5814 x2.X.n178 VSS 0.0147f
C5815 x2.X.n179 VSS 0.0371f
C5816 x2.X.t14 VSS 0.00586f
C5817 x2.X.t3 VSS 0.00586f
C5818 x2.X.n180 VSS 0.0147f
C5819 x2.X.n181 VSS 0.0371f
C5820 x2.X.t9 VSS 0.00586f
C5821 x2.X.t4 VSS 0.00586f
C5822 x2.X.n182 VSS 0.0147f
C5823 x2.X.n183 VSS 0.0365f
C5824 VDD.t99 VSS 5.58e-19
C5825 VDD.t60 VSS 5.58e-19
C5826 VDD.n0 VSS 0.00121f
C5827 VDD.n1 VSS 0.00102f
C5828 VDD.n2 VSS 0.00167f
C5829 VDD.t11 VSS 5.58e-19
C5830 VDD.t7 VSS 5.58e-19
C5831 VDD.n3 VSS 0.00121f
C5832 VDD.n4 VSS 0.00102f
C5833 VDD.n5 VSS 0.00167f
C5834 VDD.t289 VSS 5.58e-19
C5835 VDD.t205 VSS 5.58e-19
C5836 VDD.n6 VSS 0.00121f
C5837 VDD.n7 VSS 0.00102f
C5838 VDD.n8 VSS 0.00167f
C5839 VDD.t421 VSS 5.58e-19
C5840 VDD.t653 VSS 5.58e-19
C5841 VDD.n9 VSS 0.00121f
C5842 VDD.n10 VSS 0.00102f
C5843 VDD.n11 VSS 0.00167f
C5844 VDD.t93 VSS 5.58e-19
C5845 VDD.t138 VSS 5.58e-19
C5846 VDD.n12 VSS 0.00121f
C5847 VDD.n13 VSS 0.0014f
C5848 VDD.t174 VSS 5.58e-19
C5849 VDD.t279 VSS 5.58e-19
C5850 VDD.n14 VSS 0.00121f
C5851 VDD.n15 VSS 0.00102f
C5852 VDD.n16 VSS 0.00167f
C5853 VDD.t662 VSS 5.58e-19
C5854 VDD.t26 VSS 5.58e-19
C5855 VDD.n17 VSS 0.00121f
C5856 VDD.n18 VSS 0.00141f
C5857 VDD.n19 VSS 0.00101f
C5858 VDD.t661 VSS 0.00437f
C5859 VDD.t25 VSS 0.00537f
C5860 VDD.n20 VSS 0.0049f
C5861 VDD.n21 VSS 0.00102f
C5862 VDD.n22 VSS 0.00187f
C5863 VDD.n23 VSS 0.0025f
C5864 VDD.n24 VSS 0.00259f
C5865 VDD.n25 VSS 0.0084f
C5866 VDD.n26 VSS 0.00101f
C5867 VDD.n27 VSS 0.0011f
C5868 VDD.n28 VSS 0.00285f
C5869 VDD.t689 VSS 0.00131f
C5870 VDD.t688 VSS 0.00537f
C5871 VDD.n29 VSS 0.00793f
C5872 VDD.n30 VSS 0.00102f
C5873 VDD.n31 VSS 0.00188f
C5874 VDD.n32 VSS 0.00289f
C5875 VDD.n33 VSS 0.00285f
C5876 VDD.t27 VSS 0.00537f
C5877 VDD.n34 VSS 0.00537f
C5878 VDD.n35 VSS 0.00101f
C5879 VDD.n36 VSS 0.0014f
C5880 VDD.n37 VSS 0.00285f
C5881 VDD.t437 VSS 0.00537f
C5882 VDD.n38 VSS 0.0049f
C5883 VDD.n39 VSS 0.00101f
C5884 VDD.n40 VSS 0.00172f
C5885 VDD.n41 VSS 0.00285f
C5886 VDD.t153 VSS 0.00992f
C5887 VDD.n42 VSS 0.007f
C5888 VDD.n43 VSS 0.00177f
C5889 VDD.n44 VSS 0.00164f
C5890 VDD.n45 VSS 0.00285f
C5891 VDD.n46 VSS 0.00183f
C5892 VDD.t154 VSS 5.02e-19
C5893 VDD.t506 VSS 5.29e-19
C5894 VDD.n47 VSS 0.0011f
C5895 VDD.n48 VSS 0.00261f
C5896 VDD.n49 VSS 0.00274f
C5897 VDD.n50 VSS 0.00139f
C5898 VDD.n51 VSS 1.26e-19
C5899 VDD.t540 VSS 0.00138f
C5900 VDD.t759 VSS 5.9e-19
C5901 VDD.n52 VSS 0.00258f
C5902 VDD.n53 VSS 2.16e-19
C5903 VDD.n54 VSS 6.27e-19
C5904 VDD.n55 VSS 0.00131f
C5905 VDD.n56 VSS 2.16e-19
C5906 VDD.n57 VSS 0.00359f
C5907 VDD.n58 VSS 4.92e-19
C5908 VDD.n59 VSS 9.75e-19
C5909 VDD.t766 VSS 5.82e-19
C5910 VDD.n60 VSS 0.00292f
C5911 VDD.t504 VSS 0.00174f
C5912 VDD.n61 VSS 0.00159f
C5913 VDD.n62 VSS 2.13e-19
C5914 VDD.n63 VSS 8.62e-19
C5915 VDD.n64 VSS 1.59e-19
C5916 VDD.n65 VSS 2.64e-19
C5917 VDD.n66 VSS 0.00143f
C5918 VDD.t505 VSS 0.0124f
C5919 VDD.t681 VSS 0.00502f
C5920 VDD.n67 VSS 0.0063f
C5921 VDD.n68 VSS 0.00107f
C5922 VDD.n69 VSS 0.00163f
C5923 VDD.n70 VSS 0.0027f
C5924 VDD.t316 VSS 8.96e-19
C5925 VDD.t152 VSS 0.00201f
C5926 VDD.n71 VSS 0.00323f
C5927 VDD.n72 VSS 0.00423f
C5928 VDD.t315 VSS 0.00525f
C5929 VDD.n73 VSS 0.00572f
C5930 VDD.n74 VSS 0.00101f
C5931 VDD.n75 VSS 9.47e-19
C5932 VDD.n76 VSS 0.00285f
C5933 VDD.t151 VSS 0.00537f
C5934 VDD.n77 VSS 0.00764f
C5935 VDD.n78 VSS 0.00101f
C5936 VDD.n79 VSS 0.00102f
C5937 VDD.n80 VSS 0.00285f
C5938 VDD.n81 VSS 0.0084f
C5939 VDD.n82 VSS 0.00101f
C5940 VDD.n83 VSS 0.00172f
C5941 VDD.n84 VSS 0.00285f
C5942 VDD.t438 VSS 0.00537f
C5943 VDD.n85 VSS 0.0049f
C5944 VDD.n86 VSS 0.00101f
C5945 VDD.n87 VSS 0.00172f
C5946 VDD.n88 VSS 0.00285f
C5947 VDD.t28 VSS 0.00537f
C5948 VDD.n89 VSS 0.00589f
C5949 VDD.n90 VSS 0.00101f
C5950 VDD.n91 VSS 0.00172f
C5951 VDD.n92 VSS 0.00285f
C5952 VDD.t119 VSS 0.00537f
C5953 VDD.n93 VSS 0.0056f
C5954 VDD.n94 VSS 0.00101f
C5955 VDD.n95 VSS 0.00122f
C5956 VDD.n96 VSS 0.00285f
C5957 VDD.t120 VSS 7.06e-19
C5958 VDD.t542 VSS 5.29e-19
C5959 VDD.n97 VSS 0.00129f
C5960 VDD.t541 VSS 0.00537f
C5961 VDD.n98 VSS 0.00706f
C5962 VDD.n99 VSS 0.00102f
C5963 VDD.n100 VSS 0.00189f
C5964 VDD.n101 VSS 0.00234f
C5965 VDD.n102 VSS 0.00285f
C5966 VDD.n103 VSS 0.00618f
C5967 VDD.n104 VSS 0.00101f
C5968 VDD.n105 VSS 0.00152f
C5969 VDD.n106 VSS 0.00285f
C5970 VDD.t312 VSS 0.00537f
C5971 VDD.t313 VSS 0.00537f
C5972 VDD.n107 VSS 0.0042f
C5973 VDD.n108 VSS 0.00101f
C5974 VDD.n109 VSS 0.0016f
C5975 VDD.n110 VSS 0.00285f
C5976 VDD.t314 VSS 0.00243f
C5977 VDD.n111 VSS 0.00251f
C5978 VDD.n112 VSS 0.00817f
C5979 VDD.n113 VSS 9.18e-19
C5980 VDD.n114 VSS 0.00212f
C5981 VDD.n115 VSS 0.00285f
C5982 VDD.n116 VSS 0.00197f
C5983 VDD.n117 VSS 3.68e-19
C5984 VDD.n118 VSS 0.00165f
C5985 VDD.n119 VSS 5e-19
C5986 VDD.n120 VSS 9.34e-20
C5987 VDD.n121 VSS 0.00531f
C5988 VDD.n122 VSS 9.92e-19
C5989 VDD.t33 VSS 0.00543f
C5990 VDD.n123 VSS 0.00192f
C5991 VDD.n124 VSS 5.16e-19
C5992 VDD.n125 VSS 3.9e-19
C5993 VDD.n126 VSS 0.00169f
C5994 VDD.n127 VSS 0.00118f
C5995 VDD.n128 VSS 0.00116f
C5996 VDD.n129 VSS 0.00152f
C5997 VDD.t34 VSS 8.48e-19
C5998 VDD.t118 VSS -4.69e-19
C5999 VDD.n130 VSS 0.00333f
C6000 VDD.n131 VSS 6.2e-19
C6001 VDD.n132 VSS 0.00135f
C6002 VDD.n133 VSS 5e-19
C6003 VDD.t117 VSS 0.00432f
C6004 VDD.n134 VSS 0.0021f
C6005 VDD.n135 VSS 0.00455f
C6006 VDD.n136 VSS 6.04e-19
C6007 VDD.n137 VSS 3.9e-19
C6008 VDD.n138 VSS 1.3e-19
C6009 VDD.n139 VSS 2.64e-19
C6010 VDD.n140 VSS 0.00143f
C6011 VDD.n141 VSS 0.00858f
C6012 VDD.n142 VSS 9.12e-19
C6013 VDD.n143 VSS 0.00151f
C6014 VDD.n144 VSS 0.00284f
C6015 VDD.t121 VSS 0.00537f
C6016 VDD.n145 VSS 0.00776f
C6017 VDD.n146 VSS 0.00101f
C6018 VDD.n147 VSS 0.00172f
C6019 VDD.n148 VSS 0.00285f
C6020 VDD.t122 VSS 7.86e-19
C6021 VDD.t197 VSS -2.51e-19
C6022 VDD.n149 VSS 0.00362f
C6023 VDD.n150 VSS 0.00382f
C6024 VDD.t196 VSS 0.00537f
C6025 VDD.n151 VSS 0.00554f
C6026 VDD.n152 VSS 0.00101f
C6027 VDD.n153 VSS 9.18e-19
C6028 VDD.n154 VSS 0.00285f
C6029 VDD.n155 VSS 0.00214f
C6030 VDD.n156 VSS 9.77e-19
C6031 VDD.n157 VSS 0.00101f
C6032 VDD.n158 VSS 0.00817f
C6033 VDD.t278 VSS 0.00537f
C6034 VDD.n159 VSS 0.0049f
C6035 VDD.t173 VSS 0.00437f
C6036 VDD.n160 VSS 0.00101f
C6037 VDD.n161 VSS 0.0014f
C6038 VDD.n162 VSS 0.00187f
C6039 VDD.n163 VSS 0.0025f
C6040 VDD.n164 VSS 0.00259f
C6041 VDD.n165 VSS 0.0084f
C6042 VDD.n166 VSS 0.00101f
C6043 VDD.n167 VSS 0.0011f
C6044 VDD.n168 VSS 0.00285f
C6045 VDD.t283 VSS 0.00131f
C6046 VDD.t282 VSS 0.00537f
C6047 VDD.n169 VSS 0.00793f
C6048 VDD.n170 VSS 0.00102f
C6049 VDD.n171 VSS 0.00188f
C6050 VDD.n172 VSS 0.00289f
C6051 VDD.n173 VSS 0.00285f
C6052 VDD.t280 VSS 0.00537f
C6053 VDD.n174 VSS 0.00537f
C6054 VDD.n175 VSS 0.00101f
C6055 VDD.n176 VSS 0.0014f
C6056 VDD.n177 VSS 0.00285f
C6057 VDD.t208 VSS 0.00537f
C6058 VDD.n178 VSS 0.0049f
C6059 VDD.n179 VSS 0.00101f
C6060 VDD.n180 VSS 0.00172f
C6061 VDD.n181 VSS 0.00285f
C6062 VDD.t441 VSS 0.00992f
C6063 VDD.n182 VSS 0.007f
C6064 VDD.n183 VSS 0.00177f
C6065 VDD.n184 VSS 0.00164f
C6066 VDD.n185 VSS 0.00285f
C6067 VDD.n186 VSS 0.00183f
C6068 VDD.t442 VSS 5.02e-19
C6069 VDD.t503 VSS 5.29e-19
C6070 VDD.n187 VSS 0.0011f
C6071 VDD.n188 VSS 0.00261f
C6072 VDD.n189 VSS 0.00274f
C6073 VDD.n190 VSS 0.00135f
C6074 VDD.n191 VSS 1.26e-19
C6075 VDD.t519 VSS 0.00138f
C6076 VDD.t767 VSS 5.9e-19
C6077 VDD.n192 VSS 0.00258f
C6078 VDD.n193 VSS 2.16e-19
C6079 VDD.n194 VSS 6.27e-19
C6080 VDD.n195 VSS 0.00131f
C6081 VDD.n196 VSS 2.16e-19
C6082 VDD.n197 VSS 0.00359f
C6083 VDD.n198 VSS 4.92e-19
C6084 VDD.n199 VSS 9.75e-19
C6085 VDD.t769 VSS 5.82e-19
C6086 VDD.n200 VSS 0.00292f
C6087 VDD.t501 VSS 0.00175f
C6088 VDD.n201 VSS 0.00161f
C6089 VDD.n202 VSS 2.15e-19
C6090 VDD.n203 VSS 8.62e-19
C6091 VDD.n204 VSS 1.59e-19
C6092 VDD.n205 VSS 2.64e-19
C6093 VDD.n206 VSS 0.00143f
C6094 VDD.t502 VSS 0.0124f
C6095 VDD.t709 VSS 0.00502f
C6096 VDD.n207 VSS 0.0063f
C6097 VDD.n208 VSS 9.56e-19
C6098 VDD.n209 VSS 0.00163f
C6099 VDD.n210 VSS 0.0027f
C6100 VDD.t361 VSS 8.96e-19
C6101 VDD.t444 VSS 0.00201f
C6102 VDD.n211 VSS 0.00323f
C6103 VDD.n212 VSS 0.00423f
C6104 VDD.t360 VSS 0.00525f
C6105 VDD.n213 VSS 0.00572f
C6106 VDD.n214 VSS 0.00101f
C6107 VDD.n215 VSS 9.47e-19
C6108 VDD.n216 VSS 0.00285f
C6109 VDD.t443 VSS 0.00537f
C6110 VDD.n217 VSS 0.00764f
C6111 VDD.n218 VSS 0.00101f
C6112 VDD.n219 VSS 0.00102f
C6113 VDD.n220 VSS 0.00285f
C6114 VDD.n221 VSS 0.0084f
C6115 VDD.n222 VSS 0.00101f
C6116 VDD.n223 VSS 0.00172f
C6117 VDD.n224 VSS 0.00285f
C6118 VDD.t209 VSS 0.00537f
C6119 VDD.n225 VSS 0.0049f
C6120 VDD.n226 VSS 0.00101f
C6121 VDD.n227 VSS 0.00172f
C6122 VDD.n228 VSS 0.00285f
C6123 VDD.t281 VSS 0.00537f
C6124 VDD.n229 VSS 0.00589f
C6125 VDD.n230 VSS 0.00101f
C6126 VDD.n231 VSS 0.00172f
C6127 VDD.n232 VSS 0.00285f
C6128 VDD.t586 VSS 0.00537f
C6129 VDD.n233 VSS 0.0056f
C6130 VDD.n234 VSS 0.00101f
C6131 VDD.n235 VSS 0.00122f
C6132 VDD.n236 VSS 0.00285f
C6133 VDD.t587 VSS 7.06e-19
C6134 VDD.t521 VSS 5.29e-19
C6135 VDD.n237 VSS 0.00129f
C6136 VDD.t520 VSS 0.00537f
C6137 VDD.n238 VSS 0.00706f
C6138 VDD.n239 VSS 0.00102f
C6139 VDD.n240 VSS 0.00189f
C6140 VDD.n241 VSS 0.00234f
C6141 VDD.n242 VSS 0.00285f
C6142 VDD.n243 VSS 0.00618f
C6143 VDD.n244 VSS 0.00101f
C6144 VDD.n245 VSS 0.00152f
C6145 VDD.n246 VSS 0.00285f
C6146 VDD.t424 VSS 0.00537f
C6147 VDD.t358 VSS 0.00537f
C6148 VDD.n247 VSS 0.0042f
C6149 VDD.n248 VSS 0.00101f
C6150 VDD.n249 VSS 0.0016f
C6151 VDD.n250 VSS 0.00285f
C6152 VDD.t359 VSS 0.00243f
C6153 VDD.n251 VSS 0.00251f
C6154 VDD.n252 VSS 0.00922f
C6155 VDD.n253 VSS 0.00102f
C6156 VDD.n254 VSS 0.00214f
C6157 VDD.n255 VSS 0.00261f
C6158 VDD.n256 VSS 0.00119f
C6159 VDD.n257 VSS 0.00833f
C6160 VDD.n258 VSS 0.00199f
C6161 VDD.n259 VSS 0.00186f
C6162 VDD.n260 VSS 5e-19
C6163 VDD.t594 VSS 0.00432f
C6164 VDD.n261 VSS 0.00181f
C6165 VDD.n262 VSS 0.00642f
C6166 VDD.n263 VSS 6.04e-19
C6167 VDD.n264 VSS 3.9e-19
C6168 VDD.n265 VSS 3.68e-19
C6169 VDD.n266 VSS 2.5e-19
C6170 VDD.n267 VSS 0.00128f
C6171 VDD.n268 VSS 0.00807f
C6172 VDD.t595 VSS 8.48e-19
C6173 VDD.t589 VSS -4.69e-19
C6174 VDD.n269 VSS 0.00333f
C6175 VDD.n270 VSS 0.00188f
C6176 VDD.t588 VSS 0.00537f
C6177 VDD.n271 VSS 0.00566f
C6178 VDD.n272 VSS 9.12e-19
C6179 VDD.n273 VSS 0.00173f
C6180 VDD.n274 VSS 0.00158f
C6181 VDD.n275 VSS 0.00858f
C6182 VDD.n276 VSS 0.00101f
C6183 VDD.n277 VSS 0.00165f
C6184 VDD.n278 VSS 0.00285f
C6185 VDD.t584 VSS 0.00537f
C6186 VDD.n279 VSS 0.00776f
C6187 VDD.n280 VSS 0.00101f
C6188 VDD.n281 VSS 0.00172f
C6189 VDD.n282 VSS 0.00285f
C6190 VDD.t585 VSS 7.86e-19
C6191 VDD.t271 VSS -2.51e-19
C6192 VDD.n283 VSS 0.00362f
C6193 VDD.n284 VSS 0.00382f
C6194 VDD.t270 VSS 0.00537f
C6195 VDD.n285 VSS 0.00554f
C6196 VDD.n286 VSS 0.00101f
C6197 VDD.n287 VSS 9.18e-19
C6198 VDD.n288 VSS 0.00285f
C6199 VDD.n289 VSS 9.77e-19
C6200 VDD.n290 VSS 0.00214f
C6201 VDD.n291 VSS 0.00167f
C6202 VDD.n292 VSS 0.00101f
C6203 VDD.n293 VSS 0.00817f
C6204 VDD.n294 VSS 0.00101f
C6205 VDD.t92 VSS 0.00437f
C6206 VDD.t137 VSS 0.00537f
C6207 VDD.n295 VSS 0.0049f
C6208 VDD.n296 VSS 0.00102f
C6209 VDD.n297 VSS 0.00187f
C6210 VDD.n298 VSS 0.0025f
C6211 VDD.n299 VSS 0.00259f
C6212 VDD.n300 VSS 0.0084f
C6213 VDD.n301 VSS 0.00101f
C6214 VDD.n302 VSS 0.0011f
C6215 VDD.n303 VSS 0.00285f
C6216 VDD.t345 VSS 0.00131f
C6217 VDD.t344 VSS 0.00537f
C6218 VDD.n304 VSS 0.00793f
C6219 VDD.n305 VSS 0.00102f
C6220 VDD.n306 VSS 0.00188f
C6221 VDD.n307 VSS 0.00289f
C6222 VDD.n308 VSS 0.00285f
C6223 VDD.t135 VSS 0.00537f
C6224 VDD.n309 VSS 0.00537f
C6225 VDD.n310 VSS 0.00101f
C6226 VDD.n311 VSS 0.0014f
C6227 VDD.n312 VSS 0.00285f
C6228 VDD.t683 VSS 0.00537f
C6229 VDD.n313 VSS 0.0049f
C6230 VDD.n314 VSS 0.00101f
C6231 VDD.n315 VSS 0.00172f
C6232 VDD.n316 VSS 0.00285f
C6233 VDD.t559 VSS 0.00992f
C6234 VDD.n317 VSS 0.007f
C6235 VDD.n318 VSS 0.00102f
C6236 VDD.n319 VSS 0.00164f
C6237 VDD.n320 VSS 0.00285f
C6238 VDD.n321 VSS 0.00183f
C6239 VDD.t560 VSS 5.02e-19
C6240 VDD.t494 VSS 5.29e-19
C6241 VDD.n322 VSS 0.0011f
C6242 VDD.n323 VSS 0.00261f
C6243 VDD.n324 VSS 0.00274f
C6244 VDD.n325 VSS 0.00135f
C6245 VDD.n326 VSS 1.26e-19
C6246 VDD.t513 VSS 0.00138f
C6247 VDD.t772 VSS 5.9e-19
C6248 VDD.n327 VSS 0.00258f
C6249 VDD.n328 VSS 2.16e-19
C6250 VDD.n329 VSS 6.27e-19
C6251 VDD.n330 VSS 0.00131f
C6252 VDD.n331 VSS 2.16e-19
C6253 VDD.n332 VSS 0.00359f
C6254 VDD.n333 VSS 4.92e-19
C6255 VDD.n334 VSS 9.75e-19
C6256 VDD.t770 VSS 5.82e-19
C6257 VDD.n335 VSS 0.00292f
C6258 VDD.t492 VSS 0.00175f
C6259 VDD.n336 VSS 0.00161f
C6260 VDD.n337 VSS 2.15e-19
C6261 VDD.n338 VSS 8.62e-19
C6262 VDD.n339 VSS 1.59e-19
C6263 VDD.n340 VSS 2.64e-19
C6264 VDD.n341 VSS 0.00143f
C6265 VDD.t493 VSS 0.0124f
C6266 VDD.t189 VSS 0.00502f
C6267 VDD.n342 VSS 0.0063f
C6268 VDD.n343 VSS 9.56e-19
C6269 VDD.n344 VSS 0.00163f
C6270 VDD.n345 VSS 0.0027f
C6271 VDD.t108 VSS 8.96e-19
C6272 VDD.t562 VSS 0.00201f
C6273 VDD.n346 VSS 0.00323f
C6274 VDD.n347 VSS 0.00423f
C6275 VDD.t107 VSS 0.00525f
C6276 VDD.n348 VSS 0.00572f
C6277 VDD.n349 VSS 0.00101f
C6278 VDD.n350 VSS 9.47e-19
C6279 VDD.n351 VSS 0.00285f
C6280 VDD.t561 VSS 0.00537f
C6281 VDD.n352 VSS 0.00764f
C6282 VDD.n353 VSS 0.00101f
C6283 VDD.n354 VSS 0.00102f
C6284 VDD.n355 VSS 0.00285f
C6285 VDD.n356 VSS 0.0084f
C6286 VDD.n357 VSS 0.00101f
C6287 VDD.n358 VSS 0.00172f
C6288 VDD.n359 VSS 0.00285f
C6289 VDD.t682 VSS 0.00537f
C6290 VDD.n360 VSS 0.0049f
C6291 VDD.n361 VSS 0.00101f
C6292 VDD.n362 VSS 0.00172f
C6293 VDD.n363 VSS 0.00285f
C6294 VDD.t136 VSS 0.00537f
C6295 VDD.n364 VSS 0.00589f
C6296 VDD.n365 VSS 0.00101f
C6297 VDD.n366 VSS 0.00172f
C6298 VDD.n367 VSS 0.00285f
C6299 VDD.t294 VSS 0.00537f
C6300 VDD.n368 VSS 0.0056f
C6301 VDD.n369 VSS 0.00101f
C6302 VDD.n370 VSS 0.00122f
C6303 VDD.n371 VSS 0.00285f
C6304 VDD.t295 VSS 7.06e-19
C6305 VDD.t515 VSS 5.29e-19
C6306 VDD.n372 VSS 0.00129f
C6307 VDD.t514 VSS 0.00537f
C6308 VDD.n373 VSS 0.00706f
C6309 VDD.n374 VSS 0.00102f
C6310 VDD.n375 VSS 0.00189f
C6311 VDD.n376 VSS 0.00234f
C6312 VDD.n377 VSS 0.00285f
C6313 VDD.n378 VSS 0.00618f
C6314 VDD.n379 VSS 0.00101f
C6315 VDD.n380 VSS 0.00152f
C6316 VDD.n381 VSS 0.00285f
C6317 VDD.t445 VSS 0.00537f
C6318 VDD.t105 VSS 0.00537f
C6319 VDD.n382 VSS 0.0042f
C6320 VDD.n383 VSS 0.00101f
C6321 VDD.n384 VSS 0.0016f
C6322 VDD.n385 VSS 0.00285f
C6323 VDD.t106 VSS 0.00243f
C6324 VDD.n386 VSS 0.00251f
C6325 VDD.n387 VSS 0.00817f
C6326 VDD.n388 VSS 9.18e-19
C6327 VDD.n389 VSS 0.00212f
C6328 VDD.n390 VSS 0.00285f
C6329 VDD.n391 VSS 0.00197f
C6330 VDD.n392 VSS 3.68e-19
C6331 VDD.n393 VSS 0.00165f
C6332 VDD.n394 VSS 5e-19
C6333 VDD.n395 VSS 9.34e-20
C6334 VDD.n396 VSS 0.00531f
C6335 VDD.n397 VSS 9.92e-19
C6336 VDD.t12 VSS 0.00543f
C6337 VDD.n398 VSS 0.00192f
C6338 VDD.n399 VSS 5.16e-19
C6339 VDD.n400 VSS 3.9e-19
C6340 VDD.n401 VSS 0.00169f
C6341 VDD.n402 VSS 0.00118f
C6342 VDD.n403 VSS 0.00116f
C6343 VDD.n404 VSS 0.00152f
C6344 VDD.t13 VSS 8.48e-19
C6345 VDD.t293 VSS -4.69e-19
C6346 VDD.n405 VSS 0.00333f
C6347 VDD.n406 VSS 6.2e-19
C6348 VDD.n407 VSS 0.00133f
C6349 VDD.n408 VSS 3.68e-19
C6350 VDD.n409 VSS 4.94e-19
C6351 VDD.n410 VSS 9.34e-20
C6352 VDD.t292 VSS 0.00432f
C6353 VDD.n411 VSS 0.00204f
C6354 VDD.n412 VSS 9.92e-19
C6355 VDD.n413 VSS 0.00362f
C6356 VDD.n414 VSS 5.16e-19
C6357 VDD.n415 VSS 4.33e-20
C6358 VDD.n416 VSS 1.3e-19
C6359 VDD.n417 VSS 2.64e-19
C6360 VDD.n418 VSS 0.00143f
C6361 VDD.n419 VSS 0.00858f
C6362 VDD.n420 VSS 9.12e-19
C6363 VDD.n421 VSS 0.00151f
C6364 VDD.n422 VSS 0.00284f
C6365 VDD.t290 VSS 0.00537f
C6366 VDD.n423 VSS 0.00776f
C6367 VDD.n424 VSS 0.00101f
C6368 VDD.n425 VSS 0.00172f
C6369 VDD.n426 VSS 0.00285f
C6370 VDD.t291 VSS 7.86e-19
C6371 VDD.t5 VSS -2.51e-19
C6372 VDD.n427 VSS 0.00362f
C6373 VDD.n428 VSS 0.00382f
C6374 VDD.t4 VSS 0.00537f
C6375 VDD.n429 VSS 0.00554f
C6376 VDD.n430 VSS 0.00101f
C6377 VDD.n431 VSS 9.18e-19
C6378 VDD.n432 VSS 0.00285f
C6379 VDD.n433 VSS 0.00214f
C6380 VDD.n434 VSS 9.77e-19
C6381 VDD.n435 VSS 0.00101f
C6382 VDD.n436 VSS 0.00817f
C6383 VDD.t652 VSS 0.00537f
C6384 VDD.n437 VSS 0.0049f
C6385 VDD.t420 VSS 0.00437f
C6386 VDD.n438 VSS 0.00101f
C6387 VDD.n439 VSS 0.0014f
C6388 VDD.n440 VSS 0.00187f
C6389 VDD.n441 VSS 0.0025f
C6390 VDD.n442 VSS 0.00259f
C6391 VDD.n443 VSS 0.0084f
C6392 VDD.n444 VSS 0.00101f
C6393 VDD.n445 VSS 0.0011f
C6394 VDD.n446 VSS 0.00285f
C6395 VDD.t566 VSS 0.00131f
C6396 VDD.t565 VSS 0.00537f
C6397 VDD.n447 VSS 0.00793f
C6398 VDD.n448 VSS 0.00102f
C6399 VDD.n449 VSS 0.00188f
C6400 VDD.n450 VSS 0.00289f
C6401 VDD.n451 VSS 0.00285f
C6402 VDD.t650 VSS 0.00537f
C6403 VDD.n452 VSS 0.00537f
C6404 VDD.n453 VSS 0.00101f
C6405 VDD.n454 VSS 0.0014f
C6406 VDD.n455 VSS 0.00285f
C6407 VDD.t199 VSS 0.00537f
C6408 VDD.n456 VSS 0.0049f
C6409 VDD.n457 VSS 0.00101f
C6410 VDD.n458 VSS 0.00172f
C6411 VDD.n459 VSS 0.00285f
C6412 VDD.t725 VSS 0.00992f
C6413 VDD.n460 VSS 0.007f
C6414 VDD.n461 VSS 9.56e-19
C6415 VDD.n462 VSS 0.00164f
C6416 VDD.n463 VSS 0.00285f
C6417 VDD.n464 VSS 0.00183f
C6418 VDD.t726 VSS 5.02e-19
C6419 VDD.t536 VSS 5.29e-19
C6420 VDD.n465 VSS 0.0011f
C6421 VDD.n466 VSS 0.00261f
C6422 VDD.n467 VSS 0.00274f
C6423 VDD.n468 VSS 0.00135f
C6424 VDD.n469 VSS 1.26e-19
C6425 VDD.t495 VSS 0.00138f
C6426 VDD.t754 VSS 5.9e-19
C6427 VDD.n470 VSS 0.00258f
C6428 VDD.n471 VSS 2.16e-19
C6429 VDD.n472 VSS 6.27e-19
C6430 VDD.n473 VSS 0.00131f
C6431 VDD.n474 VSS 2.16e-19
C6432 VDD.n475 VSS 0.00359f
C6433 VDD.n476 VSS 4.92e-19
C6434 VDD.n477 VSS 9.75e-19
C6435 VDD.t755 VSS 5.82e-19
C6436 VDD.n478 VSS 0.00292f
C6437 VDD.t534 VSS 0.00175f
C6438 VDD.n479 VSS 0.00161f
C6439 VDD.n480 VSS 2.15e-19
C6440 VDD.n481 VSS 8.62e-19
C6441 VDD.n482 VSS 1.59e-19
C6442 VDD.n483 VSS 2.64e-19
C6443 VDD.n484 VSS 0.00143f
C6444 VDD.t535 VSS 0.0124f
C6445 VDD.t311 VSS 0.00502f
C6446 VDD.n485 VSS 0.0063f
C6447 VDD.n486 VSS 0.00107f
C6448 VDD.n487 VSS 0.00163f
C6449 VDD.n488 VSS 0.0027f
C6450 VDD.t436 VSS 8.96e-19
C6451 VDD.t724 VSS 0.00201f
C6452 VDD.n489 VSS 0.00323f
C6453 VDD.n490 VSS 0.00423f
C6454 VDD.t435 VSS 0.00525f
C6455 VDD.n491 VSS 0.00572f
C6456 VDD.n492 VSS 0.00101f
C6457 VDD.n493 VSS 9.47e-19
C6458 VDD.n494 VSS 0.00285f
C6459 VDD.t723 VSS 0.00537f
C6460 VDD.n495 VSS 0.00764f
C6461 VDD.n496 VSS 0.00101f
C6462 VDD.n497 VSS 0.00102f
C6463 VDD.n498 VSS 0.00285f
C6464 VDD.n499 VSS 0.0084f
C6465 VDD.n500 VSS 0.00101f
C6466 VDD.n501 VSS 0.00172f
C6467 VDD.n502 VSS 0.00285f
C6468 VDD.t198 VSS 0.00537f
C6469 VDD.n503 VSS 0.0049f
C6470 VDD.n504 VSS 0.00101f
C6471 VDD.n505 VSS 0.00172f
C6472 VDD.n506 VSS 0.00285f
C6473 VDD.t651 VSS 0.00537f
C6474 VDD.n507 VSS 0.00589f
C6475 VDD.n508 VSS 0.00101f
C6476 VDD.n509 VSS 0.00172f
C6477 VDD.n510 VSS 0.00285f
C6478 VDD.t734 VSS 0.00537f
C6479 VDD.n511 VSS 0.0056f
C6480 VDD.n512 VSS 0.00101f
C6481 VDD.n513 VSS 0.00122f
C6482 VDD.n514 VSS 0.00285f
C6483 VDD.t735 VSS 7.06e-19
C6484 VDD.t497 VSS 5.29e-19
C6485 VDD.n515 VSS 0.00129f
C6486 VDD.t496 VSS 0.00537f
C6487 VDD.n516 VSS 0.00706f
C6488 VDD.n517 VSS 0.00102f
C6489 VDD.n518 VSS 0.00189f
C6490 VDD.n519 VSS 0.00234f
C6491 VDD.n520 VSS 0.00285f
C6492 VDD.n521 VSS 0.00618f
C6493 VDD.n522 VSS 0.00101f
C6494 VDD.n523 VSS 0.00152f
C6495 VDD.n524 VSS 0.00285f
C6496 VDD.t476 VSS 0.00537f
C6497 VDD.t433 VSS 0.00537f
C6498 VDD.n525 VSS 0.0042f
C6499 VDD.n526 VSS 0.00101f
C6500 VDD.n527 VSS 0.0016f
C6501 VDD.n528 VSS 0.00285f
C6502 VDD.t434 VSS 0.00243f
C6503 VDD.n529 VSS 0.00251f
C6504 VDD.n530 VSS 0.00916f
C6505 VDD.n531 VSS 0.00101f
C6506 VDD.n532 VSS 0.00249f
C6507 VDD.n533 VSS 0.00285f
C6508 VDD.t29 VSS 0.00437f
C6509 VDD.n534 VSS 0.00723f
C6510 VDD.n535 VSS 9.18e-19
C6511 VDD.n536 VSS 0.00362f
C6512 VDD.n537 VSS 0.00285f
C6513 VDD.n538 VSS 0.00188f
C6514 VDD.t30 VSS 8.48e-19
C6515 VDD.t733 VSS -4.69e-19
C6516 VDD.n539 VSS 0.00333f
C6517 VDD.n540 VSS 6.2e-19
C6518 VDD.n541 VSS 1.08e-19
C6519 VDD.n542 VSS 0.00139f
C6520 VDD.n543 VSS 5e-19
C6521 VDD.n544 VSS 9.34e-20
C6522 VDD.n545 VSS 0.00344f
C6523 VDD.n546 VSS 9.92e-19
C6524 VDD.t732 VSS 0.00537f
C6525 VDD.n547 VSS 0.00222f
C6526 VDD.n548 VSS 5.11e-19
C6527 VDD.n549 VSS 3.9e-19
C6528 VDD.n550 VSS 0.00169f
C6529 VDD.n551 VSS 0.00143f
C6530 VDD.n552 VSS 0.00858f
C6531 VDD.n553 VSS 0.00101f
C6532 VDD.n554 VSS 0.00152f
C6533 VDD.n555 VSS 0.00259f
C6534 VDD.t730 VSS 0.00537f
C6535 VDD.n556 VSS 0.00776f
C6536 VDD.n557 VSS 0.00101f
C6537 VDD.n558 VSS 0.00172f
C6538 VDD.n559 VSS 0.00285f
C6539 VDD.t731 VSS 7.86e-19
C6540 VDD.t626 VSS -2.51e-19
C6541 VDD.n560 VSS 0.00362f
C6542 VDD.n561 VSS 0.00382f
C6543 VDD.t625 VSS 0.00537f
C6544 VDD.n562 VSS 0.00554f
C6545 VDD.n563 VSS 0.00101f
C6546 VDD.n564 VSS 9.18e-19
C6547 VDD.n565 VSS 0.00285f
C6548 VDD.n566 VSS 0.00214f
C6549 VDD.n567 VSS 9.77e-19
C6550 VDD.n568 VSS 0.00101f
C6551 VDD.n569 VSS 0.00817f
C6552 VDD.t204 VSS 0.00537f
C6553 VDD.n570 VSS 0.0049f
C6554 VDD.t288 VSS 0.00437f
C6555 VDD.n571 VSS 0.00101f
C6556 VDD.n572 VSS 0.0014f
C6557 VDD.n573 VSS 0.00187f
C6558 VDD.n574 VSS 0.0025f
C6559 VDD.n575 VSS 0.00259f
C6560 VDD.n576 VSS 0.0084f
C6561 VDD.n577 VSS 0.00101f
C6562 VDD.n578 VSS 0.0011f
C6563 VDD.n579 VSS 0.00285f
C6564 VDD.t266 VSS 0.00131f
C6565 VDD.t265 VSS 0.00537f
C6566 VDD.n580 VSS 0.00793f
C6567 VDD.n581 VSS 0.00102f
C6568 VDD.n582 VSS 0.00188f
C6569 VDD.n583 VSS 0.00289f
C6570 VDD.n584 VSS 0.00285f
C6571 VDD.t206 VSS 0.00537f
C6572 VDD.n585 VSS 0.00537f
C6573 VDD.n586 VSS 0.00101f
C6574 VDD.n587 VSS 0.0014f
C6575 VDD.n588 VSS 0.00285f
C6576 VDD.t148 VSS 0.00537f
C6577 VDD.n589 VSS 0.0049f
C6578 VDD.n590 VSS 0.00101f
C6579 VDD.n591 VSS 0.00172f
C6580 VDD.n592 VSS 0.00285f
C6581 VDD.t41 VSS 0.00992f
C6582 VDD.n593 VSS 0.007f
C6583 VDD.n594 VSS 0.00116f
C6584 VDD.n595 VSS 0.00164f
C6585 VDD.n596 VSS 0.00285f
C6586 VDD.n597 VSS 0.00183f
C6587 VDD.t42 VSS 5.02e-19
C6588 VDD.t527 VSS 5.29e-19
C6589 VDD.n598 VSS 0.0011f
C6590 VDD.n599 VSS 0.00261f
C6591 VDD.n600 VSS 0.00274f
C6592 VDD.n601 VSS 0.00135f
C6593 VDD.n602 VSS 1.26e-19
C6594 VDD.t537 VSS 0.00138f
C6595 VDD.t760 VSS 5.9e-19
C6596 VDD.n603 VSS 0.00258f
C6597 VDD.n604 VSS 2.16e-19
C6598 VDD.n605 VSS 6.27e-19
C6599 VDD.n606 VSS 0.00131f
C6600 VDD.n607 VSS 2.16e-19
C6601 VDD.n608 VSS 0.00359f
C6602 VDD.n609 VSS 4.92e-19
C6603 VDD.n610 VSS 9.75e-19
C6604 VDD.t758 VSS 5.82e-19
C6605 VDD.n611 VSS 0.00292f
C6606 VDD.t525 VSS 0.00175f
C6607 VDD.n612 VSS 0.00161f
C6608 VDD.n613 VSS 2.15e-19
C6609 VDD.n614 VSS 8.62e-19
C6610 VDD.n615 VSS 1.59e-19
C6611 VDD.n616 VSS 2.64e-19
C6612 VDD.n617 VSS 0.00143f
C6613 VDD.t526 VSS 0.0124f
C6614 VDD.t579 VSS 0.00502f
C6615 VDD.n618 VSS 0.0063f
C6616 VDD.n619 VSS 0.00107f
C6617 VDD.n620 VSS 0.00163f
C6618 VDD.n621 VSS 0.0027f
C6619 VDD.t635 VSS 8.96e-19
C6620 VDD.t40 VSS 0.00201f
C6621 VDD.n622 VSS 0.00323f
C6622 VDD.n623 VSS 0.00423f
C6623 VDD.t634 VSS 0.00525f
C6624 VDD.n624 VSS 0.00572f
C6625 VDD.n625 VSS 0.00101f
C6626 VDD.n626 VSS 9.47e-19
C6627 VDD.n627 VSS 0.00285f
C6628 VDD.t39 VSS 0.00537f
C6629 VDD.n628 VSS 0.00764f
C6630 VDD.n629 VSS 0.00101f
C6631 VDD.n630 VSS 0.00102f
C6632 VDD.n631 VSS 0.00285f
C6633 VDD.n632 VSS 0.0084f
C6634 VDD.n633 VSS 0.00101f
C6635 VDD.n634 VSS 0.00172f
C6636 VDD.n635 VSS 0.00285f
C6637 VDD.t149 VSS 0.00537f
C6638 VDD.n636 VSS 0.0049f
C6639 VDD.n637 VSS 0.00101f
C6640 VDD.n638 VSS 0.00172f
C6641 VDD.n639 VSS 0.00285f
C6642 VDD.t207 VSS 0.00537f
C6643 VDD.n640 VSS 0.00589f
C6644 VDD.n641 VSS 0.00101f
C6645 VDD.n642 VSS 0.00172f
C6646 VDD.n643 VSS 0.00285f
C6647 VDD.t80 VSS 0.00537f
C6648 VDD.n644 VSS 0.0056f
C6649 VDD.n645 VSS 0.00101f
C6650 VDD.n646 VSS 0.00122f
C6651 VDD.n647 VSS 0.00285f
C6652 VDD.t81 VSS 7.06e-19
C6653 VDD.t539 VSS 5.29e-19
C6654 VDD.n648 VSS 0.00129f
C6655 VDD.t538 VSS 0.00537f
C6656 VDD.n649 VSS 0.00706f
C6657 VDD.n650 VSS 0.00102f
C6658 VDD.n651 VSS 0.00189f
C6659 VDD.n652 VSS 0.00234f
C6660 VDD.n653 VSS 0.00285f
C6661 VDD.n654 VSS 0.00618f
C6662 VDD.n655 VSS 0.00101f
C6663 VDD.n656 VSS 0.00152f
C6664 VDD.n657 VSS 0.00285f
C6665 VDD.t339 VSS 0.00537f
C6666 VDD.t636 VSS 0.00537f
C6667 VDD.n658 VSS 0.0042f
C6668 VDD.n659 VSS 0.00101f
C6669 VDD.n660 VSS 0.0016f
C6670 VDD.n661 VSS 0.00285f
C6671 VDD.t637 VSS 0.00243f
C6672 VDD.n662 VSS 0.00251f
C6673 VDD.n663 VSS 0.00916f
C6674 VDD.n664 VSS 0.00101f
C6675 VDD.n665 VSS 0.00249f
C6676 VDD.n666 VSS 0.00285f
C6677 VDD.t479 VSS 0.00543f
C6678 VDD.n667 VSS 0.00723f
C6679 VDD.n668 VSS 0.00102f
C6680 VDD.n669 VSS 0.00364f
C6681 VDD.n670 VSS 0.00261f
C6682 VDD.n671 VSS 0.00143f
C6683 VDD.n672 VSS 0.00188f
C6684 VDD.t480 VSS 8.48e-19
C6685 VDD.t83 VSS -4.69e-19
C6686 VDD.n673 VSS 0.00333f
C6687 VDD.n674 VSS 6.2e-19
C6688 VDD.n675 VSS 0.00133f
C6689 VDD.n676 VSS 3.68e-19
C6690 VDD.n677 VSS 4.94e-19
C6691 VDD.n678 VSS 9.34e-20
C6692 VDD.t82 VSS 0.00432f
C6693 VDD.n679 VSS 0.00204f
C6694 VDD.n680 VSS 9.92e-19
C6695 VDD.n681 VSS 0.00362f
C6696 VDD.n682 VSS 5.16e-19
C6697 VDD.n683 VSS 4.33e-20
C6698 VDD.n684 VSS 1.3e-19
C6699 VDD.n685 VSS 2.64e-19
C6700 VDD.n686 VSS 0.00143f
C6701 VDD.n687 VSS 0.00858f
C6702 VDD.n688 VSS 9.12e-19
C6703 VDD.n689 VSS 0.00151f
C6704 VDD.n690 VSS 0.00284f
C6705 VDD.t84 VSS 0.00537f
C6706 VDD.n691 VSS 0.00776f
C6707 VDD.n692 VSS 0.00101f
C6708 VDD.n693 VSS 0.00172f
C6709 VDD.n694 VSS 0.00285f
C6710 VDD.t85 VSS 7.86e-19
C6711 VDD.t191 VSS -2.51e-19
C6712 VDD.n695 VSS 0.00362f
C6713 VDD.n696 VSS 0.00382f
C6714 VDD.t190 VSS 0.00537f
C6715 VDD.n697 VSS 0.00554f
C6716 VDD.n698 VSS 0.00101f
C6717 VDD.n699 VSS 9.18e-19
C6718 VDD.n700 VSS 0.00285f
C6719 VDD.n701 VSS 0.00214f
C6720 VDD.n702 VSS 9.77e-19
C6721 VDD.n703 VSS 0.00101f
C6722 VDD.n704 VSS 0.00817f
C6723 VDD.t6 VSS 0.00537f
C6724 VDD.n705 VSS 0.0049f
C6725 VDD.t10 VSS 0.00437f
C6726 VDD.n706 VSS 0.00101f
C6727 VDD.n707 VSS 0.0014f
C6728 VDD.n708 VSS 0.00187f
C6729 VDD.n709 VSS 0.0025f
C6730 VDD.n710 VSS 0.00259f
C6731 VDD.n711 VSS 0.0084f
C6732 VDD.n712 VSS 0.00101f
C6733 VDD.n713 VSS 0.0011f
C6734 VDD.n714 VSS 0.00285f
C6735 VDD.t69 VSS 0.00131f
C6736 VDD.t68 VSS 0.00537f
C6737 VDD.n715 VSS 0.00793f
C6738 VDD.n716 VSS 0.00102f
C6739 VDD.n717 VSS 0.00188f
C6740 VDD.n718 VSS 0.00289f
C6741 VDD.n719 VSS 0.00285f
C6742 VDD.t8 VSS 0.00537f
C6743 VDD.n720 VSS 0.00537f
C6744 VDD.n721 VSS 0.00101f
C6745 VDD.n722 VSS 0.0014f
C6746 VDD.n723 VSS 0.00285f
C6747 VDD.t297 VSS 0.00537f
C6748 VDD.n724 VSS 0.0049f
C6749 VDD.n725 VSS 0.00101f
C6750 VDD.n726 VSS 0.00172f
C6751 VDD.n727 VSS 0.00285f
C6752 VDD.t64 VSS 0.00992f
C6753 VDD.n728 VSS 0.007f
C6754 VDD.n729 VSS 9.56e-19
C6755 VDD.n730 VSS 0.00164f
C6756 VDD.n731 VSS 0.00285f
C6757 VDD.n732 VSS 0.00183f
C6758 VDD.t65 VSS 5.02e-19
C6759 VDD.t509 VSS 5.29e-19
C6760 VDD.n733 VSS 0.0011f
C6761 VDD.n734 VSS 0.00261f
C6762 VDD.n735 VSS 0.00274f
C6763 VDD.n736 VSS 0.00135f
C6764 VDD.n737 VSS 1.26e-19
C6765 VDD.t528 VSS 0.00138f
C6766 VDD.t762 VSS 5.9e-19
C6767 VDD.n738 VSS 0.00258f
C6768 VDD.n739 VSS 2.16e-19
C6769 VDD.n740 VSS 6.27e-19
C6770 VDD.n741 VSS 0.00131f
C6771 VDD.n742 VSS 2.16e-19
C6772 VDD.n743 VSS 0.00359f
C6773 VDD.n744 VSS 4.92e-19
C6774 VDD.n745 VSS 9.75e-19
C6775 VDD.t764 VSS 5.82e-19
C6776 VDD.n746 VSS 0.00292f
C6777 VDD.t507 VSS 0.00175f
C6778 VDD.n747 VSS 0.00161f
C6779 VDD.n748 VSS 2.15e-19
C6780 VDD.n749 VSS 8.62e-19
C6781 VDD.n750 VSS 1.59e-19
C6782 VDD.n751 VSS 2.64e-19
C6783 VDD.n752 VSS 0.00143f
C6784 VDD.t508 VSS 0.0124f
C6785 VDD.t72 VSS 0.00502f
C6786 VDD.n753 VSS 0.0063f
C6787 VDD.n754 VSS 1e-18
C6788 VDD.n755 VSS 0.00163f
C6789 VDD.n756 VSS 0.0027f
C6790 VDD.t20 VSS 8.96e-19
C6791 VDD.t63 VSS 0.00201f
C6792 VDD.n757 VSS 0.00323f
C6793 VDD.n758 VSS 0.00423f
C6794 VDD.t19 VSS 0.00525f
C6795 VDD.n759 VSS 0.00572f
C6796 VDD.n760 VSS 0.00101f
C6797 VDD.n761 VSS 9.47e-19
C6798 VDD.n762 VSS 0.00285f
C6799 VDD.t62 VSS 0.00537f
C6800 VDD.n763 VSS 0.00764f
C6801 VDD.n764 VSS 0.00101f
C6802 VDD.n765 VSS 0.00102f
C6803 VDD.n766 VSS 0.00285f
C6804 VDD.n767 VSS 0.0084f
C6805 VDD.n768 VSS 0.00101f
C6806 VDD.n769 VSS 0.00172f
C6807 VDD.n770 VSS 0.00285f
C6808 VDD.t298 VSS 0.00537f
C6809 VDD.n771 VSS 0.0049f
C6810 VDD.n772 VSS 0.00101f
C6811 VDD.n773 VSS 0.00172f
C6812 VDD.n774 VSS 0.00285f
C6813 VDD.t9 VSS 0.00537f
C6814 VDD.n775 VSS 0.00589f
C6815 VDD.n776 VSS 0.00101f
C6816 VDD.n777 VSS 0.00172f
C6817 VDD.n778 VSS 0.00285f
C6818 VDD.t713 VSS 0.00537f
C6819 VDD.n779 VSS 0.0056f
C6820 VDD.n780 VSS 0.00101f
C6821 VDD.n781 VSS 0.00122f
C6822 VDD.n782 VSS 0.00285f
C6823 VDD.t714 VSS 7.06e-19
C6824 VDD.t530 VSS 5.29e-19
C6825 VDD.n783 VSS 0.00129f
C6826 VDD.t529 VSS 0.00537f
C6827 VDD.n784 VSS 0.00706f
C6828 VDD.n785 VSS 0.00102f
C6829 VDD.n786 VSS 0.00189f
C6830 VDD.n787 VSS 0.00234f
C6831 VDD.n788 VSS 0.00285f
C6832 VDD.n789 VSS 0.00618f
C6833 VDD.n790 VSS 0.00101f
C6834 VDD.n791 VSS 0.00152f
C6835 VDD.n792 VSS 0.00285f
C6836 VDD.t104 VSS 0.00537f
C6837 VDD.t21 VSS 0.00537f
C6838 VDD.n793 VSS 0.0042f
C6839 VDD.n794 VSS 0.00101f
C6840 VDD.n795 VSS 0.0016f
C6841 VDD.n796 VSS 0.00285f
C6842 VDD.t22 VSS 0.00243f
C6843 VDD.n797 VSS 0.00251f
C6844 VDD.n798 VSS 0.00817f
C6845 VDD.n799 VSS 9.18e-19
C6846 VDD.n800 VSS 0.00212f
C6847 VDD.n801 VSS 0.00285f
C6848 VDD.n802 VSS 0.00197f
C6849 VDD.n803 VSS 3.68e-19
C6850 VDD.n804 VSS 0.0016f
C6851 VDD.n805 VSS 5e-19
C6852 VDD.n806 VSS 9.34e-20
C6853 VDD.n807 VSS 0.00531f
C6854 VDD.n808 VSS 9.92e-19
C6855 VDD.t17 VSS 0.00432f
C6856 VDD.n809 VSS 0.00192f
C6857 VDD.n810 VSS 4.12e-19
C6858 VDD.n811 VSS 3.9e-19
C6859 VDD.n812 VSS 0.00169f
C6860 VDD.n813 VSS 0.00141f
C6861 VDD.n814 VSS 0.00116f
C6862 VDD.n815 VSS 0.00152f
C6863 VDD.t18 VSS 8.48e-19
C6864 VDD.t712 VSS -4.69e-19
C6865 VDD.n816 VSS 0.00333f
C6866 VDD.n817 VSS 6.2e-19
C6867 VDD.n818 VSS 8.66e-20
C6868 VDD.n819 VSS 4.94e-19
C6869 VDD.n820 VSS 9.34e-20
C6870 VDD.n821 VSS 0.00338f
C6871 VDD.n822 VSS 9.92e-19
C6872 VDD.t711 VSS 0.00543f
C6873 VDD.n823 VSS 0.00227f
C6874 VDD.n824 VSS 5.16e-19
C6875 VDD.n825 VSS 4.33e-20
C6876 VDD.n826 VSS 0.0014f
C6877 VDD.n827 VSS 3.68e-19
C6878 VDD.n828 VSS 2.64e-19
C6879 VDD.n829 VSS 0.00143f
C6880 VDD.n830 VSS 0.00858f
C6881 VDD.n831 VSS 0.00102f
C6882 VDD.n832 VSS 0.00153f
C6883 VDD.n833 VSS 0.00261f
C6884 VDD.t715 VSS 0.00537f
C6885 VDD.n834 VSS 0.00776f
C6886 VDD.n835 VSS 0.00101f
C6887 VDD.n836 VSS 0.00172f
C6888 VDD.n837 VSS 0.00285f
C6889 VDD.t716 VSS 7.86e-19
C6890 VDD.t451 VSS -2.51e-19
C6891 VDD.n838 VSS 0.00362f
C6892 VDD.n839 VSS 0.00382f
C6893 VDD.t450 VSS 0.00537f
C6894 VDD.n840 VSS 0.00554f
C6895 VDD.n841 VSS 0.00101f
C6896 VDD.n842 VSS 9.18e-19
C6897 VDD.n843 VSS 0.00285f
C6898 VDD.n844 VSS 0.00214f
C6899 VDD.n845 VSS 9.77e-19
C6900 VDD.n846 VSS 0.00101f
C6901 VDD.n847 VSS 0.00817f
C6902 VDD.t59 VSS 0.00537f
C6903 VDD.n848 VSS 0.0049f
C6904 VDD.t98 VSS 0.00437f
C6905 VDD.n849 VSS 0.00101f
C6906 VDD.n850 VSS 0.0014f
C6907 VDD.n851 VSS 0.00187f
C6908 VDD.n852 VSS 0.0025f
C6909 VDD.n853 VSS 0.00259f
C6910 VDD.n854 VSS 0.0084f
C6911 VDD.n855 VSS 0.00101f
C6912 VDD.n856 VSS 0.0011f
C6913 VDD.n857 VSS 0.00285f
C6914 VDD.t349 VSS 0.00131f
C6915 VDD.t348 VSS 0.00537f
C6916 VDD.n858 VSS 0.00793f
C6917 VDD.n859 VSS 0.00102f
C6918 VDD.n860 VSS 0.00188f
C6919 VDD.n861 VSS 0.00289f
C6920 VDD.n862 VSS 0.00285f
C6921 VDD.t58 VSS 0.00537f
C6922 VDD.n863 VSS 0.00537f
C6923 VDD.n864 VSS 0.00101f
C6924 VDD.n865 VSS 0.0014f
C6925 VDD.n866 VSS 0.00285f
C6926 VDD.t49 VSS 0.00537f
C6927 VDD.n867 VSS 0.0049f
C6928 VDD.n868 VSS 0.00101f
C6929 VDD.n869 VSS 0.00172f
C6930 VDD.n870 VSS 0.00285f
C6931 VDD.t337 VSS 0.00992f
C6932 VDD.n871 VSS 0.007f
C6933 VDD.n872 VSS 9.56e-19
C6934 VDD.n873 VSS 0.00164f
C6935 VDD.n874 VSS 0.00285f
C6936 VDD.n875 VSS 0.00183f
C6937 VDD.t338 VSS 5.02e-19
C6938 VDD.t551 VSS 5.29e-19
C6939 VDD.n876 VSS 0.0011f
C6940 VDD.n877 VSS 0.00261f
C6941 VDD.n878 VSS 0.00274f
C6942 VDD.n879 VSS 0.00135f
C6943 VDD.n880 VSS 1.26e-19
C6944 VDD.t531 VSS 0.00138f
C6945 VDD.t761 VSS 5.9e-19
C6946 VDD.n881 VSS 0.00258f
C6947 VDD.n882 VSS 2.16e-19
C6948 VDD.n883 VSS 6.27e-19
C6949 VDD.n884 VSS 0.00131f
C6950 VDD.n885 VSS 2.16e-19
C6951 VDD.n886 VSS 0.00359f
C6952 VDD.n887 VSS 4.92e-19
C6953 VDD.n888 VSS 9.75e-19
C6954 VDD.t771 VSS 5.82e-19
C6955 VDD.n889 VSS 0.00292f
C6956 VDD.t549 VSS 0.00175f
C6957 VDD.n890 VSS 0.00161f
C6958 VDD.n891 VSS 2.15e-19
C6959 VDD.n892 VSS 8.62e-19
C6960 VDD.n893 VSS 1.59e-19
C6961 VDD.n894 VSS 2.64e-19
C6962 VDD.n895 VSS 0.00143f
C6963 VDD.t550 VSS 0.0124f
C6964 VDD.t481 VSS 0.00502f
C6965 VDD.n896 VSS 0.0063f
C6966 VDD.n897 VSS 9.56e-19
C6967 VDD.n898 VSS 0.00163f
C6968 VDD.n899 VSS 0.0027f
C6969 VDD.t318 VSS 8.96e-19
C6970 VDD.t336 VSS 0.00201f
C6971 VDD.n900 VSS 0.00323f
C6972 VDD.n901 VSS 0.00423f
C6973 VDD.t317 VSS 0.00525f
C6974 VDD.n902 VSS 0.00572f
C6975 VDD.n903 VSS 0.00101f
C6976 VDD.n904 VSS 9.47e-19
C6977 VDD.n905 VSS 0.00285f
C6978 VDD.t335 VSS 0.00537f
C6979 VDD.n906 VSS 0.00764f
C6980 VDD.n907 VSS 0.00101f
C6981 VDD.n908 VSS 0.00102f
C6982 VDD.n909 VSS 0.00285f
C6983 VDD.n910 VSS 0.0084f
C6984 VDD.n911 VSS 0.00101f
C6985 VDD.n912 VSS 0.00172f
C6986 VDD.n913 VSS 0.00285f
C6987 VDD.t48 VSS 0.00537f
C6988 VDD.n914 VSS 0.0049f
C6989 VDD.n915 VSS 0.00101f
C6990 VDD.n916 VSS 0.00172f
C6991 VDD.n917 VSS 0.00285f
C6992 VDD.t61 VSS 0.00537f
C6993 VDD.n918 VSS 0.00589f
C6994 VDD.n919 VSS 0.00101f
C6995 VDD.n920 VSS 0.00172f
C6996 VDD.n921 VSS 0.00285f
C6997 VDD.t181 VSS 0.00537f
C6998 VDD.n922 VSS 0.0056f
C6999 VDD.n923 VSS 0.00101f
C7000 VDD.n924 VSS 0.00122f
C7001 VDD.n925 VSS 0.00285f
C7002 VDD.t182 VSS 7.06e-19
C7003 VDD.t533 VSS 5.29e-19
C7004 VDD.n926 VSS 0.00129f
C7005 VDD.t532 VSS 0.00537f
C7006 VDD.n927 VSS 0.00706f
C7007 VDD.n928 VSS 0.00102f
C7008 VDD.n929 VSS 0.00189f
C7009 VDD.n930 VSS 0.00234f
C7010 VDD.n931 VSS 0.00285f
C7011 VDD.n932 VSS 0.00618f
C7012 VDD.n933 VSS 0.00101f
C7013 VDD.n934 VSS 0.00152f
C7014 VDD.n935 VSS 0.00285f
C7015 VDD.t47 VSS 0.00537f
C7016 VDD.t319 VSS 0.00537f
C7017 VDD.n936 VSS 0.0042f
C7018 VDD.n937 VSS 0.00101f
C7019 VDD.n938 VSS 0.00111f
C7020 VDD.n939 VSS 0.00285f
C7021 VDD.t320 VSS 0.00245f
C7022 VDD.n940 VSS 0.00381f
C7023 VDD.n941 VSS 0.00799f
C7024 VDD.n942 VSS 9.16e-19
C7025 VDD.n943 VSS 0.00132f
C7026 VDD.n944 VSS 4.79e-19
C7027 VDD.n945 VSS 0.00281f
C7028 VDD.n946 VSS 0.00143f
C7029 VDD.n947 VSS 0.00126f
C7030 VDD.n948 VSS 3.71e-19
C7031 VDD.n949 VSS 4.81e-19
C7032 VDD.n950 VSS 9.6e-20
C7033 VDD.n951 VSS 0.00496f
C7034 VDD.n952 VSS 9.92e-19
C7035 VDD.t601 VSS 0.00566f
C7036 VDD.n953 VSS 0.00227f
C7037 VDD.n954 VSS 5.71e-19
C7038 VDD.n955 VSS 1.53e-19
C7039 VDD.n956 VSS 0.00168f
C7040 VDD.n957 VSS 3.71e-19
C7041 VDD.n958 VSS 2.64e-19
C7042 VDD.n959 VSS 0.00119f
C7043 VDD.n960 VSS 0.00121f
C7044 VDD.n961 VSS 0.00159f
C7045 VDD.t602 VSS 8.48e-19
C7046 VDD.t184 VSS -4.69e-19
C7047 VDD.n962 VSS 0.00333f
C7048 VDD.n963 VSS 6.01e-19
C7049 VDD.n964 VSS 0.0013f
C7050 VDD.n965 VSS 3.71e-19
C7051 VDD.n966 VSS 5.03e-19
C7052 VDD.n967 VSS 9.6e-20
C7053 VDD.t183 VSS 0.00426f
C7054 VDD.n968 VSS 0.00198f
C7055 VDD.n969 VSS 9.92e-19
C7056 VDD.n970 VSS 0.00367f
C7057 VDD.n971 VSS 5.54e-19
C7058 VDD.n972 VSS 6.53e-20
C7059 VDD.n973 VSS 1.53e-19
C7060 VDD.n974 VSS 2.64e-19
C7061 VDD.n975 VSS 0.00143f
C7062 VDD.n976 VSS 0.00858f
C7063 VDD.n977 VSS 9.33e-19
C7064 VDD.n978 VSS 0.00153f
C7065 VDD.n979 VSS 0.00282f
C7066 VDD.t179 VSS 0.00537f
C7067 VDD.n980 VSS 0.00776f
C7068 VDD.n981 VSS 0.00104f
C7069 VDD.n982 VSS 0.00175f
C7070 VDD.n983 VSS 0.00285f
C7071 VDD.t180 VSS 7.86e-19
C7072 VDD.t176 VSS -2.51e-19
C7073 VDD.n984 VSS 0.00362f
C7074 VDD.n985 VSS 0.00384f
C7075 VDD.t175 VSS 0.00616f
C7076 VDD.n986 VSS 0.00554f
C7077 VDD.n987 VSS 0.00104f
C7078 VDD.n988 VSS 9.34e-19
C7079 VDD.n989 VSS 0.00285f
C7080 VDD.n990 VSS 0.0129f
C7081 VDD.n991 VSS 0.0017f
C7082 VDD.n992 VSS 0.00214f
C7083 VDD.n993 VSS 0.00285f
C7084 VDD.t111 VSS 5.58e-19
C7085 VDD.t211 VSS 5.58e-19
C7086 VDD.n994 VSS 0.00121f
C7087 VDD.n995 VSS 0.0025f
C7088 VDD.n996 VSS 0.00187f
C7089 VDD.n997 VSS 0.00102f
C7090 VDD.n998 VSS 0.00791f
C7091 VDD.n999 VSS 0.00102f
C7092 VDD.n1000 VSS 0.00188f
C7093 VDD.n1001 VSS 0.00285f
C7094 VDD.n1002 VSS 0.00172f
C7095 VDD.n1003 VSS 0.00101f
C7096 VDD.t50 VSS 0.00535f
C7097 VDD.n1004 VSS 0.00102f
C7098 VDD.n1005 VSS 0.00189f
C7099 VDD.n1006 VSS 0.00285f
C7100 VDD.n1007 VSS 0.00172f
C7101 VDD.n1008 VSS 0.00101f
C7102 VDD.n1009 VSS 0.00762f
C7103 VDD.n1010 VSS 0.00101f
C7104 VDD.t53 VSS 0.00201f
C7105 VDD.t668 VSS 8.96e-19
C7106 VDD.n1011 VSS 0.00323f
C7107 VDD.n1012 VSS 0.00423f
C7108 VDD.n1013 VSS 0.00285f
C7109 VDD.n1014 VSS 0.00172f
C7110 VDD.n1015 VSS 0.00101f
C7111 VDD.n1016 VSS 0.00558f
C7112 VDD.n1017 VSS 0.00101f
C7113 VDD.n1018 VSS 0.00122f
C7114 VDD.n1019 VSS 0.00285f
C7115 VDD.t381 VSS 5.29e-19
C7116 VDD.t645 VSS 7.06e-19
C7117 VDD.n1020 VSS 0.00129f
C7118 VDD.n1021 VSS 0.00102f
C7119 VDD.n1022 VSS 0.0016f
C7120 VDD.n1023 VSS 0.00101f
C7121 VDD.t547 VSS 0.0129f
C7122 VDD.n1024 VSS 0.00199f
C7123 VDD.t666 VSS 0.00243f
C7124 VDD.n1025 VSS 0.00251f
C7125 VDD.n1026 VSS 0.00143f
C7126 VDD.t757 VSS 8.03e-19
C7127 VDD.n1027 VSS 0.0026f
C7128 VDD.t546 VSS 0.00148f
C7129 VDD.n1028 VSS 0.00165f
C7130 VDD.n1029 VSS 0.00285f
C7131 VDD.n1030 VSS 9.18e-19
C7132 VDD.n1031 VSS 0.00101f
C7133 VDD.n1032 VSS 0.00101f
C7134 VDD.n1033 VSS 0.0014f
C7135 VDD.t3 VSS -2.51e-19
C7136 VDD.t649 VSS 7.86e-19
C7137 VDD.n1034 VSS 0.00362f
C7138 VDD.n1035 VSS 0.00382f
C7139 VDD.n1036 VSS 0.00285f
C7140 VDD.t157 VSS 5.58e-19
C7141 VDD.t578 VSS 5.58e-19
C7142 VDD.n1037 VSS 0.00121f
C7143 VDD.n1038 VSS 0.0011f
C7144 VDD.n1039 VSS 0.00101f
C7145 VDD.t66 VSS 0.00535f
C7146 VDD.n1040 VSS 0.00101f
C7147 VDD.t67 VSS 0.00131f
C7148 VDD.n1041 VSS 0.00289f
C7149 VDD.n1042 VSS 0.00172f
C7150 VDD.n1043 VSS 0.00285f
C7151 VDD.t203 VSS 5.29e-19
C7152 VDD.t193 VSS 5.02e-19
C7153 VDD.n1044 VSS 0.0011f
C7154 VDD.n1045 VSS 0.00257f
C7155 VDD.n1046 VSS 0.00189f
C7156 VDD.n1047 VSS 0.00102f
C7157 VDD.n1048 VSS 0.00101f
C7158 VDD.n1049 VSS 0.00547f
C7159 VDD.n1050 VSS 0.00101f
C7160 VDD.n1051 VSS 0.00172f
C7161 VDD.n1052 VSS 0.00285f
C7162 VDD.t195 VSS 0.00201f
C7163 VDD.t328 VSS 8.96e-19
C7164 VDD.n1053 VSS 0.00323f
C7165 VDD.n1054 VSS 0.00423f
C7166 VDD.n1055 VSS 0.00101f
C7167 VDD.t423 VSS 0.00535f
C7168 VDD.n1056 VSS 0.00101f
C7169 VDD.n1057 VSS 0.00172f
C7170 VDD.n1058 VSS 0.00102f
C7171 VDD.n1059 VSS 0.00285f
C7172 VDD.n1060 VSS 0.00122f
C7173 VDD.n1061 VSS 0.00101f
C7174 VDD.t490 VSS 0.00535f
C7175 VDD.n1062 VSS 0.00101f
C7176 VDD.t491 VSS 5.29e-19
C7177 VDD.t570 VSS 7.06e-19
C7178 VDD.n1063 VSS 0.00129f
C7179 VDD.n1064 VSS 0.00234f
C7180 VDD.n1065 VSS 0.0016f
C7181 VDD.n1066 VSS 0.00143f
C7182 VDD.n1067 VSS 0.00199f
C7183 VDD.t330 VSS 0.00243f
C7184 VDD.n1068 VSS 0.00251f
C7185 VDD.n1069 VSS 0.00774f
C7186 VDD.n1070 VSS 0.00101f
C7187 VDD.n1071 VSS 0.00172f
C7188 VDD.n1072 VSS 0.00173f
C7189 VDD.n1073 VSS 0.00214f
C7190 VDD.t656 VSS -2.51e-19
C7191 VDD.t568 VSS 7.86e-19
C7192 VDD.n1074 VSS 0.00362f
C7193 VDD.n1075 VSS 0.00382f
C7194 VDD.n1076 VSS 0.00101f
C7195 VDD.t274 VSS 0.00535f
C7196 VDD.n1077 VSS 0.00102f
C7197 VDD.n1078 VSS 0.00187f
C7198 VDD.n1079 VSS 0.00167f
C7199 VDD.n1080 VSS 0.00285f
C7200 VDD.t264 VSS 0.00131f
C7201 VDD.n1081 VSS 0.00289f
C7202 VDD.n1082 VSS 0.00188f
C7203 VDD.n1083 VSS 0.00102f
C7204 VDD.t116 VSS 0.00535f
C7205 VDD.n1084 VSS 0.00101f
C7206 VDD.n1085 VSS 0.00172f
C7207 VDD.n1086 VSS 0.00285f
C7208 VDD.t32 VSS 5.29e-19
C7209 VDD.t457 VSS 5.02e-19
C7210 VDD.n1087 VSS 0.0011f
C7211 VDD.n1088 VSS 0.00257f
C7212 VDD.n1089 VSS 0.00189f
C7213 VDD.n1090 VSS 0.00102f
C7214 VDD.n1091 VSS 0.00547f
C7215 VDD.n1092 VSS 0.00101f
C7216 VDD.n1093 VSS 0.00172f
C7217 VDD.n1094 VSS 0.00285f
C7218 VDD.t459 VSS 0.00201f
C7219 VDD.t722 VSS 8.96e-19
C7220 VDD.n1095 VSS 0.00323f
C7221 VDD.n1096 VSS 0.00423f
C7222 VDD.n1097 VSS 0.00101f
C7223 VDD.t702 VSS 0.00535f
C7224 VDD.n1098 VSS 0.00101f
C7225 VDD.n1099 VSS 0.00172f
C7226 VDD.n1100 VSS 0.00102f
C7227 VDD.n1101 VSS 0.00285f
C7228 VDD.n1102 VSS 0.00122f
C7229 VDD.n1103 VSS 0.00101f
C7230 VDD.t146 VSS 0.00535f
C7231 VDD.n1104 VSS 0.00101f
C7232 VDD.t147 VSS 5.29e-19
C7233 VDD.t643 VSS 7.06e-19
C7234 VDD.n1105 VSS 0.00129f
C7235 VDD.n1106 VSS 0.00234f
C7236 VDD.n1107 VSS 0.0016f
C7237 VDD.n1108 VSS 0.00143f
C7238 VDD.n1109 VSS 0.00199f
C7239 VDD.t720 VSS 0.00243f
C7240 VDD.n1110 VSS 0.00251f
C7241 VDD.n1111 VSS 0.00774f
C7242 VDD.n1112 VSS 0.00101f
C7243 VDD.n1113 VSS 0.00172f
C7244 VDD.n1114 VSS 0.00173f
C7245 VDD.n1115 VSS 0.00214f
C7246 VDD.t752 VSS -2.51e-19
C7247 VDD.t641 VSS 7.86e-19
C7248 VDD.n1116 VSS 0.00362f
C7249 VDD.n1117 VSS 0.00382f
C7250 VDD.n1118 VSS 0.00101f
C7251 VDD.t200 VSS 0.00535f
C7252 VDD.n1119 VSS 0.00102f
C7253 VDD.n1120 VSS 0.00187f
C7254 VDD.n1121 VSS 0.00167f
C7255 VDD.n1122 VSS 0.00285f
C7256 VDD.t564 VSS 0.00131f
C7257 VDD.n1123 VSS 0.00289f
C7258 VDD.n1124 VSS 0.00188f
C7259 VDD.n1125 VSS 0.00102f
C7260 VDD.t141 VSS 0.00535f
C7261 VDD.n1126 VSS 0.00101f
C7262 VDD.n1127 VSS 0.00172f
C7263 VDD.n1128 VSS 0.00285f
C7264 VDD.t89 VSS 5.29e-19
C7265 VDD.t334 VSS 5.02e-19
C7266 VDD.n1129 VSS 0.0011f
C7267 VDD.n1130 VSS 0.00257f
C7268 VDD.n1131 VSS 0.00189f
C7269 VDD.n1132 VSS 0.00102f
C7270 VDD.n1133 VSS 0.00547f
C7271 VDD.n1134 VSS 0.00101f
C7272 VDD.n1135 VSS 0.00172f
C7273 VDD.n1136 VSS 0.00285f
C7274 VDD.t332 VSS 0.00201f
C7275 VDD.t674 VSS 8.96e-19
C7276 VDD.n1137 VSS 0.00323f
C7277 VDD.n1138 VSS 0.00423f
C7278 VDD.n1139 VSS 0.00101f
C7279 VDD.t96 VSS 0.00535f
C7280 VDD.n1140 VSS 0.00101f
C7281 VDD.n1141 VSS 0.00172f
C7282 VDD.n1142 VSS 0.00102f
C7283 VDD.n1143 VSS 0.00285f
C7284 VDD.n1144 VSS 0.00122f
C7285 VDD.n1145 VSS 0.00101f
C7286 VDD.t144 VSS 0.00535f
C7287 VDD.n1146 VSS 0.00101f
C7288 VDD.t145 VSS 5.29e-19
C7289 VDD.t622 VSS 7.06e-19
C7290 VDD.n1147 VSS 0.00129f
C7291 VDD.n1148 VSS 0.00234f
C7292 VDD.n1149 VSS 0.0016f
C7293 VDD.n1150 VSS 0.00143f
C7294 VDD.n1151 VSS 0.00199f
C7295 VDD.t676 VSS 0.00243f
C7296 VDD.n1152 VSS 0.00251f
C7297 VDD.n1153 VSS 0.00774f
C7298 VDD.n1154 VSS 0.00101f
C7299 VDD.n1155 VSS 0.00172f
C7300 VDD.n1156 VSS 0.00173f
C7301 VDD.n1157 VSS 0.00214f
C7302 VDD.t377 VSS -2.51e-19
C7303 VDD.t620 VSS 7.86e-19
C7304 VDD.n1158 VSS 0.00362f
C7305 VDD.n1159 VSS 0.00382f
C7306 VDD.n1160 VSS 0.00101f
C7307 VDD.t663 VSS 0.00535f
C7308 VDD.n1161 VSS 0.00102f
C7309 VDD.n1162 VSS 0.00187f
C7310 VDD.n1163 VSS 0.00167f
C7311 VDD.n1164 VSS 0.00285f
C7312 VDD.t343 VSS 0.00131f
C7313 VDD.n1165 VSS 0.00289f
C7314 VDD.n1166 VSS 0.00188f
C7315 VDD.n1167 VSS 0.00102f
C7316 VDD.t326 VSS 0.00535f
C7317 VDD.n1168 VSS 0.00101f
C7318 VDD.n1169 VSS 0.00172f
C7319 VDD.n1170 VSS 0.00285f
C7320 VDD.t629 VSS 5.29e-19
C7321 VDD.t708 VSS 5.02e-19
C7322 VDD.n1171 VSS 0.0011f
C7323 VDD.n1172 VSS 0.00257f
C7324 VDD.n1173 VSS 0.00189f
C7325 VDD.n1174 VSS 0.00102f
C7326 VDD.n1175 VSS 0.00547f
C7327 VDD.n1176 VSS 0.00101f
C7328 VDD.n1177 VSS 0.00172f
C7329 VDD.n1178 VSS 0.00285f
C7330 VDD.t706 VSS 0.00201f
C7331 VDD.t574 VSS 8.96e-19
C7332 VDD.n1179 VSS 0.00323f
C7333 VDD.n1180 VSS 0.00423f
C7334 VDD.n1181 VSS 0.00101f
C7335 VDD.t186 VSS 0.00535f
C7336 VDD.n1182 VSS 0.00101f
C7337 VDD.n1183 VSS 0.00172f
C7338 VDD.n1184 VSS 0.00102f
C7339 VDD.n1185 VSS 0.00285f
C7340 VDD.n1186 VSS 0.00122f
C7341 VDD.n1187 VSS 0.00101f
C7342 VDD.t90 VSS 0.00535f
C7343 VDD.n1188 VSS 0.00101f
C7344 VDD.t91 VSS 5.29e-19
C7345 VDD.t304 VSS 7.06e-19
C7346 VDD.n1189 VSS 0.00129f
C7347 VDD.n1190 VSS 0.00234f
C7348 VDD.n1191 VSS 0.0016f
C7349 VDD.n1192 VSS 0.00143f
C7350 VDD.n1193 VSS 0.00199f
C7351 VDD.t576 VSS 0.00243f
C7352 VDD.n1194 VSS 0.00251f
C7353 VDD.n1195 VSS 0.00774f
C7354 VDD.n1196 VSS 0.00101f
C7355 VDD.n1197 VSS 0.00172f
C7356 VDD.n1198 VSS 0.00173f
C7357 VDD.n1199 VSS 0.00214f
C7358 VDD.t718 VSS -2.51e-19
C7359 VDD.t308 VSS 7.86e-19
C7360 VDD.n1200 VSS 0.00362f
C7361 VDD.n1201 VSS 0.00382f
C7362 VDD.n1202 VSS 0.00101f
C7363 VDD.t669 VSS 0.00535f
C7364 VDD.n1203 VSS 0.00102f
C7365 VDD.n1204 VSS 0.00187f
C7366 VDD.n1205 VSS 0.00167f
C7367 VDD.n1206 VSS 0.00285f
C7368 VDD.t131 VSS 0.00131f
C7369 VDD.n1207 VSS 0.00289f
C7370 VDD.n1208 VSS 0.00188f
C7371 VDD.n1209 VSS 0.00102f
C7372 VDD.t580 VSS 0.00535f
C7373 VDD.n1210 VSS 0.00101f
C7374 VDD.n1211 VSS 0.00172f
C7375 VDD.n1212 VSS 0.00285f
C7376 VDD.t36 VSS 5.29e-19
C7377 VDD.t254 VSS 5.02e-19
C7378 VDD.n1213 VSS 0.0011f
C7379 VDD.n1214 VSS 0.00257f
C7380 VDD.n1215 VSS 0.00189f
C7381 VDD.n1216 VSS 0.00102f
C7382 VDD.n1217 VSS 0.00547f
C7383 VDD.n1218 VSS 0.00101f
C7384 VDD.n1219 VSS 0.00172f
C7385 VDD.n1220 VSS 0.00285f
C7386 VDD.t252 VSS 0.00201f
C7387 VDD.t737 VSS 8.96e-19
C7388 VDD.n1221 VSS 0.00323f
C7389 VDD.n1222 VSS 0.00423f
C7390 VDD.n1223 VSS 0.00101f
C7391 VDD.t729 VSS 0.00535f
C7392 VDD.n1224 VSS 0.00101f
C7393 VDD.n1225 VSS 0.00172f
C7394 VDD.n1226 VSS 0.00102f
C7395 VDD.n1227 VSS 0.00285f
C7396 VDD.n1228 VSS 0.00122f
C7397 VDD.n1229 VSS 0.00101f
C7398 VDD.t596 VSS 0.00535f
C7399 VDD.n1230 VSS 0.00101f
C7400 VDD.t597 VSS 5.29e-19
C7401 VDD.t258 VSS 7.06e-19
C7402 VDD.n1231 VSS 0.00129f
C7403 VDD.n1232 VSS 0.00234f
C7404 VDD.n1233 VSS 0.0016f
C7405 VDD.n1234 VSS 0.00143f
C7406 VDD.n1235 VSS 0.00199f
C7407 VDD.t739 VSS 0.00243f
C7408 VDD.n1236 VSS 0.00251f
C7409 VDD.n1237 VSS 0.00774f
C7410 VDD.n1238 VSS 0.00101f
C7411 VDD.n1239 VSS 0.00172f
C7412 VDD.n1240 VSS 0.00173f
C7413 VDD.n1241 VSS 0.00214f
C7414 VDD.t310 VSS -2.51e-19
C7415 VDD.t262 VSS 7.86e-19
C7416 VDD.n1242 VSS 0.00362f
C7417 VDD.n1243 VSS 0.00382f
C7418 VDD.n1244 VSS 0.00101f
C7419 VDD.t418 VSS 0.00535f
C7420 VDD.n1245 VSS 0.00102f
C7421 VDD.n1246 VSS 0.00187f
C7422 VDD.n1247 VSS 0.00167f
C7423 VDD.n1248 VSS 0.00285f
C7424 VDD.t593 VSS 0.00131f
C7425 VDD.n1249 VSS 0.00289f
C7426 VDD.n1250 VSS 0.00188f
C7427 VDD.n1251 VSS 0.00102f
C7428 VDD.t129 VSS 0.00535f
C7429 VDD.n1252 VSS 0.00101f
C7430 VDD.n1253 VSS 0.00172f
C7431 VDD.n1254 VSS 0.00285f
C7432 VDD.t600 VSS 5.29e-19
C7433 VDD.t371 VSS 5.02e-19
C7434 VDD.n1255 VSS 0.0011f
C7435 VDD.n1256 VSS 0.00257f
C7436 VDD.n1257 VSS 0.00189f
C7437 VDD.n1258 VSS 0.00102f
C7438 VDD.n1259 VSS 0.00547f
C7439 VDD.n1260 VSS 0.00101f
C7440 VDD.n1261 VSS 0.00172f
C7441 VDD.n1262 VSS 0.00285f
C7442 VDD.t373 VSS 0.00201f
C7443 VDD.t55 VSS 8.96e-19
C7444 VDD.n1263 VSS 0.00323f
C7445 VDD.n1264 VSS 0.00423f
C7446 VDD.n1265 VSS 0.00101f
C7447 VDD.t741 VSS 0.00535f
C7448 VDD.n1266 VSS 0.00101f
C7449 VDD.n1267 VSS 0.00172f
C7450 VDD.n1268 VSS 0.00102f
C7451 VDD.n1269 VSS 0.00285f
C7452 VDD.n1270 VSS 0.00122f
C7453 VDD.n1271 VSS 0.00101f
C7454 VDD.t630 VSS 0.00535f
C7455 VDD.n1272 VSS 0.00101f
C7456 VDD.t631 VSS 5.29e-19
C7457 VDD.t166 VSS 7.06e-19
C7458 VDD.n1273 VSS 0.00129f
C7459 VDD.n1274 VSS 0.00234f
C7460 VDD.n1275 VSS 0.0016f
C7461 VDD.n1276 VSS 0.00143f
C7462 VDD.n1277 VSS 0.00199f
C7463 VDD.t57 VSS 0.00243f
C7464 VDD.n1278 VSS 0.00251f
C7465 VDD.n1279 VSS 0.00774f
C7466 VDD.n1280 VSS 0.00101f
C7467 VDD.n1281 VSS 0.00172f
C7468 VDD.n1282 VSS 0.00173f
C7469 VDD.n1283 VSS 0.00182f
C7470 VDD.t604 VSS -2.51e-19
C7471 VDD.t164 VSS 7.86e-19
C7472 VDD.n1284 VSS 0.00362f
C7473 VDD.n1285 VSS 0.00382f
C7474 VDD.n1286 VSS 0.0128f
C7475 VDD.t603 VSS 0.00614f
C7476 VDD.t163 VSS 0.00535f
C7477 VDD.n1287 VSS 0.00553f
C7478 VDD.n1288 VSS 0.00101f
C7479 VDD.n1289 VSS 9.18e-19
C7480 VDD.n1290 VSS 0.00674f
C7481 VDD.n1291 VSS 0.00285f
C7482 VDD.n1292 VSS 2.64e-19
C7483 VDD.t768 VSS 8.03e-19
C7484 VDD.n1293 VSS 0.0026f
C7485 VDD.t510 VSS 0.00148f
C7486 VDD.t168 VSS -4.69e-19
C7487 VDD.t512 VSS 8.48e-19
C7488 VDD.n1294 VSS 0.00333f
C7489 VDD.n1295 VSS 0.00185f
C7490 VDD.n1296 VSS 0.00315f
C7491 VDD.n1297 VSS 3.68e-19
C7492 VDD.n1298 VSS 6.99e-19
C7493 VDD.n1299 VSS 0.00141f
C7494 VDD.n1300 VSS 0.0026f
C7495 VDD.n1301 VSS 0.00285f
C7496 VDD.n1302 VSS 0.00165f
C7497 VDD.n1303 VSS 6.26e-19
C7498 VDD.n1304 VSS 0.00855f
C7499 VDD.t167 VSS 0.00884f
C7500 VDD.t511 VSS 0.0129f
C7501 VDD.n1305 VSS 0.011f
C7502 VDD.t56 VSS 0.00535f
C7503 VDD.n1306 VSS 0.00617f
C7504 VDD.t710 VSS 0.00535f
C7505 VDD.n1307 VSS 0.00419f
C7506 VDD.n1308 VSS 0.00101f
C7507 VDD.n1309 VSS 7.23e-19
C7508 VDD.n1310 VSS 0.00247f
C7509 VDD.n1311 VSS 0.00284f
C7510 VDD.n1312 VSS 0.00285f
C7511 VDD.n1313 VSS 0.00285f
C7512 VDD.n1314 VSS 0.00285f
C7513 VDD.n1315 VSS 0.00152f
C7514 VDD.n1316 VSS 0.00189f
C7515 VDD.n1317 VSS 0.00102f
C7516 VDD.n1318 VSS 0.00704f
C7517 VDD.t165 VSS 0.00535f
C7518 VDD.n1319 VSS 0.00558f
C7519 VDD.n1320 VSS 0.00489f
C7520 VDD.t126 VSS 0.00535f
C7521 VDD.n1321 VSS 0.00588f
C7522 VDD.n1322 VSS 0.00101f
C7523 VDD.n1323 VSS 0.00172f
C7524 VDD.n1324 VSS 0.00285f
C7525 VDD.n1325 VSS 0.00285f
C7526 VDD.n1326 VSS 0.00285f
C7527 VDD.n1327 VSS 0.00172f
C7528 VDD.n1328 VSS 0.00101f
C7529 VDD.n1329 VSS 0.00838f
C7530 VDD.t372 VSS 0.00535f
C7531 VDD.n1330 VSS 0.00762f
C7532 VDD.t215 VSS 0.005f
C7533 VDD.t54 VSS 0.00524f
C7534 VDD.n1331 VSS 0.0057f
C7535 VDD.n1332 VSS 0.00101f
C7536 VDD.n1333 VSS 9.47e-19
C7537 VDD.n1334 VSS 0.00285f
C7538 VDD.n1335 VSS 0.00285f
C7539 VDD.n1336 VSS 0.00285f
C7540 VDD.n1337 VSS 0.0011f
C7541 VDD.n1338 VSS 0.00101f
C7542 VDD.n1339 VSS 0.00617f
C7543 VDD.t599 VSS 0.00535f
C7544 VDD.n1340 VSS 0.00617f
C7545 VDD.t370 VSS 0.00535f
C7546 VDD.n1341 VSS 0.00489f
C7547 VDD.t740 VSS 0.00535f
C7548 VDD.n1342 VSS 0.00698f
C7549 VDD.n1343 VSS 0.00101f
C7550 VDD.n1344 VSS 0.00164f
C7551 VDD.n1345 VSS 0.00285f
C7552 VDD.n1346 VSS 0.00285f
C7553 VDD.n1347 VSS 0.00285f
C7554 VDD.n1348 VSS 0.0014f
C7555 VDD.n1349 VSS 0.00101f
C7556 VDD.n1350 VSS 0.00535f
C7557 VDD.t592 VSS 0.00535f
C7558 VDD.n1351 VSS 0.00791f
C7559 VDD.n1352 VSS 0.00489f
C7560 VDD.t127 VSS 0.00535f
C7561 VDD.n1353 VSS 0.00838f
C7562 VDD.n1354 VSS 0.00101f
C7563 VDD.n1355 VSS 0.0011f
C7564 VDD.n1356 VSS 0.00285f
C7565 VDD.t128 VSS 5.58e-19
C7566 VDD.t419 VSS 5.58e-19
C7567 VDD.n1357 VSS 0.00121f
C7568 VDD.n1358 VSS 0.0025f
C7569 VDD.n1359 VSS 0.00285f
C7570 VDD.n1360 VSS 0.00169f
C7571 VDD.n1361 VSS 0.0014f
C7572 VDD.n1362 VSS 0.00101f
C7573 VDD.n1363 VSS 0.00716f
C7574 VDD.t309 VSS 0.00535f
C7575 VDD.t261 VSS 0.00535f
C7576 VDD.n1364 VSS 0.00553f
C7577 VDD.n1365 VSS 0.00101f
C7578 VDD.n1366 VSS 9.18e-19
C7579 VDD.n1367 VSS 0.00285f
C7580 VDD.n1368 VSS 0.00285f
C7581 VDD.n1369 VSS 2.64e-19
C7582 VDD.t773 VSS 8.03e-19
C7583 VDD.n1370 VSS 0.0026f
C7584 VDD.t498 VSS 0.00148f
C7585 VDD.t260 VSS -4.69e-19
C7586 VDD.t500 VSS 8.48e-19
C7587 VDD.n1371 VSS 0.00333f
C7588 VDD.n1372 VSS 0.00189f
C7589 VDD.n1373 VSS 0.00328f
C7590 VDD.n1374 VSS 3.68e-19
C7591 VDD.n1375 VSS 7.03e-19
C7592 VDD.n1376 VSS 0.00143f
C7593 VDD.n1377 VSS 0.00261f
C7594 VDD.n1378 VSS 0.00285f
C7595 VDD.n1379 VSS 0.00165f
C7596 VDD.n1380 VSS 6.26e-19
C7597 VDD.n1381 VSS 0.00855f
C7598 VDD.t259 VSS 0.00884f
C7599 VDD.t499 VSS 0.0129f
C7600 VDD.n1382 VSS 0.011f
C7601 VDD.t738 VSS 0.00535f
C7602 VDD.n1383 VSS 0.00617f
C7603 VDD.t248 VSS 0.00535f
C7604 VDD.n1384 VSS 0.00419f
C7605 VDD.n1385 VSS 0.00101f
C7606 VDD.n1386 VSS 7.23e-19
C7607 VDD.n1387 VSS 0.00247f
C7608 VDD.n1388 VSS 0.00284f
C7609 VDD.n1389 VSS 0.00285f
C7610 VDD.n1390 VSS 0.00285f
C7611 VDD.n1391 VSS 0.00285f
C7612 VDD.n1392 VSS 0.00152f
C7613 VDD.n1393 VSS 0.00189f
C7614 VDD.n1394 VSS 0.00102f
C7615 VDD.n1395 VSS 0.00704f
C7616 VDD.t257 VSS 0.00535f
C7617 VDD.n1396 VSS 0.00558f
C7618 VDD.n1397 VSS 0.00489f
C7619 VDD.t583 VSS 0.00535f
C7620 VDD.n1398 VSS 0.00588f
C7621 VDD.n1399 VSS 0.00101f
C7622 VDD.n1400 VSS 0.00172f
C7623 VDD.n1401 VSS 0.00285f
C7624 VDD.n1402 VSS 0.00285f
C7625 VDD.n1403 VSS 0.00285f
C7626 VDD.n1404 VSS 0.00172f
C7627 VDD.n1405 VSS 0.00101f
C7628 VDD.n1406 VSS 0.00838f
C7629 VDD.t251 VSS 0.00535f
C7630 VDD.n1407 VSS 0.00762f
C7631 VDD.t139 VSS 0.005f
C7632 VDD.t736 VSS 0.00524f
C7633 VDD.n1408 VSS 0.0057f
C7634 VDD.n1409 VSS 0.00101f
C7635 VDD.n1410 VSS 9.47e-19
C7636 VDD.n1411 VSS 0.00285f
C7637 VDD.n1412 VSS 0.00285f
C7638 VDD.n1413 VSS 0.00285f
C7639 VDD.n1414 VSS 0.0011f
C7640 VDD.n1415 VSS 0.00101f
C7641 VDD.n1416 VSS 0.00617f
C7642 VDD.t35 VSS 0.00535f
C7643 VDD.n1417 VSS 0.00617f
C7644 VDD.t253 VSS 0.00535f
C7645 VDD.n1418 VSS 0.00489f
C7646 VDD.t728 VSS 0.00535f
C7647 VDD.n1419 VSS 0.00698f
C7648 VDD.n1420 VSS 0.00101f
C7649 VDD.n1421 VSS 0.00164f
C7650 VDD.n1422 VSS 0.00285f
C7651 VDD.n1423 VSS 0.00285f
C7652 VDD.n1424 VSS 0.00285f
C7653 VDD.n1425 VSS 0.0014f
C7654 VDD.n1426 VSS 0.00101f
C7655 VDD.n1427 VSS 0.00535f
C7656 VDD.t130 VSS 0.00535f
C7657 VDD.n1428 VSS 0.00791f
C7658 VDD.n1429 VSS 0.00489f
C7659 VDD.t581 VSS 0.00535f
C7660 VDD.n1430 VSS 0.00838f
C7661 VDD.n1431 VSS 0.00101f
C7662 VDD.n1432 VSS 0.0011f
C7663 VDD.n1433 VSS 0.00285f
C7664 VDD.t582 VSS 5.58e-19
C7665 VDD.t670 VSS 5.58e-19
C7666 VDD.n1434 VSS 0.00121f
C7667 VDD.n1435 VSS 0.0025f
C7668 VDD.n1436 VSS 0.00285f
C7669 VDD.n1437 VSS 0.00169f
C7670 VDD.n1438 VSS 0.0014f
C7671 VDD.n1439 VSS 0.00101f
C7672 VDD.n1440 VSS 0.00716f
C7673 VDD.t717 VSS 0.00535f
C7674 VDD.t307 VSS 0.00535f
C7675 VDD.n1441 VSS 0.00553f
C7676 VDD.n1442 VSS 0.00101f
C7677 VDD.n1443 VSS 9.18e-19
C7678 VDD.n1444 VSS 0.00285f
C7679 VDD.n1445 VSS 0.00285f
C7680 VDD.n1446 VSS 2.64e-19
C7681 VDD.t753 VSS 8.03e-19
C7682 VDD.n1447 VSS 0.0026f
C7683 VDD.t552 VSS 0.00148f
C7684 VDD.t306 VSS -4.69e-19
C7685 VDD.t554 VSS 8.48e-19
C7686 VDD.n1448 VSS 0.00333f
C7687 VDD.n1449 VSS 0.00189f
C7688 VDD.n1450 VSS 0.00329f
C7689 VDD.n1451 VSS 3.68e-19
C7690 VDD.n1452 VSS 7.03e-19
C7691 VDD.n1453 VSS 0.00143f
C7692 VDD.n1454 VSS 0.00261f
C7693 VDD.n1455 VSS 0.00285f
C7694 VDD.n1456 VSS 0.00165f
C7695 VDD.n1457 VSS 6.26e-19
C7696 VDD.n1458 VSS 0.00855f
C7697 VDD.t305 VSS 0.00884f
C7698 VDD.t553 VSS 0.0129f
C7699 VDD.n1459 VSS 0.011f
C7700 VDD.t575 VSS 0.00535f
C7701 VDD.n1460 VSS 0.00617f
C7702 VDD.t727 VSS 0.00535f
C7703 VDD.n1461 VSS 0.00419f
C7704 VDD.n1462 VSS 0.00101f
C7705 VDD.n1463 VSS 7.23e-19
C7706 VDD.n1464 VSS 0.00247f
C7707 VDD.n1465 VSS 0.00284f
C7708 VDD.n1466 VSS 0.00285f
C7709 VDD.n1467 VSS 0.00285f
C7710 VDD.n1468 VSS 0.00285f
C7711 VDD.n1469 VSS 0.00152f
C7712 VDD.n1470 VSS 0.00189f
C7713 VDD.n1471 VSS 0.00102f
C7714 VDD.n1472 VSS 0.00704f
C7715 VDD.t303 VSS 0.00535f
C7716 VDD.n1473 VSS 0.00558f
C7717 VDD.n1474 VSS 0.00489f
C7718 VDD.t323 VSS 0.00535f
C7719 VDD.n1475 VSS 0.00588f
C7720 VDD.n1476 VSS 0.00101f
C7721 VDD.n1477 VSS 0.00172f
C7722 VDD.n1478 VSS 0.00285f
C7723 VDD.n1479 VSS 0.00285f
C7724 VDD.n1480 VSS 0.00285f
C7725 VDD.n1481 VSS 0.00172f
C7726 VDD.n1482 VSS 0.00101f
C7727 VDD.n1483 VSS 0.00838f
C7728 VDD.t705 VSS 0.00535f
C7729 VDD.n1484 VSS 0.00762f
C7730 VDD.t150 VSS 0.005f
C7731 VDD.t573 VSS 0.00524f
C7732 VDD.n1485 VSS 0.0057f
C7733 VDD.n1486 VSS 0.00101f
C7734 VDD.n1487 VSS 9.47e-19
C7735 VDD.n1488 VSS 0.00285f
C7736 VDD.n1489 VSS 0.00285f
C7737 VDD.n1490 VSS 0.00285f
C7738 VDD.n1491 VSS 0.0011f
C7739 VDD.n1492 VSS 0.00101f
C7740 VDD.n1493 VSS 0.00617f
C7741 VDD.t628 VSS 0.00535f
C7742 VDD.n1494 VSS 0.00617f
C7743 VDD.t707 VSS 0.00535f
C7744 VDD.n1495 VSS 0.00489f
C7745 VDD.t185 VSS 0.00535f
C7746 VDD.n1496 VSS 0.00698f
C7747 VDD.n1497 VSS 0.00101f
C7748 VDD.n1498 VSS 0.00164f
C7749 VDD.n1499 VSS 0.00285f
C7750 VDD.n1500 VSS 0.00285f
C7751 VDD.n1501 VSS 0.00285f
C7752 VDD.n1502 VSS 0.0014f
C7753 VDD.n1503 VSS 0.00101f
C7754 VDD.n1504 VSS 0.00535f
C7755 VDD.t342 VSS 0.00535f
C7756 VDD.n1505 VSS 0.00791f
C7757 VDD.n1506 VSS 0.00489f
C7758 VDD.t324 VSS 0.00535f
C7759 VDD.n1507 VSS 0.00838f
C7760 VDD.n1508 VSS 0.00101f
C7761 VDD.n1509 VSS 0.0011f
C7762 VDD.n1510 VSS 0.00285f
C7763 VDD.t325 VSS 5.58e-19
C7764 VDD.t664 VSS 5.58e-19
C7765 VDD.n1511 VSS 0.00121f
C7766 VDD.n1512 VSS 0.0025f
C7767 VDD.n1513 VSS 0.00285f
C7768 VDD.n1514 VSS 0.00169f
C7769 VDD.n1515 VSS 0.0014f
C7770 VDD.n1516 VSS 0.00101f
C7771 VDD.n1517 VSS 0.00716f
C7772 VDD.t376 VSS 0.00535f
C7773 VDD.t619 VSS 0.00535f
C7774 VDD.n1518 VSS 0.00553f
C7775 VDD.n1519 VSS 0.00101f
C7776 VDD.n1520 VSS 9.18e-19
C7777 VDD.n1521 VSS 0.00285f
C7778 VDD.n1522 VSS 0.00285f
C7779 VDD.n1523 VSS 2.64e-19
C7780 VDD.t756 VSS 8.03e-19
C7781 VDD.n1524 VSS 0.0026f
C7782 VDD.t543 VSS 0.00148f
C7783 VDD.t618 VSS -4.69e-19
C7784 VDD.t545 VSS 8.48e-19
C7785 VDD.n1525 VSS 0.00333f
C7786 VDD.n1526 VSS 0.00189f
C7787 VDD.n1527 VSS 0.00329f
C7788 VDD.n1528 VSS 3.68e-19
C7789 VDD.n1529 VSS 7.03e-19
C7790 VDD.n1530 VSS 0.00143f
C7791 VDD.n1531 VSS 0.00261f
C7792 VDD.n1532 VSS 0.00285f
C7793 VDD.n1533 VSS 0.00165f
C7794 VDD.n1534 VSS 6.26e-19
C7795 VDD.n1535 VSS 0.00855f
C7796 VDD.t617 VSS 0.00884f
C7797 VDD.t544 VSS 0.0129f
C7798 VDD.n1536 VSS 0.011f
C7799 VDD.t675 VSS 0.00535f
C7800 VDD.n1537 VSS 0.00617f
C7801 VDD.t123 VSS 0.00535f
C7802 VDD.n1538 VSS 0.00419f
C7803 VDD.n1539 VSS 0.00101f
C7804 VDD.n1540 VSS 7.04e-19
C7805 VDD.n1541 VSS 0.00247f
C7806 VDD.n1542 VSS 0.00284f
C7807 VDD.n1543 VSS 0.00285f
C7808 VDD.n1544 VSS 0.00285f
C7809 VDD.n1545 VSS 0.00285f
C7810 VDD.n1546 VSS 0.00152f
C7811 VDD.n1547 VSS 0.00189f
C7812 VDD.n1548 VSS 0.00102f
C7813 VDD.n1549 VSS 0.00704f
C7814 VDD.t621 VSS 0.00535f
C7815 VDD.n1550 VSS 0.00558f
C7816 VDD.n1551 VSS 0.00489f
C7817 VDD.t140 VSS 0.00535f
C7818 VDD.n1552 VSS 0.00588f
C7819 VDD.n1553 VSS 0.00101f
C7820 VDD.n1554 VSS 0.00172f
C7821 VDD.n1555 VSS 0.00285f
C7822 VDD.n1556 VSS 0.00285f
C7823 VDD.n1557 VSS 0.00285f
C7824 VDD.n1558 VSS 0.00172f
C7825 VDD.n1559 VSS 0.00101f
C7826 VDD.n1560 VSS 0.00838f
C7827 VDD.t331 VSS 0.00535f
C7828 VDD.n1561 VSS 0.00762f
C7829 VDD.t214 VSS 0.005f
C7830 VDD.t673 VSS 0.00524f
C7831 VDD.n1562 VSS 0.0057f
C7832 VDD.n1563 VSS 0.00101f
C7833 VDD.n1564 VSS 9.47e-19
C7834 VDD.n1565 VSS 0.00285f
C7835 VDD.n1566 VSS 0.00285f
C7836 VDD.n1567 VSS 0.00285f
C7837 VDD.n1568 VSS 0.0011f
C7838 VDD.n1569 VSS 0.00101f
C7839 VDD.n1570 VSS 0.00617f
C7840 VDD.t88 VSS 0.00535f
C7841 VDD.n1571 VSS 0.00617f
C7842 VDD.t333 VSS 0.00535f
C7843 VDD.n1572 VSS 0.00489f
C7844 VDD.t97 VSS 0.00535f
C7845 VDD.n1573 VSS 0.00698f
C7846 VDD.n1574 VSS 0.00101f
C7847 VDD.n1575 VSS 0.00164f
C7848 VDD.n1576 VSS 0.00285f
C7849 VDD.n1577 VSS 0.00285f
C7850 VDD.n1578 VSS 0.00285f
C7851 VDD.n1579 VSS 0.0014f
C7852 VDD.n1580 VSS 0.00101f
C7853 VDD.n1581 VSS 0.00535f
C7854 VDD.t563 VSS 0.00535f
C7855 VDD.n1582 VSS 0.00791f
C7856 VDD.n1583 VSS 0.00489f
C7857 VDD.t142 VSS 0.00535f
C7858 VDD.n1584 VSS 0.00838f
C7859 VDD.n1585 VSS 0.00101f
C7860 VDD.n1586 VSS 0.0011f
C7861 VDD.n1587 VSS 0.00285f
C7862 VDD.t143 VSS 5.58e-19
C7863 VDD.t201 VSS 5.58e-19
C7864 VDD.n1588 VSS 0.00121f
C7865 VDD.n1589 VSS 0.0025f
C7866 VDD.n1590 VSS 0.00285f
C7867 VDD.n1591 VSS 0.00169f
C7868 VDD.n1592 VSS 0.0014f
C7869 VDD.n1593 VSS 0.00101f
C7870 VDD.n1594 VSS 0.00716f
C7871 VDD.t751 VSS 0.00535f
C7872 VDD.t640 VSS 0.00535f
C7873 VDD.n1595 VSS 0.00553f
C7874 VDD.n1596 VSS 0.00101f
C7875 VDD.n1597 VSS 9.18e-19
C7876 VDD.n1598 VSS 0.00285f
C7877 VDD.n1599 VSS 0.00285f
C7878 VDD.n1600 VSS 2.64e-19
C7879 VDD.t763 VSS 8.03e-19
C7880 VDD.n1601 VSS 0.0026f
C7881 VDD.t522 VSS 0.00148f
C7882 VDD.t639 VSS -4.69e-19
C7883 VDD.t524 VSS 8.48e-19
C7884 VDD.n1602 VSS 0.00333f
C7885 VDD.n1603 VSS 0.00189f
C7886 VDD.n1604 VSS 0.00328f
C7887 VDD.n1605 VSS 3.68e-19
C7888 VDD.n1606 VSS 7.03e-19
C7889 VDD.n1607 VSS 0.00143f
C7890 VDD.n1608 VSS 0.00261f
C7891 VDD.n1609 VSS 0.00285f
C7892 VDD.n1610 VSS 0.00165f
C7893 VDD.n1611 VSS 6.26e-19
C7894 VDD.n1612 VSS 0.00855f
C7895 VDD.t638 VSS 0.00884f
C7896 VDD.t523 VSS 0.0129f
C7897 VDD.n1613 VSS 0.011f
C7898 VDD.t719 VSS 0.00535f
C7899 VDD.n1614 VSS 0.00617f
C7900 VDD.t296 VSS 0.00535f
C7901 VDD.n1615 VSS 0.00419f
C7902 VDD.n1616 VSS 0.00101f
C7903 VDD.n1617 VSS 7.23e-19
C7904 VDD.n1618 VSS 0.00247f
C7905 VDD.n1619 VSS 0.00284f
C7906 VDD.n1620 VSS 0.00285f
C7907 VDD.n1621 VSS 0.00285f
C7908 VDD.n1622 VSS 0.00285f
C7909 VDD.n1623 VSS 0.00152f
C7910 VDD.n1624 VSS 0.00189f
C7911 VDD.n1625 VSS 0.00102f
C7912 VDD.n1626 VSS 0.00704f
C7913 VDD.t642 VSS 0.00535f
C7914 VDD.n1627 VSS 0.00558f
C7915 VDD.n1628 VSS 0.00489f
C7916 VDD.t115 VSS 0.00535f
C7917 VDD.n1629 VSS 0.00588f
C7918 VDD.n1630 VSS 0.00101f
C7919 VDD.n1631 VSS 0.00172f
C7920 VDD.n1632 VSS 0.00285f
C7921 VDD.n1633 VSS 0.00285f
C7922 VDD.n1634 VSS 0.00285f
C7923 VDD.n1635 VSS 0.00172f
C7924 VDD.n1636 VSS 0.00101f
C7925 VDD.n1637 VSS 0.00838f
C7926 VDD.t458 VSS 0.00535f
C7927 VDD.n1638 VSS 0.00762f
C7928 VDD.t742 VSS 0.005f
C7929 VDD.t721 VSS 0.00524f
C7930 VDD.n1639 VSS 0.0057f
C7931 VDD.n1640 VSS 0.00101f
C7932 VDD.n1641 VSS 9.47e-19
C7933 VDD.n1642 VSS 0.00285f
C7934 VDD.n1643 VSS 0.00285f
C7935 VDD.n1644 VSS 0.00285f
C7936 VDD.n1645 VSS 0.0011f
C7937 VDD.n1646 VSS 0.00101f
C7938 VDD.n1647 VSS 0.00617f
C7939 VDD.t31 VSS 0.00535f
C7940 VDD.n1648 VSS 0.00617f
C7941 VDD.t456 VSS 0.00535f
C7942 VDD.n1649 VSS 0.00489f
C7943 VDD.t703 VSS 0.00535f
C7944 VDD.n1650 VSS 0.00698f
C7945 VDD.n1651 VSS 0.00101f
C7946 VDD.n1652 VSS 0.00164f
C7947 VDD.n1653 VSS 0.00285f
C7948 VDD.n1654 VSS 0.00285f
C7949 VDD.n1655 VSS 0.00285f
C7950 VDD.n1656 VSS 0.0014f
C7951 VDD.n1657 VSS 0.00101f
C7952 VDD.n1658 VSS 0.00535f
C7953 VDD.t263 VSS 0.00535f
C7954 VDD.n1659 VSS 0.00791f
C7955 VDD.n1660 VSS 0.00489f
C7956 VDD.t113 VSS 0.00535f
C7957 VDD.n1661 VSS 0.00838f
C7958 VDD.n1662 VSS 0.00101f
C7959 VDD.n1663 VSS 0.0011f
C7960 VDD.n1664 VSS 0.00285f
C7961 VDD.t114 VSS 5.58e-19
C7962 VDD.t275 VSS 5.58e-19
C7963 VDD.n1665 VSS 0.00121f
C7964 VDD.n1666 VSS 0.0025f
C7965 VDD.n1667 VSS 0.00285f
C7966 VDD.n1668 VSS 0.00169f
C7967 VDD.n1669 VSS 0.0014f
C7968 VDD.n1670 VSS 0.00101f
C7969 VDD.n1671 VSS 0.00716f
C7970 VDD.t655 VSS 0.00535f
C7971 VDD.t567 VSS 0.00535f
C7972 VDD.n1672 VSS 0.00553f
C7973 VDD.n1673 VSS 0.00101f
C7974 VDD.n1674 VSS 9.18e-19
C7975 VDD.n1675 VSS 0.00285f
C7976 VDD.n1676 VSS 0.00285f
C7977 VDD.n1677 VSS 2.64e-19
C7978 VDD.t765 VSS 8.03e-19
C7979 VDD.n1678 VSS 0.0026f
C7980 VDD.t516 VSS 0.00148f
C7981 VDD.t572 VSS -4.69e-19
C7982 VDD.t518 VSS 8.48e-19
C7983 VDD.n1679 VSS 0.00333f
C7984 VDD.n1680 VSS 0.00189f
C7985 VDD.n1681 VSS 0.00328f
C7986 VDD.n1682 VSS 3.68e-19
C7987 VDD.n1683 VSS 7.03e-19
C7988 VDD.n1684 VSS 0.00143f
C7989 VDD.n1685 VSS 0.00261f
C7990 VDD.n1686 VSS 0.00285f
C7991 VDD.n1687 VSS 0.00165f
C7992 VDD.n1688 VSS 6.26e-19
C7993 VDD.n1689 VSS 0.00855f
C7994 VDD.t571 VSS 0.00884f
C7995 VDD.t517 VSS 0.0129f
C7996 VDD.n1690 VSS 0.011f
C7997 VDD.t329 VSS 0.00535f
C7998 VDD.n1691 VSS 0.00617f
C7999 VDD.t704 VSS 0.00535f
C8000 VDD.n1692 VSS 0.00419f
C8001 VDD.n1693 VSS 0.00101f
C8002 VDD.n1694 VSS 6.94e-19
C8003 VDD.n1695 VSS 0.00247f
C8004 VDD.n1696 VSS 0.00284f
C8005 VDD.n1697 VSS 0.00285f
C8006 VDD.n1698 VSS 0.00285f
C8007 VDD.n1699 VSS 0.00285f
C8008 VDD.n1700 VSS 0.00152f
C8009 VDD.n1701 VSS 0.00189f
C8010 VDD.n1702 VSS 0.00102f
C8011 VDD.n1703 VSS 0.00704f
C8012 VDD.t569 VSS 0.00535f
C8013 VDD.n1704 VSS 0.00558f
C8014 VDD.n1705 VSS 0.00489f
C8015 VDD.t158 VSS 0.00535f
C8016 VDD.n1706 VSS 0.00588f
C8017 VDD.n1707 VSS 0.00101f
C8018 VDD.n1708 VSS 0.00172f
C8019 VDD.n1709 VSS 0.00285f
C8020 VDD.n1710 VSS 0.00285f
C8021 VDD.n1711 VSS 0.00285f
C8022 VDD.n1712 VSS 0.00172f
C8023 VDD.n1713 VSS 0.00101f
C8024 VDD.n1714 VSS 0.00838f
C8025 VDD.t194 VSS 0.00535f
C8026 VDD.n1715 VSS 0.00762f
C8027 VDD.t654 VSS 0.005f
C8028 VDD.t327 VSS 0.00524f
C8029 VDD.n1716 VSS 0.0057f
C8030 VDD.n1717 VSS 0.00101f
C8031 VDD.n1718 VSS 9.47e-19
C8032 VDD.n1719 VSS 0.00285f
C8033 VDD.n1720 VSS 0.00285f
C8034 VDD.n1721 VSS 0.00285f
C8035 VDD.n1722 VSS 0.0011f
C8036 VDD.n1723 VSS 0.00101f
C8037 VDD.n1724 VSS 0.00617f
C8038 VDD.t202 VSS 0.00535f
C8039 VDD.n1725 VSS 0.00617f
C8040 VDD.t192 VSS 0.00535f
C8041 VDD.n1726 VSS 0.00535f
C8042 VDD.t155 VSS 0.00535f
C8043 VDD.n1727 VSS 0.00489f
C8044 VDD.t422 VSS 0.00535f
C8045 VDD.n1728 VSS 0.00698f
C8046 VDD.n1729 VSS 0.00101f
C8047 VDD.n1730 VSS 0.00164f
C8048 VDD.n1731 VSS 0.00285f
C8049 VDD.n1732 VSS 0.00285f
C8050 VDD.n1733 VSS 0.00285f
C8051 VDD.n1734 VSS 0.00285f
C8052 VDD.n1735 VSS 0.0014f
C8053 VDD.n1736 VSS 0.00188f
C8054 VDD.n1737 VSS 0.00102f
C8055 VDD.n1738 VSS 0.00791f
C8056 VDD.n1739 VSS 0.00838f
C8057 VDD.t156 VSS 0.00535f
C8058 VDD.t577 VSS 0.00535f
C8059 VDD.n1740 VSS 0.00489f
C8060 VDD.n1741 VSS 0.00102f
C8061 VDD.n1742 VSS 0.00187f
C8062 VDD.n1743 VSS 0.0025f
C8063 VDD.n1744 VSS 0.00285f
C8064 VDD.n1745 VSS 0.00169f
C8065 VDD.n1746 VSS 0.00214f
C8066 VDD.n1747 VSS 0.00167f
C8067 VDD.n1748 VSS 0.00101f
C8068 VDD.n1749 VSS 0.00716f
C8069 VDD.t2 VSS 0.00535f
C8070 VDD.n1750 VSS 0.00553f
C8071 VDD.t648 VSS 0.00535f
C8072 VDD.n1751 VSS 0.00774f
C8073 VDD.t646 VSS 0.00884f
C8074 VDD.n1752 VSS 0.00855f
C8075 VDD.n1753 VSS 6.26e-19
C8076 VDD.n1754 VSS 0.00101f
C8077 VDD.n1755 VSS 0.00172f
C8078 VDD.n1756 VSS 0.00285f
C8079 VDD.n1757 VSS 0.00285f
C8080 VDD.n1758 VSS 0.00261f
C8081 VDD.n1759 VSS 0.00173f
C8082 VDD.t647 VSS -4.69e-19
C8083 VDD.t548 VSS 8.48e-19
C8084 VDD.n1760 VSS 0.00333f
C8085 VDD.n1761 VSS 0.00189f
C8086 VDD.n1762 VSS 0.00329f
C8087 VDD.n1763 VSS 7.03e-19
C8088 VDD.n1764 VSS 3.68e-19
C8089 VDD.n1765 VSS 2.64e-19
C8090 VDD.n1766 VSS 0.00143f
C8091 VDD.n1767 VSS 0.00285f
C8092 VDD.n1768 VSS 0.00284f
C8093 VDD.n1769 VSS 0.00247f
C8094 VDD.n1770 VSS 8.78e-19
C8095 VDD.n1771 VSS 0.011f
C8096 VDD.t665 VSS 0.00535f
C8097 VDD.n1772 VSS 0.00419f
C8098 VDD.t16 VSS 0.00535f
C8099 VDD.t644 VSS 0.00535f
C8100 VDD.n1773 VSS 0.00704f
C8101 VDD.t380 VSS 0.00535f
C8102 VDD.n1774 VSS 0.00617f
C8103 VDD.n1775 VSS 0.00101f
C8104 VDD.n1776 VSS 0.00152f
C8105 VDD.n1777 VSS 0.00189f
C8106 VDD.n1778 VSS 0.00234f
C8107 VDD.n1779 VSS 0.00285f
C8108 VDD.n1780 VSS 0.00285f
C8109 VDD.n1781 VSS 0.00285f
C8110 VDD.n1782 VSS 0.00285f
C8111 VDD.n1783 VSS 0.00172f
C8112 VDD.n1784 VSS 0.00101f
C8113 VDD.n1785 VSS 0.00588f
C8114 VDD.t112 VSS 0.00535f
C8115 VDD.n1786 VSS 0.00489f
C8116 VDD.t428 VSS 0.00535f
C8117 VDD.t52 VSS 0.00535f
C8118 VDD.n1787 VSS 0.00838f
C8119 VDD.n1788 VSS 0.00101f
C8120 VDD.n1789 VSS 0.00172f
C8121 VDD.n1790 VSS 0.00102f
C8122 VDD.n1791 VSS 0.00285f
C8123 VDD.n1792 VSS 0.00285f
C8124 VDD.n1793 VSS 9.47e-19
C8125 VDD.n1794 VSS 0.00101f
C8126 VDD.n1795 VSS 0.0057f
C8127 VDD.t667 VSS 0.00524f
C8128 VDD.t73 VSS 0.005f
C8129 VDD.n1796 VSS 0.00547f
C8130 VDD.n1797 VSS 0.00617f
C8131 VDD.t477 VSS 0.00535f
C8132 VDD.n1798 VSS 0.00617f
C8133 VDD.n1799 VSS 0.00101f
C8134 VDD.n1800 VSS 0.0011f
C8135 VDD.n1801 VSS 0.00285f
C8136 VDD.t478 VSS 5.29e-19
C8137 VDD.t51 VSS 5.02e-19
C8138 VDD.n1802 VSS 0.0011f
C8139 VDD.n1803 VSS 0.00257f
C8140 VDD.n1804 VSS 0.00285f
C8141 VDD.n1805 VSS 0.00285f
C8142 VDD.n1806 VSS 0.00164f
C8143 VDD.n1807 VSS 0.00101f
C8144 VDD.n1808 VSS 0.00698f
C8145 VDD.t427 VSS 0.00535f
C8146 VDD.n1809 VSS 0.00489f
C8147 VDD.t109 VSS 0.00535f
C8148 VDD.t284 VSS 0.00535f
C8149 VDD.n1810 VSS 0.00535f
C8150 VDD.n1811 VSS 0.00101f
C8151 VDD.n1812 VSS 0.0014f
C8152 VDD.n1813 VSS 0.00285f
C8153 VDD.t285 VSS 0.00131f
C8154 VDD.n1814 VSS 0.00289f
C8155 VDD.n1815 VSS 0.00285f
C8156 VDD.n1816 VSS 0.00285f
C8157 VDD.n1817 VSS 0.0011f
C8158 VDD.n1818 VSS 0.00101f
C8159 VDD.n1819 VSS 0.00838f
C8160 VDD.t110 VSS 0.00535f
C8161 VDD.n1820 VSS 0.00489f
C8162 VDD.t210 VSS 0.00535f
C8163 VDD.n1821 VSS 9.81e-19
C8164 VDD.n1822 VSS 0.0014f
C8165 VDD.n1823 VSS 0.00169f
C8166 VDD.n1824 VSS 0.00285f
C8167 VDD.t485 VSS 7.16e-19
C8168 VDD.t44 VSS 2.33e-19
C8169 VDD.n1825 VSS 0.00366f
C8170 VDD.n1826 VSS 0.00285f
C8171 VDD.n1827 VSS 0.00101f
C8172 VDD.t467 VSS 0.00541f
C8173 VDD.n1828 VSS 0.00101f
C8174 VDD.n1829 VSS 0.00172f
C8175 VDD.n1830 VSS 8.81e-19
C8176 VDD.n1831 VSS 0.00285f
C8177 VDD.n1832 VSS 0.00172f
C8178 VDD.n1833 VSS 0.00101f
C8179 VDD.t482 VSS 0.00541f
C8180 VDD.n1834 VSS 0.00101f
C8181 VDD.t483 VSS 3.94e-19
C8182 VDD.t178 VSS 5.02e-19
C8183 VDD.n1835 VSS 0.00103f
C8184 VDD.n1836 VSS 0.0024f
C8185 VDD.n1837 VSS 0.0115f
C8186 VDD.n1838 VSS 0.00146f
C8187 VDD.n1839 VSS 0.00101f
C8188 VDD.n1840 VSS 0.0108f
C8189 VDD.n1841 VSS 0.00101f
C8190 VDD.n1842 VSS 0.00146f
C8191 VDD.n1843 VSS 0.00101f
C8192 VDD.n1844 VSS 0.0108f
C8193 VDD.n1845 VSS 0.00101f
C8194 VDD.n1846 VSS 8.62e-19
C8195 VDD.n1847 VSS 0.00285f
C8196 VDD.t432 VSS 5.02e-19
C8197 VDD.t75 VSS 3.94e-19
C8198 VDD.n1848 VSS 0.00103f
C8199 VDD.n1849 VSS 0.00204f
C8200 VDD.n1850 VSS 0.00101f
C8201 VDD.n1851 VSS 0.00101f
C8202 VDD.n1852 VSS 0.00953f
C8203 VDD.n1853 VSS 0.00101f
C8204 VDD.n1854 VSS 8.62e-19
C8205 VDD.n1855 VSS 7.87e-19
C8206 VDD.n1856 VSS 8.62e-19
C8207 VDD.n1857 VSS 0.00285f
C8208 VDD.n1858 VSS 8.62e-19
C8209 VDD.n1859 VSS 0.00101f
C8210 VDD.t429 VSS 0.00541f
C8211 VDD.n1860 VSS 0.00101f
C8212 VDD.n1861 VSS 8.62e-19
C8213 VDD.t170 VSS 7.16e-19
C8214 VDD.t430 VSS 2.33e-19
C8215 VDD.n1862 VSS 0.00366f
C8216 VDD.n1863 VSS 8.62e-19
C8217 VDD.n1864 VSS 0.00285f
C8218 VDD.t687 VSS 7.16e-19
C8219 VDD.t300 VSS 2.33e-19
C8220 VDD.n1865 VSS 0.00366f
C8221 VDD.n1866 VSS 0.00285f
C8222 VDD.n1867 VSS 0.00112f
C8223 VDD.n1868 VSS 0.00145f
C8224 VDD.n1869 VSS 0.00101f
C8225 VDD.t464 VSS 0.00541f
C8226 VDD.n1870 VSS 0.00101f
C8227 VDD.n1871 VSS 0.00172f
C8228 VDD.n1872 VSS 8.81e-19
C8229 VDD.n1873 VSS 0.00285f
C8230 VDD.n1874 VSS 0.00172f
C8231 VDD.n1875 VSS 0.00101f
C8232 VDD.t356 VSS 0.00541f
C8233 VDD.n1876 VSS 0.00101f
C8234 VDD.t357 VSS 3.94e-19
C8235 VDD.t160 VSS 5.02e-19
C8236 VDD.n1877 VSS 0.00103f
C8237 VDD.n1878 VSS 0.0024f
C8238 VDD.n1879 VSS 0.0115f
C8239 VDD.n1880 VSS 0.00146f
C8240 VDD.n1881 VSS 0.00101f
C8241 VDD.n1882 VSS 0.0108f
C8242 VDD.n1883 VSS 0.00101f
C8243 VDD.n1884 VSS 0.00146f
C8244 VDD.n1885 VSS 9.9e-19
C8245 VDD.n1886 VSS 0.0108f
C8246 VDD.n1887 VSS 9.92e-19
C8247 VDD.n1888 VSS 8.62e-19
C8248 VDD.n1889 VSS 0.00285f
C8249 VDD.t672 VSS 5.02e-19
C8250 VDD.t172 VSS 3.94e-19
C8251 VDD.n1890 VSS 0.00103f
C8252 VDD.n1891 VSS 0.00204f
C8253 VDD.n1892 VSS 0.00101f
C8254 VDD.n1893 VSS 0.00101f
C8255 VDD.n1894 VSS 0.00953f
C8256 VDD.n1895 VSS 0.00101f
C8257 VDD.n1896 VSS 8.62e-19
C8258 VDD.n1897 VSS 7.87e-19
C8259 VDD.n1898 VSS 8.62e-19
C8260 VDD.n1899 VSS 0.00285f
C8261 VDD.n1900 VSS 8.62e-19
C8262 VDD.n1901 VSS 0.00101f
C8263 VDD.t100 VSS 0.00541f
C8264 VDD.n1902 VSS 0.00101f
C8265 VDD.n1903 VSS 8.62e-19
C8266 VDD.t487 VSS 7.16e-19
C8267 VDD.t101 VSS 2.33e-19
C8268 VDD.n1904 VSS 0.00366f
C8269 VDD.n1905 VSS 8.62e-19
C8270 VDD.n1906 VSS 0.00285f
C8271 VDD.t353 VSS 7.16e-19
C8272 VDD.t447 VSS 2.33e-19
C8273 VDD.n1907 VSS 0.00366f
C8274 VDD.n1908 VSS 0.00285f
C8275 VDD.n1909 VSS 0.00112f
C8276 VDD.n1910 VSS 0.00145f
C8277 VDD.n1911 VSS 0.00101f
C8278 VDD.n1912 VSS 0.00101f
C8279 VDD.t465 VSS 0.00541f
C8280 VDD.n1913 VSS 0.00101f
C8281 VDD.n1914 VSS 0.00172f
C8282 VDD.n1915 VSS 8.81e-19
C8283 VDD.n1916 VSS 0.00285f
C8284 VDD.n1917 VSS 0.00172f
C8285 VDD.n1918 VSS 0.00101f
C8286 VDD.t679 VSS 0.00541f
C8287 VDD.n1919 VSS 0.00101f
C8288 VDD.t680 VSS 3.94e-19
C8289 VDD.t591 VSS 5.02e-19
C8290 VDD.n1920 VSS 0.00103f
C8291 VDD.n1921 VSS 0.0024f
C8292 VDD.n1922 VSS 0.0115f
C8293 VDD.n1923 VSS 0.00546f
C8294 VDD.n1924 VSS 0.00349f
C8295 VDD.n1925 VSS 0.00553f
C8296 VDD.n1926 VSS 0.00101f
C8297 VDD.n1927 VSS 0.00129f
C8298 VDD.n1928 VSS 0.00285f
C8299 VDD.n1929 VSS 0.00172f
C8300 VDD.t556 VSS 5.02e-19
C8301 VDD.t426 VSS 3.94e-19
C8302 VDD.n1930 VSS 0.00103f
C8303 VDD.n1931 VSS 0.0024f
C8304 VDD.n1932 VSS 0.00101f
C8305 VDD.n1933 VSS 0.00635f
C8306 VDD.n1934 VSS 0.00101f
C8307 VDD.n1935 VSS 0.00172f
C8308 VDD.n1936 VSS 0.00258f
C8309 VDD.n1937 VSS 8.81e-19
C8310 VDD.n1938 VSS 0.00101f
C8311 VDD.n1939 VSS 0.0108f
C8312 VDD.n1940 VSS 0.00101f
C8313 VDD.n1941 VSS 0.00145f
C8314 VDD.t678 VSS 7.16e-19
C8315 VDD.t658 VSS 2.33e-19
C8316 VDD.n1942 VSS 0.00366f
C8317 VDD.n1943 VSS 0.00285f
C8318 VDD.n1944 VSS 0.00285f
C8319 VDD.n1945 VSS 8.44e-19
C8320 VDD.n1946 VSS 0.00101f
C8321 VDD.t632 VSS 0.00541f
C8322 VDD.n1947 VSS 0.00101f
C8323 VDD.n1948 VSS 8.62e-19
C8324 VDD.n1949 VSS 0.00285f
C8325 VDD.n1950 VSS 8.62e-19
C8326 VDD.n1951 VSS 0.00101f
C8327 VDD.t86 VSS 0.00541f
C8328 VDD.n1952 VSS 0.00101f
C8329 VDD.n1953 VSS 8.06e-19
C8330 VDD.n1954 VSS 8.62e-19
C8331 VDD.n1955 VSS 0.0115f
C8332 VDD.n1956 VSS 8.7e-19
C8333 VDD.n1957 VSS 0.00101f
C8334 VDD.n1958 VSS 0.0108f
C8335 VDD.n1959 VSS 0.00101f
C8336 VDD.n1960 VSS 0.00146f
C8337 VDD.n1961 VSS 0.00101f
C8338 VDD.n1962 VSS 0.00988f
C8339 VDD.n1963 VSS 9.23e-19
C8340 VDD.n1964 VSS 1.59e-19
C8341 VDD.n1965 VSS 9.34e-20
C8342 VDD.n1966 VSS 0.00535f
C8343 VDD.n1967 VSS 5e-19
C8344 VDD.n1968 VSS 1.59e-19
C8345 VDD.n1969 VSS 0.00118f
C8346 VDD.n1970 VSS 1.87e-20
C8347 VDD.n1971 VSS 4.18e-19
C8348 VDD.n1972 VSS 1e-18
C8349 VDD.n1973 VSS 9.34e-20
C8350 VDD.n1974 VSS 1.59e-19
C8351 VDD.t322 VSS 5.02e-19
C8352 VDD.t385 VSS 3.94e-19
C8353 VDD.n1975 VSS 0.00103f
C8354 VDD.n1976 VSS 1.59e-19
C8355 VDD.n1977 VSS 2.64e-19
C8356 VDD.n1978 VSS 1.59e-19
C8357 VDD.n1979 VSS 5e-19
C8358 VDD.n1980 VSS 0.00447f
C8359 VDD.n1981 VSS 4.18e-19
C8360 VDD.n1982 VSS 1.87e-20
C8361 VDD.n1983 VSS 0.00141f
C8362 VDD.n1984 VSS 1.59e-19
C8363 VDD.n1985 VSS 9.34e-20
C8364 VDD.n1986 VSS 0.00535f
C8365 VDD.n1987 VSS 5e-19
C8366 VDD.n1988 VSS 1.59e-19
C8367 VDD.n1989 VSS 0.00118f
C8368 VDD.n1990 VSS 1.87e-20
C8369 VDD.n1991 VSS 4.18e-19
C8370 VDD.n1992 VSS 1e-18
C8371 VDD.n1993 VSS 9.34e-20
C8372 VDD.n1994 VSS 1.59e-19
C8373 VDD.n1995 VSS 1.59e-19
C8374 VDD.n1996 VSS 2.64e-19
C8375 VDD.n1997 VSS 1.59e-19
C8376 VDD.n1998 VSS 5e-19
C8377 VDD.n1999 VSS 0.00188f
C8378 VDD.n2000 VSS 4.18e-19
C8379 VDD.n2001 VSS 1.87e-20
C8380 VDD.n2002 VSS 0.00115f
C8381 VDD.t133 VSS 7.16e-19
C8382 VDD.t24 VSS 2.33e-19
C8383 VDD.n2003 VSS 0.00366f
C8384 VDD.n2004 VSS 1.59e-19
C8385 VDD.n2005 VSS 9.34e-20
C8386 VDD.n2006 VSS 0.0108f
C8387 VDD.n2007 VSS 0.00101f
C8388 VDD.n2008 VSS 1.59e-19
C8389 VDD.n2009 VSS 8.62e-19
C8390 VDD.n2010 VSS 0.00101f
C8391 VDD.t382 VSS 0.00541f
C8392 VDD.n2011 VSS 0.00101f
C8393 VDD.n2012 VSS 8.62e-19
C8394 VDD.t383 VSS 7.16e-19
C8395 VDD.t287 VSS 2.33e-19
C8396 VDD.n2013 VSS 0.00366f
C8397 VDD.n2014 VSS 8.44e-19
C8398 VDD.n2015 VSS 0.00237f
C8399 VDD.n2016 VSS 0.00285f
C8400 VDD.n2017 VSS 8.62e-19
C8401 VDD.n2018 VSS 0.00101f
C8402 VDD.t439 VSS 0.00541f
C8403 VDD.n2019 VSS 0.00101f
C8404 VDD.n2020 VSS 8.06e-19
C8405 VDD.n2021 VSS 8.62e-19
C8406 VDD.n2022 VSS 0.0115f
C8407 VDD.n2023 VSS 8.7e-19
C8408 VDD.n2024 VSS 0.00101f
C8409 VDD.n2025 VSS 0.0108f
C8410 VDD.n2026 VSS 0.00101f
C8411 VDD.n2027 VSS 0.00146f
C8412 VDD.n2028 VSS 0.00101f
C8413 VDD.n2029 VSS 0.00988f
C8414 VDD.n2030 VSS 9.23e-19
C8415 VDD.n2031 VSS 1.59e-19
C8416 VDD.n2032 VSS 9.34e-20
C8417 VDD.n2033 VSS 0.00535f
C8418 VDD.n2034 VSS 5e-19
C8419 VDD.n2035 VSS 1.59e-19
C8420 VDD.n2036 VSS 0.00118f
C8421 VDD.n2037 VSS 1.87e-20
C8422 VDD.n2038 VSS 4.18e-19
C8423 VDD.n2039 VSS 1e-18
C8424 VDD.n2040 VSS 9.34e-20
C8425 VDD.n2041 VSS 1.59e-19
C8426 VDD.t302 VSS 5.02e-19
C8427 VDD.t162 VSS 3.94e-19
C8428 VDD.n2042 VSS 0.00103f
C8429 VDD.n2043 VSS 1.59e-19
C8430 VDD.n2044 VSS 2.64e-19
C8431 VDD.n2045 VSS 1.59e-19
C8432 VDD.n2046 VSS 5e-19
C8433 VDD.n2047 VSS 0.00447f
C8434 VDD.n2048 VSS 4.18e-19
C8435 VDD.n2049 VSS 1.87e-20
C8436 VDD.n2050 VSS 0.00141f
C8437 VDD.n2051 VSS 1.59e-19
C8438 VDD.n2052 VSS 9.34e-20
C8439 VDD.n2053 VSS 0.00535f
C8440 VDD.n2054 VSS 5e-19
C8441 VDD.n2055 VSS 1.59e-19
C8442 VDD.n2056 VSS 0.00118f
C8443 VDD.n2057 VSS 1.87e-20
C8444 VDD.n2058 VSS 4.18e-19
C8445 VDD.n2059 VSS 1e-18
C8446 VDD.n2060 VSS 9.34e-20
C8447 VDD.n2061 VSS 1.59e-19
C8448 VDD.n2062 VSS 1.59e-19
C8449 VDD.n2063 VSS 2.64e-19
C8450 VDD.n2064 VSS 1.59e-19
C8451 VDD.n2065 VSS 5e-19
C8452 VDD.n2066 VSS 0.00188f
C8453 VDD.n2067 VSS 4.18e-19
C8454 VDD.n2068 VSS 1.87e-20
C8455 VDD.n2069 VSS 0.00115f
C8456 VDD.t489 VSS 7.16e-19
C8457 VDD.t277 VSS 2.33e-19
C8458 VDD.n2070 VSS 0.00366f
C8459 VDD.n2071 VSS 1.59e-19
C8460 VDD.n2072 VSS 9.34e-20
C8461 VDD.n2073 VSS 0.0138f
C8462 VDD.n2074 VSS 0.00125f
C8463 VDD.n2075 VSS 1.59e-19
C8464 VDD.n2076 VSS 1.59e-19
C8465 VDD.n2077 VSS 0.00126f
C8466 VDD.n2078 VSS 1.59e-19
C8467 VDD.n2079 VSS 9.34e-20
C8468 VDD.t340 VSS 0.00441f
C8469 VDD.n2080 VSS 4.72e-19
C8470 VDD.t125 VSS 7.16e-19
C8471 VDD.t341 VSS 2.33e-19
C8472 VDD.n2081 VSS 0.00366f
C8473 VDD.n2082 VSS 2.06e-19
C8474 VDD.n2083 VSS 2.64e-19
C8475 VDD.n2084 VSS 1.59e-19
C8476 VDD.n2085 VSS 1.59e-19
C8477 VDD.n2086 VSS 4.72e-19
C8478 VDD.n2087 VSS 9.34e-20
C8479 VDD.n2088 VSS 0.00318f
C8480 VDD.n2089 VSS 4.45e-19
C8481 VDD.n2090 VSS 6e-19
C8482 VDD.n2091 VSS 2.64e-19
C8483 VDD.n2092 VSS 1.59e-19
C8484 VDD.n2093 VSS 0.00133f
C8485 VDD.n2094 VSS 9.34e-20
C8486 VDD.n2095 VSS 0.00506f
C8487 VDD.n2096 VSS 4.72e-19
C8488 VDD.n2097 VSS 1.59e-19
C8489 VDD.n2098 VSS 0.00126f
C8490 VDD.n2099 VSS 6e-19
C8491 VDD.n2100 VSS 4.45e-19
C8492 VDD.t598 VSS 6.47e-19
C8493 VDD.n2101 VSS 9.34e-20
C8494 VDD.n2102 VSS 1.59e-19
C8495 VDD.n2103 VSS 6e-19
C8496 VDD.n2104 VSS 1.59e-19
C8497 VDD.n2105 VSS 2.64e-19
C8498 VDD.n2106 VSS 1.59e-19
C8499 VDD.n2107 VSS 4.72e-19
C8500 VDD.n2108 VSS 0.004f
C8501 VDD.n2109 VSS 4.45e-19
C8502 VDD.n2110 VSS 2.25e-19
C8503 VDD.n2111 VSS 2.64e-19
C8504 VDD.n2112 VSS 1.59e-19
C8505 VDD.n2113 VSS 0.00133f
C8506 VDD.n2114 VSS 9.34e-20
C8507 VDD.n2115 VSS 0.00506f
C8508 VDD.n2116 VSS 4.72e-19
C8509 VDD.n2117 VSS 1.59e-19
C8510 VDD.n2118 VSS 8.03e-19
C8511 VDD.n2119 VSS 5.05e-19
C8512 VDD.n2120 VSS 0.0108f
C8513 VDD.n2121 VSS 0.00101f
C8514 VDD.n2122 VSS 0.00146f
C8515 VDD.n2123 VSS 0.00101f
C8516 VDD.n2124 VSS 0.0107f
C8517 VDD.n2125 VSS 1e-18
C8518 VDD.n2126 VSS 1.59e-19
C8519 VDD.n2127 VSS 9.34e-20
C8520 VDD.n2128 VSS 0.00453f
C8521 VDD.n2129 VSS 4.23e-19
C8522 VDD.n2130 VSS 1.59e-19
C8523 VDD.n2131 VSS 0.0014f
C8524 VDD.n2132 VSS 2.81e-19
C8525 VDD.n2133 VSS 4.94e-19
C8526 VDD.n2134 VSS 1e-18
C8527 VDD.n2135 VSS 9.34e-20
C8528 VDD.n2136 VSS 1.59e-19
C8529 VDD.t103 VSS 5.02e-19
C8530 VDD.t660 VSS 3.94e-19
C8531 VDD.n2137 VSS 0.00103f
C8532 VDD.n2138 VSS 1.59e-19
C8533 VDD.n2139 VSS 2.64e-19
C8534 VDD.n2140 VSS 1.59e-19
C8535 VDD.n2141 VSS 4.23e-19
C8536 VDD.n2142 VSS 9.41e-19
C8537 VDD.n2143 VSS 4.94e-19
C8538 VDD.n2144 VSS 2.81e-19
C8539 VDD.n2145 VSS 0.00119f
C8540 VDD.n2146 VSS 1.59e-19
C8541 VDD.n2147 VSS 9.34e-20
C8542 VDD.n2148 VSS 0.00453f
C8543 VDD.n2149 VSS 4.23e-19
C8544 VDD.n2150 VSS 1.59e-19
C8545 VDD.n2151 VSS 0.0014f
C8546 VDD.n2152 VSS 2.81e-19
C8547 VDD.n2153 VSS 4.94e-19
C8548 VDD.n2154 VSS 1e-18
C8549 VDD.n2155 VSS 9.34e-20
C8550 VDD.n2156 VSS 1.59e-19
C8551 VDD.n2157 VSS 1.59e-19
C8552 VDD.n2158 VSS 2.64e-19
C8553 VDD.n2159 VSS 1.59e-19
C8554 VDD.n2160 VSS 4.23e-19
C8555 VDD.n2161 VSS 0.00353f
C8556 VDD.n2162 VSS 4.94e-19
C8557 VDD.n2163 VSS 2.81e-19
C8558 VDD.n2164 VSS 0.00115f
C8559 VDD.t379 VSS 7.16e-19
C8560 VDD.t188 VSS 2.33e-19
C8561 VDD.n2165 VSS 0.00366f
C8562 VDD.n2166 VSS 1.59e-19
C8563 VDD.n2167 VSS 9.34e-20
C8564 VDD.n2168 VSS 0.00994f
C8565 VDD.n2169 VSS 9.29e-19
C8566 VDD.n2170 VSS 1.59e-19
C8567 VDD.n2171 VSS 6.66e-19
C8568 VDD.n2172 VSS 5.05e-19
C8569 VDD.n2173 VSS 4.45e-19
C8570 VDD.n2174 VSS 6e-19
C8571 VDD.n2175 VSS 1.59e-19
C8572 VDD.n2176 VSS 2.64e-19
C8573 VDD.t347 VSS 7.16e-19
C8574 VDD.t624 VSS 2.33e-19
C8575 VDD.n2177 VSS 0.00366f
C8576 VDD.n2178 VSS 1.59e-19
C8577 VDD.n2179 VSS 0.00133f
C8578 VDD.n2180 VSS 9.34e-20
C8579 VDD.t346 VSS 0.00441f
C8580 VDD.n2181 VSS 4.72e-19
C8581 VDD.n2182 VSS 1.59e-19
C8582 VDD.n2183 VSS 0.00126f
C8583 VDD.n2184 VSS 6e-19
C8584 VDD.n2185 VSS 4.45e-19
C8585 VDD.n2186 VSS 1e-18
C8586 VDD.n2187 VSS 9.34e-20
C8587 VDD.n2188 VSS 1.59e-19
C8588 VDD.n2189 VSS 6e-19
C8589 VDD.n2190 VSS 1.59e-19
C8590 VDD.n2191 VSS 2.64e-19
C8591 VDD.n2192 VSS 1.59e-19
C8592 VDD.n2193 VSS 4.72e-19
C8593 VDD.n2194 VSS 0.00476f
C8594 VDD.n2195 VSS 4.45e-19
C8595 VDD.n2196 VSS 6e-19
C8596 VDD.n2197 VSS 2.64e-19
C8597 VDD.n2198 VSS 1.59e-19
C8598 VDD.n2199 VSS 0.00133f
C8599 VDD.n2200 VSS 9.34e-20
C8600 VDD.t354 VSS 0.00441f
C8601 VDD.n2201 VSS 4.72e-19
C8602 VDD.n2202 VSS 1.59e-19
C8603 VDD.n2203 VSS 0.00126f
C8604 VDD.n2204 VSS 2.25e-19
C8605 VDD.n2205 VSS 4.45e-19
C8606 VDD.n2206 VSS 1e-18
C8607 VDD.n2207 VSS 9.34e-20
C8608 VDD.n2208 VSS 1.59e-19
C8609 VDD.t15 VSS 3.94e-19
C8610 VDD.t355 VSS 5.02e-19
C8611 VDD.n2209 VSS 0.00103f
C8612 VDD.n2210 VSS 0.00208f
C8613 VDD.n2211 VSS 4.31e-19
C8614 VDD.n2212 VSS 1.59e-19
C8615 VDD.n2213 VSS 2.64e-19
C8616 VDD.n2214 VSS 1.59e-19
C8617 VDD.n2215 VSS 4.72e-19
C8618 VDD.n2216 VSS 0.00541f
C8619 VDD.n2217 VSS 5.05e-19
C8620 VDD.n2218 VSS 8.03e-19
C8621 VDD.n2219 VSS 2.64e-19
C8622 VDD.n2220 VSS 1.59e-19
C8623 VDD.n2221 VSS 1.59e-19
C8624 VDD.n2222 VSS 4.18e-19
C8625 VDD.n2223 VSS 9.34e-20
C8626 VDD.n2224 VSS 0.002f
C8627 VDD.n2225 VSS 5e-19
C8628 VDD.n2226 VSS 3e-19
C8629 VDD.n2227 VSS 0.00118f
C8630 VDD.t453 VSS 5.02e-19
C8631 VDD.t256 VSS 3.94e-19
C8632 VDD.n2228 VSS 0.00103f
C8633 VDD.n2229 VSS 1.59e-19
C8634 VDD.n2230 VSS 9.34e-20
C8635 VDD.t452 VSS 0.00441f
C8636 VDD.n2231 VSS 4.18e-19
C8637 VDD.n2232 VSS 1.59e-19
C8638 VDD.n2233 VSS 0.00141f
C8639 VDD.n2234 VSS 3e-19
C8640 VDD.n2235 VSS 5e-19
C8641 VDD.n2236 VSS 1e-18
C8642 VDD.n2237 VSS 9.34e-20
C8643 VDD.n2238 VSS 1.59e-19
C8644 VDD.n2239 VSS 1.59e-19
C8645 VDD.n2240 VSS 2.64e-19
C8646 VDD.n2241 VSS 1.59e-19
C8647 VDD.n2242 VSS 4.18e-19
C8648 VDD.n2243 VSS 0.00282f
C8649 VDD.n2244 VSS 5e-19
C8650 VDD.n2245 VSS 3e-19
C8651 VDD.n2246 VSS 0.00118f
C8652 VDD.n2247 VSS 1.59e-19
C8653 VDD.n2248 VSS 9.34e-20
C8654 VDD.t684 VSS 0.00441f
C8655 VDD.n2249 VSS 4.18e-19
C8656 VDD.n2250 VSS 1.59e-19
C8657 VDD.n2251 VSS 0.00141f
C8658 VDD.n2252 VSS 3e-19
C8659 VDD.n2253 VSS 5e-19
C8660 VDD.n2254 VSS 0.00516f
C8661 VDD.n2255 VSS 9.34e-20
C8662 VDD.n2256 VSS 1.59e-19
C8663 VDD.t685 VSS 7.16e-19
C8664 VDD.t213 VSS 2.33e-19
C8665 VDD.n2257 VSS 0.00366f
C8666 VDD.n2258 VSS 1.59e-19
C8667 VDD.n2259 VSS 0.00824f
C8668 VDD.n2260 VSS 2.64e-19
C8669 VDD.n2261 VSS 0.00115f
C8670 VDD.n2262 VSS 1.87e-20
C8671 VDD.n2263 VSS 0.00253f
C8672 VDD.n2264 VSS 5.44e-19
C8673 VDD.n2265 VSS 4.18e-19
C8674 VDD.n2266 VSS 0.00427f
C8675 VDD.t212 VSS 0.00171f
C8676 VDD.n2267 VSS 0.00365f
C8677 VDD.n2268 VSS 0.00194f
C8678 VDD.n2269 VSS 1e-18
C8679 VDD.n2270 VSS 9.34e-20
C8680 VDD.n2271 VSS 1.59e-19
C8681 VDD.n2272 VSS 5.53e-19
C8682 VDD.n2273 VSS 5.53e-19
C8683 VDD.n2274 VSS 0.00118f
C8684 VDD.n2275 VSS 2.64e-19
C8685 VDD.n2276 VSS 0.00141f
C8686 VDD.n2277 VSS 3e-19
C8687 VDD.n2278 VSS 5e-19
C8688 VDD.n2279 VSS 0.00347f
C8689 VDD.n2280 VSS 1e-18
C8690 VDD.t473 VSS 0.00441f
C8691 VDD.n2281 VSS 0.00259f
C8692 VDD.n2282 VSS 4.18e-19
C8693 VDD.n2283 VSS 5.53e-19
C8694 VDD.n2284 VSS 5.53e-19
C8695 VDD.n2285 VSS 1.59e-19
C8696 VDD.n2286 VSS 2.64e-19
C8697 VDD.n2287 VSS 0.00141f
C8698 VDD.n2288 VSS 0.00118f
C8699 VDD.n2289 VSS 5.53e-19
C8700 VDD.n2290 VSS 5.53e-19
C8701 VDD.n2291 VSS 1.59e-19
C8702 VDD.n2292 VSS 9.34e-20
C8703 VDD.n2293 VSS 1e-18
C8704 VDD.n2294 VSS 0.00447f
C8705 VDD.n2295 VSS 0.00535f
C8706 VDD.n2296 VSS 5e-19
C8707 VDD.n2297 VSS 3e-19
C8708 VDD.n2298 VSS 0.00141f
C8709 VDD.n2299 VSS 2.64e-19
C8710 VDD.n2300 VSS 0.00118f
C8711 VDD.n2301 VSS 5.53e-19
C8712 VDD.n2302 VSS 5.53e-19
C8713 VDD.n2303 VSS 4.18e-19
C8714 VDD.n2304 VSS 0.00435f
C8715 VDD.t37 VSS 0.00441f
C8716 VDD.n2305 VSS 0.00106f
C8717 VDD.n2306 VSS 0.00318f
C8718 VDD.n2307 VSS 1e-18
C8719 VDD.n2308 VSS 9.34e-20
C8720 VDD.n2309 VSS 1.59e-19
C8721 VDD.n2310 VSS 5.53e-19
C8722 VDD.n2311 VSS 5.53e-19
C8723 VDD.n2312 VSS 0.00118f
C8724 VDD.n2313 VSS 2.64e-19
C8725 VDD.n2314 VSS 0.00141f
C8726 VDD.n2315 VSS 3e-19
C8727 VDD.n2316 VSS 5e-19
C8728 VDD.n2317 VSS 0.00224f
C8729 VDD.n2318 VSS 1e-18
C8730 VDD.t255 VSS 0.00441f
C8731 VDD.n2319 VSS 0.00341f
C8732 VDD.n2320 VSS 4.18e-19
C8733 VDD.n2321 VSS 1.31e-19
C8734 VDD.n2322 VSS 0.00208f
C8735 VDD.n2323 VSS 4.31e-19
C8736 VDD.n2324 VSS 1.59e-19
C8737 VDD.n2325 VSS 2.64e-19
C8738 VDD.n2326 VSS 0.00141f
C8739 VDD.n2327 VSS 0.00118f
C8740 VDD.n2328 VSS 5.53e-19
C8741 VDD.n2329 VSS 5.53e-19
C8742 VDD.n2330 VSS 1.59e-19
C8743 VDD.n2331 VSS 9.34e-20
C8744 VDD.n2332 VSS 1e-18
C8745 VDD.n2333 VSS 0.00447f
C8746 VDD.n2334 VSS 0.0108f
C8747 VDD.n2335 VSS 0.00101f
C8748 VDD.n2336 VSS 0.00146f
C8749 VDD.n2337 VSS 0.00101f
C8750 VDD.n2338 VSS 0.0108f
C8751 VDD.n2339 VSS 0.00101f
C8752 VDD.n2340 VSS 0.0105f
C8753 VDD.n2341 VSS 9.78e-19
C8754 VDD.n2342 VSS 0.0014f
C8755 VDD.n2343 VSS 0.00146f
C8756 VDD.n2344 VSS 0.00146f
C8757 VDD.n2345 VSS 0.00101f
C8758 VDD.n2346 VSS 0.0108f
C8759 VDD.n2347 VSS 0.0108f
C8760 VDD.n2348 VSS 0.0108f
C8761 VDD.n2349 VSS 0.00101f
C8762 VDD.n2350 VSS 0.00146f
C8763 VDD.n2351 VSS 0.00144f
C8764 VDD.n2352 VSS 7.79e-19
C8765 VDD.n2353 VSS 5.05e-19
C8766 VDD.n2354 VSS 0.00541f
C8767 VDD.n2355 VSS 1e-18
C8768 VDD.n2356 VSS 0.00535f
C8769 VDD.n2357 VSS 5e-19
C8770 VDD.n2358 VSS 3e-19
C8771 VDD.n2359 VSS 7.14e-19
C8772 VDD.n2360 VSS 0.0101f
C8773 VDD.n2361 VSS 2.06e-19
C8774 VDD.n2362 VSS 1.59e-19
C8775 VDD.n2363 VSS 9.34e-20
C8776 VDD.n2364 VSS 1e-18
C8777 VDD.n2365 VSS 0.00506f
C8778 VDD.n2366 VSS 0.00476f
C8779 VDD.n2367 VSS 4.45e-19
C8780 VDD.n2368 VSS 6e-19
C8781 VDD.n2369 VSS 6e-19
C8782 VDD.n2370 VSS 0.00126f
C8783 VDD.n2371 VSS 2.64e-19
C8784 VDD.n2372 VSS 0.00133f
C8785 VDD.n2373 VSS 2.06e-19
C8786 VDD.n2374 VSS 4.72e-19
C8787 VDD.n2375 VSS 0.00141f
C8788 VDD.t14 VSS 0.00441f
C8789 VDD.n2376 VSS 0.004f
C8790 VDD.n2377 VSS 0.00165f
C8791 VDD.n2378 VSS 1e-18
C8792 VDD.n2379 VSS 9.34e-20
C8793 VDD.n2380 VSS 1.59e-19
C8794 VDD.n2381 VSS 2.06e-19
C8795 VDD.n2382 VSS 0.00133f
C8796 VDD.n2383 VSS 2.64e-19
C8797 VDD.n2384 VSS 0.00126f
C8798 VDD.n2385 VSS 6e-19
C8799 VDD.n2386 VSS 6e-19
C8800 VDD.n2387 VSS 4.45e-19
C8801 VDD.n2388 VSS 0.00376f
C8802 VDD.n2389 VSS 8.23e-19
C8803 VDD.t350 VSS 6.47e-19
C8804 VDD.n2390 VSS 0.00459f
C8805 VDD.n2391 VSS 4.72e-19
C8806 VDD.n2392 VSS 2.06e-19
C8807 VDD.n2393 VSS 1.59e-19
C8808 VDD.n2394 VSS 6e-19
C8809 VDD.n2395 VSS 0.00126f
C8810 VDD.n2396 VSS 0.00133f
C8811 VDD.n2397 VSS 2.06e-19
C8812 VDD.n2398 VSS 1.59e-19
C8813 VDD.n2399 VSS 9.34e-20
C8814 VDD.n2400 VSS 1e-18
C8815 VDD.n2401 VSS 0.00506f
C8816 VDD.n2402 VSS 0.00476f
C8817 VDD.n2403 VSS 4.45e-19
C8818 VDD.n2404 VSS 6e-19
C8819 VDD.n2405 VSS 6e-19
C8820 VDD.n2406 VSS 0.00126f
C8821 VDD.n2407 VSS 2.64e-19
C8822 VDD.n2408 VSS 0.00133f
C8823 VDD.n2409 VSS 2.06e-19
C8824 VDD.n2410 VSS 4.72e-19
C8825 VDD.n2411 VSS 0.00224f
C8826 VDD.t466 VSS 0.00441f
C8827 VDD.n2412 VSS 0.00318f
C8828 VDD.n2413 VSS 0.00288f
C8829 VDD.n2414 VSS 1e-18
C8830 VDD.n2415 VSS 9.34e-20
C8831 VDD.n2416 VSS 1.59e-19
C8832 VDD.n2417 VSS 2.06e-19
C8833 VDD.n2418 VSS 0.00133f
C8834 VDD.n2419 VSS 2.64e-19
C8835 VDD.n2420 VSS 0.00126f
C8836 VDD.n2421 VSS 6e-19
C8837 VDD.n2422 VSS 6e-19
C8838 VDD.n2423 VSS 4.45e-19
C8839 VDD.n2424 VSS 0.00253f
C8840 VDD.n2425 VSS 1e-18
C8841 VDD.t623 VSS 0.00441f
C8842 VDD.n2426 VSS 0.00388f
C8843 VDD.n2427 VSS 4.72e-19
C8844 VDD.n2428 VSS 2.06e-19
C8845 VDD.n2429 VSS 1.22e-19
C8846 VDD.n2430 VSS 0.00205f
C8847 VDD.n2431 VSS 5.81e-19
C8848 VDD.n2432 VSS 0.00126f
C8849 VDD.n2433 VSS 2.48e-19
C8850 VDD.n2434 VSS 2.64e-19
C8851 VDD.n2435 VSS 0.00133f
C8852 VDD.n2436 VSS 2.06e-19
C8853 VDD.n2437 VSS 1.59e-19
C8854 VDD.n2438 VSS 9.34e-20
C8855 VDD.n2439 VSS 1e-18
C8856 VDD.n2440 VSS 0.00541f
C8857 VDD.n2441 VSS 0.0102f
C8858 VDD.n2442 VSS 9.5e-19
C8859 VDD.n2443 VSS 0.00125f
C8860 VDD.n2444 VSS 0.00123f
C8861 VDD.n2445 VSS 5.93e-19
C8862 VDD.n2446 VSS 0.00276f
C8863 VDD.n2447 VSS 2.64e-19
C8864 VDD.n2448 VSS 2.79e-19
C8865 VDD.n2449 VSS 2.81e-19
C8866 VDD.n2450 VSS 5.05e-19
C8867 VDD.n2451 VSS 0.00541f
C8868 VDD.n2452 VSS 1e-18
C8869 VDD.t187 VSS 0.00176f
C8870 VDD.n2453 VSS 0.00106f
C8871 VDD.n2454 VSS 4.23e-19
C8872 VDD.n2455 VSS 5.62e-19
C8873 VDD.n2456 VSS 0.00255f
C8874 VDD.n2457 VSS 1.59e-19
C8875 VDD.n2458 VSS 2.64e-19
C8876 VDD.n2459 VSS 0.0014f
C8877 VDD.n2460 VSS 0.00119f
C8878 VDD.n2461 VSS 5.62e-19
C8879 VDD.n2462 VSS 5.62e-19
C8880 VDD.n2463 VSS 1.59e-19
C8881 VDD.n2464 VSS 9.34e-20
C8882 VDD.n2465 VSS 1e-18
C8883 VDD.n2466 VSS 0.00206f
C8884 VDD.t378 VSS 0.00441f
C8885 VDD.n2467 VSS 0.00335f
C8886 VDD.n2468 VSS 4.94e-19
C8887 VDD.n2469 VSS 2.81e-19
C8888 VDD.n2470 VSS 0.0014f
C8889 VDD.n2471 VSS 2.64e-19
C8890 VDD.n2472 VSS 0.00119f
C8891 VDD.n2473 VSS 5.62e-19
C8892 VDD.n2474 VSS 5.62e-19
C8893 VDD.n2475 VSS 4.23e-19
C8894 VDD.n2476 VSS 0.00271f
C8895 VDD.t470 VSS 0.00441f
C8896 VDD.n2477 VSS 0.00271f
C8897 VDD.n2478 VSS 1e-18
C8898 VDD.n2479 VSS 9.34e-20
C8899 VDD.n2480 VSS 1.59e-19
C8900 VDD.n2481 VSS 5.62e-19
C8901 VDD.n2482 VSS 5.62e-19
C8902 VDD.n2483 VSS 0.00119f
C8903 VDD.n2484 VSS 2.64e-19
C8904 VDD.n2485 VSS 0.0014f
C8905 VDD.n2486 VSS 2.81e-19
C8906 VDD.n2487 VSS 4.94e-19
C8907 VDD.n2488 VSS 0.00529f
C8908 VDD.n2489 VSS 1e-18
C8909 VDD.t627 VSS 0.00441f
C8910 VDD.n2490 VSS 0.00447f
C8911 VDD.n2491 VSS 4.23e-19
C8912 VDD.n2492 VSS 5.62e-19
C8913 VDD.n2493 VSS 5.62e-19
C8914 VDD.n2494 VSS 1.59e-19
C8915 VDD.n2495 VSS 2.64e-19
C8916 VDD.n2496 VSS 0.0014f
C8917 VDD.n2497 VSS 0.00119f
C8918 VDD.n2498 VSS 5.62e-19
C8919 VDD.n2499 VSS 5.62e-19
C8920 VDD.n2500 VSS 1.59e-19
C8921 VDD.n2501 VSS 9.34e-20
C8922 VDD.n2502 VSS 1e-18
C8923 VDD.n2503 VSS 0.00329f
C8924 VDD.t102 VSS 0.00441f
C8925 VDD.n2504 VSS 0.00212f
C8926 VDD.n2505 VSS 4.94e-19
C8927 VDD.n2506 VSS 2.81e-19
C8928 VDD.n2507 VSS 0.0014f
C8929 VDD.n2508 VSS 2.64e-19
C8930 VDD.n2509 VSS 0.00119f
C8931 VDD.n2510 VSS 4.31e-19
C8932 VDD.n2511 VSS 0.00208f
C8933 VDD.n2512 VSS 1.5e-19
C8934 VDD.n2513 VSS 4.23e-19
C8935 VDD.n2514 VSS 0.00353f
C8936 VDD.t659 VSS 0.00441f
C8937 VDD.n2515 VSS 0.00188f
C8938 VDD.n2516 VSS 1e-18
C8939 VDD.n2517 VSS 9.34e-20
C8940 VDD.n2518 VSS 1.59e-19
C8941 VDD.n2519 VSS 5.62e-19
C8942 VDD.n2520 VSS 5.62e-19
C8943 VDD.n2521 VSS 0.00119f
C8944 VDD.n2522 VSS 2.64e-19
C8945 VDD.n2523 VSS 7.14e-19
C8946 VDD.n2524 VSS 2.81e-19
C8947 VDD.n2525 VSS 4.94e-19
C8948 VDD.n2526 VSS 0.00529f
C8949 VDD.n2527 VSS 1e-18
C8950 VDD.n2528 VSS 0.00541f
C8951 VDD.n2529 VSS 5.05e-19
C8952 VDD.n2530 VSS 7.84e-19
C8953 VDD.n2531 VSS 0.00143f
C8954 VDD.n2532 VSS 0.00146f
C8955 VDD.n2533 VSS 0.00101f
C8956 VDD.n2534 VSS 0.0108f
C8957 VDD.n2535 VSS 0.0108f
C8958 VDD.n2536 VSS 0.0108f
C8959 VDD.n2537 VSS 0.00101f
C8960 VDD.n2538 VSS 0.00146f
C8961 VDD.n2539 VSS 0.00146f
C8962 VDD.n2540 VSS 0.0014f
C8963 VDD.n2541 VSS 9.78e-19
C8964 VDD.n2542 VSS 0.0105f
C8965 VDD.n2543 VSS 0.00541f
C8966 VDD.n2544 VSS 1e-18
C8967 VDD.n2545 VSS 9.34e-20
C8968 VDD.n2546 VSS 1.59e-19
C8969 VDD.n2547 VSS 2.06e-19
C8970 VDD.n2548 VSS 0.0101f
C8971 VDD.n2549 VSS 2.64e-19
C8972 VDD.n2550 VSS 0.00126f
C8973 VDD.n2551 VSS 6e-19
C8974 VDD.n2552 VSS 6e-19
C8975 VDD.n2553 VSS 4.45e-19
C8976 VDD.n2554 VSS 0.00476f
C8977 VDD.n2555 VSS 1e-18
C8978 VDD.t374 VSS 0.00441f
C8979 VDD.n2556 VSS 0.00141f
C8980 VDD.n2557 VSS 4.72e-19
C8981 VDD.n2558 VSS 2.06e-19
C8982 VDD.n2559 VSS 1.59e-19
C8983 VDD.t375 VSS 3.94e-19
C8984 VDD.t455 VSS 5.02e-19
C8985 VDD.n2560 VSS 0.00103f
C8986 VDD.n2561 VSS 0.00208f
C8987 VDD.n2562 VSS 4.31e-19
C8988 VDD.n2563 VSS 0.00126f
C8989 VDD.n2564 VSS 0.00133f
C8990 VDD.n2565 VSS 2.06e-19
C8991 VDD.n2566 VSS 1.59e-19
C8992 VDD.n2567 VSS 9.34e-20
C8993 VDD.n2568 VSS 1e-18
C8994 VDD.n2569 VSS 0.00165f
C8995 VDD.t454 VSS 0.00441f
C8996 VDD.n2570 VSS 8.23e-19
C8997 VDD.n2571 VSS 0.00376f
C8998 VDD.n2572 VSS 4.45e-19
C8999 VDD.n2573 VSS 6e-19
C9000 VDD.n2574 VSS 6e-19
C9001 VDD.n2575 VSS 0.00126f
C9002 VDD.n2576 VSS 2.64e-19
C9003 VDD.n2577 VSS 0.00133f
C9004 VDD.n2578 VSS 2.06e-19
C9005 VDD.n2579 VSS 4.72e-19
C9006 VDD.n2580 VSS 0.00459f
C9007 VDD.n2581 VSS 0.00476f
C9008 VDD.n2582 VSS 1e-18
C9009 VDD.n2583 VSS 9.34e-20
C9010 VDD.n2584 VSS 1.59e-19
C9011 VDD.n2585 VSS 2.06e-19
C9012 VDD.n2586 VSS 0.00133f
C9013 VDD.n2587 VSS 2.64e-19
C9014 VDD.n2588 VSS 0.00126f
C9015 VDD.n2589 VSS 6e-19
C9016 VDD.n2590 VSS 6e-19
C9017 VDD.n2591 VSS 4.45e-19
C9018 VDD.n2592 VSS 0.00476f
C9019 VDD.n2593 VSS 1e-18
C9020 VDD.t471 VSS 0.00441f
C9021 VDD.n2594 VSS 0.00224f
C9022 VDD.n2595 VSS 4.72e-19
C9023 VDD.n2596 VSS 2.06e-19
C9024 VDD.n2597 VSS 1.59e-19
C9025 VDD.n2598 VSS 6e-19
C9026 VDD.n2599 VSS 0.00126f
C9027 VDD.n2600 VSS 0.00133f
C9028 VDD.n2601 VSS 2.06e-19
C9029 VDD.n2602 VSS 1.59e-19
C9030 VDD.n2603 VSS 9.34e-20
C9031 VDD.n2604 VSS 1e-18
C9032 VDD.n2605 VSS 0.00288f
C9033 VDD.t124 VSS 0.00441f
C9034 VDD.n2606 VSS 0.00388f
C9035 VDD.n2607 VSS 1e-18
C9036 VDD.n2608 VSS 0.00253f
C9037 VDD.n2609 VSS 4.45e-19
C9038 VDD.n2610 VSS 6e-19
C9039 VDD.n2611 VSS 6e-19
C9040 VDD.n2612 VSS 0.00126f
C9041 VDD.n2613 VSS 0.00133f
C9042 VDD.n2614 VSS 2.64e-19
C9043 VDD.n2615 VSS 1.22e-19
C9044 VDD.n2616 VSS 0.00205f
C9045 VDD.n2617 VSS 5.81e-19
C9046 VDD.n2618 VSS 6e-19
C9047 VDD.n2619 VSS 4.45e-19
C9048 VDD.n2620 VSS 1e-18
C9049 VDD.n2621 VSS 0.00906f
C9050 VDD.n2622 VSS 8e-19
C9051 VDD.n2623 VSS 2.06e-19
C9052 VDD.n2624 VSS 0.00133f
C9053 VDD.n2625 VSS 2.64e-19
C9054 VDD.n2626 VSS 2.48e-19
C9055 VDD.n2627 VSS 0.00119f
C9056 VDD.n2628 VSS 0.00156f
C9057 VDD.n2629 VSS 8.31e-19
C9058 VDD.n2630 VSS 0.00273f
C9059 VDD.n2631 VSS 2.64e-19
C9060 VDD.n2632 VSS 2.79e-19
C9061 VDD.n2633 VSS 1.87e-20
C9062 VDD.n2634 VSS 5.05e-19
C9063 VDD.n2635 VSS 0.00541f
C9064 VDD.n2636 VSS 1e-18
C9065 VDD.t276 VSS 0.00259f
C9066 VDD.n2637 VSS 0.00271f
C9067 VDD.n2638 VSS 5e-19
C9068 VDD.n2639 VSS 6.94e-19
C9069 VDD.n2640 VSS 6.75e-19
C9070 VDD.n2641 VSS 0.00214f
C9071 VDD.n2642 VSS 2.81e-20
C9072 VDD.n2643 VSS 2.64e-19
C9073 VDD.n2644 VSS 0.00118f
C9074 VDD.n2645 VSS 0.00141f
C9075 VDD.n2646 VSS 6.94e-19
C9076 VDD.n2647 VSS 6.94e-19
C9077 VDD.n2648 VSS 1.59e-19
C9078 VDD.n2649 VSS 9.34e-20
C9079 VDD.n2650 VSS 1e-18
C9080 VDD.n2651 VSS 0.00371f
C9081 VDD.t488 VSS 0.00441f
C9082 VDD.n2652 VSS 0.00171f
C9083 VDD.n2653 VSS 4.18e-19
C9084 VDD.n2654 VSS 1.87e-20
C9085 VDD.n2655 VSS 0.00118f
C9086 VDD.n2656 VSS 2.64e-19
C9087 VDD.n2657 VSS 0.00141f
C9088 VDD.n2658 VSS 6.94e-19
C9089 VDD.n2659 VSS 6.94e-19
C9090 VDD.n2660 VSS 5e-19
C9091 VDD.n2661 VSS 0.00435f
C9092 VDD.t475 VSS 0.00441f
C9093 VDD.n2662 VSS 0.00106f
C9094 VDD.n2663 VSS 1e-18
C9095 VDD.n2664 VSS 9.34e-20
C9096 VDD.n2665 VSS 1.59e-19
C9097 VDD.n2666 VSS 6.94e-19
C9098 VDD.n2667 VSS 6.94e-19
C9099 VDD.n2668 VSS 0.00141f
C9100 VDD.n2669 VSS 2.64e-19
C9101 VDD.n2670 VSS 0.00118f
C9102 VDD.n2671 VSS 1.87e-20
C9103 VDD.n2672 VSS 4.18e-19
C9104 VDD.n2673 VSS 0.00447f
C9105 VDD.n2674 VSS 1e-18
C9106 VDD.n2675 VSS 0.00535f
C9107 VDD.n2676 VSS 5e-19
C9108 VDD.n2677 VSS 6.94e-19
C9109 VDD.n2678 VSS 6.94e-19
C9110 VDD.n2679 VSS 1.59e-19
C9111 VDD.n2680 VSS 2.64e-19
C9112 VDD.n2681 VSS 0.00118f
C9113 VDD.n2682 VSS 0.00141f
C9114 VDD.n2683 VSS 6.94e-19
C9115 VDD.n2684 VSS 6.94e-19
C9116 VDD.n2685 VSS 1.59e-19
C9117 VDD.n2686 VSS 9.34e-20
C9118 VDD.n2687 VSS 7.65e-19
C9119 VDD.t272 VSS 9.41e-19
C9120 VDD.n2688 VSS 0.00424f
C9121 VDD.t301 VSS 0.00441f
C9122 VDD.n2689 VSS 4.71e-19
C9123 VDD.n2690 VSS 4.18e-19
C9124 VDD.n2691 VSS 1.87e-20
C9125 VDD.n2692 VSS 0.00118f
C9126 VDD.n2693 VSS 2.64e-19
C9127 VDD.n2694 VSS 0.00141f
C9128 VDD.n2695 VSS 4.31e-19
C9129 VDD.n2696 VSS 0.00208f
C9130 VDD.n2697 VSS 4.12e-19
C9131 VDD.n2698 VSS 5e-19
C9132 VDD.n2699 VSS 0.00518f
C9133 VDD.t161 VSS 0.00441f
C9134 VDD.n2700 VSS 2.35e-19
C9135 VDD.n2701 VSS 1e-18
C9136 VDD.n2702 VSS 9.34e-20
C9137 VDD.n2703 VSS 1.59e-19
C9138 VDD.n2704 VSS 6.94e-19
C9139 VDD.n2705 VSS 6.94e-19
C9140 VDD.n2706 VSS 0.00141f
C9141 VDD.n2707 VSS 2.64e-19
C9142 VDD.n2708 VSS 7.14e-19
C9143 VDD.n2709 VSS 1.87e-20
C9144 VDD.n2710 VSS 4.18e-19
C9145 VDD.n2711 VSS 0.00447f
C9146 VDD.n2712 VSS 1e-18
C9147 VDD.n2713 VSS 0.00541f
C9148 VDD.n2714 VSS 5.05e-19
C9149 VDD.n2715 VSS 8.43e-19
C9150 VDD.n2716 VSS 0.00132f
C9151 VDD.n2717 VSS 0.00146f
C9152 VDD.n2718 VSS 0.00101f
C9153 VDD.n2719 VSS 0.0108f
C9154 VDD.n2720 VSS 0.0108f
C9155 VDD.n2721 VSS 0.0108f
C9156 VDD.n2722 VSS 0.00101f
C9157 VDD.n2723 VSS 0.00146f
C9158 VDD.n2724 VSS 0.00146f
C9159 VDD.n2725 VSS 0.00119f
C9160 VDD.n2726 VSS 0.00146f
C9161 VDD.n2727 VSS 0.00101f
C9162 VDD.n2728 VSS 0.0108f
C9163 VDD.n2729 VSS 0.0108f
C9164 VDD.n2730 VSS 0.00565f
C9165 VDD.t76 VSS 0.00541f
C9166 VDD.n2731 VSS 0.00859f
C9167 VDD.n2732 VSS 0.00101f
C9168 VDD.n2733 VSS 8.62e-19
C9169 VDD.t77 VSS 3.94e-19
C9170 VDD.t440 VSS 5.02e-19
C9171 VDD.n2734 VSS 0.00103f
C9172 VDD.n2735 VSS 0.00202f
C9173 VDD.n2736 VSS 4.31e-19
C9174 VDD.n2737 VSS 8.62e-19
C9175 VDD.n2738 VSS 0.00285f
C9176 VDD.n2739 VSS 0.00285f
C9177 VDD.n2740 VSS 0.00285f
C9178 VDD.n2741 VSS 8.62e-19
C9179 VDD.n2742 VSS 8.62e-19
C9180 VDD.n2743 VSS 0.00101f
C9181 VDD.n2744 VSS 0.00424f
C9182 VDD.t38 VSS 0.00541f
C9183 VDD.n2745 VSS 0.00859f
C9184 VDD.n2746 VSS 0.00606f
C9185 VDD.t472 VSS 0.00541f
C9186 VDD.n2747 VSS 0.00941f
C9187 VDD.n2748 VSS 0.00101f
C9188 VDD.n2749 VSS 8.62e-19
C9189 VDD.n2750 VSS 8.62e-19
C9190 VDD.n2751 VSS 8.62e-19
C9191 VDD.n2752 VSS 0.00285f
C9192 VDD.n2753 VSS 0.00285f
C9193 VDD.n2754 VSS 0.00168f
C9194 VDD.n2755 VSS 0.00285f
C9195 VDD.n2756 VSS 5.06e-19
C9196 VDD.n2757 VSS 8.62e-19
C9197 VDD.n2758 VSS 0.00101f
C9198 VDD.n2759 VSS 0.00618f
C9199 VDD.n2760 VSS 0.00565f
C9200 VDD.t286 VSS 0.00141f
C9201 VDD.n2761 VSS 0.00941f
C9202 VDD.n2762 VSS 0.00101f
C9203 VDD.n2763 VSS 0.00113f
C9204 VDD.n2764 VSS 0.0013f
C9205 VDD.n2765 VSS 8.31e-19
C9206 VDD.n2766 VSS 0.00273f
C9207 VDD.n2767 VSS 2.64e-19
C9208 VDD.n2768 VSS 2.79e-19
C9209 VDD.n2769 VSS 1.87e-20
C9210 VDD.n2770 VSS 5.05e-19
C9211 VDD.n2771 VSS 0.00541f
C9212 VDD.n2772 VSS 1e-18
C9213 VDD.t23 VSS 0.00259f
C9214 VDD.n2773 VSS 0.00271f
C9215 VDD.n2774 VSS 5e-19
C9216 VDD.n2775 VSS 6.94e-19
C9217 VDD.n2776 VSS 6.75e-19
C9218 VDD.n2777 VSS 0.00214f
C9219 VDD.n2778 VSS 2.81e-20
C9220 VDD.n2779 VSS 2.64e-19
C9221 VDD.n2780 VSS 0.00118f
C9222 VDD.n2781 VSS 0.00141f
C9223 VDD.n2782 VSS 6.94e-19
C9224 VDD.n2783 VSS 6.94e-19
C9225 VDD.n2784 VSS 1.59e-19
C9226 VDD.n2785 VSS 9.34e-20
C9227 VDD.n2786 VSS 1e-18
C9228 VDD.n2787 VSS 0.00371f
C9229 VDD.t132 VSS 0.00441f
C9230 VDD.n2788 VSS 0.00171f
C9231 VDD.n2789 VSS 4.18e-19
C9232 VDD.n2790 VSS 1.87e-20
C9233 VDD.n2791 VSS 0.00118f
C9234 VDD.n2792 VSS 2.64e-19
C9235 VDD.n2793 VSS 0.00141f
C9236 VDD.n2794 VSS 6.94e-19
C9237 VDD.n2795 VSS 6.94e-19
C9238 VDD.n2796 VSS 5e-19
C9239 VDD.n2797 VSS 0.00435f
C9240 VDD.t468 VSS 0.00441f
C9241 VDD.n2798 VSS 0.00106f
C9242 VDD.n2799 VSS 1e-18
C9243 VDD.n2800 VSS 9.34e-20
C9244 VDD.n2801 VSS 1.59e-19
C9245 VDD.n2802 VSS 6.94e-19
C9246 VDD.n2803 VSS 6.94e-19
C9247 VDD.n2804 VSS 0.00141f
C9248 VDD.n2805 VSS 2.64e-19
C9249 VDD.n2806 VSS 0.00118f
C9250 VDD.n2807 VSS 1.87e-20
C9251 VDD.n2808 VSS 4.18e-19
C9252 VDD.n2809 VSS 0.00447f
C9253 VDD.n2810 VSS 1e-18
C9254 VDD.n2811 VSS 0.00535f
C9255 VDD.n2812 VSS 5e-19
C9256 VDD.n2813 VSS 6.94e-19
C9257 VDD.n2814 VSS 6.94e-19
C9258 VDD.n2815 VSS 1.59e-19
C9259 VDD.n2816 VSS 2.64e-19
C9260 VDD.n2817 VSS 0.00118f
C9261 VDD.n2818 VSS 0.00141f
C9262 VDD.n2819 VSS 6.94e-19
C9263 VDD.n2820 VSS 6.94e-19
C9264 VDD.n2821 VSS 1.59e-19
C9265 VDD.n2822 VSS 9.34e-20
C9266 VDD.n2823 VSS 7.65e-19
C9267 VDD.t351 VSS 9.41e-19
C9268 VDD.n2824 VSS 0.00424f
C9269 VDD.t321 VSS 0.00441f
C9270 VDD.n2825 VSS 4.71e-19
C9271 VDD.n2826 VSS 4.18e-19
C9272 VDD.n2827 VSS 1.87e-20
C9273 VDD.n2828 VSS 0.00118f
C9274 VDD.n2829 VSS 2.64e-19
C9275 VDD.n2830 VSS 0.00141f
C9276 VDD.n2831 VSS 4.31e-19
C9277 VDD.n2832 VSS 0.00208f
C9278 VDD.n2833 VSS 4.12e-19
C9279 VDD.n2834 VSS 5e-19
C9280 VDD.n2835 VSS 0.00518f
C9281 VDD.t384 VSS 0.00441f
C9282 VDD.n2836 VSS 2.35e-19
C9283 VDD.n2837 VSS 1e-18
C9284 VDD.n2838 VSS 9.34e-20
C9285 VDD.n2839 VSS 1.59e-19
C9286 VDD.n2840 VSS 6.94e-19
C9287 VDD.n2841 VSS 6.94e-19
C9288 VDD.n2842 VSS 0.00141f
C9289 VDD.n2843 VSS 2.64e-19
C9290 VDD.n2844 VSS 7.14e-19
C9291 VDD.n2845 VSS 1.87e-20
C9292 VDD.n2846 VSS 4.18e-19
C9293 VDD.n2847 VSS 0.00447f
C9294 VDD.n2848 VSS 1e-18
C9295 VDD.n2849 VSS 0.00541f
C9296 VDD.n2850 VSS 5.05e-19
C9297 VDD.n2851 VSS 8.43e-19
C9298 VDD.n2852 VSS 0.00132f
C9299 VDD.n2853 VSS 0.00146f
C9300 VDD.n2854 VSS 0.00101f
C9301 VDD.n2855 VSS 0.0108f
C9302 VDD.n2856 VSS 0.0108f
C9303 VDD.n2857 VSS 0.0108f
C9304 VDD.n2858 VSS 0.00101f
C9305 VDD.n2859 VSS 0.00146f
C9306 VDD.n2860 VSS 0.00146f
C9307 VDD.n2861 VSS 0.00119f
C9308 VDD.n2862 VSS 0.00146f
C9309 VDD.n2863 VSS 0.00101f
C9310 VDD.n2864 VSS 0.0108f
C9311 VDD.n2865 VSS 0.0108f
C9312 VDD.n2866 VSS 0.00565f
C9313 VDD.t267 VSS 0.00541f
C9314 VDD.n2867 VSS 0.00859f
C9315 VDD.n2868 VSS 0.00101f
C9316 VDD.n2869 VSS 8.62e-19
C9317 VDD.t268 VSS 3.94e-19
C9318 VDD.t87 VSS 5.02e-19
C9319 VDD.n2870 VSS 0.00103f
C9320 VDD.n2871 VSS 0.00202f
C9321 VDD.n2872 VSS 4.31e-19
C9322 VDD.n2873 VSS 8.62e-19
C9323 VDD.n2874 VSS 0.00285f
C9324 VDD.n2875 VSS 0.00285f
C9325 VDD.n2876 VSS 0.00285f
C9326 VDD.n2877 VSS 8.62e-19
C9327 VDD.n2878 VSS 8.62e-19
C9328 VDD.n2879 VSS 0.00101f
C9329 VDD.n2880 VSS 0.00424f
C9330 VDD.t134 VSS 0.00541f
C9331 VDD.n2881 VSS 0.00859f
C9332 VDD.n2882 VSS 0.00606f
C9333 VDD.t469 VSS 0.00541f
C9334 VDD.n2883 VSS 0.00941f
C9335 VDD.n2884 VSS 0.00101f
C9336 VDD.n2885 VSS 8.62e-19
C9337 VDD.n2886 VSS 8.62e-19
C9338 VDD.n2887 VSS 0.00285f
C9339 VDD.n2888 VSS 0.00285f
C9340 VDD.n2889 VSS 8.62e-19
C9341 VDD.t633 VSS 7.16e-19
C9342 VDD.t449 VSS 2.33e-19
C9343 VDD.n2890 VSS 0.00366f
C9344 VDD.n2891 VSS 0.00237f
C9345 VDD.n2892 VSS 5.06e-19
C9346 VDD.n2893 VSS 8.62e-19
C9347 VDD.n2894 VSS 0.00101f
C9348 VDD.n2895 VSS 0.00618f
C9349 VDD.n2896 VSS 0.00565f
C9350 VDD.t448 VSS 0.00141f
C9351 VDD.n2897 VSS 0.00941f
C9352 VDD.n2898 VSS 0.00101f
C9353 VDD.n2899 VSS 0.00113f
C9354 VDD.n2900 VSS 8.62e-19
C9355 VDD.n2901 VSS 0.00168f
C9356 VDD.n2902 VSS 0.00304f
C9357 VDD.n2903 VSS 0.00171f
C9358 VDD.n2904 VSS 0.00101f
C9359 VDD.n2905 VSS 0.00823f
C9360 VDD.t657 VSS 0.00365f
C9361 VDD.n2906 VSS 0.00559f
C9362 VDD.t677 VSS 0.00541f
C9363 VDD.t474 VSS 0.00541f
C9364 VDD.n2907 VSS 0.00606f
C9365 VDD.n2908 VSS 0.00101f
C9366 VDD.n2909 VSS 0.00172f
C9367 VDD.n2910 VSS 0.00285f
C9368 VDD.n2911 VSS 0.00285f
C9369 VDD.n2912 VSS 0.00285f
C9370 VDD.n2913 VSS 0.00172f
C9371 VDD.n2914 VSS 0.00101f
C9372 VDD.n2915 VSS 0.0108f
C9373 VDD.n2916 VSS 0.00623f
C9374 VDD.t461 VSS 0.00506f
C9375 VDD.t555 VSS 0.00459f
C9376 VDD.t425 VSS 0.00541f
C9377 VDD.n2917 VSS 0.00565f
C9378 VDD.n2918 VSS 0.00101f
C9379 VDD.n2919 VSS 0.00129f
C9380 VDD.n2920 VSS 0.00285f
C9381 VDD.n2921 VSS 0.00285f
C9382 VDD.n2922 VSS 0.00214f
C9383 VDD.n2923 VSS 0.00583f
C9384 VDD.n2924 VSS 0.00349f
C9385 VDD.n2925 VSS 0.0409f
C9386 VDD.n2926 VSS 0.0409f
C9387 VDD.n2927 VSS 0.00553f
C9388 VDD.n2928 VSS 0.0108f
C9389 VDD.n2929 VSS 0.00101f
C9390 VDD.n2930 VSS 0.00172f
C9391 VDD.n2931 VSS 0.00129f
C9392 VDD.n2932 VSS 0.00285f
C9393 VDD.n2933 VSS 0.00285f
C9394 VDD.n2934 VSS 0.00129f
C9395 VDD.n2935 VSS 0.00101f
C9396 VDD.n2936 VSS 0.00565f
C9397 VDD.t590 VSS 0.00459f
C9398 VDD.t273 VSS 0.00506f
C9399 VDD.n2937 VSS 0.00623f
C9400 VDD.n2938 VSS 0.00635f
C9401 VDD.n2939 VSS 0.0108f
C9402 VDD.n2940 VSS 0.00101f
C9403 VDD.n2941 VSS 0.00172f
C9404 VDD.n2942 VSS 0.00285f
C9405 VDD.n2943 VSS 0.00285f
C9406 VDD.n2944 VSS 0.00285f
C9407 VDD.n2945 VSS 0.00172f
C9408 VDD.n2946 VSS 0.00101f
C9409 VDD.n2947 VSS 0.00606f
C9410 VDD.t352 VSS 0.00541f
C9411 VDD.n2948 VSS 0.00641f
C9412 VDD.t446 VSS 0.00376f
C9413 VDD.n2949 VSS 0.0105f
C9414 VDD.n2950 VSS 0.0108f
C9415 VDD.n2951 VSS 0.00706f
C9416 VDD.n2952 VSS 0.00101f
C9417 VDD.n2953 VSS 0.00171f
C9418 VDD.n2954 VSS 0.00168f
C9419 VDD.n2955 VSS 0.00301f
C9420 VDD.n2956 VSS 0.00258f
C9421 VDD.n2957 VSS 5.25e-19
C9422 VDD.n2958 VSS 0.00235f
C9423 VDD.n2959 VSS 8.44e-19
C9424 VDD.n2960 VSS 0.00101f
C9425 VDD.n2961 VSS 8.23e-19
C9426 VDD.n2962 VSS 0.00559f
C9427 VDD.t486 VSS 0.00541f
C9428 VDD.t463 VSS 0.00541f
C9429 VDD.n2963 VSS 0.00606f
C9430 VDD.n2964 VSS 0.00101f
C9431 VDD.n2965 VSS 8.62e-19
C9432 VDD.n2966 VSS 8.62e-19
C9433 VDD.n2967 VSS 8.62e-19
C9434 VDD.n2968 VSS 0.00285f
C9435 VDD.n2969 VSS 0.00285f
C9436 VDD.n2970 VSS 0.00285f
C9437 VDD.n2971 VSS 8.62e-19
C9438 VDD.n2972 VSS 8.62e-19
C9439 VDD.n2973 VSS 0.00101f
C9440 VDD.n2974 VSS 0.00847f
C9441 VDD.t249 VSS 0.00541f
C9442 VDD.n2975 VSS 0.00424f
C9443 VDD.t671 VSS 0.00541f
C9444 VDD.n2976 VSS 0.00871f
C9445 VDD.t171 VSS 0.00541f
C9446 VDD.n2977 VSS 0.00565f
C9447 VDD.n2978 VSS 0.00101f
C9448 VDD.n2979 VSS 4.31e-19
C9449 VDD.n2980 VSS 8.62e-19
C9450 VDD.n2981 VSS 0.00285f
C9451 VDD.n2982 VSS 0.00214f
C9452 VDD.n2983 VSS 8.72e-19
C9453 VDD.n2984 VSS 0.0012f
C9454 VDD.n2985 VSS 0.00146f
C9455 VDD.n2986 VSS 0.00131f
C9456 VDD.n2987 VSS 0.0108f
C9457 VDD.n2988 VSS 0.0108f
C9458 VDD.n2989 VSS 0.0108f
C9459 VDD.n2990 VSS 0.00101f
C9460 VDD.n2991 VSS 0.00146f
C9461 VDD.n2992 VSS 0.00146f
C9462 VDD.n2993 VSS 0.00146f
C9463 VDD.n2994 VSS 0.00101f
C9464 VDD.n2995 VSS 0.0108f
C9465 VDD.n2996 VSS 0.0108f
C9466 VDD.n2997 VSS 0.00553f
C9467 VDD.n2998 VSS 0.0108f
C9468 VDD.n2999 VSS 0.00101f
C9469 VDD.n3000 VSS 0.00172f
C9470 VDD.n3001 VSS 0.00129f
C9471 VDD.n3002 VSS 0.00285f
C9472 VDD.n3003 VSS 0.00285f
C9473 VDD.n3004 VSS 0.00129f
C9474 VDD.n3005 VSS 0.00101f
C9475 VDD.n3006 VSS 0.00565f
C9476 VDD.t159 VSS 0.00459f
C9477 VDD.t269 VSS 0.00506f
C9478 VDD.n3007 VSS 0.00623f
C9479 VDD.n3008 VSS 0.00635f
C9480 VDD.n3009 VSS 0.0108f
C9481 VDD.n3010 VSS 0.00101f
C9482 VDD.n3011 VSS 0.00172f
C9483 VDD.n3012 VSS 0.00285f
C9484 VDD.n3013 VSS 0.00285f
C9485 VDD.n3014 VSS 0.00285f
C9486 VDD.n3015 VSS 0.00172f
C9487 VDD.n3016 VSS 0.00101f
C9488 VDD.n3017 VSS 0.00606f
C9489 VDD.t686 VSS 0.00541f
C9490 VDD.n3018 VSS 0.00641f
C9491 VDD.t299 VSS 0.00376f
C9492 VDD.n3019 VSS 0.00706f
C9493 VDD.n3020 VSS 0.0105f
C9494 VDD.n3021 VSS 0.0108f
C9495 VDD.n3022 VSS 0.00101f
C9496 VDD.n3023 VSS 0.00101f
C9497 VDD.n3024 VSS 0.00171f
C9498 VDD.n3025 VSS 0.00168f
C9499 VDD.n3026 VSS 0.00301f
C9500 VDD.n3027 VSS 0.00258f
C9501 VDD.n3028 VSS 5.25e-19
C9502 VDD.n3029 VSS 0.00235f
C9503 VDD.n3030 VSS 8.44e-19
C9504 VDD.n3031 VSS 0.00101f
C9505 VDD.n3032 VSS 8.23e-19
C9506 VDD.n3033 VSS 0.00559f
C9507 VDD.t169 VSS 0.00541f
C9508 VDD.t462 VSS 0.00541f
C9509 VDD.n3034 VSS 0.00606f
C9510 VDD.n3035 VSS 0.00101f
C9511 VDD.n3036 VSS 8.62e-19
C9512 VDD.n3037 VSS 8.62e-19
C9513 VDD.n3038 VSS 8.62e-19
C9514 VDD.n3039 VSS 0.00285f
C9515 VDD.n3040 VSS 0.00285f
C9516 VDD.n3041 VSS 0.00285f
C9517 VDD.n3042 VSS 8.62e-19
C9518 VDD.n3043 VSS 8.62e-19
C9519 VDD.n3044 VSS 0.00101f
C9520 VDD.n3045 VSS 0.00847f
C9521 VDD.t250 VSS 0.00541f
C9522 VDD.n3046 VSS 0.00424f
C9523 VDD.t431 VSS 0.00541f
C9524 VDD.n3047 VSS 0.00871f
C9525 VDD.t74 VSS 0.00541f
C9526 VDD.n3048 VSS 0.00565f
C9527 VDD.n3049 VSS 0.00101f
C9528 VDD.n3050 VSS 4.31e-19
C9529 VDD.n3051 VSS 8.62e-19
C9530 VDD.n3052 VSS 0.00285f
C9531 VDD.n3053 VSS 0.00214f
C9532 VDD.n3054 VSS 8.72e-19
C9533 VDD.n3055 VSS 0.0012f
C9534 VDD.n3056 VSS 0.00146f
C9535 VDD.n3057 VSS 0.00101f
C9536 VDD.n3058 VSS 0.0108f
C9537 VDD.n3059 VSS 0.0108f
C9538 VDD.n3060 VSS 0.0108f
C9539 VDD.n3061 VSS 0.00101f
C9540 VDD.n3062 VSS 0.00146f
C9541 VDD.n3063 VSS 0.00146f
C9542 VDD.n3064 VSS 0.00146f
C9543 VDD.n3065 VSS 0.00101f
C9544 VDD.n3066 VSS 0.0108f
C9545 VDD.n3067 VSS 0.0108f
C9546 VDD.n3068 VSS 0.00553f
C9547 VDD.n3069 VSS 0.0108f
C9548 VDD.n3070 VSS 0.00101f
C9549 VDD.n3071 VSS 0.00172f
C9550 VDD.n3072 VSS 0.00129f
C9551 VDD.n3073 VSS 0.00285f
C9552 VDD.n3074 VSS 0.00285f
C9553 VDD.n3075 VSS 0.00129f
C9554 VDD.n3076 VSS 0.00101f
C9555 VDD.n3077 VSS 0.00565f
C9556 VDD.t177 VSS 0.00459f
C9557 VDD.t460 VSS 0.00506f
C9558 VDD.n3078 VSS 0.00623f
C9559 VDD.n3079 VSS 0.00635f
C9560 VDD.n3080 VSS 0.0108f
C9561 VDD.n3081 VSS 0.00101f
C9562 VDD.n3082 VSS 0.00172f
C9563 VDD.n3083 VSS 0.00285f
C9564 VDD.n3084 VSS 0.00285f
C9565 VDD.n3085 VSS 0.00285f
C9566 VDD.n3086 VSS 0.00172f
C9567 VDD.n3087 VSS 0.00101f
C9568 VDD.n3088 VSS 0.00606f
C9569 VDD.t484 VSS 0.00541f
C9570 VDD.n3089 VSS 0.00641f
C9571 VDD.t43 VSS 0.00376f
C9572 VDD.n3090 VSS 0.0118f
C9573 VDD.n3091 VSS 0.00171f
C9574 VDD.n3092 VSS 0.00168f
C9575 VDD.n3093 VSS 0.00285f
C9576 VDD.t558 VSS 7.4e-19
C9577 VDD.t79 VSS 7.4e-19
C9578 VDD.n3094 VSS 0.00179f
C9579 VDD.n3095 VSS 0.00339f
C9580 VDD.n3096 VSS 0.00187f
C9581 VDD.n3097 VSS 0.00102f
C9582 VDD.n3098 VSS 0.00101f
C9583 VDD.n3099 VSS 0.00285f
C9584 VDD.t369 VSS 8.73e-19
C9585 VDD.t71 VSS 8.73e-19
C9586 VDD.n3100 VSS 0.00199f
C9587 VDD.n3101 VSS 0.0031f
C9588 VDD.n3102 VSS 0.00101f
C9589 VDD.t362 VSS 0.00535f
C9590 VDD.n3103 VSS 0.00101f
C9591 VDD.n3104 VSS 9.56e-19
C9592 VDD.t363 VSS 8.73e-19
C9593 VDD.t367 VSS 8.73e-19
C9594 VDD.n3105 VSS 0.00207f
C9595 VDD.n3106 VSS 0.00355f
C9596 VDD.n3107 VSS 9.18e-19
C9597 VDD.t365 VSS 0.00365f
C9598 VDD.n3108 VSS 0.0061f
C9599 VDD.n3109 VSS 0.00101f
C9600 VDD.t615 VSS 0.00535f
C9601 VDD.n3110 VSS 0.00101f
C9602 VDD.t610 VSS 8.73e-19
C9603 VDD.t616 VSS 8.73e-19
C9604 VDD.n3111 VSS 0.00198f
C9605 VDD.n3112 VSS 0.00239f
C9606 VDD.t614 VSS 0.00346f
C9607 VDD.n3113 VSS 0.00337f
C9608 VDD.n3114 VSS 0.00285f
C9609 VDD.t612 VSS 8.73e-19
C9610 VDD.t606 VSS 8.73e-19
C9611 VDD.n3115 VSS 0.00198f
C9612 VDD.n3116 VSS 0.00239f
C9613 VDD.n3117 VSS 0.00101f
C9614 VDD.t607 VSS 0.00535f
C9615 VDD.n3118 VSS 0.00101f
C9616 VDD.t417 VSS 8.73e-19
C9617 VDD.t608 VSS 8.73e-19
C9618 VDD.n3119 VSS 0.00198f
C9619 VDD.n3120 VSS 0.00239f
C9620 VDD.n3121 VSS 0.00111f
C9621 VDD.n3122 VSS 0.00285f
C9622 VDD.t411 VSS 8.73e-19
C9623 VDD.t397 VSS 8.73e-19
C9624 VDD.n3123 VSS 0.00198f
C9625 VDD.n3124 VSS 0.00239f
C9626 VDD.n3125 VSS 0.00101f
C9627 VDD.t386 VSS 0.00535f
C9628 VDD.n3126 VSS 0.00101f
C9629 VDD.t387 VSS 8.73e-19
C9630 VDD.t401 VSS 8.73e-19
C9631 VDD.n3127 VSS 0.00198f
C9632 VDD.n3128 VSS 0.00239f
C9633 VDD.n3129 VSS 0.00141f
C9634 VDD.n3130 VSS 0.00285f
C9635 VDD.t389 VSS 8.73e-19
C9636 VDD.t405 VSS 8.73e-19
C9637 VDD.n3131 VSS 0.00198f
C9638 VDD.n3132 VSS 0.00239f
C9639 VDD.n3133 VSS 0.00101f
C9640 VDD.t406 VSS 0.00535f
C9641 VDD.n3134 VSS 0.00101f
C9642 VDD.n3135 VSS 0.00144f
C9643 VDD.t407 VSS 8.73e-19
C9644 VDD.t391 VSS 8.73e-19
C9645 VDD.n3136 VSS 0.00198f
C9646 VDD.n3137 VSS 0.00239f
C9647 VDD.n3138 VSS 0.00285f
C9648 VDD.n3139 VSS 0.00129f
C9649 VDD.t409 VSS 8.73e-19
C9650 VDD.t395 VSS 8.73e-19
C9651 VDD.n3140 VSS 0.00198f
C9652 VDD.n3141 VSS 0.00239f
C9653 VDD.n3142 VSS 0.00101f
C9654 VDD.t402 VSS 0.00535f
C9655 VDD.n3143 VSS 0.00101f
C9656 VDD.n3144 VSS 0.00114f
C9657 VDD.t413 VSS 8.73e-19
C9658 VDD.t399 VSS 8.73e-19
C9659 VDD.n3145 VSS 0.00198f
C9660 VDD.n3146 VSS 0.00239f
C9661 VDD.n3147 VSS 0.00285f
C9662 VDD.n3148 VSS 9.93e-19
C9663 VDD.t415 VSS 8.73e-19
C9664 VDD.t403 VSS 8.73e-19
C9665 VDD.n3149 VSS 0.00198f
C9666 VDD.n3150 VSS 0.00239f
C9667 VDD.n3151 VSS 0.00101f
C9668 VDD.t393 VSS 0.00324f
C9669 VDD.n3152 VSS 0.00275f
C9670 VDD.n3153 VSS 0.00285f
C9671 VDD.t95 VSS 7.4e-19
C9672 VDD.t46 VSS 7.4e-19
C9673 VDD.n3154 VSS 0.00179f
C9674 VDD.n3155 VSS 0.00339f
C9675 VDD.n3156 VSS 0.00187f
C9676 VDD.n3157 VSS 0.00102f
C9677 VDD.n3158 VSS 0.00101f
C9678 VDD.n3159 VSS 0.00285f
C9679 VDD.t750 VSS 8.73e-19
C9680 VDD.t1 VSS 8.73e-19
C9681 VDD.n3160 VSS 0.00199f
C9682 VDD.n3161 VSS 0.0031f
C9683 VDD.n3162 VSS 0.00101f
C9684 VDD.t747 VSS 0.00535f
C9685 VDD.n3163 VSS 0.00101f
C9686 VDD.n3164 VSS 9.56e-19
C9687 VDD.t748 VSS 8.73e-19
C9688 VDD.t746 VSS 8.73e-19
C9689 VDD.n3165 VSS 0.00207f
C9690 VDD.n3166 VSS 0.00355f
C9691 VDD.n3167 VSS 9.18e-19
C9692 VDD.t744 VSS 0.00365f
C9693 VDD.n3168 VSS 0.0061f
C9694 VDD.n3169 VSS 0.00101f
C9695 VDD.t696 VSS 0.00535f
C9696 VDD.n3170 VSS 0.00101f
C9697 VDD.t693 VSS 8.73e-19
C9698 VDD.t697 VSS 8.73e-19
C9699 VDD.n3171 VSS 0.00198f
C9700 VDD.n3172 VSS 0.00239f
C9701 VDD.t691 VSS 0.00346f
C9702 VDD.n3173 VSS 0.00337f
C9703 VDD.n3174 VSS 0.00285f
C9704 VDD.t695 VSS 8.73e-19
C9705 VDD.t699 VSS 8.73e-19
C9706 VDD.n3175 VSS 0.00198f
C9707 VDD.n3176 VSS 0.00239f
C9708 VDD.n3177 VSS 0.00101f
C9709 VDD.t700 VSS 0.00535f
C9710 VDD.n3178 VSS 0.00101f
C9711 VDD.t225 VSS 8.73e-19
C9712 VDD.t701 VSS 8.73e-19
C9713 VDD.n3179 VSS 0.00198f
C9714 VDD.n3180 VSS 0.00239f
C9715 VDD.n3181 VSS 0.00111f
C9716 VDD.n3182 VSS 0.00285f
C9717 VDD.t229 VSS 8.73e-19
C9718 VDD.t241 VSS 8.73e-19
C9719 VDD.n3183 VSS 0.00198f
C9720 VDD.n3184 VSS 0.00239f
C9721 VDD.n3185 VSS 0.00101f
C9722 VDD.t216 VSS 0.00535f
C9723 VDD.n3186 VSS 0.00101f
C9724 VDD.t217 VSS 8.73e-19
C9725 VDD.t239 VSS 8.73e-19
C9726 VDD.n3187 VSS 0.00198f
C9727 VDD.n3188 VSS 0.00239f
C9728 VDD.n3189 VSS 0.00141f
C9729 VDD.n3190 VSS 0.00285f
C9730 VDD.t219 VSS 8.73e-19
C9731 VDD.t245 VSS 8.73e-19
C9732 VDD.n3191 VSS 0.00198f
C9733 VDD.n3192 VSS 0.00239f
C9734 VDD.n3193 VSS 0.00101f
C9735 VDD.t222 VSS 0.00535f
C9736 VDD.n3194 VSS 0.00101f
C9737 VDD.n3195 VSS 0.00144f
C9738 VDD.t223 VSS 8.73e-19
C9739 VDD.t235 VSS 8.73e-19
C9740 VDD.n3196 VSS 0.00198f
C9741 VDD.n3197 VSS 0.00239f
C9742 VDD.n3198 VSS 0.00285f
C9743 VDD.n3199 VSS 0.00129f
C9744 VDD.t227 VSS 8.73e-19
C9745 VDD.t237 VSS 8.73e-19
C9746 VDD.n3200 VSS 0.00198f
C9747 VDD.n3201 VSS 0.00239f
C9748 VDD.n3202 VSS 0.00101f
C9749 VDD.t246 VSS 0.00535f
C9750 VDD.n3203 VSS 0.00101f
C9751 VDD.n3204 VSS 0.00114f
C9752 VDD.t231 VSS 8.73e-19
C9753 VDD.t243 VSS 8.73e-19
C9754 VDD.n3205 VSS 0.00198f
C9755 VDD.n3206 VSS 0.00239f
C9756 VDD.n3207 VSS 0.293f
C9757 VDD.n3208 VSS 9.93e-19
C9758 VDD.t221 VSS 8.73e-19
C9759 VDD.t247 VSS 8.73e-19
C9760 VDD.n3209 VSS 0.00198f
C9761 VDD.n3210 VSS 0.00239f
C9762 VDD.n3211 VSS 0.00101f
C9763 VDD.t233 VSS 0.00324f
C9764 VDD.n3212 VSS 0.00275f
C9765 VDD.n3213 VSS 0.0275f
C9766 VDD.n3214 VSS 0.00803f
C9767 VDD.t232 VSS 0.0057f
C9768 VDD.n3215 VSS 0.00489f
C9769 VDD.t220 VSS 0.00535f
C9770 VDD.n3216 VSS 0.00489f
C9771 VDD.n3217 VSS 0.00101f
C9772 VDD.n3218 VSS 0.00144f
C9773 VDD.n3219 VSS 0.00285f
C9774 VDD.n3220 VSS 0.00285f
C9775 VDD.n3221 VSS 0.00285f
C9776 VDD.n3222 VSS 0.00129f
C9777 VDD.n3223 VSS 0.00101f
C9778 VDD.n3224 VSS 0.00489f
C9779 VDD.t230 VSS 0.00512f
C9780 VDD.t242 VSS 0.00512f
C9781 VDD.n3225 VSS 0.00489f
C9782 VDD.t226 VSS 0.00535f
C9783 VDD.n3226 VSS 0.00489f
C9784 VDD.t236 VSS 0.00535f
C9785 VDD.n3227 VSS 0.00489f
C9786 VDD.n3228 VSS 0.00101f
C9787 VDD.n3229 VSS 0.00114f
C9788 VDD.n3230 VSS 0.00285f
C9789 VDD.n3231 VSS 0.00285f
C9790 VDD.n3232 VSS 0.00157f
C9791 VDD.n3233 VSS 0.00285f
C9792 VDD.n3234 VSS 0.00285f
C9793 VDD.n3235 VSS 9.93e-19
C9794 VDD.n3236 VSS 0.00101f
C9795 VDD.n3237 VSS 0.00489f
C9796 VDD.t234 VSS 0.00535f
C9797 VDD.n3238 VSS 0.00489f
C9798 VDD.t218 VSS 0.00535f
C9799 VDD.n3239 VSS 0.00489f
C9800 VDD.t244 VSS 0.00535f
C9801 VDD.n3240 VSS 0.00489f
C9802 VDD.n3241 VSS 0.00101f
C9803 VDD.n3242 VSS 8.81e-19
C9804 VDD.n3243 VSS 0.00156f
C9805 VDD.n3244 VSS 0.00285f
C9806 VDD.n3245 VSS 0.00285f
C9807 VDD.n3246 VSS 0.00285f
C9808 VDD.n3247 VSS 0.00103f
C9809 VDD.n3248 VSS 0.00101f
C9810 VDD.n3249 VSS 0.00489f
C9811 VDD.t238 VSS 0.00535f
C9812 VDD.n3250 VSS 0.00489f
C9813 VDD.t228 VSS 0.00535f
C9814 VDD.t224 VSS 0.00977f
C9815 VDD.t240 VSS 0.00535f
C9816 VDD.n3251 VSS 0.00489f
C9817 VDD.n3252 VSS 0.00101f
C9818 VDD.n3253 VSS 0.00118f
C9819 VDD.n3254 VSS 0.00126f
C9820 VDD.n3255 VSS 0.00285f
C9821 VDD.n3256 VSS 0.00285f
C9822 VDD.n3257 VSS 0.00285f
C9823 VDD.n3258 VSS 0.00133f
C9824 VDD.n3259 VSS 0.00101f
C9825 VDD.n3260 VSS 0.00489f
C9826 VDD.t694 VSS 0.00535f
C9827 VDD.n3261 VSS 0.00489f
C9828 VDD.t698 VSS 0.00535f
C9829 VDD.n3262 VSS 0.00489f
C9830 VDD.t692 VSS 0.00535f
C9831 VDD.n3263 VSS 0.00489f
C9832 VDD.n3264 VSS 0.00101f
C9833 VDD.n3265 VSS 0.00148f
C9834 VDD.n3266 VSS 9.56e-19
C9835 VDD.n3267 VSS 0.00285f
C9836 VDD.n3268 VSS 0.00168f
C9837 VDD.n3269 VSS 0.00285f
C9838 VDD.n3270 VSS 0.00157f
C9839 VDD.n3271 VSS 0.00101f
C9840 VDD.n3272 VSS 0.00489f
C9841 VDD.t690 VSS 0.00535f
C9842 VDD.n3273 VSS 0.00372f
C9843 VDD.n3274 VSS 0.00489f
C9844 VDD.t743 VSS 0.00535f
C9845 VDD.n3275 VSS 0.00884f
C9846 VDD.n3276 VSS 0.00101f
C9847 VDD.n3277 VSS 8.72e-19
C9848 VDD.n3278 VSS 0.00214f
C9849 VDD.n3279 VSS 0.00285f
C9850 VDD.n3280 VSS 0.00285f
C9851 VDD.n3281 VSS 0.00285f
C9852 VDD.n3282 VSS 0.0012f
C9853 VDD.n3283 VSS 0.00187f
C9854 VDD.n3284 VSS 0.00102f
C9855 VDD.n3285 VSS 0.00489f
C9856 VDD.t745 VSS 0.00535f
C9857 VDD.n3286 VSS 0.00489f
C9858 VDD.t749 VSS 0.00535f
C9859 VDD.n3287 VSS 0.00372f
C9860 VDD.t0 VSS 0.00535f
C9861 VDD.n3288 VSS 0.00489f
C9862 VDD.n3289 VSS 0.00101f
C9863 VDD.n3290 VSS 9.09e-19
C9864 VDD.n3291 VSS 0.00101f
C9865 VDD.n3292 VSS 0.00214f
C9866 VDD.n3293 VSS 0.00214f
C9867 VDD.n3294 VSS 0.00127f
C9868 VDD.n3295 VSS 0.00101f
C9869 VDD.n3296 VSS 0.00721f
C9870 VDD.t94 VSS 0.00535f
C9871 VDD.n3297 VSS 0.00512f
C9872 VDD.t45 VSS 0.00535f
C9873 VDD.n3298 VSS 0.00378f
C9874 VDD.n3299 VSS 0.00101f
C9875 VDD.n3300 VSS 7.12e-19
C9876 VDD.n3301 VSS 0.00214f
C9877 VDD.n3302 VSS 0.0259f
C9878 VDD.n3303 VSS 0.0163f
C9879 VDD.n3304 VSS 0.00803f
C9880 VDD.t392 VSS 0.0057f
C9881 VDD.n3305 VSS 0.00489f
C9882 VDD.t414 VSS 0.00535f
C9883 VDD.n3306 VSS 0.00489f
C9884 VDD.n3307 VSS 0.00101f
C9885 VDD.n3308 VSS 0.00144f
C9886 VDD.n3309 VSS 0.00285f
C9887 VDD.n3310 VSS 0.00285f
C9888 VDD.n3311 VSS 0.00285f
C9889 VDD.n3312 VSS 0.00129f
C9890 VDD.n3313 VSS 0.00101f
C9891 VDD.n3314 VSS 0.00489f
C9892 VDD.t412 VSS 0.00512f
C9893 VDD.t398 VSS 0.00512f
C9894 VDD.n3315 VSS 0.00489f
C9895 VDD.t408 VSS 0.00535f
C9896 VDD.n3316 VSS 0.00489f
C9897 VDD.t394 VSS 0.00535f
C9898 VDD.n3317 VSS 0.00489f
C9899 VDD.n3318 VSS 0.00101f
C9900 VDD.n3319 VSS 0.00114f
C9901 VDD.n3320 VSS 0.00285f
C9902 VDD.n3321 VSS 0.00285f
C9903 VDD.n3322 VSS 0.00157f
C9904 VDD.n3323 VSS 0.00285f
C9905 VDD.n3324 VSS 0.00285f
C9906 VDD.n3325 VSS 9.93e-19
C9907 VDD.n3326 VSS 0.00101f
C9908 VDD.n3327 VSS 0.00489f
C9909 VDD.t390 VSS 0.00535f
C9910 VDD.n3328 VSS 0.00489f
C9911 VDD.t388 VSS 0.00535f
C9912 VDD.n3329 VSS 0.00489f
C9913 VDD.t404 VSS 0.00535f
C9914 VDD.n3330 VSS 0.00489f
C9915 VDD.n3331 VSS 0.00101f
C9916 VDD.n3332 VSS 8.81e-19
C9917 VDD.n3333 VSS 0.00156f
C9918 VDD.n3334 VSS 0.00285f
C9919 VDD.n3335 VSS 0.00285f
C9920 VDD.n3336 VSS 0.00285f
C9921 VDD.n3337 VSS 0.00103f
C9922 VDD.n3338 VSS 0.00101f
C9923 VDD.n3339 VSS 0.00489f
C9924 VDD.t400 VSS 0.00535f
C9925 VDD.n3340 VSS 0.00489f
C9926 VDD.t410 VSS 0.00535f
C9927 VDD.t416 VSS 0.00977f
C9928 VDD.t396 VSS 0.00535f
C9929 VDD.n3341 VSS 0.00489f
C9930 VDD.n3342 VSS 0.00101f
C9931 VDD.n3343 VSS 0.00118f
C9932 VDD.n3344 VSS 0.00126f
C9933 VDD.n3345 VSS 0.00285f
C9934 VDD.n3346 VSS 0.00285f
C9935 VDD.n3347 VSS 0.00285f
C9936 VDD.n3348 VSS 0.00133f
C9937 VDD.n3349 VSS 0.00101f
C9938 VDD.n3350 VSS 0.00489f
C9939 VDD.t611 VSS 0.00535f
C9940 VDD.n3351 VSS 0.00489f
C9941 VDD.t605 VSS 0.00535f
C9942 VDD.n3352 VSS 0.00489f
C9943 VDD.t609 VSS 0.00535f
C9944 VDD.n3353 VSS 0.00489f
C9945 VDD.n3354 VSS 0.00101f
C9946 VDD.n3355 VSS 0.00148f
C9947 VDD.n3356 VSS 9.56e-19
C9948 VDD.n3357 VSS 0.00285f
C9949 VDD.n3358 VSS 0.00168f
C9950 VDD.n3359 VSS 0.00285f
C9951 VDD.n3360 VSS 0.00157f
C9952 VDD.n3361 VSS 0.00101f
C9953 VDD.n3362 VSS 0.00489f
C9954 VDD.t613 VSS 0.00535f
C9955 VDD.n3363 VSS 0.00372f
C9956 VDD.n3364 VSS 0.00489f
C9957 VDD.t364 VSS 0.00535f
C9958 VDD.n3365 VSS 0.00884f
C9959 VDD.n3366 VSS 0.00101f
C9960 VDD.n3367 VSS 8.72e-19
C9961 VDD.n3368 VSS 0.00214f
C9962 VDD.n3369 VSS 0.00285f
C9963 VDD.n3370 VSS 0.00285f
C9964 VDD.n3371 VSS 0.00285f
C9965 VDD.n3372 VSS 0.0012f
C9966 VDD.n3373 VSS 0.00187f
C9967 VDD.n3374 VSS 0.00102f
C9968 VDD.n3375 VSS 0.00489f
C9969 VDD.t366 VSS 0.00535f
C9970 VDD.n3376 VSS 0.00489f
C9971 VDD.t368 VSS 0.00535f
C9972 VDD.n3377 VSS 0.00372f
C9973 VDD.t70 VSS 0.00535f
C9974 VDD.n3378 VSS 0.00489f
C9975 VDD.n3379 VSS 0.00101f
C9976 VDD.n3380 VSS 9.09e-19
C9977 VDD.n3381 VSS 0.00101f
C9978 VDD.n3382 VSS 0.00214f
C9979 VDD.n3383 VSS 0.00214f
C9980 VDD.n3384 VSS 0.00127f
C9981 VDD.n3385 VSS 0.00101f
C9982 VDD.n3386 VSS 0.00721f
C9983 VDD.t557 VSS 0.00535f
C9984 VDD.n3387 VSS 0.00512f
C9985 VDD.t78 VSS 0.00535f
C9986 VDD.n3388 VSS 0.00378f
C9987 VDD.n3389 VSS 0.00101f
C9988 VDD.n3390 VSS 7.12e-19
C9989 VDD.n3391 VSS 0.00214f
C9990 VDD.n3392 VSS 0.182f
C9991 VDD.n3393 VSS 0.0931f
C9992 VDD.n3394 VSS 0.0797f
.ends

