magic
tech sky130A
magscale 1 2
timestamp 1699323028
<< error_p >>
rect 916 1676 974 1682
rect 916 1642 928 1676
rect 916 1636 974 1642
<< nwell >>
rect 836 1776 1054 1856
rect 370 1687 1054 1776
rect 370 748 1040 1687
rect 370 500 1042 748
<< pmos >>
rect 930 1723 960 1807
<< pdiff >>
rect 872 1795 930 1807
rect 872 1735 884 1795
rect 918 1735 930 1795
rect 872 1723 930 1735
rect 960 1723 1018 1807
<< pdiffc >>
rect 884 1735 918 1795
<< nsubdiff >>
rect 440 600 978 614
rect 440 566 488 600
rect 522 566 568 600
rect 602 566 648 600
rect 682 566 728 600
rect 762 566 808 600
rect 842 566 888 600
rect 922 566 978 600
rect 440 546 978 566
<< nsubdiffcont >>
rect 488 566 522 600
rect 568 566 602 600
rect 648 566 682 600
rect 728 566 762 600
rect 808 566 842 600
rect 888 566 922 600
<< poly >>
rect 930 1807 960 1835
rect 930 1692 960 1723
rect 912 1676 978 1692
rect 912 1642 928 1676
rect 962 1642 978 1676
rect 912 1626 978 1642
<< polycont >>
rect 928 1642 962 1676
<< locali >>
rect 884 1795 918 1811
rect 884 1719 918 1735
rect 912 1642 928 1676
rect 962 1642 978 1676
rect 372 600 1042 614
rect 372 566 488 600
rect 524 566 568 600
rect 604 566 648 600
rect 684 566 728 600
rect 764 566 808 600
rect 844 566 888 600
rect 924 566 1042 600
rect 372 548 1042 566
<< viali >>
rect 884 1735 918 1795
rect 928 1642 962 1676
rect 490 566 522 600
rect 522 566 524 600
rect 570 566 602 600
rect 602 566 604 600
rect 650 566 682 600
rect 682 566 684 600
rect 730 566 762 600
rect 762 566 764 600
rect 810 566 842 600
rect 842 566 844 600
rect 890 566 922 600
rect 922 566 924 600
<< metal1 >>
rect 878 1796 924 1807
rect 855 1732 862 1796
rect 926 1732 934 1796
rect 855 1731 934 1732
rect 878 1723 924 1731
rect 916 1676 974 1682
rect 916 1642 928 1676
rect 962 1642 974 1676
rect 916 1636 974 1642
rect 372 606 1042 614
rect 372 554 480 606
rect 532 554 560 606
rect 612 554 640 606
rect 692 554 720 606
rect 772 554 800 606
rect 852 554 880 606
rect 932 554 1042 606
rect 372 548 1042 554
<< via1 >>
rect 862 1795 926 1796
rect 862 1735 884 1795
rect 884 1735 918 1795
rect 918 1735 926 1795
rect 862 1732 926 1735
rect 480 600 532 606
rect 480 566 490 600
rect 490 566 524 600
rect 524 566 532 600
rect 480 554 532 566
rect 560 600 612 606
rect 560 566 570 600
rect 570 566 604 600
rect 604 566 612 600
rect 560 554 612 566
rect 640 600 692 606
rect 640 566 650 600
rect 650 566 684 600
rect 684 566 692 600
rect 640 554 692 566
rect 720 600 772 606
rect 720 566 730 600
rect 730 566 764 600
rect 764 566 772 600
rect 720 554 772 566
rect 800 600 852 606
rect 800 566 810 600
rect 810 566 844 600
rect 844 566 852 600
rect 800 554 852 566
rect 880 600 932 606
rect 880 566 890 600
rect 890 566 924 600
rect 924 566 932 600
rect 880 554 932 566
<< metal2 >>
rect 852 1732 862 1796
rect 926 1732 935 1796
rect 855 1731 934 1732
rect 372 608 1042 614
rect 372 552 476 608
rect 532 552 556 608
rect 612 552 636 608
rect 692 552 716 608
rect 772 552 796 608
rect 852 552 876 608
rect 932 552 1042 608
rect 372 548 1042 552
<< via2 >>
rect 862 1732 926 1796
rect 476 606 532 608
rect 476 554 480 606
rect 480 554 532 606
rect 476 552 532 554
rect 556 606 612 608
rect 556 554 560 606
rect 560 554 612 606
rect 556 552 612 554
rect 636 606 692 608
rect 636 554 640 606
rect 640 554 692 606
rect 636 552 692 554
rect 716 606 772 608
rect 716 554 720 606
rect 720 554 772 606
rect 716 552 772 554
rect 796 606 852 608
rect 796 554 800 606
rect 800 554 852 606
rect 796 552 852 554
rect 876 606 932 608
rect 876 554 880 606
rect 880 554 932 606
rect 876 552 932 554
<< metal3 >>
rect 852 1796 935 1801
rect 852 1775 862 1796
rect 369 1773 862 1775
rect 926 1775 935 1796
rect 926 1773 1041 1775
rect 369 1709 473 1773
rect 537 1709 553 1773
rect 617 1709 633 1773
rect 697 1709 713 1773
rect 777 1709 793 1773
rect 857 1732 862 1773
rect 857 1709 873 1732
rect 937 1709 1041 1773
rect 369 1707 1041 1709
rect 369 1553 435 1707
rect 369 1489 370 1553
rect 434 1489 435 1553
rect 369 1473 435 1489
rect 369 1409 370 1473
rect 434 1409 435 1473
rect 369 1393 435 1409
rect 369 1329 370 1393
rect 434 1329 435 1393
rect 369 1313 435 1329
rect 369 1249 370 1313
rect 434 1249 435 1313
rect 369 1233 435 1249
rect 369 1169 370 1233
rect 434 1169 435 1233
rect 369 1153 435 1169
rect 369 1089 370 1153
rect 434 1089 435 1153
rect 369 1073 435 1089
rect 369 1009 370 1073
rect 434 1009 435 1073
rect 369 993 435 1009
rect 369 929 370 993
rect 434 929 435 993
rect 369 913 435 929
rect 369 849 370 913
rect 434 849 435 913
rect 369 833 435 849
rect 369 769 370 833
rect 434 769 435 833
rect 369 679 435 769
rect 495 675 555 1707
rect 615 615 675 1645
rect 735 675 795 1707
rect 855 615 915 1645
rect 975 1553 1041 1707
rect 975 1489 976 1553
rect 1040 1489 1041 1553
rect 975 1473 1041 1489
rect 975 1409 976 1473
rect 1040 1409 1041 1473
rect 975 1393 1041 1409
rect 975 1329 976 1393
rect 1040 1329 1041 1393
rect 975 1313 1041 1329
rect 975 1249 976 1313
rect 1040 1249 1041 1313
rect 975 1233 1041 1249
rect 975 1169 976 1233
rect 1040 1169 1041 1233
rect 975 1153 1041 1169
rect 975 1089 976 1153
rect 1040 1089 1041 1153
rect 975 1073 1041 1089
rect 975 1009 976 1073
rect 1040 1009 1041 1073
rect 975 993 1041 1009
rect 975 929 976 993
rect 1040 929 1041 993
rect 975 913 1041 929
rect 975 849 976 913
rect 1040 849 1041 913
rect 975 833 1041 849
rect 975 769 976 833
rect 1040 769 1041 833
rect 975 679 1041 769
rect 369 613 1041 615
rect 369 549 473 613
rect 537 549 553 613
rect 617 549 633 613
rect 697 549 713 613
rect 777 549 793 613
rect 857 549 873 613
rect 937 549 1041 613
rect 369 547 1041 549
<< via3 >>
rect 473 1709 537 1773
rect 553 1709 617 1773
rect 633 1709 697 1773
rect 713 1709 777 1773
rect 793 1709 857 1773
rect 873 1732 926 1773
rect 926 1732 937 1773
rect 873 1709 937 1732
rect 370 1489 434 1553
rect 370 1409 434 1473
rect 370 1329 434 1393
rect 370 1249 434 1313
rect 370 1169 434 1233
rect 370 1089 434 1153
rect 370 1009 434 1073
rect 370 929 434 993
rect 370 849 434 913
rect 370 769 434 833
rect 976 1489 1040 1553
rect 976 1409 1040 1473
rect 976 1329 1040 1393
rect 976 1249 1040 1313
rect 976 1169 1040 1233
rect 976 1089 1040 1153
rect 976 1009 1040 1073
rect 976 929 1040 993
rect 976 849 1040 913
rect 976 769 1040 833
rect 473 608 537 613
rect 473 552 476 608
rect 476 552 532 608
rect 532 552 537 608
rect 473 549 537 552
rect 553 608 617 613
rect 553 552 556 608
rect 556 552 612 608
rect 612 552 617 608
rect 553 549 617 552
rect 633 608 697 613
rect 633 552 636 608
rect 636 552 692 608
rect 692 552 697 608
rect 633 549 697 552
rect 713 608 777 613
rect 713 552 716 608
rect 716 552 772 608
rect 772 552 777 608
rect 713 549 777 552
rect 793 608 857 613
rect 793 552 796 608
rect 796 552 852 608
rect 852 552 857 608
rect 793 549 857 552
rect 873 608 937 613
rect 873 552 876 608
rect 876 552 932 608
rect 932 552 937 608
rect 873 549 937 552
<< metal4 >>
rect 369 1773 1041 1775
rect 369 1709 473 1773
rect 537 1709 553 1773
rect 617 1709 633 1773
rect 697 1709 713 1773
rect 777 1709 793 1773
rect 857 1709 873 1773
rect 937 1709 1041 1773
rect 369 1707 1041 1709
rect 369 1553 435 1707
rect 369 1489 370 1553
rect 434 1489 435 1553
rect 369 1473 435 1489
rect 369 1409 370 1473
rect 434 1409 435 1473
rect 369 1393 435 1409
rect 369 1329 370 1393
rect 434 1329 435 1393
rect 369 1313 435 1329
rect 369 1249 370 1313
rect 434 1249 435 1313
rect 369 1233 435 1249
rect 369 1169 370 1233
rect 434 1169 435 1233
rect 369 1153 435 1169
rect 369 1089 370 1153
rect 434 1089 435 1153
rect 369 1073 435 1089
rect 369 1009 370 1073
rect 434 1009 435 1073
rect 369 993 435 1009
rect 369 929 370 993
rect 434 929 435 993
rect 369 913 435 929
rect 369 849 370 913
rect 434 849 435 913
rect 369 833 435 849
rect 369 769 370 833
rect 434 769 435 833
rect 369 679 435 769
rect 495 615 555 1645
rect 615 675 675 1707
rect 735 615 795 1645
rect 855 675 915 1707
rect 975 1553 1041 1707
rect 975 1489 976 1553
rect 1040 1489 1041 1553
rect 975 1473 1041 1489
rect 975 1409 976 1473
rect 1040 1409 1041 1473
rect 975 1393 1041 1409
rect 975 1329 976 1393
rect 1040 1329 1041 1393
rect 975 1313 1041 1329
rect 975 1249 976 1313
rect 1040 1249 1041 1313
rect 975 1233 1041 1249
rect 975 1169 976 1233
rect 1040 1169 1041 1233
rect 975 1153 1041 1169
rect 975 1089 976 1153
rect 1040 1089 1041 1153
rect 975 1073 1041 1089
rect 975 1009 976 1073
rect 1040 1009 1041 1073
rect 975 993 1041 1009
rect 975 929 976 993
rect 1040 929 1041 993
rect 975 913 1041 929
rect 975 849 976 913
rect 1040 849 1041 913
rect 975 833 1041 849
rect 975 769 976 833
rect 1040 769 1041 833
rect 975 679 1041 769
rect 369 614 1041 615
rect 369 613 1042 614
rect 369 549 473 613
rect 537 549 553 613
rect 617 549 633 613
rect 697 549 713 613
rect 777 549 793 613
rect 857 549 873 613
rect 937 549 1042 613
rect 369 547 1042 549
rect 372 546 1042 547
<< labels >>
flabel metal1 928 1642 962 1676 0 FreeSans 320 0 0 0 SW
port 1 nsew
flabel nwell 372 546 1042 614 0 FreeSans 320 0 0 0 VDD
flabel pdiff 960 1723 1018 1807 0 FreeSans 320 0 0 0 delay_signal
port 2 nsew
flabel metal4 372 546 473 615 0 FreeSans 320 0 0 0 VDD
port 6 nsew
<< end >>
