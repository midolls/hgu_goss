magic
tech sky130A
magscale 1 2
timestamp 1699343576
<< nmoslvt >>
rect -35 -42 35 42
<< ndiff >>
rect -93 30 -35 42
rect -93 -30 -81 30
rect -47 -30 -35 30
rect -93 -42 -35 -30
rect 35 30 93 42
rect 35 -30 47 30
rect 81 -30 93 30
rect 35 -42 93 -30
<< ndiffc >>
rect -81 -30 -47 30
rect 47 -30 81 30
<< poly >>
rect -35 42 35 68
rect -35 -68 35 -42
<< locali >>
rect -81 30 -47 46
rect -81 -46 -47 -30
rect 47 30 81 46
rect 47 -46 81 -30
<< viali >>
rect -81 -30 -47 30
rect 47 -30 81 30
<< metal1 >>
rect -87 30 -41 42
rect -87 -30 -81 30
rect -47 -30 -41 30
rect -87 -42 -41 -30
rect 41 30 87 42
rect 41 -30 47 30
rect 81 -30 87 30
rect 41 -42 87 -30
<< properties >>
string FIXED_BBOX -178 -199 178 199
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 0.420 l 0.350 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
