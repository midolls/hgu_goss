magic
tech sky130A
magscale 1 2
timestamp 1699484509
<< error_p >>
rect -281 589 -263 757
rect -113 589 -79 769
rect -113 586 -95 589
rect -79 586 141 589
rect -113 550 141 586
rect -125 538 141 550
rect -129 522 -43 538
rect -33 522 -17 538
rect 17 522 33 538
rect 63 522 79 538
rect 113 522 129 538
rect -125 502 -43 522
rect -263 -407 62 -383
rect -263 -476 71 -407
rect -399 -637 71 -476
rect -399 -703 -263 -637
rect -231 -644 -224 -637
rect -219 -644 71 -637
rect -231 -645 71 -644
rect -219 -661 71 -645
rect -196 -680 107 -671
rect 204 -680 224 -671
rect -196 -703 224 -680
rect -231 -705 224 -703
rect -231 -707 23 -705
rect -232 -716 -219 -707
rect 240 -716 260 -707
rect -232 -741 260 -716
<< nwell >>
rect -263 589 263 769
rect -263 538 -113 589
rect -79 538 263 589
rect -263 -620 263 538
rect 62 -637 263 -620
rect -263 -644 263 -637
rect -263 -645 -231 -644
rect -224 -645 -219 -644
rect -263 -661 -219 -645
rect 71 -661 263 -644
rect -263 -703 263 -661
rect -263 -707 -231 -703
rect -224 -707 263 -703
rect -219 -716 240 -707
<< pmos >>
rect -63 -550 -33 550
rect 33 -550 63 550
<< pdiff >>
rect -125 -538 -113 550
rect -79 -538 -63 550
rect -125 -550 -63 -538
rect -33 538 33 550
rect -33 -538 -17 538
rect 17 -538 33 538
rect -33 -550 33 -538
rect 63 538 125 550
rect 63 -538 79 538
rect 113 -538 125 538
rect 63 -550 125 -538
<< pdiffc >>
rect -113 -538 -79 538
rect -17 -538 17 538
rect 79 -538 113 538
<< nsubdiff >>
rect -171 699 -121 733
rect -71 699 -25 733
rect 25 699 71 733
rect 121 699 224 733
rect 190 637 224 699
rect 190 -671 224 -595
rect -196 -705 -121 -671
rect -71 -705 -25 -671
rect 25 -705 71 -671
rect 121 -705 224 -671
<< nsubdiffcont >>
rect -121 699 -71 733
rect -25 699 25 733
rect 71 699 121 733
rect 190 -595 224 637
rect -121 -705 -71 -671
rect -25 -705 25 -671
rect 71 -705 121 -671
<< poly >>
rect -63 550 -33 576
rect 33 550 63 576
rect -63 -576 -33 -550
rect 33 -576 63 -550
<< locali >>
rect -171 699 -121 733
rect -71 699 -25 733
rect 25 699 71 733
rect 121 699 224 733
rect 190 637 224 699
rect -113 -554 -79 -538
rect -17 -554 17 -538
rect 79 -554 113 -538
rect 190 -671 224 -595
rect -196 -705 -121 -671
rect -71 -705 -25 -671
rect 25 -705 71 -671
rect 121 -705 224 -671
<< viali >>
rect -113 -538 -79 538
rect -17 -538 17 538
rect 79 -538 113 538
<< metal1 >>
rect -119 -538 -113 550
rect -79 -538 -73 550
rect -119 -550 -73 -538
rect -23 538 23 550
rect -23 -538 -17 538
rect 17 -538 23 538
rect -23 -550 23 -538
rect 73 538 119 550
rect 73 -538 79 538
rect 113 -538 119 538
rect 73 -550 119 -538
<< properties >>
string FIXED_BBOX -210 -716 210 716
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.5 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
