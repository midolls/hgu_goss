magic
tech sky130A
timestamp 1698470214
<< pwell >>
rect -1309 572 -1294 584
use hgu_cdac_unit  x1
timestamp 1698470058
transform -1 0 -791 0 -1 926
box 343 299 679 913
use hgu_cdac_unit  x2
timestamp 1698470058
transform 1 0 -1813 0 1 294
box 343 299 679 913
<< labels >>
flabel pwell -1309 572 -1294 584 0 FreeSans 80 0 0 0 SUB
port 1 nsew
<< end >>
