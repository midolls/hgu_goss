magic
tech sky130A
magscale 1 2
timestamp 1697885093
<< nwell >>
rect 2532 94 2608 112
<< psubdiff >>
rect 826 -336 1338 -324
rect 826 -370 868 -336
rect 902 -370 968 -336
rect 1002 -370 1068 -336
rect 1102 -370 1168 -336
rect 1202 -370 1268 -336
rect 1302 -370 1338 -336
rect 826 -382 1338 -370
rect 2028 -336 2540 -324
rect 2028 -370 2070 -336
rect 2104 -370 2170 -336
rect 2204 -370 2270 -336
rect 2304 -370 2370 -336
rect 2404 -370 2470 -336
rect 2504 -370 2540 -336
rect 2028 -382 2540 -370
rect 544 -816 2834 -792
rect 544 -850 568 -816
rect 602 -850 668 -816
rect 702 -850 768 -816
rect 802 -850 868 -816
rect 902 -850 968 -816
rect 1002 -850 1068 -816
rect 1102 -850 1168 -816
rect 1202 -850 1268 -816
rect 1302 -850 1368 -816
rect 1402 -850 1468 -816
rect 1502 -850 1568 -816
rect 1602 -850 1668 -816
rect 1702 -850 1768 -816
rect 1802 -850 1868 -816
rect 1902 -850 1968 -816
rect 2002 -850 2068 -816
rect 2102 -850 2168 -816
rect 2202 -850 2268 -816
rect 2302 -850 2368 -816
rect 2402 -850 2468 -816
rect 2502 -850 2568 -816
rect 2602 -850 2668 -816
rect 2702 -850 2768 -816
rect 2802 -850 2834 -816
rect 544 -976 2834 -850
rect 544 -1010 568 -976
rect 602 -1010 668 -976
rect 702 -980 2834 -976
rect 702 -1010 1568 -980
rect 544 -1014 1568 -1010
rect 1602 -1014 1668 -980
rect 1702 -1014 1768 -980
rect 1802 -1014 2834 -980
rect 544 -1034 2834 -1014
rect 764 -1038 2834 -1034
rect 764 -1062 1516 -1038
rect 764 -1096 770 -1062
rect 804 -1096 868 -1062
rect 902 -1096 968 -1062
rect 1002 -1096 1068 -1062
rect 1102 -1096 1168 -1062
rect 1202 -1096 1268 -1062
rect 1302 -1096 1368 -1062
rect 1402 -1096 1468 -1062
rect 1502 -1096 1516 -1062
rect 764 -1120 1516 -1096
rect 1860 -1062 2834 -1038
rect 1860 -1096 1868 -1062
rect 1902 -1096 1968 -1062
rect 2002 -1096 2068 -1062
rect 2102 -1096 2168 -1062
rect 2202 -1096 2268 -1062
rect 2302 -1096 2368 -1062
rect 2402 -1096 2468 -1062
rect 2502 -1096 2568 -1062
rect 2602 -1096 2668 -1062
rect 2702 -1096 2768 -1062
rect 2802 -1096 2834 -1062
rect 1860 -1120 2834 -1096
<< nsubdiff >>
rect 762 412 2624 428
rect 762 378 802 412
rect 836 378 958 412
rect 992 378 1114 412
rect 1148 378 1270 412
rect 1304 378 1426 412
rect 1460 378 1582 412
rect 1616 378 1738 412
rect 1772 378 1894 412
rect 1928 378 2050 412
rect 2084 378 2206 412
rect 2240 378 2362 412
rect 2396 378 2518 412
rect 2552 378 2624 412
rect 762 364 2624 378
rect 758 -1792 2440 -1776
rect 758 -1826 818 -1792
rect 852 -1826 958 -1792
rect 992 -1826 1114 -1792
rect 1148 -1826 1270 -1792
rect 1304 -1826 1426 -1792
rect 1460 -1826 1582 -1792
rect 1616 -1826 1738 -1792
rect 1772 -1826 1894 -1792
rect 1928 -1826 2050 -1792
rect 2084 -1826 2206 -1792
rect 2240 -1826 2362 -1792
rect 2396 -1826 2440 -1792
rect 758 -1840 2440 -1826
<< psubdiffcont >>
rect 868 -370 902 -336
rect 968 -370 1002 -336
rect 1068 -370 1102 -336
rect 1168 -370 1202 -336
rect 1268 -370 1302 -336
rect 2070 -370 2104 -336
rect 2170 -370 2204 -336
rect 2270 -370 2304 -336
rect 2370 -370 2404 -336
rect 2470 -370 2504 -336
rect 568 -850 602 -816
rect 668 -850 702 -816
rect 768 -850 802 -816
rect 868 -850 902 -816
rect 968 -850 1002 -816
rect 1068 -850 1102 -816
rect 1168 -850 1202 -816
rect 1268 -850 1302 -816
rect 1368 -850 1402 -816
rect 1468 -850 1502 -816
rect 1568 -850 1602 -816
rect 1668 -850 1702 -816
rect 1768 -850 1802 -816
rect 1868 -850 1902 -816
rect 1968 -850 2002 -816
rect 2068 -850 2102 -816
rect 2168 -850 2202 -816
rect 2268 -850 2302 -816
rect 2368 -850 2402 -816
rect 2468 -850 2502 -816
rect 2568 -850 2602 -816
rect 2668 -850 2702 -816
rect 2768 -850 2802 -816
rect 568 -1010 602 -976
rect 668 -1010 702 -976
rect 1568 -1014 1602 -980
rect 1668 -1014 1702 -980
rect 1768 -1014 1802 -980
rect 770 -1096 804 -1062
rect 868 -1096 902 -1062
rect 968 -1096 1002 -1062
rect 1068 -1096 1102 -1062
rect 1168 -1096 1202 -1062
rect 1268 -1096 1302 -1062
rect 1368 -1096 1402 -1062
rect 1468 -1096 1502 -1062
rect 1868 -1096 1902 -1062
rect 1968 -1096 2002 -1062
rect 2068 -1096 2102 -1062
rect 2168 -1096 2202 -1062
rect 2268 -1096 2302 -1062
rect 2368 -1096 2402 -1062
rect 2468 -1096 2502 -1062
rect 2568 -1096 2602 -1062
rect 2668 -1096 2702 -1062
rect 2768 -1096 2802 -1062
<< nsubdiffcont >>
rect 802 378 836 412
rect 958 378 992 412
rect 1114 378 1148 412
rect 1270 378 1304 412
rect 1426 378 1460 412
rect 1582 378 1616 412
rect 1738 378 1772 412
rect 1894 378 1928 412
rect 2050 378 2084 412
rect 2206 378 2240 412
rect 2362 378 2396 412
rect 2518 378 2552 412
rect 818 -1826 852 -1792
rect 958 -1826 992 -1792
rect 1114 -1826 1148 -1792
rect 1270 -1826 1304 -1792
rect 1426 -1826 1460 -1792
rect 1582 -1826 1616 -1792
rect 1738 -1826 1772 -1792
rect 1894 -1826 1928 -1792
rect 2050 -1826 2084 -1792
rect 2206 -1826 2240 -1792
rect 2362 -1826 2396 -1792
<< poly >>
rect 1040 24 1074 96
rect 1040 8 1106 24
rect 1040 -26 1056 8
rect 1090 -26 1106 8
rect 1040 -42 1106 -26
rect 1248 -22 1278 110
rect 1416 64 1566 94
rect 1248 -38 1328 -22
rect 1040 -132 1074 -42
rect 1248 -72 1278 -38
rect 1312 -72 1328 -38
rect 1248 -88 1328 -72
rect 1248 -152 1278 -88
rect 1416 -446 1446 64
rect 1624 22 1654 78
rect 1536 -8 1654 22
rect 1712 22 1742 78
rect 1800 64 1950 94
rect 1712 -8 1830 22
rect 1536 -26 1566 -8
rect 1488 -38 1566 -26
rect 1488 -72 1504 -38
rect 1538 -72 1566 -38
rect 1488 -84 1566 -72
rect 1536 -154 1566 -84
rect 1800 -94 1830 -8
rect 1800 -106 1878 -94
rect 1800 -140 1828 -106
rect 1862 -140 1878 -106
rect 1800 -152 1878 -140
rect 1800 -160 1830 -152
rect 1650 -398 1716 -384
rect 1650 -432 1666 -398
rect 1700 -432 1716 -398
rect 1650 -446 1716 -432
rect 1920 -446 1950 64
rect 2088 -86 2118 110
rect 2292 24 2322 96
rect 2256 8 2322 24
rect 2256 -26 2272 8
rect 2306 -26 2322 8
rect 2256 -42 2322 -26
rect 2036 -102 2118 -86
rect 2036 -136 2052 -102
rect 2086 -136 2118 -102
rect 2292 -132 2322 -42
rect 2036 -152 2118 -136
rect 1416 -476 1524 -446
rect 1842 -476 1950 -446
rect 534 -1522 564 -1292
rect 622 -1456 652 -1292
rect 768 -1306 852 -1290
rect 768 -1340 784 -1306
rect 818 -1340 852 -1306
rect 768 -1356 852 -1340
rect 622 -1472 704 -1456
rect 622 -1506 654 -1472
rect 688 -1506 704 -1472
rect 622 -1522 704 -1506
rect 822 -1522 852 -1356
rect 1216 -1394 1248 -1312
rect 1422 -1394 1452 -1292
rect 1592 -1300 1658 -1286
rect 1592 -1334 1608 -1300
rect 1642 -1334 1658 -1300
rect 1592 -1348 1658 -1334
rect 1716 -1300 1782 -1286
rect 1716 -1334 1732 -1300
rect 1766 -1334 1782 -1300
rect 1716 -1348 1782 -1334
rect 1216 -1408 1314 -1394
rect 1216 -1442 1264 -1408
rect 1298 -1442 1314 -1408
rect 1216 -1456 1314 -1442
rect 1422 -1408 1506 -1394
rect 1422 -1442 1456 -1408
rect 1490 -1442 1506 -1408
rect 1422 -1456 1506 -1442
rect 1716 -1404 1782 -1390
rect 1920 -1394 1950 -1292
rect 2124 -1394 2156 -1312
rect 1716 -1438 1732 -1404
rect 1766 -1438 1782 -1404
rect 1716 -1452 1782 -1438
rect 1872 -1408 1950 -1394
rect 1872 -1442 1888 -1408
rect 1922 -1442 1950 -1408
rect 1216 -1508 1248 -1456
rect 1422 -1522 1452 -1456
rect 1592 -1472 1658 -1458
rect 1592 -1506 1608 -1472
rect 1642 -1506 1658 -1472
rect 1592 -1520 1658 -1506
rect 1628 -1532 1658 -1520
rect 1716 -1522 1746 -1452
rect 1872 -1456 1950 -1442
rect 2060 -1408 2156 -1394
rect 2060 -1442 2076 -1408
rect 2110 -1442 2156 -1408
rect 2060 -1456 2156 -1442
rect 1920 -1522 1950 -1456
rect 2124 -1508 2156 -1456
rect 482 -1768 564 -1752
rect 482 -1802 498 -1768
rect 532 -1802 564 -1768
rect 482 -1818 564 -1802
<< polycont >>
rect 1056 -26 1090 8
rect 1278 -72 1312 -38
rect 1504 -72 1538 -38
rect 1828 -140 1862 -106
rect 1666 -432 1700 -398
rect 2272 -26 2306 8
rect 2052 -136 2086 -102
rect 784 -1340 818 -1306
rect 654 -1506 688 -1472
rect 1608 -1334 1642 -1300
rect 1732 -1334 1766 -1300
rect 1264 -1442 1298 -1408
rect 1456 -1442 1490 -1408
rect 1732 -1438 1766 -1404
rect 1888 -1442 1922 -1408
rect 1608 -1506 1642 -1472
rect 2076 -1442 2110 -1408
rect 498 -1802 532 -1768
<< locali >>
rect 762 412 2624 428
rect 762 378 802 412
rect 836 378 958 412
rect 992 378 1114 412
rect 1148 378 1270 412
rect 1304 378 1426 412
rect 1460 378 1582 412
rect 1616 378 1738 412
rect 1772 378 1894 412
rect 1928 378 2050 412
rect 2084 378 2206 412
rect 2240 378 2362 412
rect 2396 378 2518 412
rect 2552 378 2624 412
rect 762 364 2624 378
rect 898 298 932 364
rect 1090 300 1124 364
rect 1290 298 1324 364
rect 1490 296 1524 364
rect 1666 290 1700 364
rect 1842 308 1876 364
rect 2042 298 2076 364
rect 2242 298 2276 364
rect 2434 308 2468 364
rect 1040 -26 1056 8
rect 1090 -26 1106 8
rect 2256 -26 2272 8
rect 2306 -26 2322 8
rect 1262 -72 1278 -38
rect 1312 -72 1328 -38
rect 1488 -72 1504 -38
rect 1538 -72 1554 -38
rect 1812 -140 1828 -106
rect 1862 -140 1878 -106
rect 2036 -136 2052 -102
rect 2086 -136 2102 -102
rect 898 -324 932 -218
rect 1090 -324 1124 -228
rect 1290 -324 1324 -240
rect 2042 -324 2076 -176
rect 2242 -324 2276 -266
rect 2434 -324 2468 -262
rect 826 -336 1338 -324
rect 826 -370 868 -336
rect 902 -370 968 -336
rect 1002 -370 1068 -336
rect 1102 -370 1168 -336
rect 1202 -370 1268 -336
rect 1302 -370 1338 -336
rect 826 -382 1338 -370
rect 2028 -336 2540 -324
rect 2028 -370 2070 -336
rect 2104 -370 2170 -336
rect 2204 -370 2270 -336
rect 2304 -370 2370 -336
rect 2404 -370 2470 -336
rect 2504 -370 2540 -336
rect 2028 -382 2540 -370
rect 1650 -432 1666 -398
rect 1700 -432 1716 -398
rect 1570 -792 1604 -690
rect 1762 -792 1796 -690
rect 544 -816 2834 -792
rect 544 -850 568 -816
rect 602 -850 668 -816
rect 702 -850 768 -816
rect 802 -850 868 -816
rect 902 -850 968 -816
rect 1002 -850 1068 -816
rect 1102 -850 1168 -816
rect 1202 -850 1268 -816
rect 1302 -850 1368 -816
rect 1402 -850 1468 -816
rect 1502 -850 1568 -816
rect 1602 -850 1668 -816
rect 1702 -850 1768 -816
rect 1802 -850 1868 -816
rect 1902 -850 1968 -816
rect 2002 -850 2068 -816
rect 2102 -850 2168 -816
rect 2202 -850 2268 -816
rect 2302 -850 2368 -816
rect 2402 -850 2468 -816
rect 2502 -850 2568 -816
rect 2602 -850 2668 -816
rect 2702 -850 2768 -816
rect 2802 -850 2834 -816
rect 544 -976 2834 -850
rect 544 -1010 568 -976
rect 602 -1010 668 -976
rect 702 -980 2834 -976
rect 702 -1010 1568 -980
rect 544 -1014 1568 -1010
rect 1602 -1014 1668 -980
rect 1702 -1014 1768 -980
rect 1802 -1014 2834 -980
rect 544 -1034 2834 -1014
rect 664 -1112 698 -1034
rect 764 -1038 2834 -1034
rect 764 -1062 1516 -1038
rect 764 -1096 770 -1062
rect 804 -1096 868 -1062
rect 902 -1096 968 -1062
rect 1002 -1096 1068 -1062
rect 1102 -1096 1168 -1062
rect 1202 -1096 1268 -1062
rect 1302 -1096 1368 -1062
rect 1402 -1096 1468 -1062
rect 1502 -1096 1516 -1062
rect 1670 -1094 1704 -1038
rect 1860 -1062 2834 -1038
rect 764 -1120 1516 -1096
rect 1860 -1096 1868 -1062
rect 1902 -1096 1968 -1062
rect 2002 -1096 2068 -1062
rect 2102 -1096 2168 -1062
rect 2202 -1096 2268 -1062
rect 2302 -1096 2368 -1062
rect 2402 -1096 2468 -1062
rect 2502 -1096 2568 -1062
rect 2602 -1096 2668 -1062
rect 2702 -1096 2768 -1062
rect 2802 -1096 2834 -1062
rect 1860 -1120 2834 -1096
rect 776 -1196 810 -1120
rect 1072 -1176 1106 -1120
rect 1264 -1180 1298 -1120
rect 1464 -1182 1498 -1120
rect 1874 -1182 1908 -1120
rect 2074 -1180 2108 -1120
rect 2266 -1180 2300 -1120
rect 768 -1340 784 -1306
rect 818 -1340 834 -1306
rect 1592 -1334 1608 -1300
rect 1642 -1334 1658 -1300
rect 1716 -1334 1732 -1300
rect 1766 -1334 1782 -1300
rect 1248 -1442 1264 -1408
rect 1298 -1442 1314 -1408
rect 1440 -1442 1456 -1408
rect 1490 -1442 1506 -1408
rect 1716 -1438 1732 -1404
rect 1766 -1438 1782 -1404
rect 1872 -1442 1888 -1408
rect 1922 -1442 1938 -1408
rect 2060 -1442 2076 -1408
rect 2110 -1442 2126 -1408
rect 488 -1506 654 -1472
rect 688 -1506 704 -1472
rect 1592 -1506 1608 -1472
rect 1642 -1506 1658 -1472
rect 488 -1550 522 -1506
rect 482 -1802 498 -1768
rect 532 -1802 548 -1768
rect 776 -1776 810 -1716
rect 1072 -1776 1106 -1642
rect 1264 -1776 1298 -1642
rect 1464 -1776 1498 -1720
rect 1670 -1776 1704 -1660
rect 1874 -1776 1908 -1716
rect 2074 -1776 2108 -1720
rect 2266 -1776 2300 -1720
rect 758 -1792 2440 -1776
rect 758 -1826 818 -1792
rect 852 -1826 958 -1792
rect 992 -1826 1114 -1792
rect 1148 -1826 1270 -1792
rect 1304 -1826 1426 -1792
rect 1460 -1826 1582 -1792
rect 1616 -1826 1738 -1792
rect 1772 -1826 1894 -1792
rect 1928 -1826 2050 -1792
rect 2084 -1826 2206 -1792
rect 2240 -1826 2362 -1792
rect 2396 -1826 2440 -1792
rect 758 -1840 2440 -1826
<< viali >>
rect 802 378 836 412
rect 958 378 992 412
rect 1114 378 1148 412
rect 1270 378 1304 412
rect 1426 378 1460 412
rect 1582 378 1616 412
rect 1738 378 1772 412
rect 1894 378 1928 412
rect 2050 378 2084 412
rect 2206 378 2240 412
rect 2362 378 2396 412
rect 2518 378 2552 412
rect 1056 -26 1090 8
rect 2272 -26 2306 8
rect 1278 -72 1312 -38
rect 1504 -72 1538 -38
rect 1828 -140 1862 -106
rect 2052 -136 2086 -102
rect 868 -370 902 -336
rect 968 -370 1002 -336
rect 1068 -370 1102 -336
rect 1168 -370 1202 -336
rect 1268 -370 1302 -336
rect 2070 -370 2104 -336
rect 2170 -370 2204 -336
rect 2270 -370 2304 -336
rect 2370 -370 2404 -336
rect 2470 -370 2504 -336
rect 1666 -432 1700 -398
rect 568 -850 602 -816
rect 668 -850 702 -816
rect 768 -850 802 -816
rect 868 -850 902 -816
rect 968 -850 1002 -816
rect 1068 -850 1102 -816
rect 1168 -850 1202 -816
rect 1268 -850 1302 -816
rect 1368 -850 1402 -816
rect 1468 -850 1502 -816
rect 1568 -850 1602 -816
rect 1668 -850 1702 -816
rect 1768 -850 1802 -816
rect 1868 -850 1902 -816
rect 1968 -850 2002 -816
rect 2068 -850 2102 -816
rect 2168 -850 2202 -816
rect 2268 -850 2302 -816
rect 2368 -850 2402 -816
rect 2468 -850 2502 -816
rect 2568 -850 2602 -816
rect 2668 -850 2702 -816
rect 2768 -850 2802 -816
rect 568 -1010 602 -976
rect 668 -1010 702 -976
rect 1568 -1014 1602 -980
rect 1668 -1014 1702 -980
rect 1768 -1014 1802 -980
rect 770 -1096 804 -1062
rect 868 -1096 902 -1062
rect 968 -1096 1002 -1062
rect 1068 -1096 1102 -1062
rect 1168 -1096 1202 -1062
rect 1268 -1096 1302 -1062
rect 1368 -1096 1402 -1062
rect 1468 -1096 1502 -1062
rect 1868 -1096 1902 -1062
rect 1968 -1096 2002 -1062
rect 2068 -1096 2102 -1062
rect 2168 -1096 2202 -1062
rect 2268 -1096 2302 -1062
rect 2368 -1096 2402 -1062
rect 2468 -1096 2502 -1062
rect 2568 -1096 2602 -1062
rect 2668 -1096 2702 -1062
rect 2768 -1096 2802 -1062
rect 784 -1340 818 -1306
rect 1608 -1334 1642 -1300
rect 1732 -1334 1766 -1300
rect 1264 -1442 1298 -1408
rect 1456 -1442 1490 -1408
rect 1732 -1438 1766 -1404
rect 1888 -1442 1922 -1408
rect 2076 -1442 2110 -1408
rect 654 -1506 688 -1472
rect 1608 -1506 1642 -1472
rect 498 -1802 532 -1768
rect 818 -1826 852 -1792
rect 958 -1826 992 -1792
rect 1114 -1826 1148 -1792
rect 1270 -1826 1304 -1792
rect 1426 -1826 1460 -1792
rect 1582 -1826 1616 -1792
rect 1738 -1826 1772 -1792
rect 1894 -1826 1928 -1792
rect 2050 -1826 2084 -1792
rect 2206 -1826 2240 -1792
rect 2362 -1826 2396 -1792
<< metal1 >>
rect 762 422 2834 428
rect 762 412 2776 422
rect 762 378 802 412
rect 836 378 958 412
rect 992 378 1114 412
rect 1148 378 1270 412
rect 1304 378 1426 412
rect 1460 378 1582 412
rect 1616 378 1738 412
rect 1772 378 1894 412
rect 1928 378 2050 412
rect 2084 378 2206 412
rect 2240 378 2362 412
rect 2396 378 2518 412
rect 2552 378 2776 412
rect 762 370 2776 378
rect 2828 370 2834 422
rect 762 364 2834 370
rect 802 100 836 150
rect 994 100 1028 142
rect 802 66 1028 100
rect 802 -60 836 66
rect 1042 16 1106 22
rect 1042 -36 1048 16
rect 1100 8 1106 16
rect 1202 8 1236 152
rect 1100 -26 1236 8
rect 1100 -36 1106 -26
rect 1042 -42 1106 -36
rect 802 -72 878 -60
rect 802 -124 814 -72
rect 866 -102 878 -72
rect 866 -124 1028 -102
rect 802 -136 1028 -124
rect 802 -188 836 -136
rect 994 -178 1028 -136
rect 1202 -220 1236 -26
rect 1264 -28 1328 -22
rect 1264 -80 1270 -28
rect 1322 -80 1328 -28
rect 1264 -86 1328 -80
rect 1486 -28 1550 -22
rect 1486 -80 1492 -28
rect 1544 -80 1550 -28
rect 1486 -86 1550 -80
rect 1578 -86 1612 112
rect 1754 -18 1788 110
rect 1724 -24 1788 -18
rect 1724 -76 1730 -24
rect 1782 -76 1788 -24
rect 1724 -82 1788 -76
rect 1578 -92 1642 -86
rect 1578 -144 1584 -92
rect 1636 -144 1642 -92
rect 1578 -150 1642 -144
rect 1578 -184 1612 -150
rect 1754 -180 1788 -82
rect 2130 8 2164 142
rect 2338 100 2372 142
rect 2530 112 2564 142
rect 2530 100 2608 112
rect 2338 66 2544 100
rect 2530 48 2544 66
rect 2596 48 2608 100
rect 2530 36 2608 48
rect 2256 16 2320 22
rect 2256 8 2262 16
rect 2130 -26 2262 8
rect 1816 -92 1880 -86
rect 1816 -144 1822 -92
rect 1874 -144 1880 -92
rect 1816 -150 1880 -144
rect 2036 -92 2100 -86
rect 2036 -144 2042 -92
rect 2094 -144 2100 -92
rect 2036 -150 2100 -144
rect 2130 -178 2164 -26
rect 2256 -36 2262 -26
rect 2314 -36 2320 16
rect 2256 -42 2320 -36
rect 2530 -102 2564 36
rect 2338 -136 2564 -102
rect 2338 -178 2372 -136
rect 2530 -178 2564 -136
rect 826 -336 1338 -324
rect 826 -370 868 -336
rect 902 -370 968 -336
rect 1002 -370 1068 -336
rect 1102 -370 1168 -336
rect 1202 -370 1268 -336
rect 1302 -370 1338 -336
rect 2028 -336 2540 -324
rect 548 -470 640 -380
rect 826 -382 1338 -370
rect 1490 -440 1524 -376
rect 690 -474 1524 -440
rect 1650 -388 1714 -382
rect 1650 -440 1656 -388
rect 1708 -440 1714 -388
rect 1650 -446 1714 -440
rect 1842 -440 1876 -366
rect 2028 -370 2070 -336
rect 2104 -370 2170 -336
rect 2204 -370 2270 -336
rect 2304 -370 2370 -336
rect 2404 -370 2470 -336
rect 2504 -370 2540 -336
rect 2028 -382 2540 -370
rect 1842 -474 2676 -440
rect 2726 -468 2818 -378
rect 690 -502 724 -474
rect 882 -502 916 -474
rect 1074 -502 1108 -474
rect 1266 -648 1300 -474
rect 2066 -514 2100 -474
rect 2258 -514 2292 -474
rect 2450 -516 2484 -474
rect 2642 -514 2676 -474
rect 594 -730 628 -690
rect 786 -730 820 -690
rect 978 -730 1012 -690
rect 1170 -730 1204 -690
rect 1362 -730 1396 -690
rect 1474 -730 1508 -694
rect 1666 -730 1700 -690
rect 1970 -730 2004 -690
rect 2162 -730 2196 -690
rect 2354 -730 2388 -690
rect 2546 -730 2580 -690
rect 2738 -730 2772 -690
rect 594 -764 2772 -730
rect 544 -816 2834 -792
rect 544 -850 568 -816
rect 602 -850 668 -816
rect 702 -850 768 -816
rect 802 -850 868 -816
rect 902 -850 968 -816
rect 1002 -850 1068 -816
rect 1102 -850 1168 -816
rect 1202 -850 1268 -816
rect 1302 -850 1368 -816
rect 1402 -850 1468 -816
rect 1502 -850 1568 -816
rect 1602 -850 1668 -816
rect 1702 -850 1768 -816
rect 1802 -850 1868 -816
rect 1902 -850 1968 -816
rect 2002 -850 2068 -816
rect 2102 -850 2168 -816
rect 2202 -850 2268 -816
rect 2302 -850 2368 -816
rect 2402 -850 2468 -816
rect 2502 -850 2568 -816
rect 2602 -850 2668 -816
rect 2702 -850 2768 -816
rect 2802 -850 2834 -816
rect 544 -976 2834 -850
rect 544 -1010 568 -976
rect 602 -1010 668 -976
rect 702 -980 2834 -976
rect 702 -1010 1568 -980
rect 544 -1014 1568 -1010
rect 1602 -1014 1668 -980
rect 1702 -1014 1768 -980
rect 1802 -1014 2834 -980
rect 544 -1034 2834 -1014
rect 764 -1038 2834 -1034
rect 764 -1062 1516 -1038
rect 764 -1096 770 -1062
rect 804 -1096 868 -1062
rect 902 -1096 968 -1062
rect 1002 -1096 1068 -1062
rect 1102 -1096 1168 -1062
rect 1202 -1096 1268 -1062
rect 1302 -1096 1368 -1062
rect 1402 -1096 1468 -1062
rect 1502 -1096 1516 -1062
rect 764 -1120 1516 -1096
rect 1860 -1062 2834 -1038
rect 1860 -1096 1868 -1062
rect 1902 -1096 1968 -1062
rect 2002 -1096 2068 -1062
rect 2102 -1096 2168 -1062
rect 2202 -1096 2268 -1062
rect 2302 -1096 2368 -1062
rect 2402 -1096 2468 -1062
rect 2502 -1096 2568 -1062
rect 2602 -1096 2668 -1062
rect 2702 -1096 2768 -1062
rect 2802 -1096 2834 -1062
rect 1860 -1120 2834 -1096
rect 970 -1186 1016 -1174
rect 970 -1254 976 -1186
rect 1010 -1254 1016 -1186
rect 488 -1306 522 -1256
rect 768 -1306 830 -1300
rect 488 -1340 784 -1306
rect 818 -1340 830 -1306
rect 576 -1600 610 -1340
rect 768 -1346 830 -1340
rect 864 -1438 898 -1258
rect 970 -1266 1016 -1254
rect 1162 -1186 1208 -1174
rect 1162 -1254 1168 -1186
rect 1202 -1254 1208 -1186
rect 1576 -1232 1582 -1226
rect 1752 -1232 1758 -1226
rect 1792 -1232 1798 -1226
rect 1162 -1266 1208 -1254
rect 976 -1294 1010 -1266
rect 1168 -1294 1202 -1266
rect 976 -1328 1202 -1294
rect 864 -1444 928 -1438
rect 640 -1458 704 -1456
rect 638 -1462 704 -1458
rect 638 -1512 646 -1462
rect 640 -1514 646 -1512
rect 698 -1514 704 -1462
rect 640 -1520 704 -1514
rect 864 -1496 870 -1444
rect 922 -1496 928 -1444
rect 864 -1502 928 -1496
rect 976 -1490 1010 -1328
rect 1252 -1408 1310 -1402
rect 1382 -1408 1416 -1254
rect 1532 -1260 1616 -1232
rect 1752 -1260 1840 -1232
rect 1252 -1442 1264 -1408
rect 1298 -1442 1416 -1408
rect 1252 -1448 1310 -1442
rect 864 -1556 898 -1502
rect 976 -1524 1202 -1490
rect 976 -1553 1010 -1524
rect 1168 -1553 1202 -1524
rect 970 -1609 1016 -1553
rect 970 -1709 976 -1609
rect 1010 -1709 1016 -1609
rect 482 -1758 546 -1752
rect 482 -1810 488 -1758
rect 540 -1768 546 -1758
rect 664 -1768 698 -1720
rect 970 -1721 1016 -1709
rect 1162 -1565 1208 -1553
rect 1162 -1709 1168 -1565
rect 1202 -1709 1208 -1565
rect 1382 -1597 1416 -1442
rect 1444 -1408 1502 -1402
rect 1532 -1404 1566 -1260
rect 1594 -1294 1658 -1288
rect 1594 -1346 1600 -1294
rect 1652 -1346 1658 -1294
rect 1594 -1352 1658 -1346
rect 1714 -1294 1778 -1288
rect 1714 -1346 1720 -1294
rect 1772 -1346 1778 -1294
rect 1714 -1352 1778 -1346
rect 1720 -1404 1778 -1398
rect 1532 -1408 1732 -1404
rect 1444 -1442 1456 -1408
rect 1490 -1438 1732 -1408
rect 1766 -1438 1778 -1404
rect 1490 -1442 1566 -1438
rect 1444 -1448 1502 -1442
rect 1532 -1552 1566 -1442
rect 1720 -1444 1778 -1438
rect 1806 -1408 1840 -1260
rect 1876 -1408 1934 -1402
rect 1806 -1442 1888 -1408
rect 1922 -1442 1934 -1408
rect 1596 -1472 1654 -1466
rect 1806 -1472 1840 -1442
rect 1876 -1448 1934 -1442
rect 1962 -1408 1996 -1254
rect 2170 -1294 2204 -1266
rect 2362 -1294 2396 -1254
rect 2170 -1328 2396 -1294
rect 2064 -1408 2122 -1402
rect 1962 -1442 2076 -1408
rect 2110 -1442 2122 -1408
rect 1596 -1506 1608 -1472
rect 1642 -1506 1840 -1472
rect 1596 -1512 1654 -1506
rect 1806 -1552 1840 -1506
rect 1532 -1586 1616 -1552
rect 1752 -1586 1840 -1552
rect 1962 -1597 1996 -1442
rect 2064 -1448 2122 -1442
rect 2362 -1490 2396 -1328
rect 2170 -1524 2396 -1490
rect 2170 -1558 2204 -1524
rect 2362 -1609 2396 -1524
rect 1162 -1721 1208 -1709
rect 540 -1802 698 -1768
rect 758 -1782 2828 -1776
rect 758 -1792 2770 -1782
rect 540 -1810 546 -1802
rect 482 -1816 546 -1810
rect 758 -1826 818 -1792
rect 852 -1826 958 -1792
rect 992 -1826 1114 -1792
rect 1148 -1826 1270 -1792
rect 1304 -1826 1426 -1792
rect 1460 -1826 1582 -1792
rect 1616 -1826 1738 -1792
rect 1772 -1826 1894 -1792
rect 1928 -1826 2050 -1792
rect 2084 -1826 2206 -1792
rect 2240 -1826 2362 -1792
rect 2396 -1826 2770 -1792
rect 758 -1834 2770 -1826
rect 2822 -1834 2828 -1782
rect 758 -1840 2828 -1834
<< via1 >>
rect 2776 370 2828 422
rect 1048 8 1100 16
rect 1048 -26 1056 8
rect 1056 -26 1090 8
rect 1090 -26 1100 8
rect 1048 -36 1100 -26
rect 814 -124 866 -72
rect 1270 -38 1322 -28
rect 1270 -72 1278 -38
rect 1278 -72 1312 -38
rect 1312 -72 1322 -38
rect 1270 -80 1322 -72
rect 1492 -38 1544 -28
rect 1492 -72 1504 -38
rect 1504 -72 1538 -38
rect 1538 -72 1544 -38
rect 1492 -80 1544 -72
rect 1730 -76 1782 -24
rect 1584 -144 1636 -92
rect 2544 48 2596 100
rect 2262 8 2314 16
rect 2262 -26 2272 8
rect 2272 -26 2306 8
rect 2306 -26 2314 8
rect 1822 -106 1874 -92
rect 1822 -140 1828 -106
rect 1828 -140 1862 -106
rect 1862 -140 1874 -106
rect 1822 -144 1874 -140
rect 2042 -102 2094 -92
rect 2042 -136 2052 -102
rect 2052 -136 2086 -102
rect 2086 -136 2094 -102
rect 2042 -144 2094 -136
rect 2262 -36 2314 -26
rect 1656 -398 1708 -388
rect 1656 -432 1666 -398
rect 1666 -432 1700 -398
rect 1700 -432 1708 -398
rect 1656 -440 1708 -432
rect 646 -1472 698 -1462
rect 646 -1506 654 -1472
rect 654 -1506 688 -1472
rect 688 -1506 698 -1472
rect 646 -1514 698 -1506
rect 870 -1496 922 -1444
rect 488 -1768 540 -1758
rect 1600 -1300 1652 -1294
rect 1600 -1334 1608 -1300
rect 1608 -1334 1642 -1300
rect 1642 -1334 1652 -1300
rect 1600 -1346 1652 -1334
rect 1720 -1300 1772 -1294
rect 1720 -1334 1732 -1300
rect 1732 -1334 1766 -1300
rect 1766 -1334 1772 -1300
rect 1720 -1346 1772 -1334
rect 488 -1802 498 -1768
rect 498 -1802 532 -1768
rect 532 -1802 540 -1768
rect 488 -1810 540 -1802
rect 2770 -1834 2822 -1782
<< metal2 >>
rect 2770 422 2834 428
rect 2770 370 2776 422
rect 2828 370 2834 422
rect 2770 364 2834 370
rect 488 102 564 112
rect 488 46 498 102
rect 554 46 564 102
rect 488 36 564 46
rect 488 -1752 516 36
rect 670 -60 698 112
rect 2532 102 2608 112
rect 2532 46 2542 102
rect 2598 46 2608 102
rect 2532 36 2608 46
rect 1042 16 1106 22
rect 1042 -36 1048 16
rect 1100 -36 1106 16
rect 2256 16 2320 22
rect 1042 -42 1106 -36
rect 1264 -24 1550 -22
rect 1724 -24 1788 -18
rect 1264 -28 1730 -24
rect 658 -70 734 -60
rect 658 -126 668 -70
rect 724 -126 734 -70
rect 658 -136 734 -126
rect 802 -70 878 -60
rect 802 -126 812 -70
rect 868 -126 878 -70
rect 802 -136 878 -126
rect 670 -1456 698 -136
rect 1062 -982 1090 -42
rect 1264 -80 1270 -28
rect 1322 -56 1492 -28
rect 1322 -80 1328 -56
rect 1264 -86 1328 -80
rect 1486 -80 1492 -56
rect 1544 -58 1730 -28
rect 1544 -80 1550 -58
rect 1486 -86 1550 -80
rect 1724 -76 1730 -58
rect 1782 -76 1788 -24
rect 2256 -36 2262 16
rect 2314 -36 2320 16
rect 2256 -42 2320 -36
rect 1724 -82 1788 -76
rect 1578 -92 1642 -86
rect 1578 -144 1584 -92
rect 1636 -116 1642 -92
rect 1816 -92 1880 -86
rect 1816 -116 1822 -92
rect 1636 -144 1822 -116
rect 1874 -116 1880 -92
rect 2036 -92 2100 -86
rect 2036 -116 2042 -92
rect 1874 -144 2042 -116
rect 2094 -144 2100 -92
rect 1578 -150 2100 -144
rect 1650 -388 1714 -382
rect 1650 -440 1656 -388
rect 1708 -440 1714 -388
rect 1650 -446 1714 -440
rect 2272 -982 2300 -42
rect 1062 -1010 1618 -982
rect 1590 -1288 1618 -1010
rect 1744 -1012 2300 -982
rect 1744 -1288 1772 -1012
rect 1590 -1294 1658 -1288
rect 1590 -1346 1600 -1294
rect 1652 -1346 1658 -1294
rect 1590 -1352 1658 -1346
rect 1714 -1294 1784 -1288
rect 1714 -1346 1720 -1294
rect 1772 -1346 1784 -1294
rect 1714 -1352 1784 -1346
rect 864 -1444 928 -1438
rect 640 -1462 704 -1456
rect 640 -1514 646 -1462
rect 698 -1514 704 -1462
rect 864 -1496 870 -1444
rect 922 -1496 928 -1444
rect 864 -1502 928 -1496
rect 640 -1520 704 -1514
rect 482 -1758 546 -1752
rect 482 -1810 488 -1758
rect 540 -1810 546 -1758
rect 482 -1816 546 -1810
rect 670 -1816 698 -1520
rect 2800 -1776 2828 364
rect 2764 -1782 2828 -1776
rect 2764 -1834 2770 -1782
rect 2822 -1834 2828 -1782
rect 2764 -1840 2828 -1834
<< via2 >>
rect 498 46 554 102
rect 2542 100 2598 102
rect 2542 48 2544 100
rect 2544 48 2596 100
rect 2596 48 2598 100
rect 2542 46 2598 48
rect 668 -126 724 -70
rect 812 -72 868 -70
rect 812 -124 814 -72
rect 814 -124 866 -72
rect 866 -124 868 -72
rect 812 -126 868 -124
<< metal3 >>
rect 488 104 564 112
rect 2532 104 2608 112
rect 488 102 2608 104
rect 488 46 498 102
rect 554 46 2542 102
rect 2598 46 2608 102
rect 488 44 2608 46
rect 488 36 564 44
rect 2532 36 2608 44
rect 658 -66 734 -60
rect 802 -66 878 -60
rect 488 -70 2608 -66
rect 488 -126 668 -70
rect 724 -126 812 -70
rect 868 -126 2608 -70
rect 658 -136 734 -126
rect 802 -136 878 -126
use sky130_fd_pr__nfet_01v8_HNLS5R  XM1
timestamp 1697527592
transform 1 0 1683 0 1 -602
box -221 -126 221 156
use sky130_fd_pr__nfet_01v8_lvt_Y5HS5Z  XM2
timestamp 1697708322
transform 1 0 995 0 1 -602
box -417 -126 413 188
use sky130_fd_pr__nfet_01v8_lvt_Y5HS5Z  XM3
timestamp 1697708322
transform -1 0 2371 0 1 -602
box -417 -126 413 188
use sky130_fd_pr__nfet_01v8_648S5X  XM4
timestamp 1697700693
transform 1 0 1551 0 1 -278
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_648S5X  XM5
timestamp 1697700693
transform 1 0 1815 0 1 -278
box -73 -126 73 126
use sky130_fd_pr__pfet_01v8_XGS3BL  XM6
timestamp 1697700693
transform 1 0 1639 0 1 209
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM7
timestamp 1697700693
transform 1 0 1727 0 1 209
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM8
timestamp 1697700693
transform 1 0 1551 0 1 209
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM9
timestamp 1697700693
transform 1 0 1463 0 1 209
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM10
timestamp 1697700693
transform 1 0 1815 0 1 209
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM11
timestamp 1697700693
transform 1 0 1903 0 1 209
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_MQX2PY  XM12
timestamp 1697710383
transform 1 0 2103 0 1 225
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_L7T3GD  XM13
timestamp 1697710383
transform 1 0 2103 0 1 -220
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_MQP8BZ  XM14
timestamp 1697710383
transform 1 0 2403 0 1 225
box -311 -303 311 303
use sky130_fd_pr__nfet_01v8_PK34ES  XM15
timestamp 1697705701
transform 1 0 2403 0 1 -224
box -173 -72 173 92
use sky130_fd_pr__pfet_01v8_MQX2PY  XM16
timestamp 1697710383
transform -1 0 1731 0 -1 -1637
box -211 -303 211 303
use sky130_fd_pr__pfet_01v8_MQX2PY  XM17
timestamp 1697710383
transform -1 0 1643 0 -1 -1637
box -211 -303 211 303
use sky130_fd_pr__pfet_01v8_MQX2PY  XM18
timestamp 1697710383
transform 1 0 1263 0 1 225
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_9NW3WL  XM19
timestamp 1697452276
transform -1 0 1643 0 -1 -1176
box -73 -110 73 110
use sky130_fd_pr__nfet_01v8_L7T3GD  XM20
timestamp 1697710383
transform -1 0 1263 0 1 -220
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_MQP8BZ  XM21
timestamp 1697710383
transform -1 0 963 0 1 225
box -311 -303 311 303
use sky130_fd_pr__nfet_01v8_PK34ES  XM22
timestamp 1697705701
transform 1 0 963 0 1 -224
box -173 -72 173 92
use sky130_fd_pr__nfet_01v8_9NW3WL  XM23
timestamp 1697452276
transform -1 0 1731 0 -1 -1176
box -73 -110 73 110
use sky130_fd_pr__pfet_01v8_MQX2PY  XM24
timestamp 1697710383
transform 1 0 637 0 -1 -1637
box -211 -303 211 303
use sky130_fd_pr__pfet_01v8_MQX2PY  XM25
timestamp 1697710383
transform 1 0 549 0 -1 -1637
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_9NW3WL  XM26
timestamp 1697452276
transform 1 0 637 0 -1 -1182
box -73 -110 73 110
use sky130_fd_pr__nfet_01v8_9NW3WL  XM27
timestamp 1697452276
transform 1 0 549 0 -1 -1182
box -73 -110 73 110
use sky130_fd_pr__pfet_01v8_MQX2PY  XM28
timestamp 1697710383
transform 1 0 837 0 -1 -1637
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_L7T3GD  XM29
timestamp 1697710383
transform 1 0 837 0 -1 -1224
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_MQX2PY  XM30
timestamp 1697710383
transform -1 0 1437 0 -1 -1637
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_L7T3GD  XM31
timestamp 1697710383
transform -1 0 1437 0 -1 -1224
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_MQP8BZ  XM32
timestamp 1697710383
transform -1 0 1137 0 -1 -1637
box -311 -303 311 303
use sky130_fd_pr__nfet_01v8_PK34ES  XM33
timestamp 1697705701
transform -1 0 1137 0 -1 -1220
box -173 -72 173 92
use sky130_fd_pr__pfet_01v8_MQX2PY  XM34
timestamp 1697710383
transform 1 0 1935 0 -1 -1637
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_L7T3GD  XM35
timestamp 1697710383
transform 1 0 1935 0 -1 -1224
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_MQP8BZ  XM36
timestamp 1697710383
transform 1 0 2235 0 -1 -1637
box -311 -303 311 303
use sky130_fd_pr__nfet_01v8_PK34ES  XM37
timestamp 1697705701
transform 1 0 2235 0 -1 -1220
box -173 -72 173 92
<< labels >>
flabel space 1578 -92 1612 121 0 FreeSans 288 0 0 0 X
flabel space 1754 -24 1788 121 0 FreeSans 288 0 0 0 Y
flabel space 2130 -190 2164 153 0 FreeSans 288 0 0 0 X_inv
flabel space 2530 -190 2564 48 0 FreeSans 288 0 0 0 X_drive
flabel metal1 2726 -468 2818 -378 0 FreeSans 288 0 0 0 cdac_vn
port 1 nsew
flabel metal1 548 -470 640 -380 0 FreeSans 288 0 0 0 cdac_vp
port 2 nsew
flabel space 1202 -220 1236 153 0 FreeSans 240 0 0 0 Y_inv
flabel space 802 -72 836 153 0 FreeSans 240 0 0 0 Y_drive
flabel space 864 -1444 898 -1254 0 FreeSans 240 0 0 0 ready
port 3 nsew
flabel metal1 2362 -1609 2396 -1254 0 FreeSans 240 0 0 0 comp_outp
port 5 nsew
flabel metal1 976 -1609 1010 -1254 0 FreeSans 240 0 0 0 comp_outn
port 6 nsew
flabel metal1 1806 -1586 1840 -1232 0 FreeSans 240 0 0 0 RS_p
flabel metal1 1532 -1586 1566 -1232 0 FreeSans 240 0 0 0 RS_n
flabel via1 1656 -440 1708 -388 0 FreeSans 240 0 0 0 clk
port 7 nsew
flabel metal1 836 364 958 428 0 FreeSans 240 0 0 0 VDD
port 8 nsew
flabel metal1 702 -980 2834 -850 0 FreeSans 240 0 0 0 VSS
port 9 nsew
<< end >>
