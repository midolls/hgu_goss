* NGSPICE file created from hgu_cdac_unit.ext - technology: sky130A

.subckt hgu_cdac_unit CBOT CTOP SUB
C0 CTOP CBOT 5.11f
.ends

