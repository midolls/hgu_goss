magic
tech sky130A
magscale 1 2
timestamp 1706708240
<< nwell >>
rect 116 1595 1020 1994
rect 392 606 1020 977
<< pwell >>
rect 155 1355 425 1537
rect 472 1355 658 1537
rect 748 1355 934 1537
rect 368 1317 402 1355
rect 472 1351 493 1355
rect 748 1351 769 1355
rect 459 1317 493 1351
rect 735 1317 769 1351
rect 643 1221 677 1255
rect 919 1221 953 1255
rect 643 1217 664 1221
rect 919 1217 940 1221
rect 478 1035 664 1217
rect 754 1035 940 1217
<< scnmos >>
rect 233 1381 263 1511
rect 317 1381 347 1511
rect 550 1381 580 1511
rect 826 1381 856 1511
rect 556 1061 586 1191
rect 832 1061 862 1191
<< scpmoshvt >>
rect 233 1631 263 1831
rect 317 1631 347 1831
rect 550 1631 580 1831
rect 826 1631 856 1831
rect 556 741 586 941
rect 832 741 862 941
<< ndiff >>
rect 181 1495 233 1511
rect 181 1461 189 1495
rect 223 1461 233 1495
rect 181 1427 233 1461
rect 181 1393 189 1427
rect 223 1393 233 1427
rect 181 1381 233 1393
rect 263 1381 317 1511
rect 347 1495 399 1511
rect 347 1461 357 1495
rect 391 1461 399 1495
rect 347 1427 399 1461
rect 347 1393 357 1427
rect 391 1393 399 1427
rect 347 1381 399 1393
rect 498 1499 550 1511
rect 498 1465 506 1499
rect 540 1465 550 1499
rect 498 1431 550 1465
rect 498 1397 506 1431
rect 540 1397 550 1431
rect 498 1381 550 1397
rect 580 1499 632 1511
rect 580 1465 590 1499
rect 624 1465 632 1499
rect 580 1431 632 1465
rect 580 1397 590 1431
rect 624 1397 632 1431
rect 580 1381 632 1397
rect 774 1499 826 1511
rect 774 1465 782 1499
rect 816 1465 826 1499
rect 774 1431 826 1465
rect 774 1397 782 1431
rect 816 1397 826 1431
rect 774 1381 826 1397
rect 856 1499 908 1511
rect 856 1465 866 1499
rect 900 1465 908 1499
rect 856 1431 908 1465
rect 856 1397 866 1431
rect 900 1397 908 1431
rect 856 1381 908 1397
rect 504 1175 556 1191
rect 504 1141 512 1175
rect 546 1141 556 1175
rect 504 1107 556 1141
rect 504 1073 512 1107
rect 546 1073 556 1107
rect 504 1061 556 1073
rect 586 1175 638 1191
rect 586 1141 596 1175
rect 630 1141 638 1175
rect 586 1107 638 1141
rect 586 1073 596 1107
rect 630 1073 638 1107
rect 586 1061 638 1073
rect 780 1175 832 1191
rect 780 1141 788 1175
rect 822 1141 832 1175
rect 780 1107 832 1141
rect 780 1073 788 1107
rect 822 1073 832 1107
rect 780 1061 832 1073
rect 862 1175 914 1191
rect 862 1141 872 1175
rect 906 1141 914 1175
rect 862 1107 914 1141
rect 862 1073 872 1107
rect 906 1073 914 1107
rect 862 1061 914 1073
<< pdiff >>
rect 181 1819 233 1831
rect 181 1785 189 1819
rect 223 1785 233 1819
rect 181 1751 233 1785
rect 181 1717 189 1751
rect 223 1717 233 1751
rect 181 1683 233 1717
rect 181 1649 189 1683
rect 223 1649 233 1683
rect 181 1631 233 1649
rect 263 1819 317 1831
rect 263 1785 273 1819
rect 307 1785 317 1819
rect 263 1751 317 1785
rect 263 1717 273 1751
rect 307 1717 317 1751
rect 263 1683 317 1717
rect 263 1649 273 1683
rect 307 1649 317 1683
rect 263 1631 317 1649
rect 347 1819 399 1831
rect 347 1785 357 1819
rect 391 1785 399 1819
rect 347 1751 399 1785
rect 347 1717 357 1751
rect 391 1717 399 1751
rect 347 1683 399 1717
rect 347 1649 357 1683
rect 391 1649 399 1683
rect 347 1631 399 1649
rect 498 1819 550 1831
rect 498 1785 506 1819
rect 540 1785 550 1819
rect 498 1751 550 1785
rect 498 1717 506 1751
rect 540 1717 550 1751
rect 498 1683 550 1717
rect 498 1649 506 1683
rect 540 1649 550 1683
rect 498 1631 550 1649
rect 580 1819 632 1831
rect 580 1785 590 1819
rect 624 1785 632 1819
rect 580 1751 632 1785
rect 580 1717 590 1751
rect 624 1717 632 1751
rect 580 1683 632 1717
rect 580 1649 590 1683
rect 624 1649 632 1683
rect 580 1631 632 1649
rect 774 1819 826 1831
rect 774 1785 782 1819
rect 816 1785 826 1819
rect 774 1751 826 1785
rect 774 1717 782 1751
rect 816 1717 826 1751
rect 774 1683 826 1717
rect 774 1649 782 1683
rect 816 1649 826 1683
rect 774 1631 826 1649
rect 856 1819 908 1831
rect 856 1785 866 1819
rect 900 1785 908 1819
rect 856 1751 908 1785
rect 856 1717 866 1751
rect 900 1717 908 1751
rect 856 1683 908 1717
rect 856 1649 866 1683
rect 900 1649 908 1683
rect 856 1631 908 1649
rect 504 923 556 941
rect 504 889 512 923
rect 546 889 556 923
rect 504 855 556 889
rect 504 821 512 855
rect 546 821 556 855
rect 504 787 556 821
rect 504 753 512 787
rect 546 753 556 787
rect 504 741 556 753
rect 586 923 638 941
rect 586 889 596 923
rect 630 889 638 923
rect 586 855 638 889
rect 586 821 596 855
rect 630 821 638 855
rect 586 787 638 821
rect 586 753 596 787
rect 630 753 638 787
rect 586 741 638 753
rect 780 923 832 941
rect 780 889 788 923
rect 822 889 832 923
rect 780 855 832 889
rect 780 821 788 855
rect 822 821 832 855
rect 780 787 832 821
rect 780 753 788 787
rect 822 753 832 787
rect 780 741 832 753
rect 862 923 914 941
rect 862 889 872 923
rect 906 889 914 923
rect 862 855 914 889
rect 862 821 872 855
rect 906 821 914 855
rect 862 787 914 821
rect 862 753 872 787
rect 906 753 914 787
rect 862 741 914 753
<< ndiffc >>
rect 189 1461 223 1495
rect 189 1393 223 1427
rect 357 1461 391 1495
rect 357 1393 391 1427
rect 506 1465 540 1499
rect 506 1397 540 1431
rect 590 1465 624 1499
rect 590 1397 624 1431
rect 782 1465 816 1499
rect 782 1397 816 1431
rect 866 1465 900 1499
rect 866 1397 900 1431
rect 512 1141 546 1175
rect 512 1073 546 1107
rect 596 1141 630 1175
rect 596 1073 630 1107
rect 788 1141 822 1175
rect 788 1073 822 1107
rect 872 1141 906 1175
rect 872 1073 906 1107
<< pdiffc >>
rect 189 1785 223 1819
rect 189 1717 223 1751
rect 189 1649 223 1683
rect 273 1785 307 1819
rect 273 1717 307 1751
rect 273 1649 307 1683
rect 357 1785 391 1819
rect 357 1717 391 1751
rect 357 1649 391 1683
rect 506 1785 540 1819
rect 506 1717 540 1751
rect 506 1649 540 1683
rect 590 1785 624 1819
rect 590 1717 624 1751
rect 590 1649 624 1683
rect 782 1785 816 1819
rect 782 1717 816 1751
rect 782 1649 816 1683
rect 866 1785 900 1819
rect 866 1717 900 1751
rect 866 1649 900 1683
rect 512 889 546 923
rect 512 821 546 855
rect 512 753 546 787
rect 596 889 630 923
rect 596 821 630 855
rect 596 753 630 787
rect 788 889 822 923
rect 788 821 822 855
rect 788 753 822 787
rect 872 889 906 923
rect 872 821 906 855
rect 872 753 906 787
<< psubdiff >>
rect 154 1310 982 1326
rect 154 1308 644 1310
rect 154 1306 554 1308
rect 154 1304 274 1306
rect 154 1270 186 1304
rect 220 1272 274 1304
rect 308 1302 458 1306
rect 308 1272 368 1302
rect 220 1270 368 1272
rect 154 1268 368 1270
rect 402 1272 458 1302
rect 492 1274 554 1306
rect 588 1276 644 1308
rect 678 1308 982 1310
rect 678 1276 740 1308
rect 588 1274 740 1276
rect 774 1306 982 1308
rect 774 1274 832 1306
rect 492 1272 832 1274
rect 866 1304 982 1306
rect 866 1272 920 1304
rect 402 1270 920 1272
rect 954 1270 982 1304
rect 402 1268 982 1270
rect 154 1246 982 1268
<< nsubdiff >>
rect 154 1940 982 1950
rect 154 1938 556 1940
rect 154 1904 184 1938
rect 218 1936 462 1938
rect 218 1904 276 1936
rect 154 1902 276 1904
rect 310 1902 366 1936
rect 400 1904 462 1936
rect 496 1906 556 1938
rect 590 1938 826 1940
rect 590 1906 646 1938
rect 496 1904 646 1906
rect 680 1904 736 1938
rect 770 1906 826 1938
rect 860 1938 982 1940
rect 860 1906 918 1938
rect 770 1904 918 1906
rect 952 1904 982 1938
rect 400 1902 982 1904
rect 154 1896 982 1902
rect 430 646 460 680
rect 494 646 552 680
rect 586 646 644 680
rect 678 678 982 680
rect 678 646 734 678
rect 430 644 734 646
rect 768 644 826 678
rect 860 644 918 678
rect 952 644 982 678
<< psubdiffcont >>
rect 186 1270 220 1304
rect 274 1272 308 1306
rect 368 1268 402 1302
rect 458 1272 492 1306
rect 554 1274 588 1308
rect 644 1276 678 1310
rect 740 1274 774 1308
rect 832 1272 866 1306
rect 920 1270 954 1304
<< nsubdiffcont >>
rect 184 1904 218 1938
rect 276 1902 310 1936
rect 366 1902 400 1936
rect 462 1904 496 1938
rect 556 1906 590 1940
rect 646 1904 680 1938
rect 736 1904 770 1938
rect 826 1906 860 1940
rect 918 1904 952 1938
rect 460 646 494 680
rect 552 646 586 680
rect 644 646 678 680
rect 734 644 768 678
rect 826 644 860 678
rect 918 644 952 678
<< poly >>
rect 233 1831 263 1857
rect 317 1831 347 1857
rect 550 1831 580 1857
rect 826 1831 856 1857
rect 233 1599 263 1631
rect 175 1583 263 1599
rect 175 1549 192 1583
rect 226 1549 263 1583
rect 175 1533 263 1549
rect 233 1511 263 1533
rect 317 1599 347 1631
rect 550 1599 580 1631
rect 826 1599 856 1631
rect 317 1583 409 1599
rect 317 1549 360 1583
rect 394 1549 409 1583
rect 317 1533 409 1549
rect 494 1583 580 1599
rect 494 1549 510 1583
rect 544 1549 580 1583
rect 494 1533 580 1549
rect 770 1583 856 1599
rect 770 1549 786 1583
rect 820 1549 856 1583
rect 770 1533 856 1549
rect 317 1511 347 1533
rect 550 1511 580 1533
rect 826 1511 856 1533
rect 233 1355 263 1381
rect 317 1355 347 1381
rect 550 1355 580 1381
rect 826 1355 856 1381
rect 556 1191 586 1217
rect 832 1191 862 1217
rect 556 1039 586 1061
rect 832 1039 862 1061
rect 556 1023 642 1039
rect 556 989 592 1023
rect 626 989 642 1023
rect 556 973 642 989
rect 832 1023 918 1039
rect 832 989 868 1023
rect 902 989 918 1023
rect 832 973 918 989
rect 556 941 586 973
rect 832 941 862 973
rect 556 715 586 741
rect 832 715 862 741
<< polycont >>
rect 192 1549 226 1583
rect 360 1549 394 1583
rect 510 1549 544 1583
rect 786 1549 820 1583
rect 592 989 626 1023
rect 868 989 902 1023
<< locali >>
rect 154 1940 982 1950
rect 154 1938 556 1940
rect 154 1904 184 1938
rect 218 1936 462 1938
rect 218 1904 276 1936
rect 154 1902 276 1904
rect 310 1902 366 1936
rect 400 1904 462 1936
rect 496 1906 556 1938
rect 590 1938 826 1940
rect 590 1906 646 1938
rect 496 1904 646 1906
rect 680 1904 736 1938
rect 770 1906 826 1938
rect 860 1938 982 1940
rect 860 1906 918 1938
rect 770 1904 918 1906
rect 952 1904 982 1938
rect 400 1902 982 1904
rect 154 1895 982 1902
rect 154 1861 183 1895
rect 217 1861 275 1895
rect 309 1861 367 1895
rect 401 1861 459 1895
rect 493 1861 551 1895
rect 585 1861 643 1895
rect 677 1861 735 1895
rect 769 1861 827 1895
rect 861 1861 919 1895
rect 953 1861 982 1895
rect 171 1819 223 1861
rect 171 1785 189 1819
rect 171 1751 223 1785
rect 171 1717 189 1751
rect 171 1683 223 1717
rect 171 1649 189 1683
rect 171 1633 223 1649
rect 257 1819 323 1827
rect 257 1785 273 1819
rect 307 1785 323 1819
rect 257 1751 323 1785
rect 257 1717 273 1751
rect 307 1730 323 1751
rect 257 1696 276 1717
rect 310 1696 323 1730
rect 257 1683 323 1696
rect 257 1649 273 1683
rect 307 1649 323 1683
rect 257 1631 323 1649
rect 357 1819 413 1861
rect 391 1785 413 1819
rect 357 1751 413 1785
rect 391 1717 413 1751
rect 357 1683 413 1717
rect 391 1649 413 1683
rect 357 1633 413 1649
rect 498 1819 540 1861
rect 498 1785 506 1819
rect 498 1751 540 1785
rect 498 1717 506 1751
rect 498 1683 540 1717
rect 498 1649 506 1683
rect 498 1633 540 1649
rect 574 1819 640 1827
rect 574 1785 590 1819
rect 624 1785 640 1819
rect 574 1751 640 1785
rect 574 1717 590 1751
rect 624 1717 640 1751
rect 574 1683 640 1717
rect 574 1649 590 1683
rect 624 1649 640 1683
rect 574 1631 640 1649
rect 774 1819 816 1861
rect 774 1785 782 1819
rect 774 1751 816 1785
rect 774 1717 782 1751
rect 774 1683 816 1717
rect 774 1649 782 1683
rect 774 1633 816 1649
rect 850 1819 916 1827
rect 850 1785 866 1819
rect 900 1785 916 1819
rect 850 1751 916 1785
rect 850 1717 866 1751
rect 900 1717 916 1751
rect 850 1683 916 1717
rect 850 1649 866 1683
rect 900 1649 916 1683
rect 850 1631 916 1649
rect 175 1586 242 1599
rect 175 1552 184 1586
rect 218 1583 242 1586
rect 175 1549 192 1552
rect 226 1549 242 1583
rect 276 1511 310 1631
rect 344 1594 411 1599
rect 344 1549 360 1594
rect 394 1549 411 1594
rect 494 1592 560 1597
rect 494 1558 508 1592
rect 542 1583 560 1592
rect 494 1549 510 1558
rect 544 1549 560 1583
rect 594 1592 640 1631
rect 770 1592 836 1597
rect 594 1583 836 1592
rect 594 1552 786 1583
rect 344 1545 411 1549
rect 171 1495 310 1511
rect 171 1461 189 1495
rect 223 1461 310 1495
rect 171 1427 310 1461
rect 171 1393 189 1427
rect 223 1393 310 1427
rect 171 1385 310 1393
rect 351 1495 413 1511
rect 351 1461 357 1495
rect 391 1461 413 1495
rect 351 1427 413 1461
rect 351 1393 357 1427
rect 391 1393 413 1427
rect 351 1351 413 1393
rect 494 1499 540 1515
rect 594 1511 640 1552
rect 770 1549 786 1552
rect 820 1549 836 1583
rect 870 1590 916 1631
rect 870 1556 876 1590
rect 910 1556 916 1590
rect 494 1465 506 1499
rect 494 1431 540 1465
rect 494 1397 506 1431
rect 494 1351 540 1397
rect 574 1499 640 1511
rect 574 1465 590 1499
rect 624 1465 640 1499
rect 574 1431 640 1465
rect 574 1397 590 1431
rect 624 1397 640 1431
rect 574 1385 640 1397
rect 770 1499 816 1515
rect 870 1511 916 1556
rect 770 1465 782 1499
rect 770 1431 816 1465
rect 770 1397 782 1431
rect 770 1351 816 1397
rect 850 1499 916 1511
rect 850 1465 866 1499
rect 900 1465 916 1499
rect 850 1431 916 1465
rect 850 1397 866 1431
rect 900 1397 916 1431
rect 850 1385 916 1397
rect 154 1317 183 1351
rect 217 1317 275 1351
rect 309 1317 367 1351
rect 401 1317 459 1351
rect 493 1317 551 1351
rect 585 1317 643 1351
rect 677 1317 735 1351
rect 769 1317 827 1351
rect 861 1317 919 1351
rect 953 1317 982 1351
rect 154 1310 982 1317
rect 154 1308 644 1310
rect 154 1306 554 1308
rect 154 1304 274 1306
rect 154 1270 186 1304
rect 220 1272 274 1304
rect 308 1302 458 1306
rect 308 1272 368 1302
rect 220 1270 368 1272
rect 154 1268 368 1270
rect 402 1272 458 1302
rect 492 1274 554 1306
rect 588 1276 644 1308
rect 678 1308 982 1310
rect 678 1276 740 1308
rect 588 1274 740 1276
rect 774 1306 982 1308
rect 774 1274 832 1306
rect 492 1272 832 1274
rect 866 1304 982 1306
rect 866 1272 920 1304
rect 402 1270 920 1272
rect 954 1270 982 1304
rect 402 1268 982 1270
rect 154 1255 982 1268
rect 154 1246 459 1255
rect 430 1221 459 1246
rect 493 1221 551 1255
rect 585 1221 643 1255
rect 677 1221 735 1255
rect 769 1221 827 1255
rect 861 1221 919 1255
rect 953 1221 982 1255
rect 496 1175 562 1187
rect 496 1141 512 1175
rect 546 1141 562 1175
rect 496 1107 562 1141
rect 496 1073 512 1107
rect 546 1073 562 1107
rect 496 1061 562 1073
rect 596 1175 642 1221
rect 630 1141 642 1175
rect 596 1107 642 1141
rect 630 1073 642 1107
rect 496 1014 542 1061
rect 596 1057 642 1073
rect 772 1175 838 1187
rect 772 1141 788 1175
rect 822 1141 838 1175
rect 772 1107 838 1141
rect 772 1073 788 1107
rect 822 1073 838 1107
rect 772 1061 838 1073
rect 872 1175 918 1221
rect 906 1141 918 1175
rect 872 1107 918 1141
rect 906 1073 918 1107
rect 530 980 542 1014
rect 496 941 542 980
rect 576 989 592 1023
rect 626 1018 642 1023
rect 772 1018 818 1061
rect 872 1057 918 1073
rect 626 989 818 1018
rect 576 978 818 989
rect 576 975 642 978
rect 772 941 818 978
rect 852 989 868 1023
rect 902 1014 918 1023
rect 852 980 872 989
rect 906 980 918 1014
rect 852 975 918 980
rect 496 923 562 941
rect 496 889 512 923
rect 546 889 562 923
rect 496 855 562 889
rect 496 821 512 855
rect 546 821 562 855
rect 496 787 562 821
rect 496 753 512 787
rect 546 753 562 787
rect 496 745 562 753
rect 596 923 638 939
rect 630 889 638 923
rect 596 855 638 889
rect 630 821 638 855
rect 596 787 638 821
rect 630 753 638 787
rect 596 711 638 753
rect 772 923 838 941
rect 772 889 788 923
rect 822 889 838 923
rect 772 855 838 889
rect 772 821 788 855
rect 822 821 838 855
rect 772 787 838 821
rect 772 753 788 787
rect 822 753 838 787
rect 772 745 838 753
rect 872 923 914 939
rect 906 889 914 923
rect 872 855 914 889
rect 906 821 914 855
rect 872 787 914 821
rect 906 753 914 787
rect 872 711 914 753
rect 430 677 459 711
rect 493 680 551 711
rect 585 680 643 711
rect 677 680 735 711
rect 494 677 551 680
rect 586 677 643 680
rect 678 678 735 680
rect 769 678 827 711
rect 861 678 919 711
rect 430 646 460 677
rect 494 646 552 677
rect 586 646 644 677
rect 678 646 734 678
rect 769 677 826 678
rect 861 677 918 678
rect 953 677 982 711
rect 430 644 734 646
rect 768 644 826 677
rect 860 644 918 677
rect 952 644 982 677
<< viali >>
rect 183 1861 217 1895
rect 275 1861 309 1895
rect 367 1861 401 1895
rect 459 1861 493 1895
rect 551 1861 585 1895
rect 643 1861 677 1895
rect 735 1861 769 1895
rect 827 1861 861 1895
rect 919 1861 953 1895
rect 276 1717 307 1730
rect 307 1717 310 1730
rect 276 1696 310 1717
rect 184 1583 218 1586
rect 184 1552 192 1583
rect 192 1552 218 1583
rect 360 1583 394 1594
rect 360 1560 394 1583
rect 508 1583 542 1592
rect 508 1558 510 1583
rect 510 1558 542 1583
rect 876 1556 910 1590
rect 183 1317 217 1351
rect 275 1317 309 1351
rect 367 1317 401 1351
rect 459 1317 493 1351
rect 551 1317 585 1351
rect 643 1317 677 1351
rect 735 1317 769 1351
rect 827 1317 861 1351
rect 919 1317 953 1351
rect 459 1221 493 1255
rect 551 1221 585 1255
rect 643 1221 677 1255
rect 735 1221 769 1255
rect 827 1221 861 1255
rect 919 1221 953 1255
rect 496 980 530 1014
rect 872 989 902 1014
rect 902 989 906 1014
rect 872 980 906 989
rect 459 680 493 711
rect 551 680 585 711
rect 643 680 677 711
rect 459 677 460 680
rect 460 677 493 680
rect 551 677 552 680
rect 552 677 585 680
rect 643 677 644 680
rect 644 677 677 680
rect 735 678 769 711
rect 827 678 861 711
rect 919 678 953 711
rect 735 677 768 678
rect 768 677 769 678
rect 827 677 860 678
rect 860 677 861 678
rect 919 677 952 678
rect 952 677 953 678
<< metal1 >>
rect 974 1926 1278 1946
rect 154 1895 1278 1926
rect 154 1861 183 1895
rect 217 1861 275 1895
rect 309 1861 367 1895
rect 401 1861 459 1895
rect 493 1861 551 1895
rect 585 1861 643 1895
rect 677 1861 735 1895
rect 769 1861 827 1895
rect 861 1861 919 1895
rect 953 1861 1278 1895
rect 154 1832 1278 1861
rect 154 1830 982 1832
rect 258 1740 328 1756
rect 258 1730 552 1740
rect 258 1696 276 1730
rect 310 1696 552 1730
rect 258 1690 552 1696
rect 258 1682 328 1690
rect 66 1586 238 1602
rect 66 1552 184 1586
rect 218 1552 238 1586
rect 66 1536 238 1552
rect 342 1598 408 1606
rect 500 1598 552 1690
rect 342 1546 348 1598
rect 400 1546 408 1598
rect 494 1592 558 1598
rect 494 1558 508 1592
rect 542 1558 558 1592
rect 494 1546 558 1558
rect 854 1592 932 1602
rect 342 1542 408 1546
rect 854 1540 868 1592
rect 920 1540 932 1592
rect 854 1536 932 1540
rect 106 1382 460 1384
rect 106 1351 982 1382
rect 106 1317 183 1351
rect 217 1317 275 1351
rect 309 1317 367 1351
rect 401 1317 459 1351
rect 493 1317 551 1351
rect 585 1317 643 1351
rect 677 1317 735 1351
rect 769 1317 827 1351
rect 861 1317 919 1351
rect 953 1317 982 1351
rect 106 1255 982 1317
rect 106 1221 459 1255
rect 493 1221 551 1255
rect 585 1221 643 1255
rect 677 1221 735 1255
rect 769 1221 827 1255
rect 861 1221 919 1255
rect 953 1221 982 1255
rect 106 1190 982 1221
rect 854 1026 922 1030
rect 144 1024 542 1026
rect 144 972 352 1024
rect 404 1014 542 1024
rect 404 980 496 1014
rect 530 980 542 1014
rect 404 972 542 980
rect 144 968 542 972
rect 854 974 860 1026
rect 914 974 922 1026
rect 854 968 922 974
rect 144 966 432 968
rect 1076 742 1278 1832
rect 430 711 1278 742
rect 430 677 459 711
rect 493 677 551 711
rect 585 677 643 711
rect 677 677 735 711
rect 769 677 827 711
rect 861 677 919 711
rect 953 677 1278 711
rect 430 646 1278 677
rect 734 644 768 646
rect 972 644 1278 646
<< via1 >>
rect 348 1594 400 1598
rect 348 1560 360 1594
rect 360 1560 394 1594
rect 394 1560 400 1594
rect 348 1546 400 1560
rect 868 1590 920 1592
rect 868 1556 876 1590
rect 876 1556 910 1590
rect 910 1556 920 1590
rect 868 1540 920 1556
rect 352 972 404 1024
rect 860 1014 914 1026
rect 860 980 872 1014
rect 872 980 906 1014
rect 906 980 914 1014
rect 860 974 914 980
<< metal2 >>
rect 342 1598 408 1606
rect 342 1546 348 1598
rect 400 1566 408 1598
rect 854 1592 928 1602
rect 400 1546 414 1566
rect 342 1024 414 1546
rect 342 972 352 1024
rect 404 972 414 1024
rect 342 968 414 972
rect 854 1540 868 1592
rect 920 1540 928 1592
rect 854 1026 928 1540
rect 854 974 860 1026
rect 914 974 928 1026
rect 854 968 928 974
<< labels >>
flabel metal1 144 966 352 1026 0 FreeSans 320 0 0 0 ring_osil
port 1 nsew
flabel metal1 1076 644 1278 1946 0 FreeSans 320 0 0 0 vdd
port 2 nsew
flabel metal1 66 1536 184 1602 0 FreeSans 320 0 0 0 en
port 0 nsew
flabel metal1 106 1190 460 1384 0 FreeSans 320 0 0 0 gnd
port 5 nsew
flabel locali 276 1419 310 1453 0 FreeSans 250 0 0 0 x5.Y
flabel locali 276 1487 310 1521 0 FreeSans 250 0 0 0 x5.Y
flabel locali 276 1555 310 1589 0 FreeSans 250 0 0 0 x5.Y
flabel locali 368 1555 402 1589 0 FreeSans 250 0 0 0 x5.B
flabel locali 184 1555 218 1589 0 FreeSans 250 0 0 0 x5.A
flabel nwell 368 1861 402 1895 0 FreeSans 200 0 0 0 x5.VPB
flabel pwell 368 1317 402 1351 0 FreeSans 200 0 0 0 x5.VNB
flabel metal1 368 1317 402 1351 0 FreeSans 200 0 0 0 x5.VGND
flabel metal1 368 1861 402 1895 0 FreeSans 200 0 0 0 x5.VPWR
rlabel comment 430 1334 430 1334 6 x5.nand2_1
rlabel metal1 154 1286 430 1382 1 x5.VGND
rlabel metal1 154 1830 430 1926 1 x5.VPWR
flabel locali 508 915 542 949 0 FreeSans 340 0 0 0 x4.Y
flabel locali 508 983 542 1017 0 FreeSans 340 0 0 0 x4.Y
flabel locali 600 983 634 1017 0 FreeSans 340 0 0 0 x4.A
flabel nwell 643 677 677 711 0 FreeSans 200 0 0 0 x4.VPB
flabel pwell 643 1221 677 1255 0 FreeSans 200 0 0 0 x4.VNB
flabel metal1 643 1221 677 1255 0 FreeSans 200 0 0 0 x4.VGND
flabel metal1 643 677 677 711 0 FreeSans 200 0 0 0 x4.VPWR
rlabel comment 706 1238 706 1238 8 x4.inv_1
rlabel metal1 430 1190 706 1286 5 x4.VGND
rlabel metal1 430 646 706 742 5 x4.VPWR
flabel locali 784 915 818 949 0 FreeSans 340 0 0 0 x3.Y
flabel locali 784 983 818 1017 0 FreeSans 340 0 0 0 x3.Y
flabel locali 876 983 910 1017 0 FreeSans 340 0 0 0 x3.A
flabel nwell 919 677 953 711 0 FreeSans 200 0 0 0 x3.VPB
flabel pwell 919 1221 953 1255 0 FreeSans 200 0 0 0 x3.VNB
flabel metal1 919 1221 953 1255 0 FreeSans 200 0 0 0 x3.VGND
flabel metal1 919 677 953 711 0 FreeSans 200 0 0 0 x3.VPWR
rlabel comment 982 1238 982 1238 8 x3.inv_1
rlabel metal1 706 1190 982 1286 5 x3.VGND
rlabel metal1 706 646 982 742 5 x3.VPWR
flabel locali 870 1623 904 1657 0 FreeSans 340 0 0 0 x2.Y
flabel locali 870 1555 904 1589 0 FreeSans 340 0 0 0 x2.Y
flabel locali 778 1555 812 1589 0 FreeSans 340 0 0 0 x2.A
flabel nwell 735 1861 769 1895 0 FreeSans 200 0 0 0 x2.VPB
flabel pwell 735 1317 769 1351 0 FreeSans 200 0 0 0 x2.VNB
flabel metal1 735 1317 769 1351 0 FreeSans 200 0 0 0 x2.VGND
flabel metal1 735 1861 769 1895 0 FreeSans 200 0 0 0 x2.VPWR
rlabel comment 706 1334 706 1334 4 x2.inv_1
rlabel metal1 706 1286 982 1382 1 x2.VGND
rlabel metal1 706 1830 982 1926 1 x2.VPWR
flabel locali 594 1623 628 1657 0 FreeSans 340 0 0 0 x1.Y
flabel locali 594 1555 628 1589 0 FreeSans 340 0 0 0 x1.Y
flabel locali 502 1555 536 1589 0 FreeSans 340 0 0 0 x1.A
flabel nwell 459 1861 493 1895 0 FreeSans 200 0 0 0 x1.VPB
flabel pwell 459 1317 493 1351 0 FreeSans 200 0 0 0 x1.VNB
flabel metal1 459 1317 493 1351 0 FreeSans 200 0 0 0 x1.VGND
flabel metal1 459 1861 493 1895 0 FreeSans 200 0 0 0 x1.VPWR
rlabel comment 430 1334 430 1334 4 x1.inv_1
rlabel metal1 430 1286 706 1382 1 x1.VGND
rlabel metal1 430 1830 706 1926 1 x1.VPWR
<< end >>
