* NGSPICE file created from hgu_cdac_cap_16.ext - technology: sky130A

.subckt hgu_cdac_cap_16 SUB
C0 x1[8].CTOP x1[9].CTOP 40.4f
C1 x1[9].CTOP x1[9].CBOT 40.4f
.ends

