magic
tech sky130A
magscale 1 2
timestamp 1698238152
<< pwell >>
rect 1732 2020 1758 2052
rect 1732 998 1758 1030
<< metal3 >>
rect 1412 2692 2084 2694
rect 1412 2628 1516 2692
rect 1580 2628 1596 2692
rect 1660 2628 1676 2692
rect 1740 2628 1756 2692
rect 1820 2628 1836 2692
rect 1900 2628 1916 2692
rect 1980 2628 2084 2692
rect 1412 2626 2084 2628
rect 1412 2580 1478 2626
rect 1412 2516 1413 2580
rect 1477 2516 1478 2580
rect 1412 2500 1478 2516
rect 1412 2436 1413 2500
rect 1477 2436 1478 2500
rect 1412 2420 1478 2436
rect 1412 2356 1413 2420
rect 1477 2356 1478 2420
rect 1412 2340 1478 2356
rect 1412 2276 1413 2340
rect 1477 2276 1478 2340
rect 1412 2260 1478 2276
rect 1412 2196 1413 2260
rect 1477 2196 1478 2260
rect 1412 2180 1478 2196
rect 1412 2116 1413 2180
rect 1477 2116 1478 2180
rect 1412 2100 1478 2116
rect 1412 2036 1413 2100
rect 1477 2036 1478 2100
rect 1412 2020 1478 2036
rect 1412 1956 1413 2020
rect 1477 1956 1478 2020
rect 1412 1940 1478 1956
rect 1412 1876 1413 1940
rect 1477 1876 1478 1940
rect 1412 1860 1478 1876
rect 1412 1796 1413 1860
rect 1477 1796 1478 1860
rect 1412 1732 1478 1796
rect 1538 1732 1598 2626
rect 1658 1672 1718 2566
rect 1778 1732 1838 2626
rect 2018 2580 2084 2626
rect 1898 1672 1958 2566
rect 2018 2516 2019 2580
rect 2083 2516 2084 2580
rect 2018 2500 2084 2516
rect 2018 2436 2019 2500
rect 2083 2436 2084 2500
rect 2018 2420 2084 2436
rect 2018 2356 2019 2420
rect 2083 2356 2084 2420
rect 2018 2340 2084 2356
rect 2018 2276 2019 2340
rect 2083 2276 2084 2340
rect 2018 2260 2084 2276
rect 2018 2196 2019 2260
rect 2083 2196 2084 2260
rect 2018 2180 2084 2196
rect 2018 2116 2019 2180
rect 2083 2116 2084 2180
rect 2018 2100 2084 2116
rect 2018 2036 2019 2100
rect 2083 2036 2084 2100
rect 2018 2020 2084 2036
rect 2018 1956 2019 2020
rect 2083 1956 2084 2020
rect 2018 1940 2084 1956
rect 2018 1876 2019 1940
rect 2083 1876 2084 1940
rect 2018 1860 2084 1876
rect 2018 1796 2019 1860
rect 2083 1796 2084 1860
rect 2018 1732 2084 1796
rect 1412 1670 2084 1672
rect 1412 1606 1516 1670
rect 1580 1606 1596 1670
rect 1660 1606 1676 1670
rect 1740 1606 1756 1670
rect 1820 1606 1836 1670
rect 1900 1606 1916 1670
rect 1980 1606 2084 1670
rect 1412 1604 2084 1606
rect 1412 1558 1478 1604
rect 1412 1494 1413 1558
rect 1477 1494 1478 1558
rect 1412 1478 1478 1494
rect 1412 1414 1413 1478
rect 1477 1414 1478 1478
rect 1412 1398 1478 1414
rect 1412 1334 1413 1398
rect 1477 1334 1478 1398
rect 1412 1318 1478 1334
rect 1412 1254 1413 1318
rect 1477 1254 1478 1318
rect 1412 1238 1478 1254
rect 1412 1174 1413 1238
rect 1477 1174 1478 1238
rect 1412 1158 1478 1174
rect 1412 1094 1413 1158
rect 1477 1094 1478 1158
rect 1412 1078 1478 1094
rect 1412 1014 1413 1078
rect 1477 1014 1478 1078
rect 1412 998 1478 1014
rect 1412 934 1413 998
rect 1477 934 1478 998
rect 1412 918 1478 934
rect 1412 854 1413 918
rect 1477 854 1478 918
rect 1412 838 1478 854
rect 1412 774 1413 838
rect 1477 774 1478 838
rect 1412 710 1478 774
rect 1538 710 1598 1604
rect 1658 650 1718 1544
rect 1778 710 1838 1604
rect 2018 1558 2084 1604
rect 1898 650 1958 1544
rect 2018 1494 2019 1558
rect 2083 1494 2084 1558
rect 2018 1478 2084 1494
rect 2018 1414 2019 1478
rect 2083 1414 2084 1478
rect 2018 1398 2084 1414
rect 2018 1334 2019 1398
rect 2083 1334 2084 1398
rect 2018 1318 2084 1334
rect 2018 1254 2019 1318
rect 2083 1254 2084 1318
rect 2018 1238 2084 1254
rect 2018 1174 2019 1238
rect 2083 1174 2084 1238
rect 2018 1158 2084 1174
rect 2018 1094 2019 1158
rect 2083 1094 2084 1158
rect 2018 1078 2084 1094
rect 2018 1014 2019 1078
rect 2083 1014 2084 1078
rect 2018 998 2084 1014
rect 2018 934 2019 998
rect 2083 934 2084 998
rect 2018 918 2084 934
rect 2018 854 2019 918
rect 2083 854 2084 918
rect 2018 838 2084 854
rect 2018 774 2019 838
rect 2083 774 2084 838
rect 2018 710 2084 774
rect 1538 648 1958 650
rect 1538 584 1596 648
rect 1660 584 1676 648
rect 1740 584 1756 648
rect 1820 584 1836 648
rect 1900 584 1958 648
rect 1538 582 1958 584
<< via3 >>
rect 1516 2628 1580 2692
rect 1596 2628 1660 2692
rect 1676 2628 1740 2692
rect 1756 2628 1820 2692
rect 1836 2628 1900 2692
rect 1916 2628 1980 2692
rect 1413 2516 1477 2580
rect 1413 2436 1477 2500
rect 1413 2356 1477 2420
rect 1413 2276 1477 2340
rect 1413 2196 1477 2260
rect 1413 2116 1477 2180
rect 1413 2036 1477 2100
rect 1413 1956 1477 2020
rect 1413 1876 1477 1940
rect 1413 1796 1477 1860
rect 2019 2516 2083 2580
rect 2019 2436 2083 2500
rect 2019 2356 2083 2420
rect 2019 2276 2083 2340
rect 2019 2196 2083 2260
rect 2019 2116 2083 2180
rect 2019 2036 2083 2100
rect 2019 1956 2083 2020
rect 2019 1876 2083 1940
rect 2019 1796 2083 1860
rect 1516 1606 1580 1670
rect 1596 1606 1660 1670
rect 1676 1606 1740 1670
rect 1756 1606 1820 1670
rect 1836 1606 1900 1670
rect 1916 1606 1980 1670
rect 1413 1494 1477 1558
rect 1413 1414 1477 1478
rect 1413 1334 1477 1398
rect 1413 1254 1477 1318
rect 1413 1174 1477 1238
rect 1413 1094 1477 1158
rect 1413 1014 1477 1078
rect 1413 934 1477 998
rect 1413 854 1477 918
rect 1413 774 1477 838
rect 2019 1494 2083 1558
rect 2019 1414 2083 1478
rect 2019 1334 2083 1398
rect 2019 1254 2083 1318
rect 2019 1174 2083 1238
rect 2019 1094 2083 1158
rect 2019 1014 2083 1078
rect 2019 934 2083 998
rect 2019 854 2083 918
rect 2019 774 2083 838
rect 1596 584 1660 648
rect 1676 584 1740 648
rect 1756 584 1820 648
rect 1836 584 1900 648
<< metal4 >>
rect 1412 2692 2084 2694
rect 1412 2628 1516 2692
rect 1580 2628 1596 2692
rect 1660 2628 1676 2692
rect 1740 2628 1756 2692
rect 1820 2628 1836 2692
rect 1900 2628 1916 2692
rect 1980 2628 2084 2692
rect 1412 2626 2084 2628
rect 1412 2580 1478 2626
rect 1412 2516 1413 2580
rect 1477 2516 1478 2580
rect 1412 2500 1478 2516
rect 1412 2436 1413 2500
rect 1477 2436 1478 2500
rect 1412 2420 1478 2436
rect 1412 2356 1413 2420
rect 1477 2356 1478 2420
rect 1412 2340 1478 2356
rect 1412 2276 1413 2340
rect 1477 2276 1478 2340
rect 1412 2260 1478 2276
rect 1412 2196 1413 2260
rect 1477 2196 1478 2260
rect 1412 2180 1478 2196
rect 1412 2116 1413 2180
rect 1477 2116 1478 2180
rect 1412 2100 1478 2116
rect 1412 2036 1413 2100
rect 1477 2036 1478 2100
rect 1412 2020 1478 2036
rect 1412 1956 1413 2020
rect 1477 1956 1478 2020
rect 1412 1940 1478 1956
rect 1412 1876 1413 1940
rect 1477 1876 1478 1940
rect 1412 1860 1478 1876
rect 1412 1796 1413 1860
rect 1477 1796 1478 1860
rect 1412 1732 1478 1796
rect 1538 1672 1598 2566
rect 1658 1732 1718 2626
rect 1778 1672 1838 2566
rect 1898 1732 1958 2626
rect 2018 2580 2084 2626
rect 2018 2516 2019 2580
rect 2083 2516 2084 2580
rect 2018 2500 2084 2516
rect 2018 2436 2019 2500
rect 2083 2436 2084 2500
rect 2018 2420 2084 2436
rect 2018 2356 2019 2420
rect 2083 2356 2084 2420
rect 2018 2340 2084 2356
rect 2018 2276 2019 2340
rect 2083 2276 2084 2340
rect 2018 2260 2084 2276
rect 2018 2196 2019 2260
rect 2083 2196 2084 2260
rect 2018 2180 2084 2196
rect 2018 2116 2019 2180
rect 2083 2116 2084 2180
rect 2018 2100 2084 2116
rect 2018 2036 2019 2100
rect 2083 2036 2084 2100
rect 2018 2020 2084 2036
rect 2018 1956 2019 2020
rect 2083 1956 2084 2020
rect 2018 1940 2084 1956
rect 2018 1876 2019 1940
rect 2083 1876 2084 1940
rect 2018 1860 2084 1876
rect 2018 1796 2019 1860
rect 2083 1796 2084 1860
rect 2018 1732 2084 1796
rect 1412 1670 2084 1672
rect 1412 1606 1516 1670
rect 1580 1606 1596 1670
rect 1660 1606 1676 1670
rect 1740 1606 1756 1670
rect 1820 1606 1836 1670
rect 1900 1606 1916 1670
rect 1980 1606 2084 1670
rect 1412 1604 2084 1606
rect 1412 1558 1478 1604
rect 1412 1494 1413 1558
rect 1477 1494 1478 1558
rect 1412 1478 1478 1494
rect 1412 1414 1413 1478
rect 1477 1414 1478 1478
rect 1412 1398 1478 1414
rect 1412 1334 1413 1398
rect 1477 1334 1478 1398
rect 1412 1318 1478 1334
rect 1412 1254 1413 1318
rect 1477 1254 1478 1318
rect 1412 1238 1478 1254
rect 1412 1174 1413 1238
rect 1477 1174 1478 1238
rect 1412 1158 1478 1174
rect 1412 1094 1413 1158
rect 1477 1094 1478 1158
rect 1412 1078 1478 1094
rect 1412 1014 1413 1078
rect 1477 1014 1478 1078
rect 1412 998 1478 1014
rect 1412 934 1413 998
rect 1477 934 1478 998
rect 1412 918 1478 934
rect 1412 854 1413 918
rect 1477 854 1478 918
rect 1412 838 1478 854
rect 1412 774 1413 838
rect 1477 774 1478 838
rect 1412 710 1478 774
rect 1538 650 1598 1544
rect 1658 710 1718 1604
rect 1778 650 1838 1544
rect 1898 710 1958 1604
rect 2018 1558 2084 1604
rect 2018 1494 2019 1558
rect 2083 1494 2084 1558
rect 2018 1478 2084 1494
rect 2018 1414 2019 1478
rect 2083 1414 2084 1478
rect 2018 1398 2084 1414
rect 2018 1334 2019 1398
rect 2083 1334 2084 1398
rect 2018 1318 2084 1334
rect 2018 1254 2019 1318
rect 2083 1254 2084 1318
rect 2018 1238 2084 1254
rect 2018 1174 2019 1238
rect 2083 1174 2084 1238
rect 2018 1158 2084 1174
rect 2018 1094 2019 1158
rect 2083 1094 2084 1158
rect 2018 1078 2084 1094
rect 2018 1014 2019 1078
rect 2083 1014 2084 1078
rect 2018 998 2084 1014
rect 2018 934 2019 998
rect 2083 934 2084 998
rect 2018 918 2084 934
rect 2018 854 2019 918
rect 2083 854 2084 918
rect 2018 838 2084 854
rect 2018 774 2019 838
rect 2083 774 2084 838
rect 2018 710 2084 774
rect 1538 648 1958 650
rect 1538 584 1596 648
rect 1660 584 1676 648
rect 1740 584 1756 648
rect 1820 584 1836 648
rect 1900 584 1958 648
rect 1538 582 1958 584
<< labels >>
flabel space 1732 2022 1758 2054 0 FreeSans 160 0 0 0 hgu_cdac_unit_0.SUB
flabel metal4 1674 2354 1700 2386 0 FreeSans 320 0 0 0 hgu_cdac_unit_0.C1
flabel metal4 1792 1764 1818 1796 0 FreeSans 320 0 0 0 hgu_cdac_unit_0.C0
flabel space 1732 1000 1758 1032 0 FreeSans 160 0 0 0 hgu_cdac_unit_1.SUB
flabel metal4 1674 1332 1700 1364 0 FreeSans 320 0 0 0 hgu_cdac_unit_1.C1
flabel metal4 1792 742 1818 774 0 FreeSans 320 0 0 0 hgu_cdac_unit_1.C0
<< end >>
