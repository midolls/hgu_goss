magic
tech sky130A
magscale 1 2
timestamp 1699610509
<< nwell >>
rect 948 3799 1858 5355
rect 948 297 1858 1853
<< nmos >>
rect 1148 2961 1178 3511
rect 1244 2961 1274 3511
rect 1340 2961 1370 3511
rect 1436 2961 1466 3511
rect 1532 2961 1562 3511
rect 1628 2961 1658 3511
rect 1148 2141 1178 2691
rect 1244 2141 1274 2691
rect 1340 2141 1370 2691
rect 1436 2141 1466 2691
rect 1532 2141 1562 2691
rect 1628 2141 1658 2691
<< pmos >>
rect 1148 4036 1178 5136
rect 1244 4036 1274 5136
rect 1340 4036 1370 5136
rect 1436 4036 1466 5136
rect 1532 4036 1562 5136
rect 1628 4036 1658 5136
rect 1148 516 1178 1616
rect 1244 516 1274 1616
rect 1340 516 1370 1616
rect 1436 516 1466 1616
rect 1532 516 1562 1616
rect 1628 516 1658 1616
<< ndiff >>
rect 1086 3499 1148 3511
rect 1086 2973 1098 3499
rect 1132 2973 1148 3499
rect 1086 2961 1148 2973
rect 1178 3499 1244 3511
rect 1178 2973 1194 3499
rect 1228 2973 1244 3499
rect 1178 2961 1244 2973
rect 1274 3499 1340 3511
rect 1274 2973 1290 3499
rect 1324 2973 1340 3499
rect 1274 2961 1340 2973
rect 1370 3499 1436 3511
rect 1370 2973 1386 3499
rect 1420 2973 1436 3499
rect 1370 2961 1436 2973
rect 1466 3499 1532 3511
rect 1466 2973 1482 3499
rect 1516 2973 1532 3499
rect 1466 2961 1532 2973
rect 1562 3499 1628 3511
rect 1562 2973 1578 3499
rect 1612 2973 1628 3499
rect 1562 2961 1628 2973
rect 1658 3499 1720 3511
rect 1658 2973 1674 3499
rect 1708 2973 1720 3499
rect 1658 2961 1720 2973
rect 1086 2679 1148 2691
rect 1086 2153 1098 2679
rect 1132 2153 1148 2679
rect 1086 2141 1148 2153
rect 1178 2679 1244 2691
rect 1178 2153 1194 2679
rect 1228 2153 1244 2679
rect 1178 2141 1244 2153
rect 1274 2679 1340 2691
rect 1274 2153 1290 2679
rect 1324 2153 1340 2679
rect 1274 2141 1340 2153
rect 1370 2679 1436 2691
rect 1370 2153 1386 2679
rect 1420 2153 1436 2679
rect 1370 2141 1436 2153
rect 1466 2679 1532 2691
rect 1466 2153 1482 2679
rect 1516 2153 1532 2679
rect 1466 2141 1532 2153
rect 1562 2679 1628 2691
rect 1562 2153 1578 2679
rect 1612 2153 1628 2679
rect 1562 2141 1628 2153
rect 1658 2679 1720 2691
rect 1658 2153 1674 2679
rect 1708 2153 1720 2679
rect 1658 2141 1720 2153
<< pdiff >>
rect 1086 5124 1148 5136
rect 1086 4048 1098 5124
rect 1132 4048 1148 5124
rect 1086 4036 1148 4048
rect 1178 5124 1244 5136
rect 1178 4048 1194 5124
rect 1228 4048 1244 5124
rect 1178 4036 1244 4048
rect 1274 5124 1340 5136
rect 1274 4048 1290 5124
rect 1324 4048 1340 5124
rect 1274 4036 1340 4048
rect 1370 5124 1436 5136
rect 1370 4048 1386 5124
rect 1420 4048 1436 5124
rect 1370 4036 1436 4048
rect 1466 5124 1532 5136
rect 1466 4048 1482 5124
rect 1516 4048 1532 5124
rect 1466 4036 1532 4048
rect 1562 5124 1628 5136
rect 1562 4048 1578 5124
rect 1612 4048 1628 5124
rect 1562 4036 1628 4048
rect 1658 5124 1720 5136
rect 1658 4048 1674 5124
rect 1708 4048 1720 5124
rect 1658 4036 1720 4048
rect 1086 1604 1148 1616
rect 1086 528 1098 1604
rect 1132 528 1148 1604
rect 1086 516 1148 528
rect 1178 1604 1244 1616
rect 1178 528 1194 1604
rect 1228 528 1244 1604
rect 1178 516 1244 528
rect 1274 1604 1340 1616
rect 1274 528 1290 1604
rect 1324 528 1340 1604
rect 1274 516 1340 528
rect 1370 1604 1436 1616
rect 1370 528 1386 1604
rect 1420 528 1436 1604
rect 1370 516 1436 528
rect 1466 1604 1532 1616
rect 1466 528 1482 1604
rect 1516 528 1532 1604
rect 1466 516 1532 528
rect 1562 1604 1628 1616
rect 1562 528 1578 1604
rect 1612 528 1628 1604
rect 1562 516 1628 528
rect 1658 1604 1720 1616
rect 1658 528 1674 1604
rect 1708 528 1720 1604
rect 1658 516 1720 528
<< ndiffc >>
rect 1098 2973 1132 3499
rect 1194 2973 1228 3499
rect 1290 2973 1324 3499
rect 1386 2973 1420 3499
rect 1482 2973 1516 3499
rect 1578 2973 1612 3499
rect 1674 2973 1708 3499
rect 1098 2153 1132 2679
rect 1194 2153 1228 2679
rect 1290 2153 1324 2679
rect 1386 2153 1420 2679
rect 1482 2153 1516 2679
rect 1578 2153 1612 2679
rect 1674 2153 1708 2679
<< pdiffc >>
rect 1098 4048 1132 5124
rect 1194 4048 1228 5124
rect 1290 4048 1324 5124
rect 1386 4048 1420 5124
rect 1482 4048 1516 5124
rect 1578 4048 1612 5124
rect 1674 4048 1708 5124
rect 1098 528 1132 1604
rect 1194 528 1228 1604
rect 1290 528 1324 1604
rect 1386 528 1420 1604
rect 1482 528 1516 1604
rect 1578 528 1612 1604
rect 1674 528 1708 1604
<< psubdiff >>
rect 984 3684 1090 3718
rect 1140 3684 1186 3718
rect 1236 3684 1282 3718
rect 1332 3684 1378 3718
rect 1428 3684 1474 3718
rect 1524 3684 1570 3718
rect 1620 3684 1666 3718
rect 1716 3684 1822 3718
rect 984 3611 1018 3684
rect 1788 3611 1822 3684
rect 984 2843 1018 2905
rect 1788 2843 1822 2905
rect 984 2809 1090 2843
rect 1140 2809 1186 2843
rect 1236 2809 1282 2843
rect 1332 2809 1378 2843
rect 1428 2809 1474 2843
rect 1524 2809 1570 2843
rect 1620 2809 1666 2843
rect 1716 2809 1822 2843
rect 984 2747 1018 2809
rect 1788 2747 1822 2809
rect 984 1968 1018 2041
rect 1788 1968 1822 2041
rect 984 1934 1090 1968
rect 1140 1934 1186 1968
rect 1236 1934 1282 1968
rect 1332 1934 1378 1968
rect 1428 1934 1474 1968
rect 1524 1934 1570 1968
rect 1620 1934 1666 1968
rect 1716 1934 1822 1968
<< nsubdiff >>
rect 984 5285 1090 5319
rect 1140 5285 1186 5319
rect 1236 5285 1282 5319
rect 1332 5285 1378 5319
rect 1428 5285 1474 5319
rect 1524 5285 1570 5319
rect 1620 5285 1666 5319
rect 1716 5285 1819 5319
rect 984 5223 1018 5285
rect 1785 5223 1819 5285
rect 984 3869 1018 3992
rect 1785 3869 1819 3991
rect 984 3835 1090 3869
rect 1140 3835 1186 3869
rect 1236 3835 1282 3869
rect 1332 3835 1378 3869
rect 1428 3835 1474 3869
rect 1524 3835 1570 3869
rect 1620 3835 1666 3869
rect 1716 3835 1819 3869
rect 984 1783 1090 1817
rect 1140 1783 1186 1817
rect 1236 1783 1282 1817
rect 1332 1783 1378 1817
rect 1428 1783 1474 1817
rect 1524 1783 1570 1817
rect 1620 1783 1666 1817
rect 1716 1783 1819 1817
rect 984 1660 1018 1783
rect 1785 1661 1819 1783
rect 984 367 1018 429
rect 1785 367 1819 429
rect 984 333 1090 367
rect 1140 333 1186 367
rect 1236 333 1282 367
rect 1332 333 1378 367
rect 1428 333 1474 367
rect 1524 333 1570 367
rect 1620 333 1666 367
rect 1716 333 1819 367
<< psubdiffcont >>
rect 1090 3684 1140 3718
rect 1186 3684 1236 3718
rect 1282 3684 1332 3718
rect 1378 3684 1428 3718
rect 1474 3684 1524 3718
rect 1570 3684 1620 3718
rect 1666 3684 1716 3718
rect 984 2905 1018 3611
rect 1788 2905 1822 3611
rect 1090 2809 1140 2843
rect 1186 2809 1236 2843
rect 1282 2809 1332 2843
rect 1378 2809 1428 2843
rect 1474 2809 1524 2843
rect 1570 2809 1620 2843
rect 1666 2809 1716 2843
rect 984 2041 1018 2747
rect 1788 2041 1822 2747
rect 1090 1934 1140 1968
rect 1186 1934 1236 1968
rect 1282 1934 1332 1968
rect 1378 1934 1428 1968
rect 1474 1934 1524 1968
rect 1570 1934 1620 1968
rect 1666 1934 1716 1968
<< nsubdiffcont >>
rect 1090 5285 1140 5319
rect 1186 5285 1236 5319
rect 1282 5285 1332 5319
rect 1378 5285 1428 5319
rect 1474 5285 1524 5319
rect 1570 5285 1620 5319
rect 1666 5285 1716 5319
rect 984 3992 1018 5223
rect 1785 3991 1819 5223
rect 1090 3835 1140 3869
rect 1186 3835 1236 3869
rect 1282 3835 1332 3869
rect 1378 3835 1428 3869
rect 1474 3835 1524 3869
rect 1570 3835 1620 3869
rect 1666 3835 1716 3869
rect 1090 1783 1140 1817
rect 1186 1783 1236 1817
rect 1282 1783 1332 1817
rect 1378 1783 1428 1817
rect 1474 1783 1524 1817
rect 1570 1783 1620 1817
rect 1666 1783 1716 1817
rect 984 429 1018 1660
rect 1785 429 1819 1661
rect 1090 333 1140 367
rect 1186 333 1236 367
rect 1282 333 1332 367
rect 1378 333 1428 367
rect 1474 333 1524 367
rect 1570 333 1620 367
rect 1666 333 1716 367
<< poly >>
rect 1148 5162 1466 5192
rect 1148 5136 1178 5162
rect 1244 5136 1274 5162
rect 1340 5136 1370 5162
rect 1436 5136 1466 5162
rect 1532 5162 1658 5192
rect 1532 5136 1562 5162
rect 1628 5136 1658 5162
rect 1148 4010 1178 4036
rect 1244 4010 1274 4036
rect 1340 4010 1370 4036
rect 1436 4010 1466 4036
rect 1532 4010 1562 4036
rect 1628 4010 1658 4036
rect 1148 3979 1475 4010
rect 1440 3966 1475 3979
rect 1628 3989 1694 4010
rect 1440 3950 1507 3966
rect 1440 3916 1457 3950
rect 1491 3916 1507 3950
rect 1628 3955 1644 3989
rect 1678 3955 1694 3989
rect 1628 3943 1694 3955
rect 1440 3900 1507 3916
rect 1476 3631 1543 3647
rect 1476 3611 1493 3631
rect 1436 3597 1493 3611
rect 1527 3597 1543 3631
rect 1436 3581 1543 3597
rect 1617 3626 1684 3642
rect 1617 3592 1633 3626
rect 1667 3592 1684 3626
rect 1436 3568 1466 3581
rect 1617 3576 1684 3592
rect 1148 3537 1466 3568
rect 1148 3511 1178 3537
rect 1244 3511 1274 3537
rect 1340 3511 1370 3537
rect 1436 3511 1466 3537
rect 1532 3511 1562 3537
rect 1628 3511 1658 3576
rect 1148 2935 1178 2961
rect 1244 2935 1274 2961
rect 1340 2935 1370 2961
rect 1436 2935 1466 2961
rect 1532 2935 1562 2961
rect 1628 2935 1658 2961
rect 1532 2905 1658 2935
rect 1532 2717 1658 2747
rect 1148 2691 1178 2717
rect 1244 2691 1274 2717
rect 1340 2691 1370 2717
rect 1436 2691 1466 2717
rect 1532 2691 1562 2717
rect 1628 2691 1658 2717
rect 1148 2115 1178 2141
rect 1244 2115 1274 2141
rect 1340 2115 1370 2141
rect 1436 2115 1466 2141
rect 1532 2115 1562 2141
rect 1148 2084 1466 2115
rect 1436 2071 1466 2084
rect 1628 2076 1658 2141
rect 1436 2055 1543 2071
rect 1436 2041 1493 2055
rect 1476 2021 1493 2041
rect 1527 2021 1543 2055
rect 1476 2005 1543 2021
rect 1617 2060 1684 2076
rect 1617 2026 1633 2060
rect 1667 2026 1684 2060
rect 1617 2010 1684 2026
rect 1440 1736 1507 1752
rect 1440 1702 1457 1736
rect 1491 1702 1507 1736
rect 1440 1686 1507 1702
rect 1628 1697 1694 1709
rect 1440 1673 1475 1686
rect 1148 1642 1475 1673
rect 1628 1663 1644 1697
rect 1678 1663 1694 1697
rect 1628 1642 1694 1663
rect 1148 1616 1178 1642
rect 1244 1616 1274 1642
rect 1340 1616 1370 1642
rect 1436 1616 1466 1642
rect 1532 1616 1562 1642
rect 1628 1616 1658 1642
rect 1148 491 1178 516
rect 1244 491 1274 516
rect 1340 491 1370 516
rect 1436 491 1466 516
rect 1148 460 1475 491
rect 1532 490 1562 516
rect 1628 490 1658 516
rect 1532 460 1658 490
<< polycont >>
rect 1457 3916 1491 3950
rect 1644 3955 1678 3989
rect 1493 3597 1527 3631
rect 1633 3592 1667 3626
rect 1493 2021 1527 2055
rect 1633 2026 1667 2060
rect 1457 1702 1491 1736
rect 1644 1663 1678 1697
<< locali >>
rect 984 5285 1090 5319
rect 1140 5285 1186 5319
rect 1236 5285 1282 5319
rect 1332 5285 1378 5319
rect 1428 5285 1474 5319
rect 1524 5285 1570 5319
rect 1620 5285 1666 5319
rect 1716 5285 1819 5319
rect 984 5223 1018 5285
rect 1785 5223 1819 5285
rect 1098 5124 1132 5140
rect 1098 4032 1132 4048
rect 1194 5124 1228 5140
rect 1194 4032 1228 4048
rect 1290 5124 1324 5140
rect 1290 4032 1324 4048
rect 1386 5124 1420 5140
rect 1386 4032 1420 4048
rect 1482 5124 1516 5140
rect 1482 4032 1516 4048
rect 1578 5124 1612 5140
rect 1578 4032 1612 4048
rect 1674 5124 1708 5140
rect 1674 4032 1708 4048
rect 984 3872 1018 3992
rect 1628 3955 1644 3989
rect 1678 3955 1694 3989
rect 1441 3916 1457 3950
rect 1491 3916 1507 3950
rect 1785 3869 1819 3991
rect 1018 3838 1090 3869
rect 984 3835 1090 3838
rect 1140 3835 1186 3869
rect 1236 3835 1282 3869
rect 1332 3835 1378 3869
rect 1428 3835 1474 3869
rect 1524 3835 1570 3869
rect 1620 3835 1666 3869
rect 1716 3835 1819 3869
rect 984 3684 1090 3718
rect 1140 3684 1186 3718
rect 1236 3684 1282 3718
rect 1332 3684 1378 3718
rect 1428 3684 1474 3718
rect 1524 3684 1570 3718
rect 1620 3684 1666 3718
rect 1716 3684 1822 3718
rect 984 3611 1018 3684
rect 1477 3597 1493 3631
rect 1527 3597 1543 3631
rect 1633 3626 1667 3642
rect 1633 3576 1667 3592
rect 1788 3611 1822 3684
rect 1098 3499 1132 3515
rect 1098 2957 1132 2973
rect 1194 3499 1228 3515
rect 1194 2957 1228 2973
rect 1290 3499 1324 3515
rect 1290 2957 1324 2973
rect 1386 3499 1420 3515
rect 1386 2957 1420 2973
rect 1482 3499 1516 3515
rect 1482 2957 1516 2973
rect 1578 3499 1612 3515
rect 1578 2957 1612 2973
rect 1674 3499 1708 3515
rect 1674 2957 1708 2973
rect 984 2843 1018 2905
rect 1788 2843 1822 2905
rect 984 2809 1090 2843
rect 1140 2809 1186 2843
rect 1236 2809 1282 2843
rect 1332 2809 1378 2843
rect 1428 2809 1474 2843
rect 1524 2809 1570 2843
rect 1620 2809 1666 2843
rect 1716 2809 1822 2843
rect 984 2747 1018 2809
rect 1788 2747 1822 2809
rect 1098 2679 1132 2695
rect 1098 2137 1132 2153
rect 1194 2679 1228 2695
rect 1194 2137 1228 2153
rect 1290 2679 1324 2695
rect 1290 2137 1324 2153
rect 1386 2679 1420 2695
rect 1386 2137 1420 2153
rect 1482 2679 1516 2695
rect 1482 2137 1516 2153
rect 1578 2679 1612 2695
rect 1578 2137 1612 2153
rect 1674 2679 1708 2695
rect 1674 2137 1708 2153
rect 1633 2060 1667 2076
rect 984 1968 1018 2041
rect 1477 2021 1493 2055
rect 1527 2021 1543 2055
rect 1633 2010 1667 2026
rect 1788 1968 1822 2041
rect 984 1934 1090 1968
rect 1140 1934 1186 1968
rect 1236 1934 1282 1968
rect 1332 1934 1378 1968
rect 1428 1934 1474 1968
rect 1524 1934 1570 1968
rect 1620 1934 1666 1968
rect 1716 1934 1822 1968
rect 1018 1783 1090 1817
rect 1140 1783 1186 1817
rect 1236 1783 1282 1817
rect 1332 1783 1378 1817
rect 1428 1783 1474 1817
rect 1524 1783 1570 1817
rect 1620 1783 1666 1817
rect 1716 1783 1819 1817
rect 984 1660 1018 1783
rect 1441 1702 1457 1736
rect 1491 1702 1507 1736
rect 1628 1663 1644 1697
rect 1678 1663 1694 1697
rect 1785 1661 1819 1783
rect 1098 1604 1132 1620
rect 1098 512 1132 528
rect 1194 1604 1228 1620
rect 1194 512 1228 528
rect 1290 1604 1324 1620
rect 1290 512 1324 528
rect 1386 1604 1420 1620
rect 1386 512 1420 528
rect 1482 1604 1516 1620
rect 1482 512 1516 528
rect 1578 1604 1612 1620
rect 1578 512 1612 528
rect 1674 1604 1708 1620
rect 1674 512 1708 528
rect 984 367 1018 429
rect 1785 367 1819 429
rect 984 333 1090 367
rect 1140 333 1186 367
rect 1236 333 1282 367
rect 1332 333 1378 367
rect 1428 333 1474 367
rect 1524 333 1570 367
rect 1620 333 1666 367
rect 1716 333 1819 367
<< viali >>
rect 1098 4048 1132 5124
rect 1194 4048 1228 5124
rect 1290 4048 1324 5124
rect 1386 4048 1420 5124
rect 1482 4048 1516 5124
rect 1578 4048 1612 5124
rect 1674 4048 1708 5124
rect 1644 3955 1678 3989
rect 1457 3916 1491 3950
rect 984 3838 1018 3872
rect 1493 3597 1527 3631
rect 1633 3592 1667 3626
rect 1098 2973 1132 3499
rect 1194 2973 1228 3499
rect 1290 2973 1324 3499
rect 1386 2973 1420 3499
rect 1482 2973 1516 3499
rect 1578 2973 1612 3499
rect 1674 2973 1708 3499
rect 1098 2153 1132 2679
rect 1194 2153 1228 2679
rect 1290 2153 1324 2679
rect 1386 2153 1420 2679
rect 1482 2153 1516 2679
rect 1578 2153 1612 2679
rect 1674 2153 1708 2679
rect 1493 2021 1527 2055
rect 1633 2026 1667 2060
rect 984 1783 1018 1817
rect 1457 1702 1491 1736
rect 1644 1663 1678 1697
rect 1098 528 1132 1604
rect 1194 528 1228 1604
rect 1290 528 1324 1604
rect 1386 528 1420 1604
rect 1482 528 1516 1604
rect 1578 528 1612 1604
rect 1674 528 1708 1604
<< metal1 >>
rect 1098 5175 1708 5209
rect 1098 5136 1132 5175
rect 1674 5136 1708 5175
rect 1092 5124 1138 5136
rect 1092 4048 1098 5124
rect 1132 4048 1138 5124
rect 1092 4036 1138 4048
rect 1188 5124 1234 5136
rect 1188 4048 1194 5124
rect 1228 4048 1234 5124
rect 1188 4036 1234 4048
rect 1284 5124 1330 5136
rect 1284 4048 1290 5124
rect 1324 4048 1330 5124
rect 1284 4036 1330 4048
rect 1380 5124 1426 5136
rect 1380 4048 1386 5124
rect 1420 4048 1426 5124
rect 1380 4036 1426 4048
rect 1476 5124 1522 5136
rect 1476 4048 1482 5124
rect 1516 4048 1522 5124
rect 1476 4036 1522 4048
rect 1572 5124 1618 5136
rect 1572 4048 1578 5124
rect 1612 4048 1618 5124
rect 1572 4036 1618 4048
rect 1668 5124 1714 5136
rect 1668 4048 1674 5124
rect 1708 4070 1714 5124
rect 1708 4048 1799 4070
rect 1668 4036 1799 4048
rect 1194 4002 1228 4036
rect 1386 4002 1420 4036
rect 1194 3974 1420 4002
rect 1635 4002 1687 4008
rect 751 3903 877 3913
rect 751 3797 761 3903
rect 867 3879 877 3903
rect 867 3872 1030 3879
rect 867 3838 984 3872
rect 1018 3838 1030 3872
rect 867 3831 1030 3838
rect 867 3797 877 3831
rect 751 3787 877 3797
rect 1289 3573 1323 3974
rect 1448 3959 1500 3965
rect 1631 3955 1635 3989
rect 1687 3955 1691 3989
rect 1444 3916 1448 3950
rect 1500 3916 1504 3950
rect 1635 3944 1687 3950
rect 1448 3901 1500 3907
rect 1484 3640 1536 3646
rect 1633 3635 1667 3639
rect 1480 3597 1484 3631
rect 1536 3597 1540 3631
rect 1484 3582 1536 3588
rect 1618 3583 1624 3635
rect 1676 3583 1682 3635
rect 1633 3579 1667 3583
rect 1194 3539 1420 3573
rect 1194 3511 1228 3539
rect 1386 3511 1420 3539
rect 1765 3511 1799 4036
rect 1092 3499 1138 3511
rect 1092 2973 1098 3499
rect 1132 2973 1138 3499
rect 1092 2961 1138 2973
rect 1188 3499 1234 3511
rect 1188 2973 1194 3499
rect 1228 2973 1234 3499
rect 1188 2961 1234 2973
rect 1284 3499 1330 3511
rect 1284 2973 1290 3499
rect 1324 2973 1330 3499
rect 1284 2961 1330 2973
rect 1380 3499 1426 3511
rect 1380 2973 1386 3499
rect 1420 2973 1426 3499
rect 1380 2961 1426 2973
rect 1476 3499 1522 3511
rect 1476 2973 1482 3499
rect 1516 2973 1522 3499
rect 1476 2961 1522 2973
rect 1572 3499 1618 3511
rect 1572 2973 1578 3499
rect 1612 2973 1618 3499
rect 1572 2961 1618 2973
rect 1668 3499 1799 3511
rect 1668 2973 1674 3499
rect 1708 3476 1799 3499
rect 1708 2973 1714 3476
rect 1668 2961 1714 2973
rect 1098 2922 1132 2961
rect 1290 2922 1324 2961
rect 1482 2922 1516 2961
rect 1578 2922 1612 2961
rect 1674 2922 1708 2961
rect 1098 2888 1708 2922
rect 1098 2730 1708 2764
rect 1098 2691 1132 2730
rect 1290 2691 1324 2730
rect 1482 2691 1516 2730
rect 1578 2691 1612 2730
rect 1674 2691 1708 2730
rect 1092 2679 1138 2691
rect 1092 2153 1098 2679
rect 1132 2153 1138 2679
rect 1092 2141 1138 2153
rect 1188 2679 1234 2691
rect 1188 2153 1194 2679
rect 1228 2153 1234 2679
rect 1188 2141 1234 2153
rect 1284 2679 1330 2691
rect 1284 2153 1290 2679
rect 1324 2153 1330 2679
rect 1284 2141 1330 2153
rect 1380 2679 1426 2691
rect 1380 2153 1386 2679
rect 1420 2153 1426 2679
rect 1380 2141 1426 2153
rect 1476 2679 1522 2691
rect 1476 2153 1482 2679
rect 1516 2153 1522 2679
rect 1476 2141 1522 2153
rect 1572 2679 1618 2691
rect 1572 2153 1578 2679
rect 1612 2153 1618 2679
rect 1572 2141 1618 2153
rect 1668 2679 1714 2691
rect 1668 2153 1674 2679
rect 1708 2175 1714 2679
rect 1708 2153 1785 2175
rect 1668 2141 1785 2153
rect 1194 2113 1228 2141
rect 1386 2113 1420 2141
rect 1194 2079 1420 2113
rect 748 1847 874 1857
rect 748 1741 758 1847
rect 864 1829 874 1847
rect 864 1817 1030 1829
rect 864 1783 984 1817
rect 1018 1783 1030 1817
rect 864 1771 1030 1783
rect 864 1741 874 1771
rect 748 1731 874 1741
rect 1289 1678 1323 2079
rect 1484 2064 1536 2070
rect 1633 2069 1667 2073
rect 1480 2021 1484 2055
rect 1536 2021 1540 2055
rect 1618 2017 1624 2069
rect 1676 2017 1682 2069
rect 1633 2013 1667 2017
rect 1484 2006 1536 2012
rect 1448 1745 1500 1751
rect 1444 1702 1448 1736
rect 1500 1702 1504 1736
rect 1635 1702 1687 1708
rect 1448 1687 1500 1693
rect 1194 1650 1420 1678
rect 1631 1663 1635 1697
rect 1687 1663 1691 1697
rect 1194 1616 1228 1650
rect 1386 1616 1420 1650
rect 1635 1644 1687 1650
rect 1751 1616 1785 2141
rect 1092 1604 1138 1616
rect 1092 528 1098 1604
rect 1132 528 1138 1604
rect 1092 516 1138 528
rect 1188 1604 1234 1616
rect 1188 528 1194 1604
rect 1228 528 1234 1604
rect 1188 516 1234 528
rect 1284 1604 1330 1616
rect 1284 528 1290 1604
rect 1324 528 1330 1604
rect 1284 516 1330 528
rect 1380 1604 1426 1616
rect 1380 528 1386 1604
rect 1420 528 1426 1604
rect 1380 516 1426 528
rect 1476 1604 1522 1616
rect 1476 528 1482 1604
rect 1516 528 1522 1604
rect 1476 516 1522 528
rect 1572 1604 1618 1616
rect 1572 528 1578 1604
rect 1612 528 1618 1604
rect 1572 516 1618 528
rect 1668 1604 1785 1616
rect 1668 528 1674 1604
rect 1708 1582 1785 1604
rect 1708 528 1714 1582
rect 1668 516 1714 528
rect 1098 477 1132 516
rect 1674 477 1708 516
rect 1098 443 1708 477
<< via1 >>
rect 1635 3989 1687 4002
rect 761 3797 867 3903
rect 1448 3950 1500 3959
rect 1635 3955 1644 3989
rect 1644 3955 1678 3989
rect 1678 3955 1687 3989
rect 1635 3950 1687 3955
rect 1448 3916 1457 3950
rect 1457 3916 1491 3950
rect 1491 3916 1500 3950
rect 1448 3907 1500 3916
rect 1484 3631 1536 3640
rect 1484 3597 1493 3631
rect 1493 3597 1527 3631
rect 1527 3597 1536 3631
rect 1484 3588 1536 3597
rect 1624 3626 1676 3635
rect 1624 3592 1633 3626
rect 1633 3592 1667 3626
rect 1667 3592 1676 3626
rect 1624 3583 1676 3592
rect 758 1741 864 1847
rect 1484 2055 1536 2064
rect 1484 2021 1493 2055
rect 1493 2021 1527 2055
rect 1527 2021 1536 2055
rect 1484 2012 1536 2021
rect 1624 2060 1676 2069
rect 1624 2026 1633 2060
rect 1633 2026 1667 2060
rect 1667 2026 1676 2060
rect 1624 2017 1676 2026
rect 1448 1736 1500 1745
rect 1448 1702 1457 1736
rect 1457 1702 1491 1736
rect 1491 1702 1500 1736
rect 1448 1693 1500 1702
rect 1635 1697 1687 1702
rect 1635 1663 1644 1697
rect 1644 1663 1678 1697
rect 1678 1663 1687 1697
rect 1635 1650 1687 1663
<< metal2 >>
rect 1629 4002 1694 4009
rect 1442 3959 1506 3965
rect 741 3787 751 3913
rect 877 3787 887 3913
rect 1442 3907 1448 3959
rect 1500 3907 1506 3959
rect 1629 3950 1635 4002
rect 1687 3972 1694 4002
rect 1687 3950 1701 3972
rect 1629 3944 1701 3950
rect 1442 3901 1506 3907
rect 1442 3738 1476 3901
rect 1667 3873 1701 3944
rect 1508 3864 1564 3873
rect 1508 3799 1564 3808
rect 1673 3864 1729 3873
rect 1673 3799 1729 3808
rect 1406 3682 1415 3738
rect 1471 3682 1480 3738
rect 1508 3646 1542 3799
rect 1570 3682 1580 3738
rect 1636 3721 1645 3738
rect 1636 3682 1660 3721
rect 1478 3640 1542 3646
rect 1626 3641 1660 3682
rect 1478 3588 1484 3640
rect 1536 3588 1542 3640
rect 1478 3582 1542 3588
rect 1618 3635 1682 3641
rect 1618 3583 1624 3635
rect 1676 3583 1682 3635
rect 1618 3577 1682 3583
rect 1478 2064 1542 2070
rect 1478 2012 1484 2064
rect 1536 2012 1542 2064
rect 1478 2006 1542 2012
rect 1618 2069 1682 2075
rect 1618 2017 1624 2069
rect 1676 2017 1682 2069
rect 1618 2011 1682 2017
rect 1406 1915 1415 1971
rect 1471 1915 1480 1971
rect 738 1731 748 1857
rect 874 1731 884 1857
rect 1442 1751 1476 1915
rect 1508 1853 1542 2006
rect 1626 1971 1660 2011
rect 1570 1915 1580 1971
rect 1636 1934 1660 1971
rect 1636 1915 1645 1934
rect 1508 1844 1564 1853
rect 1508 1779 1564 1788
rect 1673 1844 1729 1853
rect 1673 1779 1729 1788
rect 1442 1745 1506 1751
rect 1442 1693 1448 1745
rect 1500 1693 1506 1745
rect 1667 1708 1701 1779
rect 1442 1687 1506 1693
rect 1629 1702 1701 1708
rect 1629 1650 1635 1702
rect 1687 1680 1701 1702
rect 1687 1650 1694 1680
rect 1629 1643 1694 1650
<< via2 >>
rect 751 3903 877 3913
rect 751 3797 761 3903
rect 761 3797 867 3903
rect 867 3797 877 3903
rect 751 3787 877 3797
rect 1508 3808 1564 3864
rect 1673 3808 1729 3864
rect 1415 3682 1471 3738
rect 1580 3682 1636 3738
rect 1415 1915 1471 1971
rect 748 1847 874 1857
rect 748 1741 758 1847
rect 758 1741 864 1847
rect 864 1741 874 1847
rect 748 1731 874 1741
rect 1580 1915 1636 1971
rect 1508 1788 1564 1844
rect 1673 1788 1729 1844
<< metal3 >>
rect 735 3780 741 3920
rect 887 3780 893 3920
rect 1503 3864 1734 3869
rect 1503 3808 1508 3864
rect 1564 3808 1673 3864
rect 1729 3808 1734 3864
rect 1503 3803 1734 3808
rect 1406 3738 1641 3743
rect 1406 3682 1415 3738
rect 1471 3682 1580 3738
rect 1636 3682 1641 3738
rect 1406 3677 1641 3682
rect 1410 1971 1641 1977
rect 1410 1915 1415 1971
rect 1471 1915 1580 1971
rect 1636 1915 1641 1971
rect 1410 1909 1641 1915
rect 732 1724 738 1864
rect 884 1724 890 1864
rect 1503 1844 1734 1849
rect 1503 1788 1508 1844
rect 1564 1788 1673 1844
rect 1729 1788 1734 1844
rect 1503 1783 1734 1788
<< via3 >>
rect 741 3913 887 3920
rect 741 3787 751 3913
rect 751 3787 877 3913
rect 877 3787 887 3913
rect 741 3780 887 3787
rect 738 1857 884 1864
rect 738 1731 748 1857
rect 748 1731 874 1857
rect 874 1731 884 1857
rect 738 1724 884 1731
<< metal4 >>
rect 711 3920 917 3935
rect 711 3780 741 3920
rect 887 3780 917 3920
rect 711 1864 917 3780
rect 711 1724 738 1864
rect 884 1724 917 1864
rect 711 1688 917 1724
<< labels >>
flabel metal1 1293 3796 1316 3825 0 FreeSans 320 0 0 0 vip
port 3 nsew
flabel metal2 1632 3650 1656 3672 0 FreeSans 320 0 0 0 sw_n
port 8 nsew
flabel metal2 1674 3886 1698 3916 0 FreeSans 320 0 0 0 sw
port 10 nsew
flabel metal1 1770 3739 1795 3781 0 FreeSans 320 0 0 0 tah_vp
port 12 nsew
flabel metal1 1756 1869 1780 1907 0 FreeSans 320 0 0 0 tah_vn
port 14 nsew
flabel metal1 1292 1862 1320 1901 0 FreeSans 320 0 0 0 vin
port 16 nsew
flabel space 1008 2817 1042 2835 0 FreeSans 320 0 0 0 VSS
port 20 nsew
flabel metal4 744 2724 881 2933 0 FreeSans 640 0 0 0 VDD
port 24 nsew
flabel metal2 1674 1728 1695 1760 0 FreeSans 320 0 0 0 sw
port 27 nsew
flabel metal2 1631 1982 1656 2002 0 FreeSans 320 0 0 0 sw_n
port 29 nsew
<< end >>
