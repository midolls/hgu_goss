magic
tech sky130A
magscale 1 2
timestamp 1697716041
<< nwell >>
rect -162 -118 162 118
<< pmos >>
rect -63 -80 -33 80
rect 33 -80 63 80
<< pdiff >>
rect -125 32 -63 80
rect -125 -68 -113 32
rect -79 -68 -63 32
rect -125 -80 -63 -68
rect -33 -19 33 80
rect -33 -68 -17 -19
rect 17 -68 33 -19
rect -33 -80 33 -68
rect 63 32 125 80
rect 63 -68 79 32
rect 113 -68 125 32
rect 63 -80 125 -68
<< pdiffc >>
rect -113 -68 -79 32
rect -17 -68 17 -19
rect 79 -68 113 32
<< poly >>
rect -63 80 -33 106
rect 33 80 63 110
rect -63 -111 -33 -80
rect 33 -106 63 -80
rect -81 -127 -15 -111
rect -81 -161 -65 -127
rect -31 -161 -15 -127
rect -81 -177 -15 -161
<< polycont >>
rect -65 -161 -31 -127
<< locali >>
rect -113 32 -79 48
rect 79 32 113 48
rect -113 -84 -79 -68
rect -17 -19 17 -3
rect -17 -84 17 -68
rect 79 -84 113 -68
rect -81 -161 -65 -127
rect -31 -161 -15 -127
<< viali >>
rect -113 -68 -79 32
rect -17 -68 17 -19
rect 79 -68 113 32
<< metal1 >>
rect -113 38 -79 48
rect 79 38 113 48
rect -119 32 -73 38
rect -119 -68 -113 32
rect -79 -68 -73 32
rect 73 32 119 38
rect -17 -7 17 -3
rect -119 -80 -73 -68
rect -23 -19 23 -7
rect -23 -68 -17 -19
rect 17 -68 23 -19
rect -23 -80 23 -68
rect 73 -68 79 32
rect 113 -68 119 32
rect 73 -80 119 -68
<< properties >>
string FIXED_BBOX -210 -246 210 246
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.8 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
